VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sky130_osu_ring_oscillator_mpr2aa_8_b0r1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2aa_8_b0r1 ;
  SIZE 96.725 BY 12.465 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 33.02 0 33.37 2.96 ;
      LAYER li1 ;
        RECT 33.05 1.87 33.225 2.38 ;
        RECT 33.05 3.9 33.225 5.16 ;
        RECT 33.05 3.69 33.22 5.16 ;
      LAYER met2 ;
        RECT 33.02 2.595 33.37 2.945 ;
        RECT 33.05 2.58 33.345 2.96 ;
      LAYER met1 ;
        RECT 33.05 2.625 33.37 2.915 ;
        RECT 32.99 2.18 33.285 2.41 ;
        RECT 32.99 3.66 33.28 3.89 ;
        RECT 33.05 2.18 33.22 3.89 ;
      LAYER via1 ;
        RECT 33.12 2.695 33.27 2.845 ;
      LAYER via2 ;
        RECT 33.095 2.67 33.295 2.87 ;
      LAYER mcon ;
        RECT 33.05 3.69 33.22 3.86 ;
        RECT 33.05 2.21 33.225 2.38 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 48.8 0 49.15 2.96 ;
      LAYER li1 ;
        RECT 48.83 1.87 49.005 2.38 ;
        RECT 48.83 3.9 49.005 5.16 ;
        RECT 48.83 3.69 49 5.16 ;
      LAYER met2 ;
        RECT 48.8 2.595 49.15 2.945 ;
        RECT 48.83 2.58 49.125 2.96 ;
      LAYER met1 ;
        RECT 48.83 2.625 49.15 2.915 ;
        RECT 48.77 2.18 49.065 2.41 ;
        RECT 48.77 3.66 49.06 3.89 ;
        RECT 48.83 2.18 49 3.89 ;
      LAYER via1 ;
        RECT 48.9 2.695 49.05 2.845 ;
      LAYER via2 ;
        RECT 48.875 2.67 49.075 2.87 ;
      LAYER mcon ;
        RECT 48.83 3.69 49 3.86 ;
        RECT 48.83 2.21 49.005 2.38 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 64.575 0 64.925 2.96 ;
      LAYER li1 ;
        RECT 64.605 1.87 64.78 2.38 ;
        RECT 64.605 3.9 64.78 5.16 ;
        RECT 64.605 3.69 64.775 5.16 ;
      LAYER met2 ;
        RECT 64.575 2.595 64.925 2.945 ;
        RECT 64.605 2.58 64.9 2.96 ;
      LAYER met1 ;
        RECT 64.605 2.625 64.925 2.915 ;
        RECT 64.545 2.18 64.84 2.41 ;
        RECT 64.545 3.66 64.835 3.89 ;
        RECT 64.605 2.18 64.775 3.89 ;
      LAYER via1 ;
        RECT 64.675 2.695 64.825 2.845 ;
      LAYER via2 ;
        RECT 64.65 2.67 64.85 2.87 ;
      LAYER mcon ;
        RECT 64.605 3.69 64.775 3.86 ;
        RECT 64.605 2.21 64.78 2.38 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 80.36 0 80.71 2.96 ;
      LAYER li1 ;
        RECT 80.39 1.87 80.565 2.38 ;
        RECT 80.39 3.9 80.565 5.16 ;
        RECT 80.39 3.69 80.56 5.16 ;
      LAYER met2 ;
        RECT 80.36 2.595 80.71 2.945 ;
        RECT 80.39 2.58 80.685 2.96 ;
      LAYER met1 ;
        RECT 80.39 2.625 80.71 2.915 ;
        RECT 80.33 2.18 80.625 2.41 ;
        RECT 80.33 3.66 80.62 3.89 ;
        RECT 80.39 2.18 80.56 3.89 ;
      LAYER via1 ;
        RECT 80.46 2.695 80.61 2.845 ;
      LAYER via2 ;
        RECT 80.435 2.67 80.635 2.87 ;
      LAYER mcon ;
        RECT 80.39 3.69 80.56 3.86 ;
        RECT 80.39 2.21 80.565 2.38 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 96.145 0 96.495 2.96 ;
      LAYER li1 ;
        RECT 96.175 1.87 96.35 2.38 ;
        RECT 96.175 3.9 96.35 5.16 ;
        RECT 96.175 3.69 96.345 5.16 ;
      LAYER met2 ;
        RECT 96.145 2.595 96.495 2.945 ;
        RECT 96.175 2.58 96.47 2.96 ;
      LAYER met1 ;
        RECT 96.175 2.625 96.495 2.915 ;
        RECT 96.115 2.18 96.41 2.41 ;
        RECT 96.115 3.66 96.405 3.89 ;
        RECT 96.175 2.18 96.345 3.89 ;
      LAYER via1 ;
        RECT 96.245 2.695 96.395 2.845 ;
      LAYER via2 ;
        RECT 96.22 2.67 96.42 2.87 ;
      LAYER mcon ;
        RECT 96.175 3.69 96.345 3.86 ;
        RECT 96.175 2.21 96.35 2.38 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 28.895 2.955 29.065 4.225 ;
        RECT 28.895 8.235 29.065 9.505 ;
        RECT 24.115 8.235 24.285 9.505 ;
      LAYER met2 ;
        RECT 28.815 8.14 29.165 8.49 ;
        RECT 28.81 4 29.16 4.35 ;
        RECT 28.885 4 29.06 8.49 ;
      LAYER met1 ;
        RECT 28.81 4.055 29.295 4.225 ;
        RECT 28.81 4 29.16 4.35 ;
        RECT 28.815 8.235 29.295 8.405 ;
        RECT 28.815 8.14 29.165 8.49 ;
        RECT 24.35 8.23 29.165 8.4 ;
        RECT 24.055 8.235 24.515 8.405 ;
        RECT 24.055 8.205 24.345 8.435 ;
      LAYER via1 ;
        RECT 28.91 4.1 29.06 4.25 ;
        RECT 28.915 8.24 29.065 8.39 ;
      LAYER mcon ;
        RECT 24.115 8.235 24.285 8.405 ;
        RECT 28.895 8.235 29.065 8.405 ;
        RECT 28.895 4.055 29.065 4.225 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 44.675 2.955 44.845 4.225 ;
        RECT 44.675 8.235 44.845 9.505 ;
        RECT 39.895 8.235 40.065 9.505 ;
      LAYER met2 ;
        RECT 44.595 8.14 44.945 8.49 ;
        RECT 44.59 4 44.94 4.35 ;
        RECT 44.665 4 44.84 8.49 ;
      LAYER met1 ;
        RECT 44.59 4.055 45.075 4.225 ;
        RECT 44.59 4 44.94 4.35 ;
        RECT 44.595 8.235 45.075 8.405 ;
        RECT 44.595 8.14 44.945 8.49 ;
        RECT 40.13 8.23 44.945 8.4 ;
        RECT 39.835 8.235 40.295 8.405 ;
        RECT 39.835 8.205 40.125 8.435 ;
      LAYER via1 ;
        RECT 44.69 4.1 44.84 4.25 ;
        RECT 44.695 8.24 44.845 8.39 ;
      LAYER mcon ;
        RECT 39.895 8.235 40.065 8.405 ;
        RECT 44.675 8.235 44.845 8.405 ;
        RECT 44.675 4.055 44.845 4.225 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 60.45 2.955 60.62 4.225 ;
        RECT 60.45 8.235 60.62 9.505 ;
        RECT 55.67 8.235 55.84 9.505 ;
      LAYER met2 ;
        RECT 60.37 8.14 60.72 8.49 ;
        RECT 60.365 4 60.715 4.35 ;
        RECT 60.44 4 60.615 8.49 ;
      LAYER met1 ;
        RECT 60.365 4.055 60.85 4.225 ;
        RECT 60.365 4 60.715 4.35 ;
        RECT 60.37 8.235 60.85 8.405 ;
        RECT 60.37 8.14 60.72 8.49 ;
        RECT 55.905 8.23 60.72 8.4 ;
        RECT 55.61 8.235 56.07 8.405 ;
        RECT 55.61 8.205 55.9 8.435 ;
      LAYER via1 ;
        RECT 60.465 4.1 60.615 4.25 ;
        RECT 60.47 8.24 60.62 8.39 ;
      LAYER mcon ;
        RECT 55.67 8.235 55.84 8.405 ;
        RECT 60.45 8.235 60.62 8.405 ;
        RECT 60.45 4.055 60.62 4.225 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 76.235 2.955 76.405 4.225 ;
        RECT 76.235 8.235 76.405 9.505 ;
        RECT 71.455 8.235 71.625 9.505 ;
      LAYER met2 ;
        RECT 76.155 8.14 76.505 8.49 ;
        RECT 76.15 4 76.5 4.35 ;
        RECT 76.225 4 76.4 8.49 ;
      LAYER met1 ;
        RECT 76.15 4.055 76.635 4.225 ;
        RECT 76.15 4 76.5 4.35 ;
        RECT 76.155 8.235 76.635 8.405 ;
        RECT 76.155 8.14 76.505 8.49 ;
        RECT 71.69 8.23 76.505 8.4 ;
        RECT 71.395 8.235 71.855 8.405 ;
        RECT 71.395 8.205 71.685 8.435 ;
      LAYER via1 ;
        RECT 76.25 4.1 76.4 4.25 ;
        RECT 76.255 8.24 76.405 8.39 ;
      LAYER mcon ;
        RECT 71.455 8.235 71.625 8.405 ;
        RECT 76.235 8.235 76.405 8.405 ;
        RECT 76.235 4.055 76.405 4.225 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 92.02 2.955 92.19 4.225 ;
        RECT 92.02 8.235 92.19 9.505 ;
        RECT 87.24 8.235 87.41 9.505 ;
      LAYER met2 ;
        RECT 91.94 8.14 92.29 8.49 ;
        RECT 91.935 4 92.285 4.35 ;
        RECT 92.01 4 92.185 8.49 ;
      LAYER met1 ;
        RECT 91.935 4.055 92.42 4.225 ;
        RECT 91.935 4 92.285 4.35 ;
        RECT 91.94 8.235 92.42 8.405 ;
        RECT 91.94 8.14 92.29 8.49 ;
        RECT 87.475 8.23 92.29 8.4 ;
        RECT 87.18 8.235 87.64 8.405 ;
        RECT 87.18 8.205 87.47 8.435 ;
      LAYER via1 ;
        RECT 92.035 4.1 92.185 4.25 ;
        RECT 92.04 8.24 92.19 8.39 ;
      LAYER mcon ;
        RECT 87.24 8.235 87.41 8.405 ;
        RECT 92.02 8.235 92.19 8.405 ;
        RECT 92.02 4.055 92.19 4.225 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 15.225 8.235 15.395 9.505 ;
      LAYER met1 ;
        RECT 15.165 8.235 15.625 8.405 ;
        RECT 15.17 8.2 15.46 8.43 ;
        RECT 15.165 8.205 15.455 8.435 ;
      LAYER mcon ;
        RECT 15.225 8.235 15.395 8.405 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 5.53 96.72 7.03 ;
        RECT 17.75 5.43 96.72 7.03 ;
        RECT 80.875 5.425 96.64 7.03 ;
        RECT 95.75 5.425 95.92 7.76 ;
        RECT 95.745 4.7 95.915 7.03 ;
        RECT 91.84 5.425 95.575 7.035 ;
        RECT 94.755 4.695 94.925 7.765 ;
        RECT 92.01 4.695 92.18 7.765 ;
        RECT 90.215 4.93 90.385 7.03 ;
        RECT 87.06 5.425 89.81 7.035 ;
        RECT 89.255 4.93 89.425 7.035 ;
        RECT 87.23 5.425 87.4 7.765 ;
        RECT 86.815 4.93 86.985 7.03 ;
        RECT 85.815 4.93 85.985 7.03 ;
        RECT 84.855 4.93 85.025 7.03 ;
        RECT 82.415 4.93 82.585 7.03 ;
        RECT 65.09 5.425 80.855 7.03 ;
        RECT 79.965 5.425 80.135 7.76 ;
        RECT 79.96 4.7 80.13 7.03 ;
        RECT 76.055 5.425 79.79 7.035 ;
        RECT 78.97 4.695 79.14 7.765 ;
        RECT 76.225 4.695 76.395 7.765 ;
        RECT 74.43 4.93 74.6 7.03 ;
        RECT 71.275 5.425 74.025 7.035 ;
        RECT 73.47 4.93 73.64 7.035 ;
        RECT 71.445 5.425 71.615 7.765 ;
        RECT 71.03 4.93 71.2 7.03 ;
        RECT 70.03 4.93 70.2 7.03 ;
        RECT 69.07 4.93 69.24 7.03 ;
        RECT 66.63 4.93 66.8 7.03 ;
        RECT 49.305 5.425 65.07 7.03 ;
        RECT 64.18 5.425 64.35 7.76 ;
        RECT 64.175 4.7 64.345 7.03 ;
        RECT 60.27 5.425 64.005 7.035 ;
        RECT 63.185 4.695 63.355 7.765 ;
        RECT 60.44 4.695 60.61 7.765 ;
        RECT 58.645 4.93 58.815 7.03 ;
        RECT 55.49 5.425 58.24 7.035 ;
        RECT 57.685 4.93 57.855 7.035 ;
        RECT 55.66 5.425 55.83 7.765 ;
        RECT 55.245 4.93 55.415 7.03 ;
        RECT 54.245 4.93 54.415 7.03 ;
        RECT 53.285 4.93 53.455 7.03 ;
        RECT 50.845 4.93 51.015 7.03 ;
        RECT 33.53 5.425 49.295 7.03 ;
        RECT 48.405 5.425 48.575 7.76 ;
        RECT 48.4 4.7 48.57 7.03 ;
        RECT 44.495 5.425 48.23 7.035 ;
        RECT 47.41 4.695 47.58 7.765 ;
        RECT 44.665 4.695 44.835 7.765 ;
        RECT 42.87 4.93 43.04 7.03 ;
        RECT 39.715 5.425 42.465 7.035 ;
        RECT 41.91 4.93 42.08 7.035 ;
        RECT 39.885 5.425 40.055 7.765 ;
        RECT 39.47 4.93 39.64 7.03 ;
        RECT 38.47 4.93 38.64 7.03 ;
        RECT 37.51 4.93 37.68 7.03 ;
        RECT 35.07 4.93 35.24 7.03 ;
        RECT 17.75 5.425 33.515 7.03 ;
        RECT 32.625 5.425 32.795 7.76 ;
        RECT 32.62 4.7 32.79 7.03 ;
        RECT 28.715 5.425 32.45 7.035 ;
        RECT 31.63 4.695 31.8 7.765 ;
        RECT 28.885 4.695 29.055 7.765 ;
        RECT 27.09 4.93 27.26 7.03 ;
        RECT 23.935 5.425 26.685 7.035 ;
        RECT 26.13 4.93 26.3 7.035 ;
        RECT 24.105 5.425 24.275 7.765 ;
        RECT 23.69 4.93 23.86 7.03 ;
        RECT 22.69 4.93 22.86 7.03 ;
        RECT 21.73 4.93 21.9 7.03 ;
        RECT 19.29 4.93 19.46 7.03 ;
        RECT 15.045 5.53 17.795 7.035 ;
        RECT 17.03 10.045 17.205 10.595 ;
        RECT 17.03 7.305 17.205 8.445 ;
        RECT 17.03 5.53 17.2 10.595 ;
        RECT 15.215 5.53 15.385 7.765 ;
      LAYER met1 ;
        RECT 0 5.53 96.72 7.03 ;
        RECT 17.75 5.43 96.72 7.03 ;
        RECT 80.875 5.425 96.655 7.03 ;
        RECT 91.84 5.425 95.575 7.035 ;
        RECT 81.125 5.275 90.785 7.03 ;
        RECT 87.06 5.275 89.81 7.035 ;
        RECT 65.09 5.425 80.87 7.03 ;
        RECT 76.055 5.425 79.79 7.035 ;
        RECT 65.34 5.275 75 7.03 ;
        RECT 71.275 5.275 74.025 7.035 ;
        RECT 17.75 5.425 65.085 7.03 ;
        RECT 60.27 5.425 64.005 7.035 ;
        RECT 49.555 5.275 59.215 7.03 ;
        RECT 55.49 5.275 58.24 7.035 ;
        RECT 44.495 5.425 48.23 7.035 ;
        RECT 33.78 5.275 43.44 7.03 ;
        RECT 39.715 5.275 42.465 7.035 ;
        RECT 28.715 5.425 32.45 7.035 ;
        RECT 18 5.275 27.66 7.03 ;
        RECT 23.935 5.275 26.685 7.035 ;
        RECT 15.045 5.53 17.795 7.035 ;
        RECT 16.97 8.945 17.26 9.175 ;
        RECT 16.8 8.975 17.26 9.145 ;
      LAYER mcon ;
        RECT 17.03 8.975 17.2 9.145 ;
        RECT 17.335 6.835 17.505 7.005 ;
        RECT 18.145 5.43 18.315 5.6 ;
        RECT 18.605 5.43 18.775 5.6 ;
        RECT 19.065 5.43 19.235 5.6 ;
        RECT 19.525 5.43 19.695 5.6 ;
        RECT 19.985 5.43 20.155 5.6 ;
        RECT 20.445 5.43 20.615 5.6 ;
        RECT 20.905 5.43 21.075 5.6 ;
        RECT 21.365 5.43 21.535 5.6 ;
        RECT 21.825 5.43 21.995 5.6 ;
        RECT 22.285 5.43 22.455 5.6 ;
        RECT 22.745 5.43 22.915 5.6 ;
        RECT 23.205 5.43 23.375 5.6 ;
        RECT 23.665 5.43 23.835 5.6 ;
        RECT 24.125 5.43 24.295 5.6 ;
        RECT 24.585 5.43 24.755 5.6 ;
        RECT 25.045 5.43 25.215 5.6 ;
        RECT 25.505 5.43 25.675 5.6 ;
        RECT 25.965 5.43 26.135 5.6 ;
        RECT 26.225 6.835 26.395 7.005 ;
        RECT 26.425 5.43 26.595 5.6 ;
        RECT 26.885 5.43 27.055 5.6 ;
        RECT 27.345 5.43 27.515 5.6 ;
        RECT 31.005 6.835 31.175 7.005 ;
        RECT 31.005 5.455 31.175 5.625 ;
        RECT 31.71 6.835 31.88 7.005 ;
        RECT 31.71 5.455 31.88 5.625 ;
        RECT 32.7 5.46 32.87 5.63 ;
        RECT 32.705 6.83 32.875 7 ;
        RECT 33.925 5.43 34.095 5.6 ;
        RECT 34.385 5.43 34.555 5.6 ;
        RECT 34.845 5.43 35.015 5.6 ;
        RECT 35.305 5.43 35.475 5.6 ;
        RECT 35.765 5.43 35.935 5.6 ;
        RECT 36.225 5.43 36.395 5.6 ;
        RECT 36.685 5.43 36.855 5.6 ;
        RECT 37.145 5.43 37.315 5.6 ;
        RECT 37.605 5.43 37.775 5.6 ;
        RECT 38.065 5.43 38.235 5.6 ;
        RECT 38.525 5.43 38.695 5.6 ;
        RECT 38.985 5.43 39.155 5.6 ;
        RECT 39.445 5.43 39.615 5.6 ;
        RECT 39.905 5.43 40.075 5.6 ;
        RECT 40.365 5.43 40.535 5.6 ;
        RECT 40.825 5.43 40.995 5.6 ;
        RECT 41.285 5.43 41.455 5.6 ;
        RECT 41.745 5.43 41.915 5.6 ;
        RECT 42.005 6.835 42.175 7.005 ;
        RECT 42.205 5.43 42.375 5.6 ;
        RECT 42.665 5.43 42.835 5.6 ;
        RECT 43.125 5.43 43.295 5.6 ;
        RECT 46.785 6.835 46.955 7.005 ;
        RECT 46.785 5.455 46.955 5.625 ;
        RECT 47.49 6.835 47.66 7.005 ;
        RECT 47.49 5.455 47.66 5.625 ;
        RECT 48.48 5.46 48.65 5.63 ;
        RECT 48.485 6.83 48.655 7 ;
        RECT 49.7 5.43 49.87 5.6 ;
        RECT 50.16 5.43 50.33 5.6 ;
        RECT 50.62 5.43 50.79 5.6 ;
        RECT 51.08 5.43 51.25 5.6 ;
        RECT 51.54 5.43 51.71 5.6 ;
        RECT 52 5.43 52.17 5.6 ;
        RECT 52.46 5.43 52.63 5.6 ;
        RECT 52.92 5.43 53.09 5.6 ;
        RECT 53.38 5.43 53.55 5.6 ;
        RECT 53.84 5.43 54.01 5.6 ;
        RECT 54.3 5.43 54.47 5.6 ;
        RECT 54.76 5.43 54.93 5.6 ;
        RECT 55.22 5.43 55.39 5.6 ;
        RECT 55.68 5.43 55.85 5.6 ;
        RECT 56.14 5.43 56.31 5.6 ;
        RECT 56.6 5.43 56.77 5.6 ;
        RECT 57.06 5.43 57.23 5.6 ;
        RECT 57.52 5.43 57.69 5.6 ;
        RECT 57.78 6.835 57.95 7.005 ;
        RECT 57.98 5.43 58.15 5.6 ;
        RECT 58.44 5.43 58.61 5.6 ;
        RECT 58.9 5.43 59.07 5.6 ;
        RECT 62.56 6.835 62.73 7.005 ;
        RECT 62.56 5.455 62.73 5.625 ;
        RECT 63.265 6.835 63.435 7.005 ;
        RECT 63.265 5.455 63.435 5.625 ;
        RECT 64.255 5.46 64.425 5.63 ;
        RECT 64.26 6.83 64.43 7 ;
        RECT 65.485 5.43 65.655 5.6 ;
        RECT 65.945 5.43 66.115 5.6 ;
        RECT 66.405 5.43 66.575 5.6 ;
        RECT 66.865 5.43 67.035 5.6 ;
        RECT 67.325 5.43 67.495 5.6 ;
        RECT 67.785 5.43 67.955 5.6 ;
        RECT 68.245 5.43 68.415 5.6 ;
        RECT 68.705 5.43 68.875 5.6 ;
        RECT 69.165 5.43 69.335 5.6 ;
        RECT 69.625 5.43 69.795 5.6 ;
        RECT 70.085 5.43 70.255 5.6 ;
        RECT 70.545 5.43 70.715 5.6 ;
        RECT 71.005 5.43 71.175 5.6 ;
        RECT 71.465 5.43 71.635 5.6 ;
        RECT 71.925 5.43 72.095 5.6 ;
        RECT 72.385 5.43 72.555 5.6 ;
        RECT 72.845 5.43 73.015 5.6 ;
        RECT 73.305 5.43 73.475 5.6 ;
        RECT 73.565 6.835 73.735 7.005 ;
        RECT 73.765 5.43 73.935 5.6 ;
        RECT 74.225 5.43 74.395 5.6 ;
        RECT 74.685 5.43 74.855 5.6 ;
        RECT 78.345 6.835 78.515 7.005 ;
        RECT 78.345 5.455 78.515 5.625 ;
        RECT 79.05 6.835 79.22 7.005 ;
        RECT 79.05 5.455 79.22 5.625 ;
        RECT 80.04 5.46 80.21 5.63 ;
        RECT 80.045 6.83 80.215 7 ;
        RECT 81.27 5.43 81.44 5.6 ;
        RECT 81.73 5.43 81.9 5.6 ;
        RECT 82.19 5.43 82.36 5.6 ;
        RECT 82.65 5.43 82.82 5.6 ;
        RECT 83.11 5.43 83.28 5.6 ;
        RECT 83.57 5.43 83.74 5.6 ;
        RECT 84.03 5.43 84.2 5.6 ;
        RECT 84.49 5.43 84.66 5.6 ;
        RECT 84.95 5.43 85.12 5.6 ;
        RECT 85.41 5.43 85.58 5.6 ;
        RECT 85.87 5.43 86.04 5.6 ;
        RECT 86.33 5.43 86.5 5.6 ;
        RECT 86.79 5.43 86.96 5.6 ;
        RECT 87.25 5.43 87.42 5.6 ;
        RECT 87.71 5.43 87.88 5.6 ;
        RECT 88.17 5.43 88.34 5.6 ;
        RECT 88.63 5.43 88.8 5.6 ;
        RECT 89.09 5.43 89.26 5.6 ;
        RECT 89.35 6.835 89.52 7.005 ;
        RECT 89.55 5.43 89.72 5.6 ;
        RECT 90.01 5.43 90.18 5.6 ;
        RECT 90.47 5.43 90.64 5.6 ;
        RECT 94.13 6.835 94.3 7.005 ;
        RECT 94.13 5.455 94.3 5.625 ;
        RECT 94.835 6.835 95.005 7.005 ;
        RECT 94.835 5.455 95.005 5.625 ;
        RECT 95.825 5.46 95.995 5.63 ;
        RECT 95.83 6.83 96 7 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 90.015 4.27 90.345 5 ;
        RECT 74.23 4.27 74.56 5 ;
        RECT 58.445 4.27 58.775 5 ;
        RECT 42.67 4.27 43 5 ;
        RECT 26.89 4.27 27.22 5 ;
      LAYER li1 ;
        RECT 20.02 10.86 96.725 12.465 ;
        RECT 95.75 10.23 95.92 12.465 ;
        RECT 94.755 10.235 94.925 12.465 ;
        RECT 92.01 10.235 92.18 12.465 ;
        RECT 87.23 10.235 87.4 12.465 ;
        RECT 79.965 10.23 80.135 12.465 ;
        RECT 78.97 10.235 79.14 12.465 ;
        RECT 76.225 10.235 76.395 12.465 ;
        RECT 71.445 10.235 71.615 12.465 ;
        RECT 64.18 10.23 64.35 12.465 ;
        RECT 63.185 10.235 63.355 12.465 ;
        RECT 60.44 10.235 60.61 12.465 ;
        RECT 55.66 10.235 55.83 12.465 ;
        RECT 48.405 10.23 48.575 12.465 ;
        RECT 47.41 10.235 47.58 12.465 ;
        RECT 44.665 10.235 44.835 12.465 ;
        RECT 39.885 10.235 40.055 12.465 ;
        RECT 32.625 10.23 32.795 12.465 ;
        RECT 31.63 10.235 31.8 12.465 ;
        RECT 28.885 10.235 29.055 12.465 ;
        RECT 24.105 10.235 24.275 12.465 ;
        RECT 0.03 10.86 96.725 12.46 ;
        RECT 15.215 10.235 15.385 12.46 ;
        RECT 0 0 96.72 1.6 ;
        RECT 95.745 0 95.915 2.23 ;
        RECT 94.755 0 94.925 2.225 ;
        RECT 92.01 0 92.18 2.225 ;
        RECT 81.125 2.71 90.955 2.88 ;
        RECT 81.24 0 90.955 2.88 ;
        RECT 81.24 0 90.84 2.885 ;
        RECT 89.255 0 89.425 3.38 ;
        RECT 87.295 0 87.465 3.38 ;
        RECT 84.855 0 85.025 3.38 ;
        RECT 83.895 0 84.065 3.38 ;
        RECT 83.375 0 83.545 3.38 ;
        RECT 82.415 0 82.585 3.38 ;
        RECT 81.455 0 81.625 3.38 ;
        RECT 79.96 0 80.13 2.23 ;
        RECT 78.97 0 79.14 2.225 ;
        RECT 76.225 0 76.395 2.225 ;
        RECT 65.34 2.71 75.17 2.88 ;
        RECT 65.455 0 75.17 2.88 ;
        RECT 65.455 0 75.055 2.885 ;
        RECT 73.47 0 73.64 3.38 ;
        RECT 71.51 0 71.68 3.38 ;
        RECT 69.07 0 69.24 3.38 ;
        RECT 68.11 0 68.28 3.38 ;
        RECT 67.59 0 67.76 3.38 ;
        RECT 66.63 0 66.8 3.38 ;
        RECT 65.67 0 65.84 3.38 ;
        RECT 64.175 0 64.345 2.23 ;
        RECT 63.185 0 63.355 2.225 ;
        RECT 60.44 0 60.61 2.225 ;
        RECT 49.555 2.71 59.385 2.88 ;
        RECT 49.67 0 59.385 2.88 ;
        RECT 49.67 0 59.27 2.885 ;
        RECT 57.685 0 57.855 3.38 ;
        RECT 55.725 0 55.895 3.38 ;
        RECT 53.285 0 53.455 3.38 ;
        RECT 52.325 0 52.495 3.38 ;
        RECT 51.805 0 51.975 3.38 ;
        RECT 50.845 0 51.015 3.38 ;
        RECT 49.885 0 50.055 3.38 ;
        RECT 48.4 0 48.57 2.23 ;
        RECT 47.41 0 47.58 2.225 ;
        RECT 44.665 0 44.835 2.225 ;
        RECT 33.78 2.71 43.61 2.88 ;
        RECT 33.895 0 43.61 2.88 ;
        RECT 33.895 0 43.495 2.885 ;
        RECT 41.91 0 42.08 3.38 ;
        RECT 39.95 0 40.12 3.38 ;
        RECT 37.51 0 37.68 3.38 ;
        RECT 36.55 0 36.72 3.38 ;
        RECT 36.03 0 36.2 3.38 ;
        RECT 35.07 0 35.24 3.38 ;
        RECT 34.11 0 34.28 3.38 ;
        RECT 32.62 0 32.79 2.23 ;
        RECT 31.63 0 31.8 2.225 ;
        RECT 28.885 0 29.055 2.225 ;
        RECT 18 2.71 27.83 2.88 ;
        RECT 18.115 0 27.83 2.88 ;
        RECT 18.115 0 27.715 2.885 ;
        RECT 26.13 0 26.3 3.38 ;
        RECT 24.17 0 24.34 3.38 ;
        RECT 21.73 0 21.9 3.38 ;
        RECT 20.77 0 20.94 3.38 ;
        RECT 20.25 0 20.42 3.38 ;
        RECT 19.29 0 19.46 3.38 ;
        RECT 18.33 0 18.5 3.38 ;
        RECT 90.04 3.87 90.37 4.34 ;
        RECT 90.005 3.87 90.37 4.2 ;
        RECT 90 3.87 90.37 4.125 ;
        RECT 89.975 3.87 90.37 4.12 ;
        RECT 88.195 3.87 88.425 4.225 ;
        RECT 88.14 3.87 88.425 4.2 ;
        RECT 88.125 3.87 88.425 4.16 ;
        RECT 88.08 3.87 88.425 4.15 ;
        RECT 88.015 3.87 88.425 4.12 ;
        RECT 88.245 8.365 88.415 10.315 ;
        RECT 88.185 10.145 88.355 10.595 ;
        RECT 88.185 7.305 88.355 8.535 ;
        RECT 74.255 3.87 74.585 4.34 ;
        RECT 74.22 3.87 74.585 4.2 ;
        RECT 74.215 3.87 74.585 4.125 ;
        RECT 74.19 3.87 74.585 4.12 ;
        RECT 72.41 3.87 72.64 4.225 ;
        RECT 72.355 3.87 72.64 4.2 ;
        RECT 72.34 3.87 72.64 4.16 ;
        RECT 72.295 3.87 72.64 4.15 ;
        RECT 72.23 3.87 72.64 4.12 ;
        RECT 72.46 8.365 72.63 10.315 ;
        RECT 72.4 10.145 72.57 10.595 ;
        RECT 72.4 7.305 72.57 8.535 ;
        RECT 58.47 3.87 58.8 4.34 ;
        RECT 58.435 3.87 58.8 4.2 ;
        RECT 58.43 3.87 58.8 4.125 ;
        RECT 58.405 3.87 58.8 4.12 ;
        RECT 56.625 3.87 56.855 4.225 ;
        RECT 56.57 3.87 56.855 4.2 ;
        RECT 56.555 3.87 56.855 4.16 ;
        RECT 56.51 3.87 56.855 4.15 ;
        RECT 56.445 3.87 56.855 4.12 ;
        RECT 56.675 8.365 56.845 10.315 ;
        RECT 56.615 10.145 56.785 10.595 ;
        RECT 56.615 7.305 56.785 8.535 ;
        RECT 42.695 3.87 43.025 4.34 ;
        RECT 42.66 3.87 43.025 4.2 ;
        RECT 42.655 3.87 43.025 4.125 ;
        RECT 42.63 3.87 43.025 4.12 ;
        RECT 40.85 3.87 41.08 4.225 ;
        RECT 40.795 3.87 41.08 4.2 ;
        RECT 40.78 3.87 41.08 4.16 ;
        RECT 40.735 3.87 41.08 4.15 ;
        RECT 40.67 3.87 41.08 4.12 ;
        RECT 40.9 8.365 41.07 10.315 ;
        RECT 40.84 10.145 41.01 10.595 ;
        RECT 40.84 7.305 41.01 8.535 ;
        RECT 26.915 3.87 27.245 4.34 ;
        RECT 26.88 3.87 27.245 4.2 ;
        RECT 26.875 3.87 27.245 4.125 ;
        RECT 26.85 3.87 27.245 4.12 ;
        RECT 25.07 3.87 25.3 4.225 ;
        RECT 25.015 3.87 25.3 4.2 ;
        RECT 25 3.87 25.3 4.16 ;
        RECT 24.955 3.87 25.3 4.15 ;
        RECT 24.89 3.87 25.3 4.12 ;
        RECT 25.12 8.365 25.29 10.315 ;
        RECT 25.06 10.145 25.23 10.595 ;
        RECT 25.06 7.305 25.23 8.535 ;
      LAYER met2 ;
        RECT 90.02 4.055 90.345 4.575 ;
        RECT 74.235 4.055 74.56 4.575 ;
        RECT 58.45 4.055 58.775 4.575 ;
        RECT 42.675 4.055 43 4.575 ;
        RECT 26.895 4.055 27.22 4.575 ;
      LAYER met1 ;
        RECT 20.02 10.86 96.725 12.465 ;
        RECT 88.185 8.575 88.475 8.805 ;
        RECT 88.01 8.605 88.475 8.775 ;
        RECT 87.81 8.6 88.18 8.77 ;
        RECT 87.81 8.6 87.98 12.465 ;
        RECT 72.4 8.575 72.69 8.805 ;
        RECT 72.225 8.605 72.69 8.775 ;
        RECT 72.025 8.6 72.395 8.77 ;
        RECT 72.025 8.6 72.195 12.465 ;
        RECT 56.615 8.575 56.905 8.805 ;
        RECT 56.44 8.605 56.905 8.775 ;
        RECT 56.24 8.6 56.61 8.77 ;
        RECT 56.24 8.6 56.41 12.465 ;
        RECT 40.84 8.575 41.13 8.805 ;
        RECT 40.665 8.605 41.13 8.775 ;
        RECT 40.465 8.6 40.835 8.77 ;
        RECT 40.465 8.6 40.635 12.465 ;
        RECT 25.06 8.575 25.35 8.805 ;
        RECT 24.885 8.605 25.35 8.775 ;
        RECT 24.685 8.6 25.055 8.77 ;
        RECT 24.685 8.6 24.855 12.465 ;
        RECT 0.03 10.86 96.725 12.46 ;
        RECT 0 0 96.72 1.6 ;
        RECT 81.125 2.555 90.955 3.035 ;
        RECT 81.24 0 90.955 3.035 ;
        RECT 90.63 0 90.805 4.315 ;
        RECT 89.815 4.275 90.805 4.315 ;
        RECT 89.985 4.14 90.805 4.315 ;
        RECT 89.985 4.03 90.345 4.575 ;
        RECT 89.335 4.37 90.345 4.535 ;
        RECT 89.945 4.215 90.345 4.535 ;
        RECT 89.655 4.365 90.345 4.535 ;
        RECT 89.92 4.235 90.345 4.535 ;
        RECT 89.675 4.36 90.345 4.535 ;
        RECT 89.91 4.245 90.345 4.535 ;
        RECT 89.705 4.355 90.345 4.535 ;
        RECT 89.89 4.25 90.345 4.535 ;
        RECT 89.71 4.34 90.345 4.535 ;
        RECT 89.88 4.26 90.345 4.535 ;
        RECT 89.74 4.335 90.345 4.535 ;
        RECT 89.865 4.265 90.345 4.535 ;
        RECT 89.755 4.3 90.345 4.535 ;
        RECT 89.4 4.37 89.625 4.555 ;
        RECT 88.815 4.365 89.57 4.37 ;
        RECT 88.8 4.36 89.555 4.365 ;
        RECT 88.78 4.355 89.525 4.36 ;
        RECT 88.73 4.34 89.505 4.355 ;
        RECT 88.71 4.335 89.44 4.34 ;
        RECT 88.595 4.3 89.415 4.335 ;
        RECT 89.035 4.37 90.345 4.52 ;
        RECT 88.45 4.245 89.27 4.3 ;
        RECT 88.225 4.235 89.04 4.255 ;
        RECT 88.865 4.37 90.345 4.43 ;
        RECT 88.225 4.215 88.99 4.255 ;
        RECT 88.225 4.2 88.9 4.255 ;
        RECT 88.85 4.37 90.345 4.38 ;
        RECT 88.225 4.18 88.85 4.255 ;
        RECT 88.83 4.37 90.345 4.375 ;
        RECT 88.225 4.175 88.79 4.255 ;
        RECT 88.225 4.16 88.77 4.255 ;
        RECT 88.225 4.14 88.725 4.255 ;
        RECT 88.225 4.135 88.645 4.255 ;
        RECT 88.225 4.08 88.625 4.255 ;
        RECT 88.225 4.015 88.46 4.255 ;
        RECT 65.34 2.555 75.17 3.035 ;
        RECT 65.455 0 75.17 3.035 ;
        RECT 74.845 0 75.02 4.315 ;
        RECT 74.03 4.275 75.02 4.315 ;
        RECT 74.2 4.14 75.02 4.315 ;
        RECT 74.2 4.03 74.56 4.575 ;
        RECT 73.55 4.37 74.56 4.535 ;
        RECT 74.16 4.215 74.56 4.535 ;
        RECT 73.87 4.365 74.56 4.535 ;
        RECT 74.135 4.235 74.56 4.535 ;
        RECT 73.89 4.36 74.56 4.535 ;
        RECT 74.125 4.245 74.56 4.535 ;
        RECT 73.92 4.355 74.56 4.535 ;
        RECT 74.105 4.25 74.56 4.535 ;
        RECT 73.925 4.34 74.56 4.535 ;
        RECT 74.095 4.26 74.56 4.535 ;
        RECT 73.955 4.335 74.56 4.535 ;
        RECT 74.08 4.265 74.56 4.535 ;
        RECT 73.97 4.3 74.56 4.535 ;
        RECT 73.615 4.37 73.84 4.555 ;
        RECT 73.03 4.365 73.785 4.37 ;
        RECT 73.015 4.36 73.77 4.365 ;
        RECT 72.995 4.355 73.74 4.36 ;
        RECT 72.945 4.34 73.72 4.355 ;
        RECT 72.925 4.335 73.655 4.34 ;
        RECT 72.81 4.3 73.63 4.335 ;
        RECT 73.25 4.37 74.56 4.52 ;
        RECT 72.665 4.245 73.485 4.3 ;
        RECT 72.44 4.235 73.255 4.255 ;
        RECT 73.08 4.37 74.56 4.43 ;
        RECT 72.44 4.215 73.205 4.255 ;
        RECT 72.44 4.2 73.115 4.255 ;
        RECT 73.065 4.37 74.56 4.38 ;
        RECT 72.44 4.18 73.065 4.255 ;
        RECT 73.045 4.37 74.56 4.375 ;
        RECT 72.44 4.175 73.005 4.255 ;
        RECT 72.44 4.16 72.985 4.255 ;
        RECT 72.44 4.14 72.94 4.255 ;
        RECT 72.44 4.135 72.86 4.255 ;
        RECT 72.44 4.08 72.84 4.255 ;
        RECT 72.44 4.015 72.675 4.255 ;
        RECT 49.555 2.555 59.385 3.035 ;
        RECT 49.67 0 59.385 3.035 ;
        RECT 59.06 0 59.235 4.315 ;
        RECT 58.245 4.275 59.235 4.315 ;
        RECT 58.415 4.14 59.235 4.315 ;
        RECT 58.415 4.03 58.775 4.575 ;
        RECT 57.765 4.37 58.775 4.535 ;
        RECT 58.375 4.215 58.775 4.535 ;
        RECT 58.085 4.365 58.775 4.535 ;
        RECT 58.35 4.235 58.775 4.535 ;
        RECT 58.105 4.36 58.775 4.535 ;
        RECT 58.34 4.245 58.775 4.535 ;
        RECT 58.135 4.355 58.775 4.535 ;
        RECT 58.32 4.25 58.775 4.535 ;
        RECT 58.14 4.34 58.775 4.535 ;
        RECT 58.31 4.26 58.775 4.535 ;
        RECT 58.17 4.335 58.775 4.535 ;
        RECT 58.295 4.265 58.775 4.535 ;
        RECT 58.185 4.3 58.775 4.535 ;
        RECT 57.83 4.37 58.055 4.555 ;
        RECT 57.245 4.365 58 4.37 ;
        RECT 57.23 4.36 57.985 4.365 ;
        RECT 57.21 4.355 57.955 4.36 ;
        RECT 57.16 4.34 57.935 4.355 ;
        RECT 57.14 4.335 57.87 4.34 ;
        RECT 57.025 4.3 57.845 4.335 ;
        RECT 57.465 4.37 58.775 4.52 ;
        RECT 56.88 4.245 57.7 4.3 ;
        RECT 56.655 4.235 57.47 4.255 ;
        RECT 57.295 4.37 58.775 4.43 ;
        RECT 56.655 4.215 57.42 4.255 ;
        RECT 56.655 4.2 57.33 4.255 ;
        RECT 57.28 4.37 58.775 4.38 ;
        RECT 56.655 4.18 57.28 4.255 ;
        RECT 57.26 4.37 58.775 4.375 ;
        RECT 56.655 4.175 57.22 4.255 ;
        RECT 56.655 4.16 57.2 4.255 ;
        RECT 56.655 4.14 57.155 4.255 ;
        RECT 56.655 4.135 57.075 4.255 ;
        RECT 56.655 4.08 57.055 4.255 ;
        RECT 56.655 4.015 56.89 4.255 ;
        RECT 33.78 2.555 43.61 3.035 ;
        RECT 33.895 0 43.61 3.035 ;
        RECT 43.285 0 43.46 4.315 ;
        RECT 42.47 4.275 43.46 4.315 ;
        RECT 42.64 4.14 43.46 4.315 ;
        RECT 42.64 4.03 43 4.575 ;
        RECT 41.99 4.37 43 4.535 ;
        RECT 42.6 4.215 43 4.535 ;
        RECT 42.31 4.365 43 4.535 ;
        RECT 42.575 4.235 43 4.535 ;
        RECT 42.33 4.36 43 4.535 ;
        RECT 42.565 4.245 43 4.535 ;
        RECT 42.36 4.355 43 4.535 ;
        RECT 42.545 4.25 43 4.535 ;
        RECT 42.365 4.34 43 4.535 ;
        RECT 42.535 4.26 43 4.535 ;
        RECT 42.395 4.335 43 4.535 ;
        RECT 42.52 4.265 43 4.535 ;
        RECT 42.41 4.3 43 4.535 ;
        RECT 42.055 4.37 42.28 4.555 ;
        RECT 41.47 4.365 42.225 4.37 ;
        RECT 41.455 4.36 42.21 4.365 ;
        RECT 41.435 4.355 42.18 4.36 ;
        RECT 41.385 4.34 42.16 4.355 ;
        RECT 41.365 4.335 42.095 4.34 ;
        RECT 41.25 4.3 42.07 4.335 ;
        RECT 41.69 4.37 43 4.52 ;
        RECT 41.105 4.245 41.925 4.3 ;
        RECT 40.88 4.235 41.695 4.255 ;
        RECT 41.52 4.37 43 4.43 ;
        RECT 40.88 4.215 41.645 4.255 ;
        RECT 40.88 4.2 41.555 4.255 ;
        RECT 41.505 4.37 43 4.38 ;
        RECT 40.88 4.18 41.505 4.255 ;
        RECT 41.485 4.37 43 4.375 ;
        RECT 40.88 4.175 41.445 4.255 ;
        RECT 40.88 4.16 41.425 4.255 ;
        RECT 40.88 4.14 41.38 4.255 ;
        RECT 40.88 4.135 41.3 4.255 ;
        RECT 40.88 4.08 41.28 4.255 ;
        RECT 40.88 4.015 41.115 4.255 ;
        RECT 18 2.555 27.83 3.035 ;
        RECT 18.115 0 27.83 3.035 ;
        RECT 27.505 0 27.68 4.315 ;
        RECT 26.69 4.275 27.68 4.315 ;
        RECT 26.86 4.14 27.68 4.315 ;
        RECT 26.86 4.03 27.22 4.575 ;
        RECT 26.21 4.37 27.22 4.535 ;
        RECT 26.82 4.215 27.22 4.535 ;
        RECT 26.53 4.365 27.22 4.535 ;
        RECT 26.795 4.235 27.22 4.535 ;
        RECT 26.55 4.36 27.22 4.535 ;
        RECT 26.785 4.245 27.22 4.535 ;
        RECT 26.58 4.355 27.22 4.535 ;
        RECT 26.765 4.25 27.22 4.535 ;
        RECT 26.585 4.34 27.22 4.535 ;
        RECT 26.755 4.26 27.22 4.535 ;
        RECT 26.615 4.335 27.22 4.535 ;
        RECT 26.74 4.265 27.22 4.535 ;
        RECT 26.63 4.3 27.22 4.535 ;
        RECT 26.275 4.37 26.5 4.555 ;
        RECT 25.69 4.365 26.445 4.37 ;
        RECT 25.675 4.36 26.43 4.365 ;
        RECT 25.655 4.355 26.4 4.36 ;
        RECT 25.605 4.34 26.38 4.355 ;
        RECT 25.585 4.335 26.315 4.34 ;
        RECT 25.47 4.3 26.29 4.335 ;
        RECT 25.91 4.37 27.22 4.52 ;
        RECT 25.325 4.245 26.145 4.3 ;
        RECT 25.1 4.235 25.915 4.255 ;
        RECT 25.74 4.37 27.22 4.43 ;
        RECT 25.1 4.215 25.865 4.255 ;
        RECT 25.1 4.2 25.775 4.255 ;
        RECT 25.725 4.37 27.22 4.38 ;
        RECT 25.1 4.18 25.725 4.255 ;
        RECT 25.705 4.37 27.22 4.375 ;
        RECT 25.1 4.175 25.665 4.255 ;
        RECT 25.1 4.16 25.645 4.255 ;
        RECT 25.1 4.14 25.6 4.255 ;
        RECT 25.1 4.135 25.52 4.255 ;
        RECT 25.1 4.08 25.5 4.255 ;
        RECT 25.1 4.015 25.335 4.255 ;
      LAYER via1 ;
        RECT 26.97 4.155 27.12 4.305 ;
        RECT 42.75 4.155 42.9 4.305 ;
        RECT 58.525 4.155 58.675 4.305 ;
        RECT 74.31 4.155 74.46 4.305 ;
        RECT 90.095 4.155 90.245 4.305 ;
      LAYER via2 ;
        RECT 26.955 4.335 27.155 4.535 ;
        RECT 42.735 4.335 42.935 4.535 ;
        RECT 58.51 4.335 58.71 4.535 ;
        RECT 74.295 4.335 74.495 4.535 ;
        RECT 90.08 4.335 90.28 4.535 ;
      LAYER mcon ;
        RECT 15.295 10.895 15.465 11.065 ;
        RECT 15.975 10.895 16.145 11.065 ;
        RECT 16.655 10.895 16.825 11.065 ;
        RECT 17.335 10.895 17.505 11.065 ;
        RECT 18.145 2.71 18.315 2.88 ;
        RECT 18.605 2.71 18.775 2.88 ;
        RECT 19.065 2.71 19.235 2.88 ;
        RECT 19.525 2.71 19.695 2.88 ;
        RECT 19.985 2.71 20.155 2.88 ;
        RECT 20.445 2.71 20.615 2.88 ;
        RECT 20.905 2.71 21.075 2.88 ;
        RECT 21.365 2.71 21.535 2.88 ;
        RECT 21.825 2.71 21.995 2.88 ;
        RECT 22.285 2.71 22.455 2.88 ;
        RECT 22.745 2.71 22.915 2.88 ;
        RECT 23.205 2.71 23.375 2.88 ;
        RECT 23.665 2.71 23.835 2.88 ;
        RECT 24.125 2.71 24.295 2.88 ;
        RECT 24.185 10.895 24.355 11.065 ;
        RECT 24.585 2.71 24.755 2.88 ;
        RECT 24.865 10.895 25.035 11.065 ;
        RECT 25.045 2.71 25.215 2.88 ;
        RECT 25.12 8.605 25.29 8.775 ;
        RECT 25.13 4.055 25.3 4.225 ;
        RECT 25.505 2.71 25.675 2.88 ;
        RECT 25.545 10.895 25.715 11.065 ;
        RECT 25.965 2.71 26.135 2.88 ;
        RECT 26.225 10.895 26.395 11.065 ;
        RECT 26.425 2.71 26.595 2.88 ;
        RECT 26.885 2.71 27.055 2.88 ;
        RECT 26.975 4.17 27.145 4.34 ;
        RECT 27.345 2.71 27.515 2.88 ;
        RECT 28.965 10.895 29.135 11.065 ;
        RECT 28.965 1.395 29.135 1.565 ;
        RECT 29.645 10.895 29.815 11.065 ;
        RECT 29.645 1.395 29.815 1.565 ;
        RECT 30.325 10.895 30.495 11.065 ;
        RECT 30.325 1.395 30.495 1.565 ;
        RECT 31.005 10.895 31.175 11.065 ;
        RECT 31.005 1.395 31.175 1.565 ;
        RECT 31.71 10.895 31.88 11.065 ;
        RECT 31.71 1.395 31.88 1.565 ;
        RECT 32.7 1.4 32.87 1.57 ;
        RECT 32.705 10.89 32.875 11.06 ;
        RECT 33.925 2.71 34.095 2.88 ;
        RECT 34.385 2.71 34.555 2.88 ;
        RECT 34.845 2.71 35.015 2.88 ;
        RECT 35.305 2.71 35.475 2.88 ;
        RECT 35.765 2.71 35.935 2.88 ;
        RECT 36.225 2.71 36.395 2.88 ;
        RECT 36.685 2.71 36.855 2.88 ;
        RECT 37.145 2.71 37.315 2.88 ;
        RECT 37.605 2.71 37.775 2.88 ;
        RECT 38.065 2.71 38.235 2.88 ;
        RECT 38.525 2.71 38.695 2.88 ;
        RECT 38.985 2.71 39.155 2.88 ;
        RECT 39.445 2.71 39.615 2.88 ;
        RECT 39.905 2.71 40.075 2.88 ;
        RECT 39.965 10.895 40.135 11.065 ;
        RECT 40.365 2.71 40.535 2.88 ;
        RECT 40.645 10.895 40.815 11.065 ;
        RECT 40.825 2.71 40.995 2.88 ;
        RECT 40.9 8.605 41.07 8.775 ;
        RECT 40.91 4.055 41.08 4.225 ;
        RECT 41.285 2.71 41.455 2.88 ;
        RECT 41.325 10.895 41.495 11.065 ;
        RECT 41.745 2.71 41.915 2.88 ;
        RECT 42.005 10.895 42.175 11.065 ;
        RECT 42.205 2.71 42.375 2.88 ;
        RECT 42.665 2.71 42.835 2.88 ;
        RECT 42.755 4.17 42.925 4.34 ;
        RECT 43.125 2.71 43.295 2.88 ;
        RECT 44.745 10.895 44.915 11.065 ;
        RECT 44.745 1.395 44.915 1.565 ;
        RECT 45.425 10.895 45.595 11.065 ;
        RECT 45.425 1.395 45.595 1.565 ;
        RECT 46.105 10.895 46.275 11.065 ;
        RECT 46.105 1.395 46.275 1.565 ;
        RECT 46.785 10.895 46.955 11.065 ;
        RECT 46.785 1.395 46.955 1.565 ;
        RECT 47.49 10.895 47.66 11.065 ;
        RECT 47.49 1.395 47.66 1.565 ;
        RECT 48.48 1.4 48.65 1.57 ;
        RECT 48.485 10.89 48.655 11.06 ;
        RECT 49.7 2.71 49.87 2.88 ;
        RECT 50.16 2.71 50.33 2.88 ;
        RECT 50.62 2.71 50.79 2.88 ;
        RECT 51.08 2.71 51.25 2.88 ;
        RECT 51.54 2.71 51.71 2.88 ;
        RECT 52 2.71 52.17 2.88 ;
        RECT 52.46 2.71 52.63 2.88 ;
        RECT 52.92 2.71 53.09 2.88 ;
        RECT 53.38 2.71 53.55 2.88 ;
        RECT 53.84 2.71 54.01 2.88 ;
        RECT 54.3 2.71 54.47 2.88 ;
        RECT 54.76 2.71 54.93 2.88 ;
        RECT 55.22 2.71 55.39 2.88 ;
        RECT 55.68 2.71 55.85 2.88 ;
        RECT 55.74 10.895 55.91 11.065 ;
        RECT 56.14 2.71 56.31 2.88 ;
        RECT 56.42 10.895 56.59 11.065 ;
        RECT 56.6 2.71 56.77 2.88 ;
        RECT 56.675 8.605 56.845 8.775 ;
        RECT 56.685 4.055 56.855 4.225 ;
        RECT 57.06 2.71 57.23 2.88 ;
        RECT 57.1 10.895 57.27 11.065 ;
        RECT 57.52 2.71 57.69 2.88 ;
        RECT 57.78 10.895 57.95 11.065 ;
        RECT 57.98 2.71 58.15 2.88 ;
        RECT 58.44 2.71 58.61 2.88 ;
        RECT 58.53 4.17 58.7 4.34 ;
        RECT 58.9 2.71 59.07 2.88 ;
        RECT 60.52 10.895 60.69 11.065 ;
        RECT 60.52 1.395 60.69 1.565 ;
        RECT 61.2 10.895 61.37 11.065 ;
        RECT 61.2 1.395 61.37 1.565 ;
        RECT 61.88 10.895 62.05 11.065 ;
        RECT 61.88 1.395 62.05 1.565 ;
        RECT 62.56 10.895 62.73 11.065 ;
        RECT 62.56 1.395 62.73 1.565 ;
        RECT 63.265 10.895 63.435 11.065 ;
        RECT 63.265 1.395 63.435 1.565 ;
        RECT 64.255 1.4 64.425 1.57 ;
        RECT 64.26 10.89 64.43 11.06 ;
        RECT 65.485 2.71 65.655 2.88 ;
        RECT 65.945 2.71 66.115 2.88 ;
        RECT 66.405 2.71 66.575 2.88 ;
        RECT 66.865 2.71 67.035 2.88 ;
        RECT 67.325 2.71 67.495 2.88 ;
        RECT 67.785 2.71 67.955 2.88 ;
        RECT 68.245 2.71 68.415 2.88 ;
        RECT 68.705 2.71 68.875 2.88 ;
        RECT 69.165 2.71 69.335 2.88 ;
        RECT 69.625 2.71 69.795 2.88 ;
        RECT 70.085 2.71 70.255 2.88 ;
        RECT 70.545 2.71 70.715 2.88 ;
        RECT 71.005 2.71 71.175 2.88 ;
        RECT 71.465 2.71 71.635 2.88 ;
        RECT 71.525 10.895 71.695 11.065 ;
        RECT 71.925 2.71 72.095 2.88 ;
        RECT 72.205 10.895 72.375 11.065 ;
        RECT 72.385 2.71 72.555 2.88 ;
        RECT 72.46 8.605 72.63 8.775 ;
        RECT 72.47 4.055 72.64 4.225 ;
        RECT 72.845 2.71 73.015 2.88 ;
        RECT 72.885 10.895 73.055 11.065 ;
        RECT 73.305 2.71 73.475 2.88 ;
        RECT 73.565 10.895 73.735 11.065 ;
        RECT 73.765 2.71 73.935 2.88 ;
        RECT 74.225 2.71 74.395 2.88 ;
        RECT 74.315 4.17 74.485 4.34 ;
        RECT 74.685 2.71 74.855 2.88 ;
        RECT 76.305 10.895 76.475 11.065 ;
        RECT 76.305 1.395 76.475 1.565 ;
        RECT 76.985 10.895 77.155 11.065 ;
        RECT 76.985 1.395 77.155 1.565 ;
        RECT 77.665 10.895 77.835 11.065 ;
        RECT 77.665 1.395 77.835 1.565 ;
        RECT 78.345 10.895 78.515 11.065 ;
        RECT 78.345 1.395 78.515 1.565 ;
        RECT 79.05 10.895 79.22 11.065 ;
        RECT 79.05 1.395 79.22 1.565 ;
        RECT 80.04 1.4 80.21 1.57 ;
        RECT 80.045 10.89 80.215 11.06 ;
        RECT 81.27 2.71 81.44 2.88 ;
        RECT 81.73 2.71 81.9 2.88 ;
        RECT 82.19 2.71 82.36 2.88 ;
        RECT 82.65 2.71 82.82 2.88 ;
        RECT 83.11 2.71 83.28 2.88 ;
        RECT 83.57 2.71 83.74 2.88 ;
        RECT 84.03 2.71 84.2 2.88 ;
        RECT 84.49 2.71 84.66 2.88 ;
        RECT 84.95 2.71 85.12 2.88 ;
        RECT 85.41 2.71 85.58 2.88 ;
        RECT 85.87 2.71 86.04 2.88 ;
        RECT 86.33 2.71 86.5 2.88 ;
        RECT 86.79 2.71 86.96 2.88 ;
        RECT 87.25 2.71 87.42 2.88 ;
        RECT 87.31 10.895 87.48 11.065 ;
        RECT 87.71 2.71 87.88 2.88 ;
        RECT 87.99 10.895 88.16 11.065 ;
        RECT 88.17 2.71 88.34 2.88 ;
        RECT 88.245 8.605 88.415 8.775 ;
        RECT 88.255 4.055 88.425 4.225 ;
        RECT 88.63 2.71 88.8 2.88 ;
        RECT 88.67 10.895 88.84 11.065 ;
        RECT 89.09 2.71 89.26 2.88 ;
        RECT 89.35 10.895 89.52 11.065 ;
        RECT 89.55 2.71 89.72 2.88 ;
        RECT 90.01 2.71 90.18 2.88 ;
        RECT 90.1 4.17 90.27 4.34 ;
        RECT 90.47 2.71 90.64 2.88 ;
        RECT 92.09 10.895 92.26 11.065 ;
        RECT 92.09 1.395 92.26 1.565 ;
        RECT 92.77 10.895 92.94 11.065 ;
        RECT 92.77 1.395 92.94 1.565 ;
        RECT 93.45 10.895 93.62 11.065 ;
        RECT 93.45 1.395 93.62 1.565 ;
        RECT 94.13 10.895 94.3 11.065 ;
        RECT 94.13 1.395 94.3 1.565 ;
        RECT 94.835 10.895 95.005 11.065 ;
        RECT 94.835 1.395 95.005 1.565 ;
        RECT 95.825 1.4 95.995 1.57 ;
        RECT 95.83 10.89 96 11.06 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 96.095 7.215 96.445 12.46 ;
      RECT 96.095 7.215 96.45 7.57 ;
      RECT 88.515 9.325 88.885 9.695 ;
      RECT 88.555 9.005 88.89 9.37 ;
      RECT 88.555 9.005 88.94 9.315 ;
      RECT 88.555 9.005 91.345 9.31 ;
      RECT 91.04 4.145 91.345 9.31 ;
      RECT 91.005 4.145 91.375 4.515 ;
      RECT 86.375 3.145 86.705 4.04 ;
      RECT 85.495 3.31 85.825 4.04 ;
      RECT 86.37 3.145 86.74 3.945 ;
      RECT 89.535 3.145 89.865 3.875 ;
      RECT 89.495 3.03 89.675 3.68 ;
      RECT 85.505 3.145 89.865 3.515 ;
      RECT 85.995 4.83 86.325 5.16 ;
      RECT 84.79 4.845 86.325 5.145 ;
      RECT 84.79 3.725 85.09 5.145 ;
      RECT 84.535 3.71 84.865 4.04 ;
      RECT 80.31 7.215 80.66 12.46 ;
      RECT 80.31 7.215 80.665 7.57 ;
      RECT 72.73 9.325 73.1 9.695 ;
      RECT 72.77 9.005 73.105 9.37 ;
      RECT 72.77 9.005 73.155 9.315 ;
      RECT 72.77 9.005 75.56 9.31 ;
      RECT 75.255 4.145 75.56 9.31 ;
      RECT 75.22 4.145 75.59 4.515 ;
      RECT 70.59 3.145 70.92 4.04 ;
      RECT 69.71 3.31 70.04 4.04 ;
      RECT 70.585 3.145 70.955 3.945 ;
      RECT 73.75 3.145 74.08 3.875 ;
      RECT 73.71 3.03 73.89 3.68 ;
      RECT 69.72 3.145 74.08 3.515 ;
      RECT 70.21 4.83 70.54 5.16 ;
      RECT 69.005 4.845 70.54 5.145 ;
      RECT 69.005 3.725 69.305 5.145 ;
      RECT 68.75 3.71 69.08 4.04 ;
      RECT 64.525 7.215 64.875 12.46 ;
      RECT 64.525 7.215 64.88 7.57 ;
      RECT 56.945 9.325 57.315 9.695 ;
      RECT 56.985 9.005 57.32 9.37 ;
      RECT 56.985 9.005 57.37 9.315 ;
      RECT 56.985 9.005 59.775 9.31 ;
      RECT 59.47 4.145 59.775 9.31 ;
      RECT 59.435 4.145 59.805 4.515 ;
      RECT 54.805 3.145 55.135 4.04 ;
      RECT 53.925 3.31 54.255 4.04 ;
      RECT 54.8 3.145 55.17 3.945 ;
      RECT 57.965 3.145 58.295 3.875 ;
      RECT 57.925 3.03 58.105 3.68 ;
      RECT 53.935 3.145 58.295 3.515 ;
      RECT 54.425 4.83 54.755 5.16 ;
      RECT 53.22 4.845 54.755 5.145 ;
      RECT 53.22 3.725 53.52 5.145 ;
      RECT 52.965 3.71 53.295 4.04 ;
      RECT 48.75 7.215 49.1 12.46 ;
      RECT 48.75 7.215 49.105 7.57 ;
      RECT 41.17 9.325 41.54 9.695 ;
      RECT 41.21 9.005 41.545 9.37 ;
      RECT 41.21 9.005 41.595 9.315 ;
      RECT 41.21 9.005 44 9.31 ;
      RECT 43.695 4.145 44 9.31 ;
      RECT 43.66 4.145 44.03 4.515 ;
      RECT 39.03 3.145 39.36 4.04 ;
      RECT 38.15 3.31 38.48 4.04 ;
      RECT 39.025 3.145 39.395 3.945 ;
      RECT 42.19 3.145 42.52 3.875 ;
      RECT 42.15 3.03 42.33 3.68 ;
      RECT 38.16 3.145 42.52 3.515 ;
      RECT 38.65 4.83 38.98 5.16 ;
      RECT 37.445 4.845 38.98 5.145 ;
      RECT 37.445 3.725 37.745 5.145 ;
      RECT 37.19 3.71 37.52 4.04 ;
      RECT 32.97 7.215 33.32 12.46 ;
      RECT 32.97 7.215 33.325 7.57 ;
      RECT 25.39 9.325 25.76 9.695 ;
      RECT 25.43 9.005 25.765 9.37 ;
      RECT 25.43 9.005 25.815 9.315 ;
      RECT 25.43 9.005 28.22 9.31 ;
      RECT 27.915 4.145 28.22 9.31 ;
      RECT 27.88 4.145 28.25 4.515 ;
      RECT 23.25 3.145 23.58 4.04 ;
      RECT 22.37 3.31 22.7 4.04 ;
      RECT 23.245 3.145 23.615 3.945 ;
      RECT 26.41 3.145 26.74 3.875 ;
      RECT 26.37 3.03 26.55 3.68 ;
      RECT 22.38 3.145 26.74 3.515 ;
      RECT 22.87 4.83 23.2 5.16 ;
      RECT 21.665 4.845 23.2 5.145 ;
      RECT 21.665 3.725 21.965 5.145 ;
      RECT 21.41 3.71 21.74 4.04 ;
      RECT 87.935 3.87 88.265 4.6 ;
      RECT 83.815 3.71 84.145 4.44 ;
      RECT 82.815 3.15 83.145 3.88 ;
      RECT 81.375 3.87 81.705 4.6 ;
      RECT 72.15 3.87 72.48 4.6 ;
      RECT 68.03 3.71 68.36 4.44 ;
      RECT 67.03 3.15 67.36 3.88 ;
      RECT 65.59 3.87 65.92 4.6 ;
      RECT 56.365 3.87 56.695 4.6 ;
      RECT 52.245 3.71 52.575 4.44 ;
      RECT 51.245 3.15 51.575 3.88 ;
      RECT 49.805 3.87 50.135 4.6 ;
      RECT 40.59 3.87 40.92 4.6 ;
      RECT 36.47 3.71 36.8 4.44 ;
      RECT 35.47 3.15 35.8 3.88 ;
      RECT 34.03 3.87 34.36 4.6 ;
      RECT 24.81 3.87 25.14 4.6 ;
      RECT 20.69 3.71 21.02 4.44 ;
      RECT 19.69 3.15 20.02 3.88 ;
      RECT 18.25 3.87 18.58 4.6 ;
    LAYER via2 ;
      RECT 96.18 7.3 96.38 7.5 ;
      RECT 91.09 4.23 91.29 4.43 ;
      RECT 89.6 3.61 89.8 3.81 ;
      RECT 88.6 9.41 88.8 9.61 ;
      RECT 88 4.335 88.2 4.535 ;
      RECT 86.44 3.775 86.64 3.975 ;
      RECT 86.06 4.895 86.26 5.095 ;
      RECT 85.56 3.775 85.76 3.975 ;
      RECT 84.6 3.775 84.8 3.975 ;
      RECT 83.88 3.775 84.08 3.975 ;
      RECT 82.88 3.215 83.08 3.415 ;
      RECT 81.44 4.335 81.64 4.535 ;
      RECT 80.395 7.3 80.595 7.5 ;
      RECT 75.305 4.23 75.505 4.43 ;
      RECT 73.815 3.61 74.015 3.81 ;
      RECT 72.815 9.41 73.015 9.61 ;
      RECT 72.215 4.335 72.415 4.535 ;
      RECT 70.655 3.775 70.855 3.975 ;
      RECT 70.275 4.895 70.475 5.095 ;
      RECT 69.775 3.775 69.975 3.975 ;
      RECT 68.815 3.775 69.015 3.975 ;
      RECT 68.095 3.775 68.295 3.975 ;
      RECT 67.095 3.215 67.295 3.415 ;
      RECT 65.655 4.335 65.855 4.535 ;
      RECT 64.61 7.3 64.81 7.5 ;
      RECT 59.52 4.23 59.72 4.43 ;
      RECT 58.03 3.61 58.23 3.81 ;
      RECT 57.03 9.41 57.23 9.61 ;
      RECT 56.43 4.335 56.63 4.535 ;
      RECT 54.87 3.775 55.07 3.975 ;
      RECT 54.49 4.895 54.69 5.095 ;
      RECT 53.99 3.775 54.19 3.975 ;
      RECT 53.03 3.775 53.23 3.975 ;
      RECT 52.31 3.775 52.51 3.975 ;
      RECT 51.31 3.215 51.51 3.415 ;
      RECT 49.87 4.335 50.07 4.535 ;
      RECT 48.835 7.3 49.035 7.5 ;
      RECT 43.745 4.23 43.945 4.43 ;
      RECT 42.255 3.61 42.455 3.81 ;
      RECT 41.255 9.41 41.455 9.61 ;
      RECT 40.655 4.335 40.855 4.535 ;
      RECT 39.095 3.775 39.295 3.975 ;
      RECT 38.715 4.895 38.915 5.095 ;
      RECT 38.215 3.775 38.415 3.975 ;
      RECT 37.255 3.775 37.455 3.975 ;
      RECT 36.535 3.775 36.735 3.975 ;
      RECT 35.535 3.215 35.735 3.415 ;
      RECT 34.095 4.335 34.295 4.535 ;
      RECT 33.055 7.3 33.255 7.5 ;
      RECT 27.965 4.23 28.165 4.43 ;
      RECT 26.475 3.61 26.675 3.81 ;
      RECT 25.475 9.41 25.675 9.61 ;
      RECT 24.875 4.335 25.075 4.535 ;
      RECT 23.315 3.775 23.515 3.975 ;
      RECT 22.935 4.895 23.135 5.095 ;
      RECT 22.435 3.775 22.635 3.975 ;
      RECT 21.475 3.775 21.675 3.975 ;
      RECT 20.755 3.775 20.955 3.975 ;
      RECT 19.755 3.215 19.955 3.415 ;
      RECT 18.315 4.335 18.515 4.535 ;
    LAYER met2 ;
      RECT 16.23 10.685 96.35 10.855 ;
      RECT 96.18 9.56 96.35 10.855 ;
      RECT 16.23 8.54 16.4 10.855 ;
      RECT 96.15 9.56 96.5 9.91 ;
      RECT 16.165 8.54 16.455 8.89 ;
      RECT 96.14 7.215 96.42 7.585 ;
      RECT 96.095 7.215 96.45 7.57 ;
      RECT 92.99 8.505 93.31 8.83 ;
      RECT 93.02 7.98 93.19 8.83 ;
      RECT 93.02 7.98 93.195 8.33 ;
      RECT 93.02 7.98 93.995 8.155 ;
      RECT 93.82 3.26 93.995 8.155 ;
      RECT 93.765 3.26 94.115 3.61 ;
      RECT 93.79 8.94 94.115 9.265 ;
      RECT 92.675 9.03 94.115 9.2 ;
      RECT 92.675 3.69 92.835 9.2 ;
      RECT 92.99 3.66 93.31 3.98 ;
      RECT 92.675 3.69 93.31 3.86 ;
      RECT 82.76 3.215 83.02 3.475 ;
      RECT 82.815 3.175 83.12 3.455 ;
      RECT 82.815 2.715 82.99 3.475 ;
      RECT 91.33 2.635 91.68 2.985 ;
      RECT 82.815 2.715 91.68 2.89 ;
      RECT 91.005 4.145 91.375 4.515 ;
      RECT 91.09 3.53 91.26 4.515 ;
      RECT 87.11 3.75 87.345 4.01 ;
      RECT 90.255 3.53 90.42 3.79 ;
      RECT 90.16 3.52 90.175 3.79 ;
      RECT 90.255 3.53 91.26 3.71 ;
      RECT 88.76 3.09 88.8 3.23 ;
      RECT 90.175 3.525 90.255 3.79 ;
      RECT 90.12 3.52 90.16 3.756 ;
      RECT 90.106 3.52 90.12 3.756 ;
      RECT 90.02 3.525 90.106 3.758 ;
      RECT 89.975 3.532 90.02 3.76 ;
      RECT 89.945 3.532 89.975 3.762 ;
      RECT 89.92 3.527 89.945 3.764 ;
      RECT 89.89 3.523 89.92 3.773 ;
      RECT 89.88 3.52 89.89 3.785 ;
      RECT 89.875 3.52 89.88 3.793 ;
      RECT 89.87 3.52 89.875 3.798 ;
      RECT 89.86 3.519 89.87 3.808 ;
      RECT 89.855 3.518 89.86 3.818 ;
      RECT 89.84 3.517 89.855 3.823 ;
      RECT 89.812 3.514 89.84 3.85 ;
      RECT 89.726 3.506 89.812 3.85 ;
      RECT 89.64 3.495 89.726 3.85 ;
      RECT 89.6 3.48 89.64 3.85 ;
      RECT 89.56 3.454 89.6 3.85 ;
      RECT 89.555 3.436 89.56 3.662 ;
      RECT 89.545 3.432 89.555 3.652 ;
      RECT 89.53 3.422 89.545 3.639 ;
      RECT 89.51 3.406 89.53 3.624 ;
      RECT 89.495 3.391 89.51 3.609 ;
      RECT 89.485 3.38 89.495 3.599 ;
      RECT 89.46 3.364 89.485 3.588 ;
      RECT 89.455 3.351 89.46 3.578 ;
      RECT 89.45 3.347 89.455 3.573 ;
      RECT 89.395 3.333 89.45 3.551 ;
      RECT 89.356 3.314 89.395 3.515 ;
      RECT 89.27 3.288 89.356 3.468 ;
      RECT 89.266 3.27 89.27 3.434 ;
      RECT 89.18 3.251 89.266 3.412 ;
      RECT 89.175 3.233 89.18 3.39 ;
      RECT 89.17 3.231 89.175 3.388 ;
      RECT 89.16 3.23 89.17 3.383 ;
      RECT 89.1 3.217 89.16 3.369 ;
      RECT 89.055 3.195 89.1 3.348 ;
      RECT 88.995 3.172 89.055 3.327 ;
      RECT 88.931 3.147 88.995 3.302 ;
      RECT 88.845 3.117 88.931 3.271 ;
      RECT 88.83 3.097 88.845 3.25 ;
      RECT 88.8 3.092 88.83 3.241 ;
      RECT 88.747 3.09 88.76 3.23 ;
      RECT 88.661 3.09 88.747 3.232 ;
      RECT 88.575 3.09 88.661 3.234 ;
      RECT 88.555 3.09 88.575 3.238 ;
      RECT 88.51 3.092 88.555 3.249 ;
      RECT 88.47 3.102 88.51 3.265 ;
      RECT 88.466 3.111 88.47 3.273 ;
      RECT 88.38 3.131 88.466 3.289 ;
      RECT 88.37 3.15 88.38 3.307 ;
      RECT 88.365 3.152 88.37 3.31 ;
      RECT 88.355 3.156 88.365 3.313 ;
      RECT 88.335 3.161 88.355 3.323 ;
      RECT 88.305 3.171 88.335 3.343 ;
      RECT 88.3 3.178 88.305 3.357 ;
      RECT 88.29 3.182 88.3 3.364 ;
      RECT 88.275 3.19 88.29 3.375 ;
      RECT 88.265 3.2 88.275 3.386 ;
      RECT 88.255 3.207 88.265 3.394 ;
      RECT 88.23 3.22 88.255 3.409 ;
      RECT 88.166 3.256 88.23 3.448 ;
      RECT 88.08 3.319 88.166 3.512 ;
      RECT 88.045 3.37 88.08 3.565 ;
      RECT 88.04 3.387 88.045 3.582 ;
      RECT 88.025 3.396 88.04 3.589 ;
      RECT 88.005 3.411 88.025 3.603 ;
      RECT 88 3.422 88.005 3.613 ;
      RECT 87.98 3.435 88 3.623 ;
      RECT 87.975 3.445 87.98 3.633 ;
      RECT 87.96 3.45 87.975 3.642 ;
      RECT 87.95 3.46 87.96 3.653 ;
      RECT 87.92 3.477 87.95 3.67 ;
      RECT 87.91 3.495 87.92 3.688 ;
      RECT 87.895 3.506 87.91 3.699 ;
      RECT 87.855 3.53 87.895 3.715 ;
      RECT 87.82 3.564 87.855 3.732 ;
      RECT 87.79 3.587 87.82 3.744 ;
      RECT 87.775 3.597 87.79 3.753 ;
      RECT 87.735 3.607 87.775 3.764 ;
      RECT 87.715 3.618 87.735 3.776 ;
      RECT 87.71 3.622 87.715 3.783 ;
      RECT 87.695 3.626 87.71 3.788 ;
      RECT 87.685 3.631 87.695 3.793 ;
      RECT 87.68 3.634 87.685 3.796 ;
      RECT 87.65 3.64 87.68 3.803 ;
      RECT 87.615 3.65 87.65 3.817 ;
      RECT 87.555 3.665 87.615 3.837 ;
      RECT 87.5 3.685 87.555 3.861 ;
      RECT 87.471 3.7 87.5 3.879 ;
      RECT 87.385 3.72 87.471 3.904 ;
      RECT 87.38 3.735 87.385 3.924 ;
      RECT 87.37 3.738 87.38 3.925 ;
      RECT 87.345 3.745 87.37 4.01 ;
      RECT 80.34 8.94 80.69 9.29 ;
      RECT 89.165 8.895 89.515 9.245 ;
      RECT 80.34 8.97 89.515 9.17 ;
      RECT 87.76 4.98 87.77 5.17 ;
      RECT 86.02 4.855 86.3 5.135 ;
      RECT 89.065 3.795 89.07 4.28 ;
      RECT 88.96 3.795 89.02 4.055 ;
      RECT 89.285 4.765 89.29 4.84 ;
      RECT 89.275 4.632 89.285 4.875 ;
      RECT 89.265 4.467 89.275 4.896 ;
      RECT 89.26 4.337 89.265 4.912 ;
      RECT 89.25 4.227 89.26 4.928 ;
      RECT 89.245 4.126 89.25 4.945 ;
      RECT 89.24 4.108 89.245 4.955 ;
      RECT 89.235 4.09 89.24 4.965 ;
      RECT 89.225 4.065 89.235 4.98 ;
      RECT 89.22 4.045 89.225 4.995 ;
      RECT 89.2 3.795 89.22 5.02 ;
      RECT 89.185 3.795 89.2 5.053 ;
      RECT 89.155 3.795 89.185 5.075 ;
      RECT 89.135 3.795 89.155 5.089 ;
      RECT 89.115 3.795 89.135 4.605 ;
      RECT 89.13 4.672 89.135 5.094 ;
      RECT 89.125 4.702 89.13 5.096 ;
      RECT 89.12 4.715 89.125 5.099 ;
      RECT 89.115 4.725 89.12 5.103 ;
      RECT 89.11 3.795 89.115 4.523 ;
      RECT 89.11 4.735 89.115 5.105 ;
      RECT 89.105 3.795 89.11 4.5 ;
      RECT 89.095 4.757 89.11 5.105 ;
      RECT 89.09 3.795 89.105 4.445 ;
      RECT 89.085 4.782 89.095 5.105 ;
      RECT 89.085 3.795 89.09 4.39 ;
      RECT 89.075 3.795 89.085 4.338 ;
      RECT 89.08 4.795 89.085 5.106 ;
      RECT 89.075 4.807 89.08 5.107 ;
      RECT 89.07 3.795 89.075 4.298 ;
      RECT 89.07 4.82 89.075 5.108 ;
      RECT 89.055 4.835 89.07 5.109 ;
      RECT 89.06 3.795 89.065 4.26 ;
      RECT 89.055 3.795 89.06 4.225 ;
      RECT 89.05 3.795 89.055 4.2 ;
      RECT 89.045 4.862 89.055 5.111 ;
      RECT 89.04 3.795 89.05 4.158 ;
      RECT 89.04 4.88 89.045 5.112 ;
      RECT 89.035 3.795 89.04 4.118 ;
      RECT 89.035 4.887 89.04 5.113 ;
      RECT 89.03 3.795 89.035 4.09 ;
      RECT 89.025 4.905 89.035 5.114 ;
      RECT 89.02 3.795 89.03 4.07 ;
      RECT 89.015 4.925 89.025 5.116 ;
      RECT 89.005 4.942 89.015 5.117 ;
      RECT 88.97 4.965 89.005 5.12 ;
      RECT 88.915 4.983 88.97 5.126 ;
      RECT 88.829 4.991 88.915 5.135 ;
      RECT 88.743 5.002 88.829 5.146 ;
      RECT 88.657 5.012 88.743 5.157 ;
      RECT 88.571 5.022 88.657 5.169 ;
      RECT 88.485 5.032 88.571 5.18 ;
      RECT 88.465 5.038 88.485 5.186 ;
      RECT 88.385 5.04 88.465 5.19 ;
      RECT 88.38 5.039 88.385 5.195 ;
      RECT 88.372 5.038 88.38 5.195 ;
      RECT 88.286 5.034 88.372 5.193 ;
      RECT 88.2 5.026 88.286 5.19 ;
      RECT 88.114 5.017 88.2 5.186 ;
      RECT 88.028 5.009 88.114 5.183 ;
      RECT 87.942 5.001 88.028 5.179 ;
      RECT 87.856 4.992 87.942 5.176 ;
      RECT 87.77 4.984 87.856 5.172 ;
      RECT 87.715 4.977 87.76 5.17 ;
      RECT 87.63 4.97 87.715 5.168 ;
      RECT 87.556 4.962 87.63 5.164 ;
      RECT 87.47 4.954 87.556 5.161 ;
      RECT 87.467 4.95 87.47 5.159 ;
      RECT 87.381 4.946 87.467 5.158 ;
      RECT 87.295 4.938 87.381 5.155 ;
      RECT 87.21 4.933 87.295 5.152 ;
      RECT 87.124 4.93 87.21 5.149 ;
      RECT 87.038 4.928 87.124 5.146 ;
      RECT 86.952 4.925 87.038 5.143 ;
      RECT 86.866 4.922 86.952 5.14 ;
      RECT 86.78 4.919 86.866 5.137 ;
      RECT 86.704 4.917 86.78 5.134 ;
      RECT 86.618 4.914 86.704 5.131 ;
      RECT 86.532 4.911 86.618 5.129 ;
      RECT 86.446 4.909 86.532 5.126 ;
      RECT 86.36 4.906 86.446 5.123 ;
      RECT 86.3 4.897 86.36 5.121 ;
      RECT 88.81 4.515 88.885 4.775 ;
      RECT 88.79 4.495 88.795 4.775 ;
      RECT 88.11 4.28 88.215 4.575 ;
      RECT 82.555 4.255 82.625 4.515 ;
      RECT 88.45 4.13 88.455 4.501 ;
      RECT 88.44 4.185 88.445 4.501 ;
      RECT 88.745 3.355 88.805 3.615 ;
      RECT 88.8 4.51 88.81 4.775 ;
      RECT 88.795 4.5 88.8 4.775 ;
      RECT 88.715 4.447 88.79 4.775 ;
      RECT 88.74 3.355 88.745 3.635 ;
      RECT 88.73 3.355 88.74 3.655 ;
      RECT 88.715 3.355 88.73 3.685 ;
      RECT 88.7 3.355 88.715 3.728 ;
      RECT 88.695 4.39 88.715 4.775 ;
      RECT 88.685 3.355 88.7 3.765 ;
      RECT 88.68 4.37 88.695 4.775 ;
      RECT 88.68 3.355 88.685 3.788 ;
      RECT 88.67 3.355 88.68 3.813 ;
      RECT 88.64 4.337 88.68 4.775 ;
      RECT 88.645 3.355 88.67 3.863 ;
      RECT 88.64 3.355 88.645 3.918 ;
      RECT 88.635 3.355 88.64 3.96 ;
      RECT 88.625 4.3 88.64 4.775 ;
      RECT 88.63 3.355 88.635 4.003 ;
      RECT 88.625 3.355 88.63 4.068 ;
      RECT 88.62 3.355 88.625 4.09 ;
      RECT 88.62 4.288 88.625 4.64 ;
      RECT 88.615 3.355 88.62 4.158 ;
      RECT 88.615 4.28 88.62 4.623 ;
      RECT 88.61 3.355 88.615 4.203 ;
      RECT 88.605 4.262 88.615 4.6 ;
      RECT 88.605 3.355 88.61 4.24 ;
      RECT 88.595 3.355 88.605 4.58 ;
      RECT 88.59 3.355 88.595 4.563 ;
      RECT 88.585 3.355 88.59 4.548 ;
      RECT 88.58 3.355 88.585 4.533 ;
      RECT 88.56 3.355 88.58 4.523 ;
      RECT 88.555 3.355 88.56 4.513 ;
      RECT 88.545 3.355 88.555 4.509 ;
      RECT 88.54 3.632 88.545 4.508 ;
      RECT 88.535 3.655 88.54 4.507 ;
      RECT 88.53 3.685 88.535 4.506 ;
      RECT 88.525 3.712 88.53 4.505 ;
      RECT 88.52 3.74 88.525 4.505 ;
      RECT 88.515 3.767 88.52 4.505 ;
      RECT 88.51 3.787 88.515 4.505 ;
      RECT 88.505 3.815 88.51 4.505 ;
      RECT 88.495 3.857 88.505 4.505 ;
      RECT 88.485 3.902 88.495 4.504 ;
      RECT 88.48 3.955 88.485 4.503 ;
      RECT 88.475 3.987 88.48 4.502 ;
      RECT 88.47 4.007 88.475 4.501 ;
      RECT 88.465 4.045 88.47 4.501 ;
      RECT 88.46 4.067 88.465 4.501 ;
      RECT 88.455 4.092 88.46 4.501 ;
      RECT 88.445 4.157 88.45 4.501 ;
      RECT 88.43 4.217 88.44 4.501 ;
      RECT 88.415 4.227 88.43 4.501 ;
      RECT 88.395 4.237 88.415 4.501 ;
      RECT 88.365 4.242 88.395 4.498 ;
      RECT 88.305 4.252 88.365 4.495 ;
      RECT 88.285 4.261 88.305 4.5 ;
      RECT 88.26 4.267 88.285 4.513 ;
      RECT 88.24 4.272 88.26 4.528 ;
      RECT 88.215 4.277 88.24 4.575 ;
      RECT 88.086 4.279 88.11 4.575 ;
      RECT 88 4.274 88.086 4.575 ;
      RECT 87.96 4.271 88 4.575 ;
      RECT 87.91 4.273 87.96 4.555 ;
      RECT 87.88 4.277 87.91 4.555 ;
      RECT 87.801 4.287 87.88 4.555 ;
      RECT 87.715 4.302 87.801 4.556 ;
      RECT 87.665 4.312 87.715 4.557 ;
      RECT 87.657 4.315 87.665 4.557 ;
      RECT 87.571 4.317 87.657 4.558 ;
      RECT 87.485 4.321 87.571 4.558 ;
      RECT 87.399 4.325 87.485 4.559 ;
      RECT 87.313 4.328 87.399 4.56 ;
      RECT 87.227 4.332 87.313 4.56 ;
      RECT 87.141 4.336 87.227 4.561 ;
      RECT 87.055 4.339 87.141 4.562 ;
      RECT 86.969 4.343 87.055 4.562 ;
      RECT 86.883 4.347 86.969 4.563 ;
      RECT 86.797 4.351 86.883 4.564 ;
      RECT 86.711 4.354 86.797 4.564 ;
      RECT 86.625 4.358 86.711 4.565 ;
      RECT 86.595 4.36 86.625 4.565 ;
      RECT 86.509 4.363 86.595 4.566 ;
      RECT 86.423 4.367 86.509 4.567 ;
      RECT 86.337 4.371 86.423 4.568 ;
      RECT 86.251 4.374 86.337 4.568 ;
      RECT 86.165 4.378 86.251 4.569 ;
      RECT 86.13 4.383 86.165 4.57 ;
      RECT 86.075 4.393 86.13 4.577 ;
      RECT 86.05 4.405 86.075 4.587 ;
      RECT 86.015 4.418 86.05 4.595 ;
      RECT 85.975 4.435 86.015 4.618 ;
      RECT 85.955 4.448 85.975 4.645 ;
      RECT 85.925 4.46 85.955 4.673 ;
      RECT 85.92 4.468 85.925 4.693 ;
      RECT 85.915 4.471 85.92 4.703 ;
      RECT 85.865 4.483 85.915 4.737 ;
      RECT 85.855 4.498 85.865 4.77 ;
      RECT 85.845 4.504 85.855 4.783 ;
      RECT 85.835 4.511 85.845 4.795 ;
      RECT 85.81 4.524 85.835 4.813 ;
      RECT 85.795 4.539 85.81 4.835 ;
      RECT 85.785 4.547 85.795 4.851 ;
      RECT 85.77 4.556 85.785 4.866 ;
      RECT 85.76 4.566 85.77 4.88 ;
      RECT 85.741 4.579 85.76 4.897 ;
      RECT 85.655 4.624 85.741 4.962 ;
      RECT 85.64 4.669 85.655 5.02 ;
      RECT 85.635 4.678 85.64 5.033 ;
      RECT 85.625 4.685 85.635 5.038 ;
      RECT 85.62 4.69 85.625 5.042 ;
      RECT 85.6 4.7 85.62 5.049 ;
      RECT 85.575 4.72 85.6 5.063 ;
      RECT 85.54 4.745 85.575 5.083 ;
      RECT 85.525 4.768 85.54 5.098 ;
      RECT 85.515 4.778 85.525 5.103 ;
      RECT 85.505 4.786 85.515 5.11 ;
      RECT 85.495 4.795 85.505 5.116 ;
      RECT 85.475 4.807 85.495 5.118 ;
      RECT 85.465 4.82 85.475 5.12 ;
      RECT 85.44 4.835 85.465 5.123 ;
      RECT 85.42 4.852 85.44 5.127 ;
      RECT 85.38 4.88 85.42 5.133 ;
      RECT 85.315 4.927 85.38 5.142 ;
      RECT 85.3 4.96 85.315 5.15 ;
      RECT 85.295 4.967 85.3 5.152 ;
      RECT 85.245 4.992 85.295 5.157 ;
      RECT 85.23 5.016 85.245 5.164 ;
      RECT 85.18 5.021 85.23 5.165 ;
      RECT 85.094 5.025 85.18 5.165 ;
      RECT 85.008 5.025 85.094 5.165 ;
      RECT 84.922 5.025 85.008 5.166 ;
      RECT 84.836 5.025 84.922 5.166 ;
      RECT 84.75 5.025 84.836 5.166 ;
      RECT 84.684 5.025 84.75 5.166 ;
      RECT 84.598 5.025 84.684 5.167 ;
      RECT 84.512 5.025 84.598 5.167 ;
      RECT 84.426 5.026 84.512 5.168 ;
      RECT 84.34 5.026 84.426 5.168 ;
      RECT 84.254 5.026 84.34 5.168 ;
      RECT 84.168 5.026 84.254 5.169 ;
      RECT 84.082 5.026 84.168 5.169 ;
      RECT 83.996 5.027 84.082 5.17 ;
      RECT 83.91 5.027 83.996 5.17 ;
      RECT 83.89 5.027 83.91 5.17 ;
      RECT 83.804 5.027 83.89 5.17 ;
      RECT 83.718 5.027 83.804 5.17 ;
      RECT 83.632 5.028 83.718 5.17 ;
      RECT 83.546 5.028 83.632 5.17 ;
      RECT 83.46 5.028 83.546 5.17 ;
      RECT 83.374 5.029 83.46 5.17 ;
      RECT 83.288 5.029 83.374 5.17 ;
      RECT 83.202 5.029 83.288 5.17 ;
      RECT 83.116 5.029 83.202 5.17 ;
      RECT 83.03 5.03 83.116 5.17 ;
      RECT 82.98 5.027 83.03 5.17 ;
      RECT 82.97 5.025 82.98 5.169 ;
      RECT 82.966 5.025 82.97 5.168 ;
      RECT 82.88 5.02 82.966 5.163 ;
      RECT 82.858 5.013 82.88 5.157 ;
      RECT 82.772 5.004 82.858 5.151 ;
      RECT 82.686 4.991 82.772 5.142 ;
      RECT 82.6 4.977 82.686 5.132 ;
      RECT 82.555 4.967 82.6 5.125 ;
      RECT 82.535 4.255 82.555 4.533 ;
      RECT 82.535 4.96 82.555 5.121 ;
      RECT 82.505 4.255 82.535 4.555 ;
      RECT 82.495 4.927 82.535 5.118 ;
      RECT 82.49 4.255 82.505 4.575 ;
      RECT 82.49 4.892 82.495 5.116 ;
      RECT 82.485 4.255 82.49 4.7 ;
      RECT 82.485 4.852 82.49 5.116 ;
      RECT 82.475 4.255 82.485 5.116 ;
      RECT 82.4 4.255 82.475 5.11 ;
      RECT 82.37 4.255 82.4 5.1 ;
      RECT 82.365 4.255 82.37 5.092 ;
      RECT 82.36 4.297 82.365 5.085 ;
      RECT 82.35 4.366 82.36 5.076 ;
      RECT 82.345 4.436 82.35 5.028 ;
      RECT 82.34 4.5 82.345 4.925 ;
      RECT 82.335 4.535 82.34 4.88 ;
      RECT 82.333 4.572 82.335 4.772 ;
      RECT 82.33 4.58 82.333 4.765 ;
      RECT 82.325 4.645 82.33 4.708 ;
      RECT 86.4 3.735 86.68 4.015 ;
      RECT 86.39 3.735 86.68 3.878 ;
      RECT 86.345 3.6 86.605 3.86 ;
      RECT 86.345 3.715 86.66 3.86 ;
      RECT 86.345 3.685 86.655 3.86 ;
      RECT 86.345 3.672 86.645 3.86 ;
      RECT 86.345 3.662 86.64 3.86 ;
      RECT 82.32 3.645 82.58 3.905 ;
      RECT 86.09 3.195 86.35 3.455 ;
      RECT 86.08 3.22 86.35 3.415 ;
      RECT 86.075 3.22 86.08 3.414 ;
      RECT 86.005 3.215 86.075 3.406 ;
      RECT 85.92 3.202 86.005 3.389 ;
      RECT 85.916 3.194 85.92 3.379 ;
      RECT 85.83 3.187 85.916 3.369 ;
      RECT 85.821 3.179 85.83 3.359 ;
      RECT 85.735 3.172 85.821 3.347 ;
      RECT 85.715 3.163 85.735 3.333 ;
      RECT 85.66 3.158 85.715 3.325 ;
      RECT 85.65 3.152 85.66 3.319 ;
      RECT 85.63 3.15 85.65 3.315 ;
      RECT 85.622 3.149 85.63 3.311 ;
      RECT 85.536 3.141 85.622 3.3 ;
      RECT 85.45 3.127 85.536 3.28 ;
      RECT 85.39 3.115 85.45 3.265 ;
      RECT 85.38 3.11 85.39 3.26 ;
      RECT 85.33 3.11 85.38 3.262 ;
      RECT 85.283 3.112 85.33 3.266 ;
      RECT 85.197 3.119 85.283 3.271 ;
      RECT 85.111 3.127 85.197 3.277 ;
      RECT 85.025 3.136 85.111 3.283 ;
      RECT 84.966 3.142 85.025 3.288 ;
      RECT 84.88 3.147 84.966 3.294 ;
      RECT 84.805 3.152 84.88 3.3 ;
      RECT 84.766 3.154 84.805 3.305 ;
      RECT 84.68 3.151 84.766 3.31 ;
      RECT 84.595 3.149 84.68 3.317 ;
      RECT 84.563 3.148 84.595 3.32 ;
      RECT 84.477 3.147 84.563 3.321 ;
      RECT 84.391 3.146 84.477 3.322 ;
      RECT 84.305 3.145 84.391 3.322 ;
      RECT 84.219 3.144 84.305 3.323 ;
      RECT 84.133 3.143 84.219 3.324 ;
      RECT 84.047 3.142 84.133 3.325 ;
      RECT 83.961 3.141 84.047 3.325 ;
      RECT 83.875 3.14 83.961 3.326 ;
      RECT 83.825 3.14 83.875 3.327 ;
      RECT 83.811 3.141 83.825 3.327 ;
      RECT 83.725 3.148 83.811 3.328 ;
      RECT 83.651 3.159 83.725 3.329 ;
      RECT 83.565 3.168 83.651 3.33 ;
      RECT 83.53 3.175 83.565 3.345 ;
      RECT 83.505 3.178 83.53 3.375 ;
      RECT 83.48 3.187 83.505 3.404 ;
      RECT 83.47 3.198 83.48 3.424 ;
      RECT 83.46 3.206 83.47 3.438 ;
      RECT 83.455 3.212 83.46 3.448 ;
      RECT 83.43 3.229 83.455 3.465 ;
      RECT 83.415 3.251 83.43 3.493 ;
      RECT 83.385 3.277 83.415 3.523 ;
      RECT 83.365 3.306 83.385 3.553 ;
      RECT 83.36 3.321 83.365 3.57 ;
      RECT 83.34 3.336 83.36 3.585 ;
      RECT 83.33 3.354 83.34 3.603 ;
      RECT 83.32 3.365 83.33 3.618 ;
      RECT 83.27 3.397 83.32 3.644 ;
      RECT 83.265 3.427 83.27 3.664 ;
      RECT 83.255 3.44 83.265 3.67 ;
      RECT 83.246 3.45 83.255 3.678 ;
      RECT 83.235 3.461 83.246 3.686 ;
      RECT 83.23 3.471 83.235 3.692 ;
      RECT 83.215 3.492 83.23 3.699 ;
      RECT 83.2 3.522 83.215 3.707 ;
      RECT 83.165 3.552 83.2 3.713 ;
      RECT 83.14 3.57 83.165 3.72 ;
      RECT 83.09 3.578 83.14 3.729 ;
      RECT 83.065 3.583 83.09 3.738 ;
      RECT 83.01 3.589 83.065 3.748 ;
      RECT 83.005 3.594 83.01 3.756 ;
      RECT 82.991 3.597 83.005 3.758 ;
      RECT 82.905 3.609 82.991 3.77 ;
      RECT 82.895 3.621 82.905 3.783 ;
      RECT 82.81 3.634 82.895 3.795 ;
      RECT 82.766 3.651 82.81 3.809 ;
      RECT 82.68 3.668 82.766 3.825 ;
      RECT 82.65 3.682 82.68 3.839 ;
      RECT 82.64 3.687 82.65 3.844 ;
      RECT 82.58 3.69 82.64 3.853 ;
      RECT 85.47 3.96 85.73 4.22 ;
      RECT 85.47 3.96 85.75 4.073 ;
      RECT 85.47 3.96 85.775 4.04 ;
      RECT 85.47 3.96 85.78 4.02 ;
      RECT 85.52 3.735 85.8 4.015 ;
      RECT 85.075 4.47 85.335 4.73 ;
      RECT 85.065 4.327 85.26 4.668 ;
      RECT 85.06 4.435 85.275 4.66 ;
      RECT 85.055 4.485 85.335 4.65 ;
      RECT 85.045 4.562 85.335 4.635 ;
      RECT 85.065 4.41 85.275 4.668 ;
      RECT 85.075 4.285 85.26 4.73 ;
      RECT 85.075 4.18 85.24 4.73 ;
      RECT 85.085 4.167 85.24 4.73 ;
      RECT 85.085 4.125 85.23 4.73 ;
      RECT 85.09 4.05 85.23 4.73 ;
      RECT 85.12 3.7 85.23 4.73 ;
      RECT 85.125 3.43 85.25 4.053 ;
      RECT 85.095 4.005 85.25 4.053 ;
      RECT 85.11 3.807 85.23 4.73 ;
      RECT 85.1 3.917 85.25 4.053 ;
      RECT 85.125 3.43 85.265 3.91 ;
      RECT 85.125 3.43 85.285 3.785 ;
      RECT 85.09 3.43 85.35 3.69 ;
      RECT 84.56 3.735 84.84 4.015 ;
      RECT 84.545 3.735 84.84 3.995 ;
      RECT 82.6 4.6 82.86 4.86 ;
      RECT 84.385 4.455 84.645 4.715 ;
      RECT 84.365 4.475 84.645 4.69 ;
      RECT 84.322 4.475 84.365 4.689 ;
      RECT 84.236 4.476 84.322 4.686 ;
      RECT 84.15 4.477 84.236 4.682 ;
      RECT 84.075 4.479 84.15 4.679 ;
      RECT 84.052 4.48 84.075 4.677 ;
      RECT 83.966 4.481 84.052 4.675 ;
      RECT 83.88 4.482 83.966 4.672 ;
      RECT 83.856 4.483 83.88 4.67 ;
      RECT 83.77 4.485 83.856 4.667 ;
      RECT 83.685 4.487 83.77 4.668 ;
      RECT 83.628 4.488 83.685 4.674 ;
      RECT 83.542 4.49 83.628 4.684 ;
      RECT 83.456 4.493 83.542 4.697 ;
      RECT 83.37 4.495 83.456 4.709 ;
      RECT 83.356 4.496 83.37 4.716 ;
      RECT 83.27 4.497 83.356 4.724 ;
      RECT 83.23 4.499 83.27 4.733 ;
      RECT 83.221 4.5 83.23 4.736 ;
      RECT 83.135 4.508 83.221 4.742 ;
      RECT 83.115 4.517 83.135 4.75 ;
      RECT 83.03 4.532 83.115 4.758 ;
      RECT 82.97 4.555 83.03 4.769 ;
      RECT 82.96 4.567 82.97 4.774 ;
      RECT 82.92 4.577 82.96 4.778 ;
      RECT 82.865 4.594 82.92 4.786 ;
      RECT 82.86 4.604 82.865 4.79 ;
      RECT 83.926 3.735 83.985 4.132 ;
      RECT 83.84 3.735 84.045 4.123 ;
      RECT 83.835 3.765 84.045 4.118 ;
      RECT 83.801 3.765 84.045 4.116 ;
      RECT 83.715 3.765 84.045 4.11 ;
      RECT 83.67 3.765 84.065 4.088 ;
      RECT 83.67 3.765 84.085 4.043 ;
      RECT 83.63 3.765 84.085 4.033 ;
      RECT 83.84 3.735 84.12 4.015 ;
      RECT 83.575 3.735 83.835 3.995 ;
      RECT 81.4 4.295 81.68 4.575 ;
      RECT 81.37 4.257 81.625 4.56 ;
      RECT 81.365 4.258 81.625 4.558 ;
      RECT 81.36 4.259 81.625 4.552 ;
      RECT 81.355 4.262 81.625 4.545 ;
      RECT 81.35 4.295 81.68 4.538 ;
      RECT 81.32 4.265 81.625 4.525 ;
      RECT 81.32 4.292 81.645 4.525 ;
      RECT 81.32 4.282 81.64 4.525 ;
      RECT 81.32 4.267 81.635 4.525 ;
      RECT 81.4 4.254 81.615 4.575 ;
      RECT 81.486 4.252 81.615 4.575 ;
      RECT 81.572 4.25 81.6 4.575 ;
      RECT 80.355 7.215 80.635 7.585 ;
      RECT 80.31 7.215 80.665 7.57 ;
      RECT 77.205 8.505 77.525 8.83 ;
      RECT 77.235 7.98 77.405 8.83 ;
      RECT 77.235 7.98 77.41 8.33 ;
      RECT 77.235 7.98 78.21 8.155 ;
      RECT 78.035 3.26 78.21 8.155 ;
      RECT 77.98 3.26 78.33 3.61 ;
      RECT 78.005 8.94 78.33 9.265 ;
      RECT 76.89 9.03 78.33 9.2 ;
      RECT 76.89 3.69 77.05 9.2 ;
      RECT 77.205 3.66 77.525 3.98 ;
      RECT 76.89 3.69 77.525 3.86 ;
      RECT 66.975 3.215 67.235 3.475 ;
      RECT 67.03 3.175 67.335 3.455 ;
      RECT 67.03 2.715 67.205 3.475 ;
      RECT 75.545 2.635 75.895 2.985 ;
      RECT 67.03 2.715 75.895 2.89 ;
      RECT 75.22 4.145 75.59 4.515 ;
      RECT 75.305 3.53 75.475 4.515 ;
      RECT 71.325 3.75 71.56 4.01 ;
      RECT 74.47 3.53 74.635 3.79 ;
      RECT 74.375 3.52 74.39 3.79 ;
      RECT 74.47 3.53 75.475 3.71 ;
      RECT 72.975 3.09 73.015 3.23 ;
      RECT 74.39 3.525 74.47 3.79 ;
      RECT 74.335 3.52 74.375 3.756 ;
      RECT 74.321 3.52 74.335 3.756 ;
      RECT 74.235 3.525 74.321 3.758 ;
      RECT 74.19 3.532 74.235 3.76 ;
      RECT 74.16 3.532 74.19 3.762 ;
      RECT 74.135 3.527 74.16 3.764 ;
      RECT 74.105 3.523 74.135 3.773 ;
      RECT 74.095 3.52 74.105 3.785 ;
      RECT 74.09 3.52 74.095 3.793 ;
      RECT 74.085 3.52 74.09 3.798 ;
      RECT 74.075 3.519 74.085 3.808 ;
      RECT 74.07 3.518 74.075 3.818 ;
      RECT 74.055 3.517 74.07 3.823 ;
      RECT 74.027 3.514 74.055 3.85 ;
      RECT 73.941 3.506 74.027 3.85 ;
      RECT 73.855 3.495 73.941 3.85 ;
      RECT 73.815 3.48 73.855 3.85 ;
      RECT 73.775 3.454 73.815 3.85 ;
      RECT 73.77 3.436 73.775 3.662 ;
      RECT 73.76 3.432 73.77 3.652 ;
      RECT 73.745 3.422 73.76 3.639 ;
      RECT 73.725 3.406 73.745 3.624 ;
      RECT 73.71 3.391 73.725 3.609 ;
      RECT 73.7 3.38 73.71 3.599 ;
      RECT 73.675 3.364 73.7 3.588 ;
      RECT 73.67 3.351 73.675 3.578 ;
      RECT 73.665 3.347 73.67 3.573 ;
      RECT 73.61 3.333 73.665 3.551 ;
      RECT 73.571 3.314 73.61 3.515 ;
      RECT 73.485 3.288 73.571 3.468 ;
      RECT 73.481 3.27 73.485 3.434 ;
      RECT 73.395 3.251 73.481 3.412 ;
      RECT 73.39 3.233 73.395 3.39 ;
      RECT 73.385 3.231 73.39 3.388 ;
      RECT 73.375 3.23 73.385 3.383 ;
      RECT 73.315 3.217 73.375 3.369 ;
      RECT 73.27 3.195 73.315 3.348 ;
      RECT 73.21 3.172 73.27 3.327 ;
      RECT 73.146 3.147 73.21 3.302 ;
      RECT 73.06 3.117 73.146 3.271 ;
      RECT 73.045 3.097 73.06 3.25 ;
      RECT 73.015 3.092 73.045 3.241 ;
      RECT 72.962 3.09 72.975 3.23 ;
      RECT 72.876 3.09 72.962 3.232 ;
      RECT 72.79 3.09 72.876 3.234 ;
      RECT 72.77 3.09 72.79 3.238 ;
      RECT 72.725 3.092 72.77 3.249 ;
      RECT 72.685 3.102 72.725 3.265 ;
      RECT 72.681 3.111 72.685 3.273 ;
      RECT 72.595 3.131 72.681 3.289 ;
      RECT 72.585 3.15 72.595 3.307 ;
      RECT 72.58 3.152 72.585 3.31 ;
      RECT 72.57 3.156 72.58 3.313 ;
      RECT 72.55 3.161 72.57 3.323 ;
      RECT 72.52 3.171 72.55 3.343 ;
      RECT 72.515 3.178 72.52 3.357 ;
      RECT 72.505 3.182 72.515 3.364 ;
      RECT 72.49 3.19 72.505 3.375 ;
      RECT 72.48 3.2 72.49 3.386 ;
      RECT 72.47 3.207 72.48 3.394 ;
      RECT 72.445 3.22 72.47 3.409 ;
      RECT 72.381 3.256 72.445 3.448 ;
      RECT 72.295 3.319 72.381 3.512 ;
      RECT 72.26 3.37 72.295 3.565 ;
      RECT 72.255 3.387 72.26 3.582 ;
      RECT 72.24 3.396 72.255 3.589 ;
      RECT 72.22 3.411 72.24 3.603 ;
      RECT 72.215 3.422 72.22 3.613 ;
      RECT 72.195 3.435 72.215 3.623 ;
      RECT 72.19 3.445 72.195 3.633 ;
      RECT 72.175 3.45 72.19 3.642 ;
      RECT 72.165 3.46 72.175 3.653 ;
      RECT 72.135 3.477 72.165 3.67 ;
      RECT 72.125 3.495 72.135 3.688 ;
      RECT 72.11 3.506 72.125 3.699 ;
      RECT 72.07 3.53 72.11 3.715 ;
      RECT 72.035 3.564 72.07 3.732 ;
      RECT 72.005 3.587 72.035 3.744 ;
      RECT 71.99 3.597 72.005 3.753 ;
      RECT 71.95 3.607 71.99 3.764 ;
      RECT 71.93 3.618 71.95 3.776 ;
      RECT 71.925 3.622 71.93 3.783 ;
      RECT 71.91 3.626 71.925 3.788 ;
      RECT 71.9 3.631 71.91 3.793 ;
      RECT 71.895 3.634 71.9 3.796 ;
      RECT 71.865 3.64 71.895 3.803 ;
      RECT 71.83 3.65 71.865 3.817 ;
      RECT 71.77 3.665 71.83 3.837 ;
      RECT 71.715 3.685 71.77 3.861 ;
      RECT 71.686 3.7 71.715 3.879 ;
      RECT 71.6 3.72 71.686 3.904 ;
      RECT 71.595 3.735 71.6 3.924 ;
      RECT 71.585 3.738 71.595 3.925 ;
      RECT 71.56 3.745 71.585 4.01 ;
      RECT 64.555 8.94 64.905 9.29 ;
      RECT 73.38 8.895 73.73 9.245 ;
      RECT 64.555 8.97 73.73 9.17 ;
      RECT 71.975 4.98 71.985 5.17 ;
      RECT 70.235 4.855 70.515 5.135 ;
      RECT 73.28 3.795 73.285 4.28 ;
      RECT 73.175 3.795 73.235 4.055 ;
      RECT 73.5 4.765 73.505 4.84 ;
      RECT 73.49 4.632 73.5 4.875 ;
      RECT 73.48 4.467 73.49 4.896 ;
      RECT 73.475 4.337 73.48 4.912 ;
      RECT 73.465 4.227 73.475 4.928 ;
      RECT 73.46 4.126 73.465 4.945 ;
      RECT 73.455 4.108 73.46 4.955 ;
      RECT 73.45 4.09 73.455 4.965 ;
      RECT 73.44 4.065 73.45 4.98 ;
      RECT 73.435 4.045 73.44 4.995 ;
      RECT 73.415 3.795 73.435 5.02 ;
      RECT 73.4 3.795 73.415 5.053 ;
      RECT 73.37 3.795 73.4 5.075 ;
      RECT 73.35 3.795 73.37 5.089 ;
      RECT 73.33 3.795 73.35 4.605 ;
      RECT 73.345 4.672 73.35 5.094 ;
      RECT 73.34 4.702 73.345 5.096 ;
      RECT 73.335 4.715 73.34 5.099 ;
      RECT 73.33 4.725 73.335 5.103 ;
      RECT 73.325 3.795 73.33 4.523 ;
      RECT 73.325 4.735 73.33 5.105 ;
      RECT 73.32 3.795 73.325 4.5 ;
      RECT 73.31 4.757 73.325 5.105 ;
      RECT 73.305 3.795 73.32 4.445 ;
      RECT 73.3 4.782 73.31 5.105 ;
      RECT 73.3 3.795 73.305 4.39 ;
      RECT 73.29 3.795 73.3 4.338 ;
      RECT 73.295 4.795 73.3 5.106 ;
      RECT 73.29 4.807 73.295 5.107 ;
      RECT 73.285 3.795 73.29 4.298 ;
      RECT 73.285 4.82 73.29 5.108 ;
      RECT 73.27 4.835 73.285 5.109 ;
      RECT 73.275 3.795 73.28 4.26 ;
      RECT 73.27 3.795 73.275 4.225 ;
      RECT 73.265 3.795 73.27 4.2 ;
      RECT 73.26 4.862 73.27 5.111 ;
      RECT 73.255 3.795 73.265 4.158 ;
      RECT 73.255 4.88 73.26 5.112 ;
      RECT 73.25 3.795 73.255 4.118 ;
      RECT 73.25 4.887 73.255 5.113 ;
      RECT 73.245 3.795 73.25 4.09 ;
      RECT 73.24 4.905 73.25 5.114 ;
      RECT 73.235 3.795 73.245 4.07 ;
      RECT 73.23 4.925 73.24 5.116 ;
      RECT 73.22 4.942 73.23 5.117 ;
      RECT 73.185 4.965 73.22 5.12 ;
      RECT 73.13 4.983 73.185 5.126 ;
      RECT 73.044 4.991 73.13 5.135 ;
      RECT 72.958 5.002 73.044 5.146 ;
      RECT 72.872 5.012 72.958 5.157 ;
      RECT 72.786 5.022 72.872 5.169 ;
      RECT 72.7 5.032 72.786 5.18 ;
      RECT 72.68 5.038 72.7 5.186 ;
      RECT 72.6 5.04 72.68 5.19 ;
      RECT 72.595 5.039 72.6 5.195 ;
      RECT 72.587 5.038 72.595 5.195 ;
      RECT 72.501 5.034 72.587 5.193 ;
      RECT 72.415 5.026 72.501 5.19 ;
      RECT 72.329 5.017 72.415 5.186 ;
      RECT 72.243 5.009 72.329 5.183 ;
      RECT 72.157 5.001 72.243 5.179 ;
      RECT 72.071 4.992 72.157 5.176 ;
      RECT 71.985 4.984 72.071 5.172 ;
      RECT 71.93 4.977 71.975 5.17 ;
      RECT 71.845 4.97 71.93 5.168 ;
      RECT 71.771 4.962 71.845 5.164 ;
      RECT 71.685 4.954 71.771 5.161 ;
      RECT 71.682 4.95 71.685 5.159 ;
      RECT 71.596 4.946 71.682 5.158 ;
      RECT 71.51 4.938 71.596 5.155 ;
      RECT 71.425 4.933 71.51 5.152 ;
      RECT 71.339 4.93 71.425 5.149 ;
      RECT 71.253 4.928 71.339 5.146 ;
      RECT 71.167 4.925 71.253 5.143 ;
      RECT 71.081 4.922 71.167 5.14 ;
      RECT 70.995 4.919 71.081 5.137 ;
      RECT 70.919 4.917 70.995 5.134 ;
      RECT 70.833 4.914 70.919 5.131 ;
      RECT 70.747 4.911 70.833 5.129 ;
      RECT 70.661 4.909 70.747 5.126 ;
      RECT 70.575 4.906 70.661 5.123 ;
      RECT 70.515 4.897 70.575 5.121 ;
      RECT 73.025 4.515 73.1 4.775 ;
      RECT 73.005 4.495 73.01 4.775 ;
      RECT 72.325 4.28 72.43 4.575 ;
      RECT 66.77 4.255 66.84 4.515 ;
      RECT 72.665 4.13 72.67 4.501 ;
      RECT 72.655 4.185 72.66 4.501 ;
      RECT 72.96 3.355 73.02 3.615 ;
      RECT 73.015 4.51 73.025 4.775 ;
      RECT 73.01 4.5 73.015 4.775 ;
      RECT 72.93 4.447 73.005 4.775 ;
      RECT 72.955 3.355 72.96 3.635 ;
      RECT 72.945 3.355 72.955 3.655 ;
      RECT 72.93 3.355 72.945 3.685 ;
      RECT 72.915 3.355 72.93 3.728 ;
      RECT 72.91 4.39 72.93 4.775 ;
      RECT 72.9 3.355 72.915 3.765 ;
      RECT 72.895 4.37 72.91 4.775 ;
      RECT 72.895 3.355 72.9 3.788 ;
      RECT 72.885 3.355 72.895 3.813 ;
      RECT 72.855 4.337 72.895 4.775 ;
      RECT 72.86 3.355 72.885 3.863 ;
      RECT 72.855 3.355 72.86 3.918 ;
      RECT 72.85 3.355 72.855 3.96 ;
      RECT 72.84 4.3 72.855 4.775 ;
      RECT 72.845 3.355 72.85 4.003 ;
      RECT 72.84 3.355 72.845 4.068 ;
      RECT 72.835 3.355 72.84 4.09 ;
      RECT 72.835 4.288 72.84 4.64 ;
      RECT 72.83 3.355 72.835 4.158 ;
      RECT 72.83 4.28 72.835 4.623 ;
      RECT 72.825 3.355 72.83 4.203 ;
      RECT 72.82 4.262 72.83 4.6 ;
      RECT 72.82 3.355 72.825 4.24 ;
      RECT 72.81 3.355 72.82 4.58 ;
      RECT 72.805 3.355 72.81 4.563 ;
      RECT 72.8 3.355 72.805 4.548 ;
      RECT 72.795 3.355 72.8 4.533 ;
      RECT 72.775 3.355 72.795 4.523 ;
      RECT 72.77 3.355 72.775 4.513 ;
      RECT 72.76 3.355 72.77 4.509 ;
      RECT 72.755 3.632 72.76 4.508 ;
      RECT 72.75 3.655 72.755 4.507 ;
      RECT 72.745 3.685 72.75 4.506 ;
      RECT 72.74 3.712 72.745 4.505 ;
      RECT 72.735 3.74 72.74 4.505 ;
      RECT 72.73 3.767 72.735 4.505 ;
      RECT 72.725 3.787 72.73 4.505 ;
      RECT 72.72 3.815 72.725 4.505 ;
      RECT 72.71 3.857 72.72 4.505 ;
      RECT 72.7 3.902 72.71 4.504 ;
      RECT 72.695 3.955 72.7 4.503 ;
      RECT 72.69 3.987 72.695 4.502 ;
      RECT 72.685 4.007 72.69 4.501 ;
      RECT 72.68 4.045 72.685 4.501 ;
      RECT 72.675 4.067 72.68 4.501 ;
      RECT 72.67 4.092 72.675 4.501 ;
      RECT 72.66 4.157 72.665 4.501 ;
      RECT 72.645 4.217 72.655 4.501 ;
      RECT 72.63 4.227 72.645 4.501 ;
      RECT 72.61 4.237 72.63 4.501 ;
      RECT 72.58 4.242 72.61 4.498 ;
      RECT 72.52 4.252 72.58 4.495 ;
      RECT 72.5 4.261 72.52 4.5 ;
      RECT 72.475 4.267 72.5 4.513 ;
      RECT 72.455 4.272 72.475 4.528 ;
      RECT 72.43 4.277 72.455 4.575 ;
      RECT 72.301 4.279 72.325 4.575 ;
      RECT 72.215 4.274 72.301 4.575 ;
      RECT 72.175 4.271 72.215 4.575 ;
      RECT 72.125 4.273 72.175 4.555 ;
      RECT 72.095 4.277 72.125 4.555 ;
      RECT 72.016 4.287 72.095 4.555 ;
      RECT 71.93 4.302 72.016 4.556 ;
      RECT 71.88 4.312 71.93 4.557 ;
      RECT 71.872 4.315 71.88 4.557 ;
      RECT 71.786 4.317 71.872 4.558 ;
      RECT 71.7 4.321 71.786 4.558 ;
      RECT 71.614 4.325 71.7 4.559 ;
      RECT 71.528 4.328 71.614 4.56 ;
      RECT 71.442 4.332 71.528 4.56 ;
      RECT 71.356 4.336 71.442 4.561 ;
      RECT 71.27 4.339 71.356 4.562 ;
      RECT 71.184 4.343 71.27 4.562 ;
      RECT 71.098 4.347 71.184 4.563 ;
      RECT 71.012 4.351 71.098 4.564 ;
      RECT 70.926 4.354 71.012 4.564 ;
      RECT 70.84 4.358 70.926 4.565 ;
      RECT 70.81 4.36 70.84 4.565 ;
      RECT 70.724 4.363 70.81 4.566 ;
      RECT 70.638 4.367 70.724 4.567 ;
      RECT 70.552 4.371 70.638 4.568 ;
      RECT 70.466 4.374 70.552 4.568 ;
      RECT 70.38 4.378 70.466 4.569 ;
      RECT 70.345 4.383 70.38 4.57 ;
      RECT 70.29 4.393 70.345 4.577 ;
      RECT 70.265 4.405 70.29 4.587 ;
      RECT 70.23 4.418 70.265 4.595 ;
      RECT 70.19 4.435 70.23 4.618 ;
      RECT 70.17 4.448 70.19 4.645 ;
      RECT 70.14 4.46 70.17 4.673 ;
      RECT 70.135 4.468 70.14 4.693 ;
      RECT 70.13 4.471 70.135 4.703 ;
      RECT 70.08 4.483 70.13 4.737 ;
      RECT 70.07 4.498 70.08 4.77 ;
      RECT 70.06 4.504 70.07 4.783 ;
      RECT 70.05 4.511 70.06 4.795 ;
      RECT 70.025 4.524 70.05 4.813 ;
      RECT 70.01 4.539 70.025 4.835 ;
      RECT 70 4.547 70.01 4.851 ;
      RECT 69.985 4.556 70 4.866 ;
      RECT 69.975 4.566 69.985 4.88 ;
      RECT 69.956 4.579 69.975 4.897 ;
      RECT 69.87 4.624 69.956 4.962 ;
      RECT 69.855 4.669 69.87 5.02 ;
      RECT 69.85 4.678 69.855 5.033 ;
      RECT 69.84 4.685 69.85 5.038 ;
      RECT 69.835 4.69 69.84 5.042 ;
      RECT 69.815 4.7 69.835 5.049 ;
      RECT 69.79 4.72 69.815 5.063 ;
      RECT 69.755 4.745 69.79 5.083 ;
      RECT 69.74 4.768 69.755 5.098 ;
      RECT 69.73 4.778 69.74 5.103 ;
      RECT 69.72 4.786 69.73 5.11 ;
      RECT 69.71 4.795 69.72 5.116 ;
      RECT 69.69 4.807 69.71 5.118 ;
      RECT 69.68 4.82 69.69 5.12 ;
      RECT 69.655 4.835 69.68 5.123 ;
      RECT 69.635 4.852 69.655 5.127 ;
      RECT 69.595 4.88 69.635 5.133 ;
      RECT 69.53 4.927 69.595 5.142 ;
      RECT 69.515 4.96 69.53 5.15 ;
      RECT 69.51 4.967 69.515 5.152 ;
      RECT 69.46 4.992 69.51 5.157 ;
      RECT 69.445 5.016 69.46 5.164 ;
      RECT 69.395 5.021 69.445 5.165 ;
      RECT 69.309 5.025 69.395 5.165 ;
      RECT 69.223 5.025 69.309 5.165 ;
      RECT 69.137 5.025 69.223 5.166 ;
      RECT 69.051 5.025 69.137 5.166 ;
      RECT 68.965 5.025 69.051 5.166 ;
      RECT 68.899 5.025 68.965 5.166 ;
      RECT 68.813 5.025 68.899 5.167 ;
      RECT 68.727 5.025 68.813 5.167 ;
      RECT 68.641 5.026 68.727 5.168 ;
      RECT 68.555 5.026 68.641 5.168 ;
      RECT 68.469 5.026 68.555 5.168 ;
      RECT 68.383 5.026 68.469 5.169 ;
      RECT 68.297 5.026 68.383 5.169 ;
      RECT 68.211 5.027 68.297 5.17 ;
      RECT 68.125 5.027 68.211 5.17 ;
      RECT 68.105 5.027 68.125 5.17 ;
      RECT 68.019 5.027 68.105 5.17 ;
      RECT 67.933 5.027 68.019 5.17 ;
      RECT 67.847 5.028 67.933 5.17 ;
      RECT 67.761 5.028 67.847 5.17 ;
      RECT 67.675 5.028 67.761 5.17 ;
      RECT 67.589 5.029 67.675 5.17 ;
      RECT 67.503 5.029 67.589 5.17 ;
      RECT 67.417 5.029 67.503 5.17 ;
      RECT 67.331 5.029 67.417 5.17 ;
      RECT 67.245 5.03 67.331 5.17 ;
      RECT 67.195 5.027 67.245 5.17 ;
      RECT 67.185 5.025 67.195 5.169 ;
      RECT 67.181 5.025 67.185 5.168 ;
      RECT 67.095 5.02 67.181 5.163 ;
      RECT 67.073 5.013 67.095 5.157 ;
      RECT 66.987 5.004 67.073 5.151 ;
      RECT 66.901 4.991 66.987 5.142 ;
      RECT 66.815 4.977 66.901 5.132 ;
      RECT 66.77 4.967 66.815 5.125 ;
      RECT 66.75 4.255 66.77 4.533 ;
      RECT 66.75 4.96 66.77 5.121 ;
      RECT 66.72 4.255 66.75 4.555 ;
      RECT 66.71 4.927 66.75 5.118 ;
      RECT 66.705 4.255 66.72 4.575 ;
      RECT 66.705 4.892 66.71 5.116 ;
      RECT 66.7 4.255 66.705 4.7 ;
      RECT 66.7 4.852 66.705 5.116 ;
      RECT 66.69 4.255 66.7 5.116 ;
      RECT 66.615 4.255 66.69 5.11 ;
      RECT 66.585 4.255 66.615 5.1 ;
      RECT 66.58 4.255 66.585 5.092 ;
      RECT 66.575 4.297 66.58 5.085 ;
      RECT 66.565 4.366 66.575 5.076 ;
      RECT 66.56 4.436 66.565 5.028 ;
      RECT 66.555 4.5 66.56 4.925 ;
      RECT 66.55 4.535 66.555 4.88 ;
      RECT 66.548 4.572 66.55 4.772 ;
      RECT 66.545 4.58 66.548 4.765 ;
      RECT 66.54 4.645 66.545 4.708 ;
      RECT 70.615 3.735 70.895 4.015 ;
      RECT 70.605 3.735 70.895 3.878 ;
      RECT 70.56 3.6 70.82 3.86 ;
      RECT 70.56 3.715 70.875 3.86 ;
      RECT 70.56 3.685 70.87 3.86 ;
      RECT 70.56 3.672 70.86 3.86 ;
      RECT 70.56 3.662 70.855 3.86 ;
      RECT 66.535 3.645 66.795 3.905 ;
      RECT 70.305 3.195 70.565 3.455 ;
      RECT 70.295 3.22 70.565 3.415 ;
      RECT 70.29 3.22 70.295 3.414 ;
      RECT 70.22 3.215 70.29 3.406 ;
      RECT 70.135 3.202 70.22 3.389 ;
      RECT 70.131 3.194 70.135 3.379 ;
      RECT 70.045 3.187 70.131 3.369 ;
      RECT 70.036 3.179 70.045 3.359 ;
      RECT 69.95 3.172 70.036 3.347 ;
      RECT 69.93 3.163 69.95 3.333 ;
      RECT 69.875 3.158 69.93 3.325 ;
      RECT 69.865 3.152 69.875 3.319 ;
      RECT 69.845 3.15 69.865 3.315 ;
      RECT 69.837 3.149 69.845 3.311 ;
      RECT 69.751 3.141 69.837 3.3 ;
      RECT 69.665 3.127 69.751 3.28 ;
      RECT 69.605 3.115 69.665 3.265 ;
      RECT 69.595 3.11 69.605 3.26 ;
      RECT 69.545 3.11 69.595 3.262 ;
      RECT 69.498 3.112 69.545 3.266 ;
      RECT 69.412 3.119 69.498 3.271 ;
      RECT 69.326 3.127 69.412 3.277 ;
      RECT 69.24 3.136 69.326 3.283 ;
      RECT 69.181 3.142 69.24 3.288 ;
      RECT 69.095 3.147 69.181 3.294 ;
      RECT 69.02 3.152 69.095 3.3 ;
      RECT 68.981 3.154 69.02 3.305 ;
      RECT 68.895 3.151 68.981 3.31 ;
      RECT 68.81 3.149 68.895 3.317 ;
      RECT 68.778 3.148 68.81 3.32 ;
      RECT 68.692 3.147 68.778 3.321 ;
      RECT 68.606 3.146 68.692 3.322 ;
      RECT 68.52 3.145 68.606 3.322 ;
      RECT 68.434 3.144 68.52 3.323 ;
      RECT 68.348 3.143 68.434 3.324 ;
      RECT 68.262 3.142 68.348 3.325 ;
      RECT 68.176 3.141 68.262 3.325 ;
      RECT 68.09 3.14 68.176 3.326 ;
      RECT 68.04 3.14 68.09 3.327 ;
      RECT 68.026 3.141 68.04 3.327 ;
      RECT 67.94 3.148 68.026 3.328 ;
      RECT 67.866 3.159 67.94 3.329 ;
      RECT 67.78 3.168 67.866 3.33 ;
      RECT 67.745 3.175 67.78 3.345 ;
      RECT 67.72 3.178 67.745 3.375 ;
      RECT 67.695 3.187 67.72 3.404 ;
      RECT 67.685 3.198 67.695 3.424 ;
      RECT 67.675 3.206 67.685 3.438 ;
      RECT 67.67 3.212 67.675 3.448 ;
      RECT 67.645 3.229 67.67 3.465 ;
      RECT 67.63 3.251 67.645 3.493 ;
      RECT 67.6 3.277 67.63 3.523 ;
      RECT 67.58 3.306 67.6 3.553 ;
      RECT 67.575 3.321 67.58 3.57 ;
      RECT 67.555 3.336 67.575 3.585 ;
      RECT 67.545 3.354 67.555 3.603 ;
      RECT 67.535 3.365 67.545 3.618 ;
      RECT 67.485 3.397 67.535 3.644 ;
      RECT 67.48 3.427 67.485 3.664 ;
      RECT 67.47 3.44 67.48 3.67 ;
      RECT 67.461 3.45 67.47 3.678 ;
      RECT 67.45 3.461 67.461 3.686 ;
      RECT 67.445 3.471 67.45 3.692 ;
      RECT 67.43 3.492 67.445 3.699 ;
      RECT 67.415 3.522 67.43 3.707 ;
      RECT 67.38 3.552 67.415 3.713 ;
      RECT 67.355 3.57 67.38 3.72 ;
      RECT 67.305 3.578 67.355 3.729 ;
      RECT 67.28 3.583 67.305 3.738 ;
      RECT 67.225 3.589 67.28 3.748 ;
      RECT 67.22 3.594 67.225 3.756 ;
      RECT 67.206 3.597 67.22 3.758 ;
      RECT 67.12 3.609 67.206 3.77 ;
      RECT 67.11 3.621 67.12 3.783 ;
      RECT 67.025 3.634 67.11 3.795 ;
      RECT 66.981 3.651 67.025 3.809 ;
      RECT 66.895 3.668 66.981 3.825 ;
      RECT 66.865 3.682 66.895 3.839 ;
      RECT 66.855 3.687 66.865 3.844 ;
      RECT 66.795 3.69 66.855 3.853 ;
      RECT 69.685 3.96 69.945 4.22 ;
      RECT 69.685 3.96 69.965 4.073 ;
      RECT 69.685 3.96 69.99 4.04 ;
      RECT 69.685 3.96 69.995 4.02 ;
      RECT 69.735 3.735 70.015 4.015 ;
      RECT 69.29 4.47 69.55 4.73 ;
      RECT 69.28 4.327 69.475 4.668 ;
      RECT 69.275 4.435 69.49 4.66 ;
      RECT 69.27 4.485 69.55 4.65 ;
      RECT 69.26 4.562 69.55 4.635 ;
      RECT 69.28 4.41 69.49 4.668 ;
      RECT 69.29 4.285 69.475 4.73 ;
      RECT 69.29 4.18 69.455 4.73 ;
      RECT 69.3 4.167 69.455 4.73 ;
      RECT 69.3 4.125 69.445 4.73 ;
      RECT 69.305 4.05 69.445 4.73 ;
      RECT 69.335 3.7 69.445 4.73 ;
      RECT 69.34 3.43 69.465 4.053 ;
      RECT 69.31 4.005 69.465 4.053 ;
      RECT 69.325 3.807 69.445 4.73 ;
      RECT 69.315 3.917 69.465 4.053 ;
      RECT 69.34 3.43 69.48 3.91 ;
      RECT 69.34 3.43 69.5 3.785 ;
      RECT 69.305 3.43 69.565 3.69 ;
      RECT 68.775 3.735 69.055 4.015 ;
      RECT 68.76 3.735 69.055 3.995 ;
      RECT 66.815 4.6 67.075 4.86 ;
      RECT 68.6 4.455 68.86 4.715 ;
      RECT 68.58 4.475 68.86 4.69 ;
      RECT 68.537 4.475 68.58 4.689 ;
      RECT 68.451 4.476 68.537 4.686 ;
      RECT 68.365 4.477 68.451 4.682 ;
      RECT 68.29 4.479 68.365 4.679 ;
      RECT 68.267 4.48 68.29 4.677 ;
      RECT 68.181 4.481 68.267 4.675 ;
      RECT 68.095 4.482 68.181 4.672 ;
      RECT 68.071 4.483 68.095 4.67 ;
      RECT 67.985 4.485 68.071 4.667 ;
      RECT 67.9 4.487 67.985 4.668 ;
      RECT 67.843 4.488 67.9 4.674 ;
      RECT 67.757 4.49 67.843 4.684 ;
      RECT 67.671 4.493 67.757 4.697 ;
      RECT 67.585 4.495 67.671 4.709 ;
      RECT 67.571 4.496 67.585 4.716 ;
      RECT 67.485 4.497 67.571 4.724 ;
      RECT 67.445 4.499 67.485 4.733 ;
      RECT 67.436 4.5 67.445 4.736 ;
      RECT 67.35 4.508 67.436 4.742 ;
      RECT 67.33 4.517 67.35 4.75 ;
      RECT 67.245 4.532 67.33 4.758 ;
      RECT 67.185 4.555 67.245 4.769 ;
      RECT 67.175 4.567 67.185 4.774 ;
      RECT 67.135 4.577 67.175 4.778 ;
      RECT 67.08 4.594 67.135 4.786 ;
      RECT 67.075 4.604 67.08 4.79 ;
      RECT 68.141 3.735 68.2 4.132 ;
      RECT 68.055 3.735 68.26 4.123 ;
      RECT 68.05 3.765 68.26 4.118 ;
      RECT 68.016 3.765 68.26 4.116 ;
      RECT 67.93 3.765 68.26 4.11 ;
      RECT 67.885 3.765 68.28 4.088 ;
      RECT 67.885 3.765 68.3 4.043 ;
      RECT 67.845 3.765 68.3 4.033 ;
      RECT 68.055 3.735 68.335 4.015 ;
      RECT 67.79 3.735 68.05 3.995 ;
      RECT 65.615 4.295 65.895 4.575 ;
      RECT 65.585 4.257 65.84 4.56 ;
      RECT 65.58 4.258 65.84 4.558 ;
      RECT 65.575 4.259 65.84 4.552 ;
      RECT 65.57 4.262 65.84 4.545 ;
      RECT 65.565 4.295 65.895 4.538 ;
      RECT 65.535 4.265 65.84 4.525 ;
      RECT 65.535 4.292 65.86 4.525 ;
      RECT 65.535 4.282 65.855 4.525 ;
      RECT 65.535 4.267 65.85 4.525 ;
      RECT 65.615 4.254 65.83 4.575 ;
      RECT 65.701 4.252 65.83 4.575 ;
      RECT 65.787 4.25 65.815 4.575 ;
      RECT 64.57 7.215 64.85 7.585 ;
      RECT 64.525 7.215 64.88 7.57 ;
      RECT 61.42 8.505 61.74 8.83 ;
      RECT 61.45 7.98 61.62 8.83 ;
      RECT 61.45 7.98 61.625 8.33 ;
      RECT 61.45 7.98 62.425 8.155 ;
      RECT 62.25 3.26 62.425 8.155 ;
      RECT 62.195 3.26 62.545 3.61 ;
      RECT 62.22 8.94 62.545 9.265 ;
      RECT 61.105 9.03 62.545 9.2 ;
      RECT 61.105 3.69 61.265 9.2 ;
      RECT 61.42 3.66 61.74 3.98 ;
      RECT 61.105 3.69 61.74 3.86 ;
      RECT 51.19 3.215 51.45 3.475 ;
      RECT 51.245 3.175 51.55 3.455 ;
      RECT 51.245 2.715 51.42 3.475 ;
      RECT 59.76 2.635 60.11 2.985 ;
      RECT 51.245 2.715 60.11 2.89 ;
      RECT 59.435 4.145 59.805 4.515 ;
      RECT 59.52 3.53 59.69 4.515 ;
      RECT 55.54 3.75 55.775 4.01 ;
      RECT 58.685 3.53 58.85 3.79 ;
      RECT 58.59 3.52 58.605 3.79 ;
      RECT 58.685 3.53 59.69 3.71 ;
      RECT 57.19 3.09 57.23 3.23 ;
      RECT 58.605 3.525 58.685 3.79 ;
      RECT 58.55 3.52 58.59 3.756 ;
      RECT 58.536 3.52 58.55 3.756 ;
      RECT 58.45 3.525 58.536 3.758 ;
      RECT 58.405 3.532 58.45 3.76 ;
      RECT 58.375 3.532 58.405 3.762 ;
      RECT 58.35 3.527 58.375 3.764 ;
      RECT 58.32 3.523 58.35 3.773 ;
      RECT 58.31 3.52 58.32 3.785 ;
      RECT 58.305 3.52 58.31 3.793 ;
      RECT 58.3 3.52 58.305 3.798 ;
      RECT 58.29 3.519 58.3 3.808 ;
      RECT 58.285 3.518 58.29 3.818 ;
      RECT 58.27 3.517 58.285 3.823 ;
      RECT 58.242 3.514 58.27 3.85 ;
      RECT 58.156 3.506 58.242 3.85 ;
      RECT 58.07 3.495 58.156 3.85 ;
      RECT 58.03 3.48 58.07 3.85 ;
      RECT 57.99 3.454 58.03 3.85 ;
      RECT 57.985 3.436 57.99 3.662 ;
      RECT 57.975 3.432 57.985 3.652 ;
      RECT 57.96 3.422 57.975 3.639 ;
      RECT 57.94 3.406 57.96 3.624 ;
      RECT 57.925 3.391 57.94 3.609 ;
      RECT 57.915 3.38 57.925 3.599 ;
      RECT 57.89 3.364 57.915 3.588 ;
      RECT 57.885 3.351 57.89 3.578 ;
      RECT 57.88 3.347 57.885 3.573 ;
      RECT 57.825 3.333 57.88 3.551 ;
      RECT 57.786 3.314 57.825 3.515 ;
      RECT 57.7 3.288 57.786 3.468 ;
      RECT 57.696 3.27 57.7 3.434 ;
      RECT 57.61 3.251 57.696 3.412 ;
      RECT 57.605 3.233 57.61 3.39 ;
      RECT 57.6 3.231 57.605 3.388 ;
      RECT 57.59 3.23 57.6 3.383 ;
      RECT 57.53 3.217 57.59 3.369 ;
      RECT 57.485 3.195 57.53 3.348 ;
      RECT 57.425 3.172 57.485 3.327 ;
      RECT 57.361 3.147 57.425 3.302 ;
      RECT 57.275 3.117 57.361 3.271 ;
      RECT 57.26 3.097 57.275 3.25 ;
      RECT 57.23 3.092 57.26 3.241 ;
      RECT 57.177 3.09 57.19 3.23 ;
      RECT 57.091 3.09 57.177 3.232 ;
      RECT 57.005 3.09 57.091 3.234 ;
      RECT 56.985 3.09 57.005 3.238 ;
      RECT 56.94 3.092 56.985 3.249 ;
      RECT 56.9 3.102 56.94 3.265 ;
      RECT 56.896 3.111 56.9 3.273 ;
      RECT 56.81 3.131 56.896 3.289 ;
      RECT 56.8 3.15 56.81 3.307 ;
      RECT 56.795 3.152 56.8 3.31 ;
      RECT 56.785 3.156 56.795 3.313 ;
      RECT 56.765 3.161 56.785 3.323 ;
      RECT 56.735 3.171 56.765 3.343 ;
      RECT 56.73 3.178 56.735 3.357 ;
      RECT 56.72 3.182 56.73 3.364 ;
      RECT 56.705 3.19 56.72 3.375 ;
      RECT 56.695 3.2 56.705 3.386 ;
      RECT 56.685 3.207 56.695 3.394 ;
      RECT 56.66 3.22 56.685 3.409 ;
      RECT 56.596 3.256 56.66 3.448 ;
      RECT 56.51 3.319 56.596 3.512 ;
      RECT 56.475 3.37 56.51 3.565 ;
      RECT 56.47 3.387 56.475 3.582 ;
      RECT 56.455 3.396 56.47 3.589 ;
      RECT 56.435 3.411 56.455 3.603 ;
      RECT 56.43 3.422 56.435 3.613 ;
      RECT 56.41 3.435 56.43 3.623 ;
      RECT 56.405 3.445 56.41 3.633 ;
      RECT 56.39 3.45 56.405 3.642 ;
      RECT 56.38 3.46 56.39 3.653 ;
      RECT 56.35 3.477 56.38 3.67 ;
      RECT 56.34 3.495 56.35 3.688 ;
      RECT 56.325 3.506 56.34 3.699 ;
      RECT 56.285 3.53 56.325 3.715 ;
      RECT 56.25 3.564 56.285 3.732 ;
      RECT 56.22 3.587 56.25 3.744 ;
      RECT 56.205 3.597 56.22 3.753 ;
      RECT 56.165 3.607 56.205 3.764 ;
      RECT 56.145 3.618 56.165 3.776 ;
      RECT 56.14 3.622 56.145 3.783 ;
      RECT 56.125 3.626 56.14 3.788 ;
      RECT 56.115 3.631 56.125 3.793 ;
      RECT 56.11 3.634 56.115 3.796 ;
      RECT 56.08 3.64 56.11 3.803 ;
      RECT 56.045 3.65 56.08 3.817 ;
      RECT 55.985 3.665 56.045 3.837 ;
      RECT 55.93 3.685 55.985 3.861 ;
      RECT 55.901 3.7 55.93 3.879 ;
      RECT 55.815 3.72 55.901 3.904 ;
      RECT 55.81 3.735 55.815 3.924 ;
      RECT 55.8 3.738 55.81 3.925 ;
      RECT 55.775 3.745 55.8 4.01 ;
      RECT 48.825 8.945 49.175 9.295 ;
      RECT 57.65 8.9 58 9.25 ;
      RECT 48.825 8.975 58 9.175 ;
      RECT 56.19 4.98 56.2 5.17 ;
      RECT 54.45 4.855 54.73 5.135 ;
      RECT 57.495 3.795 57.5 4.28 ;
      RECT 57.39 3.795 57.45 4.055 ;
      RECT 57.715 4.765 57.72 4.84 ;
      RECT 57.705 4.632 57.715 4.875 ;
      RECT 57.695 4.467 57.705 4.896 ;
      RECT 57.69 4.337 57.695 4.912 ;
      RECT 57.68 4.227 57.69 4.928 ;
      RECT 57.675 4.126 57.68 4.945 ;
      RECT 57.67 4.108 57.675 4.955 ;
      RECT 57.665 4.09 57.67 4.965 ;
      RECT 57.655 4.065 57.665 4.98 ;
      RECT 57.65 4.045 57.655 4.995 ;
      RECT 57.63 3.795 57.65 5.02 ;
      RECT 57.615 3.795 57.63 5.053 ;
      RECT 57.585 3.795 57.615 5.075 ;
      RECT 57.565 3.795 57.585 5.089 ;
      RECT 57.545 3.795 57.565 4.605 ;
      RECT 57.56 4.672 57.565 5.094 ;
      RECT 57.555 4.702 57.56 5.096 ;
      RECT 57.55 4.715 57.555 5.099 ;
      RECT 57.545 4.725 57.55 5.103 ;
      RECT 57.54 3.795 57.545 4.523 ;
      RECT 57.54 4.735 57.545 5.105 ;
      RECT 57.535 3.795 57.54 4.5 ;
      RECT 57.525 4.757 57.54 5.105 ;
      RECT 57.52 3.795 57.535 4.445 ;
      RECT 57.515 4.782 57.525 5.105 ;
      RECT 57.515 3.795 57.52 4.39 ;
      RECT 57.505 3.795 57.515 4.338 ;
      RECT 57.51 4.795 57.515 5.106 ;
      RECT 57.505 4.807 57.51 5.107 ;
      RECT 57.5 3.795 57.505 4.298 ;
      RECT 57.5 4.82 57.505 5.108 ;
      RECT 57.485 4.835 57.5 5.109 ;
      RECT 57.49 3.795 57.495 4.26 ;
      RECT 57.485 3.795 57.49 4.225 ;
      RECT 57.48 3.795 57.485 4.2 ;
      RECT 57.475 4.862 57.485 5.111 ;
      RECT 57.47 3.795 57.48 4.158 ;
      RECT 57.47 4.88 57.475 5.112 ;
      RECT 57.465 3.795 57.47 4.118 ;
      RECT 57.465 4.887 57.47 5.113 ;
      RECT 57.46 3.795 57.465 4.09 ;
      RECT 57.455 4.905 57.465 5.114 ;
      RECT 57.45 3.795 57.46 4.07 ;
      RECT 57.445 4.925 57.455 5.116 ;
      RECT 57.435 4.942 57.445 5.117 ;
      RECT 57.4 4.965 57.435 5.12 ;
      RECT 57.345 4.983 57.4 5.126 ;
      RECT 57.259 4.991 57.345 5.135 ;
      RECT 57.173 5.002 57.259 5.146 ;
      RECT 57.087 5.012 57.173 5.157 ;
      RECT 57.001 5.022 57.087 5.169 ;
      RECT 56.915 5.032 57.001 5.18 ;
      RECT 56.895 5.038 56.915 5.186 ;
      RECT 56.815 5.04 56.895 5.19 ;
      RECT 56.81 5.039 56.815 5.195 ;
      RECT 56.802 5.038 56.81 5.195 ;
      RECT 56.716 5.034 56.802 5.193 ;
      RECT 56.63 5.026 56.716 5.19 ;
      RECT 56.544 5.017 56.63 5.186 ;
      RECT 56.458 5.009 56.544 5.183 ;
      RECT 56.372 5.001 56.458 5.179 ;
      RECT 56.286 4.992 56.372 5.176 ;
      RECT 56.2 4.984 56.286 5.172 ;
      RECT 56.145 4.977 56.19 5.17 ;
      RECT 56.06 4.97 56.145 5.168 ;
      RECT 55.986 4.962 56.06 5.164 ;
      RECT 55.9 4.954 55.986 5.161 ;
      RECT 55.897 4.95 55.9 5.159 ;
      RECT 55.811 4.946 55.897 5.158 ;
      RECT 55.725 4.938 55.811 5.155 ;
      RECT 55.64 4.933 55.725 5.152 ;
      RECT 55.554 4.93 55.64 5.149 ;
      RECT 55.468 4.928 55.554 5.146 ;
      RECT 55.382 4.925 55.468 5.143 ;
      RECT 55.296 4.922 55.382 5.14 ;
      RECT 55.21 4.919 55.296 5.137 ;
      RECT 55.134 4.917 55.21 5.134 ;
      RECT 55.048 4.914 55.134 5.131 ;
      RECT 54.962 4.911 55.048 5.129 ;
      RECT 54.876 4.909 54.962 5.126 ;
      RECT 54.79 4.906 54.876 5.123 ;
      RECT 54.73 4.897 54.79 5.121 ;
      RECT 57.24 4.515 57.315 4.775 ;
      RECT 57.22 4.495 57.225 4.775 ;
      RECT 56.54 4.28 56.645 4.575 ;
      RECT 50.985 4.255 51.055 4.515 ;
      RECT 56.88 4.13 56.885 4.501 ;
      RECT 56.87 4.185 56.875 4.501 ;
      RECT 57.175 3.355 57.235 3.615 ;
      RECT 57.23 4.51 57.24 4.775 ;
      RECT 57.225 4.5 57.23 4.775 ;
      RECT 57.145 4.447 57.22 4.775 ;
      RECT 57.17 3.355 57.175 3.635 ;
      RECT 57.16 3.355 57.17 3.655 ;
      RECT 57.145 3.355 57.16 3.685 ;
      RECT 57.13 3.355 57.145 3.728 ;
      RECT 57.125 4.39 57.145 4.775 ;
      RECT 57.115 3.355 57.13 3.765 ;
      RECT 57.11 4.37 57.125 4.775 ;
      RECT 57.11 3.355 57.115 3.788 ;
      RECT 57.1 3.355 57.11 3.813 ;
      RECT 57.07 4.337 57.11 4.775 ;
      RECT 57.075 3.355 57.1 3.863 ;
      RECT 57.07 3.355 57.075 3.918 ;
      RECT 57.065 3.355 57.07 3.96 ;
      RECT 57.055 4.3 57.07 4.775 ;
      RECT 57.06 3.355 57.065 4.003 ;
      RECT 57.055 3.355 57.06 4.068 ;
      RECT 57.05 3.355 57.055 4.09 ;
      RECT 57.05 4.288 57.055 4.64 ;
      RECT 57.045 3.355 57.05 4.158 ;
      RECT 57.045 4.28 57.05 4.623 ;
      RECT 57.04 3.355 57.045 4.203 ;
      RECT 57.035 4.262 57.045 4.6 ;
      RECT 57.035 3.355 57.04 4.24 ;
      RECT 57.025 3.355 57.035 4.58 ;
      RECT 57.02 3.355 57.025 4.563 ;
      RECT 57.015 3.355 57.02 4.548 ;
      RECT 57.01 3.355 57.015 4.533 ;
      RECT 56.99 3.355 57.01 4.523 ;
      RECT 56.985 3.355 56.99 4.513 ;
      RECT 56.975 3.355 56.985 4.509 ;
      RECT 56.97 3.632 56.975 4.508 ;
      RECT 56.965 3.655 56.97 4.507 ;
      RECT 56.96 3.685 56.965 4.506 ;
      RECT 56.955 3.712 56.96 4.505 ;
      RECT 56.95 3.74 56.955 4.505 ;
      RECT 56.945 3.767 56.95 4.505 ;
      RECT 56.94 3.787 56.945 4.505 ;
      RECT 56.935 3.815 56.94 4.505 ;
      RECT 56.925 3.857 56.935 4.505 ;
      RECT 56.915 3.902 56.925 4.504 ;
      RECT 56.91 3.955 56.915 4.503 ;
      RECT 56.905 3.987 56.91 4.502 ;
      RECT 56.9 4.007 56.905 4.501 ;
      RECT 56.895 4.045 56.9 4.501 ;
      RECT 56.89 4.067 56.895 4.501 ;
      RECT 56.885 4.092 56.89 4.501 ;
      RECT 56.875 4.157 56.88 4.501 ;
      RECT 56.86 4.217 56.87 4.501 ;
      RECT 56.845 4.227 56.86 4.501 ;
      RECT 56.825 4.237 56.845 4.501 ;
      RECT 56.795 4.242 56.825 4.498 ;
      RECT 56.735 4.252 56.795 4.495 ;
      RECT 56.715 4.261 56.735 4.5 ;
      RECT 56.69 4.267 56.715 4.513 ;
      RECT 56.67 4.272 56.69 4.528 ;
      RECT 56.645 4.277 56.67 4.575 ;
      RECT 56.516 4.279 56.54 4.575 ;
      RECT 56.43 4.274 56.516 4.575 ;
      RECT 56.39 4.271 56.43 4.575 ;
      RECT 56.34 4.273 56.39 4.555 ;
      RECT 56.31 4.277 56.34 4.555 ;
      RECT 56.231 4.287 56.31 4.555 ;
      RECT 56.145 4.302 56.231 4.556 ;
      RECT 56.095 4.312 56.145 4.557 ;
      RECT 56.087 4.315 56.095 4.557 ;
      RECT 56.001 4.317 56.087 4.558 ;
      RECT 55.915 4.321 56.001 4.558 ;
      RECT 55.829 4.325 55.915 4.559 ;
      RECT 55.743 4.328 55.829 4.56 ;
      RECT 55.657 4.332 55.743 4.56 ;
      RECT 55.571 4.336 55.657 4.561 ;
      RECT 55.485 4.339 55.571 4.562 ;
      RECT 55.399 4.343 55.485 4.562 ;
      RECT 55.313 4.347 55.399 4.563 ;
      RECT 55.227 4.351 55.313 4.564 ;
      RECT 55.141 4.354 55.227 4.564 ;
      RECT 55.055 4.358 55.141 4.565 ;
      RECT 55.025 4.36 55.055 4.565 ;
      RECT 54.939 4.363 55.025 4.566 ;
      RECT 54.853 4.367 54.939 4.567 ;
      RECT 54.767 4.371 54.853 4.568 ;
      RECT 54.681 4.374 54.767 4.568 ;
      RECT 54.595 4.378 54.681 4.569 ;
      RECT 54.56 4.383 54.595 4.57 ;
      RECT 54.505 4.393 54.56 4.577 ;
      RECT 54.48 4.405 54.505 4.587 ;
      RECT 54.445 4.418 54.48 4.595 ;
      RECT 54.405 4.435 54.445 4.618 ;
      RECT 54.385 4.448 54.405 4.645 ;
      RECT 54.355 4.46 54.385 4.673 ;
      RECT 54.35 4.468 54.355 4.693 ;
      RECT 54.345 4.471 54.35 4.703 ;
      RECT 54.295 4.483 54.345 4.737 ;
      RECT 54.285 4.498 54.295 4.77 ;
      RECT 54.275 4.504 54.285 4.783 ;
      RECT 54.265 4.511 54.275 4.795 ;
      RECT 54.24 4.524 54.265 4.813 ;
      RECT 54.225 4.539 54.24 4.835 ;
      RECT 54.215 4.547 54.225 4.851 ;
      RECT 54.2 4.556 54.215 4.866 ;
      RECT 54.19 4.566 54.2 4.88 ;
      RECT 54.171 4.579 54.19 4.897 ;
      RECT 54.085 4.624 54.171 4.962 ;
      RECT 54.07 4.669 54.085 5.02 ;
      RECT 54.065 4.678 54.07 5.033 ;
      RECT 54.055 4.685 54.065 5.038 ;
      RECT 54.05 4.69 54.055 5.042 ;
      RECT 54.03 4.7 54.05 5.049 ;
      RECT 54.005 4.72 54.03 5.063 ;
      RECT 53.97 4.745 54.005 5.083 ;
      RECT 53.955 4.768 53.97 5.098 ;
      RECT 53.945 4.778 53.955 5.103 ;
      RECT 53.935 4.786 53.945 5.11 ;
      RECT 53.925 4.795 53.935 5.116 ;
      RECT 53.905 4.807 53.925 5.118 ;
      RECT 53.895 4.82 53.905 5.12 ;
      RECT 53.87 4.835 53.895 5.123 ;
      RECT 53.85 4.852 53.87 5.127 ;
      RECT 53.81 4.88 53.85 5.133 ;
      RECT 53.745 4.927 53.81 5.142 ;
      RECT 53.73 4.96 53.745 5.15 ;
      RECT 53.725 4.967 53.73 5.152 ;
      RECT 53.675 4.992 53.725 5.157 ;
      RECT 53.66 5.016 53.675 5.164 ;
      RECT 53.61 5.021 53.66 5.165 ;
      RECT 53.524 5.025 53.61 5.165 ;
      RECT 53.438 5.025 53.524 5.165 ;
      RECT 53.352 5.025 53.438 5.166 ;
      RECT 53.266 5.025 53.352 5.166 ;
      RECT 53.18 5.025 53.266 5.166 ;
      RECT 53.114 5.025 53.18 5.166 ;
      RECT 53.028 5.025 53.114 5.167 ;
      RECT 52.942 5.025 53.028 5.167 ;
      RECT 52.856 5.026 52.942 5.168 ;
      RECT 52.77 5.026 52.856 5.168 ;
      RECT 52.684 5.026 52.77 5.168 ;
      RECT 52.598 5.026 52.684 5.169 ;
      RECT 52.512 5.026 52.598 5.169 ;
      RECT 52.426 5.027 52.512 5.17 ;
      RECT 52.34 5.027 52.426 5.17 ;
      RECT 52.32 5.027 52.34 5.17 ;
      RECT 52.234 5.027 52.32 5.17 ;
      RECT 52.148 5.027 52.234 5.17 ;
      RECT 52.062 5.028 52.148 5.17 ;
      RECT 51.976 5.028 52.062 5.17 ;
      RECT 51.89 5.028 51.976 5.17 ;
      RECT 51.804 5.029 51.89 5.17 ;
      RECT 51.718 5.029 51.804 5.17 ;
      RECT 51.632 5.029 51.718 5.17 ;
      RECT 51.546 5.029 51.632 5.17 ;
      RECT 51.46 5.03 51.546 5.17 ;
      RECT 51.41 5.027 51.46 5.17 ;
      RECT 51.4 5.025 51.41 5.169 ;
      RECT 51.396 5.025 51.4 5.168 ;
      RECT 51.31 5.02 51.396 5.163 ;
      RECT 51.288 5.013 51.31 5.157 ;
      RECT 51.202 5.004 51.288 5.151 ;
      RECT 51.116 4.991 51.202 5.142 ;
      RECT 51.03 4.977 51.116 5.132 ;
      RECT 50.985 4.967 51.03 5.125 ;
      RECT 50.965 4.255 50.985 4.533 ;
      RECT 50.965 4.96 50.985 5.121 ;
      RECT 50.935 4.255 50.965 4.555 ;
      RECT 50.925 4.927 50.965 5.118 ;
      RECT 50.92 4.255 50.935 4.575 ;
      RECT 50.92 4.892 50.925 5.116 ;
      RECT 50.915 4.255 50.92 4.7 ;
      RECT 50.915 4.852 50.92 5.116 ;
      RECT 50.905 4.255 50.915 5.116 ;
      RECT 50.83 4.255 50.905 5.11 ;
      RECT 50.8 4.255 50.83 5.1 ;
      RECT 50.795 4.255 50.8 5.092 ;
      RECT 50.79 4.297 50.795 5.085 ;
      RECT 50.78 4.366 50.79 5.076 ;
      RECT 50.775 4.436 50.78 5.028 ;
      RECT 50.77 4.5 50.775 4.925 ;
      RECT 50.765 4.535 50.77 4.88 ;
      RECT 50.763 4.572 50.765 4.772 ;
      RECT 50.76 4.58 50.763 4.765 ;
      RECT 50.755 4.645 50.76 4.708 ;
      RECT 54.83 3.735 55.11 4.015 ;
      RECT 54.82 3.735 55.11 3.878 ;
      RECT 54.775 3.6 55.035 3.86 ;
      RECT 54.775 3.715 55.09 3.86 ;
      RECT 54.775 3.685 55.085 3.86 ;
      RECT 54.775 3.672 55.075 3.86 ;
      RECT 54.775 3.662 55.07 3.86 ;
      RECT 50.75 3.645 51.01 3.905 ;
      RECT 54.52 3.195 54.78 3.455 ;
      RECT 54.51 3.22 54.78 3.415 ;
      RECT 54.505 3.22 54.51 3.414 ;
      RECT 54.435 3.215 54.505 3.406 ;
      RECT 54.35 3.202 54.435 3.389 ;
      RECT 54.346 3.194 54.35 3.379 ;
      RECT 54.26 3.187 54.346 3.369 ;
      RECT 54.251 3.179 54.26 3.359 ;
      RECT 54.165 3.172 54.251 3.347 ;
      RECT 54.145 3.163 54.165 3.333 ;
      RECT 54.09 3.158 54.145 3.325 ;
      RECT 54.08 3.152 54.09 3.319 ;
      RECT 54.06 3.15 54.08 3.315 ;
      RECT 54.052 3.149 54.06 3.311 ;
      RECT 53.966 3.141 54.052 3.3 ;
      RECT 53.88 3.127 53.966 3.28 ;
      RECT 53.82 3.115 53.88 3.265 ;
      RECT 53.81 3.11 53.82 3.26 ;
      RECT 53.76 3.11 53.81 3.262 ;
      RECT 53.713 3.112 53.76 3.266 ;
      RECT 53.627 3.119 53.713 3.271 ;
      RECT 53.541 3.127 53.627 3.277 ;
      RECT 53.455 3.136 53.541 3.283 ;
      RECT 53.396 3.142 53.455 3.288 ;
      RECT 53.31 3.147 53.396 3.294 ;
      RECT 53.235 3.152 53.31 3.3 ;
      RECT 53.196 3.154 53.235 3.305 ;
      RECT 53.11 3.151 53.196 3.31 ;
      RECT 53.025 3.149 53.11 3.317 ;
      RECT 52.993 3.148 53.025 3.32 ;
      RECT 52.907 3.147 52.993 3.321 ;
      RECT 52.821 3.146 52.907 3.322 ;
      RECT 52.735 3.145 52.821 3.322 ;
      RECT 52.649 3.144 52.735 3.323 ;
      RECT 52.563 3.143 52.649 3.324 ;
      RECT 52.477 3.142 52.563 3.325 ;
      RECT 52.391 3.141 52.477 3.325 ;
      RECT 52.305 3.14 52.391 3.326 ;
      RECT 52.255 3.14 52.305 3.327 ;
      RECT 52.241 3.141 52.255 3.327 ;
      RECT 52.155 3.148 52.241 3.328 ;
      RECT 52.081 3.159 52.155 3.329 ;
      RECT 51.995 3.168 52.081 3.33 ;
      RECT 51.96 3.175 51.995 3.345 ;
      RECT 51.935 3.178 51.96 3.375 ;
      RECT 51.91 3.187 51.935 3.404 ;
      RECT 51.9 3.198 51.91 3.424 ;
      RECT 51.89 3.206 51.9 3.438 ;
      RECT 51.885 3.212 51.89 3.448 ;
      RECT 51.86 3.229 51.885 3.465 ;
      RECT 51.845 3.251 51.86 3.493 ;
      RECT 51.815 3.277 51.845 3.523 ;
      RECT 51.795 3.306 51.815 3.553 ;
      RECT 51.79 3.321 51.795 3.57 ;
      RECT 51.77 3.336 51.79 3.585 ;
      RECT 51.76 3.354 51.77 3.603 ;
      RECT 51.75 3.365 51.76 3.618 ;
      RECT 51.7 3.397 51.75 3.644 ;
      RECT 51.695 3.427 51.7 3.664 ;
      RECT 51.685 3.44 51.695 3.67 ;
      RECT 51.676 3.45 51.685 3.678 ;
      RECT 51.665 3.461 51.676 3.686 ;
      RECT 51.66 3.471 51.665 3.692 ;
      RECT 51.645 3.492 51.66 3.699 ;
      RECT 51.63 3.522 51.645 3.707 ;
      RECT 51.595 3.552 51.63 3.713 ;
      RECT 51.57 3.57 51.595 3.72 ;
      RECT 51.52 3.578 51.57 3.729 ;
      RECT 51.495 3.583 51.52 3.738 ;
      RECT 51.44 3.589 51.495 3.748 ;
      RECT 51.435 3.594 51.44 3.756 ;
      RECT 51.421 3.597 51.435 3.758 ;
      RECT 51.335 3.609 51.421 3.77 ;
      RECT 51.325 3.621 51.335 3.783 ;
      RECT 51.24 3.634 51.325 3.795 ;
      RECT 51.196 3.651 51.24 3.809 ;
      RECT 51.11 3.668 51.196 3.825 ;
      RECT 51.08 3.682 51.11 3.839 ;
      RECT 51.07 3.687 51.08 3.844 ;
      RECT 51.01 3.69 51.07 3.853 ;
      RECT 53.9 3.96 54.16 4.22 ;
      RECT 53.9 3.96 54.18 4.073 ;
      RECT 53.9 3.96 54.205 4.04 ;
      RECT 53.9 3.96 54.21 4.02 ;
      RECT 53.95 3.735 54.23 4.015 ;
      RECT 53.505 4.47 53.765 4.73 ;
      RECT 53.495 4.327 53.69 4.668 ;
      RECT 53.49 4.435 53.705 4.66 ;
      RECT 53.485 4.485 53.765 4.65 ;
      RECT 53.475 4.562 53.765 4.635 ;
      RECT 53.495 4.41 53.705 4.668 ;
      RECT 53.505 4.285 53.69 4.73 ;
      RECT 53.505 4.18 53.67 4.73 ;
      RECT 53.515 4.167 53.67 4.73 ;
      RECT 53.515 4.125 53.66 4.73 ;
      RECT 53.52 4.05 53.66 4.73 ;
      RECT 53.55 3.7 53.66 4.73 ;
      RECT 53.555 3.43 53.68 4.053 ;
      RECT 53.525 4.005 53.68 4.053 ;
      RECT 53.54 3.807 53.66 4.73 ;
      RECT 53.53 3.917 53.68 4.053 ;
      RECT 53.555 3.43 53.695 3.91 ;
      RECT 53.555 3.43 53.715 3.785 ;
      RECT 53.52 3.43 53.78 3.69 ;
      RECT 52.99 3.735 53.27 4.015 ;
      RECT 52.975 3.735 53.27 3.995 ;
      RECT 51.03 4.6 51.29 4.86 ;
      RECT 52.815 4.455 53.075 4.715 ;
      RECT 52.795 4.475 53.075 4.69 ;
      RECT 52.752 4.475 52.795 4.689 ;
      RECT 52.666 4.476 52.752 4.686 ;
      RECT 52.58 4.477 52.666 4.682 ;
      RECT 52.505 4.479 52.58 4.679 ;
      RECT 52.482 4.48 52.505 4.677 ;
      RECT 52.396 4.481 52.482 4.675 ;
      RECT 52.31 4.482 52.396 4.672 ;
      RECT 52.286 4.483 52.31 4.67 ;
      RECT 52.2 4.485 52.286 4.667 ;
      RECT 52.115 4.487 52.2 4.668 ;
      RECT 52.058 4.488 52.115 4.674 ;
      RECT 51.972 4.49 52.058 4.684 ;
      RECT 51.886 4.493 51.972 4.697 ;
      RECT 51.8 4.495 51.886 4.709 ;
      RECT 51.786 4.496 51.8 4.716 ;
      RECT 51.7 4.497 51.786 4.724 ;
      RECT 51.66 4.499 51.7 4.733 ;
      RECT 51.651 4.5 51.66 4.736 ;
      RECT 51.565 4.508 51.651 4.742 ;
      RECT 51.545 4.517 51.565 4.75 ;
      RECT 51.46 4.532 51.545 4.758 ;
      RECT 51.4 4.555 51.46 4.769 ;
      RECT 51.39 4.567 51.4 4.774 ;
      RECT 51.35 4.577 51.39 4.778 ;
      RECT 51.295 4.594 51.35 4.786 ;
      RECT 51.29 4.604 51.295 4.79 ;
      RECT 52.356 3.735 52.415 4.132 ;
      RECT 52.27 3.735 52.475 4.123 ;
      RECT 52.265 3.765 52.475 4.118 ;
      RECT 52.231 3.765 52.475 4.116 ;
      RECT 52.145 3.765 52.475 4.11 ;
      RECT 52.1 3.765 52.495 4.088 ;
      RECT 52.1 3.765 52.515 4.043 ;
      RECT 52.06 3.765 52.515 4.033 ;
      RECT 52.27 3.735 52.55 4.015 ;
      RECT 52.005 3.735 52.265 3.995 ;
      RECT 49.83 4.295 50.11 4.575 ;
      RECT 49.8 4.257 50.055 4.56 ;
      RECT 49.795 4.258 50.055 4.558 ;
      RECT 49.79 4.259 50.055 4.552 ;
      RECT 49.785 4.262 50.055 4.545 ;
      RECT 49.78 4.295 50.11 4.538 ;
      RECT 49.75 4.265 50.055 4.525 ;
      RECT 49.75 4.292 50.075 4.525 ;
      RECT 49.75 4.282 50.07 4.525 ;
      RECT 49.75 4.267 50.065 4.525 ;
      RECT 49.83 4.254 50.045 4.575 ;
      RECT 49.916 4.252 50.045 4.575 ;
      RECT 50.002 4.25 50.03 4.575 ;
      RECT 48.795 7.215 49.075 7.585 ;
      RECT 48.75 7.215 49.105 7.57 ;
      RECT 45.645 8.505 45.965 8.83 ;
      RECT 45.675 7.98 45.845 8.83 ;
      RECT 45.675 7.98 45.85 8.33 ;
      RECT 45.675 7.98 46.65 8.155 ;
      RECT 46.475 3.26 46.65 8.155 ;
      RECT 46.42 3.26 46.77 3.61 ;
      RECT 46.445 8.94 46.77 9.265 ;
      RECT 45.33 9.03 46.77 9.2 ;
      RECT 45.33 3.69 45.49 9.2 ;
      RECT 45.645 3.66 45.965 3.98 ;
      RECT 45.33 3.69 45.965 3.86 ;
      RECT 35.415 3.215 35.675 3.475 ;
      RECT 35.47 3.175 35.775 3.455 ;
      RECT 35.47 2.715 35.645 3.475 ;
      RECT 43.985 2.635 44.335 2.985 ;
      RECT 35.47 2.715 44.335 2.89 ;
      RECT 43.66 4.145 44.03 4.515 ;
      RECT 43.745 3.53 43.915 4.515 ;
      RECT 39.765 3.75 40 4.01 ;
      RECT 42.91 3.53 43.075 3.79 ;
      RECT 42.815 3.52 42.83 3.79 ;
      RECT 42.91 3.53 43.915 3.71 ;
      RECT 41.415 3.09 41.455 3.23 ;
      RECT 42.83 3.525 42.91 3.79 ;
      RECT 42.775 3.52 42.815 3.756 ;
      RECT 42.761 3.52 42.775 3.756 ;
      RECT 42.675 3.525 42.761 3.758 ;
      RECT 42.63 3.532 42.675 3.76 ;
      RECT 42.6 3.532 42.63 3.762 ;
      RECT 42.575 3.527 42.6 3.764 ;
      RECT 42.545 3.523 42.575 3.773 ;
      RECT 42.535 3.52 42.545 3.785 ;
      RECT 42.53 3.52 42.535 3.793 ;
      RECT 42.525 3.52 42.53 3.798 ;
      RECT 42.515 3.519 42.525 3.808 ;
      RECT 42.51 3.518 42.515 3.818 ;
      RECT 42.495 3.517 42.51 3.823 ;
      RECT 42.467 3.514 42.495 3.85 ;
      RECT 42.381 3.506 42.467 3.85 ;
      RECT 42.295 3.495 42.381 3.85 ;
      RECT 42.255 3.48 42.295 3.85 ;
      RECT 42.215 3.454 42.255 3.85 ;
      RECT 42.21 3.436 42.215 3.662 ;
      RECT 42.2 3.432 42.21 3.652 ;
      RECT 42.185 3.422 42.2 3.639 ;
      RECT 42.165 3.406 42.185 3.624 ;
      RECT 42.15 3.391 42.165 3.609 ;
      RECT 42.14 3.38 42.15 3.599 ;
      RECT 42.115 3.364 42.14 3.588 ;
      RECT 42.11 3.351 42.115 3.578 ;
      RECT 42.105 3.347 42.11 3.573 ;
      RECT 42.05 3.333 42.105 3.551 ;
      RECT 42.011 3.314 42.05 3.515 ;
      RECT 41.925 3.288 42.011 3.468 ;
      RECT 41.921 3.27 41.925 3.434 ;
      RECT 41.835 3.251 41.921 3.412 ;
      RECT 41.83 3.233 41.835 3.39 ;
      RECT 41.825 3.231 41.83 3.388 ;
      RECT 41.815 3.23 41.825 3.383 ;
      RECT 41.755 3.217 41.815 3.369 ;
      RECT 41.71 3.195 41.755 3.348 ;
      RECT 41.65 3.172 41.71 3.327 ;
      RECT 41.586 3.147 41.65 3.302 ;
      RECT 41.5 3.117 41.586 3.271 ;
      RECT 41.485 3.097 41.5 3.25 ;
      RECT 41.455 3.092 41.485 3.241 ;
      RECT 41.402 3.09 41.415 3.23 ;
      RECT 41.316 3.09 41.402 3.232 ;
      RECT 41.23 3.09 41.316 3.234 ;
      RECT 41.21 3.09 41.23 3.238 ;
      RECT 41.165 3.092 41.21 3.249 ;
      RECT 41.125 3.102 41.165 3.265 ;
      RECT 41.121 3.111 41.125 3.273 ;
      RECT 41.035 3.131 41.121 3.289 ;
      RECT 41.025 3.15 41.035 3.307 ;
      RECT 41.02 3.152 41.025 3.31 ;
      RECT 41.01 3.156 41.02 3.313 ;
      RECT 40.99 3.161 41.01 3.323 ;
      RECT 40.96 3.171 40.99 3.343 ;
      RECT 40.955 3.178 40.96 3.357 ;
      RECT 40.945 3.182 40.955 3.364 ;
      RECT 40.93 3.19 40.945 3.375 ;
      RECT 40.92 3.2 40.93 3.386 ;
      RECT 40.91 3.207 40.92 3.394 ;
      RECT 40.885 3.22 40.91 3.409 ;
      RECT 40.821 3.256 40.885 3.448 ;
      RECT 40.735 3.319 40.821 3.512 ;
      RECT 40.7 3.37 40.735 3.565 ;
      RECT 40.695 3.387 40.7 3.582 ;
      RECT 40.68 3.396 40.695 3.589 ;
      RECT 40.66 3.411 40.68 3.603 ;
      RECT 40.655 3.422 40.66 3.613 ;
      RECT 40.635 3.435 40.655 3.623 ;
      RECT 40.63 3.445 40.635 3.633 ;
      RECT 40.615 3.45 40.63 3.642 ;
      RECT 40.605 3.46 40.615 3.653 ;
      RECT 40.575 3.477 40.605 3.67 ;
      RECT 40.565 3.495 40.575 3.688 ;
      RECT 40.55 3.506 40.565 3.699 ;
      RECT 40.51 3.53 40.55 3.715 ;
      RECT 40.475 3.564 40.51 3.732 ;
      RECT 40.445 3.587 40.475 3.744 ;
      RECT 40.43 3.597 40.445 3.753 ;
      RECT 40.39 3.607 40.43 3.764 ;
      RECT 40.37 3.618 40.39 3.776 ;
      RECT 40.365 3.622 40.37 3.783 ;
      RECT 40.35 3.626 40.365 3.788 ;
      RECT 40.34 3.631 40.35 3.793 ;
      RECT 40.335 3.634 40.34 3.796 ;
      RECT 40.305 3.64 40.335 3.803 ;
      RECT 40.27 3.65 40.305 3.817 ;
      RECT 40.21 3.665 40.27 3.837 ;
      RECT 40.155 3.685 40.21 3.861 ;
      RECT 40.126 3.7 40.155 3.879 ;
      RECT 40.04 3.72 40.126 3.904 ;
      RECT 40.035 3.735 40.04 3.924 ;
      RECT 40.025 3.738 40.035 3.925 ;
      RECT 40 3.745 40.025 4.01 ;
      RECT 33.045 8.94 33.395 9.29 ;
      RECT 41.87 8.895 42.22 9.245 ;
      RECT 33.045 8.97 42.22 9.17 ;
      RECT 40.415 4.98 40.425 5.17 ;
      RECT 38.675 4.855 38.955 5.135 ;
      RECT 41.72 3.795 41.725 4.28 ;
      RECT 41.615 3.795 41.675 4.055 ;
      RECT 41.94 4.765 41.945 4.84 ;
      RECT 41.93 4.632 41.94 4.875 ;
      RECT 41.92 4.467 41.93 4.896 ;
      RECT 41.915 4.337 41.92 4.912 ;
      RECT 41.905 4.227 41.915 4.928 ;
      RECT 41.9 4.126 41.905 4.945 ;
      RECT 41.895 4.108 41.9 4.955 ;
      RECT 41.89 4.09 41.895 4.965 ;
      RECT 41.88 4.065 41.89 4.98 ;
      RECT 41.875 4.045 41.88 4.995 ;
      RECT 41.855 3.795 41.875 5.02 ;
      RECT 41.84 3.795 41.855 5.053 ;
      RECT 41.81 3.795 41.84 5.075 ;
      RECT 41.79 3.795 41.81 5.089 ;
      RECT 41.77 3.795 41.79 4.605 ;
      RECT 41.785 4.672 41.79 5.094 ;
      RECT 41.78 4.702 41.785 5.096 ;
      RECT 41.775 4.715 41.78 5.099 ;
      RECT 41.77 4.725 41.775 5.103 ;
      RECT 41.765 3.795 41.77 4.523 ;
      RECT 41.765 4.735 41.77 5.105 ;
      RECT 41.76 3.795 41.765 4.5 ;
      RECT 41.75 4.757 41.765 5.105 ;
      RECT 41.745 3.795 41.76 4.445 ;
      RECT 41.74 4.782 41.75 5.105 ;
      RECT 41.74 3.795 41.745 4.39 ;
      RECT 41.73 3.795 41.74 4.338 ;
      RECT 41.735 4.795 41.74 5.106 ;
      RECT 41.73 4.807 41.735 5.107 ;
      RECT 41.725 3.795 41.73 4.298 ;
      RECT 41.725 4.82 41.73 5.108 ;
      RECT 41.71 4.835 41.725 5.109 ;
      RECT 41.715 3.795 41.72 4.26 ;
      RECT 41.71 3.795 41.715 4.225 ;
      RECT 41.705 3.795 41.71 4.2 ;
      RECT 41.7 4.862 41.71 5.111 ;
      RECT 41.695 3.795 41.705 4.158 ;
      RECT 41.695 4.88 41.7 5.112 ;
      RECT 41.69 3.795 41.695 4.118 ;
      RECT 41.69 4.887 41.695 5.113 ;
      RECT 41.685 3.795 41.69 4.09 ;
      RECT 41.68 4.905 41.69 5.114 ;
      RECT 41.675 3.795 41.685 4.07 ;
      RECT 41.67 4.925 41.68 5.116 ;
      RECT 41.66 4.942 41.67 5.117 ;
      RECT 41.625 4.965 41.66 5.12 ;
      RECT 41.57 4.983 41.625 5.126 ;
      RECT 41.484 4.991 41.57 5.135 ;
      RECT 41.398 5.002 41.484 5.146 ;
      RECT 41.312 5.012 41.398 5.157 ;
      RECT 41.226 5.022 41.312 5.169 ;
      RECT 41.14 5.032 41.226 5.18 ;
      RECT 41.12 5.038 41.14 5.186 ;
      RECT 41.04 5.04 41.12 5.19 ;
      RECT 41.035 5.039 41.04 5.195 ;
      RECT 41.027 5.038 41.035 5.195 ;
      RECT 40.941 5.034 41.027 5.193 ;
      RECT 40.855 5.026 40.941 5.19 ;
      RECT 40.769 5.017 40.855 5.186 ;
      RECT 40.683 5.009 40.769 5.183 ;
      RECT 40.597 5.001 40.683 5.179 ;
      RECT 40.511 4.992 40.597 5.176 ;
      RECT 40.425 4.984 40.511 5.172 ;
      RECT 40.37 4.977 40.415 5.17 ;
      RECT 40.285 4.97 40.37 5.168 ;
      RECT 40.211 4.962 40.285 5.164 ;
      RECT 40.125 4.954 40.211 5.161 ;
      RECT 40.122 4.95 40.125 5.159 ;
      RECT 40.036 4.946 40.122 5.158 ;
      RECT 39.95 4.938 40.036 5.155 ;
      RECT 39.865 4.933 39.95 5.152 ;
      RECT 39.779 4.93 39.865 5.149 ;
      RECT 39.693 4.928 39.779 5.146 ;
      RECT 39.607 4.925 39.693 5.143 ;
      RECT 39.521 4.922 39.607 5.14 ;
      RECT 39.435 4.919 39.521 5.137 ;
      RECT 39.359 4.917 39.435 5.134 ;
      RECT 39.273 4.914 39.359 5.131 ;
      RECT 39.187 4.911 39.273 5.129 ;
      RECT 39.101 4.909 39.187 5.126 ;
      RECT 39.015 4.906 39.101 5.123 ;
      RECT 38.955 4.897 39.015 5.121 ;
      RECT 41.465 4.515 41.54 4.775 ;
      RECT 41.445 4.495 41.45 4.775 ;
      RECT 40.765 4.28 40.87 4.575 ;
      RECT 35.21 4.255 35.28 4.515 ;
      RECT 41.105 4.13 41.11 4.501 ;
      RECT 41.095 4.185 41.1 4.501 ;
      RECT 41.4 3.355 41.46 3.615 ;
      RECT 41.455 4.51 41.465 4.775 ;
      RECT 41.45 4.5 41.455 4.775 ;
      RECT 41.37 4.447 41.445 4.775 ;
      RECT 41.395 3.355 41.4 3.635 ;
      RECT 41.385 3.355 41.395 3.655 ;
      RECT 41.37 3.355 41.385 3.685 ;
      RECT 41.355 3.355 41.37 3.728 ;
      RECT 41.35 4.39 41.37 4.775 ;
      RECT 41.34 3.355 41.355 3.765 ;
      RECT 41.335 4.37 41.35 4.775 ;
      RECT 41.335 3.355 41.34 3.788 ;
      RECT 41.325 3.355 41.335 3.813 ;
      RECT 41.295 4.337 41.335 4.775 ;
      RECT 41.3 3.355 41.325 3.863 ;
      RECT 41.295 3.355 41.3 3.918 ;
      RECT 41.29 3.355 41.295 3.96 ;
      RECT 41.28 4.3 41.295 4.775 ;
      RECT 41.285 3.355 41.29 4.003 ;
      RECT 41.28 3.355 41.285 4.068 ;
      RECT 41.275 3.355 41.28 4.09 ;
      RECT 41.275 4.288 41.28 4.64 ;
      RECT 41.27 3.355 41.275 4.158 ;
      RECT 41.27 4.28 41.275 4.623 ;
      RECT 41.265 3.355 41.27 4.203 ;
      RECT 41.26 4.262 41.27 4.6 ;
      RECT 41.26 3.355 41.265 4.24 ;
      RECT 41.25 3.355 41.26 4.58 ;
      RECT 41.245 3.355 41.25 4.563 ;
      RECT 41.24 3.355 41.245 4.548 ;
      RECT 41.235 3.355 41.24 4.533 ;
      RECT 41.215 3.355 41.235 4.523 ;
      RECT 41.21 3.355 41.215 4.513 ;
      RECT 41.2 3.355 41.21 4.509 ;
      RECT 41.195 3.632 41.2 4.508 ;
      RECT 41.19 3.655 41.195 4.507 ;
      RECT 41.185 3.685 41.19 4.506 ;
      RECT 41.18 3.712 41.185 4.505 ;
      RECT 41.175 3.74 41.18 4.505 ;
      RECT 41.17 3.767 41.175 4.505 ;
      RECT 41.165 3.787 41.17 4.505 ;
      RECT 41.16 3.815 41.165 4.505 ;
      RECT 41.15 3.857 41.16 4.505 ;
      RECT 41.14 3.902 41.15 4.504 ;
      RECT 41.135 3.955 41.14 4.503 ;
      RECT 41.13 3.987 41.135 4.502 ;
      RECT 41.125 4.007 41.13 4.501 ;
      RECT 41.12 4.045 41.125 4.501 ;
      RECT 41.115 4.067 41.12 4.501 ;
      RECT 41.11 4.092 41.115 4.501 ;
      RECT 41.1 4.157 41.105 4.501 ;
      RECT 41.085 4.217 41.095 4.501 ;
      RECT 41.07 4.227 41.085 4.501 ;
      RECT 41.05 4.237 41.07 4.501 ;
      RECT 41.02 4.242 41.05 4.498 ;
      RECT 40.96 4.252 41.02 4.495 ;
      RECT 40.94 4.261 40.96 4.5 ;
      RECT 40.915 4.267 40.94 4.513 ;
      RECT 40.895 4.272 40.915 4.528 ;
      RECT 40.87 4.277 40.895 4.575 ;
      RECT 40.741 4.279 40.765 4.575 ;
      RECT 40.655 4.274 40.741 4.575 ;
      RECT 40.615 4.271 40.655 4.575 ;
      RECT 40.565 4.273 40.615 4.555 ;
      RECT 40.535 4.277 40.565 4.555 ;
      RECT 40.456 4.287 40.535 4.555 ;
      RECT 40.37 4.302 40.456 4.556 ;
      RECT 40.32 4.312 40.37 4.557 ;
      RECT 40.312 4.315 40.32 4.557 ;
      RECT 40.226 4.317 40.312 4.558 ;
      RECT 40.14 4.321 40.226 4.558 ;
      RECT 40.054 4.325 40.14 4.559 ;
      RECT 39.968 4.328 40.054 4.56 ;
      RECT 39.882 4.332 39.968 4.56 ;
      RECT 39.796 4.336 39.882 4.561 ;
      RECT 39.71 4.339 39.796 4.562 ;
      RECT 39.624 4.343 39.71 4.562 ;
      RECT 39.538 4.347 39.624 4.563 ;
      RECT 39.452 4.351 39.538 4.564 ;
      RECT 39.366 4.354 39.452 4.564 ;
      RECT 39.28 4.358 39.366 4.565 ;
      RECT 39.25 4.36 39.28 4.565 ;
      RECT 39.164 4.363 39.25 4.566 ;
      RECT 39.078 4.367 39.164 4.567 ;
      RECT 38.992 4.371 39.078 4.568 ;
      RECT 38.906 4.374 38.992 4.568 ;
      RECT 38.82 4.378 38.906 4.569 ;
      RECT 38.785 4.383 38.82 4.57 ;
      RECT 38.73 4.393 38.785 4.577 ;
      RECT 38.705 4.405 38.73 4.587 ;
      RECT 38.67 4.418 38.705 4.595 ;
      RECT 38.63 4.435 38.67 4.618 ;
      RECT 38.61 4.448 38.63 4.645 ;
      RECT 38.58 4.46 38.61 4.673 ;
      RECT 38.575 4.468 38.58 4.693 ;
      RECT 38.57 4.471 38.575 4.703 ;
      RECT 38.52 4.483 38.57 4.737 ;
      RECT 38.51 4.498 38.52 4.77 ;
      RECT 38.5 4.504 38.51 4.783 ;
      RECT 38.49 4.511 38.5 4.795 ;
      RECT 38.465 4.524 38.49 4.813 ;
      RECT 38.45 4.539 38.465 4.835 ;
      RECT 38.44 4.547 38.45 4.851 ;
      RECT 38.425 4.556 38.44 4.866 ;
      RECT 38.415 4.566 38.425 4.88 ;
      RECT 38.396 4.579 38.415 4.897 ;
      RECT 38.31 4.624 38.396 4.962 ;
      RECT 38.295 4.669 38.31 5.02 ;
      RECT 38.29 4.678 38.295 5.033 ;
      RECT 38.28 4.685 38.29 5.038 ;
      RECT 38.275 4.69 38.28 5.042 ;
      RECT 38.255 4.7 38.275 5.049 ;
      RECT 38.23 4.72 38.255 5.063 ;
      RECT 38.195 4.745 38.23 5.083 ;
      RECT 38.18 4.768 38.195 5.098 ;
      RECT 38.17 4.778 38.18 5.103 ;
      RECT 38.16 4.786 38.17 5.11 ;
      RECT 38.15 4.795 38.16 5.116 ;
      RECT 38.13 4.807 38.15 5.118 ;
      RECT 38.12 4.82 38.13 5.12 ;
      RECT 38.095 4.835 38.12 5.123 ;
      RECT 38.075 4.852 38.095 5.127 ;
      RECT 38.035 4.88 38.075 5.133 ;
      RECT 37.97 4.927 38.035 5.142 ;
      RECT 37.955 4.96 37.97 5.15 ;
      RECT 37.95 4.967 37.955 5.152 ;
      RECT 37.9 4.992 37.95 5.157 ;
      RECT 37.885 5.016 37.9 5.164 ;
      RECT 37.835 5.021 37.885 5.165 ;
      RECT 37.749 5.025 37.835 5.165 ;
      RECT 37.663 5.025 37.749 5.165 ;
      RECT 37.577 5.025 37.663 5.166 ;
      RECT 37.491 5.025 37.577 5.166 ;
      RECT 37.405 5.025 37.491 5.166 ;
      RECT 37.339 5.025 37.405 5.166 ;
      RECT 37.253 5.025 37.339 5.167 ;
      RECT 37.167 5.025 37.253 5.167 ;
      RECT 37.081 5.026 37.167 5.168 ;
      RECT 36.995 5.026 37.081 5.168 ;
      RECT 36.909 5.026 36.995 5.168 ;
      RECT 36.823 5.026 36.909 5.169 ;
      RECT 36.737 5.026 36.823 5.169 ;
      RECT 36.651 5.027 36.737 5.17 ;
      RECT 36.565 5.027 36.651 5.17 ;
      RECT 36.545 5.027 36.565 5.17 ;
      RECT 36.459 5.027 36.545 5.17 ;
      RECT 36.373 5.027 36.459 5.17 ;
      RECT 36.287 5.028 36.373 5.17 ;
      RECT 36.201 5.028 36.287 5.17 ;
      RECT 36.115 5.028 36.201 5.17 ;
      RECT 36.029 5.029 36.115 5.17 ;
      RECT 35.943 5.029 36.029 5.17 ;
      RECT 35.857 5.029 35.943 5.17 ;
      RECT 35.771 5.029 35.857 5.17 ;
      RECT 35.685 5.03 35.771 5.17 ;
      RECT 35.635 5.027 35.685 5.17 ;
      RECT 35.625 5.025 35.635 5.169 ;
      RECT 35.621 5.025 35.625 5.168 ;
      RECT 35.535 5.02 35.621 5.163 ;
      RECT 35.513 5.013 35.535 5.157 ;
      RECT 35.427 5.004 35.513 5.151 ;
      RECT 35.341 4.991 35.427 5.142 ;
      RECT 35.255 4.977 35.341 5.132 ;
      RECT 35.21 4.967 35.255 5.125 ;
      RECT 35.19 4.255 35.21 4.533 ;
      RECT 35.19 4.96 35.21 5.121 ;
      RECT 35.16 4.255 35.19 4.555 ;
      RECT 35.15 4.927 35.19 5.118 ;
      RECT 35.145 4.255 35.16 4.575 ;
      RECT 35.145 4.892 35.15 5.116 ;
      RECT 35.14 4.255 35.145 4.7 ;
      RECT 35.14 4.852 35.145 5.116 ;
      RECT 35.13 4.255 35.14 5.116 ;
      RECT 35.055 4.255 35.13 5.11 ;
      RECT 35.025 4.255 35.055 5.1 ;
      RECT 35.02 4.255 35.025 5.092 ;
      RECT 35.015 4.297 35.02 5.085 ;
      RECT 35.005 4.366 35.015 5.076 ;
      RECT 35 4.436 35.005 5.028 ;
      RECT 34.995 4.5 35 4.925 ;
      RECT 34.99 4.535 34.995 4.88 ;
      RECT 34.988 4.572 34.99 4.772 ;
      RECT 34.985 4.58 34.988 4.765 ;
      RECT 34.98 4.645 34.985 4.708 ;
      RECT 39.055 3.735 39.335 4.015 ;
      RECT 39.045 3.735 39.335 3.878 ;
      RECT 39 3.6 39.26 3.86 ;
      RECT 39 3.715 39.315 3.86 ;
      RECT 39 3.685 39.31 3.86 ;
      RECT 39 3.672 39.3 3.86 ;
      RECT 39 3.662 39.295 3.86 ;
      RECT 34.975 3.645 35.235 3.905 ;
      RECT 38.745 3.195 39.005 3.455 ;
      RECT 38.735 3.22 39.005 3.415 ;
      RECT 38.73 3.22 38.735 3.414 ;
      RECT 38.66 3.215 38.73 3.406 ;
      RECT 38.575 3.202 38.66 3.389 ;
      RECT 38.571 3.194 38.575 3.379 ;
      RECT 38.485 3.187 38.571 3.369 ;
      RECT 38.476 3.179 38.485 3.359 ;
      RECT 38.39 3.172 38.476 3.347 ;
      RECT 38.37 3.163 38.39 3.333 ;
      RECT 38.315 3.158 38.37 3.325 ;
      RECT 38.305 3.152 38.315 3.319 ;
      RECT 38.285 3.15 38.305 3.315 ;
      RECT 38.277 3.149 38.285 3.311 ;
      RECT 38.191 3.141 38.277 3.3 ;
      RECT 38.105 3.127 38.191 3.28 ;
      RECT 38.045 3.115 38.105 3.265 ;
      RECT 38.035 3.11 38.045 3.26 ;
      RECT 37.985 3.11 38.035 3.262 ;
      RECT 37.938 3.112 37.985 3.266 ;
      RECT 37.852 3.119 37.938 3.271 ;
      RECT 37.766 3.127 37.852 3.277 ;
      RECT 37.68 3.136 37.766 3.283 ;
      RECT 37.621 3.142 37.68 3.288 ;
      RECT 37.535 3.147 37.621 3.294 ;
      RECT 37.46 3.152 37.535 3.3 ;
      RECT 37.421 3.154 37.46 3.305 ;
      RECT 37.335 3.151 37.421 3.31 ;
      RECT 37.25 3.149 37.335 3.317 ;
      RECT 37.218 3.148 37.25 3.32 ;
      RECT 37.132 3.147 37.218 3.321 ;
      RECT 37.046 3.146 37.132 3.322 ;
      RECT 36.96 3.145 37.046 3.322 ;
      RECT 36.874 3.144 36.96 3.323 ;
      RECT 36.788 3.143 36.874 3.324 ;
      RECT 36.702 3.142 36.788 3.325 ;
      RECT 36.616 3.141 36.702 3.325 ;
      RECT 36.53 3.14 36.616 3.326 ;
      RECT 36.48 3.14 36.53 3.327 ;
      RECT 36.466 3.141 36.48 3.327 ;
      RECT 36.38 3.148 36.466 3.328 ;
      RECT 36.306 3.159 36.38 3.329 ;
      RECT 36.22 3.168 36.306 3.33 ;
      RECT 36.185 3.175 36.22 3.345 ;
      RECT 36.16 3.178 36.185 3.375 ;
      RECT 36.135 3.187 36.16 3.404 ;
      RECT 36.125 3.198 36.135 3.424 ;
      RECT 36.115 3.206 36.125 3.438 ;
      RECT 36.11 3.212 36.115 3.448 ;
      RECT 36.085 3.229 36.11 3.465 ;
      RECT 36.07 3.251 36.085 3.493 ;
      RECT 36.04 3.277 36.07 3.523 ;
      RECT 36.02 3.306 36.04 3.553 ;
      RECT 36.015 3.321 36.02 3.57 ;
      RECT 35.995 3.336 36.015 3.585 ;
      RECT 35.985 3.354 35.995 3.603 ;
      RECT 35.975 3.365 35.985 3.618 ;
      RECT 35.925 3.397 35.975 3.644 ;
      RECT 35.92 3.427 35.925 3.664 ;
      RECT 35.91 3.44 35.92 3.67 ;
      RECT 35.901 3.45 35.91 3.678 ;
      RECT 35.89 3.461 35.901 3.686 ;
      RECT 35.885 3.471 35.89 3.692 ;
      RECT 35.87 3.492 35.885 3.699 ;
      RECT 35.855 3.522 35.87 3.707 ;
      RECT 35.82 3.552 35.855 3.713 ;
      RECT 35.795 3.57 35.82 3.72 ;
      RECT 35.745 3.578 35.795 3.729 ;
      RECT 35.72 3.583 35.745 3.738 ;
      RECT 35.665 3.589 35.72 3.748 ;
      RECT 35.66 3.594 35.665 3.756 ;
      RECT 35.646 3.597 35.66 3.758 ;
      RECT 35.56 3.609 35.646 3.77 ;
      RECT 35.55 3.621 35.56 3.783 ;
      RECT 35.465 3.634 35.55 3.795 ;
      RECT 35.421 3.651 35.465 3.809 ;
      RECT 35.335 3.668 35.421 3.825 ;
      RECT 35.305 3.682 35.335 3.839 ;
      RECT 35.295 3.687 35.305 3.844 ;
      RECT 35.235 3.69 35.295 3.853 ;
      RECT 38.125 3.96 38.385 4.22 ;
      RECT 38.125 3.96 38.405 4.073 ;
      RECT 38.125 3.96 38.43 4.04 ;
      RECT 38.125 3.96 38.435 4.02 ;
      RECT 38.175 3.735 38.455 4.015 ;
      RECT 37.73 4.47 37.99 4.73 ;
      RECT 37.72 4.327 37.915 4.668 ;
      RECT 37.715 4.435 37.93 4.66 ;
      RECT 37.71 4.485 37.99 4.65 ;
      RECT 37.7 4.562 37.99 4.635 ;
      RECT 37.72 4.41 37.93 4.668 ;
      RECT 37.73 4.285 37.915 4.73 ;
      RECT 37.73 4.18 37.895 4.73 ;
      RECT 37.74 4.167 37.895 4.73 ;
      RECT 37.74 4.125 37.885 4.73 ;
      RECT 37.745 4.05 37.885 4.73 ;
      RECT 37.775 3.7 37.885 4.73 ;
      RECT 37.78 3.43 37.905 4.053 ;
      RECT 37.75 4.005 37.905 4.053 ;
      RECT 37.765 3.807 37.885 4.73 ;
      RECT 37.755 3.917 37.905 4.053 ;
      RECT 37.78 3.43 37.92 3.91 ;
      RECT 37.78 3.43 37.94 3.785 ;
      RECT 37.745 3.43 38.005 3.69 ;
      RECT 37.215 3.735 37.495 4.015 ;
      RECT 37.2 3.735 37.495 3.995 ;
      RECT 35.255 4.6 35.515 4.86 ;
      RECT 37.04 4.455 37.3 4.715 ;
      RECT 37.02 4.475 37.3 4.69 ;
      RECT 36.977 4.475 37.02 4.689 ;
      RECT 36.891 4.476 36.977 4.686 ;
      RECT 36.805 4.477 36.891 4.682 ;
      RECT 36.73 4.479 36.805 4.679 ;
      RECT 36.707 4.48 36.73 4.677 ;
      RECT 36.621 4.481 36.707 4.675 ;
      RECT 36.535 4.482 36.621 4.672 ;
      RECT 36.511 4.483 36.535 4.67 ;
      RECT 36.425 4.485 36.511 4.667 ;
      RECT 36.34 4.487 36.425 4.668 ;
      RECT 36.283 4.488 36.34 4.674 ;
      RECT 36.197 4.49 36.283 4.684 ;
      RECT 36.111 4.493 36.197 4.697 ;
      RECT 36.025 4.495 36.111 4.709 ;
      RECT 36.011 4.496 36.025 4.716 ;
      RECT 35.925 4.497 36.011 4.724 ;
      RECT 35.885 4.499 35.925 4.733 ;
      RECT 35.876 4.5 35.885 4.736 ;
      RECT 35.79 4.508 35.876 4.742 ;
      RECT 35.77 4.517 35.79 4.75 ;
      RECT 35.685 4.532 35.77 4.758 ;
      RECT 35.625 4.555 35.685 4.769 ;
      RECT 35.615 4.567 35.625 4.774 ;
      RECT 35.575 4.577 35.615 4.778 ;
      RECT 35.52 4.594 35.575 4.786 ;
      RECT 35.515 4.604 35.52 4.79 ;
      RECT 36.581 3.735 36.64 4.132 ;
      RECT 36.495 3.735 36.7 4.123 ;
      RECT 36.49 3.765 36.7 4.118 ;
      RECT 36.456 3.765 36.7 4.116 ;
      RECT 36.37 3.765 36.7 4.11 ;
      RECT 36.325 3.765 36.72 4.088 ;
      RECT 36.325 3.765 36.74 4.043 ;
      RECT 36.285 3.765 36.74 4.033 ;
      RECT 36.495 3.735 36.775 4.015 ;
      RECT 36.23 3.735 36.49 3.995 ;
      RECT 34.055 4.295 34.335 4.575 ;
      RECT 34.025 4.257 34.28 4.56 ;
      RECT 34.02 4.258 34.28 4.558 ;
      RECT 34.015 4.259 34.28 4.552 ;
      RECT 34.01 4.262 34.28 4.545 ;
      RECT 34.005 4.295 34.335 4.538 ;
      RECT 33.975 4.265 34.28 4.525 ;
      RECT 33.975 4.292 34.3 4.525 ;
      RECT 33.975 4.282 34.295 4.525 ;
      RECT 33.975 4.267 34.29 4.525 ;
      RECT 34.055 4.254 34.27 4.575 ;
      RECT 34.141 4.252 34.27 4.575 ;
      RECT 34.227 4.25 34.255 4.575 ;
      RECT 33.015 7.215 33.295 7.585 ;
      RECT 32.97 7.215 33.325 7.57 ;
      RECT 29.865 8.505 30.185 8.83 ;
      RECT 29.895 7.98 30.065 8.83 ;
      RECT 29.895 7.98 30.07 8.33 ;
      RECT 29.895 7.98 30.87 8.155 ;
      RECT 30.695 3.26 30.87 8.155 ;
      RECT 30.64 3.26 30.99 3.61 ;
      RECT 30.665 8.94 30.99 9.265 ;
      RECT 29.55 9.03 30.99 9.2 ;
      RECT 29.55 3.69 29.71 9.2 ;
      RECT 29.865 3.66 30.185 3.98 ;
      RECT 29.55 3.69 30.185 3.86 ;
      RECT 19.635 3.215 19.895 3.475 ;
      RECT 19.69 3.175 19.995 3.455 ;
      RECT 19.69 2.715 19.865 3.475 ;
      RECT 28.205 2.635 28.555 2.985 ;
      RECT 19.69 2.715 28.555 2.89 ;
      RECT 27.88 4.145 28.25 4.515 ;
      RECT 27.965 3.53 28.135 4.515 ;
      RECT 23.985 3.75 24.22 4.01 ;
      RECT 27.13 3.53 27.295 3.79 ;
      RECT 27.035 3.52 27.05 3.79 ;
      RECT 27.13 3.53 28.135 3.71 ;
      RECT 25.635 3.09 25.675 3.23 ;
      RECT 27.05 3.525 27.13 3.79 ;
      RECT 26.995 3.52 27.035 3.756 ;
      RECT 26.981 3.52 26.995 3.756 ;
      RECT 26.895 3.525 26.981 3.758 ;
      RECT 26.85 3.532 26.895 3.76 ;
      RECT 26.82 3.532 26.85 3.762 ;
      RECT 26.795 3.527 26.82 3.764 ;
      RECT 26.765 3.523 26.795 3.773 ;
      RECT 26.755 3.52 26.765 3.785 ;
      RECT 26.75 3.52 26.755 3.793 ;
      RECT 26.745 3.52 26.75 3.798 ;
      RECT 26.735 3.519 26.745 3.808 ;
      RECT 26.73 3.518 26.735 3.818 ;
      RECT 26.715 3.517 26.73 3.823 ;
      RECT 26.687 3.514 26.715 3.85 ;
      RECT 26.601 3.506 26.687 3.85 ;
      RECT 26.515 3.495 26.601 3.85 ;
      RECT 26.475 3.48 26.515 3.85 ;
      RECT 26.435 3.454 26.475 3.85 ;
      RECT 26.43 3.436 26.435 3.662 ;
      RECT 26.42 3.432 26.43 3.652 ;
      RECT 26.405 3.422 26.42 3.639 ;
      RECT 26.385 3.406 26.405 3.624 ;
      RECT 26.37 3.391 26.385 3.609 ;
      RECT 26.36 3.38 26.37 3.599 ;
      RECT 26.335 3.364 26.36 3.588 ;
      RECT 26.33 3.351 26.335 3.578 ;
      RECT 26.325 3.347 26.33 3.573 ;
      RECT 26.27 3.333 26.325 3.551 ;
      RECT 26.231 3.314 26.27 3.515 ;
      RECT 26.145 3.288 26.231 3.468 ;
      RECT 26.141 3.27 26.145 3.434 ;
      RECT 26.055 3.251 26.141 3.412 ;
      RECT 26.05 3.233 26.055 3.39 ;
      RECT 26.045 3.231 26.05 3.388 ;
      RECT 26.035 3.23 26.045 3.383 ;
      RECT 25.975 3.217 26.035 3.369 ;
      RECT 25.93 3.195 25.975 3.348 ;
      RECT 25.87 3.172 25.93 3.327 ;
      RECT 25.806 3.147 25.87 3.302 ;
      RECT 25.72 3.117 25.806 3.271 ;
      RECT 25.705 3.097 25.72 3.25 ;
      RECT 25.675 3.092 25.705 3.241 ;
      RECT 25.622 3.09 25.635 3.23 ;
      RECT 25.536 3.09 25.622 3.232 ;
      RECT 25.45 3.09 25.536 3.234 ;
      RECT 25.43 3.09 25.45 3.238 ;
      RECT 25.385 3.092 25.43 3.249 ;
      RECT 25.345 3.102 25.385 3.265 ;
      RECT 25.341 3.111 25.345 3.273 ;
      RECT 25.255 3.131 25.341 3.289 ;
      RECT 25.245 3.15 25.255 3.307 ;
      RECT 25.24 3.152 25.245 3.31 ;
      RECT 25.23 3.156 25.24 3.313 ;
      RECT 25.21 3.161 25.23 3.323 ;
      RECT 25.18 3.171 25.21 3.343 ;
      RECT 25.175 3.178 25.18 3.357 ;
      RECT 25.165 3.182 25.175 3.364 ;
      RECT 25.15 3.19 25.165 3.375 ;
      RECT 25.14 3.2 25.15 3.386 ;
      RECT 25.13 3.207 25.14 3.394 ;
      RECT 25.105 3.22 25.13 3.409 ;
      RECT 25.041 3.256 25.105 3.448 ;
      RECT 24.955 3.319 25.041 3.512 ;
      RECT 24.92 3.37 24.955 3.565 ;
      RECT 24.915 3.387 24.92 3.582 ;
      RECT 24.9 3.396 24.915 3.589 ;
      RECT 24.88 3.411 24.9 3.603 ;
      RECT 24.875 3.422 24.88 3.613 ;
      RECT 24.855 3.435 24.875 3.623 ;
      RECT 24.85 3.445 24.855 3.633 ;
      RECT 24.835 3.45 24.85 3.642 ;
      RECT 24.825 3.46 24.835 3.653 ;
      RECT 24.795 3.477 24.825 3.67 ;
      RECT 24.785 3.495 24.795 3.688 ;
      RECT 24.77 3.506 24.785 3.699 ;
      RECT 24.73 3.53 24.77 3.715 ;
      RECT 24.695 3.564 24.73 3.732 ;
      RECT 24.665 3.587 24.695 3.744 ;
      RECT 24.65 3.597 24.665 3.753 ;
      RECT 24.61 3.607 24.65 3.764 ;
      RECT 24.59 3.618 24.61 3.776 ;
      RECT 24.585 3.622 24.59 3.783 ;
      RECT 24.57 3.626 24.585 3.788 ;
      RECT 24.56 3.631 24.57 3.793 ;
      RECT 24.555 3.634 24.56 3.796 ;
      RECT 24.525 3.64 24.555 3.803 ;
      RECT 24.49 3.65 24.525 3.817 ;
      RECT 24.43 3.665 24.49 3.837 ;
      RECT 24.375 3.685 24.43 3.861 ;
      RECT 24.346 3.7 24.375 3.879 ;
      RECT 24.26 3.72 24.346 3.904 ;
      RECT 24.255 3.735 24.26 3.924 ;
      RECT 24.245 3.738 24.255 3.925 ;
      RECT 24.22 3.745 24.245 4.01 ;
      RECT 16.54 9.28 16.83 9.63 ;
      RECT 16.54 9.37 17.945 9.54 ;
      RECT 17.775 8.97 17.945 9.54 ;
      RECT 26.06 8.89 26.41 9.24 ;
      RECT 17.775 8.97 26.41 9.14 ;
      RECT 24.635 4.98 24.645 5.17 ;
      RECT 22.895 4.855 23.175 5.135 ;
      RECT 25.94 3.795 25.945 4.28 ;
      RECT 25.835 3.795 25.895 4.055 ;
      RECT 26.16 4.765 26.165 4.84 ;
      RECT 26.15 4.632 26.16 4.875 ;
      RECT 26.14 4.467 26.15 4.896 ;
      RECT 26.135 4.337 26.14 4.912 ;
      RECT 26.125 4.227 26.135 4.928 ;
      RECT 26.12 4.126 26.125 4.945 ;
      RECT 26.115 4.108 26.12 4.955 ;
      RECT 26.11 4.09 26.115 4.965 ;
      RECT 26.1 4.065 26.11 4.98 ;
      RECT 26.095 4.045 26.1 4.995 ;
      RECT 26.075 3.795 26.095 5.02 ;
      RECT 26.06 3.795 26.075 5.053 ;
      RECT 26.03 3.795 26.06 5.075 ;
      RECT 26.01 3.795 26.03 5.089 ;
      RECT 25.99 3.795 26.01 4.605 ;
      RECT 26.005 4.672 26.01 5.094 ;
      RECT 26 4.702 26.005 5.096 ;
      RECT 25.995 4.715 26 5.099 ;
      RECT 25.99 4.725 25.995 5.103 ;
      RECT 25.985 3.795 25.99 4.523 ;
      RECT 25.985 4.735 25.99 5.105 ;
      RECT 25.98 3.795 25.985 4.5 ;
      RECT 25.97 4.757 25.985 5.105 ;
      RECT 25.965 3.795 25.98 4.445 ;
      RECT 25.96 4.782 25.97 5.105 ;
      RECT 25.96 3.795 25.965 4.39 ;
      RECT 25.95 3.795 25.96 4.338 ;
      RECT 25.955 4.795 25.96 5.106 ;
      RECT 25.95 4.807 25.955 5.107 ;
      RECT 25.945 3.795 25.95 4.298 ;
      RECT 25.945 4.82 25.95 5.108 ;
      RECT 25.93 4.835 25.945 5.109 ;
      RECT 25.935 3.795 25.94 4.26 ;
      RECT 25.93 3.795 25.935 4.225 ;
      RECT 25.925 3.795 25.93 4.2 ;
      RECT 25.92 4.862 25.93 5.111 ;
      RECT 25.915 3.795 25.925 4.158 ;
      RECT 25.915 4.88 25.92 5.112 ;
      RECT 25.91 3.795 25.915 4.118 ;
      RECT 25.91 4.887 25.915 5.113 ;
      RECT 25.905 3.795 25.91 4.09 ;
      RECT 25.9 4.905 25.91 5.114 ;
      RECT 25.895 3.795 25.905 4.07 ;
      RECT 25.89 4.925 25.9 5.116 ;
      RECT 25.88 4.942 25.89 5.117 ;
      RECT 25.845 4.965 25.88 5.12 ;
      RECT 25.79 4.983 25.845 5.126 ;
      RECT 25.704 4.991 25.79 5.135 ;
      RECT 25.618 5.002 25.704 5.146 ;
      RECT 25.532 5.012 25.618 5.157 ;
      RECT 25.446 5.022 25.532 5.169 ;
      RECT 25.36 5.032 25.446 5.18 ;
      RECT 25.34 5.038 25.36 5.186 ;
      RECT 25.26 5.04 25.34 5.19 ;
      RECT 25.255 5.039 25.26 5.195 ;
      RECT 25.247 5.038 25.255 5.195 ;
      RECT 25.161 5.034 25.247 5.193 ;
      RECT 25.075 5.026 25.161 5.19 ;
      RECT 24.989 5.017 25.075 5.186 ;
      RECT 24.903 5.009 24.989 5.183 ;
      RECT 24.817 5.001 24.903 5.179 ;
      RECT 24.731 4.992 24.817 5.176 ;
      RECT 24.645 4.984 24.731 5.172 ;
      RECT 24.59 4.977 24.635 5.17 ;
      RECT 24.505 4.97 24.59 5.168 ;
      RECT 24.431 4.962 24.505 5.164 ;
      RECT 24.345 4.954 24.431 5.161 ;
      RECT 24.342 4.95 24.345 5.159 ;
      RECT 24.256 4.946 24.342 5.158 ;
      RECT 24.17 4.938 24.256 5.155 ;
      RECT 24.085 4.933 24.17 5.152 ;
      RECT 23.999 4.93 24.085 5.149 ;
      RECT 23.913 4.928 23.999 5.146 ;
      RECT 23.827 4.925 23.913 5.143 ;
      RECT 23.741 4.922 23.827 5.14 ;
      RECT 23.655 4.919 23.741 5.137 ;
      RECT 23.579 4.917 23.655 5.134 ;
      RECT 23.493 4.914 23.579 5.131 ;
      RECT 23.407 4.911 23.493 5.129 ;
      RECT 23.321 4.909 23.407 5.126 ;
      RECT 23.235 4.906 23.321 5.123 ;
      RECT 23.175 4.897 23.235 5.121 ;
      RECT 25.685 4.515 25.76 4.775 ;
      RECT 25.665 4.495 25.67 4.775 ;
      RECT 24.985 4.28 25.09 4.575 ;
      RECT 19.43 4.255 19.5 4.515 ;
      RECT 25.325 4.13 25.33 4.501 ;
      RECT 25.315 4.185 25.32 4.501 ;
      RECT 25.62 3.355 25.68 3.615 ;
      RECT 25.675 4.51 25.685 4.775 ;
      RECT 25.67 4.5 25.675 4.775 ;
      RECT 25.59 4.447 25.665 4.775 ;
      RECT 25.615 3.355 25.62 3.635 ;
      RECT 25.605 3.355 25.615 3.655 ;
      RECT 25.59 3.355 25.605 3.685 ;
      RECT 25.575 3.355 25.59 3.728 ;
      RECT 25.57 4.39 25.59 4.775 ;
      RECT 25.56 3.355 25.575 3.765 ;
      RECT 25.555 4.37 25.57 4.775 ;
      RECT 25.555 3.355 25.56 3.788 ;
      RECT 25.545 3.355 25.555 3.813 ;
      RECT 25.515 4.337 25.555 4.775 ;
      RECT 25.52 3.355 25.545 3.863 ;
      RECT 25.515 3.355 25.52 3.918 ;
      RECT 25.51 3.355 25.515 3.96 ;
      RECT 25.5 4.3 25.515 4.775 ;
      RECT 25.505 3.355 25.51 4.003 ;
      RECT 25.5 3.355 25.505 4.068 ;
      RECT 25.495 3.355 25.5 4.09 ;
      RECT 25.495 4.288 25.5 4.64 ;
      RECT 25.49 3.355 25.495 4.158 ;
      RECT 25.49 4.28 25.495 4.623 ;
      RECT 25.485 3.355 25.49 4.203 ;
      RECT 25.48 4.262 25.49 4.6 ;
      RECT 25.48 3.355 25.485 4.24 ;
      RECT 25.47 3.355 25.48 4.58 ;
      RECT 25.465 3.355 25.47 4.563 ;
      RECT 25.46 3.355 25.465 4.548 ;
      RECT 25.455 3.355 25.46 4.533 ;
      RECT 25.435 3.355 25.455 4.523 ;
      RECT 25.43 3.355 25.435 4.513 ;
      RECT 25.42 3.355 25.43 4.509 ;
      RECT 25.415 3.632 25.42 4.508 ;
      RECT 25.41 3.655 25.415 4.507 ;
      RECT 25.405 3.685 25.41 4.506 ;
      RECT 25.4 3.712 25.405 4.505 ;
      RECT 25.395 3.74 25.4 4.505 ;
      RECT 25.39 3.767 25.395 4.505 ;
      RECT 25.385 3.787 25.39 4.505 ;
      RECT 25.38 3.815 25.385 4.505 ;
      RECT 25.37 3.857 25.38 4.505 ;
      RECT 25.36 3.902 25.37 4.504 ;
      RECT 25.355 3.955 25.36 4.503 ;
      RECT 25.35 3.987 25.355 4.502 ;
      RECT 25.345 4.007 25.35 4.501 ;
      RECT 25.34 4.045 25.345 4.501 ;
      RECT 25.335 4.067 25.34 4.501 ;
      RECT 25.33 4.092 25.335 4.501 ;
      RECT 25.32 4.157 25.325 4.501 ;
      RECT 25.305 4.217 25.315 4.501 ;
      RECT 25.29 4.227 25.305 4.501 ;
      RECT 25.27 4.237 25.29 4.501 ;
      RECT 25.24 4.242 25.27 4.498 ;
      RECT 25.18 4.252 25.24 4.495 ;
      RECT 25.16 4.261 25.18 4.5 ;
      RECT 25.135 4.267 25.16 4.513 ;
      RECT 25.115 4.272 25.135 4.528 ;
      RECT 25.09 4.277 25.115 4.575 ;
      RECT 24.961 4.279 24.985 4.575 ;
      RECT 24.875 4.274 24.961 4.575 ;
      RECT 24.835 4.271 24.875 4.575 ;
      RECT 24.785 4.273 24.835 4.555 ;
      RECT 24.755 4.277 24.785 4.555 ;
      RECT 24.676 4.287 24.755 4.555 ;
      RECT 24.59 4.302 24.676 4.556 ;
      RECT 24.54 4.312 24.59 4.557 ;
      RECT 24.532 4.315 24.54 4.557 ;
      RECT 24.446 4.317 24.532 4.558 ;
      RECT 24.36 4.321 24.446 4.558 ;
      RECT 24.274 4.325 24.36 4.559 ;
      RECT 24.188 4.328 24.274 4.56 ;
      RECT 24.102 4.332 24.188 4.56 ;
      RECT 24.016 4.336 24.102 4.561 ;
      RECT 23.93 4.339 24.016 4.562 ;
      RECT 23.844 4.343 23.93 4.562 ;
      RECT 23.758 4.347 23.844 4.563 ;
      RECT 23.672 4.351 23.758 4.564 ;
      RECT 23.586 4.354 23.672 4.564 ;
      RECT 23.5 4.358 23.586 4.565 ;
      RECT 23.47 4.36 23.5 4.565 ;
      RECT 23.384 4.363 23.47 4.566 ;
      RECT 23.298 4.367 23.384 4.567 ;
      RECT 23.212 4.371 23.298 4.568 ;
      RECT 23.126 4.374 23.212 4.568 ;
      RECT 23.04 4.378 23.126 4.569 ;
      RECT 23.005 4.383 23.04 4.57 ;
      RECT 22.95 4.393 23.005 4.577 ;
      RECT 22.925 4.405 22.95 4.587 ;
      RECT 22.89 4.418 22.925 4.595 ;
      RECT 22.85 4.435 22.89 4.618 ;
      RECT 22.83 4.448 22.85 4.645 ;
      RECT 22.8 4.46 22.83 4.673 ;
      RECT 22.795 4.468 22.8 4.693 ;
      RECT 22.79 4.471 22.795 4.703 ;
      RECT 22.74 4.483 22.79 4.737 ;
      RECT 22.73 4.498 22.74 4.77 ;
      RECT 22.72 4.504 22.73 4.783 ;
      RECT 22.71 4.511 22.72 4.795 ;
      RECT 22.685 4.524 22.71 4.813 ;
      RECT 22.67 4.539 22.685 4.835 ;
      RECT 22.66 4.547 22.67 4.851 ;
      RECT 22.645 4.556 22.66 4.866 ;
      RECT 22.635 4.566 22.645 4.88 ;
      RECT 22.616 4.579 22.635 4.897 ;
      RECT 22.53 4.624 22.616 4.962 ;
      RECT 22.515 4.669 22.53 5.02 ;
      RECT 22.51 4.678 22.515 5.033 ;
      RECT 22.5 4.685 22.51 5.038 ;
      RECT 22.495 4.69 22.5 5.042 ;
      RECT 22.475 4.7 22.495 5.049 ;
      RECT 22.45 4.72 22.475 5.063 ;
      RECT 22.415 4.745 22.45 5.083 ;
      RECT 22.4 4.768 22.415 5.098 ;
      RECT 22.39 4.778 22.4 5.103 ;
      RECT 22.38 4.786 22.39 5.11 ;
      RECT 22.37 4.795 22.38 5.116 ;
      RECT 22.35 4.807 22.37 5.118 ;
      RECT 22.34 4.82 22.35 5.12 ;
      RECT 22.315 4.835 22.34 5.123 ;
      RECT 22.295 4.852 22.315 5.127 ;
      RECT 22.255 4.88 22.295 5.133 ;
      RECT 22.19 4.927 22.255 5.142 ;
      RECT 22.175 4.96 22.19 5.15 ;
      RECT 22.17 4.967 22.175 5.152 ;
      RECT 22.12 4.992 22.17 5.157 ;
      RECT 22.105 5.016 22.12 5.164 ;
      RECT 22.055 5.021 22.105 5.165 ;
      RECT 21.969 5.025 22.055 5.165 ;
      RECT 21.883 5.025 21.969 5.165 ;
      RECT 21.797 5.025 21.883 5.166 ;
      RECT 21.711 5.025 21.797 5.166 ;
      RECT 21.625 5.025 21.711 5.166 ;
      RECT 21.559 5.025 21.625 5.166 ;
      RECT 21.473 5.025 21.559 5.167 ;
      RECT 21.387 5.025 21.473 5.167 ;
      RECT 21.301 5.026 21.387 5.168 ;
      RECT 21.215 5.026 21.301 5.168 ;
      RECT 21.129 5.026 21.215 5.168 ;
      RECT 21.043 5.026 21.129 5.169 ;
      RECT 20.957 5.026 21.043 5.169 ;
      RECT 20.871 5.027 20.957 5.17 ;
      RECT 20.785 5.027 20.871 5.17 ;
      RECT 20.765 5.027 20.785 5.17 ;
      RECT 20.679 5.027 20.765 5.17 ;
      RECT 20.593 5.027 20.679 5.17 ;
      RECT 20.507 5.028 20.593 5.17 ;
      RECT 20.421 5.028 20.507 5.17 ;
      RECT 20.335 5.028 20.421 5.17 ;
      RECT 20.249 5.029 20.335 5.17 ;
      RECT 20.163 5.029 20.249 5.17 ;
      RECT 20.077 5.029 20.163 5.17 ;
      RECT 19.991 5.029 20.077 5.17 ;
      RECT 19.905 5.03 19.991 5.17 ;
      RECT 19.855 5.027 19.905 5.17 ;
      RECT 19.845 5.025 19.855 5.169 ;
      RECT 19.841 5.025 19.845 5.168 ;
      RECT 19.755 5.02 19.841 5.163 ;
      RECT 19.733 5.013 19.755 5.157 ;
      RECT 19.647 5.004 19.733 5.151 ;
      RECT 19.561 4.991 19.647 5.142 ;
      RECT 19.475 4.977 19.561 5.132 ;
      RECT 19.43 4.967 19.475 5.125 ;
      RECT 19.41 4.255 19.43 4.533 ;
      RECT 19.41 4.96 19.43 5.121 ;
      RECT 19.38 4.255 19.41 4.555 ;
      RECT 19.37 4.927 19.41 5.118 ;
      RECT 19.365 4.255 19.38 4.575 ;
      RECT 19.365 4.892 19.37 5.116 ;
      RECT 19.36 4.255 19.365 4.7 ;
      RECT 19.36 4.852 19.365 5.116 ;
      RECT 19.35 4.255 19.36 5.116 ;
      RECT 19.275 4.255 19.35 5.11 ;
      RECT 19.245 4.255 19.275 5.1 ;
      RECT 19.24 4.255 19.245 5.092 ;
      RECT 19.235 4.297 19.24 5.085 ;
      RECT 19.225 4.366 19.235 5.076 ;
      RECT 19.22 4.436 19.225 5.028 ;
      RECT 19.215 4.5 19.22 4.925 ;
      RECT 19.21 4.535 19.215 4.88 ;
      RECT 19.208 4.572 19.21 4.772 ;
      RECT 19.205 4.58 19.208 4.765 ;
      RECT 19.2 4.645 19.205 4.708 ;
      RECT 23.275 3.735 23.555 4.015 ;
      RECT 23.265 3.735 23.555 3.878 ;
      RECT 23.22 3.6 23.48 3.86 ;
      RECT 23.22 3.715 23.535 3.86 ;
      RECT 23.22 3.685 23.53 3.86 ;
      RECT 23.22 3.672 23.52 3.86 ;
      RECT 23.22 3.662 23.515 3.86 ;
      RECT 19.195 3.645 19.455 3.905 ;
      RECT 22.965 3.195 23.225 3.455 ;
      RECT 22.955 3.22 23.225 3.415 ;
      RECT 22.95 3.22 22.955 3.414 ;
      RECT 22.88 3.215 22.95 3.406 ;
      RECT 22.795 3.202 22.88 3.389 ;
      RECT 22.791 3.194 22.795 3.379 ;
      RECT 22.705 3.187 22.791 3.369 ;
      RECT 22.696 3.179 22.705 3.359 ;
      RECT 22.61 3.172 22.696 3.347 ;
      RECT 22.59 3.163 22.61 3.333 ;
      RECT 22.535 3.158 22.59 3.325 ;
      RECT 22.525 3.152 22.535 3.319 ;
      RECT 22.505 3.15 22.525 3.315 ;
      RECT 22.497 3.149 22.505 3.311 ;
      RECT 22.411 3.141 22.497 3.3 ;
      RECT 22.325 3.127 22.411 3.28 ;
      RECT 22.265 3.115 22.325 3.265 ;
      RECT 22.255 3.11 22.265 3.26 ;
      RECT 22.205 3.11 22.255 3.262 ;
      RECT 22.158 3.112 22.205 3.266 ;
      RECT 22.072 3.119 22.158 3.271 ;
      RECT 21.986 3.127 22.072 3.277 ;
      RECT 21.9 3.136 21.986 3.283 ;
      RECT 21.841 3.142 21.9 3.288 ;
      RECT 21.755 3.147 21.841 3.294 ;
      RECT 21.68 3.152 21.755 3.3 ;
      RECT 21.641 3.154 21.68 3.305 ;
      RECT 21.555 3.151 21.641 3.31 ;
      RECT 21.47 3.149 21.555 3.317 ;
      RECT 21.438 3.148 21.47 3.32 ;
      RECT 21.352 3.147 21.438 3.321 ;
      RECT 21.266 3.146 21.352 3.322 ;
      RECT 21.18 3.145 21.266 3.322 ;
      RECT 21.094 3.144 21.18 3.323 ;
      RECT 21.008 3.143 21.094 3.324 ;
      RECT 20.922 3.142 21.008 3.325 ;
      RECT 20.836 3.141 20.922 3.325 ;
      RECT 20.75 3.14 20.836 3.326 ;
      RECT 20.7 3.14 20.75 3.327 ;
      RECT 20.686 3.141 20.7 3.327 ;
      RECT 20.6 3.148 20.686 3.328 ;
      RECT 20.526 3.159 20.6 3.329 ;
      RECT 20.44 3.168 20.526 3.33 ;
      RECT 20.405 3.175 20.44 3.345 ;
      RECT 20.38 3.178 20.405 3.375 ;
      RECT 20.355 3.187 20.38 3.404 ;
      RECT 20.345 3.198 20.355 3.424 ;
      RECT 20.335 3.206 20.345 3.438 ;
      RECT 20.33 3.212 20.335 3.448 ;
      RECT 20.305 3.229 20.33 3.465 ;
      RECT 20.29 3.251 20.305 3.493 ;
      RECT 20.26 3.277 20.29 3.523 ;
      RECT 20.24 3.306 20.26 3.553 ;
      RECT 20.235 3.321 20.24 3.57 ;
      RECT 20.215 3.336 20.235 3.585 ;
      RECT 20.205 3.354 20.215 3.603 ;
      RECT 20.195 3.365 20.205 3.618 ;
      RECT 20.145 3.397 20.195 3.644 ;
      RECT 20.14 3.427 20.145 3.664 ;
      RECT 20.13 3.44 20.14 3.67 ;
      RECT 20.121 3.45 20.13 3.678 ;
      RECT 20.11 3.461 20.121 3.686 ;
      RECT 20.105 3.471 20.11 3.692 ;
      RECT 20.09 3.492 20.105 3.699 ;
      RECT 20.075 3.522 20.09 3.707 ;
      RECT 20.04 3.552 20.075 3.713 ;
      RECT 20.015 3.57 20.04 3.72 ;
      RECT 19.965 3.578 20.015 3.729 ;
      RECT 19.94 3.583 19.965 3.738 ;
      RECT 19.885 3.589 19.94 3.748 ;
      RECT 19.88 3.594 19.885 3.756 ;
      RECT 19.866 3.597 19.88 3.758 ;
      RECT 19.78 3.609 19.866 3.77 ;
      RECT 19.77 3.621 19.78 3.783 ;
      RECT 19.685 3.634 19.77 3.795 ;
      RECT 19.641 3.651 19.685 3.809 ;
      RECT 19.555 3.668 19.641 3.825 ;
      RECT 19.525 3.682 19.555 3.839 ;
      RECT 19.515 3.687 19.525 3.844 ;
      RECT 19.455 3.69 19.515 3.853 ;
      RECT 22.345 3.96 22.605 4.22 ;
      RECT 22.345 3.96 22.625 4.073 ;
      RECT 22.345 3.96 22.65 4.04 ;
      RECT 22.345 3.96 22.655 4.02 ;
      RECT 22.395 3.735 22.675 4.015 ;
      RECT 21.95 4.47 22.21 4.73 ;
      RECT 21.94 4.327 22.135 4.668 ;
      RECT 21.935 4.435 22.15 4.66 ;
      RECT 21.93 4.485 22.21 4.65 ;
      RECT 21.92 4.562 22.21 4.635 ;
      RECT 21.94 4.41 22.15 4.668 ;
      RECT 21.95 4.285 22.135 4.73 ;
      RECT 21.95 4.18 22.115 4.73 ;
      RECT 21.96 4.167 22.115 4.73 ;
      RECT 21.96 4.125 22.105 4.73 ;
      RECT 21.965 4.05 22.105 4.73 ;
      RECT 21.995 3.7 22.105 4.73 ;
      RECT 22 3.43 22.125 4.053 ;
      RECT 21.97 4.005 22.125 4.053 ;
      RECT 21.985 3.807 22.105 4.73 ;
      RECT 21.975 3.917 22.125 4.053 ;
      RECT 22 3.43 22.14 3.91 ;
      RECT 22 3.43 22.16 3.785 ;
      RECT 21.965 3.43 22.225 3.69 ;
      RECT 21.435 3.735 21.715 4.015 ;
      RECT 21.42 3.735 21.715 3.995 ;
      RECT 19.475 4.6 19.735 4.86 ;
      RECT 21.26 4.455 21.52 4.715 ;
      RECT 21.24 4.475 21.52 4.69 ;
      RECT 21.197 4.475 21.24 4.689 ;
      RECT 21.111 4.476 21.197 4.686 ;
      RECT 21.025 4.477 21.111 4.682 ;
      RECT 20.95 4.479 21.025 4.679 ;
      RECT 20.927 4.48 20.95 4.677 ;
      RECT 20.841 4.481 20.927 4.675 ;
      RECT 20.755 4.482 20.841 4.672 ;
      RECT 20.731 4.483 20.755 4.67 ;
      RECT 20.645 4.485 20.731 4.667 ;
      RECT 20.56 4.487 20.645 4.668 ;
      RECT 20.503 4.488 20.56 4.674 ;
      RECT 20.417 4.49 20.503 4.684 ;
      RECT 20.331 4.493 20.417 4.697 ;
      RECT 20.245 4.495 20.331 4.709 ;
      RECT 20.231 4.496 20.245 4.716 ;
      RECT 20.145 4.497 20.231 4.724 ;
      RECT 20.105 4.499 20.145 4.733 ;
      RECT 20.096 4.5 20.105 4.736 ;
      RECT 20.01 4.508 20.096 4.742 ;
      RECT 19.99 4.517 20.01 4.75 ;
      RECT 19.905 4.532 19.99 4.758 ;
      RECT 19.845 4.555 19.905 4.769 ;
      RECT 19.835 4.567 19.845 4.774 ;
      RECT 19.795 4.577 19.835 4.778 ;
      RECT 19.74 4.594 19.795 4.786 ;
      RECT 19.735 4.604 19.74 4.79 ;
      RECT 20.801 3.735 20.86 4.132 ;
      RECT 20.715 3.735 20.92 4.123 ;
      RECT 20.71 3.765 20.92 4.118 ;
      RECT 20.676 3.765 20.92 4.116 ;
      RECT 20.59 3.765 20.92 4.11 ;
      RECT 20.545 3.765 20.94 4.088 ;
      RECT 20.545 3.765 20.96 4.043 ;
      RECT 20.505 3.765 20.96 4.033 ;
      RECT 20.715 3.735 20.995 4.015 ;
      RECT 20.45 3.735 20.71 3.995 ;
      RECT 18.275 4.295 18.555 4.575 ;
      RECT 18.245 4.257 18.5 4.56 ;
      RECT 18.24 4.258 18.5 4.558 ;
      RECT 18.235 4.259 18.5 4.552 ;
      RECT 18.23 4.262 18.5 4.545 ;
      RECT 18.225 4.295 18.555 4.538 ;
      RECT 18.195 4.265 18.5 4.525 ;
      RECT 18.195 4.292 18.52 4.525 ;
      RECT 18.195 4.282 18.515 4.525 ;
      RECT 18.195 4.267 18.51 4.525 ;
      RECT 18.275 4.254 18.49 4.575 ;
      RECT 18.361 4.252 18.49 4.575 ;
      RECT 18.447 4.25 18.475 4.575 ;
      RECT 88.515 9.325 88.885 9.695 ;
      RECT 72.73 9.325 73.1 9.695 ;
      RECT 56.945 9.325 57.315 9.695 ;
      RECT 41.17 9.325 41.54 9.695 ;
      RECT 25.39 9.325 25.76 9.695 ;
    LAYER via1 ;
      RECT 96.25 9.66 96.4 9.81 ;
      RECT 96.205 7.325 96.355 7.475 ;
      RECT 93.88 9.025 94.03 9.175 ;
      RECT 93.865 3.36 94.015 3.51 ;
      RECT 93.075 3.745 93.225 3.895 ;
      RECT 93.075 8.61 93.225 8.76 ;
      RECT 91.43 2.735 91.58 2.885 ;
      RECT 91.115 4.255 91.265 4.405 ;
      RECT 90.215 3.585 90.365 3.735 ;
      RECT 89.265 8.995 89.415 9.145 ;
      RECT 89.015 3.85 89.165 4 ;
      RECT 88.68 4.57 88.83 4.72 ;
      RECT 88.625 9.435 88.775 9.585 ;
      RECT 88.6 3.41 88.75 3.56 ;
      RECT 87.165 3.805 87.315 3.955 ;
      RECT 86.4 3.655 86.55 3.805 ;
      RECT 86.145 3.25 86.295 3.4 ;
      RECT 85.525 4.015 85.675 4.165 ;
      RECT 85.145 3.485 85.295 3.635 ;
      RECT 85.13 4.525 85.28 4.675 ;
      RECT 84.6 3.79 84.75 3.94 ;
      RECT 84.44 4.51 84.59 4.66 ;
      RECT 83.63 3.79 83.78 3.94 ;
      RECT 82.815 3.27 82.965 3.42 ;
      RECT 82.655 4.655 82.805 4.805 ;
      RECT 82.42 4.31 82.57 4.46 ;
      RECT 82.375 3.7 82.525 3.85 ;
      RECT 81.375 4.32 81.525 4.47 ;
      RECT 80.44 9.04 80.59 9.19 ;
      RECT 80.42 7.325 80.57 7.475 ;
      RECT 78.095 9.025 78.245 9.175 ;
      RECT 78.08 3.36 78.23 3.51 ;
      RECT 77.29 3.745 77.44 3.895 ;
      RECT 77.29 8.61 77.44 8.76 ;
      RECT 75.645 2.735 75.795 2.885 ;
      RECT 75.33 4.255 75.48 4.405 ;
      RECT 74.43 3.585 74.58 3.735 ;
      RECT 73.48 8.995 73.63 9.145 ;
      RECT 73.23 3.85 73.38 4 ;
      RECT 72.895 4.57 73.045 4.72 ;
      RECT 72.84 9.435 72.99 9.585 ;
      RECT 72.815 3.41 72.965 3.56 ;
      RECT 71.38 3.805 71.53 3.955 ;
      RECT 70.615 3.655 70.765 3.805 ;
      RECT 70.36 3.25 70.51 3.4 ;
      RECT 69.74 4.015 69.89 4.165 ;
      RECT 69.36 3.485 69.51 3.635 ;
      RECT 69.345 4.525 69.495 4.675 ;
      RECT 68.815 3.79 68.965 3.94 ;
      RECT 68.655 4.51 68.805 4.66 ;
      RECT 67.845 3.79 67.995 3.94 ;
      RECT 67.03 3.27 67.18 3.42 ;
      RECT 66.87 4.655 67.02 4.805 ;
      RECT 66.635 4.31 66.785 4.46 ;
      RECT 66.59 3.7 66.74 3.85 ;
      RECT 65.59 4.32 65.74 4.47 ;
      RECT 64.655 9.04 64.805 9.19 ;
      RECT 64.635 7.325 64.785 7.475 ;
      RECT 62.31 9.025 62.46 9.175 ;
      RECT 62.295 3.36 62.445 3.51 ;
      RECT 61.505 3.745 61.655 3.895 ;
      RECT 61.505 8.61 61.655 8.76 ;
      RECT 59.86 2.735 60.01 2.885 ;
      RECT 59.545 4.255 59.695 4.405 ;
      RECT 58.645 3.585 58.795 3.735 ;
      RECT 57.75 9 57.9 9.15 ;
      RECT 57.445 3.85 57.595 4 ;
      RECT 57.11 4.57 57.26 4.72 ;
      RECT 57.055 9.435 57.205 9.585 ;
      RECT 57.03 3.41 57.18 3.56 ;
      RECT 55.595 3.805 55.745 3.955 ;
      RECT 54.83 3.655 54.98 3.805 ;
      RECT 54.575 3.25 54.725 3.4 ;
      RECT 53.955 4.015 54.105 4.165 ;
      RECT 53.575 3.485 53.725 3.635 ;
      RECT 53.56 4.525 53.71 4.675 ;
      RECT 53.03 3.79 53.18 3.94 ;
      RECT 52.87 4.51 53.02 4.66 ;
      RECT 52.06 3.79 52.21 3.94 ;
      RECT 51.245 3.27 51.395 3.42 ;
      RECT 51.085 4.655 51.235 4.805 ;
      RECT 50.85 4.31 51 4.46 ;
      RECT 50.805 3.7 50.955 3.85 ;
      RECT 49.805 4.32 49.955 4.47 ;
      RECT 48.925 9.045 49.075 9.195 ;
      RECT 48.86 7.325 49.01 7.475 ;
      RECT 46.535 9.025 46.685 9.175 ;
      RECT 46.52 3.36 46.67 3.51 ;
      RECT 45.73 3.745 45.88 3.895 ;
      RECT 45.73 8.61 45.88 8.76 ;
      RECT 44.085 2.735 44.235 2.885 ;
      RECT 43.77 4.255 43.92 4.405 ;
      RECT 42.87 3.585 43.02 3.735 ;
      RECT 41.97 8.995 42.12 9.145 ;
      RECT 41.67 3.85 41.82 4 ;
      RECT 41.335 4.57 41.485 4.72 ;
      RECT 41.28 9.435 41.43 9.585 ;
      RECT 41.255 3.41 41.405 3.56 ;
      RECT 39.82 3.805 39.97 3.955 ;
      RECT 39.055 3.655 39.205 3.805 ;
      RECT 38.8 3.25 38.95 3.4 ;
      RECT 38.18 4.015 38.33 4.165 ;
      RECT 37.8 3.485 37.95 3.635 ;
      RECT 37.785 4.525 37.935 4.675 ;
      RECT 37.255 3.79 37.405 3.94 ;
      RECT 37.095 4.51 37.245 4.66 ;
      RECT 36.285 3.79 36.435 3.94 ;
      RECT 35.47 3.27 35.62 3.42 ;
      RECT 35.31 4.655 35.46 4.805 ;
      RECT 35.075 4.31 35.225 4.46 ;
      RECT 35.03 3.7 35.18 3.85 ;
      RECT 34.03 4.32 34.18 4.47 ;
      RECT 33.145 9.04 33.295 9.19 ;
      RECT 33.08 7.325 33.23 7.475 ;
      RECT 30.755 9.025 30.905 9.175 ;
      RECT 30.74 3.36 30.89 3.51 ;
      RECT 29.95 3.745 30.1 3.895 ;
      RECT 29.95 8.61 30.1 8.76 ;
      RECT 28.305 2.735 28.455 2.885 ;
      RECT 27.99 4.255 28.14 4.405 ;
      RECT 27.09 3.585 27.24 3.735 ;
      RECT 26.16 8.99 26.31 9.14 ;
      RECT 25.89 3.85 26.04 4 ;
      RECT 25.555 4.57 25.705 4.72 ;
      RECT 25.5 9.435 25.65 9.585 ;
      RECT 25.475 3.41 25.625 3.56 ;
      RECT 24.04 3.805 24.19 3.955 ;
      RECT 23.275 3.655 23.425 3.805 ;
      RECT 23.02 3.25 23.17 3.4 ;
      RECT 22.4 4.015 22.55 4.165 ;
      RECT 22.02 3.485 22.17 3.635 ;
      RECT 22.005 4.525 22.155 4.675 ;
      RECT 21.475 3.79 21.625 3.94 ;
      RECT 21.315 4.51 21.465 4.66 ;
      RECT 20.505 3.79 20.655 3.94 ;
      RECT 19.69 3.27 19.84 3.42 ;
      RECT 19.53 4.655 19.68 4.805 ;
      RECT 19.295 4.31 19.445 4.46 ;
      RECT 19.25 3.7 19.4 3.85 ;
      RECT 18.25 4.32 18.4 4.47 ;
      RECT 16.61 9.38 16.76 9.53 ;
      RECT 16.235 8.64 16.385 8.79 ;
    LAYER met1 ;
      RECT 96.12 10.05 96.415 10.28 ;
      RECT 96.18 9.56 96.355 10.28 ;
      RECT 96.15 9.56 96.5 9.91 ;
      RECT 96.18 8.57 96.35 10.28 ;
      RECT 96.12 8.57 96.41 8.8 ;
      RECT 96.14 7.215 96.42 7.585 ;
      RECT 96.095 7.215 96.445 7.565 ;
      RECT 95.125 10.055 95.42 10.285 ;
      RECT 95.185 8.575 95.355 10.285 ;
      RECT 95.125 8.575 95.415 8.805 ;
      RECT 95.125 8.61 95.98 8.77 ;
      RECT 95.81 8.2 95.98 8.77 ;
      RECT 95.125 8.605 95.52 8.77 ;
      RECT 95.75 8.2 96.04 8.43 ;
      RECT 95.75 8.23 96.21 8.4 ;
      RECT 95.71 4.03 96.035 4.26 ;
      RECT 95.71 4.06 96.205 4.23 ;
      RECT 95.71 3.69 95.9 4.26 ;
      RECT 95.125 3.655 95.415 3.885 ;
      RECT 95.125 3.69 95.9 3.86 ;
      RECT 95.185 2.175 95.355 3.885 ;
      RECT 95.125 2.175 95.42 2.405 ;
      RECT 94.755 4.025 95.045 4.255 ;
      RECT 94.755 4.055 95.215 4.225 ;
      RECT 94.82 2.95 94.985 4.255 ;
      RECT 93.335 2.915 93.625 3.145 ;
      RECT 93.335 2.95 94.985 3.12 ;
      RECT 93.395 2.175 93.565 3.145 ;
      RECT 93.335 2.175 93.625 2.405 ;
      RECT 93.335 10.055 93.625 10.285 ;
      RECT 93.395 9.315 93.565 10.285 ;
      RECT 93.395 9.405 94.985 9.575 ;
      RECT 94.815 8.205 94.985 9.575 ;
      RECT 93.335 9.315 93.625 9.545 ;
      RECT 94.755 8.205 95.045 8.435 ;
      RECT 94.755 8.235 95.215 8.405 ;
      RECT 93.765 3.26 94.115 3.61 ;
      RECT 91.43 3.32 94.115 3.49 ;
      RECT 93.595 3.315 94.115 3.49 ;
      RECT 91.43 2.635 91.6 3.49 ;
      RECT 91.33 2.635 91.68 2.985 ;
      RECT 93.79 8.94 94.115 9.265 ;
      RECT 89.165 8.895 89.515 9.245 ;
      RECT 93.765 8.945 94.115 9.175 ;
      RECT 88.985 8.945 89.515 9.175 ;
      RECT 93.595 8.97 94.115 9.145 ;
      RECT 88.815 8.975 89.515 9.145 ;
      RECT 88.985 8.97 94.115 9.14 ;
      RECT 92.99 3.66 93.31 3.98 ;
      RECT 92.965 3.655 93.255 3.885 ;
      RECT 92.89 3.685 93.31 3.86 ;
      RECT 92.79 3.685 93.31 3.855 ;
      RECT 92.99 8.54 93.31 8.83 ;
      RECT 92.965 8.575 93.31 8.805 ;
      RECT 92.79 8.605 93.31 8.775 ;
      RECT 89.625 3.76 89.81 3.97 ;
      RECT 89.615 3.765 89.825 3.963 ;
      RECT 89.615 3.765 89.911 3.94 ;
      RECT 89.615 3.765 89.97 3.915 ;
      RECT 89.615 3.765 90.025 3.895 ;
      RECT 89.615 3.765 90.035 3.883 ;
      RECT 89.615 3.765 90.23 3.822 ;
      RECT 89.615 3.765 90.26 3.805 ;
      RECT 89.615 3.765 90.28 3.795 ;
      RECT 90.16 3.53 90.42 3.79 ;
      RECT 90.145 3.62 90.16 3.837 ;
      RECT 89.68 3.752 90.42 3.79 ;
      RECT 90.131 3.631 90.145 3.843 ;
      RECT 89.72 3.745 90.42 3.79 ;
      RECT 90.045 3.671 90.131 3.862 ;
      RECT 89.97 3.732 90.42 3.79 ;
      RECT 90.04 3.707 90.045 3.879 ;
      RECT 90.025 3.717 90.42 3.79 ;
      RECT 90.035 3.712 90.04 3.881 ;
      RECT 88.96 3.795 89.065 4.055 ;
      RECT 89.775 3.32 89.78 3.545 ;
      RECT 89.905 3.32 89.96 3.53 ;
      RECT 89.96 3.325 89.97 3.523 ;
      RECT 89.866 3.32 89.905 3.533 ;
      RECT 89.78 3.32 89.866 3.54 ;
      RECT 89.76 3.325 89.775 3.546 ;
      RECT 89.75 3.365 89.76 3.548 ;
      RECT 89.72 3.375 89.75 3.55 ;
      RECT 89.715 3.38 89.72 3.552 ;
      RECT 89.69 3.385 89.715 3.554 ;
      RECT 89.675 3.39 89.69 3.556 ;
      RECT 89.66 3.392 89.675 3.558 ;
      RECT 89.655 3.397 89.66 3.56 ;
      RECT 89.605 3.405 89.655 3.563 ;
      RECT 89.58 3.414 89.605 3.568 ;
      RECT 89.57 3.421 89.58 3.573 ;
      RECT 89.565 3.424 89.57 3.577 ;
      RECT 89.545 3.427 89.565 3.586 ;
      RECT 89.515 3.435 89.545 3.606 ;
      RECT 89.486 3.448 89.515 3.628 ;
      RECT 89.4 3.482 89.486 3.672 ;
      RECT 89.395 3.508 89.4 3.71 ;
      RECT 89.39 3.512 89.395 3.719 ;
      RECT 89.355 3.525 89.39 3.752 ;
      RECT 89.345 3.539 89.355 3.79 ;
      RECT 89.34 3.543 89.345 3.803 ;
      RECT 89.335 3.547 89.34 3.808 ;
      RECT 89.325 3.555 89.335 3.82 ;
      RECT 89.32 3.562 89.325 3.835 ;
      RECT 89.295 3.575 89.32 3.86 ;
      RECT 89.255 3.604 89.295 3.915 ;
      RECT 89.24 3.629 89.255 3.97 ;
      RECT 89.23 3.64 89.24 3.993 ;
      RECT 89.225 3.647 89.23 4.005 ;
      RECT 89.22 3.651 89.225 4.013 ;
      RECT 89.165 3.679 89.22 4.055 ;
      RECT 89.145 3.715 89.165 4.055 ;
      RECT 89.13 3.73 89.145 4.055 ;
      RECT 89.075 3.762 89.13 4.055 ;
      RECT 89.065 3.792 89.075 4.055 ;
      RECT 88.675 3.407 88.86 3.645 ;
      RECT 88.66 3.409 88.87 3.64 ;
      RECT 88.545 3.355 88.805 3.615 ;
      RECT 88.54 3.392 88.805 3.569 ;
      RECT 88.535 3.402 88.805 3.566 ;
      RECT 88.53 3.442 88.87 3.56 ;
      RECT 88.525 3.475 88.87 3.55 ;
      RECT 88.535 3.417 88.885 3.488 ;
      RECT 88.832 4.515 88.845 5.045 ;
      RECT 88.746 4.515 88.845 5.044 ;
      RECT 88.746 4.515 88.85 5.043 ;
      RECT 88.66 4.515 88.85 5.041 ;
      RECT 88.655 4.515 88.85 5.038 ;
      RECT 88.655 4.515 88.86 5.036 ;
      RECT 88.65 4.807 88.86 5.033 ;
      RECT 88.65 4.817 88.865 5.03 ;
      RECT 88.65 4.885 88.87 5.026 ;
      RECT 88.64 4.89 88.87 5.025 ;
      RECT 88.64 4.982 88.875 5.022 ;
      RECT 88.625 4.515 88.885 4.775 ;
      RECT 88.555 10.055 88.845 10.285 ;
      RECT 88.615 9.315 88.785 10.285 ;
      RECT 88.53 9.34 88.87 9.685 ;
      RECT 88.555 9.315 88.845 9.685 ;
      RECT 87.855 3.505 87.9 5.04 ;
      RECT 88.055 3.505 88.085 3.72 ;
      RECT 86.43 3.245 86.55 3.455 ;
      RECT 86.09 3.195 86.35 3.455 ;
      RECT 86.09 3.24 86.385 3.445 ;
      RECT 88.095 3.521 88.1 3.575 ;
      RECT 88.09 3.514 88.095 3.708 ;
      RECT 88.085 3.508 88.09 3.715 ;
      RECT 88.04 3.505 88.055 3.728 ;
      RECT 88.035 3.505 88.04 3.75 ;
      RECT 88.03 3.505 88.035 3.798 ;
      RECT 88.025 3.505 88.03 3.818 ;
      RECT 88.015 3.505 88.025 3.925 ;
      RECT 88.01 3.505 88.015 3.988 ;
      RECT 88.005 3.505 88.01 4.045 ;
      RECT 88 3.505 88.005 4.053 ;
      RECT 87.985 3.505 88 4.16 ;
      RECT 87.975 3.505 87.985 4.295 ;
      RECT 87.965 3.505 87.975 4.405 ;
      RECT 87.955 3.505 87.965 4.462 ;
      RECT 87.95 3.505 87.955 4.502 ;
      RECT 87.945 3.505 87.95 4.538 ;
      RECT 87.935 3.505 87.945 4.578 ;
      RECT 87.93 3.505 87.935 4.62 ;
      RECT 87.91 3.505 87.93 4.685 ;
      RECT 87.915 4.83 87.92 5.01 ;
      RECT 87.91 4.812 87.915 5.018 ;
      RECT 87.905 3.505 87.91 4.748 ;
      RECT 87.905 4.792 87.91 5.025 ;
      RECT 87.9 3.505 87.905 5.035 ;
      RECT 87.845 3.505 87.855 3.805 ;
      RECT 87.85 4.052 87.855 5.04 ;
      RECT 87.845 4.117 87.85 5.04 ;
      RECT 87.84 3.506 87.845 3.795 ;
      RECT 87.835 4.182 87.845 5.04 ;
      RECT 87.83 3.507 87.84 3.785 ;
      RECT 87.82 4.295 87.835 5.04 ;
      RECT 87.825 3.508 87.83 3.775 ;
      RECT 87.805 3.509 87.825 3.753 ;
      RECT 87.81 4.392 87.82 5.04 ;
      RECT 87.805 4.467 87.81 5.04 ;
      RECT 87.795 3.508 87.805 3.73 ;
      RECT 87.8 4.51 87.805 5.04 ;
      RECT 87.795 4.537 87.8 5.04 ;
      RECT 87.785 3.506 87.795 3.718 ;
      RECT 87.79 4.58 87.795 5.04 ;
      RECT 87.785 4.607 87.79 5.04 ;
      RECT 87.775 3.505 87.785 3.705 ;
      RECT 87.78 4.622 87.785 5.04 ;
      RECT 87.74 4.68 87.78 5.04 ;
      RECT 87.77 3.504 87.775 3.69 ;
      RECT 87.765 3.502 87.77 3.683 ;
      RECT 87.755 3.499 87.765 3.673 ;
      RECT 87.75 3.496 87.755 3.658 ;
      RECT 87.735 3.492 87.75 3.651 ;
      RECT 87.73 4.735 87.74 5.04 ;
      RECT 87.73 3.489 87.735 3.646 ;
      RECT 87.715 3.485 87.73 3.64 ;
      RECT 87.725 4.752 87.73 5.04 ;
      RECT 87.715 4.815 87.725 5.04 ;
      RECT 87.635 3.47 87.715 3.62 ;
      RECT 87.71 4.822 87.715 5.035 ;
      RECT 87.705 4.83 87.71 5.025 ;
      RECT 87.625 3.456 87.635 3.604 ;
      RECT 87.61 3.452 87.625 3.602 ;
      RECT 87.6 3.447 87.61 3.598 ;
      RECT 87.575 3.44 87.6 3.59 ;
      RECT 87.57 3.435 87.575 3.585 ;
      RECT 87.56 3.435 87.57 3.583 ;
      RECT 87.55 3.433 87.56 3.581 ;
      RECT 87.52 3.425 87.55 3.575 ;
      RECT 87.505 3.417 87.52 3.568 ;
      RECT 87.485 3.412 87.505 3.561 ;
      RECT 87.48 3.408 87.485 3.556 ;
      RECT 87.45 3.401 87.48 3.55 ;
      RECT 87.425 3.392 87.45 3.54 ;
      RECT 87.395 3.385 87.425 3.532 ;
      RECT 87.37 3.375 87.395 3.523 ;
      RECT 87.355 3.367 87.37 3.517 ;
      RECT 87.33 3.362 87.355 3.512 ;
      RECT 87.32 3.358 87.33 3.507 ;
      RECT 87.3 3.353 87.32 3.502 ;
      RECT 87.265 3.348 87.3 3.495 ;
      RECT 87.205 3.343 87.265 3.488 ;
      RECT 87.192 3.339 87.205 3.486 ;
      RECT 87.106 3.334 87.192 3.483 ;
      RECT 87.02 3.324 87.106 3.479 ;
      RECT 86.979 3.317 87.02 3.476 ;
      RECT 86.893 3.31 86.979 3.473 ;
      RECT 86.807 3.3 86.893 3.469 ;
      RECT 86.721 3.29 86.807 3.464 ;
      RECT 86.635 3.28 86.721 3.46 ;
      RECT 86.625 3.265 86.635 3.458 ;
      RECT 86.615 3.25 86.625 3.458 ;
      RECT 86.55 3.245 86.615 3.457 ;
      RECT 86.385 3.242 86.43 3.45 ;
      RECT 87.63 4.147 87.635 4.338 ;
      RECT 87.625 4.142 87.63 4.345 ;
      RECT 87.611 4.14 87.625 4.351 ;
      RECT 87.525 4.14 87.611 4.353 ;
      RECT 87.521 4.14 87.525 4.356 ;
      RECT 87.435 4.14 87.521 4.374 ;
      RECT 87.425 4.145 87.435 4.393 ;
      RECT 87.415 4.2 87.425 4.397 ;
      RECT 87.39 4.215 87.415 4.404 ;
      RECT 87.35 4.235 87.39 4.417 ;
      RECT 87.345 4.247 87.35 4.427 ;
      RECT 87.33 4.253 87.345 4.432 ;
      RECT 87.325 4.258 87.33 4.436 ;
      RECT 87.305 4.265 87.325 4.441 ;
      RECT 87.235 4.29 87.305 4.458 ;
      RECT 87.195 4.318 87.235 4.478 ;
      RECT 87.19 4.328 87.195 4.486 ;
      RECT 87.17 4.335 87.19 4.488 ;
      RECT 87.165 4.342 87.17 4.491 ;
      RECT 87.135 4.35 87.165 4.494 ;
      RECT 87.13 4.355 87.135 4.498 ;
      RECT 87.056 4.359 87.13 4.506 ;
      RECT 86.97 4.368 87.056 4.522 ;
      RECT 86.966 4.373 86.97 4.531 ;
      RECT 86.88 4.378 86.966 4.541 ;
      RECT 86.84 4.386 86.88 4.553 ;
      RECT 86.79 4.392 86.84 4.56 ;
      RECT 86.705 4.401 86.79 4.575 ;
      RECT 86.63 4.412 86.705 4.593 ;
      RECT 86.595 4.419 86.63 4.603 ;
      RECT 86.52 4.427 86.595 4.608 ;
      RECT 86.465 4.436 86.52 4.608 ;
      RECT 86.44 4.441 86.465 4.606 ;
      RECT 86.43 4.444 86.44 4.604 ;
      RECT 86.395 4.446 86.43 4.602 ;
      RECT 86.365 4.448 86.395 4.598 ;
      RECT 86.32 4.447 86.365 4.594 ;
      RECT 86.3 4.442 86.32 4.591 ;
      RECT 86.25 4.427 86.3 4.588 ;
      RECT 86.24 4.412 86.25 4.583 ;
      RECT 86.19 4.397 86.24 4.573 ;
      RECT 86.14 4.372 86.19 4.553 ;
      RECT 86.13 4.357 86.14 4.535 ;
      RECT 86.125 4.355 86.13 4.529 ;
      RECT 86.105 4.35 86.125 4.524 ;
      RECT 86.1 4.342 86.105 4.518 ;
      RECT 86.085 4.336 86.1 4.511 ;
      RECT 86.08 4.331 86.085 4.503 ;
      RECT 86.06 4.326 86.08 4.495 ;
      RECT 86.045 4.319 86.06 4.488 ;
      RECT 86.03 4.313 86.045 4.479 ;
      RECT 86.025 4.307 86.03 4.472 ;
      RECT 85.98 4.282 86.025 4.458 ;
      RECT 85.965 4.252 85.98 4.44 ;
      RECT 85.95 4.235 85.965 4.431 ;
      RECT 85.925 4.215 85.95 4.419 ;
      RECT 85.885 4.185 85.925 4.399 ;
      RECT 85.875 4.155 85.885 4.384 ;
      RECT 85.86 4.145 85.875 4.377 ;
      RECT 85.805 4.11 85.86 4.356 ;
      RECT 85.79 4.073 85.805 4.335 ;
      RECT 85.78 4.06 85.79 4.327 ;
      RECT 85.73 4.03 85.78 4.309 ;
      RECT 85.715 3.96 85.73 4.29 ;
      RECT 85.67 3.96 85.715 4.273 ;
      RECT 85.645 3.96 85.67 4.255 ;
      RECT 85.635 3.96 85.645 4.248 ;
      RECT 85.556 3.96 85.635 4.241 ;
      RECT 85.47 3.96 85.556 4.233 ;
      RECT 85.455 3.992 85.47 4.228 ;
      RECT 85.38 4.002 85.455 4.224 ;
      RECT 85.36 4.012 85.38 4.219 ;
      RECT 85.335 4.012 85.36 4.216 ;
      RECT 85.325 4.002 85.335 4.215 ;
      RECT 85.315 3.975 85.325 4.214 ;
      RECT 85.275 3.97 85.315 4.212 ;
      RECT 85.23 3.97 85.275 4.208 ;
      RECT 85.205 3.97 85.23 4.203 ;
      RECT 85.155 3.97 85.205 4.19 ;
      RECT 85.115 3.975 85.125 4.175 ;
      RECT 85.125 3.97 85.155 4.18 ;
      RECT 87.11 3.75 87.37 4.01 ;
      RECT 87.105 3.772 87.37 3.968 ;
      RECT 86.345 3.6 86.565 3.965 ;
      RECT 86.327 3.687 86.565 3.964 ;
      RECT 86.31 3.692 86.565 3.961 ;
      RECT 86.31 3.692 86.585 3.96 ;
      RECT 86.28 3.702 86.585 3.958 ;
      RECT 86.275 3.717 86.585 3.954 ;
      RECT 86.275 3.717 86.59 3.953 ;
      RECT 86.27 3.775 86.59 3.951 ;
      RECT 86.27 3.775 86.6 3.948 ;
      RECT 86.265 3.84 86.6 3.943 ;
      RECT 86.345 3.6 86.605 3.86 ;
      RECT 85.09 3.43 85.35 3.69 ;
      RECT 85.09 3.473 85.436 3.664 ;
      RECT 85.09 3.473 85.48 3.663 ;
      RECT 85.09 3.473 85.5 3.661 ;
      RECT 85.09 3.473 85.6 3.66 ;
      RECT 85.09 3.473 85.62 3.658 ;
      RECT 85.09 3.473 85.63 3.653 ;
      RECT 85.5 3.44 85.69 3.65 ;
      RECT 85.5 3.442 85.695 3.648 ;
      RECT 85.49 3.447 85.7 3.64 ;
      RECT 85.436 3.471 85.7 3.64 ;
      RECT 85.48 3.465 85.49 3.662 ;
      RECT 85.49 3.445 85.695 3.648 ;
      RECT 84.445 4.505 84.65 4.735 ;
      RECT 84.385 4.455 84.44 4.715 ;
      RECT 84.445 4.455 84.645 4.735 ;
      RECT 85.415 4.77 85.42 4.797 ;
      RECT 85.405 4.68 85.415 4.802 ;
      RECT 85.4 4.602 85.405 4.808 ;
      RECT 85.39 4.592 85.4 4.815 ;
      RECT 85.385 4.582 85.39 4.821 ;
      RECT 85.375 4.577 85.385 4.823 ;
      RECT 85.36 4.569 85.375 4.831 ;
      RECT 85.345 4.56 85.36 4.843 ;
      RECT 85.335 4.552 85.345 4.853 ;
      RECT 85.3 4.47 85.335 4.871 ;
      RECT 85.265 4.47 85.3 4.89 ;
      RECT 85.25 4.47 85.265 4.898 ;
      RECT 85.195 4.47 85.25 4.898 ;
      RECT 85.161 4.47 85.195 4.889 ;
      RECT 85.075 4.47 85.161 4.865 ;
      RECT 85.065 4.53 85.075 4.847 ;
      RECT 85.025 4.532 85.065 4.838 ;
      RECT 85.02 4.534 85.025 4.828 ;
      RECT 85 4.536 85.02 4.823 ;
      RECT 84.99 4.539 85 4.818 ;
      RECT 84.98 4.54 84.99 4.813 ;
      RECT 84.956 4.541 84.98 4.805 ;
      RECT 84.87 4.546 84.956 4.783 ;
      RECT 84.815 4.545 84.87 4.756 ;
      RECT 84.8 4.538 84.815 4.743 ;
      RECT 84.765 4.533 84.8 4.739 ;
      RECT 84.71 4.525 84.765 4.738 ;
      RECT 84.65 4.512 84.71 4.736 ;
      RECT 84.44 4.455 84.445 4.723 ;
      RECT 84.515 3.825 84.7 4.035 ;
      RECT 84.505 3.83 84.715 4.028 ;
      RECT 84.545 3.735 84.805 3.995 ;
      RECT 84.5 3.892 84.805 3.918 ;
      RECT 83.845 3.685 83.85 4.485 ;
      RECT 83.79 3.735 83.82 4.485 ;
      RECT 83.78 3.735 83.785 4.045 ;
      RECT 83.765 3.735 83.77 4.04 ;
      RECT 83.31 3.78 83.325 3.995 ;
      RECT 83.24 3.78 83.325 3.99 ;
      RECT 84.505 3.36 84.575 3.57 ;
      RECT 84.575 3.367 84.585 3.565 ;
      RECT 84.471 3.36 84.505 3.577 ;
      RECT 84.385 3.36 84.471 3.601 ;
      RECT 84.375 3.365 84.385 3.62 ;
      RECT 84.37 3.377 84.375 3.623 ;
      RECT 84.355 3.392 84.37 3.627 ;
      RECT 84.35 3.41 84.355 3.631 ;
      RECT 84.31 3.42 84.35 3.64 ;
      RECT 84.295 3.427 84.31 3.652 ;
      RECT 84.28 3.432 84.295 3.657 ;
      RECT 84.265 3.435 84.28 3.662 ;
      RECT 84.255 3.437 84.265 3.666 ;
      RECT 84.22 3.444 84.255 3.674 ;
      RECT 84.185 3.452 84.22 3.688 ;
      RECT 84.175 3.458 84.185 3.697 ;
      RECT 84.17 3.46 84.175 3.699 ;
      RECT 84.15 3.463 84.17 3.705 ;
      RECT 84.12 3.47 84.15 3.716 ;
      RECT 84.11 3.476 84.12 3.723 ;
      RECT 84.085 3.479 84.11 3.73 ;
      RECT 84.075 3.483 84.085 3.738 ;
      RECT 84.07 3.484 84.075 3.76 ;
      RECT 84.065 3.485 84.07 3.775 ;
      RECT 84.06 3.486 84.065 3.79 ;
      RECT 84.055 3.487 84.06 3.805 ;
      RECT 84.05 3.488 84.055 3.835 ;
      RECT 84.04 3.49 84.05 3.868 ;
      RECT 84.025 3.494 84.04 3.915 ;
      RECT 84.015 3.497 84.025 3.96 ;
      RECT 84.01 3.5 84.015 3.988 ;
      RECT 84 3.502 84.01 4.015 ;
      RECT 83.995 3.505 84 4.05 ;
      RECT 83.965 3.51 83.995 4.108 ;
      RECT 83.96 3.515 83.965 4.193 ;
      RECT 83.955 3.517 83.96 4.228 ;
      RECT 83.95 3.519 83.955 4.31 ;
      RECT 83.945 3.521 83.95 4.398 ;
      RECT 83.935 3.523 83.945 4.48 ;
      RECT 83.92 3.537 83.935 4.485 ;
      RECT 83.885 3.582 83.92 4.485 ;
      RECT 83.875 3.622 83.885 4.485 ;
      RECT 83.86 3.65 83.875 4.485 ;
      RECT 83.855 3.667 83.86 4.485 ;
      RECT 83.85 3.675 83.855 4.485 ;
      RECT 83.84 3.69 83.845 4.485 ;
      RECT 83.835 3.697 83.84 4.485 ;
      RECT 83.825 3.717 83.835 4.485 ;
      RECT 83.82 3.73 83.825 4.485 ;
      RECT 83.785 3.735 83.79 4.07 ;
      RECT 83.77 4.125 83.79 4.485 ;
      RECT 83.77 3.735 83.78 4.043 ;
      RECT 83.765 4.165 83.77 4.485 ;
      RECT 83.715 3.735 83.765 4.038 ;
      RECT 83.76 4.202 83.765 4.485 ;
      RECT 83.75 4.225 83.76 4.485 ;
      RECT 83.745 4.27 83.75 4.485 ;
      RECT 83.735 4.28 83.745 4.478 ;
      RECT 83.661 3.735 83.715 4.032 ;
      RECT 83.575 3.735 83.661 4.025 ;
      RECT 83.526 3.782 83.575 4.018 ;
      RECT 83.44 3.79 83.526 4.011 ;
      RECT 83.425 3.787 83.44 4.006 ;
      RECT 83.411 3.78 83.425 4.005 ;
      RECT 83.325 3.78 83.411 4 ;
      RECT 83.23 3.785 83.24 3.985 ;
      RECT 82.82 3.215 82.835 3.615 ;
      RECT 83.015 3.215 83.02 3.475 ;
      RECT 82.76 3.215 82.805 3.475 ;
      RECT 83.215 4.52 83.22 4.725 ;
      RECT 83.21 4.51 83.215 4.73 ;
      RECT 83.205 4.497 83.21 4.735 ;
      RECT 83.2 4.477 83.205 4.735 ;
      RECT 83.175 4.43 83.2 4.735 ;
      RECT 83.14 4.345 83.175 4.735 ;
      RECT 83.135 4.282 83.14 4.735 ;
      RECT 83.13 4.267 83.135 4.735 ;
      RECT 83.115 4.227 83.13 4.735 ;
      RECT 83.11 4.202 83.115 4.735 ;
      RECT 83.1 4.185 83.11 4.735 ;
      RECT 83.065 4.107 83.1 4.735 ;
      RECT 83.06 4.05 83.065 4.735 ;
      RECT 83.055 4.037 83.06 4.735 ;
      RECT 83.045 4.015 83.055 4.735 ;
      RECT 83.035 3.98 83.045 4.735 ;
      RECT 83.025 3.95 83.035 4.735 ;
      RECT 83.015 3.865 83.025 4.378 ;
      RECT 83.022 4.51 83.025 4.735 ;
      RECT 83.02 4.52 83.022 4.735 ;
      RECT 83.01 4.53 83.02 4.73 ;
      RECT 83.005 3.215 83.015 3.61 ;
      RECT 83.01 3.742 83.015 4.353 ;
      RECT 83.005 3.64 83.01 4.336 ;
      RECT 82.995 3.215 83.005 4.312 ;
      RECT 82.99 3.215 82.995 4.283 ;
      RECT 82.985 3.215 82.99 4.273 ;
      RECT 82.965 3.215 82.985 4.235 ;
      RECT 82.96 3.215 82.965 4.193 ;
      RECT 82.955 3.215 82.96 4.173 ;
      RECT 82.925 3.215 82.955 4.123 ;
      RECT 82.915 3.215 82.925 4.07 ;
      RECT 82.91 3.215 82.915 4.043 ;
      RECT 82.905 3.215 82.91 4.028 ;
      RECT 82.895 3.215 82.905 4.005 ;
      RECT 82.885 3.215 82.895 3.98 ;
      RECT 82.88 3.215 82.885 3.92 ;
      RECT 82.87 3.215 82.88 3.858 ;
      RECT 82.865 3.215 82.87 3.778 ;
      RECT 82.86 3.215 82.865 3.743 ;
      RECT 82.855 3.215 82.86 3.718 ;
      RECT 82.85 3.215 82.855 3.703 ;
      RECT 82.845 3.215 82.85 3.673 ;
      RECT 82.84 3.215 82.845 3.65 ;
      RECT 82.835 3.215 82.84 3.623 ;
      RECT 82.805 3.215 82.82 3.61 ;
      RECT 81.96 4.75 82.145 4.96 ;
      RECT 81.95 4.755 82.16 4.953 ;
      RECT 81.95 4.755 82.18 4.925 ;
      RECT 81.95 4.755 82.195 4.904 ;
      RECT 81.95 4.755 82.21 4.902 ;
      RECT 81.95 4.755 82.22 4.901 ;
      RECT 81.95 4.755 82.25 4.898 ;
      RECT 82.6 4.6 82.86 4.86 ;
      RECT 82.56 4.647 82.86 4.843 ;
      RECT 82.551 4.655 82.56 4.846 ;
      RECT 82.145 4.748 82.86 4.843 ;
      RECT 82.465 4.673 82.551 4.853 ;
      RECT 82.16 4.745 82.86 4.843 ;
      RECT 82.406 4.695 82.465 4.865 ;
      RECT 82.18 4.741 82.86 4.843 ;
      RECT 82.32 4.707 82.406 4.876 ;
      RECT 82.195 4.737 82.86 4.843 ;
      RECT 82.265 4.72 82.32 4.888 ;
      RECT 82.21 4.735 82.86 4.843 ;
      RECT 82.25 4.726 82.265 4.894 ;
      RECT 82.22 4.731 82.86 4.843 ;
      RECT 82.365 4.255 82.625 4.515 ;
      RECT 82.365 4.275 82.735 4.485 ;
      RECT 82.365 4.28 82.745 4.48 ;
      RECT 82.556 3.694 82.635 3.925 ;
      RECT 82.47 3.697 82.685 3.92 ;
      RECT 82.465 3.697 82.685 3.915 ;
      RECT 82.465 3.702 82.695 3.913 ;
      RECT 82.44 3.702 82.695 3.91 ;
      RECT 82.44 3.71 82.705 3.908 ;
      RECT 82.32 3.645 82.58 3.905 ;
      RECT 82.32 3.692 82.63 3.905 ;
      RECT 81.575 4.265 81.58 4.525 ;
      RECT 81.405 4.035 81.41 4.525 ;
      RECT 81.29 4.275 81.295 4.5 ;
      RECT 82 3.37 82.005 3.58 ;
      RECT 82.005 3.375 82.02 3.575 ;
      RECT 81.94 3.37 82 3.588 ;
      RECT 81.925 3.37 81.94 3.598 ;
      RECT 81.875 3.37 81.925 3.615 ;
      RECT 81.855 3.37 81.875 3.638 ;
      RECT 81.84 3.37 81.855 3.65 ;
      RECT 81.82 3.37 81.84 3.66 ;
      RECT 81.81 3.375 81.82 3.669 ;
      RECT 81.805 3.385 81.81 3.674 ;
      RECT 81.8 3.397 81.805 3.678 ;
      RECT 81.79 3.42 81.8 3.683 ;
      RECT 81.785 3.435 81.79 3.687 ;
      RECT 81.78 3.452 81.785 3.69 ;
      RECT 81.775 3.46 81.78 3.693 ;
      RECT 81.765 3.465 81.775 3.697 ;
      RECT 81.76 3.472 81.765 3.702 ;
      RECT 81.75 3.477 81.76 3.706 ;
      RECT 81.725 3.489 81.75 3.717 ;
      RECT 81.705 3.506 81.725 3.733 ;
      RECT 81.68 3.523 81.705 3.755 ;
      RECT 81.645 3.546 81.68 3.813 ;
      RECT 81.625 3.568 81.645 3.875 ;
      RECT 81.62 3.578 81.625 3.91 ;
      RECT 81.61 3.585 81.62 3.948 ;
      RECT 81.605 3.592 81.61 3.968 ;
      RECT 81.6 3.603 81.605 4.005 ;
      RECT 81.595 3.611 81.6 4.07 ;
      RECT 81.585 3.622 81.595 4.123 ;
      RECT 81.58 3.64 81.585 4.193 ;
      RECT 81.575 3.65 81.58 4.23 ;
      RECT 81.57 3.66 81.575 4.525 ;
      RECT 81.565 3.672 81.57 4.525 ;
      RECT 81.56 3.682 81.565 4.525 ;
      RECT 81.55 3.692 81.56 4.525 ;
      RECT 81.54 3.715 81.55 4.525 ;
      RECT 81.525 3.75 81.54 4.525 ;
      RECT 81.485 3.812 81.525 4.525 ;
      RECT 81.48 3.865 81.485 4.525 ;
      RECT 81.455 3.9 81.48 4.525 ;
      RECT 81.44 3.945 81.455 4.525 ;
      RECT 81.435 3.967 81.44 4.525 ;
      RECT 81.425 3.98 81.435 4.525 ;
      RECT 81.415 4.005 81.425 4.525 ;
      RECT 81.41 4.027 81.415 4.525 ;
      RECT 81.385 4.065 81.405 4.525 ;
      RECT 81.345 4.122 81.385 4.525 ;
      RECT 81.34 4.172 81.345 4.525 ;
      RECT 81.335 4.19 81.34 4.525 ;
      RECT 81.33 4.202 81.335 4.525 ;
      RECT 81.32 4.22 81.33 4.525 ;
      RECT 81.31 4.24 81.32 4.5 ;
      RECT 81.305 4.257 81.31 4.5 ;
      RECT 81.295 4.27 81.305 4.5 ;
      RECT 81.265 4.28 81.29 4.5 ;
      RECT 81.255 4.287 81.265 4.5 ;
      RECT 81.24 4.297 81.255 4.495 ;
      RECT 80.335 10.05 80.63 10.28 ;
      RECT 80.395 8.57 80.565 10.28 ;
      RECT 80.34 8.94 80.69 9.29 ;
      RECT 80.335 8.57 80.625 8.8 ;
      RECT 80.355 7.215 80.635 7.585 ;
      RECT 80.31 7.215 80.66 7.565 ;
      RECT 79.34 10.055 79.635 10.285 ;
      RECT 79.4 8.575 79.57 10.285 ;
      RECT 79.34 8.575 79.63 8.805 ;
      RECT 79.34 8.61 80.195 8.77 ;
      RECT 80.025 8.2 80.195 8.77 ;
      RECT 79.34 8.605 79.735 8.77 ;
      RECT 79.965 8.2 80.255 8.43 ;
      RECT 79.965 8.23 80.425 8.4 ;
      RECT 79.925 4.03 80.25 4.26 ;
      RECT 79.925 4.06 80.42 4.23 ;
      RECT 79.925 3.69 80.115 4.26 ;
      RECT 79.34 3.655 79.63 3.885 ;
      RECT 79.34 3.69 80.115 3.86 ;
      RECT 79.4 2.175 79.57 3.885 ;
      RECT 79.34 2.175 79.635 2.405 ;
      RECT 78.97 4.025 79.26 4.255 ;
      RECT 78.97 4.055 79.43 4.225 ;
      RECT 79.035 2.95 79.2 4.255 ;
      RECT 77.55 2.915 77.84 3.145 ;
      RECT 77.55 2.95 79.2 3.12 ;
      RECT 77.61 2.175 77.78 3.145 ;
      RECT 77.55 2.175 77.84 2.405 ;
      RECT 77.55 10.055 77.84 10.285 ;
      RECT 77.61 9.315 77.78 10.285 ;
      RECT 77.61 9.405 79.2 9.575 ;
      RECT 79.03 8.205 79.2 9.575 ;
      RECT 77.55 9.315 77.84 9.545 ;
      RECT 78.97 8.205 79.26 8.435 ;
      RECT 78.97 8.235 79.43 8.405 ;
      RECT 77.98 3.26 78.33 3.61 ;
      RECT 75.645 3.32 78.33 3.49 ;
      RECT 77.81 3.315 78.33 3.49 ;
      RECT 75.645 2.635 75.815 3.49 ;
      RECT 75.545 2.635 75.895 2.985 ;
      RECT 78.005 8.94 78.33 9.265 ;
      RECT 73.38 8.895 73.73 9.245 ;
      RECT 77.98 8.945 78.33 9.175 ;
      RECT 73.2 8.945 73.73 9.175 ;
      RECT 77.81 8.97 78.33 9.145 ;
      RECT 73.03 8.975 73.73 9.145 ;
      RECT 73.2 8.97 78.33 9.14 ;
      RECT 77.205 3.66 77.525 3.98 ;
      RECT 77.18 3.655 77.47 3.885 ;
      RECT 77.105 3.685 77.525 3.86 ;
      RECT 77.005 3.685 77.525 3.855 ;
      RECT 77.205 8.54 77.525 8.83 ;
      RECT 77.18 8.575 77.525 8.805 ;
      RECT 77.005 8.605 77.525 8.775 ;
      RECT 73.84 3.76 74.025 3.97 ;
      RECT 73.83 3.765 74.04 3.963 ;
      RECT 73.83 3.765 74.126 3.94 ;
      RECT 73.83 3.765 74.185 3.915 ;
      RECT 73.83 3.765 74.24 3.895 ;
      RECT 73.83 3.765 74.25 3.883 ;
      RECT 73.83 3.765 74.445 3.822 ;
      RECT 73.83 3.765 74.475 3.805 ;
      RECT 73.83 3.765 74.495 3.795 ;
      RECT 74.375 3.53 74.635 3.79 ;
      RECT 74.36 3.62 74.375 3.837 ;
      RECT 73.895 3.752 74.635 3.79 ;
      RECT 74.346 3.631 74.36 3.843 ;
      RECT 73.935 3.745 74.635 3.79 ;
      RECT 74.26 3.671 74.346 3.862 ;
      RECT 74.185 3.732 74.635 3.79 ;
      RECT 74.255 3.707 74.26 3.879 ;
      RECT 74.24 3.717 74.635 3.79 ;
      RECT 74.25 3.712 74.255 3.881 ;
      RECT 73.175 3.795 73.28 4.055 ;
      RECT 73.99 3.32 73.995 3.545 ;
      RECT 74.12 3.32 74.175 3.53 ;
      RECT 74.175 3.325 74.185 3.523 ;
      RECT 74.081 3.32 74.12 3.533 ;
      RECT 73.995 3.32 74.081 3.54 ;
      RECT 73.975 3.325 73.99 3.546 ;
      RECT 73.965 3.365 73.975 3.548 ;
      RECT 73.935 3.375 73.965 3.55 ;
      RECT 73.93 3.38 73.935 3.552 ;
      RECT 73.905 3.385 73.93 3.554 ;
      RECT 73.89 3.39 73.905 3.556 ;
      RECT 73.875 3.392 73.89 3.558 ;
      RECT 73.87 3.397 73.875 3.56 ;
      RECT 73.82 3.405 73.87 3.563 ;
      RECT 73.795 3.414 73.82 3.568 ;
      RECT 73.785 3.421 73.795 3.573 ;
      RECT 73.78 3.424 73.785 3.577 ;
      RECT 73.76 3.427 73.78 3.586 ;
      RECT 73.73 3.435 73.76 3.606 ;
      RECT 73.701 3.448 73.73 3.628 ;
      RECT 73.615 3.482 73.701 3.672 ;
      RECT 73.61 3.508 73.615 3.71 ;
      RECT 73.605 3.512 73.61 3.719 ;
      RECT 73.57 3.525 73.605 3.752 ;
      RECT 73.56 3.539 73.57 3.79 ;
      RECT 73.555 3.543 73.56 3.803 ;
      RECT 73.55 3.547 73.555 3.808 ;
      RECT 73.54 3.555 73.55 3.82 ;
      RECT 73.535 3.562 73.54 3.835 ;
      RECT 73.51 3.575 73.535 3.86 ;
      RECT 73.47 3.604 73.51 3.915 ;
      RECT 73.455 3.629 73.47 3.97 ;
      RECT 73.445 3.64 73.455 3.993 ;
      RECT 73.44 3.647 73.445 4.005 ;
      RECT 73.435 3.651 73.44 4.013 ;
      RECT 73.38 3.679 73.435 4.055 ;
      RECT 73.36 3.715 73.38 4.055 ;
      RECT 73.345 3.73 73.36 4.055 ;
      RECT 73.29 3.762 73.345 4.055 ;
      RECT 73.28 3.792 73.29 4.055 ;
      RECT 72.89 3.407 73.075 3.645 ;
      RECT 72.875 3.409 73.085 3.64 ;
      RECT 72.76 3.355 73.02 3.615 ;
      RECT 72.755 3.392 73.02 3.569 ;
      RECT 72.75 3.402 73.02 3.566 ;
      RECT 72.745 3.442 73.085 3.56 ;
      RECT 72.74 3.475 73.085 3.55 ;
      RECT 72.75 3.417 73.1 3.488 ;
      RECT 73.047 4.515 73.06 5.045 ;
      RECT 72.961 4.515 73.06 5.044 ;
      RECT 72.961 4.515 73.065 5.043 ;
      RECT 72.875 4.515 73.065 5.041 ;
      RECT 72.87 4.515 73.065 5.038 ;
      RECT 72.87 4.515 73.075 5.036 ;
      RECT 72.865 4.807 73.075 5.033 ;
      RECT 72.865 4.817 73.08 5.03 ;
      RECT 72.865 4.885 73.085 5.026 ;
      RECT 72.855 4.89 73.085 5.025 ;
      RECT 72.855 4.982 73.09 5.022 ;
      RECT 72.84 4.515 73.1 4.775 ;
      RECT 72.77 10.055 73.06 10.285 ;
      RECT 72.83 9.315 73 10.285 ;
      RECT 72.745 9.34 73.085 9.685 ;
      RECT 72.77 9.315 73.06 9.685 ;
      RECT 72.07 3.505 72.115 5.04 ;
      RECT 72.27 3.505 72.3 3.72 ;
      RECT 70.645 3.245 70.765 3.455 ;
      RECT 70.305 3.195 70.565 3.455 ;
      RECT 70.305 3.24 70.6 3.445 ;
      RECT 72.31 3.521 72.315 3.575 ;
      RECT 72.305 3.514 72.31 3.708 ;
      RECT 72.3 3.508 72.305 3.715 ;
      RECT 72.255 3.505 72.27 3.728 ;
      RECT 72.25 3.505 72.255 3.75 ;
      RECT 72.245 3.505 72.25 3.798 ;
      RECT 72.24 3.505 72.245 3.818 ;
      RECT 72.23 3.505 72.24 3.925 ;
      RECT 72.225 3.505 72.23 3.988 ;
      RECT 72.22 3.505 72.225 4.045 ;
      RECT 72.215 3.505 72.22 4.053 ;
      RECT 72.2 3.505 72.215 4.16 ;
      RECT 72.19 3.505 72.2 4.295 ;
      RECT 72.18 3.505 72.19 4.405 ;
      RECT 72.17 3.505 72.18 4.462 ;
      RECT 72.165 3.505 72.17 4.502 ;
      RECT 72.16 3.505 72.165 4.538 ;
      RECT 72.15 3.505 72.16 4.578 ;
      RECT 72.145 3.505 72.15 4.62 ;
      RECT 72.125 3.505 72.145 4.685 ;
      RECT 72.13 4.83 72.135 5.01 ;
      RECT 72.125 4.812 72.13 5.018 ;
      RECT 72.12 3.505 72.125 4.748 ;
      RECT 72.12 4.792 72.125 5.025 ;
      RECT 72.115 3.505 72.12 5.035 ;
      RECT 72.06 3.505 72.07 3.805 ;
      RECT 72.065 4.052 72.07 5.04 ;
      RECT 72.06 4.117 72.065 5.04 ;
      RECT 72.055 3.506 72.06 3.795 ;
      RECT 72.05 4.182 72.06 5.04 ;
      RECT 72.045 3.507 72.055 3.785 ;
      RECT 72.035 4.295 72.05 5.04 ;
      RECT 72.04 3.508 72.045 3.775 ;
      RECT 72.02 3.509 72.04 3.753 ;
      RECT 72.025 4.392 72.035 5.04 ;
      RECT 72.02 4.467 72.025 5.04 ;
      RECT 72.01 3.508 72.02 3.73 ;
      RECT 72.015 4.51 72.02 5.04 ;
      RECT 72.01 4.537 72.015 5.04 ;
      RECT 72 3.506 72.01 3.718 ;
      RECT 72.005 4.58 72.01 5.04 ;
      RECT 72 4.607 72.005 5.04 ;
      RECT 71.99 3.505 72 3.705 ;
      RECT 71.995 4.622 72 5.04 ;
      RECT 71.955 4.68 71.995 5.04 ;
      RECT 71.985 3.504 71.99 3.69 ;
      RECT 71.98 3.502 71.985 3.683 ;
      RECT 71.97 3.499 71.98 3.673 ;
      RECT 71.965 3.496 71.97 3.658 ;
      RECT 71.95 3.492 71.965 3.651 ;
      RECT 71.945 4.735 71.955 5.04 ;
      RECT 71.945 3.489 71.95 3.646 ;
      RECT 71.93 3.485 71.945 3.64 ;
      RECT 71.94 4.752 71.945 5.04 ;
      RECT 71.93 4.815 71.94 5.04 ;
      RECT 71.85 3.47 71.93 3.62 ;
      RECT 71.925 4.822 71.93 5.035 ;
      RECT 71.92 4.83 71.925 5.025 ;
      RECT 71.84 3.456 71.85 3.604 ;
      RECT 71.825 3.452 71.84 3.602 ;
      RECT 71.815 3.447 71.825 3.598 ;
      RECT 71.79 3.44 71.815 3.59 ;
      RECT 71.785 3.435 71.79 3.585 ;
      RECT 71.775 3.435 71.785 3.583 ;
      RECT 71.765 3.433 71.775 3.581 ;
      RECT 71.735 3.425 71.765 3.575 ;
      RECT 71.72 3.417 71.735 3.568 ;
      RECT 71.7 3.412 71.72 3.561 ;
      RECT 71.695 3.408 71.7 3.556 ;
      RECT 71.665 3.401 71.695 3.55 ;
      RECT 71.64 3.392 71.665 3.54 ;
      RECT 71.61 3.385 71.64 3.532 ;
      RECT 71.585 3.375 71.61 3.523 ;
      RECT 71.57 3.367 71.585 3.517 ;
      RECT 71.545 3.362 71.57 3.512 ;
      RECT 71.535 3.358 71.545 3.507 ;
      RECT 71.515 3.353 71.535 3.502 ;
      RECT 71.48 3.348 71.515 3.495 ;
      RECT 71.42 3.343 71.48 3.488 ;
      RECT 71.407 3.339 71.42 3.486 ;
      RECT 71.321 3.334 71.407 3.483 ;
      RECT 71.235 3.324 71.321 3.479 ;
      RECT 71.194 3.317 71.235 3.476 ;
      RECT 71.108 3.31 71.194 3.473 ;
      RECT 71.022 3.3 71.108 3.469 ;
      RECT 70.936 3.29 71.022 3.464 ;
      RECT 70.85 3.28 70.936 3.46 ;
      RECT 70.84 3.265 70.85 3.458 ;
      RECT 70.83 3.25 70.84 3.458 ;
      RECT 70.765 3.245 70.83 3.457 ;
      RECT 70.6 3.242 70.645 3.45 ;
      RECT 71.845 4.147 71.85 4.338 ;
      RECT 71.84 4.142 71.845 4.345 ;
      RECT 71.826 4.14 71.84 4.351 ;
      RECT 71.74 4.14 71.826 4.353 ;
      RECT 71.736 4.14 71.74 4.356 ;
      RECT 71.65 4.14 71.736 4.374 ;
      RECT 71.64 4.145 71.65 4.393 ;
      RECT 71.63 4.2 71.64 4.397 ;
      RECT 71.605 4.215 71.63 4.404 ;
      RECT 71.565 4.235 71.605 4.417 ;
      RECT 71.56 4.247 71.565 4.427 ;
      RECT 71.545 4.253 71.56 4.432 ;
      RECT 71.54 4.258 71.545 4.436 ;
      RECT 71.52 4.265 71.54 4.441 ;
      RECT 71.45 4.29 71.52 4.458 ;
      RECT 71.41 4.318 71.45 4.478 ;
      RECT 71.405 4.328 71.41 4.486 ;
      RECT 71.385 4.335 71.405 4.488 ;
      RECT 71.38 4.342 71.385 4.491 ;
      RECT 71.35 4.35 71.38 4.494 ;
      RECT 71.345 4.355 71.35 4.498 ;
      RECT 71.271 4.359 71.345 4.506 ;
      RECT 71.185 4.368 71.271 4.522 ;
      RECT 71.181 4.373 71.185 4.531 ;
      RECT 71.095 4.378 71.181 4.541 ;
      RECT 71.055 4.386 71.095 4.553 ;
      RECT 71.005 4.392 71.055 4.56 ;
      RECT 70.92 4.401 71.005 4.575 ;
      RECT 70.845 4.412 70.92 4.593 ;
      RECT 70.81 4.419 70.845 4.603 ;
      RECT 70.735 4.427 70.81 4.608 ;
      RECT 70.68 4.436 70.735 4.608 ;
      RECT 70.655 4.441 70.68 4.606 ;
      RECT 70.645 4.444 70.655 4.604 ;
      RECT 70.61 4.446 70.645 4.602 ;
      RECT 70.58 4.448 70.61 4.598 ;
      RECT 70.535 4.447 70.58 4.594 ;
      RECT 70.515 4.442 70.535 4.591 ;
      RECT 70.465 4.427 70.515 4.588 ;
      RECT 70.455 4.412 70.465 4.583 ;
      RECT 70.405 4.397 70.455 4.573 ;
      RECT 70.355 4.372 70.405 4.553 ;
      RECT 70.345 4.357 70.355 4.535 ;
      RECT 70.34 4.355 70.345 4.529 ;
      RECT 70.32 4.35 70.34 4.524 ;
      RECT 70.315 4.342 70.32 4.518 ;
      RECT 70.3 4.336 70.315 4.511 ;
      RECT 70.295 4.331 70.3 4.503 ;
      RECT 70.275 4.326 70.295 4.495 ;
      RECT 70.26 4.319 70.275 4.488 ;
      RECT 70.245 4.313 70.26 4.479 ;
      RECT 70.24 4.307 70.245 4.472 ;
      RECT 70.195 4.282 70.24 4.458 ;
      RECT 70.18 4.252 70.195 4.44 ;
      RECT 70.165 4.235 70.18 4.431 ;
      RECT 70.14 4.215 70.165 4.419 ;
      RECT 70.1 4.185 70.14 4.399 ;
      RECT 70.09 4.155 70.1 4.384 ;
      RECT 70.075 4.145 70.09 4.377 ;
      RECT 70.02 4.11 70.075 4.356 ;
      RECT 70.005 4.073 70.02 4.335 ;
      RECT 69.995 4.06 70.005 4.327 ;
      RECT 69.945 4.03 69.995 4.309 ;
      RECT 69.93 3.96 69.945 4.29 ;
      RECT 69.885 3.96 69.93 4.273 ;
      RECT 69.86 3.96 69.885 4.255 ;
      RECT 69.85 3.96 69.86 4.248 ;
      RECT 69.771 3.96 69.85 4.241 ;
      RECT 69.685 3.96 69.771 4.233 ;
      RECT 69.67 3.992 69.685 4.228 ;
      RECT 69.595 4.002 69.67 4.224 ;
      RECT 69.575 4.012 69.595 4.219 ;
      RECT 69.55 4.012 69.575 4.216 ;
      RECT 69.54 4.002 69.55 4.215 ;
      RECT 69.53 3.975 69.54 4.214 ;
      RECT 69.49 3.97 69.53 4.212 ;
      RECT 69.445 3.97 69.49 4.208 ;
      RECT 69.42 3.97 69.445 4.203 ;
      RECT 69.37 3.97 69.42 4.19 ;
      RECT 69.33 3.975 69.34 4.175 ;
      RECT 69.34 3.97 69.37 4.18 ;
      RECT 71.325 3.75 71.585 4.01 ;
      RECT 71.32 3.772 71.585 3.968 ;
      RECT 70.56 3.6 70.78 3.965 ;
      RECT 70.542 3.687 70.78 3.964 ;
      RECT 70.525 3.692 70.78 3.961 ;
      RECT 70.525 3.692 70.8 3.96 ;
      RECT 70.495 3.702 70.8 3.958 ;
      RECT 70.49 3.717 70.8 3.954 ;
      RECT 70.49 3.717 70.805 3.953 ;
      RECT 70.485 3.775 70.805 3.951 ;
      RECT 70.485 3.775 70.815 3.948 ;
      RECT 70.48 3.84 70.815 3.943 ;
      RECT 70.56 3.6 70.82 3.86 ;
      RECT 69.305 3.43 69.565 3.69 ;
      RECT 69.305 3.473 69.651 3.664 ;
      RECT 69.305 3.473 69.695 3.663 ;
      RECT 69.305 3.473 69.715 3.661 ;
      RECT 69.305 3.473 69.815 3.66 ;
      RECT 69.305 3.473 69.835 3.658 ;
      RECT 69.305 3.473 69.845 3.653 ;
      RECT 69.715 3.44 69.905 3.65 ;
      RECT 69.715 3.442 69.91 3.648 ;
      RECT 69.705 3.447 69.915 3.64 ;
      RECT 69.651 3.471 69.915 3.64 ;
      RECT 69.695 3.465 69.705 3.662 ;
      RECT 69.705 3.445 69.91 3.648 ;
      RECT 68.66 4.505 68.865 4.735 ;
      RECT 68.6 4.455 68.655 4.715 ;
      RECT 68.66 4.455 68.86 4.735 ;
      RECT 69.63 4.77 69.635 4.797 ;
      RECT 69.62 4.68 69.63 4.802 ;
      RECT 69.615 4.602 69.62 4.808 ;
      RECT 69.605 4.592 69.615 4.815 ;
      RECT 69.6 4.582 69.605 4.821 ;
      RECT 69.59 4.577 69.6 4.823 ;
      RECT 69.575 4.569 69.59 4.831 ;
      RECT 69.56 4.56 69.575 4.843 ;
      RECT 69.55 4.552 69.56 4.853 ;
      RECT 69.515 4.47 69.55 4.871 ;
      RECT 69.48 4.47 69.515 4.89 ;
      RECT 69.465 4.47 69.48 4.898 ;
      RECT 69.41 4.47 69.465 4.898 ;
      RECT 69.376 4.47 69.41 4.889 ;
      RECT 69.29 4.47 69.376 4.865 ;
      RECT 69.28 4.53 69.29 4.847 ;
      RECT 69.24 4.532 69.28 4.838 ;
      RECT 69.235 4.534 69.24 4.828 ;
      RECT 69.215 4.536 69.235 4.823 ;
      RECT 69.205 4.539 69.215 4.818 ;
      RECT 69.195 4.54 69.205 4.813 ;
      RECT 69.171 4.541 69.195 4.805 ;
      RECT 69.085 4.546 69.171 4.783 ;
      RECT 69.03 4.545 69.085 4.756 ;
      RECT 69.015 4.538 69.03 4.743 ;
      RECT 68.98 4.533 69.015 4.739 ;
      RECT 68.925 4.525 68.98 4.738 ;
      RECT 68.865 4.512 68.925 4.736 ;
      RECT 68.655 4.455 68.66 4.723 ;
      RECT 68.73 3.825 68.915 4.035 ;
      RECT 68.72 3.83 68.93 4.028 ;
      RECT 68.76 3.735 69.02 3.995 ;
      RECT 68.715 3.892 69.02 3.918 ;
      RECT 68.06 3.685 68.065 4.485 ;
      RECT 68.005 3.735 68.035 4.485 ;
      RECT 67.995 3.735 68 4.045 ;
      RECT 67.98 3.735 67.985 4.04 ;
      RECT 67.525 3.78 67.54 3.995 ;
      RECT 67.455 3.78 67.54 3.99 ;
      RECT 68.72 3.36 68.79 3.57 ;
      RECT 68.79 3.367 68.8 3.565 ;
      RECT 68.686 3.36 68.72 3.577 ;
      RECT 68.6 3.36 68.686 3.601 ;
      RECT 68.59 3.365 68.6 3.62 ;
      RECT 68.585 3.377 68.59 3.623 ;
      RECT 68.57 3.392 68.585 3.627 ;
      RECT 68.565 3.41 68.57 3.631 ;
      RECT 68.525 3.42 68.565 3.64 ;
      RECT 68.51 3.427 68.525 3.652 ;
      RECT 68.495 3.432 68.51 3.657 ;
      RECT 68.48 3.435 68.495 3.662 ;
      RECT 68.47 3.437 68.48 3.666 ;
      RECT 68.435 3.444 68.47 3.674 ;
      RECT 68.4 3.452 68.435 3.688 ;
      RECT 68.39 3.458 68.4 3.697 ;
      RECT 68.385 3.46 68.39 3.699 ;
      RECT 68.365 3.463 68.385 3.705 ;
      RECT 68.335 3.47 68.365 3.716 ;
      RECT 68.325 3.476 68.335 3.723 ;
      RECT 68.3 3.479 68.325 3.73 ;
      RECT 68.29 3.483 68.3 3.738 ;
      RECT 68.285 3.484 68.29 3.76 ;
      RECT 68.28 3.485 68.285 3.775 ;
      RECT 68.275 3.486 68.28 3.79 ;
      RECT 68.27 3.487 68.275 3.805 ;
      RECT 68.265 3.488 68.27 3.835 ;
      RECT 68.255 3.49 68.265 3.868 ;
      RECT 68.24 3.494 68.255 3.915 ;
      RECT 68.23 3.497 68.24 3.96 ;
      RECT 68.225 3.5 68.23 3.988 ;
      RECT 68.215 3.502 68.225 4.015 ;
      RECT 68.21 3.505 68.215 4.05 ;
      RECT 68.18 3.51 68.21 4.108 ;
      RECT 68.175 3.515 68.18 4.193 ;
      RECT 68.17 3.517 68.175 4.228 ;
      RECT 68.165 3.519 68.17 4.31 ;
      RECT 68.16 3.521 68.165 4.398 ;
      RECT 68.15 3.523 68.16 4.48 ;
      RECT 68.135 3.537 68.15 4.485 ;
      RECT 68.1 3.582 68.135 4.485 ;
      RECT 68.09 3.622 68.1 4.485 ;
      RECT 68.075 3.65 68.09 4.485 ;
      RECT 68.07 3.667 68.075 4.485 ;
      RECT 68.065 3.675 68.07 4.485 ;
      RECT 68.055 3.69 68.06 4.485 ;
      RECT 68.05 3.697 68.055 4.485 ;
      RECT 68.04 3.717 68.05 4.485 ;
      RECT 68.035 3.73 68.04 4.485 ;
      RECT 68 3.735 68.005 4.07 ;
      RECT 67.985 4.125 68.005 4.485 ;
      RECT 67.985 3.735 67.995 4.043 ;
      RECT 67.98 4.165 67.985 4.485 ;
      RECT 67.93 3.735 67.98 4.038 ;
      RECT 67.975 4.202 67.98 4.485 ;
      RECT 67.965 4.225 67.975 4.485 ;
      RECT 67.96 4.27 67.965 4.485 ;
      RECT 67.95 4.28 67.96 4.478 ;
      RECT 67.876 3.735 67.93 4.032 ;
      RECT 67.79 3.735 67.876 4.025 ;
      RECT 67.741 3.782 67.79 4.018 ;
      RECT 67.655 3.79 67.741 4.011 ;
      RECT 67.64 3.787 67.655 4.006 ;
      RECT 67.626 3.78 67.64 4.005 ;
      RECT 67.54 3.78 67.626 4 ;
      RECT 67.445 3.785 67.455 3.985 ;
      RECT 67.035 3.215 67.05 3.615 ;
      RECT 67.23 3.215 67.235 3.475 ;
      RECT 66.975 3.215 67.02 3.475 ;
      RECT 67.43 4.52 67.435 4.725 ;
      RECT 67.425 4.51 67.43 4.73 ;
      RECT 67.42 4.497 67.425 4.735 ;
      RECT 67.415 4.477 67.42 4.735 ;
      RECT 67.39 4.43 67.415 4.735 ;
      RECT 67.355 4.345 67.39 4.735 ;
      RECT 67.35 4.282 67.355 4.735 ;
      RECT 67.345 4.267 67.35 4.735 ;
      RECT 67.33 4.227 67.345 4.735 ;
      RECT 67.325 4.202 67.33 4.735 ;
      RECT 67.315 4.185 67.325 4.735 ;
      RECT 67.28 4.107 67.315 4.735 ;
      RECT 67.275 4.05 67.28 4.735 ;
      RECT 67.27 4.037 67.275 4.735 ;
      RECT 67.26 4.015 67.27 4.735 ;
      RECT 67.25 3.98 67.26 4.735 ;
      RECT 67.24 3.95 67.25 4.735 ;
      RECT 67.23 3.865 67.24 4.378 ;
      RECT 67.237 4.51 67.24 4.735 ;
      RECT 67.235 4.52 67.237 4.735 ;
      RECT 67.225 4.53 67.235 4.73 ;
      RECT 67.22 3.215 67.23 3.61 ;
      RECT 67.225 3.742 67.23 4.353 ;
      RECT 67.22 3.64 67.225 4.336 ;
      RECT 67.21 3.215 67.22 4.312 ;
      RECT 67.205 3.215 67.21 4.283 ;
      RECT 67.2 3.215 67.205 4.273 ;
      RECT 67.18 3.215 67.2 4.235 ;
      RECT 67.175 3.215 67.18 4.193 ;
      RECT 67.17 3.215 67.175 4.173 ;
      RECT 67.14 3.215 67.17 4.123 ;
      RECT 67.13 3.215 67.14 4.07 ;
      RECT 67.125 3.215 67.13 4.043 ;
      RECT 67.12 3.215 67.125 4.028 ;
      RECT 67.11 3.215 67.12 4.005 ;
      RECT 67.1 3.215 67.11 3.98 ;
      RECT 67.095 3.215 67.1 3.92 ;
      RECT 67.085 3.215 67.095 3.858 ;
      RECT 67.08 3.215 67.085 3.778 ;
      RECT 67.075 3.215 67.08 3.743 ;
      RECT 67.07 3.215 67.075 3.718 ;
      RECT 67.065 3.215 67.07 3.703 ;
      RECT 67.06 3.215 67.065 3.673 ;
      RECT 67.055 3.215 67.06 3.65 ;
      RECT 67.05 3.215 67.055 3.623 ;
      RECT 67.02 3.215 67.035 3.61 ;
      RECT 66.175 4.75 66.36 4.96 ;
      RECT 66.165 4.755 66.375 4.953 ;
      RECT 66.165 4.755 66.395 4.925 ;
      RECT 66.165 4.755 66.41 4.904 ;
      RECT 66.165 4.755 66.425 4.902 ;
      RECT 66.165 4.755 66.435 4.901 ;
      RECT 66.165 4.755 66.465 4.898 ;
      RECT 66.815 4.6 67.075 4.86 ;
      RECT 66.775 4.647 67.075 4.843 ;
      RECT 66.766 4.655 66.775 4.846 ;
      RECT 66.36 4.748 67.075 4.843 ;
      RECT 66.68 4.673 66.766 4.853 ;
      RECT 66.375 4.745 67.075 4.843 ;
      RECT 66.621 4.695 66.68 4.865 ;
      RECT 66.395 4.741 67.075 4.843 ;
      RECT 66.535 4.707 66.621 4.876 ;
      RECT 66.41 4.737 67.075 4.843 ;
      RECT 66.48 4.72 66.535 4.888 ;
      RECT 66.425 4.735 67.075 4.843 ;
      RECT 66.465 4.726 66.48 4.894 ;
      RECT 66.435 4.731 67.075 4.843 ;
      RECT 66.58 4.255 66.84 4.515 ;
      RECT 66.58 4.275 66.95 4.485 ;
      RECT 66.58 4.28 66.96 4.48 ;
      RECT 66.771 3.694 66.85 3.925 ;
      RECT 66.685 3.697 66.9 3.92 ;
      RECT 66.68 3.697 66.9 3.915 ;
      RECT 66.68 3.702 66.91 3.913 ;
      RECT 66.655 3.702 66.91 3.91 ;
      RECT 66.655 3.71 66.92 3.908 ;
      RECT 66.535 3.645 66.795 3.905 ;
      RECT 66.535 3.692 66.845 3.905 ;
      RECT 65.79 4.265 65.795 4.525 ;
      RECT 65.62 4.035 65.625 4.525 ;
      RECT 65.505 4.275 65.51 4.5 ;
      RECT 66.215 3.37 66.22 3.58 ;
      RECT 66.22 3.375 66.235 3.575 ;
      RECT 66.155 3.37 66.215 3.588 ;
      RECT 66.14 3.37 66.155 3.598 ;
      RECT 66.09 3.37 66.14 3.615 ;
      RECT 66.07 3.37 66.09 3.638 ;
      RECT 66.055 3.37 66.07 3.65 ;
      RECT 66.035 3.37 66.055 3.66 ;
      RECT 66.025 3.375 66.035 3.669 ;
      RECT 66.02 3.385 66.025 3.674 ;
      RECT 66.015 3.397 66.02 3.678 ;
      RECT 66.005 3.42 66.015 3.683 ;
      RECT 66 3.435 66.005 3.687 ;
      RECT 65.995 3.452 66 3.69 ;
      RECT 65.99 3.46 65.995 3.693 ;
      RECT 65.98 3.465 65.99 3.697 ;
      RECT 65.975 3.472 65.98 3.702 ;
      RECT 65.965 3.477 65.975 3.706 ;
      RECT 65.94 3.489 65.965 3.717 ;
      RECT 65.92 3.506 65.94 3.733 ;
      RECT 65.895 3.523 65.92 3.755 ;
      RECT 65.86 3.546 65.895 3.813 ;
      RECT 65.84 3.568 65.86 3.875 ;
      RECT 65.835 3.578 65.84 3.91 ;
      RECT 65.825 3.585 65.835 3.948 ;
      RECT 65.82 3.592 65.825 3.968 ;
      RECT 65.815 3.603 65.82 4.005 ;
      RECT 65.81 3.611 65.815 4.07 ;
      RECT 65.8 3.622 65.81 4.123 ;
      RECT 65.795 3.64 65.8 4.193 ;
      RECT 65.79 3.65 65.795 4.23 ;
      RECT 65.785 3.66 65.79 4.525 ;
      RECT 65.78 3.672 65.785 4.525 ;
      RECT 65.775 3.682 65.78 4.525 ;
      RECT 65.765 3.692 65.775 4.525 ;
      RECT 65.755 3.715 65.765 4.525 ;
      RECT 65.74 3.75 65.755 4.525 ;
      RECT 65.7 3.812 65.74 4.525 ;
      RECT 65.695 3.865 65.7 4.525 ;
      RECT 65.67 3.9 65.695 4.525 ;
      RECT 65.655 3.945 65.67 4.525 ;
      RECT 65.65 3.967 65.655 4.525 ;
      RECT 65.64 3.98 65.65 4.525 ;
      RECT 65.63 4.005 65.64 4.525 ;
      RECT 65.625 4.027 65.63 4.525 ;
      RECT 65.6 4.065 65.62 4.525 ;
      RECT 65.56 4.122 65.6 4.525 ;
      RECT 65.555 4.172 65.56 4.525 ;
      RECT 65.55 4.19 65.555 4.525 ;
      RECT 65.545 4.202 65.55 4.525 ;
      RECT 65.535 4.22 65.545 4.525 ;
      RECT 65.525 4.24 65.535 4.5 ;
      RECT 65.52 4.257 65.525 4.5 ;
      RECT 65.51 4.27 65.52 4.5 ;
      RECT 65.48 4.28 65.505 4.5 ;
      RECT 65.47 4.287 65.48 4.5 ;
      RECT 65.455 4.297 65.47 4.495 ;
      RECT 64.55 10.05 64.845 10.28 ;
      RECT 64.61 8.57 64.78 10.28 ;
      RECT 64.555 8.94 64.905 9.29 ;
      RECT 64.55 8.57 64.84 8.8 ;
      RECT 64.57 7.215 64.85 7.585 ;
      RECT 64.525 7.215 64.875 7.565 ;
      RECT 63.555 10.055 63.85 10.285 ;
      RECT 63.615 8.575 63.785 10.285 ;
      RECT 63.555 8.575 63.845 8.805 ;
      RECT 63.555 8.61 64.41 8.77 ;
      RECT 64.24 8.2 64.41 8.77 ;
      RECT 63.555 8.605 63.95 8.77 ;
      RECT 64.18 8.2 64.47 8.43 ;
      RECT 64.18 8.23 64.64 8.4 ;
      RECT 64.14 4.03 64.465 4.26 ;
      RECT 64.14 4.06 64.635 4.23 ;
      RECT 64.14 3.69 64.33 4.26 ;
      RECT 63.555 3.655 63.845 3.885 ;
      RECT 63.555 3.69 64.33 3.86 ;
      RECT 63.615 2.175 63.785 3.885 ;
      RECT 63.555 2.175 63.85 2.405 ;
      RECT 63.185 4.025 63.475 4.255 ;
      RECT 63.185 4.055 63.645 4.225 ;
      RECT 63.25 2.95 63.415 4.255 ;
      RECT 61.765 2.915 62.055 3.145 ;
      RECT 61.765 2.95 63.415 3.12 ;
      RECT 61.825 2.175 61.995 3.145 ;
      RECT 61.765 2.175 62.055 2.405 ;
      RECT 61.765 10.055 62.055 10.285 ;
      RECT 61.825 9.315 61.995 10.285 ;
      RECT 61.825 9.405 63.415 9.575 ;
      RECT 63.245 8.205 63.415 9.575 ;
      RECT 61.765 9.315 62.055 9.545 ;
      RECT 63.185 8.205 63.475 8.435 ;
      RECT 63.185 8.235 63.645 8.405 ;
      RECT 62.195 3.26 62.545 3.61 ;
      RECT 59.86 3.32 62.545 3.49 ;
      RECT 62.025 3.315 62.545 3.49 ;
      RECT 59.86 2.635 60.03 3.49 ;
      RECT 59.76 2.635 60.11 2.985 ;
      RECT 62.22 8.94 62.545 9.265 ;
      RECT 57.65 8.9 58 9.25 ;
      RECT 62.195 8.945 62.545 9.175 ;
      RECT 57.415 8.945 58 9.175 ;
      RECT 62.025 8.97 62.545 9.145 ;
      RECT 57.245 8.975 58 9.145 ;
      RECT 57.415 8.97 62.545 9.14 ;
      RECT 61.42 3.66 61.74 3.98 ;
      RECT 61.395 3.655 61.685 3.885 ;
      RECT 61.32 3.685 61.74 3.86 ;
      RECT 61.22 3.685 61.74 3.855 ;
      RECT 61.42 8.54 61.74 8.83 ;
      RECT 61.395 8.575 61.74 8.805 ;
      RECT 61.22 8.605 61.74 8.775 ;
      RECT 58.055 3.76 58.24 3.97 ;
      RECT 58.045 3.765 58.255 3.963 ;
      RECT 58.045 3.765 58.341 3.94 ;
      RECT 58.045 3.765 58.4 3.915 ;
      RECT 58.045 3.765 58.455 3.895 ;
      RECT 58.045 3.765 58.465 3.883 ;
      RECT 58.045 3.765 58.66 3.822 ;
      RECT 58.045 3.765 58.69 3.805 ;
      RECT 58.045 3.765 58.71 3.795 ;
      RECT 58.59 3.53 58.85 3.79 ;
      RECT 58.575 3.62 58.59 3.837 ;
      RECT 58.11 3.752 58.85 3.79 ;
      RECT 58.561 3.631 58.575 3.843 ;
      RECT 58.15 3.745 58.85 3.79 ;
      RECT 58.475 3.671 58.561 3.862 ;
      RECT 58.4 3.732 58.85 3.79 ;
      RECT 58.47 3.707 58.475 3.879 ;
      RECT 58.455 3.717 58.85 3.79 ;
      RECT 58.465 3.712 58.47 3.881 ;
      RECT 57.39 3.795 57.495 4.055 ;
      RECT 58.205 3.32 58.21 3.545 ;
      RECT 58.335 3.32 58.39 3.53 ;
      RECT 58.39 3.325 58.4 3.523 ;
      RECT 58.296 3.32 58.335 3.533 ;
      RECT 58.21 3.32 58.296 3.54 ;
      RECT 58.19 3.325 58.205 3.546 ;
      RECT 58.18 3.365 58.19 3.548 ;
      RECT 58.15 3.375 58.18 3.55 ;
      RECT 58.145 3.38 58.15 3.552 ;
      RECT 58.12 3.385 58.145 3.554 ;
      RECT 58.105 3.39 58.12 3.556 ;
      RECT 58.09 3.392 58.105 3.558 ;
      RECT 58.085 3.397 58.09 3.56 ;
      RECT 58.035 3.405 58.085 3.563 ;
      RECT 58.01 3.414 58.035 3.568 ;
      RECT 58 3.421 58.01 3.573 ;
      RECT 57.995 3.424 58 3.577 ;
      RECT 57.975 3.427 57.995 3.586 ;
      RECT 57.945 3.435 57.975 3.606 ;
      RECT 57.916 3.448 57.945 3.628 ;
      RECT 57.83 3.482 57.916 3.672 ;
      RECT 57.825 3.508 57.83 3.71 ;
      RECT 57.82 3.512 57.825 3.719 ;
      RECT 57.785 3.525 57.82 3.752 ;
      RECT 57.775 3.539 57.785 3.79 ;
      RECT 57.77 3.543 57.775 3.803 ;
      RECT 57.765 3.547 57.77 3.808 ;
      RECT 57.755 3.555 57.765 3.82 ;
      RECT 57.75 3.562 57.755 3.835 ;
      RECT 57.725 3.575 57.75 3.86 ;
      RECT 57.685 3.604 57.725 3.915 ;
      RECT 57.67 3.629 57.685 3.97 ;
      RECT 57.66 3.64 57.67 3.993 ;
      RECT 57.655 3.647 57.66 4.005 ;
      RECT 57.65 3.651 57.655 4.013 ;
      RECT 57.595 3.679 57.65 4.055 ;
      RECT 57.575 3.715 57.595 4.055 ;
      RECT 57.56 3.73 57.575 4.055 ;
      RECT 57.505 3.762 57.56 4.055 ;
      RECT 57.495 3.792 57.505 4.055 ;
      RECT 57.105 3.407 57.29 3.645 ;
      RECT 57.09 3.409 57.3 3.64 ;
      RECT 56.975 3.355 57.235 3.615 ;
      RECT 56.97 3.392 57.235 3.569 ;
      RECT 56.965 3.402 57.235 3.566 ;
      RECT 56.96 3.442 57.3 3.56 ;
      RECT 56.955 3.475 57.3 3.55 ;
      RECT 56.965 3.417 57.315 3.488 ;
      RECT 57.262 4.515 57.275 5.045 ;
      RECT 57.176 4.515 57.275 5.044 ;
      RECT 57.176 4.515 57.28 5.043 ;
      RECT 57.09 4.515 57.28 5.041 ;
      RECT 57.085 4.515 57.28 5.038 ;
      RECT 57.085 4.515 57.29 5.036 ;
      RECT 57.08 4.807 57.29 5.033 ;
      RECT 57.08 4.817 57.295 5.03 ;
      RECT 57.08 4.885 57.3 5.026 ;
      RECT 57.07 4.89 57.3 5.025 ;
      RECT 57.07 4.982 57.305 5.022 ;
      RECT 57.055 4.515 57.315 4.775 ;
      RECT 56.985 10.055 57.275 10.285 ;
      RECT 57.045 9.315 57.215 10.285 ;
      RECT 56.96 9.34 57.3 9.685 ;
      RECT 56.985 9.315 57.275 9.685 ;
      RECT 56.285 3.505 56.33 5.04 ;
      RECT 56.485 3.505 56.515 3.72 ;
      RECT 54.86 3.245 54.98 3.455 ;
      RECT 54.52 3.195 54.78 3.455 ;
      RECT 54.52 3.24 54.815 3.445 ;
      RECT 56.525 3.521 56.53 3.575 ;
      RECT 56.52 3.514 56.525 3.708 ;
      RECT 56.515 3.508 56.52 3.715 ;
      RECT 56.47 3.505 56.485 3.728 ;
      RECT 56.465 3.505 56.47 3.75 ;
      RECT 56.46 3.505 56.465 3.798 ;
      RECT 56.455 3.505 56.46 3.818 ;
      RECT 56.445 3.505 56.455 3.925 ;
      RECT 56.44 3.505 56.445 3.988 ;
      RECT 56.435 3.505 56.44 4.045 ;
      RECT 56.43 3.505 56.435 4.053 ;
      RECT 56.415 3.505 56.43 4.16 ;
      RECT 56.405 3.505 56.415 4.295 ;
      RECT 56.395 3.505 56.405 4.405 ;
      RECT 56.385 3.505 56.395 4.462 ;
      RECT 56.38 3.505 56.385 4.502 ;
      RECT 56.375 3.505 56.38 4.538 ;
      RECT 56.365 3.505 56.375 4.578 ;
      RECT 56.36 3.505 56.365 4.62 ;
      RECT 56.34 3.505 56.36 4.685 ;
      RECT 56.345 4.83 56.35 5.01 ;
      RECT 56.34 4.812 56.345 5.018 ;
      RECT 56.335 3.505 56.34 4.748 ;
      RECT 56.335 4.792 56.34 5.025 ;
      RECT 56.33 3.505 56.335 5.035 ;
      RECT 56.275 3.505 56.285 3.805 ;
      RECT 56.28 4.052 56.285 5.04 ;
      RECT 56.275 4.117 56.28 5.04 ;
      RECT 56.27 3.506 56.275 3.795 ;
      RECT 56.265 4.182 56.275 5.04 ;
      RECT 56.26 3.507 56.27 3.785 ;
      RECT 56.25 4.295 56.265 5.04 ;
      RECT 56.255 3.508 56.26 3.775 ;
      RECT 56.235 3.509 56.255 3.753 ;
      RECT 56.24 4.392 56.25 5.04 ;
      RECT 56.235 4.467 56.24 5.04 ;
      RECT 56.225 3.508 56.235 3.73 ;
      RECT 56.23 4.51 56.235 5.04 ;
      RECT 56.225 4.537 56.23 5.04 ;
      RECT 56.215 3.506 56.225 3.718 ;
      RECT 56.22 4.58 56.225 5.04 ;
      RECT 56.215 4.607 56.22 5.04 ;
      RECT 56.205 3.505 56.215 3.705 ;
      RECT 56.21 4.622 56.215 5.04 ;
      RECT 56.17 4.68 56.21 5.04 ;
      RECT 56.2 3.504 56.205 3.69 ;
      RECT 56.195 3.502 56.2 3.683 ;
      RECT 56.185 3.499 56.195 3.673 ;
      RECT 56.18 3.496 56.185 3.658 ;
      RECT 56.165 3.492 56.18 3.651 ;
      RECT 56.16 4.735 56.17 5.04 ;
      RECT 56.16 3.489 56.165 3.646 ;
      RECT 56.145 3.485 56.16 3.64 ;
      RECT 56.155 4.752 56.16 5.04 ;
      RECT 56.145 4.815 56.155 5.04 ;
      RECT 56.065 3.47 56.145 3.62 ;
      RECT 56.14 4.822 56.145 5.035 ;
      RECT 56.135 4.83 56.14 5.025 ;
      RECT 56.055 3.456 56.065 3.604 ;
      RECT 56.04 3.452 56.055 3.602 ;
      RECT 56.03 3.447 56.04 3.598 ;
      RECT 56.005 3.44 56.03 3.59 ;
      RECT 56 3.435 56.005 3.585 ;
      RECT 55.99 3.435 56 3.583 ;
      RECT 55.98 3.433 55.99 3.581 ;
      RECT 55.95 3.425 55.98 3.575 ;
      RECT 55.935 3.417 55.95 3.568 ;
      RECT 55.915 3.412 55.935 3.561 ;
      RECT 55.91 3.408 55.915 3.556 ;
      RECT 55.88 3.401 55.91 3.55 ;
      RECT 55.855 3.392 55.88 3.54 ;
      RECT 55.825 3.385 55.855 3.532 ;
      RECT 55.8 3.375 55.825 3.523 ;
      RECT 55.785 3.367 55.8 3.517 ;
      RECT 55.76 3.362 55.785 3.512 ;
      RECT 55.75 3.358 55.76 3.507 ;
      RECT 55.73 3.353 55.75 3.502 ;
      RECT 55.695 3.348 55.73 3.495 ;
      RECT 55.635 3.343 55.695 3.488 ;
      RECT 55.622 3.339 55.635 3.486 ;
      RECT 55.536 3.334 55.622 3.483 ;
      RECT 55.45 3.324 55.536 3.479 ;
      RECT 55.409 3.317 55.45 3.476 ;
      RECT 55.323 3.31 55.409 3.473 ;
      RECT 55.237 3.3 55.323 3.469 ;
      RECT 55.151 3.29 55.237 3.464 ;
      RECT 55.065 3.28 55.151 3.46 ;
      RECT 55.055 3.265 55.065 3.458 ;
      RECT 55.045 3.25 55.055 3.458 ;
      RECT 54.98 3.245 55.045 3.457 ;
      RECT 54.815 3.242 54.86 3.45 ;
      RECT 56.06 4.147 56.065 4.338 ;
      RECT 56.055 4.142 56.06 4.345 ;
      RECT 56.041 4.14 56.055 4.351 ;
      RECT 55.955 4.14 56.041 4.353 ;
      RECT 55.951 4.14 55.955 4.356 ;
      RECT 55.865 4.14 55.951 4.374 ;
      RECT 55.855 4.145 55.865 4.393 ;
      RECT 55.845 4.2 55.855 4.397 ;
      RECT 55.82 4.215 55.845 4.404 ;
      RECT 55.78 4.235 55.82 4.417 ;
      RECT 55.775 4.247 55.78 4.427 ;
      RECT 55.76 4.253 55.775 4.432 ;
      RECT 55.755 4.258 55.76 4.436 ;
      RECT 55.735 4.265 55.755 4.441 ;
      RECT 55.665 4.29 55.735 4.458 ;
      RECT 55.625 4.318 55.665 4.478 ;
      RECT 55.62 4.328 55.625 4.486 ;
      RECT 55.6 4.335 55.62 4.488 ;
      RECT 55.595 4.342 55.6 4.491 ;
      RECT 55.565 4.35 55.595 4.494 ;
      RECT 55.56 4.355 55.565 4.498 ;
      RECT 55.486 4.359 55.56 4.506 ;
      RECT 55.4 4.368 55.486 4.522 ;
      RECT 55.396 4.373 55.4 4.531 ;
      RECT 55.31 4.378 55.396 4.541 ;
      RECT 55.27 4.386 55.31 4.553 ;
      RECT 55.22 4.392 55.27 4.56 ;
      RECT 55.135 4.401 55.22 4.575 ;
      RECT 55.06 4.412 55.135 4.593 ;
      RECT 55.025 4.419 55.06 4.603 ;
      RECT 54.95 4.427 55.025 4.608 ;
      RECT 54.895 4.436 54.95 4.608 ;
      RECT 54.87 4.441 54.895 4.606 ;
      RECT 54.86 4.444 54.87 4.604 ;
      RECT 54.825 4.446 54.86 4.602 ;
      RECT 54.795 4.448 54.825 4.598 ;
      RECT 54.75 4.447 54.795 4.594 ;
      RECT 54.73 4.442 54.75 4.591 ;
      RECT 54.68 4.427 54.73 4.588 ;
      RECT 54.67 4.412 54.68 4.583 ;
      RECT 54.62 4.397 54.67 4.573 ;
      RECT 54.57 4.372 54.62 4.553 ;
      RECT 54.56 4.357 54.57 4.535 ;
      RECT 54.555 4.355 54.56 4.529 ;
      RECT 54.535 4.35 54.555 4.524 ;
      RECT 54.53 4.342 54.535 4.518 ;
      RECT 54.515 4.336 54.53 4.511 ;
      RECT 54.51 4.331 54.515 4.503 ;
      RECT 54.49 4.326 54.51 4.495 ;
      RECT 54.475 4.319 54.49 4.488 ;
      RECT 54.46 4.313 54.475 4.479 ;
      RECT 54.455 4.307 54.46 4.472 ;
      RECT 54.41 4.282 54.455 4.458 ;
      RECT 54.395 4.252 54.41 4.44 ;
      RECT 54.38 4.235 54.395 4.431 ;
      RECT 54.355 4.215 54.38 4.419 ;
      RECT 54.315 4.185 54.355 4.399 ;
      RECT 54.305 4.155 54.315 4.384 ;
      RECT 54.29 4.145 54.305 4.377 ;
      RECT 54.235 4.11 54.29 4.356 ;
      RECT 54.22 4.073 54.235 4.335 ;
      RECT 54.21 4.06 54.22 4.327 ;
      RECT 54.16 4.03 54.21 4.309 ;
      RECT 54.145 3.96 54.16 4.29 ;
      RECT 54.1 3.96 54.145 4.273 ;
      RECT 54.075 3.96 54.1 4.255 ;
      RECT 54.065 3.96 54.075 4.248 ;
      RECT 53.986 3.96 54.065 4.241 ;
      RECT 53.9 3.96 53.986 4.233 ;
      RECT 53.885 3.992 53.9 4.228 ;
      RECT 53.81 4.002 53.885 4.224 ;
      RECT 53.79 4.012 53.81 4.219 ;
      RECT 53.765 4.012 53.79 4.216 ;
      RECT 53.755 4.002 53.765 4.215 ;
      RECT 53.745 3.975 53.755 4.214 ;
      RECT 53.705 3.97 53.745 4.212 ;
      RECT 53.66 3.97 53.705 4.208 ;
      RECT 53.635 3.97 53.66 4.203 ;
      RECT 53.585 3.97 53.635 4.19 ;
      RECT 53.545 3.975 53.555 4.175 ;
      RECT 53.555 3.97 53.585 4.18 ;
      RECT 55.54 3.75 55.8 4.01 ;
      RECT 55.535 3.772 55.8 3.968 ;
      RECT 54.775 3.6 54.995 3.965 ;
      RECT 54.757 3.687 54.995 3.964 ;
      RECT 54.74 3.692 54.995 3.961 ;
      RECT 54.74 3.692 55.015 3.96 ;
      RECT 54.71 3.702 55.015 3.958 ;
      RECT 54.705 3.717 55.015 3.954 ;
      RECT 54.705 3.717 55.02 3.953 ;
      RECT 54.7 3.775 55.02 3.951 ;
      RECT 54.7 3.775 55.03 3.948 ;
      RECT 54.695 3.84 55.03 3.943 ;
      RECT 54.775 3.6 55.035 3.86 ;
      RECT 53.52 3.43 53.78 3.69 ;
      RECT 53.52 3.473 53.866 3.664 ;
      RECT 53.52 3.473 53.91 3.663 ;
      RECT 53.52 3.473 53.93 3.661 ;
      RECT 53.52 3.473 54.03 3.66 ;
      RECT 53.52 3.473 54.05 3.658 ;
      RECT 53.52 3.473 54.06 3.653 ;
      RECT 53.93 3.44 54.12 3.65 ;
      RECT 53.93 3.442 54.125 3.648 ;
      RECT 53.92 3.447 54.13 3.64 ;
      RECT 53.866 3.471 54.13 3.64 ;
      RECT 53.91 3.465 53.92 3.662 ;
      RECT 53.92 3.445 54.125 3.648 ;
      RECT 52.875 4.505 53.08 4.735 ;
      RECT 52.815 4.455 52.87 4.715 ;
      RECT 52.875 4.455 53.075 4.735 ;
      RECT 53.845 4.77 53.85 4.797 ;
      RECT 53.835 4.68 53.845 4.802 ;
      RECT 53.83 4.602 53.835 4.808 ;
      RECT 53.82 4.592 53.83 4.815 ;
      RECT 53.815 4.582 53.82 4.821 ;
      RECT 53.805 4.577 53.815 4.823 ;
      RECT 53.79 4.569 53.805 4.831 ;
      RECT 53.775 4.56 53.79 4.843 ;
      RECT 53.765 4.552 53.775 4.853 ;
      RECT 53.73 4.47 53.765 4.871 ;
      RECT 53.695 4.47 53.73 4.89 ;
      RECT 53.68 4.47 53.695 4.898 ;
      RECT 53.625 4.47 53.68 4.898 ;
      RECT 53.591 4.47 53.625 4.889 ;
      RECT 53.505 4.47 53.591 4.865 ;
      RECT 53.495 4.53 53.505 4.847 ;
      RECT 53.455 4.532 53.495 4.838 ;
      RECT 53.45 4.534 53.455 4.828 ;
      RECT 53.43 4.536 53.45 4.823 ;
      RECT 53.42 4.539 53.43 4.818 ;
      RECT 53.41 4.54 53.42 4.813 ;
      RECT 53.386 4.541 53.41 4.805 ;
      RECT 53.3 4.546 53.386 4.783 ;
      RECT 53.245 4.545 53.3 4.756 ;
      RECT 53.23 4.538 53.245 4.743 ;
      RECT 53.195 4.533 53.23 4.739 ;
      RECT 53.14 4.525 53.195 4.738 ;
      RECT 53.08 4.512 53.14 4.736 ;
      RECT 52.87 4.455 52.875 4.723 ;
      RECT 52.945 3.825 53.13 4.035 ;
      RECT 52.935 3.83 53.145 4.028 ;
      RECT 52.975 3.735 53.235 3.995 ;
      RECT 52.93 3.892 53.235 3.918 ;
      RECT 52.275 3.685 52.28 4.485 ;
      RECT 52.22 3.735 52.25 4.485 ;
      RECT 52.21 3.735 52.215 4.045 ;
      RECT 52.195 3.735 52.2 4.04 ;
      RECT 51.74 3.78 51.755 3.995 ;
      RECT 51.67 3.78 51.755 3.99 ;
      RECT 52.935 3.36 53.005 3.57 ;
      RECT 53.005 3.367 53.015 3.565 ;
      RECT 52.901 3.36 52.935 3.577 ;
      RECT 52.815 3.36 52.901 3.601 ;
      RECT 52.805 3.365 52.815 3.62 ;
      RECT 52.8 3.377 52.805 3.623 ;
      RECT 52.785 3.392 52.8 3.627 ;
      RECT 52.78 3.41 52.785 3.631 ;
      RECT 52.74 3.42 52.78 3.64 ;
      RECT 52.725 3.427 52.74 3.652 ;
      RECT 52.71 3.432 52.725 3.657 ;
      RECT 52.695 3.435 52.71 3.662 ;
      RECT 52.685 3.437 52.695 3.666 ;
      RECT 52.65 3.444 52.685 3.674 ;
      RECT 52.615 3.452 52.65 3.688 ;
      RECT 52.605 3.458 52.615 3.697 ;
      RECT 52.6 3.46 52.605 3.699 ;
      RECT 52.58 3.463 52.6 3.705 ;
      RECT 52.55 3.47 52.58 3.716 ;
      RECT 52.54 3.476 52.55 3.723 ;
      RECT 52.515 3.479 52.54 3.73 ;
      RECT 52.505 3.483 52.515 3.738 ;
      RECT 52.5 3.484 52.505 3.76 ;
      RECT 52.495 3.485 52.5 3.775 ;
      RECT 52.49 3.486 52.495 3.79 ;
      RECT 52.485 3.487 52.49 3.805 ;
      RECT 52.48 3.488 52.485 3.835 ;
      RECT 52.47 3.49 52.48 3.868 ;
      RECT 52.455 3.494 52.47 3.915 ;
      RECT 52.445 3.497 52.455 3.96 ;
      RECT 52.44 3.5 52.445 3.988 ;
      RECT 52.43 3.502 52.44 4.015 ;
      RECT 52.425 3.505 52.43 4.05 ;
      RECT 52.395 3.51 52.425 4.108 ;
      RECT 52.39 3.515 52.395 4.193 ;
      RECT 52.385 3.517 52.39 4.228 ;
      RECT 52.38 3.519 52.385 4.31 ;
      RECT 52.375 3.521 52.38 4.398 ;
      RECT 52.365 3.523 52.375 4.48 ;
      RECT 52.35 3.537 52.365 4.485 ;
      RECT 52.315 3.582 52.35 4.485 ;
      RECT 52.305 3.622 52.315 4.485 ;
      RECT 52.29 3.65 52.305 4.485 ;
      RECT 52.285 3.667 52.29 4.485 ;
      RECT 52.28 3.675 52.285 4.485 ;
      RECT 52.27 3.69 52.275 4.485 ;
      RECT 52.265 3.697 52.27 4.485 ;
      RECT 52.255 3.717 52.265 4.485 ;
      RECT 52.25 3.73 52.255 4.485 ;
      RECT 52.215 3.735 52.22 4.07 ;
      RECT 52.2 4.125 52.22 4.485 ;
      RECT 52.2 3.735 52.21 4.043 ;
      RECT 52.195 4.165 52.2 4.485 ;
      RECT 52.145 3.735 52.195 4.038 ;
      RECT 52.19 4.202 52.195 4.485 ;
      RECT 52.18 4.225 52.19 4.485 ;
      RECT 52.175 4.27 52.18 4.485 ;
      RECT 52.165 4.28 52.175 4.478 ;
      RECT 52.091 3.735 52.145 4.032 ;
      RECT 52.005 3.735 52.091 4.025 ;
      RECT 51.956 3.782 52.005 4.018 ;
      RECT 51.87 3.79 51.956 4.011 ;
      RECT 51.855 3.787 51.87 4.006 ;
      RECT 51.841 3.78 51.855 4.005 ;
      RECT 51.755 3.78 51.841 4 ;
      RECT 51.66 3.785 51.67 3.985 ;
      RECT 51.25 3.215 51.265 3.615 ;
      RECT 51.445 3.215 51.45 3.475 ;
      RECT 51.19 3.215 51.235 3.475 ;
      RECT 51.645 4.52 51.65 4.725 ;
      RECT 51.64 4.51 51.645 4.73 ;
      RECT 51.635 4.497 51.64 4.735 ;
      RECT 51.63 4.477 51.635 4.735 ;
      RECT 51.605 4.43 51.63 4.735 ;
      RECT 51.57 4.345 51.605 4.735 ;
      RECT 51.565 4.282 51.57 4.735 ;
      RECT 51.56 4.267 51.565 4.735 ;
      RECT 51.545 4.227 51.56 4.735 ;
      RECT 51.54 4.202 51.545 4.735 ;
      RECT 51.53 4.185 51.54 4.735 ;
      RECT 51.495 4.107 51.53 4.735 ;
      RECT 51.49 4.05 51.495 4.735 ;
      RECT 51.485 4.037 51.49 4.735 ;
      RECT 51.475 4.015 51.485 4.735 ;
      RECT 51.465 3.98 51.475 4.735 ;
      RECT 51.455 3.95 51.465 4.735 ;
      RECT 51.445 3.865 51.455 4.378 ;
      RECT 51.452 4.51 51.455 4.735 ;
      RECT 51.45 4.52 51.452 4.735 ;
      RECT 51.44 4.53 51.45 4.73 ;
      RECT 51.435 3.215 51.445 3.61 ;
      RECT 51.44 3.742 51.445 4.353 ;
      RECT 51.435 3.64 51.44 4.336 ;
      RECT 51.425 3.215 51.435 4.312 ;
      RECT 51.42 3.215 51.425 4.283 ;
      RECT 51.415 3.215 51.42 4.273 ;
      RECT 51.395 3.215 51.415 4.235 ;
      RECT 51.39 3.215 51.395 4.193 ;
      RECT 51.385 3.215 51.39 4.173 ;
      RECT 51.355 3.215 51.385 4.123 ;
      RECT 51.345 3.215 51.355 4.07 ;
      RECT 51.34 3.215 51.345 4.043 ;
      RECT 51.335 3.215 51.34 4.028 ;
      RECT 51.325 3.215 51.335 4.005 ;
      RECT 51.315 3.215 51.325 3.98 ;
      RECT 51.31 3.215 51.315 3.92 ;
      RECT 51.3 3.215 51.31 3.858 ;
      RECT 51.295 3.215 51.3 3.778 ;
      RECT 51.29 3.215 51.295 3.743 ;
      RECT 51.285 3.215 51.29 3.718 ;
      RECT 51.28 3.215 51.285 3.703 ;
      RECT 51.275 3.215 51.28 3.673 ;
      RECT 51.27 3.215 51.275 3.65 ;
      RECT 51.265 3.215 51.27 3.623 ;
      RECT 51.235 3.215 51.25 3.61 ;
      RECT 50.39 4.75 50.575 4.96 ;
      RECT 50.38 4.755 50.59 4.953 ;
      RECT 50.38 4.755 50.61 4.925 ;
      RECT 50.38 4.755 50.625 4.904 ;
      RECT 50.38 4.755 50.64 4.902 ;
      RECT 50.38 4.755 50.65 4.901 ;
      RECT 50.38 4.755 50.68 4.898 ;
      RECT 51.03 4.6 51.29 4.86 ;
      RECT 50.99 4.647 51.29 4.843 ;
      RECT 50.981 4.655 50.99 4.846 ;
      RECT 50.575 4.748 51.29 4.843 ;
      RECT 50.895 4.673 50.981 4.853 ;
      RECT 50.59 4.745 51.29 4.843 ;
      RECT 50.836 4.695 50.895 4.865 ;
      RECT 50.61 4.741 51.29 4.843 ;
      RECT 50.75 4.707 50.836 4.876 ;
      RECT 50.625 4.737 51.29 4.843 ;
      RECT 50.695 4.72 50.75 4.888 ;
      RECT 50.64 4.735 51.29 4.843 ;
      RECT 50.68 4.726 50.695 4.894 ;
      RECT 50.65 4.731 51.29 4.843 ;
      RECT 50.795 4.255 51.055 4.515 ;
      RECT 50.795 4.275 51.165 4.485 ;
      RECT 50.795 4.28 51.175 4.48 ;
      RECT 50.986 3.694 51.065 3.925 ;
      RECT 50.9 3.697 51.115 3.92 ;
      RECT 50.895 3.697 51.115 3.915 ;
      RECT 50.895 3.702 51.125 3.913 ;
      RECT 50.87 3.702 51.125 3.91 ;
      RECT 50.87 3.71 51.135 3.908 ;
      RECT 50.75 3.645 51.01 3.905 ;
      RECT 50.75 3.692 51.06 3.905 ;
      RECT 50.005 4.265 50.01 4.525 ;
      RECT 49.835 4.035 49.84 4.525 ;
      RECT 49.72 4.275 49.725 4.5 ;
      RECT 50.43 3.37 50.435 3.58 ;
      RECT 50.435 3.375 50.45 3.575 ;
      RECT 50.37 3.37 50.43 3.588 ;
      RECT 50.355 3.37 50.37 3.598 ;
      RECT 50.305 3.37 50.355 3.615 ;
      RECT 50.285 3.37 50.305 3.638 ;
      RECT 50.27 3.37 50.285 3.65 ;
      RECT 50.25 3.37 50.27 3.66 ;
      RECT 50.24 3.375 50.25 3.669 ;
      RECT 50.235 3.385 50.24 3.674 ;
      RECT 50.23 3.397 50.235 3.678 ;
      RECT 50.22 3.42 50.23 3.683 ;
      RECT 50.215 3.435 50.22 3.687 ;
      RECT 50.21 3.452 50.215 3.69 ;
      RECT 50.205 3.46 50.21 3.693 ;
      RECT 50.195 3.465 50.205 3.697 ;
      RECT 50.19 3.472 50.195 3.702 ;
      RECT 50.18 3.477 50.19 3.706 ;
      RECT 50.155 3.489 50.18 3.717 ;
      RECT 50.135 3.506 50.155 3.733 ;
      RECT 50.11 3.523 50.135 3.755 ;
      RECT 50.075 3.546 50.11 3.813 ;
      RECT 50.055 3.568 50.075 3.875 ;
      RECT 50.05 3.578 50.055 3.91 ;
      RECT 50.04 3.585 50.05 3.948 ;
      RECT 50.035 3.592 50.04 3.968 ;
      RECT 50.03 3.603 50.035 4.005 ;
      RECT 50.025 3.611 50.03 4.07 ;
      RECT 50.015 3.622 50.025 4.123 ;
      RECT 50.01 3.64 50.015 4.193 ;
      RECT 50.005 3.65 50.01 4.23 ;
      RECT 50 3.66 50.005 4.525 ;
      RECT 49.995 3.672 50 4.525 ;
      RECT 49.99 3.682 49.995 4.525 ;
      RECT 49.98 3.692 49.99 4.525 ;
      RECT 49.97 3.715 49.98 4.525 ;
      RECT 49.955 3.75 49.97 4.525 ;
      RECT 49.915 3.812 49.955 4.525 ;
      RECT 49.91 3.865 49.915 4.525 ;
      RECT 49.885 3.9 49.91 4.525 ;
      RECT 49.87 3.945 49.885 4.525 ;
      RECT 49.865 3.967 49.87 4.525 ;
      RECT 49.855 3.98 49.865 4.525 ;
      RECT 49.845 4.005 49.855 4.525 ;
      RECT 49.84 4.027 49.845 4.525 ;
      RECT 49.815 4.065 49.835 4.525 ;
      RECT 49.775 4.122 49.815 4.525 ;
      RECT 49.77 4.172 49.775 4.525 ;
      RECT 49.765 4.19 49.77 4.525 ;
      RECT 49.76 4.202 49.765 4.525 ;
      RECT 49.75 4.22 49.76 4.525 ;
      RECT 49.74 4.24 49.75 4.5 ;
      RECT 49.735 4.257 49.74 4.5 ;
      RECT 49.725 4.27 49.735 4.5 ;
      RECT 49.695 4.28 49.72 4.5 ;
      RECT 49.685 4.287 49.695 4.5 ;
      RECT 49.67 4.297 49.685 4.495 ;
      RECT 48.775 10.05 49.07 10.28 ;
      RECT 48.835 8.57 49.005 10.28 ;
      RECT 48.82 8.945 49.175 9.3 ;
      RECT 48.775 8.57 49.065 8.8 ;
      RECT 48.795 7.215 49.075 7.585 ;
      RECT 48.75 7.215 49.1 7.565 ;
      RECT 47.78 10.055 48.075 10.285 ;
      RECT 47.84 8.575 48.01 10.285 ;
      RECT 47.78 8.575 48.07 8.805 ;
      RECT 47.78 8.61 48.635 8.77 ;
      RECT 48.465 8.2 48.635 8.77 ;
      RECT 47.78 8.605 48.175 8.77 ;
      RECT 48.405 8.2 48.695 8.43 ;
      RECT 48.405 8.23 48.865 8.4 ;
      RECT 48.365 4.03 48.69 4.26 ;
      RECT 48.365 4.06 48.86 4.23 ;
      RECT 48.365 3.69 48.555 4.26 ;
      RECT 47.78 3.655 48.07 3.885 ;
      RECT 47.78 3.69 48.555 3.86 ;
      RECT 47.84 2.175 48.01 3.885 ;
      RECT 47.78 2.175 48.075 2.405 ;
      RECT 47.41 4.025 47.7 4.255 ;
      RECT 47.41 4.055 47.87 4.225 ;
      RECT 47.475 2.95 47.64 4.255 ;
      RECT 45.99 2.915 46.28 3.145 ;
      RECT 45.99 2.95 47.64 3.12 ;
      RECT 46.05 2.175 46.22 3.145 ;
      RECT 45.99 2.175 46.28 2.405 ;
      RECT 45.99 10.055 46.28 10.285 ;
      RECT 46.05 9.315 46.22 10.285 ;
      RECT 46.05 9.405 47.64 9.575 ;
      RECT 47.47 8.205 47.64 9.575 ;
      RECT 45.99 9.315 46.28 9.545 ;
      RECT 47.41 8.205 47.7 8.435 ;
      RECT 47.41 8.235 47.87 8.405 ;
      RECT 46.42 3.26 46.77 3.61 ;
      RECT 44.085 3.32 46.77 3.49 ;
      RECT 46.25 3.315 46.77 3.49 ;
      RECT 44.085 2.635 44.255 3.49 ;
      RECT 43.985 2.635 44.335 2.985 ;
      RECT 46.445 8.94 46.77 9.265 ;
      RECT 41.87 8.895 42.22 9.245 ;
      RECT 46.42 8.945 46.77 9.175 ;
      RECT 41.64 8.945 42.22 9.175 ;
      RECT 46.25 8.97 46.77 9.145 ;
      RECT 41.47 8.975 42.22 9.145 ;
      RECT 41.64 8.97 46.77 9.14 ;
      RECT 45.645 3.66 45.965 3.98 ;
      RECT 45.62 3.655 45.91 3.885 ;
      RECT 45.545 3.685 45.965 3.86 ;
      RECT 45.445 3.685 45.965 3.855 ;
      RECT 45.645 8.54 45.965 8.83 ;
      RECT 45.62 8.575 45.965 8.805 ;
      RECT 45.445 8.605 45.965 8.775 ;
      RECT 42.28 3.76 42.465 3.97 ;
      RECT 42.27 3.765 42.48 3.963 ;
      RECT 42.27 3.765 42.566 3.94 ;
      RECT 42.27 3.765 42.625 3.915 ;
      RECT 42.27 3.765 42.68 3.895 ;
      RECT 42.27 3.765 42.69 3.883 ;
      RECT 42.27 3.765 42.885 3.822 ;
      RECT 42.27 3.765 42.915 3.805 ;
      RECT 42.27 3.765 42.935 3.795 ;
      RECT 42.815 3.53 43.075 3.79 ;
      RECT 42.8 3.62 42.815 3.837 ;
      RECT 42.335 3.752 43.075 3.79 ;
      RECT 42.786 3.631 42.8 3.843 ;
      RECT 42.375 3.745 43.075 3.79 ;
      RECT 42.7 3.671 42.786 3.862 ;
      RECT 42.625 3.732 43.075 3.79 ;
      RECT 42.695 3.707 42.7 3.879 ;
      RECT 42.68 3.717 43.075 3.79 ;
      RECT 42.69 3.712 42.695 3.881 ;
      RECT 41.615 3.795 41.72 4.055 ;
      RECT 42.43 3.32 42.435 3.545 ;
      RECT 42.56 3.32 42.615 3.53 ;
      RECT 42.615 3.325 42.625 3.523 ;
      RECT 42.521 3.32 42.56 3.533 ;
      RECT 42.435 3.32 42.521 3.54 ;
      RECT 42.415 3.325 42.43 3.546 ;
      RECT 42.405 3.365 42.415 3.548 ;
      RECT 42.375 3.375 42.405 3.55 ;
      RECT 42.37 3.38 42.375 3.552 ;
      RECT 42.345 3.385 42.37 3.554 ;
      RECT 42.33 3.39 42.345 3.556 ;
      RECT 42.315 3.392 42.33 3.558 ;
      RECT 42.31 3.397 42.315 3.56 ;
      RECT 42.26 3.405 42.31 3.563 ;
      RECT 42.235 3.414 42.26 3.568 ;
      RECT 42.225 3.421 42.235 3.573 ;
      RECT 42.22 3.424 42.225 3.577 ;
      RECT 42.2 3.427 42.22 3.586 ;
      RECT 42.17 3.435 42.2 3.606 ;
      RECT 42.141 3.448 42.17 3.628 ;
      RECT 42.055 3.482 42.141 3.672 ;
      RECT 42.05 3.508 42.055 3.71 ;
      RECT 42.045 3.512 42.05 3.719 ;
      RECT 42.01 3.525 42.045 3.752 ;
      RECT 42 3.539 42.01 3.79 ;
      RECT 41.995 3.543 42 3.803 ;
      RECT 41.99 3.547 41.995 3.808 ;
      RECT 41.98 3.555 41.99 3.82 ;
      RECT 41.975 3.562 41.98 3.835 ;
      RECT 41.95 3.575 41.975 3.86 ;
      RECT 41.91 3.604 41.95 3.915 ;
      RECT 41.895 3.629 41.91 3.97 ;
      RECT 41.885 3.64 41.895 3.993 ;
      RECT 41.88 3.647 41.885 4.005 ;
      RECT 41.875 3.651 41.88 4.013 ;
      RECT 41.82 3.679 41.875 4.055 ;
      RECT 41.8 3.715 41.82 4.055 ;
      RECT 41.785 3.73 41.8 4.055 ;
      RECT 41.73 3.762 41.785 4.055 ;
      RECT 41.72 3.792 41.73 4.055 ;
      RECT 41.33 3.407 41.515 3.645 ;
      RECT 41.315 3.409 41.525 3.64 ;
      RECT 41.2 3.355 41.46 3.615 ;
      RECT 41.195 3.392 41.46 3.569 ;
      RECT 41.19 3.402 41.46 3.566 ;
      RECT 41.185 3.442 41.525 3.56 ;
      RECT 41.18 3.475 41.525 3.55 ;
      RECT 41.19 3.417 41.54 3.488 ;
      RECT 41.487 4.515 41.5 5.045 ;
      RECT 41.401 4.515 41.5 5.044 ;
      RECT 41.401 4.515 41.505 5.043 ;
      RECT 41.315 4.515 41.505 5.041 ;
      RECT 41.31 4.515 41.505 5.038 ;
      RECT 41.31 4.515 41.515 5.036 ;
      RECT 41.305 4.807 41.515 5.033 ;
      RECT 41.305 4.817 41.52 5.03 ;
      RECT 41.305 4.885 41.525 5.026 ;
      RECT 41.295 4.89 41.525 5.025 ;
      RECT 41.295 4.982 41.53 5.022 ;
      RECT 41.28 4.515 41.54 4.775 ;
      RECT 41.21 10.055 41.5 10.285 ;
      RECT 41.27 9.315 41.44 10.285 ;
      RECT 41.185 9.34 41.525 9.685 ;
      RECT 41.21 9.315 41.5 9.685 ;
      RECT 40.51 3.505 40.555 5.04 ;
      RECT 40.71 3.505 40.74 3.72 ;
      RECT 39.085 3.245 39.205 3.455 ;
      RECT 38.745 3.195 39.005 3.455 ;
      RECT 38.745 3.24 39.04 3.445 ;
      RECT 40.75 3.521 40.755 3.575 ;
      RECT 40.745 3.514 40.75 3.708 ;
      RECT 40.74 3.508 40.745 3.715 ;
      RECT 40.695 3.505 40.71 3.728 ;
      RECT 40.69 3.505 40.695 3.75 ;
      RECT 40.685 3.505 40.69 3.798 ;
      RECT 40.68 3.505 40.685 3.818 ;
      RECT 40.67 3.505 40.68 3.925 ;
      RECT 40.665 3.505 40.67 3.988 ;
      RECT 40.66 3.505 40.665 4.045 ;
      RECT 40.655 3.505 40.66 4.053 ;
      RECT 40.64 3.505 40.655 4.16 ;
      RECT 40.63 3.505 40.64 4.295 ;
      RECT 40.62 3.505 40.63 4.405 ;
      RECT 40.61 3.505 40.62 4.462 ;
      RECT 40.605 3.505 40.61 4.502 ;
      RECT 40.6 3.505 40.605 4.538 ;
      RECT 40.59 3.505 40.6 4.578 ;
      RECT 40.585 3.505 40.59 4.62 ;
      RECT 40.565 3.505 40.585 4.685 ;
      RECT 40.57 4.83 40.575 5.01 ;
      RECT 40.565 4.812 40.57 5.018 ;
      RECT 40.56 3.505 40.565 4.748 ;
      RECT 40.56 4.792 40.565 5.025 ;
      RECT 40.555 3.505 40.56 5.035 ;
      RECT 40.5 3.505 40.51 3.805 ;
      RECT 40.505 4.052 40.51 5.04 ;
      RECT 40.5 4.117 40.505 5.04 ;
      RECT 40.495 3.506 40.5 3.795 ;
      RECT 40.49 4.182 40.5 5.04 ;
      RECT 40.485 3.507 40.495 3.785 ;
      RECT 40.475 4.295 40.49 5.04 ;
      RECT 40.48 3.508 40.485 3.775 ;
      RECT 40.46 3.509 40.48 3.753 ;
      RECT 40.465 4.392 40.475 5.04 ;
      RECT 40.46 4.467 40.465 5.04 ;
      RECT 40.45 3.508 40.46 3.73 ;
      RECT 40.455 4.51 40.46 5.04 ;
      RECT 40.45 4.537 40.455 5.04 ;
      RECT 40.44 3.506 40.45 3.718 ;
      RECT 40.445 4.58 40.45 5.04 ;
      RECT 40.44 4.607 40.445 5.04 ;
      RECT 40.43 3.505 40.44 3.705 ;
      RECT 40.435 4.622 40.44 5.04 ;
      RECT 40.395 4.68 40.435 5.04 ;
      RECT 40.425 3.504 40.43 3.69 ;
      RECT 40.42 3.502 40.425 3.683 ;
      RECT 40.41 3.499 40.42 3.673 ;
      RECT 40.405 3.496 40.41 3.658 ;
      RECT 40.39 3.492 40.405 3.651 ;
      RECT 40.385 4.735 40.395 5.04 ;
      RECT 40.385 3.489 40.39 3.646 ;
      RECT 40.37 3.485 40.385 3.64 ;
      RECT 40.38 4.752 40.385 5.04 ;
      RECT 40.37 4.815 40.38 5.04 ;
      RECT 40.29 3.47 40.37 3.62 ;
      RECT 40.365 4.822 40.37 5.035 ;
      RECT 40.36 4.83 40.365 5.025 ;
      RECT 40.28 3.456 40.29 3.604 ;
      RECT 40.265 3.452 40.28 3.602 ;
      RECT 40.255 3.447 40.265 3.598 ;
      RECT 40.23 3.44 40.255 3.59 ;
      RECT 40.225 3.435 40.23 3.585 ;
      RECT 40.215 3.435 40.225 3.583 ;
      RECT 40.205 3.433 40.215 3.581 ;
      RECT 40.175 3.425 40.205 3.575 ;
      RECT 40.16 3.417 40.175 3.568 ;
      RECT 40.14 3.412 40.16 3.561 ;
      RECT 40.135 3.408 40.14 3.556 ;
      RECT 40.105 3.401 40.135 3.55 ;
      RECT 40.08 3.392 40.105 3.54 ;
      RECT 40.05 3.385 40.08 3.532 ;
      RECT 40.025 3.375 40.05 3.523 ;
      RECT 40.01 3.367 40.025 3.517 ;
      RECT 39.985 3.362 40.01 3.512 ;
      RECT 39.975 3.358 39.985 3.507 ;
      RECT 39.955 3.353 39.975 3.502 ;
      RECT 39.92 3.348 39.955 3.495 ;
      RECT 39.86 3.343 39.92 3.488 ;
      RECT 39.847 3.339 39.86 3.486 ;
      RECT 39.761 3.334 39.847 3.483 ;
      RECT 39.675 3.324 39.761 3.479 ;
      RECT 39.634 3.317 39.675 3.476 ;
      RECT 39.548 3.31 39.634 3.473 ;
      RECT 39.462 3.3 39.548 3.469 ;
      RECT 39.376 3.29 39.462 3.464 ;
      RECT 39.29 3.28 39.376 3.46 ;
      RECT 39.28 3.265 39.29 3.458 ;
      RECT 39.27 3.25 39.28 3.458 ;
      RECT 39.205 3.245 39.27 3.457 ;
      RECT 39.04 3.242 39.085 3.45 ;
      RECT 40.285 4.147 40.29 4.338 ;
      RECT 40.28 4.142 40.285 4.345 ;
      RECT 40.266 4.14 40.28 4.351 ;
      RECT 40.18 4.14 40.266 4.353 ;
      RECT 40.176 4.14 40.18 4.356 ;
      RECT 40.09 4.14 40.176 4.374 ;
      RECT 40.08 4.145 40.09 4.393 ;
      RECT 40.07 4.2 40.08 4.397 ;
      RECT 40.045 4.215 40.07 4.404 ;
      RECT 40.005 4.235 40.045 4.417 ;
      RECT 40 4.247 40.005 4.427 ;
      RECT 39.985 4.253 40 4.432 ;
      RECT 39.98 4.258 39.985 4.436 ;
      RECT 39.96 4.265 39.98 4.441 ;
      RECT 39.89 4.29 39.96 4.458 ;
      RECT 39.85 4.318 39.89 4.478 ;
      RECT 39.845 4.328 39.85 4.486 ;
      RECT 39.825 4.335 39.845 4.488 ;
      RECT 39.82 4.342 39.825 4.491 ;
      RECT 39.79 4.35 39.82 4.494 ;
      RECT 39.785 4.355 39.79 4.498 ;
      RECT 39.711 4.359 39.785 4.506 ;
      RECT 39.625 4.368 39.711 4.522 ;
      RECT 39.621 4.373 39.625 4.531 ;
      RECT 39.535 4.378 39.621 4.541 ;
      RECT 39.495 4.386 39.535 4.553 ;
      RECT 39.445 4.392 39.495 4.56 ;
      RECT 39.36 4.401 39.445 4.575 ;
      RECT 39.285 4.412 39.36 4.593 ;
      RECT 39.25 4.419 39.285 4.603 ;
      RECT 39.175 4.427 39.25 4.608 ;
      RECT 39.12 4.436 39.175 4.608 ;
      RECT 39.095 4.441 39.12 4.606 ;
      RECT 39.085 4.444 39.095 4.604 ;
      RECT 39.05 4.446 39.085 4.602 ;
      RECT 39.02 4.448 39.05 4.598 ;
      RECT 38.975 4.447 39.02 4.594 ;
      RECT 38.955 4.442 38.975 4.591 ;
      RECT 38.905 4.427 38.955 4.588 ;
      RECT 38.895 4.412 38.905 4.583 ;
      RECT 38.845 4.397 38.895 4.573 ;
      RECT 38.795 4.372 38.845 4.553 ;
      RECT 38.785 4.357 38.795 4.535 ;
      RECT 38.78 4.355 38.785 4.529 ;
      RECT 38.76 4.35 38.78 4.524 ;
      RECT 38.755 4.342 38.76 4.518 ;
      RECT 38.74 4.336 38.755 4.511 ;
      RECT 38.735 4.331 38.74 4.503 ;
      RECT 38.715 4.326 38.735 4.495 ;
      RECT 38.7 4.319 38.715 4.488 ;
      RECT 38.685 4.313 38.7 4.479 ;
      RECT 38.68 4.307 38.685 4.472 ;
      RECT 38.635 4.282 38.68 4.458 ;
      RECT 38.62 4.252 38.635 4.44 ;
      RECT 38.605 4.235 38.62 4.431 ;
      RECT 38.58 4.215 38.605 4.419 ;
      RECT 38.54 4.185 38.58 4.399 ;
      RECT 38.53 4.155 38.54 4.384 ;
      RECT 38.515 4.145 38.53 4.377 ;
      RECT 38.46 4.11 38.515 4.356 ;
      RECT 38.445 4.073 38.46 4.335 ;
      RECT 38.435 4.06 38.445 4.327 ;
      RECT 38.385 4.03 38.435 4.309 ;
      RECT 38.37 3.96 38.385 4.29 ;
      RECT 38.325 3.96 38.37 4.273 ;
      RECT 38.3 3.96 38.325 4.255 ;
      RECT 38.29 3.96 38.3 4.248 ;
      RECT 38.211 3.96 38.29 4.241 ;
      RECT 38.125 3.96 38.211 4.233 ;
      RECT 38.11 3.992 38.125 4.228 ;
      RECT 38.035 4.002 38.11 4.224 ;
      RECT 38.015 4.012 38.035 4.219 ;
      RECT 37.99 4.012 38.015 4.216 ;
      RECT 37.98 4.002 37.99 4.215 ;
      RECT 37.97 3.975 37.98 4.214 ;
      RECT 37.93 3.97 37.97 4.212 ;
      RECT 37.885 3.97 37.93 4.208 ;
      RECT 37.86 3.97 37.885 4.203 ;
      RECT 37.81 3.97 37.86 4.19 ;
      RECT 37.77 3.975 37.78 4.175 ;
      RECT 37.78 3.97 37.81 4.18 ;
      RECT 39.765 3.75 40.025 4.01 ;
      RECT 39.76 3.772 40.025 3.968 ;
      RECT 39 3.6 39.22 3.965 ;
      RECT 38.982 3.687 39.22 3.964 ;
      RECT 38.965 3.692 39.22 3.961 ;
      RECT 38.965 3.692 39.24 3.96 ;
      RECT 38.935 3.702 39.24 3.958 ;
      RECT 38.93 3.717 39.24 3.954 ;
      RECT 38.93 3.717 39.245 3.953 ;
      RECT 38.925 3.775 39.245 3.951 ;
      RECT 38.925 3.775 39.255 3.948 ;
      RECT 38.92 3.84 39.255 3.943 ;
      RECT 39 3.6 39.26 3.86 ;
      RECT 37.745 3.43 38.005 3.69 ;
      RECT 37.745 3.473 38.091 3.664 ;
      RECT 37.745 3.473 38.135 3.663 ;
      RECT 37.745 3.473 38.155 3.661 ;
      RECT 37.745 3.473 38.255 3.66 ;
      RECT 37.745 3.473 38.275 3.658 ;
      RECT 37.745 3.473 38.285 3.653 ;
      RECT 38.155 3.44 38.345 3.65 ;
      RECT 38.155 3.442 38.35 3.648 ;
      RECT 38.145 3.447 38.355 3.64 ;
      RECT 38.091 3.471 38.355 3.64 ;
      RECT 38.135 3.465 38.145 3.662 ;
      RECT 38.145 3.445 38.35 3.648 ;
      RECT 37.1 4.505 37.305 4.735 ;
      RECT 37.04 4.455 37.095 4.715 ;
      RECT 37.1 4.455 37.3 4.735 ;
      RECT 38.07 4.77 38.075 4.797 ;
      RECT 38.06 4.68 38.07 4.802 ;
      RECT 38.055 4.602 38.06 4.808 ;
      RECT 38.045 4.592 38.055 4.815 ;
      RECT 38.04 4.582 38.045 4.821 ;
      RECT 38.03 4.577 38.04 4.823 ;
      RECT 38.015 4.569 38.03 4.831 ;
      RECT 38 4.56 38.015 4.843 ;
      RECT 37.99 4.552 38 4.853 ;
      RECT 37.955 4.47 37.99 4.871 ;
      RECT 37.92 4.47 37.955 4.89 ;
      RECT 37.905 4.47 37.92 4.898 ;
      RECT 37.85 4.47 37.905 4.898 ;
      RECT 37.816 4.47 37.85 4.889 ;
      RECT 37.73 4.47 37.816 4.865 ;
      RECT 37.72 4.53 37.73 4.847 ;
      RECT 37.68 4.532 37.72 4.838 ;
      RECT 37.675 4.534 37.68 4.828 ;
      RECT 37.655 4.536 37.675 4.823 ;
      RECT 37.645 4.539 37.655 4.818 ;
      RECT 37.635 4.54 37.645 4.813 ;
      RECT 37.611 4.541 37.635 4.805 ;
      RECT 37.525 4.546 37.611 4.783 ;
      RECT 37.47 4.545 37.525 4.756 ;
      RECT 37.455 4.538 37.47 4.743 ;
      RECT 37.42 4.533 37.455 4.739 ;
      RECT 37.365 4.525 37.42 4.738 ;
      RECT 37.305 4.512 37.365 4.736 ;
      RECT 37.095 4.455 37.1 4.723 ;
      RECT 37.17 3.825 37.355 4.035 ;
      RECT 37.16 3.83 37.37 4.028 ;
      RECT 37.2 3.735 37.46 3.995 ;
      RECT 37.155 3.892 37.46 3.918 ;
      RECT 36.5 3.685 36.505 4.485 ;
      RECT 36.445 3.735 36.475 4.485 ;
      RECT 36.435 3.735 36.44 4.045 ;
      RECT 36.42 3.735 36.425 4.04 ;
      RECT 35.965 3.78 35.98 3.995 ;
      RECT 35.895 3.78 35.98 3.99 ;
      RECT 37.16 3.36 37.23 3.57 ;
      RECT 37.23 3.367 37.24 3.565 ;
      RECT 37.126 3.36 37.16 3.577 ;
      RECT 37.04 3.36 37.126 3.601 ;
      RECT 37.03 3.365 37.04 3.62 ;
      RECT 37.025 3.377 37.03 3.623 ;
      RECT 37.01 3.392 37.025 3.627 ;
      RECT 37.005 3.41 37.01 3.631 ;
      RECT 36.965 3.42 37.005 3.64 ;
      RECT 36.95 3.427 36.965 3.652 ;
      RECT 36.935 3.432 36.95 3.657 ;
      RECT 36.92 3.435 36.935 3.662 ;
      RECT 36.91 3.437 36.92 3.666 ;
      RECT 36.875 3.444 36.91 3.674 ;
      RECT 36.84 3.452 36.875 3.688 ;
      RECT 36.83 3.458 36.84 3.697 ;
      RECT 36.825 3.46 36.83 3.699 ;
      RECT 36.805 3.463 36.825 3.705 ;
      RECT 36.775 3.47 36.805 3.716 ;
      RECT 36.765 3.476 36.775 3.723 ;
      RECT 36.74 3.479 36.765 3.73 ;
      RECT 36.73 3.483 36.74 3.738 ;
      RECT 36.725 3.484 36.73 3.76 ;
      RECT 36.72 3.485 36.725 3.775 ;
      RECT 36.715 3.486 36.72 3.79 ;
      RECT 36.71 3.487 36.715 3.805 ;
      RECT 36.705 3.488 36.71 3.835 ;
      RECT 36.695 3.49 36.705 3.868 ;
      RECT 36.68 3.494 36.695 3.915 ;
      RECT 36.67 3.497 36.68 3.96 ;
      RECT 36.665 3.5 36.67 3.988 ;
      RECT 36.655 3.502 36.665 4.015 ;
      RECT 36.65 3.505 36.655 4.05 ;
      RECT 36.62 3.51 36.65 4.108 ;
      RECT 36.615 3.515 36.62 4.193 ;
      RECT 36.61 3.517 36.615 4.228 ;
      RECT 36.605 3.519 36.61 4.31 ;
      RECT 36.6 3.521 36.605 4.398 ;
      RECT 36.59 3.523 36.6 4.48 ;
      RECT 36.575 3.537 36.59 4.485 ;
      RECT 36.54 3.582 36.575 4.485 ;
      RECT 36.53 3.622 36.54 4.485 ;
      RECT 36.515 3.65 36.53 4.485 ;
      RECT 36.51 3.667 36.515 4.485 ;
      RECT 36.505 3.675 36.51 4.485 ;
      RECT 36.495 3.69 36.5 4.485 ;
      RECT 36.49 3.697 36.495 4.485 ;
      RECT 36.48 3.717 36.49 4.485 ;
      RECT 36.475 3.73 36.48 4.485 ;
      RECT 36.44 3.735 36.445 4.07 ;
      RECT 36.425 4.125 36.445 4.485 ;
      RECT 36.425 3.735 36.435 4.043 ;
      RECT 36.42 4.165 36.425 4.485 ;
      RECT 36.37 3.735 36.42 4.038 ;
      RECT 36.415 4.202 36.42 4.485 ;
      RECT 36.405 4.225 36.415 4.485 ;
      RECT 36.4 4.27 36.405 4.485 ;
      RECT 36.39 4.28 36.4 4.478 ;
      RECT 36.316 3.735 36.37 4.032 ;
      RECT 36.23 3.735 36.316 4.025 ;
      RECT 36.181 3.782 36.23 4.018 ;
      RECT 36.095 3.79 36.181 4.011 ;
      RECT 36.08 3.787 36.095 4.006 ;
      RECT 36.066 3.78 36.08 4.005 ;
      RECT 35.98 3.78 36.066 4 ;
      RECT 35.885 3.785 35.895 3.985 ;
      RECT 35.475 3.215 35.49 3.615 ;
      RECT 35.67 3.215 35.675 3.475 ;
      RECT 35.415 3.215 35.46 3.475 ;
      RECT 35.87 4.52 35.875 4.725 ;
      RECT 35.865 4.51 35.87 4.73 ;
      RECT 35.86 4.497 35.865 4.735 ;
      RECT 35.855 4.477 35.86 4.735 ;
      RECT 35.83 4.43 35.855 4.735 ;
      RECT 35.795 4.345 35.83 4.735 ;
      RECT 35.79 4.282 35.795 4.735 ;
      RECT 35.785 4.267 35.79 4.735 ;
      RECT 35.77 4.227 35.785 4.735 ;
      RECT 35.765 4.202 35.77 4.735 ;
      RECT 35.755 4.185 35.765 4.735 ;
      RECT 35.72 4.107 35.755 4.735 ;
      RECT 35.715 4.05 35.72 4.735 ;
      RECT 35.71 4.037 35.715 4.735 ;
      RECT 35.7 4.015 35.71 4.735 ;
      RECT 35.69 3.98 35.7 4.735 ;
      RECT 35.68 3.95 35.69 4.735 ;
      RECT 35.67 3.865 35.68 4.378 ;
      RECT 35.677 4.51 35.68 4.735 ;
      RECT 35.675 4.52 35.677 4.735 ;
      RECT 35.665 4.53 35.675 4.73 ;
      RECT 35.66 3.215 35.67 3.61 ;
      RECT 35.665 3.742 35.67 4.353 ;
      RECT 35.66 3.64 35.665 4.336 ;
      RECT 35.65 3.215 35.66 4.312 ;
      RECT 35.645 3.215 35.65 4.283 ;
      RECT 35.64 3.215 35.645 4.273 ;
      RECT 35.62 3.215 35.64 4.235 ;
      RECT 35.615 3.215 35.62 4.193 ;
      RECT 35.61 3.215 35.615 4.173 ;
      RECT 35.58 3.215 35.61 4.123 ;
      RECT 35.57 3.215 35.58 4.07 ;
      RECT 35.565 3.215 35.57 4.043 ;
      RECT 35.56 3.215 35.565 4.028 ;
      RECT 35.55 3.215 35.56 4.005 ;
      RECT 35.54 3.215 35.55 3.98 ;
      RECT 35.535 3.215 35.54 3.92 ;
      RECT 35.525 3.215 35.535 3.858 ;
      RECT 35.52 3.215 35.525 3.778 ;
      RECT 35.515 3.215 35.52 3.743 ;
      RECT 35.51 3.215 35.515 3.718 ;
      RECT 35.505 3.215 35.51 3.703 ;
      RECT 35.5 3.215 35.505 3.673 ;
      RECT 35.495 3.215 35.5 3.65 ;
      RECT 35.49 3.215 35.495 3.623 ;
      RECT 35.46 3.215 35.475 3.61 ;
      RECT 34.615 4.75 34.8 4.96 ;
      RECT 34.605 4.755 34.815 4.953 ;
      RECT 34.605 4.755 34.835 4.925 ;
      RECT 34.605 4.755 34.85 4.904 ;
      RECT 34.605 4.755 34.865 4.902 ;
      RECT 34.605 4.755 34.875 4.901 ;
      RECT 34.605 4.755 34.905 4.898 ;
      RECT 35.255 4.6 35.515 4.86 ;
      RECT 35.215 4.647 35.515 4.843 ;
      RECT 35.206 4.655 35.215 4.846 ;
      RECT 34.8 4.748 35.515 4.843 ;
      RECT 35.12 4.673 35.206 4.853 ;
      RECT 34.815 4.745 35.515 4.843 ;
      RECT 35.061 4.695 35.12 4.865 ;
      RECT 34.835 4.741 35.515 4.843 ;
      RECT 34.975 4.707 35.061 4.876 ;
      RECT 34.85 4.737 35.515 4.843 ;
      RECT 34.92 4.72 34.975 4.888 ;
      RECT 34.865 4.735 35.515 4.843 ;
      RECT 34.905 4.726 34.92 4.894 ;
      RECT 34.875 4.731 35.515 4.843 ;
      RECT 35.02 4.255 35.28 4.515 ;
      RECT 35.02 4.275 35.39 4.485 ;
      RECT 35.02 4.28 35.4 4.48 ;
      RECT 35.211 3.694 35.29 3.925 ;
      RECT 35.125 3.697 35.34 3.92 ;
      RECT 35.12 3.697 35.34 3.915 ;
      RECT 35.12 3.702 35.35 3.913 ;
      RECT 35.095 3.702 35.35 3.91 ;
      RECT 35.095 3.71 35.36 3.908 ;
      RECT 34.975 3.645 35.235 3.905 ;
      RECT 34.975 3.692 35.285 3.905 ;
      RECT 34.23 4.265 34.235 4.525 ;
      RECT 34.06 4.035 34.065 4.525 ;
      RECT 33.945 4.275 33.95 4.5 ;
      RECT 34.655 3.37 34.66 3.58 ;
      RECT 34.66 3.375 34.675 3.575 ;
      RECT 34.595 3.37 34.655 3.588 ;
      RECT 34.58 3.37 34.595 3.598 ;
      RECT 34.53 3.37 34.58 3.615 ;
      RECT 34.51 3.37 34.53 3.638 ;
      RECT 34.495 3.37 34.51 3.65 ;
      RECT 34.475 3.37 34.495 3.66 ;
      RECT 34.465 3.375 34.475 3.669 ;
      RECT 34.46 3.385 34.465 3.674 ;
      RECT 34.455 3.397 34.46 3.678 ;
      RECT 34.445 3.42 34.455 3.683 ;
      RECT 34.44 3.435 34.445 3.687 ;
      RECT 34.435 3.452 34.44 3.69 ;
      RECT 34.43 3.46 34.435 3.693 ;
      RECT 34.42 3.465 34.43 3.697 ;
      RECT 34.415 3.472 34.42 3.702 ;
      RECT 34.405 3.477 34.415 3.706 ;
      RECT 34.38 3.489 34.405 3.717 ;
      RECT 34.36 3.506 34.38 3.733 ;
      RECT 34.335 3.523 34.36 3.755 ;
      RECT 34.3 3.546 34.335 3.813 ;
      RECT 34.28 3.568 34.3 3.875 ;
      RECT 34.275 3.578 34.28 3.91 ;
      RECT 34.265 3.585 34.275 3.948 ;
      RECT 34.26 3.592 34.265 3.968 ;
      RECT 34.255 3.603 34.26 4.005 ;
      RECT 34.25 3.611 34.255 4.07 ;
      RECT 34.24 3.622 34.25 4.123 ;
      RECT 34.235 3.64 34.24 4.193 ;
      RECT 34.23 3.65 34.235 4.23 ;
      RECT 34.225 3.66 34.23 4.525 ;
      RECT 34.22 3.672 34.225 4.525 ;
      RECT 34.215 3.682 34.22 4.525 ;
      RECT 34.205 3.692 34.215 4.525 ;
      RECT 34.195 3.715 34.205 4.525 ;
      RECT 34.18 3.75 34.195 4.525 ;
      RECT 34.14 3.812 34.18 4.525 ;
      RECT 34.135 3.865 34.14 4.525 ;
      RECT 34.11 3.9 34.135 4.525 ;
      RECT 34.095 3.945 34.11 4.525 ;
      RECT 34.09 3.967 34.095 4.525 ;
      RECT 34.08 3.98 34.09 4.525 ;
      RECT 34.07 4.005 34.08 4.525 ;
      RECT 34.065 4.027 34.07 4.525 ;
      RECT 34.04 4.065 34.06 4.525 ;
      RECT 34 4.122 34.04 4.525 ;
      RECT 33.995 4.172 34 4.525 ;
      RECT 33.99 4.19 33.995 4.525 ;
      RECT 33.985 4.202 33.99 4.525 ;
      RECT 33.975 4.22 33.985 4.525 ;
      RECT 33.965 4.24 33.975 4.5 ;
      RECT 33.96 4.257 33.965 4.5 ;
      RECT 33.95 4.27 33.96 4.5 ;
      RECT 33.92 4.28 33.945 4.5 ;
      RECT 33.91 4.287 33.92 4.5 ;
      RECT 33.895 4.297 33.91 4.495 ;
      RECT 32.995 10.05 33.29 10.28 ;
      RECT 33.055 8.57 33.225 10.28 ;
      RECT 33.045 8.94 33.395 9.29 ;
      RECT 32.995 8.57 33.285 8.8 ;
      RECT 33.015 7.215 33.295 7.585 ;
      RECT 32.97 7.215 33.32 7.565 ;
      RECT 32 10.055 32.295 10.285 ;
      RECT 32.06 8.575 32.23 10.285 ;
      RECT 32 8.575 32.29 8.805 ;
      RECT 32 8.61 32.855 8.77 ;
      RECT 32.685 8.2 32.855 8.77 ;
      RECT 32 8.605 32.395 8.77 ;
      RECT 32.625 8.2 32.915 8.43 ;
      RECT 32.625 8.23 33.085 8.4 ;
      RECT 32.585 4.03 32.91 4.26 ;
      RECT 32.585 4.06 33.08 4.23 ;
      RECT 32.585 3.69 32.775 4.26 ;
      RECT 32 3.655 32.29 3.885 ;
      RECT 32 3.69 32.775 3.86 ;
      RECT 32.06 2.175 32.23 3.885 ;
      RECT 32 2.175 32.295 2.405 ;
      RECT 31.63 4.025 31.92 4.255 ;
      RECT 31.63 4.055 32.09 4.225 ;
      RECT 31.695 2.95 31.86 4.255 ;
      RECT 30.21 2.915 30.5 3.145 ;
      RECT 30.21 2.95 31.86 3.12 ;
      RECT 30.27 2.175 30.44 3.145 ;
      RECT 30.21 2.175 30.5 2.405 ;
      RECT 30.21 10.055 30.5 10.285 ;
      RECT 30.27 9.315 30.44 10.285 ;
      RECT 30.27 9.405 31.86 9.575 ;
      RECT 31.69 8.205 31.86 9.575 ;
      RECT 30.21 9.315 30.5 9.545 ;
      RECT 31.63 8.205 31.92 8.435 ;
      RECT 31.63 8.235 32.09 8.405 ;
      RECT 30.64 3.26 30.99 3.61 ;
      RECT 28.305 3.32 30.99 3.49 ;
      RECT 30.47 3.315 30.99 3.49 ;
      RECT 28.305 2.635 28.475 3.49 ;
      RECT 28.205 2.635 28.555 2.985 ;
      RECT 30.665 8.94 30.99 9.265 ;
      RECT 26.06 8.89 26.41 9.24 ;
      RECT 30.64 8.945 30.99 9.175 ;
      RECT 25.86 8.945 26.41 9.175 ;
      RECT 30.47 8.97 30.99 9.145 ;
      RECT 25.69 8.975 26.41 9.145 ;
      RECT 25.86 8.97 30.99 9.14 ;
      RECT 29.865 3.66 30.185 3.98 ;
      RECT 29.84 3.655 30.13 3.885 ;
      RECT 29.765 3.685 30.185 3.86 ;
      RECT 29.665 3.685 30.185 3.855 ;
      RECT 29.865 8.54 30.185 8.83 ;
      RECT 29.84 8.575 30.185 8.805 ;
      RECT 29.665 8.605 30.185 8.775 ;
      RECT 26.5 3.76 26.685 3.97 ;
      RECT 26.49 3.765 26.7 3.963 ;
      RECT 26.49 3.765 26.786 3.94 ;
      RECT 26.49 3.765 26.845 3.915 ;
      RECT 26.49 3.765 26.9 3.895 ;
      RECT 26.49 3.765 26.91 3.883 ;
      RECT 26.49 3.765 27.105 3.822 ;
      RECT 26.49 3.765 27.135 3.805 ;
      RECT 26.49 3.765 27.155 3.795 ;
      RECT 27.035 3.53 27.295 3.79 ;
      RECT 27.02 3.62 27.035 3.837 ;
      RECT 26.555 3.752 27.295 3.79 ;
      RECT 27.006 3.631 27.02 3.843 ;
      RECT 26.595 3.745 27.295 3.79 ;
      RECT 26.92 3.671 27.006 3.862 ;
      RECT 26.845 3.732 27.295 3.79 ;
      RECT 26.915 3.707 26.92 3.879 ;
      RECT 26.9 3.717 27.295 3.79 ;
      RECT 26.91 3.712 26.915 3.881 ;
      RECT 25.835 3.795 25.94 4.055 ;
      RECT 26.65 3.32 26.655 3.545 ;
      RECT 26.78 3.32 26.835 3.53 ;
      RECT 26.835 3.325 26.845 3.523 ;
      RECT 26.741 3.32 26.78 3.533 ;
      RECT 26.655 3.32 26.741 3.54 ;
      RECT 26.635 3.325 26.65 3.546 ;
      RECT 26.625 3.365 26.635 3.548 ;
      RECT 26.595 3.375 26.625 3.55 ;
      RECT 26.59 3.38 26.595 3.552 ;
      RECT 26.565 3.385 26.59 3.554 ;
      RECT 26.55 3.39 26.565 3.556 ;
      RECT 26.535 3.392 26.55 3.558 ;
      RECT 26.53 3.397 26.535 3.56 ;
      RECT 26.48 3.405 26.53 3.563 ;
      RECT 26.455 3.414 26.48 3.568 ;
      RECT 26.445 3.421 26.455 3.573 ;
      RECT 26.44 3.424 26.445 3.577 ;
      RECT 26.42 3.427 26.44 3.586 ;
      RECT 26.39 3.435 26.42 3.606 ;
      RECT 26.361 3.448 26.39 3.628 ;
      RECT 26.275 3.482 26.361 3.672 ;
      RECT 26.27 3.508 26.275 3.71 ;
      RECT 26.265 3.512 26.27 3.719 ;
      RECT 26.23 3.525 26.265 3.752 ;
      RECT 26.22 3.539 26.23 3.79 ;
      RECT 26.215 3.543 26.22 3.803 ;
      RECT 26.21 3.547 26.215 3.808 ;
      RECT 26.2 3.555 26.21 3.82 ;
      RECT 26.195 3.562 26.2 3.835 ;
      RECT 26.17 3.575 26.195 3.86 ;
      RECT 26.13 3.604 26.17 3.915 ;
      RECT 26.115 3.629 26.13 3.97 ;
      RECT 26.105 3.64 26.115 3.993 ;
      RECT 26.1 3.647 26.105 4.005 ;
      RECT 26.095 3.651 26.1 4.013 ;
      RECT 26.04 3.679 26.095 4.055 ;
      RECT 26.02 3.715 26.04 4.055 ;
      RECT 26.005 3.73 26.02 4.055 ;
      RECT 25.95 3.762 26.005 4.055 ;
      RECT 25.94 3.792 25.95 4.055 ;
      RECT 25.55 3.407 25.735 3.645 ;
      RECT 25.535 3.409 25.745 3.64 ;
      RECT 25.42 3.355 25.68 3.615 ;
      RECT 25.415 3.392 25.68 3.569 ;
      RECT 25.41 3.402 25.68 3.566 ;
      RECT 25.405 3.442 25.745 3.56 ;
      RECT 25.4 3.475 25.745 3.55 ;
      RECT 25.41 3.417 25.76 3.488 ;
      RECT 25.707 4.515 25.72 5.045 ;
      RECT 25.621 4.515 25.72 5.044 ;
      RECT 25.621 4.515 25.725 5.043 ;
      RECT 25.535 4.515 25.725 5.041 ;
      RECT 25.53 4.515 25.725 5.038 ;
      RECT 25.53 4.515 25.735 5.036 ;
      RECT 25.525 4.807 25.735 5.033 ;
      RECT 25.525 4.817 25.74 5.03 ;
      RECT 25.525 4.885 25.745 5.026 ;
      RECT 25.515 4.89 25.745 5.025 ;
      RECT 25.515 4.982 25.75 5.022 ;
      RECT 25.5 4.515 25.76 4.775 ;
      RECT 25.43 10.055 25.72 10.285 ;
      RECT 25.49 9.315 25.66 10.285 ;
      RECT 25.405 9.34 25.745 9.685 ;
      RECT 25.43 9.315 25.72 9.685 ;
      RECT 24.73 3.505 24.775 5.04 ;
      RECT 24.93 3.505 24.96 3.72 ;
      RECT 23.305 3.245 23.425 3.455 ;
      RECT 22.965 3.195 23.225 3.455 ;
      RECT 22.965 3.24 23.26 3.445 ;
      RECT 24.97 3.521 24.975 3.575 ;
      RECT 24.965 3.514 24.97 3.708 ;
      RECT 24.96 3.508 24.965 3.715 ;
      RECT 24.915 3.505 24.93 3.728 ;
      RECT 24.91 3.505 24.915 3.75 ;
      RECT 24.905 3.505 24.91 3.798 ;
      RECT 24.9 3.505 24.905 3.818 ;
      RECT 24.89 3.505 24.9 3.925 ;
      RECT 24.885 3.505 24.89 3.988 ;
      RECT 24.88 3.505 24.885 4.045 ;
      RECT 24.875 3.505 24.88 4.053 ;
      RECT 24.86 3.505 24.875 4.16 ;
      RECT 24.85 3.505 24.86 4.295 ;
      RECT 24.84 3.505 24.85 4.405 ;
      RECT 24.83 3.505 24.84 4.462 ;
      RECT 24.825 3.505 24.83 4.502 ;
      RECT 24.82 3.505 24.825 4.538 ;
      RECT 24.81 3.505 24.82 4.578 ;
      RECT 24.805 3.505 24.81 4.62 ;
      RECT 24.785 3.505 24.805 4.685 ;
      RECT 24.79 4.83 24.795 5.01 ;
      RECT 24.785 4.812 24.79 5.018 ;
      RECT 24.78 3.505 24.785 4.748 ;
      RECT 24.78 4.792 24.785 5.025 ;
      RECT 24.775 3.505 24.78 5.035 ;
      RECT 24.72 3.505 24.73 3.805 ;
      RECT 24.725 4.052 24.73 5.04 ;
      RECT 24.72 4.117 24.725 5.04 ;
      RECT 24.715 3.506 24.72 3.795 ;
      RECT 24.71 4.182 24.72 5.04 ;
      RECT 24.705 3.507 24.715 3.785 ;
      RECT 24.695 4.295 24.71 5.04 ;
      RECT 24.7 3.508 24.705 3.775 ;
      RECT 24.68 3.509 24.7 3.753 ;
      RECT 24.685 4.392 24.695 5.04 ;
      RECT 24.68 4.467 24.685 5.04 ;
      RECT 24.67 3.508 24.68 3.73 ;
      RECT 24.675 4.51 24.68 5.04 ;
      RECT 24.67 4.537 24.675 5.04 ;
      RECT 24.66 3.506 24.67 3.718 ;
      RECT 24.665 4.58 24.67 5.04 ;
      RECT 24.66 4.607 24.665 5.04 ;
      RECT 24.65 3.505 24.66 3.705 ;
      RECT 24.655 4.622 24.66 5.04 ;
      RECT 24.615 4.68 24.655 5.04 ;
      RECT 24.645 3.504 24.65 3.69 ;
      RECT 24.64 3.502 24.645 3.683 ;
      RECT 24.63 3.499 24.64 3.673 ;
      RECT 24.625 3.496 24.63 3.658 ;
      RECT 24.61 3.492 24.625 3.651 ;
      RECT 24.605 4.735 24.615 5.04 ;
      RECT 24.605 3.489 24.61 3.646 ;
      RECT 24.59 3.485 24.605 3.64 ;
      RECT 24.6 4.752 24.605 5.04 ;
      RECT 24.59 4.815 24.6 5.04 ;
      RECT 24.51 3.47 24.59 3.62 ;
      RECT 24.585 4.822 24.59 5.035 ;
      RECT 24.58 4.83 24.585 5.025 ;
      RECT 24.5 3.456 24.51 3.604 ;
      RECT 24.485 3.452 24.5 3.602 ;
      RECT 24.475 3.447 24.485 3.598 ;
      RECT 24.45 3.44 24.475 3.59 ;
      RECT 24.445 3.435 24.45 3.585 ;
      RECT 24.435 3.435 24.445 3.583 ;
      RECT 24.425 3.433 24.435 3.581 ;
      RECT 24.395 3.425 24.425 3.575 ;
      RECT 24.38 3.417 24.395 3.568 ;
      RECT 24.36 3.412 24.38 3.561 ;
      RECT 24.355 3.408 24.36 3.556 ;
      RECT 24.325 3.401 24.355 3.55 ;
      RECT 24.3 3.392 24.325 3.54 ;
      RECT 24.27 3.385 24.3 3.532 ;
      RECT 24.245 3.375 24.27 3.523 ;
      RECT 24.23 3.367 24.245 3.517 ;
      RECT 24.205 3.362 24.23 3.512 ;
      RECT 24.195 3.358 24.205 3.507 ;
      RECT 24.175 3.353 24.195 3.502 ;
      RECT 24.14 3.348 24.175 3.495 ;
      RECT 24.08 3.343 24.14 3.488 ;
      RECT 24.067 3.339 24.08 3.486 ;
      RECT 23.981 3.334 24.067 3.483 ;
      RECT 23.895 3.324 23.981 3.479 ;
      RECT 23.854 3.317 23.895 3.476 ;
      RECT 23.768 3.31 23.854 3.473 ;
      RECT 23.682 3.3 23.768 3.469 ;
      RECT 23.596 3.29 23.682 3.464 ;
      RECT 23.51 3.28 23.596 3.46 ;
      RECT 23.5 3.265 23.51 3.458 ;
      RECT 23.49 3.25 23.5 3.458 ;
      RECT 23.425 3.245 23.49 3.457 ;
      RECT 23.26 3.242 23.305 3.45 ;
      RECT 24.505 4.147 24.51 4.338 ;
      RECT 24.5 4.142 24.505 4.345 ;
      RECT 24.486 4.14 24.5 4.351 ;
      RECT 24.4 4.14 24.486 4.353 ;
      RECT 24.396 4.14 24.4 4.356 ;
      RECT 24.31 4.14 24.396 4.374 ;
      RECT 24.3 4.145 24.31 4.393 ;
      RECT 24.29 4.2 24.3 4.397 ;
      RECT 24.265 4.215 24.29 4.404 ;
      RECT 24.225 4.235 24.265 4.417 ;
      RECT 24.22 4.247 24.225 4.427 ;
      RECT 24.205 4.253 24.22 4.432 ;
      RECT 24.2 4.258 24.205 4.436 ;
      RECT 24.18 4.265 24.2 4.441 ;
      RECT 24.11 4.29 24.18 4.458 ;
      RECT 24.07 4.318 24.11 4.478 ;
      RECT 24.065 4.328 24.07 4.486 ;
      RECT 24.045 4.335 24.065 4.488 ;
      RECT 24.04 4.342 24.045 4.491 ;
      RECT 24.01 4.35 24.04 4.494 ;
      RECT 24.005 4.355 24.01 4.498 ;
      RECT 23.931 4.359 24.005 4.506 ;
      RECT 23.845 4.368 23.931 4.522 ;
      RECT 23.841 4.373 23.845 4.531 ;
      RECT 23.755 4.378 23.841 4.541 ;
      RECT 23.715 4.386 23.755 4.553 ;
      RECT 23.665 4.392 23.715 4.56 ;
      RECT 23.58 4.401 23.665 4.575 ;
      RECT 23.505 4.412 23.58 4.593 ;
      RECT 23.47 4.419 23.505 4.603 ;
      RECT 23.395 4.427 23.47 4.608 ;
      RECT 23.34 4.436 23.395 4.608 ;
      RECT 23.315 4.441 23.34 4.606 ;
      RECT 23.305 4.444 23.315 4.604 ;
      RECT 23.27 4.446 23.305 4.602 ;
      RECT 23.24 4.448 23.27 4.598 ;
      RECT 23.195 4.447 23.24 4.594 ;
      RECT 23.175 4.442 23.195 4.591 ;
      RECT 23.125 4.427 23.175 4.588 ;
      RECT 23.115 4.412 23.125 4.583 ;
      RECT 23.065 4.397 23.115 4.573 ;
      RECT 23.015 4.372 23.065 4.553 ;
      RECT 23.005 4.357 23.015 4.535 ;
      RECT 23 4.355 23.005 4.529 ;
      RECT 22.98 4.35 23 4.524 ;
      RECT 22.975 4.342 22.98 4.518 ;
      RECT 22.96 4.336 22.975 4.511 ;
      RECT 22.955 4.331 22.96 4.503 ;
      RECT 22.935 4.326 22.955 4.495 ;
      RECT 22.92 4.319 22.935 4.488 ;
      RECT 22.905 4.313 22.92 4.479 ;
      RECT 22.9 4.307 22.905 4.472 ;
      RECT 22.855 4.282 22.9 4.458 ;
      RECT 22.84 4.252 22.855 4.44 ;
      RECT 22.825 4.235 22.84 4.431 ;
      RECT 22.8 4.215 22.825 4.419 ;
      RECT 22.76 4.185 22.8 4.399 ;
      RECT 22.75 4.155 22.76 4.384 ;
      RECT 22.735 4.145 22.75 4.377 ;
      RECT 22.68 4.11 22.735 4.356 ;
      RECT 22.665 4.073 22.68 4.335 ;
      RECT 22.655 4.06 22.665 4.327 ;
      RECT 22.605 4.03 22.655 4.309 ;
      RECT 22.59 3.96 22.605 4.29 ;
      RECT 22.545 3.96 22.59 4.273 ;
      RECT 22.52 3.96 22.545 4.255 ;
      RECT 22.51 3.96 22.52 4.248 ;
      RECT 22.431 3.96 22.51 4.241 ;
      RECT 22.345 3.96 22.431 4.233 ;
      RECT 22.33 3.992 22.345 4.228 ;
      RECT 22.255 4.002 22.33 4.224 ;
      RECT 22.235 4.012 22.255 4.219 ;
      RECT 22.21 4.012 22.235 4.216 ;
      RECT 22.2 4.002 22.21 4.215 ;
      RECT 22.19 3.975 22.2 4.214 ;
      RECT 22.15 3.97 22.19 4.212 ;
      RECT 22.105 3.97 22.15 4.208 ;
      RECT 22.08 3.97 22.105 4.203 ;
      RECT 22.03 3.97 22.08 4.19 ;
      RECT 21.99 3.975 22 4.175 ;
      RECT 22 3.97 22.03 4.18 ;
      RECT 23.985 3.75 24.245 4.01 ;
      RECT 23.98 3.772 24.245 3.968 ;
      RECT 23.22 3.6 23.44 3.965 ;
      RECT 23.202 3.687 23.44 3.964 ;
      RECT 23.185 3.692 23.44 3.961 ;
      RECT 23.185 3.692 23.46 3.96 ;
      RECT 23.155 3.702 23.46 3.958 ;
      RECT 23.15 3.717 23.46 3.954 ;
      RECT 23.15 3.717 23.465 3.953 ;
      RECT 23.145 3.775 23.465 3.951 ;
      RECT 23.145 3.775 23.475 3.948 ;
      RECT 23.14 3.84 23.475 3.943 ;
      RECT 23.22 3.6 23.48 3.86 ;
      RECT 21.965 3.43 22.225 3.69 ;
      RECT 21.965 3.473 22.311 3.664 ;
      RECT 21.965 3.473 22.355 3.663 ;
      RECT 21.965 3.473 22.375 3.661 ;
      RECT 21.965 3.473 22.475 3.66 ;
      RECT 21.965 3.473 22.495 3.658 ;
      RECT 21.965 3.473 22.505 3.653 ;
      RECT 22.375 3.44 22.565 3.65 ;
      RECT 22.375 3.442 22.57 3.648 ;
      RECT 22.365 3.447 22.575 3.64 ;
      RECT 22.311 3.471 22.575 3.64 ;
      RECT 22.355 3.465 22.365 3.662 ;
      RECT 22.365 3.445 22.57 3.648 ;
      RECT 21.32 4.505 21.525 4.735 ;
      RECT 21.26 4.455 21.315 4.715 ;
      RECT 21.32 4.455 21.52 4.735 ;
      RECT 22.29 4.77 22.295 4.797 ;
      RECT 22.28 4.68 22.29 4.802 ;
      RECT 22.275 4.602 22.28 4.808 ;
      RECT 22.265 4.592 22.275 4.815 ;
      RECT 22.26 4.582 22.265 4.821 ;
      RECT 22.25 4.577 22.26 4.823 ;
      RECT 22.235 4.569 22.25 4.831 ;
      RECT 22.22 4.56 22.235 4.843 ;
      RECT 22.21 4.552 22.22 4.853 ;
      RECT 22.175 4.47 22.21 4.871 ;
      RECT 22.14 4.47 22.175 4.89 ;
      RECT 22.125 4.47 22.14 4.898 ;
      RECT 22.07 4.47 22.125 4.898 ;
      RECT 22.036 4.47 22.07 4.889 ;
      RECT 21.95 4.47 22.036 4.865 ;
      RECT 21.94 4.53 21.95 4.847 ;
      RECT 21.9 4.532 21.94 4.838 ;
      RECT 21.895 4.534 21.9 4.828 ;
      RECT 21.875 4.536 21.895 4.823 ;
      RECT 21.865 4.539 21.875 4.818 ;
      RECT 21.855 4.54 21.865 4.813 ;
      RECT 21.831 4.541 21.855 4.805 ;
      RECT 21.745 4.546 21.831 4.783 ;
      RECT 21.69 4.545 21.745 4.756 ;
      RECT 21.675 4.538 21.69 4.743 ;
      RECT 21.64 4.533 21.675 4.739 ;
      RECT 21.585 4.525 21.64 4.738 ;
      RECT 21.525 4.512 21.585 4.736 ;
      RECT 21.315 4.455 21.32 4.723 ;
      RECT 21.39 3.825 21.575 4.035 ;
      RECT 21.38 3.83 21.59 4.028 ;
      RECT 21.42 3.735 21.68 3.995 ;
      RECT 21.375 3.892 21.68 3.918 ;
      RECT 20.72 3.685 20.725 4.485 ;
      RECT 20.665 3.735 20.695 4.485 ;
      RECT 20.655 3.735 20.66 4.045 ;
      RECT 20.64 3.735 20.645 4.04 ;
      RECT 20.185 3.78 20.2 3.995 ;
      RECT 20.115 3.78 20.2 3.99 ;
      RECT 21.38 3.36 21.45 3.57 ;
      RECT 21.45 3.367 21.46 3.565 ;
      RECT 21.346 3.36 21.38 3.577 ;
      RECT 21.26 3.36 21.346 3.601 ;
      RECT 21.25 3.365 21.26 3.62 ;
      RECT 21.245 3.377 21.25 3.623 ;
      RECT 21.23 3.392 21.245 3.627 ;
      RECT 21.225 3.41 21.23 3.631 ;
      RECT 21.185 3.42 21.225 3.64 ;
      RECT 21.17 3.427 21.185 3.652 ;
      RECT 21.155 3.432 21.17 3.657 ;
      RECT 21.14 3.435 21.155 3.662 ;
      RECT 21.13 3.437 21.14 3.666 ;
      RECT 21.095 3.444 21.13 3.674 ;
      RECT 21.06 3.452 21.095 3.688 ;
      RECT 21.05 3.458 21.06 3.697 ;
      RECT 21.045 3.46 21.05 3.699 ;
      RECT 21.025 3.463 21.045 3.705 ;
      RECT 20.995 3.47 21.025 3.716 ;
      RECT 20.985 3.476 20.995 3.723 ;
      RECT 20.96 3.479 20.985 3.73 ;
      RECT 20.95 3.483 20.96 3.738 ;
      RECT 20.945 3.484 20.95 3.76 ;
      RECT 20.94 3.485 20.945 3.775 ;
      RECT 20.935 3.486 20.94 3.79 ;
      RECT 20.93 3.487 20.935 3.805 ;
      RECT 20.925 3.488 20.93 3.835 ;
      RECT 20.915 3.49 20.925 3.868 ;
      RECT 20.9 3.494 20.915 3.915 ;
      RECT 20.89 3.497 20.9 3.96 ;
      RECT 20.885 3.5 20.89 3.988 ;
      RECT 20.875 3.502 20.885 4.015 ;
      RECT 20.87 3.505 20.875 4.05 ;
      RECT 20.84 3.51 20.87 4.108 ;
      RECT 20.835 3.515 20.84 4.193 ;
      RECT 20.83 3.517 20.835 4.228 ;
      RECT 20.825 3.519 20.83 4.31 ;
      RECT 20.82 3.521 20.825 4.398 ;
      RECT 20.81 3.523 20.82 4.48 ;
      RECT 20.795 3.537 20.81 4.485 ;
      RECT 20.76 3.582 20.795 4.485 ;
      RECT 20.75 3.622 20.76 4.485 ;
      RECT 20.735 3.65 20.75 4.485 ;
      RECT 20.73 3.667 20.735 4.485 ;
      RECT 20.725 3.675 20.73 4.485 ;
      RECT 20.715 3.69 20.72 4.485 ;
      RECT 20.71 3.697 20.715 4.485 ;
      RECT 20.7 3.717 20.71 4.485 ;
      RECT 20.695 3.73 20.7 4.485 ;
      RECT 20.66 3.735 20.665 4.07 ;
      RECT 20.645 4.125 20.665 4.485 ;
      RECT 20.645 3.735 20.655 4.043 ;
      RECT 20.64 4.165 20.645 4.485 ;
      RECT 20.59 3.735 20.64 4.038 ;
      RECT 20.635 4.202 20.64 4.485 ;
      RECT 20.625 4.225 20.635 4.485 ;
      RECT 20.62 4.27 20.625 4.485 ;
      RECT 20.61 4.28 20.62 4.478 ;
      RECT 20.536 3.735 20.59 4.032 ;
      RECT 20.45 3.735 20.536 4.025 ;
      RECT 20.401 3.782 20.45 4.018 ;
      RECT 20.315 3.79 20.401 4.011 ;
      RECT 20.3 3.787 20.315 4.006 ;
      RECT 20.286 3.78 20.3 4.005 ;
      RECT 20.2 3.78 20.286 4 ;
      RECT 20.105 3.785 20.115 3.985 ;
      RECT 19.695 3.215 19.71 3.615 ;
      RECT 19.89 3.215 19.895 3.475 ;
      RECT 19.635 3.215 19.68 3.475 ;
      RECT 20.09 4.52 20.095 4.725 ;
      RECT 20.085 4.51 20.09 4.73 ;
      RECT 20.08 4.497 20.085 4.735 ;
      RECT 20.075 4.477 20.08 4.735 ;
      RECT 20.05 4.43 20.075 4.735 ;
      RECT 20.015 4.345 20.05 4.735 ;
      RECT 20.01 4.282 20.015 4.735 ;
      RECT 20.005 4.267 20.01 4.735 ;
      RECT 19.99 4.227 20.005 4.735 ;
      RECT 19.985 4.202 19.99 4.735 ;
      RECT 19.975 4.185 19.985 4.735 ;
      RECT 19.94 4.107 19.975 4.735 ;
      RECT 19.935 4.05 19.94 4.735 ;
      RECT 19.93 4.037 19.935 4.735 ;
      RECT 19.92 4.015 19.93 4.735 ;
      RECT 19.91 3.98 19.92 4.735 ;
      RECT 19.9 3.95 19.91 4.735 ;
      RECT 19.89 3.865 19.9 4.378 ;
      RECT 19.897 4.51 19.9 4.735 ;
      RECT 19.895 4.52 19.897 4.735 ;
      RECT 19.885 4.53 19.895 4.73 ;
      RECT 19.88 3.215 19.89 3.61 ;
      RECT 19.885 3.742 19.89 4.353 ;
      RECT 19.88 3.64 19.885 4.336 ;
      RECT 19.87 3.215 19.88 4.312 ;
      RECT 19.865 3.215 19.87 4.283 ;
      RECT 19.86 3.215 19.865 4.273 ;
      RECT 19.84 3.215 19.86 4.235 ;
      RECT 19.835 3.215 19.84 4.193 ;
      RECT 19.83 3.215 19.835 4.173 ;
      RECT 19.8 3.215 19.83 4.123 ;
      RECT 19.79 3.215 19.8 4.07 ;
      RECT 19.785 3.215 19.79 4.043 ;
      RECT 19.78 3.215 19.785 4.028 ;
      RECT 19.77 3.215 19.78 4.005 ;
      RECT 19.76 3.215 19.77 3.98 ;
      RECT 19.755 3.215 19.76 3.92 ;
      RECT 19.745 3.215 19.755 3.858 ;
      RECT 19.74 3.215 19.745 3.778 ;
      RECT 19.735 3.215 19.74 3.743 ;
      RECT 19.73 3.215 19.735 3.718 ;
      RECT 19.725 3.215 19.73 3.703 ;
      RECT 19.72 3.215 19.725 3.673 ;
      RECT 19.715 3.215 19.72 3.65 ;
      RECT 19.71 3.215 19.715 3.623 ;
      RECT 19.68 3.215 19.695 3.61 ;
      RECT 18.835 4.75 19.02 4.96 ;
      RECT 18.825 4.755 19.035 4.953 ;
      RECT 18.825 4.755 19.055 4.925 ;
      RECT 18.825 4.755 19.07 4.904 ;
      RECT 18.825 4.755 19.085 4.902 ;
      RECT 18.825 4.755 19.095 4.901 ;
      RECT 18.825 4.755 19.125 4.898 ;
      RECT 19.475 4.6 19.735 4.86 ;
      RECT 19.435 4.647 19.735 4.843 ;
      RECT 19.426 4.655 19.435 4.846 ;
      RECT 19.02 4.748 19.735 4.843 ;
      RECT 19.34 4.673 19.426 4.853 ;
      RECT 19.035 4.745 19.735 4.843 ;
      RECT 19.281 4.695 19.34 4.865 ;
      RECT 19.055 4.741 19.735 4.843 ;
      RECT 19.195 4.707 19.281 4.876 ;
      RECT 19.07 4.737 19.735 4.843 ;
      RECT 19.14 4.72 19.195 4.888 ;
      RECT 19.085 4.735 19.735 4.843 ;
      RECT 19.125 4.726 19.14 4.894 ;
      RECT 19.095 4.731 19.735 4.843 ;
      RECT 19.24 4.255 19.5 4.515 ;
      RECT 19.24 4.275 19.61 4.485 ;
      RECT 19.24 4.28 19.62 4.48 ;
      RECT 19.431 3.694 19.51 3.925 ;
      RECT 19.345 3.697 19.56 3.92 ;
      RECT 19.34 3.697 19.56 3.915 ;
      RECT 19.34 3.702 19.57 3.913 ;
      RECT 19.315 3.702 19.57 3.91 ;
      RECT 19.315 3.71 19.58 3.908 ;
      RECT 19.195 3.645 19.455 3.905 ;
      RECT 19.195 3.692 19.505 3.905 ;
      RECT 18.45 4.265 18.455 4.525 ;
      RECT 18.28 4.035 18.285 4.525 ;
      RECT 18.165 4.275 18.17 4.5 ;
      RECT 18.875 3.37 18.88 3.58 ;
      RECT 18.88 3.375 18.895 3.575 ;
      RECT 18.815 3.37 18.875 3.588 ;
      RECT 18.8 3.37 18.815 3.598 ;
      RECT 18.75 3.37 18.8 3.615 ;
      RECT 18.73 3.37 18.75 3.638 ;
      RECT 18.715 3.37 18.73 3.65 ;
      RECT 18.695 3.37 18.715 3.66 ;
      RECT 18.685 3.375 18.695 3.669 ;
      RECT 18.68 3.385 18.685 3.674 ;
      RECT 18.675 3.397 18.68 3.678 ;
      RECT 18.665 3.42 18.675 3.683 ;
      RECT 18.66 3.435 18.665 3.687 ;
      RECT 18.655 3.452 18.66 3.69 ;
      RECT 18.65 3.46 18.655 3.693 ;
      RECT 18.64 3.465 18.65 3.697 ;
      RECT 18.635 3.472 18.64 3.702 ;
      RECT 18.625 3.477 18.635 3.706 ;
      RECT 18.6 3.489 18.625 3.717 ;
      RECT 18.58 3.506 18.6 3.733 ;
      RECT 18.555 3.523 18.58 3.755 ;
      RECT 18.52 3.546 18.555 3.813 ;
      RECT 18.5 3.568 18.52 3.875 ;
      RECT 18.495 3.578 18.5 3.91 ;
      RECT 18.485 3.585 18.495 3.948 ;
      RECT 18.48 3.592 18.485 3.968 ;
      RECT 18.475 3.603 18.48 4.005 ;
      RECT 18.47 3.611 18.475 4.07 ;
      RECT 18.46 3.622 18.47 4.123 ;
      RECT 18.455 3.64 18.46 4.193 ;
      RECT 18.45 3.65 18.455 4.23 ;
      RECT 18.445 3.66 18.45 4.525 ;
      RECT 18.44 3.672 18.445 4.525 ;
      RECT 18.435 3.682 18.44 4.525 ;
      RECT 18.425 3.692 18.435 4.525 ;
      RECT 18.415 3.715 18.425 4.525 ;
      RECT 18.4 3.75 18.415 4.525 ;
      RECT 18.36 3.812 18.4 4.525 ;
      RECT 18.355 3.865 18.36 4.525 ;
      RECT 18.33 3.9 18.355 4.525 ;
      RECT 18.315 3.945 18.33 4.525 ;
      RECT 18.31 3.967 18.315 4.525 ;
      RECT 18.3 3.98 18.31 4.525 ;
      RECT 18.29 4.005 18.3 4.525 ;
      RECT 18.285 4.027 18.29 4.525 ;
      RECT 18.26 4.065 18.28 4.525 ;
      RECT 18.22 4.122 18.26 4.525 ;
      RECT 18.215 4.172 18.22 4.525 ;
      RECT 18.21 4.19 18.215 4.525 ;
      RECT 18.205 4.202 18.21 4.525 ;
      RECT 18.195 4.22 18.205 4.525 ;
      RECT 18.185 4.24 18.195 4.5 ;
      RECT 18.18 4.257 18.185 4.5 ;
      RECT 18.17 4.27 18.18 4.5 ;
      RECT 18.14 4.28 18.165 4.5 ;
      RECT 18.13 4.287 18.14 4.5 ;
      RECT 18.115 4.297 18.13 4.495 ;
      RECT 16.54 10.055 16.83 10.285 ;
      RECT 16.6 9.31 16.77 10.285 ;
      RECT 16.51 9.31 16.86 9.6 ;
      RECT 16.135 8.57 16.485 8.86 ;
      RECT 15.995 8.605 16.485 8.775 ;
      RECT 91.005 4.145 91.375 4.515 ;
      RECT 75.22 4.145 75.59 4.515 ;
      RECT 59.435 4.145 59.805 4.515 ;
      RECT 43.66 4.145 44.03 4.515 ;
      RECT 27.88 4.145 28.25 4.515 ;
    LAYER mcon ;
      RECT 96.185 7.3 96.355 7.47 ;
      RECT 96.18 8.6 96.35 8.77 ;
      RECT 96.18 10.08 96.35 10.25 ;
      RECT 95.81 8.23 95.98 8.4 ;
      RECT 95.805 4.06 95.975 4.23 ;
      RECT 95.185 2.205 95.355 2.375 ;
      RECT 95.185 3.685 95.355 3.855 ;
      RECT 95.185 8.605 95.355 8.775 ;
      RECT 95.185 10.085 95.355 10.255 ;
      RECT 94.815 4.055 94.985 4.225 ;
      RECT 94.815 8.235 94.985 8.405 ;
      RECT 93.825 3.315 93.995 3.485 ;
      RECT 93.825 8.975 93.995 9.145 ;
      RECT 93.395 2.205 93.565 2.375 ;
      RECT 93.395 2.945 93.565 3.115 ;
      RECT 93.395 9.345 93.565 9.515 ;
      RECT 93.395 10.085 93.565 10.255 ;
      RECT 93.025 3.685 93.195 3.855 ;
      RECT 93.025 8.605 93.195 8.775 ;
      RECT 89.78 3.34 89.95 3.51 ;
      RECT 89.635 3.78 89.805 3.95 ;
      RECT 89.045 8.975 89.215 9.145 ;
      RECT 89.025 3.82 89.195 3.99 ;
      RECT 88.68 3.455 88.85 3.625 ;
      RECT 88.67 4.815 88.84 4.985 ;
      RECT 88.615 9.345 88.785 9.515 ;
      RECT 88.615 10.085 88.785 10.255 ;
      RECT 87.905 3.53 88.075 3.7 ;
      RECT 87.725 4.845 87.895 5.015 ;
      RECT 87.445 4.16 87.615 4.33 ;
      RECT 87.125 3.785 87.295 3.955 ;
      RECT 86.435 3.265 86.605 3.435 ;
      RECT 86.36 3.735 86.53 3.905 ;
      RECT 85.51 3.46 85.68 3.63 ;
      RECT 85.17 4.655 85.34 4.825 ;
      RECT 85.135 3.99 85.305 4.16 ;
      RECT 84.525 3.845 84.695 4.015 ;
      RECT 84.455 4.545 84.625 4.715 ;
      RECT 84.395 3.38 84.565 3.55 ;
      RECT 83.755 4.295 83.925 4.465 ;
      RECT 83.25 3.8 83.42 3.97 ;
      RECT 83.03 4.545 83.2 4.715 ;
      RECT 82.825 3.425 82.995 3.595 ;
      RECT 82.555 4.295 82.725 4.465 ;
      RECT 82.515 3.725 82.685 3.895 ;
      RECT 81.97 4.77 82.14 4.94 ;
      RECT 81.83 3.39 82 3.56 ;
      RECT 81.26 4.31 81.43 4.48 ;
      RECT 80.4 7.3 80.57 7.47 ;
      RECT 80.395 8.6 80.565 8.77 ;
      RECT 80.395 10.08 80.565 10.25 ;
      RECT 80.025 8.23 80.195 8.4 ;
      RECT 80.02 4.06 80.19 4.23 ;
      RECT 79.4 2.205 79.57 2.375 ;
      RECT 79.4 3.685 79.57 3.855 ;
      RECT 79.4 8.605 79.57 8.775 ;
      RECT 79.4 10.085 79.57 10.255 ;
      RECT 79.03 4.055 79.2 4.225 ;
      RECT 79.03 8.235 79.2 8.405 ;
      RECT 78.04 3.315 78.21 3.485 ;
      RECT 78.04 8.975 78.21 9.145 ;
      RECT 77.61 2.205 77.78 2.375 ;
      RECT 77.61 2.945 77.78 3.115 ;
      RECT 77.61 9.345 77.78 9.515 ;
      RECT 77.61 10.085 77.78 10.255 ;
      RECT 77.24 3.685 77.41 3.855 ;
      RECT 77.24 8.605 77.41 8.775 ;
      RECT 73.995 3.34 74.165 3.51 ;
      RECT 73.85 3.78 74.02 3.95 ;
      RECT 73.26 8.975 73.43 9.145 ;
      RECT 73.24 3.82 73.41 3.99 ;
      RECT 72.895 3.455 73.065 3.625 ;
      RECT 72.885 4.815 73.055 4.985 ;
      RECT 72.83 9.345 73 9.515 ;
      RECT 72.83 10.085 73 10.255 ;
      RECT 72.12 3.53 72.29 3.7 ;
      RECT 71.94 4.845 72.11 5.015 ;
      RECT 71.66 4.16 71.83 4.33 ;
      RECT 71.34 3.785 71.51 3.955 ;
      RECT 70.65 3.265 70.82 3.435 ;
      RECT 70.575 3.735 70.745 3.905 ;
      RECT 69.725 3.46 69.895 3.63 ;
      RECT 69.385 4.655 69.555 4.825 ;
      RECT 69.35 3.99 69.52 4.16 ;
      RECT 68.74 3.845 68.91 4.015 ;
      RECT 68.67 4.545 68.84 4.715 ;
      RECT 68.61 3.38 68.78 3.55 ;
      RECT 67.97 4.295 68.14 4.465 ;
      RECT 67.465 3.8 67.635 3.97 ;
      RECT 67.245 4.545 67.415 4.715 ;
      RECT 67.04 3.425 67.21 3.595 ;
      RECT 66.77 4.295 66.94 4.465 ;
      RECT 66.73 3.725 66.9 3.895 ;
      RECT 66.185 4.77 66.355 4.94 ;
      RECT 66.045 3.39 66.215 3.56 ;
      RECT 65.475 4.31 65.645 4.48 ;
      RECT 64.615 7.3 64.785 7.47 ;
      RECT 64.61 8.6 64.78 8.77 ;
      RECT 64.61 10.08 64.78 10.25 ;
      RECT 64.24 8.23 64.41 8.4 ;
      RECT 64.235 4.06 64.405 4.23 ;
      RECT 63.615 2.205 63.785 2.375 ;
      RECT 63.615 3.685 63.785 3.855 ;
      RECT 63.615 8.605 63.785 8.775 ;
      RECT 63.615 10.085 63.785 10.255 ;
      RECT 63.245 4.055 63.415 4.225 ;
      RECT 63.245 8.235 63.415 8.405 ;
      RECT 62.255 3.315 62.425 3.485 ;
      RECT 62.255 8.975 62.425 9.145 ;
      RECT 61.825 2.205 61.995 2.375 ;
      RECT 61.825 2.945 61.995 3.115 ;
      RECT 61.825 9.345 61.995 9.515 ;
      RECT 61.825 10.085 61.995 10.255 ;
      RECT 61.455 3.685 61.625 3.855 ;
      RECT 61.455 8.605 61.625 8.775 ;
      RECT 58.21 3.34 58.38 3.51 ;
      RECT 58.065 3.78 58.235 3.95 ;
      RECT 57.475 8.975 57.645 9.145 ;
      RECT 57.455 3.82 57.625 3.99 ;
      RECT 57.11 3.455 57.28 3.625 ;
      RECT 57.1 4.815 57.27 4.985 ;
      RECT 57.045 9.345 57.215 9.515 ;
      RECT 57.045 10.085 57.215 10.255 ;
      RECT 56.335 3.53 56.505 3.7 ;
      RECT 56.155 4.845 56.325 5.015 ;
      RECT 55.875 4.16 56.045 4.33 ;
      RECT 55.555 3.785 55.725 3.955 ;
      RECT 54.865 3.265 55.035 3.435 ;
      RECT 54.79 3.735 54.96 3.905 ;
      RECT 53.94 3.46 54.11 3.63 ;
      RECT 53.6 4.655 53.77 4.825 ;
      RECT 53.565 3.99 53.735 4.16 ;
      RECT 52.955 3.845 53.125 4.015 ;
      RECT 52.885 4.545 53.055 4.715 ;
      RECT 52.825 3.38 52.995 3.55 ;
      RECT 52.185 4.295 52.355 4.465 ;
      RECT 51.68 3.8 51.85 3.97 ;
      RECT 51.46 4.545 51.63 4.715 ;
      RECT 51.255 3.425 51.425 3.595 ;
      RECT 50.985 4.295 51.155 4.465 ;
      RECT 50.945 3.725 51.115 3.895 ;
      RECT 50.4 4.77 50.57 4.94 ;
      RECT 50.26 3.39 50.43 3.56 ;
      RECT 49.69 4.31 49.86 4.48 ;
      RECT 48.84 7.3 49.01 7.47 ;
      RECT 48.835 8.6 49.005 8.77 ;
      RECT 48.835 10.08 49.005 10.25 ;
      RECT 48.465 8.23 48.635 8.4 ;
      RECT 48.46 4.06 48.63 4.23 ;
      RECT 47.84 2.205 48.01 2.375 ;
      RECT 47.84 3.685 48.01 3.855 ;
      RECT 47.84 8.605 48.01 8.775 ;
      RECT 47.84 10.085 48.01 10.255 ;
      RECT 47.47 4.055 47.64 4.225 ;
      RECT 47.47 8.235 47.64 8.405 ;
      RECT 46.48 3.315 46.65 3.485 ;
      RECT 46.48 8.975 46.65 9.145 ;
      RECT 46.05 2.205 46.22 2.375 ;
      RECT 46.05 2.945 46.22 3.115 ;
      RECT 46.05 9.345 46.22 9.515 ;
      RECT 46.05 10.085 46.22 10.255 ;
      RECT 45.68 3.685 45.85 3.855 ;
      RECT 45.68 8.605 45.85 8.775 ;
      RECT 42.435 3.34 42.605 3.51 ;
      RECT 42.29 3.78 42.46 3.95 ;
      RECT 41.7 8.975 41.87 9.145 ;
      RECT 41.68 3.82 41.85 3.99 ;
      RECT 41.335 3.455 41.505 3.625 ;
      RECT 41.325 4.815 41.495 4.985 ;
      RECT 41.27 9.345 41.44 9.515 ;
      RECT 41.27 10.085 41.44 10.255 ;
      RECT 40.56 3.53 40.73 3.7 ;
      RECT 40.38 4.845 40.55 5.015 ;
      RECT 40.1 4.16 40.27 4.33 ;
      RECT 39.78 3.785 39.95 3.955 ;
      RECT 39.09 3.265 39.26 3.435 ;
      RECT 39.015 3.735 39.185 3.905 ;
      RECT 38.165 3.46 38.335 3.63 ;
      RECT 37.825 4.655 37.995 4.825 ;
      RECT 37.79 3.99 37.96 4.16 ;
      RECT 37.18 3.845 37.35 4.015 ;
      RECT 37.11 4.545 37.28 4.715 ;
      RECT 37.05 3.38 37.22 3.55 ;
      RECT 36.41 4.295 36.58 4.465 ;
      RECT 35.905 3.8 36.075 3.97 ;
      RECT 35.685 4.545 35.855 4.715 ;
      RECT 35.48 3.425 35.65 3.595 ;
      RECT 35.21 4.295 35.38 4.465 ;
      RECT 35.17 3.725 35.34 3.895 ;
      RECT 34.625 4.77 34.795 4.94 ;
      RECT 34.485 3.39 34.655 3.56 ;
      RECT 33.915 4.31 34.085 4.48 ;
      RECT 33.06 7.3 33.23 7.47 ;
      RECT 33.055 8.6 33.225 8.77 ;
      RECT 33.055 10.08 33.225 10.25 ;
      RECT 32.685 8.23 32.855 8.4 ;
      RECT 32.68 4.06 32.85 4.23 ;
      RECT 32.06 2.205 32.23 2.375 ;
      RECT 32.06 3.685 32.23 3.855 ;
      RECT 32.06 8.605 32.23 8.775 ;
      RECT 32.06 10.085 32.23 10.255 ;
      RECT 31.69 4.055 31.86 4.225 ;
      RECT 31.69 8.235 31.86 8.405 ;
      RECT 30.7 3.315 30.87 3.485 ;
      RECT 30.7 8.975 30.87 9.145 ;
      RECT 30.27 2.205 30.44 2.375 ;
      RECT 30.27 2.945 30.44 3.115 ;
      RECT 30.27 9.345 30.44 9.515 ;
      RECT 30.27 10.085 30.44 10.255 ;
      RECT 29.9 3.685 30.07 3.855 ;
      RECT 29.9 8.605 30.07 8.775 ;
      RECT 26.655 3.34 26.825 3.51 ;
      RECT 26.51 3.78 26.68 3.95 ;
      RECT 25.92 8.975 26.09 9.145 ;
      RECT 25.9 3.82 26.07 3.99 ;
      RECT 25.555 3.455 25.725 3.625 ;
      RECT 25.545 4.815 25.715 4.985 ;
      RECT 25.49 9.345 25.66 9.515 ;
      RECT 25.49 10.085 25.66 10.255 ;
      RECT 24.78 3.53 24.95 3.7 ;
      RECT 24.6 4.845 24.77 5.015 ;
      RECT 24.32 4.16 24.49 4.33 ;
      RECT 24 3.785 24.17 3.955 ;
      RECT 23.31 3.265 23.48 3.435 ;
      RECT 23.235 3.735 23.405 3.905 ;
      RECT 22.385 3.46 22.555 3.63 ;
      RECT 22.045 4.655 22.215 4.825 ;
      RECT 22.01 3.99 22.18 4.16 ;
      RECT 21.4 3.845 21.57 4.015 ;
      RECT 21.33 4.545 21.5 4.715 ;
      RECT 21.27 3.38 21.44 3.55 ;
      RECT 20.63 4.295 20.8 4.465 ;
      RECT 20.125 3.8 20.295 3.97 ;
      RECT 19.905 4.545 20.075 4.715 ;
      RECT 19.7 3.425 19.87 3.595 ;
      RECT 19.43 4.295 19.6 4.465 ;
      RECT 19.39 3.725 19.56 3.895 ;
      RECT 18.845 4.77 19.015 4.94 ;
      RECT 18.705 3.39 18.875 3.56 ;
      RECT 18.135 4.31 18.305 4.48 ;
      RECT 16.6 9.345 16.77 9.515 ;
      RECT 16.6 10.085 16.77 10.255 ;
      RECT 16.23 8.605 16.4 8.775 ;
    LAYER li1 ;
      RECT 96.18 7.3 96.35 8.77 ;
      RECT 96.18 7.3 96.355 8.56 ;
      RECT 95.81 9.25 96.28 9.42 ;
      RECT 95.81 8.23 95.98 9.42 ;
      RECT 95.805 3.04 95.975 4.23 ;
      RECT 95.805 3.04 96.275 3.21 ;
      RECT 95.185 3.895 95.36 5.155 ;
      RECT 95.185 3.685 95.355 5.155 ;
      RECT 95.185 7.305 95.355 8.775 ;
      RECT 95.185 7.305 95.36 8.565 ;
      RECT 94.815 3.035 94.985 4.225 ;
      RECT 94.815 3.035 95.285 3.205 ;
      RECT 94.815 9.255 95.285 9.425 ;
      RECT 94.815 8.235 94.985 9.425 ;
      RECT 93.825 4.015 94 5.155 ;
      RECT 93.825 1.865 93.995 5.155 ;
      RECT 93.825 1.865 94 2.415 ;
      RECT 93.825 10.045 94 10.595 ;
      RECT 93.825 7.305 93.995 10.595 ;
      RECT 93.825 7.305 94 8.445 ;
      RECT 93.395 3.895 93.57 5.155 ;
      RECT 93.395 2.945 93.565 5.155 ;
      RECT 93.395 7.305 93.565 9.515 ;
      RECT 93.395 7.305 93.57 8.565 ;
      RECT 92.965 3.925 93.135 5.155 ;
      RECT 93.025 2.145 93.195 4.095 ;
      RECT 92.965 1.865 93.135 2.315 ;
      RECT 92.965 10.145 93.135 10.595 ;
      RECT 93.025 8.365 93.195 10.315 ;
      RECT 92.965 7.305 93.135 8.535 ;
      RECT 92.44 3.895 92.615 5.155 ;
      RECT 92.44 1.865 92.61 5.155 ;
      RECT 92.44 3.365 92.85 3.695 ;
      RECT 92.44 2.525 92.85 2.855 ;
      RECT 92.44 1.865 92.615 2.355 ;
      RECT 92.44 10.105 92.615 10.595 ;
      RECT 92.44 7.305 92.61 10.595 ;
      RECT 92.44 9.605 92.85 9.935 ;
      RECT 92.44 8.765 92.85 9.095 ;
      RECT 92.44 7.305 92.615 8.565 ;
      RECT 89.78 3.27 90.51 3.51 ;
      RECT 90.322 3.065 90.51 3.51 ;
      RECT 90.15 3.077 90.525 3.504 ;
      RECT 90.065 3.092 90.545 3.489 ;
      RECT 90.065 3.107 90.55 3.479 ;
      RECT 90.02 3.127 90.565 3.471 ;
      RECT 89.997 3.162 90.58 3.425 ;
      RECT 89.911 3.185 90.585 3.385 ;
      RECT 89.911 3.203 90.595 3.355 ;
      RECT 89.78 3.272 90.6 3.318 ;
      RECT 89.825 3.215 90.595 3.355 ;
      RECT 89.911 3.167 90.58 3.425 ;
      RECT 89.997 3.136 90.565 3.471 ;
      RECT 90.02 3.117 90.55 3.479 ;
      RECT 90.065 3.09 90.525 3.504 ;
      RECT 90.15 3.072 90.51 3.51 ;
      RECT 90.236 3.066 90.51 3.51 ;
      RECT 90.322 3.061 90.455 3.51 ;
      RECT 90.408 3.056 90.455 3.51 ;
      RECT 89.97 4.67 89.975 4.683 ;
      RECT 89.965 4.565 89.97 4.688 ;
      RECT 89.94 4.425 89.965 4.703 ;
      RECT 89.905 4.376 89.94 4.735 ;
      RECT 89.9 4.344 89.905 4.755 ;
      RECT 89.895 4.335 89.9 4.755 ;
      RECT 89.815 4.3 89.895 4.755 ;
      RECT 89.752 4.27 89.815 4.755 ;
      RECT 89.666 4.258 89.752 4.755 ;
      RECT 89.58 4.244 89.666 4.755 ;
      RECT 89.5 4.231 89.58 4.741 ;
      RECT 89.465 4.223 89.5 4.721 ;
      RECT 89.455 4.22 89.465 4.712 ;
      RECT 89.425 4.215 89.455 4.699 ;
      RECT 89.375 4.19 89.425 4.675 ;
      RECT 89.361 4.164 89.375 4.657 ;
      RECT 89.275 4.124 89.361 4.633 ;
      RECT 89.23 4.072 89.275 4.602 ;
      RECT 89.22 4.047 89.23 4.589 ;
      RECT 89.215 3.828 89.22 3.85 ;
      RECT 89.21 4.03 89.22 4.585 ;
      RECT 89.21 3.826 89.215 3.94 ;
      RECT 89.2 3.822 89.21 4.581 ;
      RECT 89.156 3.82 89.2 4.569 ;
      RECT 89.07 3.82 89.156 4.54 ;
      RECT 89.04 3.82 89.07 4.513 ;
      RECT 89.025 3.82 89.04 4.501 ;
      RECT 88.985 3.832 89.025 4.486 ;
      RECT 88.965 3.851 88.985 4.465 ;
      RECT 88.955 3.861 88.965 4.449 ;
      RECT 88.945 3.867 88.955 4.438 ;
      RECT 88.925 3.877 88.945 4.421 ;
      RECT 88.92 3.886 88.925 4.408 ;
      RECT 88.915 3.89 88.92 4.358 ;
      RECT 88.905 3.896 88.915 4.275 ;
      RECT 88.9 3.9 88.905 4.189 ;
      RECT 88.895 3.92 88.9 4.126 ;
      RECT 88.89 3.943 88.895 4.073 ;
      RECT 88.885 3.961 88.89 4.018 ;
      RECT 89.495 3.78 89.665 4.04 ;
      RECT 89.665 3.745 89.71 4.026 ;
      RECT 89.626 3.747 89.715 4.009 ;
      RECT 89.515 3.764 89.801 3.98 ;
      RECT 89.515 3.779 89.805 3.952 ;
      RECT 89.515 3.76 89.715 4.009 ;
      RECT 89.54 3.748 89.665 4.04 ;
      RECT 89.626 3.746 89.71 4.026 ;
      RECT 89.045 10.045 89.22 10.595 ;
      RECT 89.045 7.305 89.215 10.595 ;
      RECT 89.045 7.305 89.22 8.445 ;
      RECT 88.68 3.135 88.85 3.625 ;
      RECT 88.68 3.135 88.885 3.605 ;
      RECT 88.815 3.055 88.925 3.565 ;
      RECT 88.796 3.059 88.945 3.535 ;
      RECT 88.71 3.067 88.965 3.518 ;
      RECT 88.71 3.073 88.97 3.508 ;
      RECT 88.71 3.082 88.99 3.496 ;
      RECT 88.685 3.107 89.02 3.474 ;
      RECT 88.685 3.127 89.025 3.454 ;
      RECT 88.68 3.14 89.035 3.434 ;
      RECT 88.68 3.207 89.04 3.415 ;
      RECT 88.68 3.34 89.045 3.402 ;
      RECT 88.675 3.145 89.035 3.235 ;
      RECT 88.685 3.102 88.99 3.496 ;
      RECT 88.796 3.057 88.925 3.565 ;
      RECT 88.67 4.81 88.97 5.065 ;
      RECT 88.755 4.776 88.97 5.065 ;
      RECT 88.755 4.779 88.975 4.925 ;
      RECT 88.69 4.8 88.975 4.925 ;
      RECT 88.725 4.79 88.97 5.065 ;
      RECT 88.72 4.795 88.975 4.925 ;
      RECT 88.755 4.774 88.956 5.065 ;
      RECT 88.841 4.765 88.956 5.065 ;
      RECT 88.841 4.759 88.87 5.065 ;
      RECT 88.615 7.305 88.785 9.515 ;
      RECT 88.615 7.305 88.79 8.565 ;
      RECT 88.33 4.4 88.34 4.89 ;
      RECT 87.99 4.335 88 4.635 ;
      RECT 88.505 4.507 88.51 4.726 ;
      RECT 88.495 4.487 88.505 4.743 ;
      RECT 88.485 4.467 88.495 4.773 ;
      RECT 88.48 4.457 88.485 4.788 ;
      RECT 88.475 4.453 88.48 4.793 ;
      RECT 88.46 4.445 88.475 4.8 ;
      RECT 88.42 4.425 88.46 4.825 ;
      RECT 88.395 4.407 88.42 4.858 ;
      RECT 88.39 4.405 88.395 4.871 ;
      RECT 88.37 4.402 88.39 4.875 ;
      RECT 88.34 4.4 88.37 4.885 ;
      RECT 88.27 4.402 88.33 4.886 ;
      RECT 88.25 4.402 88.27 4.88 ;
      RECT 88.225 4.4 88.25 4.877 ;
      RECT 88.19 4.395 88.225 4.873 ;
      RECT 88.17 4.389 88.19 4.86 ;
      RECT 88.16 4.386 88.17 4.848 ;
      RECT 88.14 4.383 88.16 4.833 ;
      RECT 88.12 4.379 88.14 4.815 ;
      RECT 88.115 4.376 88.12 4.805 ;
      RECT 88.11 4.375 88.115 4.803 ;
      RECT 88.1 4.372 88.11 4.795 ;
      RECT 88.09 4.366 88.1 4.778 ;
      RECT 88.08 4.36 88.09 4.76 ;
      RECT 88.07 4.354 88.08 4.748 ;
      RECT 88.06 4.348 88.07 4.728 ;
      RECT 88.055 4.344 88.06 4.713 ;
      RECT 88.05 4.342 88.055 4.705 ;
      RECT 88.045 4.34 88.05 4.698 ;
      RECT 88.04 4.338 88.045 4.688 ;
      RECT 88.035 4.336 88.04 4.682 ;
      RECT 88.025 4.335 88.035 4.672 ;
      RECT 88.015 4.335 88.025 4.663 ;
      RECT 88 4.335 88.015 4.648 ;
      RECT 87.96 4.335 87.99 4.632 ;
      RECT 87.94 4.337 87.96 4.627 ;
      RECT 87.935 4.342 87.94 4.625 ;
      RECT 87.905 4.35 87.935 4.623 ;
      RECT 87.875 4.365 87.905 4.622 ;
      RECT 87.83 4.387 87.875 4.627 ;
      RECT 87.825 4.402 87.83 4.631 ;
      RECT 87.81 4.407 87.825 4.633 ;
      RECT 87.805 4.411 87.81 4.635 ;
      RECT 87.745 4.434 87.805 4.644 ;
      RECT 87.725 4.46 87.745 4.657 ;
      RECT 87.715 4.467 87.725 4.661 ;
      RECT 87.7 4.474 87.715 4.664 ;
      RECT 87.68 4.484 87.7 4.667 ;
      RECT 87.675 4.492 87.68 4.67 ;
      RECT 87.63 4.497 87.675 4.677 ;
      RECT 87.62 4.5 87.63 4.684 ;
      RECT 87.61 4.5 87.62 4.688 ;
      RECT 87.575 4.502 87.61 4.7 ;
      RECT 87.555 4.505 87.575 4.713 ;
      RECT 87.515 4.508 87.555 4.724 ;
      RECT 87.5 4.51 87.515 4.737 ;
      RECT 87.49 4.51 87.5 4.742 ;
      RECT 87.465 4.511 87.49 4.75 ;
      RECT 87.455 4.513 87.465 4.755 ;
      RECT 87.45 4.514 87.455 4.758 ;
      RECT 87.425 4.512 87.45 4.761 ;
      RECT 87.41 4.51 87.425 4.762 ;
      RECT 87.39 4.507 87.41 4.764 ;
      RECT 87.37 4.502 87.39 4.764 ;
      RECT 87.31 4.497 87.37 4.761 ;
      RECT 87.275 4.472 87.31 4.757 ;
      RECT 87.265 4.449 87.275 4.755 ;
      RECT 87.235 4.426 87.265 4.755 ;
      RECT 87.225 4.405 87.235 4.755 ;
      RECT 87.2 4.387 87.225 4.753 ;
      RECT 87.185 4.365 87.2 4.75 ;
      RECT 87.17 4.347 87.185 4.748 ;
      RECT 87.15 4.337 87.17 4.746 ;
      RECT 87.135 4.332 87.15 4.745 ;
      RECT 87.12 4.33 87.135 4.744 ;
      RECT 87.09 4.331 87.12 4.742 ;
      RECT 87.07 4.334 87.09 4.74 ;
      RECT 87.013 4.338 87.07 4.74 ;
      RECT 86.927 4.347 87.013 4.74 ;
      RECT 86.841 4.358 86.927 4.74 ;
      RECT 86.755 4.369 86.841 4.74 ;
      RECT 86.735 4.376 86.755 4.748 ;
      RECT 86.725 4.379 86.735 4.755 ;
      RECT 86.66 4.384 86.725 4.773 ;
      RECT 86.63 4.391 86.66 4.798 ;
      RECT 86.62 4.394 86.63 4.805 ;
      RECT 86.575 4.398 86.62 4.81 ;
      RECT 86.545 4.403 86.575 4.815 ;
      RECT 86.544 4.405 86.545 4.815 ;
      RECT 86.458 4.411 86.544 4.815 ;
      RECT 86.372 4.422 86.458 4.815 ;
      RECT 86.286 4.434 86.372 4.815 ;
      RECT 86.2 4.445 86.286 4.815 ;
      RECT 86.185 4.452 86.2 4.81 ;
      RECT 86.18 4.454 86.185 4.804 ;
      RECT 86.16 4.465 86.18 4.799 ;
      RECT 86.15 4.483 86.16 4.793 ;
      RECT 86.145 4.495 86.15 4.593 ;
      RECT 88.44 3.248 88.46 3.335 ;
      RECT 88.435 3.183 88.44 3.367 ;
      RECT 88.425 3.15 88.435 3.372 ;
      RECT 88.42 3.13 88.425 3.378 ;
      RECT 88.39 3.13 88.42 3.395 ;
      RECT 88.341 3.13 88.39 3.431 ;
      RECT 88.255 3.13 88.341 3.489 ;
      RECT 88.226 3.14 88.255 3.538 ;
      RECT 88.14 3.182 88.226 3.591 ;
      RECT 88.12 3.22 88.14 3.638 ;
      RECT 88.095 3.237 88.12 3.658 ;
      RECT 88.085 3.251 88.095 3.678 ;
      RECT 88.08 3.257 88.085 3.688 ;
      RECT 88.075 3.261 88.08 3.695 ;
      RECT 88.025 3.281 88.075 3.7 ;
      RECT 87.96 3.325 88.025 3.7 ;
      RECT 87.935 3.375 87.96 3.7 ;
      RECT 87.925 3.405 87.935 3.7 ;
      RECT 87.92 3.432 87.925 3.7 ;
      RECT 87.915 3.45 87.92 3.7 ;
      RECT 87.905 3.492 87.915 3.7 ;
      RECT 87.66 10.105 87.835 10.595 ;
      RECT 87.66 7.305 87.83 10.595 ;
      RECT 87.66 9.605 88.07 9.935 ;
      RECT 87.66 8.765 88.07 9.095 ;
      RECT 87.66 7.305 87.835 8.565 ;
      RECT 87.735 4.85 87.925 5.075 ;
      RECT 87.725 4.851 87.93 5.07 ;
      RECT 87.725 4.853 87.94 5.05 ;
      RECT 87.725 4.857 87.945 5.035 ;
      RECT 87.725 4.844 87.895 5.07 ;
      RECT 87.725 4.847 87.92 5.07 ;
      RECT 87.735 4.843 87.895 5.075 ;
      RECT 87.821 4.841 87.895 5.075 ;
      RECT 87.445 4.092 87.615 4.33 ;
      RECT 87.445 4.092 87.701 4.244 ;
      RECT 87.445 4.092 87.705 4.154 ;
      RECT 87.495 3.865 87.715 4.133 ;
      RECT 87.49 3.882 87.72 4.106 ;
      RECT 87.455 4.04 87.72 4.106 ;
      RECT 87.475 3.89 87.615 4.33 ;
      RECT 87.465 3.972 87.725 4.089 ;
      RECT 87.46 4.02 87.725 4.089 ;
      RECT 87.465 3.93 87.72 4.106 ;
      RECT 87.49 3.867 87.715 4.133 ;
      RECT 87.055 3.842 87.225 4.04 ;
      RECT 87.055 3.842 87.27 4.015 ;
      RECT 87.125 3.785 87.295 3.973 ;
      RECT 87.1 3.8 87.295 3.973 ;
      RECT 86.715 3.846 86.745 4.04 ;
      RECT 86.71 3.818 86.715 4.04 ;
      RECT 86.68 3.792 86.71 4.042 ;
      RECT 86.655 3.75 86.68 4.045 ;
      RECT 86.645 3.722 86.655 4.047 ;
      RECT 86.61 3.702 86.645 4.049 ;
      RECT 86.545 3.687 86.61 4.055 ;
      RECT 86.495 3.685 86.545 4.061 ;
      RECT 86.472 3.687 86.495 4.066 ;
      RECT 86.386 3.698 86.472 4.072 ;
      RECT 86.3 3.716 86.386 4.082 ;
      RECT 86.285 3.727 86.3 4.088 ;
      RECT 86.215 3.75 86.285 4.094 ;
      RECT 86.16 3.782 86.215 4.102 ;
      RECT 86.12 3.805 86.16 4.108 ;
      RECT 86.106 3.818 86.12 4.111 ;
      RECT 86.02 3.84 86.106 4.117 ;
      RECT 86.005 3.865 86.02 4.123 ;
      RECT 85.965 3.88 86.005 4.127 ;
      RECT 85.915 3.895 85.965 4.132 ;
      RECT 85.89 3.902 85.915 4.136 ;
      RECT 85.83 3.897 85.89 4.14 ;
      RECT 85.815 3.888 85.83 4.144 ;
      RECT 85.745 3.878 85.815 4.14 ;
      RECT 85.72 3.87 85.74 4.13 ;
      RECT 85.661 3.87 85.72 4.108 ;
      RECT 85.575 3.87 85.661 4.065 ;
      RECT 85.74 3.87 85.745 4.135 ;
      RECT 86.435 3.101 86.605 3.435 ;
      RECT 86.405 3.101 86.605 3.43 ;
      RECT 86.345 3.068 86.405 3.418 ;
      RECT 86.345 3.124 86.615 3.413 ;
      RECT 86.32 3.124 86.615 3.407 ;
      RECT 86.315 3.065 86.345 3.404 ;
      RECT 86.3 3.071 86.435 3.402 ;
      RECT 86.295 3.079 86.52 3.39 ;
      RECT 86.295 3.131 86.63 3.343 ;
      RECT 86.28 3.087 86.52 3.338 ;
      RECT 86.28 3.157 86.64 3.279 ;
      RECT 86.25 3.107 86.605 3.24 ;
      RECT 86.25 3.197 86.65 3.236 ;
      RECT 86.3 3.076 86.52 3.402 ;
      RECT 85.64 3.406 85.695 3.67 ;
      RECT 85.64 3.406 85.76 3.669 ;
      RECT 85.64 3.406 85.785 3.668 ;
      RECT 85.64 3.406 85.85 3.667 ;
      RECT 85.785 3.372 85.865 3.666 ;
      RECT 85.6 3.416 86.01 3.665 ;
      RECT 85.64 3.413 86.01 3.665 ;
      RECT 85.6 3.421 86.015 3.658 ;
      RECT 85.585 3.423 86.015 3.657 ;
      RECT 85.585 3.43 86.02 3.653 ;
      RECT 85.565 3.429 86.015 3.649 ;
      RECT 85.565 3.437 86.025 3.648 ;
      RECT 85.56 3.434 86.02 3.644 ;
      RECT 85.56 3.447 86.035 3.643 ;
      RECT 85.545 3.437 86.025 3.642 ;
      RECT 85.51 3.45 86.035 3.635 ;
      RECT 85.695 3.405 86.005 3.665 ;
      RECT 85.695 3.39 85.955 3.665 ;
      RECT 85.76 3.377 85.89 3.665 ;
      RECT 85.305 4.466 85.32 4.859 ;
      RECT 85.27 4.471 85.32 4.858 ;
      RECT 85.305 4.47 85.365 4.857 ;
      RECT 85.25 4.481 85.365 4.856 ;
      RECT 85.265 4.477 85.365 4.856 ;
      RECT 85.23 4.487 85.44 4.853 ;
      RECT 85.23 4.506 85.485 4.851 ;
      RECT 85.23 4.513 85.49 4.848 ;
      RECT 85.215 4.49 85.44 4.845 ;
      RECT 85.195 4.495 85.44 4.838 ;
      RECT 85.19 4.499 85.44 4.834 ;
      RECT 85.19 4.516 85.5 4.833 ;
      RECT 85.17 4.51 85.485 4.829 ;
      RECT 85.17 4.519 85.505 4.823 ;
      RECT 85.165 4.525 85.505 4.595 ;
      RECT 85.23 4.485 85.365 4.853 ;
      RECT 85.105 3.848 85.305 4.16 ;
      RECT 85.18 3.826 85.305 4.16 ;
      RECT 85.12 3.845 85.31 4.145 ;
      RECT 85.09 3.856 85.31 4.143 ;
      RECT 85.105 3.851 85.315 4.109 ;
      RECT 85.09 3.955 85.32 4.076 ;
      RECT 85.12 3.827 85.305 4.16 ;
      RECT 85.18 3.805 85.28 4.16 ;
      RECT 85.205 3.802 85.28 4.16 ;
      RECT 85.205 3.797 85.225 4.16 ;
      RECT 84.61 3.865 84.785 4.04 ;
      RECT 84.605 3.865 84.785 4.038 ;
      RECT 84.58 3.865 84.785 4.033 ;
      RECT 84.525 3.845 84.695 4.023 ;
      RECT 84.525 3.852 84.76 4.023 ;
      RECT 84.61 4.532 84.625 4.715 ;
      RECT 84.6 4.51 84.61 4.715 ;
      RECT 84.585 4.49 84.6 4.715 ;
      RECT 84.575 4.465 84.585 4.715 ;
      RECT 84.545 4.43 84.575 4.715 ;
      RECT 84.51 4.37 84.545 4.715 ;
      RECT 84.505 4.332 84.51 4.715 ;
      RECT 84.455 4.283 84.505 4.715 ;
      RECT 84.445 4.233 84.455 4.703 ;
      RECT 84.43 4.212 84.445 4.663 ;
      RECT 84.41 4.18 84.43 4.613 ;
      RECT 84.385 4.136 84.41 4.553 ;
      RECT 84.38 4.108 84.385 4.508 ;
      RECT 84.375 4.099 84.38 4.494 ;
      RECT 84.37 4.092 84.375 4.481 ;
      RECT 84.365 4.087 84.37 4.47 ;
      RECT 84.36 4.072 84.365 4.46 ;
      RECT 84.355 4.05 84.36 4.447 ;
      RECT 84.345 4.01 84.355 4.422 ;
      RECT 84.32 3.94 84.345 4.378 ;
      RECT 84.315 3.88 84.32 4.343 ;
      RECT 84.3 3.86 84.315 4.31 ;
      RECT 84.295 3.86 84.3 4.285 ;
      RECT 84.265 3.86 84.295 4.24 ;
      RECT 84.22 3.86 84.265 4.18 ;
      RECT 84.145 3.86 84.22 4.128 ;
      RECT 84.14 3.86 84.145 4.093 ;
      RECT 84.135 3.86 84.14 4.083 ;
      RECT 84.13 3.86 84.135 4.063 ;
      RECT 84.395 3.08 84.565 3.55 ;
      RECT 84.34 3.073 84.535 3.534 ;
      RECT 84.34 3.087 84.57 3.533 ;
      RECT 84.325 3.088 84.57 3.514 ;
      RECT 84.32 3.106 84.57 3.5 ;
      RECT 84.325 3.089 84.575 3.498 ;
      RECT 84.31 3.12 84.575 3.483 ;
      RECT 84.325 3.095 84.58 3.468 ;
      RECT 84.305 3.135 84.58 3.465 ;
      RECT 84.32 3.107 84.585 3.45 ;
      RECT 84.32 3.119 84.59 3.43 ;
      RECT 84.305 3.135 84.595 3.413 ;
      RECT 84.305 3.145 84.6 3.268 ;
      RECT 84.3 3.145 84.6 3.225 ;
      RECT 84.3 3.16 84.605 3.203 ;
      RECT 84.395 3.07 84.535 3.55 ;
      RECT 84.395 3.068 84.505 3.55 ;
      RECT 84.481 3.065 84.505 3.55 ;
      RECT 84.14 4.732 84.145 4.778 ;
      RECT 84.13 4.58 84.14 4.802 ;
      RECT 84.125 4.425 84.13 4.827 ;
      RECT 84.11 4.387 84.125 4.838 ;
      RECT 84.105 4.37 84.11 4.845 ;
      RECT 84.095 4.358 84.105 4.852 ;
      RECT 84.09 4.349 84.095 4.854 ;
      RECT 84.085 4.347 84.09 4.858 ;
      RECT 84.04 4.338 84.085 4.873 ;
      RECT 84.035 4.33 84.04 4.887 ;
      RECT 84.03 4.327 84.035 4.891 ;
      RECT 84.015 4.322 84.03 4.899 ;
      RECT 83.96 4.312 84.015 4.91 ;
      RECT 83.925 4.3 83.96 4.911 ;
      RECT 83.916 4.295 83.925 4.905 ;
      RECT 83.83 4.295 83.916 4.895 ;
      RECT 83.8 4.295 83.83 4.873 ;
      RECT 83.79 4.295 83.795 4.853 ;
      RECT 83.785 4.295 83.79 4.815 ;
      RECT 83.78 4.295 83.785 4.773 ;
      RECT 83.775 4.295 83.78 4.733 ;
      RECT 83.77 4.295 83.775 4.663 ;
      RECT 83.76 4.295 83.77 4.585 ;
      RECT 83.755 4.295 83.76 4.485 ;
      RECT 83.795 4.295 83.8 4.855 ;
      RECT 83.29 4.377 83.38 4.855 ;
      RECT 83.275 4.38 83.395 4.853 ;
      RECT 83.29 4.379 83.395 4.853 ;
      RECT 83.255 4.386 83.42 4.843 ;
      RECT 83.275 4.38 83.42 4.843 ;
      RECT 83.24 4.392 83.42 4.831 ;
      RECT 83.275 4.383 83.47 4.824 ;
      RECT 83.226 4.4 83.47 4.822 ;
      RECT 83.255 4.39 83.48 4.81 ;
      RECT 83.226 4.411 83.51 4.801 ;
      RECT 83.14 4.435 83.51 4.795 ;
      RECT 83.14 4.448 83.55 4.778 ;
      RECT 83.135 4.47 83.55 4.771 ;
      RECT 83.105 4.485 83.55 4.761 ;
      RECT 83.1 4.496 83.55 4.751 ;
      RECT 83.07 4.509 83.55 4.742 ;
      RECT 83.055 4.527 83.55 4.731 ;
      RECT 83.03 4.54 83.55 4.721 ;
      RECT 83.29 4.376 83.3 4.855 ;
      RECT 83.336 3.8 83.375 4.045 ;
      RECT 83.25 3.8 83.385 4.043 ;
      RECT 83.135 3.825 83.385 4.04 ;
      RECT 83.135 3.825 83.39 4.038 ;
      RECT 83.135 3.825 83.405 4.033 ;
      RECT 83.241 3.8 83.42 4.013 ;
      RECT 83.155 3.808 83.42 4.013 ;
      RECT 82.825 3.16 82.995 3.595 ;
      RECT 82.815 3.194 82.995 3.578 ;
      RECT 82.895 3.13 83.065 3.565 ;
      RECT 82.8 3.205 83.065 3.543 ;
      RECT 82.895 3.14 83.07 3.533 ;
      RECT 82.825 3.192 83.1 3.518 ;
      RECT 82.785 3.218 83.1 3.503 ;
      RECT 82.785 3.26 83.11 3.483 ;
      RECT 82.78 3.285 83.115 3.465 ;
      RECT 82.78 3.295 83.12 3.45 ;
      RECT 82.775 3.232 83.1 3.448 ;
      RECT 82.775 3.305 83.125 3.433 ;
      RECT 82.77 3.242 83.1 3.43 ;
      RECT 82.765 3.326 83.13 3.413 ;
      RECT 82.765 3.358 83.135 3.393 ;
      RECT 82.76 3.272 83.11 3.385 ;
      RECT 82.765 3.257 83.1 3.413 ;
      RECT 82.78 3.227 83.1 3.465 ;
      RECT 82.625 3.814 82.85 4.07 ;
      RECT 82.625 3.847 82.87 4.06 ;
      RECT 82.59 3.847 82.87 4.058 ;
      RECT 82.59 3.86 82.875 4.048 ;
      RECT 82.59 3.88 82.885 4.04 ;
      RECT 82.59 3.977 82.89 4.033 ;
      RECT 82.57 3.725 82.7 4.023 ;
      RECT 82.525 3.88 82.885 3.965 ;
      RECT 82.515 3.725 82.7 3.91 ;
      RECT 82.515 3.757 82.786 3.91 ;
      RECT 82.48 4.287 82.5 4.465 ;
      RECT 82.445 4.24 82.48 4.465 ;
      RECT 82.43 4.18 82.445 4.465 ;
      RECT 82.405 4.127 82.43 4.465 ;
      RECT 82.39 4.08 82.405 4.465 ;
      RECT 82.37 4.057 82.39 4.465 ;
      RECT 82.345 4.022 82.37 4.465 ;
      RECT 82.335 3.868 82.345 4.465 ;
      RECT 82.305 3.863 82.335 4.456 ;
      RECT 82.3 3.86 82.305 4.446 ;
      RECT 82.285 3.86 82.3 4.42 ;
      RECT 82.28 3.86 82.285 4.383 ;
      RECT 82.255 3.86 82.28 4.335 ;
      RECT 82.235 3.86 82.255 4.26 ;
      RECT 82.225 3.86 82.235 4.22 ;
      RECT 82.22 3.86 82.225 4.195 ;
      RECT 82.215 3.86 82.22 4.178 ;
      RECT 82.21 3.86 82.215 4.16 ;
      RECT 82.205 3.861 82.21 4.15 ;
      RECT 82.195 3.863 82.205 4.118 ;
      RECT 82.185 3.865 82.195 4.085 ;
      RECT 82.175 3.868 82.185 4.058 ;
      RECT 82.5 4.295 82.725 4.465 ;
      RECT 81.83 3.107 82 3.56 ;
      RECT 81.83 3.107 82.09 3.526 ;
      RECT 81.83 3.107 82.12 3.51 ;
      RECT 81.83 3.107 82.15 3.483 ;
      RECT 82.086 3.085 82.165 3.465 ;
      RECT 81.865 3.092 82.17 3.45 ;
      RECT 81.865 3.1 82.18 3.413 ;
      RECT 81.825 3.127 82.18 3.385 ;
      RECT 81.81 3.14 82.18 3.35 ;
      RECT 81.83 3.115 82.2 3.34 ;
      RECT 81.805 3.18 82.2 3.31 ;
      RECT 81.805 3.21 82.205 3.293 ;
      RECT 81.8 3.24 82.205 3.28 ;
      RECT 81.865 3.089 82.165 3.465 ;
      RECT 82 3.086 82.086 3.544 ;
      RECT 81.951 3.087 82.165 3.465 ;
      RECT 82.095 4.747 82.14 4.94 ;
      RECT 82.085 4.717 82.095 4.94 ;
      RECT 82.08 4.702 82.085 4.94 ;
      RECT 82.04 4.612 82.08 4.94 ;
      RECT 82.035 4.525 82.04 4.94 ;
      RECT 82.025 4.495 82.035 4.94 ;
      RECT 82.02 4.455 82.025 4.94 ;
      RECT 82.01 4.417 82.02 4.94 ;
      RECT 82.005 4.382 82.01 4.94 ;
      RECT 81.985 4.335 82.005 4.94 ;
      RECT 81.97 4.26 81.985 4.94 ;
      RECT 81.965 4.215 81.97 4.935 ;
      RECT 81.96 4.195 81.965 4.908 ;
      RECT 81.955 4.175 81.96 4.893 ;
      RECT 81.95 4.15 81.955 4.873 ;
      RECT 81.945 4.128 81.95 4.858 ;
      RECT 81.94 4.106 81.945 4.84 ;
      RECT 81.935 4.085 81.94 4.83 ;
      RECT 81.925 4.057 81.935 4.8 ;
      RECT 81.915 4.02 81.925 4.768 ;
      RECT 81.905 3.98 81.915 4.735 ;
      RECT 81.895 3.958 81.905 4.705 ;
      RECT 81.865 3.91 81.895 4.637 ;
      RECT 81.85 3.87 81.865 4.564 ;
      RECT 81.84 3.87 81.85 4.53 ;
      RECT 81.835 3.87 81.84 4.505 ;
      RECT 81.83 3.87 81.835 4.49 ;
      RECT 81.825 3.87 81.83 4.468 ;
      RECT 81.82 3.87 81.825 4.455 ;
      RECT 81.805 3.87 81.82 4.42 ;
      RECT 81.785 3.87 81.805 4.36 ;
      RECT 81.775 3.87 81.785 4.31 ;
      RECT 81.755 3.87 81.775 4.258 ;
      RECT 81.735 3.87 81.755 4.215 ;
      RECT 81.725 3.87 81.735 4.203 ;
      RECT 81.695 3.87 81.725 4.19 ;
      RECT 81.665 3.891 81.695 4.17 ;
      RECT 81.655 3.919 81.665 4.15 ;
      RECT 81.64 3.936 81.655 4.118 ;
      RECT 81.635 3.95 81.64 4.085 ;
      RECT 81.63 3.958 81.635 4.058 ;
      RECT 81.625 3.966 81.63 4.02 ;
      RECT 81.63 4.49 81.635 4.825 ;
      RECT 81.595 4.477 81.63 4.824 ;
      RECT 81.525 4.417 81.595 4.823 ;
      RECT 81.445 4.36 81.525 4.822 ;
      RECT 81.31 4.32 81.445 4.821 ;
      RECT 81.31 4.507 81.645 4.81 ;
      RECT 81.27 4.507 81.645 4.8 ;
      RECT 81.27 4.525 81.65 4.795 ;
      RECT 81.27 4.615 81.655 4.785 ;
      RECT 81.265 4.31 81.43 4.765 ;
      RECT 81.26 4.31 81.43 4.508 ;
      RECT 81.26 4.467 81.625 4.508 ;
      RECT 81.26 4.455 81.62 4.508 ;
      RECT 80.395 7.3 80.565 8.77 ;
      RECT 80.395 7.3 80.57 8.56 ;
      RECT 80.025 9.25 80.495 9.42 ;
      RECT 80.025 8.23 80.195 9.42 ;
      RECT 80.02 3.04 80.19 4.23 ;
      RECT 80.02 3.04 80.49 3.21 ;
      RECT 79.4 3.895 79.575 5.155 ;
      RECT 79.4 3.685 79.57 5.155 ;
      RECT 79.4 7.305 79.57 8.775 ;
      RECT 79.4 7.305 79.575 8.565 ;
      RECT 79.03 3.035 79.2 4.225 ;
      RECT 79.03 3.035 79.5 3.205 ;
      RECT 79.03 9.255 79.5 9.425 ;
      RECT 79.03 8.235 79.2 9.425 ;
      RECT 78.04 4.015 78.215 5.155 ;
      RECT 78.04 1.865 78.21 5.155 ;
      RECT 78.04 1.865 78.215 2.415 ;
      RECT 78.04 10.045 78.215 10.595 ;
      RECT 78.04 7.305 78.21 10.595 ;
      RECT 78.04 7.305 78.215 8.445 ;
      RECT 77.61 3.895 77.785 5.155 ;
      RECT 77.61 2.945 77.78 5.155 ;
      RECT 77.61 7.305 77.78 9.515 ;
      RECT 77.61 7.305 77.785 8.565 ;
      RECT 77.18 3.925 77.35 5.155 ;
      RECT 77.24 2.145 77.41 4.095 ;
      RECT 77.18 1.865 77.35 2.315 ;
      RECT 77.18 10.145 77.35 10.595 ;
      RECT 77.24 8.365 77.41 10.315 ;
      RECT 77.18 7.305 77.35 8.535 ;
      RECT 76.655 3.895 76.83 5.155 ;
      RECT 76.655 1.865 76.825 5.155 ;
      RECT 76.655 3.365 77.065 3.695 ;
      RECT 76.655 2.525 77.065 2.855 ;
      RECT 76.655 1.865 76.83 2.355 ;
      RECT 76.655 10.105 76.83 10.595 ;
      RECT 76.655 7.305 76.825 10.595 ;
      RECT 76.655 9.605 77.065 9.935 ;
      RECT 76.655 8.765 77.065 9.095 ;
      RECT 76.655 7.305 76.83 8.565 ;
      RECT 73.995 3.27 74.725 3.51 ;
      RECT 74.537 3.065 74.725 3.51 ;
      RECT 74.365 3.077 74.74 3.504 ;
      RECT 74.28 3.092 74.76 3.489 ;
      RECT 74.28 3.107 74.765 3.479 ;
      RECT 74.235 3.127 74.78 3.471 ;
      RECT 74.212 3.162 74.795 3.425 ;
      RECT 74.126 3.185 74.8 3.385 ;
      RECT 74.126 3.203 74.81 3.355 ;
      RECT 73.995 3.272 74.815 3.318 ;
      RECT 74.04 3.215 74.81 3.355 ;
      RECT 74.126 3.167 74.795 3.425 ;
      RECT 74.212 3.136 74.78 3.471 ;
      RECT 74.235 3.117 74.765 3.479 ;
      RECT 74.28 3.09 74.74 3.504 ;
      RECT 74.365 3.072 74.725 3.51 ;
      RECT 74.451 3.066 74.725 3.51 ;
      RECT 74.537 3.061 74.67 3.51 ;
      RECT 74.623 3.056 74.67 3.51 ;
      RECT 74.185 4.67 74.19 4.683 ;
      RECT 74.18 4.565 74.185 4.688 ;
      RECT 74.155 4.425 74.18 4.703 ;
      RECT 74.12 4.376 74.155 4.735 ;
      RECT 74.115 4.344 74.12 4.755 ;
      RECT 74.11 4.335 74.115 4.755 ;
      RECT 74.03 4.3 74.11 4.755 ;
      RECT 73.967 4.27 74.03 4.755 ;
      RECT 73.881 4.258 73.967 4.755 ;
      RECT 73.795 4.244 73.881 4.755 ;
      RECT 73.715 4.231 73.795 4.741 ;
      RECT 73.68 4.223 73.715 4.721 ;
      RECT 73.67 4.22 73.68 4.712 ;
      RECT 73.64 4.215 73.67 4.699 ;
      RECT 73.59 4.19 73.64 4.675 ;
      RECT 73.576 4.164 73.59 4.657 ;
      RECT 73.49 4.124 73.576 4.633 ;
      RECT 73.445 4.072 73.49 4.602 ;
      RECT 73.435 4.047 73.445 4.589 ;
      RECT 73.43 3.828 73.435 3.85 ;
      RECT 73.425 4.03 73.435 4.585 ;
      RECT 73.425 3.826 73.43 3.94 ;
      RECT 73.415 3.822 73.425 4.581 ;
      RECT 73.371 3.82 73.415 4.569 ;
      RECT 73.285 3.82 73.371 4.54 ;
      RECT 73.255 3.82 73.285 4.513 ;
      RECT 73.24 3.82 73.255 4.501 ;
      RECT 73.2 3.832 73.24 4.486 ;
      RECT 73.18 3.851 73.2 4.465 ;
      RECT 73.17 3.861 73.18 4.449 ;
      RECT 73.16 3.867 73.17 4.438 ;
      RECT 73.14 3.877 73.16 4.421 ;
      RECT 73.135 3.886 73.14 4.408 ;
      RECT 73.13 3.89 73.135 4.358 ;
      RECT 73.12 3.896 73.13 4.275 ;
      RECT 73.115 3.9 73.12 4.189 ;
      RECT 73.11 3.92 73.115 4.126 ;
      RECT 73.105 3.943 73.11 4.073 ;
      RECT 73.1 3.961 73.105 4.018 ;
      RECT 73.71 3.78 73.88 4.04 ;
      RECT 73.88 3.745 73.925 4.026 ;
      RECT 73.841 3.747 73.93 4.009 ;
      RECT 73.73 3.764 74.016 3.98 ;
      RECT 73.73 3.779 74.02 3.952 ;
      RECT 73.73 3.76 73.93 4.009 ;
      RECT 73.755 3.748 73.88 4.04 ;
      RECT 73.841 3.746 73.925 4.026 ;
      RECT 73.26 10.045 73.435 10.595 ;
      RECT 73.26 7.305 73.43 10.595 ;
      RECT 73.26 7.305 73.435 8.445 ;
      RECT 72.895 3.135 73.065 3.625 ;
      RECT 72.895 3.135 73.1 3.605 ;
      RECT 73.03 3.055 73.14 3.565 ;
      RECT 73.011 3.059 73.16 3.535 ;
      RECT 72.925 3.067 73.18 3.518 ;
      RECT 72.925 3.073 73.185 3.508 ;
      RECT 72.925 3.082 73.205 3.496 ;
      RECT 72.9 3.107 73.235 3.474 ;
      RECT 72.9 3.127 73.24 3.454 ;
      RECT 72.895 3.14 73.25 3.434 ;
      RECT 72.895 3.207 73.255 3.415 ;
      RECT 72.895 3.34 73.26 3.402 ;
      RECT 72.89 3.145 73.25 3.235 ;
      RECT 72.9 3.102 73.205 3.496 ;
      RECT 73.011 3.057 73.14 3.565 ;
      RECT 72.885 4.81 73.185 5.065 ;
      RECT 72.97 4.776 73.185 5.065 ;
      RECT 72.97 4.779 73.19 4.925 ;
      RECT 72.905 4.8 73.19 4.925 ;
      RECT 72.94 4.79 73.185 5.065 ;
      RECT 72.935 4.795 73.19 4.925 ;
      RECT 72.97 4.774 73.171 5.065 ;
      RECT 73.056 4.765 73.171 5.065 ;
      RECT 73.056 4.759 73.085 5.065 ;
      RECT 72.83 7.305 73 9.515 ;
      RECT 72.83 7.305 73.005 8.565 ;
      RECT 72.545 4.4 72.555 4.89 ;
      RECT 72.205 4.335 72.215 4.635 ;
      RECT 72.72 4.507 72.725 4.726 ;
      RECT 72.71 4.487 72.72 4.743 ;
      RECT 72.7 4.467 72.71 4.773 ;
      RECT 72.695 4.457 72.7 4.788 ;
      RECT 72.69 4.453 72.695 4.793 ;
      RECT 72.675 4.445 72.69 4.8 ;
      RECT 72.635 4.425 72.675 4.825 ;
      RECT 72.61 4.407 72.635 4.858 ;
      RECT 72.605 4.405 72.61 4.871 ;
      RECT 72.585 4.402 72.605 4.875 ;
      RECT 72.555 4.4 72.585 4.885 ;
      RECT 72.485 4.402 72.545 4.886 ;
      RECT 72.465 4.402 72.485 4.88 ;
      RECT 72.44 4.4 72.465 4.877 ;
      RECT 72.405 4.395 72.44 4.873 ;
      RECT 72.385 4.389 72.405 4.86 ;
      RECT 72.375 4.386 72.385 4.848 ;
      RECT 72.355 4.383 72.375 4.833 ;
      RECT 72.335 4.379 72.355 4.815 ;
      RECT 72.33 4.376 72.335 4.805 ;
      RECT 72.325 4.375 72.33 4.803 ;
      RECT 72.315 4.372 72.325 4.795 ;
      RECT 72.305 4.366 72.315 4.778 ;
      RECT 72.295 4.36 72.305 4.76 ;
      RECT 72.285 4.354 72.295 4.748 ;
      RECT 72.275 4.348 72.285 4.728 ;
      RECT 72.27 4.344 72.275 4.713 ;
      RECT 72.265 4.342 72.27 4.705 ;
      RECT 72.26 4.34 72.265 4.698 ;
      RECT 72.255 4.338 72.26 4.688 ;
      RECT 72.25 4.336 72.255 4.682 ;
      RECT 72.24 4.335 72.25 4.672 ;
      RECT 72.23 4.335 72.24 4.663 ;
      RECT 72.215 4.335 72.23 4.648 ;
      RECT 72.175 4.335 72.205 4.632 ;
      RECT 72.155 4.337 72.175 4.627 ;
      RECT 72.15 4.342 72.155 4.625 ;
      RECT 72.12 4.35 72.15 4.623 ;
      RECT 72.09 4.365 72.12 4.622 ;
      RECT 72.045 4.387 72.09 4.627 ;
      RECT 72.04 4.402 72.045 4.631 ;
      RECT 72.025 4.407 72.04 4.633 ;
      RECT 72.02 4.411 72.025 4.635 ;
      RECT 71.96 4.434 72.02 4.644 ;
      RECT 71.94 4.46 71.96 4.657 ;
      RECT 71.93 4.467 71.94 4.661 ;
      RECT 71.915 4.474 71.93 4.664 ;
      RECT 71.895 4.484 71.915 4.667 ;
      RECT 71.89 4.492 71.895 4.67 ;
      RECT 71.845 4.497 71.89 4.677 ;
      RECT 71.835 4.5 71.845 4.684 ;
      RECT 71.825 4.5 71.835 4.688 ;
      RECT 71.79 4.502 71.825 4.7 ;
      RECT 71.77 4.505 71.79 4.713 ;
      RECT 71.73 4.508 71.77 4.724 ;
      RECT 71.715 4.51 71.73 4.737 ;
      RECT 71.705 4.51 71.715 4.742 ;
      RECT 71.68 4.511 71.705 4.75 ;
      RECT 71.67 4.513 71.68 4.755 ;
      RECT 71.665 4.514 71.67 4.758 ;
      RECT 71.64 4.512 71.665 4.761 ;
      RECT 71.625 4.51 71.64 4.762 ;
      RECT 71.605 4.507 71.625 4.764 ;
      RECT 71.585 4.502 71.605 4.764 ;
      RECT 71.525 4.497 71.585 4.761 ;
      RECT 71.49 4.472 71.525 4.757 ;
      RECT 71.48 4.449 71.49 4.755 ;
      RECT 71.45 4.426 71.48 4.755 ;
      RECT 71.44 4.405 71.45 4.755 ;
      RECT 71.415 4.387 71.44 4.753 ;
      RECT 71.4 4.365 71.415 4.75 ;
      RECT 71.385 4.347 71.4 4.748 ;
      RECT 71.365 4.337 71.385 4.746 ;
      RECT 71.35 4.332 71.365 4.745 ;
      RECT 71.335 4.33 71.35 4.744 ;
      RECT 71.305 4.331 71.335 4.742 ;
      RECT 71.285 4.334 71.305 4.74 ;
      RECT 71.228 4.338 71.285 4.74 ;
      RECT 71.142 4.347 71.228 4.74 ;
      RECT 71.056 4.358 71.142 4.74 ;
      RECT 70.97 4.369 71.056 4.74 ;
      RECT 70.95 4.376 70.97 4.748 ;
      RECT 70.94 4.379 70.95 4.755 ;
      RECT 70.875 4.384 70.94 4.773 ;
      RECT 70.845 4.391 70.875 4.798 ;
      RECT 70.835 4.394 70.845 4.805 ;
      RECT 70.79 4.398 70.835 4.81 ;
      RECT 70.76 4.403 70.79 4.815 ;
      RECT 70.759 4.405 70.76 4.815 ;
      RECT 70.673 4.411 70.759 4.815 ;
      RECT 70.587 4.422 70.673 4.815 ;
      RECT 70.501 4.434 70.587 4.815 ;
      RECT 70.415 4.445 70.501 4.815 ;
      RECT 70.4 4.452 70.415 4.81 ;
      RECT 70.395 4.454 70.4 4.804 ;
      RECT 70.375 4.465 70.395 4.799 ;
      RECT 70.365 4.483 70.375 4.793 ;
      RECT 70.36 4.495 70.365 4.593 ;
      RECT 72.655 3.248 72.675 3.335 ;
      RECT 72.65 3.183 72.655 3.367 ;
      RECT 72.64 3.15 72.65 3.372 ;
      RECT 72.635 3.13 72.64 3.378 ;
      RECT 72.605 3.13 72.635 3.395 ;
      RECT 72.556 3.13 72.605 3.431 ;
      RECT 72.47 3.13 72.556 3.489 ;
      RECT 72.441 3.14 72.47 3.538 ;
      RECT 72.355 3.182 72.441 3.591 ;
      RECT 72.335 3.22 72.355 3.638 ;
      RECT 72.31 3.237 72.335 3.658 ;
      RECT 72.3 3.251 72.31 3.678 ;
      RECT 72.295 3.257 72.3 3.688 ;
      RECT 72.29 3.261 72.295 3.695 ;
      RECT 72.24 3.281 72.29 3.7 ;
      RECT 72.175 3.325 72.24 3.7 ;
      RECT 72.15 3.375 72.175 3.7 ;
      RECT 72.14 3.405 72.15 3.7 ;
      RECT 72.135 3.432 72.14 3.7 ;
      RECT 72.13 3.45 72.135 3.7 ;
      RECT 72.12 3.492 72.13 3.7 ;
      RECT 71.875 10.105 72.05 10.595 ;
      RECT 71.875 7.305 72.045 10.595 ;
      RECT 71.875 9.605 72.285 9.935 ;
      RECT 71.875 8.765 72.285 9.095 ;
      RECT 71.875 7.305 72.05 8.565 ;
      RECT 71.95 4.85 72.14 5.075 ;
      RECT 71.94 4.851 72.145 5.07 ;
      RECT 71.94 4.853 72.155 5.05 ;
      RECT 71.94 4.857 72.16 5.035 ;
      RECT 71.94 4.844 72.11 5.07 ;
      RECT 71.94 4.847 72.135 5.07 ;
      RECT 71.95 4.843 72.11 5.075 ;
      RECT 72.036 4.841 72.11 5.075 ;
      RECT 71.66 4.092 71.83 4.33 ;
      RECT 71.66 4.092 71.916 4.244 ;
      RECT 71.66 4.092 71.92 4.154 ;
      RECT 71.71 3.865 71.93 4.133 ;
      RECT 71.705 3.882 71.935 4.106 ;
      RECT 71.67 4.04 71.935 4.106 ;
      RECT 71.69 3.89 71.83 4.33 ;
      RECT 71.68 3.972 71.94 4.089 ;
      RECT 71.675 4.02 71.94 4.089 ;
      RECT 71.68 3.93 71.935 4.106 ;
      RECT 71.705 3.867 71.93 4.133 ;
      RECT 71.27 3.842 71.44 4.04 ;
      RECT 71.27 3.842 71.485 4.015 ;
      RECT 71.34 3.785 71.51 3.973 ;
      RECT 71.315 3.8 71.51 3.973 ;
      RECT 70.93 3.846 70.96 4.04 ;
      RECT 70.925 3.818 70.93 4.04 ;
      RECT 70.895 3.792 70.925 4.042 ;
      RECT 70.87 3.75 70.895 4.045 ;
      RECT 70.86 3.722 70.87 4.047 ;
      RECT 70.825 3.702 70.86 4.049 ;
      RECT 70.76 3.687 70.825 4.055 ;
      RECT 70.71 3.685 70.76 4.061 ;
      RECT 70.687 3.687 70.71 4.066 ;
      RECT 70.601 3.698 70.687 4.072 ;
      RECT 70.515 3.716 70.601 4.082 ;
      RECT 70.5 3.727 70.515 4.088 ;
      RECT 70.43 3.75 70.5 4.094 ;
      RECT 70.375 3.782 70.43 4.102 ;
      RECT 70.335 3.805 70.375 4.108 ;
      RECT 70.321 3.818 70.335 4.111 ;
      RECT 70.235 3.84 70.321 4.117 ;
      RECT 70.22 3.865 70.235 4.123 ;
      RECT 70.18 3.88 70.22 4.127 ;
      RECT 70.13 3.895 70.18 4.132 ;
      RECT 70.105 3.902 70.13 4.136 ;
      RECT 70.045 3.897 70.105 4.14 ;
      RECT 70.03 3.888 70.045 4.144 ;
      RECT 69.96 3.878 70.03 4.14 ;
      RECT 69.935 3.87 69.955 4.13 ;
      RECT 69.876 3.87 69.935 4.108 ;
      RECT 69.79 3.87 69.876 4.065 ;
      RECT 69.955 3.87 69.96 4.135 ;
      RECT 70.65 3.101 70.82 3.435 ;
      RECT 70.62 3.101 70.82 3.43 ;
      RECT 70.56 3.068 70.62 3.418 ;
      RECT 70.56 3.124 70.83 3.413 ;
      RECT 70.535 3.124 70.83 3.407 ;
      RECT 70.53 3.065 70.56 3.404 ;
      RECT 70.515 3.071 70.65 3.402 ;
      RECT 70.51 3.079 70.735 3.39 ;
      RECT 70.51 3.131 70.845 3.343 ;
      RECT 70.495 3.087 70.735 3.338 ;
      RECT 70.495 3.157 70.855 3.279 ;
      RECT 70.465 3.107 70.82 3.24 ;
      RECT 70.465 3.197 70.865 3.236 ;
      RECT 70.515 3.076 70.735 3.402 ;
      RECT 69.855 3.406 69.91 3.67 ;
      RECT 69.855 3.406 69.975 3.669 ;
      RECT 69.855 3.406 70 3.668 ;
      RECT 69.855 3.406 70.065 3.667 ;
      RECT 70 3.372 70.08 3.666 ;
      RECT 69.815 3.416 70.225 3.665 ;
      RECT 69.855 3.413 70.225 3.665 ;
      RECT 69.815 3.421 70.23 3.658 ;
      RECT 69.8 3.423 70.23 3.657 ;
      RECT 69.8 3.43 70.235 3.653 ;
      RECT 69.78 3.429 70.23 3.649 ;
      RECT 69.78 3.437 70.24 3.648 ;
      RECT 69.775 3.434 70.235 3.644 ;
      RECT 69.775 3.447 70.25 3.643 ;
      RECT 69.76 3.437 70.24 3.642 ;
      RECT 69.725 3.45 70.25 3.635 ;
      RECT 69.91 3.405 70.22 3.665 ;
      RECT 69.91 3.39 70.17 3.665 ;
      RECT 69.975 3.377 70.105 3.665 ;
      RECT 69.52 4.466 69.535 4.859 ;
      RECT 69.485 4.471 69.535 4.858 ;
      RECT 69.52 4.47 69.58 4.857 ;
      RECT 69.465 4.481 69.58 4.856 ;
      RECT 69.48 4.477 69.58 4.856 ;
      RECT 69.445 4.487 69.655 4.853 ;
      RECT 69.445 4.506 69.7 4.851 ;
      RECT 69.445 4.513 69.705 4.848 ;
      RECT 69.43 4.49 69.655 4.845 ;
      RECT 69.41 4.495 69.655 4.838 ;
      RECT 69.405 4.499 69.655 4.834 ;
      RECT 69.405 4.516 69.715 4.833 ;
      RECT 69.385 4.51 69.7 4.829 ;
      RECT 69.385 4.519 69.72 4.823 ;
      RECT 69.38 4.525 69.72 4.595 ;
      RECT 69.445 4.485 69.58 4.853 ;
      RECT 69.32 3.848 69.52 4.16 ;
      RECT 69.395 3.826 69.52 4.16 ;
      RECT 69.335 3.845 69.525 4.145 ;
      RECT 69.305 3.856 69.525 4.143 ;
      RECT 69.32 3.851 69.53 4.109 ;
      RECT 69.305 3.955 69.535 4.076 ;
      RECT 69.335 3.827 69.52 4.16 ;
      RECT 69.395 3.805 69.495 4.16 ;
      RECT 69.42 3.802 69.495 4.16 ;
      RECT 69.42 3.797 69.44 4.16 ;
      RECT 68.825 3.865 69 4.04 ;
      RECT 68.82 3.865 69 4.038 ;
      RECT 68.795 3.865 69 4.033 ;
      RECT 68.74 3.845 68.91 4.023 ;
      RECT 68.74 3.852 68.975 4.023 ;
      RECT 68.825 4.532 68.84 4.715 ;
      RECT 68.815 4.51 68.825 4.715 ;
      RECT 68.8 4.49 68.815 4.715 ;
      RECT 68.79 4.465 68.8 4.715 ;
      RECT 68.76 4.43 68.79 4.715 ;
      RECT 68.725 4.37 68.76 4.715 ;
      RECT 68.72 4.332 68.725 4.715 ;
      RECT 68.67 4.283 68.72 4.715 ;
      RECT 68.66 4.233 68.67 4.703 ;
      RECT 68.645 4.212 68.66 4.663 ;
      RECT 68.625 4.18 68.645 4.613 ;
      RECT 68.6 4.136 68.625 4.553 ;
      RECT 68.595 4.108 68.6 4.508 ;
      RECT 68.59 4.099 68.595 4.494 ;
      RECT 68.585 4.092 68.59 4.481 ;
      RECT 68.58 4.087 68.585 4.47 ;
      RECT 68.575 4.072 68.58 4.46 ;
      RECT 68.57 4.05 68.575 4.447 ;
      RECT 68.56 4.01 68.57 4.422 ;
      RECT 68.535 3.94 68.56 4.378 ;
      RECT 68.53 3.88 68.535 4.343 ;
      RECT 68.515 3.86 68.53 4.31 ;
      RECT 68.51 3.86 68.515 4.285 ;
      RECT 68.48 3.86 68.51 4.24 ;
      RECT 68.435 3.86 68.48 4.18 ;
      RECT 68.36 3.86 68.435 4.128 ;
      RECT 68.355 3.86 68.36 4.093 ;
      RECT 68.35 3.86 68.355 4.083 ;
      RECT 68.345 3.86 68.35 4.063 ;
      RECT 68.61 3.08 68.78 3.55 ;
      RECT 68.555 3.073 68.75 3.534 ;
      RECT 68.555 3.087 68.785 3.533 ;
      RECT 68.54 3.088 68.785 3.514 ;
      RECT 68.535 3.106 68.785 3.5 ;
      RECT 68.54 3.089 68.79 3.498 ;
      RECT 68.525 3.12 68.79 3.483 ;
      RECT 68.54 3.095 68.795 3.468 ;
      RECT 68.52 3.135 68.795 3.465 ;
      RECT 68.535 3.107 68.8 3.45 ;
      RECT 68.535 3.119 68.805 3.43 ;
      RECT 68.52 3.135 68.81 3.413 ;
      RECT 68.52 3.145 68.815 3.268 ;
      RECT 68.515 3.145 68.815 3.225 ;
      RECT 68.515 3.16 68.82 3.203 ;
      RECT 68.61 3.07 68.75 3.55 ;
      RECT 68.61 3.068 68.72 3.55 ;
      RECT 68.696 3.065 68.72 3.55 ;
      RECT 68.355 4.732 68.36 4.778 ;
      RECT 68.345 4.58 68.355 4.802 ;
      RECT 68.34 4.425 68.345 4.827 ;
      RECT 68.325 4.387 68.34 4.838 ;
      RECT 68.32 4.37 68.325 4.845 ;
      RECT 68.31 4.358 68.32 4.852 ;
      RECT 68.305 4.349 68.31 4.854 ;
      RECT 68.3 4.347 68.305 4.858 ;
      RECT 68.255 4.338 68.3 4.873 ;
      RECT 68.25 4.33 68.255 4.887 ;
      RECT 68.245 4.327 68.25 4.891 ;
      RECT 68.23 4.322 68.245 4.899 ;
      RECT 68.175 4.312 68.23 4.91 ;
      RECT 68.14 4.3 68.175 4.911 ;
      RECT 68.131 4.295 68.14 4.905 ;
      RECT 68.045 4.295 68.131 4.895 ;
      RECT 68.015 4.295 68.045 4.873 ;
      RECT 68.005 4.295 68.01 4.853 ;
      RECT 68 4.295 68.005 4.815 ;
      RECT 67.995 4.295 68 4.773 ;
      RECT 67.99 4.295 67.995 4.733 ;
      RECT 67.985 4.295 67.99 4.663 ;
      RECT 67.975 4.295 67.985 4.585 ;
      RECT 67.97 4.295 67.975 4.485 ;
      RECT 68.01 4.295 68.015 4.855 ;
      RECT 67.505 4.377 67.595 4.855 ;
      RECT 67.49 4.38 67.61 4.853 ;
      RECT 67.505 4.379 67.61 4.853 ;
      RECT 67.47 4.386 67.635 4.843 ;
      RECT 67.49 4.38 67.635 4.843 ;
      RECT 67.455 4.392 67.635 4.831 ;
      RECT 67.49 4.383 67.685 4.824 ;
      RECT 67.441 4.4 67.685 4.822 ;
      RECT 67.47 4.39 67.695 4.81 ;
      RECT 67.441 4.411 67.725 4.801 ;
      RECT 67.355 4.435 67.725 4.795 ;
      RECT 67.355 4.448 67.765 4.778 ;
      RECT 67.35 4.47 67.765 4.771 ;
      RECT 67.32 4.485 67.765 4.761 ;
      RECT 67.315 4.496 67.765 4.751 ;
      RECT 67.285 4.509 67.765 4.742 ;
      RECT 67.27 4.527 67.765 4.731 ;
      RECT 67.245 4.54 67.765 4.721 ;
      RECT 67.505 4.376 67.515 4.855 ;
      RECT 67.551 3.8 67.59 4.045 ;
      RECT 67.465 3.8 67.6 4.043 ;
      RECT 67.35 3.825 67.6 4.04 ;
      RECT 67.35 3.825 67.605 4.038 ;
      RECT 67.35 3.825 67.62 4.033 ;
      RECT 67.456 3.8 67.635 4.013 ;
      RECT 67.37 3.808 67.635 4.013 ;
      RECT 67.04 3.16 67.21 3.595 ;
      RECT 67.03 3.194 67.21 3.578 ;
      RECT 67.11 3.13 67.28 3.565 ;
      RECT 67.015 3.205 67.28 3.543 ;
      RECT 67.11 3.14 67.285 3.533 ;
      RECT 67.04 3.192 67.315 3.518 ;
      RECT 67 3.218 67.315 3.503 ;
      RECT 67 3.26 67.325 3.483 ;
      RECT 66.995 3.285 67.33 3.465 ;
      RECT 66.995 3.295 67.335 3.45 ;
      RECT 66.99 3.232 67.315 3.448 ;
      RECT 66.99 3.305 67.34 3.433 ;
      RECT 66.985 3.242 67.315 3.43 ;
      RECT 66.98 3.326 67.345 3.413 ;
      RECT 66.98 3.358 67.35 3.393 ;
      RECT 66.975 3.272 67.325 3.385 ;
      RECT 66.98 3.257 67.315 3.413 ;
      RECT 66.995 3.227 67.315 3.465 ;
      RECT 66.84 3.814 67.065 4.07 ;
      RECT 66.84 3.847 67.085 4.06 ;
      RECT 66.805 3.847 67.085 4.058 ;
      RECT 66.805 3.86 67.09 4.048 ;
      RECT 66.805 3.88 67.1 4.04 ;
      RECT 66.805 3.977 67.105 4.033 ;
      RECT 66.785 3.725 66.915 4.023 ;
      RECT 66.74 3.88 67.1 3.965 ;
      RECT 66.73 3.725 66.915 3.91 ;
      RECT 66.73 3.757 67.001 3.91 ;
      RECT 66.695 4.287 66.715 4.465 ;
      RECT 66.66 4.24 66.695 4.465 ;
      RECT 66.645 4.18 66.66 4.465 ;
      RECT 66.62 4.127 66.645 4.465 ;
      RECT 66.605 4.08 66.62 4.465 ;
      RECT 66.585 4.057 66.605 4.465 ;
      RECT 66.56 4.022 66.585 4.465 ;
      RECT 66.55 3.868 66.56 4.465 ;
      RECT 66.52 3.863 66.55 4.456 ;
      RECT 66.515 3.86 66.52 4.446 ;
      RECT 66.5 3.86 66.515 4.42 ;
      RECT 66.495 3.86 66.5 4.383 ;
      RECT 66.47 3.86 66.495 4.335 ;
      RECT 66.45 3.86 66.47 4.26 ;
      RECT 66.44 3.86 66.45 4.22 ;
      RECT 66.435 3.86 66.44 4.195 ;
      RECT 66.43 3.86 66.435 4.178 ;
      RECT 66.425 3.86 66.43 4.16 ;
      RECT 66.42 3.861 66.425 4.15 ;
      RECT 66.41 3.863 66.42 4.118 ;
      RECT 66.4 3.865 66.41 4.085 ;
      RECT 66.39 3.868 66.4 4.058 ;
      RECT 66.715 4.295 66.94 4.465 ;
      RECT 66.045 3.107 66.215 3.56 ;
      RECT 66.045 3.107 66.305 3.526 ;
      RECT 66.045 3.107 66.335 3.51 ;
      RECT 66.045 3.107 66.365 3.483 ;
      RECT 66.301 3.085 66.38 3.465 ;
      RECT 66.08 3.092 66.385 3.45 ;
      RECT 66.08 3.1 66.395 3.413 ;
      RECT 66.04 3.127 66.395 3.385 ;
      RECT 66.025 3.14 66.395 3.35 ;
      RECT 66.045 3.115 66.415 3.34 ;
      RECT 66.02 3.18 66.415 3.31 ;
      RECT 66.02 3.21 66.42 3.293 ;
      RECT 66.015 3.24 66.42 3.28 ;
      RECT 66.08 3.089 66.38 3.465 ;
      RECT 66.215 3.086 66.301 3.544 ;
      RECT 66.166 3.087 66.38 3.465 ;
      RECT 66.31 4.747 66.355 4.94 ;
      RECT 66.3 4.717 66.31 4.94 ;
      RECT 66.295 4.702 66.3 4.94 ;
      RECT 66.255 4.612 66.295 4.94 ;
      RECT 66.25 4.525 66.255 4.94 ;
      RECT 66.24 4.495 66.25 4.94 ;
      RECT 66.235 4.455 66.24 4.94 ;
      RECT 66.225 4.417 66.235 4.94 ;
      RECT 66.22 4.382 66.225 4.94 ;
      RECT 66.2 4.335 66.22 4.94 ;
      RECT 66.185 4.26 66.2 4.94 ;
      RECT 66.18 4.215 66.185 4.935 ;
      RECT 66.175 4.195 66.18 4.908 ;
      RECT 66.17 4.175 66.175 4.893 ;
      RECT 66.165 4.15 66.17 4.873 ;
      RECT 66.16 4.128 66.165 4.858 ;
      RECT 66.155 4.106 66.16 4.84 ;
      RECT 66.15 4.085 66.155 4.83 ;
      RECT 66.14 4.057 66.15 4.8 ;
      RECT 66.13 4.02 66.14 4.768 ;
      RECT 66.12 3.98 66.13 4.735 ;
      RECT 66.11 3.958 66.12 4.705 ;
      RECT 66.08 3.91 66.11 4.637 ;
      RECT 66.065 3.87 66.08 4.564 ;
      RECT 66.055 3.87 66.065 4.53 ;
      RECT 66.05 3.87 66.055 4.505 ;
      RECT 66.045 3.87 66.05 4.49 ;
      RECT 66.04 3.87 66.045 4.468 ;
      RECT 66.035 3.87 66.04 4.455 ;
      RECT 66.02 3.87 66.035 4.42 ;
      RECT 66 3.87 66.02 4.36 ;
      RECT 65.99 3.87 66 4.31 ;
      RECT 65.97 3.87 65.99 4.258 ;
      RECT 65.95 3.87 65.97 4.215 ;
      RECT 65.94 3.87 65.95 4.203 ;
      RECT 65.91 3.87 65.94 4.19 ;
      RECT 65.88 3.891 65.91 4.17 ;
      RECT 65.87 3.919 65.88 4.15 ;
      RECT 65.855 3.936 65.87 4.118 ;
      RECT 65.85 3.95 65.855 4.085 ;
      RECT 65.845 3.958 65.85 4.058 ;
      RECT 65.84 3.966 65.845 4.02 ;
      RECT 65.845 4.49 65.85 4.825 ;
      RECT 65.81 4.477 65.845 4.824 ;
      RECT 65.74 4.417 65.81 4.823 ;
      RECT 65.66 4.36 65.74 4.822 ;
      RECT 65.525 4.32 65.66 4.821 ;
      RECT 65.525 4.507 65.86 4.81 ;
      RECT 65.485 4.507 65.86 4.8 ;
      RECT 65.485 4.525 65.865 4.795 ;
      RECT 65.485 4.615 65.87 4.785 ;
      RECT 65.48 4.31 65.645 4.765 ;
      RECT 65.475 4.31 65.645 4.508 ;
      RECT 65.475 4.467 65.84 4.508 ;
      RECT 65.475 4.455 65.835 4.508 ;
      RECT 64.61 7.3 64.78 8.77 ;
      RECT 64.61 7.3 64.785 8.56 ;
      RECT 64.24 9.25 64.71 9.42 ;
      RECT 64.24 8.23 64.41 9.42 ;
      RECT 64.235 3.04 64.405 4.23 ;
      RECT 64.235 3.04 64.705 3.21 ;
      RECT 63.615 3.895 63.79 5.155 ;
      RECT 63.615 3.685 63.785 5.155 ;
      RECT 63.615 7.305 63.785 8.775 ;
      RECT 63.615 7.305 63.79 8.565 ;
      RECT 63.245 3.035 63.415 4.225 ;
      RECT 63.245 3.035 63.715 3.205 ;
      RECT 63.245 9.255 63.715 9.425 ;
      RECT 63.245 8.235 63.415 9.425 ;
      RECT 62.255 4.015 62.43 5.155 ;
      RECT 62.255 1.865 62.425 5.155 ;
      RECT 62.255 1.865 62.43 2.415 ;
      RECT 62.255 10.045 62.43 10.595 ;
      RECT 62.255 7.305 62.425 10.595 ;
      RECT 62.255 7.305 62.43 8.445 ;
      RECT 61.825 3.895 62 5.155 ;
      RECT 61.825 2.945 61.995 5.155 ;
      RECT 61.825 7.305 61.995 9.515 ;
      RECT 61.825 7.305 62 8.565 ;
      RECT 61.395 3.925 61.565 5.155 ;
      RECT 61.455 2.145 61.625 4.095 ;
      RECT 61.395 1.865 61.565 2.315 ;
      RECT 61.395 10.145 61.565 10.595 ;
      RECT 61.455 8.365 61.625 10.315 ;
      RECT 61.395 7.305 61.565 8.535 ;
      RECT 60.87 3.895 61.045 5.155 ;
      RECT 60.87 1.865 61.04 5.155 ;
      RECT 60.87 3.365 61.28 3.695 ;
      RECT 60.87 2.525 61.28 2.855 ;
      RECT 60.87 1.865 61.045 2.355 ;
      RECT 60.87 10.105 61.045 10.595 ;
      RECT 60.87 7.305 61.04 10.595 ;
      RECT 60.87 9.605 61.28 9.935 ;
      RECT 60.87 8.765 61.28 9.095 ;
      RECT 60.87 7.305 61.045 8.565 ;
      RECT 58.21 3.27 58.94 3.51 ;
      RECT 58.752 3.065 58.94 3.51 ;
      RECT 58.58 3.077 58.955 3.504 ;
      RECT 58.495 3.092 58.975 3.489 ;
      RECT 58.495 3.107 58.98 3.479 ;
      RECT 58.45 3.127 58.995 3.471 ;
      RECT 58.427 3.162 59.01 3.425 ;
      RECT 58.341 3.185 59.015 3.385 ;
      RECT 58.341 3.203 59.025 3.355 ;
      RECT 58.21 3.272 59.03 3.318 ;
      RECT 58.255 3.215 59.025 3.355 ;
      RECT 58.341 3.167 59.01 3.425 ;
      RECT 58.427 3.136 58.995 3.471 ;
      RECT 58.45 3.117 58.98 3.479 ;
      RECT 58.495 3.09 58.955 3.504 ;
      RECT 58.58 3.072 58.94 3.51 ;
      RECT 58.666 3.066 58.94 3.51 ;
      RECT 58.752 3.061 58.885 3.51 ;
      RECT 58.838 3.056 58.885 3.51 ;
      RECT 58.4 4.67 58.405 4.683 ;
      RECT 58.395 4.565 58.4 4.688 ;
      RECT 58.37 4.425 58.395 4.703 ;
      RECT 58.335 4.376 58.37 4.735 ;
      RECT 58.33 4.344 58.335 4.755 ;
      RECT 58.325 4.335 58.33 4.755 ;
      RECT 58.245 4.3 58.325 4.755 ;
      RECT 58.182 4.27 58.245 4.755 ;
      RECT 58.096 4.258 58.182 4.755 ;
      RECT 58.01 4.244 58.096 4.755 ;
      RECT 57.93 4.231 58.01 4.741 ;
      RECT 57.895 4.223 57.93 4.721 ;
      RECT 57.885 4.22 57.895 4.712 ;
      RECT 57.855 4.215 57.885 4.699 ;
      RECT 57.805 4.19 57.855 4.675 ;
      RECT 57.791 4.164 57.805 4.657 ;
      RECT 57.705 4.124 57.791 4.633 ;
      RECT 57.66 4.072 57.705 4.602 ;
      RECT 57.65 4.047 57.66 4.589 ;
      RECT 57.645 3.828 57.65 3.85 ;
      RECT 57.64 4.03 57.65 4.585 ;
      RECT 57.64 3.826 57.645 3.94 ;
      RECT 57.63 3.822 57.64 4.581 ;
      RECT 57.586 3.82 57.63 4.569 ;
      RECT 57.5 3.82 57.586 4.54 ;
      RECT 57.47 3.82 57.5 4.513 ;
      RECT 57.455 3.82 57.47 4.501 ;
      RECT 57.415 3.832 57.455 4.486 ;
      RECT 57.395 3.851 57.415 4.465 ;
      RECT 57.385 3.861 57.395 4.449 ;
      RECT 57.375 3.867 57.385 4.438 ;
      RECT 57.355 3.877 57.375 4.421 ;
      RECT 57.35 3.886 57.355 4.408 ;
      RECT 57.345 3.89 57.35 4.358 ;
      RECT 57.335 3.896 57.345 4.275 ;
      RECT 57.33 3.9 57.335 4.189 ;
      RECT 57.325 3.92 57.33 4.126 ;
      RECT 57.32 3.943 57.325 4.073 ;
      RECT 57.315 3.961 57.32 4.018 ;
      RECT 57.925 3.78 58.095 4.04 ;
      RECT 58.095 3.745 58.14 4.026 ;
      RECT 58.056 3.747 58.145 4.009 ;
      RECT 57.945 3.764 58.231 3.98 ;
      RECT 57.945 3.779 58.235 3.952 ;
      RECT 57.945 3.76 58.145 4.009 ;
      RECT 57.97 3.748 58.095 4.04 ;
      RECT 58.056 3.746 58.14 4.026 ;
      RECT 57.475 10.045 57.65 10.595 ;
      RECT 57.475 7.305 57.645 10.595 ;
      RECT 57.475 7.305 57.65 8.445 ;
      RECT 57.11 3.135 57.28 3.625 ;
      RECT 57.11 3.135 57.315 3.605 ;
      RECT 57.245 3.055 57.355 3.565 ;
      RECT 57.226 3.059 57.375 3.535 ;
      RECT 57.14 3.067 57.395 3.518 ;
      RECT 57.14 3.073 57.4 3.508 ;
      RECT 57.14 3.082 57.42 3.496 ;
      RECT 57.115 3.107 57.45 3.474 ;
      RECT 57.115 3.127 57.455 3.454 ;
      RECT 57.11 3.14 57.465 3.434 ;
      RECT 57.11 3.207 57.47 3.415 ;
      RECT 57.11 3.34 57.475 3.402 ;
      RECT 57.105 3.145 57.465 3.235 ;
      RECT 57.115 3.102 57.42 3.496 ;
      RECT 57.226 3.057 57.355 3.565 ;
      RECT 57.1 4.81 57.4 5.065 ;
      RECT 57.185 4.776 57.4 5.065 ;
      RECT 57.185 4.779 57.405 4.925 ;
      RECT 57.12 4.8 57.405 4.925 ;
      RECT 57.155 4.79 57.4 5.065 ;
      RECT 57.15 4.795 57.405 4.925 ;
      RECT 57.185 4.774 57.386 5.065 ;
      RECT 57.271 4.765 57.386 5.065 ;
      RECT 57.271 4.759 57.3 5.065 ;
      RECT 57.045 7.305 57.215 9.515 ;
      RECT 57.045 7.305 57.22 8.565 ;
      RECT 56.76 4.4 56.77 4.89 ;
      RECT 56.42 4.335 56.43 4.635 ;
      RECT 56.935 4.507 56.94 4.726 ;
      RECT 56.925 4.487 56.935 4.743 ;
      RECT 56.915 4.467 56.925 4.773 ;
      RECT 56.91 4.457 56.915 4.788 ;
      RECT 56.905 4.453 56.91 4.793 ;
      RECT 56.89 4.445 56.905 4.8 ;
      RECT 56.85 4.425 56.89 4.825 ;
      RECT 56.825 4.407 56.85 4.858 ;
      RECT 56.82 4.405 56.825 4.871 ;
      RECT 56.8 4.402 56.82 4.875 ;
      RECT 56.77 4.4 56.8 4.885 ;
      RECT 56.7 4.402 56.76 4.886 ;
      RECT 56.68 4.402 56.7 4.88 ;
      RECT 56.655 4.4 56.68 4.877 ;
      RECT 56.62 4.395 56.655 4.873 ;
      RECT 56.6 4.389 56.62 4.86 ;
      RECT 56.59 4.386 56.6 4.848 ;
      RECT 56.57 4.383 56.59 4.833 ;
      RECT 56.55 4.379 56.57 4.815 ;
      RECT 56.545 4.376 56.55 4.805 ;
      RECT 56.54 4.375 56.545 4.803 ;
      RECT 56.53 4.372 56.54 4.795 ;
      RECT 56.52 4.366 56.53 4.778 ;
      RECT 56.51 4.36 56.52 4.76 ;
      RECT 56.5 4.354 56.51 4.748 ;
      RECT 56.49 4.348 56.5 4.728 ;
      RECT 56.485 4.344 56.49 4.713 ;
      RECT 56.48 4.342 56.485 4.705 ;
      RECT 56.475 4.34 56.48 4.698 ;
      RECT 56.47 4.338 56.475 4.688 ;
      RECT 56.465 4.336 56.47 4.682 ;
      RECT 56.455 4.335 56.465 4.672 ;
      RECT 56.445 4.335 56.455 4.663 ;
      RECT 56.43 4.335 56.445 4.648 ;
      RECT 56.39 4.335 56.42 4.632 ;
      RECT 56.37 4.337 56.39 4.627 ;
      RECT 56.365 4.342 56.37 4.625 ;
      RECT 56.335 4.35 56.365 4.623 ;
      RECT 56.305 4.365 56.335 4.622 ;
      RECT 56.26 4.387 56.305 4.627 ;
      RECT 56.255 4.402 56.26 4.631 ;
      RECT 56.24 4.407 56.255 4.633 ;
      RECT 56.235 4.411 56.24 4.635 ;
      RECT 56.175 4.434 56.235 4.644 ;
      RECT 56.155 4.46 56.175 4.657 ;
      RECT 56.145 4.467 56.155 4.661 ;
      RECT 56.13 4.474 56.145 4.664 ;
      RECT 56.11 4.484 56.13 4.667 ;
      RECT 56.105 4.492 56.11 4.67 ;
      RECT 56.06 4.497 56.105 4.677 ;
      RECT 56.05 4.5 56.06 4.684 ;
      RECT 56.04 4.5 56.05 4.688 ;
      RECT 56.005 4.502 56.04 4.7 ;
      RECT 55.985 4.505 56.005 4.713 ;
      RECT 55.945 4.508 55.985 4.724 ;
      RECT 55.93 4.51 55.945 4.737 ;
      RECT 55.92 4.51 55.93 4.742 ;
      RECT 55.895 4.511 55.92 4.75 ;
      RECT 55.885 4.513 55.895 4.755 ;
      RECT 55.88 4.514 55.885 4.758 ;
      RECT 55.855 4.512 55.88 4.761 ;
      RECT 55.84 4.51 55.855 4.762 ;
      RECT 55.82 4.507 55.84 4.764 ;
      RECT 55.8 4.502 55.82 4.764 ;
      RECT 55.74 4.497 55.8 4.761 ;
      RECT 55.705 4.472 55.74 4.757 ;
      RECT 55.695 4.449 55.705 4.755 ;
      RECT 55.665 4.426 55.695 4.755 ;
      RECT 55.655 4.405 55.665 4.755 ;
      RECT 55.63 4.387 55.655 4.753 ;
      RECT 55.615 4.365 55.63 4.75 ;
      RECT 55.6 4.347 55.615 4.748 ;
      RECT 55.58 4.337 55.6 4.746 ;
      RECT 55.565 4.332 55.58 4.745 ;
      RECT 55.55 4.33 55.565 4.744 ;
      RECT 55.52 4.331 55.55 4.742 ;
      RECT 55.5 4.334 55.52 4.74 ;
      RECT 55.443 4.338 55.5 4.74 ;
      RECT 55.357 4.347 55.443 4.74 ;
      RECT 55.271 4.358 55.357 4.74 ;
      RECT 55.185 4.369 55.271 4.74 ;
      RECT 55.165 4.376 55.185 4.748 ;
      RECT 55.155 4.379 55.165 4.755 ;
      RECT 55.09 4.384 55.155 4.773 ;
      RECT 55.06 4.391 55.09 4.798 ;
      RECT 55.05 4.394 55.06 4.805 ;
      RECT 55.005 4.398 55.05 4.81 ;
      RECT 54.975 4.403 55.005 4.815 ;
      RECT 54.974 4.405 54.975 4.815 ;
      RECT 54.888 4.411 54.974 4.815 ;
      RECT 54.802 4.422 54.888 4.815 ;
      RECT 54.716 4.434 54.802 4.815 ;
      RECT 54.63 4.445 54.716 4.815 ;
      RECT 54.615 4.452 54.63 4.81 ;
      RECT 54.61 4.454 54.615 4.804 ;
      RECT 54.59 4.465 54.61 4.799 ;
      RECT 54.58 4.483 54.59 4.793 ;
      RECT 54.575 4.495 54.58 4.593 ;
      RECT 56.87 3.248 56.89 3.335 ;
      RECT 56.865 3.183 56.87 3.367 ;
      RECT 56.855 3.15 56.865 3.372 ;
      RECT 56.85 3.13 56.855 3.378 ;
      RECT 56.82 3.13 56.85 3.395 ;
      RECT 56.771 3.13 56.82 3.431 ;
      RECT 56.685 3.13 56.771 3.489 ;
      RECT 56.656 3.14 56.685 3.538 ;
      RECT 56.57 3.182 56.656 3.591 ;
      RECT 56.55 3.22 56.57 3.638 ;
      RECT 56.525 3.237 56.55 3.658 ;
      RECT 56.515 3.251 56.525 3.678 ;
      RECT 56.51 3.257 56.515 3.688 ;
      RECT 56.505 3.261 56.51 3.695 ;
      RECT 56.455 3.281 56.505 3.7 ;
      RECT 56.39 3.325 56.455 3.7 ;
      RECT 56.365 3.375 56.39 3.7 ;
      RECT 56.355 3.405 56.365 3.7 ;
      RECT 56.35 3.432 56.355 3.7 ;
      RECT 56.345 3.45 56.35 3.7 ;
      RECT 56.335 3.492 56.345 3.7 ;
      RECT 56.09 10.105 56.265 10.595 ;
      RECT 56.09 7.305 56.26 10.595 ;
      RECT 56.09 9.605 56.5 9.935 ;
      RECT 56.09 8.765 56.5 9.095 ;
      RECT 56.09 7.305 56.265 8.565 ;
      RECT 56.165 4.85 56.355 5.075 ;
      RECT 56.155 4.851 56.36 5.07 ;
      RECT 56.155 4.853 56.37 5.05 ;
      RECT 56.155 4.857 56.375 5.035 ;
      RECT 56.155 4.844 56.325 5.07 ;
      RECT 56.155 4.847 56.35 5.07 ;
      RECT 56.165 4.843 56.325 5.075 ;
      RECT 56.251 4.841 56.325 5.075 ;
      RECT 55.875 4.092 56.045 4.33 ;
      RECT 55.875 4.092 56.131 4.244 ;
      RECT 55.875 4.092 56.135 4.154 ;
      RECT 55.925 3.865 56.145 4.133 ;
      RECT 55.92 3.882 56.15 4.106 ;
      RECT 55.885 4.04 56.15 4.106 ;
      RECT 55.905 3.89 56.045 4.33 ;
      RECT 55.895 3.972 56.155 4.089 ;
      RECT 55.89 4.02 56.155 4.089 ;
      RECT 55.895 3.93 56.15 4.106 ;
      RECT 55.92 3.867 56.145 4.133 ;
      RECT 55.485 3.842 55.655 4.04 ;
      RECT 55.485 3.842 55.7 4.015 ;
      RECT 55.555 3.785 55.725 3.973 ;
      RECT 55.53 3.8 55.725 3.973 ;
      RECT 55.145 3.846 55.175 4.04 ;
      RECT 55.14 3.818 55.145 4.04 ;
      RECT 55.11 3.792 55.14 4.042 ;
      RECT 55.085 3.75 55.11 4.045 ;
      RECT 55.075 3.722 55.085 4.047 ;
      RECT 55.04 3.702 55.075 4.049 ;
      RECT 54.975 3.687 55.04 4.055 ;
      RECT 54.925 3.685 54.975 4.061 ;
      RECT 54.902 3.687 54.925 4.066 ;
      RECT 54.816 3.698 54.902 4.072 ;
      RECT 54.73 3.716 54.816 4.082 ;
      RECT 54.715 3.727 54.73 4.088 ;
      RECT 54.645 3.75 54.715 4.094 ;
      RECT 54.59 3.782 54.645 4.102 ;
      RECT 54.55 3.805 54.59 4.108 ;
      RECT 54.536 3.818 54.55 4.111 ;
      RECT 54.45 3.84 54.536 4.117 ;
      RECT 54.435 3.865 54.45 4.123 ;
      RECT 54.395 3.88 54.435 4.127 ;
      RECT 54.345 3.895 54.395 4.132 ;
      RECT 54.32 3.902 54.345 4.136 ;
      RECT 54.26 3.897 54.32 4.14 ;
      RECT 54.245 3.888 54.26 4.144 ;
      RECT 54.175 3.878 54.245 4.14 ;
      RECT 54.15 3.87 54.17 4.13 ;
      RECT 54.091 3.87 54.15 4.108 ;
      RECT 54.005 3.87 54.091 4.065 ;
      RECT 54.17 3.87 54.175 4.135 ;
      RECT 54.865 3.101 55.035 3.435 ;
      RECT 54.835 3.101 55.035 3.43 ;
      RECT 54.775 3.068 54.835 3.418 ;
      RECT 54.775 3.124 55.045 3.413 ;
      RECT 54.75 3.124 55.045 3.407 ;
      RECT 54.745 3.065 54.775 3.404 ;
      RECT 54.73 3.071 54.865 3.402 ;
      RECT 54.725 3.079 54.95 3.39 ;
      RECT 54.725 3.131 55.06 3.343 ;
      RECT 54.71 3.087 54.95 3.338 ;
      RECT 54.71 3.157 55.07 3.279 ;
      RECT 54.68 3.107 55.035 3.24 ;
      RECT 54.68 3.197 55.08 3.236 ;
      RECT 54.73 3.076 54.95 3.402 ;
      RECT 54.07 3.406 54.125 3.67 ;
      RECT 54.07 3.406 54.19 3.669 ;
      RECT 54.07 3.406 54.215 3.668 ;
      RECT 54.07 3.406 54.28 3.667 ;
      RECT 54.215 3.372 54.295 3.666 ;
      RECT 54.03 3.416 54.44 3.665 ;
      RECT 54.07 3.413 54.44 3.665 ;
      RECT 54.03 3.421 54.445 3.658 ;
      RECT 54.015 3.423 54.445 3.657 ;
      RECT 54.015 3.43 54.45 3.653 ;
      RECT 53.995 3.429 54.445 3.649 ;
      RECT 53.995 3.437 54.455 3.648 ;
      RECT 53.99 3.434 54.45 3.644 ;
      RECT 53.99 3.447 54.465 3.643 ;
      RECT 53.975 3.437 54.455 3.642 ;
      RECT 53.94 3.45 54.465 3.635 ;
      RECT 54.125 3.405 54.435 3.665 ;
      RECT 54.125 3.39 54.385 3.665 ;
      RECT 54.19 3.377 54.32 3.665 ;
      RECT 53.735 4.466 53.75 4.859 ;
      RECT 53.7 4.471 53.75 4.858 ;
      RECT 53.735 4.47 53.795 4.857 ;
      RECT 53.68 4.481 53.795 4.856 ;
      RECT 53.695 4.477 53.795 4.856 ;
      RECT 53.66 4.487 53.87 4.853 ;
      RECT 53.66 4.506 53.915 4.851 ;
      RECT 53.66 4.513 53.92 4.848 ;
      RECT 53.645 4.49 53.87 4.845 ;
      RECT 53.625 4.495 53.87 4.838 ;
      RECT 53.62 4.499 53.87 4.834 ;
      RECT 53.62 4.516 53.93 4.833 ;
      RECT 53.6 4.51 53.915 4.829 ;
      RECT 53.6 4.519 53.935 4.823 ;
      RECT 53.595 4.525 53.935 4.595 ;
      RECT 53.66 4.485 53.795 4.853 ;
      RECT 53.535 3.848 53.735 4.16 ;
      RECT 53.61 3.826 53.735 4.16 ;
      RECT 53.55 3.845 53.74 4.145 ;
      RECT 53.52 3.856 53.74 4.143 ;
      RECT 53.535 3.851 53.745 4.109 ;
      RECT 53.52 3.955 53.75 4.076 ;
      RECT 53.55 3.827 53.735 4.16 ;
      RECT 53.61 3.805 53.71 4.16 ;
      RECT 53.635 3.802 53.71 4.16 ;
      RECT 53.635 3.797 53.655 4.16 ;
      RECT 53.04 3.865 53.215 4.04 ;
      RECT 53.035 3.865 53.215 4.038 ;
      RECT 53.01 3.865 53.215 4.033 ;
      RECT 52.955 3.845 53.125 4.023 ;
      RECT 52.955 3.852 53.19 4.023 ;
      RECT 53.04 4.532 53.055 4.715 ;
      RECT 53.03 4.51 53.04 4.715 ;
      RECT 53.015 4.49 53.03 4.715 ;
      RECT 53.005 4.465 53.015 4.715 ;
      RECT 52.975 4.43 53.005 4.715 ;
      RECT 52.94 4.37 52.975 4.715 ;
      RECT 52.935 4.332 52.94 4.715 ;
      RECT 52.885 4.283 52.935 4.715 ;
      RECT 52.875 4.233 52.885 4.703 ;
      RECT 52.86 4.212 52.875 4.663 ;
      RECT 52.84 4.18 52.86 4.613 ;
      RECT 52.815 4.136 52.84 4.553 ;
      RECT 52.81 4.108 52.815 4.508 ;
      RECT 52.805 4.099 52.81 4.494 ;
      RECT 52.8 4.092 52.805 4.481 ;
      RECT 52.795 4.087 52.8 4.47 ;
      RECT 52.79 4.072 52.795 4.46 ;
      RECT 52.785 4.05 52.79 4.447 ;
      RECT 52.775 4.01 52.785 4.422 ;
      RECT 52.75 3.94 52.775 4.378 ;
      RECT 52.745 3.88 52.75 4.343 ;
      RECT 52.73 3.86 52.745 4.31 ;
      RECT 52.725 3.86 52.73 4.285 ;
      RECT 52.695 3.86 52.725 4.24 ;
      RECT 52.65 3.86 52.695 4.18 ;
      RECT 52.575 3.86 52.65 4.128 ;
      RECT 52.57 3.86 52.575 4.093 ;
      RECT 52.565 3.86 52.57 4.083 ;
      RECT 52.56 3.86 52.565 4.063 ;
      RECT 52.825 3.08 52.995 3.55 ;
      RECT 52.77 3.073 52.965 3.534 ;
      RECT 52.77 3.087 53 3.533 ;
      RECT 52.755 3.088 53 3.514 ;
      RECT 52.75 3.106 53 3.5 ;
      RECT 52.755 3.089 53.005 3.498 ;
      RECT 52.74 3.12 53.005 3.483 ;
      RECT 52.755 3.095 53.01 3.468 ;
      RECT 52.735 3.135 53.01 3.465 ;
      RECT 52.75 3.107 53.015 3.45 ;
      RECT 52.75 3.119 53.02 3.43 ;
      RECT 52.735 3.135 53.025 3.413 ;
      RECT 52.735 3.145 53.03 3.268 ;
      RECT 52.73 3.145 53.03 3.225 ;
      RECT 52.73 3.16 53.035 3.203 ;
      RECT 52.825 3.07 52.965 3.55 ;
      RECT 52.825 3.068 52.935 3.55 ;
      RECT 52.911 3.065 52.935 3.55 ;
      RECT 52.57 4.732 52.575 4.778 ;
      RECT 52.56 4.58 52.57 4.802 ;
      RECT 52.555 4.425 52.56 4.827 ;
      RECT 52.54 4.387 52.555 4.838 ;
      RECT 52.535 4.37 52.54 4.845 ;
      RECT 52.525 4.358 52.535 4.852 ;
      RECT 52.52 4.349 52.525 4.854 ;
      RECT 52.515 4.347 52.52 4.858 ;
      RECT 52.47 4.338 52.515 4.873 ;
      RECT 52.465 4.33 52.47 4.887 ;
      RECT 52.46 4.327 52.465 4.891 ;
      RECT 52.445 4.322 52.46 4.899 ;
      RECT 52.39 4.312 52.445 4.91 ;
      RECT 52.355 4.3 52.39 4.911 ;
      RECT 52.346 4.295 52.355 4.905 ;
      RECT 52.26 4.295 52.346 4.895 ;
      RECT 52.23 4.295 52.26 4.873 ;
      RECT 52.22 4.295 52.225 4.853 ;
      RECT 52.215 4.295 52.22 4.815 ;
      RECT 52.21 4.295 52.215 4.773 ;
      RECT 52.205 4.295 52.21 4.733 ;
      RECT 52.2 4.295 52.205 4.663 ;
      RECT 52.19 4.295 52.2 4.585 ;
      RECT 52.185 4.295 52.19 4.485 ;
      RECT 52.225 4.295 52.23 4.855 ;
      RECT 51.72 4.377 51.81 4.855 ;
      RECT 51.705 4.38 51.825 4.853 ;
      RECT 51.72 4.379 51.825 4.853 ;
      RECT 51.685 4.386 51.85 4.843 ;
      RECT 51.705 4.38 51.85 4.843 ;
      RECT 51.67 4.392 51.85 4.831 ;
      RECT 51.705 4.383 51.9 4.824 ;
      RECT 51.656 4.4 51.9 4.822 ;
      RECT 51.685 4.39 51.91 4.81 ;
      RECT 51.656 4.411 51.94 4.801 ;
      RECT 51.57 4.435 51.94 4.795 ;
      RECT 51.57 4.448 51.98 4.778 ;
      RECT 51.565 4.47 51.98 4.771 ;
      RECT 51.535 4.485 51.98 4.761 ;
      RECT 51.53 4.496 51.98 4.751 ;
      RECT 51.5 4.509 51.98 4.742 ;
      RECT 51.485 4.527 51.98 4.731 ;
      RECT 51.46 4.54 51.98 4.721 ;
      RECT 51.72 4.376 51.73 4.855 ;
      RECT 51.766 3.8 51.805 4.045 ;
      RECT 51.68 3.8 51.815 4.043 ;
      RECT 51.565 3.825 51.815 4.04 ;
      RECT 51.565 3.825 51.82 4.038 ;
      RECT 51.565 3.825 51.835 4.033 ;
      RECT 51.671 3.8 51.85 4.013 ;
      RECT 51.585 3.808 51.85 4.013 ;
      RECT 51.255 3.16 51.425 3.595 ;
      RECT 51.245 3.194 51.425 3.578 ;
      RECT 51.325 3.13 51.495 3.565 ;
      RECT 51.23 3.205 51.495 3.543 ;
      RECT 51.325 3.14 51.5 3.533 ;
      RECT 51.255 3.192 51.53 3.518 ;
      RECT 51.215 3.218 51.53 3.503 ;
      RECT 51.215 3.26 51.54 3.483 ;
      RECT 51.21 3.285 51.545 3.465 ;
      RECT 51.21 3.295 51.55 3.45 ;
      RECT 51.205 3.232 51.53 3.448 ;
      RECT 51.205 3.305 51.555 3.433 ;
      RECT 51.2 3.242 51.53 3.43 ;
      RECT 51.195 3.326 51.56 3.413 ;
      RECT 51.195 3.358 51.565 3.393 ;
      RECT 51.19 3.272 51.54 3.385 ;
      RECT 51.195 3.257 51.53 3.413 ;
      RECT 51.21 3.227 51.53 3.465 ;
      RECT 51.055 3.814 51.28 4.07 ;
      RECT 51.055 3.847 51.3 4.06 ;
      RECT 51.02 3.847 51.3 4.058 ;
      RECT 51.02 3.86 51.305 4.048 ;
      RECT 51.02 3.88 51.315 4.04 ;
      RECT 51.02 3.977 51.32 4.033 ;
      RECT 51 3.725 51.13 4.023 ;
      RECT 50.955 3.88 51.315 3.965 ;
      RECT 50.945 3.725 51.13 3.91 ;
      RECT 50.945 3.757 51.216 3.91 ;
      RECT 50.91 4.287 50.93 4.465 ;
      RECT 50.875 4.24 50.91 4.465 ;
      RECT 50.86 4.18 50.875 4.465 ;
      RECT 50.835 4.127 50.86 4.465 ;
      RECT 50.82 4.08 50.835 4.465 ;
      RECT 50.8 4.057 50.82 4.465 ;
      RECT 50.775 4.022 50.8 4.465 ;
      RECT 50.765 3.868 50.775 4.465 ;
      RECT 50.735 3.863 50.765 4.456 ;
      RECT 50.73 3.86 50.735 4.446 ;
      RECT 50.715 3.86 50.73 4.42 ;
      RECT 50.71 3.86 50.715 4.383 ;
      RECT 50.685 3.86 50.71 4.335 ;
      RECT 50.665 3.86 50.685 4.26 ;
      RECT 50.655 3.86 50.665 4.22 ;
      RECT 50.65 3.86 50.655 4.195 ;
      RECT 50.645 3.86 50.65 4.178 ;
      RECT 50.64 3.86 50.645 4.16 ;
      RECT 50.635 3.861 50.64 4.15 ;
      RECT 50.625 3.863 50.635 4.118 ;
      RECT 50.615 3.865 50.625 4.085 ;
      RECT 50.605 3.868 50.615 4.058 ;
      RECT 50.93 4.295 51.155 4.465 ;
      RECT 50.26 3.107 50.43 3.56 ;
      RECT 50.26 3.107 50.52 3.526 ;
      RECT 50.26 3.107 50.55 3.51 ;
      RECT 50.26 3.107 50.58 3.483 ;
      RECT 50.516 3.085 50.595 3.465 ;
      RECT 50.295 3.092 50.6 3.45 ;
      RECT 50.295 3.1 50.61 3.413 ;
      RECT 50.255 3.127 50.61 3.385 ;
      RECT 50.24 3.14 50.61 3.35 ;
      RECT 50.26 3.115 50.63 3.34 ;
      RECT 50.235 3.18 50.63 3.31 ;
      RECT 50.235 3.21 50.635 3.293 ;
      RECT 50.23 3.24 50.635 3.28 ;
      RECT 50.295 3.089 50.595 3.465 ;
      RECT 50.43 3.086 50.516 3.544 ;
      RECT 50.381 3.087 50.595 3.465 ;
      RECT 50.525 4.747 50.57 4.94 ;
      RECT 50.515 4.717 50.525 4.94 ;
      RECT 50.51 4.702 50.515 4.94 ;
      RECT 50.47 4.612 50.51 4.94 ;
      RECT 50.465 4.525 50.47 4.94 ;
      RECT 50.455 4.495 50.465 4.94 ;
      RECT 50.45 4.455 50.455 4.94 ;
      RECT 50.44 4.417 50.45 4.94 ;
      RECT 50.435 4.382 50.44 4.94 ;
      RECT 50.415 4.335 50.435 4.94 ;
      RECT 50.4 4.26 50.415 4.94 ;
      RECT 50.395 4.215 50.4 4.935 ;
      RECT 50.39 4.195 50.395 4.908 ;
      RECT 50.385 4.175 50.39 4.893 ;
      RECT 50.38 4.15 50.385 4.873 ;
      RECT 50.375 4.128 50.38 4.858 ;
      RECT 50.37 4.106 50.375 4.84 ;
      RECT 50.365 4.085 50.37 4.83 ;
      RECT 50.355 4.057 50.365 4.8 ;
      RECT 50.345 4.02 50.355 4.768 ;
      RECT 50.335 3.98 50.345 4.735 ;
      RECT 50.325 3.958 50.335 4.705 ;
      RECT 50.295 3.91 50.325 4.637 ;
      RECT 50.28 3.87 50.295 4.564 ;
      RECT 50.27 3.87 50.28 4.53 ;
      RECT 50.265 3.87 50.27 4.505 ;
      RECT 50.26 3.87 50.265 4.49 ;
      RECT 50.255 3.87 50.26 4.468 ;
      RECT 50.25 3.87 50.255 4.455 ;
      RECT 50.235 3.87 50.25 4.42 ;
      RECT 50.215 3.87 50.235 4.36 ;
      RECT 50.205 3.87 50.215 4.31 ;
      RECT 50.185 3.87 50.205 4.258 ;
      RECT 50.165 3.87 50.185 4.215 ;
      RECT 50.155 3.87 50.165 4.203 ;
      RECT 50.125 3.87 50.155 4.19 ;
      RECT 50.095 3.891 50.125 4.17 ;
      RECT 50.085 3.919 50.095 4.15 ;
      RECT 50.07 3.936 50.085 4.118 ;
      RECT 50.065 3.95 50.07 4.085 ;
      RECT 50.06 3.958 50.065 4.058 ;
      RECT 50.055 3.966 50.06 4.02 ;
      RECT 50.06 4.49 50.065 4.825 ;
      RECT 50.025 4.477 50.06 4.824 ;
      RECT 49.955 4.417 50.025 4.823 ;
      RECT 49.875 4.36 49.955 4.822 ;
      RECT 49.74 4.32 49.875 4.821 ;
      RECT 49.74 4.507 50.075 4.81 ;
      RECT 49.7 4.507 50.075 4.8 ;
      RECT 49.7 4.525 50.08 4.795 ;
      RECT 49.7 4.615 50.085 4.785 ;
      RECT 49.695 4.31 49.86 4.765 ;
      RECT 49.69 4.31 49.86 4.508 ;
      RECT 49.69 4.467 50.055 4.508 ;
      RECT 49.69 4.455 50.05 4.508 ;
      RECT 48.835 7.3 49.005 8.77 ;
      RECT 48.835 7.3 49.01 8.56 ;
      RECT 48.465 9.25 48.935 9.42 ;
      RECT 48.465 8.23 48.635 9.42 ;
      RECT 48.46 3.04 48.63 4.23 ;
      RECT 48.46 3.04 48.93 3.21 ;
      RECT 47.84 3.895 48.015 5.155 ;
      RECT 47.84 3.685 48.01 5.155 ;
      RECT 47.84 7.305 48.01 8.775 ;
      RECT 47.84 7.305 48.015 8.565 ;
      RECT 47.47 3.035 47.64 4.225 ;
      RECT 47.47 3.035 47.94 3.205 ;
      RECT 47.47 9.255 47.94 9.425 ;
      RECT 47.47 8.235 47.64 9.425 ;
      RECT 46.48 4.015 46.655 5.155 ;
      RECT 46.48 1.865 46.65 5.155 ;
      RECT 46.48 1.865 46.655 2.415 ;
      RECT 46.48 10.045 46.655 10.595 ;
      RECT 46.48 7.305 46.65 10.595 ;
      RECT 46.48 7.305 46.655 8.445 ;
      RECT 46.05 3.895 46.225 5.155 ;
      RECT 46.05 2.945 46.22 5.155 ;
      RECT 46.05 7.305 46.22 9.515 ;
      RECT 46.05 7.305 46.225 8.565 ;
      RECT 45.62 3.925 45.79 5.155 ;
      RECT 45.68 2.145 45.85 4.095 ;
      RECT 45.62 1.865 45.79 2.315 ;
      RECT 45.62 10.145 45.79 10.595 ;
      RECT 45.68 8.365 45.85 10.315 ;
      RECT 45.62 7.305 45.79 8.535 ;
      RECT 45.095 3.895 45.27 5.155 ;
      RECT 45.095 1.865 45.265 5.155 ;
      RECT 45.095 3.365 45.505 3.695 ;
      RECT 45.095 2.525 45.505 2.855 ;
      RECT 45.095 1.865 45.27 2.355 ;
      RECT 45.095 10.105 45.27 10.595 ;
      RECT 45.095 7.305 45.265 10.595 ;
      RECT 45.095 9.605 45.505 9.935 ;
      RECT 45.095 8.765 45.505 9.095 ;
      RECT 45.095 7.305 45.27 8.565 ;
      RECT 42.435 3.27 43.165 3.51 ;
      RECT 42.977 3.065 43.165 3.51 ;
      RECT 42.805 3.077 43.18 3.504 ;
      RECT 42.72 3.092 43.2 3.489 ;
      RECT 42.72 3.107 43.205 3.479 ;
      RECT 42.675 3.127 43.22 3.471 ;
      RECT 42.652 3.162 43.235 3.425 ;
      RECT 42.566 3.185 43.24 3.385 ;
      RECT 42.566 3.203 43.25 3.355 ;
      RECT 42.435 3.272 43.255 3.318 ;
      RECT 42.48 3.215 43.25 3.355 ;
      RECT 42.566 3.167 43.235 3.425 ;
      RECT 42.652 3.136 43.22 3.471 ;
      RECT 42.675 3.117 43.205 3.479 ;
      RECT 42.72 3.09 43.18 3.504 ;
      RECT 42.805 3.072 43.165 3.51 ;
      RECT 42.891 3.066 43.165 3.51 ;
      RECT 42.977 3.061 43.11 3.51 ;
      RECT 43.063 3.056 43.11 3.51 ;
      RECT 42.625 4.67 42.63 4.683 ;
      RECT 42.62 4.565 42.625 4.688 ;
      RECT 42.595 4.425 42.62 4.703 ;
      RECT 42.56 4.376 42.595 4.735 ;
      RECT 42.555 4.344 42.56 4.755 ;
      RECT 42.55 4.335 42.555 4.755 ;
      RECT 42.47 4.3 42.55 4.755 ;
      RECT 42.407 4.27 42.47 4.755 ;
      RECT 42.321 4.258 42.407 4.755 ;
      RECT 42.235 4.244 42.321 4.755 ;
      RECT 42.155 4.231 42.235 4.741 ;
      RECT 42.12 4.223 42.155 4.721 ;
      RECT 42.11 4.22 42.12 4.712 ;
      RECT 42.08 4.215 42.11 4.699 ;
      RECT 42.03 4.19 42.08 4.675 ;
      RECT 42.016 4.164 42.03 4.657 ;
      RECT 41.93 4.124 42.016 4.633 ;
      RECT 41.885 4.072 41.93 4.602 ;
      RECT 41.875 4.047 41.885 4.589 ;
      RECT 41.87 3.828 41.875 3.85 ;
      RECT 41.865 4.03 41.875 4.585 ;
      RECT 41.865 3.826 41.87 3.94 ;
      RECT 41.855 3.822 41.865 4.581 ;
      RECT 41.811 3.82 41.855 4.569 ;
      RECT 41.725 3.82 41.811 4.54 ;
      RECT 41.695 3.82 41.725 4.513 ;
      RECT 41.68 3.82 41.695 4.501 ;
      RECT 41.64 3.832 41.68 4.486 ;
      RECT 41.62 3.851 41.64 4.465 ;
      RECT 41.61 3.861 41.62 4.449 ;
      RECT 41.6 3.867 41.61 4.438 ;
      RECT 41.58 3.877 41.6 4.421 ;
      RECT 41.575 3.886 41.58 4.408 ;
      RECT 41.57 3.89 41.575 4.358 ;
      RECT 41.56 3.896 41.57 4.275 ;
      RECT 41.555 3.9 41.56 4.189 ;
      RECT 41.55 3.92 41.555 4.126 ;
      RECT 41.545 3.943 41.55 4.073 ;
      RECT 41.54 3.961 41.545 4.018 ;
      RECT 42.15 3.78 42.32 4.04 ;
      RECT 42.32 3.745 42.365 4.026 ;
      RECT 42.281 3.747 42.37 4.009 ;
      RECT 42.17 3.764 42.456 3.98 ;
      RECT 42.17 3.779 42.46 3.952 ;
      RECT 42.17 3.76 42.37 4.009 ;
      RECT 42.195 3.748 42.32 4.04 ;
      RECT 42.281 3.746 42.365 4.026 ;
      RECT 41.7 10.045 41.875 10.595 ;
      RECT 41.7 7.305 41.87 10.595 ;
      RECT 41.7 7.305 41.875 8.445 ;
      RECT 41.335 3.135 41.505 3.625 ;
      RECT 41.335 3.135 41.54 3.605 ;
      RECT 41.47 3.055 41.58 3.565 ;
      RECT 41.451 3.059 41.6 3.535 ;
      RECT 41.365 3.067 41.62 3.518 ;
      RECT 41.365 3.073 41.625 3.508 ;
      RECT 41.365 3.082 41.645 3.496 ;
      RECT 41.34 3.107 41.675 3.474 ;
      RECT 41.34 3.127 41.68 3.454 ;
      RECT 41.335 3.14 41.69 3.434 ;
      RECT 41.335 3.207 41.695 3.415 ;
      RECT 41.335 3.34 41.7 3.402 ;
      RECT 41.33 3.145 41.69 3.235 ;
      RECT 41.34 3.102 41.645 3.496 ;
      RECT 41.451 3.057 41.58 3.565 ;
      RECT 41.325 4.81 41.625 5.065 ;
      RECT 41.41 4.776 41.625 5.065 ;
      RECT 41.41 4.779 41.63 4.925 ;
      RECT 41.345 4.8 41.63 4.925 ;
      RECT 41.38 4.79 41.625 5.065 ;
      RECT 41.375 4.795 41.63 4.925 ;
      RECT 41.41 4.774 41.611 5.065 ;
      RECT 41.496 4.765 41.611 5.065 ;
      RECT 41.496 4.759 41.525 5.065 ;
      RECT 41.27 7.305 41.44 9.515 ;
      RECT 41.27 7.305 41.445 8.565 ;
      RECT 40.985 4.4 40.995 4.89 ;
      RECT 40.645 4.335 40.655 4.635 ;
      RECT 41.16 4.507 41.165 4.726 ;
      RECT 41.15 4.487 41.16 4.743 ;
      RECT 41.14 4.467 41.15 4.773 ;
      RECT 41.135 4.457 41.14 4.788 ;
      RECT 41.13 4.453 41.135 4.793 ;
      RECT 41.115 4.445 41.13 4.8 ;
      RECT 41.075 4.425 41.115 4.825 ;
      RECT 41.05 4.407 41.075 4.858 ;
      RECT 41.045 4.405 41.05 4.871 ;
      RECT 41.025 4.402 41.045 4.875 ;
      RECT 40.995 4.4 41.025 4.885 ;
      RECT 40.925 4.402 40.985 4.886 ;
      RECT 40.905 4.402 40.925 4.88 ;
      RECT 40.88 4.4 40.905 4.877 ;
      RECT 40.845 4.395 40.88 4.873 ;
      RECT 40.825 4.389 40.845 4.86 ;
      RECT 40.815 4.386 40.825 4.848 ;
      RECT 40.795 4.383 40.815 4.833 ;
      RECT 40.775 4.379 40.795 4.815 ;
      RECT 40.77 4.376 40.775 4.805 ;
      RECT 40.765 4.375 40.77 4.803 ;
      RECT 40.755 4.372 40.765 4.795 ;
      RECT 40.745 4.366 40.755 4.778 ;
      RECT 40.735 4.36 40.745 4.76 ;
      RECT 40.725 4.354 40.735 4.748 ;
      RECT 40.715 4.348 40.725 4.728 ;
      RECT 40.71 4.344 40.715 4.713 ;
      RECT 40.705 4.342 40.71 4.705 ;
      RECT 40.7 4.34 40.705 4.698 ;
      RECT 40.695 4.338 40.7 4.688 ;
      RECT 40.69 4.336 40.695 4.682 ;
      RECT 40.68 4.335 40.69 4.672 ;
      RECT 40.67 4.335 40.68 4.663 ;
      RECT 40.655 4.335 40.67 4.648 ;
      RECT 40.615 4.335 40.645 4.632 ;
      RECT 40.595 4.337 40.615 4.627 ;
      RECT 40.59 4.342 40.595 4.625 ;
      RECT 40.56 4.35 40.59 4.623 ;
      RECT 40.53 4.365 40.56 4.622 ;
      RECT 40.485 4.387 40.53 4.627 ;
      RECT 40.48 4.402 40.485 4.631 ;
      RECT 40.465 4.407 40.48 4.633 ;
      RECT 40.46 4.411 40.465 4.635 ;
      RECT 40.4 4.434 40.46 4.644 ;
      RECT 40.38 4.46 40.4 4.657 ;
      RECT 40.37 4.467 40.38 4.661 ;
      RECT 40.355 4.474 40.37 4.664 ;
      RECT 40.335 4.484 40.355 4.667 ;
      RECT 40.33 4.492 40.335 4.67 ;
      RECT 40.285 4.497 40.33 4.677 ;
      RECT 40.275 4.5 40.285 4.684 ;
      RECT 40.265 4.5 40.275 4.688 ;
      RECT 40.23 4.502 40.265 4.7 ;
      RECT 40.21 4.505 40.23 4.713 ;
      RECT 40.17 4.508 40.21 4.724 ;
      RECT 40.155 4.51 40.17 4.737 ;
      RECT 40.145 4.51 40.155 4.742 ;
      RECT 40.12 4.511 40.145 4.75 ;
      RECT 40.11 4.513 40.12 4.755 ;
      RECT 40.105 4.514 40.11 4.758 ;
      RECT 40.08 4.512 40.105 4.761 ;
      RECT 40.065 4.51 40.08 4.762 ;
      RECT 40.045 4.507 40.065 4.764 ;
      RECT 40.025 4.502 40.045 4.764 ;
      RECT 39.965 4.497 40.025 4.761 ;
      RECT 39.93 4.472 39.965 4.757 ;
      RECT 39.92 4.449 39.93 4.755 ;
      RECT 39.89 4.426 39.92 4.755 ;
      RECT 39.88 4.405 39.89 4.755 ;
      RECT 39.855 4.387 39.88 4.753 ;
      RECT 39.84 4.365 39.855 4.75 ;
      RECT 39.825 4.347 39.84 4.748 ;
      RECT 39.805 4.337 39.825 4.746 ;
      RECT 39.79 4.332 39.805 4.745 ;
      RECT 39.775 4.33 39.79 4.744 ;
      RECT 39.745 4.331 39.775 4.742 ;
      RECT 39.725 4.334 39.745 4.74 ;
      RECT 39.668 4.338 39.725 4.74 ;
      RECT 39.582 4.347 39.668 4.74 ;
      RECT 39.496 4.358 39.582 4.74 ;
      RECT 39.41 4.369 39.496 4.74 ;
      RECT 39.39 4.376 39.41 4.748 ;
      RECT 39.38 4.379 39.39 4.755 ;
      RECT 39.315 4.384 39.38 4.773 ;
      RECT 39.285 4.391 39.315 4.798 ;
      RECT 39.275 4.394 39.285 4.805 ;
      RECT 39.23 4.398 39.275 4.81 ;
      RECT 39.2 4.403 39.23 4.815 ;
      RECT 39.199 4.405 39.2 4.815 ;
      RECT 39.113 4.411 39.199 4.815 ;
      RECT 39.027 4.422 39.113 4.815 ;
      RECT 38.941 4.434 39.027 4.815 ;
      RECT 38.855 4.445 38.941 4.815 ;
      RECT 38.84 4.452 38.855 4.81 ;
      RECT 38.835 4.454 38.84 4.804 ;
      RECT 38.815 4.465 38.835 4.799 ;
      RECT 38.805 4.483 38.815 4.793 ;
      RECT 38.8 4.495 38.805 4.593 ;
      RECT 41.095 3.248 41.115 3.335 ;
      RECT 41.09 3.183 41.095 3.367 ;
      RECT 41.08 3.15 41.09 3.372 ;
      RECT 41.075 3.13 41.08 3.378 ;
      RECT 41.045 3.13 41.075 3.395 ;
      RECT 40.996 3.13 41.045 3.431 ;
      RECT 40.91 3.13 40.996 3.489 ;
      RECT 40.881 3.14 40.91 3.538 ;
      RECT 40.795 3.182 40.881 3.591 ;
      RECT 40.775 3.22 40.795 3.638 ;
      RECT 40.75 3.237 40.775 3.658 ;
      RECT 40.74 3.251 40.75 3.678 ;
      RECT 40.735 3.257 40.74 3.688 ;
      RECT 40.73 3.261 40.735 3.695 ;
      RECT 40.68 3.281 40.73 3.7 ;
      RECT 40.615 3.325 40.68 3.7 ;
      RECT 40.59 3.375 40.615 3.7 ;
      RECT 40.58 3.405 40.59 3.7 ;
      RECT 40.575 3.432 40.58 3.7 ;
      RECT 40.57 3.45 40.575 3.7 ;
      RECT 40.56 3.492 40.57 3.7 ;
      RECT 40.315 10.105 40.49 10.595 ;
      RECT 40.315 7.305 40.485 10.595 ;
      RECT 40.315 9.605 40.725 9.935 ;
      RECT 40.315 8.765 40.725 9.095 ;
      RECT 40.315 7.305 40.49 8.565 ;
      RECT 40.39 4.85 40.58 5.075 ;
      RECT 40.38 4.851 40.585 5.07 ;
      RECT 40.38 4.853 40.595 5.05 ;
      RECT 40.38 4.857 40.6 5.035 ;
      RECT 40.38 4.844 40.55 5.07 ;
      RECT 40.38 4.847 40.575 5.07 ;
      RECT 40.39 4.843 40.55 5.075 ;
      RECT 40.476 4.841 40.55 5.075 ;
      RECT 40.1 4.092 40.27 4.33 ;
      RECT 40.1 4.092 40.356 4.244 ;
      RECT 40.1 4.092 40.36 4.154 ;
      RECT 40.15 3.865 40.37 4.133 ;
      RECT 40.145 3.882 40.375 4.106 ;
      RECT 40.11 4.04 40.375 4.106 ;
      RECT 40.13 3.89 40.27 4.33 ;
      RECT 40.12 3.972 40.38 4.089 ;
      RECT 40.115 4.02 40.38 4.089 ;
      RECT 40.12 3.93 40.375 4.106 ;
      RECT 40.145 3.867 40.37 4.133 ;
      RECT 39.71 3.842 39.88 4.04 ;
      RECT 39.71 3.842 39.925 4.015 ;
      RECT 39.78 3.785 39.95 3.973 ;
      RECT 39.755 3.8 39.95 3.973 ;
      RECT 39.37 3.846 39.4 4.04 ;
      RECT 39.365 3.818 39.37 4.04 ;
      RECT 39.335 3.792 39.365 4.042 ;
      RECT 39.31 3.75 39.335 4.045 ;
      RECT 39.3 3.722 39.31 4.047 ;
      RECT 39.265 3.702 39.3 4.049 ;
      RECT 39.2 3.687 39.265 4.055 ;
      RECT 39.15 3.685 39.2 4.061 ;
      RECT 39.127 3.687 39.15 4.066 ;
      RECT 39.041 3.698 39.127 4.072 ;
      RECT 38.955 3.716 39.041 4.082 ;
      RECT 38.94 3.727 38.955 4.088 ;
      RECT 38.87 3.75 38.94 4.094 ;
      RECT 38.815 3.782 38.87 4.102 ;
      RECT 38.775 3.805 38.815 4.108 ;
      RECT 38.761 3.818 38.775 4.111 ;
      RECT 38.675 3.84 38.761 4.117 ;
      RECT 38.66 3.865 38.675 4.123 ;
      RECT 38.62 3.88 38.66 4.127 ;
      RECT 38.57 3.895 38.62 4.132 ;
      RECT 38.545 3.902 38.57 4.136 ;
      RECT 38.485 3.897 38.545 4.14 ;
      RECT 38.47 3.888 38.485 4.144 ;
      RECT 38.4 3.878 38.47 4.14 ;
      RECT 38.375 3.87 38.395 4.13 ;
      RECT 38.316 3.87 38.375 4.108 ;
      RECT 38.23 3.87 38.316 4.065 ;
      RECT 38.395 3.87 38.4 4.135 ;
      RECT 39.09 3.101 39.26 3.435 ;
      RECT 39.06 3.101 39.26 3.43 ;
      RECT 39 3.068 39.06 3.418 ;
      RECT 39 3.124 39.27 3.413 ;
      RECT 38.975 3.124 39.27 3.407 ;
      RECT 38.97 3.065 39 3.404 ;
      RECT 38.955 3.071 39.09 3.402 ;
      RECT 38.95 3.079 39.175 3.39 ;
      RECT 38.95 3.131 39.285 3.343 ;
      RECT 38.935 3.087 39.175 3.338 ;
      RECT 38.935 3.157 39.295 3.279 ;
      RECT 38.905 3.107 39.26 3.24 ;
      RECT 38.905 3.197 39.305 3.236 ;
      RECT 38.955 3.076 39.175 3.402 ;
      RECT 38.295 3.406 38.35 3.67 ;
      RECT 38.295 3.406 38.415 3.669 ;
      RECT 38.295 3.406 38.44 3.668 ;
      RECT 38.295 3.406 38.505 3.667 ;
      RECT 38.44 3.372 38.52 3.666 ;
      RECT 38.255 3.416 38.665 3.665 ;
      RECT 38.295 3.413 38.665 3.665 ;
      RECT 38.255 3.421 38.67 3.658 ;
      RECT 38.24 3.423 38.67 3.657 ;
      RECT 38.24 3.43 38.675 3.653 ;
      RECT 38.22 3.429 38.67 3.649 ;
      RECT 38.22 3.437 38.68 3.648 ;
      RECT 38.215 3.434 38.675 3.644 ;
      RECT 38.215 3.447 38.69 3.643 ;
      RECT 38.2 3.437 38.68 3.642 ;
      RECT 38.165 3.45 38.69 3.635 ;
      RECT 38.35 3.405 38.66 3.665 ;
      RECT 38.35 3.39 38.61 3.665 ;
      RECT 38.415 3.377 38.545 3.665 ;
      RECT 37.96 4.466 37.975 4.859 ;
      RECT 37.925 4.471 37.975 4.858 ;
      RECT 37.96 4.47 38.02 4.857 ;
      RECT 37.905 4.481 38.02 4.856 ;
      RECT 37.92 4.477 38.02 4.856 ;
      RECT 37.885 4.487 38.095 4.853 ;
      RECT 37.885 4.506 38.14 4.851 ;
      RECT 37.885 4.513 38.145 4.848 ;
      RECT 37.87 4.49 38.095 4.845 ;
      RECT 37.85 4.495 38.095 4.838 ;
      RECT 37.845 4.499 38.095 4.834 ;
      RECT 37.845 4.516 38.155 4.833 ;
      RECT 37.825 4.51 38.14 4.829 ;
      RECT 37.825 4.519 38.16 4.823 ;
      RECT 37.82 4.525 38.16 4.595 ;
      RECT 37.885 4.485 38.02 4.853 ;
      RECT 37.76 3.848 37.96 4.16 ;
      RECT 37.835 3.826 37.96 4.16 ;
      RECT 37.775 3.845 37.965 4.145 ;
      RECT 37.745 3.856 37.965 4.143 ;
      RECT 37.76 3.851 37.97 4.109 ;
      RECT 37.745 3.955 37.975 4.076 ;
      RECT 37.775 3.827 37.96 4.16 ;
      RECT 37.835 3.805 37.935 4.16 ;
      RECT 37.86 3.802 37.935 4.16 ;
      RECT 37.86 3.797 37.88 4.16 ;
      RECT 37.265 3.865 37.44 4.04 ;
      RECT 37.26 3.865 37.44 4.038 ;
      RECT 37.235 3.865 37.44 4.033 ;
      RECT 37.18 3.845 37.35 4.023 ;
      RECT 37.18 3.852 37.415 4.023 ;
      RECT 37.265 4.532 37.28 4.715 ;
      RECT 37.255 4.51 37.265 4.715 ;
      RECT 37.24 4.49 37.255 4.715 ;
      RECT 37.23 4.465 37.24 4.715 ;
      RECT 37.2 4.43 37.23 4.715 ;
      RECT 37.165 4.37 37.2 4.715 ;
      RECT 37.16 4.332 37.165 4.715 ;
      RECT 37.11 4.283 37.16 4.715 ;
      RECT 37.1 4.233 37.11 4.703 ;
      RECT 37.085 4.212 37.1 4.663 ;
      RECT 37.065 4.18 37.085 4.613 ;
      RECT 37.04 4.136 37.065 4.553 ;
      RECT 37.035 4.108 37.04 4.508 ;
      RECT 37.03 4.099 37.035 4.494 ;
      RECT 37.025 4.092 37.03 4.481 ;
      RECT 37.02 4.087 37.025 4.47 ;
      RECT 37.015 4.072 37.02 4.46 ;
      RECT 37.01 4.05 37.015 4.447 ;
      RECT 37 4.01 37.01 4.422 ;
      RECT 36.975 3.94 37 4.378 ;
      RECT 36.97 3.88 36.975 4.343 ;
      RECT 36.955 3.86 36.97 4.31 ;
      RECT 36.95 3.86 36.955 4.285 ;
      RECT 36.92 3.86 36.95 4.24 ;
      RECT 36.875 3.86 36.92 4.18 ;
      RECT 36.8 3.86 36.875 4.128 ;
      RECT 36.795 3.86 36.8 4.093 ;
      RECT 36.79 3.86 36.795 4.083 ;
      RECT 36.785 3.86 36.79 4.063 ;
      RECT 37.05 3.08 37.22 3.55 ;
      RECT 36.995 3.073 37.19 3.534 ;
      RECT 36.995 3.087 37.225 3.533 ;
      RECT 36.98 3.088 37.225 3.514 ;
      RECT 36.975 3.106 37.225 3.5 ;
      RECT 36.98 3.089 37.23 3.498 ;
      RECT 36.965 3.12 37.23 3.483 ;
      RECT 36.98 3.095 37.235 3.468 ;
      RECT 36.96 3.135 37.235 3.465 ;
      RECT 36.975 3.107 37.24 3.45 ;
      RECT 36.975 3.119 37.245 3.43 ;
      RECT 36.96 3.135 37.25 3.413 ;
      RECT 36.96 3.145 37.255 3.268 ;
      RECT 36.955 3.145 37.255 3.225 ;
      RECT 36.955 3.16 37.26 3.203 ;
      RECT 37.05 3.07 37.19 3.55 ;
      RECT 37.05 3.068 37.16 3.55 ;
      RECT 37.136 3.065 37.16 3.55 ;
      RECT 36.795 4.732 36.8 4.778 ;
      RECT 36.785 4.58 36.795 4.802 ;
      RECT 36.78 4.425 36.785 4.827 ;
      RECT 36.765 4.387 36.78 4.838 ;
      RECT 36.76 4.37 36.765 4.845 ;
      RECT 36.75 4.358 36.76 4.852 ;
      RECT 36.745 4.349 36.75 4.854 ;
      RECT 36.74 4.347 36.745 4.858 ;
      RECT 36.695 4.338 36.74 4.873 ;
      RECT 36.69 4.33 36.695 4.887 ;
      RECT 36.685 4.327 36.69 4.891 ;
      RECT 36.67 4.322 36.685 4.899 ;
      RECT 36.615 4.312 36.67 4.91 ;
      RECT 36.58 4.3 36.615 4.911 ;
      RECT 36.571 4.295 36.58 4.905 ;
      RECT 36.485 4.295 36.571 4.895 ;
      RECT 36.455 4.295 36.485 4.873 ;
      RECT 36.445 4.295 36.45 4.853 ;
      RECT 36.44 4.295 36.445 4.815 ;
      RECT 36.435 4.295 36.44 4.773 ;
      RECT 36.43 4.295 36.435 4.733 ;
      RECT 36.425 4.295 36.43 4.663 ;
      RECT 36.415 4.295 36.425 4.585 ;
      RECT 36.41 4.295 36.415 4.485 ;
      RECT 36.45 4.295 36.455 4.855 ;
      RECT 35.945 4.377 36.035 4.855 ;
      RECT 35.93 4.38 36.05 4.853 ;
      RECT 35.945 4.379 36.05 4.853 ;
      RECT 35.91 4.386 36.075 4.843 ;
      RECT 35.93 4.38 36.075 4.843 ;
      RECT 35.895 4.392 36.075 4.831 ;
      RECT 35.93 4.383 36.125 4.824 ;
      RECT 35.881 4.4 36.125 4.822 ;
      RECT 35.91 4.39 36.135 4.81 ;
      RECT 35.881 4.411 36.165 4.801 ;
      RECT 35.795 4.435 36.165 4.795 ;
      RECT 35.795 4.448 36.205 4.778 ;
      RECT 35.79 4.47 36.205 4.771 ;
      RECT 35.76 4.485 36.205 4.761 ;
      RECT 35.755 4.496 36.205 4.751 ;
      RECT 35.725 4.509 36.205 4.742 ;
      RECT 35.71 4.527 36.205 4.731 ;
      RECT 35.685 4.54 36.205 4.721 ;
      RECT 35.945 4.376 35.955 4.855 ;
      RECT 35.991 3.8 36.03 4.045 ;
      RECT 35.905 3.8 36.04 4.043 ;
      RECT 35.79 3.825 36.04 4.04 ;
      RECT 35.79 3.825 36.045 4.038 ;
      RECT 35.79 3.825 36.06 4.033 ;
      RECT 35.896 3.8 36.075 4.013 ;
      RECT 35.81 3.808 36.075 4.013 ;
      RECT 35.48 3.16 35.65 3.595 ;
      RECT 35.47 3.194 35.65 3.578 ;
      RECT 35.55 3.13 35.72 3.565 ;
      RECT 35.455 3.205 35.72 3.543 ;
      RECT 35.55 3.14 35.725 3.533 ;
      RECT 35.48 3.192 35.755 3.518 ;
      RECT 35.44 3.218 35.755 3.503 ;
      RECT 35.44 3.26 35.765 3.483 ;
      RECT 35.435 3.285 35.77 3.465 ;
      RECT 35.435 3.295 35.775 3.45 ;
      RECT 35.43 3.232 35.755 3.448 ;
      RECT 35.43 3.305 35.78 3.433 ;
      RECT 35.425 3.242 35.755 3.43 ;
      RECT 35.42 3.326 35.785 3.413 ;
      RECT 35.42 3.358 35.79 3.393 ;
      RECT 35.415 3.272 35.765 3.385 ;
      RECT 35.42 3.257 35.755 3.413 ;
      RECT 35.435 3.227 35.755 3.465 ;
      RECT 35.28 3.814 35.505 4.07 ;
      RECT 35.28 3.847 35.525 4.06 ;
      RECT 35.245 3.847 35.525 4.058 ;
      RECT 35.245 3.86 35.53 4.048 ;
      RECT 35.245 3.88 35.54 4.04 ;
      RECT 35.245 3.977 35.545 4.033 ;
      RECT 35.225 3.725 35.355 4.023 ;
      RECT 35.18 3.88 35.54 3.965 ;
      RECT 35.17 3.725 35.355 3.91 ;
      RECT 35.17 3.757 35.441 3.91 ;
      RECT 35.135 4.287 35.155 4.465 ;
      RECT 35.1 4.24 35.135 4.465 ;
      RECT 35.085 4.18 35.1 4.465 ;
      RECT 35.06 4.127 35.085 4.465 ;
      RECT 35.045 4.08 35.06 4.465 ;
      RECT 35.025 4.057 35.045 4.465 ;
      RECT 35 4.022 35.025 4.465 ;
      RECT 34.99 3.868 35 4.465 ;
      RECT 34.96 3.863 34.99 4.456 ;
      RECT 34.955 3.86 34.96 4.446 ;
      RECT 34.94 3.86 34.955 4.42 ;
      RECT 34.935 3.86 34.94 4.383 ;
      RECT 34.91 3.86 34.935 4.335 ;
      RECT 34.89 3.86 34.91 4.26 ;
      RECT 34.88 3.86 34.89 4.22 ;
      RECT 34.875 3.86 34.88 4.195 ;
      RECT 34.87 3.86 34.875 4.178 ;
      RECT 34.865 3.86 34.87 4.16 ;
      RECT 34.86 3.861 34.865 4.15 ;
      RECT 34.85 3.863 34.86 4.118 ;
      RECT 34.84 3.865 34.85 4.085 ;
      RECT 34.83 3.868 34.84 4.058 ;
      RECT 35.155 4.295 35.38 4.465 ;
      RECT 34.485 3.107 34.655 3.56 ;
      RECT 34.485 3.107 34.745 3.526 ;
      RECT 34.485 3.107 34.775 3.51 ;
      RECT 34.485 3.107 34.805 3.483 ;
      RECT 34.741 3.085 34.82 3.465 ;
      RECT 34.52 3.092 34.825 3.45 ;
      RECT 34.52 3.1 34.835 3.413 ;
      RECT 34.48 3.127 34.835 3.385 ;
      RECT 34.465 3.14 34.835 3.35 ;
      RECT 34.485 3.115 34.855 3.34 ;
      RECT 34.46 3.18 34.855 3.31 ;
      RECT 34.46 3.21 34.86 3.293 ;
      RECT 34.455 3.24 34.86 3.28 ;
      RECT 34.52 3.089 34.82 3.465 ;
      RECT 34.655 3.086 34.741 3.544 ;
      RECT 34.606 3.087 34.82 3.465 ;
      RECT 34.75 4.747 34.795 4.94 ;
      RECT 34.74 4.717 34.75 4.94 ;
      RECT 34.735 4.702 34.74 4.94 ;
      RECT 34.695 4.612 34.735 4.94 ;
      RECT 34.69 4.525 34.695 4.94 ;
      RECT 34.68 4.495 34.69 4.94 ;
      RECT 34.675 4.455 34.68 4.94 ;
      RECT 34.665 4.417 34.675 4.94 ;
      RECT 34.66 4.382 34.665 4.94 ;
      RECT 34.64 4.335 34.66 4.94 ;
      RECT 34.625 4.26 34.64 4.94 ;
      RECT 34.62 4.215 34.625 4.935 ;
      RECT 34.615 4.195 34.62 4.908 ;
      RECT 34.61 4.175 34.615 4.893 ;
      RECT 34.605 4.15 34.61 4.873 ;
      RECT 34.6 4.128 34.605 4.858 ;
      RECT 34.595 4.106 34.6 4.84 ;
      RECT 34.59 4.085 34.595 4.83 ;
      RECT 34.58 4.057 34.59 4.8 ;
      RECT 34.57 4.02 34.58 4.768 ;
      RECT 34.56 3.98 34.57 4.735 ;
      RECT 34.55 3.958 34.56 4.705 ;
      RECT 34.52 3.91 34.55 4.637 ;
      RECT 34.505 3.87 34.52 4.564 ;
      RECT 34.495 3.87 34.505 4.53 ;
      RECT 34.49 3.87 34.495 4.505 ;
      RECT 34.485 3.87 34.49 4.49 ;
      RECT 34.48 3.87 34.485 4.468 ;
      RECT 34.475 3.87 34.48 4.455 ;
      RECT 34.46 3.87 34.475 4.42 ;
      RECT 34.44 3.87 34.46 4.36 ;
      RECT 34.43 3.87 34.44 4.31 ;
      RECT 34.41 3.87 34.43 4.258 ;
      RECT 34.39 3.87 34.41 4.215 ;
      RECT 34.38 3.87 34.39 4.203 ;
      RECT 34.35 3.87 34.38 4.19 ;
      RECT 34.32 3.891 34.35 4.17 ;
      RECT 34.31 3.919 34.32 4.15 ;
      RECT 34.295 3.936 34.31 4.118 ;
      RECT 34.29 3.95 34.295 4.085 ;
      RECT 34.285 3.958 34.29 4.058 ;
      RECT 34.28 3.966 34.285 4.02 ;
      RECT 34.285 4.49 34.29 4.825 ;
      RECT 34.25 4.477 34.285 4.824 ;
      RECT 34.18 4.417 34.25 4.823 ;
      RECT 34.1 4.36 34.18 4.822 ;
      RECT 33.965 4.32 34.1 4.821 ;
      RECT 33.965 4.507 34.3 4.81 ;
      RECT 33.925 4.507 34.3 4.8 ;
      RECT 33.925 4.525 34.305 4.795 ;
      RECT 33.925 4.615 34.31 4.785 ;
      RECT 33.92 4.31 34.085 4.765 ;
      RECT 33.915 4.31 34.085 4.508 ;
      RECT 33.915 4.467 34.28 4.508 ;
      RECT 33.915 4.455 34.275 4.508 ;
      RECT 33.055 7.3 33.225 8.77 ;
      RECT 33.055 7.3 33.23 8.56 ;
      RECT 32.685 9.25 33.155 9.42 ;
      RECT 32.685 8.23 32.855 9.42 ;
      RECT 32.68 3.04 32.85 4.23 ;
      RECT 32.68 3.04 33.15 3.21 ;
      RECT 32.06 3.895 32.235 5.155 ;
      RECT 32.06 3.685 32.23 5.155 ;
      RECT 32.06 7.305 32.23 8.775 ;
      RECT 32.06 7.305 32.235 8.565 ;
      RECT 31.69 3.035 31.86 4.225 ;
      RECT 31.69 3.035 32.16 3.205 ;
      RECT 31.69 9.255 32.16 9.425 ;
      RECT 31.69 8.235 31.86 9.425 ;
      RECT 30.7 4.015 30.875 5.155 ;
      RECT 30.7 1.865 30.87 5.155 ;
      RECT 30.7 1.865 30.875 2.415 ;
      RECT 30.7 10.045 30.875 10.595 ;
      RECT 30.7 7.305 30.87 10.595 ;
      RECT 30.7 7.305 30.875 8.445 ;
      RECT 30.27 3.895 30.445 5.155 ;
      RECT 30.27 2.945 30.44 5.155 ;
      RECT 30.27 7.305 30.44 9.515 ;
      RECT 30.27 7.305 30.445 8.565 ;
      RECT 29.84 3.925 30.01 5.155 ;
      RECT 29.9 2.145 30.07 4.095 ;
      RECT 29.84 1.865 30.01 2.315 ;
      RECT 29.84 10.145 30.01 10.595 ;
      RECT 29.9 8.365 30.07 10.315 ;
      RECT 29.84 7.305 30.01 8.535 ;
      RECT 29.315 3.895 29.49 5.155 ;
      RECT 29.315 1.865 29.485 5.155 ;
      RECT 29.315 3.365 29.725 3.695 ;
      RECT 29.315 2.525 29.725 2.855 ;
      RECT 29.315 1.865 29.49 2.355 ;
      RECT 29.315 10.105 29.49 10.595 ;
      RECT 29.315 7.305 29.485 10.595 ;
      RECT 29.315 9.605 29.725 9.935 ;
      RECT 29.315 8.765 29.725 9.095 ;
      RECT 29.315 7.305 29.49 8.565 ;
      RECT 26.655 3.27 27.385 3.51 ;
      RECT 27.197 3.065 27.385 3.51 ;
      RECT 27.025 3.077 27.4 3.504 ;
      RECT 26.94 3.092 27.42 3.489 ;
      RECT 26.94 3.107 27.425 3.479 ;
      RECT 26.895 3.127 27.44 3.471 ;
      RECT 26.872 3.162 27.455 3.425 ;
      RECT 26.786 3.185 27.46 3.385 ;
      RECT 26.786 3.203 27.47 3.355 ;
      RECT 26.655 3.272 27.475 3.318 ;
      RECT 26.7 3.215 27.47 3.355 ;
      RECT 26.786 3.167 27.455 3.425 ;
      RECT 26.872 3.136 27.44 3.471 ;
      RECT 26.895 3.117 27.425 3.479 ;
      RECT 26.94 3.09 27.4 3.504 ;
      RECT 27.025 3.072 27.385 3.51 ;
      RECT 27.111 3.066 27.385 3.51 ;
      RECT 27.197 3.061 27.33 3.51 ;
      RECT 27.283 3.056 27.33 3.51 ;
      RECT 26.845 4.67 26.85 4.683 ;
      RECT 26.84 4.565 26.845 4.688 ;
      RECT 26.815 4.425 26.84 4.703 ;
      RECT 26.78 4.376 26.815 4.735 ;
      RECT 26.775 4.344 26.78 4.755 ;
      RECT 26.77 4.335 26.775 4.755 ;
      RECT 26.69 4.3 26.77 4.755 ;
      RECT 26.627 4.27 26.69 4.755 ;
      RECT 26.541 4.258 26.627 4.755 ;
      RECT 26.455 4.244 26.541 4.755 ;
      RECT 26.375 4.231 26.455 4.741 ;
      RECT 26.34 4.223 26.375 4.721 ;
      RECT 26.33 4.22 26.34 4.712 ;
      RECT 26.3 4.215 26.33 4.699 ;
      RECT 26.25 4.19 26.3 4.675 ;
      RECT 26.236 4.164 26.25 4.657 ;
      RECT 26.15 4.124 26.236 4.633 ;
      RECT 26.105 4.072 26.15 4.602 ;
      RECT 26.095 4.047 26.105 4.589 ;
      RECT 26.09 3.828 26.095 3.85 ;
      RECT 26.085 4.03 26.095 4.585 ;
      RECT 26.085 3.826 26.09 3.94 ;
      RECT 26.075 3.822 26.085 4.581 ;
      RECT 26.031 3.82 26.075 4.569 ;
      RECT 25.945 3.82 26.031 4.54 ;
      RECT 25.915 3.82 25.945 4.513 ;
      RECT 25.9 3.82 25.915 4.501 ;
      RECT 25.86 3.832 25.9 4.486 ;
      RECT 25.84 3.851 25.86 4.465 ;
      RECT 25.83 3.861 25.84 4.449 ;
      RECT 25.82 3.867 25.83 4.438 ;
      RECT 25.8 3.877 25.82 4.421 ;
      RECT 25.795 3.886 25.8 4.408 ;
      RECT 25.79 3.89 25.795 4.358 ;
      RECT 25.78 3.896 25.79 4.275 ;
      RECT 25.775 3.9 25.78 4.189 ;
      RECT 25.77 3.92 25.775 4.126 ;
      RECT 25.765 3.943 25.77 4.073 ;
      RECT 25.76 3.961 25.765 4.018 ;
      RECT 26.37 3.78 26.54 4.04 ;
      RECT 26.54 3.745 26.585 4.026 ;
      RECT 26.501 3.747 26.59 4.009 ;
      RECT 26.39 3.764 26.676 3.98 ;
      RECT 26.39 3.779 26.68 3.952 ;
      RECT 26.39 3.76 26.59 4.009 ;
      RECT 26.415 3.748 26.54 4.04 ;
      RECT 26.501 3.746 26.585 4.026 ;
      RECT 25.92 10.045 26.095 10.595 ;
      RECT 25.92 7.305 26.09 10.595 ;
      RECT 25.92 7.305 26.095 8.445 ;
      RECT 25.555 3.135 25.725 3.625 ;
      RECT 25.555 3.135 25.76 3.605 ;
      RECT 25.69 3.055 25.8 3.565 ;
      RECT 25.671 3.059 25.82 3.535 ;
      RECT 25.585 3.067 25.84 3.518 ;
      RECT 25.585 3.073 25.845 3.508 ;
      RECT 25.585 3.082 25.865 3.496 ;
      RECT 25.56 3.107 25.895 3.474 ;
      RECT 25.56 3.127 25.9 3.454 ;
      RECT 25.555 3.14 25.91 3.434 ;
      RECT 25.555 3.207 25.915 3.415 ;
      RECT 25.555 3.34 25.92 3.402 ;
      RECT 25.55 3.145 25.91 3.235 ;
      RECT 25.56 3.102 25.865 3.496 ;
      RECT 25.671 3.057 25.8 3.565 ;
      RECT 25.545 4.81 25.845 5.065 ;
      RECT 25.63 4.776 25.845 5.065 ;
      RECT 25.63 4.779 25.85 4.925 ;
      RECT 25.565 4.8 25.85 4.925 ;
      RECT 25.6 4.79 25.845 5.065 ;
      RECT 25.595 4.795 25.85 4.925 ;
      RECT 25.63 4.774 25.831 5.065 ;
      RECT 25.716 4.765 25.831 5.065 ;
      RECT 25.716 4.759 25.745 5.065 ;
      RECT 25.49 7.305 25.66 9.515 ;
      RECT 25.49 7.305 25.665 8.565 ;
      RECT 25.205 4.4 25.215 4.89 ;
      RECT 24.865 4.335 24.875 4.635 ;
      RECT 25.38 4.507 25.385 4.726 ;
      RECT 25.37 4.487 25.38 4.743 ;
      RECT 25.36 4.467 25.37 4.773 ;
      RECT 25.355 4.457 25.36 4.788 ;
      RECT 25.35 4.453 25.355 4.793 ;
      RECT 25.335 4.445 25.35 4.8 ;
      RECT 25.295 4.425 25.335 4.825 ;
      RECT 25.27 4.407 25.295 4.858 ;
      RECT 25.265 4.405 25.27 4.871 ;
      RECT 25.245 4.402 25.265 4.875 ;
      RECT 25.215 4.4 25.245 4.885 ;
      RECT 25.145 4.402 25.205 4.886 ;
      RECT 25.125 4.402 25.145 4.88 ;
      RECT 25.1 4.4 25.125 4.877 ;
      RECT 25.065 4.395 25.1 4.873 ;
      RECT 25.045 4.389 25.065 4.86 ;
      RECT 25.035 4.386 25.045 4.848 ;
      RECT 25.015 4.383 25.035 4.833 ;
      RECT 24.995 4.379 25.015 4.815 ;
      RECT 24.99 4.376 24.995 4.805 ;
      RECT 24.985 4.375 24.99 4.803 ;
      RECT 24.975 4.372 24.985 4.795 ;
      RECT 24.965 4.366 24.975 4.778 ;
      RECT 24.955 4.36 24.965 4.76 ;
      RECT 24.945 4.354 24.955 4.748 ;
      RECT 24.935 4.348 24.945 4.728 ;
      RECT 24.93 4.344 24.935 4.713 ;
      RECT 24.925 4.342 24.93 4.705 ;
      RECT 24.92 4.34 24.925 4.698 ;
      RECT 24.915 4.338 24.92 4.688 ;
      RECT 24.91 4.336 24.915 4.682 ;
      RECT 24.9 4.335 24.91 4.672 ;
      RECT 24.89 4.335 24.9 4.663 ;
      RECT 24.875 4.335 24.89 4.648 ;
      RECT 24.835 4.335 24.865 4.632 ;
      RECT 24.815 4.337 24.835 4.627 ;
      RECT 24.81 4.342 24.815 4.625 ;
      RECT 24.78 4.35 24.81 4.623 ;
      RECT 24.75 4.365 24.78 4.622 ;
      RECT 24.705 4.387 24.75 4.627 ;
      RECT 24.7 4.402 24.705 4.631 ;
      RECT 24.685 4.407 24.7 4.633 ;
      RECT 24.68 4.411 24.685 4.635 ;
      RECT 24.62 4.434 24.68 4.644 ;
      RECT 24.6 4.46 24.62 4.657 ;
      RECT 24.59 4.467 24.6 4.661 ;
      RECT 24.575 4.474 24.59 4.664 ;
      RECT 24.555 4.484 24.575 4.667 ;
      RECT 24.55 4.492 24.555 4.67 ;
      RECT 24.505 4.497 24.55 4.677 ;
      RECT 24.495 4.5 24.505 4.684 ;
      RECT 24.485 4.5 24.495 4.688 ;
      RECT 24.45 4.502 24.485 4.7 ;
      RECT 24.43 4.505 24.45 4.713 ;
      RECT 24.39 4.508 24.43 4.724 ;
      RECT 24.375 4.51 24.39 4.737 ;
      RECT 24.365 4.51 24.375 4.742 ;
      RECT 24.34 4.511 24.365 4.75 ;
      RECT 24.33 4.513 24.34 4.755 ;
      RECT 24.325 4.514 24.33 4.758 ;
      RECT 24.3 4.512 24.325 4.761 ;
      RECT 24.285 4.51 24.3 4.762 ;
      RECT 24.265 4.507 24.285 4.764 ;
      RECT 24.245 4.502 24.265 4.764 ;
      RECT 24.185 4.497 24.245 4.761 ;
      RECT 24.15 4.472 24.185 4.757 ;
      RECT 24.14 4.449 24.15 4.755 ;
      RECT 24.11 4.426 24.14 4.755 ;
      RECT 24.1 4.405 24.11 4.755 ;
      RECT 24.075 4.387 24.1 4.753 ;
      RECT 24.06 4.365 24.075 4.75 ;
      RECT 24.045 4.347 24.06 4.748 ;
      RECT 24.025 4.337 24.045 4.746 ;
      RECT 24.01 4.332 24.025 4.745 ;
      RECT 23.995 4.33 24.01 4.744 ;
      RECT 23.965 4.331 23.995 4.742 ;
      RECT 23.945 4.334 23.965 4.74 ;
      RECT 23.888 4.338 23.945 4.74 ;
      RECT 23.802 4.347 23.888 4.74 ;
      RECT 23.716 4.358 23.802 4.74 ;
      RECT 23.63 4.369 23.716 4.74 ;
      RECT 23.61 4.376 23.63 4.748 ;
      RECT 23.6 4.379 23.61 4.755 ;
      RECT 23.535 4.384 23.6 4.773 ;
      RECT 23.505 4.391 23.535 4.798 ;
      RECT 23.495 4.394 23.505 4.805 ;
      RECT 23.45 4.398 23.495 4.81 ;
      RECT 23.42 4.403 23.45 4.815 ;
      RECT 23.419 4.405 23.42 4.815 ;
      RECT 23.333 4.411 23.419 4.815 ;
      RECT 23.247 4.422 23.333 4.815 ;
      RECT 23.161 4.434 23.247 4.815 ;
      RECT 23.075 4.445 23.161 4.815 ;
      RECT 23.06 4.452 23.075 4.81 ;
      RECT 23.055 4.454 23.06 4.804 ;
      RECT 23.035 4.465 23.055 4.799 ;
      RECT 23.025 4.483 23.035 4.793 ;
      RECT 23.02 4.495 23.025 4.593 ;
      RECT 25.315 3.248 25.335 3.335 ;
      RECT 25.31 3.183 25.315 3.367 ;
      RECT 25.3 3.15 25.31 3.372 ;
      RECT 25.295 3.13 25.3 3.378 ;
      RECT 25.265 3.13 25.295 3.395 ;
      RECT 25.216 3.13 25.265 3.431 ;
      RECT 25.13 3.13 25.216 3.489 ;
      RECT 25.101 3.14 25.13 3.538 ;
      RECT 25.015 3.182 25.101 3.591 ;
      RECT 24.995 3.22 25.015 3.638 ;
      RECT 24.97 3.237 24.995 3.658 ;
      RECT 24.96 3.251 24.97 3.678 ;
      RECT 24.955 3.257 24.96 3.688 ;
      RECT 24.95 3.261 24.955 3.695 ;
      RECT 24.9 3.281 24.95 3.7 ;
      RECT 24.835 3.325 24.9 3.7 ;
      RECT 24.81 3.375 24.835 3.7 ;
      RECT 24.8 3.405 24.81 3.7 ;
      RECT 24.795 3.432 24.8 3.7 ;
      RECT 24.79 3.45 24.795 3.7 ;
      RECT 24.78 3.492 24.79 3.7 ;
      RECT 24.535 10.105 24.71 10.595 ;
      RECT 24.535 7.305 24.705 10.595 ;
      RECT 24.535 9.605 24.945 9.935 ;
      RECT 24.535 8.765 24.945 9.095 ;
      RECT 24.535 7.305 24.71 8.565 ;
      RECT 24.61 4.85 24.8 5.075 ;
      RECT 24.6 4.851 24.805 5.07 ;
      RECT 24.6 4.853 24.815 5.05 ;
      RECT 24.6 4.857 24.82 5.035 ;
      RECT 24.6 4.844 24.77 5.07 ;
      RECT 24.6 4.847 24.795 5.07 ;
      RECT 24.61 4.843 24.77 5.075 ;
      RECT 24.696 4.841 24.77 5.075 ;
      RECT 24.32 4.092 24.49 4.33 ;
      RECT 24.32 4.092 24.576 4.244 ;
      RECT 24.32 4.092 24.58 4.154 ;
      RECT 24.37 3.865 24.59 4.133 ;
      RECT 24.365 3.882 24.595 4.106 ;
      RECT 24.33 4.04 24.595 4.106 ;
      RECT 24.35 3.89 24.49 4.33 ;
      RECT 24.34 3.972 24.6 4.089 ;
      RECT 24.335 4.02 24.6 4.089 ;
      RECT 24.34 3.93 24.595 4.106 ;
      RECT 24.365 3.867 24.59 4.133 ;
      RECT 23.93 3.842 24.1 4.04 ;
      RECT 23.93 3.842 24.145 4.015 ;
      RECT 24 3.785 24.17 3.973 ;
      RECT 23.975 3.8 24.17 3.973 ;
      RECT 23.59 3.846 23.62 4.04 ;
      RECT 23.585 3.818 23.59 4.04 ;
      RECT 23.555 3.792 23.585 4.042 ;
      RECT 23.53 3.75 23.555 4.045 ;
      RECT 23.52 3.722 23.53 4.047 ;
      RECT 23.485 3.702 23.52 4.049 ;
      RECT 23.42 3.687 23.485 4.055 ;
      RECT 23.37 3.685 23.42 4.061 ;
      RECT 23.347 3.687 23.37 4.066 ;
      RECT 23.261 3.698 23.347 4.072 ;
      RECT 23.175 3.716 23.261 4.082 ;
      RECT 23.16 3.727 23.175 4.088 ;
      RECT 23.09 3.75 23.16 4.094 ;
      RECT 23.035 3.782 23.09 4.102 ;
      RECT 22.995 3.805 23.035 4.108 ;
      RECT 22.981 3.818 22.995 4.111 ;
      RECT 22.895 3.84 22.981 4.117 ;
      RECT 22.88 3.865 22.895 4.123 ;
      RECT 22.84 3.88 22.88 4.127 ;
      RECT 22.79 3.895 22.84 4.132 ;
      RECT 22.765 3.902 22.79 4.136 ;
      RECT 22.705 3.897 22.765 4.14 ;
      RECT 22.69 3.888 22.705 4.144 ;
      RECT 22.62 3.878 22.69 4.14 ;
      RECT 22.595 3.87 22.615 4.13 ;
      RECT 22.536 3.87 22.595 4.108 ;
      RECT 22.45 3.87 22.536 4.065 ;
      RECT 22.615 3.87 22.62 4.135 ;
      RECT 23.31 3.101 23.48 3.435 ;
      RECT 23.28 3.101 23.48 3.43 ;
      RECT 23.22 3.068 23.28 3.418 ;
      RECT 23.22 3.124 23.49 3.413 ;
      RECT 23.195 3.124 23.49 3.407 ;
      RECT 23.19 3.065 23.22 3.404 ;
      RECT 23.175 3.071 23.31 3.402 ;
      RECT 23.17 3.079 23.395 3.39 ;
      RECT 23.17 3.131 23.505 3.343 ;
      RECT 23.155 3.087 23.395 3.338 ;
      RECT 23.155 3.157 23.515 3.279 ;
      RECT 23.125 3.107 23.48 3.24 ;
      RECT 23.125 3.197 23.525 3.236 ;
      RECT 23.175 3.076 23.395 3.402 ;
      RECT 22.515 3.406 22.57 3.67 ;
      RECT 22.515 3.406 22.635 3.669 ;
      RECT 22.515 3.406 22.66 3.668 ;
      RECT 22.515 3.406 22.725 3.667 ;
      RECT 22.66 3.372 22.74 3.666 ;
      RECT 22.475 3.416 22.885 3.665 ;
      RECT 22.515 3.413 22.885 3.665 ;
      RECT 22.475 3.421 22.89 3.658 ;
      RECT 22.46 3.423 22.89 3.657 ;
      RECT 22.46 3.43 22.895 3.653 ;
      RECT 22.44 3.429 22.89 3.649 ;
      RECT 22.44 3.437 22.9 3.648 ;
      RECT 22.435 3.434 22.895 3.644 ;
      RECT 22.435 3.447 22.91 3.643 ;
      RECT 22.42 3.437 22.9 3.642 ;
      RECT 22.385 3.45 22.91 3.635 ;
      RECT 22.57 3.405 22.88 3.665 ;
      RECT 22.57 3.39 22.83 3.665 ;
      RECT 22.635 3.377 22.765 3.665 ;
      RECT 22.18 4.466 22.195 4.859 ;
      RECT 22.145 4.471 22.195 4.858 ;
      RECT 22.18 4.47 22.24 4.857 ;
      RECT 22.125 4.481 22.24 4.856 ;
      RECT 22.14 4.477 22.24 4.856 ;
      RECT 22.105 4.487 22.315 4.853 ;
      RECT 22.105 4.506 22.36 4.851 ;
      RECT 22.105 4.513 22.365 4.848 ;
      RECT 22.09 4.49 22.315 4.845 ;
      RECT 22.07 4.495 22.315 4.838 ;
      RECT 22.065 4.499 22.315 4.834 ;
      RECT 22.065 4.516 22.375 4.833 ;
      RECT 22.045 4.51 22.36 4.829 ;
      RECT 22.045 4.519 22.38 4.823 ;
      RECT 22.04 4.525 22.38 4.595 ;
      RECT 22.105 4.485 22.24 4.853 ;
      RECT 21.98 3.848 22.18 4.16 ;
      RECT 22.055 3.826 22.18 4.16 ;
      RECT 21.995 3.845 22.185 4.145 ;
      RECT 21.965 3.856 22.185 4.143 ;
      RECT 21.98 3.851 22.19 4.109 ;
      RECT 21.965 3.955 22.195 4.076 ;
      RECT 21.995 3.827 22.18 4.16 ;
      RECT 22.055 3.805 22.155 4.16 ;
      RECT 22.08 3.802 22.155 4.16 ;
      RECT 22.08 3.797 22.1 4.16 ;
      RECT 21.485 3.865 21.66 4.04 ;
      RECT 21.48 3.865 21.66 4.038 ;
      RECT 21.455 3.865 21.66 4.033 ;
      RECT 21.4 3.845 21.57 4.023 ;
      RECT 21.4 3.852 21.635 4.023 ;
      RECT 21.485 4.532 21.5 4.715 ;
      RECT 21.475 4.51 21.485 4.715 ;
      RECT 21.46 4.49 21.475 4.715 ;
      RECT 21.45 4.465 21.46 4.715 ;
      RECT 21.42 4.43 21.45 4.715 ;
      RECT 21.385 4.37 21.42 4.715 ;
      RECT 21.38 4.332 21.385 4.715 ;
      RECT 21.33 4.283 21.38 4.715 ;
      RECT 21.32 4.233 21.33 4.703 ;
      RECT 21.305 4.212 21.32 4.663 ;
      RECT 21.285 4.18 21.305 4.613 ;
      RECT 21.26 4.136 21.285 4.553 ;
      RECT 21.255 4.108 21.26 4.508 ;
      RECT 21.25 4.099 21.255 4.494 ;
      RECT 21.245 4.092 21.25 4.481 ;
      RECT 21.24 4.087 21.245 4.47 ;
      RECT 21.235 4.072 21.24 4.46 ;
      RECT 21.23 4.05 21.235 4.447 ;
      RECT 21.22 4.01 21.23 4.422 ;
      RECT 21.195 3.94 21.22 4.378 ;
      RECT 21.19 3.88 21.195 4.343 ;
      RECT 21.175 3.86 21.19 4.31 ;
      RECT 21.17 3.86 21.175 4.285 ;
      RECT 21.14 3.86 21.17 4.24 ;
      RECT 21.095 3.86 21.14 4.18 ;
      RECT 21.02 3.86 21.095 4.128 ;
      RECT 21.015 3.86 21.02 4.093 ;
      RECT 21.01 3.86 21.015 4.083 ;
      RECT 21.005 3.86 21.01 4.063 ;
      RECT 21.27 3.08 21.44 3.55 ;
      RECT 21.215 3.073 21.41 3.534 ;
      RECT 21.215 3.087 21.445 3.533 ;
      RECT 21.2 3.088 21.445 3.514 ;
      RECT 21.195 3.106 21.445 3.5 ;
      RECT 21.2 3.089 21.45 3.498 ;
      RECT 21.185 3.12 21.45 3.483 ;
      RECT 21.2 3.095 21.455 3.468 ;
      RECT 21.18 3.135 21.455 3.465 ;
      RECT 21.195 3.107 21.46 3.45 ;
      RECT 21.195 3.119 21.465 3.43 ;
      RECT 21.18 3.135 21.47 3.413 ;
      RECT 21.18 3.145 21.475 3.268 ;
      RECT 21.175 3.145 21.475 3.225 ;
      RECT 21.175 3.16 21.48 3.203 ;
      RECT 21.27 3.07 21.41 3.55 ;
      RECT 21.27 3.068 21.38 3.55 ;
      RECT 21.356 3.065 21.38 3.55 ;
      RECT 21.015 4.732 21.02 4.778 ;
      RECT 21.005 4.58 21.015 4.802 ;
      RECT 21 4.425 21.005 4.827 ;
      RECT 20.985 4.387 21 4.838 ;
      RECT 20.98 4.37 20.985 4.845 ;
      RECT 20.97 4.358 20.98 4.852 ;
      RECT 20.965 4.349 20.97 4.854 ;
      RECT 20.96 4.347 20.965 4.858 ;
      RECT 20.915 4.338 20.96 4.873 ;
      RECT 20.91 4.33 20.915 4.887 ;
      RECT 20.905 4.327 20.91 4.891 ;
      RECT 20.89 4.322 20.905 4.899 ;
      RECT 20.835 4.312 20.89 4.91 ;
      RECT 20.8 4.3 20.835 4.911 ;
      RECT 20.791 4.295 20.8 4.905 ;
      RECT 20.705 4.295 20.791 4.895 ;
      RECT 20.675 4.295 20.705 4.873 ;
      RECT 20.665 4.295 20.67 4.853 ;
      RECT 20.66 4.295 20.665 4.815 ;
      RECT 20.655 4.295 20.66 4.773 ;
      RECT 20.65 4.295 20.655 4.733 ;
      RECT 20.645 4.295 20.65 4.663 ;
      RECT 20.635 4.295 20.645 4.585 ;
      RECT 20.63 4.295 20.635 4.485 ;
      RECT 20.67 4.295 20.675 4.855 ;
      RECT 20.165 4.377 20.255 4.855 ;
      RECT 20.15 4.38 20.27 4.853 ;
      RECT 20.165 4.379 20.27 4.853 ;
      RECT 20.13 4.386 20.295 4.843 ;
      RECT 20.15 4.38 20.295 4.843 ;
      RECT 20.115 4.392 20.295 4.831 ;
      RECT 20.15 4.383 20.345 4.824 ;
      RECT 20.101 4.4 20.345 4.822 ;
      RECT 20.13 4.39 20.355 4.81 ;
      RECT 20.101 4.411 20.385 4.801 ;
      RECT 20.015 4.435 20.385 4.795 ;
      RECT 20.015 4.448 20.425 4.778 ;
      RECT 20.01 4.47 20.425 4.771 ;
      RECT 19.98 4.485 20.425 4.761 ;
      RECT 19.975 4.496 20.425 4.751 ;
      RECT 19.945 4.509 20.425 4.742 ;
      RECT 19.93 4.527 20.425 4.731 ;
      RECT 19.905 4.54 20.425 4.721 ;
      RECT 20.165 4.376 20.175 4.855 ;
      RECT 20.211 3.8 20.25 4.045 ;
      RECT 20.125 3.8 20.26 4.043 ;
      RECT 20.01 3.825 20.26 4.04 ;
      RECT 20.01 3.825 20.265 4.038 ;
      RECT 20.01 3.825 20.28 4.033 ;
      RECT 20.116 3.8 20.295 4.013 ;
      RECT 20.03 3.808 20.295 4.013 ;
      RECT 19.7 3.16 19.87 3.595 ;
      RECT 19.69 3.194 19.87 3.578 ;
      RECT 19.77 3.13 19.94 3.565 ;
      RECT 19.675 3.205 19.94 3.543 ;
      RECT 19.77 3.14 19.945 3.533 ;
      RECT 19.7 3.192 19.975 3.518 ;
      RECT 19.66 3.218 19.975 3.503 ;
      RECT 19.66 3.26 19.985 3.483 ;
      RECT 19.655 3.285 19.99 3.465 ;
      RECT 19.655 3.295 19.995 3.45 ;
      RECT 19.65 3.232 19.975 3.448 ;
      RECT 19.65 3.305 20 3.433 ;
      RECT 19.645 3.242 19.975 3.43 ;
      RECT 19.64 3.326 20.005 3.413 ;
      RECT 19.64 3.358 20.01 3.393 ;
      RECT 19.635 3.272 19.985 3.385 ;
      RECT 19.64 3.257 19.975 3.413 ;
      RECT 19.655 3.227 19.975 3.465 ;
      RECT 19.5 3.814 19.725 4.07 ;
      RECT 19.5 3.847 19.745 4.06 ;
      RECT 19.465 3.847 19.745 4.058 ;
      RECT 19.465 3.86 19.75 4.048 ;
      RECT 19.465 3.88 19.76 4.04 ;
      RECT 19.465 3.977 19.765 4.033 ;
      RECT 19.445 3.725 19.575 4.023 ;
      RECT 19.4 3.88 19.76 3.965 ;
      RECT 19.39 3.725 19.575 3.91 ;
      RECT 19.39 3.757 19.661 3.91 ;
      RECT 19.355 4.287 19.375 4.465 ;
      RECT 19.32 4.24 19.355 4.465 ;
      RECT 19.305 4.18 19.32 4.465 ;
      RECT 19.28 4.127 19.305 4.465 ;
      RECT 19.265 4.08 19.28 4.465 ;
      RECT 19.245 4.057 19.265 4.465 ;
      RECT 19.22 4.022 19.245 4.465 ;
      RECT 19.21 3.868 19.22 4.465 ;
      RECT 19.18 3.863 19.21 4.456 ;
      RECT 19.175 3.86 19.18 4.446 ;
      RECT 19.16 3.86 19.175 4.42 ;
      RECT 19.155 3.86 19.16 4.383 ;
      RECT 19.13 3.86 19.155 4.335 ;
      RECT 19.11 3.86 19.13 4.26 ;
      RECT 19.1 3.86 19.11 4.22 ;
      RECT 19.095 3.86 19.1 4.195 ;
      RECT 19.09 3.86 19.095 4.178 ;
      RECT 19.085 3.86 19.09 4.16 ;
      RECT 19.08 3.861 19.085 4.15 ;
      RECT 19.07 3.863 19.08 4.118 ;
      RECT 19.06 3.865 19.07 4.085 ;
      RECT 19.05 3.868 19.06 4.058 ;
      RECT 19.375 4.295 19.6 4.465 ;
      RECT 18.705 3.107 18.875 3.56 ;
      RECT 18.705 3.107 18.965 3.526 ;
      RECT 18.705 3.107 18.995 3.51 ;
      RECT 18.705 3.107 19.025 3.483 ;
      RECT 18.961 3.085 19.04 3.465 ;
      RECT 18.74 3.092 19.045 3.45 ;
      RECT 18.74 3.1 19.055 3.413 ;
      RECT 18.7 3.127 19.055 3.385 ;
      RECT 18.685 3.14 19.055 3.35 ;
      RECT 18.705 3.115 19.075 3.34 ;
      RECT 18.68 3.18 19.075 3.31 ;
      RECT 18.68 3.21 19.08 3.293 ;
      RECT 18.675 3.24 19.08 3.28 ;
      RECT 18.74 3.089 19.04 3.465 ;
      RECT 18.875 3.086 18.961 3.544 ;
      RECT 18.826 3.087 19.04 3.465 ;
      RECT 18.97 4.747 19.015 4.94 ;
      RECT 18.96 4.717 18.97 4.94 ;
      RECT 18.955 4.702 18.96 4.94 ;
      RECT 18.915 4.612 18.955 4.94 ;
      RECT 18.91 4.525 18.915 4.94 ;
      RECT 18.9 4.495 18.91 4.94 ;
      RECT 18.895 4.455 18.9 4.94 ;
      RECT 18.885 4.417 18.895 4.94 ;
      RECT 18.88 4.382 18.885 4.94 ;
      RECT 18.86 4.335 18.88 4.94 ;
      RECT 18.845 4.26 18.86 4.94 ;
      RECT 18.84 4.215 18.845 4.935 ;
      RECT 18.835 4.195 18.84 4.908 ;
      RECT 18.83 4.175 18.835 4.893 ;
      RECT 18.825 4.15 18.83 4.873 ;
      RECT 18.82 4.128 18.825 4.858 ;
      RECT 18.815 4.106 18.82 4.84 ;
      RECT 18.81 4.085 18.815 4.83 ;
      RECT 18.8 4.057 18.81 4.8 ;
      RECT 18.79 4.02 18.8 4.768 ;
      RECT 18.78 3.98 18.79 4.735 ;
      RECT 18.77 3.958 18.78 4.705 ;
      RECT 18.74 3.91 18.77 4.637 ;
      RECT 18.725 3.87 18.74 4.564 ;
      RECT 18.715 3.87 18.725 4.53 ;
      RECT 18.71 3.87 18.715 4.505 ;
      RECT 18.705 3.87 18.71 4.49 ;
      RECT 18.7 3.87 18.705 4.468 ;
      RECT 18.695 3.87 18.7 4.455 ;
      RECT 18.68 3.87 18.695 4.42 ;
      RECT 18.66 3.87 18.68 4.36 ;
      RECT 18.65 3.87 18.66 4.31 ;
      RECT 18.63 3.87 18.65 4.258 ;
      RECT 18.61 3.87 18.63 4.215 ;
      RECT 18.6 3.87 18.61 4.203 ;
      RECT 18.57 3.87 18.6 4.19 ;
      RECT 18.54 3.891 18.57 4.17 ;
      RECT 18.53 3.919 18.54 4.15 ;
      RECT 18.515 3.936 18.53 4.118 ;
      RECT 18.51 3.95 18.515 4.085 ;
      RECT 18.505 3.958 18.51 4.058 ;
      RECT 18.5 3.966 18.505 4.02 ;
      RECT 18.505 4.49 18.51 4.825 ;
      RECT 18.47 4.477 18.505 4.824 ;
      RECT 18.4 4.417 18.47 4.823 ;
      RECT 18.32 4.36 18.4 4.822 ;
      RECT 18.185 4.32 18.32 4.821 ;
      RECT 18.185 4.507 18.52 4.81 ;
      RECT 18.145 4.507 18.52 4.8 ;
      RECT 18.145 4.525 18.525 4.795 ;
      RECT 18.145 4.615 18.53 4.785 ;
      RECT 18.14 4.31 18.305 4.765 ;
      RECT 18.135 4.31 18.305 4.508 ;
      RECT 18.135 4.467 18.5 4.508 ;
      RECT 18.135 4.455 18.495 4.508 ;
      RECT 16.6 7.305 16.77 9.515 ;
      RECT 16.6 7.305 16.775 8.565 ;
      RECT 16.17 10.145 16.34 10.595 ;
      RECT 16.23 8.365 16.4 10.315 ;
      RECT 16.17 7.305 16.34 8.535 ;
      RECT 15.645 10.105 15.82 10.595 ;
      RECT 15.645 7.305 15.815 10.595 ;
      RECT 15.645 9.605 16.055 9.935 ;
      RECT 15.645 8.765 16.055 9.095 ;
      RECT 15.645 7.305 15.82 8.565 ;
      RECT 96.18 10.08 96.355 10.59 ;
      RECT 95.185 1.865 95.36 2.375 ;
      RECT 95.185 10.085 95.36 10.595 ;
      RECT 93.395 1.865 93.57 2.375 ;
      RECT 93.395 10.085 93.57 10.595 ;
      RECT 91.005 4.145 91.375 4.515 ;
      RECT 88.615 10.085 88.79 10.595 ;
      RECT 80.395 10.08 80.57 10.59 ;
      RECT 79.4 1.865 79.575 2.375 ;
      RECT 79.4 10.085 79.575 10.595 ;
      RECT 77.61 1.865 77.785 2.375 ;
      RECT 77.61 10.085 77.785 10.595 ;
      RECT 75.22 4.145 75.59 4.515 ;
      RECT 72.83 10.085 73.005 10.595 ;
      RECT 64.61 10.08 64.785 10.59 ;
      RECT 63.615 1.865 63.79 2.375 ;
      RECT 63.615 10.085 63.79 10.595 ;
      RECT 61.825 1.865 62 2.375 ;
      RECT 61.825 10.085 62 10.595 ;
      RECT 59.435 4.145 59.805 4.515 ;
      RECT 57.045 10.085 57.22 10.595 ;
      RECT 48.835 10.08 49.01 10.59 ;
      RECT 47.84 1.865 48.015 2.375 ;
      RECT 47.84 10.085 48.015 10.595 ;
      RECT 46.05 1.865 46.225 2.375 ;
      RECT 46.05 10.085 46.225 10.595 ;
      RECT 43.66 4.145 44.03 4.515 ;
      RECT 41.27 10.085 41.445 10.595 ;
      RECT 33.055 10.08 33.23 10.59 ;
      RECT 32.06 1.865 32.235 2.375 ;
      RECT 32.06 10.085 32.235 10.595 ;
      RECT 30.27 1.865 30.445 2.375 ;
      RECT 30.27 10.085 30.445 10.595 ;
      RECT 27.88 4.145 28.25 4.515 ;
      RECT 25.49 10.085 25.665 10.595 ;
      RECT 16.6 10.085 16.775 10.595 ;
  END
END sky130_osu_ring_oscillator_mpr2aa_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2aa_8_b0r2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2aa_8_b0r2 ;
  SIZE 96.775 BY 12.46 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 33.05 0 33.43 3.06 ;
      LAYER li1 ;
        RECT 33.095 1.865 33.27 2.375 ;
        RECT 33.095 3.895 33.27 5.155 ;
        RECT 33.095 3.685 33.265 5.155 ;
      LAYER met2 ;
        RECT 33.05 2.68 33.43 3.06 ;
      LAYER met1 ;
        RECT 33.095 2.725 33.415 3.015 ;
        RECT 33.035 2.175 33.33 2.405 ;
        RECT 33.035 3.655 33.325 3.885 ;
        RECT 33.095 2.175 33.265 3.885 ;
      LAYER via1 ;
        RECT 33.165 2.795 33.315 2.945 ;
      LAYER via2 ;
        RECT 33.14 2.77 33.34 2.97 ;
      LAYER mcon ;
        RECT 33.095 3.685 33.265 3.855 ;
        RECT 33.095 2.205 33.27 2.375 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 48.83 0 49.21 3.06 ;
      LAYER li1 ;
        RECT 48.875 1.865 49.05 2.375 ;
        RECT 48.875 3.895 49.05 5.155 ;
        RECT 48.875 3.685 49.045 5.155 ;
      LAYER met2 ;
        RECT 48.83 2.68 49.21 3.06 ;
      LAYER met1 ;
        RECT 48.875 2.725 49.195 3.015 ;
        RECT 48.815 2.175 49.11 2.405 ;
        RECT 48.815 3.655 49.105 3.885 ;
        RECT 48.875 2.175 49.045 3.885 ;
      LAYER via1 ;
        RECT 48.945 2.795 49.095 2.945 ;
      LAYER via2 ;
        RECT 48.92 2.77 49.12 2.97 ;
      LAYER mcon ;
        RECT 48.875 3.685 49.045 3.855 ;
        RECT 48.875 2.205 49.05 2.375 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 64.605 0 64.985 3.06 ;
      LAYER li1 ;
        RECT 64.65 1.865 64.825 2.375 ;
        RECT 64.65 3.895 64.825 5.155 ;
        RECT 64.65 3.685 64.82 5.155 ;
      LAYER met2 ;
        RECT 64.605 2.68 64.985 3.06 ;
      LAYER met1 ;
        RECT 64.65 2.725 64.97 3.015 ;
        RECT 64.59 2.175 64.885 2.405 ;
        RECT 64.59 3.655 64.88 3.885 ;
        RECT 64.65 2.175 64.82 3.885 ;
      LAYER via1 ;
        RECT 64.72 2.795 64.87 2.945 ;
      LAYER via2 ;
        RECT 64.695 2.77 64.895 2.97 ;
      LAYER mcon ;
        RECT 64.65 3.685 64.82 3.855 ;
        RECT 64.65 2.205 64.825 2.375 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 80.39 0 80.77 3.06 ;
      LAYER li1 ;
        RECT 80.435 1.865 80.61 2.375 ;
        RECT 80.435 3.895 80.61 5.155 ;
        RECT 80.435 3.685 80.605 5.155 ;
      LAYER met2 ;
        RECT 80.39 2.68 80.77 3.06 ;
      LAYER met1 ;
        RECT 80.435 2.725 80.755 3.015 ;
        RECT 80.375 2.175 80.67 2.405 ;
        RECT 80.375 3.655 80.665 3.885 ;
        RECT 80.435 2.175 80.605 3.885 ;
      LAYER via1 ;
        RECT 80.505 2.795 80.655 2.945 ;
      LAYER via2 ;
        RECT 80.48 2.77 80.68 2.97 ;
      LAYER mcon ;
        RECT 80.435 3.685 80.605 3.855 ;
        RECT 80.435 2.205 80.61 2.375 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 96.175 0 96.555 3.06 ;
      LAYER li1 ;
        RECT 96.22 1.865 96.395 2.375 ;
        RECT 96.22 3.895 96.395 5.155 ;
        RECT 96.22 3.685 96.39 5.155 ;
      LAYER met2 ;
        RECT 96.175 2.68 96.555 3.06 ;
      LAYER met1 ;
        RECT 96.22 2.725 96.54 3.015 ;
        RECT 96.16 2.175 96.455 2.405 ;
        RECT 96.16 3.655 96.45 3.885 ;
        RECT 96.22 2.175 96.39 3.885 ;
      LAYER via1 ;
        RECT 96.29 2.795 96.44 2.945 ;
      LAYER via2 ;
        RECT 96.265 2.77 96.465 2.97 ;
      LAYER mcon ;
        RECT 96.22 3.685 96.39 3.855 ;
        RECT 96.22 2.205 96.395 2.375 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 28.945 2.955 29.115 4.225 ;
        RECT 28.945 8.235 29.115 9.505 ;
        RECT 24.165 8.235 24.335 9.505 ;
      LAYER met2 ;
        RECT 28.865 8.14 29.215 8.49 ;
        RECT 28.86 4 29.21 4.35 ;
        RECT 28.935 4 29.11 8.49 ;
      LAYER met1 ;
        RECT 28.86 4.055 29.345 4.225 ;
        RECT 28.86 4 29.21 4.35 ;
        RECT 28.865 8.235 29.345 8.405 ;
        RECT 28.865 8.14 29.215 8.49 ;
        RECT 24.4 8.23 29.215 8.4 ;
        RECT 24.105 8.235 24.565 8.405 ;
        RECT 24.105 8.205 24.395 8.435 ;
      LAYER via1 ;
        RECT 28.96 4.1 29.11 4.25 ;
        RECT 28.965 8.24 29.115 8.39 ;
      LAYER mcon ;
        RECT 24.165 8.235 24.335 8.405 ;
        RECT 28.945 8.235 29.115 8.405 ;
        RECT 28.945 4.055 29.115 4.225 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 44.725 2.955 44.895 4.225 ;
        RECT 44.725 8.235 44.895 9.505 ;
        RECT 39.945 8.235 40.115 9.505 ;
      LAYER met2 ;
        RECT 44.645 8.14 44.995 8.49 ;
        RECT 44.64 4 44.99 4.35 ;
        RECT 44.715 4 44.89 8.49 ;
      LAYER met1 ;
        RECT 44.64 4.055 45.125 4.225 ;
        RECT 44.64 4 44.99 4.35 ;
        RECT 44.645 8.235 45.125 8.405 ;
        RECT 44.645 8.14 44.995 8.49 ;
        RECT 40.18 8.23 44.995 8.4 ;
        RECT 39.885 8.235 40.345 8.405 ;
        RECT 39.885 8.205 40.175 8.435 ;
      LAYER via1 ;
        RECT 44.74 4.1 44.89 4.25 ;
        RECT 44.745 8.24 44.895 8.39 ;
      LAYER mcon ;
        RECT 39.945 8.235 40.115 8.405 ;
        RECT 44.725 8.235 44.895 8.405 ;
        RECT 44.725 4.055 44.895 4.225 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 60.5 2.955 60.67 4.225 ;
        RECT 60.5 8.235 60.67 9.505 ;
        RECT 55.72 8.235 55.89 9.505 ;
      LAYER met2 ;
        RECT 60.42 8.14 60.77 8.49 ;
        RECT 60.415 4 60.765 4.35 ;
        RECT 60.49 4 60.665 8.49 ;
      LAYER met1 ;
        RECT 60.415 4.055 60.9 4.225 ;
        RECT 60.415 4 60.765 4.35 ;
        RECT 60.42 8.235 60.9 8.405 ;
        RECT 60.42 8.14 60.77 8.49 ;
        RECT 55.955 8.23 60.77 8.4 ;
        RECT 55.66 8.235 56.12 8.405 ;
        RECT 55.66 8.205 55.95 8.435 ;
      LAYER via1 ;
        RECT 60.515 4.1 60.665 4.25 ;
        RECT 60.52 8.24 60.67 8.39 ;
      LAYER mcon ;
        RECT 55.72 8.235 55.89 8.405 ;
        RECT 60.5 8.235 60.67 8.405 ;
        RECT 60.5 4.055 60.67 4.225 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 76.285 2.955 76.455 4.225 ;
        RECT 76.285 8.235 76.455 9.505 ;
        RECT 71.505 8.235 71.675 9.505 ;
      LAYER met2 ;
        RECT 76.205 8.14 76.555 8.49 ;
        RECT 76.2 4 76.55 4.35 ;
        RECT 76.275 4 76.45 8.49 ;
      LAYER met1 ;
        RECT 76.2 4.055 76.685 4.225 ;
        RECT 76.2 4 76.55 4.35 ;
        RECT 76.205 8.235 76.685 8.405 ;
        RECT 76.205 8.14 76.555 8.49 ;
        RECT 71.74 8.23 76.555 8.4 ;
        RECT 71.445 8.235 71.905 8.405 ;
        RECT 71.445 8.205 71.735 8.435 ;
      LAYER via1 ;
        RECT 76.3 4.1 76.45 4.25 ;
        RECT 76.305 8.24 76.455 8.39 ;
      LAYER mcon ;
        RECT 71.505 8.235 71.675 8.405 ;
        RECT 76.285 8.235 76.455 8.405 ;
        RECT 76.285 4.055 76.455 4.225 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 92.07 2.955 92.24 4.225 ;
        RECT 92.07 8.235 92.24 9.505 ;
        RECT 87.29 8.235 87.46 9.505 ;
      LAYER met2 ;
        RECT 91.99 8.14 92.34 8.49 ;
        RECT 91.985 4 92.335 4.35 ;
        RECT 92.06 4 92.235 8.49 ;
      LAYER met1 ;
        RECT 91.985 4.055 92.47 4.225 ;
        RECT 91.985 4 92.335 4.35 ;
        RECT 91.99 8.235 92.47 8.405 ;
        RECT 91.99 8.14 92.34 8.49 ;
        RECT 87.525 8.23 92.34 8.4 ;
        RECT 87.23 8.235 87.69 8.405 ;
        RECT 87.23 8.205 87.52 8.435 ;
      LAYER via1 ;
        RECT 92.085 4.1 92.235 4.25 ;
        RECT 92.09 8.24 92.24 8.39 ;
      LAYER mcon ;
        RECT 87.29 8.235 87.46 8.405 ;
        RECT 92.07 8.235 92.24 8.405 ;
        RECT 92.07 4.055 92.24 4.225 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 15.29 8.235 15.46 9.505 ;
      LAYER met1 ;
        RECT 15.175 8.235 15.69 8.405 ;
        RECT 15.23 8.205 15.52 8.435 ;
        RECT 15.175 8.2 15.465 8.43 ;
      LAYER mcon ;
        RECT 15.29 8.235 15.46 8.405 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.005 5.43 96.77 7.03 ;
        RECT 91.89 5.43 96.615 7.035 ;
        RECT 91.89 5.425 96.61 7.035 ;
        RECT 95.795 5.425 95.965 7.765 ;
        RECT 95.79 4.695 95.96 7.035 ;
        RECT 94.805 4.695 94.975 7.765 ;
        RECT 92.06 4.695 92.23 7.765 ;
        RECT 90.265 4.93 90.435 7.03 ;
        RECT 87.11 5.43 89.86 7.035 ;
        RECT 89.305 4.93 89.475 7.035 ;
        RECT 87.28 5.43 87.45 7.765 ;
        RECT 86.865 4.93 87.035 7.03 ;
        RECT 85.865 4.93 86.035 7.03 ;
        RECT 84.905 4.93 85.075 7.03 ;
        RECT 82.465 4.93 82.635 7.03 ;
        RECT 76.105 5.43 80.83 7.035 ;
        RECT 76.105 5.425 80.825 7.035 ;
        RECT 80.01 5.425 80.18 7.765 ;
        RECT 80.005 4.695 80.175 7.035 ;
        RECT 79.02 4.695 79.19 7.765 ;
        RECT 76.275 4.695 76.445 7.765 ;
        RECT 74.48 4.93 74.65 7.03 ;
        RECT 71.325 5.43 74.075 7.035 ;
        RECT 73.52 4.93 73.69 7.035 ;
        RECT 71.495 5.43 71.665 7.765 ;
        RECT 71.08 4.93 71.25 7.03 ;
        RECT 70.08 4.93 70.25 7.03 ;
        RECT 69.12 4.93 69.29 7.03 ;
        RECT 66.68 4.93 66.85 7.03 ;
        RECT 60.32 5.43 65.225 7.035 ;
        RECT 60.32 5.425 65.04 7.035 ;
        RECT 64.225 5.425 64.395 7.765 ;
        RECT 64.22 4.695 64.39 7.035 ;
        RECT 63.235 4.695 63.405 7.765 ;
        RECT 60.49 4.695 60.66 7.765 ;
        RECT 58.695 4.93 58.865 7.03 ;
        RECT 55.54 5.43 58.29 7.035 ;
        RECT 57.735 4.93 57.905 7.035 ;
        RECT 55.71 5.43 55.88 7.765 ;
        RECT 55.295 4.93 55.465 7.03 ;
        RECT 54.295 4.93 54.465 7.03 ;
        RECT 53.335 4.93 53.505 7.03 ;
        RECT 50.895 4.93 51.065 7.03 ;
        RECT 44.545 5.43 49.27 7.035 ;
        RECT 44.545 5.425 49.265 7.035 ;
        RECT 48.45 5.425 48.62 7.765 ;
        RECT 48.445 4.695 48.615 7.035 ;
        RECT 47.46 4.695 47.63 7.765 ;
        RECT 44.715 4.695 44.885 7.765 ;
        RECT 42.92 4.93 43.09 7.03 ;
        RECT 39.765 5.43 42.515 7.035 ;
        RECT 41.96 4.93 42.13 7.035 ;
        RECT 39.935 5.43 40.105 7.765 ;
        RECT 39.52 4.93 39.69 7.03 ;
        RECT 38.52 4.93 38.69 7.03 ;
        RECT 37.56 4.93 37.73 7.03 ;
        RECT 35.12 4.93 35.29 7.03 ;
        RECT 28.765 5.43 33.49 7.035 ;
        RECT 28.765 5.425 33.485 7.035 ;
        RECT 32.67 5.425 32.84 7.765 ;
        RECT 32.665 4.695 32.835 7.035 ;
        RECT 31.68 4.695 31.85 7.765 ;
        RECT 28.935 4.695 29.105 7.765 ;
        RECT 27.14 4.93 27.31 7.03 ;
        RECT 23.985 5.43 26.735 7.035 ;
        RECT 26.18 4.93 26.35 7.035 ;
        RECT 24.155 5.43 24.325 7.765 ;
        RECT 23.74 4.93 23.91 7.03 ;
        RECT 22.74 4.93 22.91 7.03 ;
        RECT 21.78 4.93 21.95 7.03 ;
        RECT 19.34 4.93 19.51 7.03 ;
        RECT 15.11 5.43 17.86 7.035 ;
        RECT 17.095 10.045 17.27 10.595 ;
        RECT 17.095 7.305 17.27 8.445 ;
        RECT 17.095 5.43 17.265 10.595 ;
        RECT 15.28 5.43 15.45 7.765 ;
      LAYER met1 ;
        RECT 0.005 5.43 96.77 7.03 ;
        RECT 91.89 5.43 96.615 7.035 ;
        RECT 91.89 5.425 96.61 7.035 ;
        RECT 81.175 5.275 90.835 7.03 ;
        RECT 87.11 5.275 89.86 7.035 ;
        RECT 76.105 5.43 80.83 7.035 ;
        RECT 76.105 5.425 80.825 7.035 ;
        RECT 65.39 5.275 75.05 7.03 ;
        RECT 71.325 5.275 74.075 7.035 ;
        RECT 60.32 5.43 65.225 7.035 ;
        RECT 60.32 5.425 65.04 7.035 ;
        RECT 49.605 5.275 59.265 7.03 ;
        RECT 55.54 5.275 58.29 7.035 ;
        RECT 44.545 5.43 49.27 7.035 ;
        RECT 44.545 5.425 49.265 7.035 ;
        RECT 33.83 5.275 43.49 7.03 ;
        RECT 39.765 5.275 42.515 7.035 ;
        RECT 28.765 5.43 33.49 7.035 ;
        RECT 28.765 5.425 33.485 7.035 ;
        RECT 18.05 5.275 27.71 7.03 ;
        RECT 23.985 5.275 26.735 7.035 ;
        RECT 15.11 5.43 17.86 7.035 ;
        RECT 17.035 8.945 17.325 9.175 ;
        RECT 16.865 8.975 17.325 9.145 ;
      LAYER mcon ;
        RECT 17.095 8.975 17.265 9.145 ;
        RECT 17.4 6.835 17.57 7.005 ;
        RECT 18.195 5.43 18.365 5.6 ;
        RECT 18.655 5.43 18.825 5.6 ;
        RECT 19.115 5.43 19.285 5.6 ;
        RECT 19.575 5.43 19.745 5.6 ;
        RECT 20.035 5.43 20.205 5.6 ;
        RECT 20.495 5.43 20.665 5.6 ;
        RECT 20.955 5.43 21.125 5.6 ;
        RECT 21.415 5.43 21.585 5.6 ;
        RECT 21.875 5.43 22.045 5.6 ;
        RECT 22.335 5.43 22.505 5.6 ;
        RECT 22.795 5.43 22.965 5.6 ;
        RECT 23.255 5.43 23.425 5.6 ;
        RECT 23.715 5.43 23.885 5.6 ;
        RECT 24.175 5.43 24.345 5.6 ;
        RECT 24.635 5.43 24.805 5.6 ;
        RECT 25.095 5.43 25.265 5.6 ;
        RECT 25.555 5.43 25.725 5.6 ;
        RECT 26.015 5.43 26.185 5.6 ;
        RECT 26.275 6.835 26.445 7.005 ;
        RECT 26.475 5.43 26.645 5.6 ;
        RECT 26.935 5.43 27.105 5.6 ;
        RECT 27.395 5.43 27.565 5.6 ;
        RECT 31.055 6.835 31.225 7.005 ;
        RECT 31.055 5.455 31.225 5.625 ;
        RECT 31.76 6.835 31.93 7.005 ;
        RECT 31.76 5.455 31.93 5.625 ;
        RECT 32.745 5.455 32.915 5.625 ;
        RECT 32.75 6.835 32.92 7.005 ;
        RECT 33.975 5.43 34.145 5.6 ;
        RECT 34.435 5.43 34.605 5.6 ;
        RECT 34.895 5.43 35.065 5.6 ;
        RECT 35.355 5.43 35.525 5.6 ;
        RECT 35.815 5.43 35.985 5.6 ;
        RECT 36.275 5.43 36.445 5.6 ;
        RECT 36.735 5.43 36.905 5.6 ;
        RECT 37.195 5.43 37.365 5.6 ;
        RECT 37.655 5.43 37.825 5.6 ;
        RECT 38.115 5.43 38.285 5.6 ;
        RECT 38.575 5.43 38.745 5.6 ;
        RECT 39.035 5.43 39.205 5.6 ;
        RECT 39.495 5.43 39.665 5.6 ;
        RECT 39.955 5.43 40.125 5.6 ;
        RECT 40.415 5.43 40.585 5.6 ;
        RECT 40.875 5.43 41.045 5.6 ;
        RECT 41.335 5.43 41.505 5.6 ;
        RECT 41.795 5.43 41.965 5.6 ;
        RECT 42.055 6.835 42.225 7.005 ;
        RECT 42.255 5.43 42.425 5.6 ;
        RECT 42.715 5.43 42.885 5.6 ;
        RECT 43.175 5.43 43.345 5.6 ;
        RECT 46.835 6.835 47.005 7.005 ;
        RECT 46.835 5.455 47.005 5.625 ;
        RECT 47.54 6.835 47.71 7.005 ;
        RECT 47.54 5.455 47.71 5.625 ;
        RECT 48.525 5.455 48.695 5.625 ;
        RECT 48.53 6.835 48.7 7.005 ;
        RECT 49.75 5.43 49.92 5.6 ;
        RECT 50.21 5.43 50.38 5.6 ;
        RECT 50.67 5.43 50.84 5.6 ;
        RECT 51.13 5.43 51.3 5.6 ;
        RECT 51.59 5.43 51.76 5.6 ;
        RECT 52.05 5.43 52.22 5.6 ;
        RECT 52.51 5.43 52.68 5.6 ;
        RECT 52.97 5.43 53.14 5.6 ;
        RECT 53.43 5.43 53.6 5.6 ;
        RECT 53.89 5.43 54.06 5.6 ;
        RECT 54.35 5.43 54.52 5.6 ;
        RECT 54.81 5.43 54.98 5.6 ;
        RECT 55.27 5.43 55.44 5.6 ;
        RECT 55.73 5.43 55.9 5.6 ;
        RECT 56.19 5.43 56.36 5.6 ;
        RECT 56.65 5.43 56.82 5.6 ;
        RECT 57.11 5.43 57.28 5.6 ;
        RECT 57.57 5.43 57.74 5.6 ;
        RECT 57.83 6.835 58 7.005 ;
        RECT 58.03 5.43 58.2 5.6 ;
        RECT 58.49 5.43 58.66 5.6 ;
        RECT 58.95 5.43 59.12 5.6 ;
        RECT 62.61 6.835 62.78 7.005 ;
        RECT 62.61 5.455 62.78 5.625 ;
        RECT 63.315 6.835 63.485 7.005 ;
        RECT 63.315 5.455 63.485 5.625 ;
        RECT 64.3 5.455 64.47 5.625 ;
        RECT 64.305 6.835 64.475 7.005 ;
        RECT 65.535 5.43 65.705 5.6 ;
        RECT 65.995 5.43 66.165 5.6 ;
        RECT 66.455 5.43 66.625 5.6 ;
        RECT 66.915 5.43 67.085 5.6 ;
        RECT 67.375 5.43 67.545 5.6 ;
        RECT 67.835 5.43 68.005 5.6 ;
        RECT 68.295 5.43 68.465 5.6 ;
        RECT 68.755 5.43 68.925 5.6 ;
        RECT 69.215 5.43 69.385 5.6 ;
        RECT 69.675 5.43 69.845 5.6 ;
        RECT 70.135 5.43 70.305 5.6 ;
        RECT 70.595 5.43 70.765 5.6 ;
        RECT 71.055 5.43 71.225 5.6 ;
        RECT 71.515 5.43 71.685 5.6 ;
        RECT 71.975 5.43 72.145 5.6 ;
        RECT 72.435 5.43 72.605 5.6 ;
        RECT 72.895 5.43 73.065 5.6 ;
        RECT 73.355 5.43 73.525 5.6 ;
        RECT 73.615 6.835 73.785 7.005 ;
        RECT 73.815 5.43 73.985 5.6 ;
        RECT 74.275 5.43 74.445 5.6 ;
        RECT 74.735 5.43 74.905 5.6 ;
        RECT 78.395 6.835 78.565 7.005 ;
        RECT 78.395 5.455 78.565 5.625 ;
        RECT 79.1 6.835 79.27 7.005 ;
        RECT 79.1 5.455 79.27 5.625 ;
        RECT 80.085 5.455 80.255 5.625 ;
        RECT 80.09 6.835 80.26 7.005 ;
        RECT 81.32 5.43 81.49 5.6 ;
        RECT 81.78 5.43 81.95 5.6 ;
        RECT 82.24 5.43 82.41 5.6 ;
        RECT 82.7 5.43 82.87 5.6 ;
        RECT 83.16 5.43 83.33 5.6 ;
        RECT 83.62 5.43 83.79 5.6 ;
        RECT 84.08 5.43 84.25 5.6 ;
        RECT 84.54 5.43 84.71 5.6 ;
        RECT 85 5.43 85.17 5.6 ;
        RECT 85.46 5.43 85.63 5.6 ;
        RECT 85.92 5.43 86.09 5.6 ;
        RECT 86.38 5.43 86.55 5.6 ;
        RECT 86.84 5.43 87.01 5.6 ;
        RECT 87.3 5.43 87.47 5.6 ;
        RECT 87.76 5.43 87.93 5.6 ;
        RECT 88.22 5.43 88.39 5.6 ;
        RECT 88.68 5.43 88.85 5.6 ;
        RECT 89.14 5.43 89.31 5.6 ;
        RECT 89.4 6.835 89.57 7.005 ;
        RECT 89.6 5.43 89.77 5.6 ;
        RECT 90.06 5.43 90.23 5.6 ;
        RECT 90.52 5.43 90.69 5.6 ;
        RECT 94.18 6.835 94.35 7.005 ;
        RECT 94.18 5.455 94.35 5.625 ;
        RECT 94.885 6.835 95.055 7.005 ;
        RECT 94.885 5.455 95.055 5.625 ;
        RECT 95.87 5.455 96.04 5.625 ;
        RECT 95.875 6.835 96.045 7.005 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 90.065 4.27 90.395 5 ;
        RECT 74.28 4.27 74.61 5 ;
        RECT 58.495 4.27 58.825 5 ;
        RECT 42.72 4.27 43.05 5 ;
        RECT 26.94 4.27 27.27 5 ;
      LAYER li1 ;
        RECT 0.005 0 96.775 1.6 ;
        RECT 95.79 0 95.96 2.225 ;
        RECT 94.805 0 94.975 2.225 ;
        RECT 92.06 0 92.23 2.225 ;
        RECT 81.175 0 91.005 2.885 ;
        RECT 89.305 0 89.475 3.38 ;
        RECT 87.345 0 87.515 3.38 ;
        RECT 84.905 0 85.075 3.38 ;
        RECT 83.945 0 84.115 3.38 ;
        RECT 83.425 0 83.595 3.38 ;
        RECT 82.465 0 82.635 3.38 ;
        RECT 81.505 0 81.675 3.38 ;
        RECT 80.005 0 80.175 2.225 ;
        RECT 79.02 0 79.19 2.225 ;
        RECT 76.275 0 76.445 2.225 ;
        RECT 65.39 0 75.22 2.885 ;
        RECT 73.52 0 73.69 3.38 ;
        RECT 71.56 0 71.73 3.38 ;
        RECT 69.12 0 69.29 3.38 ;
        RECT 68.16 0 68.33 3.38 ;
        RECT 67.64 0 67.81 3.38 ;
        RECT 66.68 0 66.85 3.38 ;
        RECT 65.72 0 65.89 3.38 ;
        RECT 64.22 0 64.39 2.225 ;
        RECT 63.235 0 63.405 2.225 ;
        RECT 60.49 0 60.66 2.225 ;
        RECT 49.605 0 59.435 2.885 ;
        RECT 57.735 0 57.905 3.38 ;
        RECT 55.775 0 55.945 3.38 ;
        RECT 53.335 0 53.505 3.38 ;
        RECT 52.375 0 52.545 3.38 ;
        RECT 51.855 0 52.025 3.38 ;
        RECT 50.895 0 51.065 3.38 ;
        RECT 49.935 0 50.105 3.38 ;
        RECT 48.445 0 48.615 2.225 ;
        RECT 47.46 0 47.63 2.225 ;
        RECT 44.715 0 44.885 2.225 ;
        RECT 33.83 0 43.66 2.885 ;
        RECT 41.96 0 42.13 3.38 ;
        RECT 40 0 40.17 3.38 ;
        RECT 37.56 0 37.73 3.38 ;
        RECT 36.6 0 36.77 3.38 ;
        RECT 36.08 0 36.25 3.38 ;
        RECT 35.12 0 35.29 3.38 ;
        RECT 34.16 0 34.33 3.38 ;
        RECT 32.665 0 32.835 2.225 ;
        RECT 31.68 0 31.85 2.225 ;
        RECT 28.935 0 29.105 2.225 ;
        RECT 18.05 0 27.88 2.885 ;
        RECT 26.18 0 26.35 3.38 ;
        RECT 24.22 0 24.39 3.38 ;
        RECT 21.78 0 21.95 3.38 ;
        RECT 20.82 0 20.99 3.38 ;
        RECT 20.3 0 20.47 3.38 ;
        RECT 19.34 0 19.51 3.38 ;
        RECT 18.38 0 18.55 3.38 ;
        RECT 0 10.86 96.775 12.46 ;
        RECT 95.795 10.235 95.965 12.46 ;
        RECT 94.805 10.235 94.975 12.46 ;
        RECT 92.06 10.235 92.23 12.46 ;
        RECT 87.28 10.235 87.45 12.46 ;
        RECT 80.01 10.235 80.18 12.46 ;
        RECT 79.02 10.235 79.19 12.46 ;
        RECT 76.275 10.235 76.445 12.46 ;
        RECT 71.495 10.235 71.665 12.46 ;
        RECT 64.225 10.235 64.395 12.46 ;
        RECT 63.235 10.235 63.405 12.46 ;
        RECT 60.49 10.235 60.66 12.46 ;
        RECT 55.71 10.235 55.88 12.46 ;
        RECT 48.45 10.235 48.62 12.46 ;
        RECT 47.46 10.235 47.63 12.46 ;
        RECT 44.715 10.235 44.885 12.46 ;
        RECT 39.935 10.235 40.105 12.46 ;
        RECT 32.67 10.235 32.84 12.46 ;
        RECT 31.68 10.235 31.85 12.46 ;
        RECT 28.935 10.235 29.105 12.46 ;
        RECT 24.155 10.235 24.325 12.46 ;
        RECT 15.28 10.235 15.45 12.46 ;
        RECT 90.075 3.87 90.435 4.645 ;
        RECT 90.025 3.87 90.435 4.17 ;
        RECT 88.06 3.87 88.475 4.225 ;
        RECT 88.295 8.365 88.465 10.315 ;
        RECT 88.235 10.145 88.405 10.595 ;
        RECT 88.235 7.305 88.405 8.535 ;
        RECT 74.29 3.87 74.65 4.645 ;
        RECT 74.24 3.87 74.65 4.17 ;
        RECT 72.275 3.87 72.69 4.225 ;
        RECT 72.51 8.365 72.68 10.315 ;
        RECT 72.45 10.145 72.62 10.595 ;
        RECT 72.45 7.305 72.62 8.535 ;
        RECT 58.505 3.87 58.865 4.645 ;
        RECT 58.455 3.87 58.865 4.17 ;
        RECT 56.49 3.87 56.905 4.225 ;
        RECT 56.725 8.365 56.895 10.315 ;
        RECT 56.665 10.145 56.835 10.595 ;
        RECT 56.665 7.305 56.835 8.535 ;
        RECT 42.73 3.87 43.09 4.645 ;
        RECT 42.68 3.87 43.09 4.17 ;
        RECT 40.715 3.87 41.13 4.225 ;
        RECT 40.95 8.365 41.12 10.315 ;
        RECT 40.89 10.145 41.06 10.595 ;
        RECT 40.89 7.305 41.06 8.535 ;
        RECT 26.95 3.87 27.31 4.645 ;
        RECT 26.9 3.87 27.31 4.17 ;
        RECT 24.935 3.87 25.35 4.225 ;
        RECT 25.17 8.365 25.34 10.315 ;
        RECT 25.11 10.145 25.28 10.595 ;
        RECT 25.11 7.305 25.28 8.535 ;
      LAYER met2 ;
        RECT 90.06 4.07 90.435 4.645 ;
        RECT 90.09 3.945 90.435 4.645 ;
        RECT 74.275 4.07 74.65 4.645 ;
        RECT 74.305 3.945 74.65 4.645 ;
        RECT 58.49 4.07 58.865 4.645 ;
        RECT 58.52 3.945 58.865 4.645 ;
        RECT 42.715 4.07 43.09 4.645 ;
        RECT 42.745 3.945 43.09 4.645 ;
        RECT 26.935 4.07 27.31 4.645 ;
        RECT 26.965 3.945 27.31 4.645 ;
      LAYER met1 ;
        RECT 0.005 0 96.775 1.6 ;
        RECT 81.175 0 91.005 2.885 ;
        RECT 81.175 0 90.835 3.035 ;
        RECT 90.615 0 90.8 4.33 ;
        RECT 89.93 4.165 90.8 4.33 ;
        RECT 90.025 4.145 90.8 4.33 ;
        RECT 90.075 4.075 90.435 4.745 ;
        RECT 90.09 4.07 90.435 4.745 ;
        RECT 90.025 4.075 90.435 4.72 ;
        RECT 89.215 4.26 90.435 4.57 ;
        RECT 88.27 4.235 89.285 4.26 ;
        RECT 89.175 4.26 90.435 4.565 ;
        RECT 89.11 4.26 90.435 4.51 ;
        RECT 88.27 4.215 89.135 4.26 ;
        RECT 89.075 4.26 90.435 4.475 ;
        RECT 88.915 4.26 90.435 4.425 ;
        RECT 88.27 4.195 89.02 4.26 ;
        RECT 88.9 4.26 90.435 4.38 ;
        RECT 88.79 4.26 90.435 4.375 ;
        RECT 88.27 4.165 88.895 4.26 ;
        RECT 88.27 4.13 88.805 4.26 ;
        RECT 88.675 4.26 90.435 4.345 ;
        RECT 88.27 4.075 88.7 4.26 ;
        RECT 88.27 4.05 88.675 4.26 ;
        RECT 88.61 4.26 90.8 4.31 ;
        RECT 88.47 4.26 90.8 4.29 ;
        RECT 88.27 4.035 88.515 4.26 ;
        RECT 88.27 4.02 88.5 4.26 ;
        RECT 65.39 0 75.22 2.885 ;
        RECT 65.39 0 75.05 3.035 ;
        RECT 74.83 0 75.015 4.33 ;
        RECT 74.145 4.165 75.015 4.33 ;
        RECT 74.24 4.145 75.015 4.33 ;
        RECT 74.29 4.075 74.65 4.745 ;
        RECT 74.305 4.07 74.65 4.745 ;
        RECT 74.24 4.075 74.65 4.72 ;
        RECT 73.43 4.26 74.65 4.57 ;
        RECT 72.485 4.235 73.5 4.26 ;
        RECT 73.39 4.26 74.65 4.565 ;
        RECT 73.325 4.26 74.65 4.51 ;
        RECT 72.485 4.215 73.35 4.26 ;
        RECT 73.29 4.26 74.65 4.475 ;
        RECT 73.13 4.26 74.65 4.425 ;
        RECT 72.485 4.195 73.235 4.26 ;
        RECT 73.115 4.26 74.65 4.38 ;
        RECT 73.005 4.26 74.65 4.375 ;
        RECT 72.485 4.165 73.11 4.26 ;
        RECT 72.485 4.13 73.02 4.26 ;
        RECT 72.89 4.26 74.65 4.345 ;
        RECT 72.485 4.075 72.915 4.26 ;
        RECT 72.485 4.05 72.89 4.26 ;
        RECT 72.825 4.26 75.015 4.31 ;
        RECT 72.685 4.26 75.015 4.29 ;
        RECT 72.485 4.035 72.73 4.26 ;
        RECT 72.485 4.02 72.715 4.26 ;
        RECT 49.605 0 59.435 2.885 ;
        RECT 49.605 0 59.265 3.035 ;
        RECT 59.045 0 59.23 4.33 ;
        RECT 58.36 4.165 59.23 4.33 ;
        RECT 58.455 4.145 59.23 4.33 ;
        RECT 58.505 4.075 58.865 4.745 ;
        RECT 58.52 4.07 58.865 4.745 ;
        RECT 58.455 4.075 58.865 4.72 ;
        RECT 57.645 4.26 58.865 4.57 ;
        RECT 56.7 4.235 57.715 4.26 ;
        RECT 57.605 4.26 58.865 4.565 ;
        RECT 57.54 4.26 58.865 4.51 ;
        RECT 56.7 4.215 57.565 4.26 ;
        RECT 57.505 4.26 58.865 4.475 ;
        RECT 57.345 4.26 58.865 4.425 ;
        RECT 56.7 4.195 57.45 4.26 ;
        RECT 57.33 4.26 58.865 4.38 ;
        RECT 57.22 4.26 58.865 4.375 ;
        RECT 56.7 4.165 57.325 4.26 ;
        RECT 56.7 4.13 57.235 4.26 ;
        RECT 57.105 4.26 58.865 4.345 ;
        RECT 56.7 4.075 57.13 4.26 ;
        RECT 56.7 4.05 57.105 4.26 ;
        RECT 57.04 4.26 59.23 4.31 ;
        RECT 56.9 4.26 59.23 4.29 ;
        RECT 56.7 4.035 56.945 4.26 ;
        RECT 56.7 4.02 56.93 4.26 ;
        RECT 33.83 0 43.66 2.885 ;
        RECT 33.83 0 43.49 3.035 ;
        RECT 43.27 0 43.455 4.33 ;
        RECT 42.585 4.165 43.455 4.33 ;
        RECT 42.68 4.145 43.455 4.33 ;
        RECT 42.73 4.075 43.09 4.745 ;
        RECT 42.745 4.07 43.09 4.745 ;
        RECT 42.68 4.075 43.09 4.72 ;
        RECT 41.87 4.26 43.09 4.57 ;
        RECT 40.925 4.235 41.94 4.26 ;
        RECT 41.83 4.26 43.09 4.565 ;
        RECT 41.765 4.26 43.09 4.51 ;
        RECT 40.925 4.215 41.79 4.26 ;
        RECT 41.73 4.26 43.09 4.475 ;
        RECT 41.57 4.26 43.09 4.425 ;
        RECT 40.925 4.195 41.675 4.26 ;
        RECT 41.555 4.26 43.09 4.38 ;
        RECT 41.445 4.26 43.09 4.375 ;
        RECT 40.925 4.165 41.55 4.26 ;
        RECT 40.925 4.13 41.46 4.26 ;
        RECT 41.33 4.26 43.09 4.345 ;
        RECT 40.925 4.075 41.355 4.26 ;
        RECT 40.925 4.05 41.33 4.26 ;
        RECT 41.265 4.26 43.455 4.31 ;
        RECT 41.125 4.26 43.455 4.29 ;
        RECT 40.925 4.035 41.17 4.26 ;
        RECT 40.925 4.02 41.155 4.26 ;
        RECT 18.05 0 27.88 2.885 ;
        RECT 18.05 0 27.71 3.035 ;
        RECT 27.49 0 27.675 4.33 ;
        RECT 26.805 4.165 27.675 4.33 ;
        RECT 26.9 4.145 27.675 4.33 ;
        RECT 26.95 4.075 27.31 4.745 ;
        RECT 26.965 4.07 27.31 4.745 ;
        RECT 26.9 4.075 27.31 4.72 ;
        RECT 26.09 4.26 27.31 4.57 ;
        RECT 25.145 4.235 26.16 4.26 ;
        RECT 26.05 4.26 27.31 4.565 ;
        RECT 25.985 4.26 27.31 4.51 ;
        RECT 25.145 4.215 26.01 4.26 ;
        RECT 25.95 4.26 27.31 4.475 ;
        RECT 25.79 4.26 27.31 4.425 ;
        RECT 25.145 4.195 25.895 4.26 ;
        RECT 25.775 4.26 27.31 4.38 ;
        RECT 25.665 4.26 27.31 4.375 ;
        RECT 25.145 4.165 25.77 4.26 ;
        RECT 25.145 4.13 25.68 4.26 ;
        RECT 25.55 4.26 27.31 4.345 ;
        RECT 25.145 4.075 25.575 4.26 ;
        RECT 25.145 4.05 25.55 4.26 ;
        RECT 25.485 4.26 27.675 4.31 ;
        RECT 25.345 4.26 27.675 4.29 ;
        RECT 25.145 4.035 25.39 4.26 ;
        RECT 25.145 4.02 25.375 4.26 ;
        RECT 0 10.86 96.775 12.46 ;
        RECT 88.235 8.575 88.525 8.805 ;
        RECT 88.06 8.605 88.525 8.775 ;
        RECT 87.86 8.6 88.23 8.77 ;
        RECT 87.86 8.6 88.03 12.46 ;
        RECT 72.45 8.575 72.74 8.805 ;
        RECT 72.275 8.605 72.74 8.775 ;
        RECT 72.075 8.6 72.445 8.77 ;
        RECT 72.075 8.6 72.245 12.46 ;
        RECT 56.665 8.575 56.955 8.805 ;
        RECT 56.49 8.605 56.955 8.775 ;
        RECT 56.29 8.6 56.66 8.77 ;
        RECT 56.29 8.6 56.46 12.46 ;
        RECT 40.89 8.575 41.18 8.805 ;
        RECT 40.715 8.605 41.18 8.775 ;
        RECT 40.515 8.6 40.885 8.77 ;
        RECT 40.515 8.6 40.685 12.46 ;
        RECT 25.11 8.575 25.4 8.805 ;
        RECT 24.935 8.605 25.4 8.775 ;
        RECT 24.735 8.6 25.105 8.77 ;
        RECT 24.735 8.6 24.905 12.46 ;
      LAYER via1 ;
        RECT 27.02 4.155 27.17 4.305 ;
        RECT 42.8 4.155 42.95 4.305 ;
        RECT 58.575 4.155 58.725 4.305 ;
        RECT 74.36 4.155 74.51 4.305 ;
        RECT 90.145 4.155 90.295 4.305 ;
      LAYER via2 ;
        RECT 27.005 4.335 27.205 4.535 ;
        RECT 42.785 4.335 42.985 4.535 ;
        RECT 58.56 4.335 58.76 4.535 ;
        RECT 74.345 4.335 74.545 4.535 ;
        RECT 90.13 4.335 90.33 4.535 ;
      LAYER mcon ;
        RECT 15.36 10.895 15.53 11.065 ;
        RECT 16.04 10.895 16.21 11.065 ;
        RECT 16.72 10.895 16.89 11.065 ;
        RECT 17.4 10.895 17.57 11.065 ;
        RECT 18.195 2.71 18.365 2.88 ;
        RECT 18.655 2.71 18.825 2.88 ;
        RECT 19.115 2.71 19.285 2.88 ;
        RECT 19.575 2.71 19.745 2.88 ;
        RECT 20.035 2.71 20.205 2.88 ;
        RECT 20.495 2.71 20.665 2.88 ;
        RECT 20.955 2.71 21.125 2.88 ;
        RECT 21.415 2.71 21.585 2.88 ;
        RECT 21.875 2.71 22.045 2.88 ;
        RECT 22.335 2.71 22.505 2.88 ;
        RECT 22.795 2.71 22.965 2.88 ;
        RECT 23.255 2.71 23.425 2.88 ;
        RECT 23.715 2.71 23.885 2.88 ;
        RECT 24.175 2.71 24.345 2.88 ;
        RECT 24.235 10.895 24.405 11.065 ;
        RECT 24.635 2.71 24.805 2.88 ;
        RECT 24.915 10.895 25.085 11.065 ;
        RECT 25.095 2.71 25.265 2.88 ;
        RECT 25.17 8.605 25.34 8.775 ;
        RECT 25.18 4.055 25.35 4.225 ;
        RECT 25.555 2.71 25.725 2.88 ;
        RECT 25.595 10.895 25.765 11.065 ;
        RECT 26.015 2.71 26.185 2.88 ;
        RECT 26.275 10.895 26.445 11.065 ;
        RECT 26.475 2.71 26.645 2.88 ;
        RECT 26.935 2.71 27.105 2.88 ;
        RECT 27.025 4.17 27.195 4.34 ;
        RECT 27.395 2.71 27.565 2.88 ;
        RECT 29.015 10.895 29.185 11.065 ;
        RECT 29.015 1.395 29.185 1.565 ;
        RECT 29.695 10.895 29.865 11.065 ;
        RECT 29.695 1.395 29.865 1.565 ;
        RECT 30.375 10.895 30.545 11.065 ;
        RECT 30.375 1.395 30.545 1.565 ;
        RECT 31.055 10.895 31.225 11.065 ;
        RECT 31.055 1.395 31.225 1.565 ;
        RECT 31.76 10.895 31.93 11.065 ;
        RECT 31.76 1.395 31.93 1.565 ;
        RECT 32.745 1.395 32.915 1.565 ;
        RECT 32.75 10.895 32.92 11.065 ;
        RECT 33.975 2.71 34.145 2.88 ;
        RECT 34.435 2.71 34.605 2.88 ;
        RECT 34.895 2.71 35.065 2.88 ;
        RECT 35.355 2.71 35.525 2.88 ;
        RECT 35.815 2.71 35.985 2.88 ;
        RECT 36.275 2.71 36.445 2.88 ;
        RECT 36.735 2.71 36.905 2.88 ;
        RECT 37.195 2.71 37.365 2.88 ;
        RECT 37.655 2.71 37.825 2.88 ;
        RECT 38.115 2.71 38.285 2.88 ;
        RECT 38.575 2.71 38.745 2.88 ;
        RECT 39.035 2.71 39.205 2.88 ;
        RECT 39.495 2.71 39.665 2.88 ;
        RECT 39.955 2.71 40.125 2.88 ;
        RECT 40.015 10.895 40.185 11.065 ;
        RECT 40.415 2.71 40.585 2.88 ;
        RECT 40.695 10.895 40.865 11.065 ;
        RECT 40.875 2.71 41.045 2.88 ;
        RECT 40.95 8.605 41.12 8.775 ;
        RECT 40.96 4.055 41.13 4.225 ;
        RECT 41.335 2.71 41.505 2.88 ;
        RECT 41.375 10.895 41.545 11.065 ;
        RECT 41.795 2.71 41.965 2.88 ;
        RECT 42.055 10.895 42.225 11.065 ;
        RECT 42.255 2.71 42.425 2.88 ;
        RECT 42.715 2.71 42.885 2.88 ;
        RECT 42.805 4.17 42.975 4.34 ;
        RECT 43.175 2.71 43.345 2.88 ;
        RECT 44.795 10.895 44.965 11.065 ;
        RECT 44.795 1.395 44.965 1.565 ;
        RECT 45.475 10.895 45.645 11.065 ;
        RECT 45.475 1.395 45.645 1.565 ;
        RECT 46.155 10.895 46.325 11.065 ;
        RECT 46.155 1.395 46.325 1.565 ;
        RECT 46.835 10.895 47.005 11.065 ;
        RECT 46.835 1.395 47.005 1.565 ;
        RECT 47.54 10.895 47.71 11.065 ;
        RECT 47.54 1.395 47.71 1.565 ;
        RECT 48.525 1.395 48.695 1.565 ;
        RECT 48.53 10.895 48.7 11.065 ;
        RECT 49.75 2.71 49.92 2.88 ;
        RECT 50.21 2.71 50.38 2.88 ;
        RECT 50.67 2.71 50.84 2.88 ;
        RECT 51.13 2.71 51.3 2.88 ;
        RECT 51.59 2.71 51.76 2.88 ;
        RECT 52.05 2.71 52.22 2.88 ;
        RECT 52.51 2.71 52.68 2.88 ;
        RECT 52.97 2.71 53.14 2.88 ;
        RECT 53.43 2.71 53.6 2.88 ;
        RECT 53.89 2.71 54.06 2.88 ;
        RECT 54.35 2.71 54.52 2.88 ;
        RECT 54.81 2.71 54.98 2.88 ;
        RECT 55.27 2.71 55.44 2.88 ;
        RECT 55.73 2.71 55.9 2.88 ;
        RECT 55.79 10.895 55.96 11.065 ;
        RECT 56.19 2.71 56.36 2.88 ;
        RECT 56.47 10.895 56.64 11.065 ;
        RECT 56.65 2.71 56.82 2.88 ;
        RECT 56.725 8.605 56.895 8.775 ;
        RECT 56.735 4.055 56.905 4.225 ;
        RECT 57.11 2.71 57.28 2.88 ;
        RECT 57.15 10.895 57.32 11.065 ;
        RECT 57.57 2.71 57.74 2.88 ;
        RECT 57.83 10.895 58 11.065 ;
        RECT 58.03 2.71 58.2 2.88 ;
        RECT 58.49 2.71 58.66 2.88 ;
        RECT 58.58 4.17 58.75 4.34 ;
        RECT 58.95 2.71 59.12 2.88 ;
        RECT 60.57 10.895 60.74 11.065 ;
        RECT 60.57 1.395 60.74 1.565 ;
        RECT 61.25 10.895 61.42 11.065 ;
        RECT 61.25 1.395 61.42 1.565 ;
        RECT 61.93 10.895 62.1 11.065 ;
        RECT 61.93 1.395 62.1 1.565 ;
        RECT 62.61 10.895 62.78 11.065 ;
        RECT 62.61 1.395 62.78 1.565 ;
        RECT 63.315 10.895 63.485 11.065 ;
        RECT 63.315 1.395 63.485 1.565 ;
        RECT 64.3 1.395 64.47 1.565 ;
        RECT 64.305 10.895 64.475 11.065 ;
        RECT 65.535 2.71 65.705 2.88 ;
        RECT 65.995 2.71 66.165 2.88 ;
        RECT 66.455 2.71 66.625 2.88 ;
        RECT 66.915 2.71 67.085 2.88 ;
        RECT 67.375 2.71 67.545 2.88 ;
        RECT 67.835 2.71 68.005 2.88 ;
        RECT 68.295 2.71 68.465 2.88 ;
        RECT 68.755 2.71 68.925 2.88 ;
        RECT 69.215 2.71 69.385 2.88 ;
        RECT 69.675 2.71 69.845 2.88 ;
        RECT 70.135 2.71 70.305 2.88 ;
        RECT 70.595 2.71 70.765 2.88 ;
        RECT 71.055 2.71 71.225 2.88 ;
        RECT 71.515 2.71 71.685 2.88 ;
        RECT 71.575 10.895 71.745 11.065 ;
        RECT 71.975 2.71 72.145 2.88 ;
        RECT 72.255 10.895 72.425 11.065 ;
        RECT 72.435 2.71 72.605 2.88 ;
        RECT 72.51 8.605 72.68 8.775 ;
        RECT 72.52 4.055 72.69 4.225 ;
        RECT 72.895 2.71 73.065 2.88 ;
        RECT 72.935 10.895 73.105 11.065 ;
        RECT 73.355 2.71 73.525 2.88 ;
        RECT 73.615 10.895 73.785 11.065 ;
        RECT 73.815 2.71 73.985 2.88 ;
        RECT 74.275 2.71 74.445 2.88 ;
        RECT 74.365 4.17 74.535 4.34 ;
        RECT 74.735 2.71 74.905 2.88 ;
        RECT 76.355 10.895 76.525 11.065 ;
        RECT 76.355 1.395 76.525 1.565 ;
        RECT 77.035 10.895 77.205 11.065 ;
        RECT 77.035 1.395 77.205 1.565 ;
        RECT 77.715 10.895 77.885 11.065 ;
        RECT 77.715 1.395 77.885 1.565 ;
        RECT 78.395 10.895 78.565 11.065 ;
        RECT 78.395 1.395 78.565 1.565 ;
        RECT 79.1 10.895 79.27 11.065 ;
        RECT 79.1 1.395 79.27 1.565 ;
        RECT 80.085 1.395 80.255 1.565 ;
        RECT 80.09 10.895 80.26 11.065 ;
        RECT 81.32 2.71 81.49 2.88 ;
        RECT 81.78 2.71 81.95 2.88 ;
        RECT 82.24 2.71 82.41 2.88 ;
        RECT 82.7 2.71 82.87 2.88 ;
        RECT 83.16 2.71 83.33 2.88 ;
        RECT 83.62 2.71 83.79 2.88 ;
        RECT 84.08 2.71 84.25 2.88 ;
        RECT 84.54 2.71 84.71 2.88 ;
        RECT 85 2.71 85.17 2.88 ;
        RECT 85.46 2.71 85.63 2.88 ;
        RECT 85.92 2.71 86.09 2.88 ;
        RECT 86.38 2.71 86.55 2.88 ;
        RECT 86.84 2.71 87.01 2.88 ;
        RECT 87.3 2.71 87.47 2.88 ;
        RECT 87.36 10.895 87.53 11.065 ;
        RECT 87.76 2.71 87.93 2.88 ;
        RECT 88.04 10.895 88.21 11.065 ;
        RECT 88.22 2.71 88.39 2.88 ;
        RECT 88.295 8.605 88.465 8.775 ;
        RECT 88.305 4.055 88.475 4.225 ;
        RECT 88.68 2.71 88.85 2.88 ;
        RECT 88.72 10.895 88.89 11.065 ;
        RECT 89.14 2.71 89.31 2.88 ;
        RECT 89.4 10.895 89.57 11.065 ;
        RECT 89.6 2.71 89.77 2.88 ;
        RECT 90.06 2.71 90.23 2.88 ;
        RECT 90.15 4.17 90.32 4.34 ;
        RECT 90.52 2.71 90.69 2.88 ;
        RECT 92.14 10.895 92.31 11.065 ;
        RECT 92.14 1.395 92.31 1.565 ;
        RECT 92.82 10.895 92.99 11.065 ;
        RECT 92.82 1.395 92.99 1.565 ;
        RECT 93.5 10.895 93.67 11.065 ;
        RECT 93.5 1.395 93.67 1.565 ;
        RECT 94.18 10.895 94.35 11.065 ;
        RECT 94.18 1.395 94.35 1.565 ;
        RECT 94.885 10.895 95.055 11.065 ;
        RECT 94.885 1.395 95.055 1.565 ;
        RECT 95.87 1.395 96.04 1.565 ;
        RECT 95.875 10.895 96.045 11.065 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 88.565 9.325 88.935 9.695 ;
      RECT 88.605 9.005 88.935 9.695 ;
      RECT 88.605 9.005 91.395 9.31 ;
      RECT 91.09 4.145 91.395 9.31 ;
      RECT 91.055 4.145 91.425 4.515 ;
      RECT 86.425 3.145 86.755 4.04 ;
      RECT 85.545 3.31 85.875 4.04 ;
      RECT 86.42 3.145 86.79 3.945 ;
      RECT 89.585 3.145 89.915 3.875 ;
      RECT 89.545 3.03 89.725 3.68 ;
      RECT 85.555 3.145 89.915 3.515 ;
      RECT 86.045 4.83 86.375 5.16 ;
      RECT 84.84 4.845 86.375 5.145 ;
      RECT 84.84 3.725 85.14 5.145 ;
      RECT 84.585 3.71 84.915 4.04 ;
      RECT 72.78 9.325 73.15 9.695 ;
      RECT 72.82 9.005 73.15 9.695 ;
      RECT 72.82 9.005 75.61 9.31 ;
      RECT 75.305 4.145 75.61 9.31 ;
      RECT 75.27 4.145 75.64 4.515 ;
      RECT 70.64 3.145 70.97 4.04 ;
      RECT 69.76 3.31 70.09 4.04 ;
      RECT 70.635 3.145 71.005 3.945 ;
      RECT 73.8 3.145 74.13 3.875 ;
      RECT 73.76 3.03 73.94 3.68 ;
      RECT 69.77 3.145 74.13 3.515 ;
      RECT 70.26 4.83 70.59 5.16 ;
      RECT 69.055 4.845 70.59 5.145 ;
      RECT 69.055 3.725 69.355 5.145 ;
      RECT 68.8 3.71 69.13 4.04 ;
      RECT 56.995 9.325 57.365 9.695 ;
      RECT 57.035 9.005 57.365 9.695 ;
      RECT 57.035 9.005 59.825 9.31 ;
      RECT 59.52 4.145 59.825 9.31 ;
      RECT 59.485 4.145 59.855 4.515 ;
      RECT 54.855 3.145 55.185 4.04 ;
      RECT 53.975 3.31 54.305 4.04 ;
      RECT 54.85 3.145 55.22 3.945 ;
      RECT 58.015 3.145 58.345 3.875 ;
      RECT 57.975 3.03 58.155 3.68 ;
      RECT 53.985 3.145 58.345 3.515 ;
      RECT 54.475 4.83 54.805 5.16 ;
      RECT 53.27 4.845 54.805 5.145 ;
      RECT 53.27 3.725 53.57 5.145 ;
      RECT 53.015 3.71 53.345 4.04 ;
      RECT 41.22 9.325 41.59 9.695 ;
      RECT 41.26 9.005 41.59 9.695 ;
      RECT 41.26 9.005 44.05 9.31 ;
      RECT 43.745 4.145 44.05 9.31 ;
      RECT 43.71 4.145 44.08 4.515 ;
      RECT 39.08 3.145 39.41 4.04 ;
      RECT 38.2 3.31 38.53 4.04 ;
      RECT 39.075 3.145 39.445 3.945 ;
      RECT 42.24 3.145 42.57 3.875 ;
      RECT 42.2 3.03 42.38 3.68 ;
      RECT 38.21 3.145 42.57 3.515 ;
      RECT 38.7 4.83 39.03 5.16 ;
      RECT 37.495 4.845 39.03 5.145 ;
      RECT 37.495 3.725 37.795 5.145 ;
      RECT 37.24 3.71 37.57 4.04 ;
      RECT 25.44 9.325 25.81 9.695 ;
      RECT 25.48 9.005 25.81 9.695 ;
      RECT 25.48 9.005 28.27 9.31 ;
      RECT 27.965 4.145 28.27 9.31 ;
      RECT 27.93 4.145 28.3 4.515 ;
      RECT 23.3 3.145 23.63 4.04 ;
      RECT 22.42 3.31 22.75 4.04 ;
      RECT 23.295 3.145 23.665 3.945 ;
      RECT 26.46 3.145 26.79 3.875 ;
      RECT 26.42 3.03 26.6 3.68 ;
      RECT 22.43 3.145 26.79 3.515 ;
      RECT 22.92 4.83 23.25 5.16 ;
      RECT 21.715 4.845 23.25 5.145 ;
      RECT 21.715 3.725 22.015 5.145 ;
      RECT 21.46 3.71 21.79 4.04 ;
      RECT 96.14 7.215 96.49 12.46 ;
      RECT 87.985 3.87 88.315 4.6 ;
      RECT 83.865 3.71 84.195 4.44 ;
      RECT 82.865 3.15 83.195 3.88 ;
      RECT 81.425 3.87 81.755 4.6 ;
      RECT 80.355 7.215 80.705 12.46 ;
      RECT 72.2 3.87 72.53 4.6 ;
      RECT 68.08 3.71 68.41 4.44 ;
      RECT 67.08 3.15 67.41 3.88 ;
      RECT 65.64 3.87 65.97 4.6 ;
      RECT 64.57 7.215 64.92 12.46 ;
      RECT 56.415 3.87 56.745 4.6 ;
      RECT 52.295 3.71 52.625 4.44 ;
      RECT 51.295 3.15 51.625 3.88 ;
      RECT 49.855 3.87 50.185 4.6 ;
      RECT 48.795 7.215 49.145 12.46 ;
      RECT 40.64 3.87 40.97 4.6 ;
      RECT 36.52 3.71 36.85 4.44 ;
      RECT 35.52 3.15 35.85 3.88 ;
      RECT 34.08 3.87 34.41 4.6 ;
      RECT 33.015 7.215 33.365 12.46 ;
      RECT 24.86 3.87 25.19 4.6 ;
      RECT 20.74 3.71 21.07 4.44 ;
      RECT 19.74 3.15 20.07 3.88 ;
      RECT 18.3 3.87 18.63 4.6 ;
    LAYER via2 ;
      RECT 96.225 7.3 96.425 7.5 ;
      RECT 91.14 4.23 91.34 4.43 ;
      RECT 89.65 3.61 89.85 3.81 ;
      RECT 88.65 9.41 88.85 9.61 ;
      RECT 88.05 4.335 88.25 4.535 ;
      RECT 86.49 3.775 86.69 3.975 ;
      RECT 86.11 4.895 86.31 5.095 ;
      RECT 85.61 3.775 85.81 3.975 ;
      RECT 84.65 3.775 84.85 3.975 ;
      RECT 83.93 3.775 84.13 3.975 ;
      RECT 82.93 3.215 83.13 3.415 ;
      RECT 81.49 4.335 81.69 4.535 ;
      RECT 80.44 7.3 80.64 7.5 ;
      RECT 75.355 4.23 75.555 4.43 ;
      RECT 73.865 3.61 74.065 3.81 ;
      RECT 72.865 9.41 73.065 9.61 ;
      RECT 72.265 4.335 72.465 4.535 ;
      RECT 70.705 3.775 70.905 3.975 ;
      RECT 70.325 4.895 70.525 5.095 ;
      RECT 69.825 3.775 70.025 3.975 ;
      RECT 68.865 3.775 69.065 3.975 ;
      RECT 68.145 3.775 68.345 3.975 ;
      RECT 67.145 3.215 67.345 3.415 ;
      RECT 65.705 4.335 65.905 4.535 ;
      RECT 64.655 7.3 64.855 7.5 ;
      RECT 59.57 4.23 59.77 4.43 ;
      RECT 58.08 3.61 58.28 3.81 ;
      RECT 57.08 9.41 57.28 9.61 ;
      RECT 56.48 4.335 56.68 4.535 ;
      RECT 54.92 3.775 55.12 3.975 ;
      RECT 54.54 4.895 54.74 5.095 ;
      RECT 54.04 3.775 54.24 3.975 ;
      RECT 53.08 3.775 53.28 3.975 ;
      RECT 52.36 3.775 52.56 3.975 ;
      RECT 51.36 3.215 51.56 3.415 ;
      RECT 49.92 4.335 50.12 4.535 ;
      RECT 48.88 7.3 49.08 7.5 ;
      RECT 43.795 4.23 43.995 4.43 ;
      RECT 42.305 3.61 42.505 3.81 ;
      RECT 41.305 9.41 41.505 9.61 ;
      RECT 40.705 4.335 40.905 4.535 ;
      RECT 39.145 3.775 39.345 3.975 ;
      RECT 38.765 4.895 38.965 5.095 ;
      RECT 38.265 3.775 38.465 3.975 ;
      RECT 37.305 3.775 37.505 3.975 ;
      RECT 36.585 3.775 36.785 3.975 ;
      RECT 35.585 3.215 35.785 3.415 ;
      RECT 34.145 4.335 34.345 4.535 ;
      RECT 33.1 7.3 33.3 7.5 ;
      RECT 28.015 4.23 28.215 4.43 ;
      RECT 26.525 3.61 26.725 3.81 ;
      RECT 25.525 9.41 25.725 9.61 ;
      RECT 24.925 4.335 25.125 4.535 ;
      RECT 23.365 3.775 23.565 3.975 ;
      RECT 22.985 4.895 23.185 5.095 ;
      RECT 22.485 3.775 22.685 3.975 ;
      RECT 21.525 3.775 21.725 3.975 ;
      RECT 20.805 3.775 21.005 3.975 ;
      RECT 19.805 3.215 20.005 3.415 ;
      RECT 18.365 4.335 18.565 4.535 ;
    LAYER met2 ;
      RECT 16.23 10.685 65.755 10.855 ;
      RECT 96.23 9.55 96.4 10.845 ;
      RECT 65.755 10.675 96.4 10.845 ;
      RECT 16.23 8.54 16.4 10.855 ;
      RECT 96.2 9.55 96.55 9.9 ;
      RECT 16.17 8.54 16.46 8.89 ;
      RECT 93.04 8.505 93.36 8.83 ;
      RECT 93.07 7.98 93.24 8.83 ;
      RECT 93.07 7.98 93.245 8.33 ;
      RECT 93.07 7.98 94.045 8.155 ;
      RECT 93.87 3.26 94.045 8.155 ;
      RECT 93.815 3.26 94.165 3.61 ;
      RECT 93.84 8.94 94.165 9.265 ;
      RECT 92.725 9.03 94.165 9.2 ;
      RECT 92.725 3.69 92.885 9.2 ;
      RECT 93.04 3.66 93.36 3.98 ;
      RECT 92.725 3.69 93.36 3.86 ;
      RECT 81.45 4.295 81.73 4.575 ;
      RECT 81.42 4.295 81.73 4.56 ;
      RECT 81.415 4.295 81.73 4.558 ;
      RECT 81.41 2.625 81.58 4.552 ;
      RECT 81.405 4.262 81.675 4.545 ;
      RECT 81.4 4.295 81.73 4.538 ;
      RECT 81.37 4.265 81.675 4.525 ;
      RECT 81.37 4.292 81.695 4.525 ;
      RECT 81.37 4.282 81.69 4.525 ;
      RECT 81.37 4.267 81.685 4.525 ;
      RECT 81.41 4.257 81.675 4.552 ;
      RECT 81.41 4.252 81.665 4.552 ;
      RECT 81.41 4.251 81.65 4.552 ;
      RECT 91.38 2.635 91.73 2.985 ;
      RECT 91.375 2.635 91.73 2.89 ;
      RECT 81.41 2.625 91.62 2.795 ;
      RECT 91.055 4.145 91.425 4.515 ;
      RECT 91.14 3.53 91.31 4.515 ;
      RECT 87.16 3.75 87.395 4.01 ;
      RECT 90.305 3.53 90.47 3.79 ;
      RECT 90.21 3.52 90.225 3.79 ;
      RECT 90.305 3.53 91.31 3.71 ;
      RECT 88.81 3.09 88.85 3.23 ;
      RECT 90.225 3.525 90.305 3.79 ;
      RECT 90.17 3.52 90.21 3.756 ;
      RECT 90.156 3.52 90.17 3.756 ;
      RECT 90.07 3.525 90.156 3.758 ;
      RECT 90.025 3.532 90.07 3.76 ;
      RECT 89.995 3.532 90.025 3.762 ;
      RECT 89.97 3.527 89.995 3.764 ;
      RECT 89.94 3.523 89.97 3.773 ;
      RECT 89.93 3.52 89.94 3.785 ;
      RECT 89.925 3.52 89.93 3.793 ;
      RECT 89.92 3.52 89.925 3.798 ;
      RECT 89.91 3.519 89.92 3.808 ;
      RECT 89.905 3.518 89.91 3.818 ;
      RECT 89.89 3.517 89.905 3.823 ;
      RECT 89.862 3.514 89.89 3.85 ;
      RECT 89.776 3.506 89.862 3.85 ;
      RECT 89.69 3.495 89.776 3.85 ;
      RECT 89.65 3.48 89.69 3.85 ;
      RECT 89.61 3.454 89.65 3.85 ;
      RECT 89.605 3.436 89.61 3.662 ;
      RECT 89.595 3.432 89.605 3.652 ;
      RECT 89.58 3.422 89.595 3.639 ;
      RECT 89.56 3.406 89.58 3.624 ;
      RECT 89.545 3.391 89.56 3.609 ;
      RECT 89.535 3.38 89.545 3.599 ;
      RECT 89.51 3.364 89.535 3.588 ;
      RECT 89.505 3.351 89.51 3.578 ;
      RECT 89.5 3.347 89.505 3.573 ;
      RECT 89.445 3.333 89.5 3.551 ;
      RECT 89.406 3.314 89.445 3.515 ;
      RECT 89.32 3.288 89.406 3.468 ;
      RECT 89.316 3.27 89.32 3.434 ;
      RECT 89.23 3.251 89.316 3.412 ;
      RECT 89.225 3.233 89.23 3.39 ;
      RECT 89.22 3.231 89.225 3.388 ;
      RECT 89.21 3.23 89.22 3.383 ;
      RECT 89.15 3.217 89.21 3.369 ;
      RECT 89.105 3.195 89.15 3.348 ;
      RECT 89.045 3.172 89.105 3.327 ;
      RECT 88.981 3.147 89.045 3.302 ;
      RECT 88.895 3.117 88.981 3.271 ;
      RECT 88.88 3.097 88.895 3.25 ;
      RECT 88.85 3.092 88.88 3.241 ;
      RECT 88.797 3.09 88.81 3.23 ;
      RECT 88.711 3.09 88.797 3.232 ;
      RECT 88.625 3.09 88.711 3.234 ;
      RECT 88.605 3.09 88.625 3.238 ;
      RECT 88.56 3.092 88.605 3.249 ;
      RECT 88.52 3.102 88.56 3.265 ;
      RECT 88.516 3.111 88.52 3.273 ;
      RECT 88.43 3.131 88.516 3.289 ;
      RECT 88.42 3.15 88.43 3.307 ;
      RECT 88.415 3.152 88.42 3.31 ;
      RECT 88.405 3.156 88.415 3.313 ;
      RECT 88.385 3.161 88.405 3.323 ;
      RECT 88.355 3.171 88.385 3.343 ;
      RECT 88.35 3.178 88.355 3.357 ;
      RECT 88.34 3.182 88.35 3.364 ;
      RECT 88.325 3.19 88.34 3.375 ;
      RECT 88.315 3.2 88.325 3.386 ;
      RECT 88.305 3.207 88.315 3.394 ;
      RECT 88.28 3.22 88.305 3.409 ;
      RECT 88.216 3.256 88.28 3.448 ;
      RECT 88.13 3.319 88.216 3.512 ;
      RECT 88.095 3.37 88.13 3.565 ;
      RECT 88.09 3.387 88.095 3.582 ;
      RECT 88.075 3.396 88.09 3.589 ;
      RECT 88.055 3.411 88.075 3.603 ;
      RECT 88.05 3.422 88.055 3.613 ;
      RECT 88.03 3.435 88.05 3.623 ;
      RECT 88.025 3.445 88.03 3.633 ;
      RECT 88.01 3.45 88.025 3.642 ;
      RECT 88 3.46 88.01 3.653 ;
      RECT 87.97 3.477 88 3.67 ;
      RECT 87.96 3.495 87.97 3.688 ;
      RECT 87.945 3.506 87.96 3.699 ;
      RECT 87.905 3.53 87.945 3.715 ;
      RECT 87.87 3.564 87.905 3.732 ;
      RECT 87.84 3.587 87.87 3.744 ;
      RECT 87.825 3.597 87.84 3.753 ;
      RECT 87.785 3.607 87.825 3.764 ;
      RECT 87.765 3.618 87.785 3.776 ;
      RECT 87.76 3.622 87.765 3.783 ;
      RECT 87.745 3.626 87.76 3.788 ;
      RECT 87.735 3.631 87.745 3.793 ;
      RECT 87.73 3.634 87.735 3.796 ;
      RECT 87.7 3.64 87.73 3.803 ;
      RECT 87.665 3.65 87.7 3.817 ;
      RECT 87.605 3.665 87.665 3.837 ;
      RECT 87.55 3.685 87.605 3.861 ;
      RECT 87.521 3.7 87.55 3.879 ;
      RECT 87.435 3.72 87.521 3.904 ;
      RECT 87.43 3.735 87.435 3.924 ;
      RECT 87.42 3.738 87.43 3.925 ;
      RECT 87.395 3.745 87.42 4.01 ;
      RECT 80.39 8.945 80.74 9.295 ;
      RECT 89.215 8.9 89.565 9.25 ;
      RECT 80.39 8.975 89.565 9.175 ;
      RECT 87.81 4.98 87.82 5.17 ;
      RECT 86.07 4.855 86.35 5.135 ;
      RECT 89.115 3.795 89.12 4.28 ;
      RECT 89.01 3.795 89.07 4.055 ;
      RECT 89.335 4.765 89.34 4.84 ;
      RECT 89.325 4.632 89.335 4.875 ;
      RECT 89.315 4.467 89.325 4.896 ;
      RECT 89.31 4.337 89.315 4.912 ;
      RECT 89.3 4.227 89.31 4.928 ;
      RECT 89.295 4.126 89.3 4.945 ;
      RECT 89.29 4.108 89.295 4.955 ;
      RECT 89.285 4.09 89.29 4.965 ;
      RECT 89.275 4.065 89.285 4.98 ;
      RECT 89.27 4.045 89.275 4.995 ;
      RECT 89.25 3.795 89.27 5.02 ;
      RECT 89.235 3.795 89.25 5.053 ;
      RECT 89.205 3.795 89.235 5.075 ;
      RECT 89.185 3.795 89.205 5.089 ;
      RECT 89.165 3.795 89.185 4.605 ;
      RECT 89.18 4.672 89.185 5.094 ;
      RECT 89.175 4.702 89.18 5.096 ;
      RECT 89.17 4.715 89.175 5.099 ;
      RECT 89.165 4.725 89.17 5.103 ;
      RECT 89.16 3.795 89.165 4.523 ;
      RECT 89.16 4.735 89.165 5.105 ;
      RECT 89.155 3.795 89.16 4.5 ;
      RECT 89.145 4.757 89.16 5.105 ;
      RECT 89.14 3.795 89.155 4.445 ;
      RECT 89.135 4.782 89.145 5.105 ;
      RECT 89.135 3.795 89.14 4.39 ;
      RECT 89.125 3.795 89.135 4.338 ;
      RECT 89.13 4.795 89.135 5.106 ;
      RECT 89.125 4.807 89.13 5.107 ;
      RECT 89.12 3.795 89.125 4.298 ;
      RECT 89.12 4.82 89.125 5.108 ;
      RECT 89.105 4.835 89.12 5.109 ;
      RECT 89.11 3.795 89.115 4.26 ;
      RECT 89.105 3.795 89.11 4.225 ;
      RECT 89.1 3.795 89.105 4.2 ;
      RECT 89.095 4.862 89.105 5.111 ;
      RECT 89.09 3.795 89.1 4.158 ;
      RECT 89.09 4.88 89.095 5.112 ;
      RECT 89.085 3.795 89.09 4.118 ;
      RECT 89.085 4.887 89.09 5.113 ;
      RECT 89.08 3.795 89.085 4.09 ;
      RECT 89.075 4.905 89.085 5.114 ;
      RECT 89.07 3.795 89.08 4.07 ;
      RECT 89.065 4.925 89.075 5.116 ;
      RECT 89.055 4.942 89.065 5.117 ;
      RECT 89.02 4.965 89.055 5.12 ;
      RECT 88.965 4.983 89.02 5.126 ;
      RECT 88.879 4.991 88.965 5.135 ;
      RECT 88.793 5.002 88.879 5.146 ;
      RECT 88.707 5.012 88.793 5.157 ;
      RECT 88.621 5.022 88.707 5.169 ;
      RECT 88.535 5.032 88.621 5.18 ;
      RECT 88.515 5.038 88.535 5.186 ;
      RECT 88.435 5.04 88.515 5.19 ;
      RECT 88.43 5.039 88.435 5.195 ;
      RECT 88.422 5.038 88.43 5.195 ;
      RECT 88.336 5.034 88.422 5.193 ;
      RECT 88.25 5.026 88.336 5.19 ;
      RECT 88.164 5.017 88.25 5.186 ;
      RECT 88.078 5.009 88.164 5.183 ;
      RECT 87.992 5.001 88.078 5.179 ;
      RECT 87.906 4.992 87.992 5.176 ;
      RECT 87.82 4.984 87.906 5.172 ;
      RECT 87.765 4.977 87.81 5.17 ;
      RECT 87.68 4.97 87.765 5.168 ;
      RECT 87.606 4.962 87.68 5.164 ;
      RECT 87.52 4.954 87.606 5.161 ;
      RECT 87.517 4.95 87.52 5.159 ;
      RECT 87.431 4.946 87.517 5.158 ;
      RECT 87.345 4.938 87.431 5.155 ;
      RECT 87.26 4.933 87.345 5.152 ;
      RECT 87.174 4.93 87.26 5.149 ;
      RECT 87.088 4.928 87.174 5.146 ;
      RECT 87.002 4.925 87.088 5.143 ;
      RECT 86.916 4.922 87.002 5.14 ;
      RECT 86.83 4.919 86.916 5.137 ;
      RECT 86.754 4.917 86.83 5.134 ;
      RECT 86.668 4.914 86.754 5.131 ;
      RECT 86.582 4.911 86.668 5.129 ;
      RECT 86.496 4.909 86.582 5.126 ;
      RECT 86.41 4.906 86.496 5.123 ;
      RECT 86.35 4.897 86.41 5.121 ;
      RECT 88.86 4.515 88.935 4.775 ;
      RECT 88.84 4.495 88.845 4.775 ;
      RECT 88.16 4.28 88.265 4.575 ;
      RECT 82.605 4.255 82.675 4.515 ;
      RECT 88.5 4.13 88.505 4.501 ;
      RECT 88.49 4.185 88.495 4.501 ;
      RECT 88.795 3.355 88.855 3.615 ;
      RECT 88.85 4.51 88.86 4.775 ;
      RECT 88.845 4.5 88.85 4.775 ;
      RECT 88.765 4.447 88.84 4.775 ;
      RECT 88.79 3.355 88.795 3.635 ;
      RECT 88.78 3.355 88.79 3.655 ;
      RECT 88.765 3.355 88.78 3.685 ;
      RECT 88.75 3.355 88.765 3.728 ;
      RECT 88.745 4.39 88.765 4.775 ;
      RECT 88.735 3.355 88.75 3.765 ;
      RECT 88.73 4.37 88.745 4.775 ;
      RECT 88.73 3.355 88.735 3.788 ;
      RECT 88.72 3.355 88.73 3.813 ;
      RECT 88.69 4.337 88.73 4.775 ;
      RECT 88.695 3.355 88.72 3.863 ;
      RECT 88.69 3.355 88.695 3.918 ;
      RECT 88.685 3.355 88.69 3.96 ;
      RECT 88.675 4.3 88.69 4.775 ;
      RECT 88.68 3.355 88.685 4.003 ;
      RECT 88.675 3.355 88.68 4.068 ;
      RECT 88.67 3.355 88.675 4.09 ;
      RECT 88.67 4.288 88.675 4.64 ;
      RECT 88.665 3.355 88.67 4.158 ;
      RECT 88.665 4.28 88.67 4.623 ;
      RECT 88.66 3.355 88.665 4.203 ;
      RECT 88.655 4.262 88.665 4.6 ;
      RECT 88.655 3.355 88.66 4.24 ;
      RECT 88.645 3.355 88.655 4.58 ;
      RECT 88.64 3.355 88.645 4.563 ;
      RECT 88.635 3.355 88.64 4.548 ;
      RECT 88.63 3.355 88.635 4.533 ;
      RECT 88.61 3.355 88.63 4.523 ;
      RECT 88.605 3.355 88.61 4.513 ;
      RECT 88.595 3.355 88.605 4.509 ;
      RECT 88.59 3.632 88.595 4.508 ;
      RECT 88.585 3.655 88.59 4.507 ;
      RECT 88.58 3.685 88.585 4.506 ;
      RECT 88.575 3.712 88.58 4.505 ;
      RECT 88.57 3.74 88.575 4.505 ;
      RECT 88.565 3.767 88.57 4.505 ;
      RECT 88.56 3.787 88.565 4.505 ;
      RECT 88.555 3.815 88.56 4.505 ;
      RECT 88.545 3.857 88.555 4.505 ;
      RECT 88.535 3.902 88.545 4.504 ;
      RECT 88.53 3.955 88.535 4.503 ;
      RECT 88.525 3.987 88.53 4.502 ;
      RECT 88.52 4.007 88.525 4.501 ;
      RECT 88.515 4.045 88.52 4.501 ;
      RECT 88.51 4.067 88.515 4.501 ;
      RECT 88.505 4.092 88.51 4.501 ;
      RECT 88.495 4.157 88.5 4.501 ;
      RECT 88.48 4.217 88.49 4.501 ;
      RECT 88.465 4.227 88.48 4.501 ;
      RECT 88.445 4.237 88.465 4.501 ;
      RECT 88.415 4.242 88.445 4.498 ;
      RECT 88.355 4.252 88.415 4.495 ;
      RECT 88.335 4.261 88.355 4.5 ;
      RECT 88.31 4.267 88.335 4.513 ;
      RECT 88.29 4.272 88.31 4.528 ;
      RECT 88.265 4.277 88.29 4.575 ;
      RECT 88.136 4.279 88.16 4.575 ;
      RECT 88.05 4.274 88.136 4.575 ;
      RECT 88.01 4.271 88.05 4.575 ;
      RECT 87.96 4.273 88.01 4.555 ;
      RECT 87.93 4.277 87.96 4.555 ;
      RECT 87.851 4.287 87.93 4.555 ;
      RECT 87.765 4.302 87.851 4.556 ;
      RECT 87.715 4.312 87.765 4.557 ;
      RECT 87.707 4.315 87.715 4.557 ;
      RECT 87.621 4.317 87.707 4.558 ;
      RECT 87.535 4.321 87.621 4.558 ;
      RECT 87.449 4.325 87.535 4.559 ;
      RECT 87.363 4.328 87.449 4.56 ;
      RECT 87.277 4.332 87.363 4.56 ;
      RECT 87.191 4.336 87.277 4.561 ;
      RECT 87.105 4.339 87.191 4.562 ;
      RECT 87.019 4.343 87.105 4.562 ;
      RECT 86.933 4.347 87.019 4.563 ;
      RECT 86.847 4.351 86.933 4.564 ;
      RECT 86.761 4.354 86.847 4.564 ;
      RECT 86.675 4.358 86.761 4.565 ;
      RECT 86.645 4.36 86.675 4.565 ;
      RECT 86.559 4.363 86.645 4.566 ;
      RECT 86.473 4.367 86.559 4.567 ;
      RECT 86.387 4.371 86.473 4.568 ;
      RECT 86.301 4.374 86.387 4.568 ;
      RECT 86.215 4.378 86.301 4.569 ;
      RECT 86.18 4.383 86.215 4.57 ;
      RECT 86.125 4.393 86.18 4.577 ;
      RECT 86.1 4.405 86.125 4.587 ;
      RECT 86.065 4.418 86.1 4.595 ;
      RECT 86.025 4.435 86.065 4.618 ;
      RECT 86.005 4.448 86.025 4.645 ;
      RECT 85.975 4.46 86.005 4.673 ;
      RECT 85.97 4.468 85.975 4.693 ;
      RECT 85.965 4.471 85.97 4.703 ;
      RECT 85.915 4.483 85.965 4.737 ;
      RECT 85.905 4.498 85.915 4.77 ;
      RECT 85.895 4.504 85.905 4.783 ;
      RECT 85.885 4.511 85.895 4.795 ;
      RECT 85.86 4.524 85.885 4.813 ;
      RECT 85.845 4.539 85.86 4.835 ;
      RECT 85.835 4.547 85.845 4.851 ;
      RECT 85.82 4.556 85.835 4.866 ;
      RECT 85.81 4.566 85.82 4.88 ;
      RECT 85.791 4.579 85.81 4.897 ;
      RECT 85.705 4.624 85.791 4.962 ;
      RECT 85.69 4.669 85.705 5.02 ;
      RECT 85.685 4.678 85.69 5.033 ;
      RECT 85.675 4.685 85.685 5.038 ;
      RECT 85.67 4.69 85.675 5.042 ;
      RECT 85.65 4.7 85.67 5.049 ;
      RECT 85.625 4.72 85.65 5.063 ;
      RECT 85.59 4.745 85.625 5.083 ;
      RECT 85.575 4.768 85.59 5.098 ;
      RECT 85.565 4.778 85.575 5.103 ;
      RECT 85.555 4.786 85.565 5.11 ;
      RECT 85.545 4.795 85.555 5.116 ;
      RECT 85.525 4.807 85.545 5.118 ;
      RECT 85.515 4.82 85.525 5.12 ;
      RECT 85.49 4.835 85.515 5.123 ;
      RECT 85.47 4.852 85.49 5.127 ;
      RECT 85.43 4.88 85.47 5.133 ;
      RECT 85.365 4.927 85.43 5.142 ;
      RECT 85.35 4.96 85.365 5.15 ;
      RECT 85.345 4.967 85.35 5.152 ;
      RECT 85.295 4.992 85.345 5.157 ;
      RECT 85.28 5.016 85.295 5.164 ;
      RECT 85.23 5.021 85.28 5.165 ;
      RECT 85.144 5.025 85.23 5.165 ;
      RECT 85.058 5.025 85.144 5.165 ;
      RECT 84.972 5.025 85.058 5.166 ;
      RECT 84.886 5.025 84.972 5.166 ;
      RECT 84.8 5.025 84.886 5.166 ;
      RECT 84.734 5.025 84.8 5.166 ;
      RECT 84.648 5.025 84.734 5.167 ;
      RECT 84.562 5.025 84.648 5.167 ;
      RECT 84.476 5.026 84.562 5.168 ;
      RECT 84.39 5.026 84.476 5.168 ;
      RECT 84.304 5.026 84.39 5.168 ;
      RECT 84.218 5.026 84.304 5.169 ;
      RECT 84.132 5.026 84.218 5.169 ;
      RECT 84.046 5.027 84.132 5.17 ;
      RECT 83.96 5.027 84.046 5.17 ;
      RECT 83.94 5.027 83.96 5.17 ;
      RECT 83.854 5.027 83.94 5.17 ;
      RECT 83.768 5.027 83.854 5.17 ;
      RECT 83.682 5.028 83.768 5.17 ;
      RECT 83.596 5.028 83.682 5.17 ;
      RECT 83.51 5.028 83.596 5.17 ;
      RECT 83.424 5.029 83.51 5.17 ;
      RECT 83.338 5.029 83.424 5.17 ;
      RECT 83.252 5.029 83.338 5.17 ;
      RECT 83.166 5.029 83.252 5.17 ;
      RECT 83.08 5.03 83.166 5.17 ;
      RECT 83.03 5.027 83.08 5.17 ;
      RECT 83.02 5.025 83.03 5.169 ;
      RECT 83.016 5.025 83.02 5.168 ;
      RECT 82.93 5.02 83.016 5.163 ;
      RECT 82.908 5.013 82.93 5.157 ;
      RECT 82.822 5.004 82.908 5.151 ;
      RECT 82.736 4.991 82.822 5.142 ;
      RECT 82.65 4.977 82.736 5.132 ;
      RECT 82.605 4.967 82.65 5.125 ;
      RECT 82.585 4.255 82.605 4.533 ;
      RECT 82.585 4.96 82.605 5.121 ;
      RECT 82.555 4.255 82.585 4.555 ;
      RECT 82.545 4.927 82.585 5.118 ;
      RECT 82.54 4.255 82.555 4.575 ;
      RECT 82.54 4.892 82.545 5.116 ;
      RECT 82.535 4.255 82.54 4.7 ;
      RECT 82.535 4.852 82.54 5.116 ;
      RECT 82.525 4.255 82.535 5.116 ;
      RECT 82.45 4.255 82.525 5.11 ;
      RECT 82.42 4.255 82.45 5.1 ;
      RECT 82.415 4.255 82.42 5.092 ;
      RECT 82.41 4.297 82.415 5.085 ;
      RECT 82.4 4.366 82.41 5.076 ;
      RECT 82.395 4.436 82.4 5.028 ;
      RECT 82.39 4.5 82.395 4.925 ;
      RECT 82.385 4.535 82.39 4.88 ;
      RECT 82.383 4.572 82.385 4.772 ;
      RECT 82.38 4.58 82.383 4.765 ;
      RECT 82.375 4.645 82.38 4.708 ;
      RECT 86.45 3.735 86.73 4.015 ;
      RECT 86.44 3.735 86.73 3.878 ;
      RECT 86.395 3.6 86.655 3.86 ;
      RECT 86.395 3.715 86.71 3.86 ;
      RECT 86.395 3.685 86.705 3.86 ;
      RECT 86.395 3.672 86.695 3.86 ;
      RECT 86.395 3.662 86.69 3.86 ;
      RECT 82.37 3.645 82.63 3.905 ;
      RECT 86.14 3.195 86.4 3.455 ;
      RECT 86.13 3.22 86.4 3.415 ;
      RECT 86.125 3.22 86.13 3.414 ;
      RECT 86.055 3.215 86.125 3.406 ;
      RECT 85.97 3.202 86.055 3.389 ;
      RECT 85.966 3.194 85.97 3.379 ;
      RECT 85.88 3.187 85.966 3.369 ;
      RECT 85.871 3.179 85.88 3.359 ;
      RECT 85.785 3.172 85.871 3.347 ;
      RECT 85.765 3.163 85.785 3.333 ;
      RECT 85.71 3.158 85.765 3.325 ;
      RECT 85.7 3.152 85.71 3.319 ;
      RECT 85.68 3.15 85.7 3.315 ;
      RECT 85.672 3.149 85.68 3.311 ;
      RECT 85.586 3.141 85.672 3.3 ;
      RECT 85.5 3.127 85.586 3.28 ;
      RECT 85.44 3.115 85.5 3.265 ;
      RECT 85.43 3.11 85.44 3.26 ;
      RECT 85.38 3.11 85.43 3.262 ;
      RECT 85.333 3.112 85.38 3.266 ;
      RECT 85.247 3.119 85.333 3.271 ;
      RECT 85.161 3.127 85.247 3.277 ;
      RECT 85.075 3.136 85.161 3.283 ;
      RECT 85.016 3.142 85.075 3.288 ;
      RECT 84.93 3.147 85.016 3.294 ;
      RECT 84.855 3.152 84.93 3.3 ;
      RECT 84.816 3.154 84.855 3.305 ;
      RECT 84.73 3.151 84.816 3.31 ;
      RECT 84.645 3.149 84.73 3.317 ;
      RECT 84.613 3.148 84.645 3.32 ;
      RECT 84.527 3.147 84.613 3.321 ;
      RECT 84.441 3.146 84.527 3.322 ;
      RECT 84.355 3.145 84.441 3.322 ;
      RECT 84.269 3.144 84.355 3.323 ;
      RECT 84.183 3.143 84.269 3.324 ;
      RECT 84.097 3.142 84.183 3.325 ;
      RECT 84.011 3.141 84.097 3.325 ;
      RECT 83.925 3.14 84.011 3.326 ;
      RECT 83.875 3.14 83.925 3.327 ;
      RECT 83.861 3.141 83.875 3.327 ;
      RECT 83.775 3.148 83.861 3.328 ;
      RECT 83.701 3.159 83.775 3.329 ;
      RECT 83.615 3.168 83.701 3.33 ;
      RECT 83.58 3.175 83.615 3.345 ;
      RECT 83.555 3.178 83.58 3.375 ;
      RECT 83.53 3.187 83.555 3.404 ;
      RECT 83.52 3.198 83.53 3.424 ;
      RECT 83.51 3.206 83.52 3.438 ;
      RECT 83.505 3.212 83.51 3.448 ;
      RECT 83.48 3.229 83.505 3.465 ;
      RECT 83.465 3.251 83.48 3.493 ;
      RECT 83.435 3.277 83.465 3.523 ;
      RECT 83.415 3.306 83.435 3.553 ;
      RECT 83.41 3.321 83.415 3.57 ;
      RECT 83.39 3.336 83.41 3.585 ;
      RECT 83.38 3.354 83.39 3.603 ;
      RECT 83.37 3.365 83.38 3.618 ;
      RECT 83.32 3.397 83.37 3.644 ;
      RECT 83.315 3.427 83.32 3.664 ;
      RECT 83.305 3.44 83.315 3.67 ;
      RECT 83.296 3.45 83.305 3.678 ;
      RECT 83.285 3.461 83.296 3.686 ;
      RECT 83.28 3.471 83.285 3.692 ;
      RECT 83.265 3.492 83.28 3.699 ;
      RECT 83.25 3.522 83.265 3.707 ;
      RECT 83.215 3.552 83.25 3.713 ;
      RECT 83.19 3.57 83.215 3.72 ;
      RECT 83.14 3.578 83.19 3.729 ;
      RECT 83.115 3.583 83.14 3.738 ;
      RECT 83.06 3.589 83.115 3.748 ;
      RECT 83.055 3.594 83.06 3.756 ;
      RECT 83.041 3.597 83.055 3.758 ;
      RECT 82.955 3.609 83.041 3.77 ;
      RECT 82.945 3.621 82.955 3.783 ;
      RECT 82.86 3.634 82.945 3.795 ;
      RECT 82.816 3.651 82.86 3.809 ;
      RECT 82.73 3.668 82.816 3.825 ;
      RECT 82.7 3.682 82.73 3.839 ;
      RECT 82.69 3.687 82.7 3.844 ;
      RECT 82.63 3.69 82.69 3.853 ;
      RECT 85.52 3.96 85.78 4.22 ;
      RECT 85.52 3.96 85.8 4.073 ;
      RECT 85.52 3.96 85.825 4.04 ;
      RECT 85.52 3.96 85.83 4.02 ;
      RECT 85.57 3.735 85.85 4.015 ;
      RECT 85.125 4.47 85.385 4.73 ;
      RECT 85.115 4.327 85.31 4.668 ;
      RECT 85.11 4.435 85.325 4.66 ;
      RECT 85.105 4.485 85.385 4.65 ;
      RECT 85.095 4.562 85.385 4.635 ;
      RECT 85.115 4.41 85.325 4.668 ;
      RECT 85.125 4.285 85.31 4.73 ;
      RECT 85.125 4.18 85.29 4.73 ;
      RECT 85.135 4.167 85.29 4.73 ;
      RECT 85.135 4.125 85.28 4.73 ;
      RECT 85.14 4.05 85.28 4.73 ;
      RECT 85.17 3.7 85.28 4.73 ;
      RECT 85.175 3.43 85.3 4.053 ;
      RECT 85.145 4.005 85.3 4.053 ;
      RECT 85.16 3.807 85.28 4.73 ;
      RECT 85.15 3.917 85.3 4.053 ;
      RECT 85.175 3.43 85.315 3.91 ;
      RECT 85.175 3.43 85.335 3.785 ;
      RECT 85.14 3.43 85.4 3.69 ;
      RECT 84.61 3.735 84.89 4.015 ;
      RECT 84.595 3.735 84.89 3.995 ;
      RECT 82.65 4.6 82.91 4.86 ;
      RECT 84.435 4.455 84.695 4.715 ;
      RECT 84.415 4.475 84.695 4.69 ;
      RECT 84.372 4.475 84.415 4.689 ;
      RECT 84.286 4.476 84.372 4.686 ;
      RECT 84.2 4.477 84.286 4.682 ;
      RECT 84.125 4.479 84.2 4.679 ;
      RECT 84.102 4.48 84.125 4.677 ;
      RECT 84.016 4.481 84.102 4.675 ;
      RECT 83.93 4.482 84.016 4.672 ;
      RECT 83.906 4.483 83.93 4.67 ;
      RECT 83.82 4.485 83.906 4.667 ;
      RECT 83.735 4.487 83.82 4.668 ;
      RECT 83.678 4.488 83.735 4.674 ;
      RECT 83.592 4.49 83.678 4.684 ;
      RECT 83.506 4.493 83.592 4.697 ;
      RECT 83.42 4.495 83.506 4.709 ;
      RECT 83.406 4.496 83.42 4.716 ;
      RECT 83.32 4.497 83.406 4.724 ;
      RECT 83.28 4.499 83.32 4.733 ;
      RECT 83.271 4.5 83.28 4.736 ;
      RECT 83.185 4.508 83.271 4.742 ;
      RECT 83.165 4.517 83.185 4.75 ;
      RECT 83.08 4.532 83.165 4.758 ;
      RECT 83.02 4.555 83.08 4.769 ;
      RECT 83.01 4.567 83.02 4.774 ;
      RECT 82.97 4.577 83.01 4.778 ;
      RECT 82.915 4.594 82.97 4.786 ;
      RECT 82.91 4.604 82.915 4.79 ;
      RECT 83.976 3.735 84.035 4.132 ;
      RECT 83.89 3.735 84.095 4.123 ;
      RECT 83.885 3.765 84.095 4.118 ;
      RECT 83.851 3.765 84.095 4.116 ;
      RECT 83.765 3.765 84.095 4.11 ;
      RECT 83.72 3.765 84.115 4.088 ;
      RECT 83.72 3.765 84.135 4.043 ;
      RECT 83.68 3.765 84.135 4.033 ;
      RECT 83.89 3.735 84.17 4.015 ;
      RECT 83.625 3.735 83.885 3.995 ;
      RECT 82.81 3.215 83.07 3.475 ;
      RECT 82.89 3.175 83.17 3.455 ;
      RECT 77.255 8.505 77.575 8.83 ;
      RECT 77.285 7.98 77.455 8.83 ;
      RECT 77.285 7.98 77.46 8.33 ;
      RECT 77.285 7.98 78.26 8.155 ;
      RECT 78.085 3.26 78.26 8.155 ;
      RECT 78.03 3.26 78.38 3.61 ;
      RECT 78.055 8.94 78.38 9.265 ;
      RECT 76.94 9.03 78.38 9.2 ;
      RECT 76.94 3.69 77.1 9.2 ;
      RECT 77.255 3.66 77.575 3.98 ;
      RECT 76.94 3.69 77.575 3.86 ;
      RECT 65.665 4.295 65.945 4.575 ;
      RECT 65.635 4.295 65.945 4.56 ;
      RECT 65.63 4.295 65.945 4.558 ;
      RECT 65.625 2.625 65.795 4.552 ;
      RECT 65.62 4.262 65.89 4.545 ;
      RECT 65.615 4.295 65.945 4.538 ;
      RECT 65.585 4.265 65.89 4.525 ;
      RECT 65.585 4.292 65.91 4.525 ;
      RECT 65.585 4.282 65.905 4.525 ;
      RECT 65.585 4.267 65.9 4.525 ;
      RECT 65.625 4.257 65.89 4.552 ;
      RECT 65.625 4.252 65.88 4.552 ;
      RECT 65.625 4.251 65.865 4.552 ;
      RECT 75.595 2.635 75.945 2.985 ;
      RECT 75.59 2.635 75.945 2.89 ;
      RECT 65.625 2.625 75.835 2.795 ;
      RECT 75.27 4.145 75.64 4.515 ;
      RECT 75.355 3.53 75.525 4.515 ;
      RECT 71.375 3.75 71.61 4.01 ;
      RECT 74.52 3.53 74.685 3.79 ;
      RECT 74.425 3.52 74.44 3.79 ;
      RECT 74.52 3.53 75.525 3.71 ;
      RECT 73.025 3.09 73.065 3.23 ;
      RECT 74.44 3.525 74.52 3.79 ;
      RECT 74.385 3.52 74.425 3.756 ;
      RECT 74.371 3.52 74.385 3.756 ;
      RECT 74.285 3.525 74.371 3.758 ;
      RECT 74.24 3.532 74.285 3.76 ;
      RECT 74.21 3.532 74.24 3.762 ;
      RECT 74.185 3.527 74.21 3.764 ;
      RECT 74.155 3.523 74.185 3.773 ;
      RECT 74.145 3.52 74.155 3.785 ;
      RECT 74.14 3.52 74.145 3.793 ;
      RECT 74.135 3.52 74.14 3.798 ;
      RECT 74.125 3.519 74.135 3.808 ;
      RECT 74.12 3.518 74.125 3.818 ;
      RECT 74.105 3.517 74.12 3.823 ;
      RECT 74.077 3.514 74.105 3.85 ;
      RECT 73.991 3.506 74.077 3.85 ;
      RECT 73.905 3.495 73.991 3.85 ;
      RECT 73.865 3.48 73.905 3.85 ;
      RECT 73.825 3.454 73.865 3.85 ;
      RECT 73.82 3.436 73.825 3.662 ;
      RECT 73.81 3.432 73.82 3.652 ;
      RECT 73.795 3.422 73.81 3.639 ;
      RECT 73.775 3.406 73.795 3.624 ;
      RECT 73.76 3.391 73.775 3.609 ;
      RECT 73.75 3.38 73.76 3.599 ;
      RECT 73.725 3.364 73.75 3.588 ;
      RECT 73.72 3.351 73.725 3.578 ;
      RECT 73.715 3.347 73.72 3.573 ;
      RECT 73.66 3.333 73.715 3.551 ;
      RECT 73.621 3.314 73.66 3.515 ;
      RECT 73.535 3.288 73.621 3.468 ;
      RECT 73.531 3.27 73.535 3.434 ;
      RECT 73.445 3.251 73.531 3.412 ;
      RECT 73.44 3.233 73.445 3.39 ;
      RECT 73.435 3.231 73.44 3.388 ;
      RECT 73.425 3.23 73.435 3.383 ;
      RECT 73.365 3.217 73.425 3.369 ;
      RECT 73.32 3.195 73.365 3.348 ;
      RECT 73.26 3.172 73.32 3.327 ;
      RECT 73.196 3.147 73.26 3.302 ;
      RECT 73.11 3.117 73.196 3.271 ;
      RECT 73.095 3.097 73.11 3.25 ;
      RECT 73.065 3.092 73.095 3.241 ;
      RECT 73.012 3.09 73.025 3.23 ;
      RECT 72.926 3.09 73.012 3.232 ;
      RECT 72.84 3.09 72.926 3.234 ;
      RECT 72.82 3.09 72.84 3.238 ;
      RECT 72.775 3.092 72.82 3.249 ;
      RECT 72.735 3.102 72.775 3.265 ;
      RECT 72.731 3.111 72.735 3.273 ;
      RECT 72.645 3.131 72.731 3.289 ;
      RECT 72.635 3.15 72.645 3.307 ;
      RECT 72.63 3.152 72.635 3.31 ;
      RECT 72.62 3.156 72.63 3.313 ;
      RECT 72.6 3.161 72.62 3.323 ;
      RECT 72.57 3.171 72.6 3.343 ;
      RECT 72.565 3.178 72.57 3.357 ;
      RECT 72.555 3.182 72.565 3.364 ;
      RECT 72.54 3.19 72.555 3.375 ;
      RECT 72.53 3.2 72.54 3.386 ;
      RECT 72.52 3.207 72.53 3.394 ;
      RECT 72.495 3.22 72.52 3.409 ;
      RECT 72.431 3.256 72.495 3.448 ;
      RECT 72.345 3.319 72.431 3.512 ;
      RECT 72.31 3.37 72.345 3.565 ;
      RECT 72.305 3.387 72.31 3.582 ;
      RECT 72.29 3.396 72.305 3.589 ;
      RECT 72.27 3.411 72.29 3.603 ;
      RECT 72.265 3.422 72.27 3.613 ;
      RECT 72.245 3.435 72.265 3.623 ;
      RECT 72.24 3.445 72.245 3.633 ;
      RECT 72.225 3.45 72.24 3.642 ;
      RECT 72.215 3.46 72.225 3.653 ;
      RECT 72.185 3.477 72.215 3.67 ;
      RECT 72.175 3.495 72.185 3.688 ;
      RECT 72.16 3.506 72.175 3.699 ;
      RECT 72.12 3.53 72.16 3.715 ;
      RECT 72.085 3.564 72.12 3.732 ;
      RECT 72.055 3.587 72.085 3.744 ;
      RECT 72.04 3.597 72.055 3.753 ;
      RECT 72 3.607 72.04 3.764 ;
      RECT 71.98 3.618 72 3.776 ;
      RECT 71.975 3.622 71.98 3.783 ;
      RECT 71.96 3.626 71.975 3.788 ;
      RECT 71.95 3.631 71.96 3.793 ;
      RECT 71.945 3.634 71.95 3.796 ;
      RECT 71.915 3.64 71.945 3.803 ;
      RECT 71.88 3.65 71.915 3.817 ;
      RECT 71.82 3.665 71.88 3.837 ;
      RECT 71.765 3.685 71.82 3.861 ;
      RECT 71.736 3.7 71.765 3.879 ;
      RECT 71.65 3.72 71.736 3.904 ;
      RECT 71.645 3.735 71.65 3.924 ;
      RECT 71.635 3.738 71.645 3.925 ;
      RECT 71.61 3.745 71.635 4.01 ;
      RECT 64.605 8.945 64.955 9.295 ;
      RECT 73.43 8.89 73.78 9.24 ;
      RECT 64.605 8.975 65.755 9.175 ;
      RECT 65.755 8.965 73.78 9.165 ;
      RECT 72.025 4.98 72.035 5.17 ;
      RECT 70.285 4.855 70.565 5.135 ;
      RECT 73.33 3.795 73.335 4.28 ;
      RECT 73.225 3.795 73.285 4.055 ;
      RECT 73.55 4.765 73.555 4.84 ;
      RECT 73.54 4.632 73.55 4.875 ;
      RECT 73.53 4.467 73.54 4.896 ;
      RECT 73.525 4.337 73.53 4.912 ;
      RECT 73.515 4.227 73.525 4.928 ;
      RECT 73.51 4.126 73.515 4.945 ;
      RECT 73.505 4.108 73.51 4.955 ;
      RECT 73.5 4.09 73.505 4.965 ;
      RECT 73.49 4.065 73.5 4.98 ;
      RECT 73.485 4.045 73.49 4.995 ;
      RECT 73.465 3.795 73.485 5.02 ;
      RECT 73.45 3.795 73.465 5.053 ;
      RECT 73.42 3.795 73.45 5.075 ;
      RECT 73.4 3.795 73.42 5.089 ;
      RECT 73.38 3.795 73.4 4.605 ;
      RECT 73.395 4.672 73.4 5.094 ;
      RECT 73.39 4.702 73.395 5.096 ;
      RECT 73.385 4.715 73.39 5.099 ;
      RECT 73.38 4.725 73.385 5.103 ;
      RECT 73.375 3.795 73.38 4.523 ;
      RECT 73.375 4.735 73.38 5.105 ;
      RECT 73.37 3.795 73.375 4.5 ;
      RECT 73.36 4.757 73.375 5.105 ;
      RECT 73.355 3.795 73.37 4.445 ;
      RECT 73.35 4.782 73.36 5.105 ;
      RECT 73.35 3.795 73.355 4.39 ;
      RECT 73.34 3.795 73.35 4.338 ;
      RECT 73.345 4.795 73.35 5.106 ;
      RECT 73.34 4.807 73.345 5.107 ;
      RECT 73.335 3.795 73.34 4.298 ;
      RECT 73.335 4.82 73.34 5.108 ;
      RECT 73.32 4.835 73.335 5.109 ;
      RECT 73.325 3.795 73.33 4.26 ;
      RECT 73.32 3.795 73.325 4.225 ;
      RECT 73.315 3.795 73.32 4.2 ;
      RECT 73.31 4.862 73.32 5.111 ;
      RECT 73.305 3.795 73.315 4.158 ;
      RECT 73.305 4.88 73.31 5.112 ;
      RECT 73.3 3.795 73.305 4.118 ;
      RECT 73.3 4.887 73.305 5.113 ;
      RECT 73.295 3.795 73.3 4.09 ;
      RECT 73.29 4.905 73.3 5.114 ;
      RECT 73.285 3.795 73.295 4.07 ;
      RECT 73.28 4.925 73.29 5.116 ;
      RECT 73.27 4.942 73.28 5.117 ;
      RECT 73.235 4.965 73.27 5.12 ;
      RECT 73.18 4.983 73.235 5.126 ;
      RECT 73.094 4.991 73.18 5.135 ;
      RECT 73.008 5.002 73.094 5.146 ;
      RECT 72.922 5.012 73.008 5.157 ;
      RECT 72.836 5.022 72.922 5.169 ;
      RECT 72.75 5.032 72.836 5.18 ;
      RECT 72.73 5.038 72.75 5.186 ;
      RECT 72.65 5.04 72.73 5.19 ;
      RECT 72.645 5.039 72.65 5.195 ;
      RECT 72.637 5.038 72.645 5.195 ;
      RECT 72.551 5.034 72.637 5.193 ;
      RECT 72.465 5.026 72.551 5.19 ;
      RECT 72.379 5.017 72.465 5.186 ;
      RECT 72.293 5.009 72.379 5.183 ;
      RECT 72.207 5.001 72.293 5.179 ;
      RECT 72.121 4.992 72.207 5.176 ;
      RECT 72.035 4.984 72.121 5.172 ;
      RECT 71.98 4.977 72.025 5.17 ;
      RECT 71.895 4.97 71.98 5.168 ;
      RECT 71.821 4.962 71.895 5.164 ;
      RECT 71.735 4.954 71.821 5.161 ;
      RECT 71.732 4.95 71.735 5.159 ;
      RECT 71.646 4.946 71.732 5.158 ;
      RECT 71.56 4.938 71.646 5.155 ;
      RECT 71.475 4.933 71.56 5.152 ;
      RECT 71.389 4.93 71.475 5.149 ;
      RECT 71.303 4.928 71.389 5.146 ;
      RECT 71.217 4.925 71.303 5.143 ;
      RECT 71.131 4.922 71.217 5.14 ;
      RECT 71.045 4.919 71.131 5.137 ;
      RECT 70.969 4.917 71.045 5.134 ;
      RECT 70.883 4.914 70.969 5.131 ;
      RECT 70.797 4.911 70.883 5.129 ;
      RECT 70.711 4.909 70.797 5.126 ;
      RECT 70.625 4.906 70.711 5.123 ;
      RECT 70.565 4.897 70.625 5.121 ;
      RECT 73.075 4.515 73.15 4.775 ;
      RECT 73.055 4.495 73.06 4.775 ;
      RECT 72.375 4.28 72.48 4.575 ;
      RECT 66.82 4.255 66.89 4.515 ;
      RECT 72.715 4.13 72.72 4.501 ;
      RECT 72.705 4.185 72.71 4.501 ;
      RECT 73.01 3.355 73.07 3.615 ;
      RECT 73.065 4.51 73.075 4.775 ;
      RECT 73.06 4.5 73.065 4.775 ;
      RECT 72.98 4.447 73.055 4.775 ;
      RECT 73.005 3.355 73.01 3.635 ;
      RECT 72.995 3.355 73.005 3.655 ;
      RECT 72.98 3.355 72.995 3.685 ;
      RECT 72.965 3.355 72.98 3.728 ;
      RECT 72.96 4.39 72.98 4.775 ;
      RECT 72.95 3.355 72.965 3.765 ;
      RECT 72.945 4.37 72.96 4.775 ;
      RECT 72.945 3.355 72.95 3.788 ;
      RECT 72.935 3.355 72.945 3.813 ;
      RECT 72.905 4.337 72.945 4.775 ;
      RECT 72.91 3.355 72.935 3.863 ;
      RECT 72.905 3.355 72.91 3.918 ;
      RECT 72.9 3.355 72.905 3.96 ;
      RECT 72.89 4.3 72.905 4.775 ;
      RECT 72.895 3.355 72.9 4.003 ;
      RECT 72.89 3.355 72.895 4.068 ;
      RECT 72.885 3.355 72.89 4.09 ;
      RECT 72.885 4.288 72.89 4.64 ;
      RECT 72.88 3.355 72.885 4.158 ;
      RECT 72.88 4.28 72.885 4.623 ;
      RECT 72.875 3.355 72.88 4.203 ;
      RECT 72.87 4.262 72.88 4.6 ;
      RECT 72.87 3.355 72.875 4.24 ;
      RECT 72.86 3.355 72.87 4.58 ;
      RECT 72.855 3.355 72.86 4.563 ;
      RECT 72.85 3.355 72.855 4.548 ;
      RECT 72.845 3.355 72.85 4.533 ;
      RECT 72.825 3.355 72.845 4.523 ;
      RECT 72.82 3.355 72.825 4.513 ;
      RECT 72.81 3.355 72.82 4.509 ;
      RECT 72.805 3.632 72.81 4.508 ;
      RECT 72.8 3.655 72.805 4.507 ;
      RECT 72.795 3.685 72.8 4.506 ;
      RECT 72.79 3.712 72.795 4.505 ;
      RECT 72.785 3.74 72.79 4.505 ;
      RECT 72.78 3.767 72.785 4.505 ;
      RECT 72.775 3.787 72.78 4.505 ;
      RECT 72.77 3.815 72.775 4.505 ;
      RECT 72.76 3.857 72.77 4.505 ;
      RECT 72.75 3.902 72.76 4.504 ;
      RECT 72.745 3.955 72.75 4.503 ;
      RECT 72.74 3.987 72.745 4.502 ;
      RECT 72.735 4.007 72.74 4.501 ;
      RECT 72.73 4.045 72.735 4.501 ;
      RECT 72.725 4.067 72.73 4.501 ;
      RECT 72.72 4.092 72.725 4.501 ;
      RECT 72.71 4.157 72.715 4.501 ;
      RECT 72.695 4.217 72.705 4.501 ;
      RECT 72.68 4.227 72.695 4.501 ;
      RECT 72.66 4.237 72.68 4.501 ;
      RECT 72.63 4.242 72.66 4.498 ;
      RECT 72.57 4.252 72.63 4.495 ;
      RECT 72.55 4.261 72.57 4.5 ;
      RECT 72.525 4.267 72.55 4.513 ;
      RECT 72.505 4.272 72.525 4.528 ;
      RECT 72.48 4.277 72.505 4.575 ;
      RECT 72.351 4.279 72.375 4.575 ;
      RECT 72.265 4.274 72.351 4.575 ;
      RECT 72.225 4.271 72.265 4.575 ;
      RECT 72.175 4.273 72.225 4.555 ;
      RECT 72.145 4.277 72.175 4.555 ;
      RECT 72.066 4.287 72.145 4.555 ;
      RECT 71.98 4.302 72.066 4.556 ;
      RECT 71.93 4.312 71.98 4.557 ;
      RECT 71.922 4.315 71.93 4.557 ;
      RECT 71.836 4.317 71.922 4.558 ;
      RECT 71.75 4.321 71.836 4.558 ;
      RECT 71.664 4.325 71.75 4.559 ;
      RECT 71.578 4.328 71.664 4.56 ;
      RECT 71.492 4.332 71.578 4.56 ;
      RECT 71.406 4.336 71.492 4.561 ;
      RECT 71.32 4.339 71.406 4.562 ;
      RECT 71.234 4.343 71.32 4.562 ;
      RECT 71.148 4.347 71.234 4.563 ;
      RECT 71.062 4.351 71.148 4.564 ;
      RECT 70.976 4.354 71.062 4.564 ;
      RECT 70.89 4.358 70.976 4.565 ;
      RECT 70.86 4.36 70.89 4.565 ;
      RECT 70.774 4.363 70.86 4.566 ;
      RECT 70.688 4.367 70.774 4.567 ;
      RECT 70.602 4.371 70.688 4.568 ;
      RECT 70.516 4.374 70.602 4.568 ;
      RECT 70.43 4.378 70.516 4.569 ;
      RECT 70.395 4.383 70.43 4.57 ;
      RECT 70.34 4.393 70.395 4.577 ;
      RECT 70.315 4.405 70.34 4.587 ;
      RECT 70.28 4.418 70.315 4.595 ;
      RECT 70.24 4.435 70.28 4.618 ;
      RECT 70.22 4.448 70.24 4.645 ;
      RECT 70.19 4.46 70.22 4.673 ;
      RECT 70.185 4.468 70.19 4.693 ;
      RECT 70.18 4.471 70.185 4.703 ;
      RECT 70.13 4.483 70.18 4.737 ;
      RECT 70.12 4.498 70.13 4.77 ;
      RECT 70.11 4.504 70.12 4.783 ;
      RECT 70.1 4.511 70.11 4.795 ;
      RECT 70.075 4.524 70.1 4.813 ;
      RECT 70.06 4.539 70.075 4.835 ;
      RECT 70.05 4.547 70.06 4.851 ;
      RECT 70.035 4.556 70.05 4.866 ;
      RECT 70.025 4.566 70.035 4.88 ;
      RECT 70.006 4.579 70.025 4.897 ;
      RECT 69.92 4.624 70.006 4.962 ;
      RECT 69.905 4.669 69.92 5.02 ;
      RECT 69.9 4.678 69.905 5.033 ;
      RECT 69.89 4.685 69.9 5.038 ;
      RECT 69.885 4.69 69.89 5.042 ;
      RECT 69.865 4.7 69.885 5.049 ;
      RECT 69.84 4.72 69.865 5.063 ;
      RECT 69.805 4.745 69.84 5.083 ;
      RECT 69.79 4.768 69.805 5.098 ;
      RECT 69.78 4.778 69.79 5.103 ;
      RECT 69.77 4.786 69.78 5.11 ;
      RECT 69.76 4.795 69.77 5.116 ;
      RECT 69.74 4.807 69.76 5.118 ;
      RECT 69.73 4.82 69.74 5.12 ;
      RECT 69.705 4.835 69.73 5.123 ;
      RECT 69.685 4.852 69.705 5.127 ;
      RECT 69.645 4.88 69.685 5.133 ;
      RECT 69.58 4.927 69.645 5.142 ;
      RECT 69.565 4.96 69.58 5.15 ;
      RECT 69.56 4.967 69.565 5.152 ;
      RECT 69.51 4.992 69.56 5.157 ;
      RECT 69.495 5.016 69.51 5.164 ;
      RECT 69.445 5.021 69.495 5.165 ;
      RECT 69.359 5.025 69.445 5.165 ;
      RECT 69.273 5.025 69.359 5.165 ;
      RECT 69.187 5.025 69.273 5.166 ;
      RECT 69.101 5.025 69.187 5.166 ;
      RECT 69.015 5.025 69.101 5.166 ;
      RECT 68.949 5.025 69.015 5.166 ;
      RECT 68.863 5.025 68.949 5.167 ;
      RECT 68.777 5.025 68.863 5.167 ;
      RECT 68.691 5.026 68.777 5.168 ;
      RECT 68.605 5.026 68.691 5.168 ;
      RECT 68.519 5.026 68.605 5.168 ;
      RECT 68.433 5.026 68.519 5.169 ;
      RECT 68.347 5.026 68.433 5.169 ;
      RECT 68.261 5.027 68.347 5.17 ;
      RECT 68.175 5.027 68.261 5.17 ;
      RECT 68.155 5.027 68.175 5.17 ;
      RECT 68.069 5.027 68.155 5.17 ;
      RECT 67.983 5.027 68.069 5.17 ;
      RECT 67.897 5.028 67.983 5.17 ;
      RECT 67.811 5.028 67.897 5.17 ;
      RECT 67.725 5.028 67.811 5.17 ;
      RECT 67.639 5.029 67.725 5.17 ;
      RECT 67.553 5.029 67.639 5.17 ;
      RECT 67.467 5.029 67.553 5.17 ;
      RECT 67.381 5.029 67.467 5.17 ;
      RECT 67.295 5.03 67.381 5.17 ;
      RECT 67.245 5.027 67.295 5.17 ;
      RECT 67.235 5.025 67.245 5.169 ;
      RECT 67.231 5.025 67.235 5.168 ;
      RECT 67.145 5.02 67.231 5.163 ;
      RECT 67.123 5.013 67.145 5.157 ;
      RECT 67.037 5.004 67.123 5.151 ;
      RECT 66.951 4.991 67.037 5.142 ;
      RECT 66.865 4.977 66.951 5.132 ;
      RECT 66.82 4.967 66.865 5.125 ;
      RECT 66.8 4.255 66.82 4.533 ;
      RECT 66.8 4.96 66.82 5.121 ;
      RECT 66.77 4.255 66.8 4.555 ;
      RECT 66.76 4.927 66.8 5.118 ;
      RECT 66.755 4.255 66.77 4.575 ;
      RECT 66.755 4.892 66.76 5.116 ;
      RECT 66.75 4.255 66.755 4.7 ;
      RECT 66.75 4.852 66.755 5.116 ;
      RECT 66.74 4.255 66.75 5.116 ;
      RECT 66.665 4.255 66.74 5.11 ;
      RECT 66.635 4.255 66.665 5.1 ;
      RECT 66.63 4.255 66.635 5.092 ;
      RECT 66.625 4.297 66.63 5.085 ;
      RECT 66.615 4.366 66.625 5.076 ;
      RECT 66.61 4.436 66.615 5.028 ;
      RECT 66.605 4.5 66.61 4.925 ;
      RECT 66.6 4.535 66.605 4.88 ;
      RECT 66.598 4.572 66.6 4.772 ;
      RECT 66.595 4.58 66.598 4.765 ;
      RECT 66.59 4.645 66.595 4.708 ;
      RECT 70.665 3.735 70.945 4.015 ;
      RECT 70.655 3.735 70.945 3.878 ;
      RECT 70.61 3.6 70.87 3.86 ;
      RECT 70.61 3.715 70.925 3.86 ;
      RECT 70.61 3.685 70.92 3.86 ;
      RECT 70.61 3.672 70.91 3.86 ;
      RECT 70.61 3.662 70.905 3.86 ;
      RECT 66.585 3.645 66.845 3.905 ;
      RECT 70.355 3.195 70.615 3.455 ;
      RECT 70.345 3.22 70.615 3.415 ;
      RECT 70.34 3.22 70.345 3.414 ;
      RECT 70.27 3.215 70.34 3.406 ;
      RECT 70.185 3.202 70.27 3.389 ;
      RECT 70.181 3.194 70.185 3.379 ;
      RECT 70.095 3.187 70.181 3.369 ;
      RECT 70.086 3.179 70.095 3.359 ;
      RECT 70 3.172 70.086 3.347 ;
      RECT 69.98 3.163 70 3.333 ;
      RECT 69.925 3.158 69.98 3.325 ;
      RECT 69.915 3.152 69.925 3.319 ;
      RECT 69.895 3.15 69.915 3.315 ;
      RECT 69.887 3.149 69.895 3.311 ;
      RECT 69.801 3.141 69.887 3.3 ;
      RECT 69.715 3.127 69.801 3.28 ;
      RECT 69.655 3.115 69.715 3.265 ;
      RECT 69.645 3.11 69.655 3.26 ;
      RECT 69.595 3.11 69.645 3.262 ;
      RECT 69.548 3.112 69.595 3.266 ;
      RECT 69.462 3.119 69.548 3.271 ;
      RECT 69.376 3.127 69.462 3.277 ;
      RECT 69.29 3.136 69.376 3.283 ;
      RECT 69.231 3.142 69.29 3.288 ;
      RECT 69.145 3.147 69.231 3.294 ;
      RECT 69.07 3.152 69.145 3.3 ;
      RECT 69.031 3.154 69.07 3.305 ;
      RECT 68.945 3.151 69.031 3.31 ;
      RECT 68.86 3.149 68.945 3.317 ;
      RECT 68.828 3.148 68.86 3.32 ;
      RECT 68.742 3.147 68.828 3.321 ;
      RECT 68.656 3.146 68.742 3.322 ;
      RECT 68.57 3.145 68.656 3.322 ;
      RECT 68.484 3.144 68.57 3.323 ;
      RECT 68.398 3.143 68.484 3.324 ;
      RECT 68.312 3.142 68.398 3.325 ;
      RECT 68.226 3.141 68.312 3.325 ;
      RECT 68.14 3.14 68.226 3.326 ;
      RECT 68.09 3.14 68.14 3.327 ;
      RECT 68.076 3.141 68.09 3.327 ;
      RECT 67.99 3.148 68.076 3.328 ;
      RECT 67.916 3.159 67.99 3.329 ;
      RECT 67.83 3.168 67.916 3.33 ;
      RECT 67.795 3.175 67.83 3.345 ;
      RECT 67.77 3.178 67.795 3.375 ;
      RECT 67.745 3.187 67.77 3.404 ;
      RECT 67.735 3.198 67.745 3.424 ;
      RECT 67.725 3.206 67.735 3.438 ;
      RECT 67.72 3.212 67.725 3.448 ;
      RECT 67.695 3.229 67.72 3.465 ;
      RECT 67.68 3.251 67.695 3.493 ;
      RECT 67.65 3.277 67.68 3.523 ;
      RECT 67.63 3.306 67.65 3.553 ;
      RECT 67.625 3.321 67.63 3.57 ;
      RECT 67.605 3.336 67.625 3.585 ;
      RECT 67.595 3.354 67.605 3.603 ;
      RECT 67.585 3.365 67.595 3.618 ;
      RECT 67.535 3.397 67.585 3.644 ;
      RECT 67.53 3.427 67.535 3.664 ;
      RECT 67.52 3.44 67.53 3.67 ;
      RECT 67.511 3.45 67.52 3.678 ;
      RECT 67.5 3.461 67.511 3.686 ;
      RECT 67.495 3.471 67.5 3.692 ;
      RECT 67.48 3.492 67.495 3.699 ;
      RECT 67.465 3.522 67.48 3.707 ;
      RECT 67.43 3.552 67.465 3.713 ;
      RECT 67.405 3.57 67.43 3.72 ;
      RECT 67.355 3.578 67.405 3.729 ;
      RECT 67.33 3.583 67.355 3.738 ;
      RECT 67.275 3.589 67.33 3.748 ;
      RECT 67.27 3.594 67.275 3.756 ;
      RECT 67.256 3.597 67.27 3.758 ;
      RECT 67.17 3.609 67.256 3.77 ;
      RECT 67.16 3.621 67.17 3.783 ;
      RECT 67.075 3.634 67.16 3.795 ;
      RECT 67.031 3.651 67.075 3.809 ;
      RECT 66.945 3.668 67.031 3.825 ;
      RECT 66.915 3.682 66.945 3.839 ;
      RECT 66.905 3.687 66.915 3.844 ;
      RECT 66.845 3.69 66.905 3.853 ;
      RECT 69.735 3.96 69.995 4.22 ;
      RECT 69.735 3.96 70.015 4.073 ;
      RECT 69.735 3.96 70.04 4.04 ;
      RECT 69.735 3.96 70.045 4.02 ;
      RECT 69.785 3.735 70.065 4.015 ;
      RECT 69.34 4.47 69.6 4.73 ;
      RECT 69.33 4.327 69.525 4.668 ;
      RECT 69.325 4.435 69.54 4.66 ;
      RECT 69.32 4.485 69.6 4.65 ;
      RECT 69.31 4.562 69.6 4.635 ;
      RECT 69.33 4.41 69.54 4.668 ;
      RECT 69.34 4.285 69.525 4.73 ;
      RECT 69.34 4.18 69.505 4.73 ;
      RECT 69.35 4.167 69.505 4.73 ;
      RECT 69.35 4.125 69.495 4.73 ;
      RECT 69.355 4.05 69.495 4.73 ;
      RECT 69.385 3.7 69.495 4.73 ;
      RECT 69.39 3.43 69.515 4.053 ;
      RECT 69.36 4.005 69.515 4.053 ;
      RECT 69.375 3.807 69.495 4.73 ;
      RECT 69.365 3.917 69.515 4.053 ;
      RECT 69.39 3.43 69.53 3.91 ;
      RECT 69.39 3.43 69.55 3.785 ;
      RECT 69.355 3.43 69.615 3.69 ;
      RECT 68.825 3.735 69.105 4.015 ;
      RECT 68.81 3.735 69.105 3.995 ;
      RECT 66.865 4.6 67.125 4.86 ;
      RECT 68.65 4.455 68.91 4.715 ;
      RECT 68.63 4.475 68.91 4.69 ;
      RECT 68.587 4.475 68.63 4.689 ;
      RECT 68.501 4.476 68.587 4.686 ;
      RECT 68.415 4.477 68.501 4.682 ;
      RECT 68.34 4.479 68.415 4.679 ;
      RECT 68.317 4.48 68.34 4.677 ;
      RECT 68.231 4.481 68.317 4.675 ;
      RECT 68.145 4.482 68.231 4.672 ;
      RECT 68.121 4.483 68.145 4.67 ;
      RECT 68.035 4.485 68.121 4.667 ;
      RECT 67.95 4.487 68.035 4.668 ;
      RECT 67.893 4.488 67.95 4.674 ;
      RECT 67.807 4.49 67.893 4.684 ;
      RECT 67.721 4.493 67.807 4.697 ;
      RECT 67.635 4.495 67.721 4.709 ;
      RECT 67.621 4.496 67.635 4.716 ;
      RECT 67.535 4.497 67.621 4.724 ;
      RECT 67.495 4.499 67.535 4.733 ;
      RECT 67.486 4.5 67.495 4.736 ;
      RECT 67.4 4.508 67.486 4.742 ;
      RECT 67.38 4.517 67.4 4.75 ;
      RECT 67.295 4.532 67.38 4.758 ;
      RECT 67.235 4.555 67.295 4.769 ;
      RECT 67.225 4.567 67.235 4.774 ;
      RECT 67.185 4.577 67.225 4.778 ;
      RECT 67.13 4.594 67.185 4.786 ;
      RECT 67.125 4.604 67.13 4.79 ;
      RECT 68.191 3.735 68.25 4.132 ;
      RECT 68.105 3.735 68.31 4.123 ;
      RECT 68.1 3.765 68.31 4.118 ;
      RECT 68.066 3.765 68.31 4.116 ;
      RECT 67.98 3.765 68.31 4.11 ;
      RECT 67.935 3.765 68.33 4.088 ;
      RECT 67.935 3.765 68.35 4.043 ;
      RECT 67.895 3.765 68.35 4.033 ;
      RECT 68.105 3.735 68.385 4.015 ;
      RECT 67.84 3.735 68.1 3.995 ;
      RECT 67.025 3.215 67.285 3.475 ;
      RECT 67.105 3.175 67.385 3.455 ;
      RECT 61.47 8.505 61.79 8.83 ;
      RECT 61.5 7.98 61.67 8.83 ;
      RECT 61.5 7.98 61.675 8.33 ;
      RECT 61.5 7.98 62.475 8.155 ;
      RECT 62.3 3.26 62.475 8.155 ;
      RECT 62.245 3.26 62.595 3.61 ;
      RECT 62.27 8.94 62.595 9.265 ;
      RECT 61.155 9.03 62.595 9.2 ;
      RECT 61.155 3.69 61.315 9.2 ;
      RECT 61.47 3.66 61.79 3.98 ;
      RECT 61.155 3.69 61.79 3.86 ;
      RECT 49.88 4.295 50.16 4.575 ;
      RECT 49.85 4.295 50.16 4.56 ;
      RECT 49.845 4.295 50.16 4.558 ;
      RECT 49.84 2.625 50.01 4.552 ;
      RECT 49.835 4.262 50.105 4.545 ;
      RECT 49.83 4.295 50.16 4.538 ;
      RECT 49.8 4.265 50.105 4.525 ;
      RECT 49.8 4.292 50.125 4.525 ;
      RECT 49.8 4.282 50.12 4.525 ;
      RECT 49.8 4.267 50.115 4.525 ;
      RECT 49.84 4.257 50.105 4.552 ;
      RECT 49.84 4.252 50.095 4.552 ;
      RECT 49.84 4.251 50.08 4.552 ;
      RECT 59.81 2.635 60.16 2.985 ;
      RECT 59.805 2.635 60.16 2.89 ;
      RECT 49.84 2.625 60.05 2.795 ;
      RECT 59.485 4.145 59.855 4.515 ;
      RECT 59.57 3.53 59.74 4.515 ;
      RECT 55.59 3.75 55.825 4.01 ;
      RECT 58.735 3.53 58.9 3.79 ;
      RECT 58.64 3.52 58.655 3.79 ;
      RECT 58.735 3.53 59.74 3.71 ;
      RECT 57.24 3.09 57.28 3.23 ;
      RECT 58.655 3.525 58.735 3.79 ;
      RECT 58.6 3.52 58.64 3.756 ;
      RECT 58.586 3.52 58.6 3.756 ;
      RECT 58.5 3.525 58.586 3.758 ;
      RECT 58.455 3.532 58.5 3.76 ;
      RECT 58.425 3.532 58.455 3.762 ;
      RECT 58.4 3.527 58.425 3.764 ;
      RECT 58.37 3.523 58.4 3.773 ;
      RECT 58.36 3.52 58.37 3.785 ;
      RECT 58.355 3.52 58.36 3.793 ;
      RECT 58.35 3.52 58.355 3.798 ;
      RECT 58.34 3.519 58.35 3.808 ;
      RECT 58.335 3.518 58.34 3.818 ;
      RECT 58.32 3.517 58.335 3.823 ;
      RECT 58.292 3.514 58.32 3.85 ;
      RECT 58.206 3.506 58.292 3.85 ;
      RECT 58.12 3.495 58.206 3.85 ;
      RECT 58.08 3.48 58.12 3.85 ;
      RECT 58.04 3.454 58.08 3.85 ;
      RECT 58.035 3.436 58.04 3.662 ;
      RECT 58.025 3.432 58.035 3.652 ;
      RECT 58.01 3.422 58.025 3.639 ;
      RECT 57.99 3.406 58.01 3.624 ;
      RECT 57.975 3.391 57.99 3.609 ;
      RECT 57.965 3.38 57.975 3.599 ;
      RECT 57.94 3.364 57.965 3.588 ;
      RECT 57.935 3.351 57.94 3.578 ;
      RECT 57.93 3.347 57.935 3.573 ;
      RECT 57.875 3.333 57.93 3.551 ;
      RECT 57.836 3.314 57.875 3.515 ;
      RECT 57.75 3.288 57.836 3.468 ;
      RECT 57.746 3.27 57.75 3.434 ;
      RECT 57.66 3.251 57.746 3.412 ;
      RECT 57.655 3.233 57.66 3.39 ;
      RECT 57.65 3.231 57.655 3.388 ;
      RECT 57.64 3.23 57.65 3.383 ;
      RECT 57.58 3.217 57.64 3.369 ;
      RECT 57.535 3.195 57.58 3.348 ;
      RECT 57.475 3.172 57.535 3.327 ;
      RECT 57.411 3.147 57.475 3.302 ;
      RECT 57.325 3.117 57.411 3.271 ;
      RECT 57.31 3.097 57.325 3.25 ;
      RECT 57.28 3.092 57.31 3.241 ;
      RECT 57.227 3.09 57.24 3.23 ;
      RECT 57.141 3.09 57.227 3.232 ;
      RECT 57.055 3.09 57.141 3.234 ;
      RECT 57.035 3.09 57.055 3.238 ;
      RECT 56.99 3.092 57.035 3.249 ;
      RECT 56.95 3.102 56.99 3.265 ;
      RECT 56.946 3.111 56.95 3.273 ;
      RECT 56.86 3.131 56.946 3.289 ;
      RECT 56.85 3.15 56.86 3.307 ;
      RECT 56.845 3.152 56.85 3.31 ;
      RECT 56.835 3.156 56.845 3.313 ;
      RECT 56.815 3.161 56.835 3.323 ;
      RECT 56.785 3.171 56.815 3.343 ;
      RECT 56.78 3.178 56.785 3.357 ;
      RECT 56.77 3.182 56.78 3.364 ;
      RECT 56.755 3.19 56.77 3.375 ;
      RECT 56.745 3.2 56.755 3.386 ;
      RECT 56.735 3.207 56.745 3.394 ;
      RECT 56.71 3.22 56.735 3.409 ;
      RECT 56.646 3.256 56.71 3.448 ;
      RECT 56.56 3.319 56.646 3.512 ;
      RECT 56.525 3.37 56.56 3.565 ;
      RECT 56.52 3.387 56.525 3.582 ;
      RECT 56.505 3.396 56.52 3.589 ;
      RECT 56.485 3.411 56.505 3.603 ;
      RECT 56.48 3.422 56.485 3.613 ;
      RECT 56.46 3.435 56.48 3.623 ;
      RECT 56.455 3.445 56.46 3.633 ;
      RECT 56.44 3.45 56.455 3.642 ;
      RECT 56.43 3.46 56.44 3.653 ;
      RECT 56.4 3.477 56.43 3.67 ;
      RECT 56.39 3.495 56.4 3.688 ;
      RECT 56.375 3.506 56.39 3.699 ;
      RECT 56.335 3.53 56.375 3.715 ;
      RECT 56.3 3.564 56.335 3.732 ;
      RECT 56.27 3.587 56.3 3.744 ;
      RECT 56.255 3.597 56.27 3.753 ;
      RECT 56.215 3.607 56.255 3.764 ;
      RECT 56.195 3.618 56.215 3.776 ;
      RECT 56.19 3.622 56.195 3.783 ;
      RECT 56.175 3.626 56.19 3.788 ;
      RECT 56.165 3.631 56.175 3.793 ;
      RECT 56.16 3.634 56.165 3.796 ;
      RECT 56.13 3.64 56.16 3.803 ;
      RECT 56.095 3.65 56.13 3.817 ;
      RECT 56.035 3.665 56.095 3.837 ;
      RECT 55.98 3.685 56.035 3.861 ;
      RECT 55.951 3.7 55.98 3.879 ;
      RECT 55.865 3.72 55.951 3.904 ;
      RECT 55.86 3.735 55.865 3.924 ;
      RECT 55.85 3.738 55.86 3.925 ;
      RECT 55.825 3.745 55.85 4.01 ;
      RECT 48.875 8.945 49.225 9.295 ;
      RECT 57.7 8.9 58.05 9.25 ;
      RECT 48.875 8.975 58.05 9.175 ;
      RECT 56.24 4.98 56.25 5.17 ;
      RECT 54.5 4.855 54.78 5.135 ;
      RECT 57.545 3.795 57.55 4.28 ;
      RECT 57.44 3.795 57.5 4.055 ;
      RECT 57.765 4.765 57.77 4.84 ;
      RECT 57.755 4.632 57.765 4.875 ;
      RECT 57.745 4.467 57.755 4.896 ;
      RECT 57.74 4.337 57.745 4.912 ;
      RECT 57.73 4.227 57.74 4.928 ;
      RECT 57.725 4.126 57.73 4.945 ;
      RECT 57.72 4.108 57.725 4.955 ;
      RECT 57.715 4.09 57.72 4.965 ;
      RECT 57.705 4.065 57.715 4.98 ;
      RECT 57.7 4.045 57.705 4.995 ;
      RECT 57.68 3.795 57.7 5.02 ;
      RECT 57.665 3.795 57.68 5.053 ;
      RECT 57.635 3.795 57.665 5.075 ;
      RECT 57.615 3.795 57.635 5.089 ;
      RECT 57.595 3.795 57.615 4.605 ;
      RECT 57.61 4.672 57.615 5.094 ;
      RECT 57.605 4.702 57.61 5.096 ;
      RECT 57.6 4.715 57.605 5.099 ;
      RECT 57.595 4.725 57.6 5.103 ;
      RECT 57.59 3.795 57.595 4.523 ;
      RECT 57.59 4.735 57.595 5.105 ;
      RECT 57.585 3.795 57.59 4.5 ;
      RECT 57.575 4.757 57.59 5.105 ;
      RECT 57.57 3.795 57.585 4.445 ;
      RECT 57.565 4.782 57.575 5.105 ;
      RECT 57.565 3.795 57.57 4.39 ;
      RECT 57.555 3.795 57.565 4.338 ;
      RECT 57.56 4.795 57.565 5.106 ;
      RECT 57.555 4.807 57.56 5.107 ;
      RECT 57.55 3.795 57.555 4.298 ;
      RECT 57.55 4.82 57.555 5.108 ;
      RECT 57.535 4.835 57.55 5.109 ;
      RECT 57.54 3.795 57.545 4.26 ;
      RECT 57.535 3.795 57.54 4.225 ;
      RECT 57.53 3.795 57.535 4.2 ;
      RECT 57.525 4.862 57.535 5.111 ;
      RECT 57.52 3.795 57.53 4.158 ;
      RECT 57.52 4.88 57.525 5.112 ;
      RECT 57.515 3.795 57.52 4.118 ;
      RECT 57.515 4.887 57.52 5.113 ;
      RECT 57.51 3.795 57.515 4.09 ;
      RECT 57.505 4.905 57.515 5.114 ;
      RECT 57.5 3.795 57.51 4.07 ;
      RECT 57.495 4.925 57.505 5.116 ;
      RECT 57.485 4.942 57.495 5.117 ;
      RECT 57.45 4.965 57.485 5.12 ;
      RECT 57.395 4.983 57.45 5.126 ;
      RECT 57.309 4.991 57.395 5.135 ;
      RECT 57.223 5.002 57.309 5.146 ;
      RECT 57.137 5.012 57.223 5.157 ;
      RECT 57.051 5.022 57.137 5.169 ;
      RECT 56.965 5.032 57.051 5.18 ;
      RECT 56.945 5.038 56.965 5.186 ;
      RECT 56.865 5.04 56.945 5.19 ;
      RECT 56.86 5.039 56.865 5.195 ;
      RECT 56.852 5.038 56.86 5.195 ;
      RECT 56.766 5.034 56.852 5.193 ;
      RECT 56.68 5.026 56.766 5.19 ;
      RECT 56.594 5.017 56.68 5.186 ;
      RECT 56.508 5.009 56.594 5.183 ;
      RECT 56.422 5.001 56.508 5.179 ;
      RECT 56.336 4.992 56.422 5.176 ;
      RECT 56.25 4.984 56.336 5.172 ;
      RECT 56.195 4.977 56.24 5.17 ;
      RECT 56.11 4.97 56.195 5.168 ;
      RECT 56.036 4.962 56.11 5.164 ;
      RECT 55.95 4.954 56.036 5.161 ;
      RECT 55.947 4.95 55.95 5.159 ;
      RECT 55.861 4.946 55.947 5.158 ;
      RECT 55.775 4.938 55.861 5.155 ;
      RECT 55.69 4.933 55.775 5.152 ;
      RECT 55.604 4.93 55.69 5.149 ;
      RECT 55.518 4.928 55.604 5.146 ;
      RECT 55.432 4.925 55.518 5.143 ;
      RECT 55.346 4.922 55.432 5.14 ;
      RECT 55.26 4.919 55.346 5.137 ;
      RECT 55.184 4.917 55.26 5.134 ;
      RECT 55.098 4.914 55.184 5.131 ;
      RECT 55.012 4.911 55.098 5.129 ;
      RECT 54.926 4.909 55.012 5.126 ;
      RECT 54.84 4.906 54.926 5.123 ;
      RECT 54.78 4.897 54.84 5.121 ;
      RECT 57.29 4.515 57.365 4.775 ;
      RECT 57.27 4.495 57.275 4.775 ;
      RECT 56.59 4.28 56.695 4.575 ;
      RECT 51.035 4.255 51.105 4.515 ;
      RECT 56.93 4.13 56.935 4.501 ;
      RECT 56.92 4.185 56.925 4.501 ;
      RECT 57.225 3.355 57.285 3.615 ;
      RECT 57.28 4.51 57.29 4.775 ;
      RECT 57.275 4.5 57.28 4.775 ;
      RECT 57.195 4.447 57.27 4.775 ;
      RECT 57.22 3.355 57.225 3.635 ;
      RECT 57.21 3.355 57.22 3.655 ;
      RECT 57.195 3.355 57.21 3.685 ;
      RECT 57.18 3.355 57.195 3.728 ;
      RECT 57.175 4.39 57.195 4.775 ;
      RECT 57.165 3.355 57.18 3.765 ;
      RECT 57.16 4.37 57.175 4.775 ;
      RECT 57.16 3.355 57.165 3.788 ;
      RECT 57.15 3.355 57.16 3.813 ;
      RECT 57.12 4.337 57.16 4.775 ;
      RECT 57.125 3.355 57.15 3.863 ;
      RECT 57.12 3.355 57.125 3.918 ;
      RECT 57.115 3.355 57.12 3.96 ;
      RECT 57.105 4.3 57.12 4.775 ;
      RECT 57.11 3.355 57.115 4.003 ;
      RECT 57.105 3.355 57.11 4.068 ;
      RECT 57.1 3.355 57.105 4.09 ;
      RECT 57.1 4.288 57.105 4.64 ;
      RECT 57.095 3.355 57.1 4.158 ;
      RECT 57.095 4.28 57.1 4.623 ;
      RECT 57.09 3.355 57.095 4.203 ;
      RECT 57.085 4.262 57.095 4.6 ;
      RECT 57.085 3.355 57.09 4.24 ;
      RECT 57.075 3.355 57.085 4.58 ;
      RECT 57.07 3.355 57.075 4.563 ;
      RECT 57.065 3.355 57.07 4.548 ;
      RECT 57.06 3.355 57.065 4.533 ;
      RECT 57.04 3.355 57.06 4.523 ;
      RECT 57.035 3.355 57.04 4.513 ;
      RECT 57.025 3.355 57.035 4.509 ;
      RECT 57.02 3.632 57.025 4.508 ;
      RECT 57.015 3.655 57.02 4.507 ;
      RECT 57.01 3.685 57.015 4.506 ;
      RECT 57.005 3.712 57.01 4.505 ;
      RECT 57 3.74 57.005 4.505 ;
      RECT 56.995 3.767 57 4.505 ;
      RECT 56.99 3.787 56.995 4.505 ;
      RECT 56.985 3.815 56.99 4.505 ;
      RECT 56.975 3.857 56.985 4.505 ;
      RECT 56.965 3.902 56.975 4.504 ;
      RECT 56.96 3.955 56.965 4.503 ;
      RECT 56.955 3.987 56.96 4.502 ;
      RECT 56.95 4.007 56.955 4.501 ;
      RECT 56.945 4.045 56.95 4.501 ;
      RECT 56.94 4.067 56.945 4.501 ;
      RECT 56.935 4.092 56.94 4.501 ;
      RECT 56.925 4.157 56.93 4.501 ;
      RECT 56.91 4.217 56.92 4.501 ;
      RECT 56.895 4.227 56.91 4.501 ;
      RECT 56.875 4.237 56.895 4.501 ;
      RECT 56.845 4.242 56.875 4.498 ;
      RECT 56.785 4.252 56.845 4.495 ;
      RECT 56.765 4.261 56.785 4.5 ;
      RECT 56.74 4.267 56.765 4.513 ;
      RECT 56.72 4.272 56.74 4.528 ;
      RECT 56.695 4.277 56.72 4.575 ;
      RECT 56.566 4.279 56.59 4.575 ;
      RECT 56.48 4.274 56.566 4.575 ;
      RECT 56.44 4.271 56.48 4.575 ;
      RECT 56.39 4.273 56.44 4.555 ;
      RECT 56.36 4.277 56.39 4.555 ;
      RECT 56.281 4.287 56.36 4.555 ;
      RECT 56.195 4.302 56.281 4.556 ;
      RECT 56.145 4.312 56.195 4.557 ;
      RECT 56.137 4.315 56.145 4.557 ;
      RECT 56.051 4.317 56.137 4.558 ;
      RECT 55.965 4.321 56.051 4.558 ;
      RECT 55.879 4.325 55.965 4.559 ;
      RECT 55.793 4.328 55.879 4.56 ;
      RECT 55.707 4.332 55.793 4.56 ;
      RECT 55.621 4.336 55.707 4.561 ;
      RECT 55.535 4.339 55.621 4.562 ;
      RECT 55.449 4.343 55.535 4.562 ;
      RECT 55.363 4.347 55.449 4.563 ;
      RECT 55.277 4.351 55.363 4.564 ;
      RECT 55.191 4.354 55.277 4.564 ;
      RECT 55.105 4.358 55.191 4.565 ;
      RECT 55.075 4.36 55.105 4.565 ;
      RECT 54.989 4.363 55.075 4.566 ;
      RECT 54.903 4.367 54.989 4.567 ;
      RECT 54.817 4.371 54.903 4.568 ;
      RECT 54.731 4.374 54.817 4.568 ;
      RECT 54.645 4.378 54.731 4.569 ;
      RECT 54.61 4.383 54.645 4.57 ;
      RECT 54.555 4.393 54.61 4.577 ;
      RECT 54.53 4.405 54.555 4.587 ;
      RECT 54.495 4.418 54.53 4.595 ;
      RECT 54.455 4.435 54.495 4.618 ;
      RECT 54.435 4.448 54.455 4.645 ;
      RECT 54.405 4.46 54.435 4.673 ;
      RECT 54.4 4.468 54.405 4.693 ;
      RECT 54.395 4.471 54.4 4.703 ;
      RECT 54.345 4.483 54.395 4.737 ;
      RECT 54.335 4.498 54.345 4.77 ;
      RECT 54.325 4.504 54.335 4.783 ;
      RECT 54.315 4.511 54.325 4.795 ;
      RECT 54.29 4.524 54.315 4.813 ;
      RECT 54.275 4.539 54.29 4.835 ;
      RECT 54.265 4.547 54.275 4.851 ;
      RECT 54.25 4.556 54.265 4.866 ;
      RECT 54.24 4.566 54.25 4.88 ;
      RECT 54.221 4.579 54.24 4.897 ;
      RECT 54.135 4.624 54.221 4.962 ;
      RECT 54.12 4.669 54.135 5.02 ;
      RECT 54.115 4.678 54.12 5.033 ;
      RECT 54.105 4.685 54.115 5.038 ;
      RECT 54.1 4.69 54.105 5.042 ;
      RECT 54.08 4.7 54.1 5.049 ;
      RECT 54.055 4.72 54.08 5.063 ;
      RECT 54.02 4.745 54.055 5.083 ;
      RECT 54.005 4.768 54.02 5.098 ;
      RECT 53.995 4.778 54.005 5.103 ;
      RECT 53.985 4.786 53.995 5.11 ;
      RECT 53.975 4.795 53.985 5.116 ;
      RECT 53.955 4.807 53.975 5.118 ;
      RECT 53.945 4.82 53.955 5.12 ;
      RECT 53.92 4.835 53.945 5.123 ;
      RECT 53.9 4.852 53.92 5.127 ;
      RECT 53.86 4.88 53.9 5.133 ;
      RECT 53.795 4.927 53.86 5.142 ;
      RECT 53.78 4.96 53.795 5.15 ;
      RECT 53.775 4.967 53.78 5.152 ;
      RECT 53.725 4.992 53.775 5.157 ;
      RECT 53.71 5.016 53.725 5.164 ;
      RECT 53.66 5.021 53.71 5.165 ;
      RECT 53.574 5.025 53.66 5.165 ;
      RECT 53.488 5.025 53.574 5.165 ;
      RECT 53.402 5.025 53.488 5.166 ;
      RECT 53.316 5.025 53.402 5.166 ;
      RECT 53.23 5.025 53.316 5.166 ;
      RECT 53.164 5.025 53.23 5.166 ;
      RECT 53.078 5.025 53.164 5.167 ;
      RECT 52.992 5.025 53.078 5.167 ;
      RECT 52.906 5.026 52.992 5.168 ;
      RECT 52.82 5.026 52.906 5.168 ;
      RECT 52.734 5.026 52.82 5.168 ;
      RECT 52.648 5.026 52.734 5.169 ;
      RECT 52.562 5.026 52.648 5.169 ;
      RECT 52.476 5.027 52.562 5.17 ;
      RECT 52.39 5.027 52.476 5.17 ;
      RECT 52.37 5.027 52.39 5.17 ;
      RECT 52.284 5.027 52.37 5.17 ;
      RECT 52.198 5.027 52.284 5.17 ;
      RECT 52.112 5.028 52.198 5.17 ;
      RECT 52.026 5.028 52.112 5.17 ;
      RECT 51.94 5.028 52.026 5.17 ;
      RECT 51.854 5.029 51.94 5.17 ;
      RECT 51.768 5.029 51.854 5.17 ;
      RECT 51.682 5.029 51.768 5.17 ;
      RECT 51.596 5.029 51.682 5.17 ;
      RECT 51.51 5.03 51.596 5.17 ;
      RECT 51.46 5.027 51.51 5.17 ;
      RECT 51.45 5.025 51.46 5.169 ;
      RECT 51.446 5.025 51.45 5.168 ;
      RECT 51.36 5.02 51.446 5.163 ;
      RECT 51.338 5.013 51.36 5.157 ;
      RECT 51.252 5.004 51.338 5.151 ;
      RECT 51.166 4.991 51.252 5.142 ;
      RECT 51.08 4.977 51.166 5.132 ;
      RECT 51.035 4.967 51.08 5.125 ;
      RECT 51.015 4.255 51.035 4.533 ;
      RECT 51.015 4.96 51.035 5.121 ;
      RECT 50.985 4.255 51.015 4.555 ;
      RECT 50.975 4.927 51.015 5.118 ;
      RECT 50.97 4.255 50.985 4.575 ;
      RECT 50.97 4.892 50.975 5.116 ;
      RECT 50.965 4.255 50.97 4.7 ;
      RECT 50.965 4.852 50.97 5.116 ;
      RECT 50.955 4.255 50.965 5.116 ;
      RECT 50.88 4.255 50.955 5.11 ;
      RECT 50.85 4.255 50.88 5.1 ;
      RECT 50.845 4.255 50.85 5.092 ;
      RECT 50.84 4.297 50.845 5.085 ;
      RECT 50.83 4.366 50.84 5.076 ;
      RECT 50.825 4.436 50.83 5.028 ;
      RECT 50.82 4.5 50.825 4.925 ;
      RECT 50.815 4.535 50.82 4.88 ;
      RECT 50.813 4.572 50.815 4.772 ;
      RECT 50.81 4.58 50.813 4.765 ;
      RECT 50.805 4.645 50.81 4.708 ;
      RECT 54.88 3.735 55.16 4.015 ;
      RECT 54.87 3.735 55.16 3.878 ;
      RECT 54.825 3.6 55.085 3.86 ;
      RECT 54.825 3.715 55.14 3.86 ;
      RECT 54.825 3.685 55.135 3.86 ;
      RECT 54.825 3.672 55.125 3.86 ;
      RECT 54.825 3.662 55.12 3.86 ;
      RECT 50.8 3.645 51.06 3.905 ;
      RECT 54.57 3.195 54.83 3.455 ;
      RECT 54.56 3.22 54.83 3.415 ;
      RECT 54.555 3.22 54.56 3.414 ;
      RECT 54.485 3.215 54.555 3.406 ;
      RECT 54.4 3.202 54.485 3.389 ;
      RECT 54.396 3.194 54.4 3.379 ;
      RECT 54.31 3.187 54.396 3.369 ;
      RECT 54.301 3.179 54.31 3.359 ;
      RECT 54.215 3.172 54.301 3.347 ;
      RECT 54.195 3.163 54.215 3.333 ;
      RECT 54.14 3.158 54.195 3.325 ;
      RECT 54.13 3.152 54.14 3.319 ;
      RECT 54.11 3.15 54.13 3.315 ;
      RECT 54.102 3.149 54.11 3.311 ;
      RECT 54.016 3.141 54.102 3.3 ;
      RECT 53.93 3.127 54.016 3.28 ;
      RECT 53.87 3.115 53.93 3.265 ;
      RECT 53.86 3.11 53.87 3.26 ;
      RECT 53.81 3.11 53.86 3.262 ;
      RECT 53.763 3.112 53.81 3.266 ;
      RECT 53.677 3.119 53.763 3.271 ;
      RECT 53.591 3.127 53.677 3.277 ;
      RECT 53.505 3.136 53.591 3.283 ;
      RECT 53.446 3.142 53.505 3.288 ;
      RECT 53.36 3.147 53.446 3.294 ;
      RECT 53.285 3.152 53.36 3.3 ;
      RECT 53.246 3.154 53.285 3.305 ;
      RECT 53.16 3.151 53.246 3.31 ;
      RECT 53.075 3.149 53.16 3.317 ;
      RECT 53.043 3.148 53.075 3.32 ;
      RECT 52.957 3.147 53.043 3.321 ;
      RECT 52.871 3.146 52.957 3.322 ;
      RECT 52.785 3.145 52.871 3.322 ;
      RECT 52.699 3.144 52.785 3.323 ;
      RECT 52.613 3.143 52.699 3.324 ;
      RECT 52.527 3.142 52.613 3.325 ;
      RECT 52.441 3.141 52.527 3.325 ;
      RECT 52.355 3.14 52.441 3.326 ;
      RECT 52.305 3.14 52.355 3.327 ;
      RECT 52.291 3.141 52.305 3.327 ;
      RECT 52.205 3.148 52.291 3.328 ;
      RECT 52.131 3.159 52.205 3.329 ;
      RECT 52.045 3.168 52.131 3.33 ;
      RECT 52.01 3.175 52.045 3.345 ;
      RECT 51.985 3.178 52.01 3.375 ;
      RECT 51.96 3.187 51.985 3.404 ;
      RECT 51.95 3.198 51.96 3.424 ;
      RECT 51.94 3.206 51.95 3.438 ;
      RECT 51.935 3.212 51.94 3.448 ;
      RECT 51.91 3.229 51.935 3.465 ;
      RECT 51.895 3.251 51.91 3.493 ;
      RECT 51.865 3.277 51.895 3.523 ;
      RECT 51.845 3.306 51.865 3.553 ;
      RECT 51.84 3.321 51.845 3.57 ;
      RECT 51.82 3.336 51.84 3.585 ;
      RECT 51.81 3.354 51.82 3.603 ;
      RECT 51.8 3.365 51.81 3.618 ;
      RECT 51.75 3.397 51.8 3.644 ;
      RECT 51.745 3.427 51.75 3.664 ;
      RECT 51.735 3.44 51.745 3.67 ;
      RECT 51.726 3.45 51.735 3.678 ;
      RECT 51.715 3.461 51.726 3.686 ;
      RECT 51.71 3.471 51.715 3.692 ;
      RECT 51.695 3.492 51.71 3.699 ;
      RECT 51.68 3.522 51.695 3.707 ;
      RECT 51.645 3.552 51.68 3.713 ;
      RECT 51.62 3.57 51.645 3.72 ;
      RECT 51.57 3.578 51.62 3.729 ;
      RECT 51.545 3.583 51.57 3.738 ;
      RECT 51.49 3.589 51.545 3.748 ;
      RECT 51.485 3.594 51.49 3.756 ;
      RECT 51.471 3.597 51.485 3.758 ;
      RECT 51.385 3.609 51.471 3.77 ;
      RECT 51.375 3.621 51.385 3.783 ;
      RECT 51.29 3.634 51.375 3.795 ;
      RECT 51.246 3.651 51.29 3.809 ;
      RECT 51.16 3.668 51.246 3.825 ;
      RECT 51.13 3.682 51.16 3.839 ;
      RECT 51.12 3.687 51.13 3.844 ;
      RECT 51.06 3.69 51.12 3.853 ;
      RECT 53.95 3.96 54.21 4.22 ;
      RECT 53.95 3.96 54.23 4.073 ;
      RECT 53.95 3.96 54.255 4.04 ;
      RECT 53.95 3.96 54.26 4.02 ;
      RECT 54 3.735 54.28 4.015 ;
      RECT 53.555 4.47 53.815 4.73 ;
      RECT 53.545 4.327 53.74 4.668 ;
      RECT 53.54 4.435 53.755 4.66 ;
      RECT 53.535 4.485 53.815 4.65 ;
      RECT 53.525 4.562 53.815 4.635 ;
      RECT 53.545 4.41 53.755 4.668 ;
      RECT 53.555 4.285 53.74 4.73 ;
      RECT 53.555 4.18 53.72 4.73 ;
      RECT 53.565 4.167 53.72 4.73 ;
      RECT 53.565 4.125 53.71 4.73 ;
      RECT 53.57 4.05 53.71 4.73 ;
      RECT 53.6 3.7 53.71 4.73 ;
      RECT 53.605 3.43 53.73 4.053 ;
      RECT 53.575 4.005 53.73 4.053 ;
      RECT 53.59 3.807 53.71 4.73 ;
      RECT 53.58 3.917 53.73 4.053 ;
      RECT 53.605 3.43 53.745 3.91 ;
      RECT 53.605 3.43 53.765 3.785 ;
      RECT 53.57 3.43 53.83 3.69 ;
      RECT 53.04 3.735 53.32 4.015 ;
      RECT 53.025 3.735 53.32 3.995 ;
      RECT 51.08 4.6 51.34 4.86 ;
      RECT 52.865 4.455 53.125 4.715 ;
      RECT 52.845 4.475 53.125 4.69 ;
      RECT 52.802 4.475 52.845 4.689 ;
      RECT 52.716 4.476 52.802 4.686 ;
      RECT 52.63 4.477 52.716 4.682 ;
      RECT 52.555 4.479 52.63 4.679 ;
      RECT 52.532 4.48 52.555 4.677 ;
      RECT 52.446 4.481 52.532 4.675 ;
      RECT 52.36 4.482 52.446 4.672 ;
      RECT 52.336 4.483 52.36 4.67 ;
      RECT 52.25 4.485 52.336 4.667 ;
      RECT 52.165 4.487 52.25 4.668 ;
      RECT 52.108 4.488 52.165 4.674 ;
      RECT 52.022 4.49 52.108 4.684 ;
      RECT 51.936 4.493 52.022 4.697 ;
      RECT 51.85 4.495 51.936 4.709 ;
      RECT 51.836 4.496 51.85 4.716 ;
      RECT 51.75 4.497 51.836 4.724 ;
      RECT 51.71 4.499 51.75 4.733 ;
      RECT 51.701 4.5 51.71 4.736 ;
      RECT 51.615 4.508 51.701 4.742 ;
      RECT 51.595 4.517 51.615 4.75 ;
      RECT 51.51 4.532 51.595 4.758 ;
      RECT 51.45 4.555 51.51 4.769 ;
      RECT 51.44 4.567 51.45 4.774 ;
      RECT 51.4 4.577 51.44 4.778 ;
      RECT 51.345 4.594 51.4 4.786 ;
      RECT 51.34 4.604 51.345 4.79 ;
      RECT 52.406 3.735 52.465 4.132 ;
      RECT 52.32 3.735 52.525 4.123 ;
      RECT 52.315 3.765 52.525 4.118 ;
      RECT 52.281 3.765 52.525 4.116 ;
      RECT 52.195 3.765 52.525 4.11 ;
      RECT 52.15 3.765 52.545 4.088 ;
      RECT 52.15 3.765 52.565 4.043 ;
      RECT 52.11 3.765 52.565 4.033 ;
      RECT 52.32 3.735 52.6 4.015 ;
      RECT 52.055 3.735 52.315 3.995 ;
      RECT 51.24 3.215 51.5 3.475 ;
      RECT 51.32 3.175 51.6 3.455 ;
      RECT 45.695 8.505 46.015 8.83 ;
      RECT 45.725 7.98 45.895 8.83 ;
      RECT 45.725 7.98 45.9 8.33 ;
      RECT 45.725 7.98 46.7 8.155 ;
      RECT 46.525 3.26 46.7 8.155 ;
      RECT 46.47 3.26 46.82 3.61 ;
      RECT 46.495 8.94 46.82 9.265 ;
      RECT 45.38 9.03 46.82 9.2 ;
      RECT 45.38 3.69 45.54 9.2 ;
      RECT 45.695 3.66 46.015 3.98 ;
      RECT 45.38 3.69 46.015 3.86 ;
      RECT 34.105 4.295 34.385 4.575 ;
      RECT 34.075 4.295 34.385 4.56 ;
      RECT 34.07 4.295 34.385 4.558 ;
      RECT 34.065 2.625 34.235 4.552 ;
      RECT 34.06 4.262 34.33 4.545 ;
      RECT 34.055 4.295 34.385 4.538 ;
      RECT 34.025 4.265 34.33 4.525 ;
      RECT 34.025 4.292 34.35 4.525 ;
      RECT 34.025 4.282 34.345 4.525 ;
      RECT 34.025 4.267 34.34 4.525 ;
      RECT 34.065 4.257 34.33 4.552 ;
      RECT 34.065 4.252 34.32 4.552 ;
      RECT 34.065 4.251 34.305 4.552 ;
      RECT 44.035 2.635 44.385 2.985 ;
      RECT 44.03 2.635 44.385 2.89 ;
      RECT 34.065 2.625 44.275 2.795 ;
      RECT 43.71 4.145 44.08 4.515 ;
      RECT 43.795 3.53 43.965 4.515 ;
      RECT 39.815 3.75 40.05 4.01 ;
      RECT 42.96 3.53 43.125 3.79 ;
      RECT 42.865 3.52 42.88 3.79 ;
      RECT 42.96 3.53 43.965 3.71 ;
      RECT 41.465 3.09 41.505 3.23 ;
      RECT 42.88 3.525 42.96 3.79 ;
      RECT 42.825 3.52 42.865 3.756 ;
      RECT 42.811 3.52 42.825 3.756 ;
      RECT 42.725 3.525 42.811 3.758 ;
      RECT 42.68 3.532 42.725 3.76 ;
      RECT 42.65 3.532 42.68 3.762 ;
      RECT 42.625 3.527 42.65 3.764 ;
      RECT 42.595 3.523 42.625 3.773 ;
      RECT 42.585 3.52 42.595 3.785 ;
      RECT 42.58 3.52 42.585 3.793 ;
      RECT 42.575 3.52 42.58 3.798 ;
      RECT 42.565 3.519 42.575 3.808 ;
      RECT 42.56 3.518 42.565 3.818 ;
      RECT 42.545 3.517 42.56 3.823 ;
      RECT 42.517 3.514 42.545 3.85 ;
      RECT 42.431 3.506 42.517 3.85 ;
      RECT 42.345 3.495 42.431 3.85 ;
      RECT 42.305 3.48 42.345 3.85 ;
      RECT 42.265 3.454 42.305 3.85 ;
      RECT 42.26 3.436 42.265 3.662 ;
      RECT 42.25 3.432 42.26 3.652 ;
      RECT 42.235 3.422 42.25 3.639 ;
      RECT 42.215 3.406 42.235 3.624 ;
      RECT 42.2 3.391 42.215 3.609 ;
      RECT 42.19 3.38 42.2 3.599 ;
      RECT 42.165 3.364 42.19 3.588 ;
      RECT 42.16 3.351 42.165 3.578 ;
      RECT 42.155 3.347 42.16 3.573 ;
      RECT 42.1 3.333 42.155 3.551 ;
      RECT 42.061 3.314 42.1 3.515 ;
      RECT 41.975 3.288 42.061 3.468 ;
      RECT 41.971 3.27 41.975 3.434 ;
      RECT 41.885 3.251 41.971 3.412 ;
      RECT 41.88 3.233 41.885 3.39 ;
      RECT 41.875 3.231 41.88 3.388 ;
      RECT 41.865 3.23 41.875 3.383 ;
      RECT 41.805 3.217 41.865 3.369 ;
      RECT 41.76 3.195 41.805 3.348 ;
      RECT 41.7 3.172 41.76 3.327 ;
      RECT 41.636 3.147 41.7 3.302 ;
      RECT 41.55 3.117 41.636 3.271 ;
      RECT 41.535 3.097 41.55 3.25 ;
      RECT 41.505 3.092 41.535 3.241 ;
      RECT 41.452 3.09 41.465 3.23 ;
      RECT 41.366 3.09 41.452 3.232 ;
      RECT 41.28 3.09 41.366 3.234 ;
      RECT 41.26 3.09 41.28 3.238 ;
      RECT 41.215 3.092 41.26 3.249 ;
      RECT 41.175 3.102 41.215 3.265 ;
      RECT 41.171 3.111 41.175 3.273 ;
      RECT 41.085 3.131 41.171 3.289 ;
      RECT 41.075 3.15 41.085 3.307 ;
      RECT 41.07 3.152 41.075 3.31 ;
      RECT 41.06 3.156 41.07 3.313 ;
      RECT 41.04 3.161 41.06 3.323 ;
      RECT 41.01 3.171 41.04 3.343 ;
      RECT 41.005 3.178 41.01 3.357 ;
      RECT 40.995 3.182 41.005 3.364 ;
      RECT 40.98 3.19 40.995 3.375 ;
      RECT 40.97 3.2 40.98 3.386 ;
      RECT 40.96 3.207 40.97 3.394 ;
      RECT 40.935 3.22 40.96 3.409 ;
      RECT 40.871 3.256 40.935 3.448 ;
      RECT 40.785 3.319 40.871 3.512 ;
      RECT 40.75 3.37 40.785 3.565 ;
      RECT 40.745 3.387 40.75 3.582 ;
      RECT 40.73 3.396 40.745 3.589 ;
      RECT 40.71 3.411 40.73 3.603 ;
      RECT 40.705 3.422 40.71 3.613 ;
      RECT 40.685 3.435 40.705 3.623 ;
      RECT 40.68 3.445 40.685 3.633 ;
      RECT 40.665 3.45 40.68 3.642 ;
      RECT 40.655 3.46 40.665 3.653 ;
      RECT 40.625 3.477 40.655 3.67 ;
      RECT 40.615 3.495 40.625 3.688 ;
      RECT 40.6 3.506 40.615 3.699 ;
      RECT 40.56 3.53 40.6 3.715 ;
      RECT 40.525 3.564 40.56 3.732 ;
      RECT 40.495 3.587 40.525 3.744 ;
      RECT 40.48 3.597 40.495 3.753 ;
      RECT 40.44 3.607 40.48 3.764 ;
      RECT 40.42 3.618 40.44 3.776 ;
      RECT 40.415 3.622 40.42 3.783 ;
      RECT 40.4 3.626 40.415 3.788 ;
      RECT 40.39 3.631 40.4 3.793 ;
      RECT 40.385 3.634 40.39 3.796 ;
      RECT 40.355 3.64 40.385 3.803 ;
      RECT 40.32 3.65 40.355 3.817 ;
      RECT 40.26 3.665 40.32 3.837 ;
      RECT 40.205 3.685 40.26 3.861 ;
      RECT 40.176 3.7 40.205 3.879 ;
      RECT 40.09 3.72 40.176 3.904 ;
      RECT 40.085 3.735 40.09 3.924 ;
      RECT 40.075 3.738 40.085 3.925 ;
      RECT 40.05 3.745 40.075 4.01 ;
      RECT 33.095 8.945 33.445 9.295 ;
      RECT 41.92 8.9 42.27 9.25 ;
      RECT 33.095 8.975 42.27 9.175 ;
      RECT 40.465 4.98 40.475 5.17 ;
      RECT 38.725 4.855 39.005 5.135 ;
      RECT 41.77 3.795 41.775 4.28 ;
      RECT 41.665 3.795 41.725 4.055 ;
      RECT 41.99 4.765 41.995 4.84 ;
      RECT 41.98 4.632 41.99 4.875 ;
      RECT 41.97 4.467 41.98 4.896 ;
      RECT 41.965 4.337 41.97 4.912 ;
      RECT 41.955 4.227 41.965 4.928 ;
      RECT 41.95 4.126 41.955 4.945 ;
      RECT 41.945 4.108 41.95 4.955 ;
      RECT 41.94 4.09 41.945 4.965 ;
      RECT 41.93 4.065 41.94 4.98 ;
      RECT 41.925 4.045 41.93 4.995 ;
      RECT 41.905 3.795 41.925 5.02 ;
      RECT 41.89 3.795 41.905 5.053 ;
      RECT 41.86 3.795 41.89 5.075 ;
      RECT 41.84 3.795 41.86 5.089 ;
      RECT 41.82 3.795 41.84 4.605 ;
      RECT 41.835 4.672 41.84 5.094 ;
      RECT 41.83 4.702 41.835 5.096 ;
      RECT 41.825 4.715 41.83 5.099 ;
      RECT 41.82 4.725 41.825 5.103 ;
      RECT 41.815 3.795 41.82 4.523 ;
      RECT 41.815 4.735 41.82 5.105 ;
      RECT 41.81 3.795 41.815 4.5 ;
      RECT 41.8 4.757 41.815 5.105 ;
      RECT 41.795 3.795 41.81 4.445 ;
      RECT 41.79 4.782 41.8 5.105 ;
      RECT 41.79 3.795 41.795 4.39 ;
      RECT 41.78 3.795 41.79 4.338 ;
      RECT 41.785 4.795 41.79 5.106 ;
      RECT 41.78 4.807 41.785 5.107 ;
      RECT 41.775 3.795 41.78 4.298 ;
      RECT 41.775 4.82 41.78 5.108 ;
      RECT 41.76 4.835 41.775 5.109 ;
      RECT 41.765 3.795 41.77 4.26 ;
      RECT 41.76 3.795 41.765 4.225 ;
      RECT 41.755 3.795 41.76 4.2 ;
      RECT 41.75 4.862 41.76 5.111 ;
      RECT 41.745 3.795 41.755 4.158 ;
      RECT 41.745 4.88 41.75 5.112 ;
      RECT 41.74 3.795 41.745 4.118 ;
      RECT 41.74 4.887 41.745 5.113 ;
      RECT 41.735 3.795 41.74 4.09 ;
      RECT 41.73 4.905 41.74 5.114 ;
      RECT 41.725 3.795 41.735 4.07 ;
      RECT 41.72 4.925 41.73 5.116 ;
      RECT 41.71 4.942 41.72 5.117 ;
      RECT 41.675 4.965 41.71 5.12 ;
      RECT 41.62 4.983 41.675 5.126 ;
      RECT 41.534 4.991 41.62 5.135 ;
      RECT 41.448 5.002 41.534 5.146 ;
      RECT 41.362 5.012 41.448 5.157 ;
      RECT 41.276 5.022 41.362 5.169 ;
      RECT 41.19 5.032 41.276 5.18 ;
      RECT 41.17 5.038 41.19 5.186 ;
      RECT 41.09 5.04 41.17 5.19 ;
      RECT 41.085 5.039 41.09 5.195 ;
      RECT 41.077 5.038 41.085 5.195 ;
      RECT 40.991 5.034 41.077 5.193 ;
      RECT 40.905 5.026 40.991 5.19 ;
      RECT 40.819 5.017 40.905 5.186 ;
      RECT 40.733 5.009 40.819 5.183 ;
      RECT 40.647 5.001 40.733 5.179 ;
      RECT 40.561 4.992 40.647 5.176 ;
      RECT 40.475 4.984 40.561 5.172 ;
      RECT 40.42 4.977 40.465 5.17 ;
      RECT 40.335 4.97 40.42 5.168 ;
      RECT 40.261 4.962 40.335 5.164 ;
      RECT 40.175 4.954 40.261 5.161 ;
      RECT 40.172 4.95 40.175 5.159 ;
      RECT 40.086 4.946 40.172 5.158 ;
      RECT 40 4.938 40.086 5.155 ;
      RECT 39.915 4.933 40 5.152 ;
      RECT 39.829 4.93 39.915 5.149 ;
      RECT 39.743 4.928 39.829 5.146 ;
      RECT 39.657 4.925 39.743 5.143 ;
      RECT 39.571 4.922 39.657 5.14 ;
      RECT 39.485 4.919 39.571 5.137 ;
      RECT 39.409 4.917 39.485 5.134 ;
      RECT 39.323 4.914 39.409 5.131 ;
      RECT 39.237 4.911 39.323 5.129 ;
      RECT 39.151 4.909 39.237 5.126 ;
      RECT 39.065 4.906 39.151 5.123 ;
      RECT 39.005 4.897 39.065 5.121 ;
      RECT 41.515 4.515 41.59 4.775 ;
      RECT 41.495 4.495 41.5 4.775 ;
      RECT 40.815 4.28 40.92 4.575 ;
      RECT 35.26 4.255 35.33 4.515 ;
      RECT 41.155 4.13 41.16 4.501 ;
      RECT 41.145 4.185 41.15 4.501 ;
      RECT 41.45 3.355 41.51 3.615 ;
      RECT 41.505 4.51 41.515 4.775 ;
      RECT 41.5 4.5 41.505 4.775 ;
      RECT 41.42 4.447 41.495 4.775 ;
      RECT 41.445 3.355 41.45 3.635 ;
      RECT 41.435 3.355 41.445 3.655 ;
      RECT 41.42 3.355 41.435 3.685 ;
      RECT 41.405 3.355 41.42 3.728 ;
      RECT 41.4 4.39 41.42 4.775 ;
      RECT 41.39 3.355 41.405 3.765 ;
      RECT 41.385 4.37 41.4 4.775 ;
      RECT 41.385 3.355 41.39 3.788 ;
      RECT 41.375 3.355 41.385 3.813 ;
      RECT 41.345 4.337 41.385 4.775 ;
      RECT 41.35 3.355 41.375 3.863 ;
      RECT 41.345 3.355 41.35 3.918 ;
      RECT 41.34 3.355 41.345 3.96 ;
      RECT 41.33 4.3 41.345 4.775 ;
      RECT 41.335 3.355 41.34 4.003 ;
      RECT 41.33 3.355 41.335 4.068 ;
      RECT 41.325 3.355 41.33 4.09 ;
      RECT 41.325 4.288 41.33 4.64 ;
      RECT 41.32 3.355 41.325 4.158 ;
      RECT 41.32 4.28 41.325 4.623 ;
      RECT 41.315 3.355 41.32 4.203 ;
      RECT 41.31 4.262 41.32 4.6 ;
      RECT 41.31 3.355 41.315 4.24 ;
      RECT 41.3 3.355 41.31 4.58 ;
      RECT 41.295 3.355 41.3 4.563 ;
      RECT 41.29 3.355 41.295 4.548 ;
      RECT 41.285 3.355 41.29 4.533 ;
      RECT 41.265 3.355 41.285 4.523 ;
      RECT 41.26 3.355 41.265 4.513 ;
      RECT 41.25 3.355 41.26 4.509 ;
      RECT 41.245 3.632 41.25 4.508 ;
      RECT 41.24 3.655 41.245 4.507 ;
      RECT 41.235 3.685 41.24 4.506 ;
      RECT 41.23 3.712 41.235 4.505 ;
      RECT 41.225 3.74 41.23 4.505 ;
      RECT 41.22 3.767 41.225 4.505 ;
      RECT 41.215 3.787 41.22 4.505 ;
      RECT 41.21 3.815 41.215 4.505 ;
      RECT 41.2 3.857 41.21 4.505 ;
      RECT 41.19 3.902 41.2 4.504 ;
      RECT 41.185 3.955 41.19 4.503 ;
      RECT 41.18 3.987 41.185 4.502 ;
      RECT 41.175 4.007 41.18 4.501 ;
      RECT 41.17 4.045 41.175 4.501 ;
      RECT 41.165 4.067 41.17 4.501 ;
      RECT 41.16 4.092 41.165 4.501 ;
      RECT 41.15 4.157 41.155 4.501 ;
      RECT 41.135 4.217 41.145 4.501 ;
      RECT 41.12 4.227 41.135 4.501 ;
      RECT 41.1 4.237 41.12 4.501 ;
      RECT 41.07 4.242 41.1 4.498 ;
      RECT 41.01 4.252 41.07 4.495 ;
      RECT 40.99 4.261 41.01 4.5 ;
      RECT 40.965 4.267 40.99 4.513 ;
      RECT 40.945 4.272 40.965 4.528 ;
      RECT 40.92 4.277 40.945 4.575 ;
      RECT 40.791 4.279 40.815 4.575 ;
      RECT 40.705 4.274 40.791 4.575 ;
      RECT 40.665 4.271 40.705 4.575 ;
      RECT 40.615 4.273 40.665 4.555 ;
      RECT 40.585 4.277 40.615 4.555 ;
      RECT 40.506 4.287 40.585 4.555 ;
      RECT 40.42 4.302 40.506 4.556 ;
      RECT 40.37 4.312 40.42 4.557 ;
      RECT 40.362 4.315 40.37 4.557 ;
      RECT 40.276 4.317 40.362 4.558 ;
      RECT 40.19 4.321 40.276 4.558 ;
      RECT 40.104 4.325 40.19 4.559 ;
      RECT 40.018 4.328 40.104 4.56 ;
      RECT 39.932 4.332 40.018 4.56 ;
      RECT 39.846 4.336 39.932 4.561 ;
      RECT 39.76 4.339 39.846 4.562 ;
      RECT 39.674 4.343 39.76 4.562 ;
      RECT 39.588 4.347 39.674 4.563 ;
      RECT 39.502 4.351 39.588 4.564 ;
      RECT 39.416 4.354 39.502 4.564 ;
      RECT 39.33 4.358 39.416 4.565 ;
      RECT 39.3 4.36 39.33 4.565 ;
      RECT 39.214 4.363 39.3 4.566 ;
      RECT 39.128 4.367 39.214 4.567 ;
      RECT 39.042 4.371 39.128 4.568 ;
      RECT 38.956 4.374 39.042 4.568 ;
      RECT 38.87 4.378 38.956 4.569 ;
      RECT 38.835 4.383 38.87 4.57 ;
      RECT 38.78 4.393 38.835 4.577 ;
      RECT 38.755 4.405 38.78 4.587 ;
      RECT 38.72 4.418 38.755 4.595 ;
      RECT 38.68 4.435 38.72 4.618 ;
      RECT 38.66 4.448 38.68 4.645 ;
      RECT 38.63 4.46 38.66 4.673 ;
      RECT 38.625 4.468 38.63 4.693 ;
      RECT 38.62 4.471 38.625 4.703 ;
      RECT 38.57 4.483 38.62 4.737 ;
      RECT 38.56 4.498 38.57 4.77 ;
      RECT 38.55 4.504 38.56 4.783 ;
      RECT 38.54 4.511 38.55 4.795 ;
      RECT 38.515 4.524 38.54 4.813 ;
      RECT 38.5 4.539 38.515 4.835 ;
      RECT 38.49 4.547 38.5 4.851 ;
      RECT 38.475 4.556 38.49 4.866 ;
      RECT 38.465 4.566 38.475 4.88 ;
      RECT 38.446 4.579 38.465 4.897 ;
      RECT 38.36 4.624 38.446 4.962 ;
      RECT 38.345 4.669 38.36 5.02 ;
      RECT 38.34 4.678 38.345 5.033 ;
      RECT 38.33 4.685 38.34 5.038 ;
      RECT 38.325 4.69 38.33 5.042 ;
      RECT 38.305 4.7 38.325 5.049 ;
      RECT 38.28 4.72 38.305 5.063 ;
      RECT 38.245 4.745 38.28 5.083 ;
      RECT 38.23 4.768 38.245 5.098 ;
      RECT 38.22 4.778 38.23 5.103 ;
      RECT 38.21 4.786 38.22 5.11 ;
      RECT 38.2 4.795 38.21 5.116 ;
      RECT 38.18 4.807 38.2 5.118 ;
      RECT 38.17 4.82 38.18 5.12 ;
      RECT 38.145 4.835 38.17 5.123 ;
      RECT 38.125 4.852 38.145 5.127 ;
      RECT 38.085 4.88 38.125 5.133 ;
      RECT 38.02 4.927 38.085 5.142 ;
      RECT 38.005 4.96 38.02 5.15 ;
      RECT 38 4.967 38.005 5.152 ;
      RECT 37.95 4.992 38 5.157 ;
      RECT 37.935 5.016 37.95 5.164 ;
      RECT 37.885 5.021 37.935 5.165 ;
      RECT 37.799 5.025 37.885 5.165 ;
      RECT 37.713 5.025 37.799 5.165 ;
      RECT 37.627 5.025 37.713 5.166 ;
      RECT 37.541 5.025 37.627 5.166 ;
      RECT 37.455 5.025 37.541 5.166 ;
      RECT 37.389 5.025 37.455 5.166 ;
      RECT 37.303 5.025 37.389 5.167 ;
      RECT 37.217 5.025 37.303 5.167 ;
      RECT 37.131 5.026 37.217 5.168 ;
      RECT 37.045 5.026 37.131 5.168 ;
      RECT 36.959 5.026 37.045 5.168 ;
      RECT 36.873 5.026 36.959 5.169 ;
      RECT 36.787 5.026 36.873 5.169 ;
      RECT 36.701 5.027 36.787 5.17 ;
      RECT 36.615 5.027 36.701 5.17 ;
      RECT 36.595 5.027 36.615 5.17 ;
      RECT 36.509 5.027 36.595 5.17 ;
      RECT 36.423 5.027 36.509 5.17 ;
      RECT 36.337 5.028 36.423 5.17 ;
      RECT 36.251 5.028 36.337 5.17 ;
      RECT 36.165 5.028 36.251 5.17 ;
      RECT 36.079 5.029 36.165 5.17 ;
      RECT 35.993 5.029 36.079 5.17 ;
      RECT 35.907 5.029 35.993 5.17 ;
      RECT 35.821 5.029 35.907 5.17 ;
      RECT 35.735 5.03 35.821 5.17 ;
      RECT 35.685 5.027 35.735 5.17 ;
      RECT 35.675 5.025 35.685 5.169 ;
      RECT 35.671 5.025 35.675 5.168 ;
      RECT 35.585 5.02 35.671 5.163 ;
      RECT 35.563 5.013 35.585 5.157 ;
      RECT 35.477 5.004 35.563 5.151 ;
      RECT 35.391 4.991 35.477 5.142 ;
      RECT 35.305 4.977 35.391 5.132 ;
      RECT 35.26 4.967 35.305 5.125 ;
      RECT 35.24 4.255 35.26 4.533 ;
      RECT 35.24 4.96 35.26 5.121 ;
      RECT 35.21 4.255 35.24 4.555 ;
      RECT 35.2 4.927 35.24 5.118 ;
      RECT 35.195 4.255 35.21 4.575 ;
      RECT 35.195 4.892 35.2 5.116 ;
      RECT 35.19 4.255 35.195 4.7 ;
      RECT 35.19 4.852 35.195 5.116 ;
      RECT 35.18 4.255 35.19 5.116 ;
      RECT 35.105 4.255 35.18 5.11 ;
      RECT 35.075 4.255 35.105 5.1 ;
      RECT 35.07 4.255 35.075 5.092 ;
      RECT 35.065 4.297 35.07 5.085 ;
      RECT 35.055 4.366 35.065 5.076 ;
      RECT 35.05 4.436 35.055 5.028 ;
      RECT 35.045 4.5 35.05 4.925 ;
      RECT 35.04 4.535 35.045 4.88 ;
      RECT 35.038 4.572 35.04 4.772 ;
      RECT 35.035 4.58 35.038 4.765 ;
      RECT 35.03 4.645 35.035 4.708 ;
      RECT 39.105 3.735 39.385 4.015 ;
      RECT 39.095 3.735 39.385 3.878 ;
      RECT 39.05 3.6 39.31 3.86 ;
      RECT 39.05 3.715 39.365 3.86 ;
      RECT 39.05 3.685 39.36 3.86 ;
      RECT 39.05 3.672 39.35 3.86 ;
      RECT 39.05 3.662 39.345 3.86 ;
      RECT 35.025 3.645 35.285 3.905 ;
      RECT 38.795 3.195 39.055 3.455 ;
      RECT 38.785 3.22 39.055 3.415 ;
      RECT 38.78 3.22 38.785 3.414 ;
      RECT 38.71 3.215 38.78 3.406 ;
      RECT 38.625 3.202 38.71 3.389 ;
      RECT 38.621 3.194 38.625 3.379 ;
      RECT 38.535 3.187 38.621 3.369 ;
      RECT 38.526 3.179 38.535 3.359 ;
      RECT 38.44 3.172 38.526 3.347 ;
      RECT 38.42 3.163 38.44 3.333 ;
      RECT 38.365 3.158 38.42 3.325 ;
      RECT 38.355 3.152 38.365 3.319 ;
      RECT 38.335 3.15 38.355 3.315 ;
      RECT 38.327 3.149 38.335 3.311 ;
      RECT 38.241 3.141 38.327 3.3 ;
      RECT 38.155 3.127 38.241 3.28 ;
      RECT 38.095 3.115 38.155 3.265 ;
      RECT 38.085 3.11 38.095 3.26 ;
      RECT 38.035 3.11 38.085 3.262 ;
      RECT 37.988 3.112 38.035 3.266 ;
      RECT 37.902 3.119 37.988 3.271 ;
      RECT 37.816 3.127 37.902 3.277 ;
      RECT 37.73 3.136 37.816 3.283 ;
      RECT 37.671 3.142 37.73 3.288 ;
      RECT 37.585 3.147 37.671 3.294 ;
      RECT 37.51 3.152 37.585 3.3 ;
      RECT 37.471 3.154 37.51 3.305 ;
      RECT 37.385 3.151 37.471 3.31 ;
      RECT 37.3 3.149 37.385 3.317 ;
      RECT 37.268 3.148 37.3 3.32 ;
      RECT 37.182 3.147 37.268 3.321 ;
      RECT 37.096 3.146 37.182 3.322 ;
      RECT 37.01 3.145 37.096 3.322 ;
      RECT 36.924 3.144 37.01 3.323 ;
      RECT 36.838 3.143 36.924 3.324 ;
      RECT 36.752 3.142 36.838 3.325 ;
      RECT 36.666 3.141 36.752 3.325 ;
      RECT 36.58 3.14 36.666 3.326 ;
      RECT 36.53 3.14 36.58 3.327 ;
      RECT 36.516 3.141 36.53 3.327 ;
      RECT 36.43 3.148 36.516 3.328 ;
      RECT 36.356 3.159 36.43 3.329 ;
      RECT 36.27 3.168 36.356 3.33 ;
      RECT 36.235 3.175 36.27 3.345 ;
      RECT 36.21 3.178 36.235 3.375 ;
      RECT 36.185 3.187 36.21 3.404 ;
      RECT 36.175 3.198 36.185 3.424 ;
      RECT 36.165 3.206 36.175 3.438 ;
      RECT 36.16 3.212 36.165 3.448 ;
      RECT 36.135 3.229 36.16 3.465 ;
      RECT 36.12 3.251 36.135 3.493 ;
      RECT 36.09 3.277 36.12 3.523 ;
      RECT 36.07 3.306 36.09 3.553 ;
      RECT 36.065 3.321 36.07 3.57 ;
      RECT 36.045 3.336 36.065 3.585 ;
      RECT 36.035 3.354 36.045 3.603 ;
      RECT 36.025 3.365 36.035 3.618 ;
      RECT 35.975 3.397 36.025 3.644 ;
      RECT 35.97 3.427 35.975 3.664 ;
      RECT 35.96 3.44 35.97 3.67 ;
      RECT 35.951 3.45 35.96 3.678 ;
      RECT 35.94 3.461 35.951 3.686 ;
      RECT 35.935 3.471 35.94 3.692 ;
      RECT 35.92 3.492 35.935 3.699 ;
      RECT 35.905 3.522 35.92 3.707 ;
      RECT 35.87 3.552 35.905 3.713 ;
      RECT 35.845 3.57 35.87 3.72 ;
      RECT 35.795 3.578 35.845 3.729 ;
      RECT 35.77 3.583 35.795 3.738 ;
      RECT 35.715 3.589 35.77 3.748 ;
      RECT 35.71 3.594 35.715 3.756 ;
      RECT 35.696 3.597 35.71 3.758 ;
      RECT 35.61 3.609 35.696 3.77 ;
      RECT 35.6 3.621 35.61 3.783 ;
      RECT 35.515 3.634 35.6 3.795 ;
      RECT 35.471 3.651 35.515 3.809 ;
      RECT 35.385 3.668 35.471 3.825 ;
      RECT 35.355 3.682 35.385 3.839 ;
      RECT 35.345 3.687 35.355 3.844 ;
      RECT 35.285 3.69 35.345 3.853 ;
      RECT 38.175 3.96 38.435 4.22 ;
      RECT 38.175 3.96 38.455 4.073 ;
      RECT 38.175 3.96 38.48 4.04 ;
      RECT 38.175 3.96 38.485 4.02 ;
      RECT 38.225 3.735 38.505 4.015 ;
      RECT 37.78 4.47 38.04 4.73 ;
      RECT 37.77 4.327 37.965 4.668 ;
      RECT 37.765 4.435 37.98 4.66 ;
      RECT 37.76 4.485 38.04 4.65 ;
      RECT 37.75 4.562 38.04 4.635 ;
      RECT 37.77 4.41 37.98 4.668 ;
      RECT 37.78 4.285 37.965 4.73 ;
      RECT 37.78 4.18 37.945 4.73 ;
      RECT 37.79 4.167 37.945 4.73 ;
      RECT 37.79 4.125 37.935 4.73 ;
      RECT 37.795 4.05 37.935 4.73 ;
      RECT 37.825 3.7 37.935 4.73 ;
      RECT 37.83 3.43 37.955 4.053 ;
      RECT 37.8 4.005 37.955 4.053 ;
      RECT 37.815 3.807 37.935 4.73 ;
      RECT 37.805 3.917 37.955 4.053 ;
      RECT 37.83 3.43 37.97 3.91 ;
      RECT 37.83 3.43 37.99 3.785 ;
      RECT 37.795 3.43 38.055 3.69 ;
      RECT 37.265 3.735 37.545 4.015 ;
      RECT 37.25 3.735 37.545 3.995 ;
      RECT 35.305 4.6 35.565 4.86 ;
      RECT 37.09 4.455 37.35 4.715 ;
      RECT 37.07 4.475 37.35 4.69 ;
      RECT 37.027 4.475 37.07 4.689 ;
      RECT 36.941 4.476 37.027 4.686 ;
      RECT 36.855 4.477 36.941 4.682 ;
      RECT 36.78 4.479 36.855 4.679 ;
      RECT 36.757 4.48 36.78 4.677 ;
      RECT 36.671 4.481 36.757 4.675 ;
      RECT 36.585 4.482 36.671 4.672 ;
      RECT 36.561 4.483 36.585 4.67 ;
      RECT 36.475 4.485 36.561 4.667 ;
      RECT 36.39 4.487 36.475 4.668 ;
      RECT 36.333 4.488 36.39 4.674 ;
      RECT 36.247 4.49 36.333 4.684 ;
      RECT 36.161 4.493 36.247 4.697 ;
      RECT 36.075 4.495 36.161 4.709 ;
      RECT 36.061 4.496 36.075 4.716 ;
      RECT 35.975 4.497 36.061 4.724 ;
      RECT 35.935 4.499 35.975 4.733 ;
      RECT 35.926 4.5 35.935 4.736 ;
      RECT 35.84 4.508 35.926 4.742 ;
      RECT 35.82 4.517 35.84 4.75 ;
      RECT 35.735 4.532 35.82 4.758 ;
      RECT 35.675 4.555 35.735 4.769 ;
      RECT 35.665 4.567 35.675 4.774 ;
      RECT 35.625 4.577 35.665 4.778 ;
      RECT 35.57 4.594 35.625 4.786 ;
      RECT 35.565 4.604 35.57 4.79 ;
      RECT 36.631 3.735 36.69 4.132 ;
      RECT 36.545 3.735 36.75 4.123 ;
      RECT 36.54 3.765 36.75 4.118 ;
      RECT 36.506 3.765 36.75 4.116 ;
      RECT 36.42 3.765 36.75 4.11 ;
      RECT 36.375 3.765 36.77 4.088 ;
      RECT 36.375 3.765 36.79 4.043 ;
      RECT 36.335 3.765 36.79 4.033 ;
      RECT 36.545 3.735 36.825 4.015 ;
      RECT 36.28 3.735 36.54 3.995 ;
      RECT 35.465 3.215 35.725 3.475 ;
      RECT 35.545 3.175 35.825 3.455 ;
      RECT 29.915 8.505 30.235 8.83 ;
      RECT 29.945 7.98 30.115 8.83 ;
      RECT 29.945 7.98 30.12 8.33 ;
      RECT 29.945 7.98 30.92 8.155 ;
      RECT 30.745 3.26 30.92 8.155 ;
      RECT 30.69 3.26 31.04 3.61 ;
      RECT 30.715 8.94 31.04 9.265 ;
      RECT 29.6 9.03 31.04 9.2 ;
      RECT 29.6 3.69 29.76 9.2 ;
      RECT 29.915 3.66 30.235 3.98 ;
      RECT 29.6 3.69 30.235 3.86 ;
      RECT 18.325 4.295 18.605 4.575 ;
      RECT 18.295 4.295 18.605 4.56 ;
      RECT 18.29 4.295 18.605 4.558 ;
      RECT 18.285 2.625 18.455 4.552 ;
      RECT 18.28 4.262 18.55 4.545 ;
      RECT 18.275 4.295 18.605 4.538 ;
      RECT 18.245 4.265 18.55 4.525 ;
      RECT 18.245 4.292 18.57 4.525 ;
      RECT 18.245 4.282 18.565 4.525 ;
      RECT 18.245 4.267 18.56 4.525 ;
      RECT 18.285 4.257 18.55 4.552 ;
      RECT 18.285 4.252 18.54 4.552 ;
      RECT 18.285 4.251 18.525 4.552 ;
      RECT 28.255 2.635 28.605 2.985 ;
      RECT 28.25 2.635 28.605 2.89 ;
      RECT 18.285 2.625 28.495 2.795 ;
      RECT 27.93 4.145 28.3 4.515 ;
      RECT 28.015 3.53 28.185 4.515 ;
      RECT 24.035 3.75 24.27 4.01 ;
      RECT 27.18 3.53 27.345 3.79 ;
      RECT 27.085 3.52 27.1 3.79 ;
      RECT 27.18 3.53 28.185 3.71 ;
      RECT 25.685 3.09 25.725 3.23 ;
      RECT 27.1 3.525 27.18 3.79 ;
      RECT 27.045 3.52 27.085 3.756 ;
      RECT 27.031 3.52 27.045 3.756 ;
      RECT 26.945 3.525 27.031 3.758 ;
      RECT 26.9 3.532 26.945 3.76 ;
      RECT 26.87 3.532 26.9 3.762 ;
      RECT 26.845 3.527 26.87 3.764 ;
      RECT 26.815 3.523 26.845 3.773 ;
      RECT 26.805 3.52 26.815 3.785 ;
      RECT 26.8 3.52 26.805 3.793 ;
      RECT 26.795 3.52 26.8 3.798 ;
      RECT 26.785 3.519 26.795 3.808 ;
      RECT 26.78 3.518 26.785 3.818 ;
      RECT 26.765 3.517 26.78 3.823 ;
      RECT 26.737 3.514 26.765 3.85 ;
      RECT 26.651 3.506 26.737 3.85 ;
      RECT 26.565 3.495 26.651 3.85 ;
      RECT 26.525 3.48 26.565 3.85 ;
      RECT 26.485 3.454 26.525 3.85 ;
      RECT 26.48 3.436 26.485 3.662 ;
      RECT 26.47 3.432 26.48 3.652 ;
      RECT 26.455 3.422 26.47 3.639 ;
      RECT 26.435 3.406 26.455 3.624 ;
      RECT 26.42 3.391 26.435 3.609 ;
      RECT 26.41 3.38 26.42 3.599 ;
      RECT 26.385 3.364 26.41 3.588 ;
      RECT 26.38 3.351 26.385 3.578 ;
      RECT 26.375 3.347 26.38 3.573 ;
      RECT 26.32 3.333 26.375 3.551 ;
      RECT 26.281 3.314 26.32 3.515 ;
      RECT 26.195 3.288 26.281 3.468 ;
      RECT 26.191 3.27 26.195 3.434 ;
      RECT 26.105 3.251 26.191 3.412 ;
      RECT 26.1 3.233 26.105 3.39 ;
      RECT 26.095 3.231 26.1 3.388 ;
      RECT 26.085 3.23 26.095 3.383 ;
      RECT 26.025 3.217 26.085 3.369 ;
      RECT 25.98 3.195 26.025 3.348 ;
      RECT 25.92 3.172 25.98 3.327 ;
      RECT 25.856 3.147 25.92 3.302 ;
      RECT 25.77 3.117 25.856 3.271 ;
      RECT 25.755 3.097 25.77 3.25 ;
      RECT 25.725 3.092 25.755 3.241 ;
      RECT 25.672 3.09 25.685 3.23 ;
      RECT 25.586 3.09 25.672 3.232 ;
      RECT 25.5 3.09 25.586 3.234 ;
      RECT 25.48 3.09 25.5 3.238 ;
      RECT 25.435 3.092 25.48 3.249 ;
      RECT 25.395 3.102 25.435 3.265 ;
      RECT 25.391 3.111 25.395 3.273 ;
      RECT 25.305 3.131 25.391 3.289 ;
      RECT 25.295 3.15 25.305 3.307 ;
      RECT 25.29 3.152 25.295 3.31 ;
      RECT 25.28 3.156 25.29 3.313 ;
      RECT 25.26 3.161 25.28 3.323 ;
      RECT 25.23 3.171 25.26 3.343 ;
      RECT 25.225 3.178 25.23 3.357 ;
      RECT 25.215 3.182 25.225 3.364 ;
      RECT 25.2 3.19 25.215 3.375 ;
      RECT 25.19 3.2 25.2 3.386 ;
      RECT 25.18 3.207 25.19 3.394 ;
      RECT 25.155 3.22 25.18 3.409 ;
      RECT 25.091 3.256 25.155 3.448 ;
      RECT 25.005 3.319 25.091 3.512 ;
      RECT 24.97 3.37 25.005 3.565 ;
      RECT 24.965 3.387 24.97 3.582 ;
      RECT 24.95 3.396 24.965 3.589 ;
      RECT 24.93 3.411 24.95 3.603 ;
      RECT 24.925 3.422 24.93 3.613 ;
      RECT 24.905 3.435 24.925 3.623 ;
      RECT 24.9 3.445 24.905 3.633 ;
      RECT 24.885 3.45 24.9 3.642 ;
      RECT 24.875 3.46 24.885 3.653 ;
      RECT 24.845 3.477 24.875 3.67 ;
      RECT 24.835 3.495 24.845 3.688 ;
      RECT 24.82 3.506 24.835 3.699 ;
      RECT 24.78 3.53 24.82 3.715 ;
      RECT 24.745 3.564 24.78 3.732 ;
      RECT 24.715 3.587 24.745 3.744 ;
      RECT 24.7 3.597 24.715 3.753 ;
      RECT 24.66 3.607 24.7 3.764 ;
      RECT 24.64 3.618 24.66 3.776 ;
      RECT 24.635 3.622 24.64 3.783 ;
      RECT 24.62 3.626 24.635 3.788 ;
      RECT 24.61 3.631 24.62 3.793 ;
      RECT 24.605 3.634 24.61 3.796 ;
      RECT 24.575 3.64 24.605 3.803 ;
      RECT 24.54 3.65 24.575 3.817 ;
      RECT 24.48 3.665 24.54 3.837 ;
      RECT 24.425 3.685 24.48 3.861 ;
      RECT 24.396 3.7 24.425 3.879 ;
      RECT 24.31 3.72 24.396 3.904 ;
      RECT 24.305 3.735 24.31 3.924 ;
      RECT 24.295 3.738 24.305 3.925 ;
      RECT 24.27 3.745 24.295 4.01 ;
      RECT 16.545 9.28 16.835 9.63 ;
      RECT 16.545 9.34 17.96 9.51 ;
      RECT 17.79 8.97 17.96 9.51 ;
      RECT 26.11 8.89 26.46 9.24 ;
      RECT 17.79 8.97 26.46 9.14 ;
      RECT 24.685 4.98 24.695 5.17 ;
      RECT 22.945 4.855 23.225 5.135 ;
      RECT 25.99 3.795 25.995 4.28 ;
      RECT 25.885 3.795 25.945 4.055 ;
      RECT 26.21 4.765 26.215 4.84 ;
      RECT 26.2 4.632 26.21 4.875 ;
      RECT 26.19 4.467 26.2 4.896 ;
      RECT 26.185 4.337 26.19 4.912 ;
      RECT 26.175 4.227 26.185 4.928 ;
      RECT 26.17 4.126 26.175 4.945 ;
      RECT 26.165 4.108 26.17 4.955 ;
      RECT 26.16 4.09 26.165 4.965 ;
      RECT 26.15 4.065 26.16 4.98 ;
      RECT 26.145 4.045 26.15 4.995 ;
      RECT 26.125 3.795 26.145 5.02 ;
      RECT 26.11 3.795 26.125 5.053 ;
      RECT 26.08 3.795 26.11 5.075 ;
      RECT 26.06 3.795 26.08 5.089 ;
      RECT 26.04 3.795 26.06 4.605 ;
      RECT 26.055 4.672 26.06 5.094 ;
      RECT 26.05 4.702 26.055 5.096 ;
      RECT 26.045 4.715 26.05 5.099 ;
      RECT 26.04 4.725 26.045 5.103 ;
      RECT 26.035 3.795 26.04 4.523 ;
      RECT 26.035 4.735 26.04 5.105 ;
      RECT 26.03 3.795 26.035 4.5 ;
      RECT 26.02 4.757 26.035 5.105 ;
      RECT 26.015 3.795 26.03 4.445 ;
      RECT 26.01 4.782 26.02 5.105 ;
      RECT 26.01 3.795 26.015 4.39 ;
      RECT 26 3.795 26.01 4.338 ;
      RECT 26.005 4.795 26.01 5.106 ;
      RECT 26 4.807 26.005 5.107 ;
      RECT 25.995 3.795 26 4.298 ;
      RECT 25.995 4.82 26 5.108 ;
      RECT 25.98 4.835 25.995 5.109 ;
      RECT 25.985 3.795 25.99 4.26 ;
      RECT 25.98 3.795 25.985 4.225 ;
      RECT 25.975 3.795 25.98 4.2 ;
      RECT 25.97 4.862 25.98 5.111 ;
      RECT 25.965 3.795 25.975 4.158 ;
      RECT 25.965 4.88 25.97 5.112 ;
      RECT 25.96 3.795 25.965 4.118 ;
      RECT 25.96 4.887 25.965 5.113 ;
      RECT 25.955 3.795 25.96 4.09 ;
      RECT 25.95 4.905 25.96 5.114 ;
      RECT 25.945 3.795 25.955 4.07 ;
      RECT 25.94 4.925 25.95 5.116 ;
      RECT 25.93 4.942 25.94 5.117 ;
      RECT 25.895 4.965 25.93 5.12 ;
      RECT 25.84 4.983 25.895 5.126 ;
      RECT 25.754 4.991 25.84 5.135 ;
      RECT 25.668 5.002 25.754 5.146 ;
      RECT 25.582 5.012 25.668 5.157 ;
      RECT 25.496 5.022 25.582 5.169 ;
      RECT 25.41 5.032 25.496 5.18 ;
      RECT 25.39 5.038 25.41 5.186 ;
      RECT 25.31 5.04 25.39 5.19 ;
      RECT 25.305 5.039 25.31 5.195 ;
      RECT 25.297 5.038 25.305 5.195 ;
      RECT 25.211 5.034 25.297 5.193 ;
      RECT 25.125 5.026 25.211 5.19 ;
      RECT 25.039 5.017 25.125 5.186 ;
      RECT 24.953 5.009 25.039 5.183 ;
      RECT 24.867 5.001 24.953 5.179 ;
      RECT 24.781 4.992 24.867 5.176 ;
      RECT 24.695 4.984 24.781 5.172 ;
      RECT 24.64 4.977 24.685 5.17 ;
      RECT 24.555 4.97 24.64 5.168 ;
      RECT 24.481 4.962 24.555 5.164 ;
      RECT 24.395 4.954 24.481 5.161 ;
      RECT 24.392 4.95 24.395 5.159 ;
      RECT 24.306 4.946 24.392 5.158 ;
      RECT 24.22 4.938 24.306 5.155 ;
      RECT 24.135 4.933 24.22 5.152 ;
      RECT 24.049 4.93 24.135 5.149 ;
      RECT 23.963 4.928 24.049 5.146 ;
      RECT 23.877 4.925 23.963 5.143 ;
      RECT 23.791 4.922 23.877 5.14 ;
      RECT 23.705 4.919 23.791 5.137 ;
      RECT 23.629 4.917 23.705 5.134 ;
      RECT 23.543 4.914 23.629 5.131 ;
      RECT 23.457 4.911 23.543 5.129 ;
      RECT 23.371 4.909 23.457 5.126 ;
      RECT 23.285 4.906 23.371 5.123 ;
      RECT 23.225 4.897 23.285 5.121 ;
      RECT 25.735 4.515 25.81 4.775 ;
      RECT 25.715 4.495 25.72 4.775 ;
      RECT 25.035 4.28 25.14 4.575 ;
      RECT 19.48 4.255 19.55 4.515 ;
      RECT 25.375 4.13 25.38 4.501 ;
      RECT 25.365 4.185 25.37 4.501 ;
      RECT 25.67 3.355 25.73 3.615 ;
      RECT 25.725 4.51 25.735 4.775 ;
      RECT 25.72 4.5 25.725 4.775 ;
      RECT 25.64 4.447 25.715 4.775 ;
      RECT 25.665 3.355 25.67 3.635 ;
      RECT 25.655 3.355 25.665 3.655 ;
      RECT 25.64 3.355 25.655 3.685 ;
      RECT 25.625 3.355 25.64 3.728 ;
      RECT 25.62 4.39 25.64 4.775 ;
      RECT 25.61 3.355 25.625 3.765 ;
      RECT 25.605 4.37 25.62 4.775 ;
      RECT 25.605 3.355 25.61 3.788 ;
      RECT 25.595 3.355 25.605 3.813 ;
      RECT 25.565 4.337 25.605 4.775 ;
      RECT 25.57 3.355 25.595 3.863 ;
      RECT 25.565 3.355 25.57 3.918 ;
      RECT 25.56 3.355 25.565 3.96 ;
      RECT 25.55 4.3 25.565 4.775 ;
      RECT 25.555 3.355 25.56 4.003 ;
      RECT 25.55 3.355 25.555 4.068 ;
      RECT 25.545 3.355 25.55 4.09 ;
      RECT 25.545 4.288 25.55 4.64 ;
      RECT 25.54 3.355 25.545 4.158 ;
      RECT 25.54 4.28 25.545 4.623 ;
      RECT 25.535 3.355 25.54 4.203 ;
      RECT 25.53 4.262 25.54 4.6 ;
      RECT 25.53 3.355 25.535 4.24 ;
      RECT 25.52 3.355 25.53 4.58 ;
      RECT 25.515 3.355 25.52 4.563 ;
      RECT 25.51 3.355 25.515 4.548 ;
      RECT 25.505 3.355 25.51 4.533 ;
      RECT 25.485 3.355 25.505 4.523 ;
      RECT 25.48 3.355 25.485 4.513 ;
      RECT 25.47 3.355 25.48 4.509 ;
      RECT 25.465 3.632 25.47 4.508 ;
      RECT 25.46 3.655 25.465 4.507 ;
      RECT 25.455 3.685 25.46 4.506 ;
      RECT 25.45 3.712 25.455 4.505 ;
      RECT 25.445 3.74 25.45 4.505 ;
      RECT 25.44 3.767 25.445 4.505 ;
      RECT 25.435 3.787 25.44 4.505 ;
      RECT 25.43 3.815 25.435 4.505 ;
      RECT 25.42 3.857 25.43 4.505 ;
      RECT 25.41 3.902 25.42 4.504 ;
      RECT 25.405 3.955 25.41 4.503 ;
      RECT 25.4 3.987 25.405 4.502 ;
      RECT 25.395 4.007 25.4 4.501 ;
      RECT 25.39 4.045 25.395 4.501 ;
      RECT 25.385 4.067 25.39 4.501 ;
      RECT 25.38 4.092 25.385 4.501 ;
      RECT 25.37 4.157 25.375 4.501 ;
      RECT 25.355 4.217 25.365 4.501 ;
      RECT 25.34 4.227 25.355 4.501 ;
      RECT 25.32 4.237 25.34 4.501 ;
      RECT 25.29 4.242 25.32 4.498 ;
      RECT 25.23 4.252 25.29 4.495 ;
      RECT 25.21 4.261 25.23 4.5 ;
      RECT 25.185 4.267 25.21 4.513 ;
      RECT 25.165 4.272 25.185 4.528 ;
      RECT 25.14 4.277 25.165 4.575 ;
      RECT 25.011 4.279 25.035 4.575 ;
      RECT 24.925 4.274 25.011 4.575 ;
      RECT 24.885 4.271 24.925 4.575 ;
      RECT 24.835 4.273 24.885 4.555 ;
      RECT 24.805 4.277 24.835 4.555 ;
      RECT 24.726 4.287 24.805 4.555 ;
      RECT 24.64 4.302 24.726 4.556 ;
      RECT 24.59 4.312 24.64 4.557 ;
      RECT 24.582 4.315 24.59 4.557 ;
      RECT 24.496 4.317 24.582 4.558 ;
      RECT 24.41 4.321 24.496 4.558 ;
      RECT 24.324 4.325 24.41 4.559 ;
      RECT 24.238 4.328 24.324 4.56 ;
      RECT 24.152 4.332 24.238 4.56 ;
      RECT 24.066 4.336 24.152 4.561 ;
      RECT 23.98 4.339 24.066 4.562 ;
      RECT 23.894 4.343 23.98 4.562 ;
      RECT 23.808 4.347 23.894 4.563 ;
      RECT 23.722 4.351 23.808 4.564 ;
      RECT 23.636 4.354 23.722 4.564 ;
      RECT 23.55 4.358 23.636 4.565 ;
      RECT 23.52 4.36 23.55 4.565 ;
      RECT 23.434 4.363 23.52 4.566 ;
      RECT 23.348 4.367 23.434 4.567 ;
      RECT 23.262 4.371 23.348 4.568 ;
      RECT 23.176 4.374 23.262 4.568 ;
      RECT 23.09 4.378 23.176 4.569 ;
      RECT 23.055 4.383 23.09 4.57 ;
      RECT 23 4.393 23.055 4.577 ;
      RECT 22.975 4.405 23 4.587 ;
      RECT 22.94 4.418 22.975 4.595 ;
      RECT 22.9 4.435 22.94 4.618 ;
      RECT 22.88 4.448 22.9 4.645 ;
      RECT 22.85 4.46 22.88 4.673 ;
      RECT 22.845 4.468 22.85 4.693 ;
      RECT 22.84 4.471 22.845 4.703 ;
      RECT 22.79 4.483 22.84 4.737 ;
      RECT 22.78 4.498 22.79 4.77 ;
      RECT 22.77 4.504 22.78 4.783 ;
      RECT 22.76 4.511 22.77 4.795 ;
      RECT 22.735 4.524 22.76 4.813 ;
      RECT 22.72 4.539 22.735 4.835 ;
      RECT 22.71 4.547 22.72 4.851 ;
      RECT 22.695 4.556 22.71 4.866 ;
      RECT 22.685 4.566 22.695 4.88 ;
      RECT 22.666 4.579 22.685 4.897 ;
      RECT 22.58 4.624 22.666 4.962 ;
      RECT 22.565 4.669 22.58 5.02 ;
      RECT 22.56 4.678 22.565 5.033 ;
      RECT 22.55 4.685 22.56 5.038 ;
      RECT 22.545 4.69 22.55 5.042 ;
      RECT 22.525 4.7 22.545 5.049 ;
      RECT 22.5 4.72 22.525 5.063 ;
      RECT 22.465 4.745 22.5 5.083 ;
      RECT 22.45 4.768 22.465 5.098 ;
      RECT 22.44 4.778 22.45 5.103 ;
      RECT 22.43 4.786 22.44 5.11 ;
      RECT 22.42 4.795 22.43 5.116 ;
      RECT 22.4 4.807 22.42 5.118 ;
      RECT 22.39 4.82 22.4 5.12 ;
      RECT 22.365 4.835 22.39 5.123 ;
      RECT 22.345 4.852 22.365 5.127 ;
      RECT 22.305 4.88 22.345 5.133 ;
      RECT 22.24 4.927 22.305 5.142 ;
      RECT 22.225 4.96 22.24 5.15 ;
      RECT 22.22 4.967 22.225 5.152 ;
      RECT 22.17 4.992 22.22 5.157 ;
      RECT 22.155 5.016 22.17 5.164 ;
      RECT 22.105 5.021 22.155 5.165 ;
      RECT 22.019 5.025 22.105 5.165 ;
      RECT 21.933 5.025 22.019 5.165 ;
      RECT 21.847 5.025 21.933 5.166 ;
      RECT 21.761 5.025 21.847 5.166 ;
      RECT 21.675 5.025 21.761 5.166 ;
      RECT 21.609 5.025 21.675 5.166 ;
      RECT 21.523 5.025 21.609 5.167 ;
      RECT 21.437 5.025 21.523 5.167 ;
      RECT 21.351 5.026 21.437 5.168 ;
      RECT 21.265 5.026 21.351 5.168 ;
      RECT 21.179 5.026 21.265 5.168 ;
      RECT 21.093 5.026 21.179 5.169 ;
      RECT 21.007 5.026 21.093 5.169 ;
      RECT 20.921 5.027 21.007 5.17 ;
      RECT 20.835 5.027 20.921 5.17 ;
      RECT 20.815 5.027 20.835 5.17 ;
      RECT 20.729 5.027 20.815 5.17 ;
      RECT 20.643 5.027 20.729 5.17 ;
      RECT 20.557 5.028 20.643 5.17 ;
      RECT 20.471 5.028 20.557 5.17 ;
      RECT 20.385 5.028 20.471 5.17 ;
      RECT 20.299 5.029 20.385 5.17 ;
      RECT 20.213 5.029 20.299 5.17 ;
      RECT 20.127 5.029 20.213 5.17 ;
      RECT 20.041 5.029 20.127 5.17 ;
      RECT 19.955 5.03 20.041 5.17 ;
      RECT 19.905 5.027 19.955 5.17 ;
      RECT 19.895 5.025 19.905 5.169 ;
      RECT 19.891 5.025 19.895 5.168 ;
      RECT 19.805 5.02 19.891 5.163 ;
      RECT 19.783 5.013 19.805 5.157 ;
      RECT 19.697 5.004 19.783 5.151 ;
      RECT 19.611 4.991 19.697 5.142 ;
      RECT 19.525 4.977 19.611 5.132 ;
      RECT 19.48 4.967 19.525 5.125 ;
      RECT 19.46 4.255 19.48 4.533 ;
      RECT 19.46 4.96 19.48 5.121 ;
      RECT 19.43 4.255 19.46 4.555 ;
      RECT 19.42 4.927 19.46 5.118 ;
      RECT 19.415 4.255 19.43 4.575 ;
      RECT 19.415 4.892 19.42 5.116 ;
      RECT 19.41 4.255 19.415 4.7 ;
      RECT 19.41 4.852 19.415 5.116 ;
      RECT 19.4 4.255 19.41 5.116 ;
      RECT 19.325 4.255 19.4 5.11 ;
      RECT 19.295 4.255 19.325 5.1 ;
      RECT 19.29 4.255 19.295 5.092 ;
      RECT 19.285 4.297 19.29 5.085 ;
      RECT 19.275 4.366 19.285 5.076 ;
      RECT 19.27 4.436 19.275 5.028 ;
      RECT 19.265 4.5 19.27 4.925 ;
      RECT 19.26 4.535 19.265 4.88 ;
      RECT 19.258 4.572 19.26 4.772 ;
      RECT 19.255 4.58 19.258 4.765 ;
      RECT 19.25 4.645 19.255 4.708 ;
      RECT 23.325 3.735 23.605 4.015 ;
      RECT 23.315 3.735 23.605 3.878 ;
      RECT 23.27 3.6 23.53 3.86 ;
      RECT 23.27 3.715 23.585 3.86 ;
      RECT 23.27 3.685 23.58 3.86 ;
      RECT 23.27 3.672 23.57 3.86 ;
      RECT 23.27 3.662 23.565 3.86 ;
      RECT 19.245 3.645 19.505 3.905 ;
      RECT 23.015 3.195 23.275 3.455 ;
      RECT 23.005 3.22 23.275 3.415 ;
      RECT 23 3.22 23.005 3.414 ;
      RECT 22.93 3.215 23 3.406 ;
      RECT 22.845 3.202 22.93 3.389 ;
      RECT 22.841 3.194 22.845 3.379 ;
      RECT 22.755 3.187 22.841 3.369 ;
      RECT 22.746 3.179 22.755 3.359 ;
      RECT 22.66 3.172 22.746 3.347 ;
      RECT 22.64 3.163 22.66 3.333 ;
      RECT 22.585 3.158 22.64 3.325 ;
      RECT 22.575 3.152 22.585 3.319 ;
      RECT 22.555 3.15 22.575 3.315 ;
      RECT 22.547 3.149 22.555 3.311 ;
      RECT 22.461 3.141 22.547 3.3 ;
      RECT 22.375 3.127 22.461 3.28 ;
      RECT 22.315 3.115 22.375 3.265 ;
      RECT 22.305 3.11 22.315 3.26 ;
      RECT 22.255 3.11 22.305 3.262 ;
      RECT 22.208 3.112 22.255 3.266 ;
      RECT 22.122 3.119 22.208 3.271 ;
      RECT 22.036 3.127 22.122 3.277 ;
      RECT 21.95 3.136 22.036 3.283 ;
      RECT 21.891 3.142 21.95 3.288 ;
      RECT 21.805 3.147 21.891 3.294 ;
      RECT 21.73 3.152 21.805 3.3 ;
      RECT 21.691 3.154 21.73 3.305 ;
      RECT 21.605 3.151 21.691 3.31 ;
      RECT 21.52 3.149 21.605 3.317 ;
      RECT 21.488 3.148 21.52 3.32 ;
      RECT 21.402 3.147 21.488 3.321 ;
      RECT 21.316 3.146 21.402 3.322 ;
      RECT 21.23 3.145 21.316 3.322 ;
      RECT 21.144 3.144 21.23 3.323 ;
      RECT 21.058 3.143 21.144 3.324 ;
      RECT 20.972 3.142 21.058 3.325 ;
      RECT 20.886 3.141 20.972 3.325 ;
      RECT 20.8 3.14 20.886 3.326 ;
      RECT 20.75 3.14 20.8 3.327 ;
      RECT 20.736 3.141 20.75 3.327 ;
      RECT 20.65 3.148 20.736 3.328 ;
      RECT 20.576 3.159 20.65 3.329 ;
      RECT 20.49 3.168 20.576 3.33 ;
      RECT 20.455 3.175 20.49 3.345 ;
      RECT 20.43 3.178 20.455 3.375 ;
      RECT 20.405 3.187 20.43 3.404 ;
      RECT 20.395 3.198 20.405 3.424 ;
      RECT 20.385 3.206 20.395 3.438 ;
      RECT 20.38 3.212 20.385 3.448 ;
      RECT 20.355 3.229 20.38 3.465 ;
      RECT 20.34 3.251 20.355 3.493 ;
      RECT 20.31 3.277 20.34 3.523 ;
      RECT 20.29 3.306 20.31 3.553 ;
      RECT 20.285 3.321 20.29 3.57 ;
      RECT 20.265 3.336 20.285 3.585 ;
      RECT 20.255 3.354 20.265 3.603 ;
      RECT 20.245 3.365 20.255 3.618 ;
      RECT 20.195 3.397 20.245 3.644 ;
      RECT 20.19 3.427 20.195 3.664 ;
      RECT 20.18 3.44 20.19 3.67 ;
      RECT 20.171 3.45 20.18 3.678 ;
      RECT 20.16 3.461 20.171 3.686 ;
      RECT 20.155 3.471 20.16 3.692 ;
      RECT 20.14 3.492 20.155 3.699 ;
      RECT 20.125 3.522 20.14 3.707 ;
      RECT 20.09 3.552 20.125 3.713 ;
      RECT 20.065 3.57 20.09 3.72 ;
      RECT 20.015 3.578 20.065 3.729 ;
      RECT 19.99 3.583 20.015 3.738 ;
      RECT 19.935 3.589 19.99 3.748 ;
      RECT 19.93 3.594 19.935 3.756 ;
      RECT 19.916 3.597 19.93 3.758 ;
      RECT 19.83 3.609 19.916 3.77 ;
      RECT 19.82 3.621 19.83 3.783 ;
      RECT 19.735 3.634 19.82 3.795 ;
      RECT 19.691 3.651 19.735 3.809 ;
      RECT 19.605 3.668 19.691 3.825 ;
      RECT 19.575 3.682 19.605 3.839 ;
      RECT 19.565 3.687 19.575 3.844 ;
      RECT 19.505 3.69 19.565 3.853 ;
      RECT 22.395 3.96 22.655 4.22 ;
      RECT 22.395 3.96 22.675 4.073 ;
      RECT 22.395 3.96 22.7 4.04 ;
      RECT 22.395 3.96 22.705 4.02 ;
      RECT 22.445 3.735 22.725 4.015 ;
      RECT 22 4.47 22.26 4.73 ;
      RECT 21.99 4.327 22.185 4.668 ;
      RECT 21.985 4.435 22.2 4.66 ;
      RECT 21.98 4.485 22.26 4.65 ;
      RECT 21.97 4.562 22.26 4.635 ;
      RECT 21.99 4.41 22.2 4.668 ;
      RECT 22 4.285 22.185 4.73 ;
      RECT 22 4.18 22.165 4.73 ;
      RECT 22.01 4.167 22.165 4.73 ;
      RECT 22.01 4.125 22.155 4.73 ;
      RECT 22.015 4.05 22.155 4.73 ;
      RECT 22.045 3.7 22.155 4.73 ;
      RECT 22.05 3.43 22.175 4.053 ;
      RECT 22.02 4.005 22.175 4.053 ;
      RECT 22.035 3.807 22.155 4.73 ;
      RECT 22.025 3.917 22.175 4.053 ;
      RECT 22.05 3.43 22.19 3.91 ;
      RECT 22.05 3.43 22.21 3.785 ;
      RECT 22.015 3.43 22.275 3.69 ;
      RECT 21.485 3.735 21.765 4.015 ;
      RECT 21.47 3.735 21.765 3.995 ;
      RECT 19.525 4.6 19.785 4.86 ;
      RECT 21.31 4.455 21.57 4.715 ;
      RECT 21.29 4.475 21.57 4.69 ;
      RECT 21.247 4.475 21.29 4.689 ;
      RECT 21.161 4.476 21.247 4.686 ;
      RECT 21.075 4.477 21.161 4.682 ;
      RECT 21 4.479 21.075 4.679 ;
      RECT 20.977 4.48 21 4.677 ;
      RECT 20.891 4.481 20.977 4.675 ;
      RECT 20.805 4.482 20.891 4.672 ;
      RECT 20.781 4.483 20.805 4.67 ;
      RECT 20.695 4.485 20.781 4.667 ;
      RECT 20.61 4.487 20.695 4.668 ;
      RECT 20.553 4.488 20.61 4.674 ;
      RECT 20.467 4.49 20.553 4.684 ;
      RECT 20.381 4.493 20.467 4.697 ;
      RECT 20.295 4.495 20.381 4.709 ;
      RECT 20.281 4.496 20.295 4.716 ;
      RECT 20.195 4.497 20.281 4.724 ;
      RECT 20.155 4.499 20.195 4.733 ;
      RECT 20.146 4.5 20.155 4.736 ;
      RECT 20.06 4.508 20.146 4.742 ;
      RECT 20.04 4.517 20.06 4.75 ;
      RECT 19.955 4.532 20.04 4.758 ;
      RECT 19.895 4.555 19.955 4.769 ;
      RECT 19.885 4.567 19.895 4.774 ;
      RECT 19.845 4.577 19.885 4.778 ;
      RECT 19.79 4.594 19.845 4.786 ;
      RECT 19.785 4.604 19.79 4.79 ;
      RECT 20.851 3.735 20.91 4.132 ;
      RECT 20.765 3.735 20.97 4.123 ;
      RECT 20.76 3.765 20.97 4.118 ;
      RECT 20.726 3.765 20.97 4.116 ;
      RECT 20.64 3.765 20.97 4.11 ;
      RECT 20.595 3.765 20.99 4.088 ;
      RECT 20.595 3.765 21.01 4.043 ;
      RECT 20.555 3.765 21.01 4.033 ;
      RECT 20.765 3.735 21.045 4.015 ;
      RECT 20.5 3.735 20.76 3.995 ;
      RECT 19.685 3.215 19.945 3.475 ;
      RECT 19.765 3.175 20.045 3.455 ;
      RECT 96.14 7.215 96.51 7.585 ;
      RECT 88.565 9.325 88.935 9.695 ;
      RECT 80.355 7.215 80.725 7.585 ;
      RECT 72.78 9.325 73.15 9.695 ;
      RECT 64.57 7.215 64.94 7.585 ;
      RECT 56.995 9.325 57.365 9.695 ;
      RECT 48.795 7.215 49.165 7.585 ;
      RECT 41.22 9.325 41.59 9.695 ;
      RECT 33.015 7.215 33.385 7.585 ;
      RECT 25.44 9.325 25.81 9.695 ;
    LAYER via1 ;
      RECT 96.3 9.65 96.45 9.8 ;
      RECT 96.25 7.325 96.4 7.475 ;
      RECT 93.93 9.025 94.08 9.175 ;
      RECT 93.915 3.36 94.065 3.51 ;
      RECT 93.125 3.745 93.275 3.895 ;
      RECT 93.125 8.61 93.275 8.76 ;
      RECT 91.48 2.735 91.63 2.885 ;
      RECT 91.165 4.255 91.315 4.405 ;
      RECT 90.265 3.585 90.415 3.735 ;
      RECT 89.315 9 89.465 9.15 ;
      RECT 89.065 3.85 89.215 4 ;
      RECT 88.73 4.57 88.88 4.72 ;
      RECT 88.675 9.435 88.825 9.585 ;
      RECT 88.65 3.41 88.8 3.56 ;
      RECT 87.215 3.805 87.365 3.955 ;
      RECT 86.45 3.655 86.6 3.805 ;
      RECT 86.195 3.25 86.345 3.4 ;
      RECT 85.575 4.015 85.725 4.165 ;
      RECT 85.195 3.485 85.345 3.635 ;
      RECT 85.18 4.525 85.33 4.675 ;
      RECT 84.65 3.79 84.8 3.94 ;
      RECT 84.49 4.51 84.64 4.66 ;
      RECT 83.68 3.79 83.83 3.94 ;
      RECT 82.865 3.27 83.015 3.42 ;
      RECT 82.705 4.655 82.855 4.805 ;
      RECT 82.47 4.31 82.62 4.46 ;
      RECT 82.425 3.7 82.575 3.85 ;
      RECT 81.425 4.32 81.575 4.47 ;
      RECT 80.49 9.045 80.64 9.195 ;
      RECT 80.465 7.325 80.615 7.475 ;
      RECT 78.145 9.025 78.295 9.175 ;
      RECT 78.13 3.36 78.28 3.51 ;
      RECT 77.34 3.745 77.49 3.895 ;
      RECT 77.34 8.61 77.49 8.76 ;
      RECT 75.695 2.735 75.845 2.885 ;
      RECT 75.38 4.255 75.53 4.405 ;
      RECT 74.48 3.585 74.63 3.735 ;
      RECT 73.53 8.99 73.68 9.14 ;
      RECT 73.28 3.85 73.43 4 ;
      RECT 72.945 4.57 73.095 4.72 ;
      RECT 72.89 9.435 73.04 9.585 ;
      RECT 72.865 3.41 73.015 3.56 ;
      RECT 71.43 3.805 71.58 3.955 ;
      RECT 70.665 3.655 70.815 3.805 ;
      RECT 70.41 3.25 70.56 3.4 ;
      RECT 69.79 4.015 69.94 4.165 ;
      RECT 69.41 3.485 69.56 3.635 ;
      RECT 69.395 4.525 69.545 4.675 ;
      RECT 68.865 3.79 69.015 3.94 ;
      RECT 68.705 4.51 68.855 4.66 ;
      RECT 67.895 3.79 68.045 3.94 ;
      RECT 67.08 3.27 67.23 3.42 ;
      RECT 66.92 4.655 67.07 4.805 ;
      RECT 66.685 4.31 66.835 4.46 ;
      RECT 66.64 3.7 66.79 3.85 ;
      RECT 65.64 4.32 65.79 4.47 ;
      RECT 64.705 9.045 64.855 9.195 ;
      RECT 64.68 7.325 64.83 7.475 ;
      RECT 62.36 9.025 62.51 9.175 ;
      RECT 62.345 3.36 62.495 3.51 ;
      RECT 61.555 3.745 61.705 3.895 ;
      RECT 61.555 8.61 61.705 8.76 ;
      RECT 59.91 2.735 60.06 2.885 ;
      RECT 59.595 4.255 59.745 4.405 ;
      RECT 58.695 3.585 58.845 3.735 ;
      RECT 57.8 9 57.95 9.15 ;
      RECT 57.495 3.85 57.645 4 ;
      RECT 57.16 4.57 57.31 4.72 ;
      RECT 57.105 9.435 57.255 9.585 ;
      RECT 57.08 3.41 57.23 3.56 ;
      RECT 55.645 3.805 55.795 3.955 ;
      RECT 54.88 3.655 55.03 3.805 ;
      RECT 54.625 3.25 54.775 3.4 ;
      RECT 54.005 4.015 54.155 4.165 ;
      RECT 53.625 3.485 53.775 3.635 ;
      RECT 53.61 4.525 53.76 4.675 ;
      RECT 53.08 3.79 53.23 3.94 ;
      RECT 52.92 4.51 53.07 4.66 ;
      RECT 52.11 3.79 52.26 3.94 ;
      RECT 51.295 3.27 51.445 3.42 ;
      RECT 51.135 4.655 51.285 4.805 ;
      RECT 50.9 4.31 51.05 4.46 ;
      RECT 50.855 3.7 51.005 3.85 ;
      RECT 49.855 4.32 50.005 4.47 ;
      RECT 48.975 9.045 49.125 9.195 ;
      RECT 48.905 7.325 49.055 7.475 ;
      RECT 46.585 9.025 46.735 9.175 ;
      RECT 46.57 3.36 46.72 3.51 ;
      RECT 45.78 3.745 45.93 3.895 ;
      RECT 45.78 8.61 45.93 8.76 ;
      RECT 44.135 2.735 44.285 2.885 ;
      RECT 43.82 4.255 43.97 4.405 ;
      RECT 42.92 3.585 43.07 3.735 ;
      RECT 42.02 9 42.17 9.15 ;
      RECT 41.72 3.85 41.87 4 ;
      RECT 41.385 4.57 41.535 4.72 ;
      RECT 41.33 9.435 41.48 9.585 ;
      RECT 41.305 3.41 41.455 3.56 ;
      RECT 39.87 3.805 40.02 3.955 ;
      RECT 39.105 3.655 39.255 3.805 ;
      RECT 38.85 3.25 39 3.4 ;
      RECT 38.23 4.015 38.38 4.165 ;
      RECT 37.85 3.485 38 3.635 ;
      RECT 37.835 4.525 37.985 4.675 ;
      RECT 37.305 3.79 37.455 3.94 ;
      RECT 37.145 4.51 37.295 4.66 ;
      RECT 36.335 3.79 36.485 3.94 ;
      RECT 35.52 3.27 35.67 3.42 ;
      RECT 35.36 4.655 35.51 4.805 ;
      RECT 35.125 4.31 35.275 4.46 ;
      RECT 35.08 3.7 35.23 3.85 ;
      RECT 34.08 4.32 34.23 4.47 ;
      RECT 33.195 9.045 33.345 9.195 ;
      RECT 33.125 7.325 33.275 7.475 ;
      RECT 30.805 9.025 30.955 9.175 ;
      RECT 30.79 3.36 30.94 3.51 ;
      RECT 30 3.745 30.15 3.895 ;
      RECT 30 8.61 30.15 8.76 ;
      RECT 28.355 2.735 28.505 2.885 ;
      RECT 28.04 4.255 28.19 4.405 ;
      RECT 27.14 3.585 27.29 3.735 ;
      RECT 26.21 8.99 26.36 9.14 ;
      RECT 25.94 3.85 26.09 4 ;
      RECT 25.605 4.57 25.755 4.72 ;
      RECT 25.55 9.435 25.7 9.585 ;
      RECT 25.525 3.41 25.675 3.56 ;
      RECT 24.09 3.805 24.24 3.955 ;
      RECT 23.325 3.655 23.475 3.805 ;
      RECT 23.07 3.25 23.22 3.4 ;
      RECT 22.45 4.015 22.6 4.165 ;
      RECT 22.07 3.485 22.22 3.635 ;
      RECT 22.055 4.525 22.205 4.675 ;
      RECT 21.525 3.79 21.675 3.94 ;
      RECT 21.365 4.51 21.515 4.66 ;
      RECT 20.555 3.79 20.705 3.94 ;
      RECT 19.74 3.27 19.89 3.42 ;
      RECT 19.58 4.655 19.73 4.805 ;
      RECT 19.345 4.31 19.495 4.46 ;
      RECT 19.3 3.7 19.45 3.85 ;
      RECT 18.3 4.32 18.45 4.47 ;
      RECT 16.615 9.38 16.765 9.53 ;
      RECT 16.24 8.64 16.39 8.79 ;
    LAYER met1 ;
      RECT 96.165 10.055 96.46 10.285 ;
      RECT 96.225 9.55 96.4 10.285 ;
      RECT 96.2 9.55 96.55 9.9 ;
      RECT 96.225 8.575 96.395 10.285 ;
      RECT 96.165 8.575 96.455 8.805 ;
      RECT 95.175 10.055 95.47 10.285 ;
      RECT 95.235 8.575 95.405 10.285 ;
      RECT 95.175 8.575 95.465 8.805 ;
      RECT 95.175 8.61 96.025 8.77 ;
      RECT 95.86 8.205 96.025 8.77 ;
      RECT 95.175 8.605 95.57 8.77 ;
      RECT 95.795 8.205 96.085 8.435 ;
      RECT 95.795 8.235 96.255 8.405 ;
      RECT 95.76 4.025 96.08 4.26 ;
      RECT 95.76 4.055 96.25 4.225 ;
      RECT 95.76 3.69 95.95 4.26 ;
      RECT 95.175 3.655 95.465 3.885 ;
      RECT 95.175 3.69 95.95 3.86 ;
      RECT 95.235 2.175 95.405 3.885 ;
      RECT 95.175 2.175 95.47 2.405 ;
      RECT 94.805 4.025 95.095 4.255 ;
      RECT 94.805 4.055 95.265 4.225 ;
      RECT 94.87 2.95 95.035 4.255 ;
      RECT 93.385 2.915 93.675 3.145 ;
      RECT 93.385 2.95 95.035 3.12 ;
      RECT 93.445 2.175 93.615 3.145 ;
      RECT 93.385 2.175 93.675 2.405 ;
      RECT 93.385 10.055 93.675 10.285 ;
      RECT 93.445 9.315 93.615 10.285 ;
      RECT 93.445 9.405 95.035 9.575 ;
      RECT 94.865 8.205 95.035 9.575 ;
      RECT 93.385 9.315 93.675 9.545 ;
      RECT 94.805 8.205 95.095 8.435 ;
      RECT 94.805 8.235 95.265 8.405 ;
      RECT 93.815 3.26 94.165 3.61 ;
      RECT 91.48 3.32 94.165 3.49 ;
      RECT 93.645 3.315 94.165 3.49 ;
      RECT 91.48 2.635 91.65 3.49 ;
      RECT 91.38 2.635 91.73 2.985 ;
      RECT 93.84 8.94 94.165 9.265 ;
      RECT 89.215 8.9 89.565 9.25 ;
      RECT 93.815 8.945 94.165 9.175 ;
      RECT 89.035 8.945 89.565 9.175 ;
      RECT 93.645 8.97 94.165 9.145 ;
      RECT 88.865 8.975 89.565 9.145 ;
      RECT 89.035 8.97 94.165 9.14 ;
      RECT 93.04 3.66 93.36 3.98 ;
      RECT 93.015 3.655 93.305 3.885 ;
      RECT 92.94 3.685 93.36 3.86 ;
      RECT 92.84 3.685 93.36 3.855 ;
      RECT 93.04 8.54 93.36 8.83 ;
      RECT 93.015 8.575 93.36 8.805 ;
      RECT 92.84 8.605 93.36 8.775 ;
      RECT 89.675 3.76 89.86 3.97 ;
      RECT 89.665 3.765 89.875 3.963 ;
      RECT 89.665 3.765 89.961 3.94 ;
      RECT 89.665 3.765 90.02 3.915 ;
      RECT 89.665 3.765 90.075 3.895 ;
      RECT 89.665 3.765 90.085 3.883 ;
      RECT 89.665 3.765 90.28 3.822 ;
      RECT 89.665 3.765 90.31 3.805 ;
      RECT 89.665 3.765 90.33 3.795 ;
      RECT 90.21 3.53 90.47 3.79 ;
      RECT 90.195 3.62 90.21 3.837 ;
      RECT 89.73 3.752 90.47 3.79 ;
      RECT 90.181 3.631 90.195 3.843 ;
      RECT 89.77 3.745 90.47 3.79 ;
      RECT 90.095 3.671 90.181 3.862 ;
      RECT 90.02 3.732 90.47 3.79 ;
      RECT 90.09 3.707 90.095 3.879 ;
      RECT 90.075 3.717 90.47 3.79 ;
      RECT 90.085 3.712 90.09 3.881 ;
      RECT 89.01 3.795 89.115 4.055 ;
      RECT 89.825 3.32 89.83 3.545 ;
      RECT 89.955 3.32 90.01 3.53 ;
      RECT 90.01 3.325 90.02 3.523 ;
      RECT 89.916 3.32 89.955 3.533 ;
      RECT 89.83 3.32 89.916 3.54 ;
      RECT 89.81 3.325 89.825 3.546 ;
      RECT 89.8 3.365 89.81 3.548 ;
      RECT 89.77 3.375 89.8 3.55 ;
      RECT 89.765 3.38 89.77 3.552 ;
      RECT 89.74 3.385 89.765 3.554 ;
      RECT 89.725 3.39 89.74 3.556 ;
      RECT 89.71 3.392 89.725 3.558 ;
      RECT 89.705 3.397 89.71 3.56 ;
      RECT 89.655 3.405 89.705 3.563 ;
      RECT 89.63 3.414 89.655 3.568 ;
      RECT 89.62 3.421 89.63 3.573 ;
      RECT 89.615 3.424 89.62 3.577 ;
      RECT 89.595 3.427 89.615 3.586 ;
      RECT 89.565 3.435 89.595 3.606 ;
      RECT 89.536 3.448 89.565 3.628 ;
      RECT 89.45 3.482 89.536 3.672 ;
      RECT 89.445 3.508 89.45 3.71 ;
      RECT 89.44 3.512 89.445 3.719 ;
      RECT 89.405 3.525 89.44 3.752 ;
      RECT 89.395 3.539 89.405 3.79 ;
      RECT 89.39 3.543 89.395 3.803 ;
      RECT 89.385 3.547 89.39 3.808 ;
      RECT 89.375 3.555 89.385 3.82 ;
      RECT 89.37 3.562 89.375 3.835 ;
      RECT 89.345 3.575 89.37 3.86 ;
      RECT 89.305 3.604 89.345 3.915 ;
      RECT 89.29 3.629 89.305 3.97 ;
      RECT 89.28 3.64 89.29 3.993 ;
      RECT 89.275 3.647 89.28 4.005 ;
      RECT 89.27 3.651 89.275 4.013 ;
      RECT 89.215 3.679 89.27 4.055 ;
      RECT 89.195 3.715 89.215 4.055 ;
      RECT 89.18 3.73 89.195 4.055 ;
      RECT 89.125 3.762 89.18 4.055 ;
      RECT 89.115 3.792 89.125 4.055 ;
      RECT 88.725 3.407 88.91 3.645 ;
      RECT 88.71 3.409 88.92 3.64 ;
      RECT 88.595 3.355 88.855 3.615 ;
      RECT 88.59 3.392 88.855 3.569 ;
      RECT 88.585 3.402 88.855 3.566 ;
      RECT 88.58 3.442 88.92 3.56 ;
      RECT 88.575 3.475 88.92 3.55 ;
      RECT 88.585 3.417 88.935 3.488 ;
      RECT 88.882 4.515 88.895 5.045 ;
      RECT 88.796 4.515 88.895 5.044 ;
      RECT 88.796 4.515 88.9 5.043 ;
      RECT 88.71 4.515 88.9 5.041 ;
      RECT 88.705 4.515 88.9 5.038 ;
      RECT 88.705 4.515 88.91 5.036 ;
      RECT 88.7 4.807 88.91 5.033 ;
      RECT 88.7 4.817 88.915 5.03 ;
      RECT 88.7 4.885 88.92 5.026 ;
      RECT 88.69 4.89 88.92 5.025 ;
      RECT 88.69 4.982 88.925 5.022 ;
      RECT 88.675 4.515 88.935 4.775 ;
      RECT 88.605 10.055 88.895 10.285 ;
      RECT 88.665 9.315 88.835 10.285 ;
      RECT 88.58 9.34 88.92 9.685 ;
      RECT 88.605 9.315 88.895 9.685 ;
      RECT 87.905 3.505 87.95 5.04 ;
      RECT 88.105 3.505 88.135 3.72 ;
      RECT 86.48 3.245 86.6 3.455 ;
      RECT 86.14 3.195 86.4 3.455 ;
      RECT 86.14 3.24 86.435 3.445 ;
      RECT 88.145 3.521 88.15 3.575 ;
      RECT 88.14 3.514 88.145 3.708 ;
      RECT 88.135 3.508 88.14 3.715 ;
      RECT 88.09 3.505 88.105 3.728 ;
      RECT 88.085 3.505 88.09 3.75 ;
      RECT 88.08 3.505 88.085 3.798 ;
      RECT 88.075 3.505 88.08 3.818 ;
      RECT 88.065 3.505 88.075 3.925 ;
      RECT 88.06 3.505 88.065 3.988 ;
      RECT 88.055 3.505 88.06 4.045 ;
      RECT 88.05 3.505 88.055 4.053 ;
      RECT 88.035 3.505 88.05 4.16 ;
      RECT 88.025 3.505 88.035 4.295 ;
      RECT 88.015 3.505 88.025 4.405 ;
      RECT 88.005 3.505 88.015 4.462 ;
      RECT 88 3.505 88.005 4.502 ;
      RECT 87.995 3.505 88 4.538 ;
      RECT 87.985 3.505 87.995 4.578 ;
      RECT 87.98 3.505 87.985 4.62 ;
      RECT 87.96 3.505 87.98 4.685 ;
      RECT 87.965 4.83 87.97 5.01 ;
      RECT 87.96 4.812 87.965 5.018 ;
      RECT 87.955 3.505 87.96 4.748 ;
      RECT 87.955 4.792 87.96 5.025 ;
      RECT 87.95 3.505 87.955 5.035 ;
      RECT 87.895 3.505 87.905 3.805 ;
      RECT 87.9 4.052 87.905 5.04 ;
      RECT 87.895 4.117 87.9 5.04 ;
      RECT 87.89 3.506 87.895 3.795 ;
      RECT 87.885 4.182 87.895 5.04 ;
      RECT 87.88 3.507 87.89 3.785 ;
      RECT 87.87 4.295 87.885 5.04 ;
      RECT 87.875 3.508 87.88 3.775 ;
      RECT 87.855 3.509 87.875 3.753 ;
      RECT 87.86 4.392 87.87 5.04 ;
      RECT 87.855 4.467 87.86 5.04 ;
      RECT 87.845 3.508 87.855 3.73 ;
      RECT 87.85 4.51 87.855 5.04 ;
      RECT 87.845 4.537 87.85 5.04 ;
      RECT 87.835 3.506 87.845 3.718 ;
      RECT 87.84 4.58 87.845 5.04 ;
      RECT 87.835 4.607 87.84 5.04 ;
      RECT 87.825 3.505 87.835 3.705 ;
      RECT 87.83 4.622 87.835 5.04 ;
      RECT 87.79 4.68 87.83 5.04 ;
      RECT 87.82 3.504 87.825 3.69 ;
      RECT 87.815 3.502 87.82 3.683 ;
      RECT 87.805 3.499 87.815 3.673 ;
      RECT 87.8 3.496 87.805 3.658 ;
      RECT 87.785 3.492 87.8 3.651 ;
      RECT 87.78 4.735 87.79 5.04 ;
      RECT 87.78 3.489 87.785 3.646 ;
      RECT 87.765 3.485 87.78 3.64 ;
      RECT 87.775 4.752 87.78 5.04 ;
      RECT 87.765 4.815 87.775 5.04 ;
      RECT 87.685 3.47 87.765 3.62 ;
      RECT 87.76 4.822 87.765 5.035 ;
      RECT 87.755 4.83 87.76 5.025 ;
      RECT 87.675 3.456 87.685 3.604 ;
      RECT 87.66 3.452 87.675 3.602 ;
      RECT 87.65 3.447 87.66 3.598 ;
      RECT 87.625 3.44 87.65 3.59 ;
      RECT 87.62 3.435 87.625 3.585 ;
      RECT 87.61 3.435 87.62 3.583 ;
      RECT 87.6 3.433 87.61 3.581 ;
      RECT 87.57 3.425 87.6 3.575 ;
      RECT 87.555 3.417 87.57 3.568 ;
      RECT 87.535 3.412 87.555 3.561 ;
      RECT 87.53 3.408 87.535 3.556 ;
      RECT 87.5 3.401 87.53 3.55 ;
      RECT 87.475 3.392 87.5 3.54 ;
      RECT 87.445 3.385 87.475 3.532 ;
      RECT 87.42 3.375 87.445 3.523 ;
      RECT 87.405 3.367 87.42 3.517 ;
      RECT 87.38 3.362 87.405 3.512 ;
      RECT 87.37 3.358 87.38 3.507 ;
      RECT 87.35 3.353 87.37 3.502 ;
      RECT 87.315 3.348 87.35 3.495 ;
      RECT 87.255 3.343 87.315 3.488 ;
      RECT 87.242 3.339 87.255 3.486 ;
      RECT 87.156 3.334 87.242 3.483 ;
      RECT 87.07 3.324 87.156 3.479 ;
      RECT 87.029 3.317 87.07 3.476 ;
      RECT 86.943 3.31 87.029 3.473 ;
      RECT 86.857 3.3 86.943 3.469 ;
      RECT 86.771 3.29 86.857 3.464 ;
      RECT 86.685 3.28 86.771 3.46 ;
      RECT 86.675 3.265 86.685 3.458 ;
      RECT 86.665 3.25 86.675 3.458 ;
      RECT 86.6 3.245 86.665 3.457 ;
      RECT 86.435 3.242 86.48 3.45 ;
      RECT 87.68 4.147 87.685 4.338 ;
      RECT 87.675 4.142 87.68 4.345 ;
      RECT 87.661 4.14 87.675 4.351 ;
      RECT 87.575 4.14 87.661 4.353 ;
      RECT 87.571 4.14 87.575 4.356 ;
      RECT 87.485 4.14 87.571 4.374 ;
      RECT 87.475 4.145 87.485 4.393 ;
      RECT 87.465 4.2 87.475 4.397 ;
      RECT 87.44 4.215 87.465 4.404 ;
      RECT 87.4 4.235 87.44 4.417 ;
      RECT 87.395 4.247 87.4 4.427 ;
      RECT 87.38 4.253 87.395 4.432 ;
      RECT 87.375 4.258 87.38 4.436 ;
      RECT 87.355 4.265 87.375 4.441 ;
      RECT 87.285 4.29 87.355 4.458 ;
      RECT 87.245 4.318 87.285 4.478 ;
      RECT 87.24 4.328 87.245 4.486 ;
      RECT 87.22 4.335 87.24 4.488 ;
      RECT 87.215 4.342 87.22 4.491 ;
      RECT 87.185 4.35 87.215 4.494 ;
      RECT 87.18 4.355 87.185 4.498 ;
      RECT 87.106 4.359 87.18 4.506 ;
      RECT 87.02 4.368 87.106 4.522 ;
      RECT 87.016 4.373 87.02 4.531 ;
      RECT 86.93 4.378 87.016 4.541 ;
      RECT 86.89 4.386 86.93 4.553 ;
      RECT 86.84 4.392 86.89 4.56 ;
      RECT 86.755 4.401 86.84 4.575 ;
      RECT 86.68 4.412 86.755 4.593 ;
      RECT 86.645 4.419 86.68 4.603 ;
      RECT 86.57 4.427 86.645 4.608 ;
      RECT 86.515 4.436 86.57 4.608 ;
      RECT 86.49 4.441 86.515 4.606 ;
      RECT 86.48 4.444 86.49 4.604 ;
      RECT 86.445 4.446 86.48 4.602 ;
      RECT 86.415 4.448 86.445 4.598 ;
      RECT 86.37 4.447 86.415 4.594 ;
      RECT 86.35 4.442 86.37 4.591 ;
      RECT 86.3 4.427 86.35 4.588 ;
      RECT 86.29 4.412 86.3 4.583 ;
      RECT 86.24 4.397 86.29 4.573 ;
      RECT 86.19 4.372 86.24 4.553 ;
      RECT 86.18 4.357 86.19 4.535 ;
      RECT 86.175 4.355 86.18 4.529 ;
      RECT 86.155 4.35 86.175 4.524 ;
      RECT 86.15 4.342 86.155 4.518 ;
      RECT 86.135 4.336 86.15 4.511 ;
      RECT 86.13 4.331 86.135 4.503 ;
      RECT 86.11 4.326 86.13 4.495 ;
      RECT 86.095 4.319 86.11 4.488 ;
      RECT 86.08 4.313 86.095 4.479 ;
      RECT 86.075 4.307 86.08 4.472 ;
      RECT 86.03 4.282 86.075 4.458 ;
      RECT 86.015 4.252 86.03 4.44 ;
      RECT 86 4.235 86.015 4.431 ;
      RECT 85.975 4.215 86 4.419 ;
      RECT 85.935 4.185 85.975 4.399 ;
      RECT 85.925 4.155 85.935 4.384 ;
      RECT 85.91 4.145 85.925 4.377 ;
      RECT 85.855 4.11 85.91 4.356 ;
      RECT 85.84 4.073 85.855 4.335 ;
      RECT 85.83 4.06 85.84 4.327 ;
      RECT 85.78 4.03 85.83 4.309 ;
      RECT 85.765 3.96 85.78 4.29 ;
      RECT 85.72 3.96 85.765 4.273 ;
      RECT 85.695 3.96 85.72 4.255 ;
      RECT 85.685 3.96 85.695 4.248 ;
      RECT 85.606 3.96 85.685 4.241 ;
      RECT 85.52 3.96 85.606 4.233 ;
      RECT 85.505 3.992 85.52 4.228 ;
      RECT 85.43 4.002 85.505 4.224 ;
      RECT 85.41 4.012 85.43 4.219 ;
      RECT 85.385 4.012 85.41 4.216 ;
      RECT 85.375 4.002 85.385 4.215 ;
      RECT 85.365 3.975 85.375 4.214 ;
      RECT 85.325 3.97 85.365 4.212 ;
      RECT 85.28 3.97 85.325 4.208 ;
      RECT 85.255 3.97 85.28 4.203 ;
      RECT 85.205 3.97 85.255 4.19 ;
      RECT 85.165 3.975 85.175 4.175 ;
      RECT 85.175 3.97 85.205 4.18 ;
      RECT 87.16 3.75 87.42 4.01 ;
      RECT 87.155 3.772 87.42 3.968 ;
      RECT 86.395 3.6 86.615 3.965 ;
      RECT 86.377 3.687 86.615 3.964 ;
      RECT 86.36 3.692 86.615 3.961 ;
      RECT 86.36 3.692 86.635 3.96 ;
      RECT 86.33 3.702 86.635 3.958 ;
      RECT 86.325 3.717 86.635 3.954 ;
      RECT 86.325 3.717 86.64 3.953 ;
      RECT 86.32 3.775 86.64 3.951 ;
      RECT 86.32 3.775 86.65 3.948 ;
      RECT 86.315 3.84 86.65 3.943 ;
      RECT 86.395 3.6 86.655 3.86 ;
      RECT 85.14 3.43 85.4 3.69 ;
      RECT 85.14 3.473 85.486 3.664 ;
      RECT 85.14 3.473 85.53 3.663 ;
      RECT 85.14 3.473 85.55 3.661 ;
      RECT 85.14 3.473 85.65 3.66 ;
      RECT 85.14 3.473 85.67 3.658 ;
      RECT 85.14 3.473 85.68 3.653 ;
      RECT 85.55 3.44 85.74 3.65 ;
      RECT 85.55 3.442 85.745 3.648 ;
      RECT 85.54 3.447 85.75 3.64 ;
      RECT 85.486 3.471 85.75 3.64 ;
      RECT 85.53 3.465 85.54 3.662 ;
      RECT 85.54 3.445 85.745 3.648 ;
      RECT 84.495 4.505 84.7 4.735 ;
      RECT 84.435 4.455 84.49 4.715 ;
      RECT 84.495 4.455 84.695 4.735 ;
      RECT 85.465 4.77 85.47 4.797 ;
      RECT 85.455 4.68 85.465 4.802 ;
      RECT 85.45 4.602 85.455 4.808 ;
      RECT 85.44 4.592 85.45 4.815 ;
      RECT 85.435 4.582 85.44 4.821 ;
      RECT 85.425 4.577 85.435 4.823 ;
      RECT 85.41 4.569 85.425 4.831 ;
      RECT 85.395 4.56 85.41 4.843 ;
      RECT 85.385 4.552 85.395 4.853 ;
      RECT 85.35 4.47 85.385 4.871 ;
      RECT 85.315 4.47 85.35 4.89 ;
      RECT 85.3 4.47 85.315 4.898 ;
      RECT 85.245 4.47 85.3 4.898 ;
      RECT 85.211 4.47 85.245 4.889 ;
      RECT 85.125 4.47 85.211 4.865 ;
      RECT 85.115 4.53 85.125 4.847 ;
      RECT 85.075 4.532 85.115 4.838 ;
      RECT 85.07 4.534 85.075 4.828 ;
      RECT 85.05 4.536 85.07 4.823 ;
      RECT 85.04 4.539 85.05 4.818 ;
      RECT 85.03 4.54 85.04 4.813 ;
      RECT 85.006 4.541 85.03 4.805 ;
      RECT 84.92 4.546 85.006 4.783 ;
      RECT 84.865 4.545 84.92 4.756 ;
      RECT 84.85 4.538 84.865 4.743 ;
      RECT 84.815 4.533 84.85 4.739 ;
      RECT 84.76 4.525 84.815 4.738 ;
      RECT 84.7 4.512 84.76 4.736 ;
      RECT 84.49 4.455 84.495 4.723 ;
      RECT 84.565 3.825 84.75 4.035 ;
      RECT 84.555 3.83 84.765 4.028 ;
      RECT 84.595 3.735 84.855 3.995 ;
      RECT 84.55 3.892 84.855 3.918 ;
      RECT 83.895 3.685 83.9 4.485 ;
      RECT 83.84 3.735 83.87 4.485 ;
      RECT 83.83 3.735 83.835 4.045 ;
      RECT 83.815 3.735 83.82 4.04 ;
      RECT 83.36 3.78 83.375 3.995 ;
      RECT 83.29 3.78 83.375 3.99 ;
      RECT 84.555 3.36 84.625 3.57 ;
      RECT 84.625 3.367 84.635 3.565 ;
      RECT 84.521 3.36 84.555 3.577 ;
      RECT 84.435 3.36 84.521 3.601 ;
      RECT 84.425 3.365 84.435 3.62 ;
      RECT 84.42 3.377 84.425 3.623 ;
      RECT 84.405 3.392 84.42 3.627 ;
      RECT 84.4 3.41 84.405 3.631 ;
      RECT 84.36 3.42 84.4 3.64 ;
      RECT 84.345 3.427 84.36 3.652 ;
      RECT 84.33 3.432 84.345 3.657 ;
      RECT 84.315 3.435 84.33 3.662 ;
      RECT 84.305 3.437 84.315 3.666 ;
      RECT 84.27 3.444 84.305 3.674 ;
      RECT 84.235 3.452 84.27 3.688 ;
      RECT 84.225 3.458 84.235 3.697 ;
      RECT 84.22 3.46 84.225 3.699 ;
      RECT 84.2 3.463 84.22 3.705 ;
      RECT 84.17 3.47 84.2 3.716 ;
      RECT 84.16 3.476 84.17 3.723 ;
      RECT 84.135 3.479 84.16 3.73 ;
      RECT 84.125 3.483 84.135 3.738 ;
      RECT 84.12 3.484 84.125 3.76 ;
      RECT 84.115 3.485 84.12 3.775 ;
      RECT 84.11 3.486 84.115 3.79 ;
      RECT 84.105 3.487 84.11 3.805 ;
      RECT 84.1 3.488 84.105 3.835 ;
      RECT 84.09 3.49 84.1 3.868 ;
      RECT 84.075 3.494 84.09 3.915 ;
      RECT 84.065 3.497 84.075 3.96 ;
      RECT 84.06 3.5 84.065 3.988 ;
      RECT 84.05 3.502 84.06 4.015 ;
      RECT 84.045 3.505 84.05 4.05 ;
      RECT 84.015 3.51 84.045 4.108 ;
      RECT 84.01 3.515 84.015 4.193 ;
      RECT 84.005 3.517 84.01 4.228 ;
      RECT 84 3.519 84.005 4.31 ;
      RECT 83.995 3.521 84 4.398 ;
      RECT 83.985 3.523 83.995 4.48 ;
      RECT 83.97 3.537 83.985 4.485 ;
      RECT 83.935 3.582 83.97 4.485 ;
      RECT 83.925 3.622 83.935 4.485 ;
      RECT 83.91 3.65 83.925 4.485 ;
      RECT 83.905 3.667 83.91 4.485 ;
      RECT 83.9 3.675 83.905 4.485 ;
      RECT 83.89 3.69 83.895 4.485 ;
      RECT 83.885 3.697 83.89 4.485 ;
      RECT 83.875 3.717 83.885 4.485 ;
      RECT 83.87 3.73 83.875 4.485 ;
      RECT 83.835 3.735 83.84 4.07 ;
      RECT 83.82 4.125 83.84 4.485 ;
      RECT 83.82 3.735 83.83 4.043 ;
      RECT 83.815 4.165 83.82 4.485 ;
      RECT 83.765 3.735 83.815 4.038 ;
      RECT 83.81 4.202 83.815 4.485 ;
      RECT 83.8 4.225 83.81 4.485 ;
      RECT 83.795 4.27 83.8 4.485 ;
      RECT 83.785 4.28 83.795 4.478 ;
      RECT 83.711 3.735 83.765 4.032 ;
      RECT 83.625 3.735 83.711 4.025 ;
      RECT 83.576 3.782 83.625 4.018 ;
      RECT 83.49 3.79 83.576 4.011 ;
      RECT 83.475 3.787 83.49 4.006 ;
      RECT 83.461 3.78 83.475 4.005 ;
      RECT 83.375 3.78 83.461 4 ;
      RECT 83.28 3.785 83.29 3.985 ;
      RECT 82.87 3.215 82.885 3.615 ;
      RECT 83.065 3.215 83.07 3.475 ;
      RECT 82.81 3.215 82.855 3.475 ;
      RECT 83.265 4.52 83.27 4.725 ;
      RECT 83.26 4.51 83.265 4.73 ;
      RECT 83.255 4.497 83.26 4.735 ;
      RECT 83.25 4.477 83.255 4.735 ;
      RECT 83.225 4.43 83.25 4.735 ;
      RECT 83.19 4.345 83.225 4.735 ;
      RECT 83.185 4.282 83.19 4.735 ;
      RECT 83.18 4.267 83.185 4.735 ;
      RECT 83.165 4.227 83.18 4.735 ;
      RECT 83.16 4.202 83.165 4.735 ;
      RECT 83.15 4.185 83.16 4.735 ;
      RECT 83.115 4.107 83.15 4.735 ;
      RECT 83.11 4.05 83.115 4.735 ;
      RECT 83.105 4.037 83.11 4.735 ;
      RECT 83.095 4.015 83.105 4.735 ;
      RECT 83.085 3.98 83.095 4.735 ;
      RECT 83.075 3.95 83.085 4.735 ;
      RECT 83.065 3.865 83.075 4.378 ;
      RECT 83.072 4.51 83.075 4.735 ;
      RECT 83.07 4.52 83.072 4.735 ;
      RECT 83.06 4.53 83.07 4.73 ;
      RECT 83.055 3.215 83.065 3.61 ;
      RECT 83.06 3.742 83.065 4.353 ;
      RECT 83.055 3.64 83.06 4.336 ;
      RECT 83.045 3.215 83.055 4.312 ;
      RECT 83.04 3.215 83.045 4.283 ;
      RECT 83.035 3.215 83.04 4.273 ;
      RECT 83.015 3.215 83.035 4.235 ;
      RECT 83.01 3.215 83.015 4.193 ;
      RECT 83.005 3.215 83.01 4.173 ;
      RECT 82.975 3.215 83.005 4.123 ;
      RECT 82.965 3.215 82.975 4.07 ;
      RECT 82.96 3.215 82.965 4.043 ;
      RECT 82.955 3.215 82.96 4.028 ;
      RECT 82.945 3.215 82.955 4.005 ;
      RECT 82.935 3.215 82.945 3.98 ;
      RECT 82.93 3.215 82.935 3.92 ;
      RECT 82.92 3.215 82.93 3.858 ;
      RECT 82.915 3.215 82.92 3.778 ;
      RECT 82.91 3.215 82.915 3.743 ;
      RECT 82.905 3.215 82.91 3.718 ;
      RECT 82.9 3.215 82.905 3.703 ;
      RECT 82.895 3.215 82.9 3.673 ;
      RECT 82.89 3.215 82.895 3.65 ;
      RECT 82.885 3.215 82.89 3.623 ;
      RECT 82.855 3.215 82.87 3.61 ;
      RECT 82.01 4.75 82.195 4.96 ;
      RECT 82 4.755 82.21 4.953 ;
      RECT 82 4.755 82.23 4.925 ;
      RECT 82 4.755 82.245 4.904 ;
      RECT 82 4.755 82.26 4.902 ;
      RECT 82 4.755 82.27 4.901 ;
      RECT 82 4.755 82.3 4.898 ;
      RECT 82.65 4.6 82.91 4.86 ;
      RECT 82.61 4.647 82.91 4.843 ;
      RECT 82.601 4.655 82.61 4.846 ;
      RECT 82.195 4.748 82.91 4.843 ;
      RECT 82.515 4.673 82.601 4.853 ;
      RECT 82.21 4.745 82.91 4.843 ;
      RECT 82.456 4.695 82.515 4.865 ;
      RECT 82.23 4.741 82.91 4.843 ;
      RECT 82.37 4.707 82.456 4.876 ;
      RECT 82.245 4.737 82.91 4.843 ;
      RECT 82.315 4.72 82.37 4.888 ;
      RECT 82.26 4.735 82.91 4.843 ;
      RECT 82.3 4.726 82.315 4.894 ;
      RECT 82.27 4.731 82.91 4.843 ;
      RECT 82.415 4.255 82.675 4.515 ;
      RECT 82.415 4.275 82.785 4.485 ;
      RECT 82.415 4.28 82.795 4.48 ;
      RECT 82.606 3.694 82.685 3.925 ;
      RECT 82.52 3.697 82.735 3.92 ;
      RECT 82.515 3.697 82.735 3.915 ;
      RECT 82.515 3.702 82.745 3.913 ;
      RECT 82.49 3.702 82.745 3.91 ;
      RECT 82.49 3.71 82.755 3.908 ;
      RECT 82.37 3.645 82.63 3.905 ;
      RECT 82.37 3.692 82.68 3.905 ;
      RECT 81.625 4.265 81.63 4.525 ;
      RECT 81.455 4.035 81.46 4.525 ;
      RECT 81.34 4.275 81.345 4.5 ;
      RECT 82.05 3.37 82.055 3.58 ;
      RECT 82.055 3.375 82.07 3.575 ;
      RECT 81.99 3.37 82.05 3.588 ;
      RECT 81.975 3.37 81.99 3.598 ;
      RECT 81.925 3.37 81.975 3.615 ;
      RECT 81.905 3.37 81.925 3.638 ;
      RECT 81.89 3.37 81.905 3.65 ;
      RECT 81.87 3.37 81.89 3.66 ;
      RECT 81.86 3.375 81.87 3.669 ;
      RECT 81.855 3.385 81.86 3.674 ;
      RECT 81.85 3.397 81.855 3.678 ;
      RECT 81.84 3.42 81.85 3.683 ;
      RECT 81.835 3.435 81.84 3.687 ;
      RECT 81.83 3.452 81.835 3.69 ;
      RECT 81.825 3.46 81.83 3.693 ;
      RECT 81.815 3.465 81.825 3.697 ;
      RECT 81.81 3.472 81.815 3.702 ;
      RECT 81.8 3.477 81.81 3.706 ;
      RECT 81.775 3.489 81.8 3.717 ;
      RECT 81.755 3.506 81.775 3.733 ;
      RECT 81.73 3.523 81.755 3.755 ;
      RECT 81.695 3.546 81.73 3.813 ;
      RECT 81.675 3.568 81.695 3.875 ;
      RECT 81.67 3.578 81.675 3.91 ;
      RECT 81.66 3.585 81.67 3.948 ;
      RECT 81.655 3.592 81.66 3.968 ;
      RECT 81.65 3.603 81.655 4.005 ;
      RECT 81.645 3.611 81.65 4.07 ;
      RECT 81.635 3.622 81.645 4.123 ;
      RECT 81.63 3.64 81.635 4.193 ;
      RECT 81.625 3.65 81.63 4.23 ;
      RECT 81.62 3.66 81.625 4.525 ;
      RECT 81.615 3.672 81.62 4.525 ;
      RECT 81.61 3.682 81.615 4.525 ;
      RECT 81.6 3.692 81.61 4.525 ;
      RECT 81.59 3.715 81.6 4.525 ;
      RECT 81.575 3.75 81.59 4.525 ;
      RECT 81.535 3.812 81.575 4.525 ;
      RECT 81.53 3.865 81.535 4.525 ;
      RECT 81.505 3.9 81.53 4.525 ;
      RECT 81.49 3.945 81.505 4.525 ;
      RECT 81.485 3.967 81.49 4.525 ;
      RECT 81.475 3.98 81.485 4.525 ;
      RECT 81.465 4.005 81.475 4.525 ;
      RECT 81.46 4.027 81.465 4.525 ;
      RECT 81.435 4.065 81.455 4.525 ;
      RECT 81.395 4.122 81.435 4.525 ;
      RECT 81.39 4.172 81.395 4.525 ;
      RECT 81.385 4.19 81.39 4.525 ;
      RECT 81.38 4.202 81.385 4.525 ;
      RECT 81.37 4.22 81.38 4.525 ;
      RECT 81.36 4.24 81.37 4.5 ;
      RECT 81.355 4.257 81.36 4.5 ;
      RECT 81.345 4.27 81.355 4.5 ;
      RECT 81.315 4.28 81.34 4.5 ;
      RECT 81.305 4.287 81.315 4.5 ;
      RECT 81.29 4.297 81.305 4.495 ;
      RECT 80.38 10.055 80.675 10.285 ;
      RECT 80.44 8.575 80.61 10.285 ;
      RECT 80.39 8.945 80.74 9.295 ;
      RECT 80.38 8.575 80.67 8.805 ;
      RECT 79.39 10.055 79.685 10.285 ;
      RECT 79.45 8.575 79.62 10.285 ;
      RECT 79.39 8.575 79.68 8.805 ;
      RECT 79.39 8.61 80.24 8.77 ;
      RECT 80.075 8.205 80.24 8.77 ;
      RECT 79.39 8.605 79.785 8.77 ;
      RECT 80.01 8.205 80.3 8.435 ;
      RECT 80.01 8.235 80.47 8.405 ;
      RECT 79.975 4.025 80.295 4.26 ;
      RECT 79.975 4.055 80.465 4.225 ;
      RECT 79.975 3.69 80.165 4.26 ;
      RECT 79.39 3.655 79.68 3.885 ;
      RECT 79.39 3.69 80.165 3.86 ;
      RECT 79.45 2.175 79.62 3.885 ;
      RECT 79.39 2.175 79.685 2.405 ;
      RECT 79.02 4.025 79.31 4.255 ;
      RECT 79.02 4.055 79.48 4.225 ;
      RECT 79.085 2.95 79.25 4.255 ;
      RECT 77.6 2.915 77.89 3.145 ;
      RECT 77.6 2.95 79.25 3.12 ;
      RECT 77.66 2.175 77.83 3.145 ;
      RECT 77.6 2.175 77.89 2.405 ;
      RECT 77.6 10.055 77.89 10.285 ;
      RECT 77.66 9.315 77.83 10.285 ;
      RECT 77.66 9.405 79.25 9.575 ;
      RECT 79.08 8.205 79.25 9.575 ;
      RECT 77.6 9.315 77.89 9.545 ;
      RECT 79.02 8.205 79.31 8.435 ;
      RECT 79.02 8.235 79.48 8.405 ;
      RECT 78.03 3.26 78.38 3.61 ;
      RECT 75.695 3.32 78.38 3.49 ;
      RECT 77.86 3.315 78.38 3.49 ;
      RECT 75.695 2.635 75.865 3.49 ;
      RECT 75.595 2.635 75.945 2.985 ;
      RECT 78.055 8.94 78.38 9.265 ;
      RECT 73.43 8.89 73.78 9.24 ;
      RECT 78.03 8.945 78.38 9.175 ;
      RECT 73.25 8.945 73.78 9.175 ;
      RECT 77.86 8.97 78.38 9.145 ;
      RECT 73.08 8.975 73.78 9.145 ;
      RECT 73.25 8.97 78.38 9.14 ;
      RECT 77.255 3.66 77.575 3.98 ;
      RECT 77.23 3.655 77.52 3.885 ;
      RECT 77.155 3.685 77.575 3.86 ;
      RECT 77.055 3.685 77.575 3.855 ;
      RECT 77.255 8.54 77.575 8.83 ;
      RECT 77.23 8.575 77.575 8.805 ;
      RECT 77.055 8.605 77.575 8.775 ;
      RECT 73.89 3.76 74.075 3.97 ;
      RECT 73.88 3.765 74.09 3.963 ;
      RECT 73.88 3.765 74.176 3.94 ;
      RECT 73.88 3.765 74.235 3.915 ;
      RECT 73.88 3.765 74.29 3.895 ;
      RECT 73.88 3.765 74.3 3.883 ;
      RECT 73.88 3.765 74.495 3.822 ;
      RECT 73.88 3.765 74.525 3.805 ;
      RECT 73.88 3.765 74.545 3.795 ;
      RECT 74.425 3.53 74.685 3.79 ;
      RECT 74.41 3.62 74.425 3.837 ;
      RECT 73.945 3.752 74.685 3.79 ;
      RECT 74.396 3.631 74.41 3.843 ;
      RECT 73.985 3.745 74.685 3.79 ;
      RECT 74.31 3.671 74.396 3.862 ;
      RECT 74.235 3.732 74.685 3.79 ;
      RECT 74.305 3.707 74.31 3.879 ;
      RECT 74.29 3.717 74.685 3.79 ;
      RECT 74.3 3.712 74.305 3.881 ;
      RECT 73.225 3.795 73.33 4.055 ;
      RECT 74.04 3.32 74.045 3.545 ;
      RECT 74.17 3.32 74.225 3.53 ;
      RECT 74.225 3.325 74.235 3.523 ;
      RECT 74.131 3.32 74.17 3.533 ;
      RECT 74.045 3.32 74.131 3.54 ;
      RECT 74.025 3.325 74.04 3.546 ;
      RECT 74.015 3.365 74.025 3.548 ;
      RECT 73.985 3.375 74.015 3.55 ;
      RECT 73.98 3.38 73.985 3.552 ;
      RECT 73.955 3.385 73.98 3.554 ;
      RECT 73.94 3.39 73.955 3.556 ;
      RECT 73.925 3.392 73.94 3.558 ;
      RECT 73.92 3.397 73.925 3.56 ;
      RECT 73.87 3.405 73.92 3.563 ;
      RECT 73.845 3.414 73.87 3.568 ;
      RECT 73.835 3.421 73.845 3.573 ;
      RECT 73.83 3.424 73.835 3.577 ;
      RECT 73.81 3.427 73.83 3.586 ;
      RECT 73.78 3.435 73.81 3.606 ;
      RECT 73.751 3.448 73.78 3.628 ;
      RECT 73.665 3.482 73.751 3.672 ;
      RECT 73.66 3.508 73.665 3.71 ;
      RECT 73.655 3.512 73.66 3.719 ;
      RECT 73.62 3.525 73.655 3.752 ;
      RECT 73.61 3.539 73.62 3.79 ;
      RECT 73.605 3.543 73.61 3.803 ;
      RECT 73.6 3.547 73.605 3.808 ;
      RECT 73.59 3.555 73.6 3.82 ;
      RECT 73.585 3.562 73.59 3.835 ;
      RECT 73.56 3.575 73.585 3.86 ;
      RECT 73.52 3.604 73.56 3.915 ;
      RECT 73.505 3.629 73.52 3.97 ;
      RECT 73.495 3.64 73.505 3.993 ;
      RECT 73.49 3.647 73.495 4.005 ;
      RECT 73.485 3.651 73.49 4.013 ;
      RECT 73.43 3.679 73.485 4.055 ;
      RECT 73.41 3.715 73.43 4.055 ;
      RECT 73.395 3.73 73.41 4.055 ;
      RECT 73.34 3.762 73.395 4.055 ;
      RECT 73.33 3.792 73.34 4.055 ;
      RECT 72.94 3.407 73.125 3.645 ;
      RECT 72.925 3.409 73.135 3.64 ;
      RECT 72.81 3.355 73.07 3.615 ;
      RECT 72.805 3.392 73.07 3.569 ;
      RECT 72.8 3.402 73.07 3.566 ;
      RECT 72.795 3.442 73.135 3.56 ;
      RECT 72.79 3.475 73.135 3.55 ;
      RECT 72.8 3.417 73.15 3.488 ;
      RECT 73.097 4.515 73.11 5.045 ;
      RECT 73.011 4.515 73.11 5.044 ;
      RECT 73.011 4.515 73.115 5.043 ;
      RECT 72.925 4.515 73.115 5.041 ;
      RECT 72.92 4.515 73.115 5.038 ;
      RECT 72.92 4.515 73.125 5.036 ;
      RECT 72.915 4.807 73.125 5.033 ;
      RECT 72.915 4.817 73.13 5.03 ;
      RECT 72.915 4.885 73.135 5.026 ;
      RECT 72.905 4.89 73.135 5.025 ;
      RECT 72.905 4.982 73.14 5.022 ;
      RECT 72.89 4.515 73.15 4.775 ;
      RECT 72.82 10.055 73.11 10.285 ;
      RECT 72.88 9.315 73.05 10.285 ;
      RECT 72.795 9.34 73.135 9.685 ;
      RECT 72.82 9.315 73.11 9.685 ;
      RECT 72.12 3.505 72.165 5.04 ;
      RECT 72.32 3.505 72.35 3.72 ;
      RECT 70.695 3.245 70.815 3.455 ;
      RECT 70.355 3.195 70.615 3.455 ;
      RECT 70.355 3.24 70.65 3.445 ;
      RECT 72.36 3.521 72.365 3.575 ;
      RECT 72.355 3.514 72.36 3.708 ;
      RECT 72.35 3.508 72.355 3.715 ;
      RECT 72.305 3.505 72.32 3.728 ;
      RECT 72.3 3.505 72.305 3.75 ;
      RECT 72.295 3.505 72.3 3.798 ;
      RECT 72.29 3.505 72.295 3.818 ;
      RECT 72.28 3.505 72.29 3.925 ;
      RECT 72.275 3.505 72.28 3.988 ;
      RECT 72.27 3.505 72.275 4.045 ;
      RECT 72.265 3.505 72.27 4.053 ;
      RECT 72.25 3.505 72.265 4.16 ;
      RECT 72.24 3.505 72.25 4.295 ;
      RECT 72.23 3.505 72.24 4.405 ;
      RECT 72.22 3.505 72.23 4.462 ;
      RECT 72.215 3.505 72.22 4.502 ;
      RECT 72.21 3.505 72.215 4.538 ;
      RECT 72.2 3.505 72.21 4.578 ;
      RECT 72.195 3.505 72.2 4.62 ;
      RECT 72.175 3.505 72.195 4.685 ;
      RECT 72.18 4.83 72.185 5.01 ;
      RECT 72.175 4.812 72.18 5.018 ;
      RECT 72.17 3.505 72.175 4.748 ;
      RECT 72.17 4.792 72.175 5.025 ;
      RECT 72.165 3.505 72.17 5.035 ;
      RECT 72.11 3.505 72.12 3.805 ;
      RECT 72.115 4.052 72.12 5.04 ;
      RECT 72.11 4.117 72.115 5.04 ;
      RECT 72.105 3.506 72.11 3.795 ;
      RECT 72.1 4.182 72.11 5.04 ;
      RECT 72.095 3.507 72.105 3.785 ;
      RECT 72.085 4.295 72.1 5.04 ;
      RECT 72.09 3.508 72.095 3.775 ;
      RECT 72.07 3.509 72.09 3.753 ;
      RECT 72.075 4.392 72.085 5.04 ;
      RECT 72.07 4.467 72.075 5.04 ;
      RECT 72.06 3.508 72.07 3.73 ;
      RECT 72.065 4.51 72.07 5.04 ;
      RECT 72.06 4.537 72.065 5.04 ;
      RECT 72.05 3.506 72.06 3.718 ;
      RECT 72.055 4.58 72.06 5.04 ;
      RECT 72.05 4.607 72.055 5.04 ;
      RECT 72.04 3.505 72.05 3.705 ;
      RECT 72.045 4.622 72.05 5.04 ;
      RECT 72.005 4.68 72.045 5.04 ;
      RECT 72.035 3.504 72.04 3.69 ;
      RECT 72.03 3.502 72.035 3.683 ;
      RECT 72.02 3.499 72.03 3.673 ;
      RECT 72.015 3.496 72.02 3.658 ;
      RECT 72 3.492 72.015 3.651 ;
      RECT 71.995 4.735 72.005 5.04 ;
      RECT 71.995 3.489 72 3.646 ;
      RECT 71.98 3.485 71.995 3.64 ;
      RECT 71.99 4.752 71.995 5.04 ;
      RECT 71.98 4.815 71.99 5.04 ;
      RECT 71.9 3.47 71.98 3.62 ;
      RECT 71.975 4.822 71.98 5.035 ;
      RECT 71.97 4.83 71.975 5.025 ;
      RECT 71.89 3.456 71.9 3.604 ;
      RECT 71.875 3.452 71.89 3.602 ;
      RECT 71.865 3.447 71.875 3.598 ;
      RECT 71.84 3.44 71.865 3.59 ;
      RECT 71.835 3.435 71.84 3.585 ;
      RECT 71.825 3.435 71.835 3.583 ;
      RECT 71.815 3.433 71.825 3.581 ;
      RECT 71.785 3.425 71.815 3.575 ;
      RECT 71.77 3.417 71.785 3.568 ;
      RECT 71.75 3.412 71.77 3.561 ;
      RECT 71.745 3.408 71.75 3.556 ;
      RECT 71.715 3.401 71.745 3.55 ;
      RECT 71.69 3.392 71.715 3.54 ;
      RECT 71.66 3.385 71.69 3.532 ;
      RECT 71.635 3.375 71.66 3.523 ;
      RECT 71.62 3.367 71.635 3.517 ;
      RECT 71.595 3.362 71.62 3.512 ;
      RECT 71.585 3.358 71.595 3.507 ;
      RECT 71.565 3.353 71.585 3.502 ;
      RECT 71.53 3.348 71.565 3.495 ;
      RECT 71.47 3.343 71.53 3.488 ;
      RECT 71.457 3.339 71.47 3.486 ;
      RECT 71.371 3.334 71.457 3.483 ;
      RECT 71.285 3.324 71.371 3.479 ;
      RECT 71.244 3.317 71.285 3.476 ;
      RECT 71.158 3.31 71.244 3.473 ;
      RECT 71.072 3.3 71.158 3.469 ;
      RECT 70.986 3.29 71.072 3.464 ;
      RECT 70.9 3.28 70.986 3.46 ;
      RECT 70.89 3.265 70.9 3.458 ;
      RECT 70.88 3.25 70.89 3.458 ;
      RECT 70.815 3.245 70.88 3.457 ;
      RECT 70.65 3.242 70.695 3.45 ;
      RECT 71.895 4.147 71.9 4.338 ;
      RECT 71.89 4.142 71.895 4.345 ;
      RECT 71.876 4.14 71.89 4.351 ;
      RECT 71.79 4.14 71.876 4.353 ;
      RECT 71.786 4.14 71.79 4.356 ;
      RECT 71.7 4.14 71.786 4.374 ;
      RECT 71.69 4.145 71.7 4.393 ;
      RECT 71.68 4.2 71.69 4.397 ;
      RECT 71.655 4.215 71.68 4.404 ;
      RECT 71.615 4.235 71.655 4.417 ;
      RECT 71.61 4.247 71.615 4.427 ;
      RECT 71.595 4.253 71.61 4.432 ;
      RECT 71.59 4.258 71.595 4.436 ;
      RECT 71.57 4.265 71.59 4.441 ;
      RECT 71.5 4.29 71.57 4.458 ;
      RECT 71.46 4.318 71.5 4.478 ;
      RECT 71.455 4.328 71.46 4.486 ;
      RECT 71.435 4.335 71.455 4.488 ;
      RECT 71.43 4.342 71.435 4.491 ;
      RECT 71.4 4.35 71.43 4.494 ;
      RECT 71.395 4.355 71.4 4.498 ;
      RECT 71.321 4.359 71.395 4.506 ;
      RECT 71.235 4.368 71.321 4.522 ;
      RECT 71.231 4.373 71.235 4.531 ;
      RECT 71.145 4.378 71.231 4.541 ;
      RECT 71.105 4.386 71.145 4.553 ;
      RECT 71.055 4.392 71.105 4.56 ;
      RECT 70.97 4.401 71.055 4.575 ;
      RECT 70.895 4.412 70.97 4.593 ;
      RECT 70.86 4.419 70.895 4.603 ;
      RECT 70.785 4.427 70.86 4.608 ;
      RECT 70.73 4.436 70.785 4.608 ;
      RECT 70.705 4.441 70.73 4.606 ;
      RECT 70.695 4.444 70.705 4.604 ;
      RECT 70.66 4.446 70.695 4.602 ;
      RECT 70.63 4.448 70.66 4.598 ;
      RECT 70.585 4.447 70.63 4.594 ;
      RECT 70.565 4.442 70.585 4.591 ;
      RECT 70.515 4.427 70.565 4.588 ;
      RECT 70.505 4.412 70.515 4.583 ;
      RECT 70.455 4.397 70.505 4.573 ;
      RECT 70.405 4.372 70.455 4.553 ;
      RECT 70.395 4.357 70.405 4.535 ;
      RECT 70.39 4.355 70.395 4.529 ;
      RECT 70.37 4.35 70.39 4.524 ;
      RECT 70.365 4.342 70.37 4.518 ;
      RECT 70.35 4.336 70.365 4.511 ;
      RECT 70.345 4.331 70.35 4.503 ;
      RECT 70.325 4.326 70.345 4.495 ;
      RECT 70.31 4.319 70.325 4.488 ;
      RECT 70.295 4.313 70.31 4.479 ;
      RECT 70.29 4.307 70.295 4.472 ;
      RECT 70.245 4.282 70.29 4.458 ;
      RECT 70.23 4.252 70.245 4.44 ;
      RECT 70.215 4.235 70.23 4.431 ;
      RECT 70.19 4.215 70.215 4.419 ;
      RECT 70.15 4.185 70.19 4.399 ;
      RECT 70.14 4.155 70.15 4.384 ;
      RECT 70.125 4.145 70.14 4.377 ;
      RECT 70.07 4.11 70.125 4.356 ;
      RECT 70.055 4.073 70.07 4.335 ;
      RECT 70.045 4.06 70.055 4.327 ;
      RECT 69.995 4.03 70.045 4.309 ;
      RECT 69.98 3.96 69.995 4.29 ;
      RECT 69.935 3.96 69.98 4.273 ;
      RECT 69.91 3.96 69.935 4.255 ;
      RECT 69.9 3.96 69.91 4.248 ;
      RECT 69.821 3.96 69.9 4.241 ;
      RECT 69.735 3.96 69.821 4.233 ;
      RECT 69.72 3.992 69.735 4.228 ;
      RECT 69.645 4.002 69.72 4.224 ;
      RECT 69.625 4.012 69.645 4.219 ;
      RECT 69.6 4.012 69.625 4.216 ;
      RECT 69.59 4.002 69.6 4.215 ;
      RECT 69.58 3.975 69.59 4.214 ;
      RECT 69.54 3.97 69.58 4.212 ;
      RECT 69.495 3.97 69.54 4.208 ;
      RECT 69.47 3.97 69.495 4.203 ;
      RECT 69.42 3.97 69.47 4.19 ;
      RECT 69.38 3.975 69.39 4.175 ;
      RECT 69.39 3.97 69.42 4.18 ;
      RECT 71.375 3.75 71.635 4.01 ;
      RECT 71.37 3.772 71.635 3.968 ;
      RECT 70.61 3.6 70.83 3.965 ;
      RECT 70.592 3.687 70.83 3.964 ;
      RECT 70.575 3.692 70.83 3.961 ;
      RECT 70.575 3.692 70.85 3.96 ;
      RECT 70.545 3.702 70.85 3.958 ;
      RECT 70.54 3.717 70.85 3.954 ;
      RECT 70.54 3.717 70.855 3.953 ;
      RECT 70.535 3.775 70.855 3.951 ;
      RECT 70.535 3.775 70.865 3.948 ;
      RECT 70.53 3.84 70.865 3.943 ;
      RECT 70.61 3.6 70.87 3.86 ;
      RECT 69.355 3.43 69.615 3.69 ;
      RECT 69.355 3.473 69.701 3.664 ;
      RECT 69.355 3.473 69.745 3.663 ;
      RECT 69.355 3.473 69.765 3.661 ;
      RECT 69.355 3.473 69.865 3.66 ;
      RECT 69.355 3.473 69.885 3.658 ;
      RECT 69.355 3.473 69.895 3.653 ;
      RECT 69.765 3.44 69.955 3.65 ;
      RECT 69.765 3.442 69.96 3.648 ;
      RECT 69.755 3.447 69.965 3.64 ;
      RECT 69.701 3.471 69.965 3.64 ;
      RECT 69.745 3.465 69.755 3.662 ;
      RECT 69.755 3.445 69.96 3.648 ;
      RECT 68.71 4.505 68.915 4.735 ;
      RECT 68.65 4.455 68.705 4.715 ;
      RECT 68.71 4.455 68.91 4.735 ;
      RECT 69.68 4.77 69.685 4.797 ;
      RECT 69.67 4.68 69.68 4.802 ;
      RECT 69.665 4.602 69.67 4.808 ;
      RECT 69.655 4.592 69.665 4.815 ;
      RECT 69.65 4.582 69.655 4.821 ;
      RECT 69.64 4.577 69.65 4.823 ;
      RECT 69.625 4.569 69.64 4.831 ;
      RECT 69.61 4.56 69.625 4.843 ;
      RECT 69.6 4.552 69.61 4.853 ;
      RECT 69.565 4.47 69.6 4.871 ;
      RECT 69.53 4.47 69.565 4.89 ;
      RECT 69.515 4.47 69.53 4.898 ;
      RECT 69.46 4.47 69.515 4.898 ;
      RECT 69.426 4.47 69.46 4.889 ;
      RECT 69.34 4.47 69.426 4.865 ;
      RECT 69.33 4.53 69.34 4.847 ;
      RECT 69.29 4.532 69.33 4.838 ;
      RECT 69.285 4.534 69.29 4.828 ;
      RECT 69.265 4.536 69.285 4.823 ;
      RECT 69.255 4.539 69.265 4.818 ;
      RECT 69.245 4.54 69.255 4.813 ;
      RECT 69.221 4.541 69.245 4.805 ;
      RECT 69.135 4.546 69.221 4.783 ;
      RECT 69.08 4.545 69.135 4.756 ;
      RECT 69.065 4.538 69.08 4.743 ;
      RECT 69.03 4.533 69.065 4.739 ;
      RECT 68.975 4.525 69.03 4.738 ;
      RECT 68.915 4.512 68.975 4.736 ;
      RECT 68.705 4.455 68.71 4.723 ;
      RECT 68.78 3.825 68.965 4.035 ;
      RECT 68.77 3.83 68.98 4.028 ;
      RECT 68.81 3.735 69.07 3.995 ;
      RECT 68.765 3.892 69.07 3.918 ;
      RECT 68.11 3.685 68.115 4.485 ;
      RECT 68.055 3.735 68.085 4.485 ;
      RECT 68.045 3.735 68.05 4.045 ;
      RECT 68.03 3.735 68.035 4.04 ;
      RECT 67.575 3.78 67.59 3.995 ;
      RECT 67.505 3.78 67.59 3.99 ;
      RECT 68.77 3.36 68.84 3.57 ;
      RECT 68.84 3.367 68.85 3.565 ;
      RECT 68.736 3.36 68.77 3.577 ;
      RECT 68.65 3.36 68.736 3.601 ;
      RECT 68.64 3.365 68.65 3.62 ;
      RECT 68.635 3.377 68.64 3.623 ;
      RECT 68.62 3.392 68.635 3.627 ;
      RECT 68.615 3.41 68.62 3.631 ;
      RECT 68.575 3.42 68.615 3.64 ;
      RECT 68.56 3.427 68.575 3.652 ;
      RECT 68.545 3.432 68.56 3.657 ;
      RECT 68.53 3.435 68.545 3.662 ;
      RECT 68.52 3.437 68.53 3.666 ;
      RECT 68.485 3.444 68.52 3.674 ;
      RECT 68.45 3.452 68.485 3.688 ;
      RECT 68.44 3.458 68.45 3.697 ;
      RECT 68.435 3.46 68.44 3.699 ;
      RECT 68.415 3.463 68.435 3.705 ;
      RECT 68.385 3.47 68.415 3.716 ;
      RECT 68.375 3.476 68.385 3.723 ;
      RECT 68.35 3.479 68.375 3.73 ;
      RECT 68.34 3.483 68.35 3.738 ;
      RECT 68.335 3.484 68.34 3.76 ;
      RECT 68.33 3.485 68.335 3.775 ;
      RECT 68.325 3.486 68.33 3.79 ;
      RECT 68.32 3.487 68.325 3.805 ;
      RECT 68.315 3.488 68.32 3.835 ;
      RECT 68.305 3.49 68.315 3.868 ;
      RECT 68.29 3.494 68.305 3.915 ;
      RECT 68.28 3.497 68.29 3.96 ;
      RECT 68.275 3.5 68.28 3.988 ;
      RECT 68.265 3.502 68.275 4.015 ;
      RECT 68.26 3.505 68.265 4.05 ;
      RECT 68.23 3.51 68.26 4.108 ;
      RECT 68.225 3.515 68.23 4.193 ;
      RECT 68.22 3.517 68.225 4.228 ;
      RECT 68.215 3.519 68.22 4.31 ;
      RECT 68.21 3.521 68.215 4.398 ;
      RECT 68.2 3.523 68.21 4.48 ;
      RECT 68.185 3.537 68.2 4.485 ;
      RECT 68.15 3.582 68.185 4.485 ;
      RECT 68.14 3.622 68.15 4.485 ;
      RECT 68.125 3.65 68.14 4.485 ;
      RECT 68.12 3.667 68.125 4.485 ;
      RECT 68.115 3.675 68.12 4.485 ;
      RECT 68.105 3.69 68.11 4.485 ;
      RECT 68.1 3.697 68.105 4.485 ;
      RECT 68.09 3.717 68.1 4.485 ;
      RECT 68.085 3.73 68.09 4.485 ;
      RECT 68.05 3.735 68.055 4.07 ;
      RECT 68.035 4.125 68.055 4.485 ;
      RECT 68.035 3.735 68.045 4.043 ;
      RECT 68.03 4.165 68.035 4.485 ;
      RECT 67.98 3.735 68.03 4.038 ;
      RECT 68.025 4.202 68.03 4.485 ;
      RECT 68.015 4.225 68.025 4.485 ;
      RECT 68.01 4.27 68.015 4.485 ;
      RECT 68 4.28 68.01 4.478 ;
      RECT 67.926 3.735 67.98 4.032 ;
      RECT 67.84 3.735 67.926 4.025 ;
      RECT 67.791 3.782 67.84 4.018 ;
      RECT 67.705 3.79 67.791 4.011 ;
      RECT 67.69 3.787 67.705 4.006 ;
      RECT 67.676 3.78 67.69 4.005 ;
      RECT 67.59 3.78 67.676 4 ;
      RECT 67.495 3.785 67.505 3.985 ;
      RECT 67.085 3.215 67.1 3.615 ;
      RECT 67.28 3.215 67.285 3.475 ;
      RECT 67.025 3.215 67.07 3.475 ;
      RECT 67.48 4.52 67.485 4.725 ;
      RECT 67.475 4.51 67.48 4.73 ;
      RECT 67.47 4.497 67.475 4.735 ;
      RECT 67.465 4.477 67.47 4.735 ;
      RECT 67.44 4.43 67.465 4.735 ;
      RECT 67.405 4.345 67.44 4.735 ;
      RECT 67.4 4.282 67.405 4.735 ;
      RECT 67.395 4.267 67.4 4.735 ;
      RECT 67.38 4.227 67.395 4.735 ;
      RECT 67.375 4.202 67.38 4.735 ;
      RECT 67.365 4.185 67.375 4.735 ;
      RECT 67.33 4.107 67.365 4.735 ;
      RECT 67.325 4.05 67.33 4.735 ;
      RECT 67.32 4.037 67.325 4.735 ;
      RECT 67.31 4.015 67.32 4.735 ;
      RECT 67.3 3.98 67.31 4.735 ;
      RECT 67.29 3.95 67.3 4.735 ;
      RECT 67.28 3.865 67.29 4.378 ;
      RECT 67.287 4.51 67.29 4.735 ;
      RECT 67.285 4.52 67.287 4.735 ;
      RECT 67.275 4.53 67.285 4.73 ;
      RECT 67.27 3.215 67.28 3.61 ;
      RECT 67.275 3.742 67.28 4.353 ;
      RECT 67.27 3.64 67.275 4.336 ;
      RECT 67.26 3.215 67.27 4.312 ;
      RECT 67.255 3.215 67.26 4.283 ;
      RECT 67.25 3.215 67.255 4.273 ;
      RECT 67.23 3.215 67.25 4.235 ;
      RECT 67.225 3.215 67.23 4.193 ;
      RECT 67.22 3.215 67.225 4.173 ;
      RECT 67.19 3.215 67.22 4.123 ;
      RECT 67.18 3.215 67.19 4.07 ;
      RECT 67.175 3.215 67.18 4.043 ;
      RECT 67.17 3.215 67.175 4.028 ;
      RECT 67.16 3.215 67.17 4.005 ;
      RECT 67.15 3.215 67.16 3.98 ;
      RECT 67.145 3.215 67.15 3.92 ;
      RECT 67.135 3.215 67.145 3.858 ;
      RECT 67.13 3.215 67.135 3.778 ;
      RECT 67.125 3.215 67.13 3.743 ;
      RECT 67.12 3.215 67.125 3.718 ;
      RECT 67.115 3.215 67.12 3.703 ;
      RECT 67.11 3.215 67.115 3.673 ;
      RECT 67.105 3.215 67.11 3.65 ;
      RECT 67.1 3.215 67.105 3.623 ;
      RECT 67.07 3.215 67.085 3.61 ;
      RECT 66.225 4.75 66.41 4.96 ;
      RECT 66.215 4.755 66.425 4.953 ;
      RECT 66.215 4.755 66.445 4.925 ;
      RECT 66.215 4.755 66.46 4.904 ;
      RECT 66.215 4.755 66.475 4.902 ;
      RECT 66.215 4.755 66.485 4.901 ;
      RECT 66.215 4.755 66.515 4.898 ;
      RECT 66.865 4.6 67.125 4.86 ;
      RECT 66.825 4.647 67.125 4.843 ;
      RECT 66.816 4.655 66.825 4.846 ;
      RECT 66.41 4.748 67.125 4.843 ;
      RECT 66.73 4.673 66.816 4.853 ;
      RECT 66.425 4.745 67.125 4.843 ;
      RECT 66.671 4.695 66.73 4.865 ;
      RECT 66.445 4.741 67.125 4.843 ;
      RECT 66.585 4.707 66.671 4.876 ;
      RECT 66.46 4.737 67.125 4.843 ;
      RECT 66.53 4.72 66.585 4.888 ;
      RECT 66.475 4.735 67.125 4.843 ;
      RECT 66.515 4.726 66.53 4.894 ;
      RECT 66.485 4.731 67.125 4.843 ;
      RECT 66.63 4.255 66.89 4.515 ;
      RECT 66.63 4.275 67 4.485 ;
      RECT 66.63 4.28 67.01 4.48 ;
      RECT 66.821 3.694 66.9 3.925 ;
      RECT 66.735 3.697 66.95 3.92 ;
      RECT 66.73 3.697 66.95 3.915 ;
      RECT 66.73 3.702 66.96 3.913 ;
      RECT 66.705 3.702 66.96 3.91 ;
      RECT 66.705 3.71 66.97 3.908 ;
      RECT 66.585 3.645 66.845 3.905 ;
      RECT 66.585 3.692 66.895 3.905 ;
      RECT 65.84 4.265 65.845 4.525 ;
      RECT 65.67 4.035 65.675 4.525 ;
      RECT 65.555 4.275 65.56 4.5 ;
      RECT 66.265 3.37 66.27 3.58 ;
      RECT 66.27 3.375 66.285 3.575 ;
      RECT 66.205 3.37 66.265 3.588 ;
      RECT 66.19 3.37 66.205 3.598 ;
      RECT 66.14 3.37 66.19 3.615 ;
      RECT 66.12 3.37 66.14 3.638 ;
      RECT 66.105 3.37 66.12 3.65 ;
      RECT 66.085 3.37 66.105 3.66 ;
      RECT 66.075 3.375 66.085 3.669 ;
      RECT 66.07 3.385 66.075 3.674 ;
      RECT 66.065 3.397 66.07 3.678 ;
      RECT 66.055 3.42 66.065 3.683 ;
      RECT 66.05 3.435 66.055 3.687 ;
      RECT 66.045 3.452 66.05 3.69 ;
      RECT 66.04 3.46 66.045 3.693 ;
      RECT 66.03 3.465 66.04 3.697 ;
      RECT 66.025 3.472 66.03 3.702 ;
      RECT 66.015 3.477 66.025 3.706 ;
      RECT 65.99 3.489 66.015 3.717 ;
      RECT 65.97 3.506 65.99 3.733 ;
      RECT 65.945 3.523 65.97 3.755 ;
      RECT 65.91 3.546 65.945 3.813 ;
      RECT 65.89 3.568 65.91 3.875 ;
      RECT 65.885 3.578 65.89 3.91 ;
      RECT 65.875 3.585 65.885 3.948 ;
      RECT 65.87 3.592 65.875 3.968 ;
      RECT 65.865 3.603 65.87 4.005 ;
      RECT 65.86 3.611 65.865 4.07 ;
      RECT 65.85 3.622 65.86 4.123 ;
      RECT 65.845 3.64 65.85 4.193 ;
      RECT 65.84 3.65 65.845 4.23 ;
      RECT 65.835 3.66 65.84 4.525 ;
      RECT 65.83 3.672 65.835 4.525 ;
      RECT 65.825 3.682 65.83 4.525 ;
      RECT 65.815 3.692 65.825 4.525 ;
      RECT 65.805 3.715 65.815 4.525 ;
      RECT 65.79 3.75 65.805 4.525 ;
      RECT 65.75 3.812 65.79 4.525 ;
      RECT 65.745 3.865 65.75 4.525 ;
      RECT 65.72 3.9 65.745 4.525 ;
      RECT 65.705 3.945 65.72 4.525 ;
      RECT 65.7 3.967 65.705 4.525 ;
      RECT 65.69 3.98 65.7 4.525 ;
      RECT 65.68 4.005 65.69 4.525 ;
      RECT 65.675 4.027 65.68 4.525 ;
      RECT 65.65 4.065 65.67 4.525 ;
      RECT 65.61 4.122 65.65 4.525 ;
      RECT 65.605 4.172 65.61 4.525 ;
      RECT 65.6 4.19 65.605 4.525 ;
      RECT 65.595 4.202 65.6 4.525 ;
      RECT 65.585 4.22 65.595 4.525 ;
      RECT 65.575 4.24 65.585 4.5 ;
      RECT 65.57 4.257 65.575 4.5 ;
      RECT 65.56 4.27 65.57 4.5 ;
      RECT 65.53 4.28 65.555 4.5 ;
      RECT 65.52 4.287 65.53 4.5 ;
      RECT 65.505 4.297 65.52 4.495 ;
      RECT 64.595 10.055 64.89 10.285 ;
      RECT 64.655 8.575 64.825 10.285 ;
      RECT 64.605 8.945 64.955 9.295 ;
      RECT 64.595 8.575 64.885 8.805 ;
      RECT 63.605 10.055 63.9 10.285 ;
      RECT 63.665 8.575 63.835 10.285 ;
      RECT 63.605 8.575 63.895 8.805 ;
      RECT 63.605 8.61 64.455 8.77 ;
      RECT 64.29 8.205 64.455 8.77 ;
      RECT 63.605 8.605 64 8.77 ;
      RECT 64.225 8.205 64.515 8.435 ;
      RECT 64.225 8.235 64.685 8.405 ;
      RECT 64.19 4.025 64.51 4.26 ;
      RECT 64.19 4.055 64.68 4.225 ;
      RECT 64.19 3.69 64.38 4.26 ;
      RECT 63.605 3.655 63.895 3.885 ;
      RECT 63.605 3.69 64.38 3.86 ;
      RECT 63.665 2.175 63.835 3.885 ;
      RECT 63.605 2.175 63.9 2.405 ;
      RECT 63.235 4.025 63.525 4.255 ;
      RECT 63.235 4.055 63.695 4.225 ;
      RECT 63.3 2.95 63.465 4.255 ;
      RECT 61.815 2.915 62.105 3.145 ;
      RECT 61.815 2.95 63.465 3.12 ;
      RECT 61.875 2.175 62.045 3.145 ;
      RECT 61.815 2.175 62.105 2.405 ;
      RECT 61.815 10.055 62.105 10.285 ;
      RECT 61.875 9.315 62.045 10.285 ;
      RECT 61.875 9.405 63.465 9.575 ;
      RECT 63.295 8.205 63.465 9.575 ;
      RECT 61.815 9.315 62.105 9.545 ;
      RECT 63.235 8.205 63.525 8.435 ;
      RECT 63.235 8.235 63.695 8.405 ;
      RECT 62.245 3.26 62.595 3.61 ;
      RECT 59.91 3.32 62.595 3.49 ;
      RECT 62.075 3.315 62.595 3.49 ;
      RECT 59.91 2.635 60.08 3.49 ;
      RECT 59.81 2.635 60.16 2.985 ;
      RECT 62.27 8.94 62.595 9.265 ;
      RECT 57.7 8.9 58.05 9.25 ;
      RECT 62.245 8.945 62.595 9.175 ;
      RECT 57.465 8.945 58.05 9.175 ;
      RECT 62.075 8.97 62.595 9.145 ;
      RECT 57.295 8.975 58.05 9.145 ;
      RECT 57.465 8.97 62.595 9.14 ;
      RECT 61.47 3.66 61.79 3.98 ;
      RECT 61.445 3.655 61.735 3.885 ;
      RECT 61.37 3.685 61.79 3.86 ;
      RECT 61.27 3.685 61.79 3.855 ;
      RECT 61.47 8.54 61.79 8.83 ;
      RECT 61.445 8.575 61.79 8.805 ;
      RECT 61.27 8.605 61.79 8.775 ;
      RECT 58.105 3.76 58.29 3.97 ;
      RECT 58.095 3.765 58.305 3.963 ;
      RECT 58.095 3.765 58.391 3.94 ;
      RECT 58.095 3.765 58.45 3.915 ;
      RECT 58.095 3.765 58.505 3.895 ;
      RECT 58.095 3.765 58.515 3.883 ;
      RECT 58.095 3.765 58.71 3.822 ;
      RECT 58.095 3.765 58.74 3.805 ;
      RECT 58.095 3.765 58.76 3.795 ;
      RECT 58.64 3.53 58.9 3.79 ;
      RECT 58.625 3.62 58.64 3.837 ;
      RECT 58.16 3.752 58.9 3.79 ;
      RECT 58.611 3.631 58.625 3.843 ;
      RECT 58.2 3.745 58.9 3.79 ;
      RECT 58.525 3.671 58.611 3.862 ;
      RECT 58.45 3.732 58.9 3.79 ;
      RECT 58.52 3.707 58.525 3.879 ;
      RECT 58.505 3.717 58.9 3.79 ;
      RECT 58.515 3.712 58.52 3.881 ;
      RECT 57.44 3.795 57.545 4.055 ;
      RECT 58.255 3.32 58.26 3.545 ;
      RECT 58.385 3.32 58.44 3.53 ;
      RECT 58.44 3.325 58.45 3.523 ;
      RECT 58.346 3.32 58.385 3.533 ;
      RECT 58.26 3.32 58.346 3.54 ;
      RECT 58.24 3.325 58.255 3.546 ;
      RECT 58.23 3.365 58.24 3.548 ;
      RECT 58.2 3.375 58.23 3.55 ;
      RECT 58.195 3.38 58.2 3.552 ;
      RECT 58.17 3.385 58.195 3.554 ;
      RECT 58.155 3.39 58.17 3.556 ;
      RECT 58.14 3.392 58.155 3.558 ;
      RECT 58.135 3.397 58.14 3.56 ;
      RECT 58.085 3.405 58.135 3.563 ;
      RECT 58.06 3.414 58.085 3.568 ;
      RECT 58.05 3.421 58.06 3.573 ;
      RECT 58.045 3.424 58.05 3.577 ;
      RECT 58.025 3.427 58.045 3.586 ;
      RECT 57.995 3.435 58.025 3.606 ;
      RECT 57.966 3.448 57.995 3.628 ;
      RECT 57.88 3.482 57.966 3.672 ;
      RECT 57.875 3.508 57.88 3.71 ;
      RECT 57.87 3.512 57.875 3.719 ;
      RECT 57.835 3.525 57.87 3.752 ;
      RECT 57.825 3.539 57.835 3.79 ;
      RECT 57.82 3.543 57.825 3.803 ;
      RECT 57.815 3.547 57.82 3.808 ;
      RECT 57.805 3.555 57.815 3.82 ;
      RECT 57.8 3.562 57.805 3.835 ;
      RECT 57.775 3.575 57.8 3.86 ;
      RECT 57.735 3.604 57.775 3.915 ;
      RECT 57.72 3.629 57.735 3.97 ;
      RECT 57.71 3.64 57.72 3.993 ;
      RECT 57.705 3.647 57.71 4.005 ;
      RECT 57.7 3.651 57.705 4.013 ;
      RECT 57.645 3.679 57.7 4.055 ;
      RECT 57.625 3.715 57.645 4.055 ;
      RECT 57.61 3.73 57.625 4.055 ;
      RECT 57.555 3.762 57.61 4.055 ;
      RECT 57.545 3.792 57.555 4.055 ;
      RECT 57.155 3.407 57.34 3.645 ;
      RECT 57.14 3.409 57.35 3.64 ;
      RECT 57.025 3.355 57.285 3.615 ;
      RECT 57.02 3.392 57.285 3.569 ;
      RECT 57.015 3.402 57.285 3.566 ;
      RECT 57.01 3.442 57.35 3.56 ;
      RECT 57.005 3.475 57.35 3.55 ;
      RECT 57.015 3.417 57.365 3.488 ;
      RECT 57.312 4.515 57.325 5.045 ;
      RECT 57.226 4.515 57.325 5.044 ;
      RECT 57.226 4.515 57.33 5.043 ;
      RECT 57.14 4.515 57.33 5.041 ;
      RECT 57.135 4.515 57.33 5.038 ;
      RECT 57.135 4.515 57.34 5.036 ;
      RECT 57.13 4.807 57.34 5.033 ;
      RECT 57.13 4.817 57.345 5.03 ;
      RECT 57.13 4.885 57.35 5.026 ;
      RECT 57.12 4.89 57.35 5.025 ;
      RECT 57.12 4.982 57.355 5.022 ;
      RECT 57.105 4.515 57.365 4.775 ;
      RECT 57.035 10.055 57.325 10.285 ;
      RECT 57.095 9.315 57.265 10.285 ;
      RECT 57.01 9.34 57.35 9.685 ;
      RECT 57.035 9.315 57.325 9.685 ;
      RECT 56.335 3.505 56.38 5.04 ;
      RECT 56.535 3.505 56.565 3.72 ;
      RECT 54.91 3.245 55.03 3.455 ;
      RECT 54.57 3.195 54.83 3.455 ;
      RECT 54.57 3.24 54.865 3.445 ;
      RECT 56.575 3.521 56.58 3.575 ;
      RECT 56.57 3.514 56.575 3.708 ;
      RECT 56.565 3.508 56.57 3.715 ;
      RECT 56.52 3.505 56.535 3.728 ;
      RECT 56.515 3.505 56.52 3.75 ;
      RECT 56.51 3.505 56.515 3.798 ;
      RECT 56.505 3.505 56.51 3.818 ;
      RECT 56.495 3.505 56.505 3.925 ;
      RECT 56.49 3.505 56.495 3.988 ;
      RECT 56.485 3.505 56.49 4.045 ;
      RECT 56.48 3.505 56.485 4.053 ;
      RECT 56.465 3.505 56.48 4.16 ;
      RECT 56.455 3.505 56.465 4.295 ;
      RECT 56.445 3.505 56.455 4.405 ;
      RECT 56.435 3.505 56.445 4.462 ;
      RECT 56.43 3.505 56.435 4.502 ;
      RECT 56.425 3.505 56.43 4.538 ;
      RECT 56.415 3.505 56.425 4.578 ;
      RECT 56.41 3.505 56.415 4.62 ;
      RECT 56.39 3.505 56.41 4.685 ;
      RECT 56.395 4.83 56.4 5.01 ;
      RECT 56.39 4.812 56.395 5.018 ;
      RECT 56.385 3.505 56.39 4.748 ;
      RECT 56.385 4.792 56.39 5.025 ;
      RECT 56.38 3.505 56.385 5.035 ;
      RECT 56.325 3.505 56.335 3.805 ;
      RECT 56.33 4.052 56.335 5.04 ;
      RECT 56.325 4.117 56.33 5.04 ;
      RECT 56.32 3.506 56.325 3.795 ;
      RECT 56.315 4.182 56.325 5.04 ;
      RECT 56.31 3.507 56.32 3.785 ;
      RECT 56.3 4.295 56.315 5.04 ;
      RECT 56.305 3.508 56.31 3.775 ;
      RECT 56.285 3.509 56.305 3.753 ;
      RECT 56.29 4.392 56.3 5.04 ;
      RECT 56.285 4.467 56.29 5.04 ;
      RECT 56.275 3.508 56.285 3.73 ;
      RECT 56.28 4.51 56.285 5.04 ;
      RECT 56.275 4.537 56.28 5.04 ;
      RECT 56.265 3.506 56.275 3.718 ;
      RECT 56.27 4.58 56.275 5.04 ;
      RECT 56.265 4.607 56.27 5.04 ;
      RECT 56.255 3.505 56.265 3.705 ;
      RECT 56.26 4.622 56.265 5.04 ;
      RECT 56.22 4.68 56.26 5.04 ;
      RECT 56.25 3.504 56.255 3.69 ;
      RECT 56.245 3.502 56.25 3.683 ;
      RECT 56.235 3.499 56.245 3.673 ;
      RECT 56.23 3.496 56.235 3.658 ;
      RECT 56.215 3.492 56.23 3.651 ;
      RECT 56.21 4.735 56.22 5.04 ;
      RECT 56.21 3.489 56.215 3.646 ;
      RECT 56.195 3.485 56.21 3.64 ;
      RECT 56.205 4.752 56.21 5.04 ;
      RECT 56.195 4.815 56.205 5.04 ;
      RECT 56.115 3.47 56.195 3.62 ;
      RECT 56.19 4.822 56.195 5.035 ;
      RECT 56.185 4.83 56.19 5.025 ;
      RECT 56.105 3.456 56.115 3.604 ;
      RECT 56.09 3.452 56.105 3.602 ;
      RECT 56.08 3.447 56.09 3.598 ;
      RECT 56.055 3.44 56.08 3.59 ;
      RECT 56.05 3.435 56.055 3.585 ;
      RECT 56.04 3.435 56.05 3.583 ;
      RECT 56.03 3.433 56.04 3.581 ;
      RECT 56 3.425 56.03 3.575 ;
      RECT 55.985 3.417 56 3.568 ;
      RECT 55.965 3.412 55.985 3.561 ;
      RECT 55.96 3.408 55.965 3.556 ;
      RECT 55.93 3.401 55.96 3.55 ;
      RECT 55.905 3.392 55.93 3.54 ;
      RECT 55.875 3.385 55.905 3.532 ;
      RECT 55.85 3.375 55.875 3.523 ;
      RECT 55.835 3.367 55.85 3.517 ;
      RECT 55.81 3.362 55.835 3.512 ;
      RECT 55.8 3.358 55.81 3.507 ;
      RECT 55.78 3.353 55.8 3.502 ;
      RECT 55.745 3.348 55.78 3.495 ;
      RECT 55.685 3.343 55.745 3.488 ;
      RECT 55.672 3.339 55.685 3.486 ;
      RECT 55.586 3.334 55.672 3.483 ;
      RECT 55.5 3.324 55.586 3.479 ;
      RECT 55.459 3.317 55.5 3.476 ;
      RECT 55.373 3.31 55.459 3.473 ;
      RECT 55.287 3.3 55.373 3.469 ;
      RECT 55.201 3.29 55.287 3.464 ;
      RECT 55.115 3.28 55.201 3.46 ;
      RECT 55.105 3.265 55.115 3.458 ;
      RECT 55.095 3.25 55.105 3.458 ;
      RECT 55.03 3.245 55.095 3.457 ;
      RECT 54.865 3.242 54.91 3.45 ;
      RECT 56.11 4.147 56.115 4.338 ;
      RECT 56.105 4.142 56.11 4.345 ;
      RECT 56.091 4.14 56.105 4.351 ;
      RECT 56.005 4.14 56.091 4.353 ;
      RECT 56.001 4.14 56.005 4.356 ;
      RECT 55.915 4.14 56.001 4.374 ;
      RECT 55.905 4.145 55.915 4.393 ;
      RECT 55.895 4.2 55.905 4.397 ;
      RECT 55.87 4.215 55.895 4.404 ;
      RECT 55.83 4.235 55.87 4.417 ;
      RECT 55.825 4.247 55.83 4.427 ;
      RECT 55.81 4.253 55.825 4.432 ;
      RECT 55.805 4.258 55.81 4.436 ;
      RECT 55.785 4.265 55.805 4.441 ;
      RECT 55.715 4.29 55.785 4.458 ;
      RECT 55.675 4.318 55.715 4.478 ;
      RECT 55.67 4.328 55.675 4.486 ;
      RECT 55.65 4.335 55.67 4.488 ;
      RECT 55.645 4.342 55.65 4.491 ;
      RECT 55.615 4.35 55.645 4.494 ;
      RECT 55.61 4.355 55.615 4.498 ;
      RECT 55.536 4.359 55.61 4.506 ;
      RECT 55.45 4.368 55.536 4.522 ;
      RECT 55.446 4.373 55.45 4.531 ;
      RECT 55.36 4.378 55.446 4.541 ;
      RECT 55.32 4.386 55.36 4.553 ;
      RECT 55.27 4.392 55.32 4.56 ;
      RECT 55.185 4.401 55.27 4.575 ;
      RECT 55.11 4.412 55.185 4.593 ;
      RECT 55.075 4.419 55.11 4.603 ;
      RECT 55 4.427 55.075 4.608 ;
      RECT 54.945 4.436 55 4.608 ;
      RECT 54.92 4.441 54.945 4.606 ;
      RECT 54.91 4.444 54.92 4.604 ;
      RECT 54.875 4.446 54.91 4.602 ;
      RECT 54.845 4.448 54.875 4.598 ;
      RECT 54.8 4.447 54.845 4.594 ;
      RECT 54.78 4.442 54.8 4.591 ;
      RECT 54.73 4.427 54.78 4.588 ;
      RECT 54.72 4.412 54.73 4.583 ;
      RECT 54.67 4.397 54.72 4.573 ;
      RECT 54.62 4.372 54.67 4.553 ;
      RECT 54.61 4.357 54.62 4.535 ;
      RECT 54.605 4.355 54.61 4.529 ;
      RECT 54.585 4.35 54.605 4.524 ;
      RECT 54.58 4.342 54.585 4.518 ;
      RECT 54.565 4.336 54.58 4.511 ;
      RECT 54.56 4.331 54.565 4.503 ;
      RECT 54.54 4.326 54.56 4.495 ;
      RECT 54.525 4.319 54.54 4.488 ;
      RECT 54.51 4.313 54.525 4.479 ;
      RECT 54.505 4.307 54.51 4.472 ;
      RECT 54.46 4.282 54.505 4.458 ;
      RECT 54.445 4.252 54.46 4.44 ;
      RECT 54.43 4.235 54.445 4.431 ;
      RECT 54.405 4.215 54.43 4.419 ;
      RECT 54.365 4.185 54.405 4.399 ;
      RECT 54.355 4.155 54.365 4.384 ;
      RECT 54.34 4.145 54.355 4.377 ;
      RECT 54.285 4.11 54.34 4.356 ;
      RECT 54.27 4.073 54.285 4.335 ;
      RECT 54.26 4.06 54.27 4.327 ;
      RECT 54.21 4.03 54.26 4.309 ;
      RECT 54.195 3.96 54.21 4.29 ;
      RECT 54.15 3.96 54.195 4.273 ;
      RECT 54.125 3.96 54.15 4.255 ;
      RECT 54.115 3.96 54.125 4.248 ;
      RECT 54.036 3.96 54.115 4.241 ;
      RECT 53.95 3.96 54.036 4.233 ;
      RECT 53.935 3.992 53.95 4.228 ;
      RECT 53.86 4.002 53.935 4.224 ;
      RECT 53.84 4.012 53.86 4.219 ;
      RECT 53.815 4.012 53.84 4.216 ;
      RECT 53.805 4.002 53.815 4.215 ;
      RECT 53.795 3.975 53.805 4.214 ;
      RECT 53.755 3.97 53.795 4.212 ;
      RECT 53.71 3.97 53.755 4.208 ;
      RECT 53.685 3.97 53.71 4.203 ;
      RECT 53.635 3.97 53.685 4.19 ;
      RECT 53.595 3.975 53.605 4.175 ;
      RECT 53.605 3.97 53.635 4.18 ;
      RECT 55.59 3.75 55.85 4.01 ;
      RECT 55.585 3.772 55.85 3.968 ;
      RECT 54.825 3.6 55.045 3.965 ;
      RECT 54.807 3.687 55.045 3.964 ;
      RECT 54.79 3.692 55.045 3.961 ;
      RECT 54.79 3.692 55.065 3.96 ;
      RECT 54.76 3.702 55.065 3.958 ;
      RECT 54.755 3.717 55.065 3.954 ;
      RECT 54.755 3.717 55.07 3.953 ;
      RECT 54.75 3.775 55.07 3.951 ;
      RECT 54.75 3.775 55.08 3.948 ;
      RECT 54.745 3.84 55.08 3.943 ;
      RECT 54.825 3.6 55.085 3.86 ;
      RECT 53.57 3.43 53.83 3.69 ;
      RECT 53.57 3.473 53.916 3.664 ;
      RECT 53.57 3.473 53.96 3.663 ;
      RECT 53.57 3.473 53.98 3.661 ;
      RECT 53.57 3.473 54.08 3.66 ;
      RECT 53.57 3.473 54.1 3.658 ;
      RECT 53.57 3.473 54.11 3.653 ;
      RECT 53.98 3.44 54.17 3.65 ;
      RECT 53.98 3.442 54.175 3.648 ;
      RECT 53.97 3.447 54.18 3.64 ;
      RECT 53.916 3.471 54.18 3.64 ;
      RECT 53.96 3.465 53.97 3.662 ;
      RECT 53.97 3.445 54.175 3.648 ;
      RECT 52.925 4.505 53.13 4.735 ;
      RECT 52.865 4.455 52.92 4.715 ;
      RECT 52.925 4.455 53.125 4.735 ;
      RECT 53.895 4.77 53.9 4.797 ;
      RECT 53.885 4.68 53.895 4.802 ;
      RECT 53.88 4.602 53.885 4.808 ;
      RECT 53.87 4.592 53.88 4.815 ;
      RECT 53.865 4.582 53.87 4.821 ;
      RECT 53.855 4.577 53.865 4.823 ;
      RECT 53.84 4.569 53.855 4.831 ;
      RECT 53.825 4.56 53.84 4.843 ;
      RECT 53.815 4.552 53.825 4.853 ;
      RECT 53.78 4.47 53.815 4.871 ;
      RECT 53.745 4.47 53.78 4.89 ;
      RECT 53.73 4.47 53.745 4.898 ;
      RECT 53.675 4.47 53.73 4.898 ;
      RECT 53.641 4.47 53.675 4.889 ;
      RECT 53.555 4.47 53.641 4.865 ;
      RECT 53.545 4.53 53.555 4.847 ;
      RECT 53.505 4.532 53.545 4.838 ;
      RECT 53.5 4.534 53.505 4.828 ;
      RECT 53.48 4.536 53.5 4.823 ;
      RECT 53.47 4.539 53.48 4.818 ;
      RECT 53.46 4.54 53.47 4.813 ;
      RECT 53.436 4.541 53.46 4.805 ;
      RECT 53.35 4.546 53.436 4.783 ;
      RECT 53.295 4.545 53.35 4.756 ;
      RECT 53.28 4.538 53.295 4.743 ;
      RECT 53.245 4.533 53.28 4.739 ;
      RECT 53.19 4.525 53.245 4.738 ;
      RECT 53.13 4.512 53.19 4.736 ;
      RECT 52.92 4.455 52.925 4.723 ;
      RECT 52.995 3.825 53.18 4.035 ;
      RECT 52.985 3.83 53.195 4.028 ;
      RECT 53.025 3.735 53.285 3.995 ;
      RECT 52.98 3.892 53.285 3.918 ;
      RECT 52.325 3.685 52.33 4.485 ;
      RECT 52.27 3.735 52.3 4.485 ;
      RECT 52.26 3.735 52.265 4.045 ;
      RECT 52.245 3.735 52.25 4.04 ;
      RECT 51.79 3.78 51.805 3.995 ;
      RECT 51.72 3.78 51.805 3.99 ;
      RECT 52.985 3.36 53.055 3.57 ;
      RECT 53.055 3.367 53.065 3.565 ;
      RECT 52.951 3.36 52.985 3.577 ;
      RECT 52.865 3.36 52.951 3.601 ;
      RECT 52.855 3.365 52.865 3.62 ;
      RECT 52.85 3.377 52.855 3.623 ;
      RECT 52.835 3.392 52.85 3.627 ;
      RECT 52.83 3.41 52.835 3.631 ;
      RECT 52.79 3.42 52.83 3.64 ;
      RECT 52.775 3.427 52.79 3.652 ;
      RECT 52.76 3.432 52.775 3.657 ;
      RECT 52.745 3.435 52.76 3.662 ;
      RECT 52.735 3.437 52.745 3.666 ;
      RECT 52.7 3.444 52.735 3.674 ;
      RECT 52.665 3.452 52.7 3.688 ;
      RECT 52.655 3.458 52.665 3.697 ;
      RECT 52.65 3.46 52.655 3.699 ;
      RECT 52.63 3.463 52.65 3.705 ;
      RECT 52.6 3.47 52.63 3.716 ;
      RECT 52.59 3.476 52.6 3.723 ;
      RECT 52.565 3.479 52.59 3.73 ;
      RECT 52.555 3.483 52.565 3.738 ;
      RECT 52.55 3.484 52.555 3.76 ;
      RECT 52.545 3.485 52.55 3.775 ;
      RECT 52.54 3.486 52.545 3.79 ;
      RECT 52.535 3.487 52.54 3.805 ;
      RECT 52.53 3.488 52.535 3.835 ;
      RECT 52.52 3.49 52.53 3.868 ;
      RECT 52.505 3.494 52.52 3.915 ;
      RECT 52.495 3.497 52.505 3.96 ;
      RECT 52.49 3.5 52.495 3.988 ;
      RECT 52.48 3.502 52.49 4.015 ;
      RECT 52.475 3.505 52.48 4.05 ;
      RECT 52.445 3.51 52.475 4.108 ;
      RECT 52.44 3.515 52.445 4.193 ;
      RECT 52.435 3.517 52.44 4.228 ;
      RECT 52.43 3.519 52.435 4.31 ;
      RECT 52.425 3.521 52.43 4.398 ;
      RECT 52.415 3.523 52.425 4.48 ;
      RECT 52.4 3.537 52.415 4.485 ;
      RECT 52.365 3.582 52.4 4.485 ;
      RECT 52.355 3.622 52.365 4.485 ;
      RECT 52.34 3.65 52.355 4.485 ;
      RECT 52.335 3.667 52.34 4.485 ;
      RECT 52.33 3.675 52.335 4.485 ;
      RECT 52.32 3.69 52.325 4.485 ;
      RECT 52.315 3.697 52.32 4.485 ;
      RECT 52.305 3.717 52.315 4.485 ;
      RECT 52.3 3.73 52.305 4.485 ;
      RECT 52.265 3.735 52.27 4.07 ;
      RECT 52.25 4.125 52.27 4.485 ;
      RECT 52.25 3.735 52.26 4.043 ;
      RECT 52.245 4.165 52.25 4.485 ;
      RECT 52.195 3.735 52.245 4.038 ;
      RECT 52.24 4.202 52.245 4.485 ;
      RECT 52.23 4.225 52.24 4.485 ;
      RECT 52.225 4.27 52.23 4.485 ;
      RECT 52.215 4.28 52.225 4.478 ;
      RECT 52.141 3.735 52.195 4.032 ;
      RECT 52.055 3.735 52.141 4.025 ;
      RECT 52.006 3.782 52.055 4.018 ;
      RECT 51.92 3.79 52.006 4.011 ;
      RECT 51.905 3.787 51.92 4.006 ;
      RECT 51.891 3.78 51.905 4.005 ;
      RECT 51.805 3.78 51.891 4 ;
      RECT 51.71 3.785 51.72 3.985 ;
      RECT 51.3 3.215 51.315 3.615 ;
      RECT 51.495 3.215 51.5 3.475 ;
      RECT 51.24 3.215 51.285 3.475 ;
      RECT 51.695 4.52 51.7 4.725 ;
      RECT 51.69 4.51 51.695 4.73 ;
      RECT 51.685 4.497 51.69 4.735 ;
      RECT 51.68 4.477 51.685 4.735 ;
      RECT 51.655 4.43 51.68 4.735 ;
      RECT 51.62 4.345 51.655 4.735 ;
      RECT 51.615 4.282 51.62 4.735 ;
      RECT 51.61 4.267 51.615 4.735 ;
      RECT 51.595 4.227 51.61 4.735 ;
      RECT 51.59 4.202 51.595 4.735 ;
      RECT 51.58 4.185 51.59 4.735 ;
      RECT 51.545 4.107 51.58 4.735 ;
      RECT 51.54 4.05 51.545 4.735 ;
      RECT 51.535 4.037 51.54 4.735 ;
      RECT 51.525 4.015 51.535 4.735 ;
      RECT 51.515 3.98 51.525 4.735 ;
      RECT 51.505 3.95 51.515 4.735 ;
      RECT 51.495 3.865 51.505 4.378 ;
      RECT 51.502 4.51 51.505 4.735 ;
      RECT 51.5 4.52 51.502 4.735 ;
      RECT 51.49 4.53 51.5 4.73 ;
      RECT 51.485 3.215 51.495 3.61 ;
      RECT 51.49 3.742 51.495 4.353 ;
      RECT 51.485 3.64 51.49 4.336 ;
      RECT 51.475 3.215 51.485 4.312 ;
      RECT 51.47 3.215 51.475 4.283 ;
      RECT 51.465 3.215 51.47 4.273 ;
      RECT 51.445 3.215 51.465 4.235 ;
      RECT 51.44 3.215 51.445 4.193 ;
      RECT 51.435 3.215 51.44 4.173 ;
      RECT 51.405 3.215 51.435 4.123 ;
      RECT 51.395 3.215 51.405 4.07 ;
      RECT 51.39 3.215 51.395 4.043 ;
      RECT 51.385 3.215 51.39 4.028 ;
      RECT 51.375 3.215 51.385 4.005 ;
      RECT 51.365 3.215 51.375 3.98 ;
      RECT 51.36 3.215 51.365 3.92 ;
      RECT 51.35 3.215 51.36 3.858 ;
      RECT 51.345 3.215 51.35 3.778 ;
      RECT 51.34 3.215 51.345 3.743 ;
      RECT 51.335 3.215 51.34 3.718 ;
      RECT 51.33 3.215 51.335 3.703 ;
      RECT 51.325 3.215 51.33 3.673 ;
      RECT 51.32 3.215 51.325 3.65 ;
      RECT 51.315 3.215 51.32 3.623 ;
      RECT 51.285 3.215 51.3 3.61 ;
      RECT 50.44 4.75 50.625 4.96 ;
      RECT 50.43 4.755 50.64 4.953 ;
      RECT 50.43 4.755 50.66 4.925 ;
      RECT 50.43 4.755 50.675 4.904 ;
      RECT 50.43 4.755 50.69 4.902 ;
      RECT 50.43 4.755 50.7 4.901 ;
      RECT 50.43 4.755 50.73 4.898 ;
      RECT 51.08 4.6 51.34 4.86 ;
      RECT 51.04 4.647 51.34 4.843 ;
      RECT 51.031 4.655 51.04 4.846 ;
      RECT 50.625 4.748 51.34 4.843 ;
      RECT 50.945 4.673 51.031 4.853 ;
      RECT 50.64 4.745 51.34 4.843 ;
      RECT 50.886 4.695 50.945 4.865 ;
      RECT 50.66 4.741 51.34 4.843 ;
      RECT 50.8 4.707 50.886 4.876 ;
      RECT 50.675 4.737 51.34 4.843 ;
      RECT 50.745 4.72 50.8 4.888 ;
      RECT 50.69 4.735 51.34 4.843 ;
      RECT 50.73 4.726 50.745 4.894 ;
      RECT 50.7 4.731 51.34 4.843 ;
      RECT 50.845 4.255 51.105 4.515 ;
      RECT 50.845 4.275 51.215 4.485 ;
      RECT 50.845 4.28 51.225 4.48 ;
      RECT 51.036 3.694 51.115 3.925 ;
      RECT 50.95 3.697 51.165 3.92 ;
      RECT 50.945 3.697 51.165 3.915 ;
      RECT 50.945 3.702 51.175 3.913 ;
      RECT 50.92 3.702 51.175 3.91 ;
      RECT 50.92 3.71 51.185 3.908 ;
      RECT 50.8 3.645 51.06 3.905 ;
      RECT 50.8 3.692 51.11 3.905 ;
      RECT 50.055 4.265 50.06 4.525 ;
      RECT 49.885 4.035 49.89 4.525 ;
      RECT 49.77 4.275 49.775 4.5 ;
      RECT 50.48 3.37 50.485 3.58 ;
      RECT 50.485 3.375 50.5 3.575 ;
      RECT 50.42 3.37 50.48 3.588 ;
      RECT 50.405 3.37 50.42 3.598 ;
      RECT 50.355 3.37 50.405 3.615 ;
      RECT 50.335 3.37 50.355 3.638 ;
      RECT 50.32 3.37 50.335 3.65 ;
      RECT 50.3 3.37 50.32 3.66 ;
      RECT 50.29 3.375 50.3 3.669 ;
      RECT 50.285 3.385 50.29 3.674 ;
      RECT 50.28 3.397 50.285 3.678 ;
      RECT 50.27 3.42 50.28 3.683 ;
      RECT 50.265 3.435 50.27 3.687 ;
      RECT 50.26 3.452 50.265 3.69 ;
      RECT 50.255 3.46 50.26 3.693 ;
      RECT 50.245 3.465 50.255 3.697 ;
      RECT 50.24 3.472 50.245 3.702 ;
      RECT 50.23 3.477 50.24 3.706 ;
      RECT 50.205 3.489 50.23 3.717 ;
      RECT 50.185 3.506 50.205 3.733 ;
      RECT 50.16 3.523 50.185 3.755 ;
      RECT 50.125 3.546 50.16 3.813 ;
      RECT 50.105 3.568 50.125 3.875 ;
      RECT 50.1 3.578 50.105 3.91 ;
      RECT 50.09 3.585 50.1 3.948 ;
      RECT 50.085 3.592 50.09 3.968 ;
      RECT 50.08 3.603 50.085 4.005 ;
      RECT 50.075 3.611 50.08 4.07 ;
      RECT 50.065 3.622 50.075 4.123 ;
      RECT 50.06 3.64 50.065 4.193 ;
      RECT 50.055 3.65 50.06 4.23 ;
      RECT 50.05 3.66 50.055 4.525 ;
      RECT 50.045 3.672 50.05 4.525 ;
      RECT 50.04 3.682 50.045 4.525 ;
      RECT 50.03 3.692 50.04 4.525 ;
      RECT 50.02 3.715 50.03 4.525 ;
      RECT 50.005 3.75 50.02 4.525 ;
      RECT 49.965 3.812 50.005 4.525 ;
      RECT 49.96 3.865 49.965 4.525 ;
      RECT 49.935 3.9 49.96 4.525 ;
      RECT 49.92 3.945 49.935 4.525 ;
      RECT 49.915 3.967 49.92 4.525 ;
      RECT 49.905 3.98 49.915 4.525 ;
      RECT 49.895 4.005 49.905 4.525 ;
      RECT 49.89 4.027 49.895 4.525 ;
      RECT 49.865 4.065 49.885 4.525 ;
      RECT 49.825 4.122 49.865 4.525 ;
      RECT 49.82 4.172 49.825 4.525 ;
      RECT 49.815 4.19 49.82 4.525 ;
      RECT 49.81 4.202 49.815 4.525 ;
      RECT 49.8 4.22 49.81 4.525 ;
      RECT 49.79 4.24 49.8 4.5 ;
      RECT 49.785 4.257 49.79 4.5 ;
      RECT 49.775 4.27 49.785 4.5 ;
      RECT 49.745 4.28 49.77 4.5 ;
      RECT 49.735 4.287 49.745 4.5 ;
      RECT 49.72 4.297 49.735 4.495 ;
      RECT 48.82 10.055 49.115 10.285 ;
      RECT 48.88 8.575 49.05 10.285 ;
      RECT 48.87 8.945 49.225 9.3 ;
      RECT 48.82 8.575 49.11 8.805 ;
      RECT 47.83 10.055 48.125 10.285 ;
      RECT 47.89 8.575 48.06 10.285 ;
      RECT 47.83 8.575 48.12 8.805 ;
      RECT 47.83 8.61 48.68 8.77 ;
      RECT 48.515 8.205 48.68 8.77 ;
      RECT 47.83 8.605 48.225 8.77 ;
      RECT 48.45 8.205 48.74 8.435 ;
      RECT 48.45 8.235 48.91 8.405 ;
      RECT 48.415 4.025 48.735 4.26 ;
      RECT 48.415 4.055 48.905 4.225 ;
      RECT 48.415 3.69 48.605 4.26 ;
      RECT 47.83 3.655 48.12 3.885 ;
      RECT 47.83 3.69 48.605 3.86 ;
      RECT 47.89 2.175 48.06 3.885 ;
      RECT 47.83 2.175 48.125 2.405 ;
      RECT 47.46 4.025 47.75 4.255 ;
      RECT 47.46 4.055 47.92 4.225 ;
      RECT 47.525 2.95 47.69 4.255 ;
      RECT 46.04 2.915 46.33 3.145 ;
      RECT 46.04 2.95 47.69 3.12 ;
      RECT 46.1 2.175 46.27 3.145 ;
      RECT 46.04 2.175 46.33 2.405 ;
      RECT 46.04 10.055 46.33 10.285 ;
      RECT 46.1 9.315 46.27 10.285 ;
      RECT 46.1 9.405 47.69 9.575 ;
      RECT 47.52 8.205 47.69 9.575 ;
      RECT 46.04 9.315 46.33 9.545 ;
      RECT 47.46 8.205 47.75 8.435 ;
      RECT 47.46 8.235 47.92 8.405 ;
      RECT 46.47 3.26 46.82 3.61 ;
      RECT 44.135 3.32 46.82 3.49 ;
      RECT 46.3 3.315 46.82 3.49 ;
      RECT 44.135 2.635 44.305 3.49 ;
      RECT 44.035 2.635 44.385 2.985 ;
      RECT 46.495 8.94 46.82 9.265 ;
      RECT 41.92 8.9 42.27 9.25 ;
      RECT 46.47 8.945 46.82 9.175 ;
      RECT 41.69 8.945 42.27 9.175 ;
      RECT 46.3 8.97 46.82 9.145 ;
      RECT 41.52 8.975 42.27 9.145 ;
      RECT 41.69 8.97 46.82 9.14 ;
      RECT 45.695 3.66 46.015 3.98 ;
      RECT 45.67 3.655 45.96 3.885 ;
      RECT 45.595 3.685 46.015 3.86 ;
      RECT 45.495 3.685 46.015 3.855 ;
      RECT 45.695 8.54 46.015 8.83 ;
      RECT 45.67 8.575 46.015 8.805 ;
      RECT 45.495 8.605 46.015 8.775 ;
      RECT 42.33 3.76 42.515 3.97 ;
      RECT 42.32 3.765 42.53 3.963 ;
      RECT 42.32 3.765 42.616 3.94 ;
      RECT 42.32 3.765 42.675 3.915 ;
      RECT 42.32 3.765 42.73 3.895 ;
      RECT 42.32 3.765 42.74 3.883 ;
      RECT 42.32 3.765 42.935 3.822 ;
      RECT 42.32 3.765 42.965 3.805 ;
      RECT 42.32 3.765 42.985 3.795 ;
      RECT 42.865 3.53 43.125 3.79 ;
      RECT 42.85 3.62 42.865 3.837 ;
      RECT 42.385 3.752 43.125 3.79 ;
      RECT 42.836 3.631 42.85 3.843 ;
      RECT 42.425 3.745 43.125 3.79 ;
      RECT 42.75 3.671 42.836 3.862 ;
      RECT 42.675 3.732 43.125 3.79 ;
      RECT 42.745 3.707 42.75 3.879 ;
      RECT 42.73 3.717 43.125 3.79 ;
      RECT 42.74 3.712 42.745 3.881 ;
      RECT 41.665 3.795 41.77 4.055 ;
      RECT 42.48 3.32 42.485 3.545 ;
      RECT 42.61 3.32 42.665 3.53 ;
      RECT 42.665 3.325 42.675 3.523 ;
      RECT 42.571 3.32 42.61 3.533 ;
      RECT 42.485 3.32 42.571 3.54 ;
      RECT 42.465 3.325 42.48 3.546 ;
      RECT 42.455 3.365 42.465 3.548 ;
      RECT 42.425 3.375 42.455 3.55 ;
      RECT 42.42 3.38 42.425 3.552 ;
      RECT 42.395 3.385 42.42 3.554 ;
      RECT 42.38 3.39 42.395 3.556 ;
      RECT 42.365 3.392 42.38 3.558 ;
      RECT 42.36 3.397 42.365 3.56 ;
      RECT 42.31 3.405 42.36 3.563 ;
      RECT 42.285 3.414 42.31 3.568 ;
      RECT 42.275 3.421 42.285 3.573 ;
      RECT 42.27 3.424 42.275 3.577 ;
      RECT 42.25 3.427 42.27 3.586 ;
      RECT 42.22 3.435 42.25 3.606 ;
      RECT 42.191 3.448 42.22 3.628 ;
      RECT 42.105 3.482 42.191 3.672 ;
      RECT 42.1 3.508 42.105 3.71 ;
      RECT 42.095 3.512 42.1 3.719 ;
      RECT 42.06 3.525 42.095 3.752 ;
      RECT 42.05 3.539 42.06 3.79 ;
      RECT 42.045 3.543 42.05 3.803 ;
      RECT 42.04 3.547 42.045 3.808 ;
      RECT 42.03 3.555 42.04 3.82 ;
      RECT 42.025 3.562 42.03 3.835 ;
      RECT 42 3.575 42.025 3.86 ;
      RECT 41.96 3.604 42 3.915 ;
      RECT 41.945 3.629 41.96 3.97 ;
      RECT 41.935 3.64 41.945 3.993 ;
      RECT 41.93 3.647 41.935 4.005 ;
      RECT 41.925 3.651 41.93 4.013 ;
      RECT 41.87 3.679 41.925 4.055 ;
      RECT 41.85 3.715 41.87 4.055 ;
      RECT 41.835 3.73 41.85 4.055 ;
      RECT 41.78 3.762 41.835 4.055 ;
      RECT 41.77 3.792 41.78 4.055 ;
      RECT 41.38 3.407 41.565 3.645 ;
      RECT 41.365 3.409 41.575 3.64 ;
      RECT 41.25 3.355 41.51 3.615 ;
      RECT 41.245 3.392 41.51 3.569 ;
      RECT 41.24 3.402 41.51 3.566 ;
      RECT 41.235 3.442 41.575 3.56 ;
      RECT 41.23 3.475 41.575 3.55 ;
      RECT 41.24 3.417 41.59 3.488 ;
      RECT 41.537 4.515 41.55 5.045 ;
      RECT 41.451 4.515 41.55 5.044 ;
      RECT 41.451 4.515 41.555 5.043 ;
      RECT 41.365 4.515 41.555 5.041 ;
      RECT 41.36 4.515 41.555 5.038 ;
      RECT 41.36 4.515 41.565 5.036 ;
      RECT 41.355 4.807 41.565 5.033 ;
      RECT 41.355 4.817 41.57 5.03 ;
      RECT 41.355 4.885 41.575 5.026 ;
      RECT 41.345 4.89 41.575 5.025 ;
      RECT 41.345 4.982 41.58 5.022 ;
      RECT 41.33 4.515 41.59 4.775 ;
      RECT 41.26 10.055 41.55 10.285 ;
      RECT 41.32 9.315 41.49 10.285 ;
      RECT 41.235 9.34 41.575 9.685 ;
      RECT 41.26 9.315 41.55 9.685 ;
      RECT 40.56 3.505 40.605 5.04 ;
      RECT 40.76 3.505 40.79 3.72 ;
      RECT 39.135 3.245 39.255 3.455 ;
      RECT 38.795 3.195 39.055 3.455 ;
      RECT 38.795 3.24 39.09 3.445 ;
      RECT 40.8 3.521 40.805 3.575 ;
      RECT 40.795 3.514 40.8 3.708 ;
      RECT 40.79 3.508 40.795 3.715 ;
      RECT 40.745 3.505 40.76 3.728 ;
      RECT 40.74 3.505 40.745 3.75 ;
      RECT 40.735 3.505 40.74 3.798 ;
      RECT 40.73 3.505 40.735 3.818 ;
      RECT 40.72 3.505 40.73 3.925 ;
      RECT 40.715 3.505 40.72 3.988 ;
      RECT 40.71 3.505 40.715 4.045 ;
      RECT 40.705 3.505 40.71 4.053 ;
      RECT 40.69 3.505 40.705 4.16 ;
      RECT 40.68 3.505 40.69 4.295 ;
      RECT 40.67 3.505 40.68 4.405 ;
      RECT 40.66 3.505 40.67 4.462 ;
      RECT 40.655 3.505 40.66 4.502 ;
      RECT 40.65 3.505 40.655 4.538 ;
      RECT 40.64 3.505 40.65 4.578 ;
      RECT 40.635 3.505 40.64 4.62 ;
      RECT 40.615 3.505 40.635 4.685 ;
      RECT 40.62 4.83 40.625 5.01 ;
      RECT 40.615 4.812 40.62 5.018 ;
      RECT 40.61 3.505 40.615 4.748 ;
      RECT 40.61 4.792 40.615 5.025 ;
      RECT 40.605 3.505 40.61 5.035 ;
      RECT 40.55 3.505 40.56 3.805 ;
      RECT 40.555 4.052 40.56 5.04 ;
      RECT 40.55 4.117 40.555 5.04 ;
      RECT 40.545 3.506 40.55 3.795 ;
      RECT 40.54 4.182 40.55 5.04 ;
      RECT 40.535 3.507 40.545 3.785 ;
      RECT 40.525 4.295 40.54 5.04 ;
      RECT 40.53 3.508 40.535 3.775 ;
      RECT 40.51 3.509 40.53 3.753 ;
      RECT 40.515 4.392 40.525 5.04 ;
      RECT 40.51 4.467 40.515 5.04 ;
      RECT 40.5 3.508 40.51 3.73 ;
      RECT 40.505 4.51 40.51 5.04 ;
      RECT 40.5 4.537 40.505 5.04 ;
      RECT 40.49 3.506 40.5 3.718 ;
      RECT 40.495 4.58 40.5 5.04 ;
      RECT 40.49 4.607 40.495 5.04 ;
      RECT 40.48 3.505 40.49 3.705 ;
      RECT 40.485 4.622 40.49 5.04 ;
      RECT 40.445 4.68 40.485 5.04 ;
      RECT 40.475 3.504 40.48 3.69 ;
      RECT 40.47 3.502 40.475 3.683 ;
      RECT 40.46 3.499 40.47 3.673 ;
      RECT 40.455 3.496 40.46 3.658 ;
      RECT 40.44 3.492 40.455 3.651 ;
      RECT 40.435 4.735 40.445 5.04 ;
      RECT 40.435 3.489 40.44 3.646 ;
      RECT 40.42 3.485 40.435 3.64 ;
      RECT 40.43 4.752 40.435 5.04 ;
      RECT 40.42 4.815 40.43 5.04 ;
      RECT 40.34 3.47 40.42 3.62 ;
      RECT 40.415 4.822 40.42 5.035 ;
      RECT 40.41 4.83 40.415 5.025 ;
      RECT 40.33 3.456 40.34 3.604 ;
      RECT 40.315 3.452 40.33 3.602 ;
      RECT 40.305 3.447 40.315 3.598 ;
      RECT 40.28 3.44 40.305 3.59 ;
      RECT 40.275 3.435 40.28 3.585 ;
      RECT 40.265 3.435 40.275 3.583 ;
      RECT 40.255 3.433 40.265 3.581 ;
      RECT 40.225 3.425 40.255 3.575 ;
      RECT 40.21 3.417 40.225 3.568 ;
      RECT 40.19 3.412 40.21 3.561 ;
      RECT 40.185 3.408 40.19 3.556 ;
      RECT 40.155 3.401 40.185 3.55 ;
      RECT 40.13 3.392 40.155 3.54 ;
      RECT 40.1 3.385 40.13 3.532 ;
      RECT 40.075 3.375 40.1 3.523 ;
      RECT 40.06 3.367 40.075 3.517 ;
      RECT 40.035 3.362 40.06 3.512 ;
      RECT 40.025 3.358 40.035 3.507 ;
      RECT 40.005 3.353 40.025 3.502 ;
      RECT 39.97 3.348 40.005 3.495 ;
      RECT 39.91 3.343 39.97 3.488 ;
      RECT 39.897 3.339 39.91 3.486 ;
      RECT 39.811 3.334 39.897 3.483 ;
      RECT 39.725 3.324 39.811 3.479 ;
      RECT 39.684 3.317 39.725 3.476 ;
      RECT 39.598 3.31 39.684 3.473 ;
      RECT 39.512 3.3 39.598 3.469 ;
      RECT 39.426 3.29 39.512 3.464 ;
      RECT 39.34 3.28 39.426 3.46 ;
      RECT 39.33 3.265 39.34 3.458 ;
      RECT 39.32 3.25 39.33 3.458 ;
      RECT 39.255 3.245 39.32 3.457 ;
      RECT 39.09 3.242 39.135 3.45 ;
      RECT 40.335 4.147 40.34 4.338 ;
      RECT 40.33 4.142 40.335 4.345 ;
      RECT 40.316 4.14 40.33 4.351 ;
      RECT 40.23 4.14 40.316 4.353 ;
      RECT 40.226 4.14 40.23 4.356 ;
      RECT 40.14 4.14 40.226 4.374 ;
      RECT 40.13 4.145 40.14 4.393 ;
      RECT 40.12 4.2 40.13 4.397 ;
      RECT 40.095 4.215 40.12 4.404 ;
      RECT 40.055 4.235 40.095 4.417 ;
      RECT 40.05 4.247 40.055 4.427 ;
      RECT 40.035 4.253 40.05 4.432 ;
      RECT 40.03 4.258 40.035 4.436 ;
      RECT 40.01 4.265 40.03 4.441 ;
      RECT 39.94 4.29 40.01 4.458 ;
      RECT 39.9 4.318 39.94 4.478 ;
      RECT 39.895 4.328 39.9 4.486 ;
      RECT 39.875 4.335 39.895 4.488 ;
      RECT 39.87 4.342 39.875 4.491 ;
      RECT 39.84 4.35 39.87 4.494 ;
      RECT 39.835 4.355 39.84 4.498 ;
      RECT 39.761 4.359 39.835 4.506 ;
      RECT 39.675 4.368 39.761 4.522 ;
      RECT 39.671 4.373 39.675 4.531 ;
      RECT 39.585 4.378 39.671 4.541 ;
      RECT 39.545 4.386 39.585 4.553 ;
      RECT 39.495 4.392 39.545 4.56 ;
      RECT 39.41 4.401 39.495 4.575 ;
      RECT 39.335 4.412 39.41 4.593 ;
      RECT 39.3 4.419 39.335 4.603 ;
      RECT 39.225 4.427 39.3 4.608 ;
      RECT 39.17 4.436 39.225 4.608 ;
      RECT 39.145 4.441 39.17 4.606 ;
      RECT 39.135 4.444 39.145 4.604 ;
      RECT 39.1 4.446 39.135 4.602 ;
      RECT 39.07 4.448 39.1 4.598 ;
      RECT 39.025 4.447 39.07 4.594 ;
      RECT 39.005 4.442 39.025 4.591 ;
      RECT 38.955 4.427 39.005 4.588 ;
      RECT 38.945 4.412 38.955 4.583 ;
      RECT 38.895 4.397 38.945 4.573 ;
      RECT 38.845 4.372 38.895 4.553 ;
      RECT 38.835 4.357 38.845 4.535 ;
      RECT 38.83 4.355 38.835 4.529 ;
      RECT 38.81 4.35 38.83 4.524 ;
      RECT 38.805 4.342 38.81 4.518 ;
      RECT 38.79 4.336 38.805 4.511 ;
      RECT 38.785 4.331 38.79 4.503 ;
      RECT 38.765 4.326 38.785 4.495 ;
      RECT 38.75 4.319 38.765 4.488 ;
      RECT 38.735 4.313 38.75 4.479 ;
      RECT 38.73 4.307 38.735 4.472 ;
      RECT 38.685 4.282 38.73 4.458 ;
      RECT 38.67 4.252 38.685 4.44 ;
      RECT 38.655 4.235 38.67 4.431 ;
      RECT 38.63 4.215 38.655 4.419 ;
      RECT 38.59 4.185 38.63 4.399 ;
      RECT 38.58 4.155 38.59 4.384 ;
      RECT 38.565 4.145 38.58 4.377 ;
      RECT 38.51 4.11 38.565 4.356 ;
      RECT 38.495 4.073 38.51 4.335 ;
      RECT 38.485 4.06 38.495 4.327 ;
      RECT 38.435 4.03 38.485 4.309 ;
      RECT 38.42 3.96 38.435 4.29 ;
      RECT 38.375 3.96 38.42 4.273 ;
      RECT 38.35 3.96 38.375 4.255 ;
      RECT 38.34 3.96 38.35 4.248 ;
      RECT 38.261 3.96 38.34 4.241 ;
      RECT 38.175 3.96 38.261 4.233 ;
      RECT 38.16 3.992 38.175 4.228 ;
      RECT 38.085 4.002 38.16 4.224 ;
      RECT 38.065 4.012 38.085 4.219 ;
      RECT 38.04 4.012 38.065 4.216 ;
      RECT 38.03 4.002 38.04 4.215 ;
      RECT 38.02 3.975 38.03 4.214 ;
      RECT 37.98 3.97 38.02 4.212 ;
      RECT 37.935 3.97 37.98 4.208 ;
      RECT 37.91 3.97 37.935 4.203 ;
      RECT 37.86 3.97 37.91 4.19 ;
      RECT 37.82 3.975 37.83 4.175 ;
      RECT 37.83 3.97 37.86 4.18 ;
      RECT 39.815 3.75 40.075 4.01 ;
      RECT 39.81 3.772 40.075 3.968 ;
      RECT 39.05 3.6 39.27 3.965 ;
      RECT 39.032 3.687 39.27 3.964 ;
      RECT 39.015 3.692 39.27 3.961 ;
      RECT 39.015 3.692 39.29 3.96 ;
      RECT 38.985 3.702 39.29 3.958 ;
      RECT 38.98 3.717 39.29 3.954 ;
      RECT 38.98 3.717 39.295 3.953 ;
      RECT 38.975 3.775 39.295 3.951 ;
      RECT 38.975 3.775 39.305 3.948 ;
      RECT 38.97 3.84 39.305 3.943 ;
      RECT 39.05 3.6 39.31 3.86 ;
      RECT 37.795 3.43 38.055 3.69 ;
      RECT 37.795 3.473 38.141 3.664 ;
      RECT 37.795 3.473 38.185 3.663 ;
      RECT 37.795 3.473 38.205 3.661 ;
      RECT 37.795 3.473 38.305 3.66 ;
      RECT 37.795 3.473 38.325 3.658 ;
      RECT 37.795 3.473 38.335 3.653 ;
      RECT 38.205 3.44 38.395 3.65 ;
      RECT 38.205 3.442 38.4 3.648 ;
      RECT 38.195 3.447 38.405 3.64 ;
      RECT 38.141 3.471 38.405 3.64 ;
      RECT 38.185 3.465 38.195 3.662 ;
      RECT 38.195 3.445 38.4 3.648 ;
      RECT 37.15 4.505 37.355 4.735 ;
      RECT 37.09 4.455 37.145 4.715 ;
      RECT 37.15 4.455 37.35 4.735 ;
      RECT 38.12 4.77 38.125 4.797 ;
      RECT 38.11 4.68 38.12 4.802 ;
      RECT 38.105 4.602 38.11 4.808 ;
      RECT 38.095 4.592 38.105 4.815 ;
      RECT 38.09 4.582 38.095 4.821 ;
      RECT 38.08 4.577 38.09 4.823 ;
      RECT 38.065 4.569 38.08 4.831 ;
      RECT 38.05 4.56 38.065 4.843 ;
      RECT 38.04 4.552 38.05 4.853 ;
      RECT 38.005 4.47 38.04 4.871 ;
      RECT 37.97 4.47 38.005 4.89 ;
      RECT 37.955 4.47 37.97 4.898 ;
      RECT 37.9 4.47 37.955 4.898 ;
      RECT 37.866 4.47 37.9 4.889 ;
      RECT 37.78 4.47 37.866 4.865 ;
      RECT 37.77 4.53 37.78 4.847 ;
      RECT 37.73 4.532 37.77 4.838 ;
      RECT 37.725 4.534 37.73 4.828 ;
      RECT 37.705 4.536 37.725 4.823 ;
      RECT 37.695 4.539 37.705 4.818 ;
      RECT 37.685 4.54 37.695 4.813 ;
      RECT 37.661 4.541 37.685 4.805 ;
      RECT 37.575 4.546 37.661 4.783 ;
      RECT 37.52 4.545 37.575 4.756 ;
      RECT 37.505 4.538 37.52 4.743 ;
      RECT 37.47 4.533 37.505 4.739 ;
      RECT 37.415 4.525 37.47 4.738 ;
      RECT 37.355 4.512 37.415 4.736 ;
      RECT 37.145 4.455 37.15 4.723 ;
      RECT 37.22 3.825 37.405 4.035 ;
      RECT 37.21 3.83 37.42 4.028 ;
      RECT 37.25 3.735 37.51 3.995 ;
      RECT 37.205 3.892 37.51 3.918 ;
      RECT 36.55 3.685 36.555 4.485 ;
      RECT 36.495 3.735 36.525 4.485 ;
      RECT 36.485 3.735 36.49 4.045 ;
      RECT 36.47 3.735 36.475 4.04 ;
      RECT 36.015 3.78 36.03 3.995 ;
      RECT 35.945 3.78 36.03 3.99 ;
      RECT 37.21 3.36 37.28 3.57 ;
      RECT 37.28 3.367 37.29 3.565 ;
      RECT 37.176 3.36 37.21 3.577 ;
      RECT 37.09 3.36 37.176 3.601 ;
      RECT 37.08 3.365 37.09 3.62 ;
      RECT 37.075 3.377 37.08 3.623 ;
      RECT 37.06 3.392 37.075 3.627 ;
      RECT 37.055 3.41 37.06 3.631 ;
      RECT 37.015 3.42 37.055 3.64 ;
      RECT 37 3.427 37.015 3.652 ;
      RECT 36.985 3.432 37 3.657 ;
      RECT 36.97 3.435 36.985 3.662 ;
      RECT 36.96 3.437 36.97 3.666 ;
      RECT 36.925 3.444 36.96 3.674 ;
      RECT 36.89 3.452 36.925 3.688 ;
      RECT 36.88 3.458 36.89 3.697 ;
      RECT 36.875 3.46 36.88 3.699 ;
      RECT 36.855 3.463 36.875 3.705 ;
      RECT 36.825 3.47 36.855 3.716 ;
      RECT 36.815 3.476 36.825 3.723 ;
      RECT 36.79 3.479 36.815 3.73 ;
      RECT 36.78 3.483 36.79 3.738 ;
      RECT 36.775 3.484 36.78 3.76 ;
      RECT 36.77 3.485 36.775 3.775 ;
      RECT 36.765 3.486 36.77 3.79 ;
      RECT 36.76 3.487 36.765 3.805 ;
      RECT 36.755 3.488 36.76 3.835 ;
      RECT 36.745 3.49 36.755 3.868 ;
      RECT 36.73 3.494 36.745 3.915 ;
      RECT 36.72 3.497 36.73 3.96 ;
      RECT 36.715 3.5 36.72 3.988 ;
      RECT 36.705 3.502 36.715 4.015 ;
      RECT 36.7 3.505 36.705 4.05 ;
      RECT 36.67 3.51 36.7 4.108 ;
      RECT 36.665 3.515 36.67 4.193 ;
      RECT 36.66 3.517 36.665 4.228 ;
      RECT 36.655 3.519 36.66 4.31 ;
      RECT 36.65 3.521 36.655 4.398 ;
      RECT 36.64 3.523 36.65 4.48 ;
      RECT 36.625 3.537 36.64 4.485 ;
      RECT 36.59 3.582 36.625 4.485 ;
      RECT 36.58 3.622 36.59 4.485 ;
      RECT 36.565 3.65 36.58 4.485 ;
      RECT 36.56 3.667 36.565 4.485 ;
      RECT 36.555 3.675 36.56 4.485 ;
      RECT 36.545 3.69 36.55 4.485 ;
      RECT 36.54 3.697 36.545 4.485 ;
      RECT 36.53 3.717 36.54 4.485 ;
      RECT 36.525 3.73 36.53 4.485 ;
      RECT 36.49 3.735 36.495 4.07 ;
      RECT 36.475 4.125 36.495 4.485 ;
      RECT 36.475 3.735 36.485 4.043 ;
      RECT 36.47 4.165 36.475 4.485 ;
      RECT 36.42 3.735 36.47 4.038 ;
      RECT 36.465 4.202 36.47 4.485 ;
      RECT 36.455 4.225 36.465 4.485 ;
      RECT 36.45 4.27 36.455 4.485 ;
      RECT 36.44 4.28 36.45 4.478 ;
      RECT 36.366 3.735 36.42 4.032 ;
      RECT 36.28 3.735 36.366 4.025 ;
      RECT 36.231 3.782 36.28 4.018 ;
      RECT 36.145 3.79 36.231 4.011 ;
      RECT 36.13 3.787 36.145 4.006 ;
      RECT 36.116 3.78 36.13 4.005 ;
      RECT 36.03 3.78 36.116 4 ;
      RECT 35.935 3.785 35.945 3.985 ;
      RECT 35.525 3.215 35.54 3.615 ;
      RECT 35.72 3.215 35.725 3.475 ;
      RECT 35.465 3.215 35.51 3.475 ;
      RECT 35.92 4.52 35.925 4.725 ;
      RECT 35.915 4.51 35.92 4.73 ;
      RECT 35.91 4.497 35.915 4.735 ;
      RECT 35.905 4.477 35.91 4.735 ;
      RECT 35.88 4.43 35.905 4.735 ;
      RECT 35.845 4.345 35.88 4.735 ;
      RECT 35.84 4.282 35.845 4.735 ;
      RECT 35.835 4.267 35.84 4.735 ;
      RECT 35.82 4.227 35.835 4.735 ;
      RECT 35.815 4.202 35.82 4.735 ;
      RECT 35.805 4.185 35.815 4.735 ;
      RECT 35.77 4.107 35.805 4.735 ;
      RECT 35.765 4.05 35.77 4.735 ;
      RECT 35.76 4.037 35.765 4.735 ;
      RECT 35.75 4.015 35.76 4.735 ;
      RECT 35.74 3.98 35.75 4.735 ;
      RECT 35.73 3.95 35.74 4.735 ;
      RECT 35.72 3.865 35.73 4.378 ;
      RECT 35.727 4.51 35.73 4.735 ;
      RECT 35.725 4.52 35.727 4.735 ;
      RECT 35.715 4.53 35.725 4.73 ;
      RECT 35.71 3.215 35.72 3.61 ;
      RECT 35.715 3.742 35.72 4.353 ;
      RECT 35.71 3.64 35.715 4.336 ;
      RECT 35.7 3.215 35.71 4.312 ;
      RECT 35.695 3.215 35.7 4.283 ;
      RECT 35.69 3.215 35.695 4.273 ;
      RECT 35.67 3.215 35.69 4.235 ;
      RECT 35.665 3.215 35.67 4.193 ;
      RECT 35.66 3.215 35.665 4.173 ;
      RECT 35.63 3.215 35.66 4.123 ;
      RECT 35.62 3.215 35.63 4.07 ;
      RECT 35.615 3.215 35.62 4.043 ;
      RECT 35.61 3.215 35.615 4.028 ;
      RECT 35.6 3.215 35.61 4.005 ;
      RECT 35.59 3.215 35.6 3.98 ;
      RECT 35.585 3.215 35.59 3.92 ;
      RECT 35.575 3.215 35.585 3.858 ;
      RECT 35.57 3.215 35.575 3.778 ;
      RECT 35.565 3.215 35.57 3.743 ;
      RECT 35.56 3.215 35.565 3.718 ;
      RECT 35.555 3.215 35.56 3.703 ;
      RECT 35.55 3.215 35.555 3.673 ;
      RECT 35.545 3.215 35.55 3.65 ;
      RECT 35.54 3.215 35.545 3.623 ;
      RECT 35.51 3.215 35.525 3.61 ;
      RECT 34.665 4.75 34.85 4.96 ;
      RECT 34.655 4.755 34.865 4.953 ;
      RECT 34.655 4.755 34.885 4.925 ;
      RECT 34.655 4.755 34.9 4.904 ;
      RECT 34.655 4.755 34.915 4.902 ;
      RECT 34.655 4.755 34.925 4.901 ;
      RECT 34.655 4.755 34.955 4.898 ;
      RECT 35.305 4.6 35.565 4.86 ;
      RECT 35.265 4.647 35.565 4.843 ;
      RECT 35.256 4.655 35.265 4.846 ;
      RECT 34.85 4.748 35.565 4.843 ;
      RECT 35.17 4.673 35.256 4.853 ;
      RECT 34.865 4.745 35.565 4.843 ;
      RECT 35.111 4.695 35.17 4.865 ;
      RECT 34.885 4.741 35.565 4.843 ;
      RECT 35.025 4.707 35.111 4.876 ;
      RECT 34.9 4.737 35.565 4.843 ;
      RECT 34.97 4.72 35.025 4.888 ;
      RECT 34.915 4.735 35.565 4.843 ;
      RECT 34.955 4.726 34.97 4.894 ;
      RECT 34.925 4.731 35.565 4.843 ;
      RECT 35.07 4.255 35.33 4.515 ;
      RECT 35.07 4.275 35.44 4.485 ;
      RECT 35.07 4.28 35.45 4.48 ;
      RECT 35.261 3.694 35.34 3.925 ;
      RECT 35.175 3.697 35.39 3.92 ;
      RECT 35.17 3.697 35.39 3.915 ;
      RECT 35.17 3.702 35.4 3.913 ;
      RECT 35.145 3.702 35.4 3.91 ;
      RECT 35.145 3.71 35.41 3.908 ;
      RECT 35.025 3.645 35.285 3.905 ;
      RECT 35.025 3.692 35.335 3.905 ;
      RECT 34.28 4.265 34.285 4.525 ;
      RECT 34.11 4.035 34.115 4.525 ;
      RECT 33.995 4.275 34 4.5 ;
      RECT 34.705 3.37 34.71 3.58 ;
      RECT 34.71 3.375 34.725 3.575 ;
      RECT 34.645 3.37 34.705 3.588 ;
      RECT 34.63 3.37 34.645 3.598 ;
      RECT 34.58 3.37 34.63 3.615 ;
      RECT 34.56 3.37 34.58 3.638 ;
      RECT 34.545 3.37 34.56 3.65 ;
      RECT 34.525 3.37 34.545 3.66 ;
      RECT 34.515 3.375 34.525 3.669 ;
      RECT 34.51 3.385 34.515 3.674 ;
      RECT 34.505 3.397 34.51 3.678 ;
      RECT 34.495 3.42 34.505 3.683 ;
      RECT 34.49 3.435 34.495 3.687 ;
      RECT 34.485 3.452 34.49 3.69 ;
      RECT 34.48 3.46 34.485 3.693 ;
      RECT 34.47 3.465 34.48 3.697 ;
      RECT 34.465 3.472 34.47 3.702 ;
      RECT 34.455 3.477 34.465 3.706 ;
      RECT 34.43 3.489 34.455 3.717 ;
      RECT 34.41 3.506 34.43 3.733 ;
      RECT 34.385 3.523 34.41 3.755 ;
      RECT 34.35 3.546 34.385 3.813 ;
      RECT 34.33 3.568 34.35 3.875 ;
      RECT 34.325 3.578 34.33 3.91 ;
      RECT 34.315 3.585 34.325 3.948 ;
      RECT 34.31 3.592 34.315 3.968 ;
      RECT 34.305 3.603 34.31 4.005 ;
      RECT 34.3 3.611 34.305 4.07 ;
      RECT 34.29 3.622 34.3 4.123 ;
      RECT 34.285 3.64 34.29 4.193 ;
      RECT 34.28 3.65 34.285 4.23 ;
      RECT 34.275 3.66 34.28 4.525 ;
      RECT 34.27 3.672 34.275 4.525 ;
      RECT 34.265 3.682 34.27 4.525 ;
      RECT 34.255 3.692 34.265 4.525 ;
      RECT 34.245 3.715 34.255 4.525 ;
      RECT 34.23 3.75 34.245 4.525 ;
      RECT 34.19 3.812 34.23 4.525 ;
      RECT 34.185 3.865 34.19 4.525 ;
      RECT 34.16 3.9 34.185 4.525 ;
      RECT 34.145 3.945 34.16 4.525 ;
      RECT 34.14 3.967 34.145 4.525 ;
      RECT 34.13 3.98 34.14 4.525 ;
      RECT 34.12 4.005 34.13 4.525 ;
      RECT 34.115 4.027 34.12 4.525 ;
      RECT 34.09 4.065 34.11 4.525 ;
      RECT 34.05 4.122 34.09 4.525 ;
      RECT 34.045 4.172 34.05 4.525 ;
      RECT 34.04 4.19 34.045 4.525 ;
      RECT 34.035 4.202 34.04 4.525 ;
      RECT 34.025 4.22 34.035 4.525 ;
      RECT 34.015 4.24 34.025 4.5 ;
      RECT 34.01 4.257 34.015 4.5 ;
      RECT 34 4.27 34.01 4.5 ;
      RECT 33.97 4.28 33.995 4.5 ;
      RECT 33.96 4.287 33.97 4.5 ;
      RECT 33.945 4.297 33.96 4.495 ;
      RECT 33.04 10.055 33.335 10.285 ;
      RECT 33.1 8.575 33.27 10.285 ;
      RECT 33.095 8.945 33.445 9.295 ;
      RECT 33.04 8.575 33.33 8.805 ;
      RECT 32.05 10.055 32.345 10.285 ;
      RECT 32.11 8.575 32.28 10.285 ;
      RECT 32.05 8.575 32.34 8.805 ;
      RECT 32.05 8.61 32.9 8.77 ;
      RECT 32.735 8.205 32.9 8.77 ;
      RECT 32.05 8.605 32.445 8.77 ;
      RECT 32.67 8.205 32.96 8.435 ;
      RECT 32.67 8.235 33.13 8.405 ;
      RECT 32.635 4.025 32.955 4.26 ;
      RECT 32.635 4.055 33.125 4.225 ;
      RECT 32.635 3.69 32.825 4.26 ;
      RECT 32.05 3.655 32.34 3.885 ;
      RECT 32.05 3.69 32.825 3.86 ;
      RECT 32.11 2.175 32.28 3.885 ;
      RECT 32.05 2.175 32.345 2.405 ;
      RECT 31.68 4.025 31.97 4.255 ;
      RECT 31.68 4.055 32.14 4.225 ;
      RECT 31.745 2.95 31.91 4.255 ;
      RECT 30.26 2.915 30.55 3.145 ;
      RECT 30.26 2.95 31.91 3.12 ;
      RECT 30.32 2.175 30.49 3.145 ;
      RECT 30.26 2.175 30.55 2.405 ;
      RECT 30.26 10.055 30.55 10.285 ;
      RECT 30.32 9.315 30.49 10.285 ;
      RECT 30.32 9.405 31.91 9.575 ;
      RECT 31.74 8.205 31.91 9.575 ;
      RECT 30.26 9.315 30.55 9.545 ;
      RECT 31.68 8.205 31.97 8.435 ;
      RECT 31.68 8.235 32.14 8.405 ;
      RECT 30.69 3.26 31.04 3.61 ;
      RECT 28.355 3.32 31.04 3.49 ;
      RECT 30.52 3.315 31.04 3.49 ;
      RECT 28.355 2.635 28.525 3.49 ;
      RECT 28.255 2.635 28.605 2.985 ;
      RECT 30.715 8.94 31.04 9.265 ;
      RECT 26.11 8.89 26.46 9.24 ;
      RECT 30.69 8.945 31.04 9.175 ;
      RECT 25.91 8.945 26.46 9.175 ;
      RECT 30.52 8.97 31.04 9.145 ;
      RECT 25.74 8.975 26.46 9.145 ;
      RECT 25.91 8.97 31.04 9.14 ;
      RECT 29.915 3.66 30.235 3.98 ;
      RECT 29.89 3.655 30.18 3.885 ;
      RECT 29.815 3.685 30.235 3.86 ;
      RECT 29.715 3.685 30.235 3.855 ;
      RECT 29.915 8.54 30.235 8.83 ;
      RECT 29.89 8.575 30.235 8.805 ;
      RECT 29.715 8.605 30.235 8.775 ;
      RECT 26.55 3.76 26.735 3.97 ;
      RECT 26.54 3.765 26.75 3.963 ;
      RECT 26.54 3.765 26.836 3.94 ;
      RECT 26.54 3.765 26.895 3.915 ;
      RECT 26.54 3.765 26.95 3.895 ;
      RECT 26.54 3.765 26.96 3.883 ;
      RECT 26.54 3.765 27.155 3.822 ;
      RECT 26.54 3.765 27.185 3.805 ;
      RECT 26.54 3.765 27.205 3.795 ;
      RECT 27.085 3.53 27.345 3.79 ;
      RECT 27.07 3.62 27.085 3.837 ;
      RECT 26.605 3.752 27.345 3.79 ;
      RECT 27.056 3.631 27.07 3.843 ;
      RECT 26.645 3.745 27.345 3.79 ;
      RECT 26.97 3.671 27.056 3.862 ;
      RECT 26.895 3.732 27.345 3.79 ;
      RECT 26.965 3.707 26.97 3.879 ;
      RECT 26.95 3.717 27.345 3.79 ;
      RECT 26.96 3.712 26.965 3.881 ;
      RECT 25.885 3.795 25.99 4.055 ;
      RECT 26.7 3.32 26.705 3.545 ;
      RECT 26.83 3.32 26.885 3.53 ;
      RECT 26.885 3.325 26.895 3.523 ;
      RECT 26.791 3.32 26.83 3.533 ;
      RECT 26.705 3.32 26.791 3.54 ;
      RECT 26.685 3.325 26.7 3.546 ;
      RECT 26.675 3.365 26.685 3.548 ;
      RECT 26.645 3.375 26.675 3.55 ;
      RECT 26.64 3.38 26.645 3.552 ;
      RECT 26.615 3.385 26.64 3.554 ;
      RECT 26.6 3.39 26.615 3.556 ;
      RECT 26.585 3.392 26.6 3.558 ;
      RECT 26.58 3.397 26.585 3.56 ;
      RECT 26.53 3.405 26.58 3.563 ;
      RECT 26.505 3.414 26.53 3.568 ;
      RECT 26.495 3.421 26.505 3.573 ;
      RECT 26.49 3.424 26.495 3.577 ;
      RECT 26.47 3.427 26.49 3.586 ;
      RECT 26.44 3.435 26.47 3.606 ;
      RECT 26.411 3.448 26.44 3.628 ;
      RECT 26.325 3.482 26.411 3.672 ;
      RECT 26.32 3.508 26.325 3.71 ;
      RECT 26.315 3.512 26.32 3.719 ;
      RECT 26.28 3.525 26.315 3.752 ;
      RECT 26.27 3.539 26.28 3.79 ;
      RECT 26.265 3.543 26.27 3.803 ;
      RECT 26.26 3.547 26.265 3.808 ;
      RECT 26.25 3.555 26.26 3.82 ;
      RECT 26.245 3.562 26.25 3.835 ;
      RECT 26.22 3.575 26.245 3.86 ;
      RECT 26.18 3.604 26.22 3.915 ;
      RECT 26.165 3.629 26.18 3.97 ;
      RECT 26.155 3.64 26.165 3.993 ;
      RECT 26.15 3.647 26.155 4.005 ;
      RECT 26.145 3.651 26.15 4.013 ;
      RECT 26.09 3.679 26.145 4.055 ;
      RECT 26.07 3.715 26.09 4.055 ;
      RECT 26.055 3.73 26.07 4.055 ;
      RECT 26 3.762 26.055 4.055 ;
      RECT 25.99 3.792 26 4.055 ;
      RECT 25.6 3.407 25.785 3.645 ;
      RECT 25.585 3.409 25.795 3.64 ;
      RECT 25.47 3.355 25.73 3.615 ;
      RECT 25.465 3.392 25.73 3.569 ;
      RECT 25.46 3.402 25.73 3.566 ;
      RECT 25.455 3.442 25.795 3.56 ;
      RECT 25.45 3.475 25.795 3.55 ;
      RECT 25.46 3.417 25.81 3.488 ;
      RECT 25.757 4.515 25.77 5.045 ;
      RECT 25.671 4.515 25.77 5.044 ;
      RECT 25.671 4.515 25.775 5.043 ;
      RECT 25.585 4.515 25.775 5.041 ;
      RECT 25.58 4.515 25.775 5.038 ;
      RECT 25.58 4.515 25.785 5.036 ;
      RECT 25.575 4.807 25.785 5.033 ;
      RECT 25.575 4.817 25.79 5.03 ;
      RECT 25.575 4.885 25.795 5.026 ;
      RECT 25.565 4.89 25.795 5.025 ;
      RECT 25.565 4.982 25.8 5.022 ;
      RECT 25.55 4.515 25.81 4.775 ;
      RECT 25.48 10.055 25.77 10.285 ;
      RECT 25.54 9.315 25.71 10.285 ;
      RECT 25.455 9.34 25.795 9.685 ;
      RECT 25.48 9.315 25.77 9.685 ;
      RECT 24.78 3.505 24.825 5.04 ;
      RECT 24.98 3.505 25.01 3.72 ;
      RECT 23.355 3.245 23.475 3.455 ;
      RECT 23.015 3.195 23.275 3.455 ;
      RECT 23.015 3.24 23.31 3.445 ;
      RECT 25.02 3.521 25.025 3.575 ;
      RECT 25.015 3.514 25.02 3.708 ;
      RECT 25.01 3.508 25.015 3.715 ;
      RECT 24.965 3.505 24.98 3.728 ;
      RECT 24.96 3.505 24.965 3.75 ;
      RECT 24.955 3.505 24.96 3.798 ;
      RECT 24.95 3.505 24.955 3.818 ;
      RECT 24.94 3.505 24.95 3.925 ;
      RECT 24.935 3.505 24.94 3.988 ;
      RECT 24.93 3.505 24.935 4.045 ;
      RECT 24.925 3.505 24.93 4.053 ;
      RECT 24.91 3.505 24.925 4.16 ;
      RECT 24.9 3.505 24.91 4.295 ;
      RECT 24.89 3.505 24.9 4.405 ;
      RECT 24.88 3.505 24.89 4.462 ;
      RECT 24.875 3.505 24.88 4.502 ;
      RECT 24.87 3.505 24.875 4.538 ;
      RECT 24.86 3.505 24.87 4.578 ;
      RECT 24.855 3.505 24.86 4.62 ;
      RECT 24.835 3.505 24.855 4.685 ;
      RECT 24.84 4.83 24.845 5.01 ;
      RECT 24.835 4.812 24.84 5.018 ;
      RECT 24.83 3.505 24.835 4.748 ;
      RECT 24.83 4.792 24.835 5.025 ;
      RECT 24.825 3.505 24.83 5.035 ;
      RECT 24.77 3.505 24.78 3.805 ;
      RECT 24.775 4.052 24.78 5.04 ;
      RECT 24.77 4.117 24.775 5.04 ;
      RECT 24.765 3.506 24.77 3.795 ;
      RECT 24.76 4.182 24.77 5.04 ;
      RECT 24.755 3.507 24.765 3.785 ;
      RECT 24.745 4.295 24.76 5.04 ;
      RECT 24.75 3.508 24.755 3.775 ;
      RECT 24.73 3.509 24.75 3.753 ;
      RECT 24.735 4.392 24.745 5.04 ;
      RECT 24.73 4.467 24.735 5.04 ;
      RECT 24.72 3.508 24.73 3.73 ;
      RECT 24.725 4.51 24.73 5.04 ;
      RECT 24.72 4.537 24.725 5.04 ;
      RECT 24.71 3.506 24.72 3.718 ;
      RECT 24.715 4.58 24.72 5.04 ;
      RECT 24.71 4.607 24.715 5.04 ;
      RECT 24.7 3.505 24.71 3.705 ;
      RECT 24.705 4.622 24.71 5.04 ;
      RECT 24.665 4.68 24.705 5.04 ;
      RECT 24.695 3.504 24.7 3.69 ;
      RECT 24.69 3.502 24.695 3.683 ;
      RECT 24.68 3.499 24.69 3.673 ;
      RECT 24.675 3.496 24.68 3.658 ;
      RECT 24.66 3.492 24.675 3.651 ;
      RECT 24.655 4.735 24.665 5.04 ;
      RECT 24.655 3.489 24.66 3.646 ;
      RECT 24.64 3.485 24.655 3.64 ;
      RECT 24.65 4.752 24.655 5.04 ;
      RECT 24.64 4.815 24.65 5.04 ;
      RECT 24.56 3.47 24.64 3.62 ;
      RECT 24.635 4.822 24.64 5.035 ;
      RECT 24.63 4.83 24.635 5.025 ;
      RECT 24.55 3.456 24.56 3.604 ;
      RECT 24.535 3.452 24.55 3.602 ;
      RECT 24.525 3.447 24.535 3.598 ;
      RECT 24.5 3.44 24.525 3.59 ;
      RECT 24.495 3.435 24.5 3.585 ;
      RECT 24.485 3.435 24.495 3.583 ;
      RECT 24.475 3.433 24.485 3.581 ;
      RECT 24.445 3.425 24.475 3.575 ;
      RECT 24.43 3.417 24.445 3.568 ;
      RECT 24.41 3.412 24.43 3.561 ;
      RECT 24.405 3.408 24.41 3.556 ;
      RECT 24.375 3.401 24.405 3.55 ;
      RECT 24.35 3.392 24.375 3.54 ;
      RECT 24.32 3.385 24.35 3.532 ;
      RECT 24.295 3.375 24.32 3.523 ;
      RECT 24.28 3.367 24.295 3.517 ;
      RECT 24.255 3.362 24.28 3.512 ;
      RECT 24.245 3.358 24.255 3.507 ;
      RECT 24.225 3.353 24.245 3.502 ;
      RECT 24.19 3.348 24.225 3.495 ;
      RECT 24.13 3.343 24.19 3.488 ;
      RECT 24.117 3.339 24.13 3.486 ;
      RECT 24.031 3.334 24.117 3.483 ;
      RECT 23.945 3.324 24.031 3.479 ;
      RECT 23.904 3.317 23.945 3.476 ;
      RECT 23.818 3.31 23.904 3.473 ;
      RECT 23.732 3.3 23.818 3.469 ;
      RECT 23.646 3.29 23.732 3.464 ;
      RECT 23.56 3.28 23.646 3.46 ;
      RECT 23.55 3.265 23.56 3.458 ;
      RECT 23.54 3.25 23.55 3.458 ;
      RECT 23.475 3.245 23.54 3.457 ;
      RECT 23.31 3.242 23.355 3.45 ;
      RECT 24.555 4.147 24.56 4.338 ;
      RECT 24.55 4.142 24.555 4.345 ;
      RECT 24.536 4.14 24.55 4.351 ;
      RECT 24.45 4.14 24.536 4.353 ;
      RECT 24.446 4.14 24.45 4.356 ;
      RECT 24.36 4.14 24.446 4.374 ;
      RECT 24.35 4.145 24.36 4.393 ;
      RECT 24.34 4.2 24.35 4.397 ;
      RECT 24.315 4.215 24.34 4.404 ;
      RECT 24.275 4.235 24.315 4.417 ;
      RECT 24.27 4.247 24.275 4.427 ;
      RECT 24.255 4.253 24.27 4.432 ;
      RECT 24.25 4.258 24.255 4.436 ;
      RECT 24.23 4.265 24.25 4.441 ;
      RECT 24.16 4.29 24.23 4.458 ;
      RECT 24.12 4.318 24.16 4.478 ;
      RECT 24.115 4.328 24.12 4.486 ;
      RECT 24.095 4.335 24.115 4.488 ;
      RECT 24.09 4.342 24.095 4.491 ;
      RECT 24.06 4.35 24.09 4.494 ;
      RECT 24.055 4.355 24.06 4.498 ;
      RECT 23.981 4.359 24.055 4.506 ;
      RECT 23.895 4.368 23.981 4.522 ;
      RECT 23.891 4.373 23.895 4.531 ;
      RECT 23.805 4.378 23.891 4.541 ;
      RECT 23.765 4.386 23.805 4.553 ;
      RECT 23.715 4.392 23.765 4.56 ;
      RECT 23.63 4.401 23.715 4.575 ;
      RECT 23.555 4.412 23.63 4.593 ;
      RECT 23.52 4.419 23.555 4.603 ;
      RECT 23.445 4.427 23.52 4.608 ;
      RECT 23.39 4.436 23.445 4.608 ;
      RECT 23.365 4.441 23.39 4.606 ;
      RECT 23.355 4.444 23.365 4.604 ;
      RECT 23.32 4.446 23.355 4.602 ;
      RECT 23.29 4.448 23.32 4.598 ;
      RECT 23.245 4.447 23.29 4.594 ;
      RECT 23.225 4.442 23.245 4.591 ;
      RECT 23.175 4.427 23.225 4.588 ;
      RECT 23.165 4.412 23.175 4.583 ;
      RECT 23.115 4.397 23.165 4.573 ;
      RECT 23.065 4.372 23.115 4.553 ;
      RECT 23.055 4.357 23.065 4.535 ;
      RECT 23.05 4.355 23.055 4.529 ;
      RECT 23.03 4.35 23.05 4.524 ;
      RECT 23.025 4.342 23.03 4.518 ;
      RECT 23.01 4.336 23.025 4.511 ;
      RECT 23.005 4.331 23.01 4.503 ;
      RECT 22.985 4.326 23.005 4.495 ;
      RECT 22.97 4.319 22.985 4.488 ;
      RECT 22.955 4.313 22.97 4.479 ;
      RECT 22.95 4.307 22.955 4.472 ;
      RECT 22.905 4.282 22.95 4.458 ;
      RECT 22.89 4.252 22.905 4.44 ;
      RECT 22.875 4.235 22.89 4.431 ;
      RECT 22.85 4.215 22.875 4.419 ;
      RECT 22.81 4.185 22.85 4.399 ;
      RECT 22.8 4.155 22.81 4.384 ;
      RECT 22.785 4.145 22.8 4.377 ;
      RECT 22.73 4.11 22.785 4.356 ;
      RECT 22.715 4.073 22.73 4.335 ;
      RECT 22.705 4.06 22.715 4.327 ;
      RECT 22.655 4.03 22.705 4.309 ;
      RECT 22.64 3.96 22.655 4.29 ;
      RECT 22.595 3.96 22.64 4.273 ;
      RECT 22.57 3.96 22.595 4.255 ;
      RECT 22.56 3.96 22.57 4.248 ;
      RECT 22.481 3.96 22.56 4.241 ;
      RECT 22.395 3.96 22.481 4.233 ;
      RECT 22.38 3.992 22.395 4.228 ;
      RECT 22.305 4.002 22.38 4.224 ;
      RECT 22.285 4.012 22.305 4.219 ;
      RECT 22.26 4.012 22.285 4.216 ;
      RECT 22.25 4.002 22.26 4.215 ;
      RECT 22.24 3.975 22.25 4.214 ;
      RECT 22.2 3.97 22.24 4.212 ;
      RECT 22.155 3.97 22.2 4.208 ;
      RECT 22.13 3.97 22.155 4.203 ;
      RECT 22.08 3.97 22.13 4.19 ;
      RECT 22.04 3.975 22.05 4.175 ;
      RECT 22.05 3.97 22.08 4.18 ;
      RECT 24.035 3.75 24.295 4.01 ;
      RECT 24.03 3.772 24.295 3.968 ;
      RECT 23.27 3.6 23.49 3.965 ;
      RECT 23.252 3.687 23.49 3.964 ;
      RECT 23.235 3.692 23.49 3.961 ;
      RECT 23.235 3.692 23.51 3.96 ;
      RECT 23.205 3.702 23.51 3.958 ;
      RECT 23.2 3.717 23.51 3.954 ;
      RECT 23.2 3.717 23.515 3.953 ;
      RECT 23.195 3.775 23.515 3.951 ;
      RECT 23.195 3.775 23.525 3.948 ;
      RECT 23.19 3.84 23.525 3.943 ;
      RECT 23.27 3.6 23.53 3.86 ;
      RECT 22.015 3.43 22.275 3.69 ;
      RECT 22.015 3.473 22.361 3.664 ;
      RECT 22.015 3.473 22.405 3.663 ;
      RECT 22.015 3.473 22.425 3.661 ;
      RECT 22.015 3.473 22.525 3.66 ;
      RECT 22.015 3.473 22.545 3.658 ;
      RECT 22.015 3.473 22.555 3.653 ;
      RECT 22.425 3.44 22.615 3.65 ;
      RECT 22.425 3.442 22.62 3.648 ;
      RECT 22.415 3.447 22.625 3.64 ;
      RECT 22.361 3.471 22.625 3.64 ;
      RECT 22.405 3.465 22.415 3.662 ;
      RECT 22.415 3.445 22.62 3.648 ;
      RECT 21.37 4.505 21.575 4.735 ;
      RECT 21.31 4.455 21.365 4.715 ;
      RECT 21.37 4.455 21.57 4.735 ;
      RECT 22.34 4.77 22.345 4.797 ;
      RECT 22.33 4.68 22.34 4.802 ;
      RECT 22.325 4.602 22.33 4.808 ;
      RECT 22.315 4.592 22.325 4.815 ;
      RECT 22.31 4.582 22.315 4.821 ;
      RECT 22.3 4.577 22.31 4.823 ;
      RECT 22.285 4.569 22.3 4.831 ;
      RECT 22.27 4.56 22.285 4.843 ;
      RECT 22.26 4.552 22.27 4.853 ;
      RECT 22.225 4.47 22.26 4.871 ;
      RECT 22.19 4.47 22.225 4.89 ;
      RECT 22.175 4.47 22.19 4.898 ;
      RECT 22.12 4.47 22.175 4.898 ;
      RECT 22.086 4.47 22.12 4.889 ;
      RECT 22 4.47 22.086 4.865 ;
      RECT 21.99 4.53 22 4.847 ;
      RECT 21.95 4.532 21.99 4.838 ;
      RECT 21.945 4.534 21.95 4.828 ;
      RECT 21.925 4.536 21.945 4.823 ;
      RECT 21.915 4.539 21.925 4.818 ;
      RECT 21.905 4.54 21.915 4.813 ;
      RECT 21.881 4.541 21.905 4.805 ;
      RECT 21.795 4.546 21.881 4.783 ;
      RECT 21.74 4.545 21.795 4.756 ;
      RECT 21.725 4.538 21.74 4.743 ;
      RECT 21.69 4.533 21.725 4.739 ;
      RECT 21.635 4.525 21.69 4.738 ;
      RECT 21.575 4.512 21.635 4.736 ;
      RECT 21.365 4.455 21.37 4.723 ;
      RECT 21.44 3.825 21.625 4.035 ;
      RECT 21.43 3.83 21.64 4.028 ;
      RECT 21.47 3.735 21.73 3.995 ;
      RECT 21.425 3.892 21.73 3.918 ;
      RECT 20.77 3.685 20.775 4.485 ;
      RECT 20.715 3.735 20.745 4.485 ;
      RECT 20.705 3.735 20.71 4.045 ;
      RECT 20.69 3.735 20.695 4.04 ;
      RECT 20.235 3.78 20.25 3.995 ;
      RECT 20.165 3.78 20.25 3.99 ;
      RECT 21.43 3.36 21.5 3.57 ;
      RECT 21.5 3.367 21.51 3.565 ;
      RECT 21.396 3.36 21.43 3.577 ;
      RECT 21.31 3.36 21.396 3.601 ;
      RECT 21.3 3.365 21.31 3.62 ;
      RECT 21.295 3.377 21.3 3.623 ;
      RECT 21.28 3.392 21.295 3.627 ;
      RECT 21.275 3.41 21.28 3.631 ;
      RECT 21.235 3.42 21.275 3.64 ;
      RECT 21.22 3.427 21.235 3.652 ;
      RECT 21.205 3.432 21.22 3.657 ;
      RECT 21.19 3.435 21.205 3.662 ;
      RECT 21.18 3.437 21.19 3.666 ;
      RECT 21.145 3.444 21.18 3.674 ;
      RECT 21.11 3.452 21.145 3.688 ;
      RECT 21.1 3.458 21.11 3.697 ;
      RECT 21.095 3.46 21.1 3.699 ;
      RECT 21.075 3.463 21.095 3.705 ;
      RECT 21.045 3.47 21.075 3.716 ;
      RECT 21.035 3.476 21.045 3.723 ;
      RECT 21.01 3.479 21.035 3.73 ;
      RECT 21 3.483 21.01 3.738 ;
      RECT 20.995 3.484 21 3.76 ;
      RECT 20.99 3.485 20.995 3.775 ;
      RECT 20.985 3.486 20.99 3.79 ;
      RECT 20.98 3.487 20.985 3.805 ;
      RECT 20.975 3.488 20.98 3.835 ;
      RECT 20.965 3.49 20.975 3.868 ;
      RECT 20.95 3.494 20.965 3.915 ;
      RECT 20.94 3.497 20.95 3.96 ;
      RECT 20.935 3.5 20.94 3.988 ;
      RECT 20.925 3.502 20.935 4.015 ;
      RECT 20.92 3.505 20.925 4.05 ;
      RECT 20.89 3.51 20.92 4.108 ;
      RECT 20.885 3.515 20.89 4.193 ;
      RECT 20.88 3.517 20.885 4.228 ;
      RECT 20.875 3.519 20.88 4.31 ;
      RECT 20.87 3.521 20.875 4.398 ;
      RECT 20.86 3.523 20.87 4.48 ;
      RECT 20.845 3.537 20.86 4.485 ;
      RECT 20.81 3.582 20.845 4.485 ;
      RECT 20.8 3.622 20.81 4.485 ;
      RECT 20.785 3.65 20.8 4.485 ;
      RECT 20.78 3.667 20.785 4.485 ;
      RECT 20.775 3.675 20.78 4.485 ;
      RECT 20.765 3.69 20.77 4.485 ;
      RECT 20.76 3.697 20.765 4.485 ;
      RECT 20.75 3.717 20.76 4.485 ;
      RECT 20.745 3.73 20.75 4.485 ;
      RECT 20.71 3.735 20.715 4.07 ;
      RECT 20.695 4.125 20.715 4.485 ;
      RECT 20.695 3.735 20.705 4.043 ;
      RECT 20.69 4.165 20.695 4.485 ;
      RECT 20.64 3.735 20.69 4.038 ;
      RECT 20.685 4.202 20.69 4.485 ;
      RECT 20.675 4.225 20.685 4.485 ;
      RECT 20.67 4.27 20.675 4.485 ;
      RECT 20.66 4.28 20.67 4.478 ;
      RECT 20.586 3.735 20.64 4.032 ;
      RECT 20.5 3.735 20.586 4.025 ;
      RECT 20.451 3.782 20.5 4.018 ;
      RECT 20.365 3.79 20.451 4.011 ;
      RECT 20.35 3.787 20.365 4.006 ;
      RECT 20.336 3.78 20.35 4.005 ;
      RECT 20.25 3.78 20.336 4 ;
      RECT 20.155 3.785 20.165 3.985 ;
      RECT 19.745 3.215 19.76 3.615 ;
      RECT 19.94 3.215 19.945 3.475 ;
      RECT 19.685 3.215 19.73 3.475 ;
      RECT 20.14 4.52 20.145 4.725 ;
      RECT 20.135 4.51 20.14 4.73 ;
      RECT 20.13 4.497 20.135 4.735 ;
      RECT 20.125 4.477 20.13 4.735 ;
      RECT 20.1 4.43 20.125 4.735 ;
      RECT 20.065 4.345 20.1 4.735 ;
      RECT 20.06 4.282 20.065 4.735 ;
      RECT 20.055 4.267 20.06 4.735 ;
      RECT 20.04 4.227 20.055 4.735 ;
      RECT 20.035 4.202 20.04 4.735 ;
      RECT 20.025 4.185 20.035 4.735 ;
      RECT 19.99 4.107 20.025 4.735 ;
      RECT 19.985 4.05 19.99 4.735 ;
      RECT 19.98 4.037 19.985 4.735 ;
      RECT 19.97 4.015 19.98 4.735 ;
      RECT 19.96 3.98 19.97 4.735 ;
      RECT 19.95 3.95 19.96 4.735 ;
      RECT 19.94 3.865 19.95 4.378 ;
      RECT 19.947 4.51 19.95 4.735 ;
      RECT 19.945 4.52 19.947 4.735 ;
      RECT 19.935 4.53 19.945 4.73 ;
      RECT 19.93 3.215 19.94 3.61 ;
      RECT 19.935 3.742 19.94 4.353 ;
      RECT 19.93 3.64 19.935 4.336 ;
      RECT 19.92 3.215 19.93 4.312 ;
      RECT 19.915 3.215 19.92 4.283 ;
      RECT 19.91 3.215 19.915 4.273 ;
      RECT 19.89 3.215 19.91 4.235 ;
      RECT 19.885 3.215 19.89 4.193 ;
      RECT 19.88 3.215 19.885 4.173 ;
      RECT 19.85 3.215 19.88 4.123 ;
      RECT 19.84 3.215 19.85 4.07 ;
      RECT 19.835 3.215 19.84 4.043 ;
      RECT 19.83 3.215 19.835 4.028 ;
      RECT 19.82 3.215 19.83 4.005 ;
      RECT 19.81 3.215 19.82 3.98 ;
      RECT 19.805 3.215 19.81 3.92 ;
      RECT 19.795 3.215 19.805 3.858 ;
      RECT 19.79 3.215 19.795 3.778 ;
      RECT 19.785 3.215 19.79 3.743 ;
      RECT 19.78 3.215 19.785 3.718 ;
      RECT 19.775 3.215 19.78 3.703 ;
      RECT 19.77 3.215 19.775 3.673 ;
      RECT 19.765 3.215 19.77 3.65 ;
      RECT 19.76 3.215 19.765 3.623 ;
      RECT 19.73 3.215 19.745 3.61 ;
      RECT 18.885 4.75 19.07 4.96 ;
      RECT 18.875 4.755 19.085 4.953 ;
      RECT 18.875 4.755 19.105 4.925 ;
      RECT 18.875 4.755 19.12 4.904 ;
      RECT 18.875 4.755 19.135 4.902 ;
      RECT 18.875 4.755 19.145 4.901 ;
      RECT 18.875 4.755 19.175 4.898 ;
      RECT 19.525 4.6 19.785 4.86 ;
      RECT 19.485 4.647 19.785 4.843 ;
      RECT 19.476 4.655 19.485 4.846 ;
      RECT 19.07 4.748 19.785 4.843 ;
      RECT 19.39 4.673 19.476 4.853 ;
      RECT 19.085 4.745 19.785 4.843 ;
      RECT 19.331 4.695 19.39 4.865 ;
      RECT 19.105 4.741 19.785 4.843 ;
      RECT 19.245 4.707 19.331 4.876 ;
      RECT 19.12 4.737 19.785 4.843 ;
      RECT 19.19 4.72 19.245 4.888 ;
      RECT 19.135 4.735 19.785 4.843 ;
      RECT 19.175 4.726 19.19 4.894 ;
      RECT 19.145 4.731 19.785 4.843 ;
      RECT 19.29 4.255 19.55 4.515 ;
      RECT 19.29 4.275 19.66 4.485 ;
      RECT 19.29 4.28 19.67 4.48 ;
      RECT 19.481 3.694 19.56 3.925 ;
      RECT 19.395 3.697 19.61 3.92 ;
      RECT 19.39 3.697 19.61 3.915 ;
      RECT 19.39 3.702 19.62 3.913 ;
      RECT 19.365 3.702 19.62 3.91 ;
      RECT 19.365 3.71 19.63 3.908 ;
      RECT 19.245 3.645 19.505 3.905 ;
      RECT 19.245 3.692 19.555 3.905 ;
      RECT 18.5 4.265 18.505 4.525 ;
      RECT 18.33 4.035 18.335 4.525 ;
      RECT 18.215 4.275 18.22 4.5 ;
      RECT 18.925 3.37 18.93 3.58 ;
      RECT 18.93 3.375 18.945 3.575 ;
      RECT 18.865 3.37 18.925 3.588 ;
      RECT 18.85 3.37 18.865 3.598 ;
      RECT 18.8 3.37 18.85 3.615 ;
      RECT 18.78 3.37 18.8 3.638 ;
      RECT 18.765 3.37 18.78 3.65 ;
      RECT 18.745 3.37 18.765 3.66 ;
      RECT 18.735 3.375 18.745 3.669 ;
      RECT 18.73 3.385 18.735 3.674 ;
      RECT 18.725 3.397 18.73 3.678 ;
      RECT 18.715 3.42 18.725 3.683 ;
      RECT 18.71 3.435 18.715 3.687 ;
      RECT 18.705 3.452 18.71 3.69 ;
      RECT 18.7 3.46 18.705 3.693 ;
      RECT 18.69 3.465 18.7 3.697 ;
      RECT 18.685 3.472 18.69 3.702 ;
      RECT 18.675 3.477 18.685 3.706 ;
      RECT 18.65 3.489 18.675 3.717 ;
      RECT 18.63 3.506 18.65 3.733 ;
      RECT 18.605 3.523 18.63 3.755 ;
      RECT 18.57 3.546 18.605 3.813 ;
      RECT 18.55 3.568 18.57 3.875 ;
      RECT 18.545 3.578 18.55 3.91 ;
      RECT 18.535 3.585 18.545 3.948 ;
      RECT 18.53 3.592 18.535 3.968 ;
      RECT 18.525 3.603 18.53 4.005 ;
      RECT 18.52 3.611 18.525 4.07 ;
      RECT 18.51 3.622 18.52 4.123 ;
      RECT 18.505 3.64 18.51 4.193 ;
      RECT 18.5 3.65 18.505 4.23 ;
      RECT 18.495 3.66 18.5 4.525 ;
      RECT 18.49 3.672 18.495 4.525 ;
      RECT 18.485 3.682 18.49 4.525 ;
      RECT 18.475 3.692 18.485 4.525 ;
      RECT 18.465 3.715 18.475 4.525 ;
      RECT 18.45 3.75 18.465 4.525 ;
      RECT 18.41 3.812 18.45 4.525 ;
      RECT 18.405 3.865 18.41 4.525 ;
      RECT 18.38 3.9 18.405 4.525 ;
      RECT 18.365 3.945 18.38 4.525 ;
      RECT 18.36 3.967 18.365 4.525 ;
      RECT 18.35 3.98 18.36 4.525 ;
      RECT 18.34 4.005 18.35 4.525 ;
      RECT 18.335 4.027 18.34 4.525 ;
      RECT 18.31 4.065 18.33 4.525 ;
      RECT 18.27 4.122 18.31 4.525 ;
      RECT 18.265 4.172 18.27 4.525 ;
      RECT 18.26 4.19 18.265 4.525 ;
      RECT 18.255 4.202 18.26 4.525 ;
      RECT 18.245 4.22 18.255 4.525 ;
      RECT 18.235 4.24 18.245 4.5 ;
      RECT 18.23 4.257 18.235 4.5 ;
      RECT 18.22 4.27 18.23 4.5 ;
      RECT 18.19 4.28 18.215 4.5 ;
      RECT 18.18 4.287 18.19 4.5 ;
      RECT 18.165 4.297 18.18 4.495 ;
      RECT 16.605 10.055 16.895 10.285 ;
      RECT 16.665 9.31 16.835 10.285 ;
      RECT 16.515 9.31 16.865 9.6 ;
      RECT 16.515 9.315 16.895 9.545 ;
      RECT 16.14 8.57 16.49 8.86 ;
      RECT 16.14 8.575 16.525 8.805 ;
      RECT 16.06 8.605 16.525 8.775 ;
      RECT 96.14 7.215 96.51 7.585 ;
      RECT 91.055 4.145 91.425 4.515 ;
      RECT 80.355 7.215 80.725 7.585 ;
      RECT 75.27 4.145 75.64 4.515 ;
      RECT 64.57 7.215 64.94 7.585 ;
      RECT 59.485 4.145 59.855 4.515 ;
      RECT 48.795 7.215 49.165 7.585 ;
      RECT 43.71 4.145 44.08 4.515 ;
      RECT 33.015 7.215 33.385 7.585 ;
      RECT 27.93 4.145 28.3 4.515 ;
    LAYER mcon ;
      RECT 96.23 7.305 96.4 7.475 ;
      RECT 96.225 8.605 96.395 8.775 ;
      RECT 96.225 10.085 96.395 10.255 ;
      RECT 95.855 8.235 96.025 8.405 ;
      RECT 95.85 4.055 96.02 4.225 ;
      RECT 95.235 2.205 95.405 2.375 ;
      RECT 95.235 3.685 95.405 3.855 ;
      RECT 95.235 8.605 95.405 8.775 ;
      RECT 95.235 10.085 95.405 10.255 ;
      RECT 94.865 4.055 95.035 4.225 ;
      RECT 94.865 8.235 95.035 8.405 ;
      RECT 93.875 3.315 94.045 3.485 ;
      RECT 93.875 8.975 94.045 9.145 ;
      RECT 93.445 2.205 93.615 2.375 ;
      RECT 93.445 2.945 93.615 3.115 ;
      RECT 93.445 9.345 93.615 9.515 ;
      RECT 93.445 10.085 93.615 10.255 ;
      RECT 93.075 3.685 93.245 3.855 ;
      RECT 93.075 8.605 93.245 8.775 ;
      RECT 89.83 3.34 90 3.51 ;
      RECT 89.685 3.78 89.855 3.95 ;
      RECT 89.095 8.975 89.265 9.145 ;
      RECT 89.075 3.82 89.245 3.99 ;
      RECT 88.73 3.455 88.9 3.625 ;
      RECT 88.72 4.815 88.89 4.985 ;
      RECT 88.665 9.345 88.835 9.515 ;
      RECT 88.665 10.085 88.835 10.255 ;
      RECT 87.955 3.53 88.125 3.7 ;
      RECT 87.775 4.845 87.945 5.015 ;
      RECT 87.495 4.16 87.665 4.33 ;
      RECT 87.175 3.785 87.345 3.955 ;
      RECT 86.485 3.265 86.655 3.435 ;
      RECT 86.41 3.735 86.58 3.905 ;
      RECT 85.56 3.46 85.73 3.63 ;
      RECT 85.22 4.655 85.39 4.825 ;
      RECT 85.185 3.99 85.355 4.16 ;
      RECT 84.575 3.845 84.745 4.015 ;
      RECT 84.505 4.545 84.675 4.715 ;
      RECT 84.445 3.38 84.615 3.55 ;
      RECT 83.805 4.295 83.975 4.465 ;
      RECT 83.3 3.8 83.47 3.97 ;
      RECT 83.08 4.545 83.25 4.715 ;
      RECT 82.875 3.425 83.045 3.595 ;
      RECT 82.605 4.295 82.775 4.465 ;
      RECT 82.565 3.725 82.735 3.895 ;
      RECT 82.02 4.77 82.19 4.94 ;
      RECT 81.88 3.39 82.05 3.56 ;
      RECT 81.31 4.31 81.48 4.48 ;
      RECT 80.445 7.305 80.615 7.475 ;
      RECT 80.44 8.605 80.61 8.775 ;
      RECT 80.44 10.085 80.61 10.255 ;
      RECT 80.07 8.235 80.24 8.405 ;
      RECT 80.065 4.055 80.235 4.225 ;
      RECT 79.45 2.205 79.62 2.375 ;
      RECT 79.45 3.685 79.62 3.855 ;
      RECT 79.45 8.605 79.62 8.775 ;
      RECT 79.45 10.085 79.62 10.255 ;
      RECT 79.08 4.055 79.25 4.225 ;
      RECT 79.08 8.235 79.25 8.405 ;
      RECT 78.09 3.315 78.26 3.485 ;
      RECT 78.09 8.975 78.26 9.145 ;
      RECT 77.66 2.205 77.83 2.375 ;
      RECT 77.66 2.945 77.83 3.115 ;
      RECT 77.66 9.345 77.83 9.515 ;
      RECT 77.66 10.085 77.83 10.255 ;
      RECT 77.29 3.685 77.46 3.855 ;
      RECT 77.29 8.605 77.46 8.775 ;
      RECT 74.045 3.34 74.215 3.51 ;
      RECT 73.9 3.78 74.07 3.95 ;
      RECT 73.31 8.975 73.48 9.145 ;
      RECT 73.29 3.82 73.46 3.99 ;
      RECT 72.945 3.455 73.115 3.625 ;
      RECT 72.935 4.815 73.105 4.985 ;
      RECT 72.88 9.345 73.05 9.515 ;
      RECT 72.88 10.085 73.05 10.255 ;
      RECT 72.17 3.53 72.34 3.7 ;
      RECT 71.99 4.845 72.16 5.015 ;
      RECT 71.71 4.16 71.88 4.33 ;
      RECT 71.39 3.785 71.56 3.955 ;
      RECT 70.7 3.265 70.87 3.435 ;
      RECT 70.625 3.735 70.795 3.905 ;
      RECT 69.775 3.46 69.945 3.63 ;
      RECT 69.435 4.655 69.605 4.825 ;
      RECT 69.4 3.99 69.57 4.16 ;
      RECT 68.79 3.845 68.96 4.015 ;
      RECT 68.72 4.545 68.89 4.715 ;
      RECT 68.66 3.38 68.83 3.55 ;
      RECT 68.02 4.295 68.19 4.465 ;
      RECT 67.515 3.8 67.685 3.97 ;
      RECT 67.295 4.545 67.465 4.715 ;
      RECT 67.09 3.425 67.26 3.595 ;
      RECT 66.82 4.295 66.99 4.465 ;
      RECT 66.78 3.725 66.95 3.895 ;
      RECT 66.235 4.77 66.405 4.94 ;
      RECT 66.095 3.39 66.265 3.56 ;
      RECT 65.525 4.31 65.695 4.48 ;
      RECT 64.66 7.305 64.83 7.475 ;
      RECT 64.655 8.605 64.825 8.775 ;
      RECT 64.655 10.085 64.825 10.255 ;
      RECT 64.285 8.235 64.455 8.405 ;
      RECT 64.28 4.055 64.45 4.225 ;
      RECT 63.665 2.205 63.835 2.375 ;
      RECT 63.665 3.685 63.835 3.855 ;
      RECT 63.665 8.605 63.835 8.775 ;
      RECT 63.665 10.085 63.835 10.255 ;
      RECT 63.295 4.055 63.465 4.225 ;
      RECT 63.295 8.235 63.465 8.405 ;
      RECT 62.305 3.315 62.475 3.485 ;
      RECT 62.305 8.975 62.475 9.145 ;
      RECT 61.875 2.205 62.045 2.375 ;
      RECT 61.875 2.945 62.045 3.115 ;
      RECT 61.875 9.345 62.045 9.515 ;
      RECT 61.875 10.085 62.045 10.255 ;
      RECT 61.505 3.685 61.675 3.855 ;
      RECT 61.505 8.605 61.675 8.775 ;
      RECT 58.26 3.34 58.43 3.51 ;
      RECT 58.115 3.78 58.285 3.95 ;
      RECT 57.525 8.975 57.695 9.145 ;
      RECT 57.505 3.82 57.675 3.99 ;
      RECT 57.16 3.455 57.33 3.625 ;
      RECT 57.15 4.815 57.32 4.985 ;
      RECT 57.095 9.345 57.265 9.515 ;
      RECT 57.095 10.085 57.265 10.255 ;
      RECT 56.385 3.53 56.555 3.7 ;
      RECT 56.205 4.845 56.375 5.015 ;
      RECT 55.925 4.16 56.095 4.33 ;
      RECT 55.605 3.785 55.775 3.955 ;
      RECT 54.915 3.265 55.085 3.435 ;
      RECT 54.84 3.735 55.01 3.905 ;
      RECT 53.99 3.46 54.16 3.63 ;
      RECT 53.65 4.655 53.82 4.825 ;
      RECT 53.615 3.99 53.785 4.16 ;
      RECT 53.005 3.845 53.175 4.015 ;
      RECT 52.935 4.545 53.105 4.715 ;
      RECT 52.875 3.38 53.045 3.55 ;
      RECT 52.235 4.295 52.405 4.465 ;
      RECT 51.73 3.8 51.9 3.97 ;
      RECT 51.51 4.545 51.68 4.715 ;
      RECT 51.305 3.425 51.475 3.595 ;
      RECT 51.035 4.295 51.205 4.465 ;
      RECT 50.995 3.725 51.165 3.895 ;
      RECT 50.45 4.77 50.62 4.94 ;
      RECT 50.31 3.39 50.48 3.56 ;
      RECT 49.74 4.31 49.91 4.48 ;
      RECT 48.885 7.305 49.055 7.475 ;
      RECT 48.88 8.605 49.05 8.775 ;
      RECT 48.88 10.085 49.05 10.255 ;
      RECT 48.51 8.235 48.68 8.405 ;
      RECT 48.505 4.055 48.675 4.225 ;
      RECT 47.89 2.205 48.06 2.375 ;
      RECT 47.89 3.685 48.06 3.855 ;
      RECT 47.89 8.605 48.06 8.775 ;
      RECT 47.89 10.085 48.06 10.255 ;
      RECT 47.52 4.055 47.69 4.225 ;
      RECT 47.52 8.235 47.69 8.405 ;
      RECT 46.53 3.315 46.7 3.485 ;
      RECT 46.53 8.975 46.7 9.145 ;
      RECT 46.1 2.205 46.27 2.375 ;
      RECT 46.1 2.945 46.27 3.115 ;
      RECT 46.1 9.345 46.27 9.515 ;
      RECT 46.1 10.085 46.27 10.255 ;
      RECT 45.73 3.685 45.9 3.855 ;
      RECT 45.73 8.605 45.9 8.775 ;
      RECT 42.485 3.34 42.655 3.51 ;
      RECT 42.34 3.78 42.51 3.95 ;
      RECT 41.75 8.975 41.92 9.145 ;
      RECT 41.73 3.82 41.9 3.99 ;
      RECT 41.385 3.455 41.555 3.625 ;
      RECT 41.375 4.815 41.545 4.985 ;
      RECT 41.32 9.345 41.49 9.515 ;
      RECT 41.32 10.085 41.49 10.255 ;
      RECT 40.61 3.53 40.78 3.7 ;
      RECT 40.43 4.845 40.6 5.015 ;
      RECT 40.15 4.16 40.32 4.33 ;
      RECT 39.83 3.785 40 3.955 ;
      RECT 39.14 3.265 39.31 3.435 ;
      RECT 39.065 3.735 39.235 3.905 ;
      RECT 38.215 3.46 38.385 3.63 ;
      RECT 37.875 4.655 38.045 4.825 ;
      RECT 37.84 3.99 38.01 4.16 ;
      RECT 37.23 3.845 37.4 4.015 ;
      RECT 37.16 4.545 37.33 4.715 ;
      RECT 37.1 3.38 37.27 3.55 ;
      RECT 36.46 4.295 36.63 4.465 ;
      RECT 35.955 3.8 36.125 3.97 ;
      RECT 35.735 4.545 35.905 4.715 ;
      RECT 35.53 3.425 35.7 3.595 ;
      RECT 35.26 4.295 35.43 4.465 ;
      RECT 35.22 3.725 35.39 3.895 ;
      RECT 34.675 4.77 34.845 4.94 ;
      RECT 34.535 3.39 34.705 3.56 ;
      RECT 33.965 4.31 34.135 4.48 ;
      RECT 33.105 7.305 33.275 7.475 ;
      RECT 33.1 8.605 33.27 8.775 ;
      RECT 33.1 10.085 33.27 10.255 ;
      RECT 32.73 8.235 32.9 8.405 ;
      RECT 32.725 4.055 32.895 4.225 ;
      RECT 32.11 2.205 32.28 2.375 ;
      RECT 32.11 3.685 32.28 3.855 ;
      RECT 32.11 8.605 32.28 8.775 ;
      RECT 32.11 10.085 32.28 10.255 ;
      RECT 31.74 4.055 31.91 4.225 ;
      RECT 31.74 8.235 31.91 8.405 ;
      RECT 30.75 3.315 30.92 3.485 ;
      RECT 30.75 8.975 30.92 9.145 ;
      RECT 30.32 2.205 30.49 2.375 ;
      RECT 30.32 2.945 30.49 3.115 ;
      RECT 30.32 9.345 30.49 9.515 ;
      RECT 30.32 10.085 30.49 10.255 ;
      RECT 29.95 3.685 30.12 3.855 ;
      RECT 29.95 8.605 30.12 8.775 ;
      RECT 26.705 3.34 26.875 3.51 ;
      RECT 26.56 3.78 26.73 3.95 ;
      RECT 25.97 8.975 26.14 9.145 ;
      RECT 25.95 3.82 26.12 3.99 ;
      RECT 25.605 3.455 25.775 3.625 ;
      RECT 25.595 4.815 25.765 4.985 ;
      RECT 25.54 9.345 25.71 9.515 ;
      RECT 25.54 10.085 25.71 10.255 ;
      RECT 24.83 3.53 25 3.7 ;
      RECT 24.65 4.845 24.82 5.015 ;
      RECT 24.37 4.16 24.54 4.33 ;
      RECT 24.05 3.785 24.22 3.955 ;
      RECT 23.36 3.265 23.53 3.435 ;
      RECT 23.285 3.735 23.455 3.905 ;
      RECT 22.435 3.46 22.605 3.63 ;
      RECT 22.095 4.655 22.265 4.825 ;
      RECT 22.06 3.99 22.23 4.16 ;
      RECT 21.45 3.845 21.62 4.015 ;
      RECT 21.38 4.545 21.55 4.715 ;
      RECT 21.32 3.38 21.49 3.55 ;
      RECT 20.68 4.295 20.85 4.465 ;
      RECT 20.175 3.8 20.345 3.97 ;
      RECT 19.955 4.545 20.125 4.715 ;
      RECT 19.75 3.425 19.92 3.595 ;
      RECT 19.48 4.295 19.65 4.465 ;
      RECT 19.44 3.725 19.61 3.895 ;
      RECT 18.895 4.77 19.065 4.94 ;
      RECT 18.755 3.39 18.925 3.56 ;
      RECT 18.185 4.31 18.355 4.48 ;
      RECT 16.665 9.345 16.835 9.515 ;
      RECT 16.665 10.085 16.835 10.255 ;
      RECT 16.295 8.605 16.465 8.775 ;
    LAYER li1 ;
      RECT 96.225 7.305 96.395 8.775 ;
      RECT 96.225 7.305 96.4 8.565 ;
      RECT 95.855 9.255 96.325 9.425 ;
      RECT 95.855 8.235 96.025 9.425 ;
      RECT 95.85 3.035 96.02 4.225 ;
      RECT 95.85 3.035 96.32 3.205 ;
      RECT 95.235 3.895 95.41 5.155 ;
      RECT 95.235 3.685 95.405 5.155 ;
      RECT 95.235 7.305 95.405 8.775 ;
      RECT 95.235 7.305 95.41 8.565 ;
      RECT 94.865 3.035 95.035 4.225 ;
      RECT 94.865 3.035 95.335 3.205 ;
      RECT 94.865 9.255 95.335 9.425 ;
      RECT 94.865 8.235 95.035 9.425 ;
      RECT 93.875 4.015 94.05 5.155 ;
      RECT 93.875 1.865 94.045 5.155 ;
      RECT 93.875 1.865 94.05 2.415 ;
      RECT 93.875 10.045 94.05 10.595 ;
      RECT 93.875 7.305 94.045 10.595 ;
      RECT 93.875 7.305 94.05 8.445 ;
      RECT 93.445 3.895 93.62 5.155 ;
      RECT 93.445 2.945 93.615 5.155 ;
      RECT 93.445 7.305 93.615 9.515 ;
      RECT 93.445 7.305 93.62 8.565 ;
      RECT 93.015 3.925 93.185 5.155 ;
      RECT 93.075 2.145 93.245 4.095 ;
      RECT 93.015 1.865 93.185 2.315 ;
      RECT 93.015 10.145 93.185 10.595 ;
      RECT 93.075 8.365 93.245 10.315 ;
      RECT 93.015 7.305 93.185 8.535 ;
      RECT 92.49 3.895 92.665 5.155 ;
      RECT 92.49 1.865 92.66 5.155 ;
      RECT 92.49 3.365 92.9 3.695 ;
      RECT 92.49 2.525 92.9 2.855 ;
      RECT 92.49 1.865 92.665 2.355 ;
      RECT 92.49 10.105 92.665 10.595 ;
      RECT 92.49 7.305 92.66 10.595 ;
      RECT 92.49 9.605 92.9 9.935 ;
      RECT 92.49 8.765 92.9 9.095 ;
      RECT 92.49 7.305 92.665 8.565 ;
      RECT 89.83 3.27 90.56 3.51 ;
      RECT 90.372 3.065 90.56 3.51 ;
      RECT 90.2 3.077 90.575 3.504 ;
      RECT 90.115 3.092 90.595 3.489 ;
      RECT 90.115 3.107 90.6 3.479 ;
      RECT 90.07 3.127 90.615 3.471 ;
      RECT 90.047 3.162 90.63 3.425 ;
      RECT 89.961 3.185 90.635 3.385 ;
      RECT 89.961 3.203 90.645 3.355 ;
      RECT 89.83 3.272 90.65 3.318 ;
      RECT 89.875 3.215 90.645 3.355 ;
      RECT 89.961 3.167 90.63 3.425 ;
      RECT 90.047 3.136 90.615 3.471 ;
      RECT 90.07 3.117 90.6 3.479 ;
      RECT 90.115 3.09 90.575 3.504 ;
      RECT 90.2 3.072 90.56 3.51 ;
      RECT 90.286 3.066 90.56 3.51 ;
      RECT 90.372 3.061 90.505 3.51 ;
      RECT 90.458 3.056 90.505 3.51 ;
      RECT 90.02 4.67 90.025 4.683 ;
      RECT 90.015 4.565 90.02 4.688 ;
      RECT 89.99 4.425 90.015 4.703 ;
      RECT 89.955 4.376 89.99 4.735 ;
      RECT 89.95 4.344 89.955 4.755 ;
      RECT 89.945 4.335 89.95 4.755 ;
      RECT 89.865 4.3 89.945 4.755 ;
      RECT 89.802 4.27 89.865 4.755 ;
      RECT 89.716 4.258 89.802 4.755 ;
      RECT 89.63 4.244 89.716 4.755 ;
      RECT 89.55 4.231 89.63 4.741 ;
      RECT 89.515 4.223 89.55 4.721 ;
      RECT 89.505 4.22 89.515 4.712 ;
      RECT 89.475 4.215 89.505 4.699 ;
      RECT 89.425 4.19 89.475 4.675 ;
      RECT 89.411 4.164 89.425 4.657 ;
      RECT 89.325 4.124 89.411 4.633 ;
      RECT 89.28 4.072 89.325 4.602 ;
      RECT 89.27 4.047 89.28 4.589 ;
      RECT 89.265 3.828 89.27 3.85 ;
      RECT 89.26 4.03 89.27 4.585 ;
      RECT 89.26 3.826 89.265 3.94 ;
      RECT 89.25 3.822 89.26 4.581 ;
      RECT 89.206 3.82 89.25 4.569 ;
      RECT 89.12 3.82 89.206 4.54 ;
      RECT 89.09 3.82 89.12 4.513 ;
      RECT 89.075 3.82 89.09 4.501 ;
      RECT 89.035 3.832 89.075 4.486 ;
      RECT 89.015 3.851 89.035 4.465 ;
      RECT 89.005 3.861 89.015 4.449 ;
      RECT 88.995 3.867 89.005 4.438 ;
      RECT 88.975 3.877 88.995 4.421 ;
      RECT 88.97 3.886 88.975 4.408 ;
      RECT 88.965 3.89 88.97 4.358 ;
      RECT 88.955 3.896 88.965 4.275 ;
      RECT 88.95 3.9 88.955 4.189 ;
      RECT 88.945 3.92 88.95 4.126 ;
      RECT 88.94 3.943 88.945 4.073 ;
      RECT 88.935 3.961 88.94 4.018 ;
      RECT 89.545 3.78 89.715 4.04 ;
      RECT 89.715 3.745 89.76 4.026 ;
      RECT 89.676 3.747 89.765 4.009 ;
      RECT 89.565 3.764 89.851 3.98 ;
      RECT 89.565 3.779 89.855 3.952 ;
      RECT 89.565 3.76 89.765 4.009 ;
      RECT 89.59 3.748 89.715 4.04 ;
      RECT 89.676 3.746 89.76 4.026 ;
      RECT 89.095 10.045 89.27 10.595 ;
      RECT 89.095 7.305 89.265 10.595 ;
      RECT 89.095 7.305 89.27 8.445 ;
      RECT 88.73 3.135 88.9 3.625 ;
      RECT 88.73 3.135 88.935 3.605 ;
      RECT 88.865 3.055 88.975 3.565 ;
      RECT 88.846 3.059 88.995 3.535 ;
      RECT 88.76 3.067 89.015 3.518 ;
      RECT 88.76 3.073 89.02 3.508 ;
      RECT 88.76 3.082 89.04 3.496 ;
      RECT 88.735 3.107 89.07 3.474 ;
      RECT 88.735 3.127 89.075 3.454 ;
      RECT 88.73 3.14 89.085 3.434 ;
      RECT 88.73 3.207 89.09 3.415 ;
      RECT 88.73 3.34 89.095 3.402 ;
      RECT 88.725 3.145 89.085 3.235 ;
      RECT 88.735 3.102 89.04 3.496 ;
      RECT 88.846 3.057 88.975 3.565 ;
      RECT 88.72 4.81 89.02 5.065 ;
      RECT 88.805 4.776 89.02 5.065 ;
      RECT 88.805 4.779 89.025 4.925 ;
      RECT 88.74 4.8 89.025 4.925 ;
      RECT 88.775 4.79 89.02 5.065 ;
      RECT 88.77 4.795 89.025 4.925 ;
      RECT 88.805 4.774 89.006 5.065 ;
      RECT 88.891 4.765 89.006 5.065 ;
      RECT 88.891 4.759 88.92 5.065 ;
      RECT 88.665 7.305 88.835 9.515 ;
      RECT 88.665 7.305 88.84 8.565 ;
      RECT 88.38 4.4 88.39 4.89 ;
      RECT 88.04 4.335 88.05 4.635 ;
      RECT 88.555 4.507 88.56 4.726 ;
      RECT 88.545 4.487 88.555 4.743 ;
      RECT 88.535 4.467 88.545 4.773 ;
      RECT 88.53 4.457 88.535 4.788 ;
      RECT 88.525 4.453 88.53 4.793 ;
      RECT 88.51 4.445 88.525 4.8 ;
      RECT 88.47 4.425 88.51 4.825 ;
      RECT 88.445 4.407 88.47 4.858 ;
      RECT 88.44 4.405 88.445 4.871 ;
      RECT 88.42 4.402 88.44 4.875 ;
      RECT 88.39 4.4 88.42 4.885 ;
      RECT 88.32 4.402 88.38 4.886 ;
      RECT 88.3 4.402 88.32 4.88 ;
      RECT 88.275 4.4 88.3 4.877 ;
      RECT 88.24 4.395 88.275 4.873 ;
      RECT 88.22 4.389 88.24 4.86 ;
      RECT 88.21 4.386 88.22 4.848 ;
      RECT 88.19 4.383 88.21 4.833 ;
      RECT 88.17 4.379 88.19 4.815 ;
      RECT 88.165 4.376 88.17 4.805 ;
      RECT 88.16 4.375 88.165 4.803 ;
      RECT 88.15 4.372 88.16 4.795 ;
      RECT 88.14 4.366 88.15 4.778 ;
      RECT 88.13 4.36 88.14 4.76 ;
      RECT 88.12 4.354 88.13 4.748 ;
      RECT 88.11 4.348 88.12 4.728 ;
      RECT 88.105 4.344 88.11 4.713 ;
      RECT 88.1 4.342 88.105 4.705 ;
      RECT 88.095 4.34 88.1 4.698 ;
      RECT 88.09 4.338 88.095 4.688 ;
      RECT 88.085 4.336 88.09 4.682 ;
      RECT 88.075 4.335 88.085 4.672 ;
      RECT 88.065 4.335 88.075 4.663 ;
      RECT 88.05 4.335 88.065 4.648 ;
      RECT 88.01 4.335 88.04 4.632 ;
      RECT 87.99 4.337 88.01 4.627 ;
      RECT 87.985 4.342 87.99 4.625 ;
      RECT 87.955 4.35 87.985 4.623 ;
      RECT 87.925 4.365 87.955 4.622 ;
      RECT 87.88 4.387 87.925 4.627 ;
      RECT 87.875 4.402 87.88 4.631 ;
      RECT 87.86 4.407 87.875 4.633 ;
      RECT 87.855 4.411 87.86 4.635 ;
      RECT 87.795 4.434 87.855 4.644 ;
      RECT 87.775 4.46 87.795 4.657 ;
      RECT 87.765 4.467 87.775 4.661 ;
      RECT 87.75 4.474 87.765 4.664 ;
      RECT 87.73 4.484 87.75 4.667 ;
      RECT 87.725 4.492 87.73 4.67 ;
      RECT 87.68 4.497 87.725 4.677 ;
      RECT 87.67 4.5 87.68 4.684 ;
      RECT 87.66 4.5 87.67 4.688 ;
      RECT 87.625 4.502 87.66 4.7 ;
      RECT 87.605 4.505 87.625 4.713 ;
      RECT 87.565 4.508 87.605 4.724 ;
      RECT 87.55 4.51 87.565 4.737 ;
      RECT 87.54 4.51 87.55 4.742 ;
      RECT 87.515 4.511 87.54 4.75 ;
      RECT 87.505 4.513 87.515 4.755 ;
      RECT 87.5 4.514 87.505 4.758 ;
      RECT 87.475 4.512 87.5 4.761 ;
      RECT 87.46 4.51 87.475 4.762 ;
      RECT 87.44 4.507 87.46 4.764 ;
      RECT 87.42 4.502 87.44 4.764 ;
      RECT 87.36 4.497 87.42 4.761 ;
      RECT 87.325 4.472 87.36 4.757 ;
      RECT 87.315 4.449 87.325 4.755 ;
      RECT 87.285 4.426 87.315 4.755 ;
      RECT 87.275 4.405 87.285 4.755 ;
      RECT 87.25 4.387 87.275 4.753 ;
      RECT 87.235 4.365 87.25 4.75 ;
      RECT 87.22 4.347 87.235 4.748 ;
      RECT 87.2 4.337 87.22 4.746 ;
      RECT 87.185 4.332 87.2 4.745 ;
      RECT 87.17 4.33 87.185 4.744 ;
      RECT 87.14 4.331 87.17 4.742 ;
      RECT 87.12 4.334 87.14 4.74 ;
      RECT 87.063 4.338 87.12 4.74 ;
      RECT 86.977 4.347 87.063 4.74 ;
      RECT 86.891 4.358 86.977 4.74 ;
      RECT 86.805 4.369 86.891 4.74 ;
      RECT 86.785 4.376 86.805 4.748 ;
      RECT 86.775 4.379 86.785 4.755 ;
      RECT 86.71 4.384 86.775 4.773 ;
      RECT 86.68 4.391 86.71 4.798 ;
      RECT 86.67 4.394 86.68 4.805 ;
      RECT 86.625 4.398 86.67 4.81 ;
      RECT 86.595 4.403 86.625 4.815 ;
      RECT 86.594 4.405 86.595 4.815 ;
      RECT 86.508 4.411 86.594 4.815 ;
      RECT 86.422 4.422 86.508 4.815 ;
      RECT 86.336 4.434 86.422 4.815 ;
      RECT 86.25 4.445 86.336 4.815 ;
      RECT 86.235 4.452 86.25 4.81 ;
      RECT 86.23 4.454 86.235 4.804 ;
      RECT 86.21 4.465 86.23 4.799 ;
      RECT 86.2 4.483 86.21 4.793 ;
      RECT 86.195 4.495 86.2 4.593 ;
      RECT 88.49 3.248 88.51 3.335 ;
      RECT 88.485 3.183 88.49 3.367 ;
      RECT 88.475 3.15 88.485 3.372 ;
      RECT 88.47 3.13 88.475 3.378 ;
      RECT 88.44 3.13 88.47 3.395 ;
      RECT 88.391 3.13 88.44 3.431 ;
      RECT 88.305 3.13 88.391 3.489 ;
      RECT 88.276 3.14 88.305 3.538 ;
      RECT 88.19 3.182 88.276 3.591 ;
      RECT 88.17 3.22 88.19 3.638 ;
      RECT 88.145 3.237 88.17 3.658 ;
      RECT 88.135 3.251 88.145 3.678 ;
      RECT 88.13 3.257 88.135 3.688 ;
      RECT 88.125 3.261 88.13 3.695 ;
      RECT 88.075 3.281 88.125 3.7 ;
      RECT 88.01 3.325 88.075 3.7 ;
      RECT 87.985 3.375 88.01 3.7 ;
      RECT 87.975 3.405 87.985 3.7 ;
      RECT 87.97 3.432 87.975 3.7 ;
      RECT 87.965 3.45 87.97 3.7 ;
      RECT 87.955 3.492 87.965 3.7 ;
      RECT 87.71 10.105 87.885 10.595 ;
      RECT 87.71 7.305 87.88 10.595 ;
      RECT 87.71 9.605 88.12 9.935 ;
      RECT 87.71 8.765 88.12 9.095 ;
      RECT 87.71 7.305 87.885 8.565 ;
      RECT 87.785 4.85 87.975 5.075 ;
      RECT 87.775 4.851 87.98 5.07 ;
      RECT 87.775 4.853 87.99 5.05 ;
      RECT 87.775 4.857 87.995 5.035 ;
      RECT 87.775 4.844 87.945 5.07 ;
      RECT 87.775 4.847 87.97 5.07 ;
      RECT 87.785 4.843 87.945 5.075 ;
      RECT 87.871 4.841 87.945 5.075 ;
      RECT 87.495 4.092 87.665 4.33 ;
      RECT 87.495 4.092 87.751 4.244 ;
      RECT 87.495 4.092 87.755 4.154 ;
      RECT 87.545 3.865 87.765 4.133 ;
      RECT 87.54 3.882 87.77 4.106 ;
      RECT 87.505 4.04 87.77 4.106 ;
      RECT 87.525 3.89 87.665 4.33 ;
      RECT 87.515 3.972 87.775 4.089 ;
      RECT 87.51 4.02 87.775 4.089 ;
      RECT 87.515 3.93 87.77 4.106 ;
      RECT 87.54 3.867 87.765 4.133 ;
      RECT 87.105 3.842 87.275 4.04 ;
      RECT 87.105 3.842 87.32 4.015 ;
      RECT 87.175 3.785 87.345 3.973 ;
      RECT 87.15 3.8 87.345 3.973 ;
      RECT 86.765 3.846 86.795 4.04 ;
      RECT 86.76 3.818 86.765 4.04 ;
      RECT 86.73 3.792 86.76 4.042 ;
      RECT 86.705 3.75 86.73 4.045 ;
      RECT 86.695 3.722 86.705 4.047 ;
      RECT 86.66 3.702 86.695 4.049 ;
      RECT 86.595 3.687 86.66 4.055 ;
      RECT 86.545 3.685 86.595 4.061 ;
      RECT 86.522 3.687 86.545 4.066 ;
      RECT 86.436 3.698 86.522 4.072 ;
      RECT 86.35 3.716 86.436 4.082 ;
      RECT 86.335 3.727 86.35 4.088 ;
      RECT 86.265 3.75 86.335 4.094 ;
      RECT 86.21 3.782 86.265 4.102 ;
      RECT 86.17 3.805 86.21 4.108 ;
      RECT 86.156 3.818 86.17 4.111 ;
      RECT 86.07 3.84 86.156 4.117 ;
      RECT 86.055 3.865 86.07 4.123 ;
      RECT 86.015 3.88 86.055 4.127 ;
      RECT 85.965 3.895 86.015 4.132 ;
      RECT 85.94 3.902 85.965 4.136 ;
      RECT 85.88 3.897 85.94 4.14 ;
      RECT 85.865 3.888 85.88 4.144 ;
      RECT 85.795 3.878 85.865 4.14 ;
      RECT 85.77 3.87 85.79 4.13 ;
      RECT 85.711 3.87 85.77 4.108 ;
      RECT 85.625 3.87 85.711 4.065 ;
      RECT 85.79 3.87 85.795 4.135 ;
      RECT 86.485 3.101 86.655 3.435 ;
      RECT 86.455 3.101 86.655 3.43 ;
      RECT 86.395 3.068 86.455 3.418 ;
      RECT 86.395 3.124 86.665 3.413 ;
      RECT 86.37 3.124 86.665 3.407 ;
      RECT 86.365 3.065 86.395 3.404 ;
      RECT 86.35 3.071 86.485 3.402 ;
      RECT 86.345 3.079 86.57 3.39 ;
      RECT 86.345 3.131 86.68 3.343 ;
      RECT 86.33 3.087 86.57 3.338 ;
      RECT 86.33 3.157 86.69 3.279 ;
      RECT 86.3 3.107 86.655 3.24 ;
      RECT 86.3 3.197 86.7 3.236 ;
      RECT 86.35 3.076 86.57 3.402 ;
      RECT 85.69 3.406 85.745 3.67 ;
      RECT 85.69 3.406 85.81 3.669 ;
      RECT 85.69 3.406 85.835 3.668 ;
      RECT 85.69 3.406 85.9 3.667 ;
      RECT 85.835 3.372 85.915 3.666 ;
      RECT 85.65 3.416 86.06 3.665 ;
      RECT 85.69 3.413 86.06 3.665 ;
      RECT 85.65 3.421 86.065 3.658 ;
      RECT 85.635 3.423 86.065 3.657 ;
      RECT 85.635 3.43 86.07 3.653 ;
      RECT 85.615 3.429 86.065 3.649 ;
      RECT 85.615 3.437 86.075 3.648 ;
      RECT 85.61 3.434 86.07 3.644 ;
      RECT 85.61 3.447 86.085 3.643 ;
      RECT 85.595 3.437 86.075 3.642 ;
      RECT 85.56 3.45 86.085 3.635 ;
      RECT 85.745 3.405 86.055 3.665 ;
      RECT 85.745 3.39 86.005 3.665 ;
      RECT 85.81 3.377 85.94 3.665 ;
      RECT 85.355 4.466 85.37 4.859 ;
      RECT 85.32 4.471 85.37 4.858 ;
      RECT 85.355 4.47 85.415 4.857 ;
      RECT 85.3 4.481 85.415 4.856 ;
      RECT 85.315 4.477 85.415 4.856 ;
      RECT 85.28 4.487 85.49 4.853 ;
      RECT 85.28 4.506 85.535 4.851 ;
      RECT 85.28 4.513 85.54 4.848 ;
      RECT 85.265 4.49 85.49 4.845 ;
      RECT 85.245 4.495 85.49 4.838 ;
      RECT 85.24 4.499 85.49 4.834 ;
      RECT 85.24 4.516 85.55 4.833 ;
      RECT 85.22 4.51 85.535 4.829 ;
      RECT 85.22 4.519 85.555 4.823 ;
      RECT 85.215 4.525 85.555 4.595 ;
      RECT 85.28 4.485 85.415 4.853 ;
      RECT 85.155 3.848 85.355 4.16 ;
      RECT 85.23 3.826 85.355 4.16 ;
      RECT 85.17 3.845 85.36 4.145 ;
      RECT 85.14 3.856 85.36 4.143 ;
      RECT 85.155 3.851 85.365 4.109 ;
      RECT 85.14 3.955 85.37 4.076 ;
      RECT 85.17 3.827 85.355 4.16 ;
      RECT 85.23 3.805 85.33 4.16 ;
      RECT 85.255 3.802 85.33 4.16 ;
      RECT 85.255 3.797 85.275 4.16 ;
      RECT 84.66 3.865 84.835 4.04 ;
      RECT 84.655 3.865 84.835 4.038 ;
      RECT 84.63 3.865 84.835 4.033 ;
      RECT 84.575 3.845 84.745 4.023 ;
      RECT 84.575 3.852 84.81 4.023 ;
      RECT 84.66 4.532 84.675 4.715 ;
      RECT 84.65 4.51 84.66 4.715 ;
      RECT 84.635 4.49 84.65 4.715 ;
      RECT 84.625 4.465 84.635 4.715 ;
      RECT 84.595 4.43 84.625 4.715 ;
      RECT 84.56 4.37 84.595 4.715 ;
      RECT 84.555 4.332 84.56 4.715 ;
      RECT 84.505 4.283 84.555 4.715 ;
      RECT 84.495 4.233 84.505 4.703 ;
      RECT 84.48 4.212 84.495 4.663 ;
      RECT 84.46 4.18 84.48 4.613 ;
      RECT 84.435 4.136 84.46 4.553 ;
      RECT 84.43 4.108 84.435 4.508 ;
      RECT 84.425 4.099 84.43 4.494 ;
      RECT 84.42 4.092 84.425 4.481 ;
      RECT 84.415 4.087 84.42 4.47 ;
      RECT 84.41 4.072 84.415 4.46 ;
      RECT 84.405 4.05 84.41 4.447 ;
      RECT 84.395 4.01 84.405 4.422 ;
      RECT 84.37 3.94 84.395 4.378 ;
      RECT 84.365 3.88 84.37 4.343 ;
      RECT 84.35 3.86 84.365 4.31 ;
      RECT 84.345 3.86 84.35 4.285 ;
      RECT 84.315 3.86 84.345 4.24 ;
      RECT 84.27 3.86 84.315 4.18 ;
      RECT 84.195 3.86 84.27 4.128 ;
      RECT 84.19 3.86 84.195 4.093 ;
      RECT 84.185 3.86 84.19 4.083 ;
      RECT 84.18 3.86 84.185 4.063 ;
      RECT 84.445 3.08 84.615 3.55 ;
      RECT 84.39 3.073 84.585 3.534 ;
      RECT 84.39 3.087 84.62 3.533 ;
      RECT 84.375 3.088 84.62 3.514 ;
      RECT 84.37 3.106 84.62 3.5 ;
      RECT 84.375 3.089 84.625 3.498 ;
      RECT 84.36 3.12 84.625 3.483 ;
      RECT 84.375 3.095 84.63 3.468 ;
      RECT 84.355 3.135 84.63 3.465 ;
      RECT 84.37 3.107 84.635 3.45 ;
      RECT 84.37 3.119 84.64 3.43 ;
      RECT 84.355 3.135 84.645 3.413 ;
      RECT 84.355 3.145 84.65 3.268 ;
      RECT 84.35 3.145 84.65 3.225 ;
      RECT 84.35 3.16 84.655 3.203 ;
      RECT 84.445 3.07 84.585 3.55 ;
      RECT 84.445 3.068 84.555 3.55 ;
      RECT 84.531 3.065 84.555 3.55 ;
      RECT 84.19 4.732 84.195 4.778 ;
      RECT 84.18 4.58 84.19 4.802 ;
      RECT 84.175 4.425 84.18 4.827 ;
      RECT 84.16 4.387 84.175 4.838 ;
      RECT 84.155 4.37 84.16 4.845 ;
      RECT 84.145 4.358 84.155 4.852 ;
      RECT 84.14 4.349 84.145 4.854 ;
      RECT 84.135 4.347 84.14 4.858 ;
      RECT 84.09 4.338 84.135 4.873 ;
      RECT 84.085 4.33 84.09 4.887 ;
      RECT 84.08 4.327 84.085 4.891 ;
      RECT 84.065 4.322 84.08 4.899 ;
      RECT 84.01 4.312 84.065 4.91 ;
      RECT 83.975 4.3 84.01 4.911 ;
      RECT 83.966 4.295 83.975 4.905 ;
      RECT 83.88 4.295 83.966 4.895 ;
      RECT 83.85 4.295 83.88 4.873 ;
      RECT 83.84 4.295 83.845 4.853 ;
      RECT 83.835 4.295 83.84 4.815 ;
      RECT 83.83 4.295 83.835 4.773 ;
      RECT 83.825 4.295 83.83 4.733 ;
      RECT 83.82 4.295 83.825 4.663 ;
      RECT 83.81 4.295 83.82 4.585 ;
      RECT 83.805 4.295 83.81 4.485 ;
      RECT 83.845 4.295 83.85 4.855 ;
      RECT 83.34 4.377 83.43 4.855 ;
      RECT 83.325 4.38 83.445 4.853 ;
      RECT 83.34 4.379 83.445 4.853 ;
      RECT 83.305 4.386 83.47 4.843 ;
      RECT 83.325 4.38 83.47 4.843 ;
      RECT 83.29 4.392 83.47 4.831 ;
      RECT 83.325 4.383 83.52 4.824 ;
      RECT 83.276 4.4 83.52 4.822 ;
      RECT 83.305 4.39 83.53 4.81 ;
      RECT 83.276 4.411 83.56 4.801 ;
      RECT 83.19 4.435 83.56 4.795 ;
      RECT 83.19 4.448 83.6 4.778 ;
      RECT 83.185 4.47 83.6 4.771 ;
      RECT 83.155 4.485 83.6 4.761 ;
      RECT 83.15 4.496 83.6 4.751 ;
      RECT 83.12 4.509 83.6 4.742 ;
      RECT 83.105 4.527 83.6 4.731 ;
      RECT 83.08 4.54 83.6 4.721 ;
      RECT 83.34 4.376 83.35 4.855 ;
      RECT 83.386 3.8 83.425 4.045 ;
      RECT 83.3 3.8 83.435 4.043 ;
      RECT 83.185 3.825 83.435 4.04 ;
      RECT 83.185 3.825 83.44 4.038 ;
      RECT 83.185 3.825 83.455 4.033 ;
      RECT 83.291 3.8 83.47 4.013 ;
      RECT 83.205 3.808 83.47 4.013 ;
      RECT 82.875 3.16 83.045 3.595 ;
      RECT 82.865 3.194 83.045 3.578 ;
      RECT 82.945 3.13 83.115 3.565 ;
      RECT 82.85 3.205 83.115 3.543 ;
      RECT 82.945 3.14 83.12 3.533 ;
      RECT 82.875 3.192 83.15 3.518 ;
      RECT 82.835 3.218 83.15 3.503 ;
      RECT 82.835 3.26 83.16 3.483 ;
      RECT 82.83 3.285 83.165 3.465 ;
      RECT 82.83 3.295 83.17 3.45 ;
      RECT 82.825 3.232 83.15 3.448 ;
      RECT 82.825 3.305 83.175 3.433 ;
      RECT 82.82 3.242 83.15 3.43 ;
      RECT 82.815 3.326 83.18 3.413 ;
      RECT 82.815 3.358 83.185 3.393 ;
      RECT 82.81 3.272 83.16 3.385 ;
      RECT 82.815 3.257 83.15 3.413 ;
      RECT 82.83 3.227 83.15 3.465 ;
      RECT 82.675 3.814 82.9 4.07 ;
      RECT 82.675 3.847 82.92 4.06 ;
      RECT 82.64 3.847 82.92 4.058 ;
      RECT 82.64 3.86 82.925 4.048 ;
      RECT 82.64 3.88 82.935 4.04 ;
      RECT 82.64 3.977 82.94 4.033 ;
      RECT 82.62 3.725 82.75 4.023 ;
      RECT 82.575 3.88 82.935 3.965 ;
      RECT 82.565 3.725 82.75 3.91 ;
      RECT 82.565 3.757 82.836 3.91 ;
      RECT 82.53 4.287 82.55 4.465 ;
      RECT 82.495 4.24 82.53 4.465 ;
      RECT 82.48 4.18 82.495 4.465 ;
      RECT 82.455 4.127 82.48 4.465 ;
      RECT 82.44 4.08 82.455 4.465 ;
      RECT 82.42 4.057 82.44 4.465 ;
      RECT 82.395 4.022 82.42 4.465 ;
      RECT 82.385 3.868 82.395 4.465 ;
      RECT 82.355 3.863 82.385 4.456 ;
      RECT 82.35 3.86 82.355 4.446 ;
      RECT 82.335 3.86 82.35 4.42 ;
      RECT 82.33 3.86 82.335 4.383 ;
      RECT 82.305 3.86 82.33 4.335 ;
      RECT 82.285 3.86 82.305 4.26 ;
      RECT 82.275 3.86 82.285 4.22 ;
      RECT 82.27 3.86 82.275 4.195 ;
      RECT 82.265 3.86 82.27 4.178 ;
      RECT 82.26 3.86 82.265 4.16 ;
      RECT 82.255 3.861 82.26 4.15 ;
      RECT 82.245 3.863 82.255 4.118 ;
      RECT 82.235 3.865 82.245 4.085 ;
      RECT 82.225 3.868 82.235 4.058 ;
      RECT 82.55 4.295 82.775 4.465 ;
      RECT 81.88 3.107 82.05 3.56 ;
      RECT 81.88 3.107 82.14 3.526 ;
      RECT 81.88 3.107 82.17 3.51 ;
      RECT 81.88 3.107 82.2 3.483 ;
      RECT 82.136 3.085 82.215 3.465 ;
      RECT 81.915 3.092 82.22 3.45 ;
      RECT 81.915 3.1 82.23 3.413 ;
      RECT 81.875 3.127 82.23 3.385 ;
      RECT 81.86 3.14 82.23 3.35 ;
      RECT 81.88 3.115 82.25 3.34 ;
      RECT 81.855 3.18 82.25 3.31 ;
      RECT 81.855 3.21 82.255 3.293 ;
      RECT 81.85 3.24 82.255 3.28 ;
      RECT 81.915 3.089 82.215 3.465 ;
      RECT 82.05 3.086 82.136 3.544 ;
      RECT 82.001 3.087 82.215 3.465 ;
      RECT 82.145 4.747 82.19 4.94 ;
      RECT 82.135 4.717 82.145 4.94 ;
      RECT 82.13 4.702 82.135 4.94 ;
      RECT 82.09 4.612 82.13 4.94 ;
      RECT 82.085 4.525 82.09 4.94 ;
      RECT 82.075 4.495 82.085 4.94 ;
      RECT 82.07 4.455 82.075 4.94 ;
      RECT 82.06 4.417 82.07 4.94 ;
      RECT 82.055 4.382 82.06 4.94 ;
      RECT 82.035 4.335 82.055 4.94 ;
      RECT 82.02 4.26 82.035 4.94 ;
      RECT 82.015 4.215 82.02 4.935 ;
      RECT 82.01 4.195 82.015 4.908 ;
      RECT 82.005 4.175 82.01 4.893 ;
      RECT 82 4.15 82.005 4.873 ;
      RECT 81.995 4.128 82 4.858 ;
      RECT 81.99 4.106 81.995 4.84 ;
      RECT 81.985 4.085 81.99 4.83 ;
      RECT 81.975 4.057 81.985 4.8 ;
      RECT 81.965 4.02 81.975 4.768 ;
      RECT 81.955 3.98 81.965 4.735 ;
      RECT 81.945 3.958 81.955 4.705 ;
      RECT 81.915 3.91 81.945 4.637 ;
      RECT 81.9 3.87 81.915 4.564 ;
      RECT 81.89 3.87 81.9 4.53 ;
      RECT 81.885 3.87 81.89 4.505 ;
      RECT 81.88 3.87 81.885 4.49 ;
      RECT 81.875 3.87 81.88 4.468 ;
      RECT 81.87 3.87 81.875 4.455 ;
      RECT 81.855 3.87 81.87 4.42 ;
      RECT 81.835 3.87 81.855 4.36 ;
      RECT 81.825 3.87 81.835 4.31 ;
      RECT 81.805 3.87 81.825 4.258 ;
      RECT 81.785 3.87 81.805 4.215 ;
      RECT 81.775 3.87 81.785 4.203 ;
      RECT 81.745 3.87 81.775 4.19 ;
      RECT 81.715 3.891 81.745 4.17 ;
      RECT 81.705 3.919 81.715 4.15 ;
      RECT 81.69 3.936 81.705 4.118 ;
      RECT 81.685 3.95 81.69 4.085 ;
      RECT 81.68 3.958 81.685 4.058 ;
      RECT 81.675 3.966 81.68 4.02 ;
      RECT 81.68 4.49 81.685 4.825 ;
      RECT 81.645 4.477 81.68 4.824 ;
      RECT 81.575 4.417 81.645 4.823 ;
      RECT 81.495 4.36 81.575 4.822 ;
      RECT 81.36 4.32 81.495 4.821 ;
      RECT 81.36 4.507 81.695 4.81 ;
      RECT 81.32 4.507 81.695 4.8 ;
      RECT 81.32 4.525 81.7 4.795 ;
      RECT 81.32 4.615 81.705 4.785 ;
      RECT 81.315 4.31 81.48 4.765 ;
      RECT 81.31 4.31 81.48 4.508 ;
      RECT 81.31 4.467 81.675 4.508 ;
      RECT 81.31 4.455 81.67 4.508 ;
      RECT 80.44 7.305 80.61 8.775 ;
      RECT 80.44 7.305 80.615 8.565 ;
      RECT 80.07 9.255 80.54 9.425 ;
      RECT 80.07 8.235 80.24 9.425 ;
      RECT 80.065 3.035 80.235 4.225 ;
      RECT 80.065 3.035 80.535 3.205 ;
      RECT 79.45 3.895 79.625 5.155 ;
      RECT 79.45 3.685 79.62 5.155 ;
      RECT 79.45 7.305 79.62 8.775 ;
      RECT 79.45 7.305 79.625 8.565 ;
      RECT 79.08 3.035 79.25 4.225 ;
      RECT 79.08 3.035 79.55 3.205 ;
      RECT 79.08 9.255 79.55 9.425 ;
      RECT 79.08 8.235 79.25 9.425 ;
      RECT 78.09 4.015 78.265 5.155 ;
      RECT 78.09 1.865 78.26 5.155 ;
      RECT 78.09 1.865 78.265 2.415 ;
      RECT 78.09 10.045 78.265 10.595 ;
      RECT 78.09 7.305 78.26 10.595 ;
      RECT 78.09 7.305 78.265 8.445 ;
      RECT 77.66 3.895 77.835 5.155 ;
      RECT 77.66 2.945 77.83 5.155 ;
      RECT 77.66 7.305 77.83 9.515 ;
      RECT 77.66 7.305 77.835 8.565 ;
      RECT 77.23 3.925 77.4 5.155 ;
      RECT 77.29 2.145 77.46 4.095 ;
      RECT 77.23 1.865 77.4 2.315 ;
      RECT 77.23 10.145 77.4 10.595 ;
      RECT 77.29 8.365 77.46 10.315 ;
      RECT 77.23 7.305 77.4 8.535 ;
      RECT 76.705 3.895 76.88 5.155 ;
      RECT 76.705 1.865 76.875 5.155 ;
      RECT 76.705 3.365 77.115 3.695 ;
      RECT 76.705 2.525 77.115 2.855 ;
      RECT 76.705 1.865 76.88 2.355 ;
      RECT 76.705 10.105 76.88 10.595 ;
      RECT 76.705 7.305 76.875 10.595 ;
      RECT 76.705 9.605 77.115 9.935 ;
      RECT 76.705 8.765 77.115 9.095 ;
      RECT 76.705 7.305 76.88 8.565 ;
      RECT 74.045 3.27 74.775 3.51 ;
      RECT 74.587 3.065 74.775 3.51 ;
      RECT 74.415 3.077 74.79 3.504 ;
      RECT 74.33 3.092 74.81 3.489 ;
      RECT 74.33 3.107 74.815 3.479 ;
      RECT 74.285 3.127 74.83 3.471 ;
      RECT 74.262 3.162 74.845 3.425 ;
      RECT 74.176 3.185 74.85 3.385 ;
      RECT 74.176 3.203 74.86 3.355 ;
      RECT 74.045 3.272 74.865 3.318 ;
      RECT 74.09 3.215 74.86 3.355 ;
      RECT 74.176 3.167 74.845 3.425 ;
      RECT 74.262 3.136 74.83 3.471 ;
      RECT 74.285 3.117 74.815 3.479 ;
      RECT 74.33 3.09 74.79 3.504 ;
      RECT 74.415 3.072 74.775 3.51 ;
      RECT 74.501 3.066 74.775 3.51 ;
      RECT 74.587 3.061 74.72 3.51 ;
      RECT 74.673 3.056 74.72 3.51 ;
      RECT 74.235 4.67 74.24 4.683 ;
      RECT 74.23 4.565 74.235 4.688 ;
      RECT 74.205 4.425 74.23 4.703 ;
      RECT 74.17 4.376 74.205 4.735 ;
      RECT 74.165 4.344 74.17 4.755 ;
      RECT 74.16 4.335 74.165 4.755 ;
      RECT 74.08 4.3 74.16 4.755 ;
      RECT 74.017 4.27 74.08 4.755 ;
      RECT 73.931 4.258 74.017 4.755 ;
      RECT 73.845 4.244 73.931 4.755 ;
      RECT 73.765 4.231 73.845 4.741 ;
      RECT 73.73 4.223 73.765 4.721 ;
      RECT 73.72 4.22 73.73 4.712 ;
      RECT 73.69 4.215 73.72 4.699 ;
      RECT 73.64 4.19 73.69 4.675 ;
      RECT 73.626 4.164 73.64 4.657 ;
      RECT 73.54 4.124 73.626 4.633 ;
      RECT 73.495 4.072 73.54 4.602 ;
      RECT 73.485 4.047 73.495 4.589 ;
      RECT 73.48 3.828 73.485 3.85 ;
      RECT 73.475 4.03 73.485 4.585 ;
      RECT 73.475 3.826 73.48 3.94 ;
      RECT 73.465 3.822 73.475 4.581 ;
      RECT 73.421 3.82 73.465 4.569 ;
      RECT 73.335 3.82 73.421 4.54 ;
      RECT 73.305 3.82 73.335 4.513 ;
      RECT 73.29 3.82 73.305 4.501 ;
      RECT 73.25 3.832 73.29 4.486 ;
      RECT 73.23 3.851 73.25 4.465 ;
      RECT 73.22 3.861 73.23 4.449 ;
      RECT 73.21 3.867 73.22 4.438 ;
      RECT 73.19 3.877 73.21 4.421 ;
      RECT 73.185 3.886 73.19 4.408 ;
      RECT 73.18 3.89 73.185 4.358 ;
      RECT 73.17 3.896 73.18 4.275 ;
      RECT 73.165 3.9 73.17 4.189 ;
      RECT 73.16 3.92 73.165 4.126 ;
      RECT 73.155 3.943 73.16 4.073 ;
      RECT 73.15 3.961 73.155 4.018 ;
      RECT 73.76 3.78 73.93 4.04 ;
      RECT 73.93 3.745 73.975 4.026 ;
      RECT 73.891 3.747 73.98 4.009 ;
      RECT 73.78 3.764 74.066 3.98 ;
      RECT 73.78 3.779 74.07 3.952 ;
      RECT 73.78 3.76 73.98 4.009 ;
      RECT 73.805 3.748 73.93 4.04 ;
      RECT 73.891 3.746 73.975 4.026 ;
      RECT 73.31 10.045 73.485 10.595 ;
      RECT 73.31 7.305 73.48 10.595 ;
      RECT 73.31 7.305 73.485 8.445 ;
      RECT 72.945 3.135 73.115 3.625 ;
      RECT 72.945 3.135 73.15 3.605 ;
      RECT 73.08 3.055 73.19 3.565 ;
      RECT 73.061 3.059 73.21 3.535 ;
      RECT 72.975 3.067 73.23 3.518 ;
      RECT 72.975 3.073 73.235 3.508 ;
      RECT 72.975 3.082 73.255 3.496 ;
      RECT 72.95 3.107 73.285 3.474 ;
      RECT 72.95 3.127 73.29 3.454 ;
      RECT 72.945 3.14 73.3 3.434 ;
      RECT 72.945 3.207 73.305 3.415 ;
      RECT 72.945 3.34 73.31 3.402 ;
      RECT 72.94 3.145 73.3 3.235 ;
      RECT 72.95 3.102 73.255 3.496 ;
      RECT 73.061 3.057 73.19 3.565 ;
      RECT 72.935 4.81 73.235 5.065 ;
      RECT 73.02 4.776 73.235 5.065 ;
      RECT 73.02 4.779 73.24 4.925 ;
      RECT 72.955 4.8 73.24 4.925 ;
      RECT 72.99 4.79 73.235 5.065 ;
      RECT 72.985 4.795 73.24 4.925 ;
      RECT 73.02 4.774 73.221 5.065 ;
      RECT 73.106 4.765 73.221 5.065 ;
      RECT 73.106 4.759 73.135 5.065 ;
      RECT 72.88 7.305 73.05 9.515 ;
      RECT 72.88 7.305 73.055 8.565 ;
      RECT 72.595 4.4 72.605 4.89 ;
      RECT 72.255 4.335 72.265 4.635 ;
      RECT 72.77 4.507 72.775 4.726 ;
      RECT 72.76 4.487 72.77 4.743 ;
      RECT 72.75 4.467 72.76 4.773 ;
      RECT 72.745 4.457 72.75 4.788 ;
      RECT 72.74 4.453 72.745 4.793 ;
      RECT 72.725 4.445 72.74 4.8 ;
      RECT 72.685 4.425 72.725 4.825 ;
      RECT 72.66 4.407 72.685 4.858 ;
      RECT 72.655 4.405 72.66 4.871 ;
      RECT 72.635 4.402 72.655 4.875 ;
      RECT 72.605 4.4 72.635 4.885 ;
      RECT 72.535 4.402 72.595 4.886 ;
      RECT 72.515 4.402 72.535 4.88 ;
      RECT 72.49 4.4 72.515 4.877 ;
      RECT 72.455 4.395 72.49 4.873 ;
      RECT 72.435 4.389 72.455 4.86 ;
      RECT 72.425 4.386 72.435 4.848 ;
      RECT 72.405 4.383 72.425 4.833 ;
      RECT 72.385 4.379 72.405 4.815 ;
      RECT 72.38 4.376 72.385 4.805 ;
      RECT 72.375 4.375 72.38 4.803 ;
      RECT 72.365 4.372 72.375 4.795 ;
      RECT 72.355 4.366 72.365 4.778 ;
      RECT 72.345 4.36 72.355 4.76 ;
      RECT 72.335 4.354 72.345 4.748 ;
      RECT 72.325 4.348 72.335 4.728 ;
      RECT 72.32 4.344 72.325 4.713 ;
      RECT 72.315 4.342 72.32 4.705 ;
      RECT 72.31 4.34 72.315 4.698 ;
      RECT 72.305 4.338 72.31 4.688 ;
      RECT 72.3 4.336 72.305 4.682 ;
      RECT 72.29 4.335 72.3 4.672 ;
      RECT 72.28 4.335 72.29 4.663 ;
      RECT 72.265 4.335 72.28 4.648 ;
      RECT 72.225 4.335 72.255 4.632 ;
      RECT 72.205 4.337 72.225 4.627 ;
      RECT 72.2 4.342 72.205 4.625 ;
      RECT 72.17 4.35 72.2 4.623 ;
      RECT 72.14 4.365 72.17 4.622 ;
      RECT 72.095 4.387 72.14 4.627 ;
      RECT 72.09 4.402 72.095 4.631 ;
      RECT 72.075 4.407 72.09 4.633 ;
      RECT 72.07 4.411 72.075 4.635 ;
      RECT 72.01 4.434 72.07 4.644 ;
      RECT 71.99 4.46 72.01 4.657 ;
      RECT 71.98 4.467 71.99 4.661 ;
      RECT 71.965 4.474 71.98 4.664 ;
      RECT 71.945 4.484 71.965 4.667 ;
      RECT 71.94 4.492 71.945 4.67 ;
      RECT 71.895 4.497 71.94 4.677 ;
      RECT 71.885 4.5 71.895 4.684 ;
      RECT 71.875 4.5 71.885 4.688 ;
      RECT 71.84 4.502 71.875 4.7 ;
      RECT 71.82 4.505 71.84 4.713 ;
      RECT 71.78 4.508 71.82 4.724 ;
      RECT 71.765 4.51 71.78 4.737 ;
      RECT 71.755 4.51 71.765 4.742 ;
      RECT 71.73 4.511 71.755 4.75 ;
      RECT 71.72 4.513 71.73 4.755 ;
      RECT 71.715 4.514 71.72 4.758 ;
      RECT 71.69 4.512 71.715 4.761 ;
      RECT 71.675 4.51 71.69 4.762 ;
      RECT 71.655 4.507 71.675 4.764 ;
      RECT 71.635 4.502 71.655 4.764 ;
      RECT 71.575 4.497 71.635 4.761 ;
      RECT 71.54 4.472 71.575 4.757 ;
      RECT 71.53 4.449 71.54 4.755 ;
      RECT 71.5 4.426 71.53 4.755 ;
      RECT 71.49 4.405 71.5 4.755 ;
      RECT 71.465 4.387 71.49 4.753 ;
      RECT 71.45 4.365 71.465 4.75 ;
      RECT 71.435 4.347 71.45 4.748 ;
      RECT 71.415 4.337 71.435 4.746 ;
      RECT 71.4 4.332 71.415 4.745 ;
      RECT 71.385 4.33 71.4 4.744 ;
      RECT 71.355 4.331 71.385 4.742 ;
      RECT 71.335 4.334 71.355 4.74 ;
      RECT 71.278 4.338 71.335 4.74 ;
      RECT 71.192 4.347 71.278 4.74 ;
      RECT 71.106 4.358 71.192 4.74 ;
      RECT 71.02 4.369 71.106 4.74 ;
      RECT 71 4.376 71.02 4.748 ;
      RECT 70.99 4.379 71 4.755 ;
      RECT 70.925 4.384 70.99 4.773 ;
      RECT 70.895 4.391 70.925 4.798 ;
      RECT 70.885 4.394 70.895 4.805 ;
      RECT 70.84 4.398 70.885 4.81 ;
      RECT 70.81 4.403 70.84 4.815 ;
      RECT 70.809 4.405 70.81 4.815 ;
      RECT 70.723 4.411 70.809 4.815 ;
      RECT 70.637 4.422 70.723 4.815 ;
      RECT 70.551 4.434 70.637 4.815 ;
      RECT 70.465 4.445 70.551 4.815 ;
      RECT 70.45 4.452 70.465 4.81 ;
      RECT 70.445 4.454 70.45 4.804 ;
      RECT 70.425 4.465 70.445 4.799 ;
      RECT 70.415 4.483 70.425 4.793 ;
      RECT 70.41 4.495 70.415 4.593 ;
      RECT 72.705 3.248 72.725 3.335 ;
      RECT 72.7 3.183 72.705 3.367 ;
      RECT 72.69 3.15 72.7 3.372 ;
      RECT 72.685 3.13 72.69 3.378 ;
      RECT 72.655 3.13 72.685 3.395 ;
      RECT 72.606 3.13 72.655 3.431 ;
      RECT 72.52 3.13 72.606 3.489 ;
      RECT 72.491 3.14 72.52 3.538 ;
      RECT 72.405 3.182 72.491 3.591 ;
      RECT 72.385 3.22 72.405 3.638 ;
      RECT 72.36 3.237 72.385 3.658 ;
      RECT 72.35 3.251 72.36 3.678 ;
      RECT 72.345 3.257 72.35 3.688 ;
      RECT 72.34 3.261 72.345 3.695 ;
      RECT 72.29 3.281 72.34 3.7 ;
      RECT 72.225 3.325 72.29 3.7 ;
      RECT 72.2 3.375 72.225 3.7 ;
      RECT 72.19 3.405 72.2 3.7 ;
      RECT 72.185 3.432 72.19 3.7 ;
      RECT 72.18 3.45 72.185 3.7 ;
      RECT 72.17 3.492 72.18 3.7 ;
      RECT 71.925 10.105 72.1 10.595 ;
      RECT 71.925 7.305 72.095 10.595 ;
      RECT 71.925 9.605 72.335 9.935 ;
      RECT 71.925 8.765 72.335 9.095 ;
      RECT 71.925 7.305 72.1 8.565 ;
      RECT 72 4.85 72.19 5.075 ;
      RECT 71.99 4.851 72.195 5.07 ;
      RECT 71.99 4.853 72.205 5.05 ;
      RECT 71.99 4.857 72.21 5.035 ;
      RECT 71.99 4.844 72.16 5.07 ;
      RECT 71.99 4.847 72.185 5.07 ;
      RECT 72 4.843 72.16 5.075 ;
      RECT 72.086 4.841 72.16 5.075 ;
      RECT 71.71 4.092 71.88 4.33 ;
      RECT 71.71 4.092 71.966 4.244 ;
      RECT 71.71 4.092 71.97 4.154 ;
      RECT 71.76 3.865 71.98 4.133 ;
      RECT 71.755 3.882 71.985 4.106 ;
      RECT 71.72 4.04 71.985 4.106 ;
      RECT 71.74 3.89 71.88 4.33 ;
      RECT 71.73 3.972 71.99 4.089 ;
      RECT 71.725 4.02 71.99 4.089 ;
      RECT 71.73 3.93 71.985 4.106 ;
      RECT 71.755 3.867 71.98 4.133 ;
      RECT 71.32 3.842 71.49 4.04 ;
      RECT 71.32 3.842 71.535 4.015 ;
      RECT 71.39 3.785 71.56 3.973 ;
      RECT 71.365 3.8 71.56 3.973 ;
      RECT 70.98 3.846 71.01 4.04 ;
      RECT 70.975 3.818 70.98 4.04 ;
      RECT 70.945 3.792 70.975 4.042 ;
      RECT 70.92 3.75 70.945 4.045 ;
      RECT 70.91 3.722 70.92 4.047 ;
      RECT 70.875 3.702 70.91 4.049 ;
      RECT 70.81 3.687 70.875 4.055 ;
      RECT 70.76 3.685 70.81 4.061 ;
      RECT 70.737 3.687 70.76 4.066 ;
      RECT 70.651 3.698 70.737 4.072 ;
      RECT 70.565 3.716 70.651 4.082 ;
      RECT 70.55 3.727 70.565 4.088 ;
      RECT 70.48 3.75 70.55 4.094 ;
      RECT 70.425 3.782 70.48 4.102 ;
      RECT 70.385 3.805 70.425 4.108 ;
      RECT 70.371 3.818 70.385 4.111 ;
      RECT 70.285 3.84 70.371 4.117 ;
      RECT 70.27 3.865 70.285 4.123 ;
      RECT 70.23 3.88 70.27 4.127 ;
      RECT 70.18 3.895 70.23 4.132 ;
      RECT 70.155 3.902 70.18 4.136 ;
      RECT 70.095 3.897 70.155 4.14 ;
      RECT 70.08 3.888 70.095 4.144 ;
      RECT 70.01 3.878 70.08 4.14 ;
      RECT 69.985 3.87 70.005 4.13 ;
      RECT 69.926 3.87 69.985 4.108 ;
      RECT 69.84 3.87 69.926 4.065 ;
      RECT 70.005 3.87 70.01 4.135 ;
      RECT 70.7 3.101 70.87 3.435 ;
      RECT 70.67 3.101 70.87 3.43 ;
      RECT 70.61 3.068 70.67 3.418 ;
      RECT 70.61 3.124 70.88 3.413 ;
      RECT 70.585 3.124 70.88 3.407 ;
      RECT 70.58 3.065 70.61 3.404 ;
      RECT 70.565 3.071 70.7 3.402 ;
      RECT 70.56 3.079 70.785 3.39 ;
      RECT 70.56 3.131 70.895 3.343 ;
      RECT 70.545 3.087 70.785 3.338 ;
      RECT 70.545 3.157 70.905 3.279 ;
      RECT 70.515 3.107 70.87 3.24 ;
      RECT 70.515 3.197 70.915 3.236 ;
      RECT 70.565 3.076 70.785 3.402 ;
      RECT 69.905 3.406 69.96 3.67 ;
      RECT 69.905 3.406 70.025 3.669 ;
      RECT 69.905 3.406 70.05 3.668 ;
      RECT 69.905 3.406 70.115 3.667 ;
      RECT 70.05 3.372 70.13 3.666 ;
      RECT 69.865 3.416 70.275 3.665 ;
      RECT 69.905 3.413 70.275 3.665 ;
      RECT 69.865 3.421 70.28 3.658 ;
      RECT 69.85 3.423 70.28 3.657 ;
      RECT 69.85 3.43 70.285 3.653 ;
      RECT 69.83 3.429 70.28 3.649 ;
      RECT 69.83 3.437 70.29 3.648 ;
      RECT 69.825 3.434 70.285 3.644 ;
      RECT 69.825 3.447 70.3 3.643 ;
      RECT 69.81 3.437 70.29 3.642 ;
      RECT 69.775 3.45 70.3 3.635 ;
      RECT 69.96 3.405 70.27 3.665 ;
      RECT 69.96 3.39 70.22 3.665 ;
      RECT 70.025 3.377 70.155 3.665 ;
      RECT 69.57 4.466 69.585 4.859 ;
      RECT 69.535 4.471 69.585 4.858 ;
      RECT 69.57 4.47 69.63 4.857 ;
      RECT 69.515 4.481 69.63 4.856 ;
      RECT 69.53 4.477 69.63 4.856 ;
      RECT 69.495 4.487 69.705 4.853 ;
      RECT 69.495 4.506 69.75 4.851 ;
      RECT 69.495 4.513 69.755 4.848 ;
      RECT 69.48 4.49 69.705 4.845 ;
      RECT 69.46 4.495 69.705 4.838 ;
      RECT 69.455 4.499 69.705 4.834 ;
      RECT 69.455 4.516 69.765 4.833 ;
      RECT 69.435 4.51 69.75 4.829 ;
      RECT 69.435 4.519 69.77 4.823 ;
      RECT 69.43 4.525 69.77 4.595 ;
      RECT 69.495 4.485 69.63 4.853 ;
      RECT 69.37 3.848 69.57 4.16 ;
      RECT 69.445 3.826 69.57 4.16 ;
      RECT 69.385 3.845 69.575 4.145 ;
      RECT 69.355 3.856 69.575 4.143 ;
      RECT 69.37 3.851 69.58 4.109 ;
      RECT 69.355 3.955 69.585 4.076 ;
      RECT 69.385 3.827 69.57 4.16 ;
      RECT 69.445 3.805 69.545 4.16 ;
      RECT 69.47 3.802 69.545 4.16 ;
      RECT 69.47 3.797 69.49 4.16 ;
      RECT 68.875 3.865 69.05 4.04 ;
      RECT 68.87 3.865 69.05 4.038 ;
      RECT 68.845 3.865 69.05 4.033 ;
      RECT 68.79 3.845 68.96 4.023 ;
      RECT 68.79 3.852 69.025 4.023 ;
      RECT 68.875 4.532 68.89 4.715 ;
      RECT 68.865 4.51 68.875 4.715 ;
      RECT 68.85 4.49 68.865 4.715 ;
      RECT 68.84 4.465 68.85 4.715 ;
      RECT 68.81 4.43 68.84 4.715 ;
      RECT 68.775 4.37 68.81 4.715 ;
      RECT 68.77 4.332 68.775 4.715 ;
      RECT 68.72 4.283 68.77 4.715 ;
      RECT 68.71 4.233 68.72 4.703 ;
      RECT 68.695 4.212 68.71 4.663 ;
      RECT 68.675 4.18 68.695 4.613 ;
      RECT 68.65 4.136 68.675 4.553 ;
      RECT 68.645 4.108 68.65 4.508 ;
      RECT 68.64 4.099 68.645 4.494 ;
      RECT 68.635 4.092 68.64 4.481 ;
      RECT 68.63 4.087 68.635 4.47 ;
      RECT 68.625 4.072 68.63 4.46 ;
      RECT 68.62 4.05 68.625 4.447 ;
      RECT 68.61 4.01 68.62 4.422 ;
      RECT 68.585 3.94 68.61 4.378 ;
      RECT 68.58 3.88 68.585 4.343 ;
      RECT 68.565 3.86 68.58 4.31 ;
      RECT 68.56 3.86 68.565 4.285 ;
      RECT 68.53 3.86 68.56 4.24 ;
      RECT 68.485 3.86 68.53 4.18 ;
      RECT 68.41 3.86 68.485 4.128 ;
      RECT 68.405 3.86 68.41 4.093 ;
      RECT 68.4 3.86 68.405 4.083 ;
      RECT 68.395 3.86 68.4 4.063 ;
      RECT 68.66 3.08 68.83 3.55 ;
      RECT 68.605 3.073 68.8 3.534 ;
      RECT 68.605 3.087 68.835 3.533 ;
      RECT 68.59 3.088 68.835 3.514 ;
      RECT 68.585 3.106 68.835 3.5 ;
      RECT 68.59 3.089 68.84 3.498 ;
      RECT 68.575 3.12 68.84 3.483 ;
      RECT 68.59 3.095 68.845 3.468 ;
      RECT 68.57 3.135 68.845 3.465 ;
      RECT 68.585 3.107 68.85 3.45 ;
      RECT 68.585 3.119 68.855 3.43 ;
      RECT 68.57 3.135 68.86 3.413 ;
      RECT 68.57 3.145 68.865 3.268 ;
      RECT 68.565 3.145 68.865 3.225 ;
      RECT 68.565 3.16 68.87 3.203 ;
      RECT 68.66 3.07 68.8 3.55 ;
      RECT 68.66 3.068 68.77 3.55 ;
      RECT 68.746 3.065 68.77 3.55 ;
      RECT 68.405 4.732 68.41 4.778 ;
      RECT 68.395 4.58 68.405 4.802 ;
      RECT 68.39 4.425 68.395 4.827 ;
      RECT 68.375 4.387 68.39 4.838 ;
      RECT 68.37 4.37 68.375 4.845 ;
      RECT 68.36 4.358 68.37 4.852 ;
      RECT 68.355 4.349 68.36 4.854 ;
      RECT 68.35 4.347 68.355 4.858 ;
      RECT 68.305 4.338 68.35 4.873 ;
      RECT 68.3 4.33 68.305 4.887 ;
      RECT 68.295 4.327 68.3 4.891 ;
      RECT 68.28 4.322 68.295 4.899 ;
      RECT 68.225 4.312 68.28 4.91 ;
      RECT 68.19 4.3 68.225 4.911 ;
      RECT 68.181 4.295 68.19 4.905 ;
      RECT 68.095 4.295 68.181 4.895 ;
      RECT 68.065 4.295 68.095 4.873 ;
      RECT 68.055 4.295 68.06 4.853 ;
      RECT 68.05 4.295 68.055 4.815 ;
      RECT 68.045 4.295 68.05 4.773 ;
      RECT 68.04 4.295 68.045 4.733 ;
      RECT 68.035 4.295 68.04 4.663 ;
      RECT 68.025 4.295 68.035 4.585 ;
      RECT 68.02 4.295 68.025 4.485 ;
      RECT 68.06 4.295 68.065 4.855 ;
      RECT 67.555 4.377 67.645 4.855 ;
      RECT 67.54 4.38 67.66 4.853 ;
      RECT 67.555 4.379 67.66 4.853 ;
      RECT 67.52 4.386 67.685 4.843 ;
      RECT 67.54 4.38 67.685 4.843 ;
      RECT 67.505 4.392 67.685 4.831 ;
      RECT 67.54 4.383 67.735 4.824 ;
      RECT 67.491 4.4 67.735 4.822 ;
      RECT 67.52 4.39 67.745 4.81 ;
      RECT 67.491 4.411 67.775 4.801 ;
      RECT 67.405 4.435 67.775 4.795 ;
      RECT 67.405 4.448 67.815 4.778 ;
      RECT 67.4 4.47 67.815 4.771 ;
      RECT 67.37 4.485 67.815 4.761 ;
      RECT 67.365 4.496 67.815 4.751 ;
      RECT 67.335 4.509 67.815 4.742 ;
      RECT 67.32 4.527 67.815 4.731 ;
      RECT 67.295 4.54 67.815 4.721 ;
      RECT 67.555 4.376 67.565 4.855 ;
      RECT 67.601 3.8 67.64 4.045 ;
      RECT 67.515 3.8 67.65 4.043 ;
      RECT 67.4 3.825 67.65 4.04 ;
      RECT 67.4 3.825 67.655 4.038 ;
      RECT 67.4 3.825 67.67 4.033 ;
      RECT 67.506 3.8 67.685 4.013 ;
      RECT 67.42 3.808 67.685 4.013 ;
      RECT 67.09 3.16 67.26 3.595 ;
      RECT 67.08 3.194 67.26 3.578 ;
      RECT 67.16 3.13 67.33 3.565 ;
      RECT 67.065 3.205 67.33 3.543 ;
      RECT 67.16 3.14 67.335 3.533 ;
      RECT 67.09 3.192 67.365 3.518 ;
      RECT 67.05 3.218 67.365 3.503 ;
      RECT 67.05 3.26 67.375 3.483 ;
      RECT 67.045 3.285 67.38 3.465 ;
      RECT 67.045 3.295 67.385 3.45 ;
      RECT 67.04 3.232 67.365 3.448 ;
      RECT 67.04 3.305 67.39 3.433 ;
      RECT 67.035 3.242 67.365 3.43 ;
      RECT 67.03 3.326 67.395 3.413 ;
      RECT 67.03 3.358 67.4 3.393 ;
      RECT 67.025 3.272 67.375 3.385 ;
      RECT 67.03 3.257 67.365 3.413 ;
      RECT 67.045 3.227 67.365 3.465 ;
      RECT 66.89 3.814 67.115 4.07 ;
      RECT 66.89 3.847 67.135 4.06 ;
      RECT 66.855 3.847 67.135 4.058 ;
      RECT 66.855 3.86 67.14 4.048 ;
      RECT 66.855 3.88 67.15 4.04 ;
      RECT 66.855 3.977 67.155 4.033 ;
      RECT 66.835 3.725 66.965 4.023 ;
      RECT 66.79 3.88 67.15 3.965 ;
      RECT 66.78 3.725 66.965 3.91 ;
      RECT 66.78 3.757 67.051 3.91 ;
      RECT 66.745 4.287 66.765 4.465 ;
      RECT 66.71 4.24 66.745 4.465 ;
      RECT 66.695 4.18 66.71 4.465 ;
      RECT 66.67 4.127 66.695 4.465 ;
      RECT 66.655 4.08 66.67 4.465 ;
      RECT 66.635 4.057 66.655 4.465 ;
      RECT 66.61 4.022 66.635 4.465 ;
      RECT 66.6 3.868 66.61 4.465 ;
      RECT 66.57 3.863 66.6 4.456 ;
      RECT 66.565 3.86 66.57 4.446 ;
      RECT 66.55 3.86 66.565 4.42 ;
      RECT 66.545 3.86 66.55 4.383 ;
      RECT 66.52 3.86 66.545 4.335 ;
      RECT 66.5 3.86 66.52 4.26 ;
      RECT 66.49 3.86 66.5 4.22 ;
      RECT 66.485 3.86 66.49 4.195 ;
      RECT 66.48 3.86 66.485 4.178 ;
      RECT 66.475 3.86 66.48 4.16 ;
      RECT 66.47 3.861 66.475 4.15 ;
      RECT 66.46 3.863 66.47 4.118 ;
      RECT 66.45 3.865 66.46 4.085 ;
      RECT 66.44 3.868 66.45 4.058 ;
      RECT 66.765 4.295 66.99 4.465 ;
      RECT 66.095 3.107 66.265 3.56 ;
      RECT 66.095 3.107 66.355 3.526 ;
      RECT 66.095 3.107 66.385 3.51 ;
      RECT 66.095 3.107 66.415 3.483 ;
      RECT 66.351 3.085 66.43 3.465 ;
      RECT 66.13 3.092 66.435 3.45 ;
      RECT 66.13 3.1 66.445 3.413 ;
      RECT 66.09 3.127 66.445 3.385 ;
      RECT 66.075 3.14 66.445 3.35 ;
      RECT 66.095 3.115 66.465 3.34 ;
      RECT 66.07 3.18 66.465 3.31 ;
      RECT 66.07 3.21 66.47 3.293 ;
      RECT 66.065 3.24 66.47 3.28 ;
      RECT 66.13 3.089 66.43 3.465 ;
      RECT 66.265 3.086 66.351 3.544 ;
      RECT 66.216 3.087 66.43 3.465 ;
      RECT 66.36 4.747 66.405 4.94 ;
      RECT 66.35 4.717 66.36 4.94 ;
      RECT 66.345 4.702 66.35 4.94 ;
      RECT 66.305 4.612 66.345 4.94 ;
      RECT 66.3 4.525 66.305 4.94 ;
      RECT 66.29 4.495 66.3 4.94 ;
      RECT 66.285 4.455 66.29 4.94 ;
      RECT 66.275 4.417 66.285 4.94 ;
      RECT 66.27 4.382 66.275 4.94 ;
      RECT 66.25 4.335 66.27 4.94 ;
      RECT 66.235 4.26 66.25 4.94 ;
      RECT 66.23 4.215 66.235 4.935 ;
      RECT 66.225 4.195 66.23 4.908 ;
      RECT 66.22 4.175 66.225 4.893 ;
      RECT 66.215 4.15 66.22 4.873 ;
      RECT 66.21 4.128 66.215 4.858 ;
      RECT 66.205 4.106 66.21 4.84 ;
      RECT 66.2 4.085 66.205 4.83 ;
      RECT 66.19 4.057 66.2 4.8 ;
      RECT 66.18 4.02 66.19 4.768 ;
      RECT 66.17 3.98 66.18 4.735 ;
      RECT 66.16 3.958 66.17 4.705 ;
      RECT 66.13 3.91 66.16 4.637 ;
      RECT 66.115 3.87 66.13 4.564 ;
      RECT 66.105 3.87 66.115 4.53 ;
      RECT 66.1 3.87 66.105 4.505 ;
      RECT 66.095 3.87 66.1 4.49 ;
      RECT 66.09 3.87 66.095 4.468 ;
      RECT 66.085 3.87 66.09 4.455 ;
      RECT 66.07 3.87 66.085 4.42 ;
      RECT 66.05 3.87 66.07 4.36 ;
      RECT 66.04 3.87 66.05 4.31 ;
      RECT 66.02 3.87 66.04 4.258 ;
      RECT 66 3.87 66.02 4.215 ;
      RECT 65.99 3.87 66 4.203 ;
      RECT 65.96 3.87 65.99 4.19 ;
      RECT 65.93 3.891 65.96 4.17 ;
      RECT 65.92 3.919 65.93 4.15 ;
      RECT 65.905 3.936 65.92 4.118 ;
      RECT 65.9 3.95 65.905 4.085 ;
      RECT 65.895 3.958 65.9 4.058 ;
      RECT 65.89 3.966 65.895 4.02 ;
      RECT 65.895 4.49 65.9 4.825 ;
      RECT 65.86 4.477 65.895 4.824 ;
      RECT 65.79 4.417 65.86 4.823 ;
      RECT 65.71 4.36 65.79 4.822 ;
      RECT 65.575 4.32 65.71 4.821 ;
      RECT 65.575 4.507 65.91 4.81 ;
      RECT 65.535 4.507 65.91 4.8 ;
      RECT 65.535 4.525 65.915 4.795 ;
      RECT 65.535 4.615 65.92 4.785 ;
      RECT 65.53 4.31 65.695 4.765 ;
      RECT 65.525 4.31 65.695 4.508 ;
      RECT 65.525 4.467 65.89 4.508 ;
      RECT 65.525 4.455 65.885 4.508 ;
      RECT 64.655 7.305 64.825 8.775 ;
      RECT 64.655 7.305 64.83 8.565 ;
      RECT 64.285 9.255 64.755 9.425 ;
      RECT 64.285 8.235 64.455 9.425 ;
      RECT 64.28 3.035 64.45 4.225 ;
      RECT 64.28 3.035 64.75 3.205 ;
      RECT 63.665 3.895 63.84 5.155 ;
      RECT 63.665 3.685 63.835 5.155 ;
      RECT 63.665 7.305 63.835 8.775 ;
      RECT 63.665 7.305 63.84 8.565 ;
      RECT 63.295 3.035 63.465 4.225 ;
      RECT 63.295 3.035 63.765 3.205 ;
      RECT 63.295 9.255 63.765 9.425 ;
      RECT 63.295 8.235 63.465 9.425 ;
      RECT 62.305 4.015 62.48 5.155 ;
      RECT 62.305 1.865 62.475 5.155 ;
      RECT 62.305 1.865 62.48 2.415 ;
      RECT 62.305 10.045 62.48 10.595 ;
      RECT 62.305 7.305 62.475 10.595 ;
      RECT 62.305 7.305 62.48 8.445 ;
      RECT 61.875 3.895 62.05 5.155 ;
      RECT 61.875 2.945 62.045 5.155 ;
      RECT 61.875 7.305 62.045 9.515 ;
      RECT 61.875 7.305 62.05 8.565 ;
      RECT 61.445 3.925 61.615 5.155 ;
      RECT 61.505 2.145 61.675 4.095 ;
      RECT 61.445 1.865 61.615 2.315 ;
      RECT 61.445 10.145 61.615 10.595 ;
      RECT 61.505 8.365 61.675 10.315 ;
      RECT 61.445 7.305 61.615 8.535 ;
      RECT 60.92 3.895 61.095 5.155 ;
      RECT 60.92 1.865 61.09 5.155 ;
      RECT 60.92 3.365 61.33 3.695 ;
      RECT 60.92 2.525 61.33 2.855 ;
      RECT 60.92 1.865 61.095 2.355 ;
      RECT 60.92 10.105 61.095 10.595 ;
      RECT 60.92 7.305 61.09 10.595 ;
      RECT 60.92 9.605 61.33 9.935 ;
      RECT 60.92 8.765 61.33 9.095 ;
      RECT 60.92 7.305 61.095 8.565 ;
      RECT 58.26 3.27 58.99 3.51 ;
      RECT 58.802 3.065 58.99 3.51 ;
      RECT 58.63 3.077 59.005 3.504 ;
      RECT 58.545 3.092 59.025 3.489 ;
      RECT 58.545 3.107 59.03 3.479 ;
      RECT 58.5 3.127 59.045 3.471 ;
      RECT 58.477 3.162 59.06 3.425 ;
      RECT 58.391 3.185 59.065 3.385 ;
      RECT 58.391 3.203 59.075 3.355 ;
      RECT 58.26 3.272 59.08 3.318 ;
      RECT 58.305 3.215 59.075 3.355 ;
      RECT 58.391 3.167 59.06 3.425 ;
      RECT 58.477 3.136 59.045 3.471 ;
      RECT 58.5 3.117 59.03 3.479 ;
      RECT 58.545 3.09 59.005 3.504 ;
      RECT 58.63 3.072 58.99 3.51 ;
      RECT 58.716 3.066 58.99 3.51 ;
      RECT 58.802 3.061 58.935 3.51 ;
      RECT 58.888 3.056 58.935 3.51 ;
      RECT 58.45 4.67 58.455 4.683 ;
      RECT 58.445 4.565 58.45 4.688 ;
      RECT 58.42 4.425 58.445 4.703 ;
      RECT 58.385 4.376 58.42 4.735 ;
      RECT 58.38 4.344 58.385 4.755 ;
      RECT 58.375 4.335 58.38 4.755 ;
      RECT 58.295 4.3 58.375 4.755 ;
      RECT 58.232 4.27 58.295 4.755 ;
      RECT 58.146 4.258 58.232 4.755 ;
      RECT 58.06 4.244 58.146 4.755 ;
      RECT 57.98 4.231 58.06 4.741 ;
      RECT 57.945 4.223 57.98 4.721 ;
      RECT 57.935 4.22 57.945 4.712 ;
      RECT 57.905 4.215 57.935 4.699 ;
      RECT 57.855 4.19 57.905 4.675 ;
      RECT 57.841 4.164 57.855 4.657 ;
      RECT 57.755 4.124 57.841 4.633 ;
      RECT 57.71 4.072 57.755 4.602 ;
      RECT 57.7 4.047 57.71 4.589 ;
      RECT 57.695 3.828 57.7 3.85 ;
      RECT 57.69 4.03 57.7 4.585 ;
      RECT 57.69 3.826 57.695 3.94 ;
      RECT 57.68 3.822 57.69 4.581 ;
      RECT 57.636 3.82 57.68 4.569 ;
      RECT 57.55 3.82 57.636 4.54 ;
      RECT 57.52 3.82 57.55 4.513 ;
      RECT 57.505 3.82 57.52 4.501 ;
      RECT 57.465 3.832 57.505 4.486 ;
      RECT 57.445 3.851 57.465 4.465 ;
      RECT 57.435 3.861 57.445 4.449 ;
      RECT 57.425 3.867 57.435 4.438 ;
      RECT 57.405 3.877 57.425 4.421 ;
      RECT 57.4 3.886 57.405 4.408 ;
      RECT 57.395 3.89 57.4 4.358 ;
      RECT 57.385 3.896 57.395 4.275 ;
      RECT 57.38 3.9 57.385 4.189 ;
      RECT 57.375 3.92 57.38 4.126 ;
      RECT 57.37 3.943 57.375 4.073 ;
      RECT 57.365 3.961 57.37 4.018 ;
      RECT 57.975 3.78 58.145 4.04 ;
      RECT 58.145 3.745 58.19 4.026 ;
      RECT 58.106 3.747 58.195 4.009 ;
      RECT 57.995 3.764 58.281 3.98 ;
      RECT 57.995 3.779 58.285 3.952 ;
      RECT 57.995 3.76 58.195 4.009 ;
      RECT 58.02 3.748 58.145 4.04 ;
      RECT 58.106 3.746 58.19 4.026 ;
      RECT 57.525 10.045 57.7 10.595 ;
      RECT 57.525 7.305 57.695 10.595 ;
      RECT 57.525 7.305 57.7 8.445 ;
      RECT 57.16 3.135 57.33 3.625 ;
      RECT 57.16 3.135 57.365 3.605 ;
      RECT 57.295 3.055 57.405 3.565 ;
      RECT 57.276 3.059 57.425 3.535 ;
      RECT 57.19 3.067 57.445 3.518 ;
      RECT 57.19 3.073 57.45 3.508 ;
      RECT 57.19 3.082 57.47 3.496 ;
      RECT 57.165 3.107 57.5 3.474 ;
      RECT 57.165 3.127 57.505 3.454 ;
      RECT 57.16 3.14 57.515 3.434 ;
      RECT 57.16 3.207 57.52 3.415 ;
      RECT 57.16 3.34 57.525 3.402 ;
      RECT 57.155 3.145 57.515 3.235 ;
      RECT 57.165 3.102 57.47 3.496 ;
      RECT 57.276 3.057 57.405 3.565 ;
      RECT 57.15 4.81 57.45 5.065 ;
      RECT 57.235 4.776 57.45 5.065 ;
      RECT 57.235 4.779 57.455 4.925 ;
      RECT 57.17 4.8 57.455 4.925 ;
      RECT 57.205 4.79 57.45 5.065 ;
      RECT 57.2 4.795 57.455 4.925 ;
      RECT 57.235 4.774 57.436 5.065 ;
      RECT 57.321 4.765 57.436 5.065 ;
      RECT 57.321 4.759 57.35 5.065 ;
      RECT 57.095 7.305 57.265 9.515 ;
      RECT 57.095 7.305 57.27 8.565 ;
      RECT 56.81 4.4 56.82 4.89 ;
      RECT 56.47 4.335 56.48 4.635 ;
      RECT 56.985 4.507 56.99 4.726 ;
      RECT 56.975 4.487 56.985 4.743 ;
      RECT 56.965 4.467 56.975 4.773 ;
      RECT 56.96 4.457 56.965 4.788 ;
      RECT 56.955 4.453 56.96 4.793 ;
      RECT 56.94 4.445 56.955 4.8 ;
      RECT 56.9 4.425 56.94 4.825 ;
      RECT 56.875 4.407 56.9 4.858 ;
      RECT 56.87 4.405 56.875 4.871 ;
      RECT 56.85 4.402 56.87 4.875 ;
      RECT 56.82 4.4 56.85 4.885 ;
      RECT 56.75 4.402 56.81 4.886 ;
      RECT 56.73 4.402 56.75 4.88 ;
      RECT 56.705 4.4 56.73 4.877 ;
      RECT 56.67 4.395 56.705 4.873 ;
      RECT 56.65 4.389 56.67 4.86 ;
      RECT 56.64 4.386 56.65 4.848 ;
      RECT 56.62 4.383 56.64 4.833 ;
      RECT 56.6 4.379 56.62 4.815 ;
      RECT 56.595 4.376 56.6 4.805 ;
      RECT 56.59 4.375 56.595 4.803 ;
      RECT 56.58 4.372 56.59 4.795 ;
      RECT 56.57 4.366 56.58 4.778 ;
      RECT 56.56 4.36 56.57 4.76 ;
      RECT 56.55 4.354 56.56 4.748 ;
      RECT 56.54 4.348 56.55 4.728 ;
      RECT 56.535 4.344 56.54 4.713 ;
      RECT 56.53 4.342 56.535 4.705 ;
      RECT 56.525 4.34 56.53 4.698 ;
      RECT 56.52 4.338 56.525 4.688 ;
      RECT 56.515 4.336 56.52 4.682 ;
      RECT 56.505 4.335 56.515 4.672 ;
      RECT 56.495 4.335 56.505 4.663 ;
      RECT 56.48 4.335 56.495 4.648 ;
      RECT 56.44 4.335 56.47 4.632 ;
      RECT 56.42 4.337 56.44 4.627 ;
      RECT 56.415 4.342 56.42 4.625 ;
      RECT 56.385 4.35 56.415 4.623 ;
      RECT 56.355 4.365 56.385 4.622 ;
      RECT 56.31 4.387 56.355 4.627 ;
      RECT 56.305 4.402 56.31 4.631 ;
      RECT 56.29 4.407 56.305 4.633 ;
      RECT 56.285 4.411 56.29 4.635 ;
      RECT 56.225 4.434 56.285 4.644 ;
      RECT 56.205 4.46 56.225 4.657 ;
      RECT 56.195 4.467 56.205 4.661 ;
      RECT 56.18 4.474 56.195 4.664 ;
      RECT 56.16 4.484 56.18 4.667 ;
      RECT 56.155 4.492 56.16 4.67 ;
      RECT 56.11 4.497 56.155 4.677 ;
      RECT 56.1 4.5 56.11 4.684 ;
      RECT 56.09 4.5 56.1 4.688 ;
      RECT 56.055 4.502 56.09 4.7 ;
      RECT 56.035 4.505 56.055 4.713 ;
      RECT 55.995 4.508 56.035 4.724 ;
      RECT 55.98 4.51 55.995 4.737 ;
      RECT 55.97 4.51 55.98 4.742 ;
      RECT 55.945 4.511 55.97 4.75 ;
      RECT 55.935 4.513 55.945 4.755 ;
      RECT 55.93 4.514 55.935 4.758 ;
      RECT 55.905 4.512 55.93 4.761 ;
      RECT 55.89 4.51 55.905 4.762 ;
      RECT 55.87 4.507 55.89 4.764 ;
      RECT 55.85 4.502 55.87 4.764 ;
      RECT 55.79 4.497 55.85 4.761 ;
      RECT 55.755 4.472 55.79 4.757 ;
      RECT 55.745 4.449 55.755 4.755 ;
      RECT 55.715 4.426 55.745 4.755 ;
      RECT 55.705 4.405 55.715 4.755 ;
      RECT 55.68 4.387 55.705 4.753 ;
      RECT 55.665 4.365 55.68 4.75 ;
      RECT 55.65 4.347 55.665 4.748 ;
      RECT 55.63 4.337 55.65 4.746 ;
      RECT 55.615 4.332 55.63 4.745 ;
      RECT 55.6 4.33 55.615 4.744 ;
      RECT 55.57 4.331 55.6 4.742 ;
      RECT 55.55 4.334 55.57 4.74 ;
      RECT 55.493 4.338 55.55 4.74 ;
      RECT 55.407 4.347 55.493 4.74 ;
      RECT 55.321 4.358 55.407 4.74 ;
      RECT 55.235 4.369 55.321 4.74 ;
      RECT 55.215 4.376 55.235 4.748 ;
      RECT 55.205 4.379 55.215 4.755 ;
      RECT 55.14 4.384 55.205 4.773 ;
      RECT 55.11 4.391 55.14 4.798 ;
      RECT 55.1 4.394 55.11 4.805 ;
      RECT 55.055 4.398 55.1 4.81 ;
      RECT 55.025 4.403 55.055 4.815 ;
      RECT 55.024 4.405 55.025 4.815 ;
      RECT 54.938 4.411 55.024 4.815 ;
      RECT 54.852 4.422 54.938 4.815 ;
      RECT 54.766 4.434 54.852 4.815 ;
      RECT 54.68 4.445 54.766 4.815 ;
      RECT 54.665 4.452 54.68 4.81 ;
      RECT 54.66 4.454 54.665 4.804 ;
      RECT 54.64 4.465 54.66 4.799 ;
      RECT 54.63 4.483 54.64 4.793 ;
      RECT 54.625 4.495 54.63 4.593 ;
      RECT 56.92 3.248 56.94 3.335 ;
      RECT 56.915 3.183 56.92 3.367 ;
      RECT 56.905 3.15 56.915 3.372 ;
      RECT 56.9 3.13 56.905 3.378 ;
      RECT 56.87 3.13 56.9 3.395 ;
      RECT 56.821 3.13 56.87 3.431 ;
      RECT 56.735 3.13 56.821 3.489 ;
      RECT 56.706 3.14 56.735 3.538 ;
      RECT 56.62 3.182 56.706 3.591 ;
      RECT 56.6 3.22 56.62 3.638 ;
      RECT 56.575 3.237 56.6 3.658 ;
      RECT 56.565 3.251 56.575 3.678 ;
      RECT 56.56 3.257 56.565 3.688 ;
      RECT 56.555 3.261 56.56 3.695 ;
      RECT 56.505 3.281 56.555 3.7 ;
      RECT 56.44 3.325 56.505 3.7 ;
      RECT 56.415 3.375 56.44 3.7 ;
      RECT 56.405 3.405 56.415 3.7 ;
      RECT 56.4 3.432 56.405 3.7 ;
      RECT 56.395 3.45 56.4 3.7 ;
      RECT 56.385 3.492 56.395 3.7 ;
      RECT 56.14 10.105 56.315 10.595 ;
      RECT 56.14 7.305 56.31 10.595 ;
      RECT 56.14 9.605 56.55 9.935 ;
      RECT 56.14 8.765 56.55 9.095 ;
      RECT 56.14 7.305 56.315 8.565 ;
      RECT 56.215 4.85 56.405 5.075 ;
      RECT 56.205 4.851 56.41 5.07 ;
      RECT 56.205 4.853 56.42 5.05 ;
      RECT 56.205 4.857 56.425 5.035 ;
      RECT 56.205 4.844 56.375 5.07 ;
      RECT 56.205 4.847 56.4 5.07 ;
      RECT 56.215 4.843 56.375 5.075 ;
      RECT 56.301 4.841 56.375 5.075 ;
      RECT 55.925 4.092 56.095 4.33 ;
      RECT 55.925 4.092 56.181 4.244 ;
      RECT 55.925 4.092 56.185 4.154 ;
      RECT 55.975 3.865 56.195 4.133 ;
      RECT 55.97 3.882 56.2 4.106 ;
      RECT 55.935 4.04 56.2 4.106 ;
      RECT 55.955 3.89 56.095 4.33 ;
      RECT 55.945 3.972 56.205 4.089 ;
      RECT 55.94 4.02 56.205 4.089 ;
      RECT 55.945 3.93 56.2 4.106 ;
      RECT 55.97 3.867 56.195 4.133 ;
      RECT 55.535 3.842 55.705 4.04 ;
      RECT 55.535 3.842 55.75 4.015 ;
      RECT 55.605 3.785 55.775 3.973 ;
      RECT 55.58 3.8 55.775 3.973 ;
      RECT 55.195 3.846 55.225 4.04 ;
      RECT 55.19 3.818 55.195 4.04 ;
      RECT 55.16 3.792 55.19 4.042 ;
      RECT 55.135 3.75 55.16 4.045 ;
      RECT 55.125 3.722 55.135 4.047 ;
      RECT 55.09 3.702 55.125 4.049 ;
      RECT 55.025 3.687 55.09 4.055 ;
      RECT 54.975 3.685 55.025 4.061 ;
      RECT 54.952 3.687 54.975 4.066 ;
      RECT 54.866 3.698 54.952 4.072 ;
      RECT 54.78 3.716 54.866 4.082 ;
      RECT 54.765 3.727 54.78 4.088 ;
      RECT 54.695 3.75 54.765 4.094 ;
      RECT 54.64 3.782 54.695 4.102 ;
      RECT 54.6 3.805 54.64 4.108 ;
      RECT 54.586 3.818 54.6 4.111 ;
      RECT 54.5 3.84 54.586 4.117 ;
      RECT 54.485 3.865 54.5 4.123 ;
      RECT 54.445 3.88 54.485 4.127 ;
      RECT 54.395 3.895 54.445 4.132 ;
      RECT 54.37 3.902 54.395 4.136 ;
      RECT 54.31 3.897 54.37 4.14 ;
      RECT 54.295 3.888 54.31 4.144 ;
      RECT 54.225 3.878 54.295 4.14 ;
      RECT 54.2 3.87 54.22 4.13 ;
      RECT 54.141 3.87 54.2 4.108 ;
      RECT 54.055 3.87 54.141 4.065 ;
      RECT 54.22 3.87 54.225 4.135 ;
      RECT 54.915 3.101 55.085 3.435 ;
      RECT 54.885 3.101 55.085 3.43 ;
      RECT 54.825 3.068 54.885 3.418 ;
      RECT 54.825 3.124 55.095 3.413 ;
      RECT 54.8 3.124 55.095 3.407 ;
      RECT 54.795 3.065 54.825 3.404 ;
      RECT 54.78 3.071 54.915 3.402 ;
      RECT 54.775 3.079 55 3.39 ;
      RECT 54.775 3.131 55.11 3.343 ;
      RECT 54.76 3.087 55 3.338 ;
      RECT 54.76 3.157 55.12 3.279 ;
      RECT 54.73 3.107 55.085 3.24 ;
      RECT 54.73 3.197 55.13 3.236 ;
      RECT 54.78 3.076 55 3.402 ;
      RECT 54.12 3.406 54.175 3.67 ;
      RECT 54.12 3.406 54.24 3.669 ;
      RECT 54.12 3.406 54.265 3.668 ;
      RECT 54.12 3.406 54.33 3.667 ;
      RECT 54.265 3.372 54.345 3.666 ;
      RECT 54.08 3.416 54.49 3.665 ;
      RECT 54.12 3.413 54.49 3.665 ;
      RECT 54.08 3.421 54.495 3.658 ;
      RECT 54.065 3.423 54.495 3.657 ;
      RECT 54.065 3.43 54.5 3.653 ;
      RECT 54.045 3.429 54.495 3.649 ;
      RECT 54.045 3.437 54.505 3.648 ;
      RECT 54.04 3.434 54.5 3.644 ;
      RECT 54.04 3.447 54.515 3.643 ;
      RECT 54.025 3.437 54.505 3.642 ;
      RECT 53.99 3.45 54.515 3.635 ;
      RECT 54.175 3.405 54.485 3.665 ;
      RECT 54.175 3.39 54.435 3.665 ;
      RECT 54.24 3.377 54.37 3.665 ;
      RECT 53.785 4.466 53.8 4.859 ;
      RECT 53.75 4.471 53.8 4.858 ;
      RECT 53.785 4.47 53.845 4.857 ;
      RECT 53.73 4.481 53.845 4.856 ;
      RECT 53.745 4.477 53.845 4.856 ;
      RECT 53.71 4.487 53.92 4.853 ;
      RECT 53.71 4.506 53.965 4.851 ;
      RECT 53.71 4.513 53.97 4.848 ;
      RECT 53.695 4.49 53.92 4.845 ;
      RECT 53.675 4.495 53.92 4.838 ;
      RECT 53.67 4.499 53.92 4.834 ;
      RECT 53.67 4.516 53.98 4.833 ;
      RECT 53.65 4.51 53.965 4.829 ;
      RECT 53.65 4.519 53.985 4.823 ;
      RECT 53.645 4.525 53.985 4.595 ;
      RECT 53.71 4.485 53.845 4.853 ;
      RECT 53.585 3.848 53.785 4.16 ;
      RECT 53.66 3.826 53.785 4.16 ;
      RECT 53.6 3.845 53.79 4.145 ;
      RECT 53.57 3.856 53.79 4.143 ;
      RECT 53.585 3.851 53.795 4.109 ;
      RECT 53.57 3.955 53.8 4.076 ;
      RECT 53.6 3.827 53.785 4.16 ;
      RECT 53.66 3.805 53.76 4.16 ;
      RECT 53.685 3.802 53.76 4.16 ;
      RECT 53.685 3.797 53.705 4.16 ;
      RECT 53.09 3.865 53.265 4.04 ;
      RECT 53.085 3.865 53.265 4.038 ;
      RECT 53.06 3.865 53.265 4.033 ;
      RECT 53.005 3.845 53.175 4.023 ;
      RECT 53.005 3.852 53.24 4.023 ;
      RECT 53.09 4.532 53.105 4.715 ;
      RECT 53.08 4.51 53.09 4.715 ;
      RECT 53.065 4.49 53.08 4.715 ;
      RECT 53.055 4.465 53.065 4.715 ;
      RECT 53.025 4.43 53.055 4.715 ;
      RECT 52.99 4.37 53.025 4.715 ;
      RECT 52.985 4.332 52.99 4.715 ;
      RECT 52.935 4.283 52.985 4.715 ;
      RECT 52.925 4.233 52.935 4.703 ;
      RECT 52.91 4.212 52.925 4.663 ;
      RECT 52.89 4.18 52.91 4.613 ;
      RECT 52.865 4.136 52.89 4.553 ;
      RECT 52.86 4.108 52.865 4.508 ;
      RECT 52.855 4.099 52.86 4.494 ;
      RECT 52.85 4.092 52.855 4.481 ;
      RECT 52.845 4.087 52.85 4.47 ;
      RECT 52.84 4.072 52.845 4.46 ;
      RECT 52.835 4.05 52.84 4.447 ;
      RECT 52.825 4.01 52.835 4.422 ;
      RECT 52.8 3.94 52.825 4.378 ;
      RECT 52.795 3.88 52.8 4.343 ;
      RECT 52.78 3.86 52.795 4.31 ;
      RECT 52.775 3.86 52.78 4.285 ;
      RECT 52.745 3.86 52.775 4.24 ;
      RECT 52.7 3.86 52.745 4.18 ;
      RECT 52.625 3.86 52.7 4.128 ;
      RECT 52.62 3.86 52.625 4.093 ;
      RECT 52.615 3.86 52.62 4.083 ;
      RECT 52.61 3.86 52.615 4.063 ;
      RECT 52.875 3.08 53.045 3.55 ;
      RECT 52.82 3.073 53.015 3.534 ;
      RECT 52.82 3.087 53.05 3.533 ;
      RECT 52.805 3.088 53.05 3.514 ;
      RECT 52.8 3.106 53.05 3.5 ;
      RECT 52.805 3.089 53.055 3.498 ;
      RECT 52.79 3.12 53.055 3.483 ;
      RECT 52.805 3.095 53.06 3.468 ;
      RECT 52.785 3.135 53.06 3.465 ;
      RECT 52.8 3.107 53.065 3.45 ;
      RECT 52.8 3.119 53.07 3.43 ;
      RECT 52.785 3.135 53.075 3.413 ;
      RECT 52.785 3.145 53.08 3.268 ;
      RECT 52.78 3.145 53.08 3.225 ;
      RECT 52.78 3.16 53.085 3.203 ;
      RECT 52.875 3.07 53.015 3.55 ;
      RECT 52.875 3.068 52.985 3.55 ;
      RECT 52.961 3.065 52.985 3.55 ;
      RECT 52.62 4.732 52.625 4.778 ;
      RECT 52.61 4.58 52.62 4.802 ;
      RECT 52.605 4.425 52.61 4.827 ;
      RECT 52.59 4.387 52.605 4.838 ;
      RECT 52.585 4.37 52.59 4.845 ;
      RECT 52.575 4.358 52.585 4.852 ;
      RECT 52.57 4.349 52.575 4.854 ;
      RECT 52.565 4.347 52.57 4.858 ;
      RECT 52.52 4.338 52.565 4.873 ;
      RECT 52.515 4.33 52.52 4.887 ;
      RECT 52.51 4.327 52.515 4.891 ;
      RECT 52.495 4.322 52.51 4.899 ;
      RECT 52.44 4.312 52.495 4.91 ;
      RECT 52.405 4.3 52.44 4.911 ;
      RECT 52.396 4.295 52.405 4.905 ;
      RECT 52.31 4.295 52.396 4.895 ;
      RECT 52.28 4.295 52.31 4.873 ;
      RECT 52.27 4.295 52.275 4.853 ;
      RECT 52.265 4.295 52.27 4.815 ;
      RECT 52.26 4.295 52.265 4.773 ;
      RECT 52.255 4.295 52.26 4.733 ;
      RECT 52.25 4.295 52.255 4.663 ;
      RECT 52.24 4.295 52.25 4.585 ;
      RECT 52.235 4.295 52.24 4.485 ;
      RECT 52.275 4.295 52.28 4.855 ;
      RECT 51.77 4.377 51.86 4.855 ;
      RECT 51.755 4.38 51.875 4.853 ;
      RECT 51.77 4.379 51.875 4.853 ;
      RECT 51.735 4.386 51.9 4.843 ;
      RECT 51.755 4.38 51.9 4.843 ;
      RECT 51.72 4.392 51.9 4.831 ;
      RECT 51.755 4.383 51.95 4.824 ;
      RECT 51.706 4.4 51.95 4.822 ;
      RECT 51.735 4.39 51.96 4.81 ;
      RECT 51.706 4.411 51.99 4.801 ;
      RECT 51.62 4.435 51.99 4.795 ;
      RECT 51.62 4.448 52.03 4.778 ;
      RECT 51.615 4.47 52.03 4.771 ;
      RECT 51.585 4.485 52.03 4.761 ;
      RECT 51.58 4.496 52.03 4.751 ;
      RECT 51.55 4.509 52.03 4.742 ;
      RECT 51.535 4.527 52.03 4.731 ;
      RECT 51.51 4.54 52.03 4.721 ;
      RECT 51.77 4.376 51.78 4.855 ;
      RECT 51.816 3.8 51.855 4.045 ;
      RECT 51.73 3.8 51.865 4.043 ;
      RECT 51.615 3.825 51.865 4.04 ;
      RECT 51.615 3.825 51.87 4.038 ;
      RECT 51.615 3.825 51.885 4.033 ;
      RECT 51.721 3.8 51.9 4.013 ;
      RECT 51.635 3.808 51.9 4.013 ;
      RECT 51.305 3.16 51.475 3.595 ;
      RECT 51.295 3.194 51.475 3.578 ;
      RECT 51.375 3.13 51.545 3.565 ;
      RECT 51.28 3.205 51.545 3.543 ;
      RECT 51.375 3.14 51.55 3.533 ;
      RECT 51.305 3.192 51.58 3.518 ;
      RECT 51.265 3.218 51.58 3.503 ;
      RECT 51.265 3.26 51.59 3.483 ;
      RECT 51.26 3.285 51.595 3.465 ;
      RECT 51.26 3.295 51.6 3.45 ;
      RECT 51.255 3.232 51.58 3.448 ;
      RECT 51.255 3.305 51.605 3.433 ;
      RECT 51.25 3.242 51.58 3.43 ;
      RECT 51.245 3.326 51.61 3.413 ;
      RECT 51.245 3.358 51.615 3.393 ;
      RECT 51.24 3.272 51.59 3.385 ;
      RECT 51.245 3.257 51.58 3.413 ;
      RECT 51.26 3.227 51.58 3.465 ;
      RECT 51.105 3.814 51.33 4.07 ;
      RECT 51.105 3.847 51.35 4.06 ;
      RECT 51.07 3.847 51.35 4.058 ;
      RECT 51.07 3.86 51.355 4.048 ;
      RECT 51.07 3.88 51.365 4.04 ;
      RECT 51.07 3.977 51.37 4.033 ;
      RECT 51.05 3.725 51.18 4.023 ;
      RECT 51.005 3.88 51.365 3.965 ;
      RECT 50.995 3.725 51.18 3.91 ;
      RECT 50.995 3.757 51.266 3.91 ;
      RECT 50.96 4.287 50.98 4.465 ;
      RECT 50.925 4.24 50.96 4.465 ;
      RECT 50.91 4.18 50.925 4.465 ;
      RECT 50.885 4.127 50.91 4.465 ;
      RECT 50.87 4.08 50.885 4.465 ;
      RECT 50.85 4.057 50.87 4.465 ;
      RECT 50.825 4.022 50.85 4.465 ;
      RECT 50.815 3.868 50.825 4.465 ;
      RECT 50.785 3.863 50.815 4.456 ;
      RECT 50.78 3.86 50.785 4.446 ;
      RECT 50.765 3.86 50.78 4.42 ;
      RECT 50.76 3.86 50.765 4.383 ;
      RECT 50.735 3.86 50.76 4.335 ;
      RECT 50.715 3.86 50.735 4.26 ;
      RECT 50.705 3.86 50.715 4.22 ;
      RECT 50.7 3.86 50.705 4.195 ;
      RECT 50.695 3.86 50.7 4.178 ;
      RECT 50.69 3.86 50.695 4.16 ;
      RECT 50.685 3.861 50.69 4.15 ;
      RECT 50.675 3.863 50.685 4.118 ;
      RECT 50.665 3.865 50.675 4.085 ;
      RECT 50.655 3.868 50.665 4.058 ;
      RECT 50.98 4.295 51.205 4.465 ;
      RECT 50.31 3.107 50.48 3.56 ;
      RECT 50.31 3.107 50.57 3.526 ;
      RECT 50.31 3.107 50.6 3.51 ;
      RECT 50.31 3.107 50.63 3.483 ;
      RECT 50.566 3.085 50.645 3.465 ;
      RECT 50.345 3.092 50.65 3.45 ;
      RECT 50.345 3.1 50.66 3.413 ;
      RECT 50.305 3.127 50.66 3.385 ;
      RECT 50.29 3.14 50.66 3.35 ;
      RECT 50.31 3.115 50.68 3.34 ;
      RECT 50.285 3.18 50.68 3.31 ;
      RECT 50.285 3.21 50.685 3.293 ;
      RECT 50.28 3.24 50.685 3.28 ;
      RECT 50.345 3.089 50.645 3.465 ;
      RECT 50.48 3.086 50.566 3.544 ;
      RECT 50.431 3.087 50.645 3.465 ;
      RECT 50.575 4.747 50.62 4.94 ;
      RECT 50.565 4.717 50.575 4.94 ;
      RECT 50.56 4.702 50.565 4.94 ;
      RECT 50.52 4.612 50.56 4.94 ;
      RECT 50.515 4.525 50.52 4.94 ;
      RECT 50.505 4.495 50.515 4.94 ;
      RECT 50.5 4.455 50.505 4.94 ;
      RECT 50.49 4.417 50.5 4.94 ;
      RECT 50.485 4.382 50.49 4.94 ;
      RECT 50.465 4.335 50.485 4.94 ;
      RECT 50.45 4.26 50.465 4.94 ;
      RECT 50.445 4.215 50.45 4.935 ;
      RECT 50.44 4.195 50.445 4.908 ;
      RECT 50.435 4.175 50.44 4.893 ;
      RECT 50.43 4.15 50.435 4.873 ;
      RECT 50.425 4.128 50.43 4.858 ;
      RECT 50.42 4.106 50.425 4.84 ;
      RECT 50.415 4.085 50.42 4.83 ;
      RECT 50.405 4.057 50.415 4.8 ;
      RECT 50.395 4.02 50.405 4.768 ;
      RECT 50.385 3.98 50.395 4.735 ;
      RECT 50.375 3.958 50.385 4.705 ;
      RECT 50.345 3.91 50.375 4.637 ;
      RECT 50.33 3.87 50.345 4.564 ;
      RECT 50.32 3.87 50.33 4.53 ;
      RECT 50.315 3.87 50.32 4.505 ;
      RECT 50.31 3.87 50.315 4.49 ;
      RECT 50.305 3.87 50.31 4.468 ;
      RECT 50.3 3.87 50.305 4.455 ;
      RECT 50.285 3.87 50.3 4.42 ;
      RECT 50.265 3.87 50.285 4.36 ;
      RECT 50.255 3.87 50.265 4.31 ;
      RECT 50.235 3.87 50.255 4.258 ;
      RECT 50.215 3.87 50.235 4.215 ;
      RECT 50.205 3.87 50.215 4.203 ;
      RECT 50.175 3.87 50.205 4.19 ;
      RECT 50.145 3.891 50.175 4.17 ;
      RECT 50.135 3.919 50.145 4.15 ;
      RECT 50.12 3.936 50.135 4.118 ;
      RECT 50.115 3.95 50.12 4.085 ;
      RECT 50.11 3.958 50.115 4.058 ;
      RECT 50.105 3.966 50.11 4.02 ;
      RECT 50.11 4.49 50.115 4.825 ;
      RECT 50.075 4.477 50.11 4.824 ;
      RECT 50.005 4.417 50.075 4.823 ;
      RECT 49.925 4.36 50.005 4.822 ;
      RECT 49.79 4.32 49.925 4.821 ;
      RECT 49.79 4.507 50.125 4.81 ;
      RECT 49.75 4.507 50.125 4.8 ;
      RECT 49.75 4.525 50.13 4.795 ;
      RECT 49.75 4.615 50.135 4.785 ;
      RECT 49.745 4.31 49.91 4.765 ;
      RECT 49.74 4.31 49.91 4.508 ;
      RECT 49.74 4.467 50.105 4.508 ;
      RECT 49.74 4.455 50.1 4.508 ;
      RECT 48.88 7.305 49.05 8.775 ;
      RECT 48.88 7.305 49.055 8.565 ;
      RECT 48.51 9.255 48.98 9.425 ;
      RECT 48.51 8.235 48.68 9.425 ;
      RECT 48.505 3.035 48.675 4.225 ;
      RECT 48.505 3.035 48.975 3.205 ;
      RECT 47.89 3.895 48.065 5.155 ;
      RECT 47.89 3.685 48.06 5.155 ;
      RECT 47.89 7.305 48.06 8.775 ;
      RECT 47.89 7.305 48.065 8.565 ;
      RECT 47.52 3.035 47.69 4.225 ;
      RECT 47.52 3.035 47.99 3.205 ;
      RECT 47.52 9.255 47.99 9.425 ;
      RECT 47.52 8.235 47.69 9.425 ;
      RECT 46.53 4.015 46.705 5.155 ;
      RECT 46.53 1.865 46.7 5.155 ;
      RECT 46.53 1.865 46.705 2.415 ;
      RECT 46.53 10.045 46.705 10.595 ;
      RECT 46.53 7.305 46.7 10.595 ;
      RECT 46.53 7.305 46.705 8.445 ;
      RECT 46.1 3.895 46.275 5.155 ;
      RECT 46.1 2.945 46.27 5.155 ;
      RECT 46.1 7.305 46.27 9.515 ;
      RECT 46.1 7.305 46.275 8.565 ;
      RECT 45.67 3.925 45.84 5.155 ;
      RECT 45.73 2.145 45.9 4.095 ;
      RECT 45.67 1.865 45.84 2.315 ;
      RECT 45.67 10.145 45.84 10.595 ;
      RECT 45.73 8.365 45.9 10.315 ;
      RECT 45.67 7.305 45.84 8.535 ;
      RECT 45.145 3.895 45.32 5.155 ;
      RECT 45.145 1.865 45.315 5.155 ;
      RECT 45.145 3.365 45.555 3.695 ;
      RECT 45.145 2.525 45.555 2.855 ;
      RECT 45.145 1.865 45.32 2.355 ;
      RECT 45.145 10.105 45.32 10.595 ;
      RECT 45.145 7.305 45.315 10.595 ;
      RECT 45.145 9.605 45.555 9.935 ;
      RECT 45.145 8.765 45.555 9.095 ;
      RECT 45.145 7.305 45.32 8.565 ;
      RECT 42.485 3.27 43.215 3.51 ;
      RECT 43.027 3.065 43.215 3.51 ;
      RECT 42.855 3.077 43.23 3.504 ;
      RECT 42.77 3.092 43.25 3.489 ;
      RECT 42.77 3.107 43.255 3.479 ;
      RECT 42.725 3.127 43.27 3.471 ;
      RECT 42.702 3.162 43.285 3.425 ;
      RECT 42.616 3.185 43.29 3.385 ;
      RECT 42.616 3.203 43.3 3.355 ;
      RECT 42.485 3.272 43.305 3.318 ;
      RECT 42.53 3.215 43.3 3.355 ;
      RECT 42.616 3.167 43.285 3.425 ;
      RECT 42.702 3.136 43.27 3.471 ;
      RECT 42.725 3.117 43.255 3.479 ;
      RECT 42.77 3.09 43.23 3.504 ;
      RECT 42.855 3.072 43.215 3.51 ;
      RECT 42.941 3.066 43.215 3.51 ;
      RECT 43.027 3.061 43.16 3.51 ;
      RECT 43.113 3.056 43.16 3.51 ;
      RECT 42.675 4.67 42.68 4.683 ;
      RECT 42.67 4.565 42.675 4.688 ;
      RECT 42.645 4.425 42.67 4.703 ;
      RECT 42.61 4.376 42.645 4.735 ;
      RECT 42.605 4.344 42.61 4.755 ;
      RECT 42.6 4.335 42.605 4.755 ;
      RECT 42.52 4.3 42.6 4.755 ;
      RECT 42.457 4.27 42.52 4.755 ;
      RECT 42.371 4.258 42.457 4.755 ;
      RECT 42.285 4.244 42.371 4.755 ;
      RECT 42.205 4.231 42.285 4.741 ;
      RECT 42.17 4.223 42.205 4.721 ;
      RECT 42.16 4.22 42.17 4.712 ;
      RECT 42.13 4.215 42.16 4.699 ;
      RECT 42.08 4.19 42.13 4.675 ;
      RECT 42.066 4.164 42.08 4.657 ;
      RECT 41.98 4.124 42.066 4.633 ;
      RECT 41.935 4.072 41.98 4.602 ;
      RECT 41.925 4.047 41.935 4.589 ;
      RECT 41.92 3.828 41.925 3.85 ;
      RECT 41.915 4.03 41.925 4.585 ;
      RECT 41.915 3.826 41.92 3.94 ;
      RECT 41.905 3.822 41.915 4.581 ;
      RECT 41.861 3.82 41.905 4.569 ;
      RECT 41.775 3.82 41.861 4.54 ;
      RECT 41.745 3.82 41.775 4.513 ;
      RECT 41.73 3.82 41.745 4.501 ;
      RECT 41.69 3.832 41.73 4.486 ;
      RECT 41.67 3.851 41.69 4.465 ;
      RECT 41.66 3.861 41.67 4.449 ;
      RECT 41.65 3.867 41.66 4.438 ;
      RECT 41.63 3.877 41.65 4.421 ;
      RECT 41.625 3.886 41.63 4.408 ;
      RECT 41.62 3.89 41.625 4.358 ;
      RECT 41.61 3.896 41.62 4.275 ;
      RECT 41.605 3.9 41.61 4.189 ;
      RECT 41.6 3.92 41.605 4.126 ;
      RECT 41.595 3.943 41.6 4.073 ;
      RECT 41.59 3.961 41.595 4.018 ;
      RECT 42.2 3.78 42.37 4.04 ;
      RECT 42.37 3.745 42.415 4.026 ;
      RECT 42.331 3.747 42.42 4.009 ;
      RECT 42.22 3.764 42.506 3.98 ;
      RECT 42.22 3.779 42.51 3.952 ;
      RECT 42.22 3.76 42.42 4.009 ;
      RECT 42.245 3.748 42.37 4.04 ;
      RECT 42.331 3.746 42.415 4.026 ;
      RECT 41.75 10.045 41.925 10.595 ;
      RECT 41.75 7.305 41.92 10.595 ;
      RECT 41.75 7.305 41.925 8.445 ;
      RECT 41.385 3.135 41.555 3.625 ;
      RECT 41.385 3.135 41.59 3.605 ;
      RECT 41.52 3.055 41.63 3.565 ;
      RECT 41.501 3.059 41.65 3.535 ;
      RECT 41.415 3.067 41.67 3.518 ;
      RECT 41.415 3.073 41.675 3.508 ;
      RECT 41.415 3.082 41.695 3.496 ;
      RECT 41.39 3.107 41.725 3.474 ;
      RECT 41.39 3.127 41.73 3.454 ;
      RECT 41.385 3.14 41.74 3.434 ;
      RECT 41.385 3.207 41.745 3.415 ;
      RECT 41.385 3.34 41.75 3.402 ;
      RECT 41.38 3.145 41.74 3.235 ;
      RECT 41.39 3.102 41.695 3.496 ;
      RECT 41.501 3.057 41.63 3.565 ;
      RECT 41.375 4.81 41.675 5.065 ;
      RECT 41.46 4.776 41.675 5.065 ;
      RECT 41.46 4.779 41.68 4.925 ;
      RECT 41.395 4.8 41.68 4.925 ;
      RECT 41.43 4.79 41.675 5.065 ;
      RECT 41.425 4.795 41.68 4.925 ;
      RECT 41.46 4.774 41.661 5.065 ;
      RECT 41.546 4.765 41.661 5.065 ;
      RECT 41.546 4.759 41.575 5.065 ;
      RECT 41.32 7.305 41.49 9.515 ;
      RECT 41.32 7.305 41.495 8.565 ;
      RECT 41.035 4.4 41.045 4.89 ;
      RECT 40.695 4.335 40.705 4.635 ;
      RECT 41.21 4.507 41.215 4.726 ;
      RECT 41.2 4.487 41.21 4.743 ;
      RECT 41.19 4.467 41.2 4.773 ;
      RECT 41.185 4.457 41.19 4.788 ;
      RECT 41.18 4.453 41.185 4.793 ;
      RECT 41.165 4.445 41.18 4.8 ;
      RECT 41.125 4.425 41.165 4.825 ;
      RECT 41.1 4.407 41.125 4.858 ;
      RECT 41.095 4.405 41.1 4.871 ;
      RECT 41.075 4.402 41.095 4.875 ;
      RECT 41.045 4.4 41.075 4.885 ;
      RECT 40.975 4.402 41.035 4.886 ;
      RECT 40.955 4.402 40.975 4.88 ;
      RECT 40.93 4.4 40.955 4.877 ;
      RECT 40.895 4.395 40.93 4.873 ;
      RECT 40.875 4.389 40.895 4.86 ;
      RECT 40.865 4.386 40.875 4.848 ;
      RECT 40.845 4.383 40.865 4.833 ;
      RECT 40.825 4.379 40.845 4.815 ;
      RECT 40.82 4.376 40.825 4.805 ;
      RECT 40.815 4.375 40.82 4.803 ;
      RECT 40.805 4.372 40.815 4.795 ;
      RECT 40.795 4.366 40.805 4.778 ;
      RECT 40.785 4.36 40.795 4.76 ;
      RECT 40.775 4.354 40.785 4.748 ;
      RECT 40.765 4.348 40.775 4.728 ;
      RECT 40.76 4.344 40.765 4.713 ;
      RECT 40.755 4.342 40.76 4.705 ;
      RECT 40.75 4.34 40.755 4.698 ;
      RECT 40.745 4.338 40.75 4.688 ;
      RECT 40.74 4.336 40.745 4.682 ;
      RECT 40.73 4.335 40.74 4.672 ;
      RECT 40.72 4.335 40.73 4.663 ;
      RECT 40.705 4.335 40.72 4.648 ;
      RECT 40.665 4.335 40.695 4.632 ;
      RECT 40.645 4.337 40.665 4.627 ;
      RECT 40.64 4.342 40.645 4.625 ;
      RECT 40.61 4.35 40.64 4.623 ;
      RECT 40.58 4.365 40.61 4.622 ;
      RECT 40.535 4.387 40.58 4.627 ;
      RECT 40.53 4.402 40.535 4.631 ;
      RECT 40.515 4.407 40.53 4.633 ;
      RECT 40.51 4.411 40.515 4.635 ;
      RECT 40.45 4.434 40.51 4.644 ;
      RECT 40.43 4.46 40.45 4.657 ;
      RECT 40.42 4.467 40.43 4.661 ;
      RECT 40.405 4.474 40.42 4.664 ;
      RECT 40.385 4.484 40.405 4.667 ;
      RECT 40.38 4.492 40.385 4.67 ;
      RECT 40.335 4.497 40.38 4.677 ;
      RECT 40.325 4.5 40.335 4.684 ;
      RECT 40.315 4.5 40.325 4.688 ;
      RECT 40.28 4.502 40.315 4.7 ;
      RECT 40.26 4.505 40.28 4.713 ;
      RECT 40.22 4.508 40.26 4.724 ;
      RECT 40.205 4.51 40.22 4.737 ;
      RECT 40.195 4.51 40.205 4.742 ;
      RECT 40.17 4.511 40.195 4.75 ;
      RECT 40.16 4.513 40.17 4.755 ;
      RECT 40.155 4.514 40.16 4.758 ;
      RECT 40.13 4.512 40.155 4.761 ;
      RECT 40.115 4.51 40.13 4.762 ;
      RECT 40.095 4.507 40.115 4.764 ;
      RECT 40.075 4.502 40.095 4.764 ;
      RECT 40.015 4.497 40.075 4.761 ;
      RECT 39.98 4.472 40.015 4.757 ;
      RECT 39.97 4.449 39.98 4.755 ;
      RECT 39.94 4.426 39.97 4.755 ;
      RECT 39.93 4.405 39.94 4.755 ;
      RECT 39.905 4.387 39.93 4.753 ;
      RECT 39.89 4.365 39.905 4.75 ;
      RECT 39.875 4.347 39.89 4.748 ;
      RECT 39.855 4.337 39.875 4.746 ;
      RECT 39.84 4.332 39.855 4.745 ;
      RECT 39.825 4.33 39.84 4.744 ;
      RECT 39.795 4.331 39.825 4.742 ;
      RECT 39.775 4.334 39.795 4.74 ;
      RECT 39.718 4.338 39.775 4.74 ;
      RECT 39.632 4.347 39.718 4.74 ;
      RECT 39.546 4.358 39.632 4.74 ;
      RECT 39.46 4.369 39.546 4.74 ;
      RECT 39.44 4.376 39.46 4.748 ;
      RECT 39.43 4.379 39.44 4.755 ;
      RECT 39.365 4.384 39.43 4.773 ;
      RECT 39.335 4.391 39.365 4.798 ;
      RECT 39.325 4.394 39.335 4.805 ;
      RECT 39.28 4.398 39.325 4.81 ;
      RECT 39.25 4.403 39.28 4.815 ;
      RECT 39.249 4.405 39.25 4.815 ;
      RECT 39.163 4.411 39.249 4.815 ;
      RECT 39.077 4.422 39.163 4.815 ;
      RECT 38.991 4.434 39.077 4.815 ;
      RECT 38.905 4.445 38.991 4.815 ;
      RECT 38.89 4.452 38.905 4.81 ;
      RECT 38.885 4.454 38.89 4.804 ;
      RECT 38.865 4.465 38.885 4.799 ;
      RECT 38.855 4.483 38.865 4.793 ;
      RECT 38.85 4.495 38.855 4.593 ;
      RECT 41.145 3.248 41.165 3.335 ;
      RECT 41.14 3.183 41.145 3.367 ;
      RECT 41.13 3.15 41.14 3.372 ;
      RECT 41.125 3.13 41.13 3.378 ;
      RECT 41.095 3.13 41.125 3.395 ;
      RECT 41.046 3.13 41.095 3.431 ;
      RECT 40.96 3.13 41.046 3.489 ;
      RECT 40.931 3.14 40.96 3.538 ;
      RECT 40.845 3.182 40.931 3.591 ;
      RECT 40.825 3.22 40.845 3.638 ;
      RECT 40.8 3.237 40.825 3.658 ;
      RECT 40.79 3.251 40.8 3.678 ;
      RECT 40.785 3.257 40.79 3.688 ;
      RECT 40.78 3.261 40.785 3.695 ;
      RECT 40.73 3.281 40.78 3.7 ;
      RECT 40.665 3.325 40.73 3.7 ;
      RECT 40.64 3.375 40.665 3.7 ;
      RECT 40.63 3.405 40.64 3.7 ;
      RECT 40.625 3.432 40.63 3.7 ;
      RECT 40.62 3.45 40.625 3.7 ;
      RECT 40.61 3.492 40.62 3.7 ;
      RECT 40.365 10.105 40.54 10.595 ;
      RECT 40.365 7.305 40.535 10.595 ;
      RECT 40.365 9.605 40.775 9.935 ;
      RECT 40.365 8.765 40.775 9.095 ;
      RECT 40.365 7.305 40.54 8.565 ;
      RECT 40.44 4.85 40.63 5.075 ;
      RECT 40.43 4.851 40.635 5.07 ;
      RECT 40.43 4.853 40.645 5.05 ;
      RECT 40.43 4.857 40.65 5.035 ;
      RECT 40.43 4.844 40.6 5.07 ;
      RECT 40.43 4.847 40.625 5.07 ;
      RECT 40.44 4.843 40.6 5.075 ;
      RECT 40.526 4.841 40.6 5.075 ;
      RECT 40.15 4.092 40.32 4.33 ;
      RECT 40.15 4.092 40.406 4.244 ;
      RECT 40.15 4.092 40.41 4.154 ;
      RECT 40.2 3.865 40.42 4.133 ;
      RECT 40.195 3.882 40.425 4.106 ;
      RECT 40.16 4.04 40.425 4.106 ;
      RECT 40.18 3.89 40.32 4.33 ;
      RECT 40.17 3.972 40.43 4.089 ;
      RECT 40.165 4.02 40.43 4.089 ;
      RECT 40.17 3.93 40.425 4.106 ;
      RECT 40.195 3.867 40.42 4.133 ;
      RECT 39.76 3.842 39.93 4.04 ;
      RECT 39.76 3.842 39.975 4.015 ;
      RECT 39.83 3.785 40 3.973 ;
      RECT 39.805 3.8 40 3.973 ;
      RECT 39.42 3.846 39.45 4.04 ;
      RECT 39.415 3.818 39.42 4.04 ;
      RECT 39.385 3.792 39.415 4.042 ;
      RECT 39.36 3.75 39.385 4.045 ;
      RECT 39.35 3.722 39.36 4.047 ;
      RECT 39.315 3.702 39.35 4.049 ;
      RECT 39.25 3.687 39.315 4.055 ;
      RECT 39.2 3.685 39.25 4.061 ;
      RECT 39.177 3.687 39.2 4.066 ;
      RECT 39.091 3.698 39.177 4.072 ;
      RECT 39.005 3.716 39.091 4.082 ;
      RECT 38.99 3.727 39.005 4.088 ;
      RECT 38.92 3.75 38.99 4.094 ;
      RECT 38.865 3.782 38.92 4.102 ;
      RECT 38.825 3.805 38.865 4.108 ;
      RECT 38.811 3.818 38.825 4.111 ;
      RECT 38.725 3.84 38.811 4.117 ;
      RECT 38.71 3.865 38.725 4.123 ;
      RECT 38.67 3.88 38.71 4.127 ;
      RECT 38.62 3.895 38.67 4.132 ;
      RECT 38.595 3.902 38.62 4.136 ;
      RECT 38.535 3.897 38.595 4.14 ;
      RECT 38.52 3.888 38.535 4.144 ;
      RECT 38.45 3.878 38.52 4.14 ;
      RECT 38.425 3.87 38.445 4.13 ;
      RECT 38.366 3.87 38.425 4.108 ;
      RECT 38.28 3.87 38.366 4.065 ;
      RECT 38.445 3.87 38.45 4.135 ;
      RECT 39.14 3.101 39.31 3.435 ;
      RECT 39.11 3.101 39.31 3.43 ;
      RECT 39.05 3.068 39.11 3.418 ;
      RECT 39.05 3.124 39.32 3.413 ;
      RECT 39.025 3.124 39.32 3.407 ;
      RECT 39.02 3.065 39.05 3.404 ;
      RECT 39.005 3.071 39.14 3.402 ;
      RECT 39 3.079 39.225 3.39 ;
      RECT 39 3.131 39.335 3.343 ;
      RECT 38.985 3.087 39.225 3.338 ;
      RECT 38.985 3.157 39.345 3.279 ;
      RECT 38.955 3.107 39.31 3.24 ;
      RECT 38.955 3.197 39.355 3.236 ;
      RECT 39.005 3.076 39.225 3.402 ;
      RECT 38.345 3.406 38.4 3.67 ;
      RECT 38.345 3.406 38.465 3.669 ;
      RECT 38.345 3.406 38.49 3.668 ;
      RECT 38.345 3.406 38.555 3.667 ;
      RECT 38.49 3.372 38.57 3.666 ;
      RECT 38.305 3.416 38.715 3.665 ;
      RECT 38.345 3.413 38.715 3.665 ;
      RECT 38.305 3.421 38.72 3.658 ;
      RECT 38.29 3.423 38.72 3.657 ;
      RECT 38.29 3.43 38.725 3.653 ;
      RECT 38.27 3.429 38.72 3.649 ;
      RECT 38.27 3.437 38.73 3.648 ;
      RECT 38.265 3.434 38.725 3.644 ;
      RECT 38.265 3.447 38.74 3.643 ;
      RECT 38.25 3.437 38.73 3.642 ;
      RECT 38.215 3.45 38.74 3.635 ;
      RECT 38.4 3.405 38.71 3.665 ;
      RECT 38.4 3.39 38.66 3.665 ;
      RECT 38.465 3.377 38.595 3.665 ;
      RECT 38.01 4.466 38.025 4.859 ;
      RECT 37.975 4.471 38.025 4.858 ;
      RECT 38.01 4.47 38.07 4.857 ;
      RECT 37.955 4.481 38.07 4.856 ;
      RECT 37.97 4.477 38.07 4.856 ;
      RECT 37.935 4.487 38.145 4.853 ;
      RECT 37.935 4.506 38.19 4.851 ;
      RECT 37.935 4.513 38.195 4.848 ;
      RECT 37.92 4.49 38.145 4.845 ;
      RECT 37.9 4.495 38.145 4.838 ;
      RECT 37.895 4.499 38.145 4.834 ;
      RECT 37.895 4.516 38.205 4.833 ;
      RECT 37.875 4.51 38.19 4.829 ;
      RECT 37.875 4.519 38.21 4.823 ;
      RECT 37.87 4.525 38.21 4.595 ;
      RECT 37.935 4.485 38.07 4.853 ;
      RECT 37.81 3.848 38.01 4.16 ;
      RECT 37.885 3.826 38.01 4.16 ;
      RECT 37.825 3.845 38.015 4.145 ;
      RECT 37.795 3.856 38.015 4.143 ;
      RECT 37.81 3.851 38.02 4.109 ;
      RECT 37.795 3.955 38.025 4.076 ;
      RECT 37.825 3.827 38.01 4.16 ;
      RECT 37.885 3.805 37.985 4.16 ;
      RECT 37.91 3.802 37.985 4.16 ;
      RECT 37.91 3.797 37.93 4.16 ;
      RECT 37.315 3.865 37.49 4.04 ;
      RECT 37.31 3.865 37.49 4.038 ;
      RECT 37.285 3.865 37.49 4.033 ;
      RECT 37.23 3.845 37.4 4.023 ;
      RECT 37.23 3.852 37.465 4.023 ;
      RECT 37.315 4.532 37.33 4.715 ;
      RECT 37.305 4.51 37.315 4.715 ;
      RECT 37.29 4.49 37.305 4.715 ;
      RECT 37.28 4.465 37.29 4.715 ;
      RECT 37.25 4.43 37.28 4.715 ;
      RECT 37.215 4.37 37.25 4.715 ;
      RECT 37.21 4.332 37.215 4.715 ;
      RECT 37.16 4.283 37.21 4.715 ;
      RECT 37.15 4.233 37.16 4.703 ;
      RECT 37.135 4.212 37.15 4.663 ;
      RECT 37.115 4.18 37.135 4.613 ;
      RECT 37.09 4.136 37.115 4.553 ;
      RECT 37.085 4.108 37.09 4.508 ;
      RECT 37.08 4.099 37.085 4.494 ;
      RECT 37.075 4.092 37.08 4.481 ;
      RECT 37.07 4.087 37.075 4.47 ;
      RECT 37.065 4.072 37.07 4.46 ;
      RECT 37.06 4.05 37.065 4.447 ;
      RECT 37.05 4.01 37.06 4.422 ;
      RECT 37.025 3.94 37.05 4.378 ;
      RECT 37.02 3.88 37.025 4.343 ;
      RECT 37.005 3.86 37.02 4.31 ;
      RECT 37 3.86 37.005 4.285 ;
      RECT 36.97 3.86 37 4.24 ;
      RECT 36.925 3.86 36.97 4.18 ;
      RECT 36.85 3.86 36.925 4.128 ;
      RECT 36.845 3.86 36.85 4.093 ;
      RECT 36.84 3.86 36.845 4.083 ;
      RECT 36.835 3.86 36.84 4.063 ;
      RECT 37.1 3.08 37.27 3.55 ;
      RECT 37.045 3.073 37.24 3.534 ;
      RECT 37.045 3.087 37.275 3.533 ;
      RECT 37.03 3.088 37.275 3.514 ;
      RECT 37.025 3.106 37.275 3.5 ;
      RECT 37.03 3.089 37.28 3.498 ;
      RECT 37.015 3.12 37.28 3.483 ;
      RECT 37.03 3.095 37.285 3.468 ;
      RECT 37.01 3.135 37.285 3.465 ;
      RECT 37.025 3.107 37.29 3.45 ;
      RECT 37.025 3.119 37.295 3.43 ;
      RECT 37.01 3.135 37.3 3.413 ;
      RECT 37.01 3.145 37.305 3.268 ;
      RECT 37.005 3.145 37.305 3.225 ;
      RECT 37.005 3.16 37.31 3.203 ;
      RECT 37.1 3.07 37.24 3.55 ;
      RECT 37.1 3.068 37.21 3.55 ;
      RECT 37.186 3.065 37.21 3.55 ;
      RECT 36.845 4.732 36.85 4.778 ;
      RECT 36.835 4.58 36.845 4.802 ;
      RECT 36.83 4.425 36.835 4.827 ;
      RECT 36.815 4.387 36.83 4.838 ;
      RECT 36.81 4.37 36.815 4.845 ;
      RECT 36.8 4.358 36.81 4.852 ;
      RECT 36.795 4.349 36.8 4.854 ;
      RECT 36.79 4.347 36.795 4.858 ;
      RECT 36.745 4.338 36.79 4.873 ;
      RECT 36.74 4.33 36.745 4.887 ;
      RECT 36.735 4.327 36.74 4.891 ;
      RECT 36.72 4.322 36.735 4.899 ;
      RECT 36.665 4.312 36.72 4.91 ;
      RECT 36.63 4.3 36.665 4.911 ;
      RECT 36.621 4.295 36.63 4.905 ;
      RECT 36.535 4.295 36.621 4.895 ;
      RECT 36.505 4.295 36.535 4.873 ;
      RECT 36.495 4.295 36.5 4.853 ;
      RECT 36.49 4.295 36.495 4.815 ;
      RECT 36.485 4.295 36.49 4.773 ;
      RECT 36.48 4.295 36.485 4.733 ;
      RECT 36.475 4.295 36.48 4.663 ;
      RECT 36.465 4.295 36.475 4.585 ;
      RECT 36.46 4.295 36.465 4.485 ;
      RECT 36.5 4.295 36.505 4.855 ;
      RECT 35.995 4.377 36.085 4.855 ;
      RECT 35.98 4.38 36.1 4.853 ;
      RECT 35.995 4.379 36.1 4.853 ;
      RECT 35.96 4.386 36.125 4.843 ;
      RECT 35.98 4.38 36.125 4.843 ;
      RECT 35.945 4.392 36.125 4.831 ;
      RECT 35.98 4.383 36.175 4.824 ;
      RECT 35.931 4.4 36.175 4.822 ;
      RECT 35.96 4.39 36.185 4.81 ;
      RECT 35.931 4.411 36.215 4.801 ;
      RECT 35.845 4.435 36.215 4.795 ;
      RECT 35.845 4.448 36.255 4.778 ;
      RECT 35.84 4.47 36.255 4.771 ;
      RECT 35.81 4.485 36.255 4.761 ;
      RECT 35.805 4.496 36.255 4.751 ;
      RECT 35.775 4.509 36.255 4.742 ;
      RECT 35.76 4.527 36.255 4.731 ;
      RECT 35.735 4.54 36.255 4.721 ;
      RECT 35.995 4.376 36.005 4.855 ;
      RECT 36.041 3.8 36.08 4.045 ;
      RECT 35.955 3.8 36.09 4.043 ;
      RECT 35.84 3.825 36.09 4.04 ;
      RECT 35.84 3.825 36.095 4.038 ;
      RECT 35.84 3.825 36.11 4.033 ;
      RECT 35.946 3.8 36.125 4.013 ;
      RECT 35.86 3.808 36.125 4.013 ;
      RECT 35.53 3.16 35.7 3.595 ;
      RECT 35.52 3.194 35.7 3.578 ;
      RECT 35.6 3.13 35.77 3.565 ;
      RECT 35.505 3.205 35.77 3.543 ;
      RECT 35.6 3.14 35.775 3.533 ;
      RECT 35.53 3.192 35.805 3.518 ;
      RECT 35.49 3.218 35.805 3.503 ;
      RECT 35.49 3.26 35.815 3.483 ;
      RECT 35.485 3.285 35.82 3.465 ;
      RECT 35.485 3.295 35.825 3.45 ;
      RECT 35.48 3.232 35.805 3.448 ;
      RECT 35.48 3.305 35.83 3.433 ;
      RECT 35.475 3.242 35.805 3.43 ;
      RECT 35.47 3.326 35.835 3.413 ;
      RECT 35.47 3.358 35.84 3.393 ;
      RECT 35.465 3.272 35.815 3.385 ;
      RECT 35.47 3.257 35.805 3.413 ;
      RECT 35.485 3.227 35.805 3.465 ;
      RECT 35.33 3.814 35.555 4.07 ;
      RECT 35.33 3.847 35.575 4.06 ;
      RECT 35.295 3.847 35.575 4.058 ;
      RECT 35.295 3.86 35.58 4.048 ;
      RECT 35.295 3.88 35.59 4.04 ;
      RECT 35.295 3.977 35.595 4.033 ;
      RECT 35.275 3.725 35.405 4.023 ;
      RECT 35.23 3.88 35.59 3.965 ;
      RECT 35.22 3.725 35.405 3.91 ;
      RECT 35.22 3.757 35.491 3.91 ;
      RECT 35.185 4.287 35.205 4.465 ;
      RECT 35.15 4.24 35.185 4.465 ;
      RECT 35.135 4.18 35.15 4.465 ;
      RECT 35.11 4.127 35.135 4.465 ;
      RECT 35.095 4.08 35.11 4.465 ;
      RECT 35.075 4.057 35.095 4.465 ;
      RECT 35.05 4.022 35.075 4.465 ;
      RECT 35.04 3.868 35.05 4.465 ;
      RECT 35.01 3.863 35.04 4.456 ;
      RECT 35.005 3.86 35.01 4.446 ;
      RECT 34.99 3.86 35.005 4.42 ;
      RECT 34.985 3.86 34.99 4.383 ;
      RECT 34.96 3.86 34.985 4.335 ;
      RECT 34.94 3.86 34.96 4.26 ;
      RECT 34.93 3.86 34.94 4.22 ;
      RECT 34.925 3.86 34.93 4.195 ;
      RECT 34.92 3.86 34.925 4.178 ;
      RECT 34.915 3.86 34.92 4.16 ;
      RECT 34.91 3.861 34.915 4.15 ;
      RECT 34.9 3.863 34.91 4.118 ;
      RECT 34.89 3.865 34.9 4.085 ;
      RECT 34.88 3.868 34.89 4.058 ;
      RECT 35.205 4.295 35.43 4.465 ;
      RECT 34.535 3.107 34.705 3.56 ;
      RECT 34.535 3.107 34.795 3.526 ;
      RECT 34.535 3.107 34.825 3.51 ;
      RECT 34.535 3.107 34.855 3.483 ;
      RECT 34.791 3.085 34.87 3.465 ;
      RECT 34.57 3.092 34.875 3.45 ;
      RECT 34.57 3.1 34.885 3.413 ;
      RECT 34.53 3.127 34.885 3.385 ;
      RECT 34.515 3.14 34.885 3.35 ;
      RECT 34.535 3.115 34.905 3.34 ;
      RECT 34.51 3.18 34.905 3.31 ;
      RECT 34.51 3.21 34.91 3.293 ;
      RECT 34.505 3.24 34.91 3.28 ;
      RECT 34.57 3.089 34.87 3.465 ;
      RECT 34.705 3.086 34.791 3.544 ;
      RECT 34.656 3.087 34.87 3.465 ;
      RECT 34.8 4.747 34.845 4.94 ;
      RECT 34.79 4.717 34.8 4.94 ;
      RECT 34.785 4.702 34.79 4.94 ;
      RECT 34.745 4.612 34.785 4.94 ;
      RECT 34.74 4.525 34.745 4.94 ;
      RECT 34.73 4.495 34.74 4.94 ;
      RECT 34.725 4.455 34.73 4.94 ;
      RECT 34.715 4.417 34.725 4.94 ;
      RECT 34.71 4.382 34.715 4.94 ;
      RECT 34.69 4.335 34.71 4.94 ;
      RECT 34.675 4.26 34.69 4.94 ;
      RECT 34.67 4.215 34.675 4.935 ;
      RECT 34.665 4.195 34.67 4.908 ;
      RECT 34.66 4.175 34.665 4.893 ;
      RECT 34.655 4.15 34.66 4.873 ;
      RECT 34.65 4.128 34.655 4.858 ;
      RECT 34.645 4.106 34.65 4.84 ;
      RECT 34.64 4.085 34.645 4.83 ;
      RECT 34.63 4.057 34.64 4.8 ;
      RECT 34.62 4.02 34.63 4.768 ;
      RECT 34.61 3.98 34.62 4.735 ;
      RECT 34.6 3.958 34.61 4.705 ;
      RECT 34.57 3.91 34.6 4.637 ;
      RECT 34.555 3.87 34.57 4.564 ;
      RECT 34.545 3.87 34.555 4.53 ;
      RECT 34.54 3.87 34.545 4.505 ;
      RECT 34.535 3.87 34.54 4.49 ;
      RECT 34.53 3.87 34.535 4.468 ;
      RECT 34.525 3.87 34.53 4.455 ;
      RECT 34.51 3.87 34.525 4.42 ;
      RECT 34.49 3.87 34.51 4.36 ;
      RECT 34.48 3.87 34.49 4.31 ;
      RECT 34.46 3.87 34.48 4.258 ;
      RECT 34.44 3.87 34.46 4.215 ;
      RECT 34.43 3.87 34.44 4.203 ;
      RECT 34.4 3.87 34.43 4.19 ;
      RECT 34.37 3.891 34.4 4.17 ;
      RECT 34.36 3.919 34.37 4.15 ;
      RECT 34.345 3.936 34.36 4.118 ;
      RECT 34.34 3.95 34.345 4.085 ;
      RECT 34.335 3.958 34.34 4.058 ;
      RECT 34.33 3.966 34.335 4.02 ;
      RECT 34.335 4.49 34.34 4.825 ;
      RECT 34.3 4.477 34.335 4.824 ;
      RECT 34.23 4.417 34.3 4.823 ;
      RECT 34.15 4.36 34.23 4.822 ;
      RECT 34.015 4.32 34.15 4.821 ;
      RECT 34.015 4.507 34.35 4.81 ;
      RECT 33.975 4.507 34.35 4.8 ;
      RECT 33.975 4.525 34.355 4.795 ;
      RECT 33.975 4.615 34.36 4.785 ;
      RECT 33.97 4.31 34.135 4.765 ;
      RECT 33.965 4.31 34.135 4.508 ;
      RECT 33.965 4.467 34.33 4.508 ;
      RECT 33.965 4.455 34.325 4.508 ;
      RECT 33.1 7.305 33.27 8.775 ;
      RECT 33.1 7.305 33.275 8.565 ;
      RECT 32.73 9.255 33.2 9.425 ;
      RECT 32.73 8.235 32.9 9.425 ;
      RECT 32.725 3.035 32.895 4.225 ;
      RECT 32.725 3.035 33.195 3.205 ;
      RECT 32.11 3.895 32.285 5.155 ;
      RECT 32.11 3.685 32.28 5.155 ;
      RECT 32.11 7.305 32.28 8.775 ;
      RECT 32.11 7.305 32.285 8.565 ;
      RECT 31.74 3.035 31.91 4.225 ;
      RECT 31.74 3.035 32.21 3.205 ;
      RECT 31.74 9.255 32.21 9.425 ;
      RECT 31.74 8.235 31.91 9.425 ;
      RECT 30.75 4.015 30.925 5.155 ;
      RECT 30.75 1.865 30.92 5.155 ;
      RECT 30.75 1.865 30.925 2.415 ;
      RECT 30.75 10.045 30.925 10.595 ;
      RECT 30.75 7.305 30.92 10.595 ;
      RECT 30.75 7.305 30.925 8.445 ;
      RECT 30.32 3.895 30.495 5.155 ;
      RECT 30.32 2.945 30.49 5.155 ;
      RECT 30.32 7.305 30.49 9.515 ;
      RECT 30.32 7.305 30.495 8.565 ;
      RECT 29.89 3.925 30.06 5.155 ;
      RECT 29.95 2.145 30.12 4.095 ;
      RECT 29.89 1.865 30.06 2.315 ;
      RECT 29.89 10.145 30.06 10.595 ;
      RECT 29.95 8.365 30.12 10.315 ;
      RECT 29.89 7.305 30.06 8.535 ;
      RECT 29.365 3.895 29.54 5.155 ;
      RECT 29.365 1.865 29.535 5.155 ;
      RECT 29.365 3.365 29.775 3.695 ;
      RECT 29.365 2.525 29.775 2.855 ;
      RECT 29.365 1.865 29.54 2.355 ;
      RECT 29.365 10.105 29.54 10.595 ;
      RECT 29.365 7.305 29.535 10.595 ;
      RECT 29.365 9.605 29.775 9.935 ;
      RECT 29.365 8.765 29.775 9.095 ;
      RECT 29.365 7.305 29.54 8.565 ;
      RECT 26.705 3.27 27.435 3.51 ;
      RECT 27.247 3.065 27.435 3.51 ;
      RECT 27.075 3.077 27.45 3.504 ;
      RECT 26.99 3.092 27.47 3.489 ;
      RECT 26.99 3.107 27.475 3.479 ;
      RECT 26.945 3.127 27.49 3.471 ;
      RECT 26.922 3.162 27.505 3.425 ;
      RECT 26.836 3.185 27.51 3.385 ;
      RECT 26.836 3.203 27.52 3.355 ;
      RECT 26.705 3.272 27.525 3.318 ;
      RECT 26.75 3.215 27.52 3.355 ;
      RECT 26.836 3.167 27.505 3.425 ;
      RECT 26.922 3.136 27.49 3.471 ;
      RECT 26.945 3.117 27.475 3.479 ;
      RECT 26.99 3.09 27.45 3.504 ;
      RECT 27.075 3.072 27.435 3.51 ;
      RECT 27.161 3.066 27.435 3.51 ;
      RECT 27.247 3.061 27.38 3.51 ;
      RECT 27.333 3.056 27.38 3.51 ;
      RECT 26.895 4.67 26.9 4.683 ;
      RECT 26.89 4.565 26.895 4.688 ;
      RECT 26.865 4.425 26.89 4.703 ;
      RECT 26.83 4.376 26.865 4.735 ;
      RECT 26.825 4.344 26.83 4.755 ;
      RECT 26.82 4.335 26.825 4.755 ;
      RECT 26.74 4.3 26.82 4.755 ;
      RECT 26.677 4.27 26.74 4.755 ;
      RECT 26.591 4.258 26.677 4.755 ;
      RECT 26.505 4.244 26.591 4.755 ;
      RECT 26.425 4.231 26.505 4.741 ;
      RECT 26.39 4.223 26.425 4.721 ;
      RECT 26.38 4.22 26.39 4.712 ;
      RECT 26.35 4.215 26.38 4.699 ;
      RECT 26.3 4.19 26.35 4.675 ;
      RECT 26.286 4.164 26.3 4.657 ;
      RECT 26.2 4.124 26.286 4.633 ;
      RECT 26.155 4.072 26.2 4.602 ;
      RECT 26.145 4.047 26.155 4.589 ;
      RECT 26.14 3.828 26.145 3.85 ;
      RECT 26.135 4.03 26.145 4.585 ;
      RECT 26.135 3.826 26.14 3.94 ;
      RECT 26.125 3.822 26.135 4.581 ;
      RECT 26.081 3.82 26.125 4.569 ;
      RECT 25.995 3.82 26.081 4.54 ;
      RECT 25.965 3.82 25.995 4.513 ;
      RECT 25.95 3.82 25.965 4.501 ;
      RECT 25.91 3.832 25.95 4.486 ;
      RECT 25.89 3.851 25.91 4.465 ;
      RECT 25.88 3.861 25.89 4.449 ;
      RECT 25.87 3.867 25.88 4.438 ;
      RECT 25.85 3.877 25.87 4.421 ;
      RECT 25.845 3.886 25.85 4.408 ;
      RECT 25.84 3.89 25.845 4.358 ;
      RECT 25.83 3.896 25.84 4.275 ;
      RECT 25.825 3.9 25.83 4.189 ;
      RECT 25.82 3.92 25.825 4.126 ;
      RECT 25.815 3.943 25.82 4.073 ;
      RECT 25.81 3.961 25.815 4.018 ;
      RECT 26.42 3.78 26.59 4.04 ;
      RECT 26.59 3.745 26.635 4.026 ;
      RECT 26.551 3.747 26.64 4.009 ;
      RECT 26.44 3.764 26.726 3.98 ;
      RECT 26.44 3.779 26.73 3.952 ;
      RECT 26.44 3.76 26.64 4.009 ;
      RECT 26.465 3.748 26.59 4.04 ;
      RECT 26.551 3.746 26.635 4.026 ;
      RECT 25.97 10.045 26.145 10.595 ;
      RECT 25.97 7.305 26.14 10.595 ;
      RECT 25.97 7.305 26.145 8.445 ;
      RECT 25.605 3.135 25.775 3.625 ;
      RECT 25.605 3.135 25.81 3.605 ;
      RECT 25.74 3.055 25.85 3.565 ;
      RECT 25.721 3.059 25.87 3.535 ;
      RECT 25.635 3.067 25.89 3.518 ;
      RECT 25.635 3.073 25.895 3.508 ;
      RECT 25.635 3.082 25.915 3.496 ;
      RECT 25.61 3.107 25.945 3.474 ;
      RECT 25.61 3.127 25.95 3.454 ;
      RECT 25.605 3.14 25.96 3.434 ;
      RECT 25.605 3.207 25.965 3.415 ;
      RECT 25.605 3.34 25.97 3.402 ;
      RECT 25.6 3.145 25.96 3.235 ;
      RECT 25.61 3.102 25.915 3.496 ;
      RECT 25.721 3.057 25.85 3.565 ;
      RECT 25.595 4.81 25.895 5.065 ;
      RECT 25.68 4.776 25.895 5.065 ;
      RECT 25.68 4.779 25.9 4.925 ;
      RECT 25.615 4.8 25.9 4.925 ;
      RECT 25.65 4.79 25.895 5.065 ;
      RECT 25.645 4.795 25.9 4.925 ;
      RECT 25.68 4.774 25.881 5.065 ;
      RECT 25.766 4.765 25.881 5.065 ;
      RECT 25.766 4.759 25.795 5.065 ;
      RECT 25.54 7.305 25.71 9.515 ;
      RECT 25.54 7.305 25.715 8.565 ;
      RECT 25.255 4.4 25.265 4.89 ;
      RECT 24.915 4.335 24.925 4.635 ;
      RECT 25.43 4.507 25.435 4.726 ;
      RECT 25.42 4.487 25.43 4.743 ;
      RECT 25.41 4.467 25.42 4.773 ;
      RECT 25.405 4.457 25.41 4.788 ;
      RECT 25.4 4.453 25.405 4.793 ;
      RECT 25.385 4.445 25.4 4.8 ;
      RECT 25.345 4.425 25.385 4.825 ;
      RECT 25.32 4.407 25.345 4.858 ;
      RECT 25.315 4.405 25.32 4.871 ;
      RECT 25.295 4.402 25.315 4.875 ;
      RECT 25.265 4.4 25.295 4.885 ;
      RECT 25.195 4.402 25.255 4.886 ;
      RECT 25.175 4.402 25.195 4.88 ;
      RECT 25.15 4.4 25.175 4.877 ;
      RECT 25.115 4.395 25.15 4.873 ;
      RECT 25.095 4.389 25.115 4.86 ;
      RECT 25.085 4.386 25.095 4.848 ;
      RECT 25.065 4.383 25.085 4.833 ;
      RECT 25.045 4.379 25.065 4.815 ;
      RECT 25.04 4.376 25.045 4.805 ;
      RECT 25.035 4.375 25.04 4.803 ;
      RECT 25.025 4.372 25.035 4.795 ;
      RECT 25.015 4.366 25.025 4.778 ;
      RECT 25.005 4.36 25.015 4.76 ;
      RECT 24.995 4.354 25.005 4.748 ;
      RECT 24.985 4.348 24.995 4.728 ;
      RECT 24.98 4.344 24.985 4.713 ;
      RECT 24.975 4.342 24.98 4.705 ;
      RECT 24.97 4.34 24.975 4.698 ;
      RECT 24.965 4.338 24.97 4.688 ;
      RECT 24.96 4.336 24.965 4.682 ;
      RECT 24.95 4.335 24.96 4.672 ;
      RECT 24.94 4.335 24.95 4.663 ;
      RECT 24.925 4.335 24.94 4.648 ;
      RECT 24.885 4.335 24.915 4.632 ;
      RECT 24.865 4.337 24.885 4.627 ;
      RECT 24.86 4.342 24.865 4.625 ;
      RECT 24.83 4.35 24.86 4.623 ;
      RECT 24.8 4.365 24.83 4.622 ;
      RECT 24.755 4.387 24.8 4.627 ;
      RECT 24.75 4.402 24.755 4.631 ;
      RECT 24.735 4.407 24.75 4.633 ;
      RECT 24.73 4.411 24.735 4.635 ;
      RECT 24.67 4.434 24.73 4.644 ;
      RECT 24.65 4.46 24.67 4.657 ;
      RECT 24.64 4.467 24.65 4.661 ;
      RECT 24.625 4.474 24.64 4.664 ;
      RECT 24.605 4.484 24.625 4.667 ;
      RECT 24.6 4.492 24.605 4.67 ;
      RECT 24.555 4.497 24.6 4.677 ;
      RECT 24.545 4.5 24.555 4.684 ;
      RECT 24.535 4.5 24.545 4.688 ;
      RECT 24.5 4.502 24.535 4.7 ;
      RECT 24.48 4.505 24.5 4.713 ;
      RECT 24.44 4.508 24.48 4.724 ;
      RECT 24.425 4.51 24.44 4.737 ;
      RECT 24.415 4.51 24.425 4.742 ;
      RECT 24.39 4.511 24.415 4.75 ;
      RECT 24.38 4.513 24.39 4.755 ;
      RECT 24.375 4.514 24.38 4.758 ;
      RECT 24.35 4.512 24.375 4.761 ;
      RECT 24.335 4.51 24.35 4.762 ;
      RECT 24.315 4.507 24.335 4.764 ;
      RECT 24.295 4.502 24.315 4.764 ;
      RECT 24.235 4.497 24.295 4.761 ;
      RECT 24.2 4.472 24.235 4.757 ;
      RECT 24.19 4.449 24.2 4.755 ;
      RECT 24.16 4.426 24.19 4.755 ;
      RECT 24.15 4.405 24.16 4.755 ;
      RECT 24.125 4.387 24.15 4.753 ;
      RECT 24.11 4.365 24.125 4.75 ;
      RECT 24.095 4.347 24.11 4.748 ;
      RECT 24.075 4.337 24.095 4.746 ;
      RECT 24.06 4.332 24.075 4.745 ;
      RECT 24.045 4.33 24.06 4.744 ;
      RECT 24.015 4.331 24.045 4.742 ;
      RECT 23.995 4.334 24.015 4.74 ;
      RECT 23.938 4.338 23.995 4.74 ;
      RECT 23.852 4.347 23.938 4.74 ;
      RECT 23.766 4.358 23.852 4.74 ;
      RECT 23.68 4.369 23.766 4.74 ;
      RECT 23.66 4.376 23.68 4.748 ;
      RECT 23.65 4.379 23.66 4.755 ;
      RECT 23.585 4.384 23.65 4.773 ;
      RECT 23.555 4.391 23.585 4.798 ;
      RECT 23.545 4.394 23.555 4.805 ;
      RECT 23.5 4.398 23.545 4.81 ;
      RECT 23.47 4.403 23.5 4.815 ;
      RECT 23.469 4.405 23.47 4.815 ;
      RECT 23.383 4.411 23.469 4.815 ;
      RECT 23.297 4.422 23.383 4.815 ;
      RECT 23.211 4.434 23.297 4.815 ;
      RECT 23.125 4.445 23.211 4.815 ;
      RECT 23.11 4.452 23.125 4.81 ;
      RECT 23.105 4.454 23.11 4.804 ;
      RECT 23.085 4.465 23.105 4.799 ;
      RECT 23.075 4.483 23.085 4.793 ;
      RECT 23.07 4.495 23.075 4.593 ;
      RECT 25.365 3.248 25.385 3.335 ;
      RECT 25.36 3.183 25.365 3.367 ;
      RECT 25.35 3.15 25.36 3.372 ;
      RECT 25.345 3.13 25.35 3.378 ;
      RECT 25.315 3.13 25.345 3.395 ;
      RECT 25.266 3.13 25.315 3.431 ;
      RECT 25.18 3.13 25.266 3.489 ;
      RECT 25.151 3.14 25.18 3.538 ;
      RECT 25.065 3.182 25.151 3.591 ;
      RECT 25.045 3.22 25.065 3.638 ;
      RECT 25.02 3.237 25.045 3.658 ;
      RECT 25.01 3.251 25.02 3.678 ;
      RECT 25.005 3.257 25.01 3.688 ;
      RECT 25 3.261 25.005 3.695 ;
      RECT 24.95 3.281 25 3.7 ;
      RECT 24.885 3.325 24.95 3.7 ;
      RECT 24.86 3.375 24.885 3.7 ;
      RECT 24.85 3.405 24.86 3.7 ;
      RECT 24.845 3.432 24.85 3.7 ;
      RECT 24.84 3.45 24.845 3.7 ;
      RECT 24.83 3.492 24.84 3.7 ;
      RECT 24.585 10.105 24.76 10.595 ;
      RECT 24.585 7.305 24.755 10.595 ;
      RECT 24.585 9.605 24.995 9.935 ;
      RECT 24.585 8.765 24.995 9.095 ;
      RECT 24.585 7.305 24.76 8.565 ;
      RECT 24.66 4.85 24.85 5.075 ;
      RECT 24.65 4.851 24.855 5.07 ;
      RECT 24.65 4.853 24.865 5.05 ;
      RECT 24.65 4.857 24.87 5.035 ;
      RECT 24.65 4.844 24.82 5.07 ;
      RECT 24.65 4.847 24.845 5.07 ;
      RECT 24.66 4.843 24.82 5.075 ;
      RECT 24.746 4.841 24.82 5.075 ;
      RECT 24.37 4.092 24.54 4.33 ;
      RECT 24.37 4.092 24.626 4.244 ;
      RECT 24.37 4.092 24.63 4.154 ;
      RECT 24.42 3.865 24.64 4.133 ;
      RECT 24.415 3.882 24.645 4.106 ;
      RECT 24.38 4.04 24.645 4.106 ;
      RECT 24.4 3.89 24.54 4.33 ;
      RECT 24.39 3.972 24.65 4.089 ;
      RECT 24.385 4.02 24.65 4.089 ;
      RECT 24.39 3.93 24.645 4.106 ;
      RECT 24.415 3.867 24.64 4.133 ;
      RECT 23.98 3.842 24.15 4.04 ;
      RECT 23.98 3.842 24.195 4.015 ;
      RECT 24.05 3.785 24.22 3.973 ;
      RECT 24.025 3.8 24.22 3.973 ;
      RECT 23.64 3.846 23.67 4.04 ;
      RECT 23.635 3.818 23.64 4.04 ;
      RECT 23.605 3.792 23.635 4.042 ;
      RECT 23.58 3.75 23.605 4.045 ;
      RECT 23.57 3.722 23.58 4.047 ;
      RECT 23.535 3.702 23.57 4.049 ;
      RECT 23.47 3.687 23.535 4.055 ;
      RECT 23.42 3.685 23.47 4.061 ;
      RECT 23.397 3.687 23.42 4.066 ;
      RECT 23.311 3.698 23.397 4.072 ;
      RECT 23.225 3.716 23.311 4.082 ;
      RECT 23.21 3.727 23.225 4.088 ;
      RECT 23.14 3.75 23.21 4.094 ;
      RECT 23.085 3.782 23.14 4.102 ;
      RECT 23.045 3.805 23.085 4.108 ;
      RECT 23.031 3.818 23.045 4.111 ;
      RECT 22.945 3.84 23.031 4.117 ;
      RECT 22.93 3.865 22.945 4.123 ;
      RECT 22.89 3.88 22.93 4.127 ;
      RECT 22.84 3.895 22.89 4.132 ;
      RECT 22.815 3.902 22.84 4.136 ;
      RECT 22.755 3.897 22.815 4.14 ;
      RECT 22.74 3.888 22.755 4.144 ;
      RECT 22.67 3.878 22.74 4.14 ;
      RECT 22.645 3.87 22.665 4.13 ;
      RECT 22.586 3.87 22.645 4.108 ;
      RECT 22.5 3.87 22.586 4.065 ;
      RECT 22.665 3.87 22.67 4.135 ;
      RECT 23.36 3.101 23.53 3.435 ;
      RECT 23.33 3.101 23.53 3.43 ;
      RECT 23.27 3.068 23.33 3.418 ;
      RECT 23.27 3.124 23.54 3.413 ;
      RECT 23.245 3.124 23.54 3.407 ;
      RECT 23.24 3.065 23.27 3.404 ;
      RECT 23.225 3.071 23.36 3.402 ;
      RECT 23.22 3.079 23.445 3.39 ;
      RECT 23.22 3.131 23.555 3.343 ;
      RECT 23.205 3.087 23.445 3.338 ;
      RECT 23.205 3.157 23.565 3.279 ;
      RECT 23.175 3.107 23.53 3.24 ;
      RECT 23.175 3.197 23.575 3.236 ;
      RECT 23.225 3.076 23.445 3.402 ;
      RECT 22.565 3.406 22.62 3.67 ;
      RECT 22.565 3.406 22.685 3.669 ;
      RECT 22.565 3.406 22.71 3.668 ;
      RECT 22.565 3.406 22.775 3.667 ;
      RECT 22.71 3.372 22.79 3.666 ;
      RECT 22.525 3.416 22.935 3.665 ;
      RECT 22.565 3.413 22.935 3.665 ;
      RECT 22.525 3.421 22.94 3.658 ;
      RECT 22.51 3.423 22.94 3.657 ;
      RECT 22.51 3.43 22.945 3.653 ;
      RECT 22.49 3.429 22.94 3.649 ;
      RECT 22.49 3.437 22.95 3.648 ;
      RECT 22.485 3.434 22.945 3.644 ;
      RECT 22.485 3.447 22.96 3.643 ;
      RECT 22.47 3.437 22.95 3.642 ;
      RECT 22.435 3.45 22.96 3.635 ;
      RECT 22.62 3.405 22.93 3.665 ;
      RECT 22.62 3.39 22.88 3.665 ;
      RECT 22.685 3.377 22.815 3.665 ;
      RECT 22.23 4.466 22.245 4.859 ;
      RECT 22.195 4.471 22.245 4.858 ;
      RECT 22.23 4.47 22.29 4.857 ;
      RECT 22.175 4.481 22.29 4.856 ;
      RECT 22.19 4.477 22.29 4.856 ;
      RECT 22.155 4.487 22.365 4.853 ;
      RECT 22.155 4.506 22.41 4.851 ;
      RECT 22.155 4.513 22.415 4.848 ;
      RECT 22.14 4.49 22.365 4.845 ;
      RECT 22.12 4.495 22.365 4.838 ;
      RECT 22.115 4.499 22.365 4.834 ;
      RECT 22.115 4.516 22.425 4.833 ;
      RECT 22.095 4.51 22.41 4.829 ;
      RECT 22.095 4.519 22.43 4.823 ;
      RECT 22.09 4.525 22.43 4.595 ;
      RECT 22.155 4.485 22.29 4.853 ;
      RECT 22.03 3.848 22.23 4.16 ;
      RECT 22.105 3.826 22.23 4.16 ;
      RECT 22.045 3.845 22.235 4.145 ;
      RECT 22.015 3.856 22.235 4.143 ;
      RECT 22.03 3.851 22.24 4.109 ;
      RECT 22.015 3.955 22.245 4.076 ;
      RECT 22.045 3.827 22.23 4.16 ;
      RECT 22.105 3.805 22.205 4.16 ;
      RECT 22.13 3.802 22.205 4.16 ;
      RECT 22.13 3.797 22.15 4.16 ;
      RECT 21.535 3.865 21.71 4.04 ;
      RECT 21.53 3.865 21.71 4.038 ;
      RECT 21.505 3.865 21.71 4.033 ;
      RECT 21.45 3.845 21.62 4.023 ;
      RECT 21.45 3.852 21.685 4.023 ;
      RECT 21.535 4.532 21.55 4.715 ;
      RECT 21.525 4.51 21.535 4.715 ;
      RECT 21.51 4.49 21.525 4.715 ;
      RECT 21.5 4.465 21.51 4.715 ;
      RECT 21.47 4.43 21.5 4.715 ;
      RECT 21.435 4.37 21.47 4.715 ;
      RECT 21.43 4.332 21.435 4.715 ;
      RECT 21.38 4.283 21.43 4.715 ;
      RECT 21.37 4.233 21.38 4.703 ;
      RECT 21.355 4.212 21.37 4.663 ;
      RECT 21.335 4.18 21.355 4.613 ;
      RECT 21.31 4.136 21.335 4.553 ;
      RECT 21.305 4.108 21.31 4.508 ;
      RECT 21.3 4.099 21.305 4.494 ;
      RECT 21.295 4.092 21.3 4.481 ;
      RECT 21.29 4.087 21.295 4.47 ;
      RECT 21.285 4.072 21.29 4.46 ;
      RECT 21.28 4.05 21.285 4.447 ;
      RECT 21.27 4.01 21.28 4.422 ;
      RECT 21.245 3.94 21.27 4.378 ;
      RECT 21.24 3.88 21.245 4.343 ;
      RECT 21.225 3.86 21.24 4.31 ;
      RECT 21.22 3.86 21.225 4.285 ;
      RECT 21.19 3.86 21.22 4.24 ;
      RECT 21.145 3.86 21.19 4.18 ;
      RECT 21.07 3.86 21.145 4.128 ;
      RECT 21.065 3.86 21.07 4.093 ;
      RECT 21.06 3.86 21.065 4.083 ;
      RECT 21.055 3.86 21.06 4.063 ;
      RECT 21.32 3.08 21.49 3.55 ;
      RECT 21.265 3.073 21.46 3.534 ;
      RECT 21.265 3.087 21.495 3.533 ;
      RECT 21.25 3.088 21.495 3.514 ;
      RECT 21.245 3.106 21.495 3.5 ;
      RECT 21.25 3.089 21.5 3.498 ;
      RECT 21.235 3.12 21.5 3.483 ;
      RECT 21.25 3.095 21.505 3.468 ;
      RECT 21.23 3.135 21.505 3.465 ;
      RECT 21.245 3.107 21.51 3.45 ;
      RECT 21.245 3.119 21.515 3.43 ;
      RECT 21.23 3.135 21.52 3.413 ;
      RECT 21.23 3.145 21.525 3.268 ;
      RECT 21.225 3.145 21.525 3.225 ;
      RECT 21.225 3.16 21.53 3.203 ;
      RECT 21.32 3.07 21.46 3.55 ;
      RECT 21.32 3.068 21.43 3.55 ;
      RECT 21.406 3.065 21.43 3.55 ;
      RECT 21.065 4.732 21.07 4.778 ;
      RECT 21.055 4.58 21.065 4.802 ;
      RECT 21.05 4.425 21.055 4.827 ;
      RECT 21.035 4.387 21.05 4.838 ;
      RECT 21.03 4.37 21.035 4.845 ;
      RECT 21.02 4.358 21.03 4.852 ;
      RECT 21.015 4.349 21.02 4.854 ;
      RECT 21.01 4.347 21.015 4.858 ;
      RECT 20.965 4.338 21.01 4.873 ;
      RECT 20.96 4.33 20.965 4.887 ;
      RECT 20.955 4.327 20.96 4.891 ;
      RECT 20.94 4.322 20.955 4.899 ;
      RECT 20.885 4.312 20.94 4.91 ;
      RECT 20.85 4.3 20.885 4.911 ;
      RECT 20.841 4.295 20.85 4.905 ;
      RECT 20.755 4.295 20.841 4.895 ;
      RECT 20.725 4.295 20.755 4.873 ;
      RECT 20.715 4.295 20.72 4.853 ;
      RECT 20.71 4.295 20.715 4.815 ;
      RECT 20.705 4.295 20.71 4.773 ;
      RECT 20.7 4.295 20.705 4.733 ;
      RECT 20.695 4.295 20.7 4.663 ;
      RECT 20.685 4.295 20.695 4.585 ;
      RECT 20.68 4.295 20.685 4.485 ;
      RECT 20.72 4.295 20.725 4.855 ;
      RECT 20.215 4.377 20.305 4.855 ;
      RECT 20.2 4.38 20.32 4.853 ;
      RECT 20.215 4.379 20.32 4.853 ;
      RECT 20.18 4.386 20.345 4.843 ;
      RECT 20.2 4.38 20.345 4.843 ;
      RECT 20.165 4.392 20.345 4.831 ;
      RECT 20.2 4.383 20.395 4.824 ;
      RECT 20.151 4.4 20.395 4.822 ;
      RECT 20.18 4.39 20.405 4.81 ;
      RECT 20.151 4.411 20.435 4.801 ;
      RECT 20.065 4.435 20.435 4.795 ;
      RECT 20.065 4.448 20.475 4.778 ;
      RECT 20.06 4.47 20.475 4.771 ;
      RECT 20.03 4.485 20.475 4.761 ;
      RECT 20.025 4.496 20.475 4.751 ;
      RECT 19.995 4.509 20.475 4.742 ;
      RECT 19.98 4.527 20.475 4.731 ;
      RECT 19.955 4.54 20.475 4.721 ;
      RECT 20.215 4.376 20.225 4.855 ;
      RECT 20.261 3.8 20.3 4.045 ;
      RECT 20.175 3.8 20.31 4.043 ;
      RECT 20.06 3.825 20.31 4.04 ;
      RECT 20.06 3.825 20.315 4.038 ;
      RECT 20.06 3.825 20.33 4.033 ;
      RECT 20.166 3.8 20.345 4.013 ;
      RECT 20.08 3.808 20.345 4.013 ;
      RECT 19.75 3.16 19.92 3.595 ;
      RECT 19.74 3.194 19.92 3.578 ;
      RECT 19.82 3.13 19.99 3.565 ;
      RECT 19.725 3.205 19.99 3.543 ;
      RECT 19.82 3.14 19.995 3.533 ;
      RECT 19.75 3.192 20.025 3.518 ;
      RECT 19.71 3.218 20.025 3.503 ;
      RECT 19.71 3.26 20.035 3.483 ;
      RECT 19.705 3.285 20.04 3.465 ;
      RECT 19.705 3.295 20.045 3.45 ;
      RECT 19.7 3.232 20.025 3.448 ;
      RECT 19.7 3.305 20.05 3.433 ;
      RECT 19.695 3.242 20.025 3.43 ;
      RECT 19.69 3.326 20.055 3.413 ;
      RECT 19.69 3.358 20.06 3.393 ;
      RECT 19.685 3.272 20.035 3.385 ;
      RECT 19.69 3.257 20.025 3.413 ;
      RECT 19.705 3.227 20.025 3.465 ;
      RECT 19.55 3.814 19.775 4.07 ;
      RECT 19.55 3.847 19.795 4.06 ;
      RECT 19.515 3.847 19.795 4.058 ;
      RECT 19.515 3.86 19.8 4.048 ;
      RECT 19.515 3.88 19.81 4.04 ;
      RECT 19.515 3.977 19.815 4.033 ;
      RECT 19.495 3.725 19.625 4.023 ;
      RECT 19.45 3.88 19.81 3.965 ;
      RECT 19.44 3.725 19.625 3.91 ;
      RECT 19.44 3.757 19.711 3.91 ;
      RECT 19.405 4.287 19.425 4.465 ;
      RECT 19.37 4.24 19.405 4.465 ;
      RECT 19.355 4.18 19.37 4.465 ;
      RECT 19.33 4.127 19.355 4.465 ;
      RECT 19.315 4.08 19.33 4.465 ;
      RECT 19.295 4.057 19.315 4.465 ;
      RECT 19.27 4.022 19.295 4.465 ;
      RECT 19.26 3.868 19.27 4.465 ;
      RECT 19.23 3.863 19.26 4.456 ;
      RECT 19.225 3.86 19.23 4.446 ;
      RECT 19.21 3.86 19.225 4.42 ;
      RECT 19.205 3.86 19.21 4.383 ;
      RECT 19.18 3.86 19.205 4.335 ;
      RECT 19.16 3.86 19.18 4.26 ;
      RECT 19.15 3.86 19.16 4.22 ;
      RECT 19.145 3.86 19.15 4.195 ;
      RECT 19.14 3.86 19.145 4.178 ;
      RECT 19.135 3.86 19.14 4.16 ;
      RECT 19.13 3.861 19.135 4.15 ;
      RECT 19.12 3.863 19.13 4.118 ;
      RECT 19.11 3.865 19.12 4.085 ;
      RECT 19.1 3.868 19.11 4.058 ;
      RECT 19.425 4.295 19.65 4.465 ;
      RECT 18.755 3.107 18.925 3.56 ;
      RECT 18.755 3.107 19.015 3.526 ;
      RECT 18.755 3.107 19.045 3.51 ;
      RECT 18.755 3.107 19.075 3.483 ;
      RECT 19.011 3.085 19.09 3.465 ;
      RECT 18.79 3.092 19.095 3.45 ;
      RECT 18.79 3.1 19.105 3.413 ;
      RECT 18.75 3.127 19.105 3.385 ;
      RECT 18.735 3.14 19.105 3.35 ;
      RECT 18.755 3.115 19.125 3.34 ;
      RECT 18.73 3.18 19.125 3.31 ;
      RECT 18.73 3.21 19.13 3.293 ;
      RECT 18.725 3.24 19.13 3.28 ;
      RECT 18.79 3.089 19.09 3.465 ;
      RECT 18.925 3.086 19.011 3.544 ;
      RECT 18.876 3.087 19.09 3.465 ;
      RECT 19.02 4.747 19.065 4.94 ;
      RECT 19.01 4.717 19.02 4.94 ;
      RECT 19.005 4.702 19.01 4.94 ;
      RECT 18.965 4.612 19.005 4.94 ;
      RECT 18.96 4.525 18.965 4.94 ;
      RECT 18.95 4.495 18.96 4.94 ;
      RECT 18.945 4.455 18.95 4.94 ;
      RECT 18.935 4.417 18.945 4.94 ;
      RECT 18.93 4.382 18.935 4.94 ;
      RECT 18.91 4.335 18.93 4.94 ;
      RECT 18.895 4.26 18.91 4.94 ;
      RECT 18.89 4.215 18.895 4.935 ;
      RECT 18.885 4.195 18.89 4.908 ;
      RECT 18.88 4.175 18.885 4.893 ;
      RECT 18.875 4.15 18.88 4.873 ;
      RECT 18.87 4.128 18.875 4.858 ;
      RECT 18.865 4.106 18.87 4.84 ;
      RECT 18.86 4.085 18.865 4.83 ;
      RECT 18.85 4.057 18.86 4.8 ;
      RECT 18.84 4.02 18.85 4.768 ;
      RECT 18.83 3.98 18.84 4.735 ;
      RECT 18.82 3.958 18.83 4.705 ;
      RECT 18.79 3.91 18.82 4.637 ;
      RECT 18.775 3.87 18.79 4.564 ;
      RECT 18.765 3.87 18.775 4.53 ;
      RECT 18.76 3.87 18.765 4.505 ;
      RECT 18.755 3.87 18.76 4.49 ;
      RECT 18.75 3.87 18.755 4.468 ;
      RECT 18.745 3.87 18.75 4.455 ;
      RECT 18.73 3.87 18.745 4.42 ;
      RECT 18.71 3.87 18.73 4.36 ;
      RECT 18.7 3.87 18.71 4.31 ;
      RECT 18.68 3.87 18.7 4.258 ;
      RECT 18.66 3.87 18.68 4.215 ;
      RECT 18.65 3.87 18.66 4.203 ;
      RECT 18.62 3.87 18.65 4.19 ;
      RECT 18.59 3.891 18.62 4.17 ;
      RECT 18.58 3.919 18.59 4.15 ;
      RECT 18.565 3.936 18.58 4.118 ;
      RECT 18.56 3.95 18.565 4.085 ;
      RECT 18.555 3.958 18.56 4.058 ;
      RECT 18.55 3.966 18.555 4.02 ;
      RECT 18.555 4.49 18.56 4.825 ;
      RECT 18.52 4.477 18.555 4.824 ;
      RECT 18.45 4.417 18.52 4.823 ;
      RECT 18.37 4.36 18.45 4.822 ;
      RECT 18.235 4.32 18.37 4.821 ;
      RECT 18.235 4.507 18.57 4.81 ;
      RECT 18.195 4.507 18.57 4.8 ;
      RECT 18.195 4.525 18.575 4.795 ;
      RECT 18.195 4.615 18.58 4.785 ;
      RECT 18.19 4.31 18.355 4.765 ;
      RECT 18.185 4.31 18.355 4.508 ;
      RECT 18.185 4.467 18.55 4.508 ;
      RECT 18.185 4.455 18.545 4.508 ;
      RECT 16.665 7.305 16.835 9.515 ;
      RECT 16.665 7.305 16.84 8.565 ;
      RECT 16.235 10.145 16.405 10.595 ;
      RECT 16.295 8.365 16.465 10.315 ;
      RECT 16.235 7.305 16.405 8.535 ;
      RECT 15.71 10.105 15.885 10.595 ;
      RECT 15.71 7.305 15.88 10.595 ;
      RECT 15.71 9.605 16.12 9.935 ;
      RECT 15.71 8.765 16.12 9.095 ;
      RECT 15.71 7.305 15.885 8.565 ;
      RECT 96.225 10.085 96.4 10.595 ;
      RECT 95.235 1.865 95.41 2.375 ;
      RECT 95.235 10.085 95.41 10.595 ;
      RECT 93.445 1.865 93.62 2.375 ;
      RECT 93.445 10.085 93.62 10.595 ;
      RECT 91.055 4.145 91.425 4.515 ;
      RECT 88.665 10.085 88.84 10.595 ;
      RECT 80.44 10.085 80.615 10.595 ;
      RECT 79.45 1.865 79.625 2.375 ;
      RECT 79.45 10.085 79.625 10.595 ;
      RECT 77.66 1.865 77.835 2.375 ;
      RECT 77.66 10.085 77.835 10.595 ;
      RECT 75.27 4.145 75.64 4.515 ;
      RECT 72.88 10.085 73.055 10.595 ;
      RECT 64.655 10.085 64.83 10.595 ;
      RECT 63.665 1.865 63.84 2.375 ;
      RECT 63.665 10.085 63.84 10.595 ;
      RECT 61.875 1.865 62.05 2.375 ;
      RECT 61.875 10.085 62.05 10.595 ;
      RECT 59.485 4.145 59.855 4.515 ;
      RECT 57.095 10.085 57.27 10.595 ;
      RECT 48.88 10.085 49.055 10.595 ;
      RECT 47.89 1.865 48.065 2.375 ;
      RECT 47.89 10.085 48.065 10.595 ;
      RECT 46.1 1.865 46.275 2.375 ;
      RECT 46.1 10.085 46.275 10.595 ;
      RECT 43.71 4.145 44.08 4.515 ;
      RECT 41.32 10.085 41.495 10.595 ;
      RECT 33.1 10.085 33.275 10.595 ;
      RECT 32.11 1.865 32.285 2.375 ;
      RECT 32.11 10.085 32.285 10.595 ;
      RECT 30.32 1.865 30.495 2.375 ;
      RECT 30.32 10.085 30.495 10.595 ;
      RECT 27.93 4.145 28.3 4.515 ;
      RECT 25.54 10.085 25.715 10.595 ;
      RECT 16.665 10.085 16.84 10.595 ;
  END
END sky130_osu_ring_oscillator_mpr2aa_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2at_8_b0r1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2at_8_b0r1 ;
  SIZE 107.44 BY 12.61 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 35.085 0 35.465 5.265 ;
      LAYER met2 ;
        RECT 35.1 4.9 35.45 5.25 ;
        RECT 35.13 4.885 35.42 5.265 ;
      LAYER li1 ;
        RECT 35.185 1.865 35.36 2.375 ;
        RECT 35.185 3.895 35.36 5.155 ;
        RECT 35.185 3.685 35.355 5.155 ;
      LAYER met1 ;
        RECT 35.085 4.93 35.465 5.22 ;
        RECT 35.125 2.175 35.42 2.405 ;
        RECT 35.125 3.655 35.415 3.885 ;
        RECT 35.185 2.175 35.355 3.885 ;
      LAYER via1 ;
        RECT 35.2 5 35.35 5.15 ;
      LAYER via2 ;
        RECT 35.175 4.975 35.375 5.175 ;
      LAYER mcon ;
        RECT 35.185 3.685 35.355 3.855 ;
        RECT 35.19 4.985 35.36 5.155 ;
        RECT 35.185 2.205 35.36 2.375 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 53.01 0 53.39 5.265 ;
      LAYER met2 ;
        RECT 53.025 4.9 53.375 5.25 ;
        RECT 53.055 4.885 53.345 5.265 ;
      LAYER li1 ;
        RECT 53.11 1.865 53.285 2.375 ;
        RECT 53.11 3.895 53.285 5.155 ;
        RECT 53.11 3.685 53.28 5.155 ;
      LAYER met1 ;
        RECT 53.01 4.93 53.39 5.22 ;
        RECT 53.05 2.175 53.345 2.405 ;
        RECT 53.05 3.655 53.34 3.885 ;
        RECT 53.11 2.175 53.28 3.885 ;
      LAYER via1 ;
        RECT 53.125 5 53.275 5.15 ;
      LAYER via2 ;
        RECT 53.1 4.975 53.3 5.175 ;
      LAYER mcon ;
        RECT 53.11 3.685 53.28 3.855 ;
        RECT 53.115 4.985 53.285 5.155 ;
        RECT 53.11 2.205 53.285 2.375 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 70.935 0 71.315 5.265 ;
      LAYER met2 ;
        RECT 70.95 4.9 71.3 5.25 ;
        RECT 70.98 4.885 71.27 5.265 ;
      LAYER li1 ;
        RECT 71.035 1.865 71.21 2.375 ;
        RECT 71.035 3.895 71.21 5.155 ;
        RECT 71.035 3.685 71.205 5.155 ;
      LAYER met1 ;
        RECT 70.935 4.93 71.315 5.22 ;
        RECT 70.975 2.175 71.27 2.405 ;
        RECT 70.975 3.655 71.265 3.885 ;
        RECT 71.035 2.175 71.205 3.885 ;
      LAYER via1 ;
        RECT 71.05 5 71.2 5.15 ;
      LAYER via2 ;
        RECT 71.025 4.975 71.225 5.175 ;
      LAYER mcon ;
        RECT 71.035 3.685 71.205 3.855 ;
        RECT 71.04 4.985 71.21 5.155 ;
        RECT 71.035 2.205 71.21 2.375 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 88.86 0 89.24 5.265 ;
      LAYER met2 ;
        RECT 88.875 4.9 89.225 5.25 ;
        RECT 88.905 4.885 89.195 5.265 ;
      LAYER li1 ;
        RECT 88.96 1.865 89.135 2.375 ;
        RECT 88.96 3.895 89.135 5.155 ;
        RECT 88.96 3.685 89.13 5.155 ;
      LAYER met1 ;
        RECT 88.86 4.93 89.24 5.22 ;
        RECT 88.9 2.175 89.195 2.405 ;
        RECT 88.9 3.655 89.19 3.885 ;
        RECT 88.96 2.175 89.13 3.885 ;
      LAYER via1 ;
        RECT 88.975 5 89.125 5.15 ;
      LAYER via2 ;
        RECT 88.95 4.975 89.15 5.175 ;
      LAYER mcon ;
        RECT 88.96 3.685 89.13 3.855 ;
        RECT 88.965 4.985 89.135 5.155 ;
        RECT 88.96 2.205 89.135 2.375 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 106.785 0 107.165 5.265 ;
      LAYER met2 ;
        RECT 106.8 4.9 107.15 5.25 ;
        RECT 106.83 4.885 107.12 5.265 ;
      LAYER li1 ;
        RECT 106.885 1.865 107.06 2.375 ;
        RECT 106.885 3.895 107.06 5.155 ;
        RECT 106.885 3.685 107.055 5.155 ;
      LAYER met1 ;
        RECT 106.785 4.93 107.165 5.22 ;
        RECT 106.825 2.175 107.12 2.405 ;
        RECT 106.825 3.655 107.115 3.885 ;
        RECT 106.885 2.175 107.055 3.885 ;
      LAYER via1 ;
        RECT 106.9 5 107.05 5.15 ;
      LAYER via2 ;
        RECT 106.875 4.975 107.075 5.175 ;
      LAYER mcon ;
        RECT 106.885 3.685 107.055 3.855 ;
        RECT 106.89 4.985 107.06 5.155 ;
        RECT 106.885 2.205 107.06 2.375 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 30.96 4 31.31 4.35 ;
        RECT 30.95 8.275 31.3 8.625 ;
        RECT 31.025 4 31.2 8.625 ;
      LAYER li1 ;
        RECT 31.035 2.955 31.205 4.225 ;
        RECT 31.035 8.385 31.205 9.655 ;
        RECT 26.275 8.385 26.445 9.655 ;
      LAYER met1 ;
        RECT 30.96 4.055 31.435 4.225 ;
        RECT 30.96 4 31.31 4.35 ;
        RECT 30.95 8.385 31.435 8.555 ;
        RECT 30.95 8.275 31.3 8.625 ;
        RECT 26.525 8.38 31.3 8.55 ;
        RECT 26.215 8.385 26.675 8.555 ;
        RECT 26.215 8.355 26.505 8.585 ;
      LAYER via1 ;
        RECT 31.05 8.375 31.2 8.525 ;
        RECT 31.06 4.1 31.21 4.25 ;
      LAYER mcon ;
        RECT 26.275 8.385 26.445 8.555 ;
        RECT 31.035 8.385 31.205 8.555 ;
        RECT 31.035 4.055 31.205 4.225 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 48.885 4 49.235 4.35 ;
        RECT 48.875 8.275 49.225 8.625 ;
        RECT 48.95 4 49.125 8.625 ;
      LAYER li1 ;
        RECT 48.96 2.955 49.13 4.225 ;
        RECT 48.96 8.385 49.13 9.655 ;
        RECT 44.2 8.385 44.37 9.655 ;
      LAYER met1 ;
        RECT 48.885 4.055 49.36 4.225 ;
        RECT 48.885 4 49.235 4.35 ;
        RECT 48.875 8.385 49.36 8.555 ;
        RECT 48.875 8.275 49.225 8.625 ;
        RECT 44.45 8.38 49.225 8.55 ;
        RECT 44.14 8.385 44.6 8.555 ;
        RECT 44.14 8.355 44.43 8.585 ;
      LAYER via1 ;
        RECT 48.975 8.375 49.125 8.525 ;
        RECT 48.985 4.1 49.135 4.25 ;
      LAYER mcon ;
        RECT 44.2 8.385 44.37 8.555 ;
        RECT 48.96 8.385 49.13 8.555 ;
        RECT 48.96 4.055 49.13 4.225 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 66.81 4 67.16 4.35 ;
        RECT 66.8 8.275 67.15 8.625 ;
        RECT 66.875 4 67.05 8.625 ;
      LAYER li1 ;
        RECT 66.885 2.955 67.055 4.225 ;
        RECT 66.885 8.385 67.055 9.655 ;
        RECT 62.125 8.385 62.295 9.655 ;
      LAYER met1 ;
        RECT 66.81 4.055 67.285 4.225 ;
        RECT 66.81 4 67.16 4.35 ;
        RECT 66.8 8.385 67.285 8.555 ;
        RECT 66.8 8.275 67.15 8.625 ;
        RECT 62.375 8.38 67.15 8.55 ;
        RECT 62.065 8.385 62.525 8.555 ;
        RECT 62.065 8.355 62.355 8.585 ;
      LAYER via1 ;
        RECT 66.9 8.375 67.05 8.525 ;
        RECT 66.91 4.1 67.06 4.25 ;
      LAYER mcon ;
        RECT 62.125 8.385 62.295 8.555 ;
        RECT 66.885 8.385 67.055 8.555 ;
        RECT 66.885 4.055 67.055 4.225 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 84.735 4 85.085 4.35 ;
        RECT 84.725 8.275 85.075 8.625 ;
        RECT 84.8 4 84.975 8.625 ;
      LAYER li1 ;
        RECT 84.81 2.955 84.98 4.225 ;
        RECT 84.81 8.385 84.98 9.655 ;
        RECT 80.05 8.385 80.22 9.655 ;
      LAYER met1 ;
        RECT 84.735 4.055 85.21 4.225 ;
        RECT 84.735 4 85.085 4.35 ;
        RECT 84.725 8.385 85.21 8.555 ;
        RECT 84.725 8.275 85.075 8.625 ;
        RECT 80.3 8.38 85.075 8.55 ;
        RECT 79.99 8.385 80.45 8.555 ;
        RECT 79.99 8.355 80.28 8.585 ;
      LAYER via1 ;
        RECT 84.825 8.375 84.975 8.525 ;
        RECT 84.835 4.1 84.985 4.25 ;
      LAYER mcon ;
        RECT 80.05 8.385 80.22 8.555 ;
        RECT 84.81 8.385 84.98 8.555 ;
        RECT 84.81 4.055 84.98 4.225 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 102.66 4 103.01 4.35 ;
        RECT 102.65 8.275 103 8.625 ;
        RECT 102.725 4 102.9 8.625 ;
      LAYER li1 ;
        RECT 102.735 2.955 102.905 4.225 ;
        RECT 102.735 8.385 102.905 9.655 ;
        RECT 97.975 8.385 98.145 9.655 ;
      LAYER met1 ;
        RECT 102.66 4.055 103.135 4.225 ;
        RECT 102.66 4 103.01 4.35 ;
        RECT 102.65 8.385 103.135 8.555 ;
        RECT 102.65 8.275 103 8.625 ;
        RECT 98.225 8.38 103 8.55 ;
        RECT 97.915 8.385 98.375 8.555 ;
        RECT 97.915 8.355 98.205 8.585 ;
      LAYER via1 ;
        RECT 102.75 8.375 102.9 8.525 ;
        RECT 102.76 4.1 102.91 4.25 ;
      LAYER mcon ;
        RECT 97.975 8.385 98.145 8.555 ;
        RECT 102.735 8.385 102.905 8.555 ;
        RECT 102.735 4.055 102.905 4.225 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 15.245 8.385 15.415 9.655 ;
      LAYER met1 ;
        RECT 15.185 8.385 15.645 8.555 ;
        RECT 15.19 8.35 15.48 8.58 ;
        RECT 15.185 8.355 15.475 8.585 ;
      LAYER mcon ;
        RECT 15.245 8.385 15.415 8.555 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.015 5.58 107.435 7.18 ;
        RECT 101.475 5.43 107.435 7.18 ;
        RECT 102.555 5.43 107.28 7.185 ;
        RECT 102.555 5.425 107.275 7.185 ;
        RECT 106.46 5.425 106.63 7.915 ;
        RECT 106.455 4.695 106.625 7.185 ;
        RECT 105.47 4.695 105.64 7.915 ;
        RECT 102.725 4.695 102.895 7.915 ;
        RECT 97.795 5.58 100.545 7.185 ;
        RECT 99.985 5.08 100.155 7.185 ;
        RECT 97.965 5.58 98.135 7.915 ;
        RECT 97.545 5.08 97.715 7.18 ;
        RECT 95.585 5.08 95.755 7.18 ;
        RECT 94.625 5.08 94.795 7.18 ;
        RECT 92.665 5.08 92.835 7.18 ;
        RECT 91.665 5.08 91.835 7.18 ;
        RECT 90.705 5.08 90.875 7.18 ;
        RECT 83.55 5.43 89.51 7.18 ;
        RECT 84.63 5.43 89.355 7.185 ;
        RECT 84.63 5.425 89.35 7.185 ;
        RECT 88.535 5.425 88.705 7.915 ;
        RECT 88.53 4.695 88.7 7.185 ;
        RECT 87.545 4.695 87.715 7.915 ;
        RECT 84.8 4.695 84.97 7.915 ;
        RECT 79.87 5.58 82.62 7.185 ;
        RECT 82.06 5.08 82.23 7.185 ;
        RECT 80.04 5.58 80.21 7.915 ;
        RECT 79.62 5.08 79.79 7.18 ;
        RECT 77.66 5.08 77.83 7.18 ;
        RECT 76.7 5.08 76.87 7.18 ;
        RECT 74.74 5.08 74.91 7.18 ;
        RECT 73.74 5.08 73.91 7.18 ;
        RECT 72.78 5.08 72.95 7.18 ;
        RECT 65.625 5.43 71.585 7.18 ;
        RECT 66.705 5.43 71.43 7.185 ;
        RECT 66.705 5.425 71.425 7.185 ;
        RECT 70.61 5.425 70.78 7.915 ;
        RECT 70.605 4.695 70.775 7.185 ;
        RECT 69.62 4.695 69.79 7.915 ;
        RECT 66.875 4.695 67.045 7.915 ;
        RECT 61.945 5.58 64.695 7.185 ;
        RECT 64.135 5.08 64.305 7.185 ;
        RECT 62.115 5.58 62.285 7.915 ;
        RECT 61.695 5.08 61.865 7.18 ;
        RECT 59.735 5.08 59.905 7.18 ;
        RECT 58.775 5.08 58.945 7.18 ;
        RECT 56.815 5.08 56.985 7.18 ;
        RECT 55.815 5.08 55.985 7.18 ;
        RECT 54.855 5.08 55.025 7.18 ;
        RECT 47.7 5.43 53.66 7.18 ;
        RECT 48.78 5.43 53.505 7.185 ;
        RECT 48.78 5.425 53.5 7.185 ;
        RECT 52.685 5.425 52.855 7.915 ;
        RECT 52.68 4.695 52.85 7.185 ;
        RECT 51.695 4.695 51.865 7.915 ;
        RECT 48.95 4.695 49.12 7.915 ;
        RECT 44.02 5.58 46.77 7.185 ;
        RECT 46.21 5.08 46.38 7.185 ;
        RECT 44.19 5.58 44.36 7.915 ;
        RECT 43.77 5.08 43.94 7.18 ;
        RECT 41.81 5.08 41.98 7.18 ;
        RECT 40.85 5.08 41.02 7.18 ;
        RECT 38.89 5.08 39.06 7.18 ;
        RECT 37.89 5.08 38.06 7.18 ;
        RECT 36.93 5.08 37.1 7.18 ;
        RECT 29.775 5.43 35.735 7.18 ;
        RECT 30.855 5.43 35.58 7.185 ;
        RECT 30.855 5.425 35.575 7.185 ;
        RECT 34.76 5.425 34.93 7.915 ;
        RECT 34.755 4.695 34.925 7.185 ;
        RECT 33.77 4.695 33.94 7.915 ;
        RECT 31.025 4.695 31.195 7.915 ;
        RECT 26.095 5.58 28.845 7.185 ;
        RECT 28.285 5.08 28.455 7.185 ;
        RECT 26.265 5.58 26.435 7.915 ;
        RECT 25.845 5.08 26.015 7.18 ;
        RECT 23.885 5.08 24.055 7.18 ;
        RECT 22.925 5.08 23.095 7.18 ;
        RECT 20.965 5.08 21.135 7.18 ;
        RECT 19.965 5.08 20.135 7.18 ;
        RECT 19.005 5.08 19.175 7.18 ;
        RECT 15.065 5.58 17.815 7.185 ;
        RECT 17.05 10.195 17.225 10.745 ;
        RECT 17.05 7.455 17.225 8.595 ;
        RECT 17.05 5.58 17.22 10.745 ;
        RECT 15.235 5.58 15.405 7.915 ;
      LAYER met1 ;
        RECT 0.015 5.58 107.435 7.18 ;
        RECT 89.895 5.43 107.435 7.18 ;
        RECT 102.555 5.43 107.28 7.185 ;
        RECT 102.555 5.425 107.275 7.185 ;
        RECT 89.895 5.425 101.855 7.18 ;
        RECT 97.795 5.425 100.545 7.185 ;
        RECT 71.97 5.43 89.51 7.18 ;
        RECT 84.63 5.43 89.355 7.185 ;
        RECT 84.63 5.425 89.35 7.185 ;
        RECT 71.97 5.425 83.93 7.18 ;
        RECT 79.87 5.425 82.62 7.185 ;
        RECT 54.045 5.43 71.585 7.18 ;
        RECT 66.705 5.43 71.43 7.185 ;
        RECT 66.705 5.425 71.425 7.185 ;
        RECT 54.045 5.425 66.005 7.18 ;
        RECT 61.945 5.425 64.695 7.185 ;
        RECT 36.12 5.43 53.66 7.18 ;
        RECT 48.78 5.43 53.505 7.185 ;
        RECT 48.78 5.425 53.5 7.185 ;
        RECT 36.12 5.425 48.08 7.18 ;
        RECT 44.02 5.425 46.77 7.185 ;
        RECT 18.195 5.43 35.735 7.18 ;
        RECT 30.855 5.43 35.58 7.185 ;
        RECT 30.855 5.425 35.575 7.185 ;
        RECT 18.195 5.425 30.155 7.18 ;
        RECT 26.095 5.425 28.845 7.185 ;
        RECT 15.065 5.58 17.815 7.185 ;
        RECT 16.99 9.095 17.28 9.325 ;
        RECT 16.82 9.125 17.28 9.295 ;
      LAYER mcon ;
        RECT 17.05 9.125 17.22 9.295 ;
        RECT 17.355 6.985 17.525 7.155 ;
        RECT 18.34 5.58 18.51 5.75 ;
        RECT 18.8 5.58 18.97 5.75 ;
        RECT 19.26 5.58 19.43 5.75 ;
        RECT 19.72 5.58 19.89 5.75 ;
        RECT 20.18 5.58 20.35 5.75 ;
        RECT 20.64 5.58 20.81 5.75 ;
        RECT 21.1 5.58 21.27 5.75 ;
        RECT 21.56 5.58 21.73 5.75 ;
        RECT 22.02 5.58 22.19 5.75 ;
        RECT 22.48 5.58 22.65 5.75 ;
        RECT 22.94 5.58 23.11 5.75 ;
        RECT 23.4 5.58 23.57 5.75 ;
        RECT 23.86 5.58 24.03 5.75 ;
        RECT 24.32 5.58 24.49 5.75 ;
        RECT 24.78 5.58 24.95 5.75 ;
        RECT 25.24 5.58 25.41 5.75 ;
        RECT 25.7 5.58 25.87 5.75 ;
        RECT 26.16 5.58 26.33 5.75 ;
        RECT 26.62 5.58 26.79 5.75 ;
        RECT 27.08 5.58 27.25 5.75 ;
        RECT 27.54 5.58 27.71 5.75 ;
        RECT 28 5.58 28.17 5.75 ;
        RECT 28.385 6.985 28.555 7.155 ;
        RECT 28.46 5.58 28.63 5.75 ;
        RECT 28.92 5.58 29.09 5.75 ;
        RECT 29.38 5.58 29.55 5.75 ;
        RECT 29.84 5.58 30.01 5.75 ;
        RECT 33.145 6.985 33.315 7.155 ;
        RECT 33.145 5.455 33.315 5.625 ;
        RECT 33.85 6.985 34.02 7.155 ;
        RECT 33.85 5.455 34.02 5.625 ;
        RECT 34.835 5.455 35.005 5.625 ;
        RECT 34.84 6.985 35.01 7.155 ;
        RECT 36.265 5.58 36.435 5.75 ;
        RECT 36.725 5.58 36.895 5.75 ;
        RECT 37.185 5.58 37.355 5.75 ;
        RECT 37.645 5.58 37.815 5.75 ;
        RECT 38.105 5.58 38.275 5.75 ;
        RECT 38.565 5.58 38.735 5.75 ;
        RECT 39.025 5.58 39.195 5.75 ;
        RECT 39.485 5.58 39.655 5.75 ;
        RECT 39.945 5.58 40.115 5.75 ;
        RECT 40.405 5.58 40.575 5.75 ;
        RECT 40.865 5.58 41.035 5.75 ;
        RECT 41.325 5.58 41.495 5.75 ;
        RECT 41.785 5.58 41.955 5.75 ;
        RECT 42.245 5.58 42.415 5.75 ;
        RECT 42.705 5.58 42.875 5.75 ;
        RECT 43.165 5.58 43.335 5.75 ;
        RECT 43.625 5.58 43.795 5.75 ;
        RECT 44.085 5.58 44.255 5.75 ;
        RECT 44.545 5.58 44.715 5.75 ;
        RECT 45.005 5.58 45.175 5.75 ;
        RECT 45.465 5.58 45.635 5.75 ;
        RECT 45.925 5.58 46.095 5.75 ;
        RECT 46.31 6.985 46.48 7.155 ;
        RECT 46.385 5.58 46.555 5.75 ;
        RECT 46.845 5.58 47.015 5.75 ;
        RECT 47.305 5.58 47.475 5.75 ;
        RECT 47.765 5.58 47.935 5.75 ;
        RECT 51.07 6.985 51.24 7.155 ;
        RECT 51.07 5.455 51.24 5.625 ;
        RECT 51.775 6.985 51.945 7.155 ;
        RECT 51.775 5.455 51.945 5.625 ;
        RECT 52.76 5.455 52.93 5.625 ;
        RECT 52.765 6.985 52.935 7.155 ;
        RECT 54.19 5.58 54.36 5.75 ;
        RECT 54.65 5.58 54.82 5.75 ;
        RECT 55.11 5.58 55.28 5.75 ;
        RECT 55.57 5.58 55.74 5.75 ;
        RECT 56.03 5.58 56.2 5.75 ;
        RECT 56.49 5.58 56.66 5.75 ;
        RECT 56.95 5.58 57.12 5.75 ;
        RECT 57.41 5.58 57.58 5.75 ;
        RECT 57.87 5.58 58.04 5.75 ;
        RECT 58.33 5.58 58.5 5.75 ;
        RECT 58.79 5.58 58.96 5.75 ;
        RECT 59.25 5.58 59.42 5.75 ;
        RECT 59.71 5.58 59.88 5.75 ;
        RECT 60.17 5.58 60.34 5.75 ;
        RECT 60.63 5.58 60.8 5.75 ;
        RECT 61.09 5.58 61.26 5.75 ;
        RECT 61.55 5.58 61.72 5.75 ;
        RECT 62.01 5.58 62.18 5.75 ;
        RECT 62.47 5.58 62.64 5.75 ;
        RECT 62.93 5.58 63.1 5.75 ;
        RECT 63.39 5.58 63.56 5.75 ;
        RECT 63.85 5.58 64.02 5.75 ;
        RECT 64.235 6.985 64.405 7.155 ;
        RECT 64.31 5.58 64.48 5.75 ;
        RECT 64.77 5.58 64.94 5.75 ;
        RECT 65.23 5.58 65.4 5.75 ;
        RECT 65.69 5.58 65.86 5.75 ;
        RECT 68.995 6.985 69.165 7.155 ;
        RECT 68.995 5.455 69.165 5.625 ;
        RECT 69.7 6.985 69.87 7.155 ;
        RECT 69.7 5.455 69.87 5.625 ;
        RECT 70.685 5.455 70.855 5.625 ;
        RECT 70.69 6.985 70.86 7.155 ;
        RECT 72.115 5.58 72.285 5.75 ;
        RECT 72.575 5.58 72.745 5.75 ;
        RECT 73.035 5.58 73.205 5.75 ;
        RECT 73.495 5.58 73.665 5.75 ;
        RECT 73.955 5.58 74.125 5.75 ;
        RECT 74.415 5.58 74.585 5.75 ;
        RECT 74.875 5.58 75.045 5.75 ;
        RECT 75.335 5.58 75.505 5.75 ;
        RECT 75.795 5.58 75.965 5.75 ;
        RECT 76.255 5.58 76.425 5.75 ;
        RECT 76.715 5.58 76.885 5.75 ;
        RECT 77.175 5.58 77.345 5.75 ;
        RECT 77.635 5.58 77.805 5.75 ;
        RECT 78.095 5.58 78.265 5.75 ;
        RECT 78.555 5.58 78.725 5.75 ;
        RECT 79.015 5.58 79.185 5.75 ;
        RECT 79.475 5.58 79.645 5.75 ;
        RECT 79.935 5.58 80.105 5.75 ;
        RECT 80.395 5.58 80.565 5.75 ;
        RECT 80.855 5.58 81.025 5.75 ;
        RECT 81.315 5.58 81.485 5.75 ;
        RECT 81.775 5.58 81.945 5.75 ;
        RECT 82.16 6.985 82.33 7.155 ;
        RECT 82.235 5.58 82.405 5.75 ;
        RECT 82.695 5.58 82.865 5.75 ;
        RECT 83.155 5.58 83.325 5.75 ;
        RECT 83.615 5.58 83.785 5.75 ;
        RECT 86.92 6.985 87.09 7.155 ;
        RECT 86.92 5.455 87.09 5.625 ;
        RECT 87.625 6.985 87.795 7.155 ;
        RECT 87.625 5.455 87.795 5.625 ;
        RECT 88.61 5.455 88.78 5.625 ;
        RECT 88.615 6.985 88.785 7.155 ;
        RECT 90.04 5.58 90.21 5.75 ;
        RECT 90.5 5.58 90.67 5.75 ;
        RECT 90.96 5.58 91.13 5.75 ;
        RECT 91.42 5.58 91.59 5.75 ;
        RECT 91.88 5.58 92.05 5.75 ;
        RECT 92.34 5.58 92.51 5.75 ;
        RECT 92.8 5.58 92.97 5.75 ;
        RECT 93.26 5.58 93.43 5.75 ;
        RECT 93.72 5.58 93.89 5.75 ;
        RECT 94.18 5.58 94.35 5.75 ;
        RECT 94.64 5.58 94.81 5.75 ;
        RECT 95.1 5.58 95.27 5.75 ;
        RECT 95.56 5.58 95.73 5.75 ;
        RECT 96.02 5.58 96.19 5.75 ;
        RECT 96.48 5.58 96.65 5.75 ;
        RECT 96.94 5.58 97.11 5.75 ;
        RECT 97.4 5.58 97.57 5.75 ;
        RECT 97.86 5.58 98.03 5.75 ;
        RECT 98.32 5.58 98.49 5.75 ;
        RECT 98.78 5.58 98.95 5.75 ;
        RECT 99.24 5.58 99.41 5.75 ;
        RECT 99.7 5.58 99.87 5.75 ;
        RECT 100.085 6.985 100.255 7.155 ;
        RECT 100.16 5.58 100.33 5.75 ;
        RECT 100.62 5.58 100.79 5.75 ;
        RECT 101.08 5.58 101.25 5.75 ;
        RECT 101.54 5.58 101.71 5.75 ;
        RECT 104.845 6.985 105.015 7.155 ;
        RECT 104.845 5.455 105.015 5.625 ;
        RECT 105.55 6.985 105.72 7.155 ;
        RECT 105.55 5.455 105.72 5.625 ;
        RECT 106.535 5.455 106.705 5.625 ;
        RECT 106.54 6.985 106.71 7.155 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 91.51 3.86 92.24 4.19 ;
        RECT 73.585 3.86 74.315 4.19 ;
        RECT 55.66 3.86 56.39 4.19 ;
        RECT 37.735 3.86 38.465 4.19 ;
        RECT 19.81 3.86 20.54 4.19 ;
      LAYER met2 ;
        RECT 93.185 3.93 93.445 4.19 ;
        RECT 91.86 3.9 93.205 4.175 ;
        RECT 91.855 2.5 92.2 2.845 ;
        RECT 91.86 3.885 92.15 4.49 ;
        RECT 91.95 2.5 92.12 4.49 ;
        RECT 91.815 4.41 92.075 4.67 ;
        RECT 91.855 4.165 92.265 4.49 ;
        RECT 75.26 3.93 75.52 4.19 ;
        RECT 73.935 3.9 75.28 4.175 ;
        RECT 73.93 2.5 74.275 2.845 ;
        RECT 73.935 3.885 74.225 4.49 ;
        RECT 74.025 2.5 74.195 4.49 ;
        RECT 73.89 4.41 74.15 4.67 ;
        RECT 73.93 4.165 74.34 4.49 ;
        RECT 57.335 3.93 57.595 4.19 ;
        RECT 56.01 3.9 57.355 4.175 ;
        RECT 56.005 2.5 56.35 2.845 ;
        RECT 56.01 3.885 56.3 4.49 ;
        RECT 56.1 2.5 56.27 4.49 ;
        RECT 55.965 4.41 56.225 4.67 ;
        RECT 56.005 4.165 56.415 4.49 ;
        RECT 39.41 3.93 39.67 4.19 ;
        RECT 38.085 3.9 39.43 4.175 ;
        RECT 38.08 2.5 38.425 2.845 ;
        RECT 38.085 3.885 38.375 4.49 ;
        RECT 38.175 2.5 38.345 4.49 ;
        RECT 38.04 4.41 38.3 4.67 ;
        RECT 38.08 4.165 38.49 4.49 ;
        RECT 21.485 3.93 21.745 4.19 ;
        RECT 20.16 3.9 21.505 4.175 ;
        RECT 20.155 2.5 20.5 2.845 ;
        RECT 20.16 3.885 20.45 4.49 ;
        RECT 20.25 2.5 20.42 4.49 ;
        RECT 20.115 4.41 20.375 4.67 ;
        RECT 20.155 4.165 20.565 4.49 ;
      LAYER li1 ;
        RECT 0 11.01 107.44 12.61 ;
        RECT 106.46 10.385 106.63 12.61 ;
        RECT 105.47 10.385 105.64 12.61 ;
        RECT 102.725 10.385 102.895 12.61 ;
        RECT 97.965 10.385 98.135 12.61 ;
        RECT 88.535 10.385 88.705 12.61 ;
        RECT 87.545 10.385 87.715 12.61 ;
        RECT 84.8 10.385 84.97 12.61 ;
        RECT 80.04 10.385 80.21 12.61 ;
        RECT 70.61 10.385 70.78 12.61 ;
        RECT 69.62 10.385 69.79 12.61 ;
        RECT 66.875 10.385 67.045 12.61 ;
        RECT 62.115 10.385 62.285 12.61 ;
        RECT 52.685 10.385 52.855 12.61 ;
        RECT 51.695 10.385 51.865 12.61 ;
        RECT 48.95 10.385 49.12 12.61 ;
        RECT 44.19 10.385 44.36 12.61 ;
        RECT 34.76 10.385 34.93 12.61 ;
        RECT 33.77 10.385 33.94 12.61 ;
        RECT 31.025 10.385 31.195 12.61 ;
        RECT 26.265 10.385 26.435 12.61 ;
        RECT 15.235 10.385 15.405 12.61 ;
        RECT 0.015 0 107.435 1.6 ;
        RECT 106.455 0 106.625 2.225 ;
        RECT 105.47 0 105.64 2.225 ;
        RECT 102.725 0 102.895 2.225 ;
        RECT 89.895 2.86 101.855 3.03 ;
        RECT 89.88 0 101.79 2.975 ;
        RECT 100.945 0 101.115 3.53 ;
        RECT 99.985 0 100.155 3.53 ;
        RECT 99.025 0 99.195 3.53 ;
        RECT 98.505 0 98.675 3.53 ;
        RECT 97.545 0 97.715 3.53 ;
        RECT 96.545 0 96.715 3.53 ;
        RECT 95.585 0 95.755 3.53 ;
        RECT 94.105 0 94.275 3.53 ;
        RECT 92.185 0 92.355 3.53 ;
        RECT 90.705 0 90.875 3.53 ;
        RECT 88.53 0 88.7 2.225 ;
        RECT 87.545 0 87.715 2.225 ;
        RECT 84.8 0 84.97 2.225 ;
        RECT 71.97 2.86 83.93 3.03 ;
        RECT 71.955 0 83.865 2.975 ;
        RECT 83.02 0 83.19 3.53 ;
        RECT 82.06 0 82.23 3.53 ;
        RECT 81.1 0 81.27 3.53 ;
        RECT 80.58 0 80.75 3.53 ;
        RECT 79.62 0 79.79 3.53 ;
        RECT 78.62 0 78.79 3.53 ;
        RECT 77.66 0 77.83 3.53 ;
        RECT 76.18 0 76.35 3.53 ;
        RECT 74.26 0 74.43 3.53 ;
        RECT 72.78 0 72.95 3.53 ;
        RECT 70.605 0 70.775 2.225 ;
        RECT 69.62 0 69.79 2.225 ;
        RECT 66.875 0 67.045 2.225 ;
        RECT 54.045 2.86 66.005 3.03 ;
        RECT 54.03 0 65.94 2.975 ;
        RECT 65.095 0 65.265 3.53 ;
        RECT 64.135 0 64.305 3.53 ;
        RECT 63.175 0 63.345 3.53 ;
        RECT 62.655 0 62.825 3.53 ;
        RECT 61.695 0 61.865 3.53 ;
        RECT 60.695 0 60.865 3.53 ;
        RECT 59.735 0 59.905 3.53 ;
        RECT 58.255 0 58.425 3.53 ;
        RECT 56.335 0 56.505 3.53 ;
        RECT 54.855 0 55.025 3.53 ;
        RECT 52.68 0 52.85 2.225 ;
        RECT 51.695 0 51.865 2.225 ;
        RECT 48.95 0 49.12 2.225 ;
        RECT 36.12 2.86 48.08 3.03 ;
        RECT 36.105 0 48.015 2.975 ;
        RECT 47.17 0 47.34 3.53 ;
        RECT 46.21 0 46.38 3.53 ;
        RECT 45.25 0 45.42 3.53 ;
        RECT 44.73 0 44.9 3.53 ;
        RECT 43.77 0 43.94 3.53 ;
        RECT 42.77 0 42.94 3.53 ;
        RECT 41.81 0 41.98 3.53 ;
        RECT 40.33 0 40.5 3.53 ;
        RECT 38.41 0 38.58 3.53 ;
        RECT 36.93 0 37.1 3.53 ;
        RECT 34.755 0 34.925 2.225 ;
        RECT 33.77 0 33.94 2.225 ;
        RECT 31.025 0 31.195 2.225 ;
        RECT 18.195 2.86 30.155 3.03 ;
        RECT 18.18 0 30.09 2.975 ;
        RECT 29.245 0 29.415 3.53 ;
        RECT 28.285 0 28.455 3.53 ;
        RECT 27.325 0 27.495 3.53 ;
        RECT 26.805 0 26.975 3.53 ;
        RECT 25.845 0 26.015 3.53 ;
        RECT 24.845 0 25.015 3.53 ;
        RECT 23.885 0 24.055 3.53 ;
        RECT 22.405 0 22.575 3.53 ;
        RECT 20.485 0 20.655 3.53 ;
        RECT 19.005 0 19.175 3.53 ;
        RECT 98.98 8.515 99.15 10.465 ;
        RECT 98.92 10.295 99.09 10.745 ;
        RECT 98.92 7.455 99.09 8.685 ;
        RECT 93.285 3.965 93.595 4.29 ;
        RECT 91.755 4.165 91.96 4.61 ;
        RECT 91.425 4.09 91.875 4.275 ;
        RECT 91.425 4.02 91.835 4.275 ;
        RECT 91.75 4.165 91.96 4.58 ;
        RECT 91.745 4.165 91.96 4.53 ;
        RECT 91.735 4.165 91.96 4.495 ;
        RECT 91.73 4.165 91.96 4.455 ;
        RECT 91.715 4.165 91.96 4.43 ;
        RECT 91.7 4.165 91.96 4.375 ;
        RECT 91.69 4.165 91.96 4.355 ;
        RECT 91.665 4.165 91.96 4.345 ;
        RECT 91.595 4.165 91.96 4.34 ;
        RECT 91.425 4.015 91.605 4.275 ;
        RECT 91.575 4.165 91.96 4.32 ;
        RECT 91.54 4.165 91.96 4.31 ;
        RECT 81.055 8.515 81.225 10.465 ;
        RECT 80.995 10.295 81.165 10.745 ;
        RECT 80.995 7.455 81.165 8.685 ;
        RECT 75.36 3.965 75.67 4.29 ;
        RECT 73.83 4.165 74.035 4.61 ;
        RECT 73.5 4.09 73.95 4.275 ;
        RECT 73.5 4.02 73.91 4.275 ;
        RECT 73.825 4.165 74.035 4.58 ;
        RECT 73.82 4.165 74.035 4.53 ;
        RECT 73.81 4.165 74.035 4.495 ;
        RECT 73.805 4.165 74.035 4.455 ;
        RECT 73.79 4.165 74.035 4.43 ;
        RECT 73.775 4.165 74.035 4.375 ;
        RECT 73.765 4.165 74.035 4.355 ;
        RECT 73.74 4.165 74.035 4.345 ;
        RECT 73.67 4.165 74.035 4.34 ;
        RECT 73.5 4.015 73.68 4.275 ;
        RECT 73.65 4.165 74.035 4.32 ;
        RECT 73.615 4.165 74.035 4.31 ;
        RECT 63.13 8.515 63.3 10.465 ;
        RECT 63.07 10.295 63.24 10.745 ;
        RECT 63.07 7.455 63.24 8.685 ;
        RECT 57.435 3.965 57.745 4.29 ;
        RECT 55.905 4.165 56.11 4.61 ;
        RECT 55.575 4.09 56.025 4.275 ;
        RECT 55.575 4.02 55.985 4.275 ;
        RECT 55.9 4.165 56.11 4.58 ;
        RECT 55.895 4.165 56.11 4.53 ;
        RECT 55.885 4.165 56.11 4.495 ;
        RECT 55.88 4.165 56.11 4.455 ;
        RECT 55.865 4.165 56.11 4.43 ;
        RECT 55.85 4.165 56.11 4.375 ;
        RECT 55.84 4.165 56.11 4.355 ;
        RECT 55.815 4.165 56.11 4.345 ;
        RECT 55.745 4.165 56.11 4.34 ;
        RECT 55.575 4.015 55.755 4.275 ;
        RECT 55.725 4.165 56.11 4.32 ;
        RECT 55.69 4.165 56.11 4.31 ;
        RECT 45.205 8.515 45.375 10.465 ;
        RECT 45.145 10.295 45.315 10.745 ;
        RECT 45.145 7.455 45.315 8.685 ;
        RECT 39.51 3.965 39.82 4.29 ;
        RECT 37.98 4.165 38.185 4.61 ;
        RECT 37.65 4.09 38.1 4.275 ;
        RECT 37.65 4.02 38.06 4.275 ;
        RECT 37.975 4.165 38.185 4.58 ;
        RECT 37.97 4.165 38.185 4.53 ;
        RECT 37.96 4.165 38.185 4.495 ;
        RECT 37.955 4.165 38.185 4.455 ;
        RECT 37.94 4.165 38.185 4.43 ;
        RECT 37.925 4.165 38.185 4.375 ;
        RECT 37.915 4.165 38.185 4.355 ;
        RECT 37.89 4.165 38.185 4.345 ;
        RECT 37.82 4.165 38.185 4.34 ;
        RECT 37.65 4.015 37.83 4.275 ;
        RECT 37.8 4.165 38.185 4.32 ;
        RECT 37.765 4.165 38.185 4.31 ;
        RECT 27.28 8.515 27.45 10.465 ;
        RECT 27.22 10.295 27.39 10.745 ;
        RECT 27.22 7.455 27.39 8.685 ;
        RECT 21.585 3.965 21.895 4.29 ;
        RECT 20.055 4.165 20.26 4.61 ;
        RECT 19.725 4.09 20.175 4.275 ;
        RECT 19.725 4.02 20.135 4.275 ;
        RECT 20.05 4.165 20.26 4.58 ;
        RECT 20.045 4.165 20.26 4.53 ;
        RECT 20.035 4.165 20.26 4.495 ;
        RECT 20.03 4.165 20.26 4.455 ;
        RECT 20.015 4.165 20.26 4.43 ;
        RECT 20 4.165 20.26 4.375 ;
        RECT 19.99 4.165 20.26 4.355 ;
        RECT 19.965 4.165 20.26 4.345 ;
        RECT 19.895 4.165 20.26 4.34 ;
        RECT 19.725 4.015 19.905 4.275 ;
        RECT 19.875 4.165 20.26 4.32 ;
        RECT 19.84 4.165 20.26 4.31 ;
      LAYER met1 ;
        RECT 0 11.01 107.44 12.61 ;
        RECT 98.92 8.725 99.21 8.955 ;
        RECT 98.58 8.75 99.21 8.925 ;
        RECT 98.58 8.75 98.75 12.61 ;
        RECT 80.995 8.725 81.285 8.955 ;
        RECT 80.655 8.75 81.285 8.925 ;
        RECT 80.655 8.75 80.825 12.61 ;
        RECT 63.07 8.725 63.36 8.955 ;
        RECT 62.73 8.75 63.36 8.925 ;
        RECT 62.73 8.75 62.9 12.61 ;
        RECT 45.145 8.725 45.435 8.955 ;
        RECT 44.805 8.75 45.435 8.925 ;
        RECT 44.805 8.75 44.975 12.61 ;
        RECT 27.22 8.725 27.51 8.955 ;
        RECT 26.88 8.75 27.51 8.925 ;
        RECT 26.88 8.75 27.05 12.61 ;
        RECT 0.015 0 107.435 1.6 ;
        RECT 89.895 2.705 101.855 3.185 ;
        RECT 89.88 2.58 101.79 2.975 ;
        RECT 94.31 0 101.79 3.185 ;
        RECT 90.905 0 101.79 2.3 ;
        RECT 92.875 0 94.03 3.185 ;
        RECT 89.88 2.55 92.595 2.975 ;
        RECT 90.905 0 92.595 3.185 ;
        RECT 89.88 0 101.79 2.27 ;
        RECT 89.88 0 90.625 2.975 ;
        RECT 71.97 2.705 83.93 3.185 ;
        RECT 71.955 2.58 83.865 2.975 ;
        RECT 76.385 0 83.865 3.185 ;
        RECT 72.98 0 83.865 2.3 ;
        RECT 74.95 0 76.105 3.185 ;
        RECT 71.955 2.55 74.67 2.975 ;
        RECT 72.98 0 74.67 3.185 ;
        RECT 71.955 0 83.865 2.27 ;
        RECT 71.955 0 72.7 2.975 ;
        RECT 54.045 2.705 66.005 3.185 ;
        RECT 54.03 2.58 65.94 2.975 ;
        RECT 58.46 0 65.94 3.185 ;
        RECT 55.055 0 65.94 2.3 ;
        RECT 57.025 0 58.18 3.185 ;
        RECT 54.03 2.55 56.745 2.975 ;
        RECT 55.055 0 56.745 3.185 ;
        RECT 54.03 0 65.94 2.27 ;
        RECT 54.03 0 54.775 2.975 ;
        RECT 36.12 2.705 48.08 3.185 ;
        RECT 36.105 2.58 48.015 2.975 ;
        RECT 40.535 0 48.015 3.185 ;
        RECT 37.13 0 48.015 2.3 ;
        RECT 39.1 0 40.255 3.185 ;
        RECT 36.105 2.55 38.82 2.975 ;
        RECT 37.13 0 38.82 3.185 ;
        RECT 36.105 0 48.015 2.27 ;
        RECT 36.105 0 36.85 2.975 ;
        RECT 18.195 2.705 30.155 3.185 ;
        RECT 18.18 2.58 30.09 2.975 ;
        RECT 22.61 0 30.09 3.185 ;
        RECT 19.205 0 30.09 2.3 ;
        RECT 21.175 0 22.33 3.185 ;
        RECT 18.18 2.55 20.895 2.975 ;
        RECT 19.205 0 20.895 3.185 ;
        RECT 18.18 0 30.09 2.27 ;
        RECT 18.18 0 18.925 2.975 ;
        RECT 93.185 3.945 93.485 4.165 ;
        RECT 93.185 3.93 93.445 4.19 ;
        RECT 91.815 4.41 92.075 4.67 ;
        RECT 91.72 4.41 92.075 4.64 ;
        RECT 75.26 3.945 75.56 4.165 ;
        RECT 75.26 3.93 75.52 4.19 ;
        RECT 73.89 4.41 74.15 4.67 ;
        RECT 73.795 4.41 74.15 4.64 ;
        RECT 57.335 3.945 57.635 4.165 ;
        RECT 57.335 3.93 57.595 4.19 ;
        RECT 55.965 4.41 56.225 4.67 ;
        RECT 55.87 4.41 56.225 4.64 ;
        RECT 39.41 3.945 39.71 4.165 ;
        RECT 39.41 3.93 39.67 4.19 ;
        RECT 38.04 4.41 38.3 4.67 ;
        RECT 37.945 4.41 38.3 4.64 ;
        RECT 21.485 3.945 21.785 4.165 ;
        RECT 21.485 3.93 21.745 4.19 ;
        RECT 20.115 4.41 20.375 4.67 ;
        RECT 20.02 4.41 20.375 4.64 ;
      LAYER via1 ;
        RECT 20.17 4.465 20.32 4.615 ;
        RECT 20.25 2.595 20.4 2.745 ;
        RECT 21.54 3.985 21.69 4.135 ;
        RECT 38.095 4.465 38.245 4.615 ;
        RECT 38.175 2.595 38.325 2.745 ;
        RECT 39.465 3.985 39.615 4.135 ;
        RECT 56.02 4.465 56.17 4.615 ;
        RECT 56.1 2.595 56.25 2.745 ;
        RECT 57.39 3.985 57.54 4.135 ;
        RECT 73.945 4.465 74.095 4.615 ;
        RECT 74.025 2.595 74.175 2.745 ;
        RECT 75.315 3.985 75.465 4.135 ;
        RECT 91.87 4.465 92.02 4.615 ;
        RECT 91.95 2.595 92.1 2.745 ;
        RECT 93.24 3.985 93.39 4.135 ;
      LAYER via2 ;
        RECT 20.2 3.925 20.41 4.125 ;
        RECT 38.125 3.925 38.335 4.125 ;
        RECT 56.05 3.925 56.26 4.125 ;
        RECT 73.975 3.925 74.185 4.125 ;
        RECT 91.9 3.925 92.11 4.125 ;
      LAYER mcon ;
        RECT 15.315 11.045 15.485 11.215 ;
        RECT 15.995 11.045 16.165 11.215 ;
        RECT 16.675 11.045 16.845 11.215 ;
        RECT 17.355 11.045 17.525 11.215 ;
        RECT 18.34 2.86 18.51 3.03 ;
        RECT 18.8 2.86 18.97 3.03 ;
        RECT 19.26 2.86 19.43 3.03 ;
        RECT 19.72 2.86 19.89 3.03 ;
        RECT 20.055 4.44 20.225 4.61 ;
        RECT 20.18 2.86 20.35 3.03 ;
        RECT 20.64 2.86 20.81 3.03 ;
        RECT 21.1 2.86 21.27 3.03 ;
        RECT 21.56 2.86 21.73 3.03 ;
        RECT 21.585 3.965 21.755 4.135 ;
        RECT 22.02 2.86 22.19 3.03 ;
        RECT 22.48 2.86 22.65 3.03 ;
        RECT 22.94 2.86 23.11 3.03 ;
        RECT 23.4 2.86 23.57 3.03 ;
        RECT 23.86 2.86 24.03 3.03 ;
        RECT 24.32 2.86 24.49 3.03 ;
        RECT 24.78 2.86 24.95 3.03 ;
        RECT 25.24 2.86 25.41 3.03 ;
        RECT 25.7 2.86 25.87 3.03 ;
        RECT 26.16 2.86 26.33 3.03 ;
        RECT 26.345 11.045 26.515 11.215 ;
        RECT 26.62 2.86 26.79 3.03 ;
        RECT 27.025 11.045 27.195 11.215 ;
        RECT 27.08 2.86 27.25 3.03 ;
        RECT 27.28 8.755 27.45 8.925 ;
        RECT 27.54 2.86 27.71 3.03 ;
        RECT 27.705 11.045 27.875 11.215 ;
        RECT 28 2.86 28.17 3.03 ;
        RECT 28.385 11.045 28.555 11.215 ;
        RECT 28.46 2.86 28.63 3.03 ;
        RECT 28.92 2.86 29.09 3.03 ;
        RECT 29.38 2.86 29.55 3.03 ;
        RECT 29.84 2.86 30.01 3.03 ;
        RECT 31.105 11.045 31.275 11.215 ;
        RECT 31.105 1.395 31.275 1.565 ;
        RECT 31.785 11.045 31.955 11.215 ;
        RECT 31.785 1.395 31.955 1.565 ;
        RECT 32.465 11.045 32.635 11.215 ;
        RECT 32.465 1.395 32.635 1.565 ;
        RECT 33.145 11.045 33.315 11.215 ;
        RECT 33.145 1.395 33.315 1.565 ;
        RECT 33.85 11.045 34.02 11.215 ;
        RECT 33.85 1.395 34.02 1.565 ;
        RECT 34.835 1.395 35.005 1.565 ;
        RECT 34.84 11.045 35.01 11.215 ;
        RECT 36.265 2.86 36.435 3.03 ;
        RECT 36.725 2.86 36.895 3.03 ;
        RECT 37.185 2.86 37.355 3.03 ;
        RECT 37.645 2.86 37.815 3.03 ;
        RECT 37.98 4.44 38.15 4.61 ;
        RECT 38.105 2.86 38.275 3.03 ;
        RECT 38.565 2.86 38.735 3.03 ;
        RECT 39.025 2.86 39.195 3.03 ;
        RECT 39.485 2.86 39.655 3.03 ;
        RECT 39.51 3.965 39.68 4.135 ;
        RECT 39.945 2.86 40.115 3.03 ;
        RECT 40.405 2.86 40.575 3.03 ;
        RECT 40.865 2.86 41.035 3.03 ;
        RECT 41.325 2.86 41.495 3.03 ;
        RECT 41.785 2.86 41.955 3.03 ;
        RECT 42.245 2.86 42.415 3.03 ;
        RECT 42.705 2.86 42.875 3.03 ;
        RECT 43.165 2.86 43.335 3.03 ;
        RECT 43.625 2.86 43.795 3.03 ;
        RECT 44.085 2.86 44.255 3.03 ;
        RECT 44.27 11.045 44.44 11.215 ;
        RECT 44.545 2.86 44.715 3.03 ;
        RECT 44.95 11.045 45.12 11.215 ;
        RECT 45.005 2.86 45.175 3.03 ;
        RECT 45.205 8.755 45.375 8.925 ;
        RECT 45.465 2.86 45.635 3.03 ;
        RECT 45.63 11.045 45.8 11.215 ;
        RECT 45.925 2.86 46.095 3.03 ;
        RECT 46.31 11.045 46.48 11.215 ;
        RECT 46.385 2.86 46.555 3.03 ;
        RECT 46.845 2.86 47.015 3.03 ;
        RECT 47.305 2.86 47.475 3.03 ;
        RECT 47.765 2.86 47.935 3.03 ;
        RECT 49.03 11.045 49.2 11.215 ;
        RECT 49.03 1.395 49.2 1.565 ;
        RECT 49.71 11.045 49.88 11.215 ;
        RECT 49.71 1.395 49.88 1.565 ;
        RECT 50.39 11.045 50.56 11.215 ;
        RECT 50.39 1.395 50.56 1.565 ;
        RECT 51.07 11.045 51.24 11.215 ;
        RECT 51.07 1.395 51.24 1.565 ;
        RECT 51.775 11.045 51.945 11.215 ;
        RECT 51.775 1.395 51.945 1.565 ;
        RECT 52.76 1.395 52.93 1.565 ;
        RECT 52.765 11.045 52.935 11.215 ;
        RECT 54.19 2.86 54.36 3.03 ;
        RECT 54.65 2.86 54.82 3.03 ;
        RECT 55.11 2.86 55.28 3.03 ;
        RECT 55.57 2.86 55.74 3.03 ;
        RECT 55.905 4.44 56.075 4.61 ;
        RECT 56.03 2.86 56.2 3.03 ;
        RECT 56.49 2.86 56.66 3.03 ;
        RECT 56.95 2.86 57.12 3.03 ;
        RECT 57.41 2.86 57.58 3.03 ;
        RECT 57.435 3.965 57.605 4.135 ;
        RECT 57.87 2.86 58.04 3.03 ;
        RECT 58.33 2.86 58.5 3.03 ;
        RECT 58.79 2.86 58.96 3.03 ;
        RECT 59.25 2.86 59.42 3.03 ;
        RECT 59.71 2.86 59.88 3.03 ;
        RECT 60.17 2.86 60.34 3.03 ;
        RECT 60.63 2.86 60.8 3.03 ;
        RECT 61.09 2.86 61.26 3.03 ;
        RECT 61.55 2.86 61.72 3.03 ;
        RECT 62.01 2.86 62.18 3.03 ;
        RECT 62.195 11.045 62.365 11.215 ;
        RECT 62.47 2.86 62.64 3.03 ;
        RECT 62.875 11.045 63.045 11.215 ;
        RECT 62.93 2.86 63.1 3.03 ;
        RECT 63.13 8.755 63.3 8.925 ;
        RECT 63.39 2.86 63.56 3.03 ;
        RECT 63.555 11.045 63.725 11.215 ;
        RECT 63.85 2.86 64.02 3.03 ;
        RECT 64.235 11.045 64.405 11.215 ;
        RECT 64.31 2.86 64.48 3.03 ;
        RECT 64.77 2.86 64.94 3.03 ;
        RECT 65.23 2.86 65.4 3.03 ;
        RECT 65.69 2.86 65.86 3.03 ;
        RECT 66.955 11.045 67.125 11.215 ;
        RECT 66.955 1.395 67.125 1.565 ;
        RECT 67.635 11.045 67.805 11.215 ;
        RECT 67.635 1.395 67.805 1.565 ;
        RECT 68.315 11.045 68.485 11.215 ;
        RECT 68.315 1.395 68.485 1.565 ;
        RECT 68.995 11.045 69.165 11.215 ;
        RECT 68.995 1.395 69.165 1.565 ;
        RECT 69.7 11.045 69.87 11.215 ;
        RECT 69.7 1.395 69.87 1.565 ;
        RECT 70.685 1.395 70.855 1.565 ;
        RECT 70.69 11.045 70.86 11.215 ;
        RECT 72.115 2.86 72.285 3.03 ;
        RECT 72.575 2.86 72.745 3.03 ;
        RECT 73.035 2.86 73.205 3.03 ;
        RECT 73.495 2.86 73.665 3.03 ;
        RECT 73.83 4.44 74 4.61 ;
        RECT 73.955 2.86 74.125 3.03 ;
        RECT 74.415 2.86 74.585 3.03 ;
        RECT 74.875 2.86 75.045 3.03 ;
        RECT 75.335 2.86 75.505 3.03 ;
        RECT 75.36 3.965 75.53 4.135 ;
        RECT 75.795 2.86 75.965 3.03 ;
        RECT 76.255 2.86 76.425 3.03 ;
        RECT 76.715 2.86 76.885 3.03 ;
        RECT 77.175 2.86 77.345 3.03 ;
        RECT 77.635 2.86 77.805 3.03 ;
        RECT 78.095 2.86 78.265 3.03 ;
        RECT 78.555 2.86 78.725 3.03 ;
        RECT 79.015 2.86 79.185 3.03 ;
        RECT 79.475 2.86 79.645 3.03 ;
        RECT 79.935 2.86 80.105 3.03 ;
        RECT 80.12 11.045 80.29 11.215 ;
        RECT 80.395 2.86 80.565 3.03 ;
        RECT 80.8 11.045 80.97 11.215 ;
        RECT 80.855 2.86 81.025 3.03 ;
        RECT 81.055 8.755 81.225 8.925 ;
        RECT 81.315 2.86 81.485 3.03 ;
        RECT 81.48 11.045 81.65 11.215 ;
        RECT 81.775 2.86 81.945 3.03 ;
        RECT 82.16 11.045 82.33 11.215 ;
        RECT 82.235 2.86 82.405 3.03 ;
        RECT 82.695 2.86 82.865 3.03 ;
        RECT 83.155 2.86 83.325 3.03 ;
        RECT 83.615 2.86 83.785 3.03 ;
        RECT 84.88 11.045 85.05 11.215 ;
        RECT 84.88 1.395 85.05 1.565 ;
        RECT 85.56 11.045 85.73 11.215 ;
        RECT 85.56 1.395 85.73 1.565 ;
        RECT 86.24 11.045 86.41 11.215 ;
        RECT 86.24 1.395 86.41 1.565 ;
        RECT 86.92 11.045 87.09 11.215 ;
        RECT 86.92 1.395 87.09 1.565 ;
        RECT 87.625 11.045 87.795 11.215 ;
        RECT 87.625 1.395 87.795 1.565 ;
        RECT 88.61 1.395 88.78 1.565 ;
        RECT 88.615 11.045 88.785 11.215 ;
        RECT 90.04 2.86 90.21 3.03 ;
        RECT 90.5 2.86 90.67 3.03 ;
        RECT 90.96 2.86 91.13 3.03 ;
        RECT 91.42 2.86 91.59 3.03 ;
        RECT 91.755 4.44 91.925 4.61 ;
        RECT 91.88 2.86 92.05 3.03 ;
        RECT 92.34 2.86 92.51 3.03 ;
        RECT 92.8 2.86 92.97 3.03 ;
        RECT 93.26 2.86 93.43 3.03 ;
        RECT 93.285 3.965 93.455 4.135 ;
        RECT 93.72 2.86 93.89 3.03 ;
        RECT 94.18 2.86 94.35 3.03 ;
        RECT 94.64 2.86 94.81 3.03 ;
        RECT 95.1 2.86 95.27 3.03 ;
        RECT 95.56 2.86 95.73 3.03 ;
        RECT 96.02 2.86 96.19 3.03 ;
        RECT 96.48 2.86 96.65 3.03 ;
        RECT 96.94 2.86 97.11 3.03 ;
        RECT 97.4 2.86 97.57 3.03 ;
        RECT 97.86 2.86 98.03 3.03 ;
        RECT 98.045 11.045 98.215 11.215 ;
        RECT 98.32 2.86 98.49 3.03 ;
        RECT 98.725 11.045 98.895 11.215 ;
        RECT 98.78 2.86 98.95 3.03 ;
        RECT 98.98 8.755 99.15 8.925 ;
        RECT 99.24 2.86 99.41 3.03 ;
        RECT 99.405 11.045 99.575 11.215 ;
        RECT 99.7 2.86 99.87 3.03 ;
        RECT 100.085 11.045 100.255 11.215 ;
        RECT 100.16 2.86 100.33 3.03 ;
        RECT 100.62 2.86 100.79 3.03 ;
        RECT 101.08 2.86 101.25 3.03 ;
        RECT 101.54 2.86 101.71 3.03 ;
        RECT 102.805 11.045 102.975 11.215 ;
        RECT 102.805 1.395 102.975 1.565 ;
        RECT 103.485 11.045 103.655 11.215 ;
        RECT 103.485 1.395 103.655 1.565 ;
        RECT 104.165 11.045 104.335 11.215 ;
        RECT 104.165 1.395 104.335 1.565 ;
        RECT 104.845 11.045 105.015 11.215 ;
        RECT 104.845 1.395 105.015 1.565 ;
        RECT 105.55 11.045 105.72 11.215 ;
        RECT 105.55 1.395 105.72 1.565 ;
        RECT 106.535 1.395 106.705 1.565 ;
        RECT 106.54 11.045 106.71 11.215 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 106.805 7.345 107.155 12.61 ;
      RECT 106.79 7.345 107.17 7.725 ;
      RECT 99.24 9.49 99.615 9.86 ;
      RECT 99.275 7.36 99.585 9.86 ;
      RECT 99.275 7.36 102.37 7.67 ;
      RECT 102.06 2.805 102.37 7.67 ;
      RECT 102.07 2.435 102.445 2.805 ;
      RECT 102.07 2.42 102.38 2.805 ;
      RECT 99.2 4.98 99.755 5.31 ;
      RECT 99.2 3.315 99.5 5.31 ;
      RECT 95.265 4.42 95.82 4.75 ;
      RECT 95.52 3.315 95.82 4.75 ;
      RECT 96.315 3.18 96.465 3.83 ;
      RECT 95.52 3.315 99.5 3.615 ;
      RECT 94.025 2.255 94.325 5.205 ;
      RECT 94.025 3.86 94.755 4.19 ;
      RECT 93.98 2.255 94.355 2.625 ;
      RECT 92.585 4.42 93.315 4.75 ;
      RECT 92.59 2.255 92.89 4.75 ;
      RECT 90.475 3.86 91.205 4.19 ;
      RECT 90.62 2.225 90.92 4.19 ;
      RECT 92.545 2.255 92.92 2.625 ;
      RECT 90.575 2.225 90.95 2.595 ;
      RECT 90.575 2.265 92.92 2.565 ;
      RECT 88.88 7.345 89.23 12.61 ;
      RECT 88.865 7.345 89.245 7.725 ;
      RECT 81.315 9.49 81.69 9.86 ;
      RECT 81.35 7.36 81.66 9.86 ;
      RECT 81.35 7.36 84.445 7.67 ;
      RECT 84.135 2.805 84.445 7.67 ;
      RECT 84.145 2.435 84.52 2.805 ;
      RECT 84.145 2.42 84.455 2.805 ;
      RECT 81.275 4.98 81.83 5.31 ;
      RECT 81.275 3.315 81.575 5.31 ;
      RECT 77.34 4.42 77.895 4.75 ;
      RECT 77.595 3.315 77.895 4.75 ;
      RECT 78.39 3.18 78.54 3.83 ;
      RECT 77.595 3.315 81.575 3.615 ;
      RECT 76.1 2.255 76.4 5.205 ;
      RECT 76.1 3.86 76.83 4.19 ;
      RECT 76.055 2.255 76.43 2.625 ;
      RECT 74.66 4.42 75.39 4.75 ;
      RECT 74.665 2.255 74.965 4.75 ;
      RECT 72.55 3.86 73.28 4.19 ;
      RECT 72.695 2.225 72.995 4.19 ;
      RECT 74.62 2.255 74.995 2.625 ;
      RECT 72.65 2.225 73.025 2.595 ;
      RECT 72.65 2.265 74.995 2.565 ;
      RECT 70.955 7.345 71.305 12.61 ;
      RECT 70.94 7.345 71.32 7.725 ;
      RECT 63.39 9.49 63.765 9.86 ;
      RECT 63.425 7.36 63.735 9.86 ;
      RECT 63.425 7.36 66.52 7.67 ;
      RECT 66.21 2.805 66.52 7.67 ;
      RECT 66.22 2.435 66.595 2.805 ;
      RECT 66.22 2.42 66.53 2.805 ;
      RECT 63.35 4.98 63.905 5.31 ;
      RECT 63.35 3.315 63.65 5.31 ;
      RECT 59.415 4.42 59.97 4.75 ;
      RECT 59.67 3.315 59.97 4.75 ;
      RECT 60.465 3.18 60.615 3.83 ;
      RECT 59.67 3.315 63.65 3.615 ;
      RECT 58.175 2.255 58.475 5.205 ;
      RECT 58.175 3.86 58.905 4.19 ;
      RECT 58.13 2.255 58.505 2.625 ;
      RECT 56.735 4.42 57.465 4.75 ;
      RECT 56.74 2.255 57.04 4.75 ;
      RECT 54.625 3.86 55.355 4.19 ;
      RECT 54.77 2.225 55.07 4.19 ;
      RECT 56.695 2.255 57.07 2.625 ;
      RECT 54.725 2.225 55.1 2.595 ;
      RECT 54.725 2.265 57.07 2.565 ;
      RECT 53.03 7.345 53.38 12.61 ;
      RECT 53.015 7.345 53.395 7.725 ;
      RECT 45.465 9.49 45.84 9.86 ;
      RECT 45.5 7.36 45.81 9.86 ;
      RECT 45.5 7.36 48.595 7.67 ;
      RECT 48.285 2.805 48.595 7.67 ;
      RECT 48.295 2.435 48.67 2.805 ;
      RECT 48.295 2.42 48.605 2.805 ;
      RECT 45.425 4.98 45.98 5.31 ;
      RECT 45.425 3.315 45.725 5.31 ;
      RECT 41.49 4.42 42.045 4.75 ;
      RECT 41.745 3.315 42.045 4.75 ;
      RECT 42.54 3.18 42.69 3.83 ;
      RECT 41.745 3.315 45.725 3.615 ;
      RECT 40.25 2.255 40.55 5.205 ;
      RECT 40.25 3.86 40.98 4.19 ;
      RECT 40.205 2.255 40.58 2.625 ;
      RECT 38.81 4.42 39.54 4.75 ;
      RECT 38.815 2.255 39.115 4.75 ;
      RECT 36.7 3.86 37.43 4.19 ;
      RECT 36.845 2.225 37.145 4.19 ;
      RECT 38.77 2.255 39.145 2.625 ;
      RECT 36.8 2.225 37.175 2.595 ;
      RECT 36.8 2.265 39.145 2.565 ;
      RECT 35.105 7.345 35.455 12.61 ;
      RECT 35.09 7.345 35.47 7.725 ;
      RECT 27.54 9.49 27.915 9.86 ;
      RECT 27.575 7.36 27.885 9.86 ;
      RECT 27.575 7.36 30.67 7.67 ;
      RECT 30.36 2.805 30.67 7.67 ;
      RECT 30.37 2.435 30.745 2.805 ;
      RECT 30.37 2.42 30.68 2.805 ;
      RECT 27.5 4.98 28.055 5.31 ;
      RECT 27.5 3.315 27.8 5.31 ;
      RECT 23.565 4.42 24.12 4.75 ;
      RECT 23.82 3.315 24.12 4.75 ;
      RECT 24.615 3.18 24.765 3.83 ;
      RECT 23.82 3.315 27.8 3.615 ;
      RECT 22.325 2.255 22.625 5.205 ;
      RECT 22.325 3.86 23.055 4.19 ;
      RECT 22.28 2.255 22.655 2.625 ;
      RECT 20.885 4.42 21.615 4.75 ;
      RECT 20.89 2.255 21.19 4.75 ;
      RECT 18.775 3.86 19.505 4.19 ;
      RECT 18.92 2.225 19.22 4.19 ;
      RECT 20.845 2.255 21.22 2.625 ;
      RECT 18.875 2.225 19.25 2.595 ;
      RECT 18.875 2.265 21.22 2.565 ;
      RECT 100.385 3.3 101.115 3.63 ;
      RECT 98.165 4.98 98.895 5.31 ;
      RECT 96.465 4.98 97.195 5.31 ;
      RECT 90.145 4.98 90.875 5.31 ;
      RECT 82.46 3.3 83.19 3.63 ;
      RECT 80.24 4.98 80.97 5.31 ;
      RECT 78.54 4.98 79.27 5.31 ;
      RECT 72.22 4.98 72.95 5.31 ;
      RECT 64.535 3.3 65.265 3.63 ;
      RECT 62.315 4.98 63.045 5.31 ;
      RECT 60.615 4.98 61.345 5.31 ;
      RECT 54.295 4.98 55.025 5.31 ;
      RECT 46.61 3.3 47.34 3.63 ;
      RECT 44.39 4.98 45.12 5.31 ;
      RECT 42.69 4.98 43.42 5.31 ;
      RECT 36.37 4.98 37.1 5.31 ;
      RECT 28.685 3.3 29.415 3.63 ;
      RECT 26.465 4.98 27.195 5.31 ;
      RECT 24.765 4.98 25.495 5.31 ;
      RECT 18.445 4.98 19.175 5.31 ;
    LAYER via2 ;
      RECT 106.88 7.435 107.08 7.635 ;
      RECT 102.16 2.52 102.36 2.72 ;
      RECT 100.45 3.365 100.65 3.565 ;
      RECT 99.49 5.045 99.69 5.245 ;
      RECT 99.33 9.575 99.53 9.775 ;
      RECT 98.49 5.045 98.69 5.245 ;
      RECT 96.53 5.045 96.73 5.245 ;
      RECT 95.33 4.485 95.53 4.685 ;
      RECT 94.09 3.925 94.29 4.125 ;
      RECT 94.07 2.34 94.27 2.54 ;
      RECT 92.65 4.485 92.85 4.685 ;
      RECT 92.635 2.335 92.835 2.535 ;
      RECT 90.69 3.925 90.89 4.125 ;
      RECT 90.665 2.31 90.865 2.51 ;
      RECT 90.21 5.045 90.41 5.245 ;
      RECT 88.955 7.435 89.155 7.635 ;
      RECT 84.235 2.52 84.435 2.72 ;
      RECT 82.525 3.365 82.725 3.565 ;
      RECT 81.565 5.045 81.765 5.245 ;
      RECT 81.405 9.575 81.605 9.775 ;
      RECT 80.565 5.045 80.765 5.245 ;
      RECT 78.605 5.045 78.805 5.245 ;
      RECT 77.405 4.485 77.605 4.685 ;
      RECT 76.165 3.925 76.365 4.125 ;
      RECT 76.145 2.34 76.345 2.54 ;
      RECT 74.725 4.485 74.925 4.685 ;
      RECT 74.71 2.335 74.91 2.535 ;
      RECT 72.765 3.925 72.965 4.125 ;
      RECT 72.74 2.31 72.94 2.51 ;
      RECT 72.285 5.045 72.485 5.245 ;
      RECT 71.03 7.435 71.23 7.635 ;
      RECT 66.31 2.52 66.51 2.72 ;
      RECT 64.6 3.365 64.8 3.565 ;
      RECT 63.64 5.045 63.84 5.245 ;
      RECT 63.48 9.575 63.68 9.775 ;
      RECT 62.64 5.045 62.84 5.245 ;
      RECT 60.68 5.045 60.88 5.245 ;
      RECT 59.48 4.485 59.68 4.685 ;
      RECT 58.24 3.925 58.44 4.125 ;
      RECT 58.22 2.34 58.42 2.54 ;
      RECT 56.8 4.485 57 4.685 ;
      RECT 56.785 2.335 56.985 2.535 ;
      RECT 54.84 3.925 55.04 4.125 ;
      RECT 54.815 2.31 55.015 2.51 ;
      RECT 54.36 5.045 54.56 5.245 ;
      RECT 53.105 7.435 53.305 7.635 ;
      RECT 48.385 2.52 48.585 2.72 ;
      RECT 46.675 3.365 46.875 3.565 ;
      RECT 45.715 5.045 45.915 5.245 ;
      RECT 45.555 9.575 45.755 9.775 ;
      RECT 44.715 5.045 44.915 5.245 ;
      RECT 42.755 5.045 42.955 5.245 ;
      RECT 41.555 4.485 41.755 4.685 ;
      RECT 40.315 3.925 40.515 4.125 ;
      RECT 40.295 2.34 40.495 2.54 ;
      RECT 38.875 4.485 39.075 4.685 ;
      RECT 38.86 2.335 39.06 2.535 ;
      RECT 36.915 3.925 37.115 4.125 ;
      RECT 36.89 2.31 37.09 2.51 ;
      RECT 36.435 5.045 36.635 5.245 ;
      RECT 35.18 7.435 35.38 7.635 ;
      RECT 30.46 2.52 30.66 2.72 ;
      RECT 28.75 3.365 28.95 3.565 ;
      RECT 27.79 5.045 27.99 5.245 ;
      RECT 27.63 9.575 27.83 9.775 ;
      RECT 26.79 5.045 26.99 5.245 ;
      RECT 24.83 5.045 25.03 5.245 ;
      RECT 23.63 4.485 23.83 4.685 ;
      RECT 22.39 3.925 22.59 4.125 ;
      RECT 22.37 2.34 22.57 2.54 ;
      RECT 20.95 4.485 21.15 4.685 ;
      RECT 20.935 2.335 21.135 2.535 ;
      RECT 18.99 3.925 19.19 4.125 ;
      RECT 18.965 2.31 19.165 2.51 ;
      RECT 18.51 5.045 18.71 5.245 ;
    LAYER met2 ;
      RECT 16.24 10.835 107.06 11.005 ;
      RECT 106.89 9.71 107.06 11.005 ;
      RECT 16.24 8.69 16.41 11.005 ;
      RECT 106.86 9.71 107.21 10.06 ;
      RECT 16.185 8.69 16.475 9.04 ;
      RECT 103.705 8.66 104.025 8.98 ;
      RECT 103.735 8.13 103.905 8.98 ;
      RECT 103.735 8.13 103.91 8.48 ;
      RECT 103.735 8.13 104.71 8.305 ;
      RECT 104.535 3.26 104.71 8.305 ;
      RECT 104.48 3.26 104.83 3.61 ;
      RECT 104.505 9.09 104.83 9.415 ;
      RECT 103.39 9.18 104.83 9.35 ;
      RECT 103.39 3.69 103.55 9.35 ;
      RECT 103.705 3.66 104.025 3.98 ;
      RECT 103.39 3.69 104.025 3.86 ;
      RECT 102.07 2.435 102.445 2.805 ;
      RECT 93.98 2.255 94.355 2.625 ;
      RECT 92.545 2.255 92.92 2.625 ;
      RECT 92.545 2.375 102.375 2.545 ;
      RECT 98.49 5.655 102.345 5.825 ;
      RECT 102.175 4.72 102.345 5.825 ;
      RECT 98.49 4.965 98.66 5.825 ;
      RECT 98.45 5.005 98.73 5.285 ;
      RECT 98.47 4.965 98.73 5.285 ;
      RECT 98.11 4.92 98.215 5.18 ;
      RECT 102.085 4.725 102.435 5.075 ;
      RECT 97.965 3.41 98.055 3.67 ;
      RECT 98.505 4.475 98.51 4.515 ;
      RECT 98.5 4.465 98.505 4.6 ;
      RECT 98.495 4.455 98.5 4.693 ;
      RECT 98.485 4.435 98.495 4.749 ;
      RECT 98.405 4.363 98.485 4.829 ;
      RECT 98.44 5.007 98.45 5.232 ;
      RECT 98.435 5.004 98.44 5.227 ;
      RECT 98.42 5.001 98.435 5.22 ;
      RECT 98.385 4.995 98.42 5.202 ;
      RECT 98.4 4.298 98.405 4.903 ;
      RECT 98.38 4.249 98.4 4.918 ;
      RECT 98.37 4.982 98.385 5.185 ;
      RECT 98.375 4.191 98.38 4.933 ;
      RECT 98.37 4.169 98.375 4.943 ;
      RECT 98.335 4.079 98.37 5.18 ;
      RECT 98.32 3.957 98.335 5.18 ;
      RECT 98.315 3.91 98.32 5.18 ;
      RECT 98.29 3.835 98.315 5.18 ;
      RECT 98.275 3.75 98.29 5.18 ;
      RECT 98.27 3.697 98.275 5.18 ;
      RECT 98.265 3.677 98.27 5.18 ;
      RECT 98.26 3.652 98.265 4.414 ;
      RECT 98.245 4.612 98.265 5.18 ;
      RECT 98.255 3.63 98.26 4.391 ;
      RECT 98.245 3.582 98.255 4.356 ;
      RECT 98.24 3.545 98.245 4.322 ;
      RECT 98.24 4.692 98.245 5.18 ;
      RECT 98.225 3.522 98.24 4.277 ;
      RECT 98.22 4.79 98.24 5.18 ;
      RECT 98.17 3.41 98.225 4.119 ;
      RECT 98.215 4.912 98.22 5.18 ;
      RECT 98.155 3.41 98.17 3.958 ;
      RECT 98.15 3.41 98.155 3.91 ;
      RECT 98.145 3.41 98.15 3.898 ;
      RECT 98.1 3.41 98.145 3.835 ;
      RECT 98.075 3.41 98.1 3.753 ;
      RECT 98.06 3.41 98.075 3.705 ;
      RECT 98.055 3.41 98.06 3.675 ;
      RECT 100.445 3.455 100.705 3.715 ;
      RECT 100.44 3.455 100.705 3.663 ;
      RECT 100.435 3.455 100.705 3.633 ;
      RECT 100.41 3.325 100.69 3.605 ;
      RECT 88.915 9.095 89.265 9.445 ;
      RECT 100.16 9.05 100.51 9.4 ;
      RECT 88.915 9.125 100.51 9.325 ;
      RECT 99.45 5.005 99.73 5.285 ;
      RECT 99.49 4.96 99.755 5.22 ;
      RECT 99.48 4.995 99.755 5.22 ;
      RECT 99.485 4.98 99.73 5.285 ;
      RECT 99.49 4.957 99.7 5.285 ;
      RECT 99.49 4.955 99.685 5.285 ;
      RECT 99.53 4.945 99.685 5.285 ;
      RECT 99.5 4.95 99.685 5.285 ;
      RECT 99.53 4.942 99.63 5.285 ;
      RECT 99.555 4.935 99.63 5.285 ;
      RECT 99.535 4.937 99.63 5.285 ;
      RECT 98.865 4.45 99.125 4.71 ;
      RECT 98.915 4.442 99.105 4.71 ;
      RECT 98.92 4.362 99.105 4.71 ;
      RECT 99.04 3.75 99.105 4.71 ;
      RECT 98.945 4.147 99.105 4.71 ;
      RECT 99.02 3.835 99.105 4.71 ;
      RECT 99.055 3.46 99.191 4.188 ;
      RECT 99 3.957 99.191 4.188 ;
      RECT 99.015 3.897 99.105 4.71 ;
      RECT 99.055 3.46 99.215 3.853 ;
      RECT 99.055 3.46 99.225 3.75 ;
      RECT 99.045 3.46 99.305 3.72 ;
      RECT 97.38 4.86 97.425 5.12 ;
      RECT 97.285 3.395 97.43 3.655 ;
      RECT 97.79 4.017 97.8 4.108 ;
      RECT 97.775 3.955 97.79 4.164 ;
      RECT 97.77 3.902 97.775 4.21 ;
      RECT 97.72 3.849 97.77 4.336 ;
      RECT 97.715 3.804 97.72 4.483 ;
      RECT 97.705 3.792 97.715 4.525 ;
      RECT 97.67 3.756 97.705 4.63 ;
      RECT 97.665 3.724 97.67 4.736 ;
      RECT 97.65 3.706 97.665 4.781 ;
      RECT 97.645 3.689 97.65 4.015 ;
      RECT 97.64 4.07 97.65 4.838 ;
      RECT 97.635 3.675 97.645 3.988 ;
      RECT 97.63 4.125 97.64 5.12 ;
      RECT 97.625 3.661 97.635 3.973 ;
      RECT 97.625 4.175 97.63 5.12 ;
      RECT 97.61 3.638 97.625 3.953 ;
      RECT 97.59 4.297 97.625 5.12 ;
      RECT 97.605 3.62 97.61 3.935 ;
      RECT 97.6 3.612 97.605 3.925 ;
      RECT 97.57 3.58 97.6 3.889 ;
      RECT 97.58 4.425 97.59 5.12 ;
      RECT 97.575 4.452 97.58 5.12 ;
      RECT 97.57 4.502 97.575 5.12 ;
      RECT 97.56 3.546 97.57 3.854 ;
      RECT 97.52 4.57 97.57 5.12 ;
      RECT 97.545 3.523 97.56 3.83 ;
      RECT 97.52 3.395 97.545 3.793 ;
      RECT 97.515 3.395 97.52 3.765 ;
      RECT 97.485 4.67 97.52 5.12 ;
      RECT 97.51 3.395 97.515 3.758 ;
      RECT 97.505 3.395 97.51 3.748 ;
      RECT 97.49 3.395 97.505 3.733 ;
      RECT 97.475 3.395 97.49 3.705 ;
      RECT 97.44 4.775 97.485 5.12 ;
      RECT 97.46 3.395 97.475 3.678 ;
      RECT 97.43 3.395 97.46 3.663 ;
      RECT 97.425 4.847 97.44 5.12 ;
      RECT 97.35 3.93 97.39 4.19 ;
      RECT 97.125 3.877 97.13 4.135 ;
      RECT 93.08 3.355 93.34 3.615 ;
      RECT 93.08 3.38 93.355 3.595 ;
      RECT 95.47 3.205 95.475 3.35 ;
      RECT 97.34 3.925 97.35 4.19 ;
      RECT 97.32 3.917 97.34 4.19 ;
      RECT 97.302 3.913 97.32 4.19 ;
      RECT 97.216 3.902 97.302 4.19 ;
      RECT 97.13 3.885 97.216 4.19 ;
      RECT 97.075 3.872 97.125 4.12 ;
      RECT 97.041 3.864 97.075 4.095 ;
      RECT 96.955 3.853 97.041 4.06 ;
      RECT 96.92 3.83 96.955 4.025 ;
      RECT 96.91 3.792 96.92 4.011 ;
      RECT 96.905 3.765 96.91 4.007 ;
      RECT 96.9 3.752 96.905 4.004 ;
      RECT 96.89 3.732 96.9 4 ;
      RECT 96.885 3.707 96.89 3.996 ;
      RECT 96.86 3.662 96.885 3.99 ;
      RECT 96.85 3.603 96.86 3.982 ;
      RECT 96.84 3.571 96.85 3.973 ;
      RECT 96.82 3.523 96.84 3.953 ;
      RECT 96.815 3.483 96.82 3.923 ;
      RECT 96.8 3.457 96.815 3.897 ;
      RECT 96.795 3.435 96.8 3.873 ;
      RECT 96.78 3.407 96.795 3.849 ;
      RECT 96.765 3.38 96.78 3.813 ;
      RECT 96.75 3.357 96.765 3.775 ;
      RECT 96.745 3.347 96.75 3.75 ;
      RECT 96.735 3.34 96.745 3.733 ;
      RECT 96.72 3.327 96.735 3.703 ;
      RECT 96.715 3.317 96.72 3.678 ;
      RECT 96.71 3.312 96.715 3.665 ;
      RECT 96.7 3.305 96.71 3.645 ;
      RECT 96.695 3.298 96.7 3.63 ;
      RECT 96.67 3.291 96.695 3.588 ;
      RECT 96.655 3.281 96.67 3.538 ;
      RECT 96.645 3.276 96.655 3.508 ;
      RECT 96.635 3.272 96.645 3.483 ;
      RECT 96.62 3.269 96.635 3.473 ;
      RECT 96.57 3.266 96.62 3.458 ;
      RECT 96.55 3.264 96.57 3.443 ;
      RECT 96.501 3.262 96.55 3.438 ;
      RECT 96.415 3.258 96.501 3.433 ;
      RECT 96.376 3.255 96.415 3.429 ;
      RECT 96.29 3.251 96.376 3.424 ;
      RECT 96.24 3.248 96.29 3.418 ;
      RECT 96.191 3.245 96.24 3.413 ;
      RECT 96.105 3.242 96.191 3.408 ;
      RECT 96.101 3.24 96.105 3.405 ;
      RECT 96.015 3.237 96.101 3.4 ;
      RECT 95.966 3.233 96.015 3.393 ;
      RECT 95.88 3.23 95.966 3.388 ;
      RECT 95.856 3.227 95.88 3.384 ;
      RECT 95.77 3.225 95.856 3.379 ;
      RECT 95.705 3.221 95.77 3.372 ;
      RECT 95.702 3.22 95.705 3.369 ;
      RECT 95.616 3.217 95.702 3.366 ;
      RECT 95.53 3.211 95.616 3.359 ;
      RECT 95.5 3.207 95.53 3.355 ;
      RECT 95.475 3.205 95.5 3.353 ;
      RECT 95.42 3.202 95.47 3.35 ;
      RECT 95.34 3.201 95.42 3.35 ;
      RECT 95.285 3.203 95.34 3.353 ;
      RECT 95.27 3.204 95.285 3.357 ;
      RECT 95.215 3.212 95.27 3.367 ;
      RECT 95.185 3.22 95.215 3.38 ;
      RECT 95.166 3.221 95.185 3.386 ;
      RECT 95.08 3.224 95.166 3.391 ;
      RECT 95.01 3.229 95.08 3.4 ;
      RECT 94.991 3.232 95.01 3.406 ;
      RECT 94.905 3.236 94.991 3.411 ;
      RECT 94.865 3.24 94.905 3.418 ;
      RECT 94.856 3.242 94.865 3.421 ;
      RECT 94.77 3.246 94.856 3.426 ;
      RECT 94.767 3.249 94.77 3.43 ;
      RECT 94.681 3.252 94.767 3.434 ;
      RECT 94.595 3.258 94.681 3.442 ;
      RECT 94.571 3.262 94.595 3.446 ;
      RECT 94.485 3.266 94.571 3.451 ;
      RECT 94.44 3.271 94.485 3.458 ;
      RECT 94.36 3.276 94.44 3.465 ;
      RECT 94.28 3.282 94.36 3.48 ;
      RECT 94.255 3.286 94.28 3.493 ;
      RECT 94.19 3.289 94.255 3.505 ;
      RECT 94.135 3.294 94.19 3.52 ;
      RECT 94.105 3.297 94.135 3.538 ;
      RECT 94.095 3.299 94.105 3.551 ;
      RECT 94.035 3.314 94.095 3.561 ;
      RECT 94.02 3.331 94.035 3.57 ;
      RECT 94.015 3.34 94.02 3.57 ;
      RECT 94.005 3.35 94.015 3.57 ;
      RECT 93.995 3.367 94.005 3.57 ;
      RECT 93.975 3.377 93.995 3.571 ;
      RECT 93.93 3.387 93.975 3.572 ;
      RECT 93.895 3.396 93.93 3.574 ;
      RECT 93.83 3.401 93.895 3.576 ;
      RECT 93.75 3.402 93.83 3.579 ;
      RECT 93.746 3.4 93.75 3.58 ;
      RECT 93.66 3.397 93.746 3.582 ;
      RECT 93.613 3.394 93.66 3.584 ;
      RECT 93.527 3.39 93.613 3.587 ;
      RECT 93.441 3.386 93.527 3.59 ;
      RECT 93.355 3.382 93.441 3.594 ;
      RECT 96.74 5.005 96.77 5.285 ;
      RECT 96.49 4.895 96.51 5.285 ;
      RECT 96.445 4.895 96.51 5.155 ;
      RECT 96.275 3.52 96.31 3.78 ;
      RECT 96.05 3.52 96.11 3.78 ;
      RECT 96.73 4.985 96.74 5.285 ;
      RECT 96.725 4.945 96.73 5.285 ;
      RECT 96.71 4.9 96.725 5.285 ;
      RECT 96.705 4.865 96.71 5.285 ;
      RECT 96.7 4.845 96.705 5.285 ;
      RECT 96.67 4.772 96.7 5.285 ;
      RECT 96.65 4.67 96.67 5.285 ;
      RECT 96.64 4.6 96.65 5.285 ;
      RECT 96.595 4.54 96.64 5.285 ;
      RECT 96.51 4.501 96.595 5.285 ;
      RECT 96.505 4.492 96.51 4.865 ;
      RECT 96.495 4.491 96.505 4.848 ;
      RECT 96.47 4.472 96.495 4.818 ;
      RECT 96.465 4.447 96.47 4.797 ;
      RECT 96.455 4.425 96.465 4.788 ;
      RECT 96.45 4.396 96.455 4.778 ;
      RECT 96.41 4.322 96.45 4.75 ;
      RECT 96.39 4.223 96.41 4.715 ;
      RECT 96.375 4.159 96.39 4.698 ;
      RECT 96.345 4.083 96.375 4.67 ;
      RECT 96.325 3.998 96.345 4.643 ;
      RECT 96.285 3.894 96.325 4.55 ;
      RECT 96.28 3.815 96.285 4.458 ;
      RECT 96.275 3.798 96.28 4.435 ;
      RECT 96.27 3.52 96.275 4.415 ;
      RECT 96.24 3.52 96.27 4.353 ;
      RECT 96.235 3.52 96.24 4.285 ;
      RECT 96.225 3.52 96.235 4.25 ;
      RECT 96.215 3.52 96.225 4.215 ;
      RECT 96.15 3.52 96.215 4.07 ;
      RECT 96.145 3.52 96.15 3.94 ;
      RECT 96.115 3.52 96.145 3.873 ;
      RECT 96.11 3.52 96.115 3.798 ;
      RECT 95.29 4.445 95.57 4.725 ;
      RECT 95.33 4.425 95.59 4.685 ;
      RECT 95.32 4.435 95.59 4.685 ;
      RECT 95.33 4.362 95.545 4.725 ;
      RECT 95.385 4.285 95.54 4.725 ;
      RECT 95.39 4.07 95.54 4.725 ;
      RECT 95.38 3.872 95.53 4.123 ;
      RECT 95.37 3.872 95.53 3.99 ;
      RECT 95.365 3.75 95.525 3.893 ;
      RECT 95.35 3.75 95.525 3.798 ;
      RECT 95.345 3.46 95.52 3.775 ;
      RECT 95.33 3.46 95.52 3.745 ;
      RECT 95.29 3.46 95.55 3.72 ;
      RECT 95.2 4.93 95.28 5.19 ;
      RECT 94.605 3.65 94.61 3.915 ;
      RECT 94.485 3.65 94.61 3.91 ;
      RECT 95.16 4.895 95.2 5.19 ;
      RECT 95.115 4.817 95.16 5.19 ;
      RECT 95.095 4.745 95.115 5.19 ;
      RECT 95.085 4.697 95.095 5.19 ;
      RECT 95.05 4.63 95.085 5.19 ;
      RECT 95.02 4.53 95.05 5.19 ;
      RECT 95 4.455 95.02 4.99 ;
      RECT 94.99 4.405 95 4.945 ;
      RECT 94.985 4.382 94.99 4.918 ;
      RECT 94.98 4.367 94.985 4.905 ;
      RECT 94.975 4.352 94.98 4.883 ;
      RECT 94.97 4.337 94.975 4.865 ;
      RECT 94.945 4.292 94.97 4.82 ;
      RECT 94.935 4.24 94.945 4.763 ;
      RECT 94.925 4.21 94.935 4.73 ;
      RECT 94.915 4.175 94.925 4.698 ;
      RECT 94.88 4.107 94.915 4.63 ;
      RECT 94.875 4.046 94.88 4.565 ;
      RECT 94.865 4.034 94.875 4.545 ;
      RECT 94.86 4.022 94.865 4.525 ;
      RECT 94.855 4.014 94.86 4.513 ;
      RECT 94.85 4.006 94.855 4.493 ;
      RECT 94.84 3.994 94.85 4.465 ;
      RECT 94.83 3.978 94.84 4.435 ;
      RECT 94.805 3.95 94.83 4.373 ;
      RECT 94.795 3.921 94.805 4.318 ;
      RECT 94.78 3.9 94.795 4.278 ;
      RECT 94.775 3.884 94.78 4.25 ;
      RECT 94.77 3.872 94.775 4.24 ;
      RECT 94.765 3.867 94.77 4.213 ;
      RECT 94.76 3.86 94.765 4.2 ;
      RECT 94.745 3.843 94.76 4.173 ;
      RECT 94.735 3.65 94.745 4.133 ;
      RECT 94.725 3.65 94.735 4.1 ;
      RECT 94.715 3.65 94.725 4.075 ;
      RECT 94.645 3.65 94.715 4.01 ;
      RECT 94.635 3.65 94.645 3.958 ;
      RECT 94.62 3.65 94.635 3.94 ;
      RECT 94.61 3.65 94.62 3.925 ;
      RECT 94.44 4.52 94.7 4.78 ;
      RECT 92.975 4.555 92.98 4.762 ;
      RECT 92.61 4.445 92.685 4.76 ;
      RECT 92.425 4.5 92.58 4.76 ;
      RECT 92.61 4.445 92.715 4.725 ;
      RECT 94.425 4.617 94.44 4.778 ;
      RECT 94.4 4.625 94.425 4.783 ;
      RECT 94.375 4.632 94.4 4.788 ;
      RECT 94.312 4.643 94.375 4.797 ;
      RECT 94.226 4.662 94.312 4.814 ;
      RECT 94.14 4.684 94.226 4.833 ;
      RECT 94.125 4.697 94.14 4.844 ;
      RECT 94.085 4.705 94.125 4.851 ;
      RECT 94.065 4.71 94.085 4.858 ;
      RECT 94.027 4.711 94.065 4.861 ;
      RECT 93.941 4.714 94.027 4.862 ;
      RECT 93.855 4.718 93.941 4.863 ;
      RECT 93.806 4.72 93.855 4.865 ;
      RECT 93.72 4.72 93.806 4.867 ;
      RECT 93.68 4.715 93.72 4.869 ;
      RECT 93.67 4.709 93.68 4.87 ;
      RECT 93.63 4.704 93.67 4.867 ;
      RECT 93.62 4.697 93.63 4.863 ;
      RECT 93.605 4.693 93.62 4.861 ;
      RECT 93.588 4.689 93.605 4.859 ;
      RECT 93.502 4.679 93.588 4.851 ;
      RECT 93.416 4.661 93.502 4.837 ;
      RECT 93.33 4.644 93.416 4.823 ;
      RECT 93.305 4.632 93.33 4.814 ;
      RECT 93.235 4.622 93.305 4.807 ;
      RECT 93.19 4.61 93.235 4.798 ;
      RECT 93.13 4.597 93.19 4.79 ;
      RECT 93.125 4.589 93.13 4.785 ;
      RECT 93.09 4.584 93.125 4.783 ;
      RECT 93.035 4.575 93.09 4.776 ;
      RECT 92.995 4.564 93.035 4.768 ;
      RECT 92.98 4.557 92.995 4.764 ;
      RECT 92.96 4.55 92.975 4.761 ;
      RECT 92.945 4.54 92.96 4.759 ;
      RECT 92.93 4.527 92.945 4.756 ;
      RECT 92.905 4.51 92.93 4.752 ;
      RECT 92.89 4.492 92.905 4.749 ;
      RECT 92.865 4.445 92.89 4.747 ;
      RECT 92.841 4.445 92.865 4.744 ;
      RECT 92.755 4.445 92.841 4.736 ;
      RECT 92.715 4.445 92.755 4.728 ;
      RECT 92.58 4.492 92.61 4.76 ;
      RECT 94.26 4.075 94.52 4.335 ;
      RECT 94.22 4.075 94.52 4.213 ;
      RECT 94.185 4.075 94.52 4.198 ;
      RECT 94.13 4.075 94.52 4.178 ;
      RECT 94.05 3.885 94.33 4.165 ;
      RECT 94.05 4.067 94.4 4.165 ;
      RECT 94.05 4.01 94.385 4.165 ;
      RECT 94.05 3.957 94.335 4.165 ;
      RECT 91.21 4.244 91.225 4.7 ;
      RECT 91.205 4.316 91.311 4.698 ;
      RECT 91.225 3.41 91.36 4.696 ;
      RECT 91.21 4.26 91.365 4.695 ;
      RECT 91.21 4.31 91.37 4.693 ;
      RECT 91.195 4.375 91.37 4.692 ;
      RECT 91.205 4.367 91.375 4.689 ;
      RECT 91.185 4.415 91.375 4.684 ;
      RECT 91.185 4.415 91.39 4.681 ;
      RECT 91.18 4.415 91.39 4.678 ;
      RECT 91.155 4.415 91.415 4.675 ;
      RECT 91.225 3.41 91.385 4.063 ;
      RECT 91.22 3.41 91.385 4.035 ;
      RECT 91.215 3.41 91.385 3.863 ;
      RECT 91.215 3.41 91.405 3.803 ;
      RECT 91.17 3.41 91.43 3.67 ;
      RECT 90.65 3.885 90.93 4.165 ;
      RECT 90.64 3.9 90.93 4.16 ;
      RECT 90.595 3.962 90.93 4.158 ;
      RECT 90.67 3.877 90.835 4.165 ;
      RECT 90.67 3.862 90.791 4.165 ;
      RECT 90.705 3.855 90.791 4.165 ;
      RECT 90.17 5.005 90.45 5.285 ;
      RECT 90.13 4.967 90.425 5.078 ;
      RECT 90.115 4.917 90.405 4.973 ;
      RECT 90.06 4.68 90.32 4.94 ;
      RECT 90.06 4.882 90.4 4.94 ;
      RECT 90.06 4.822 90.395 4.94 ;
      RECT 90.06 4.772 90.375 4.94 ;
      RECT 90.06 4.752 90.37 4.94 ;
      RECT 90.06 4.73 90.365 4.94 ;
      RECT 90.06 4.715 90.335 4.94 ;
      RECT 85.78 8.66 86.1 8.98 ;
      RECT 85.81 8.13 85.98 8.98 ;
      RECT 85.81 8.13 85.985 8.48 ;
      RECT 85.81 8.13 86.785 8.305 ;
      RECT 86.61 3.26 86.785 8.305 ;
      RECT 86.555 3.26 86.905 3.61 ;
      RECT 86.58 9.09 86.905 9.415 ;
      RECT 85.465 9.18 86.905 9.35 ;
      RECT 85.465 3.69 85.625 9.35 ;
      RECT 85.78 3.66 86.1 3.98 ;
      RECT 85.465 3.69 86.1 3.86 ;
      RECT 84.145 2.435 84.52 2.805 ;
      RECT 76.055 2.255 76.43 2.625 ;
      RECT 74.62 2.255 74.995 2.625 ;
      RECT 74.62 2.375 84.45 2.545 ;
      RECT 80.565 5.655 84.42 5.825 ;
      RECT 84.25 4.72 84.42 5.825 ;
      RECT 80.565 4.965 80.735 5.825 ;
      RECT 80.525 5.005 80.805 5.285 ;
      RECT 80.545 4.965 80.805 5.285 ;
      RECT 80.185 4.92 80.29 5.18 ;
      RECT 84.16 4.725 84.51 5.075 ;
      RECT 80.04 3.41 80.13 3.67 ;
      RECT 80.58 4.475 80.585 4.515 ;
      RECT 80.575 4.465 80.58 4.6 ;
      RECT 80.57 4.455 80.575 4.693 ;
      RECT 80.56 4.435 80.57 4.749 ;
      RECT 80.48 4.363 80.56 4.829 ;
      RECT 80.515 5.007 80.525 5.232 ;
      RECT 80.51 5.004 80.515 5.227 ;
      RECT 80.495 5.001 80.51 5.22 ;
      RECT 80.46 4.995 80.495 5.202 ;
      RECT 80.475 4.298 80.48 4.903 ;
      RECT 80.455 4.249 80.475 4.918 ;
      RECT 80.445 4.982 80.46 5.185 ;
      RECT 80.45 4.191 80.455 4.933 ;
      RECT 80.445 4.169 80.45 4.943 ;
      RECT 80.41 4.079 80.445 5.18 ;
      RECT 80.395 3.957 80.41 5.18 ;
      RECT 80.39 3.91 80.395 5.18 ;
      RECT 80.365 3.835 80.39 5.18 ;
      RECT 80.35 3.75 80.365 5.18 ;
      RECT 80.345 3.697 80.35 5.18 ;
      RECT 80.34 3.677 80.345 5.18 ;
      RECT 80.335 3.652 80.34 4.414 ;
      RECT 80.32 4.612 80.34 5.18 ;
      RECT 80.33 3.63 80.335 4.391 ;
      RECT 80.32 3.582 80.33 4.356 ;
      RECT 80.315 3.545 80.32 4.322 ;
      RECT 80.315 4.692 80.32 5.18 ;
      RECT 80.3 3.522 80.315 4.277 ;
      RECT 80.295 4.79 80.315 5.18 ;
      RECT 80.245 3.41 80.3 4.119 ;
      RECT 80.29 4.912 80.295 5.18 ;
      RECT 80.23 3.41 80.245 3.958 ;
      RECT 80.225 3.41 80.23 3.91 ;
      RECT 80.22 3.41 80.225 3.898 ;
      RECT 80.175 3.41 80.22 3.835 ;
      RECT 80.15 3.41 80.175 3.753 ;
      RECT 80.135 3.41 80.15 3.705 ;
      RECT 80.13 3.41 80.135 3.675 ;
      RECT 82.52 3.455 82.78 3.715 ;
      RECT 82.515 3.455 82.78 3.663 ;
      RECT 82.51 3.455 82.78 3.633 ;
      RECT 82.485 3.325 82.765 3.605 ;
      RECT 70.99 9.095 71.34 9.445 ;
      RECT 81.955 9.05 82.305 9.4 ;
      RECT 70.99 9.125 82.305 9.325 ;
      RECT 81.525 5.005 81.805 5.285 ;
      RECT 81.565 4.96 81.83 5.22 ;
      RECT 81.555 4.995 81.83 5.22 ;
      RECT 81.56 4.98 81.805 5.285 ;
      RECT 81.565 4.957 81.775 5.285 ;
      RECT 81.565 4.955 81.76 5.285 ;
      RECT 81.605 4.945 81.76 5.285 ;
      RECT 81.575 4.95 81.76 5.285 ;
      RECT 81.605 4.942 81.705 5.285 ;
      RECT 81.63 4.935 81.705 5.285 ;
      RECT 81.61 4.937 81.705 5.285 ;
      RECT 80.94 4.45 81.2 4.71 ;
      RECT 80.99 4.442 81.18 4.71 ;
      RECT 80.995 4.362 81.18 4.71 ;
      RECT 81.115 3.75 81.18 4.71 ;
      RECT 81.02 4.147 81.18 4.71 ;
      RECT 81.095 3.835 81.18 4.71 ;
      RECT 81.13 3.46 81.266 4.188 ;
      RECT 81.075 3.957 81.266 4.188 ;
      RECT 81.09 3.897 81.18 4.71 ;
      RECT 81.13 3.46 81.29 3.853 ;
      RECT 81.13 3.46 81.3 3.75 ;
      RECT 81.12 3.46 81.38 3.72 ;
      RECT 79.455 4.86 79.5 5.12 ;
      RECT 79.36 3.395 79.505 3.655 ;
      RECT 79.865 4.017 79.875 4.108 ;
      RECT 79.85 3.955 79.865 4.164 ;
      RECT 79.845 3.902 79.85 4.21 ;
      RECT 79.795 3.849 79.845 4.336 ;
      RECT 79.79 3.804 79.795 4.483 ;
      RECT 79.78 3.792 79.79 4.525 ;
      RECT 79.745 3.756 79.78 4.63 ;
      RECT 79.74 3.724 79.745 4.736 ;
      RECT 79.725 3.706 79.74 4.781 ;
      RECT 79.72 3.689 79.725 4.015 ;
      RECT 79.715 4.07 79.725 4.838 ;
      RECT 79.71 3.675 79.72 3.988 ;
      RECT 79.705 4.125 79.715 5.12 ;
      RECT 79.7 3.661 79.71 3.973 ;
      RECT 79.7 4.175 79.705 5.12 ;
      RECT 79.685 3.638 79.7 3.953 ;
      RECT 79.665 4.297 79.7 5.12 ;
      RECT 79.68 3.62 79.685 3.935 ;
      RECT 79.675 3.612 79.68 3.925 ;
      RECT 79.645 3.58 79.675 3.889 ;
      RECT 79.655 4.425 79.665 5.12 ;
      RECT 79.65 4.452 79.655 5.12 ;
      RECT 79.645 4.502 79.65 5.12 ;
      RECT 79.635 3.546 79.645 3.854 ;
      RECT 79.595 4.57 79.645 5.12 ;
      RECT 79.62 3.523 79.635 3.83 ;
      RECT 79.595 3.395 79.62 3.793 ;
      RECT 79.59 3.395 79.595 3.765 ;
      RECT 79.56 4.67 79.595 5.12 ;
      RECT 79.585 3.395 79.59 3.758 ;
      RECT 79.58 3.395 79.585 3.748 ;
      RECT 79.565 3.395 79.58 3.733 ;
      RECT 79.55 3.395 79.565 3.705 ;
      RECT 79.515 4.775 79.56 5.12 ;
      RECT 79.535 3.395 79.55 3.678 ;
      RECT 79.505 3.395 79.535 3.663 ;
      RECT 79.5 4.847 79.515 5.12 ;
      RECT 79.425 3.93 79.465 4.19 ;
      RECT 79.2 3.877 79.205 4.135 ;
      RECT 75.155 3.355 75.415 3.615 ;
      RECT 75.155 3.38 75.43 3.595 ;
      RECT 77.545 3.205 77.55 3.35 ;
      RECT 79.415 3.925 79.425 4.19 ;
      RECT 79.395 3.917 79.415 4.19 ;
      RECT 79.377 3.913 79.395 4.19 ;
      RECT 79.291 3.902 79.377 4.19 ;
      RECT 79.205 3.885 79.291 4.19 ;
      RECT 79.15 3.872 79.2 4.12 ;
      RECT 79.116 3.864 79.15 4.095 ;
      RECT 79.03 3.853 79.116 4.06 ;
      RECT 78.995 3.83 79.03 4.025 ;
      RECT 78.985 3.792 78.995 4.011 ;
      RECT 78.98 3.765 78.985 4.007 ;
      RECT 78.975 3.752 78.98 4.004 ;
      RECT 78.965 3.732 78.975 4 ;
      RECT 78.96 3.707 78.965 3.996 ;
      RECT 78.935 3.662 78.96 3.99 ;
      RECT 78.925 3.603 78.935 3.982 ;
      RECT 78.915 3.571 78.925 3.973 ;
      RECT 78.895 3.523 78.915 3.953 ;
      RECT 78.89 3.483 78.895 3.923 ;
      RECT 78.875 3.457 78.89 3.897 ;
      RECT 78.87 3.435 78.875 3.873 ;
      RECT 78.855 3.407 78.87 3.849 ;
      RECT 78.84 3.38 78.855 3.813 ;
      RECT 78.825 3.357 78.84 3.775 ;
      RECT 78.82 3.347 78.825 3.75 ;
      RECT 78.81 3.34 78.82 3.733 ;
      RECT 78.795 3.327 78.81 3.703 ;
      RECT 78.79 3.317 78.795 3.678 ;
      RECT 78.785 3.312 78.79 3.665 ;
      RECT 78.775 3.305 78.785 3.645 ;
      RECT 78.77 3.298 78.775 3.63 ;
      RECT 78.745 3.291 78.77 3.588 ;
      RECT 78.73 3.281 78.745 3.538 ;
      RECT 78.72 3.276 78.73 3.508 ;
      RECT 78.71 3.272 78.72 3.483 ;
      RECT 78.695 3.269 78.71 3.473 ;
      RECT 78.645 3.266 78.695 3.458 ;
      RECT 78.625 3.264 78.645 3.443 ;
      RECT 78.576 3.262 78.625 3.438 ;
      RECT 78.49 3.258 78.576 3.433 ;
      RECT 78.451 3.255 78.49 3.429 ;
      RECT 78.365 3.251 78.451 3.424 ;
      RECT 78.315 3.248 78.365 3.418 ;
      RECT 78.266 3.245 78.315 3.413 ;
      RECT 78.18 3.242 78.266 3.408 ;
      RECT 78.176 3.24 78.18 3.405 ;
      RECT 78.09 3.237 78.176 3.4 ;
      RECT 78.041 3.233 78.09 3.393 ;
      RECT 77.955 3.23 78.041 3.388 ;
      RECT 77.931 3.227 77.955 3.384 ;
      RECT 77.845 3.225 77.931 3.379 ;
      RECT 77.78 3.221 77.845 3.372 ;
      RECT 77.777 3.22 77.78 3.369 ;
      RECT 77.691 3.217 77.777 3.366 ;
      RECT 77.605 3.211 77.691 3.359 ;
      RECT 77.575 3.207 77.605 3.355 ;
      RECT 77.55 3.205 77.575 3.353 ;
      RECT 77.495 3.202 77.545 3.35 ;
      RECT 77.415 3.201 77.495 3.35 ;
      RECT 77.36 3.203 77.415 3.353 ;
      RECT 77.345 3.204 77.36 3.357 ;
      RECT 77.29 3.212 77.345 3.367 ;
      RECT 77.26 3.22 77.29 3.38 ;
      RECT 77.241 3.221 77.26 3.386 ;
      RECT 77.155 3.224 77.241 3.391 ;
      RECT 77.085 3.229 77.155 3.4 ;
      RECT 77.066 3.232 77.085 3.406 ;
      RECT 76.98 3.236 77.066 3.411 ;
      RECT 76.94 3.24 76.98 3.418 ;
      RECT 76.931 3.242 76.94 3.421 ;
      RECT 76.845 3.246 76.931 3.426 ;
      RECT 76.842 3.249 76.845 3.43 ;
      RECT 76.756 3.252 76.842 3.434 ;
      RECT 76.67 3.258 76.756 3.442 ;
      RECT 76.646 3.262 76.67 3.446 ;
      RECT 76.56 3.266 76.646 3.451 ;
      RECT 76.515 3.271 76.56 3.458 ;
      RECT 76.435 3.276 76.515 3.465 ;
      RECT 76.355 3.282 76.435 3.48 ;
      RECT 76.33 3.286 76.355 3.493 ;
      RECT 76.265 3.289 76.33 3.505 ;
      RECT 76.21 3.294 76.265 3.52 ;
      RECT 76.18 3.297 76.21 3.538 ;
      RECT 76.17 3.299 76.18 3.551 ;
      RECT 76.11 3.314 76.17 3.561 ;
      RECT 76.095 3.331 76.11 3.57 ;
      RECT 76.09 3.34 76.095 3.57 ;
      RECT 76.08 3.35 76.09 3.57 ;
      RECT 76.07 3.367 76.08 3.57 ;
      RECT 76.05 3.377 76.07 3.571 ;
      RECT 76.005 3.387 76.05 3.572 ;
      RECT 75.97 3.396 76.005 3.574 ;
      RECT 75.905 3.401 75.97 3.576 ;
      RECT 75.825 3.402 75.905 3.579 ;
      RECT 75.821 3.4 75.825 3.58 ;
      RECT 75.735 3.397 75.821 3.582 ;
      RECT 75.688 3.394 75.735 3.584 ;
      RECT 75.602 3.39 75.688 3.587 ;
      RECT 75.516 3.386 75.602 3.59 ;
      RECT 75.43 3.382 75.516 3.594 ;
      RECT 78.815 5.005 78.845 5.285 ;
      RECT 78.565 4.895 78.585 5.285 ;
      RECT 78.52 4.895 78.585 5.155 ;
      RECT 78.35 3.52 78.385 3.78 ;
      RECT 78.125 3.52 78.185 3.78 ;
      RECT 78.805 4.985 78.815 5.285 ;
      RECT 78.8 4.945 78.805 5.285 ;
      RECT 78.785 4.9 78.8 5.285 ;
      RECT 78.78 4.865 78.785 5.285 ;
      RECT 78.775 4.845 78.78 5.285 ;
      RECT 78.745 4.772 78.775 5.285 ;
      RECT 78.725 4.67 78.745 5.285 ;
      RECT 78.715 4.6 78.725 5.285 ;
      RECT 78.67 4.54 78.715 5.285 ;
      RECT 78.585 4.501 78.67 5.285 ;
      RECT 78.58 4.492 78.585 4.865 ;
      RECT 78.57 4.491 78.58 4.848 ;
      RECT 78.545 4.472 78.57 4.818 ;
      RECT 78.54 4.447 78.545 4.797 ;
      RECT 78.53 4.425 78.54 4.788 ;
      RECT 78.525 4.396 78.53 4.778 ;
      RECT 78.485 4.322 78.525 4.75 ;
      RECT 78.465 4.223 78.485 4.715 ;
      RECT 78.45 4.159 78.465 4.698 ;
      RECT 78.42 4.083 78.45 4.67 ;
      RECT 78.4 3.998 78.42 4.643 ;
      RECT 78.36 3.894 78.4 4.55 ;
      RECT 78.355 3.815 78.36 4.458 ;
      RECT 78.35 3.798 78.355 4.435 ;
      RECT 78.345 3.52 78.35 4.415 ;
      RECT 78.315 3.52 78.345 4.353 ;
      RECT 78.31 3.52 78.315 4.285 ;
      RECT 78.3 3.52 78.31 4.25 ;
      RECT 78.29 3.52 78.3 4.215 ;
      RECT 78.225 3.52 78.29 4.07 ;
      RECT 78.22 3.52 78.225 3.94 ;
      RECT 78.19 3.52 78.22 3.873 ;
      RECT 78.185 3.52 78.19 3.798 ;
      RECT 77.365 4.445 77.645 4.725 ;
      RECT 77.405 4.425 77.665 4.685 ;
      RECT 77.395 4.435 77.665 4.685 ;
      RECT 77.405 4.362 77.62 4.725 ;
      RECT 77.46 4.285 77.615 4.725 ;
      RECT 77.465 4.07 77.615 4.725 ;
      RECT 77.455 3.872 77.605 4.123 ;
      RECT 77.445 3.872 77.605 3.99 ;
      RECT 77.44 3.75 77.6 3.893 ;
      RECT 77.425 3.75 77.6 3.798 ;
      RECT 77.42 3.46 77.595 3.775 ;
      RECT 77.405 3.46 77.595 3.745 ;
      RECT 77.365 3.46 77.625 3.72 ;
      RECT 77.275 4.93 77.355 5.19 ;
      RECT 76.68 3.65 76.685 3.915 ;
      RECT 76.56 3.65 76.685 3.91 ;
      RECT 77.235 4.895 77.275 5.19 ;
      RECT 77.19 4.817 77.235 5.19 ;
      RECT 77.17 4.745 77.19 5.19 ;
      RECT 77.16 4.697 77.17 5.19 ;
      RECT 77.125 4.63 77.16 5.19 ;
      RECT 77.095 4.53 77.125 5.19 ;
      RECT 77.075 4.455 77.095 4.99 ;
      RECT 77.065 4.405 77.075 4.945 ;
      RECT 77.06 4.382 77.065 4.918 ;
      RECT 77.055 4.367 77.06 4.905 ;
      RECT 77.05 4.352 77.055 4.883 ;
      RECT 77.045 4.337 77.05 4.865 ;
      RECT 77.02 4.292 77.045 4.82 ;
      RECT 77.01 4.24 77.02 4.763 ;
      RECT 77 4.21 77.01 4.73 ;
      RECT 76.99 4.175 77 4.698 ;
      RECT 76.955 4.107 76.99 4.63 ;
      RECT 76.95 4.046 76.955 4.565 ;
      RECT 76.94 4.034 76.95 4.545 ;
      RECT 76.935 4.022 76.94 4.525 ;
      RECT 76.93 4.014 76.935 4.513 ;
      RECT 76.925 4.006 76.93 4.493 ;
      RECT 76.915 3.994 76.925 4.465 ;
      RECT 76.905 3.978 76.915 4.435 ;
      RECT 76.88 3.95 76.905 4.373 ;
      RECT 76.87 3.921 76.88 4.318 ;
      RECT 76.855 3.9 76.87 4.278 ;
      RECT 76.85 3.884 76.855 4.25 ;
      RECT 76.845 3.872 76.85 4.24 ;
      RECT 76.84 3.867 76.845 4.213 ;
      RECT 76.835 3.86 76.84 4.2 ;
      RECT 76.82 3.843 76.835 4.173 ;
      RECT 76.81 3.65 76.82 4.133 ;
      RECT 76.8 3.65 76.81 4.1 ;
      RECT 76.79 3.65 76.8 4.075 ;
      RECT 76.72 3.65 76.79 4.01 ;
      RECT 76.71 3.65 76.72 3.958 ;
      RECT 76.695 3.65 76.71 3.94 ;
      RECT 76.685 3.65 76.695 3.925 ;
      RECT 76.515 4.52 76.775 4.78 ;
      RECT 75.05 4.555 75.055 4.762 ;
      RECT 74.685 4.445 74.76 4.76 ;
      RECT 74.5 4.5 74.655 4.76 ;
      RECT 74.685 4.445 74.79 4.725 ;
      RECT 76.5 4.617 76.515 4.778 ;
      RECT 76.475 4.625 76.5 4.783 ;
      RECT 76.45 4.632 76.475 4.788 ;
      RECT 76.387 4.643 76.45 4.797 ;
      RECT 76.301 4.662 76.387 4.814 ;
      RECT 76.215 4.684 76.301 4.833 ;
      RECT 76.2 4.697 76.215 4.844 ;
      RECT 76.16 4.705 76.2 4.851 ;
      RECT 76.14 4.71 76.16 4.858 ;
      RECT 76.102 4.711 76.14 4.861 ;
      RECT 76.016 4.714 76.102 4.862 ;
      RECT 75.93 4.718 76.016 4.863 ;
      RECT 75.881 4.72 75.93 4.865 ;
      RECT 75.795 4.72 75.881 4.867 ;
      RECT 75.755 4.715 75.795 4.869 ;
      RECT 75.745 4.709 75.755 4.87 ;
      RECT 75.705 4.704 75.745 4.867 ;
      RECT 75.695 4.697 75.705 4.863 ;
      RECT 75.68 4.693 75.695 4.861 ;
      RECT 75.663 4.689 75.68 4.859 ;
      RECT 75.577 4.679 75.663 4.851 ;
      RECT 75.491 4.661 75.577 4.837 ;
      RECT 75.405 4.644 75.491 4.823 ;
      RECT 75.38 4.632 75.405 4.814 ;
      RECT 75.31 4.622 75.38 4.807 ;
      RECT 75.265 4.61 75.31 4.798 ;
      RECT 75.205 4.597 75.265 4.79 ;
      RECT 75.2 4.589 75.205 4.785 ;
      RECT 75.165 4.584 75.2 4.783 ;
      RECT 75.11 4.575 75.165 4.776 ;
      RECT 75.07 4.564 75.11 4.768 ;
      RECT 75.055 4.557 75.07 4.764 ;
      RECT 75.035 4.55 75.05 4.761 ;
      RECT 75.02 4.54 75.035 4.759 ;
      RECT 75.005 4.527 75.02 4.756 ;
      RECT 74.98 4.51 75.005 4.752 ;
      RECT 74.965 4.492 74.98 4.749 ;
      RECT 74.94 4.445 74.965 4.747 ;
      RECT 74.916 4.445 74.94 4.744 ;
      RECT 74.83 4.445 74.916 4.736 ;
      RECT 74.79 4.445 74.83 4.728 ;
      RECT 74.655 4.492 74.685 4.76 ;
      RECT 76.335 4.075 76.595 4.335 ;
      RECT 76.295 4.075 76.595 4.213 ;
      RECT 76.26 4.075 76.595 4.198 ;
      RECT 76.205 4.075 76.595 4.178 ;
      RECT 76.125 3.885 76.405 4.165 ;
      RECT 76.125 4.067 76.475 4.165 ;
      RECT 76.125 4.01 76.46 4.165 ;
      RECT 76.125 3.957 76.41 4.165 ;
      RECT 73.285 4.244 73.3 4.7 ;
      RECT 73.28 4.316 73.386 4.698 ;
      RECT 73.3 3.41 73.435 4.696 ;
      RECT 73.285 4.26 73.44 4.695 ;
      RECT 73.285 4.31 73.445 4.693 ;
      RECT 73.27 4.375 73.445 4.692 ;
      RECT 73.28 4.367 73.45 4.689 ;
      RECT 73.26 4.415 73.45 4.684 ;
      RECT 73.26 4.415 73.465 4.681 ;
      RECT 73.255 4.415 73.465 4.678 ;
      RECT 73.23 4.415 73.49 4.675 ;
      RECT 73.3 3.41 73.46 4.063 ;
      RECT 73.295 3.41 73.46 4.035 ;
      RECT 73.29 3.41 73.46 3.863 ;
      RECT 73.29 3.41 73.48 3.803 ;
      RECT 73.245 3.41 73.505 3.67 ;
      RECT 72.725 3.885 73.005 4.165 ;
      RECT 72.715 3.9 73.005 4.16 ;
      RECT 72.67 3.962 73.005 4.158 ;
      RECT 72.745 3.877 72.91 4.165 ;
      RECT 72.745 3.862 72.866 4.165 ;
      RECT 72.78 3.855 72.866 4.165 ;
      RECT 72.245 5.005 72.525 5.285 ;
      RECT 72.205 4.967 72.5 5.078 ;
      RECT 72.19 4.917 72.48 4.973 ;
      RECT 72.135 4.68 72.395 4.94 ;
      RECT 72.135 4.882 72.475 4.94 ;
      RECT 72.135 4.822 72.47 4.94 ;
      RECT 72.135 4.772 72.45 4.94 ;
      RECT 72.135 4.752 72.445 4.94 ;
      RECT 72.135 4.73 72.44 4.94 ;
      RECT 72.135 4.715 72.41 4.94 ;
      RECT 67.855 8.66 68.175 8.98 ;
      RECT 67.885 8.13 68.055 8.98 ;
      RECT 67.885 8.13 68.06 8.48 ;
      RECT 67.885 8.13 68.86 8.305 ;
      RECT 68.685 3.26 68.86 8.305 ;
      RECT 68.63 3.26 68.98 3.61 ;
      RECT 68.655 9.09 68.98 9.415 ;
      RECT 67.54 9.18 68.98 9.35 ;
      RECT 67.54 3.69 67.7 9.35 ;
      RECT 67.855 3.66 68.175 3.98 ;
      RECT 67.54 3.69 68.175 3.86 ;
      RECT 66.22 2.435 66.595 2.805 ;
      RECT 58.13 2.255 58.505 2.625 ;
      RECT 56.695 2.255 57.07 2.625 ;
      RECT 56.695 2.375 66.525 2.545 ;
      RECT 62.64 5.655 66.495 5.825 ;
      RECT 66.325 4.72 66.495 5.825 ;
      RECT 62.64 4.965 62.81 5.825 ;
      RECT 62.6 5.005 62.88 5.285 ;
      RECT 62.62 4.965 62.88 5.285 ;
      RECT 62.26 4.92 62.365 5.18 ;
      RECT 66.235 4.725 66.585 5.075 ;
      RECT 62.115 3.41 62.205 3.67 ;
      RECT 62.655 4.475 62.66 4.515 ;
      RECT 62.65 4.465 62.655 4.6 ;
      RECT 62.645 4.455 62.65 4.693 ;
      RECT 62.635 4.435 62.645 4.749 ;
      RECT 62.555 4.363 62.635 4.829 ;
      RECT 62.59 5.007 62.6 5.232 ;
      RECT 62.585 5.004 62.59 5.227 ;
      RECT 62.57 5.001 62.585 5.22 ;
      RECT 62.535 4.995 62.57 5.202 ;
      RECT 62.55 4.298 62.555 4.903 ;
      RECT 62.53 4.249 62.55 4.918 ;
      RECT 62.52 4.982 62.535 5.185 ;
      RECT 62.525 4.191 62.53 4.933 ;
      RECT 62.52 4.169 62.525 4.943 ;
      RECT 62.485 4.079 62.52 5.18 ;
      RECT 62.47 3.957 62.485 5.18 ;
      RECT 62.465 3.91 62.47 5.18 ;
      RECT 62.44 3.835 62.465 5.18 ;
      RECT 62.425 3.75 62.44 5.18 ;
      RECT 62.42 3.697 62.425 5.18 ;
      RECT 62.415 3.677 62.42 5.18 ;
      RECT 62.41 3.652 62.415 4.414 ;
      RECT 62.395 4.612 62.415 5.18 ;
      RECT 62.405 3.63 62.41 4.391 ;
      RECT 62.395 3.582 62.405 4.356 ;
      RECT 62.39 3.545 62.395 4.322 ;
      RECT 62.39 4.692 62.395 5.18 ;
      RECT 62.375 3.522 62.39 4.277 ;
      RECT 62.37 4.79 62.39 5.18 ;
      RECT 62.32 3.41 62.375 4.119 ;
      RECT 62.365 4.912 62.37 5.18 ;
      RECT 62.305 3.41 62.32 3.958 ;
      RECT 62.3 3.41 62.305 3.91 ;
      RECT 62.295 3.41 62.3 3.898 ;
      RECT 62.25 3.41 62.295 3.835 ;
      RECT 62.225 3.41 62.25 3.753 ;
      RECT 62.21 3.41 62.225 3.705 ;
      RECT 62.205 3.41 62.21 3.675 ;
      RECT 64.595 3.455 64.855 3.715 ;
      RECT 64.59 3.455 64.855 3.663 ;
      RECT 64.585 3.455 64.855 3.633 ;
      RECT 64.56 3.325 64.84 3.605 ;
      RECT 53.11 9.095 53.46 9.445 ;
      RECT 64.085 9.05 64.435 9.4 ;
      RECT 53.11 9.125 64.435 9.325 ;
      RECT 63.6 5.005 63.88 5.285 ;
      RECT 63.64 4.96 63.905 5.22 ;
      RECT 63.63 4.995 63.905 5.22 ;
      RECT 63.635 4.98 63.88 5.285 ;
      RECT 63.64 4.957 63.85 5.285 ;
      RECT 63.64 4.955 63.835 5.285 ;
      RECT 63.68 4.945 63.835 5.285 ;
      RECT 63.65 4.95 63.835 5.285 ;
      RECT 63.68 4.942 63.78 5.285 ;
      RECT 63.705 4.935 63.78 5.285 ;
      RECT 63.685 4.937 63.78 5.285 ;
      RECT 63.015 4.45 63.275 4.71 ;
      RECT 63.065 4.442 63.255 4.71 ;
      RECT 63.07 4.362 63.255 4.71 ;
      RECT 63.19 3.75 63.255 4.71 ;
      RECT 63.095 4.147 63.255 4.71 ;
      RECT 63.17 3.835 63.255 4.71 ;
      RECT 63.205 3.46 63.341 4.188 ;
      RECT 63.15 3.957 63.341 4.188 ;
      RECT 63.165 3.897 63.255 4.71 ;
      RECT 63.205 3.46 63.365 3.853 ;
      RECT 63.205 3.46 63.375 3.75 ;
      RECT 63.195 3.46 63.455 3.72 ;
      RECT 61.53 4.86 61.575 5.12 ;
      RECT 61.435 3.395 61.58 3.655 ;
      RECT 61.94 4.017 61.95 4.108 ;
      RECT 61.925 3.955 61.94 4.164 ;
      RECT 61.92 3.902 61.925 4.21 ;
      RECT 61.87 3.849 61.92 4.336 ;
      RECT 61.865 3.804 61.87 4.483 ;
      RECT 61.855 3.792 61.865 4.525 ;
      RECT 61.82 3.756 61.855 4.63 ;
      RECT 61.815 3.724 61.82 4.736 ;
      RECT 61.8 3.706 61.815 4.781 ;
      RECT 61.795 3.689 61.8 4.015 ;
      RECT 61.79 4.07 61.8 4.838 ;
      RECT 61.785 3.675 61.795 3.988 ;
      RECT 61.78 4.125 61.79 5.12 ;
      RECT 61.775 3.661 61.785 3.973 ;
      RECT 61.775 4.175 61.78 5.12 ;
      RECT 61.76 3.638 61.775 3.953 ;
      RECT 61.74 4.297 61.775 5.12 ;
      RECT 61.755 3.62 61.76 3.935 ;
      RECT 61.75 3.612 61.755 3.925 ;
      RECT 61.72 3.58 61.75 3.889 ;
      RECT 61.73 4.425 61.74 5.12 ;
      RECT 61.725 4.452 61.73 5.12 ;
      RECT 61.72 4.502 61.725 5.12 ;
      RECT 61.71 3.546 61.72 3.854 ;
      RECT 61.67 4.57 61.72 5.12 ;
      RECT 61.695 3.523 61.71 3.83 ;
      RECT 61.67 3.395 61.695 3.793 ;
      RECT 61.665 3.395 61.67 3.765 ;
      RECT 61.635 4.67 61.67 5.12 ;
      RECT 61.66 3.395 61.665 3.758 ;
      RECT 61.655 3.395 61.66 3.748 ;
      RECT 61.64 3.395 61.655 3.733 ;
      RECT 61.625 3.395 61.64 3.705 ;
      RECT 61.59 4.775 61.635 5.12 ;
      RECT 61.61 3.395 61.625 3.678 ;
      RECT 61.58 3.395 61.61 3.663 ;
      RECT 61.575 4.847 61.59 5.12 ;
      RECT 61.5 3.93 61.54 4.19 ;
      RECT 61.275 3.877 61.28 4.135 ;
      RECT 57.23 3.355 57.49 3.615 ;
      RECT 57.23 3.38 57.505 3.595 ;
      RECT 59.62 3.205 59.625 3.35 ;
      RECT 61.49 3.925 61.5 4.19 ;
      RECT 61.47 3.917 61.49 4.19 ;
      RECT 61.452 3.913 61.47 4.19 ;
      RECT 61.366 3.902 61.452 4.19 ;
      RECT 61.28 3.885 61.366 4.19 ;
      RECT 61.225 3.872 61.275 4.12 ;
      RECT 61.191 3.864 61.225 4.095 ;
      RECT 61.105 3.853 61.191 4.06 ;
      RECT 61.07 3.83 61.105 4.025 ;
      RECT 61.06 3.792 61.07 4.011 ;
      RECT 61.055 3.765 61.06 4.007 ;
      RECT 61.05 3.752 61.055 4.004 ;
      RECT 61.04 3.732 61.05 4 ;
      RECT 61.035 3.707 61.04 3.996 ;
      RECT 61.01 3.662 61.035 3.99 ;
      RECT 61 3.603 61.01 3.982 ;
      RECT 60.99 3.571 61 3.973 ;
      RECT 60.97 3.523 60.99 3.953 ;
      RECT 60.965 3.483 60.97 3.923 ;
      RECT 60.95 3.457 60.965 3.897 ;
      RECT 60.945 3.435 60.95 3.873 ;
      RECT 60.93 3.407 60.945 3.849 ;
      RECT 60.915 3.38 60.93 3.813 ;
      RECT 60.9 3.357 60.915 3.775 ;
      RECT 60.895 3.347 60.9 3.75 ;
      RECT 60.885 3.34 60.895 3.733 ;
      RECT 60.87 3.327 60.885 3.703 ;
      RECT 60.865 3.317 60.87 3.678 ;
      RECT 60.86 3.312 60.865 3.665 ;
      RECT 60.85 3.305 60.86 3.645 ;
      RECT 60.845 3.298 60.85 3.63 ;
      RECT 60.82 3.291 60.845 3.588 ;
      RECT 60.805 3.281 60.82 3.538 ;
      RECT 60.795 3.276 60.805 3.508 ;
      RECT 60.785 3.272 60.795 3.483 ;
      RECT 60.77 3.269 60.785 3.473 ;
      RECT 60.72 3.266 60.77 3.458 ;
      RECT 60.7 3.264 60.72 3.443 ;
      RECT 60.651 3.262 60.7 3.438 ;
      RECT 60.565 3.258 60.651 3.433 ;
      RECT 60.526 3.255 60.565 3.429 ;
      RECT 60.44 3.251 60.526 3.424 ;
      RECT 60.39 3.248 60.44 3.418 ;
      RECT 60.341 3.245 60.39 3.413 ;
      RECT 60.255 3.242 60.341 3.408 ;
      RECT 60.251 3.24 60.255 3.405 ;
      RECT 60.165 3.237 60.251 3.4 ;
      RECT 60.116 3.233 60.165 3.393 ;
      RECT 60.03 3.23 60.116 3.388 ;
      RECT 60.006 3.227 60.03 3.384 ;
      RECT 59.92 3.225 60.006 3.379 ;
      RECT 59.855 3.221 59.92 3.372 ;
      RECT 59.852 3.22 59.855 3.369 ;
      RECT 59.766 3.217 59.852 3.366 ;
      RECT 59.68 3.211 59.766 3.359 ;
      RECT 59.65 3.207 59.68 3.355 ;
      RECT 59.625 3.205 59.65 3.353 ;
      RECT 59.57 3.202 59.62 3.35 ;
      RECT 59.49 3.201 59.57 3.35 ;
      RECT 59.435 3.203 59.49 3.353 ;
      RECT 59.42 3.204 59.435 3.357 ;
      RECT 59.365 3.212 59.42 3.367 ;
      RECT 59.335 3.22 59.365 3.38 ;
      RECT 59.316 3.221 59.335 3.386 ;
      RECT 59.23 3.224 59.316 3.391 ;
      RECT 59.16 3.229 59.23 3.4 ;
      RECT 59.141 3.232 59.16 3.406 ;
      RECT 59.055 3.236 59.141 3.411 ;
      RECT 59.015 3.24 59.055 3.418 ;
      RECT 59.006 3.242 59.015 3.421 ;
      RECT 58.92 3.246 59.006 3.426 ;
      RECT 58.917 3.249 58.92 3.43 ;
      RECT 58.831 3.252 58.917 3.434 ;
      RECT 58.745 3.258 58.831 3.442 ;
      RECT 58.721 3.262 58.745 3.446 ;
      RECT 58.635 3.266 58.721 3.451 ;
      RECT 58.59 3.271 58.635 3.458 ;
      RECT 58.51 3.276 58.59 3.465 ;
      RECT 58.43 3.282 58.51 3.48 ;
      RECT 58.405 3.286 58.43 3.493 ;
      RECT 58.34 3.289 58.405 3.505 ;
      RECT 58.285 3.294 58.34 3.52 ;
      RECT 58.255 3.297 58.285 3.538 ;
      RECT 58.245 3.299 58.255 3.551 ;
      RECT 58.185 3.314 58.245 3.561 ;
      RECT 58.17 3.331 58.185 3.57 ;
      RECT 58.165 3.34 58.17 3.57 ;
      RECT 58.155 3.35 58.165 3.57 ;
      RECT 58.145 3.367 58.155 3.57 ;
      RECT 58.125 3.377 58.145 3.571 ;
      RECT 58.08 3.387 58.125 3.572 ;
      RECT 58.045 3.396 58.08 3.574 ;
      RECT 57.98 3.401 58.045 3.576 ;
      RECT 57.9 3.402 57.98 3.579 ;
      RECT 57.896 3.4 57.9 3.58 ;
      RECT 57.81 3.397 57.896 3.582 ;
      RECT 57.763 3.394 57.81 3.584 ;
      RECT 57.677 3.39 57.763 3.587 ;
      RECT 57.591 3.386 57.677 3.59 ;
      RECT 57.505 3.382 57.591 3.594 ;
      RECT 60.89 5.005 60.92 5.285 ;
      RECT 60.64 4.895 60.66 5.285 ;
      RECT 60.595 4.895 60.66 5.155 ;
      RECT 60.425 3.52 60.46 3.78 ;
      RECT 60.2 3.52 60.26 3.78 ;
      RECT 60.88 4.985 60.89 5.285 ;
      RECT 60.875 4.945 60.88 5.285 ;
      RECT 60.86 4.9 60.875 5.285 ;
      RECT 60.855 4.865 60.86 5.285 ;
      RECT 60.85 4.845 60.855 5.285 ;
      RECT 60.82 4.772 60.85 5.285 ;
      RECT 60.8 4.67 60.82 5.285 ;
      RECT 60.79 4.6 60.8 5.285 ;
      RECT 60.745 4.54 60.79 5.285 ;
      RECT 60.66 4.501 60.745 5.285 ;
      RECT 60.655 4.492 60.66 4.865 ;
      RECT 60.645 4.491 60.655 4.848 ;
      RECT 60.62 4.472 60.645 4.818 ;
      RECT 60.615 4.447 60.62 4.797 ;
      RECT 60.605 4.425 60.615 4.788 ;
      RECT 60.6 4.396 60.605 4.778 ;
      RECT 60.56 4.322 60.6 4.75 ;
      RECT 60.54 4.223 60.56 4.715 ;
      RECT 60.525 4.159 60.54 4.698 ;
      RECT 60.495 4.083 60.525 4.67 ;
      RECT 60.475 3.998 60.495 4.643 ;
      RECT 60.435 3.894 60.475 4.55 ;
      RECT 60.43 3.815 60.435 4.458 ;
      RECT 60.425 3.798 60.43 4.435 ;
      RECT 60.42 3.52 60.425 4.415 ;
      RECT 60.39 3.52 60.42 4.353 ;
      RECT 60.385 3.52 60.39 4.285 ;
      RECT 60.375 3.52 60.385 4.25 ;
      RECT 60.365 3.52 60.375 4.215 ;
      RECT 60.3 3.52 60.365 4.07 ;
      RECT 60.295 3.52 60.3 3.94 ;
      RECT 60.265 3.52 60.295 3.873 ;
      RECT 60.26 3.52 60.265 3.798 ;
      RECT 59.44 4.445 59.72 4.725 ;
      RECT 59.48 4.425 59.74 4.685 ;
      RECT 59.47 4.435 59.74 4.685 ;
      RECT 59.48 4.362 59.695 4.725 ;
      RECT 59.535 4.285 59.69 4.725 ;
      RECT 59.54 4.07 59.69 4.725 ;
      RECT 59.53 3.872 59.68 4.123 ;
      RECT 59.52 3.872 59.68 3.99 ;
      RECT 59.515 3.75 59.675 3.893 ;
      RECT 59.5 3.75 59.675 3.798 ;
      RECT 59.495 3.46 59.67 3.775 ;
      RECT 59.48 3.46 59.67 3.745 ;
      RECT 59.44 3.46 59.7 3.72 ;
      RECT 59.35 4.93 59.43 5.19 ;
      RECT 58.755 3.65 58.76 3.915 ;
      RECT 58.635 3.65 58.76 3.91 ;
      RECT 59.31 4.895 59.35 5.19 ;
      RECT 59.265 4.817 59.31 5.19 ;
      RECT 59.245 4.745 59.265 5.19 ;
      RECT 59.235 4.697 59.245 5.19 ;
      RECT 59.2 4.63 59.235 5.19 ;
      RECT 59.17 4.53 59.2 5.19 ;
      RECT 59.15 4.455 59.17 4.99 ;
      RECT 59.14 4.405 59.15 4.945 ;
      RECT 59.135 4.382 59.14 4.918 ;
      RECT 59.13 4.367 59.135 4.905 ;
      RECT 59.125 4.352 59.13 4.883 ;
      RECT 59.12 4.337 59.125 4.865 ;
      RECT 59.095 4.292 59.12 4.82 ;
      RECT 59.085 4.24 59.095 4.763 ;
      RECT 59.075 4.21 59.085 4.73 ;
      RECT 59.065 4.175 59.075 4.698 ;
      RECT 59.03 4.107 59.065 4.63 ;
      RECT 59.025 4.046 59.03 4.565 ;
      RECT 59.015 4.034 59.025 4.545 ;
      RECT 59.01 4.022 59.015 4.525 ;
      RECT 59.005 4.014 59.01 4.513 ;
      RECT 59 4.006 59.005 4.493 ;
      RECT 58.99 3.994 59 4.465 ;
      RECT 58.98 3.978 58.99 4.435 ;
      RECT 58.955 3.95 58.98 4.373 ;
      RECT 58.945 3.921 58.955 4.318 ;
      RECT 58.93 3.9 58.945 4.278 ;
      RECT 58.925 3.884 58.93 4.25 ;
      RECT 58.92 3.872 58.925 4.24 ;
      RECT 58.915 3.867 58.92 4.213 ;
      RECT 58.91 3.86 58.915 4.2 ;
      RECT 58.895 3.843 58.91 4.173 ;
      RECT 58.885 3.65 58.895 4.133 ;
      RECT 58.875 3.65 58.885 4.1 ;
      RECT 58.865 3.65 58.875 4.075 ;
      RECT 58.795 3.65 58.865 4.01 ;
      RECT 58.785 3.65 58.795 3.958 ;
      RECT 58.77 3.65 58.785 3.94 ;
      RECT 58.76 3.65 58.77 3.925 ;
      RECT 58.59 4.52 58.85 4.78 ;
      RECT 57.125 4.555 57.13 4.762 ;
      RECT 56.76 4.445 56.835 4.76 ;
      RECT 56.575 4.5 56.73 4.76 ;
      RECT 56.76 4.445 56.865 4.725 ;
      RECT 58.575 4.617 58.59 4.778 ;
      RECT 58.55 4.625 58.575 4.783 ;
      RECT 58.525 4.632 58.55 4.788 ;
      RECT 58.462 4.643 58.525 4.797 ;
      RECT 58.376 4.662 58.462 4.814 ;
      RECT 58.29 4.684 58.376 4.833 ;
      RECT 58.275 4.697 58.29 4.844 ;
      RECT 58.235 4.705 58.275 4.851 ;
      RECT 58.215 4.71 58.235 4.858 ;
      RECT 58.177 4.711 58.215 4.861 ;
      RECT 58.091 4.714 58.177 4.862 ;
      RECT 58.005 4.718 58.091 4.863 ;
      RECT 57.956 4.72 58.005 4.865 ;
      RECT 57.87 4.72 57.956 4.867 ;
      RECT 57.83 4.715 57.87 4.869 ;
      RECT 57.82 4.709 57.83 4.87 ;
      RECT 57.78 4.704 57.82 4.867 ;
      RECT 57.77 4.697 57.78 4.863 ;
      RECT 57.755 4.693 57.77 4.861 ;
      RECT 57.738 4.689 57.755 4.859 ;
      RECT 57.652 4.679 57.738 4.851 ;
      RECT 57.566 4.661 57.652 4.837 ;
      RECT 57.48 4.644 57.566 4.823 ;
      RECT 57.455 4.632 57.48 4.814 ;
      RECT 57.385 4.622 57.455 4.807 ;
      RECT 57.34 4.61 57.385 4.798 ;
      RECT 57.28 4.597 57.34 4.79 ;
      RECT 57.275 4.589 57.28 4.785 ;
      RECT 57.24 4.584 57.275 4.783 ;
      RECT 57.185 4.575 57.24 4.776 ;
      RECT 57.145 4.564 57.185 4.768 ;
      RECT 57.13 4.557 57.145 4.764 ;
      RECT 57.11 4.55 57.125 4.761 ;
      RECT 57.095 4.54 57.11 4.759 ;
      RECT 57.08 4.527 57.095 4.756 ;
      RECT 57.055 4.51 57.08 4.752 ;
      RECT 57.04 4.492 57.055 4.749 ;
      RECT 57.015 4.445 57.04 4.747 ;
      RECT 56.991 4.445 57.015 4.744 ;
      RECT 56.905 4.445 56.991 4.736 ;
      RECT 56.865 4.445 56.905 4.728 ;
      RECT 56.73 4.492 56.76 4.76 ;
      RECT 58.41 4.075 58.67 4.335 ;
      RECT 58.37 4.075 58.67 4.213 ;
      RECT 58.335 4.075 58.67 4.198 ;
      RECT 58.28 4.075 58.67 4.178 ;
      RECT 58.2 3.885 58.48 4.165 ;
      RECT 58.2 4.067 58.55 4.165 ;
      RECT 58.2 4.01 58.535 4.165 ;
      RECT 58.2 3.957 58.485 4.165 ;
      RECT 55.36 4.244 55.375 4.7 ;
      RECT 55.355 4.316 55.461 4.698 ;
      RECT 55.375 3.41 55.51 4.696 ;
      RECT 55.36 4.26 55.515 4.695 ;
      RECT 55.36 4.31 55.52 4.693 ;
      RECT 55.345 4.375 55.52 4.692 ;
      RECT 55.355 4.367 55.525 4.689 ;
      RECT 55.335 4.415 55.525 4.684 ;
      RECT 55.335 4.415 55.54 4.681 ;
      RECT 55.33 4.415 55.54 4.678 ;
      RECT 55.305 4.415 55.565 4.675 ;
      RECT 55.375 3.41 55.535 4.063 ;
      RECT 55.37 3.41 55.535 4.035 ;
      RECT 55.365 3.41 55.535 3.863 ;
      RECT 55.365 3.41 55.555 3.803 ;
      RECT 55.32 3.41 55.58 3.67 ;
      RECT 54.8 3.885 55.08 4.165 ;
      RECT 54.79 3.9 55.08 4.16 ;
      RECT 54.745 3.962 55.08 4.158 ;
      RECT 54.82 3.877 54.985 4.165 ;
      RECT 54.82 3.862 54.941 4.165 ;
      RECT 54.855 3.855 54.941 4.165 ;
      RECT 54.32 5.005 54.6 5.285 ;
      RECT 54.28 4.967 54.575 5.078 ;
      RECT 54.265 4.917 54.555 4.973 ;
      RECT 54.21 4.68 54.47 4.94 ;
      RECT 54.21 4.882 54.55 4.94 ;
      RECT 54.21 4.822 54.545 4.94 ;
      RECT 54.21 4.772 54.525 4.94 ;
      RECT 54.21 4.752 54.52 4.94 ;
      RECT 54.21 4.73 54.515 4.94 ;
      RECT 54.21 4.715 54.485 4.94 ;
      RECT 49.93 8.66 50.25 8.98 ;
      RECT 49.96 8.13 50.13 8.98 ;
      RECT 49.96 8.13 50.135 8.48 ;
      RECT 49.96 8.13 50.935 8.305 ;
      RECT 50.76 3.26 50.935 8.305 ;
      RECT 50.705 3.26 51.055 3.61 ;
      RECT 50.73 9.09 51.055 9.415 ;
      RECT 49.615 9.18 51.055 9.35 ;
      RECT 49.615 3.69 49.775 9.35 ;
      RECT 49.93 3.66 50.25 3.98 ;
      RECT 49.615 3.69 50.25 3.86 ;
      RECT 48.295 2.435 48.67 2.805 ;
      RECT 40.205 2.255 40.58 2.625 ;
      RECT 38.77 2.255 39.145 2.625 ;
      RECT 38.77 2.375 48.6 2.545 ;
      RECT 44.715 5.655 48.57 5.825 ;
      RECT 48.4 4.72 48.57 5.825 ;
      RECT 44.715 4.965 44.885 5.825 ;
      RECT 44.675 5.005 44.955 5.285 ;
      RECT 44.695 4.965 44.955 5.285 ;
      RECT 44.335 4.92 44.44 5.18 ;
      RECT 48.31 4.725 48.66 5.075 ;
      RECT 44.19 3.41 44.28 3.67 ;
      RECT 44.73 4.475 44.735 4.515 ;
      RECT 44.725 4.465 44.73 4.6 ;
      RECT 44.72 4.455 44.725 4.693 ;
      RECT 44.71 4.435 44.72 4.749 ;
      RECT 44.63 4.363 44.71 4.829 ;
      RECT 44.665 5.007 44.675 5.232 ;
      RECT 44.66 5.004 44.665 5.227 ;
      RECT 44.645 5.001 44.66 5.22 ;
      RECT 44.61 4.995 44.645 5.202 ;
      RECT 44.625 4.298 44.63 4.903 ;
      RECT 44.605 4.249 44.625 4.918 ;
      RECT 44.595 4.982 44.61 5.185 ;
      RECT 44.6 4.191 44.605 4.933 ;
      RECT 44.595 4.169 44.6 4.943 ;
      RECT 44.56 4.079 44.595 5.18 ;
      RECT 44.545 3.957 44.56 5.18 ;
      RECT 44.54 3.91 44.545 5.18 ;
      RECT 44.515 3.835 44.54 5.18 ;
      RECT 44.5 3.75 44.515 5.18 ;
      RECT 44.495 3.697 44.5 5.18 ;
      RECT 44.49 3.677 44.495 5.18 ;
      RECT 44.485 3.652 44.49 4.414 ;
      RECT 44.47 4.612 44.49 5.18 ;
      RECT 44.48 3.63 44.485 4.391 ;
      RECT 44.47 3.582 44.48 4.356 ;
      RECT 44.465 3.545 44.47 4.322 ;
      RECT 44.465 4.692 44.47 5.18 ;
      RECT 44.45 3.522 44.465 4.277 ;
      RECT 44.445 4.79 44.465 5.18 ;
      RECT 44.395 3.41 44.45 4.119 ;
      RECT 44.44 4.912 44.445 5.18 ;
      RECT 44.38 3.41 44.395 3.958 ;
      RECT 44.375 3.41 44.38 3.91 ;
      RECT 44.37 3.41 44.375 3.898 ;
      RECT 44.325 3.41 44.37 3.835 ;
      RECT 44.3 3.41 44.325 3.753 ;
      RECT 44.285 3.41 44.3 3.705 ;
      RECT 44.28 3.41 44.285 3.675 ;
      RECT 46.67 3.455 46.93 3.715 ;
      RECT 46.665 3.455 46.93 3.663 ;
      RECT 46.66 3.455 46.93 3.633 ;
      RECT 46.635 3.325 46.915 3.605 ;
      RECT 35.185 9.095 35.535 9.445 ;
      RECT 46.155 9.05 46.505 9.4 ;
      RECT 35.185 9.125 46.505 9.325 ;
      RECT 45.675 5.005 45.955 5.285 ;
      RECT 45.715 4.96 45.98 5.22 ;
      RECT 45.705 4.995 45.98 5.22 ;
      RECT 45.71 4.98 45.955 5.285 ;
      RECT 45.715 4.957 45.925 5.285 ;
      RECT 45.715 4.955 45.91 5.285 ;
      RECT 45.755 4.945 45.91 5.285 ;
      RECT 45.725 4.95 45.91 5.285 ;
      RECT 45.755 4.942 45.855 5.285 ;
      RECT 45.78 4.935 45.855 5.285 ;
      RECT 45.76 4.937 45.855 5.285 ;
      RECT 45.09 4.45 45.35 4.71 ;
      RECT 45.14 4.442 45.33 4.71 ;
      RECT 45.145 4.362 45.33 4.71 ;
      RECT 45.265 3.75 45.33 4.71 ;
      RECT 45.17 4.147 45.33 4.71 ;
      RECT 45.245 3.835 45.33 4.71 ;
      RECT 45.28 3.46 45.416 4.188 ;
      RECT 45.225 3.957 45.416 4.188 ;
      RECT 45.24 3.897 45.33 4.71 ;
      RECT 45.28 3.46 45.44 3.853 ;
      RECT 45.28 3.46 45.45 3.75 ;
      RECT 45.27 3.46 45.53 3.72 ;
      RECT 43.605 4.86 43.65 5.12 ;
      RECT 43.51 3.395 43.655 3.655 ;
      RECT 44.015 4.017 44.025 4.108 ;
      RECT 44 3.955 44.015 4.164 ;
      RECT 43.995 3.902 44 4.21 ;
      RECT 43.945 3.849 43.995 4.336 ;
      RECT 43.94 3.804 43.945 4.483 ;
      RECT 43.93 3.792 43.94 4.525 ;
      RECT 43.895 3.756 43.93 4.63 ;
      RECT 43.89 3.724 43.895 4.736 ;
      RECT 43.875 3.706 43.89 4.781 ;
      RECT 43.87 3.689 43.875 4.015 ;
      RECT 43.865 4.07 43.875 4.838 ;
      RECT 43.86 3.675 43.87 3.988 ;
      RECT 43.855 4.125 43.865 5.12 ;
      RECT 43.85 3.661 43.86 3.973 ;
      RECT 43.85 4.175 43.855 5.12 ;
      RECT 43.835 3.638 43.85 3.953 ;
      RECT 43.815 4.297 43.85 5.12 ;
      RECT 43.83 3.62 43.835 3.935 ;
      RECT 43.825 3.612 43.83 3.925 ;
      RECT 43.795 3.58 43.825 3.889 ;
      RECT 43.805 4.425 43.815 5.12 ;
      RECT 43.8 4.452 43.805 5.12 ;
      RECT 43.795 4.502 43.8 5.12 ;
      RECT 43.785 3.546 43.795 3.854 ;
      RECT 43.745 4.57 43.795 5.12 ;
      RECT 43.77 3.523 43.785 3.83 ;
      RECT 43.745 3.395 43.77 3.793 ;
      RECT 43.74 3.395 43.745 3.765 ;
      RECT 43.71 4.67 43.745 5.12 ;
      RECT 43.735 3.395 43.74 3.758 ;
      RECT 43.73 3.395 43.735 3.748 ;
      RECT 43.715 3.395 43.73 3.733 ;
      RECT 43.7 3.395 43.715 3.705 ;
      RECT 43.665 4.775 43.71 5.12 ;
      RECT 43.685 3.395 43.7 3.678 ;
      RECT 43.655 3.395 43.685 3.663 ;
      RECT 43.65 4.847 43.665 5.12 ;
      RECT 43.575 3.93 43.615 4.19 ;
      RECT 43.35 3.877 43.355 4.135 ;
      RECT 39.305 3.355 39.565 3.615 ;
      RECT 39.305 3.38 39.58 3.595 ;
      RECT 41.695 3.205 41.7 3.35 ;
      RECT 43.565 3.925 43.575 4.19 ;
      RECT 43.545 3.917 43.565 4.19 ;
      RECT 43.527 3.913 43.545 4.19 ;
      RECT 43.441 3.902 43.527 4.19 ;
      RECT 43.355 3.885 43.441 4.19 ;
      RECT 43.3 3.872 43.35 4.12 ;
      RECT 43.266 3.864 43.3 4.095 ;
      RECT 43.18 3.853 43.266 4.06 ;
      RECT 43.145 3.83 43.18 4.025 ;
      RECT 43.135 3.792 43.145 4.011 ;
      RECT 43.13 3.765 43.135 4.007 ;
      RECT 43.125 3.752 43.13 4.004 ;
      RECT 43.115 3.732 43.125 4 ;
      RECT 43.11 3.707 43.115 3.996 ;
      RECT 43.085 3.662 43.11 3.99 ;
      RECT 43.075 3.603 43.085 3.982 ;
      RECT 43.065 3.571 43.075 3.973 ;
      RECT 43.045 3.523 43.065 3.953 ;
      RECT 43.04 3.483 43.045 3.923 ;
      RECT 43.025 3.457 43.04 3.897 ;
      RECT 43.02 3.435 43.025 3.873 ;
      RECT 43.005 3.407 43.02 3.849 ;
      RECT 42.99 3.38 43.005 3.813 ;
      RECT 42.975 3.357 42.99 3.775 ;
      RECT 42.97 3.347 42.975 3.75 ;
      RECT 42.96 3.34 42.97 3.733 ;
      RECT 42.945 3.327 42.96 3.703 ;
      RECT 42.94 3.317 42.945 3.678 ;
      RECT 42.935 3.312 42.94 3.665 ;
      RECT 42.925 3.305 42.935 3.645 ;
      RECT 42.92 3.298 42.925 3.63 ;
      RECT 42.895 3.291 42.92 3.588 ;
      RECT 42.88 3.281 42.895 3.538 ;
      RECT 42.87 3.276 42.88 3.508 ;
      RECT 42.86 3.272 42.87 3.483 ;
      RECT 42.845 3.269 42.86 3.473 ;
      RECT 42.795 3.266 42.845 3.458 ;
      RECT 42.775 3.264 42.795 3.443 ;
      RECT 42.726 3.262 42.775 3.438 ;
      RECT 42.64 3.258 42.726 3.433 ;
      RECT 42.601 3.255 42.64 3.429 ;
      RECT 42.515 3.251 42.601 3.424 ;
      RECT 42.465 3.248 42.515 3.418 ;
      RECT 42.416 3.245 42.465 3.413 ;
      RECT 42.33 3.242 42.416 3.408 ;
      RECT 42.326 3.24 42.33 3.405 ;
      RECT 42.24 3.237 42.326 3.4 ;
      RECT 42.191 3.233 42.24 3.393 ;
      RECT 42.105 3.23 42.191 3.388 ;
      RECT 42.081 3.227 42.105 3.384 ;
      RECT 41.995 3.225 42.081 3.379 ;
      RECT 41.93 3.221 41.995 3.372 ;
      RECT 41.927 3.22 41.93 3.369 ;
      RECT 41.841 3.217 41.927 3.366 ;
      RECT 41.755 3.211 41.841 3.359 ;
      RECT 41.725 3.207 41.755 3.355 ;
      RECT 41.7 3.205 41.725 3.353 ;
      RECT 41.645 3.202 41.695 3.35 ;
      RECT 41.565 3.201 41.645 3.35 ;
      RECT 41.51 3.203 41.565 3.353 ;
      RECT 41.495 3.204 41.51 3.357 ;
      RECT 41.44 3.212 41.495 3.367 ;
      RECT 41.41 3.22 41.44 3.38 ;
      RECT 41.391 3.221 41.41 3.386 ;
      RECT 41.305 3.224 41.391 3.391 ;
      RECT 41.235 3.229 41.305 3.4 ;
      RECT 41.216 3.232 41.235 3.406 ;
      RECT 41.13 3.236 41.216 3.411 ;
      RECT 41.09 3.24 41.13 3.418 ;
      RECT 41.081 3.242 41.09 3.421 ;
      RECT 40.995 3.246 41.081 3.426 ;
      RECT 40.992 3.249 40.995 3.43 ;
      RECT 40.906 3.252 40.992 3.434 ;
      RECT 40.82 3.258 40.906 3.442 ;
      RECT 40.796 3.262 40.82 3.446 ;
      RECT 40.71 3.266 40.796 3.451 ;
      RECT 40.665 3.271 40.71 3.458 ;
      RECT 40.585 3.276 40.665 3.465 ;
      RECT 40.505 3.282 40.585 3.48 ;
      RECT 40.48 3.286 40.505 3.493 ;
      RECT 40.415 3.289 40.48 3.505 ;
      RECT 40.36 3.294 40.415 3.52 ;
      RECT 40.33 3.297 40.36 3.538 ;
      RECT 40.32 3.299 40.33 3.551 ;
      RECT 40.26 3.314 40.32 3.561 ;
      RECT 40.245 3.331 40.26 3.57 ;
      RECT 40.24 3.34 40.245 3.57 ;
      RECT 40.23 3.35 40.24 3.57 ;
      RECT 40.22 3.367 40.23 3.57 ;
      RECT 40.2 3.377 40.22 3.571 ;
      RECT 40.155 3.387 40.2 3.572 ;
      RECT 40.12 3.396 40.155 3.574 ;
      RECT 40.055 3.401 40.12 3.576 ;
      RECT 39.975 3.402 40.055 3.579 ;
      RECT 39.971 3.4 39.975 3.58 ;
      RECT 39.885 3.397 39.971 3.582 ;
      RECT 39.838 3.394 39.885 3.584 ;
      RECT 39.752 3.39 39.838 3.587 ;
      RECT 39.666 3.386 39.752 3.59 ;
      RECT 39.58 3.382 39.666 3.594 ;
      RECT 42.965 5.005 42.995 5.285 ;
      RECT 42.715 4.895 42.735 5.285 ;
      RECT 42.67 4.895 42.735 5.155 ;
      RECT 42.5 3.52 42.535 3.78 ;
      RECT 42.275 3.52 42.335 3.78 ;
      RECT 42.955 4.985 42.965 5.285 ;
      RECT 42.95 4.945 42.955 5.285 ;
      RECT 42.935 4.9 42.95 5.285 ;
      RECT 42.93 4.865 42.935 5.285 ;
      RECT 42.925 4.845 42.93 5.285 ;
      RECT 42.895 4.772 42.925 5.285 ;
      RECT 42.875 4.67 42.895 5.285 ;
      RECT 42.865 4.6 42.875 5.285 ;
      RECT 42.82 4.54 42.865 5.285 ;
      RECT 42.735 4.501 42.82 5.285 ;
      RECT 42.73 4.492 42.735 4.865 ;
      RECT 42.72 4.491 42.73 4.848 ;
      RECT 42.695 4.472 42.72 4.818 ;
      RECT 42.69 4.447 42.695 4.797 ;
      RECT 42.68 4.425 42.69 4.788 ;
      RECT 42.675 4.396 42.68 4.778 ;
      RECT 42.635 4.322 42.675 4.75 ;
      RECT 42.615 4.223 42.635 4.715 ;
      RECT 42.6 4.159 42.615 4.698 ;
      RECT 42.57 4.083 42.6 4.67 ;
      RECT 42.55 3.998 42.57 4.643 ;
      RECT 42.51 3.894 42.55 4.55 ;
      RECT 42.505 3.815 42.51 4.458 ;
      RECT 42.5 3.798 42.505 4.435 ;
      RECT 42.495 3.52 42.5 4.415 ;
      RECT 42.465 3.52 42.495 4.353 ;
      RECT 42.46 3.52 42.465 4.285 ;
      RECT 42.45 3.52 42.46 4.25 ;
      RECT 42.44 3.52 42.45 4.215 ;
      RECT 42.375 3.52 42.44 4.07 ;
      RECT 42.37 3.52 42.375 3.94 ;
      RECT 42.34 3.52 42.37 3.873 ;
      RECT 42.335 3.52 42.34 3.798 ;
      RECT 41.515 4.445 41.795 4.725 ;
      RECT 41.555 4.425 41.815 4.685 ;
      RECT 41.545 4.435 41.815 4.685 ;
      RECT 41.555 4.362 41.77 4.725 ;
      RECT 41.61 4.285 41.765 4.725 ;
      RECT 41.615 4.07 41.765 4.725 ;
      RECT 41.605 3.872 41.755 4.123 ;
      RECT 41.595 3.872 41.755 3.99 ;
      RECT 41.59 3.75 41.75 3.893 ;
      RECT 41.575 3.75 41.75 3.798 ;
      RECT 41.57 3.46 41.745 3.775 ;
      RECT 41.555 3.46 41.745 3.745 ;
      RECT 41.515 3.46 41.775 3.72 ;
      RECT 41.425 4.93 41.505 5.19 ;
      RECT 40.83 3.65 40.835 3.915 ;
      RECT 40.71 3.65 40.835 3.91 ;
      RECT 41.385 4.895 41.425 5.19 ;
      RECT 41.34 4.817 41.385 5.19 ;
      RECT 41.32 4.745 41.34 5.19 ;
      RECT 41.31 4.697 41.32 5.19 ;
      RECT 41.275 4.63 41.31 5.19 ;
      RECT 41.245 4.53 41.275 5.19 ;
      RECT 41.225 4.455 41.245 4.99 ;
      RECT 41.215 4.405 41.225 4.945 ;
      RECT 41.21 4.382 41.215 4.918 ;
      RECT 41.205 4.367 41.21 4.905 ;
      RECT 41.2 4.352 41.205 4.883 ;
      RECT 41.195 4.337 41.2 4.865 ;
      RECT 41.17 4.292 41.195 4.82 ;
      RECT 41.16 4.24 41.17 4.763 ;
      RECT 41.15 4.21 41.16 4.73 ;
      RECT 41.14 4.175 41.15 4.698 ;
      RECT 41.105 4.107 41.14 4.63 ;
      RECT 41.1 4.046 41.105 4.565 ;
      RECT 41.09 4.034 41.1 4.545 ;
      RECT 41.085 4.022 41.09 4.525 ;
      RECT 41.08 4.014 41.085 4.513 ;
      RECT 41.075 4.006 41.08 4.493 ;
      RECT 41.065 3.994 41.075 4.465 ;
      RECT 41.055 3.978 41.065 4.435 ;
      RECT 41.03 3.95 41.055 4.373 ;
      RECT 41.02 3.921 41.03 4.318 ;
      RECT 41.005 3.9 41.02 4.278 ;
      RECT 41 3.884 41.005 4.25 ;
      RECT 40.995 3.872 41 4.24 ;
      RECT 40.99 3.867 40.995 4.213 ;
      RECT 40.985 3.86 40.99 4.2 ;
      RECT 40.97 3.843 40.985 4.173 ;
      RECT 40.96 3.65 40.97 4.133 ;
      RECT 40.95 3.65 40.96 4.1 ;
      RECT 40.94 3.65 40.95 4.075 ;
      RECT 40.87 3.65 40.94 4.01 ;
      RECT 40.86 3.65 40.87 3.958 ;
      RECT 40.845 3.65 40.86 3.94 ;
      RECT 40.835 3.65 40.845 3.925 ;
      RECT 40.665 4.52 40.925 4.78 ;
      RECT 39.2 4.555 39.205 4.762 ;
      RECT 38.835 4.445 38.91 4.76 ;
      RECT 38.65 4.5 38.805 4.76 ;
      RECT 38.835 4.445 38.94 4.725 ;
      RECT 40.65 4.617 40.665 4.778 ;
      RECT 40.625 4.625 40.65 4.783 ;
      RECT 40.6 4.632 40.625 4.788 ;
      RECT 40.537 4.643 40.6 4.797 ;
      RECT 40.451 4.662 40.537 4.814 ;
      RECT 40.365 4.684 40.451 4.833 ;
      RECT 40.35 4.697 40.365 4.844 ;
      RECT 40.31 4.705 40.35 4.851 ;
      RECT 40.29 4.71 40.31 4.858 ;
      RECT 40.252 4.711 40.29 4.861 ;
      RECT 40.166 4.714 40.252 4.862 ;
      RECT 40.08 4.718 40.166 4.863 ;
      RECT 40.031 4.72 40.08 4.865 ;
      RECT 39.945 4.72 40.031 4.867 ;
      RECT 39.905 4.715 39.945 4.869 ;
      RECT 39.895 4.709 39.905 4.87 ;
      RECT 39.855 4.704 39.895 4.867 ;
      RECT 39.845 4.697 39.855 4.863 ;
      RECT 39.83 4.693 39.845 4.861 ;
      RECT 39.813 4.689 39.83 4.859 ;
      RECT 39.727 4.679 39.813 4.851 ;
      RECT 39.641 4.661 39.727 4.837 ;
      RECT 39.555 4.644 39.641 4.823 ;
      RECT 39.53 4.632 39.555 4.814 ;
      RECT 39.46 4.622 39.53 4.807 ;
      RECT 39.415 4.61 39.46 4.798 ;
      RECT 39.355 4.597 39.415 4.79 ;
      RECT 39.35 4.589 39.355 4.785 ;
      RECT 39.315 4.584 39.35 4.783 ;
      RECT 39.26 4.575 39.315 4.776 ;
      RECT 39.22 4.564 39.26 4.768 ;
      RECT 39.205 4.557 39.22 4.764 ;
      RECT 39.185 4.55 39.2 4.761 ;
      RECT 39.17 4.54 39.185 4.759 ;
      RECT 39.155 4.527 39.17 4.756 ;
      RECT 39.13 4.51 39.155 4.752 ;
      RECT 39.115 4.492 39.13 4.749 ;
      RECT 39.09 4.445 39.115 4.747 ;
      RECT 39.066 4.445 39.09 4.744 ;
      RECT 38.98 4.445 39.066 4.736 ;
      RECT 38.94 4.445 38.98 4.728 ;
      RECT 38.805 4.492 38.835 4.76 ;
      RECT 40.485 4.075 40.745 4.335 ;
      RECT 40.445 4.075 40.745 4.213 ;
      RECT 40.41 4.075 40.745 4.198 ;
      RECT 40.355 4.075 40.745 4.178 ;
      RECT 40.275 3.885 40.555 4.165 ;
      RECT 40.275 4.067 40.625 4.165 ;
      RECT 40.275 4.01 40.61 4.165 ;
      RECT 40.275 3.957 40.56 4.165 ;
      RECT 37.435 4.244 37.45 4.7 ;
      RECT 37.43 4.316 37.536 4.698 ;
      RECT 37.45 3.41 37.585 4.696 ;
      RECT 37.435 4.26 37.59 4.695 ;
      RECT 37.435 4.31 37.595 4.693 ;
      RECT 37.42 4.375 37.595 4.692 ;
      RECT 37.43 4.367 37.6 4.689 ;
      RECT 37.41 4.415 37.6 4.684 ;
      RECT 37.41 4.415 37.615 4.681 ;
      RECT 37.405 4.415 37.615 4.678 ;
      RECT 37.38 4.415 37.64 4.675 ;
      RECT 37.45 3.41 37.61 4.063 ;
      RECT 37.445 3.41 37.61 4.035 ;
      RECT 37.44 3.41 37.61 3.863 ;
      RECT 37.44 3.41 37.63 3.803 ;
      RECT 37.395 3.41 37.655 3.67 ;
      RECT 36.875 3.885 37.155 4.165 ;
      RECT 36.865 3.9 37.155 4.16 ;
      RECT 36.82 3.962 37.155 4.158 ;
      RECT 36.895 3.877 37.06 4.165 ;
      RECT 36.895 3.862 37.016 4.165 ;
      RECT 36.93 3.855 37.016 4.165 ;
      RECT 36.395 5.005 36.675 5.285 ;
      RECT 36.355 4.967 36.65 5.078 ;
      RECT 36.34 4.917 36.63 4.973 ;
      RECT 36.285 4.68 36.545 4.94 ;
      RECT 36.285 4.882 36.625 4.94 ;
      RECT 36.285 4.822 36.62 4.94 ;
      RECT 36.285 4.772 36.6 4.94 ;
      RECT 36.285 4.752 36.595 4.94 ;
      RECT 36.285 4.73 36.59 4.94 ;
      RECT 36.285 4.715 36.56 4.94 ;
      RECT 32.005 8.66 32.325 8.98 ;
      RECT 32.035 8.13 32.205 8.98 ;
      RECT 32.035 8.13 32.21 8.48 ;
      RECT 32.035 8.13 33.01 8.305 ;
      RECT 32.835 3.26 33.01 8.305 ;
      RECT 32.78 3.26 33.13 3.61 ;
      RECT 32.805 9.09 33.13 9.415 ;
      RECT 31.69 9.18 33.13 9.35 ;
      RECT 31.69 3.69 31.85 9.35 ;
      RECT 32.005 3.66 32.325 3.98 ;
      RECT 31.69 3.69 32.325 3.86 ;
      RECT 30.37 2.435 30.745 2.805 ;
      RECT 22.28 2.255 22.655 2.625 ;
      RECT 20.845 2.255 21.22 2.625 ;
      RECT 20.845 2.375 30.675 2.545 ;
      RECT 26.79 5.655 30.645 5.825 ;
      RECT 30.475 4.72 30.645 5.825 ;
      RECT 26.79 4.965 26.96 5.825 ;
      RECT 26.75 5.005 27.03 5.285 ;
      RECT 26.77 4.965 27.03 5.285 ;
      RECT 26.41 4.92 26.515 5.18 ;
      RECT 30.385 4.725 30.735 5.075 ;
      RECT 26.265 3.41 26.355 3.67 ;
      RECT 26.805 4.475 26.81 4.515 ;
      RECT 26.8 4.465 26.805 4.6 ;
      RECT 26.795 4.455 26.8 4.693 ;
      RECT 26.785 4.435 26.795 4.749 ;
      RECT 26.705 4.363 26.785 4.829 ;
      RECT 26.74 5.007 26.75 5.232 ;
      RECT 26.735 5.004 26.74 5.227 ;
      RECT 26.72 5.001 26.735 5.22 ;
      RECT 26.685 4.995 26.72 5.202 ;
      RECT 26.7 4.298 26.705 4.903 ;
      RECT 26.68 4.249 26.7 4.918 ;
      RECT 26.67 4.982 26.685 5.185 ;
      RECT 26.675 4.191 26.68 4.933 ;
      RECT 26.67 4.169 26.675 4.943 ;
      RECT 26.635 4.079 26.67 5.18 ;
      RECT 26.62 3.957 26.635 5.18 ;
      RECT 26.615 3.91 26.62 5.18 ;
      RECT 26.59 3.835 26.615 5.18 ;
      RECT 26.575 3.75 26.59 5.18 ;
      RECT 26.57 3.697 26.575 5.18 ;
      RECT 26.565 3.677 26.57 5.18 ;
      RECT 26.56 3.652 26.565 4.414 ;
      RECT 26.545 4.612 26.565 5.18 ;
      RECT 26.555 3.63 26.56 4.391 ;
      RECT 26.545 3.582 26.555 4.356 ;
      RECT 26.54 3.545 26.545 4.322 ;
      RECT 26.54 4.692 26.545 5.18 ;
      RECT 26.525 3.522 26.54 4.277 ;
      RECT 26.52 4.79 26.54 5.18 ;
      RECT 26.47 3.41 26.525 4.119 ;
      RECT 26.515 4.912 26.52 5.18 ;
      RECT 26.455 3.41 26.47 3.958 ;
      RECT 26.45 3.41 26.455 3.91 ;
      RECT 26.445 3.41 26.45 3.898 ;
      RECT 26.4 3.41 26.445 3.835 ;
      RECT 26.375 3.41 26.4 3.753 ;
      RECT 26.36 3.41 26.375 3.705 ;
      RECT 26.355 3.41 26.36 3.675 ;
      RECT 28.745 3.455 29.005 3.715 ;
      RECT 28.74 3.455 29.005 3.663 ;
      RECT 28.735 3.455 29.005 3.633 ;
      RECT 28.71 3.325 28.99 3.605 ;
      RECT 16.56 9.43 16.85 9.78 ;
      RECT 16.56 9.49 17.695 9.66 ;
      RECT 17.525 9.12 17.695 9.66 ;
      RECT 28.25 9.04 28.42 9.395 ;
      RECT 28.2 9.04 28.55 9.39 ;
      RECT 17.525 9.12 28.55 9.29 ;
      RECT 27.75 5.005 28.03 5.285 ;
      RECT 27.79 4.96 28.055 5.22 ;
      RECT 27.78 4.995 28.055 5.22 ;
      RECT 27.785 4.98 28.03 5.285 ;
      RECT 27.79 4.957 28 5.285 ;
      RECT 27.79 4.955 27.985 5.285 ;
      RECT 27.83 4.945 27.985 5.285 ;
      RECT 27.8 4.95 27.985 5.285 ;
      RECT 27.83 4.942 27.93 5.285 ;
      RECT 27.855 4.935 27.93 5.285 ;
      RECT 27.835 4.937 27.93 5.285 ;
      RECT 27.165 4.45 27.425 4.71 ;
      RECT 27.215 4.442 27.405 4.71 ;
      RECT 27.22 4.362 27.405 4.71 ;
      RECT 27.34 3.75 27.405 4.71 ;
      RECT 27.245 4.147 27.405 4.71 ;
      RECT 27.32 3.835 27.405 4.71 ;
      RECT 27.355 3.46 27.491 4.188 ;
      RECT 27.3 3.957 27.491 4.188 ;
      RECT 27.315 3.897 27.405 4.71 ;
      RECT 27.355 3.46 27.515 3.853 ;
      RECT 27.355 3.46 27.525 3.75 ;
      RECT 27.345 3.46 27.605 3.72 ;
      RECT 25.68 4.86 25.725 5.12 ;
      RECT 25.585 3.395 25.73 3.655 ;
      RECT 26.09 4.017 26.1 4.108 ;
      RECT 26.075 3.955 26.09 4.164 ;
      RECT 26.07 3.902 26.075 4.21 ;
      RECT 26.02 3.849 26.07 4.336 ;
      RECT 26.015 3.804 26.02 4.483 ;
      RECT 26.005 3.792 26.015 4.525 ;
      RECT 25.97 3.756 26.005 4.63 ;
      RECT 25.965 3.724 25.97 4.736 ;
      RECT 25.95 3.706 25.965 4.781 ;
      RECT 25.945 3.689 25.95 4.015 ;
      RECT 25.94 4.07 25.95 4.838 ;
      RECT 25.935 3.675 25.945 3.988 ;
      RECT 25.93 4.125 25.94 5.12 ;
      RECT 25.925 3.661 25.935 3.973 ;
      RECT 25.925 4.175 25.93 5.12 ;
      RECT 25.91 3.638 25.925 3.953 ;
      RECT 25.89 4.297 25.925 5.12 ;
      RECT 25.905 3.62 25.91 3.935 ;
      RECT 25.9 3.612 25.905 3.925 ;
      RECT 25.87 3.58 25.9 3.889 ;
      RECT 25.88 4.425 25.89 5.12 ;
      RECT 25.875 4.452 25.88 5.12 ;
      RECT 25.87 4.502 25.875 5.12 ;
      RECT 25.86 3.546 25.87 3.854 ;
      RECT 25.82 4.57 25.87 5.12 ;
      RECT 25.845 3.523 25.86 3.83 ;
      RECT 25.82 3.395 25.845 3.793 ;
      RECT 25.815 3.395 25.82 3.765 ;
      RECT 25.785 4.67 25.82 5.12 ;
      RECT 25.81 3.395 25.815 3.758 ;
      RECT 25.805 3.395 25.81 3.748 ;
      RECT 25.79 3.395 25.805 3.733 ;
      RECT 25.775 3.395 25.79 3.705 ;
      RECT 25.74 4.775 25.785 5.12 ;
      RECT 25.76 3.395 25.775 3.678 ;
      RECT 25.73 3.395 25.76 3.663 ;
      RECT 25.725 4.847 25.74 5.12 ;
      RECT 25.65 3.93 25.69 4.19 ;
      RECT 25.425 3.877 25.43 4.135 ;
      RECT 21.38 3.355 21.64 3.615 ;
      RECT 21.38 3.38 21.655 3.595 ;
      RECT 23.77 3.205 23.775 3.35 ;
      RECT 25.64 3.925 25.65 4.19 ;
      RECT 25.62 3.917 25.64 4.19 ;
      RECT 25.602 3.913 25.62 4.19 ;
      RECT 25.516 3.902 25.602 4.19 ;
      RECT 25.43 3.885 25.516 4.19 ;
      RECT 25.375 3.872 25.425 4.12 ;
      RECT 25.341 3.864 25.375 4.095 ;
      RECT 25.255 3.853 25.341 4.06 ;
      RECT 25.22 3.83 25.255 4.025 ;
      RECT 25.21 3.792 25.22 4.011 ;
      RECT 25.205 3.765 25.21 4.007 ;
      RECT 25.2 3.752 25.205 4.004 ;
      RECT 25.19 3.732 25.2 4 ;
      RECT 25.185 3.707 25.19 3.996 ;
      RECT 25.16 3.662 25.185 3.99 ;
      RECT 25.15 3.603 25.16 3.982 ;
      RECT 25.14 3.571 25.15 3.973 ;
      RECT 25.12 3.523 25.14 3.953 ;
      RECT 25.115 3.483 25.12 3.923 ;
      RECT 25.1 3.457 25.115 3.897 ;
      RECT 25.095 3.435 25.1 3.873 ;
      RECT 25.08 3.407 25.095 3.849 ;
      RECT 25.065 3.38 25.08 3.813 ;
      RECT 25.05 3.357 25.065 3.775 ;
      RECT 25.045 3.347 25.05 3.75 ;
      RECT 25.035 3.34 25.045 3.733 ;
      RECT 25.02 3.327 25.035 3.703 ;
      RECT 25.015 3.317 25.02 3.678 ;
      RECT 25.01 3.312 25.015 3.665 ;
      RECT 25 3.305 25.01 3.645 ;
      RECT 24.995 3.298 25 3.63 ;
      RECT 24.97 3.291 24.995 3.588 ;
      RECT 24.955 3.281 24.97 3.538 ;
      RECT 24.945 3.276 24.955 3.508 ;
      RECT 24.935 3.272 24.945 3.483 ;
      RECT 24.92 3.269 24.935 3.473 ;
      RECT 24.87 3.266 24.92 3.458 ;
      RECT 24.85 3.264 24.87 3.443 ;
      RECT 24.801 3.262 24.85 3.438 ;
      RECT 24.715 3.258 24.801 3.433 ;
      RECT 24.676 3.255 24.715 3.429 ;
      RECT 24.59 3.251 24.676 3.424 ;
      RECT 24.54 3.248 24.59 3.418 ;
      RECT 24.491 3.245 24.54 3.413 ;
      RECT 24.405 3.242 24.491 3.408 ;
      RECT 24.401 3.24 24.405 3.405 ;
      RECT 24.315 3.237 24.401 3.4 ;
      RECT 24.266 3.233 24.315 3.393 ;
      RECT 24.18 3.23 24.266 3.388 ;
      RECT 24.156 3.227 24.18 3.384 ;
      RECT 24.07 3.225 24.156 3.379 ;
      RECT 24.005 3.221 24.07 3.372 ;
      RECT 24.002 3.22 24.005 3.369 ;
      RECT 23.916 3.217 24.002 3.366 ;
      RECT 23.83 3.211 23.916 3.359 ;
      RECT 23.8 3.207 23.83 3.355 ;
      RECT 23.775 3.205 23.8 3.353 ;
      RECT 23.72 3.202 23.77 3.35 ;
      RECT 23.64 3.201 23.72 3.35 ;
      RECT 23.585 3.203 23.64 3.353 ;
      RECT 23.57 3.204 23.585 3.357 ;
      RECT 23.515 3.212 23.57 3.367 ;
      RECT 23.485 3.22 23.515 3.38 ;
      RECT 23.466 3.221 23.485 3.386 ;
      RECT 23.38 3.224 23.466 3.391 ;
      RECT 23.31 3.229 23.38 3.4 ;
      RECT 23.291 3.232 23.31 3.406 ;
      RECT 23.205 3.236 23.291 3.411 ;
      RECT 23.165 3.24 23.205 3.418 ;
      RECT 23.156 3.242 23.165 3.421 ;
      RECT 23.07 3.246 23.156 3.426 ;
      RECT 23.067 3.249 23.07 3.43 ;
      RECT 22.981 3.252 23.067 3.434 ;
      RECT 22.895 3.258 22.981 3.442 ;
      RECT 22.871 3.262 22.895 3.446 ;
      RECT 22.785 3.266 22.871 3.451 ;
      RECT 22.74 3.271 22.785 3.458 ;
      RECT 22.66 3.276 22.74 3.465 ;
      RECT 22.58 3.282 22.66 3.48 ;
      RECT 22.555 3.286 22.58 3.493 ;
      RECT 22.49 3.289 22.555 3.505 ;
      RECT 22.435 3.294 22.49 3.52 ;
      RECT 22.405 3.297 22.435 3.538 ;
      RECT 22.395 3.299 22.405 3.551 ;
      RECT 22.335 3.314 22.395 3.561 ;
      RECT 22.32 3.331 22.335 3.57 ;
      RECT 22.315 3.34 22.32 3.57 ;
      RECT 22.305 3.35 22.315 3.57 ;
      RECT 22.295 3.367 22.305 3.57 ;
      RECT 22.275 3.377 22.295 3.571 ;
      RECT 22.23 3.387 22.275 3.572 ;
      RECT 22.195 3.396 22.23 3.574 ;
      RECT 22.13 3.401 22.195 3.576 ;
      RECT 22.05 3.402 22.13 3.579 ;
      RECT 22.046 3.4 22.05 3.58 ;
      RECT 21.96 3.397 22.046 3.582 ;
      RECT 21.913 3.394 21.96 3.584 ;
      RECT 21.827 3.39 21.913 3.587 ;
      RECT 21.741 3.386 21.827 3.59 ;
      RECT 21.655 3.382 21.741 3.594 ;
      RECT 25.04 5.005 25.07 5.285 ;
      RECT 24.79 4.895 24.81 5.285 ;
      RECT 24.745 4.895 24.81 5.155 ;
      RECT 24.575 3.52 24.61 3.78 ;
      RECT 24.35 3.52 24.41 3.78 ;
      RECT 25.03 4.985 25.04 5.285 ;
      RECT 25.025 4.945 25.03 5.285 ;
      RECT 25.01 4.9 25.025 5.285 ;
      RECT 25.005 4.865 25.01 5.285 ;
      RECT 25 4.845 25.005 5.285 ;
      RECT 24.97 4.772 25 5.285 ;
      RECT 24.95 4.67 24.97 5.285 ;
      RECT 24.94 4.6 24.95 5.285 ;
      RECT 24.895 4.54 24.94 5.285 ;
      RECT 24.81 4.501 24.895 5.285 ;
      RECT 24.805 4.492 24.81 4.865 ;
      RECT 24.795 4.491 24.805 4.848 ;
      RECT 24.77 4.472 24.795 4.818 ;
      RECT 24.765 4.447 24.77 4.797 ;
      RECT 24.755 4.425 24.765 4.788 ;
      RECT 24.75 4.396 24.755 4.778 ;
      RECT 24.71 4.322 24.75 4.75 ;
      RECT 24.69 4.223 24.71 4.715 ;
      RECT 24.675 4.159 24.69 4.698 ;
      RECT 24.645 4.083 24.675 4.67 ;
      RECT 24.625 3.998 24.645 4.643 ;
      RECT 24.585 3.894 24.625 4.55 ;
      RECT 24.58 3.815 24.585 4.458 ;
      RECT 24.575 3.798 24.58 4.435 ;
      RECT 24.57 3.52 24.575 4.415 ;
      RECT 24.54 3.52 24.57 4.353 ;
      RECT 24.535 3.52 24.54 4.285 ;
      RECT 24.525 3.52 24.535 4.25 ;
      RECT 24.515 3.52 24.525 4.215 ;
      RECT 24.45 3.52 24.515 4.07 ;
      RECT 24.445 3.52 24.45 3.94 ;
      RECT 24.415 3.52 24.445 3.873 ;
      RECT 24.41 3.52 24.415 3.798 ;
      RECT 23.59 4.445 23.87 4.725 ;
      RECT 23.63 4.425 23.89 4.685 ;
      RECT 23.62 4.435 23.89 4.685 ;
      RECT 23.63 4.362 23.845 4.725 ;
      RECT 23.685 4.285 23.84 4.725 ;
      RECT 23.69 4.07 23.84 4.725 ;
      RECT 23.68 3.872 23.83 4.123 ;
      RECT 23.67 3.872 23.83 3.99 ;
      RECT 23.665 3.75 23.825 3.893 ;
      RECT 23.65 3.75 23.825 3.798 ;
      RECT 23.645 3.46 23.82 3.775 ;
      RECT 23.63 3.46 23.82 3.745 ;
      RECT 23.59 3.46 23.85 3.72 ;
      RECT 23.5 4.93 23.58 5.19 ;
      RECT 22.905 3.65 22.91 3.915 ;
      RECT 22.785 3.65 22.91 3.91 ;
      RECT 23.46 4.895 23.5 5.19 ;
      RECT 23.415 4.817 23.46 5.19 ;
      RECT 23.395 4.745 23.415 5.19 ;
      RECT 23.385 4.697 23.395 5.19 ;
      RECT 23.35 4.63 23.385 5.19 ;
      RECT 23.32 4.53 23.35 5.19 ;
      RECT 23.3 4.455 23.32 4.99 ;
      RECT 23.29 4.405 23.3 4.945 ;
      RECT 23.285 4.382 23.29 4.918 ;
      RECT 23.28 4.367 23.285 4.905 ;
      RECT 23.275 4.352 23.28 4.883 ;
      RECT 23.27 4.337 23.275 4.865 ;
      RECT 23.245 4.292 23.27 4.82 ;
      RECT 23.235 4.24 23.245 4.763 ;
      RECT 23.225 4.21 23.235 4.73 ;
      RECT 23.215 4.175 23.225 4.698 ;
      RECT 23.18 4.107 23.215 4.63 ;
      RECT 23.175 4.046 23.18 4.565 ;
      RECT 23.165 4.034 23.175 4.545 ;
      RECT 23.16 4.022 23.165 4.525 ;
      RECT 23.155 4.014 23.16 4.513 ;
      RECT 23.15 4.006 23.155 4.493 ;
      RECT 23.14 3.994 23.15 4.465 ;
      RECT 23.13 3.978 23.14 4.435 ;
      RECT 23.105 3.95 23.13 4.373 ;
      RECT 23.095 3.921 23.105 4.318 ;
      RECT 23.08 3.9 23.095 4.278 ;
      RECT 23.075 3.884 23.08 4.25 ;
      RECT 23.07 3.872 23.075 4.24 ;
      RECT 23.065 3.867 23.07 4.213 ;
      RECT 23.06 3.86 23.065 4.2 ;
      RECT 23.045 3.843 23.06 4.173 ;
      RECT 23.035 3.65 23.045 4.133 ;
      RECT 23.025 3.65 23.035 4.1 ;
      RECT 23.015 3.65 23.025 4.075 ;
      RECT 22.945 3.65 23.015 4.01 ;
      RECT 22.935 3.65 22.945 3.958 ;
      RECT 22.92 3.65 22.935 3.94 ;
      RECT 22.91 3.65 22.92 3.925 ;
      RECT 22.74 4.52 23 4.78 ;
      RECT 21.275 4.555 21.28 4.762 ;
      RECT 20.91 4.445 20.985 4.76 ;
      RECT 20.725 4.5 20.88 4.76 ;
      RECT 20.91 4.445 21.015 4.725 ;
      RECT 22.725 4.617 22.74 4.778 ;
      RECT 22.7 4.625 22.725 4.783 ;
      RECT 22.675 4.632 22.7 4.788 ;
      RECT 22.612 4.643 22.675 4.797 ;
      RECT 22.526 4.662 22.612 4.814 ;
      RECT 22.44 4.684 22.526 4.833 ;
      RECT 22.425 4.697 22.44 4.844 ;
      RECT 22.385 4.705 22.425 4.851 ;
      RECT 22.365 4.71 22.385 4.858 ;
      RECT 22.327 4.711 22.365 4.861 ;
      RECT 22.241 4.714 22.327 4.862 ;
      RECT 22.155 4.718 22.241 4.863 ;
      RECT 22.106 4.72 22.155 4.865 ;
      RECT 22.02 4.72 22.106 4.867 ;
      RECT 21.98 4.715 22.02 4.869 ;
      RECT 21.97 4.709 21.98 4.87 ;
      RECT 21.93 4.704 21.97 4.867 ;
      RECT 21.92 4.697 21.93 4.863 ;
      RECT 21.905 4.693 21.92 4.861 ;
      RECT 21.888 4.689 21.905 4.859 ;
      RECT 21.802 4.679 21.888 4.851 ;
      RECT 21.716 4.661 21.802 4.837 ;
      RECT 21.63 4.644 21.716 4.823 ;
      RECT 21.605 4.632 21.63 4.814 ;
      RECT 21.535 4.622 21.605 4.807 ;
      RECT 21.49 4.61 21.535 4.798 ;
      RECT 21.43 4.597 21.49 4.79 ;
      RECT 21.425 4.589 21.43 4.785 ;
      RECT 21.39 4.584 21.425 4.783 ;
      RECT 21.335 4.575 21.39 4.776 ;
      RECT 21.295 4.564 21.335 4.768 ;
      RECT 21.28 4.557 21.295 4.764 ;
      RECT 21.26 4.55 21.275 4.761 ;
      RECT 21.245 4.54 21.26 4.759 ;
      RECT 21.23 4.527 21.245 4.756 ;
      RECT 21.205 4.51 21.23 4.752 ;
      RECT 21.19 4.492 21.205 4.749 ;
      RECT 21.165 4.445 21.19 4.747 ;
      RECT 21.141 4.445 21.165 4.744 ;
      RECT 21.055 4.445 21.141 4.736 ;
      RECT 21.015 4.445 21.055 4.728 ;
      RECT 20.88 4.492 20.91 4.76 ;
      RECT 22.56 4.075 22.82 4.335 ;
      RECT 22.52 4.075 22.82 4.213 ;
      RECT 22.485 4.075 22.82 4.198 ;
      RECT 22.43 4.075 22.82 4.178 ;
      RECT 22.35 3.885 22.63 4.165 ;
      RECT 22.35 4.067 22.7 4.165 ;
      RECT 22.35 4.01 22.685 4.165 ;
      RECT 22.35 3.957 22.635 4.165 ;
      RECT 19.51 4.244 19.525 4.7 ;
      RECT 19.505 4.316 19.611 4.698 ;
      RECT 19.525 3.41 19.66 4.696 ;
      RECT 19.51 4.26 19.665 4.695 ;
      RECT 19.51 4.31 19.67 4.693 ;
      RECT 19.495 4.375 19.67 4.692 ;
      RECT 19.505 4.367 19.675 4.689 ;
      RECT 19.485 4.415 19.675 4.684 ;
      RECT 19.485 4.415 19.69 4.681 ;
      RECT 19.48 4.415 19.69 4.678 ;
      RECT 19.455 4.415 19.715 4.675 ;
      RECT 19.525 3.41 19.685 4.063 ;
      RECT 19.52 3.41 19.685 4.035 ;
      RECT 19.515 3.41 19.685 3.863 ;
      RECT 19.515 3.41 19.705 3.803 ;
      RECT 19.47 3.41 19.73 3.67 ;
      RECT 18.95 3.885 19.23 4.165 ;
      RECT 18.94 3.9 19.23 4.16 ;
      RECT 18.895 3.962 19.23 4.158 ;
      RECT 18.97 3.877 19.135 4.165 ;
      RECT 18.97 3.862 19.091 4.165 ;
      RECT 19.005 3.855 19.091 4.165 ;
      RECT 18.47 5.005 18.75 5.285 ;
      RECT 18.43 4.967 18.725 5.078 ;
      RECT 18.415 4.917 18.705 4.973 ;
      RECT 18.36 4.68 18.62 4.94 ;
      RECT 18.36 4.882 18.7 4.94 ;
      RECT 18.36 4.822 18.695 4.94 ;
      RECT 18.36 4.772 18.675 4.94 ;
      RECT 18.36 4.752 18.67 4.94 ;
      RECT 18.36 4.73 18.665 4.94 ;
      RECT 18.36 4.715 18.635 4.94 ;
      RECT 106.79 7.345 107.17 7.725 ;
      RECT 99.24 9.49 99.615 9.86 ;
      RECT 90.575 2.225 90.95 2.595 ;
      RECT 88.865 7.345 89.245 7.725 ;
      RECT 81.315 9.49 81.69 9.86 ;
      RECT 72.65 2.225 73.025 2.595 ;
      RECT 70.94 7.345 71.32 7.725 ;
      RECT 63.39 9.49 63.765 9.86 ;
      RECT 54.725 2.225 55.1 2.595 ;
      RECT 53.015 7.345 53.395 7.725 ;
      RECT 45.465 9.49 45.84 9.86 ;
      RECT 36.8 2.225 37.175 2.595 ;
      RECT 35.09 7.345 35.47 7.725 ;
      RECT 27.54 9.49 27.915 9.86 ;
      RECT 18.875 2.225 19.25 2.595 ;
    LAYER via1 ;
      RECT 106.96 9.81 107.11 9.96 ;
      RECT 106.905 7.46 107.055 7.61 ;
      RECT 104.595 9.175 104.745 9.325 ;
      RECT 104.58 3.36 104.73 3.51 ;
      RECT 103.79 3.745 103.94 3.895 ;
      RECT 103.79 8.76 103.94 8.91 ;
      RECT 102.185 2.545 102.335 2.695 ;
      RECT 102.185 4.825 102.335 4.975 ;
      RECT 100.5 3.51 100.65 3.66 ;
      RECT 100.26 9.15 100.41 9.3 ;
      RECT 99.55 5.015 99.7 5.165 ;
      RECT 99.355 9.6 99.505 9.75 ;
      RECT 99.1 3.515 99.25 3.665 ;
      RECT 98.92 4.505 99.07 4.655 ;
      RECT 98.525 5.02 98.675 5.17 ;
      RECT 98.165 4.975 98.315 5.125 ;
      RECT 98.02 3.465 98.17 3.615 ;
      RECT 97.435 4.915 97.585 5.065 ;
      RECT 97.34 3.45 97.49 3.6 ;
      RECT 97.185 3.985 97.335 4.135 ;
      RECT 96.5 4.95 96.65 5.1 ;
      RECT 96.105 3.575 96.255 3.725 ;
      RECT 95.385 4.48 95.535 4.63 ;
      RECT 95.345 3.515 95.495 3.665 ;
      RECT 95.075 4.985 95.225 5.135 ;
      RECT 94.54 3.705 94.69 3.855 ;
      RECT 94.495 4.575 94.645 4.725 ;
      RECT 94.315 4.13 94.465 4.28 ;
      RECT 93.135 3.41 93.285 3.56 ;
      RECT 92.48 4.555 92.63 4.705 ;
      RECT 91.225 3.465 91.375 3.615 ;
      RECT 91.21 4.47 91.36 4.62 ;
      RECT 90.695 3.955 90.845 4.105 ;
      RECT 90.115 4.735 90.265 4.885 ;
      RECT 89.015 9.195 89.165 9.345 ;
      RECT 88.98 7.46 89.13 7.61 ;
      RECT 86.67 9.175 86.82 9.325 ;
      RECT 86.655 3.36 86.805 3.51 ;
      RECT 85.865 3.745 86.015 3.895 ;
      RECT 85.865 8.76 86.015 8.91 ;
      RECT 84.26 2.545 84.41 2.695 ;
      RECT 84.26 4.825 84.41 4.975 ;
      RECT 82.575 3.51 82.725 3.66 ;
      RECT 82.055 9.15 82.205 9.3 ;
      RECT 81.625 5.015 81.775 5.165 ;
      RECT 81.43 9.6 81.58 9.75 ;
      RECT 81.175 3.515 81.325 3.665 ;
      RECT 80.995 4.505 81.145 4.655 ;
      RECT 80.6 5.02 80.75 5.17 ;
      RECT 80.24 4.975 80.39 5.125 ;
      RECT 80.095 3.465 80.245 3.615 ;
      RECT 79.51 4.915 79.66 5.065 ;
      RECT 79.415 3.45 79.565 3.6 ;
      RECT 79.26 3.985 79.41 4.135 ;
      RECT 78.575 4.95 78.725 5.1 ;
      RECT 78.18 3.575 78.33 3.725 ;
      RECT 77.46 4.48 77.61 4.63 ;
      RECT 77.42 3.515 77.57 3.665 ;
      RECT 77.15 4.985 77.3 5.135 ;
      RECT 76.615 3.705 76.765 3.855 ;
      RECT 76.57 4.575 76.72 4.725 ;
      RECT 76.39 4.13 76.54 4.28 ;
      RECT 75.21 3.41 75.36 3.56 ;
      RECT 74.555 4.555 74.705 4.705 ;
      RECT 73.3 3.465 73.45 3.615 ;
      RECT 73.285 4.47 73.435 4.62 ;
      RECT 72.77 3.955 72.92 4.105 ;
      RECT 72.19 4.735 72.34 4.885 ;
      RECT 71.09 9.195 71.24 9.345 ;
      RECT 71.055 7.46 71.205 7.61 ;
      RECT 68.745 9.175 68.895 9.325 ;
      RECT 68.73 3.36 68.88 3.51 ;
      RECT 67.94 3.745 68.09 3.895 ;
      RECT 67.94 8.76 68.09 8.91 ;
      RECT 66.335 2.545 66.485 2.695 ;
      RECT 66.335 4.825 66.485 4.975 ;
      RECT 64.65 3.51 64.8 3.66 ;
      RECT 64.185 9.15 64.335 9.3 ;
      RECT 63.7 5.015 63.85 5.165 ;
      RECT 63.505 9.6 63.655 9.75 ;
      RECT 63.25 3.515 63.4 3.665 ;
      RECT 63.07 4.505 63.22 4.655 ;
      RECT 62.675 5.02 62.825 5.17 ;
      RECT 62.315 4.975 62.465 5.125 ;
      RECT 62.17 3.465 62.32 3.615 ;
      RECT 61.585 4.915 61.735 5.065 ;
      RECT 61.49 3.45 61.64 3.6 ;
      RECT 61.335 3.985 61.485 4.135 ;
      RECT 60.65 4.95 60.8 5.1 ;
      RECT 60.255 3.575 60.405 3.725 ;
      RECT 59.535 4.48 59.685 4.63 ;
      RECT 59.495 3.515 59.645 3.665 ;
      RECT 59.225 4.985 59.375 5.135 ;
      RECT 58.69 3.705 58.84 3.855 ;
      RECT 58.645 4.575 58.795 4.725 ;
      RECT 58.465 4.13 58.615 4.28 ;
      RECT 57.285 3.41 57.435 3.56 ;
      RECT 56.63 4.555 56.78 4.705 ;
      RECT 55.375 3.465 55.525 3.615 ;
      RECT 55.36 4.47 55.51 4.62 ;
      RECT 54.845 3.955 54.995 4.105 ;
      RECT 54.265 4.735 54.415 4.885 ;
      RECT 53.21 9.195 53.36 9.345 ;
      RECT 53.13 7.46 53.28 7.61 ;
      RECT 50.82 9.175 50.97 9.325 ;
      RECT 50.805 3.36 50.955 3.51 ;
      RECT 50.015 3.745 50.165 3.895 ;
      RECT 50.015 8.76 50.165 8.91 ;
      RECT 48.41 2.545 48.56 2.695 ;
      RECT 48.41 4.825 48.56 4.975 ;
      RECT 46.725 3.51 46.875 3.66 ;
      RECT 46.255 9.15 46.405 9.3 ;
      RECT 45.775 5.015 45.925 5.165 ;
      RECT 45.58 9.6 45.73 9.75 ;
      RECT 45.325 3.515 45.475 3.665 ;
      RECT 45.145 4.505 45.295 4.655 ;
      RECT 44.75 5.02 44.9 5.17 ;
      RECT 44.39 4.975 44.54 5.125 ;
      RECT 44.245 3.465 44.395 3.615 ;
      RECT 43.66 4.915 43.81 5.065 ;
      RECT 43.565 3.45 43.715 3.6 ;
      RECT 43.41 3.985 43.56 4.135 ;
      RECT 42.725 4.95 42.875 5.1 ;
      RECT 42.33 3.575 42.48 3.725 ;
      RECT 41.61 4.48 41.76 4.63 ;
      RECT 41.57 3.515 41.72 3.665 ;
      RECT 41.3 4.985 41.45 5.135 ;
      RECT 40.765 3.705 40.915 3.855 ;
      RECT 40.72 4.575 40.87 4.725 ;
      RECT 40.54 4.13 40.69 4.28 ;
      RECT 39.36 3.41 39.51 3.56 ;
      RECT 38.705 4.555 38.855 4.705 ;
      RECT 37.45 3.465 37.6 3.615 ;
      RECT 37.435 4.47 37.585 4.62 ;
      RECT 36.92 3.955 37.07 4.105 ;
      RECT 36.34 4.735 36.49 4.885 ;
      RECT 35.285 9.195 35.435 9.345 ;
      RECT 35.205 7.46 35.355 7.61 ;
      RECT 32.895 9.175 33.045 9.325 ;
      RECT 32.88 3.36 33.03 3.51 ;
      RECT 32.09 3.745 32.24 3.895 ;
      RECT 32.09 8.76 32.24 8.91 ;
      RECT 30.485 2.545 30.635 2.695 ;
      RECT 30.485 4.825 30.635 4.975 ;
      RECT 28.8 3.51 28.95 3.66 ;
      RECT 28.3 9.14 28.45 9.29 ;
      RECT 27.85 5.015 28 5.165 ;
      RECT 27.655 9.6 27.805 9.75 ;
      RECT 27.4 3.515 27.55 3.665 ;
      RECT 27.22 4.505 27.37 4.655 ;
      RECT 26.825 5.02 26.975 5.17 ;
      RECT 26.465 4.975 26.615 5.125 ;
      RECT 26.32 3.465 26.47 3.615 ;
      RECT 25.735 4.915 25.885 5.065 ;
      RECT 25.64 3.45 25.79 3.6 ;
      RECT 25.485 3.985 25.635 4.135 ;
      RECT 24.8 4.95 24.95 5.1 ;
      RECT 24.405 3.575 24.555 3.725 ;
      RECT 23.685 4.48 23.835 4.63 ;
      RECT 23.645 3.515 23.795 3.665 ;
      RECT 23.375 4.985 23.525 5.135 ;
      RECT 22.84 3.705 22.99 3.855 ;
      RECT 22.795 4.575 22.945 4.725 ;
      RECT 22.615 4.13 22.765 4.28 ;
      RECT 21.435 3.41 21.585 3.56 ;
      RECT 20.78 4.555 20.93 4.705 ;
      RECT 19.525 3.465 19.675 3.615 ;
      RECT 19.51 4.47 19.66 4.62 ;
      RECT 18.995 3.955 19.145 4.105 ;
      RECT 18.415 4.735 18.565 4.885 ;
      RECT 16.63 9.53 16.78 9.68 ;
      RECT 16.255 8.79 16.405 8.94 ;
    LAYER met1 ;
      RECT 106.83 10.205 107.125 10.435 ;
      RECT 106.89 9.71 107.065 10.435 ;
      RECT 106.86 9.71 107.21 10.06 ;
      RECT 106.89 8.725 107.06 10.435 ;
      RECT 106.83 8.725 107.12 8.955 ;
      RECT 105.84 10.205 106.135 10.435 ;
      RECT 105.9 8.725 106.07 10.435 ;
      RECT 105.84 8.725 106.13 8.955 ;
      RECT 105.84 8.76 106.69 8.92 ;
      RECT 106.525 8.355 106.69 8.92 ;
      RECT 105.84 8.755 106.235 8.92 ;
      RECT 106.46 8.355 106.75 8.585 ;
      RECT 106.46 8.385 106.92 8.555 ;
      RECT 106.425 4.025 106.745 4.26 ;
      RECT 106.425 4.055 106.915 4.225 ;
      RECT 106.425 3.69 106.615 4.26 ;
      RECT 105.84 3.655 106.13 3.885 ;
      RECT 105.84 3.69 106.615 3.86 ;
      RECT 105.9 2.175 106.07 3.885 ;
      RECT 105.84 2.175 106.135 2.405 ;
      RECT 105.47 4.025 105.76 4.255 ;
      RECT 105.47 4.055 105.93 4.225 ;
      RECT 105.535 2.95 105.7 4.255 ;
      RECT 104.05 2.915 104.34 3.145 ;
      RECT 104.05 2.95 105.7 3.12 ;
      RECT 104.11 2.175 104.28 3.145 ;
      RECT 104.05 2.175 104.34 2.405 ;
      RECT 104.05 10.205 104.34 10.435 ;
      RECT 104.11 9.465 104.28 10.435 ;
      RECT 104.11 9.555 105.7 9.725 ;
      RECT 105.53 8.355 105.7 9.725 ;
      RECT 104.05 9.465 104.34 9.695 ;
      RECT 105.47 8.355 105.76 8.585 ;
      RECT 105.47 8.385 105.93 8.555 ;
      RECT 102.085 4.725 102.435 5.075 ;
      RECT 102.175 3.32 102.345 5.075 ;
      RECT 104.48 3.26 104.83 3.61 ;
      RECT 102.175 3.32 103.795 3.495 ;
      RECT 102.175 3.32 104.45 3.49 ;
      RECT 104.31 3.315 104.83 3.485 ;
      RECT 104.505 9.09 104.83 9.415 ;
      RECT 100.16 9.05 100.51 9.4 ;
      RECT 104.48 9.095 104.83 9.325 ;
      RECT 99.72 9.095 100.01 9.325 ;
      RECT 104.31 9.12 104.83 9.295 ;
      RECT 99.55 9.125 100.01 9.295 ;
      RECT 99.72 9.12 104.83 9.29 ;
      RECT 103.705 3.66 104.025 3.98 ;
      RECT 103.68 3.655 103.97 3.885 ;
      RECT 103.635 3.685 104.025 3.86 ;
      RECT 103.505 3.685 104.025 3.855 ;
      RECT 103.705 8.66 104.025 8.98 ;
      RECT 103.68 8.725 104.025 8.955 ;
      RECT 103.505 8.755 104.025 8.925 ;
      RECT 99.495 4.96 99.535 5.22 ;
      RECT 99.535 4.94 99.54 4.95 ;
      RECT 100.865 4.185 100.875 4.406 ;
      RECT 100.795 4.18 100.865 4.531 ;
      RECT 100.785 4.18 100.795 4.658 ;
      RECT 100.76 4.18 100.785 4.705 ;
      RECT 100.735 4.18 100.76 4.783 ;
      RECT 100.715 4.18 100.735 4.853 ;
      RECT 100.69 4.18 100.715 4.893 ;
      RECT 100.68 4.18 100.69 4.913 ;
      RECT 100.67 4.182 100.68 4.921 ;
      RECT 100.665 4.187 100.67 4.378 ;
      RECT 100.665 4.387 100.67 4.922 ;
      RECT 100.66 4.432 100.665 4.923 ;
      RECT 100.65 4.497 100.66 4.924 ;
      RECT 100.64 4.592 100.65 4.926 ;
      RECT 100.635 4.645 100.64 4.928 ;
      RECT 100.63 4.665 100.635 4.929 ;
      RECT 100.575 4.69 100.63 4.935 ;
      RECT 100.535 4.725 100.575 4.944 ;
      RECT 100.525 4.742 100.535 4.949 ;
      RECT 100.516 4.748 100.525 4.951 ;
      RECT 100.43 4.786 100.516 4.962 ;
      RECT 100.425 4.825 100.43 4.972 ;
      RECT 100.35 4.832 100.425 4.982 ;
      RECT 100.33 4.842 100.35 4.993 ;
      RECT 100.3 4.849 100.33 5.001 ;
      RECT 100.275 4.856 100.3 5.008 ;
      RECT 100.251 4.862 100.275 5.013 ;
      RECT 100.165 4.875 100.251 5.025 ;
      RECT 100.087 4.882 100.165 5.043 ;
      RECT 100.001 4.877 100.087 5.061 ;
      RECT 99.915 4.872 100.001 5.081 ;
      RECT 99.835 4.866 99.915 5.098 ;
      RECT 99.77 4.862 99.835 5.127 ;
      RECT 99.765 4.576 99.77 4.6 ;
      RECT 99.755 4.852 99.77 5.155 ;
      RECT 99.76 4.57 99.765 4.64 ;
      RECT 99.755 4.564 99.76 4.71 ;
      RECT 99.75 4.558 99.755 4.788 ;
      RECT 99.75 4.835 99.755 5.22 ;
      RECT 99.742 4.555 99.75 5.22 ;
      RECT 99.656 4.553 99.742 5.22 ;
      RECT 99.57 4.551 99.656 5.22 ;
      RECT 99.56 4.552 99.57 5.22 ;
      RECT 99.555 4.557 99.56 5.22 ;
      RECT 99.545 4.57 99.555 5.22 ;
      RECT 99.54 4.592 99.545 5.22 ;
      RECT 99.535 4.952 99.54 5.22 ;
      RECT 100.165 4.42 100.17 4.64 ;
      RECT 100.67 3.455 100.705 3.715 ;
      RECT 100.655 3.455 100.67 3.723 ;
      RECT 100.626 3.455 100.655 3.745 ;
      RECT 100.54 3.455 100.626 3.805 ;
      RECT 100.52 3.455 100.54 3.87 ;
      RECT 100.46 3.455 100.52 4.035 ;
      RECT 100.455 3.455 100.46 4.183 ;
      RECT 100.45 3.455 100.455 4.195 ;
      RECT 100.445 3.455 100.45 4.221 ;
      RECT 100.415 3.641 100.445 4.301 ;
      RECT 100.41 3.689 100.415 4.39 ;
      RECT 100.405 3.703 100.41 4.405 ;
      RECT 100.4 3.722 100.405 4.435 ;
      RECT 100.395 3.737 100.4 4.451 ;
      RECT 100.39 3.752 100.395 4.473 ;
      RECT 100.385 3.772 100.39 4.495 ;
      RECT 100.375 3.792 100.385 4.528 ;
      RECT 100.36 3.834 100.375 4.59 ;
      RECT 100.355 3.865 100.36 4.63 ;
      RECT 100.35 3.877 100.355 4.635 ;
      RECT 100.345 3.889 100.35 4.64 ;
      RECT 100.34 3.902 100.345 4.64 ;
      RECT 100.335 3.92 100.34 4.64 ;
      RECT 100.33 3.94 100.335 4.64 ;
      RECT 100.325 3.952 100.33 4.64 ;
      RECT 100.32 3.965 100.325 4.64 ;
      RECT 100.3 4 100.32 4.64 ;
      RECT 100.25 4.102 100.3 4.64 ;
      RECT 100.245 4.187 100.25 4.64 ;
      RECT 100.24 4.195 100.245 4.64 ;
      RECT 100.235 4.212 100.24 4.64 ;
      RECT 100.23 4.227 100.235 4.64 ;
      RECT 100.195 4.292 100.23 4.64 ;
      RECT 100.18 4.357 100.195 4.64 ;
      RECT 100.175 4.387 100.18 4.64 ;
      RECT 100.17 4.412 100.175 4.64 ;
      RECT 100.155 4.422 100.165 4.64 ;
      RECT 100.14 4.435 100.155 4.633 ;
      RECT 99.885 4.025 99.955 4.235 ;
      RECT 99.675 4.002 99.68 4.195 ;
      RECT 97.13 3.93 97.39 4.19 ;
      RECT 99.965 4.212 99.97 4.215 ;
      RECT 99.955 4.03 99.965 4.23 ;
      RECT 99.856 4.023 99.885 4.235 ;
      RECT 99.77 4.015 99.856 4.235 ;
      RECT 99.755 4.009 99.77 4.233 ;
      RECT 99.735 4.008 99.755 4.22 ;
      RECT 99.73 4.007 99.735 4.203 ;
      RECT 99.68 4.004 99.73 4.198 ;
      RECT 99.65 4.001 99.675 4.193 ;
      RECT 99.63 3.999 99.65 4.188 ;
      RECT 99.615 3.997 99.63 4.185 ;
      RECT 99.585 3.995 99.615 4.183 ;
      RECT 99.52 3.991 99.585 4.175 ;
      RECT 99.49 3.986 99.52 4.17 ;
      RECT 99.47 3.984 99.49 4.168 ;
      RECT 99.44 3.981 99.47 4.163 ;
      RECT 99.38 3.977 99.44 4.155 ;
      RECT 99.375 3.974 99.38 4.15 ;
      RECT 99.305 3.972 99.375 4.145 ;
      RECT 99.276 3.968 99.305 4.138 ;
      RECT 99.19 3.963 99.276 4.13 ;
      RECT 99.156 3.958 99.19 4.122 ;
      RECT 99.07 3.95 99.156 4.114 ;
      RECT 99.031 3.943 99.07 4.106 ;
      RECT 98.945 3.938 99.031 4.098 ;
      RECT 98.88 3.932 98.945 4.088 ;
      RECT 98.86 3.927 98.88 4.083 ;
      RECT 98.851 3.924 98.86 4.082 ;
      RECT 98.765 3.92 98.851 4.076 ;
      RECT 98.725 3.916 98.765 4.068 ;
      RECT 98.705 3.912 98.725 4.066 ;
      RECT 98.645 3.912 98.705 4.063 ;
      RECT 98.625 3.915 98.645 4.061 ;
      RECT 98.604 3.915 98.625 4.061 ;
      RECT 98.518 3.917 98.604 4.065 ;
      RECT 98.432 3.919 98.518 4.071 ;
      RECT 98.346 3.921 98.432 4.078 ;
      RECT 98.26 3.924 98.346 4.084 ;
      RECT 98.226 3.925 98.26 4.089 ;
      RECT 98.14 3.928 98.226 4.094 ;
      RECT 98.111 3.935 98.14 4.099 ;
      RECT 98.025 3.935 98.111 4.104 ;
      RECT 97.992 3.935 98.025 4.109 ;
      RECT 97.906 3.937 97.992 4.114 ;
      RECT 97.82 3.939 97.906 4.121 ;
      RECT 97.756 3.941 97.82 4.127 ;
      RECT 97.67 3.943 97.756 4.133 ;
      RECT 97.667 3.945 97.67 4.136 ;
      RECT 97.581 3.946 97.667 4.14 ;
      RECT 97.495 3.949 97.581 4.147 ;
      RECT 97.476 3.951 97.495 4.151 ;
      RECT 97.39 3.953 97.476 4.156 ;
      RECT 97.12 3.965 97.13 4.16 ;
      RECT 99.29 10.205 99.58 10.435 ;
      RECT 99.35 9.465 99.52 10.435 ;
      RECT 99.24 9.49 99.615 9.86 ;
      RECT 99.29 9.465 99.58 9.86 ;
      RECT 99.355 3.545 99.54 3.755 ;
      RECT 99.35 3.546 99.545 3.753 ;
      RECT 99.345 3.551 99.555 3.748 ;
      RECT 99.34 3.527 99.345 3.745 ;
      RECT 99.31 3.524 99.34 3.738 ;
      RECT 99.305 3.52 99.31 3.729 ;
      RECT 99.27 3.551 99.555 3.724 ;
      RECT 99.045 3.46 99.305 3.72 ;
      RECT 99.345 3.529 99.35 3.748 ;
      RECT 99.35 3.53 99.355 3.753 ;
      RECT 99.045 3.542 99.425 3.72 ;
      RECT 99.045 3.54 99.41 3.72 ;
      RECT 99.045 3.535 99.4 3.72 ;
      RECT 99 4.45 99.05 4.735 ;
      RECT 98.945 4.42 98.95 4.735 ;
      RECT 98.915 4.4 98.92 4.735 ;
      RECT 99.065 4.45 99.125 4.71 ;
      RECT 99.06 4.45 99.065 4.718 ;
      RECT 99.05 4.45 99.06 4.73 ;
      RECT 98.965 4.44 99 4.735 ;
      RECT 98.96 4.427 98.965 4.735 ;
      RECT 98.95 4.422 98.96 4.735 ;
      RECT 98.93 4.412 98.945 4.735 ;
      RECT 98.92 4.405 98.93 4.735 ;
      RECT 98.91 4.397 98.915 4.735 ;
      RECT 98.88 4.387 98.91 4.735 ;
      RECT 98.865 4.375 98.88 4.735 ;
      RECT 98.85 4.365 98.865 4.73 ;
      RECT 98.83 4.355 98.85 4.705 ;
      RECT 98.82 4.347 98.83 4.682 ;
      RECT 98.79 4.33 98.82 4.672 ;
      RECT 98.785 4.307 98.79 4.663 ;
      RECT 98.78 4.294 98.785 4.661 ;
      RECT 98.765 4.27 98.78 4.655 ;
      RECT 98.76 4.246 98.765 4.649 ;
      RECT 98.75 4.235 98.76 4.644 ;
      RECT 98.745 4.225 98.75 4.64 ;
      RECT 98.74 4.217 98.745 4.637 ;
      RECT 98.73 4.212 98.74 4.633 ;
      RECT 98.725 4.207 98.73 4.629 ;
      RECT 98.64 4.205 98.725 4.604 ;
      RECT 98.61 4.205 98.64 4.57 ;
      RECT 98.595 4.205 98.61 4.553 ;
      RECT 98.54 4.205 98.595 4.498 ;
      RECT 98.535 4.21 98.54 4.447 ;
      RECT 98.525 4.215 98.535 4.437 ;
      RECT 98.52 4.225 98.525 4.423 ;
      RECT 98.47 4.965 98.73 5.225 ;
      RECT 98.39 4.98 98.73 5.201 ;
      RECT 98.37 4.98 98.73 5.196 ;
      RECT 98.346 4.98 98.73 5.194 ;
      RECT 98.26 4.98 98.73 5.189 ;
      RECT 98.11 4.92 98.37 5.185 ;
      RECT 98.065 4.98 98.73 5.18 ;
      RECT 98.06 4.987 98.73 5.175 ;
      RECT 98.075 4.975 98.39 5.185 ;
      RECT 97.965 3.41 98.225 3.67 ;
      RECT 97.965 3.467 98.23 3.663 ;
      RECT 97.965 3.497 98.235 3.595 ;
      RECT 98.025 3.928 98.14 3.93 ;
      RECT 98.111 3.925 98.14 3.93 ;
      RECT 97.135 4.929 97.16 5.169 ;
      RECT 97.12 4.932 97.21 5.163 ;
      RECT 97.115 4.937 97.296 5.158 ;
      RECT 97.11 4.945 97.36 5.156 ;
      RECT 97.11 4.945 97.37 5.155 ;
      RECT 97.105 4.952 97.38 5.148 ;
      RECT 97.105 4.952 97.466 5.137 ;
      RECT 97.1 4.987 97.466 5.133 ;
      RECT 97.1 4.987 97.475 5.122 ;
      RECT 97.38 4.86 97.64 5.12 ;
      RECT 97.09 5.037 97.64 5.118 ;
      RECT 97.36 4.905 97.38 5.153 ;
      RECT 97.296 4.908 97.36 5.157 ;
      RECT 97.21 4.913 97.296 5.162 ;
      RECT 97.14 4.924 97.64 5.12 ;
      RECT 97.16 4.918 97.21 5.167 ;
      RECT 97.285 3.395 97.295 3.657 ;
      RECT 97.275 3.452 97.285 3.66 ;
      RECT 97.25 3.457 97.275 3.666 ;
      RECT 97.225 3.461 97.25 3.678 ;
      RECT 97.215 3.464 97.225 3.688 ;
      RECT 97.21 3.465 97.215 3.693 ;
      RECT 97.205 3.466 97.21 3.698 ;
      RECT 97.2 3.467 97.205 3.7 ;
      RECT 97.175 3.47 97.2 3.703 ;
      RECT 97.145 3.476 97.175 3.706 ;
      RECT 97.08 3.487 97.145 3.709 ;
      RECT 97.035 3.495 97.08 3.713 ;
      RECT 97.02 3.495 97.035 3.721 ;
      RECT 97.015 3.496 97.02 3.728 ;
      RECT 97.01 3.498 97.015 3.731 ;
      RECT 97.005 3.502 97.01 3.734 ;
      RECT 96.995 3.51 97.005 3.738 ;
      RECT 96.99 3.523 96.995 3.743 ;
      RECT 96.985 3.531 96.99 3.745 ;
      RECT 96.98 3.537 96.985 3.745 ;
      RECT 96.975 3.541 96.98 3.748 ;
      RECT 96.97 3.543 96.975 3.751 ;
      RECT 96.965 3.546 96.97 3.754 ;
      RECT 96.955 3.551 96.965 3.758 ;
      RECT 96.95 3.557 96.955 3.763 ;
      RECT 96.94 3.563 96.95 3.767 ;
      RECT 96.925 3.57 96.94 3.773 ;
      RECT 96.896 3.584 96.925 3.783 ;
      RECT 96.81 3.619 96.896 3.815 ;
      RECT 96.79 3.652 96.81 3.844 ;
      RECT 96.77 3.665 96.79 3.855 ;
      RECT 96.75 3.677 96.77 3.866 ;
      RECT 96.7 3.699 96.75 3.886 ;
      RECT 96.685 3.717 96.7 3.903 ;
      RECT 96.68 3.723 96.685 3.906 ;
      RECT 96.675 3.727 96.68 3.909 ;
      RECT 96.67 3.731 96.675 3.913 ;
      RECT 96.665 3.733 96.67 3.916 ;
      RECT 96.655 3.74 96.665 3.919 ;
      RECT 96.65 3.745 96.655 3.923 ;
      RECT 96.645 3.747 96.65 3.926 ;
      RECT 96.64 3.751 96.645 3.929 ;
      RECT 96.635 3.753 96.64 3.933 ;
      RECT 96.62 3.758 96.635 3.938 ;
      RECT 96.615 3.763 96.62 3.941 ;
      RECT 96.61 3.771 96.615 3.944 ;
      RECT 96.605 3.773 96.61 3.947 ;
      RECT 96.6 3.775 96.605 3.95 ;
      RECT 96.59 3.777 96.6 3.956 ;
      RECT 96.555 3.791 96.59 3.968 ;
      RECT 96.545 3.806 96.555 3.978 ;
      RECT 96.47 3.835 96.545 4.002 ;
      RECT 96.465 3.86 96.47 4.025 ;
      RECT 96.45 3.864 96.465 4.031 ;
      RECT 96.44 3.872 96.45 4.036 ;
      RECT 96.41 3.885 96.44 4.04 ;
      RECT 96.4 3.9 96.41 4.045 ;
      RECT 96.39 3.905 96.4 4.048 ;
      RECT 96.385 3.907 96.39 4.05 ;
      RECT 96.37 3.91 96.385 4.053 ;
      RECT 96.365 3.912 96.37 4.056 ;
      RECT 96.345 3.917 96.365 4.06 ;
      RECT 96.315 3.922 96.345 4.068 ;
      RECT 96.29 3.929 96.315 4.076 ;
      RECT 96.285 3.934 96.29 4.081 ;
      RECT 96.255 3.937 96.285 4.085 ;
      RECT 96.215 3.94 96.255 4.095 ;
      RECT 96.18 3.937 96.215 4.107 ;
      RECT 96.17 3.933 96.18 4.114 ;
      RECT 96.145 3.929 96.17 4.12 ;
      RECT 96.14 3.925 96.145 4.125 ;
      RECT 96.1 3.922 96.14 4.125 ;
      RECT 96.085 3.907 96.1 4.126 ;
      RECT 96.062 3.895 96.085 4.126 ;
      RECT 95.976 3.895 96.062 4.127 ;
      RECT 95.89 3.895 95.976 4.129 ;
      RECT 95.87 3.895 95.89 4.126 ;
      RECT 95.865 3.9 95.87 4.121 ;
      RECT 95.86 3.905 95.865 4.119 ;
      RECT 95.85 3.915 95.86 4.117 ;
      RECT 95.845 3.921 95.85 4.11 ;
      RECT 95.84 3.923 95.845 4.095 ;
      RECT 95.835 3.927 95.84 4.085 ;
      RECT 97.295 3.395 97.545 3.655 ;
      RECT 95.02 4.93 95.28 5.19 ;
      RECT 97.315 4.42 97.32 4.63 ;
      RECT 97.32 4.425 97.33 4.625 ;
      RECT 97.27 4.42 97.315 4.645 ;
      RECT 97.26 4.42 97.27 4.665 ;
      RECT 97.241 4.42 97.26 4.67 ;
      RECT 97.155 4.42 97.241 4.667 ;
      RECT 97.125 4.422 97.155 4.665 ;
      RECT 97.07 4.432 97.125 4.663 ;
      RECT 97.005 4.446 97.07 4.661 ;
      RECT 97 4.454 97.005 4.66 ;
      RECT 96.985 4.457 97 4.658 ;
      RECT 96.92 4.467 96.985 4.654 ;
      RECT 96.872 4.481 96.92 4.655 ;
      RECT 96.786 4.498 96.872 4.669 ;
      RECT 96.7 4.519 96.786 4.686 ;
      RECT 96.68 4.532 96.7 4.696 ;
      RECT 96.635 4.54 96.68 4.703 ;
      RECT 96.6 4.548 96.635 4.711 ;
      RECT 96.566 4.556 96.6 4.719 ;
      RECT 96.48 4.57 96.566 4.731 ;
      RECT 96.445 4.587 96.48 4.743 ;
      RECT 96.436 4.596 96.445 4.747 ;
      RECT 96.35 4.614 96.436 4.764 ;
      RECT 96.291 4.641 96.35 4.791 ;
      RECT 96.205 4.668 96.291 4.819 ;
      RECT 96.185 4.69 96.205 4.839 ;
      RECT 96.125 4.705 96.185 4.855 ;
      RECT 96.115 4.717 96.125 4.868 ;
      RECT 96.11 4.722 96.115 4.871 ;
      RECT 96.1 4.725 96.11 4.874 ;
      RECT 96.095 4.727 96.1 4.877 ;
      RECT 96.065 4.735 96.095 4.884 ;
      RECT 96.05 4.742 96.065 4.892 ;
      RECT 96.04 4.747 96.05 4.896 ;
      RECT 96.035 4.75 96.04 4.899 ;
      RECT 96.025 4.752 96.035 4.902 ;
      RECT 95.99 4.762 96.025 4.911 ;
      RECT 95.915 4.785 95.99 4.933 ;
      RECT 95.895 4.803 95.915 4.951 ;
      RECT 95.865 4.81 95.895 4.961 ;
      RECT 95.845 4.818 95.865 4.971 ;
      RECT 95.835 4.824 95.845 4.978 ;
      RECT 95.816 4.829 95.835 4.984 ;
      RECT 95.73 4.849 95.816 5.004 ;
      RECT 95.715 4.869 95.73 5.023 ;
      RECT 95.67 4.881 95.715 5.034 ;
      RECT 95.605 4.902 95.67 5.057 ;
      RECT 95.565 4.922 95.605 5.078 ;
      RECT 95.555 4.932 95.565 5.088 ;
      RECT 95.505 4.944 95.555 5.099 ;
      RECT 95.485 4.96 95.505 5.111 ;
      RECT 95.455 4.97 95.485 5.117 ;
      RECT 95.445 4.975 95.455 5.119 ;
      RECT 95.376 4.976 95.445 5.125 ;
      RECT 95.29 4.978 95.376 5.135 ;
      RECT 95.28 4.979 95.29 5.14 ;
      RECT 96.55 5.005 96.74 5.215 ;
      RECT 96.54 5.01 96.75 5.208 ;
      RECT 96.525 5.01 96.75 5.173 ;
      RECT 96.445 4.895 96.705 5.155 ;
      RECT 95.36 4.425 95.545 4.72 ;
      RECT 95.35 4.425 95.545 4.718 ;
      RECT 95.335 4.425 95.55 4.713 ;
      RECT 95.335 4.425 95.555 4.71 ;
      RECT 95.33 4.425 95.555 4.708 ;
      RECT 95.325 4.68 95.555 4.698 ;
      RECT 95.33 4.425 95.59 4.685 ;
      RECT 95.29 3.46 95.55 3.72 ;
      RECT 95.1 3.385 95.186 3.718 ;
      RECT 95.075 3.389 95.23 3.714 ;
      RECT 95.186 3.381 95.23 3.714 ;
      RECT 95.186 3.382 95.235 3.713 ;
      RECT 95.1 3.387 95.25 3.712 ;
      RECT 95.075 3.395 95.29 3.711 ;
      RECT 95.07 3.39 95.25 3.706 ;
      RECT 95.06 3.405 95.29 3.613 ;
      RECT 95.06 3.457 95.49 3.613 ;
      RECT 95.06 3.45 95.47 3.613 ;
      RECT 95.06 3.437 95.44 3.613 ;
      RECT 95.06 3.425 95.38 3.613 ;
      RECT 95.06 3.41 95.355 3.613 ;
      RECT 94.26 4.04 94.395 4.335 ;
      RECT 94.52 4.063 94.525 4.25 ;
      RECT 95.24 3.96 95.385 4.195 ;
      RECT 95.4 3.96 95.405 4.185 ;
      RECT 95.435 3.971 95.44 4.165 ;
      RECT 95.43 3.963 95.435 4.17 ;
      RECT 95.41 3.96 95.43 4.175 ;
      RECT 95.405 3.96 95.41 4.183 ;
      RECT 95.395 3.96 95.4 4.188 ;
      RECT 95.385 3.96 95.395 4.193 ;
      RECT 95.215 3.962 95.24 4.195 ;
      RECT 95.165 3.969 95.215 4.195 ;
      RECT 95.16 3.974 95.165 4.195 ;
      RECT 95.121 3.979 95.16 4.196 ;
      RECT 95.035 3.991 95.121 4.197 ;
      RECT 95.026 4.001 95.035 4.197 ;
      RECT 94.94 4.01 95.026 4.199 ;
      RECT 94.916 4.02 94.94 4.201 ;
      RECT 94.83 4.031 94.916 4.202 ;
      RECT 94.8 4.042 94.83 4.204 ;
      RECT 94.77 4.047 94.8 4.206 ;
      RECT 94.745 4.053 94.77 4.209 ;
      RECT 94.73 4.058 94.745 4.21 ;
      RECT 94.685 4.064 94.73 4.21 ;
      RECT 94.68 4.069 94.685 4.211 ;
      RECT 94.66 4.069 94.68 4.213 ;
      RECT 94.64 4.067 94.66 4.218 ;
      RECT 94.605 4.066 94.64 4.225 ;
      RECT 94.575 4.065 94.605 4.235 ;
      RECT 94.525 4.064 94.575 4.245 ;
      RECT 94.435 4.061 94.52 4.335 ;
      RECT 94.41 4.055 94.435 4.335 ;
      RECT 94.395 4.045 94.41 4.335 ;
      RECT 94.21 4.04 94.26 4.255 ;
      RECT 94.2 4.045 94.21 4.245 ;
      RECT 94.44 4.52 94.7 4.78 ;
      RECT 94.44 4.52 94.73 4.673 ;
      RECT 94.44 4.52 94.765 4.658 ;
      RECT 94.695 4.44 94.885 4.65 ;
      RECT 94.685 4.445 94.895 4.643 ;
      RECT 94.65 4.515 94.895 4.643 ;
      RECT 94.68 4.457 94.7 4.78 ;
      RECT 94.665 4.505 94.895 4.643 ;
      RECT 94.67 4.477 94.7 4.78 ;
      RECT 93.75 3.545 93.82 4.65 ;
      RECT 94.485 3.65 94.745 3.91 ;
      RECT 94.065 3.696 94.08 3.905 ;
      RECT 94.401 3.709 94.485 3.86 ;
      RECT 94.315 3.706 94.401 3.86 ;
      RECT 94.276 3.704 94.315 3.86 ;
      RECT 94.19 3.702 94.276 3.86 ;
      RECT 94.13 3.7 94.19 3.871 ;
      RECT 94.095 3.698 94.13 3.889 ;
      RECT 94.08 3.696 94.095 3.9 ;
      RECT 94.05 3.696 94.065 3.913 ;
      RECT 94.04 3.696 94.05 3.918 ;
      RECT 94.015 3.695 94.04 3.923 ;
      RECT 94 3.69 94.015 3.929 ;
      RECT 93.995 3.683 94 3.934 ;
      RECT 93.97 3.674 93.995 3.94 ;
      RECT 93.925 3.653 93.97 3.953 ;
      RECT 93.915 3.637 93.925 3.963 ;
      RECT 93.9 3.63 93.915 3.973 ;
      RECT 93.89 3.623 93.9 3.99 ;
      RECT 93.885 3.62 93.89 4.02 ;
      RECT 93.88 3.618 93.885 4.05 ;
      RECT 93.875 3.616 93.88 4.087 ;
      RECT 93.86 3.612 93.875 4.154 ;
      RECT 93.86 4.445 93.87 4.645 ;
      RECT 93.855 3.608 93.86 4.28 ;
      RECT 93.855 4.432 93.86 4.65 ;
      RECT 93.85 3.606 93.855 4.365 ;
      RECT 93.85 4.422 93.855 4.65 ;
      RECT 93.835 3.577 93.85 4.65 ;
      RECT 93.82 3.55 93.835 4.65 ;
      RECT 93.745 3.545 93.75 3.9 ;
      RECT 93.745 3.955 93.75 4.65 ;
      RECT 93.73 3.545 93.745 3.878 ;
      RECT 93.74 3.977 93.745 4.65 ;
      RECT 93.73 4.017 93.74 4.65 ;
      RECT 93.695 3.545 93.73 3.82 ;
      RECT 93.725 4.052 93.73 4.65 ;
      RECT 93.71 4.107 93.725 4.65 ;
      RECT 93.705 4.172 93.71 4.65 ;
      RECT 93.69 4.22 93.705 4.65 ;
      RECT 93.665 3.545 93.695 3.775 ;
      RECT 93.685 4.275 93.69 4.65 ;
      RECT 93.67 4.335 93.685 4.65 ;
      RECT 93.665 4.383 93.67 4.648 ;
      RECT 93.66 3.545 93.665 3.768 ;
      RECT 93.66 4.415 93.665 4.643 ;
      RECT 93.635 3.545 93.66 3.76 ;
      RECT 93.625 3.55 93.635 3.75 ;
      RECT 93.84 4.825 93.86 5.065 ;
      RECT 93.07 4.755 93.075 4.965 ;
      RECT 94.35 4.828 94.36 5.023 ;
      RECT 94.345 4.818 94.35 5.026 ;
      RECT 94.265 4.815 94.345 5.049 ;
      RECT 94.261 4.815 94.265 5.071 ;
      RECT 94.175 4.815 94.261 5.081 ;
      RECT 94.16 4.815 94.175 5.089 ;
      RECT 94.131 4.816 94.16 5.087 ;
      RECT 94.045 4.821 94.131 5.083 ;
      RECT 94.032 4.825 94.045 5.079 ;
      RECT 93.946 4.825 94.032 5.075 ;
      RECT 93.86 4.825 93.946 5.069 ;
      RECT 93.776 4.825 93.84 5.063 ;
      RECT 93.69 4.825 93.776 5.058 ;
      RECT 93.67 4.825 93.69 5.054 ;
      RECT 93.61 4.82 93.67 5.051 ;
      RECT 93.582 4.814 93.61 5.048 ;
      RECT 93.496 4.809 93.582 5.044 ;
      RECT 93.41 4.803 93.496 5.038 ;
      RECT 93.335 4.785 93.41 5.033 ;
      RECT 93.3 4.762 93.335 5.029 ;
      RECT 93.29 4.752 93.3 5.028 ;
      RECT 93.235 4.75 93.29 5.027 ;
      RECT 93.16 4.75 93.235 5.023 ;
      RECT 93.15 4.75 93.16 5.018 ;
      RECT 93.135 4.75 93.15 5.01 ;
      RECT 93.085 4.752 93.135 4.988 ;
      RECT 93.075 4.755 93.085 4.968 ;
      RECT 93.065 4.76 93.07 4.963 ;
      RECT 93.06 4.765 93.065 4.958 ;
      RECT 91.17 3.41 91.43 3.67 ;
      RECT 91.16 3.44 91.43 3.65 ;
      RECT 93.08 3.355 93.34 3.615 ;
      RECT 93.075 3.43 93.08 3.616 ;
      RECT 93.05 3.435 93.075 3.618 ;
      RECT 93.035 3.442 93.05 3.621 ;
      RECT 92.975 3.46 93.035 3.626 ;
      RECT 92.945 3.48 92.975 3.633 ;
      RECT 92.92 3.488 92.945 3.638 ;
      RECT 92.895 3.496 92.92 3.64 ;
      RECT 92.877 3.5 92.895 3.639 ;
      RECT 92.791 3.498 92.877 3.639 ;
      RECT 92.705 3.496 92.791 3.639 ;
      RECT 92.619 3.494 92.705 3.638 ;
      RECT 92.533 3.492 92.619 3.638 ;
      RECT 92.447 3.49 92.533 3.638 ;
      RECT 92.361 3.488 92.447 3.638 ;
      RECT 92.275 3.486 92.361 3.637 ;
      RECT 92.257 3.485 92.275 3.637 ;
      RECT 92.171 3.484 92.257 3.637 ;
      RECT 92.085 3.482 92.171 3.637 ;
      RECT 91.999 3.481 92.085 3.636 ;
      RECT 91.913 3.48 91.999 3.636 ;
      RECT 91.827 3.478 91.913 3.636 ;
      RECT 91.741 3.477 91.827 3.636 ;
      RECT 91.655 3.475 91.741 3.635 ;
      RECT 91.631 3.473 91.655 3.635 ;
      RECT 91.545 3.466 91.631 3.635 ;
      RECT 91.516 3.458 91.545 3.635 ;
      RECT 91.43 3.45 91.516 3.635 ;
      RECT 91.15 3.447 91.16 3.645 ;
      RECT 92.655 4.41 92.66 4.76 ;
      RECT 92.425 4.5 92.565 4.76 ;
      RECT 92.9 4.185 92.945 4.395 ;
      RECT 92.955 4.196 92.965 4.39 ;
      RECT 92.945 4.188 92.955 4.395 ;
      RECT 92.88 4.185 92.9 4.4 ;
      RECT 92.85 4.185 92.88 4.423 ;
      RECT 92.84 4.185 92.85 4.448 ;
      RECT 92.835 4.185 92.84 4.458 ;
      RECT 92.78 4.185 92.835 4.498 ;
      RECT 92.775 4.185 92.78 4.538 ;
      RECT 92.77 4.187 92.775 4.543 ;
      RECT 92.755 4.197 92.77 4.554 ;
      RECT 92.71 4.255 92.755 4.59 ;
      RECT 92.7 4.31 92.71 4.624 ;
      RECT 92.685 4.337 92.7 4.64 ;
      RECT 92.675 4.364 92.685 4.76 ;
      RECT 92.66 4.387 92.675 4.76 ;
      RECT 92.65 4.427 92.655 4.76 ;
      RECT 92.645 4.437 92.65 4.76 ;
      RECT 92.64 4.452 92.645 4.76 ;
      RECT 92.63 4.457 92.64 4.76 ;
      RECT 92.565 4.48 92.63 4.76 ;
      RECT 92.035 3.975 92.255 4.185 ;
      RECT 92.035 3.982 92.265 4.18 ;
      RECT 91.34 3.99 92.265 4.165 ;
      RECT 91.86 3.885 92.25 4.165 ;
      RECT 90.64 3.9 90.9 4.16 ;
      RECT 91.275 3.935 91.41 4.12 ;
      RECT 91.2 3.925 91.295 4.115 ;
      RECT 91.19 3.99 92.265 4.111 ;
      RECT 90.94 3.99 92.265 4.11 ;
      RECT 90.965 3.91 91.205 4.11 ;
      RECT 90.64 3.915 91.225 4.098 ;
      RECT 92.555 3.94 92.595 4.025 ;
      RECT 90.64 3.975 91.815 4.098 ;
      RECT 90.64 3.965 91.7 4.098 ;
      RECT 90.64 3.946 91.605 4.098 ;
      RECT 91.425 3.94 91.605 4.165 ;
      RECT 91.86 3.92 92.555 3.955 ;
      RECT 90.96 3.912 91.205 4.11 ;
      RECT 90.975 3.902 91.185 4.11 ;
      RECT 90.99 3.895 91.185 4.11 ;
      RECT 91.155 4.415 91.415 4.675 ;
      RECT 91.155 4.455 91.52 4.665 ;
      RECT 91.155 4.457 91.525 4.664 ;
      RECT 91.155 4.465 91.53 4.661 ;
      RECT 90.08 3.54 90.18 5.065 ;
      RECT 90.27 4.68 90.32 4.94 ;
      RECT 90.265 3.553 90.27 3.74 ;
      RECT 90.26 4.661 90.27 4.94 ;
      RECT 90.26 3.55 90.265 3.748 ;
      RECT 90.245 3.544 90.26 3.755 ;
      RECT 90.255 4.649 90.26 5.023 ;
      RECT 90.245 4.637 90.255 5.06 ;
      RECT 90.235 3.54 90.245 3.762 ;
      RECT 90.235 4.622 90.245 5.065 ;
      RECT 90.23 3.54 90.235 3.77 ;
      RECT 90.21 4.592 90.235 5.065 ;
      RECT 90.19 3.54 90.23 3.818 ;
      RECT 90.2 4.552 90.21 5.065 ;
      RECT 90.19 4.507 90.2 5.065 ;
      RECT 90.185 3.54 90.19 3.888 ;
      RECT 90.185 4.465 90.19 5.065 ;
      RECT 90.18 3.54 90.185 4.365 ;
      RECT 90.18 4.447 90.185 5.065 ;
      RECT 90.07 3.543 90.08 5.065 ;
      RECT 90.055 3.55 90.07 5.061 ;
      RECT 90.05 3.56 90.055 5.056 ;
      RECT 90.045 3.76 90.05 4.948 ;
      RECT 90.04 3.845 90.045 4.5 ;
      RECT 88.905 10.205 89.2 10.435 ;
      RECT 88.965 8.725 89.135 10.435 ;
      RECT 88.915 9.095 89.265 9.445 ;
      RECT 88.905 8.725 89.195 8.955 ;
      RECT 87.915 10.205 88.21 10.435 ;
      RECT 87.975 8.725 88.145 10.435 ;
      RECT 87.915 8.725 88.205 8.955 ;
      RECT 87.915 8.76 88.765 8.92 ;
      RECT 88.6 8.355 88.765 8.92 ;
      RECT 87.915 8.755 88.31 8.92 ;
      RECT 88.535 8.355 88.825 8.585 ;
      RECT 88.535 8.385 88.995 8.555 ;
      RECT 88.5 4.025 88.82 4.26 ;
      RECT 88.5 4.055 88.99 4.225 ;
      RECT 88.5 3.69 88.69 4.26 ;
      RECT 87.915 3.655 88.205 3.885 ;
      RECT 87.915 3.69 88.69 3.86 ;
      RECT 87.975 2.175 88.145 3.885 ;
      RECT 87.915 2.175 88.21 2.405 ;
      RECT 87.545 4.025 87.835 4.255 ;
      RECT 87.545 4.055 88.005 4.225 ;
      RECT 87.61 2.95 87.775 4.255 ;
      RECT 86.125 2.915 86.415 3.145 ;
      RECT 86.125 2.95 87.775 3.12 ;
      RECT 86.185 2.175 86.355 3.145 ;
      RECT 86.125 2.175 86.415 2.405 ;
      RECT 86.125 10.205 86.415 10.435 ;
      RECT 86.185 9.465 86.355 10.435 ;
      RECT 86.185 9.555 87.775 9.725 ;
      RECT 87.605 8.355 87.775 9.725 ;
      RECT 86.125 9.465 86.415 9.695 ;
      RECT 87.545 8.355 87.835 8.585 ;
      RECT 87.545 8.385 88.005 8.555 ;
      RECT 84.16 4.725 84.51 5.075 ;
      RECT 84.25 3.32 84.42 5.075 ;
      RECT 86.555 3.26 86.905 3.61 ;
      RECT 84.25 3.32 85.87 3.495 ;
      RECT 84.25 3.32 86.525 3.49 ;
      RECT 86.385 3.315 86.905 3.485 ;
      RECT 86.58 9.09 86.905 9.415 ;
      RECT 81.955 9.05 82.305 9.4 ;
      RECT 86.555 9.095 86.905 9.325 ;
      RECT 81.795 9.095 82.305 9.325 ;
      RECT 86.385 9.12 86.905 9.295 ;
      RECT 81.625 9.125 82.305 9.295 ;
      RECT 81.795 9.12 86.905 9.29 ;
      RECT 85.78 3.66 86.1 3.98 ;
      RECT 85.755 3.655 86.045 3.885 ;
      RECT 85.71 3.685 86.1 3.86 ;
      RECT 85.58 3.685 86.1 3.855 ;
      RECT 85.78 8.66 86.1 8.98 ;
      RECT 85.755 8.725 86.1 8.955 ;
      RECT 85.58 8.755 86.1 8.925 ;
      RECT 81.57 4.96 81.61 5.22 ;
      RECT 81.61 4.94 81.615 4.95 ;
      RECT 82.94 4.185 82.95 4.406 ;
      RECT 82.87 4.18 82.94 4.531 ;
      RECT 82.86 4.18 82.87 4.658 ;
      RECT 82.835 4.18 82.86 4.705 ;
      RECT 82.81 4.18 82.835 4.783 ;
      RECT 82.79 4.18 82.81 4.853 ;
      RECT 82.765 4.18 82.79 4.893 ;
      RECT 82.755 4.18 82.765 4.913 ;
      RECT 82.745 4.182 82.755 4.921 ;
      RECT 82.74 4.187 82.745 4.378 ;
      RECT 82.74 4.387 82.745 4.922 ;
      RECT 82.735 4.432 82.74 4.923 ;
      RECT 82.725 4.497 82.735 4.924 ;
      RECT 82.715 4.592 82.725 4.926 ;
      RECT 82.71 4.645 82.715 4.928 ;
      RECT 82.705 4.665 82.71 4.929 ;
      RECT 82.65 4.69 82.705 4.935 ;
      RECT 82.61 4.725 82.65 4.944 ;
      RECT 82.6 4.742 82.61 4.949 ;
      RECT 82.591 4.748 82.6 4.951 ;
      RECT 82.505 4.786 82.591 4.962 ;
      RECT 82.5 4.825 82.505 4.972 ;
      RECT 82.425 4.832 82.5 4.982 ;
      RECT 82.405 4.842 82.425 4.993 ;
      RECT 82.375 4.849 82.405 5.001 ;
      RECT 82.35 4.856 82.375 5.008 ;
      RECT 82.326 4.862 82.35 5.013 ;
      RECT 82.24 4.875 82.326 5.025 ;
      RECT 82.162 4.882 82.24 5.043 ;
      RECT 82.076 4.877 82.162 5.061 ;
      RECT 81.99 4.872 82.076 5.081 ;
      RECT 81.91 4.866 81.99 5.098 ;
      RECT 81.845 4.862 81.91 5.127 ;
      RECT 81.84 4.576 81.845 4.6 ;
      RECT 81.83 4.852 81.845 5.155 ;
      RECT 81.835 4.57 81.84 4.64 ;
      RECT 81.83 4.564 81.835 4.71 ;
      RECT 81.825 4.558 81.83 4.788 ;
      RECT 81.825 4.835 81.83 5.22 ;
      RECT 81.817 4.555 81.825 5.22 ;
      RECT 81.731 4.553 81.817 5.22 ;
      RECT 81.645 4.551 81.731 5.22 ;
      RECT 81.635 4.552 81.645 5.22 ;
      RECT 81.63 4.557 81.635 5.22 ;
      RECT 81.62 4.57 81.63 5.22 ;
      RECT 81.615 4.592 81.62 5.22 ;
      RECT 81.61 4.952 81.615 5.22 ;
      RECT 82.24 4.42 82.245 4.64 ;
      RECT 82.745 3.455 82.78 3.715 ;
      RECT 82.73 3.455 82.745 3.723 ;
      RECT 82.701 3.455 82.73 3.745 ;
      RECT 82.615 3.455 82.701 3.805 ;
      RECT 82.595 3.455 82.615 3.87 ;
      RECT 82.535 3.455 82.595 4.035 ;
      RECT 82.53 3.455 82.535 4.183 ;
      RECT 82.525 3.455 82.53 4.195 ;
      RECT 82.52 3.455 82.525 4.221 ;
      RECT 82.49 3.641 82.52 4.301 ;
      RECT 82.485 3.689 82.49 4.39 ;
      RECT 82.48 3.703 82.485 4.405 ;
      RECT 82.475 3.722 82.48 4.435 ;
      RECT 82.47 3.737 82.475 4.451 ;
      RECT 82.465 3.752 82.47 4.473 ;
      RECT 82.46 3.772 82.465 4.495 ;
      RECT 82.45 3.792 82.46 4.528 ;
      RECT 82.435 3.834 82.45 4.59 ;
      RECT 82.43 3.865 82.435 4.63 ;
      RECT 82.425 3.877 82.43 4.635 ;
      RECT 82.42 3.889 82.425 4.64 ;
      RECT 82.415 3.902 82.42 4.64 ;
      RECT 82.41 3.92 82.415 4.64 ;
      RECT 82.405 3.94 82.41 4.64 ;
      RECT 82.4 3.952 82.405 4.64 ;
      RECT 82.395 3.965 82.4 4.64 ;
      RECT 82.375 4 82.395 4.64 ;
      RECT 82.325 4.102 82.375 4.64 ;
      RECT 82.32 4.187 82.325 4.64 ;
      RECT 82.315 4.195 82.32 4.64 ;
      RECT 82.31 4.212 82.315 4.64 ;
      RECT 82.305 4.227 82.31 4.64 ;
      RECT 82.27 4.292 82.305 4.64 ;
      RECT 82.255 4.357 82.27 4.64 ;
      RECT 82.25 4.387 82.255 4.64 ;
      RECT 82.245 4.412 82.25 4.64 ;
      RECT 82.23 4.422 82.24 4.64 ;
      RECT 82.215 4.435 82.23 4.633 ;
      RECT 81.96 4.025 82.03 4.235 ;
      RECT 81.75 4.002 81.755 4.195 ;
      RECT 79.205 3.93 79.465 4.19 ;
      RECT 82.04 4.212 82.045 4.215 ;
      RECT 82.03 4.03 82.04 4.23 ;
      RECT 81.931 4.023 81.96 4.235 ;
      RECT 81.845 4.015 81.931 4.235 ;
      RECT 81.83 4.009 81.845 4.233 ;
      RECT 81.81 4.008 81.83 4.22 ;
      RECT 81.805 4.007 81.81 4.203 ;
      RECT 81.755 4.004 81.805 4.198 ;
      RECT 81.725 4.001 81.75 4.193 ;
      RECT 81.705 3.999 81.725 4.188 ;
      RECT 81.69 3.997 81.705 4.185 ;
      RECT 81.66 3.995 81.69 4.183 ;
      RECT 81.595 3.991 81.66 4.175 ;
      RECT 81.565 3.986 81.595 4.17 ;
      RECT 81.545 3.984 81.565 4.168 ;
      RECT 81.515 3.981 81.545 4.163 ;
      RECT 81.455 3.977 81.515 4.155 ;
      RECT 81.45 3.974 81.455 4.15 ;
      RECT 81.38 3.972 81.45 4.145 ;
      RECT 81.351 3.968 81.38 4.138 ;
      RECT 81.265 3.963 81.351 4.13 ;
      RECT 81.231 3.958 81.265 4.122 ;
      RECT 81.145 3.95 81.231 4.114 ;
      RECT 81.106 3.943 81.145 4.106 ;
      RECT 81.02 3.938 81.106 4.098 ;
      RECT 80.955 3.932 81.02 4.088 ;
      RECT 80.935 3.927 80.955 4.083 ;
      RECT 80.926 3.924 80.935 4.082 ;
      RECT 80.84 3.92 80.926 4.076 ;
      RECT 80.8 3.916 80.84 4.068 ;
      RECT 80.78 3.912 80.8 4.066 ;
      RECT 80.72 3.912 80.78 4.063 ;
      RECT 80.7 3.915 80.72 4.061 ;
      RECT 80.679 3.915 80.7 4.061 ;
      RECT 80.593 3.917 80.679 4.065 ;
      RECT 80.507 3.919 80.593 4.071 ;
      RECT 80.421 3.921 80.507 4.078 ;
      RECT 80.335 3.924 80.421 4.084 ;
      RECT 80.301 3.925 80.335 4.089 ;
      RECT 80.215 3.928 80.301 4.094 ;
      RECT 80.186 3.935 80.215 4.099 ;
      RECT 80.1 3.935 80.186 4.104 ;
      RECT 80.067 3.935 80.1 4.109 ;
      RECT 79.981 3.937 80.067 4.114 ;
      RECT 79.895 3.939 79.981 4.121 ;
      RECT 79.831 3.941 79.895 4.127 ;
      RECT 79.745 3.943 79.831 4.133 ;
      RECT 79.742 3.945 79.745 4.136 ;
      RECT 79.656 3.946 79.742 4.14 ;
      RECT 79.57 3.949 79.656 4.147 ;
      RECT 79.551 3.951 79.57 4.151 ;
      RECT 79.465 3.953 79.551 4.156 ;
      RECT 79.195 3.965 79.205 4.16 ;
      RECT 81.365 10.205 81.655 10.435 ;
      RECT 81.425 9.465 81.595 10.435 ;
      RECT 81.315 9.49 81.69 9.86 ;
      RECT 81.365 9.465 81.655 9.86 ;
      RECT 81.43 3.545 81.615 3.755 ;
      RECT 81.425 3.546 81.62 3.753 ;
      RECT 81.42 3.551 81.63 3.748 ;
      RECT 81.415 3.527 81.42 3.745 ;
      RECT 81.385 3.524 81.415 3.738 ;
      RECT 81.38 3.52 81.385 3.729 ;
      RECT 81.345 3.551 81.63 3.724 ;
      RECT 81.12 3.46 81.38 3.72 ;
      RECT 81.42 3.529 81.425 3.748 ;
      RECT 81.425 3.53 81.43 3.753 ;
      RECT 81.12 3.542 81.5 3.72 ;
      RECT 81.12 3.54 81.485 3.72 ;
      RECT 81.12 3.535 81.475 3.72 ;
      RECT 81.075 4.45 81.125 4.735 ;
      RECT 81.02 4.42 81.025 4.735 ;
      RECT 80.99 4.4 80.995 4.735 ;
      RECT 81.14 4.45 81.2 4.71 ;
      RECT 81.135 4.45 81.14 4.718 ;
      RECT 81.125 4.45 81.135 4.73 ;
      RECT 81.04 4.44 81.075 4.735 ;
      RECT 81.035 4.427 81.04 4.735 ;
      RECT 81.025 4.422 81.035 4.735 ;
      RECT 81.005 4.412 81.02 4.735 ;
      RECT 80.995 4.405 81.005 4.735 ;
      RECT 80.985 4.397 80.99 4.735 ;
      RECT 80.955 4.387 80.985 4.735 ;
      RECT 80.94 4.375 80.955 4.735 ;
      RECT 80.925 4.365 80.94 4.73 ;
      RECT 80.905 4.355 80.925 4.705 ;
      RECT 80.895 4.347 80.905 4.682 ;
      RECT 80.865 4.33 80.895 4.672 ;
      RECT 80.86 4.307 80.865 4.663 ;
      RECT 80.855 4.294 80.86 4.661 ;
      RECT 80.84 4.27 80.855 4.655 ;
      RECT 80.835 4.246 80.84 4.649 ;
      RECT 80.825 4.235 80.835 4.644 ;
      RECT 80.82 4.225 80.825 4.64 ;
      RECT 80.815 4.217 80.82 4.637 ;
      RECT 80.805 4.212 80.815 4.633 ;
      RECT 80.8 4.207 80.805 4.629 ;
      RECT 80.715 4.205 80.8 4.604 ;
      RECT 80.685 4.205 80.715 4.57 ;
      RECT 80.67 4.205 80.685 4.553 ;
      RECT 80.615 4.205 80.67 4.498 ;
      RECT 80.61 4.21 80.615 4.447 ;
      RECT 80.6 4.215 80.61 4.437 ;
      RECT 80.595 4.225 80.6 4.423 ;
      RECT 80.545 4.965 80.805 5.225 ;
      RECT 80.465 4.98 80.805 5.201 ;
      RECT 80.445 4.98 80.805 5.196 ;
      RECT 80.421 4.98 80.805 5.194 ;
      RECT 80.335 4.98 80.805 5.189 ;
      RECT 80.185 4.92 80.445 5.185 ;
      RECT 80.14 4.98 80.805 5.18 ;
      RECT 80.135 4.987 80.805 5.175 ;
      RECT 80.15 4.975 80.465 5.185 ;
      RECT 80.04 3.41 80.3 3.67 ;
      RECT 80.04 3.467 80.305 3.663 ;
      RECT 80.04 3.497 80.31 3.595 ;
      RECT 80.1 3.928 80.215 3.93 ;
      RECT 80.186 3.925 80.215 3.93 ;
      RECT 79.21 4.929 79.235 5.169 ;
      RECT 79.195 4.932 79.285 5.163 ;
      RECT 79.19 4.937 79.371 5.158 ;
      RECT 79.185 4.945 79.435 5.156 ;
      RECT 79.185 4.945 79.445 5.155 ;
      RECT 79.18 4.952 79.455 5.148 ;
      RECT 79.18 4.952 79.541 5.137 ;
      RECT 79.175 4.987 79.541 5.133 ;
      RECT 79.175 4.987 79.55 5.122 ;
      RECT 79.455 4.86 79.715 5.12 ;
      RECT 79.165 5.037 79.715 5.118 ;
      RECT 79.435 4.905 79.455 5.153 ;
      RECT 79.371 4.908 79.435 5.157 ;
      RECT 79.285 4.913 79.371 5.162 ;
      RECT 79.215 4.924 79.715 5.12 ;
      RECT 79.235 4.918 79.285 5.167 ;
      RECT 79.36 3.395 79.37 3.657 ;
      RECT 79.35 3.452 79.36 3.66 ;
      RECT 79.325 3.457 79.35 3.666 ;
      RECT 79.3 3.461 79.325 3.678 ;
      RECT 79.29 3.464 79.3 3.688 ;
      RECT 79.285 3.465 79.29 3.693 ;
      RECT 79.28 3.466 79.285 3.698 ;
      RECT 79.275 3.467 79.28 3.7 ;
      RECT 79.25 3.47 79.275 3.703 ;
      RECT 79.22 3.476 79.25 3.706 ;
      RECT 79.155 3.487 79.22 3.709 ;
      RECT 79.11 3.495 79.155 3.713 ;
      RECT 79.095 3.495 79.11 3.721 ;
      RECT 79.09 3.496 79.095 3.728 ;
      RECT 79.085 3.498 79.09 3.731 ;
      RECT 79.08 3.502 79.085 3.734 ;
      RECT 79.07 3.51 79.08 3.738 ;
      RECT 79.065 3.523 79.07 3.743 ;
      RECT 79.06 3.531 79.065 3.745 ;
      RECT 79.055 3.537 79.06 3.745 ;
      RECT 79.05 3.541 79.055 3.748 ;
      RECT 79.045 3.543 79.05 3.751 ;
      RECT 79.04 3.546 79.045 3.754 ;
      RECT 79.03 3.551 79.04 3.758 ;
      RECT 79.025 3.557 79.03 3.763 ;
      RECT 79.015 3.563 79.025 3.767 ;
      RECT 79 3.57 79.015 3.773 ;
      RECT 78.971 3.584 79 3.783 ;
      RECT 78.885 3.619 78.971 3.815 ;
      RECT 78.865 3.652 78.885 3.844 ;
      RECT 78.845 3.665 78.865 3.855 ;
      RECT 78.825 3.677 78.845 3.866 ;
      RECT 78.775 3.699 78.825 3.886 ;
      RECT 78.76 3.717 78.775 3.903 ;
      RECT 78.755 3.723 78.76 3.906 ;
      RECT 78.75 3.727 78.755 3.909 ;
      RECT 78.745 3.731 78.75 3.913 ;
      RECT 78.74 3.733 78.745 3.916 ;
      RECT 78.73 3.74 78.74 3.919 ;
      RECT 78.725 3.745 78.73 3.923 ;
      RECT 78.72 3.747 78.725 3.926 ;
      RECT 78.715 3.751 78.72 3.929 ;
      RECT 78.71 3.753 78.715 3.933 ;
      RECT 78.695 3.758 78.71 3.938 ;
      RECT 78.69 3.763 78.695 3.941 ;
      RECT 78.685 3.771 78.69 3.944 ;
      RECT 78.68 3.773 78.685 3.947 ;
      RECT 78.675 3.775 78.68 3.95 ;
      RECT 78.665 3.777 78.675 3.956 ;
      RECT 78.63 3.791 78.665 3.968 ;
      RECT 78.62 3.806 78.63 3.978 ;
      RECT 78.545 3.835 78.62 4.002 ;
      RECT 78.54 3.86 78.545 4.025 ;
      RECT 78.525 3.864 78.54 4.031 ;
      RECT 78.515 3.872 78.525 4.036 ;
      RECT 78.485 3.885 78.515 4.04 ;
      RECT 78.475 3.9 78.485 4.045 ;
      RECT 78.465 3.905 78.475 4.048 ;
      RECT 78.46 3.907 78.465 4.05 ;
      RECT 78.445 3.91 78.46 4.053 ;
      RECT 78.44 3.912 78.445 4.056 ;
      RECT 78.42 3.917 78.44 4.06 ;
      RECT 78.39 3.922 78.42 4.068 ;
      RECT 78.365 3.929 78.39 4.076 ;
      RECT 78.36 3.934 78.365 4.081 ;
      RECT 78.33 3.937 78.36 4.085 ;
      RECT 78.29 3.94 78.33 4.095 ;
      RECT 78.255 3.937 78.29 4.107 ;
      RECT 78.245 3.933 78.255 4.114 ;
      RECT 78.22 3.929 78.245 4.12 ;
      RECT 78.215 3.925 78.22 4.125 ;
      RECT 78.175 3.922 78.215 4.125 ;
      RECT 78.16 3.907 78.175 4.126 ;
      RECT 78.137 3.895 78.16 4.126 ;
      RECT 78.051 3.895 78.137 4.127 ;
      RECT 77.965 3.895 78.051 4.129 ;
      RECT 77.945 3.895 77.965 4.126 ;
      RECT 77.94 3.9 77.945 4.121 ;
      RECT 77.935 3.905 77.94 4.119 ;
      RECT 77.925 3.915 77.935 4.117 ;
      RECT 77.92 3.921 77.925 4.11 ;
      RECT 77.915 3.923 77.92 4.095 ;
      RECT 77.91 3.927 77.915 4.085 ;
      RECT 79.37 3.395 79.62 3.655 ;
      RECT 77.095 4.93 77.355 5.19 ;
      RECT 79.39 4.42 79.395 4.63 ;
      RECT 79.395 4.425 79.405 4.625 ;
      RECT 79.345 4.42 79.39 4.645 ;
      RECT 79.335 4.42 79.345 4.665 ;
      RECT 79.316 4.42 79.335 4.67 ;
      RECT 79.23 4.42 79.316 4.667 ;
      RECT 79.2 4.422 79.23 4.665 ;
      RECT 79.145 4.432 79.2 4.663 ;
      RECT 79.08 4.446 79.145 4.661 ;
      RECT 79.075 4.454 79.08 4.66 ;
      RECT 79.06 4.457 79.075 4.658 ;
      RECT 78.995 4.467 79.06 4.654 ;
      RECT 78.947 4.481 78.995 4.655 ;
      RECT 78.861 4.498 78.947 4.669 ;
      RECT 78.775 4.519 78.861 4.686 ;
      RECT 78.755 4.532 78.775 4.696 ;
      RECT 78.71 4.54 78.755 4.703 ;
      RECT 78.675 4.548 78.71 4.711 ;
      RECT 78.641 4.556 78.675 4.719 ;
      RECT 78.555 4.57 78.641 4.731 ;
      RECT 78.52 4.587 78.555 4.743 ;
      RECT 78.511 4.596 78.52 4.747 ;
      RECT 78.425 4.614 78.511 4.764 ;
      RECT 78.366 4.641 78.425 4.791 ;
      RECT 78.28 4.668 78.366 4.819 ;
      RECT 78.26 4.69 78.28 4.839 ;
      RECT 78.2 4.705 78.26 4.855 ;
      RECT 78.19 4.717 78.2 4.868 ;
      RECT 78.185 4.722 78.19 4.871 ;
      RECT 78.175 4.725 78.185 4.874 ;
      RECT 78.17 4.727 78.175 4.877 ;
      RECT 78.14 4.735 78.17 4.884 ;
      RECT 78.125 4.742 78.14 4.892 ;
      RECT 78.115 4.747 78.125 4.896 ;
      RECT 78.11 4.75 78.115 4.899 ;
      RECT 78.1 4.752 78.11 4.902 ;
      RECT 78.065 4.762 78.1 4.911 ;
      RECT 77.99 4.785 78.065 4.933 ;
      RECT 77.97 4.803 77.99 4.951 ;
      RECT 77.94 4.81 77.97 4.961 ;
      RECT 77.92 4.818 77.94 4.971 ;
      RECT 77.91 4.824 77.92 4.978 ;
      RECT 77.891 4.829 77.91 4.984 ;
      RECT 77.805 4.849 77.891 5.004 ;
      RECT 77.79 4.869 77.805 5.023 ;
      RECT 77.745 4.881 77.79 5.034 ;
      RECT 77.68 4.902 77.745 5.057 ;
      RECT 77.64 4.922 77.68 5.078 ;
      RECT 77.63 4.932 77.64 5.088 ;
      RECT 77.58 4.944 77.63 5.099 ;
      RECT 77.56 4.96 77.58 5.111 ;
      RECT 77.53 4.97 77.56 5.117 ;
      RECT 77.52 4.975 77.53 5.119 ;
      RECT 77.451 4.976 77.52 5.125 ;
      RECT 77.365 4.978 77.451 5.135 ;
      RECT 77.355 4.979 77.365 5.14 ;
      RECT 78.625 5.005 78.815 5.215 ;
      RECT 78.615 5.01 78.825 5.208 ;
      RECT 78.6 5.01 78.825 5.173 ;
      RECT 78.52 4.895 78.78 5.155 ;
      RECT 77.435 4.425 77.62 4.72 ;
      RECT 77.425 4.425 77.62 4.718 ;
      RECT 77.41 4.425 77.625 4.713 ;
      RECT 77.41 4.425 77.63 4.71 ;
      RECT 77.405 4.425 77.63 4.708 ;
      RECT 77.4 4.68 77.63 4.698 ;
      RECT 77.405 4.425 77.665 4.685 ;
      RECT 77.365 3.46 77.625 3.72 ;
      RECT 77.175 3.385 77.261 3.718 ;
      RECT 77.15 3.389 77.305 3.714 ;
      RECT 77.261 3.381 77.305 3.714 ;
      RECT 77.261 3.382 77.31 3.713 ;
      RECT 77.175 3.387 77.325 3.712 ;
      RECT 77.15 3.395 77.365 3.711 ;
      RECT 77.145 3.39 77.325 3.706 ;
      RECT 77.135 3.405 77.365 3.613 ;
      RECT 77.135 3.457 77.565 3.613 ;
      RECT 77.135 3.45 77.545 3.613 ;
      RECT 77.135 3.437 77.515 3.613 ;
      RECT 77.135 3.425 77.455 3.613 ;
      RECT 77.135 3.41 77.43 3.613 ;
      RECT 76.335 4.04 76.47 4.335 ;
      RECT 76.595 4.063 76.6 4.25 ;
      RECT 77.315 3.96 77.46 4.195 ;
      RECT 77.475 3.96 77.48 4.185 ;
      RECT 77.51 3.971 77.515 4.165 ;
      RECT 77.505 3.963 77.51 4.17 ;
      RECT 77.485 3.96 77.505 4.175 ;
      RECT 77.48 3.96 77.485 4.183 ;
      RECT 77.47 3.96 77.475 4.188 ;
      RECT 77.46 3.96 77.47 4.193 ;
      RECT 77.29 3.962 77.315 4.195 ;
      RECT 77.24 3.969 77.29 4.195 ;
      RECT 77.235 3.974 77.24 4.195 ;
      RECT 77.196 3.979 77.235 4.196 ;
      RECT 77.11 3.991 77.196 4.197 ;
      RECT 77.101 4.001 77.11 4.197 ;
      RECT 77.015 4.01 77.101 4.199 ;
      RECT 76.991 4.02 77.015 4.201 ;
      RECT 76.905 4.031 76.991 4.202 ;
      RECT 76.875 4.042 76.905 4.204 ;
      RECT 76.845 4.047 76.875 4.206 ;
      RECT 76.82 4.053 76.845 4.209 ;
      RECT 76.805 4.058 76.82 4.21 ;
      RECT 76.76 4.064 76.805 4.21 ;
      RECT 76.755 4.069 76.76 4.211 ;
      RECT 76.735 4.069 76.755 4.213 ;
      RECT 76.715 4.067 76.735 4.218 ;
      RECT 76.68 4.066 76.715 4.225 ;
      RECT 76.65 4.065 76.68 4.235 ;
      RECT 76.6 4.064 76.65 4.245 ;
      RECT 76.51 4.061 76.595 4.335 ;
      RECT 76.485 4.055 76.51 4.335 ;
      RECT 76.47 4.045 76.485 4.335 ;
      RECT 76.285 4.04 76.335 4.255 ;
      RECT 76.275 4.045 76.285 4.245 ;
      RECT 76.515 4.52 76.775 4.78 ;
      RECT 76.515 4.52 76.805 4.673 ;
      RECT 76.515 4.52 76.84 4.658 ;
      RECT 76.77 4.44 76.96 4.65 ;
      RECT 76.76 4.445 76.97 4.643 ;
      RECT 76.725 4.515 76.97 4.643 ;
      RECT 76.755 4.457 76.775 4.78 ;
      RECT 76.74 4.505 76.97 4.643 ;
      RECT 76.745 4.477 76.775 4.78 ;
      RECT 75.825 3.545 75.895 4.65 ;
      RECT 76.56 3.65 76.82 3.91 ;
      RECT 76.14 3.696 76.155 3.905 ;
      RECT 76.476 3.709 76.56 3.86 ;
      RECT 76.39 3.706 76.476 3.86 ;
      RECT 76.351 3.704 76.39 3.86 ;
      RECT 76.265 3.702 76.351 3.86 ;
      RECT 76.205 3.7 76.265 3.871 ;
      RECT 76.17 3.698 76.205 3.889 ;
      RECT 76.155 3.696 76.17 3.9 ;
      RECT 76.125 3.696 76.14 3.913 ;
      RECT 76.115 3.696 76.125 3.918 ;
      RECT 76.09 3.695 76.115 3.923 ;
      RECT 76.075 3.69 76.09 3.929 ;
      RECT 76.07 3.683 76.075 3.934 ;
      RECT 76.045 3.674 76.07 3.94 ;
      RECT 76 3.653 76.045 3.953 ;
      RECT 75.99 3.637 76 3.963 ;
      RECT 75.975 3.63 75.99 3.973 ;
      RECT 75.965 3.623 75.975 3.99 ;
      RECT 75.96 3.62 75.965 4.02 ;
      RECT 75.955 3.618 75.96 4.05 ;
      RECT 75.95 3.616 75.955 4.087 ;
      RECT 75.935 3.612 75.95 4.154 ;
      RECT 75.935 4.445 75.945 4.645 ;
      RECT 75.93 3.608 75.935 4.28 ;
      RECT 75.93 4.432 75.935 4.65 ;
      RECT 75.925 3.606 75.93 4.365 ;
      RECT 75.925 4.422 75.93 4.65 ;
      RECT 75.91 3.577 75.925 4.65 ;
      RECT 75.895 3.55 75.91 4.65 ;
      RECT 75.82 3.545 75.825 3.9 ;
      RECT 75.82 3.955 75.825 4.65 ;
      RECT 75.805 3.545 75.82 3.878 ;
      RECT 75.815 3.977 75.82 4.65 ;
      RECT 75.805 4.017 75.815 4.65 ;
      RECT 75.77 3.545 75.805 3.82 ;
      RECT 75.8 4.052 75.805 4.65 ;
      RECT 75.785 4.107 75.8 4.65 ;
      RECT 75.78 4.172 75.785 4.65 ;
      RECT 75.765 4.22 75.78 4.65 ;
      RECT 75.74 3.545 75.77 3.775 ;
      RECT 75.76 4.275 75.765 4.65 ;
      RECT 75.745 4.335 75.76 4.65 ;
      RECT 75.74 4.383 75.745 4.648 ;
      RECT 75.735 3.545 75.74 3.768 ;
      RECT 75.735 4.415 75.74 4.643 ;
      RECT 75.71 3.545 75.735 3.76 ;
      RECT 75.7 3.55 75.71 3.75 ;
      RECT 75.915 4.825 75.935 5.065 ;
      RECT 75.145 4.755 75.15 4.965 ;
      RECT 76.425 4.828 76.435 5.023 ;
      RECT 76.42 4.818 76.425 5.026 ;
      RECT 76.34 4.815 76.42 5.049 ;
      RECT 76.336 4.815 76.34 5.071 ;
      RECT 76.25 4.815 76.336 5.081 ;
      RECT 76.235 4.815 76.25 5.089 ;
      RECT 76.206 4.816 76.235 5.087 ;
      RECT 76.12 4.821 76.206 5.083 ;
      RECT 76.107 4.825 76.12 5.079 ;
      RECT 76.021 4.825 76.107 5.075 ;
      RECT 75.935 4.825 76.021 5.069 ;
      RECT 75.851 4.825 75.915 5.063 ;
      RECT 75.765 4.825 75.851 5.058 ;
      RECT 75.745 4.825 75.765 5.054 ;
      RECT 75.685 4.82 75.745 5.051 ;
      RECT 75.657 4.814 75.685 5.048 ;
      RECT 75.571 4.809 75.657 5.044 ;
      RECT 75.485 4.803 75.571 5.038 ;
      RECT 75.41 4.785 75.485 5.033 ;
      RECT 75.375 4.762 75.41 5.029 ;
      RECT 75.365 4.752 75.375 5.028 ;
      RECT 75.31 4.75 75.365 5.027 ;
      RECT 75.235 4.75 75.31 5.023 ;
      RECT 75.225 4.75 75.235 5.018 ;
      RECT 75.21 4.75 75.225 5.01 ;
      RECT 75.16 4.752 75.21 4.988 ;
      RECT 75.15 4.755 75.16 4.968 ;
      RECT 75.14 4.76 75.145 4.963 ;
      RECT 75.135 4.765 75.14 4.958 ;
      RECT 73.245 3.41 73.505 3.67 ;
      RECT 73.235 3.44 73.505 3.65 ;
      RECT 75.155 3.355 75.415 3.615 ;
      RECT 75.15 3.43 75.155 3.616 ;
      RECT 75.125 3.435 75.15 3.618 ;
      RECT 75.11 3.442 75.125 3.621 ;
      RECT 75.05 3.46 75.11 3.626 ;
      RECT 75.02 3.48 75.05 3.633 ;
      RECT 74.995 3.488 75.02 3.638 ;
      RECT 74.97 3.496 74.995 3.64 ;
      RECT 74.952 3.5 74.97 3.639 ;
      RECT 74.866 3.498 74.952 3.639 ;
      RECT 74.78 3.496 74.866 3.639 ;
      RECT 74.694 3.494 74.78 3.638 ;
      RECT 74.608 3.492 74.694 3.638 ;
      RECT 74.522 3.49 74.608 3.638 ;
      RECT 74.436 3.488 74.522 3.638 ;
      RECT 74.35 3.486 74.436 3.637 ;
      RECT 74.332 3.485 74.35 3.637 ;
      RECT 74.246 3.484 74.332 3.637 ;
      RECT 74.16 3.482 74.246 3.637 ;
      RECT 74.074 3.481 74.16 3.636 ;
      RECT 73.988 3.48 74.074 3.636 ;
      RECT 73.902 3.478 73.988 3.636 ;
      RECT 73.816 3.477 73.902 3.636 ;
      RECT 73.73 3.475 73.816 3.635 ;
      RECT 73.706 3.473 73.73 3.635 ;
      RECT 73.62 3.466 73.706 3.635 ;
      RECT 73.591 3.458 73.62 3.635 ;
      RECT 73.505 3.45 73.591 3.635 ;
      RECT 73.225 3.447 73.235 3.645 ;
      RECT 74.73 4.41 74.735 4.76 ;
      RECT 74.5 4.5 74.64 4.76 ;
      RECT 74.975 4.185 75.02 4.395 ;
      RECT 75.03 4.196 75.04 4.39 ;
      RECT 75.02 4.188 75.03 4.395 ;
      RECT 74.955 4.185 74.975 4.4 ;
      RECT 74.925 4.185 74.955 4.423 ;
      RECT 74.915 4.185 74.925 4.448 ;
      RECT 74.91 4.185 74.915 4.458 ;
      RECT 74.855 4.185 74.91 4.498 ;
      RECT 74.85 4.185 74.855 4.538 ;
      RECT 74.845 4.187 74.85 4.543 ;
      RECT 74.83 4.197 74.845 4.554 ;
      RECT 74.785 4.255 74.83 4.59 ;
      RECT 74.775 4.31 74.785 4.624 ;
      RECT 74.76 4.337 74.775 4.64 ;
      RECT 74.75 4.364 74.76 4.76 ;
      RECT 74.735 4.387 74.75 4.76 ;
      RECT 74.725 4.427 74.73 4.76 ;
      RECT 74.72 4.437 74.725 4.76 ;
      RECT 74.715 4.452 74.72 4.76 ;
      RECT 74.705 4.457 74.715 4.76 ;
      RECT 74.64 4.48 74.705 4.76 ;
      RECT 74.11 3.975 74.33 4.185 ;
      RECT 74.11 3.982 74.34 4.18 ;
      RECT 73.415 3.99 74.34 4.165 ;
      RECT 73.935 3.885 74.325 4.165 ;
      RECT 72.715 3.9 72.975 4.16 ;
      RECT 73.35 3.935 73.485 4.12 ;
      RECT 73.275 3.925 73.37 4.115 ;
      RECT 73.265 3.99 74.34 4.111 ;
      RECT 73.015 3.99 74.34 4.11 ;
      RECT 73.04 3.91 73.28 4.11 ;
      RECT 72.715 3.915 73.3 4.098 ;
      RECT 74.63 3.94 74.67 4.025 ;
      RECT 72.715 3.975 73.89 4.098 ;
      RECT 72.715 3.965 73.775 4.098 ;
      RECT 72.715 3.946 73.68 4.098 ;
      RECT 73.5 3.94 73.68 4.165 ;
      RECT 73.935 3.92 74.63 3.955 ;
      RECT 73.035 3.912 73.28 4.11 ;
      RECT 73.05 3.902 73.26 4.11 ;
      RECT 73.065 3.895 73.26 4.11 ;
      RECT 73.23 4.415 73.49 4.675 ;
      RECT 73.23 4.455 73.595 4.665 ;
      RECT 73.23 4.457 73.6 4.664 ;
      RECT 73.23 4.465 73.605 4.661 ;
      RECT 72.155 3.54 72.255 5.065 ;
      RECT 72.345 4.68 72.395 4.94 ;
      RECT 72.34 3.553 72.345 3.74 ;
      RECT 72.335 4.661 72.345 4.94 ;
      RECT 72.335 3.55 72.34 3.748 ;
      RECT 72.32 3.544 72.335 3.755 ;
      RECT 72.33 4.649 72.335 5.023 ;
      RECT 72.32 4.637 72.33 5.06 ;
      RECT 72.31 3.54 72.32 3.762 ;
      RECT 72.31 4.622 72.32 5.065 ;
      RECT 72.305 3.54 72.31 3.77 ;
      RECT 72.285 4.592 72.31 5.065 ;
      RECT 72.265 3.54 72.305 3.818 ;
      RECT 72.275 4.552 72.285 5.065 ;
      RECT 72.265 4.507 72.275 5.065 ;
      RECT 72.26 3.54 72.265 3.888 ;
      RECT 72.26 4.465 72.265 5.065 ;
      RECT 72.255 3.54 72.26 4.365 ;
      RECT 72.255 4.447 72.26 5.065 ;
      RECT 72.145 3.543 72.155 5.065 ;
      RECT 72.13 3.55 72.145 5.061 ;
      RECT 72.125 3.56 72.13 5.056 ;
      RECT 72.12 3.76 72.125 4.948 ;
      RECT 72.115 3.845 72.12 4.5 ;
      RECT 70.98 10.205 71.275 10.435 ;
      RECT 71.04 8.725 71.21 10.435 ;
      RECT 70.99 9.095 71.34 9.445 ;
      RECT 70.98 8.725 71.27 8.955 ;
      RECT 69.99 10.205 70.285 10.435 ;
      RECT 70.05 8.725 70.22 10.435 ;
      RECT 69.99 8.725 70.28 8.955 ;
      RECT 69.99 8.76 70.84 8.92 ;
      RECT 70.675 8.355 70.84 8.92 ;
      RECT 69.99 8.755 70.385 8.92 ;
      RECT 70.61 8.355 70.9 8.585 ;
      RECT 70.61 8.385 71.07 8.555 ;
      RECT 70.575 4.025 70.895 4.26 ;
      RECT 70.575 4.055 71.065 4.225 ;
      RECT 70.575 3.69 70.765 4.26 ;
      RECT 69.99 3.655 70.28 3.885 ;
      RECT 69.99 3.69 70.765 3.86 ;
      RECT 70.05 2.175 70.22 3.885 ;
      RECT 69.99 2.175 70.285 2.405 ;
      RECT 69.62 4.025 69.91 4.255 ;
      RECT 69.62 4.055 70.08 4.225 ;
      RECT 69.685 2.95 69.85 4.255 ;
      RECT 68.2 2.915 68.49 3.145 ;
      RECT 68.2 2.95 69.85 3.12 ;
      RECT 68.26 2.175 68.43 3.145 ;
      RECT 68.2 2.175 68.49 2.405 ;
      RECT 68.2 10.205 68.49 10.435 ;
      RECT 68.26 9.465 68.43 10.435 ;
      RECT 68.26 9.555 69.85 9.725 ;
      RECT 69.68 8.355 69.85 9.725 ;
      RECT 68.2 9.465 68.49 9.695 ;
      RECT 69.62 8.355 69.91 8.585 ;
      RECT 69.62 8.385 70.08 8.555 ;
      RECT 66.235 4.725 66.585 5.075 ;
      RECT 66.325 3.32 66.495 5.075 ;
      RECT 68.63 3.26 68.98 3.61 ;
      RECT 66.325 3.32 67.945 3.495 ;
      RECT 66.325 3.32 68.6 3.49 ;
      RECT 68.46 3.315 68.98 3.485 ;
      RECT 68.655 9.09 68.98 9.415 ;
      RECT 64.085 9.05 64.435 9.4 ;
      RECT 68.63 9.095 68.98 9.325 ;
      RECT 63.87 9.095 64.435 9.325 ;
      RECT 68.46 9.12 68.98 9.295 ;
      RECT 63.7 9.125 64.435 9.295 ;
      RECT 63.87 9.12 68.98 9.29 ;
      RECT 67.855 3.66 68.175 3.98 ;
      RECT 67.83 3.655 68.12 3.885 ;
      RECT 67.785 3.685 68.175 3.86 ;
      RECT 67.655 3.685 68.175 3.855 ;
      RECT 67.855 8.66 68.175 8.98 ;
      RECT 67.83 8.725 68.175 8.955 ;
      RECT 67.655 8.755 68.175 8.925 ;
      RECT 63.645 4.96 63.685 5.22 ;
      RECT 63.685 4.94 63.69 4.95 ;
      RECT 65.015 4.185 65.025 4.406 ;
      RECT 64.945 4.18 65.015 4.531 ;
      RECT 64.935 4.18 64.945 4.658 ;
      RECT 64.91 4.18 64.935 4.705 ;
      RECT 64.885 4.18 64.91 4.783 ;
      RECT 64.865 4.18 64.885 4.853 ;
      RECT 64.84 4.18 64.865 4.893 ;
      RECT 64.83 4.18 64.84 4.913 ;
      RECT 64.82 4.182 64.83 4.921 ;
      RECT 64.815 4.187 64.82 4.378 ;
      RECT 64.815 4.387 64.82 4.922 ;
      RECT 64.81 4.432 64.815 4.923 ;
      RECT 64.8 4.497 64.81 4.924 ;
      RECT 64.79 4.592 64.8 4.926 ;
      RECT 64.785 4.645 64.79 4.928 ;
      RECT 64.78 4.665 64.785 4.929 ;
      RECT 64.725 4.69 64.78 4.935 ;
      RECT 64.685 4.725 64.725 4.944 ;
      RECT 64.675 4.742 64.685 4.949 ;
      RECT 64.666 4.748 64.675 4.951 ;
      RECT 64.58 4.786 64.666 4.962 ;
      RECT 64.575 4.825 64.58 4.972 ;
      RECT 64.5 4.832 64.575 4.982 ;
      RECT 64.48 4.842 64.5 4.993 ;
      RECT 64.45 4.849 64.48 5.001 ;
      RECT 64.425 4.856 64.45 5.008 ;
      RECT 64.401 4.862 64.425 5.013 ;
      RECT 64.315 4.875 64.401 5.025 ;
      RECT 64.237 4.882 64.315 5.043 ;
      RECT 64.151 4.877 64.237 5.061 ;
      RECT 64.065 4.872 64.151 5.081 ;
      RECT 63.985 4.866 64.065 5.098 ;
      RECT 63.92 4.862 63.985 5.127 ;
      RECT 63.915 4.576 63.92 4.6 ;
      RECT 63.905 4.852 63.92 5.155 ;
      RECT 63.91 4.57 63.915 4.64 ;
      RECT 63.905 4.564 63.91 4.71 ;
      RECT 63.9 4.558 63.905 4.788 ;
      RECT 63.9 4.835 63.905 5.22 ;
      RECT 63.892 4.555 63.9 5.22 ;
      RECT 63.806 4.553 63.892 5.22 ;
      RECT 63.72 4.551 63.806 5.22 ;
      RECT 63.71 4.552 63.72 5.22 ;
      RECT 63.705 4.557 63.71 5.22 ;
      RECT 63.695 4.57 63.705 5.22 ;
      RECT 63.69 4.592 63.695 5.22 ;
      RECT 63.685 4.952 63.69 5.22 ;
      RECT 64.315 4.42 64.32 4.64 ;
      RECT 64.82 3.455 64.855 3.715 ;
      RECT 64.805 3.455 64.82 3.723 ;
      RECT 64.776 3.455 64.805 3.745 ;
      RECT 64.69 3.455 64.776 3.805 ;
      RECT 64.67 3.455 64.69 3.87 ;
      RECT 64.61 3.455 64.67 4.035 ;
      RECT 64.605 3.455 64.61 4.183 ;
      RECT 64.6 3.455 64.605 4.195 ;
      RECT 64.595 3.455 64.6 4.221 ;
      RECT 64.565 3.641 64.595 4.301 ;
      RECT 64.56 3.689 64.565 4.39 ;
      RECT 64.555 3.703 64.56 4.405 ;
      RECT 64.55 3.722 64.555 4.435 ;
      RECT 64.545 3.737 64.55 4.451 ;
      RECT 64.54 3.752 64.545 4.473 ;
      RECT 64.535 3.772 64.54 4.495 ;
      RECT 64.525 3.792 64.535 4.528 ;
      RECT 64.51 3.834 64.525 4.59 ;
      RECT 64.505 3.865 64.51 4.63 ;
      RECT 64.5 3.877 64.505 4.635 ;
      RECT 64.495 3.889 64.5 4.64 ;
      RECT 64.49 3.902 64.495 4.64 ;
      RECT 64.485 3.92 64.49 4.64 ;
      RECT 64.48 3.94 64.485 4.64 ;
      RECT 64.475 3.952 64.48 4.64 ;
      RECT 64.47 3.965 64.475 4.64 ;
      RECT 64.45 4 64.47 4.64 ;
      RECT 64.4 4.102 64.45 4.64 ;
      RECT 64.395 4.187 64.4 4.64 ;
      RECT 64.39 4.195 64.395 4.64 ;
      RECT 64.385 4.212 64.39 4.64 ;
      RECT 64.38 4.227 64.385 4.64 ;
      RECT 64.345 4.292 64.38 4.64 ;
      RECT 64.33 4.357 64.345 4.64 ;
      RECT 64.325 4.387 64.33 4.64 ;
      RECT 64.32 4.412 64.325 4.64 ;
      RECT 64.305 4.422 64.315 4.64 ;
      RECT 64.29 4.435 64.305 4.633 ;
      RECT 64.035 4.025 64.105 4.235 ;
      RECT 63.825 4.002 63.83 4.195 ;
      RECT 61.28 3.93 61.54 4.19 ;
      RECT 64.115 4.212 64.12 4.215 ;
      RECT 64.105 4.03 64.115 4.23 ;
      RECT 64.006 4.023 64.035 4.235 ;
      RECT 63.92 4.015 64.006 4.235 ;
      RECT 63.905 4.009 63.92 4.233 ;
      RECT 63.885 4.008 63.905 4.22 ;
      RECT 63.88 4.007 63.885 4.203 ;
      RECT 63.83 4.004 63.88 4.198 ;
      RECT 63.8 4.001 63.825 4.193 ;
      RECT 63.78 3.999 63.8 4.188 ;
      RECT 63.765 3.997 63.78 4.185 ;
      RECT 63.735 3.995 63.765 4.183 ;
      RECT 63.67 3.991 63.735 4.175 ;
      RECT 63.64 3.986 63.67 4.17 ;
      RECT 63.62 3.984 63.64 4.168 ;
      RECT 63.59 3.981 63.62 4.163 ;
      RECT 63.53 3.977 63.59 4.155 ;
      RECT 63.525 3.974 63.53 4.15 ;
      RECT 63.455 3.972 63.525 4.145 ;
      RECT 63.426 3.968 63.455 4.138 ;
      RECT 63.34 3.963 63.426 4.13 ;
      RECT 63.306 3.958 63.34 4.122 ;
      RECT 63.22 3.95 63.306 4.114 ;
      RECT 63.181 3.943 63.22 4.106 ;
      RECT 63.095 3.938 63.181 4.098 ;
      RECT 63.03 3.932 63.095 4.088 ;
      RECT 63.01 3.927 63.03 4.083 ;
      RECT 63.001 3.924 63.01 4.082 ;
      RECT 62.915 3.92 63.001 4.076 ;
      RECT 62.875 3.916 62.915 4.068 ;
      RECT 62.855 3.912 62.875 4.066 ;
      RECT 62.795 3.912 62.855 4.063 ;
      RECT 62.775 3.915 62.795 4.061 ;
      RECT 62.754 3.915 62.775 4.061 ;
      RECT 62.668 3.917 62.754 4.065 ;
      RECT 62.582 3.919 62.668 4.071 ;
      RECT 62.496 3.921 62.582 4.078 ;
      RECT 62.41 3.924 62.496 4.084 ;
      RECT 62.376 3.925 62.41 4.089 ;
      RECT 62.29 3.928 62.376 4.094 ;
      RECT 62.261 3.935 62.29 4.099 ;
      RECT 62.175 3.935 62.261 4.104 ;
      RECT 62.142 3.935 62.175 4.109 ;
      RECT 62.056 3.937 62.142 4.114 ;
      RECT 61.97 3.939 62.056 4.121 ;
      RECT 61.906 3.941 61.97 4.127 ;
      RECT 61.82 3.943 61.906 4.133 ;
      RECT 61.817 3.945 61.82 4.136 ;
      RECT 61.731 3.946 61.817 4.14 ;
      RECT 61.645 3.949 61.731 4.147 ;
      RECT 61.626 3.951 61.645 4.151 ;
      RECT 61.54 3.953 61.626 4.156 ;
      RECT 61.27 3.965 61.28 4.16 ;
      RECT 63.44 10.205 63.73 10.435 ;
      RECT 63.5 9.465 63.67 10.435 ;
      RECT 63.39 9.49 63.765 9.86 ;
      RECT 63.44 9.465 63.73 9.86 ;
      RECT 63.505 3.545 63.69 3.755 ;
      RECT 63.5 3.546 63.695 3.753 ;
      RECT 63.495 3.551 63.705 3.748 ;
      RECT 63.49 3.527 63.495 3.745 ;
      RECT 63.46 3.524 63.49 3.738 ;
      RECT 63.455 3.52 63.46 3.729 ;
      RECT 63.42 3.551 63.705 3.724 ;
      RECT 63.195 3.46 63.455 3.72 ;
      RECT 63.495 3.529 63.5 3.748 ;
      RECT 63.5 3.53 63.505 3.753 ;
      RECT 63.195 3.542 63.575 3.72 ;
      RECT 63.195 3.54 63.56 3.72 ;
      RECT 63.195 3.535 63.55 3.72 ;
      RECT 63.15 4.45 63.2 4.735 ;
      RECT 63.095 4.42 63.1 4.735 ;
      RECT 63.065 4.4 63.07 4.735 ;
      RECT 63.215 4.45 63.275 4.71 ;
      RECT 63.21 4.45 63.215 4.718 ;
      RECT 63.2 4.45 63.21 4.73 ;
      RECT 63.115 4.44 63.15 4.735 ;
      RECT 63.11 4.427 63.115 4.735 ;
      RECT 63.1 4.422 63.11 4.735 ;
      RECT 63.08 4.412 63.095 4.735 ;
      RECT 63.07 4.405 63.08 4.735 ;
      RECT 63.06 4.397 63.065 4.735 ;
      RECT 63.03 4.387 63.06 4.735 ;
      RECT 63.015 4.375 63.03 4.735 ;
      RECT 63 4.365 63.015 4.73 ;
      RECT 62.98 4.355 63 4.705 ;
      RECT 62.97 4.347 62.98 4.682 ;
      RECT 62.94 4.33 62.97 4.672 ;
      RECT 62.935 4.307 62.94 4.663 ;
      RECT 62.93 4.294 62.935 4.661 ;
      RECT 62.915 4.27 62.93 4.655 ;
      RECT 62.91 4.246 62.915 4.649 ;
      RECT 62.9 4.235 62.91 4.644 ;
      RECT 62.895 4.225 62.9 4.64 ;
      RECT 62.89 4.217 62.895 4.637 ;
      RECT 62.88 4.212 62.89 4.633 ;
      RECT 62.875 4.207 62.88 4.629 ;
      RECT 62.79 4.205 62.875 4.604 ;
      RECT 62.76 4.205 62.79 4.57 ;
      RECT 62.745 4.205 62.76 4.553 ;
      RECT 62.69 4.205 62.745 4.498 ;
      RECT 62.685 4.21 62.69 4.447 ;
      RECT 62.675 4.215 62.685 4.437 ;
      RECT 62.67 4.225 62.675 4.423 ;
      RECT 62.62 4.965 62.88 5.225 ;
      RECT 62.54 4.98 62.88 5.201 ;
      RECT 62.52 4.98 62.88 5.196 ;
      RECT 62.496 4.98 62.88 5.194 ;
      RECT 62.41 4.98 62.88 5.189 ;
      RECT 62.26 4.92 62.52 5.185 ;
      RECT 62.215 4.98 62.88 5.18 ;
      RECT 62.21 4.987 62.88 5.175 ;
      RECT 62.225 4.975 62.54 5.185 ;
      RECT 62.115 3.41 62.375 3.67 ;
      RECT 62.115 3.467 62.38 3.663 ;
      RECT 62.115 3.497 62.385 3.595 ;
      RECT 62.175 3.928 62.29 3.93 ;
      RECT 62.261 3.925 62.29 3.93 ;
      RECT 61.285 4.929 61.31 5.169 ;
      RECT 61.27 4.932 61.36 5.163 ;
      RECT 61.265 4.937 61.446 5.158 ;
      RECT 61.26 4.945 61.51 5.156 ;
      RECT 61.26 4.945 61.52 5.155 ;
      RECT 61.255 4.952 61.53 5.148 ;
      RECT 61.255 4.952 61.616 5.137 ;
      RECT 61.25 4.987 61.616 5.133 ;
      RECT 61.25 4.987 61.625 5.122 ;
      RECT 61.53 4.86 61.79 5.12 ;
      RECT 61.24 5.037 61.79 5.118 ;
      RECT 61.51 4.905 61.53 5.153 ;
      RECT 61.446 4.908 61.51 5.157 ;
      RECT 61.36 4.913 61.446 5.162 ;
      RECT 61.29 4.924 61.79 5.12 ;
      RECT 61.31 4.918 61.36 5.167 ;
      RECT 61.435 3.395 61.445 3.657 ;
      RECT 61.425 3.452 61.435 3.66 ;
      RECT 61.4 3.457 61.425 3.666 ;
      RECT 61.375 3.461 61.4 3.678 ;
      RECT 61.365 3.464 61.375 3.688 ;
      RECT 61.36 3.465 61.365 3.693 ;
      RECT 61.355 3.466 61.36 3.698 ;
      RECT 61.35 3.467 61.355 3.7 ;
      RECT 61.325 3.47 61.35 3.703 ;
      RECT 61.295 3.476 61.325 3.706 ;
      RECT 61.23 3.487 61.295 3.709 ;
      RECT 61.185 3.495 61.23 3.713 ;
      RECT 61.17 3.495 61.185 3.721 ;
      RECT 61.165 3.496 61.17 3.728 ;
      RECT 61.16 3.498 61.165 3.731 ;
      RECT 61.155 3.502 61.16 3.734 ;
      RECT 61.145 3.51 61.155 3.738 ;
      RECT 61.14 3.523 61.145 3.743 ;
      RECT 61.135 3.531 61.14 3.745 ;
      RECT 61.13 3.537 61.135 3.745 ;
      RECT 61.125 3.541 61.13 3.748 ;
      RECT 61.12 3.543 61.125 3.751 ;
      RECT 61.115 3.546 61.12 3.754 ;
      RECT 61.105 3.551 61.115 3.758 ;
      RECT 61.1 3.557 61.105 3.763 ;
      RECT 61.09 3.563 61.1 3.767 ;
      RECT 61.075 3.57 61.09 3.773 ;
      RECT 61.046 3.584 61.075 3.783 ;
      RECT 60.96 3.619 61.046 3.815 ;
      RECT 60.94 3.652 60.96 3.844 ;
      RECT 60.92 3.665 60.94 3.855 ;
      RECT 60.9 3.677 60.92 3.866 ;
      RECT 60.85 3.699 60.9 3.886 ;
      RECT 60.835 3.717 60.85 3.903 ;
      RECT 60.83 3.723 60.835 3.906 ;
      RECT 60.825 3.727 60.83 3.909 ;
      RECT 60.82 3.731 60.825 3.913 ;
      RECT 60.815 3.733 60.82 3.916 ;
      RECT 60.805 3.74 60.815 3.919 ;
      RECT 60.8 3.745 60.805 3.923 ;
      RECT 60.795 3.747 60.8 3.926 ;
      RECT 60.79 3.751 60.795 3.929 ;
      RECT 60.785 3.753 60.79 3.933 ;
      RECT 60.77 3.758 60.785 3.938 ;
      RECT 60.765 3.763 60.77 3.941 ;
      RECT 60.76 3.771 60.765 3.944 ;
      RECT 60.755 3.773 60.76 3.947 ;
      RECT 60.75 3.775 60.755 3.95 ;
      RECT 60.74 3.777 60.75 3.956 ;
      RECT 60.705 3.791 60.74 3.968 ;
      RECT 60.695 3.806 60.705 3.978 ;
      RECT 60.62 3.835 60.695 4.002 ;
      RECT 60.615 3.86 60.62 4.025 ;
      RECT 60.6 3.864 60.615 4.031 ;
      RECT 60.59 3.872 60.6 4.036 ;
      RECT 60.56 3.885 60.59 4.04 ;
      RECT 60.55 3.9 60.56 4.045 ;
      RECT 60.54 3.905 60.55 4.048 ;
      RECT 60.535 3.907 60.54 4.05 ;
      RECT 60.52 3.91 60.535 4.053 ;
      RECT 60.515 3.912 60.52 4.056 ;
      RECT 60.495 3.917 60.515 4.06 ;
      RECT 60.465 3.922 60.495 4.068 ;
      RECT 60.44 3.929 60.465 4.076 ;
      RECT 60.435 3.934 60.44 4.081 ;
      RECT 60.405 3.937 60.435 4.085 ;
      RECT 60.365 3.94 60.405 4.095 ;
      RECT 60.33 3.937 60.365 4.107 ;
      RECT 60.32 3.933 60.33 4.114 ;
      RECT 60.295 3.929 60.32 4.12 ;
      RECT 60.29 3.925 60.295 4.125 ;
      RECT 60.25 3.922 60.29 4.125 ;
      RECT 60.235 3.907 60.25 4.126 ;
      RECT 60.212 3.895 60.235 4.126 ;
      RECT 60.126 3.895 60.212 4.127 ;
      RECT 60.04 3.895 60.126 4.129 ;
      RECT 60.02 3.895 60.04 4.126 ;
      RECT 60.015 3.9 60.02 4.121 ;
      RECT 60.01 3.905 60.015 4.119 ;
      RECT 60 3.915 60.01 4.117 ;
      RECT 59.995 3.921 60 4.11 ;
      RECT 59.99 3.923 59.995 4.095 ;
      RECT 59.985 3.927 59.99 4.085 ;
      RECT 61.445 3.395 61.695 3.655 ;
      RECT 59.17 4.93 59.43 5.19 ;
      RECT 61.465 4.42 61.47 4.63 ;
      RECT 61.47 4.425 61.48 4.625 ;
      RECT 61.42 4.42 61.465 4.645 ;
      RECT 61.41 4.42 61.42 4.665 ;
      RECT 61.391 4.42 61.41 4.67 ;
      RECT 61.305 4.42 61.391 4.667 ;
      RECT 61.275 4.422 61.305 4.665 ;
      RECT 61.22 4.432 61.275 4.663 ;
      RECT 61.155 4.446 61.22 4.661 ;
      RECT 61.15 4.454 61.155 4.66 ;
      RECT 61.135 4.457 61.15 4.658 ;
      RECT 61.07 4.467 61.135 4.654 ;
      RECT 61.022 4.481 61.07 4.655 ;
      RECT 60.936 4.498 61.022 4.669 ;
      RECT 60.85 4.519 60.936 4.686 ;
      RECT 60.83 4.532 60.85 4.696 ;
      RECT 60.785 4.54 60.83 4.703 ;
      RECT 60.75 4.548 60.785 4.711 ;
      RECT 60.716 4.556 60.75 4.719 ;
      RECT 60.63 4.57 60.716 4.731 ;
      RECT 60.595 4.587 60.63 4.743 ;
      RECT 60.586 4.596 60.595 4.747 ;
      RECT 60.5 4.614 60.586 4.764 ;
      RECT 60.441 4.641 60.5 4.791 ;
      RECT 60.355 4.668 60.441 4.819 ;
      RECT 60.335 4.69 60.355 4.839 ;
      RECT 60.275 4.705 60.335 4.855 ;
      RECT 60.265 4.717 60.275 4.868 ;
      RECT 60.26 4.722 60.265 4.871 ;
      RECT 60.25 4.725 60.26 4.874 ;
      RECT 60.245 4.727 60.25 4.877 ;
      RECT 60.215 4.735 60.245 4.884 ;
      RECT 60.2 4.742 60.215 4.892 ;
      RECT 60.19 4.747 60.2 4.896 ;
      RECT 60.185 4.75 60.19 4.899 ;
      RECT 60.175 4.752 60.185 4.902 ;
      RECT 60.14 4.762 60.175 4.911 ;
      RECT 60.065 4.785 60.14 4.933 ;
      RECT 60.045 4.803 60.065 4.951 ;
      RECT 60.015 4.81 60.045 4.961 ;
      RECT 59.995 4.818 60.015 4.971 ;
      RECT 59.985 4.824 59.995 4.978 ;
      RECT 59.966 4.829 59.985 4.984 ;
      RECT 59.88 4.849 59.966 5.004 ;
      RECT 59.865 4.869 59.88 5.023 ;
      RECT 59.82 4.881 59.865 5.034 ;
      RECT 59.755 4.902 59.82 5.057 ;
      RECT 59.715 4.922 59.755 5.078 ;
      RECT 59.705 4.932 59.715 5.088 ;
      RECT 59.655 4.944 59.705 5.099 ;
      RECT 59.635 4.96 59.655 5.111 ;
      RECT 59.605 4.97 59.635 5.117 ;
      RECT 59.595 4.975 59.605 5.119 ;
      RECT 59.526 4.976 59.595 5.125 ;
      RECT 59.44 4.978 59.526 5.135 ;
      RECT 59.43 4.979 59.44 5.14 ;
      RECT 60.7 5.005 60.89 5.215 ;
      RECT 60.69 5.01 60.9 5.208 ;
      RECT 60.675 5.01 60.9 5.173 ;
      RECT 60.595 4.895 60.855 5.155 ;
      RECT 59.51 4.425 59.695 4.72 ;
      RECT 59.5 4.425 59.695 4.718 ;
      RECT 59.485 4.425 59.7 4.713 ;
      RECT 59.485 4.425 59.705 4.71 ;
      RECT 59.48 4.425 59.705 4.708 ;
      RECT 59.475 4.68 59.705 4.698 ;
      RECT 59.48 4.425 59.74 4.685 ;
      RECT 59.44 3.46 59.7 3.72 ;
      RECT 59.25 3.385 59.336 3.718 ;
      RECT 59.225 3.389 59.38 3.714 ;
      RECT 59.336 3.381 59.38 3.714 ;
      RECT 59.336 3.382 59.385 3.713 ;
      RECT 59.25 3.387 59.4 3.712 ;
      RECT 59.225 3.395 59.44 3.711 ;
      RECT 59.22 3.39 59.4 3.706 ;
      RECT 59.21 3.405 59.44 3.613 ;
      RECT 59.21 3.457 59.64 3.613 ;
      RECT 59.21 3.45 59.62 3.613 ;
      RECT 59.21 3.437 59.59 3.613 ;
      RECT 59.21 3.425 59.53 3.613 ;
      RECT 59.21 3.41 59.505 3.613 ;
      RECT 58.41 4.04 58.545 4.335 ;
      RECT 58.67 4.063 58.675 4.25 ;
      RECT 59.39 3.96 59.535 4.195 ;
      RECT 59.55 3.96 59.555 4.185 ;
      RECT 59.585 3.971 59.59 4.165 ;
      RECT 59.58 3.963 59.585 4.17 ;
      RECT 59.56 3.96 59.58 4.175 ;
      RECT 59.555 3.96 59.56 4.183 ;
      RECT 59.545 3.96 59.55 4.188 ;
      RECT 59.535 3.96 59.545 4.193 ;
      RECT 59.365 3.962 59.39 4.195 ;
      RECT 59.315 3.969 59.365 4.195 ;
      RECT 59.31 3.974 59.315 4.195 ;
      RECT 59.271 3.979 59.31 4.196 ;
      RECT 59.185 3.991 59.271 4.197 ;
      RECT 59.176 4.001 59.185 4.197 ;
      RECT 59.09 4.01 59.176 4.199 ;
      RECT 59.066 4.02 59.09 4.201 ;
      RECT 58.98 4.031 59.066 4.202 ;
      RECT 58.95 4.042 58.98 4.204 ;
      RECT 58.92 4.047 58.95 4.206 ;
      RECT 58.895 4.053 58.92 4.209 ;
      RECT 58.88 4.058 58.895 4.21 ;
      RECT 58.835 4.064 58.88 4.21 ;
      RECT 58.83 4.069 58.835 4.211 ;
      RECT 58.81 4.069 58.83 4.213 ;
      RECT 58.79 4.067 58.81 4.218 ;
      RECT 58.755 4.066 58.79 4.225 ;
      RECT 58.725 4.065 58.755 4.235 ;
      RECT 58.675 4.064 58.725 4.245 ;
      RECT 58.585 4.061 58.67 4.335 ;
      RECT 58.56 4.055 58.585 4.335 ;
      RECT 58.545 4.045 58.56 4.335 ;
      RECT 58.36 4.04 58.41 4.255 ;
      RECT 58.35 4.045 58.36 4.245 ;
      RECT 58.59 4.52 58.85 4.78 ;
      RECT 58.59 4.52 58.88 4.673 ;
      RECT 58.59 4.52 58.915 4.658 ;
      RECT 58.845 4.44 59.035 4.65 ;
      RECT 58.835 4.445 59.045 4.643 ;
      RECT 58.8 4.515 59.045 4.643 ;
      RECT 58.83 4.457 58.85 4.78 ;
      RECT 58.815 4.505 59.045 4.643 ;
      RECT 58.82 4.477 58.85 4.78 ;
      RECT 57.9 3.545 57.97 4.65 ;
      RECT 58.635 3.65 58.895 3.91 ;
      RECT 58.215 3.696 58.23 3.905 ;
      RECT 58.551 3.709 58.635 3.86 ;
      RECT 58.465 3.706 58.551 3.86 ;
      RECT 58.426 3.704 58.465 3.86 ;
      RECT 58.34 3.702 58.426 3.86 ;
      RECT 58.28 3.7 58.34 3.871 ;
      RECT 58.245 3.698 58.28 3.889 ;
      RECT 58.23 3.696 58.245 3.9 ;
      RECT 58.2 3.696 58.215 3.913 ;
      RECT 58.19 3.696 58.2 3.918 ;
      RECT 58.165 3.695 58.19 3.923 ;
      RECT 58.15 3.69 58.165 3.929 ;
      RECT 58.145 3.683 58.15 3.934 ;
      RECT 58.12 3.674 58.145 3.94 ;
      RECT 58.075 3.653 58.12 3.953 ;
      RECT 58.065 3.637 58.075 3.963 ;
      RECT 58.05 3.63 58.065 3.973 ;
      RECT 58.04 3.623 58.05 3.99 ;
      RECT 58.035 3.62 58.04 4.02 ;
      RECT 58.03 3.618 58.035 4.05 ;
      RECT 58.025 3.616 58.03 4.087 ;
      RECT 58.01 3.612 58.025 4.154 ;
      RECT 58.01 4.445 58.02 4.645 ;
      RECT 58.005 3.608 58.01 4.28 ;
      RECT 58.005 4.432 58.01 4.65 ;
      RECT 58 3.606 58.005 4.365 ;
      RECT 58 4.422 58.005 4.65 ;
      RECT 57.985 3.577 58 4.65 ;
      RECT 57.97 3.55 57.985 4.65 ;
      RECT 57.895 3.545 57.9 3.9 ;
      RECT 57.895 3.955 57.9 4.65 ;
      RECT 57.88 3.545 57.895 3.878 ;
      RECT 57.89 3.977 57.895 4.65 ;
      RECT 57.88 4.017 57.89 4.65 ;
      RECT 57.845 3.545 57.88 3.82 ;
      RECT 57.875 4.052 57.88 4.65 ;
      RECT 57.86 4.107 57.875 4.65 ;
      RECT 57.855 4.172 57.86 4.65 ;
      RECT 57.84 4.22 57.855 4.65 ;
      RECT 57.815 3.545 57.845 3.775 ;
      RECT 57.835 4.275 57.84 4.65 ;
      RECT 57.82 4.335 57.835 4.65 ;
      RECT 57.815 4.383 57.82 4.648 ;
      RECT 57.81 3.545 57.815 3.768 ;
      RECT 57.81 4.415 57.815 4.643 ;
      RECT 57.785 3.545 57.81 3.76 ;
      RECT 57.775 3.55 57.785 3.75 ;
      RECT 57.99 4.825 58.01 5.065 ;
      RECT 57.22 4.755 57.225 4.965 ;
      RECT 58.5 4.828 58.51 5.023 ;
      RECT 58.495 4.818 58.5 5.026 ;
      RECT 58.415 4.815 58.495 5.049 ;
      RECT 58.411 4.815 58.415 5.071 ;
      RECT 58.325 4.815 58.411 5.081 ;
      RECT 58.31 4.815 58.325 5.089 ;
      RECT 58.281 4.816 58.31 5.087 ;
      RECT 58.195 4.821 58.281 5.083 ;
      RECT 58.182 4.825 58.195 5.079 ;
      RECT 58.096 4.825 58.182 5.075 ;
      RECT 58.01 4.825 58.096 5.069 ;
      RECT 57.926 4.825 57.99 5.063 ;
      RECT 57.84 4.825 57.926 5.058 ;
      RECT 57.82 4.825 57.84 5.054 ;
      RECT 57.76 4.82 57.82 5.051 ;
      RECT 57.732 4.814 57.76 5.048 ;
      RECT 57.646 4.809 57.732 5.044 ;
      RECT 57.56 4.803 57.646 5.038 ;
      RECT 57.485 4.785 57.56 5.033 ;
      RECT 57.45 4.762 57.485 5.029 ;
      RECT 57.44 4.752 57.45 5.028 ;
      RECT 57.385 4.75 57.44 5.027 ;
      RECT 57.31 4.75 57.385 5.023 ;
      RECT 57.3 4.75 57.31 5.018 ;
      RECT 57.285 4.75 57.3 5.01 ;
      RECT 57.235 4.752 57.285 4.988 ;
      RECT 57.225 4.755 57.235 4.968 ;
      RECT 57.215 4.76 57.22 4.963 ;
      RECT 57.21 4.765 57.215 4.958 ;
      RECT 55.32 3.41 55.58 3.67 ;
      RECT 55.31 3.44 55.58 3.65 ;
      RECT 57.23 3.355 57.49 3.615 ;
      RECT 57.225 3.43 57.23 3.616 ;
      RECT 57.2 3.435 57.225 3.618 ;
      RECT 57.185 3.442 57.2 3.621 ;
      RECT 57.125 3.46 57.185 3.626 ;
      RECT 57.095 3.48 57.125 3.633 ;
      RECT 57.07 3.488 57.095 3.638 ;
      RECT 57.045 3.496 57.07 3.64 ;
      RECT 57.027 3.5 57.045 3.639 ;
      RECT 56.941 3.498 57.027 3.639 ;
      RECT 56.855 3.496 56.941 3.639 ;
      RECT 56.769 3.494 56.855 3.638 ;
      RECT 56.683 3.492 56.769 3.638 ;
      RECT 56.597 3.49 56.683 3.638 ;
      RECT 56.511 3.488 56.597 3.638 ;
      RECT 56.425 3.486 56.511 3.637 ;
      RECT 56.407 3.485 56.425 3.637 ;
      RECT 56.321 3.484 56.407 3.637 ;
      RECT 56.235 3.482 56.321 3.637 ;
      RECT 56.149 3.481 56.235 3.636 ;
      RECT 56.063 3.48 56.149 3.636 ;
      RECT 55.977 3.478 56.063 3.636 ;
      RECT 55.891 3.477 55.977 3.636 ;
      RECT 55.805 3.475 55.891 3.635 ;
      RECT 55.781 3.473 55.805 3.635 ;
      RECT 55.695 3.466 55.781 3.635 ;
      RECT 55.666 3.458 55.695 3.635 ;
      RECT 55.58 3.45 55.666 3.635 ;
      RECT 55.3 3.447 55.31 3.645 ;
      RECT 56.805 4.41 56.81 4.76 ;
      RECT 56.575 4.5 56.715 4.76 ;
      RECT 57.05 4.185 57.095 4.395 ;
      RECT 57.105 4.196 57.115 4.39 ;
      RECT 57.095 4.188 57.105 4.395 ;
      RECT 57.03 4.185 57.05 4.4 ;
      RECT 57 4.185 57.03 4.423 ;
      RECT 56.99 4.185 57 4.448 ;
      RECT 56.985 4.185 56.99 4.458 ;
      RECT 56.93 4.185 56.985 4.498 ;
      RECT 56.925 4.185 56.93 4.538 ;
      RECT 56.92 4.187 56.925 4.543 ;
      RECT 56.905 4.197 56.92 4.554 ;
      RECT 56.86 4.255 56.905 4.59 ;
      RECT 56.85 4.31 56.86 4.624 ;
      RECT 56.835 4.337 56.85 4.64 ;
      RECT 56.825 4.364 56.835 4.76 ;
      RECT 56.81 4.387 56.825 4.76 ;
      RECT 56.8 4.427 56.805 4.76 ;
      RECT 56.795 4.437 56.8 4.76 ;
      RECT 56.79 4.452 56.795 4.76 ;
      RECT 56.78 4.457 56.79 4.76 ;
      RECT 56.715 4.48 56.78 4.76 ;
      RECT 56.185 3.975 56.405 4.185 ;
      RECT 56.185 3.982 56.415 4.18 ;
      RECT 55.49 3.99 56.415 4.165 ;
      RECT 56.01 3.885 56.4 4.165 ;
      RECT 54.79 3.9 55.05 4.16 ;
      RECT 55.425 3.935 55.56 4.12 ;
      RECT 55.35 3.925 55.445 4.115 ;
      RECT 55.34 3.99 56.415 4.111 ;
      RECT 55.09 3.99 56.415 4.11 ;
      RECT 55.115 3.91 55.355 4.11 ;
      RECT 54.79 3.915 55.375 4.098 ;
      RECT 56.705 3.94 56.745 4.025 ;
      RECT 54.79 3.975 55.965 4.098 ;
      RECT 54.79 3.965 55.85 4.098 ;
      RECT 54.79 3.946 55.755 4.098 ;
      RECT 55.575 3.94 55.755 4.165 ;
      RECT 56.01 3.92 56.705 3.955 ;
      RECT 55.11 3.912 55.355 4.11 ;
      RECT 55.125 3.902 55.335 4.11 ;
      RECT 55.14 3.895 55.335 4.11 ;
      RECT 55.305 4.415 55.565 4.675 ;
      RECT 55.305 4.455 55.67 4.665 ;
      RECT 55.305 4.457 55.675 4.664 ;
      RECT 55.305 4.465 55.68 4.661 ;
      RECT 54.23 3.54 54.33 5.065 ;
      RECT 54.42 4.68 54.47 4.94 ;
      RECT 54.415 3.553 54.42 3.74 ;
      RECT 54.41 4.661 54.42 4.94 ;
      RECT 54.41 3.55 54.415 3.748 ;
      RECT 54.395 3.544 54.41 3.755 ;
      RECT 54.405 4.649 54.41 5.023 ;
      RECT 54.395 4.637 54.405 5.06 ;
      RECT 54.385 3.54 54.395 3.762 ;
      RECT 54.385 4.622 54.395 5.065 ;
      RECT 54.38 3.54 54.385 3.77 ;
      RECT 54.36 4.592 54.385 5.065 ;
      RECT 54.34 3.54 54.38 3.818 ;
      RECT 54.35 4.552 54.36 5.065 ;
      RECT 54.34 4.507 54.35 5.065 ;
      RECT 54.335 3.54 54.34 3.888 ;
      RECT 54.335 4.465 54.34 5.065 ;
      RECT 54.33 3.54 54.335 4.365 ;
      RECT 54.33 4.447 54.335 5.065 ;
      RECT 54.22 3.543 54.23 5.065 ;
      RECT 54.205 3.55 54.22 5.061 ;
      RECT 54.2 3.56 54.205 5.056 ;
      RECT 54.195 3.76 54.2 4.948 ;
      RECT 54.19 3.845 54.195 4.5 ;
      RECT 53.055 10.205 53.35 10.435 ;
      RECT 53.115 8.725 53.285 10.435 ;
      RECT 53.105 9.095 53.46 9.45 ;
      RECT 53.055 8.725 53.345 8.955 ;
      RECT 52.065 10.205 52.36 10.435 ;
      RECT 52.125 8.725 52.295 10.435 ;
      RECT 52.065 8.725 52.355 8.955 ;
      RECT 52.065 8.76 52.915 8.92 ;
      RECT 52.75 8.355 52.915 8.92 ;
      RECT 52.065 8.755 52.46 8.92 ;
      RECT 52.685 8.355 52.975 8.585 ;
      RECT 52.685 8.385 53.145 8.555 ;
      RECT 52.65 4.025 52.97 4.26 ;
      RECT 52.65 4.055 53.14 4.225 ;
      RECT 52.65 3.69 52.84 4.26 ;
      RECT 52.065 3.655 52.355 3.885 ;
      RECT 52.065 3.69 52.84 3.86 ;
      RECT 52.125 2.175 52.295 3.885 ;
      RECT 52.065 2.175 52.36 2.405 ;
      RECT 51.695 4.025 51.985 4.255 ;
      RECT 51.695 4.055 52.155 4.225 ;
      RECT 51.76 2.95 51.925 4.255 ;
      RECT 50.275 2.915 50.565 3.145 ;
      RECT 50.275 2.95 51.925 3.12 ;
      RECT 50.335 2.175 50.505 3.145 ;
      RECT 50.275 2.175 50.565 2.405 ;
      RECT 50.275 10.205 50.565 10.435 ;
      RECT 50.335 9.465 50.505 10.435 ;
      RECT 50.335 9.555 51.925 9.725 ;
      RECT 51.755 8.355 51.925 9.725 ;
      RECT 50.275 9.465 50.565 9.695 ;
      RECT 51.695 8.355 51.985 8.585 ;
      RECT 51.695 8.385 52.155 8.555 ;
      RECT 48.31 4.725 48.66 5.075 ;
      RECT 48.4 3.32 48.57 5.075 ;
      RECT 50.705 3.26 51.055 3.61 ;
      RECT 48.4 3.32 50.02 3.495 ;
      RECT 48.4 3.32 50.675 3.49 ;
      RECT 50.535 3.315 51.055 3.485 ;
      RECT 50.73 9.09 51.055 9.415 ;
      RECT 46.155 9.05 46.505 9.4 ;
      RECT 50.705 9.095 51.055 9.325 ;
      RECT 45.945 9.095 46.505 9.325 ;
      RECT 50.535 9.12 51.055 9.295 ;
      RECT 45.775 9.125 46.505 9.295 ;
      RECT 45.945 9.12 51.055 9.29 ;
      RECT 49.93 3.66 50.25 3.98 ;
      RECT 49.905 3.655 50.195 3.885 ;
      RECT 49.86 3.685 50.25 3.86 ;
      RECT 49.73 3.685 50.25 3.855 ;
      RECT 49.93 8.66 50.25 8.98 ;
      RECT 49.905 8.725 50.25 8.955 ;
      RECT 49.73 8.755 50.25 8.925 ;
      RECT 45.72 4.96 45.76 5.22 ;
      RECT 45.76 4.94 45.765 4.95 ;
      RECT 47.09 4.185 47.1 4.406 ;
      RECT 47.02 4.18 47.09 4.531 ;
      RECT 47.01 4.18 47.02 4.658 ;
      RECT 46.985 4.18 47.01 4.705 ;
      RECT 46.96 4.18 46.985 4.783 ;
      RECT 46.94 4.18 46.96 4.853 ;
      RECT 46.915 4.18 46.94 4.893 ;
      RECT 46.905 4.18 46.915 4.913 ;
      RECT 46.895 4.182 46.905 4.921 ;
      RECT 46.89 4.187 46.895 4.378 ;
      RECT 46.89 4.387 46.895 4.922 ;
      RECT 46.885 4.432 46.89 4.923 ;
      RECT 46.875 4.497 46.885 4.924 ;
      RECT 46.865 4.592 46.875 4.926 ;
      RECT 46.86 4.645 46.865 4.928 ;
      RECT 46.855 4.665 46.86 4.929 ;
      RECT 46.8 4.69 46.855 4.935 ;
      RECT 46.76 4.725 46.8 4.944 ;
      RECT 46.75 4.742 46.76 4.949 ;
      RECT 46.741 4.748 46.75 4.951 ;
      RECT 46.655 4.786 46.741 4.962 ;
      RECT 46.65 4.825 46.655 4.972 ;
      RECT 46.575 4.832 46.65 4.982 ;
      RECT 46.555 4.842 46.575 4.993 ;
      RECT 46.525 4.849 46.555 5.001 ;
      RECT 46.5 4.856 46.525 5.008 ;
      RECT 46.476 4.862 46.5 5.013 ;
      RECT 46.39 4.875 46.476 5.025 ;
      RECT 46.312 4.882 46.39 5.043 ;
      RECT 46.226 4.877 46.312 5.061 ;
      RECT 46.14 4.872 46.226 5.081 ;
      RECT 46.06 4.866 46.14 5.098 ;
      RECT 45.995 4.862 46.06 5.127 ;
      RECT 45.99 4.576 45.995 4.6 ;
      RECT 45.98 4.852 45.995 5.155 ;
      RECT 45.985 4.57 45.99 4.64 ;
      RECT 45.98 4.564 45.985 4.71 ;
      RECT 45.975 4.558 45.98 4.788 ;
      RECT 45.975 4.835 45.98 5.22 ;
      RECT 45.967 4.555 45.975 5.22 ;
      RECT 45.881 4.553 45.967 5.22 ;
      RECT 45.795 4.551 45.881 5.22 ;
      RECT 45.785 4.552 45.795 5.22 ;
      RECT 45.78 4.557 45.785 5.22 ;
      RECT 45.77 4.57 45.78 5.22 ;
      RECT 45.765 4.592 45.77 5.22 ;
      RECT 45.76 4.952 45.765 5.22 ;
      RECT 46.39 4.42 46.395 4.64 ;
      RECT 46.895 3.455 46.93 3.715 ;
      RECT 46.88 3.455 46.895 3.723 ;
      RECT 46.851 3.455 46.88 3.745 ;
      RECT 46.765 3.455 46.851 3.805 ;
      RECT 46.745 3.455 46.765 3.87 ;
      RECT 46.685 3.455 46.745 4.035 ;
      RECT 46.68 3.455 46.685 4.183 ;
      RECT 46.675 3.455 46.68 4.195 ;
      RECT 46.67 3.455 46.675 4.221 ;
      RECT 46.64 3.641 46.67 4.301 ;
      RECT 46.635 3.689 46.64 4.39 ;
      RECT 46.63 3.703 46.635 4.405 ;
      RECT 46.625 3.722 46.63 4.435 ;
      RECT 46.62 3.737 46.625 4.451 ;
      RECT 46.615 3.752 46.62 4.473 ;
      RECT 46.61 3.772 46.615 4.495 ;
      RECT 46.6 3.792 46.61 4.528 ;
      RECT 46.585 3.834 46.6 4.59 ;
      RECT 46.58 3.865 46.585 4.63 ;
      RECT 46.575 3.877 46.58 4.635 ;
      RECT 46.57 3.889 46.575 4.64 ;
      RECT 46.565 3.902 46.57 4.64 ;
      RECT 46.56 3.92 46.565 4.64 ;
      RECT 46.555 3.94 46.56 4.64 ;
      RECT 46.55 3.952 46.555 4.64 ;
      RECT 46.545 3.965 46.55 4.64 ;
      RECT 46.525 4 46.545 4.64 ;
      RECT 46.475 4.102 46.525 4.64 ;
      RECT 46.47 4.187 46.475 4.64 ;
      RECT 46.465 4.195 46.47 4.64 ;
      RECT 46.46 4.212 46.465 4.64 ;
      RECT 46.455 4.227 46.46 4.64 ;
      RECT 46.42 4.292 46.455 4.64 ;
      RECT 46.405 4.357 46.42 4.64 ;
      RECT 46.4 4.387 46.405 4.64 ;
      RECT 46.395 4.412 46.4 4.64 ;
      RECT 46.38 4.422 46.39 4.64 ;
      RECT 46.365 4.435 46.38 4.633 ;
      RECT 46.11 4.025 46.18 4.235 ;
      RECT 45.9 4.002 45.905 4.195 ;
      RECT 43.355 3.93 43.615 4.19 ;
      RECT 46.19 4.212 46.195 4.215 ;
      RECT 46.18 4.03 46.19 4.23 ;
      RECT 46.081 4.023 46.11 4.235 ;
      RECT 45.995 4.015 46.081 4.235 ;
      RECT 45.98 4.009 45.995 4.233 ;
      RECT 45.96 4.008 45.98 4.22 ;
      RECT 45.955 4.007 45.96 4.203 ;
      RECT 45.905 4.004 45.955 4.198 ;
      RECT 45.875 4.001 45.9 4.193 ;
      RECT 45.855 3.999 45.875 4.188 ;
      RECT 45.84 3.997 45.855 4.185 ;
      RECT 45.81 3.995 45.84 4.183 ;
      RECT 45.745 3.991 45.81 4.175 ;
      RECT 45.715 3.986 45.745 4.17 ;
      RECT 45.695 3.984 45.715 4.168 ;
      RECT 45.665 3.981 45.695 4.163 ;
      RECT 45.605 3.977 45.665 4.155 ;
      RECT 45.6 3.974 45.605 4.15 ;
      RECT 45.53 3.972 45.6 4.145 ;
      RECT 45.501 3.968 45.53 4.138 ;
      RECT 45.415 3.963 45.501 4.13 ;
      RECT 45.381 3.958 45.415 4.122 ;
      RECT 45.295 3.95 45.381 4.114 ;
      RECT 45.256 3.943 45.295 4.106 ;
      RECT 45.17 3.938 45.256 4.098 ;
      RECT 45.105 3.932 45.17 4.088 ;
      RECT 45.085 3.927 45.105 4.083 ;
      RECT 45.076 3.924 45.085 4.082 ;
      RECT 44.99 3.92 45.076 4.076 ;
      RECT 44.95 3.916 44.99 4.068 ;
      RECT 44.93 3.912 44.95 4.066 ;
      RECT 44.87 3.912 44.93 4.063 ;
      RECT 44.85 3.915 44.87 4.061 ;
      RECT 44.829 3.915 44.85 4.061 ;
      RECT 44.743 3.917 44.829 4.065 ;
      RECT 44.657 3.919 44.743 4.071 ;
      RECT 44.571 3.921 44.657 4.078 ;
      RECT 44.485 3.924 44.571 4.084 ;
      RECT 44.451 3.925 44.485 4.089 ;
      RECT 44.365 3.928 44.451 4.094 ;
      RECT 44.336 3.935 44.365 4.099 ;
      RECT 44.25 3.935 44.336 4.104 ;
      RECT 44.217 3.935 44.25 4.109 ;
      RECT 44.131 3.937 44.217 4.114 ;
      RECT 44.045 3.939 44.131 4.121 ;
      RECT 43.981 3.941 44.045 4.127 ;
      RECT 43.895 3.943 43.981 4.133 ;
      RECT 43.892 3.945 43.895 4.136 ;
      RECT 43.806 3.946 43.892 4.14 ;
      RECT 43.72 3.949 43.806 4.147 ;
      RECT 43.701 3.951 43.72 4.151 ;
      RECT 43.615 3.953 43.701 4.156 ;
      RECT 43.345 3.965 43.355 4.16 ;
      RECT 45.515 10.205 45.805 10.435 ;
      RECT 45.575 9.465 45.745 10.435 ;
      RECT 45.465 9.49 45.84 9.86 ;
      RECT 45.515 9.465 45.805 9.86 ;
      RECT 45.58 3.545 45.765 3.755 ;
      RECT 45.575 3.546 45.77 3.753 ;
      RECT 45.57 3.551 45.78 3.748 ;
      RECT 45.565 3.527 45.57 3.745 ;
      RECT 45.535 3.524 45.565 3.738 ;
      RECT 45.53 3.52 45.535 3.729 ;
      RECT 45.495 3.551 45.78 3.724 ;
      RECT 45.27 3.46 45.53 3.72 ;
      RECT 45.57 3.529 45.575 3.748 ;
      RECT 45.575 3.53 45.58 3.753 ;
      RECT 45.27 3.542 45.65 3.72 ;
      RECT 45.27 3.54 45.635 3.72 ;
      RECT 45.27 3.535 45.625 3.72 ;
      RECT 45.225 4.45 45.275 4.735 ;
      RECT 45.17 4.42 45.175 4.735 ;
      RECT 45.14 4.4 45.145 4.735 ;
      RECT 45.29 4.45 45.35 4.71 ;
      RECT 45.285 4.45 45.29 4.718 ;
      RECT 45.275 4.45 45.285 4.73 ;
      RECT 45.19 4.44 45.225 4.735 ;
      RECT 45.185 4.427 45.19 4.735 ;
      RECT 45.175 4.422 45.185 4.735 ;
      RECT 45.155 4.412 45.17 4.735 ;
      RECT 45.145 4.405 45.155 4.735 ;
      RECT 45.135 4.397 45.14 4.735 ;
      RECT 45.105 4.387 45.135 4.735 ;
      RECT 45.09 4.375 45.105 4.735 ;
      RECT 45.075 4.365 45.09 4.73 ;
      RECT 45.055 4.355 45.075 4.705 ;
      RECT 45.045 4.347 45.055 4.682 ;
      RECT 45.015 4.33 45.045 4.672 ;
      RECT 45.01 4.307 45.015 4.663 ;
      RECT 45.005 4.294 45.01 4.661 ;
      RECT 44.99 4.27 45.005 4.655 ;
      RECT 44.985 4.246 44.99 4.649 ;
      RECT 44.975 4.235 44.985 4.644 ;
      RECT 44.97 4.225 44.975 4.64 ;
      RECT 44.965 4.217 44.97 4.637 ;
      RECT 44.955 4.212 44.965 4.633 ;
      RECT 44.95 4.207 44.955 4.629 ;
      RECT 44.865 4.205 44.95 4.604 ;
      RECT 44.835 4.205 44.865 4.57 ;
      RECT 44.82 4.205 44.835 4.553 ;
      RECT 44.765 4.205 44.82 4.498 ;
      RECT 44.76 4.21 44.765 4.447 ;
      RECT 44.75 4.215 44.76 4.437 ;
      RECT 44.745 4.225 44.75 4.423 ;
      RECT 44.695 4.965 44.955 5.225 ;
      RECT 44.615 4.98 44.955 5.201 ;
      RECT 44.595 4.98 44.955 5.196 ;
      RECT 44.571 4.98 44.955 5.194 ;
      RECT 44.485 4.98 44.955 5.189 ;
      RECT 44.335 4.92 44.595 5.185 ;
      RECT 44.29 4.98 44.955 5.18 ;
      RECT 44.285 4.987 44.955 5.175 ;
      RECT 44.3 4.975 44.615 5.185 ;
      RECT 44.19 3.41 44.45 3.67 ;
      RECT 44.19 3.467 44.455 3.663 ;
      RECT 44.19 3.497 44.46 3.595 ;
      RECT 44.25 3.928 44.365 3.93 ;
      RECT 44.336 3.925 44.365 3.93 ;
      RECT 43.36 4.929 43.385 5.169 ;
      RECT 43.345 4.932 43.435 5.163 ;
      RECT 43.34 4.937 43.521 5.158 ;
      RECT 43.335 4.945 43.585 5.156 ;
      RECT 43.335 4.945 43.595 5.155 ;
      RECT 43.33 4.952 43.605 5.148 ;
      RECT 43.33 4.952 43.691 5.137 ;
      RECT 43.325 4.987 43.691 5.133 ;
      RECT 43.325 4.987 43.7 5.122 ;
      RECT 43.605 4.86 43.865 5.12 ;
      RECT 43.315 5.037 43.865 5.118 ;
      RECT 43.585 4.905 43.605 5.153 ;
      RECT 43.521 4.908 43.585 5.157 ;
      RECT 43.435 4.913 43.521 5.162 ;
      RECT 43.365 4.924 43.865 5.12 ;
      RECT 43.385 4.918 43.435 5.167 ;
      RECT 43.51 3.395 43.52 3.657 ;
      RECT 43.5 3.452 43.51 3.66 ;
      RECT 43.475 3.457 43.5 3.666 ;
      RECT 43.45 3.461 43.475 3.678 ;
      RECT 43.44 3.464 43.45 3.688 ;
      RECT 43.435 3.465 43.44 3.693 ;
      RECT 43.43 3.466 43.435 3.698 ;
      RECT 43.425 3.467 43.43 3.7 ;
      RECT 43.4 3.47 43.425 3.703 ;
      RECT 43.37 3.476 43.4 3.706 ;
      RECT 43.305 3.487 43.37 3.709 ;
      RECT 43.26 3.495 43.305 3.713 ;
      RECT 43.245 3.495 43.26 3.721 ;
      RECT 43.24 3.496 43.245 3.728 ;
      RECT 43.235 3.498 43.24 3.731 ;
      RECT 43.23 3.502 43.235 3.734 ;
      RECT 43.22 3.51 43.23 3.738 ;
      RECT 43.215 3.523 43.22 3.743 ;
      RECT 43.21 3.531 43.215 3.745 ;
      RECT 43.205 3.537 43.21 3.745 ;
      RECT 43.2 3.541 43.205 3.748 ;
      RECT 43.195 3.543 43.2 3.751 ;
      RECT 43.19 3.546 43.195 3.754 ;
      RECT 43.18 3.551 43.19 3.758 ;
      RECT 43.175 3.557 43.18 3.763 ;
      RECT 43.165 3.563 43.175 3.767 ;
      RECT 43.15 3.57 43.165 3.773 ;
      RECT 43.121 3.584 43.15 3.783 ;
      RECT 43.035 3.619 43.121 3.815 ;
      RECT 43.015 3.652 43.035 3.844 ;
      RECT 42.995 3.665 43.015 3.855 ;
      RECT 42.975 3.677 42.995 3.866 ;
      RECT 42.925 3.699 42.975 3.886 ;
      RECT 42.91 3.717 42.925 3.903 ;
      RECT 42.905 3.723 42.91 3.906 ;
      RECT 42.9 3.727 42.905 3.909 ;
      RECT 42.895 3.731 42.9 3.913 ;
      RECT 42.89 3.733 42.895 3.916 ;
      RECT 42.88 3.74 42.89 3.919 ;
      RECT 42.875 3.745 42.88 3.923 ;
      RECT 42.87 3.747 42.875 3.926 ;
      RECT 42.865 3.751 42.87 3.929 ;
      RECT 42.86 3.753 42.865 3.933 ;
      RECT 42.845 3.758 42.86 3.938 ;
      RECT 42.84 3.763 42.845 3.941 ;
      RECT 42.835 3.771 42.84 3.944 ;
      RECT 42.83 3.773 42.835 3.947 ;
      RECT 42.825 3.775 42.83 3.95 ;
      RECT 42.815 3.777 42.825 3.956 ;
      RECT 42.78 3.791 42.815 3.968 ;
      RECT 42.77 3.806 42.78 3.978 ;
      RECT 42.695 3.835 42.77 4.002 ;
      RECT 42.69 3.86 42.695 4.025 ;
      RECT 42.675 3.864 42.69 4.031 ;
      RECT 42.665 3.872 42.675 4.036 ;
      RECT 42.635 3.885 42.665 4.04 ;
      RECT 42.625 3.9 42.635 4.045 ;
      RECT 42.615 3.905 42.625 4.048 ;
      RECT 42.61 3.907 42.615 4.05 ;
      RECT 42.595 3.91 42.61 4.053 ;
      RECT 42.59 3.912 42.595 4.056 ;
      RECT 42.57 3.917 42.59 4.06 ;
      RECT 42.54 3.922 42.57 4.068 ;
      RECT 42.515 3.929 42.54 4.076 ;
      RECT 42.51 3.934 42.515 4.081 ;
      RECT 42.48 3.937 42.51 4.085 ;
      RECT 42.44 3.94 42.48 4.095 ;
      RECT 42.405 3.937 42.44 4.107 ;
      RECT 42.395 3.933 42.405 4.114 ;
      RECT 42.37 3.929 42.395 4.12 ;
      RECT 42.365 3.925 42.37 4.125 ;
      RECT 42.325 3.922 42.365 4.125 ;
      RECT 42.31 3.907 42.325 4.126 ;
      RECT 42.287 3.895 42.31 4.126 ;
      RECT 42.201 3.895 42.287 4.127 ;
      RECT 42.115 3.895 42.201 4.129 ;
      RECT 42.095 3.895 42.115 4.126 ;
      RECT 42.09 3.9 42.095 4.121 ;
      RECT 42.085 3.905 42.09 4.119 ;
      RECT 42.075 3.915 42.085 4.117 ;
      RECT 42.07 3.921 42.075 4.11 ;
      RECT 42.065 3.923 42.07 4.095 ;
      RECT 42.06 3.927 42.065 4.085 ;
      RECT 43.52 3.395 43.77 3.655 ;
      RECT 41.245 4.93 41.505 5.19 ;
      RECT 43.54 4.42 43.545 4.63 ;
      RECT 43.545 4.425 43.555 4.625 ;
      RECT 43.495 4.42 43.54 4.645 ;
      RECT 43.485 4.42 43.495 4.665 ;
      RECT 43.466 4.42 43.485 4.67 ;
      RECT 43.38 4.42 43.466 4.667 ;
      RECT 43.35 4.422 43.38 4.665 ;
      RECT 43.295 4.432 43.35 4.663 ;
      RECT 43.23 4.446 43.295 4.661 ;
      RECT 43.225 4.454 43.23 4.66 ;
      RECT 43.21 4.457 43.225 4.658 ;
      RECT 43.145 4.467 43.21 4.654 ;
      RECT 43.097 4.481 43.145 4.655 ;
      RECT 43.011 4.498 43.097 4.669 ;
      RECT 42.925 4.519 43.011 4.686 ;
      RECT 42.905 4.532 42.925 4.696 ;
      RECT 42.86 4.54 42.905 4.703 ;
      RECT 42.825 4.548 42.86 4.711 ;
      RECT 42.791 4.556 42.825 4.719 ;
      RECT 42.705 4.57 42.791 4.731 ;
      RECT 42.67 4.587 42.705 4.743 ;
      RECT 42.661 4.596 42.67 4.747 ;
      RECT 42.575 4.614 42.661 4.764 ;
      RECT 42.516 4.641 42.575 4.791 ;
      RECT 42.43 4.668 42.516 4.819 ;
      RECT 42.41 4.69 42.43 4.839 ;
      RECT 42.35 4.705 42.41 4.855 ;
      RECT 42.34 4.717 42.35 4.868 ;
      RECT 42.335 4.722 42.34 4.871 ;
      RECT 42.325 4.725 42.335 4.874 ;
      RECT 42.32 4.727 42.325 4.877 ;
      RECT 42.29 4.735 42.32 4.884 ;
      RECT 42.275 4.742 42.29 4.892 ;
      RECT 42.265 4.747 42.275 4.896 ;
      RECT 42.26 4.75 42.265 4.899 ;
      RECT 42.25 4.752 42.26 4.902 ;
      RECT 42.215 4.762 42.25 4.911 ;
      RECT 42.14 4.785 42.215 4.933 ;
      RECT 42.12 4.803 42.14 4.951 ;
      RECT 42.09 4.81 42.12 4.961 ;
      RECT 42.07 4.818 42.09 4.971 ;
      RECT 42.06 4.824 42.07 4.978 ;
      RECT 42.041 4.829 42.06 4.984 ;
      RECT 41.955 4.849 42.041 5.004 ;
      RECT 41.94 4.869 41.955 5.023 ;
      RECT 41.895 4.881 41.94 5.034 ;
      RECT 41.83 4.902 41.895 5.057 ;
      RECT 41.79 4.922 41.83 5.078 ;
      RECT 41.78 4.932 41.79 5.088 ;
      RECT 41.73 4.944 41.78 5.099 ;
      RECT 41.71 4.96 41.73 5.111 ;
      RECT 41.68 4.97 41.71 5.117 ;
      RECT 41.67 4.975 41.68 5.119 ;
      RECT 41.601 4.976 41.67 5.125 ;
      RECT 41.515 4.978 41.601 5.135 ;
      RECT 41.505 4.979 41.515 5.14 ;
      RECT 42.775 5.005 42.965 5.215 ;
      RECT 42.765 5.01 42.975 5.208 ;
      RECT 42.75 5.01 42.975 5.173 ;
      RECT 42.67 4.895 42.93 5.155 ;
      RECT 41.585 4.425 41.77 4.72 ;
      RECT 41.575 4.425 41.77 4.718 ;
      RECT 41.56 4.425 41.775 4.713 ;
      RECT 41.56 4.425 41.78 4.71 ;
      RECT 41.555 4.425 41.78 4.708 ;
      RECT 41.55 4.68 41.78 4.698 ;
      RECT 41.555 4.425 41.815 4.685 ;
      RECT 41.515 3.46 41.775 3.72 ;
      RECT 41.325 3.385 41.411 3.718 ;
      RECT 41.3 3.389 41.455 3.714 ;
      RECT 41.411 3.381 41.455 3.714 ;
      RECT 41.411 3.382 41.46 3.713 ;
      RECT 41.325 3.387 41.475 3.712 ;
      RECT 41.3 3.395 41.515 3.711 ;
      RECT 41.295 3.39 41.475 3.706 ;
      RECT 41.285 3.405 41.515 3.613 ;
      RECT 41.285 3.457 41.715 3.613 ;
      RECT 41.285 3.45 41.695 3.613 ;
      RECT 41.285 3.437 41.665 3.613 ;
      RECT 41.285 3.425 41.605 3.613 ;
      RECT 41.285 3.41 41.58 3.613 ;
      RECT 40.485 4.04 40.62 4.335 ;
      RECT 40.745 4.063 40.75 4.25 ;
      RECT 41.465 3.96 41.61 4.195 ;
      RECT 41.625 3.96 41.63 4.185 ;
      RECT 41.66 3.971 41.665 4.165 ;
      RECT 41.655 3.963 41.66 4.17 ;
      RECT 41.635 3.96 41.655 4.175 ;
      RECT 41.63 3.96 41.635 4.183 ;
      RECT 41.62 3.96 41.625 4.188 ;
      RECT 41.61 3.96 41.62 4.193 ;
      RECT 41.44 3.962 41.465 4.195 ;
      RECT 41.39 3.969 41.44 4.195 ;
      RECT 41.385 3.974 41.39 4.195 ;
      RECT 41.346 3.979 41.385 4.196 ;
      RECT 41.26 3.991 41.346 4.197 ;
      RECT 41.251 4.001 41.26 4.197 ;
      RECT 41.165 4.01 41.251 4.199 ;
      RECT 41.141 4.02 41.165 4.201 ;
      RECT 41.055 4.031 41.141 4.202 ;
      RECT 41.025 4.042 41.055 4.204 ;
      RECT 40.995 4.047 41.025 4.206 ;
      RECT 40.97 4.053 40.995 4.209 ;
      RECT 40.955 4.058 40.97 4.21 ;
      RECT 40.91 4.064 40.955 4.21 ;
      RECT 40.905 4.069 40.91 4.211 ;
      RECT 40.885 4.069 40.905 4.213 ;
      RECT 40.865 4.067 40.885 4.218 ;
      RECT 40.83 4.066 40.865 4.225 ;
      RECT 40.8 4.065 40.83 4.235 ;
      RECT 40.75 4.064 40.8 4.245 ;
      RECT 40.66 4.061 40.745 4.335 ;
      RECT 40.635 4.055 40.66 4.335 ;
      RECT 40.62 4.045 40.635 4.335 ;
      RECT 40.435 4.04 40.485 4.255 ;
      RECT 40.425 4.045 40.435 4.245 ;
      RECT 40.665 4.52 40.925 4.78 ;
      RECT 40.665 4.52 40.955 4.673 ;
      RECT 40.665 4.52 40.99 4.658 ;
      RECT 40.92 4.44 41.11 4.65 ;
      RECT 40.91 4.445 41.12 4.643 ;
      RECT 40.875 4.515 41.12 4.643 ;
      RECT 40.905 4.457 40.925 4.78 ;
      RECT 40.89 4.505 41.12 4.643 ;
      RECT 40.895 4.477 40.925 4.78 ;
      RECT 39.975 3.545 40.045 4.65 ;
      RECT 40.71 3.65 40.97 3.91 ;
      RECT 40.29 3.696 40.305 3.905 ;
      RECT 40.626 3.709 40.71 3.86 ;
      RECT 40.54 3.706 40.626 3.86 ;
      RECT 40.501 3.704 40.54 3.86 ;
      RECT 40.415 3.702 40.501 3.86 ;
      RECT 40.355 3.7 40.415 3.871 ;
      RECT 40.32 3.698 40.355 3.889 ;
      RECT 40.305 3.696 40.32 3.9 ;
      RECT 40.275 3.696 40.29 3.913 ;
      RECT 40.265 3.696 40.275 3.918 ;
      RECT 40.24 3.695 40.265 3.923 ;
      RECT 40.225 3.69 40.24 3.929 ;
      RECT 40.22 3.683 40.225 3.934 ;
      RECT 40.195 3.674 40.22 3.94 ;
      RECT 40.15 3.653 40.195 3.953 ;
      RECT 40.14 3.637 40.15 3.963 ;
      RECT 40.125 3.63 40.14 3.973 ;
      RECT 40.115 3.623 40.125 3.99 ;
      RECT 40.11 3.62 40.115 4.02 ;
      RECT 40.105 3.618 40.11 4.05 ;
      RECT 40.1 3.616 40.105 4.087 ;
      RECT 40.085 3.612 40.1 4.154 ;
      RECT 40.085 4.445 40.095 4.645 ;
      RECT 40.08 3.608 40.085 4.28 ;
      RECT 40.08 4.432 40.085 4.65 ;
      RECT 40.075 3.606 40.08 4.365 ;
      RECT 40.075 4.422 40.08 4.65 ;
      RECT 40.06 3.577 40.075 4.65 ;
      RECT 40.045 3.55 40.06 4.65 ;
      RECT 39.97 3.545 39.975 3.9 ;
      RECT 39.97 3.955 39.975 4.65 ;
      RECT 39.955 3.545 39.97 3.878 ;
      RECT 39.965 3.977 39.97 4.65 ;
      RECT 39.955 4.017 39.965 4.65 ;
      RECT 39.92 3.545 39.955 3.82 ;
      RECT 39.95 4.052 39.955 4.65 ;
      RECT 39.935 4.107 39.95 4.65 ;
      RECT 39.93 4.172 39.935 4.65 ;
      RECT 39.915 4.22 39.93 4.65 ;
      RECT 39.89 3.545 39.92 3.775 ;
      RECT 39.91 4.275 39.915 4.65 ;
      RECT 39.895 4.335 39.91 4.65 ;
      RECT 39.89 4.383 39.895 4.648 ;
      RECT 39.885 3.545 39.89 3.768 ;
      RECT 39.885 4.415 39.89 4.643 ;
      RECT 39.86 3.545 39.885 3.76 ;
      RECT 39.85 3.55 39.86 3.75 ;
      RECT 40.065 4.825 40.085 5.065 ;
      RECT 39.295 4.755 39.3 4.965 ;
      RECT 40.575 4.828 40.585 5.023 ;
      RECT 40.57 4.818 40.575 5.026 ;
      RECT 40.49 4.815 40.57 5.049 ;
      RECT 40.486 4.815 40.49 5.071 ;
      RECT 40.4 4.815 40.486 5.081 ;
      RECT 40.385 4.815 40.4 5.089 ;
      RECT 40.356 4.816 40.385 5.087 ;
      RECT 40.27 4.821 40.356 5.083 ;
      RECT 40.257 4.825 40.27 5.079 ;
      RECT 40.171 4.825 40.257 5.075 ;
      RECT 40.085 4.825 40.171 5.069 ;
      RECT 40.001 4.825 40.065 5.063 ;
      RECT 39.915 4.825 40.001 5.058 ;
      RECT 39.895 4.825 39.915 5.054 ;
      RECT 39.835 4.82 39.895 5.051 ;
      RECT 39.807 4.814 39.835 5.048 ;
      RECT 39.721 4.809 39.807 5.044 ;
      RECT 39.635 4.803 39.721 5.038 ;
      RECT 39.56 4.785 39.635 5.033 ;
      RECT 39.525 4.762 39.56 5.029 ;
      RECT 39.515 4.752 39.525 5.028 ;
      RECT 39.46 4.75 39.515 5.027 ;
      RECT 39.385 4.75 39.46 5.023 ;
      RECT 39.375 4.75 39.385 5.018 ;
      RECT 39.36 4.75 39.375 5.01 ;
      RECT 39.31 4.752 39.36 4.988 ;
      RECT 39.3 4.755 39.31 4.968 ;
      RECT 39.29 4.76 39.295 4.963 ;
      RECT 39.285 4.765 39.29 4.958 ;
      RECT 37.395 3.41 37.655 3.67 ;
      RECT 37.385 3.44 37.655 3.65 ;
      RECT 39.305 3.355 39.565 3.615 ;
      RECT 39.3 3.43 39.305 3.616 ;
      RECT 39.275 3.435 39.3 3.618 ;
      RECT 39.26 3.442 39.275 3.621 ;
      RECT 39.2 3.46 39.26 3.626 ;
      RECT 39.17 3.48 39.2 3.633 ;
      RECT 39.145 3.488 39.17 3.638 ;
      RECT 39.12 3.496 39.145 3.64 ;
      RECT 39.102 3.5 39.12 3.639 ;
      RECT 39.016 3.498 39.102 3.639 ;
      RECT 38.93 3.496 39.016 3.639 ;
      RECT 38.844 3.494 38.93 3.638 ;
      RECT 38.758 3.492 38.844 3.638 ;
      RECT 38.672 3.49 38.758 3.638 ;
      RECT 38.586 3.488 38.672 3.638 ;
      RECT 38.5 3.486 38.586 3.637 ;
      RECT 38.482 3.485 38.5 3.637 ;
      RECT 38.396 3.484 38.482 3.637 ;
      RECT 38.31 3.482 38.396 3.637 ;
      RECT 38.224 3.481 38.31 3.636 ;
      RECT 38.138 3.48 38.224 3.636 ;
      RECT 38.052 3.478 38.138 3.636 ;
      RECT 37.966 3.477 38.052 3.636 ;
      RECT 37.88 3.475 37.966 3.635 ;
      RECT 37.856 3.473 37.88 3.635 ;
      RECT 37.77 3.466 37.856 3.635 ;
      RECT 37.741 3.458 37.77 3.635 ;
      RECT 37.655 3.45 37.741 3.635 ;
      RECT 37.375 3.447 37.385 3.645 ;
      RECT 38.88 4.41 38.885 4.76 ;
      RECT 38.65 4.5 38.79 4.76 ;
      RECT 39.125 4.185 39.17 4.395 ;
      RECT 39.18 4.196 39.19 4.39 ;
      RECT 39.17 4.188 39.18 4.395 ;
      RECT 39.105 4.185 39.125 4.4 ;
      RECT 39.075 4.185 39.105 4.423 ;
      RECT 39.065 4.185 39.075 4.448 ;
      RECT 39.06 4.185 39.065 4.458 ;
      RECT 39.005 4.185 39.06 4.498 ;
      RECT 39 4.185 39.005 4.538 ;
      RECT 38.995 4.187 39 4.543 ;
      RECT 38.98 4.197 38.995 4.554 ;
      RECT 38.935 4.255 38.98 4.59 ;
      RECT 38.925 4.31 38.935 4.624 ;
      RECT 38.91 4.337 38.925 4.64 ;
      RECT 38.9 4.364 38.91 4.76 ;
      RECT 38.885 4.387 38.9 4.76 ;
      RECT 38.875 4.427 38.88 4.76 ;
      RECT 38.87 4.437 38.875 4.76 ;
      RECT 38.865 4.452 38.87 4.76 ;
      RECT 38.855 4.457 38.865 4.76 ;
      RECT 38.79 4.48 38.855 4.76 ;
      RECT 38.26 3.975 38.48 4.185 ;
      RECT 38.26 3.982 38.49 4.18 ;
      RECT 37.565 3.99 38.49 4.165 ;
      RECT 38.085 3.885 38.475 4.165 ;
      RECT 36.865 3.9 37.125 4.16 ;
      RECT 37.5 3.935 37.635 4.12 ;
      RECT 37.425 3.925 37.52 4.115 ;
      RECT 37.415 3.99 38.49 4.111 ;
      RECT 37.165 3.99 38.49 4.11 ;
      RECT 37.19 3.91 37.43 4.11 ;
      RECT 36.865 3.915 37.45 4.098 ;
      RECT 38.78 3.94 38.82 4.025 ;
      RECT 36.865 3.975 38.04 4.098 ;
      RECT 36.865 3.965 37.925 4.098 ;
      RECT 36.865 3.946 37.83 4.098 ;
      RECT 37.65 3.94 37.83 4.165 ;
      RECT 38.085 3.92 38.78 3.955 ;
      RECT 37.185 3.912 37.43 4.11 ;
      RECT 37.2 3.902 37.41 4.11 ;
      RECT 37.215 3.895 37.41 4.11 ;
      RECT 37.38 4.415 37.64 4.675 ;
      RECT 37.38 4.455 37.745 4.665 ;
      RECT 37.38 4.457 37.75 4.664 ;
      RECT 37.38 4.465 37.755 4.661 ;
      RECT 36.305 3.54 36.405 5.065 ;
      RECT 36.495 4.68 36.545 4.94 ;
      RECT 36.49 3.553 36.495 3.74 ;
      RECT 36.485 4.661 36.495 4.94 ;
      RECT 36.485 3.55 36.49 3.748 ;
      RECT 36.47 3.544 36.485 3.755 ;
      RECT 36.48 4.649 36.485 5.023 ;
      RECT 36.47 4.637 36.48 5.06 ;
      RECT 36.46 3.54 36.47 3.762 ;
      RECT 36.46 4.622 36.47 5.065 ;
      RECT 36.455 3.54 36.46 3.77 ;
      RECT 36.435 4.592 36.46 5.065 ;
      RECT 36.415 3.54 36.455 3.818 ;
      RECT 36.425 4.552 36.435 5.065 ;
      RECT 36.415 4.507 36.425 5.065 ;
      RECT 36.41 3.54 36.415 3.888 ;
      RECT 36.41 4.465 36.415 5.065 ;
      RECT 36.405 3.54 36.41 4.365 ;
      RECT 36.405 4.447 36.41 5.065 ;
      RECT 36.295 3.543 36.305 5.065 ;
      RECT 36.28 3.55 36.295 5.061 ;
      RECT 36.275 3.56 36.28 5.056 ;
      RECT 36.27 3.76 36.275 4.948 ;
      RECT 36.265 3.845 36.27 4.5 ;
      RECT 35.13 10.205 35.425 10.435 ;
      RECT 35.19 8.725 35.36 10.435 ;
      RECT 35.185 9.095 35.535 9.445 ;
      RECT 35.13 8.725 35.42 8.955 ;
      RECT 34.14 10.205 34.435 10.435 ;
      RECT 34.2 8.725 34.37 10.435 ;
      RECT 34.14 8.725 34.43 8.955 ;
      RECT 34.14 8.76 34.99 8.92 ;
      RECT 34.825 8.355 34.99 8.92 ;
      RECT 34.14 8.755 34.535 8.92 ;
      RECT 34.76 8.355 35.05 8.585 ;
      RECT 34.76 8.385 35.22 8.555 ;
      RECT 34.725 4.025 35.045 4.26 ;
      RECT 34.725 4.055 35.215 4.225 ;
      RECT 34.725 3.69 34.915 4.26 ;
      RECT 34.14 3.655 34.43 3.885 ;
      RECT 34.14 3.69 34.915 3.86 ;
      RECT 34.2 2.175 34.37 3.885 ;
      RECT 34.14 2.175 34.435 2.405 ;
      RECT 33.77 4.025 34.06 4.255 ;
      RECT 33.77 4.055 34.23 4.225 ;
      RECT 33.835 2.95 34 4.255 ;
      RECT 32.35 2.915 32.64 3.145 ;
      RECT 32.35 2.95 34 3.12 ;
      RECT 32.41 2.175 32.58 3.145 ;
      RECT 32.35 2.175 32.64 2.405 ;
      RECT 32.35 10.205 32.64 10.435 ;
      RECT 32.41 9.465 32.58 10.435 ;
      RECT 32.41 9.555 34 9.725 ;
      RECT 33.83 8.355 34 9.725 ;
      RECT 32.35 9.465 32.64 9.695 ;
      RECT 33.77 8.355 34.06 8.585 ;
      RECT 33.77 8.385 34.23 8.555 ;
      RECT 30.385 4.725 30.735 5.075 ;
      RECT 30.475 3.32 30.645 5.075 ;
      RECT 32.78 3.26 33.13 3.61 ;
      RECT 30.475 3.32 32.095 3.495 ;
      RECT 30.475 3.32 32.75 3.49 ;
      RECT 32.61 3.315 33.13 3.485 ;
      RECT 32.805 9.09 33.13 9.415 ;
      RECT 28.2 9.04 28.55 9.39 ;
      RECT 32.78 9.095 33.13 9.325 ;
      RECT 28.02 9.095 28.55 9.325 ;
      RECT 32.61 9.12 33.13 9.295 ;
      RECT 27.85 9.125 28.55 9.295 ;
      RECT 28.02 9.12 33.13 9.29 ;
      RECT 32.005 3.66 32.325 3.98 ;
      RECT 31.98 3.655 32.27 3.885 ;
      RECT 31.935 3.685 32.325 3.86 ;
      RECT 31.805 3.685 32.325 3.855 ;
      RECT 32.005 8.66 32.325 8.98 ;
      RECT 31.98 8.725 32.325 8.955 ;
      RECT 31.805 8.755 32.325 8.925 ;
      RECT 27.795 4.96 27.835 5.22 ;
      RECT 27.835 4.94 27.84 4.95 ;
      RECT 29.165 4.185 29.175 4.406 ;
      RECT 29.095 4.18 29.165 4.531 ;
      RECT 29.085 4.18 29.095 4.658 ;
      RECT 29.06 4.18 29.085 4.705 ;
      RECT 29.035 4.18 29.06 4.783 ;
      RECT 29.015 4.18 29.035 4.853 ;
      RECT 28.99 4.18 29.015 4.893 ;
      RECT 28.98 4.18 28.99 4.913 ;
      RECT 28.97 4.182 28.98 4.921 ;
      RECT 28.965 4.187 28.97 4.378 ;
      RECT 28.965 4.387 28.97 4.922 ;
      RECT 28.96 4.432 28.965 4.923 ;
      RECT 28.95 4.497 28.96 4.924 ;
      RECT 28.94 4.592 28.95 4.926 ;
      RECT 28.935 4.645 28.94 4.928 ;
      RECT 28.93 4.665 28.935 4.929 ;
      RECT 28.875 4.69 28.93 4.935 ;
      RECT 28.835 4.725 28.875 4.944 ;
      RECT 28.825 4.742 28.835 4.949 ;
      RECT 28.816 4.748 28.825 4.951 ;
      RECT 28.73 4.786 28.816 4.962 ;
      RECT 28.725 4.825 28.73 4.972 ;
      RECT 28.65 4.832 28.725 4.982 ;
      RECT 28.63 4.842 28.65 4.993 ;
      RECT 28.6 4.849 28.63 5.001 ;
      RECT 28.575 4.856 28.6 5.008 ;
      RECT 28.551 4.862 28.575 5.013 ;
      RECT 28.465 4.875 28.551 5.025 ;
      RECT 28.387 4.882 28.465 5.043 ;
      RECT 28.301 4.877 28.387 5.061 ;
      RECT 28.215 4.872 28.301 5.081 ;
      RECT 28.135 4.866 28.215 5.098 ;
      RECT 28.07 4.862 28.135 5.127 ;
      RECT 28.065 4.576 28.07 4.6 ;
      RECT 28.055 4.852 28.07 5.155 ;
      RECT 28.06 4.57 28.065 4.64 ;
      RECT 28.055 4.564 28.06 4.71 ;
      RECT 28.05 4.558 28.055 4.788 ;
      RECT 28.05 4.835 28.055 5.22 ;
      RECT 28.042 4.555 28.05 5.22 ;
      RECT 27.956 4.553 28.042 5.22 ;
      RECT 27.87 4.551 27.956 5.22 ;
      RECT 27.86 4.552 27.87 5.22 ;
      RECT 27.855 4.557 27.86 5.22 ;
      RECT 27.845 4.57 27.855 5.22 ;
      RECT 27.84 4.592 27.845 5.22 ;
      RECT 27.835 4.952 27.84 5.22 ;
      RECT 28.465 4.42 28.47 4.64 ;
      RECT 28.97 3.455 29.005 3.715 ;
      RECT 28.955 3.455 28.97 3.723 ;
      RECT 28.926 3.455 28.955 3.745 ;
      RECT 28.84 3.455 28.926 3.805 ;
      RECT 28.82 3.455 28.84 3.87 ;
      RECT 28.76 3.455 28.82 4.035 ;
      RECT 28.755 3.455 28.76 4.183 ;
      RECT 28.75 3.455 28.755 4.195 ;
      RECT 28.745 3.455 28.75 4.221 ;
      RECT 28.715 3.641 28.745 4.301 ;
      RECT 28.71 3.689 28.715 4.39 ;
      RECT 28.705 3.703 28.71 4.405 ;
      RECT 28.7 3.722 28.705 4.435 ;
      RECT 28.695 3.737 28.7 4.451 ;
      RECT 28.69 3.752 28.695 4.473 ;
      RECT 28.685 3.772 28.69 4.495 ;
      RECT 28.675 3.792 28.685 4.528 ;
      RECT 28.66 3.834 28.675 4.59 ;
      RECT 28.655 3.865 28.66 4.63 ;
      RECT 28.65 3.877 28.655 4.635 ;
      RECT 28.645 3.889 28.65 4.64 ;
      RECT 28.64 3.902 28.645 4.64 ;
      RECT 28.635 3.92 28.64 4.64 ;
      RECT 28.63 3.94 28.635 4.64 ;
      RECT 28.625 3.952 28.63 4.64 ;
      RECT 28.62 3.965 28.625 4.64 ;
      RECT 28.6 4 28.62 4.64 ;
      RECT 28.55 4.102 28.6 4.64 ;
      RECT 28.545 4.187 28.55 4.64 ;
      RECT 28.54 4.195 28.545 4.64 ;
      RECT 28.535 4.212 28.54 4.64 ;
      RECT 28.53 4.227 28.535 4.64 ;
      RECT 28.495 4.292 28.53 4.64 ;
      RECT 28.48 4.357 28.495 4.64 ;
      RECT 28.475 4.387 28.48 4.64 ;
      RECT 28.47 4.412 28.475 4.64 ;
      RECT 28.455 4.422 28.465 4.64 ;
      RECT 28.44 4.435 28.455 4.633 ;
      RECT 28.185 4.025 28.255 4.235 ;
      RECT 27.975 4.002 27.98 4.195 ;
      RECT 25.43 3.93 25.69 4.19 ;
      RECT 28.265 4.212 28.27 4.215 ;
      RECT 28.255 4.03 28.265 4.23 ;
      RECT 28.156 4.023 28.185 4.235 ;
      RECT 28.07 4.015 28.156 4.235 ;
      RECT 28.055 4.009 28.07 4.233 ;
      RECT 28.035 4.008 28.055 4.22 ;
      RECT 28.03 4.007 28.035 4.203 ;
      RECT 27.98 4.004 28.03 4.198 ;
      RECT 27.95 4.001 27.975 4.193 ;
      RECT 27.93 3.999 27.95 4.188 ;
      RECT 27.915 3.997 27.93 4.185 ;
      RECT 27.885 3.995 27.915 4.183 ;
      RECT 27.82 3.991 27.885 4.175 ;
      RECT 27.79 3.986 27.82 4.17 ;
      RECT 27.77 3.984 27.79 4.168 ;
      RECT 27.74 3.981 27.77 4.163 ;
      RECT 27.68 3.977 27.74 4.155 ;
      RECT 27.675 3.974 27.68 4.15 ;
      RECT 27.605 3.972 27.675 4.145 ;
      RECT 27.576 3.968 27.605 4.138 ;
      RECT 27.49 3.963 27.576 4.13 ;
      RECT 27.456 3.958 27.49 4.122 ;
      RECT 27.37 3.95 27.456 4.114 ;
      RECT 27.331 3.943 27.37 4.106 ;
      RECT 27.245 3.938 27.331 4.098 ;
      RECT 27.18 3.932 27.245 4.088 ;
      RECT 27.16 3.927 27.18 4.083 ;
      RECT 27.151 3.924 27.16 4.082 ;
      RECT 27.065 3.92 27.151 4.076 ;
      RECT 27.025 3.916 27.065 4.068 ;
      RECT 27.005 3.912 27.025 4.066 ;
      RECT 26.945 3.912 27.005 4.063 ;
      RECT 26.925 3.915 26.945 4.061 ;
      RECT 26.904 3.915 26.925 4.061 ;
      RECT 26.818 3.917 26.904 4.065 ;
      RECT 26.732 3.919 26.818 4.071 ;
      RECT 26.646 3.921 26.732 4.078 ;
      RECT 26.56 3.924 26.646 4.084 ;
      RECT 26.526 3.925 26.56 4.089 ;
      RECT 26.44 3.928 26.526 4.094 ;
      RECT 26.411 3.935 26.44 4.099 ;
      RECT 26.325 3.935 26.411 4.104 ;
      RECT 26.292 3.935 26.325 4.109 ;
      RECT 26.206 3.937 26.292 4.114 ;
      RECT 26.12 3.939 26.206 4.121 ;
      RECT 26.056 3.941 26.12 4.127 ;
      RECT 25.97 3.943 26.056 4.133 ;
      RECT 25.967 3.945 25.97 4.136 ;
      RECT 25.881 3.946 25.967 4.14 ;
      RECT 25.795 3.949 25.881 4.147 ;
      RECT 25.776 3.951 25.795 4.151 ;
      RECT 25.69 3.953 25.776 4.156 ;
      RECT 25.42 3.965 25.43 4.16 ;
      RECT 27.59 10.205 27.88 10.435 ;
      RECT 27.65 9.465 27.82 10.435 ;
      RECT 27.54 9.49 27.915 9.86 ;
      RECT 27.59 9.465 27.88 9.86 ;
      RECT 27.655 3.545 27.84 3.755 ;
      RECT 27.65 3.546 27.845 3.753 ;
      RECT 27.645 3.551 27.855 3.748 ;
      RECT 27.64 3.527 27.645 3.745 ;
      RECT 27.61 3.524 27.64 3.738 ;
      RECT 27.605 3.52 27.61 3.729 ;
      RECT 27.57 3.551 27.855 3.724 ;
      RECT 27.345 3.46 27.605 3.72 ;
      RECT 27.645 3.529 27.65 3.748 ;
      RECT 27.65 3.53 27.655 3.753 ;
      RECT 27.345 3.542 27.725 3.72 ;
      RECT 27.345 3.54 27.71 3.72 ;
      RECT 27.345 3.535 27.7 3.72 ;
      RECT 27.3 4.45 27.35 4.735 ;
      RECT 27.245 4.42 27.25 4.735 ;
      RECT 27.215 4.4 27.22 4.735 ;
      RECT 27.365 4.45 27.425 4.71 ;
      RECT 27.36 4.45 27.365 4.718 ;
      RECT 27.35 4.45 27.36 4.73 ;
      RECT 27.265 4.44 27.3 4.735 ;
      RECT 27.26 4.427 27.265 4.735 ;
      RECT 27.25 4.422 27.26 4.735 ;
      RECT 27.23 4.412 27.245 4.735 ;
      RECT 27.22 4.405 27.23 4.735 ;
      RECT 27.21 4.397 27.215 4.735 ;
      RECT 27.18 4.387 27.21 4.735 ;
      RECT 27.165 4.375 27.18 4.735 ;
      RECT 27.15 4.365 27.165 4.73 ;
      RECT 27.13 4.355 27.15 4.705 ;
      RECT 27.12 4.347 27.13 4.682 ;
      RECT 27.09 4.33 27.12 4.672 ;
      RECT 27.085 4.307 27.09 4.663 ;
      RECT 27.08 4.294 27.085 4.661 ;
      RECT 27.065 4.27 27.08 4.655 ;
      RECT 27.06 4.246 27.065 4.649 ;
      RECT 27.05 4.235 27.06 4.644 ;
      RECT 27.045 4.225 27.05 4.64 ;
      RECT 27.04 4.217 27.045 4.637 ;
      RECT 27.03 4.212 27.04 4.633 ;
      RECT 27.025 4.207 27.03 4.629 ;
      RECT 26.94 4.205 27.025 4.604 ;
      RECT 26.91 4.205 26.94 4.57 ;
      RECT 26.895 4.205 26.91 4.553 ;
      RECT 26.84 4.205 26.895 4.498 ;
      RECT 26.835 4.21 26.84 4.447 ;
      RECT 26.825 4.215 26.835 4.437 ;
      RECT 26.82 4.225 26.825 4.423 ;
      RECT 26.77 4.965 27.03 5.225 ;
      RECT 26.69 4.98 27.03 5.201 ;
      RECT 26.67 4.98 27.03 5.196 ;
      RECT 26.646 4.98 27.03 5.194 ;
      RECT 26.56 4.98 27.03 5.189 ;
      RECT 26.41 4.92 26.67 5.185 ;
      RECT 26.365 4.98 27.03 5.18 ;
      RECT 26.36 4.987 27.03 5.175 ;
      RECT 26.375 4.975 26.69 5.185 ;
      RECT 26.265 3.41 26.525 3.67 ;
      RECT 26.265 3.467 26.53 3.663 ;
      RECT 26.265 3.497 26.535 3.595 ;
      RECT 26.325 3.928 26.44 3.93 ;
      RECT 26.411 3.925 26.44 3.93 ;
      RECT 25.435 4.929 25.46 5.169 ;
      RECT 25.42 4.932 25.51 5.163 ;
      RECT 25.415 4.937 25.596 5.158 ;
      RECT 25.41 4.945 25.66 5.156 ;
      RECT 25.41 4.945 25.67 5.155 ;
      RECT 25.405 4.952 25.68 5.148 ;
      RECT 25.405 4.952 25.766 5.137 ;
      RECT 25.4 4.987 25.766 5.133 ;
      RECT 25.4 4.987 25.775 5.122 ;
      RECT 25.68 4.86 25.94 5.12 ;
      RECT 25.39 5.037 25.94 5.118 ;
      RECT 25.66 4.905 25.68 5.153 ;
      RECT 25.596 4.908 25.66 5.157 ;
      RECT 25.51 4.913 25.596 5.162 ;
      RECT 25.44 4.924 25.94 5.12 ;
      RECT 25.46 4.918 25.51 5.167 ;
      RECT 25.585 3.395 25.595 3.657 ;
      RECT 25.575 3.452 25.585 3.66 ;
      RECT 25.55 3.457 25.575 3.666 ;
      RECT 25.525 3.461 25.55 3.678 ;
      RECT 25.515 3.464 25.525 3.688 ;
      RECT 25.51 3.465 25.515 3.693 ;
      RECT 25.505 3.466 25.51 3.698 ;
      RECT 25.5 3.467 25.505 3.7 ;
      RECT 25.475 3.47 25.5 3.703 ;
      RECT 25.445 3.476 25.475 3.706 ;
      RECT 25.38 3.487 25.445 3.709 ;
      RECT 25.335 3.495 25.38 3.713 ;
      RECT 25.32 3.495 25.335 3.721 ;
      RECT 25.315 3.496 25.32 3.728 ;
      RECT 25.31 3.498 25.315 3.731 ;
      RECT 25.305 3.502 25.31 3.734 ;
      RECT 25.295 3.51 25.305 3.738 ;
      RECT 25.29 3.523 25.295 3.743 ;
      RECT 25.285 3.531 25.29 3.745 ;
      RECT 25.28 3.537 25.285 3.745 ;
      RECT 25.275 3.541 25.28 3.748 ;
      RECT 25.27 3.543 25.275 3.751 ;
      RECT 25.265 3.546 25.27 3.754 ;
      RECT 25.255 3.551 25.265 3.758 ;
      RECT 25.25 3.557 25.255 3.763 ;
      RECT 25.24 3.563 25.25 3.767 ;
      RECT 25.225 3.57 25.24 3.773 ;
      RECT 25.196 3.584 25.225 3.783 ;
      RECT 25.11 3.619 25.196 3.815 ;
      RECT 25.09 3.652 25.11 3.844 ;
      RECT 25.07 3.665 25.09 3.855 ;
      RECT 25.05 3.677 25.07 3.866 ;
      RECT 25 3.699 25.05 3.886 ;
      RECT 24.985 3.717 25 3.903 ;
      RECT 24.98 3.723 24.985 3.906 ;
      RECT 24.975 3.727 24.98 3.909 ;
      RECT 24.97 3.731 24.975 3.913 ;
      RECT 24.965 3.733 24.97 3.916 ;
      RECT 24.955 3.74 24.965 3.919 ;
      RECT 24.95 3.745 24.955 3.923 ;
      RECT 24.945 3.747 24.95 3.926 ;
      RECT 24.94 3.751 24.945 3.929 ;
      RECT 24.935 3.753 24.94 3.933 ;
      RECT 24.92 3.758 24.935 3.938 ;
      RECT 24.915 3.763 24.92 3.941 ;
      RECT 24.91 3.771 24.915 3.944 ;
      RECT 24.905 3.773 24.91 3.947 ;
      RECT 24.9 3.775 24.905 3.95 ;
      RECT 24.89 3.777 24.9 3.956 ;
      RECT 24.855 3.791 24.89 3.968 ;
      RECT 24.845 3.806 24.855 3.978 ;
      RECT 24.77 3.835 24.845 4.002 ;
      RECT 24.765 3.86 24.77 4.025 ;
      RECT 24.75 3.864 24.765 4.031 ;
      RECT 24.74 3.872 24.75 4.036 ;
      RECT 24.71 3.885 24.74 4.04 ;
      RECT 24.7 3.9 24.71 4.045 ;
      RECT 24.69 3.905 24.7 4.048 ;
      RECT 24.685 3.907 24.69 4.05 ;
      RECT 24.67 3.91 24.685 4.053 ;
      RECT 24.665 3.912 24.67 4.056 ;
      RECT 24.645 3.917 24.665 4.06 ;
      RECT 24.615 3.922 24.645 4.068 ;
      RECT 24.59 3.929 24.615 4.076 ;
      RECT 24.585 3.934 24.59 4.081 ;
      RECT 24.555 3.937 24.585 4.085 ;
      RECT 24.515 3.94 24.555 4.095 ;
      RECT 24.48 3.937 24.515 4.107 ;
      RECT 24.47 3.933 24.48 4.114 ;
      RECT 24.445 3.929 24.47 4.12 ;
      RECT 24.44 3.925 24.445 4.125 ;
      RECT 24.4 3.922 24.44 4.125 ;
      RECT 24.385 3.907 24.4 4.126 ;
      RECT 24.362 3.895 24.385 4.126 ;
      RECT 24.276 3.895 24.362 4.127 ;
      RECT 24.19 3.895 24.276 4.129 ;
      RECT 24.17 3.895 24.19 4.126 ;
      RECT 24.165 3.9 24.17 4.121 ;
      RECT 24.16 3.905 24.165 4.119 ;
      RECT 24.15 3.915 24.16 4.117 ;
      RECT 24.145 3.921 24.15 4.11 ;
      RECT 24.14 3.923 24.145 4.095 ;
      RECT 24.135 3.927 24.14 4.085 ;
      RECT 25.595 3.395 25.845 3.655 ;
      RECT 23.32 4.93 23.58 5.19 ;
      RECT 25.615 4.42 25.62 4.63 ;
      RECT 25.62 4.425 25.63 4.625 ;
      RECT 25.57 4.42 25.615 4.645 ;
      RECT 25.56 4.42 25.57 4.665 ;
      RECT 25.541 4.42 25.56 4.67 ;
      RECT 25.455 4.42 25.541 4.667 ;
      RECT 25.425 4.422 25.455 4.665 ;
      RECT 25.37 4.432 25.425 4.663 ;
      RECT 25.305 4.446 25.37 4.661 ;
      RECT 25.3 4.454 25.305 4.66 ;
      RECT 25.285 4.457 25.3 4.658 ;
      RECT 25.22 4.467 25.285 4.654 ;
      RECT 25.172 4.481 25.22 4.655 ;
      RECT 25.086 4.498 25.172 4.669 ;
      RECT 25 4.519 25.086 4.686 ;
      RECT 24.98 4.532 25 4.696 ;
      RECT 24.935 4.54 24.98 4.703 ;
      RECT 24.9 4.548 24.935 4.711 ;
      RECT 24.866 4.556 24.9 4.719 ;
      RECT 24.78 4.57 24.866 4.731 ;
      RECT 24.745 4.587 24.78 4.743 ;
      RECT 24.736 4.596 24.745 4.747 ;
      RECT 24.65 4.614 24.736 4.764 ;
      RECT 24.591 4.641 24.65 4.791 ;
      RECT 24.505 4.668 24.591 4.819 ;
      RECT 24.485 4.69 24.505 4.839 ;
      RECT 24.425 4.705 24.485 4.855 ;
      RECT 24.415 4.717 24.425 4.868 ;
      RECT 24.41 4.722 24.415 4.871 ;
      RECT 24.4 4.725 24.41 4.874 ;
      RECT 24.395 4.727 24.4 4.877 ;
      RECT 24.365 4.735 24.395 4.884 ;
      RECT 24.35 4.742 24.365 4.892 ;
      RECT 24.34 4.747 24.35 4.896 ;
      RECT 24.335 4.75 24.34 4.899 ;
      RECT 24.325 4.752 24.335 4.902 ;
      RECT 24.29 4.762 24.325 4.911 ;
      RECT 24.215 4.785 24.29 4.933 ;
      RECT 24.195 4.803 24.215 4.951 ;
      RECT 24.165 4.81 24.195 4.961 ;
      RECT 24.145 4.818 24.165 4.971 ;
      RECT 24.135 4.824 24.145 4.978 ;
      RECT 24.116 4.829 24.135 4.984 ;
      RECT 24.03 4.849 24.116 5.004 ;
      RECT 24.015 4.869 24.03 5.023 ;
      RECT 23.97 4.881 24.015 5.034 ;
      RECT 23.905 4.902 23.97 5.057 ;
      RECT 23.865 4.922 23.905 5.078 ;
      RECT 23.855 4.932 23.865 5.088 ;
      RECT 23.805 4.944 23.855 5.099 ;
      RECT 23.785 4.96 23.805 5.111 ;
      RECT 23.755 4.97 23.785 5.117 ;
      RECT 23.745 4.975 23.755 5.119 ;
      RECT 23.676 4.976 23.745 5.125 ;
      RECT 23.59 4.978 23.676 5.135 ;
      RECT 23.58 4.979 23.59 5.14 ;
      RECT 24.85 5.005 25.04 5.215 ;
      RECT 24.84 5.01 25.05 5.208 ;
      RECT 24.825 5.01 25.05 5.173 ;
      RECT 24.745 4.895 25.005 5.155 ;
      RECT 23.66 4.425 23.845 4.72 ;
      RECT 23.65 4.425 23.845 4.718 ;
      RECT 23.635 4.425 23.85 4.713 ;
      RECT 23.635 4.425 23.855 4.71 ;
      RECT 23.63 4.425 23.855 4.708 ;
      RECT 23.625 4.68 23.855 4.698 ;
      RECT 23.63 4.425 23.89 4.685 ;
      RECT 23.59 3.46 23.85 3.72 ;
      RECT 23.4 3.385 23.486 3.718 ;
      RECT 23.375 3.389 23.53 3.714 ;
      RECT 23.486 3.381 23.53 3.714 ;
      RECT 23.486 3.382 23.535 3.713 ;
      RECT 23.4 3.387 23.55 3.712 ;
      RECT 23.375 3.395 23.59 3.711 ;
      RECT 23.37 3.39 23.55 3.706 ;
      RECT 23.36 3.405 23.59 3.613 ;
      RECT 23.36 3.457 23.79 3.613 ;
      RECT 23.36 3.45 23.77 3.613 ;
      RECT 23.36 3.437 23.74 3.613 ;
      RECT 23.36 3.425 23.68 3.613 ;
      RECT 23.36 3.41 23.655 3.613 ;
      RECT 22.56 4.04 22.695 4.335 ;
      RECT 22.82 4.063 22.825 4.25 ;
      RECT 23.54 3.96 23.685 4.195 ;
      RECT 23.7 3.96 23.705 4.185 ;
      RECT 23.735 3.971 23.74 4.165 ;
      RECT 23.73 3.963 23.735 4.17 ;
      RECT 23.71 3.96 23.73 4.175 ;
      RECT 23.705 3.96 23.71 4.183 ;
      RECT 23.695 3.96 23.7 4.188 ;
      RECT 23.685 3.96 23.695 4.193 ;
      RECT 23.515 3.962 23.54 4.195 ;
      RECT 23.465 3.969 23.515 4.195 ;
      RECT 23.46 3.974 23.465 4.195 ;
      RECT 23.421 3.979 23.46 4.196 ;
      RECT 23.335 3.991 23.421 4.197 ;
      RECT 23.326 4.001 23.335 4.197 ;
      RECT 23.24 4.01 23.326 4.199 ;
      RECT 23.216 4.02 23.24 4.201 ;
      RECT 23.13 4.031 23.216 4.202 ;
      RECT 23.1 4.042 23.13 4.204 ;
      RECT 23.07 4.047 23.1 4.206 ;
      RECT 23.045 4.053 23.07 4.209 ;
      RECT 23.03 4.058 23.045 4.21 ;
      RECT 22.985 4.064 23.03 4.21 ;
      RECT 22.98 4.069 22.985 4.211 ;
      RECT 22.96 4.069 22.98 4.213 ;
      RECT 22.94 4.067 22.96 4.218 ;
      RECT 22.905 4.066 22.94 4.225 ;
      RECT 22.875 4.065 22.905 4.235 ;
      RECT 22.825 4.064 22.875 4.245 ;
      RECT 22.735 4.061 22.82 4.335 ;
      RECT 22.71 4.055 22.735 4.335 ;
      RECT 22.695 4.045 22.71 4.335 ;
      RECT 22.51 4.04 22.56 4.255 ;
      RECT 22.5 4.045 22.51 4.245 ;
      RECT 22.74 4.52 23 4.78 ;
      RECT 22.74 4.52 23.03 4.673 ;
      RECT 22.74 4.52 23.065 4.658 ;
      RECT 22.995 4.44 23.185 4.65 ;
      RECT 22.985 4.445 23.195 4.643 ;
      RECT 22.95 4.515 23.195 4.643 ;
      RECT 22.98 4.457 23 4.78 ;
      RECT 22.965 4.505 23.195 4.643 ;
      RECT 22.97 4.477 23 4.78 ;
      RECT 22.05 3.545 22.12 4.65 ;
      RECT 22.785 3.65 23.045 3.91 ;
      RECT 22.365 3.696 22.38 3.905 ;
      RECT 22.701 3.709 22.785 3.86 ;
      RECT 22.615 3.706 22.701 3.86 ;
      RECT 22.576 3.704 22.615 3.86 ;
      RECT 22.49 3.702 22.576 3.86 ;
      RECT 22.43 3.7 22.49 3.871 ;
      RECT 22.395 3.698 22.43 3.889 ;
      RECT 22.38 3.696 22.395 3.9 ;
      RECT 22.35 3.696 22.365 3.913 ;
      RECT 22.34 3.696 22.35 3.918 ;
      RECT 22.315 3.695 22.34 3.923 ;
      RECT 22.3 3.69 22.315 3.929 ;
      RECT 22.295 3.683 22.3 3.934 ;
      RECT 22.27 3.674 22.295 3.94 ;
      RECT 22.225 3.653 22.27 3.953 ;
      RECT 22.215 3.637 22.225 3.963 ;
      RECT 22.2 3.63 22.215 3.973 ;
      RECT 22.19 3.623 22.2 3.99 ;
      RECT 22.185 3.62 22.19 4.02 ;
      RECT 22.18 3.618 22.185 4.05 ;
      RECT 22.175 3.616 22.18 4.087 ;
      RECT 22.16 3.612 22.175 4.154 ;
      RECT 22.16 4.445 22.17 4.645 ;
      RECT 22.155 3.608 22.16 4.28 ;
      RECT 22.155 4.432 22.16 4.65 ;
      RECT 22.15 3.606 22.155 4.365 ;
      RECT 22.15 4.422 22.155 4.65 ;
      RECT 22.135 3.577 22.15 4.65 ;
      RECT 22.12 3.55 22.135 4.65 ;
      RECT 22.045 3.545 22.05 3.9 ;
      RECT 22.045 3.955 22.05 4.65 ;
      RECT 22.03 3.545 22.045 3.878 ;
      RECT 22.04 3.977 22.045 4.65 ;
      RECT 22.03 4.017 22.04 4.65 ;
      RECT 21.995 3.545 22.03 3.82 ;
      RECT 22.025 4.052 22.03 4.65 ;
      RECT 22.01 4.107 22.025 4.65 ;
      RECT 22.005 4.172 22.01 4.65 ;
      RECT 21.99 4.22 22.005 4.65 ;
      RECT 21.965 3.545 21.995 3.775 ;
      RECT 21.985 4.275 21.99 4.65 ;
      RECT 21.97 4.335 21.985 4.65 ;
      RECT 21.965 4.383 21.97 4.648 ;
      RECT 21.96 3.545 21.965 3.768 ;
      RECT 21.96 4.415 21.965 4.643 ;
      RECT 21.935 3.545 21.96 3.76 ;
      RECT 21.925 3.55 21.935 3.75 ;
      RECT 22.14 4.825 22.16 5.065 ;
      RECT 21.37 4.755 21.375 4.965 ;
      RECT 22.65 4.828 22.66 5.023 ;
      RECT 22.645 4.818 22.65 5.026 ;
      RECT 22.565 4.815 22.645 5.049 ;
      RECT 22.561 4.815 22.565 5.071 ;
      RECT 22.475 4.815 22.561 5.081 ;
      RECT 22.46 4.815 22.475 5.089 ;
      RECT 22.431 4.816 22.46 5.087 ;
      RECT 22.345 4.821 22.431 5.083 ;
      RECT 22.332 4.825 22.345 5.079 ;
      RECT 22.246 4.825 22.332 5.075 ;
      RECT 22.16 4.825 22.246 5.069 ;
      RECT 22.076 4.825 22.14 5.063 ;
      RECT 21.99 4.825 22.076 5.058 ;
      RECT 21.97 4.825 21.99 5.054 ;
      RECT 21.91 4.82 21.97 5.051 ;
      RECT 21.882 4.814 21.91 5.048 ;
      RECT 21.796 4.809 21.882 5.044 ;
      RECT 21.71 4.803 21.796 5.038 ;
      RECT 21.635 4.785 21.71 5.033 ;
      RECT 21.6 4.762 21.635 5.029 ;
      RECT 21.59 4.752 21.6 5.028 ;
      RECT 21.535 4.75 21.59 5.027 ;
      RECT 21.46 4.75 21.535 5.023 ;
      RECT 21.45 4.75 21.46 5.018 ;
      RECT 21.435 4.75 21.45 5.01 ;
      RECT 21.385 4.752 21.435 4.988 ;
      RECT 21.375 4.755 21.385 4.968 ;
      RECT 21.365 4.76 21.37 4.963 ;
      RECT 21.36 4.765 21.365 4.958 ;
      RECT 19.47 3.41 19.73 3.67 ;
      RECT 19.46 3.44 19.73 3.65 ;
      RECT 21.38 3.355 21.64 3.615 ;
      RECT 21.375 3.43 21.38 3.616 ;
      RECT 21.35 3.435 21.375 3.618 ;
      RECT 21.335 3.442 21.35 3.621 ;
      RECT 21.275 3.46 21.335 3.626 ;
      RECT 21.245 3.48 21.275 3.633 ;
      RECT 21.22 3.488 21.245 3.638 ;
      RECT 21.195 3.496 21.22 3.64 ;
      RECT 21.177 3.5 21.195 3.639 ;
      RECT 21.091 3.498 21.177 3.639 ;
      RECT 21.005 3.496 21.091 3.639 ;
      RECT 20.919 3.494 21.005 3.638 ;
      RECT 20.833 3.492 20.919 3.638 ;
      RECT 20.747 3.49 20.833 3.638 ;
      RECT 20.661 3.488 20.747 3.638 ;
      RECT 20.575 3.486 20.661 3.637 ;
      RECT 20.557 3.485 20.575 3.637 ;
      RECT 20.471 3.484 20.557 3.637 ;
      RECT 20.385 3.482 20.471 3.637 ;
      RECT 20.299 3.481 20.385 3.636 ;
      RECT 20.213 3.48 20.299 3.636 ;
      RECT 20.127 3.478 20.213 3.636 ;
      RECT 20.041 3.477 20.127 3.636 ;
      RECT 19.955 3.475 20.041 3.635 ;
      RECT 19.931 3.473 19.955 3.635 ;
      RECT 19.845 3.466 19.931 3.635 ;
      RECT 19.816 3.458 19.845 3.635 ;
      RECT 19.73 3.45 19.816 3.635 ;
      RECT 19.45 3.447 19.46 3.645 ;
      RECT 20.955 4.41 20.96 4.76 ;
      RECT 20.725 4.5 20.865 4.76 ;
      RECT 21.2 4.185 21.245 4.395 ;
      RECT 21.255 4.196 21.265 4.39 ;
      RECT 21.245 4.188 21.255 4.395 ;
      RECT 21.18 4.185 21.2 4.4 ;
      RECT 21.15 4.185 21.18 4.423 ;
      RECT 21.14 4.185 21.15 4.448 ;
      RECT 21.135 4.185 21.14 4.458 ;
      RECT 21.08 4.185 21.135 4.498 ;
      RECT 21.075 4.185 21.08 4.538 ;
      RECT 21.07 4.187 21.075 4.543 ;
      RECT 21.055 4.197 21.07 4.554 ;
      RECT 21.01 4.255 21.055 4.59 ;
      RECT 21 4.31 21.01 4.624 ;
      RECT 20.985 4.337 21 4.64 ;
      RECT 20.975 4.364 20.985 4.76 ;
      RECT 20.96 4.387 20.975 4.76 ;
      RECT 20.95 4.427 20.955 4.76 ;
      RECT 20.945 4.437 20.95 4.76 ;
      RECT 20.94 4.452 20.945 4.76 ;
      RECT 20.93 4.457 20.94 4.76 ;
      RECT 20.865 4.48 20.93 4.76 ;
      RECT 20.335 3.975 20.555 4.185 ;
      RECT 20.335 3.982 20.565 4.18 ;
      RECT 19.64 3.99 20.565 4.165 ;
      RECT 20.16 3.885 20.55 4.165 ;
      RECT 18.94 3.9 19.2 4.16 ;
      RECT 19.575 3.935 19.71 4.12 ;
      RECT 19.5 3.925 19.595 4.115 ;
      RECT 19.49 3.99 20.565 4.111 ;
      RECT 19.24 3.99 20.565 4.11 ;
      RECT 19.265 3.91 19.505 4.11 ;
      RECT 18.94 3.915 19.525 4.098 ;
      RECT 20.855 3.94 20.895 4.025 ;
      RECT 18.94 3.975 20.115 4.098 ;
      RECT 18.94 3.965 20 4.098 ;
      RECT 18.94 3.946 19.905 4.098 ;
      RECT 19.725 3.94 19.905 4.165 ;
      RECT 20.16 3.92 20.855 3.955 ;
      RECT 19.26 3.912 19.505 4.11 ;
      RECT 19.275 3.902 19.485 4.11 ;
      RECT 19.29 3.895 19.485 4.11 ;
      RECT 19.455 4.415 19.715 4.675 ;
      RECT 19.455 4.455 19.82 4.665 ;
      RECT 19.455 4.457 19.825 4.664 ;
      RECT 19.455 4.465 19.83 4.661 ;
      RECT 18.38 3.54 18.48 5.065 ;
      RECT 18.57 4.68 18.62 4.94 ;
      RECT 18.565 3.553 18.57 3.74 ;
      RECT 18.56 4.661 18.57 4.94 ;
      RECT 18.56 3.55 18.565 3.748 ;
      RECT 18.545 3.544 18.56 3.755 ;
      RECT 18.555 4.649 18.56 5.023 ;
      RECT 18.545 4.637 18.555 5.06 ;
      RECT 18.535 3.54 18.545 3.762 ;
      RECT 18.535 4.622 18.545 5.065 ;
      RECT 18.53 3.54 18.535 3.77 ;
      RECT 18.51 4.592 18.535 5.065 ;
      RECT 18.49 3.54 18.53 3.818 ;
      RECT 18.5 4.552 18.51 5.065 ;
      RECT 18.49 4.507 18.5 5.065 ;
      RECT 18.485 3.54 18.49 3.888 ;
      RECT 18.485 4.465 18.49 5.065 ;
      RECT 18.48 3.54 18.485 4.365 ;
      RECT 18.48 4.447 18.485 5.065 ;
      RECT 18.37 3.543 18.38 5.065 ;
      RECT 18.355 3.55 18.37 5.061 ;
      RECT 18.35 3.56 18.355 5.056 ;
      RECT 18.345 3.76 18.35 4.948 ;
      RECT 18.34 3.845 18.345 4.5 ;
      RECT 16.56 10.205 16.85 10.435 ;
      RECT 16.62 9.46 16.79 10.435 ;
      RECT 16.53 9.46 16.88 9.75 ;
      RECT 16.155 8.72 16.505 9.01 ;
      RECT 16.015 8.755 16.505 8.925 ;
      RECT 106.805 7.39 107.155 7.68 ;
      RECT 102.07 2.435 102.445 2.805 ;
      RECT 96.05 3.52 96.31 3.78 ;
      RECT 88.88 7.39 89.23 7.68 ;
      RECT 84.145 2.435 84.52 2.805 ;
      RECT 78.125 3.52 78.385 3.78 ;
      RECT 70.955 7.39 71.305 7.68 ;
      RECT 66.22 2.435 66.595 2.805 ;
      RECT 60.2 3.52 60.46 3.78 ;
      RECT 53.03 7.39 53.38 7.68 ;
      RECT 48.295 2.435 48.67 2.805 ;
      RECT 42.275 3.52 42.535 3.78 ;
      RECT 35.105 7.39 35.455 7.68 ;
      RECT 30.37 2.435 30.745 2.805 ;
      RECT 24.35 3.52 24.61 3.78 ;
    LAYER mcon ;
      RECT 106.895 7.455 107.065 7.625 ;
      RECT 106.89 8.755 107.06 8.925 ;
      RECT 106.89 10.235 107.06 10.405 ;
      RECT 106.52 8.385 106.69 8.555 ;
      RECT 106.515 4.055 106.685 4.225 ;
      RECT 105.9 2.205 106.07 2.375 ;
      RECT 105.9 3.685 106.07 3.855 ;
      RECT 105.9 8.755 106.07 8.925 ;
      RECT 105.9 10.235 106.07 10.405 ;
      RECT 105.53 4.055 105.7 4.225 ;
      RECT 105.53 8.385 105.7 8.555 ;
      RECT 104.54 3.315 104.71 3.485 ;
      RECT 104.54 9.125 104.71 9.295 ;
      RECT 104.11 2.205 104.28 2.375 ;
      RECT 104.11 2.945 104.28 3.115 ;
      RECT 104.11 9.495 104.28 9.665 ;
      RECT 104.11 10.235 104.28 10.405 ;
      RECT 103.74 3.685 103.91 3.855 ;
      RECT 103.74 8.755 103.91 8.925 ;
      RECT 100.685 4.2 100.855 4.37 ;
      RECT 100.475 3.54 100.645 3.71 ;
      RECT 100.16 4.45 100.33 4.62 ;
      RECT 99.78 9.125 99.95 9.295 ;
      RECT 99.775 4.045 99.945 4.215 ;
      RECT 99.56 4.61 99.73 4.78 ;
      RECT 99.54 5.01 99.71 5.18 ;
      RECT 99.365 3.565 99.535 3.735 ;
      RECT 99.35 9.495 99.52 9.665 ;
      RECT 99.35 10.235 99.52 10.405 ;
      RECT 98.87 4.545 99.04 4.715 ;
      RECT 98.545 4.23 98.715 4.4 ;
      RECT 98.48 5.01 98.65 5.18 ;
      RECT 98.08 4.995 98.25 5.165 ;
      RECT 98.04 3.48 98.21 3.65 ;
      RECT 97.14 3.98 97.31 4.15 ;
      RECT 97.14 4.44 97.31 4.61 ;
      RECT 97.14 4.955 97.31 5.125 ;
      RECT 97.025 3.515 97.195 3.685 ;
      RECT 96.56 5.025 96.73 5.195 ;
      RECT 96.08 3.555 96.25 3.725 ;
      RECT 95.865 3.93 96.035 4.1 ;
      RECT 95.365 4.53 95.535 4.7 ;
      RECT 95.25 3.98 95.42 4.15 ;
      RECT 95.08 3.43 95.25 3.6 ;
      RECT 94.705 4.46 94.875 4.63 ;
      RECT 94.22 4.06 94.39 4.23 ;
      RECT 94.17 4.835 94.34 5.005 ;
      RECT 93.68 4.46 93.85 4.63 ;
      RECT 93.645 3.565 93.815 3.735 ;
      RECT 93.08 4.775 93.25 4.945 ;
      RECT 92.775 4.205 92.945 4.375 ;
      RECT 92.075 3.995 92.245 4.165 ;
      RECT 91.34 4.475 91.51 4.645 ;
      RECT 91.17 3.46 91.34 3.63 ;
      RECT 90.995 3.915 91.165 4.085 ;
      RECT 90.075 3.565 90.245 3.735 ;
      RECT 90.07 4.88 90.24 5.05 ;
      RECT 88.97 7.455 89.14 7.625 ;
      RECT 88.965 8.755 89.135 8.925 ;
      RECT 88.965 10.235 89.135 10.405 ;
      RECT 88.595 8.385 88.765 8.555 ;
      RECT 88.59 4.055 88.76 4.225 ;
      RECT 87.975 2.205 88.145 2.375 ;
      RECT 87.975 3.685 88.145 3.855 ;
      RECT 87.975 8.755 88.145 8.925 ;
      RECT 87.975 10.235 88.145 10.405 ;
      RECT 87.605 4.055 87.775 4.225 ;
      RECT 87.605 8.385 87.775 8.555 ;
      RECT 86.615 3.315 86.785 3.485 ;
      RECT 86.615 9.125 86.785 9.295 ;
      RECT 86.185 2.205 86.355 2.375 ;
      RECT 86.185 2.945 86.355 3.115 ;
      RECT 86.185 9.495 86.355 9.665 ;
      RECT 86.185 10.235 86.355 10.405 ;
      RECT 85.815 3.685 85.985 3.855 ;
      RECT 85.815 8.755 85.985 8.925 ;
      RECT 82.76 4.2 82.93 4.37 ;
      RECT 82.55 3.54 82.72 3.71 ;
      RECT 82.235 4.45 82.405 4.62 ;
      RECT 81.855 9.125 82.025 9.295 ;
      RECT 81.85 4.045 82.02 4.215 ;
      RECT 81.635 4.61 81.805 4.78 ;
      RECT 81.615 5.01 81.785 5.18 ;
      RECT 81.44 3.565 81.61 3.735 ;
      RECT 81.425 9.495 81.595 9.665 ;
      RECT 81.425 10.235 81.595 10.405 ;
      RECT 80.945 4.545 81.115 4.715 ;
      RECT 80.62 4.23 80.79 4.4 ;
      RECT 80.555 5.01 80.725 5.18 ;
      RECT 80.155 4.995 80.325 5.165 ;
      RECT 80.115 3.48 80.285 3.65 ;
      RECT 79.215 3.98 79.385 4.15 ;
      RECT 79.215 4.44 79.385 4.61 ;
      RECT 79.215 4.955 79.385 5.125 ;
      RECT 79.1 3.515 79.27 3.685 ;
      RECT 78.635 5.025 78.805 5.195 ;
      RECT 78.155 3.555 78.325 3.725 ;
      RECT 77.94 3.93 78.11 4.1 ;
      RECT 77.44 4.53 77.61 4.7 ;
      RECT 77.325 3.98 77.495 4.15 ;
      RECT 77.155 3.43 77.325 3.6 ;
      RECT 76.78 4.46 76.95 4.63 ;
      RECT 76.295 4.06 76.465 4.23 ;
      RECT 76.245 4.835 76.415 5.005 ;
      RECT 75.755 4.46 75.925 4.63 ;
      RECT 75.72 3.565 75.89 3.735 ;
      RECT 75.155 4.775 75.325 4.945 ;
      RECT 74.85 4.205 75.02 4.375 ;
      RECT 74.15 3.995 74.32 4.165 ;
      RECT 73.415 4.475 73.585 4.645 ;
      RECT 73.245 3.46 73.415 3.63 ;
      RECT 73.07 3.915 73.24 4.085 ;
      RECT 72.15 3.565 72.32 3.735 ;
      RECT 72.145 4.88 72.315 5.05 ;
      RECT 71.045 7.455 71.215 7.625 ;
      RECT 71.04 8.755 71.21 8.925 ;
      RECT 71.04 10.235 71.21 10.405 ;
      RECT 70.67 8.385 70.84 8.555 ;
      RECT 70.665 4.055 70.835 4.225 ;
      RECT 70.05 2.205 70.22 2.375 ;
      RECT 70.05 3.685 70.22 3.855 ;
      RECT 70.05 8.755 70.22 8.925 ;
      RECT 70.05 10.235 70.22 10.405 ;
      RECT 69.68 4.055 69.85 4.225 ;
      RECT 69.68 8.385 69.85 8.555 ;
      RECT 68.69 3.315 68.86 3.485 ;
      RECT 68.69 9.125 68.86 9.295 ;
      RECT 68.26 2.205 68.43 2.375 ;
      RECT 68.26 2.945 68.43 3.115 ;
      RECT 68.26 9.495 68.43 9.665 ;
      RECT 68.26 10.235 68.43 10.405 ;
      RECT 67.89 3.685 68.06 3.855 ;
      RECT 67.89 8.755 68.06 8.925 ;
      RECT 64.835 4.2 65.005 4.37 ;
      RECT 64.625 3.54 64.795 3.71 ;
      RECT 64.31 4.45 64.48 4.62 ;
      RECT 63.93 9.125 64.1 9.295 ;
      RECT 63.925 4.045 64.095 4.215 ;
      RECT 63.71 4.61 63.88 4.78 ;
      RECT 63.69 5.01 63.86 5.18 ;
      RECT 63.515 3.565 63.685 3.735 ;
      RECT 63.5 9.495 63.67 9.665 ;
      RECT 63.5 10.235 63.67 10.405 ;
      RECT 63.02 4.545 63.19 4.715 ;
      RECT 62.695 4.23 62.865 4.4 ;
      RECT 62.63 5.01 62.8 5.18 ;
      RECT 62.23 4.995 62.4 5.165 ;
      RECT 62.19 3.48 62.36 3.65 ;
      RECT 61.29 3.98 61.46 4.15 ;
      RECT 61.29 4.44 61.46 4.61 ;
      RECT 61.29 4.955 61.46 5.125 ;
      RECT 61.175 3.515 61.345 3.685 ;
      RECT 60.71 5.025 60.88 5.195 ;
      RECT 60.23 3.555 60.4 3.725 ;
      RECT 60.015 3.93 60.185 4.1 ;
      RECT 59.515 4.53 59.685 4.7 ;
      RECT 59.4 3.98 59.57 4.15 ;
      RECT 59.23 3.43 59.4 3.6 ;
      RECT 58.855 4.46 59.025 4.63 ;
      RECT 58.37 4.06 58.54 4.23 ;
      RECT 58.32 4.835 58.49 5.005 ;
      RECT 57.83 4.46 58 4.63 ;
      RECT 57.795 3.565 57.965 3.735 ;
      RECT 57.23 4.775 57.4 4.945 ;
      RECT 56.925 4.205 57.095 4.375 ;
      RECT 56.225 3.995 56.395 4.165 ;
      RECT 55.49 4.475 55.66 4.645 ;
      RECT 55.32 3.46 55.49 3.63 ;
      RECT 55.145 3.915 55.315 4.085 ;
      RECT 54.225 3.565 54.395 3.735 ;
      RECT 54.22 4.88 54.39 5.05 ;
      RECT 53.12 7.455 53.29 7.625 ;
      RECT 53.115 8.755 53.285 8.925 ;
      RECT 53.115 10.235 53.285 10.405 ;
      RECT 52.745 8.385 52.915 8.555 ;
      RECT 52.74 4.055 52.91 4.225 ;
      RECT 52.125 2.205 52.295 2.375 ;
      RECT 52.125 3.685 52.295 3.855 ;
      RECT 52.125 8.755 52.295 8.925 ;
      RECT 52.125 10.235 52.295 10.405 ;
      RECT 51.755 4.055 51.925 4.225 ;
      RECT 51.755 8.385 51.925 8.555 ;
      RECT 50.765 3.315 50.935 3.485 ;
      RECT 50.765 9.125 50.935 9.295 ;
      RECT 50.335 2.205 50.505 2.375 ;
      RECT 50.335 2.945 50.505 3.115 ;
      RECT 50.335 9.495 50.505 9.665 ;
      RECT 50.335 10.235 50.505 10.405 ;
      RECT 49.965 3.685 50.135 3.855 ;
      RECT 49.965 8.755 50.135 8.925 ;
      RECT 46.91 4.2 47.08 4.37 ;
      RECT 46.7 3.54 46.87 3.71 ;
      RECT 46.385 4.45 46.555 4.62 ;
      RECT 46.005 9.125 46.175 9.295 ;
      RECT 46 4.045 46.17 4.215 ;
      RECT 45.785 4.61 45.955 4.78 ;
      RECT 45.765 5.01 45.935 5.18 ;
      RECT 45.59 3.565 45.76 3.735 ;
      RECT 45.575 9.495 45.745 9.665 ;
      RECT 45.575 10.235 45.745 10.405 ;
      RECT 45.095 4.545 45.265 4.715 ;
      RECT 44.77 4.23 44.94 4.4 ;
      RECT 44.705 5.01 44.875 5.18 ;
      RECT 44.305 4.995 44.475 5.165 ;
      RECT 44.265 3.48 44.435 3.65 ;
      RECT 43.365 3.98 43.535 4.15 ;
      RECT 43.365 4.44 43.535 4.61 ;
      RECT 43.365 4.955 43.535 5.125 ;
      RECT 43.25 3.515 43.42 3.685 ;
      RECT 42.785 5.025 42.955 5.195 ;
      RECT 42.305 3.555 42.475 3.725 ;
      RECT 42.09 3.93 42.26 4.1 ;
      RECT 41.59 4.53 41.76 4.7 ;
      RECT 41.475 3.98 41.645 4.15 ;
      RECT 41.305 3.43 41.475 3.6 ;
      RECT 40.93 4.46 41.1 4.63 ;
      RECT 40.445 4.06 40.615 4.23 ;
      RECT 40.395 4.835 40.565 5.005 ;
      RECT 39.905 4.46 40.075 4.63 ;
      RECT 39.87 3.565 40.04 3.735 ;
      RECT 39.305 4.775 39.475 4.945 ;
      RECT 39 4.205 39.17 4.375 ;
      RECT 38.3 3.995 38.47 4.165 ;
      RECT 37.565 4.475 37.735 4.645 ;
      RECT 37.395 3.46 37.565 3.63 ;
      RECT 37.22 3.915 37.39 4.085 ;
      RECT 36.3 3.565 36.47 3.735 ;
      RECT 36.295 4.88 36.465 5.05 ;
      RECT 35.195 7.455 35.365 7.625 ;
      RECT 35.19 8.755 35.36 8.925 ;
      RECT 35.19 10.235 35.36 10.405 ;
      RECT 34.82 8.385 34.99 8.555 ;
      RECT 34.815 4.055 34.985 4.225 ;
      RECT 34.2 2.205 34.37 2.375 ;
      RECT 34.2 3.685 34.37 3.855 ;
      RECT 34.2 8.755 34.37 8.925 ;
      RECT 34.2 10.235 34.37 10.405 ;
      RECT 33.83 4.055 34 4.225 ;
      RECT 33.83 8.385 34 8.555 ;
      RECT 32.84 3.315 33.01 3.485 ;
      RECT 32.84 9.125 33.01 9.295 ;
      RECT 32.41 2.205 32.58 2.375 ;
      RECT 32.41 2.945 32.58 3.115 ;
      RECT 32.41 9.495 32.58 9.665 ;
      RECT 32.41 10.235 32.58 10.405 ;
      RECT 32.04 3.685 32.21 3.855 ;
      RECT 32.04 8.755 32.21 8.925 ;
      RECT 28.985 4.2 29.155 4.37 ;
      RECT 28.775 3.54 28.945 3.71 ;
      RECT 28.46 4.45 28.63 4.62 ;
      RECT 28.08 9.125 28.25 9.295 ;
      RECT 28.075 4.045 28.245 4.215 ;
      RECT 27.86 4.61 28.03 4.78 ;
      RECT 27.84 5.01 28.01 5.18 ;
      RECT 27.665 3.565 27.835 3.735 ;
      RECT 27.65 9.495 27.82 9.665 ;
      RECT 27.65 10.235 27.82 10.405 ;
      RECT 27.17 4.545 27.34 4.715 ;
      RECT 26.845 4.23 27.015 4.4 ;
      RECT 26.78 5.01 26.95 5.18 ;
      RECT 26.38 4.995 26.55 5.165 ;
      RECT 26.34 3.48 26.51 3.65 ;
      RECT 25.44 3.98 25.61 4.15 ;
      RECT 25.44 4.44 25.61 4.61 ;
      RECT 25.44 4.955 25.61 5.125 ;
      RECT 25.325 3.515 25.495 3.685 ;
      RECT 24.86 5.025 25.03 5.195 ;
      RECT 24.38 3.555 24.55 3.725 ;
      RECT 24.165 3.93 24.335 4.1 ;
      RECT 23.665 4.53 23.835 4.7 ;
      RECT 23.55 3.98 23.72 4.15 ;
      RECT 23.38 3.43 23.55 3.6 ;
      RECT 23.005 4.46 23.175 4.63 ;
      RECT 22.52 4.06 22.69 4.23 ;
      RECT 22.47 4.835 22.64 5.005 ;
      RECT 21.98 4.46 22.15 4.63 ;
      RECT 21.945 3.565 22.115 3.735 ;
      RECT 21.38 4.775 21.55 4.945 ;
      RECT 21.075 4.205 21.245 4.375 ;
      RECT 20.375 3.995 20.545 4.165 ;
      RECT 19.64 4.475 19.81 4.645 ;
      RECT 19.47 3.46 19.64 3.63 ;
      RECT 19.295 3.915 19.465 4.085 ;
      RECT 18.375 3.565 18.545 3.735 ;
      RECT 18.37 4.88 18.54 5.05 ;
      RECT 16.62 9.495 16.79 9.665 ;
      RECT 16.62 10.235 16.79 10.405 ;
      RECT 16.25 8.755 16.42 8.925 ;
    LAYER li1 ;
      RECT 106.89 7.455 107.06 8.925 ;
      RECT 106.89 7.455 107.065 8.715 ;
      RECT 106.52 9.405 106.99 9.575 ;
      RECT 106.52 8.385 106.69 9.575 ;
      RECT 106.515 3.035 106.685 4.225 ;
      RECT 106.515 3.035 106.985 3.205 ;
      RECT 105.9 3.895 106.075 5.155 ;
      RECT 105.9 3.685 106.07 5.155 ;
      RECT 105.9 7.455 106.07 8.925 ;
      RECT 105.9 7.455 106.075 8.715 ;
      RECT 105.53 3.035 105.7 4.225 ;
      RECT 105.53 3.035 106 3.205 ;
      RECT 105.53 9.405 106 9.575 ;
      RECT 105.53 8.385 105.7 9.575 ;
      RECT 104.54 4.015 104.715 5.155 ;
      RECT 104.54 1.865 104.71 5.155 ;
      RECT 104.54 1.865 104.715 2.415 ;
      RECT 104.54 10.195 104.715 10.745 ;
      RECT 104.54 7.455 104.71 10.745 ;
      RECT 104.54 7.455 104.715 8.595 ;
      RECT 104.11 3.895 104.285 5.155 ;
      RECT 104.11 2.945 104.28 5.155 ;
      RECT 104.11 7.455 104.28 9.665 ;
      RECT 104.11 7.455 104.285 8.715 ;
      RECT 103.68 3.925 103.85 5.155 ;
      RECT 103.74 2.145 103.91 4.095 ;
      RECT 103.68 1.865 103.85 2.315 ;
      RECT 103.68 10.295 103.85 10.745 ;
      RECT 103.74 8.515 103.91 10.465 ;
      RECT 103.68 7.455 103.85 8.685 ;
      RECT 103.155 3.895 103.33 5.155 ;
      RECT 103.155 1.865 103.325 5.155 ;
      RECT 103.155 3.365 103.565 3.695 ;
      RECT 103.155 2.525 103.565 2.855 ;
      RECT 103.155 1.865 103.33 2.355 ;
      RECT 103.155 10.255 103.33 10.745 ;
      RECT 103.155 7.455 103.325 10.745 ;
      RECT 103.155 9.755 103.565 10.085 ;
      RECT 103.155 8.915 103.565 9.245 ;
      RECT 103.155 7.455 103.33 8.715 ;
      RECT 101.27 4.687 101.285 4.738 ;
      RECT 101.265 4.667 101.27 4.785 ;
      RECT 101.25 4.657 101.265 4.853 ;
      RECT 101.225 4.637 101.25 4.908 ;
      RECT 101.185 4.622 101.225 4.928 ;
      RECT 101.14 4.616 101.185 4.956 ;
      RECT 101.07 4.606 101.14 4.973 ;
      RECT 101.05 4.598 101.07 4.973 ;
      RECT 100.99 4.592 101.05 4.965 ;
      RECT 100.931 4.583 100.99 4.953 ;
      RECT 100.845 4.572 100.931 4.936 ;
      RECT 100.823 4.563 100.845 4.924 ;
      RECT 100.737 4.556 100.823 4.911 ;
      RECT 100.651 4.543 100.737 4.892 ;
      RECT 100.565 4.531 100.651 4.872 ;
      RECT 100.535 4.52 100.565 4.859 ;
      RECT 100.485 4.506 100.535 4.851 ;
      RECT 100.465 4.495 100.485 4.843 ;
      RECT 100.416 4.484 100.465 4.835 ;
      RECT 100.33 4.463 100.416 4.82 ;
      RECT 100.285 4.45 100.33 4.805 ;
      RECT 100.24 4.45 100.285 4.785 ;
      RECT 100.185 4.45 100.24 4.72 ;
      RECT 100.16 4.45 100.185 4.643 ;
      RECT 100.685 4.187 100.855 4.37 ;
      RECT 100.685 4.187 100.87 4.328 ;
      RECT 100.685 4.187 100.875 4.27 ;
      RECT 100.745 3.955 100.88 4.246 ;
      RECT 100.745 3.959 100.885 4.229 ;
      RECT 100.69 4.122 100.885 4.229 ;
      RECT 100.715 3.967 100.855 4.37 ;
      RECT 100.715 3.971 100.895 4.17 ;
      RECT 100.7 4.057 100.895 4.17 ;
      RECT 100.71 3.987 100.855 4.37 ;
      RECT 100.71 3.99 100.905 4.083 ;
      RECT 100.705 4.007 100.905 4.083 ;
      RECT 100.475 3.227 100.645 3.71 ;
      RECT 100.47 3.222 100.62 3.7 ;
      RECT 100.47 3.229 100.65 3.694 ;
      RECT 100.46 3.223 100.62 3.673 ;
      RECT 100.46 3.239 100.665 3.632 ;
      RECT 100.43 3.224 100.62 3.595 ;
      RECT 100.43 3.254 100.675 3.535 ;
      RECT 100.425 3.226 100.62 3.533 ;
      RECT 100.405 3.235 100.65 3.49 ;
      RECT 100.38 3.251 100.665 3.402 ;
      RECT 100.38 3.27 100.69 3.393 ;
      RECT 100.375 3.307 100.69 3.345 ;
      RECT 100.38 3.287 100.695 3.313 ;
      RECT 100.475 3.221 100.585 3.71 ;
      RECT 100.561 3.22 100.585 3.71 ;
      RECT 99.795 4.005 99.8 4.216 ;
      RECT 100.395 4.005 100.4 4.19 ;
      RECT 100.46 4.045 100.465 4.158 ;
      RECT 100.455 4.037 100.46 4.164 ;
      RECT 100.45 4.027 100.455 4.172 ;
      RECT 100.445 4.017 100.45 4.181 ;
      RECT 100.44 4.007 100.445 4.185 ;
      RECT 100.4 4.005 100.44 4.188 ;
      RECT 100.372 4.004 100.395 4.192 ;
      RECT 100.286 4.001 100.372 4.199 ;
      RECT 100.2 3.997 100.286 4.21 ;
      RECT 100.18 3.995 100.2 4.216 ;
      RECT 100.162 3.994 100.18 4.219 ;
      RECT 100.076 3.992 100.162 4.226 ;
      RECT 99.99 3.987 100.076 4.239 ;
      RECT 99.971 3.984 99.99 4.244 ;
      RECT 99.885 3.982 99.971 4.235 ;
      RECT 99.875 3.982 99.885 4.228 ;
      RECT 99.8 3.995 99.875 4.222 ;
      RECT 99.785 4.006 99.795 4.216 ;
      RECT 99.775 4.008 99.785 4.215 ;
      RECT 99.765 4.012 99.775 4.211 ;
      RECT 99.76 4.015 99.765 4.205 ;
      RECT 99.75 4.017 99.76 4.199 ;
      RECT 99.745 4.02 99.75 4.193 ;
      RECT 99.78 10.195 99.955 10.745 ;
      RECT 99.78 7.455 99.95 10.745 ;
      RECT 99.78 7.455 99.955 8.595 ;
      RECT 99.725 4.606 99.73 4.81 ;
      RECT 99.71 4.593 99.725 4.903 ;
      RECT 99.695 4.574 99.71 5.18 ;
      RECT 99.66 4.54 99.695 5.18 ;
      RECT 99.656 4.51 99.66 5.18 ;
      RECT 99.57 4.392 99.656 5.18 ;
      RECT 99.56 4.267 99.57 5.18 ;
      RECT 99.545 4.235 99.56 5.18 ;
      RECT 99.54 4.21 99.545 5.18 ;
      RECT 99.535 4.2 99.54 5.136 ;
      RECT 99.52 4.172 99.535 5.041 ;
      RECT 99.505 4.138 99.52 4.94 ;
      RECT 99.5 4.116 99.505 4.893 ;
      RECT 99.495 4.105 99.5 4.863 ;
      RECT 99.49 4.095 99.495 4.829 ;
      RECT 99.48 4.082 99.49 4.797 ;
      RECT 99.455 4.058 99.48 4.723 ;
      RECT 99.45 4.038 99.455 4.648 ;
      RECT 99.445 4.032 99.45 4.623 ;
      RECT 99.44 4.027 99.445 4.588 ;
      RECT 99.435 4.022 99.44 4.563 ;
      RECT 99.43 4.02 99.435 4.543 ;
      RECT 99.425 4.02 99.43 4.528 ;
      RECT 99.42 4.02 99.425 4.488 ;
      RECT 99.41 4.02 99.42 4.46 ;
      RECT 99.4 4.02 99.41 4.405 ;
      RECT 99.385 4.02 99.4 4.343 ;
      RECT 99.38 4.019 99.385 4.288 ;
      RECT 99.365 4.018 99.38 4.268 ;
      RECT 99.305 4.016 99.365 4.242 ;
      RECT 99.27 4.017 99.305 4.222 ;
      RECT 99.265 4.019 99.27 4.212 ;
      RECT 99.255 4.038 99.265 4.202 ;
      RECT 99.25 4.065 99.255 4.133 ;
      RECT 99.365 3.49 99.535 3.735 ;
      RECT 99.4 3.261 99.535 3.735 ;
      RECT 99.4 3.263 99.545 3.73 ;
      RECT 99.4 3.265 99.57 3.718 ;
      RECT 99.4 3.268 99.595 3.7 ;
      RECT 99.4 3.273 99.645 3.673 ;
      RECT 99.4 3.278 99.665 3.638 ;
      RECT 99.38 3.28 99.675 3.613 ;
      RECT 99.37 3.375 99.675 3.613 ;
      RECT 99.4 3.26 99.51 3.735 ;
      RECT 99.41 3.257 99.505 3.735 ;
      RECT 99.35 7.455 99.52 9.665 ;
      RECT 99.35 7.455 99.525 8.715 ;
      RECT 98.93 4.522 99.12 4.88 ;
      RECT 98.93 4.534 99.155 4.879 ;
      RECT 98.93 4.562 99.175 4.877 ;
      RECT 98.93 4.587 99.18 4.876 ;
      RECT 98.93 4.645 99.195 4.875 ;
      RECT 98.915 4.518 99.075 4.86 ;
      RECT 98.895 4.527 99.12 4.813 ;
      RECT 98.87 4.538 99.155 4.75 ;
      RECT 98.87 4.622 99.19 4.75 ;
      RECT 98.87 4.597 99.185 4.75 ;
      RECT 98.93 4.513 99.075 4.88 ;
      RECT 99.016 4.512 99.075 4.88 ;
      RECT 99.016 4.511 99.06 4.88 ;
      RECT 98.395 10.255 98.57 10.745 ;
      RECT 98.395 7.455 98.565 10.745 ;
      RECT 98.395 9.755 98.805 10.085 ;
      RECT 98.395 8.915 98.805 9.245 ;
      RECT 98.395 7.455 98.57 8.715 ;
      RECT 98.715 4.027 98.72 4.405 ;
      RECT 98.71 3.995 98.715 4.405 ;
      RECT 98.705 3.967 98.71 4.405 ;
      RECT 98.7 3.947 98.705 4.405 ;
      RECT 98.645 3.93 98.7 4.405 ;
      RECT 98.605 3.915 98.645 4.405 ;
      RECT 98.55 3.902 98.605 4.405 ;
      RECT 98.515 3.893 98.55 4.405 ;
      RECT 98.511 3.891 98.515 4.404 ;
      RECT 98.425 3.887 98.511 4.387 ;
      RECT 98.34 3.879 98.425 4.35 ;
      RECT 98.33 3.875 98.34 4.323 ;
      RECT 98.32 3.875 98.33 4.305 ;
      RECT 98.31 3.877 98.32 4.288 ;
      RECT 98.305 3.882 98.31 4.274 ;
      RECT 98.3 3.886 98.305 4.261 ;
      RECT 98.29 3.891 98.3 4.245 ;
      RECT 98.275 3.905 98.29 4.22 ;
      RECT 98.27 3.911 98.275 4.2 ;
      RECT 98.265 3.913 98.27 4.193 ;
      RECT 98.26 3.917 98.265 4.068 ;
      RECT 98.44 4.717 98.685 5.18 ;
      RECT 98.36 4.69 98.68 5.176 ;
      RECT 98.29 4.725 98.685 5.169 ;
      RECT 98.08 4.98 98.685 5.165 ;
      RECT 98.26 4.748 98.685 5.165 ;
      RECT 98.1 4.94 98.685 5.165 ;
      RECT 98.25 4.76 98.685 5.165 ;
      RECT 98.135 4.877 98.685 5.165 ;
      RECT 98.19 4.802 98.685 5.165 ;
      RECT 98.44 4.667 98.68 5.18 ;
      RECT 98.47 4.66 98.68 5.18 ;
      RECT 98.46 4.662 98.68 5.18 ;
      RECT 98.47 4.657 98.6 5.18 ;
      RECT 98.025 3.22 98.111 3.659 ;
      RECT 98.02 3.22 98.111 3.657 ;
      RECT 98.02 3.22 98.18 3.656 ;
      RECT 98.02 3.22 98.21 3.653 ;
      RECT 98.005 3.227 98.21 3.644 ;
      RECT 98.005 3.227 98.215 3.64 ;
      RECT 98 3.237 98.215 3.633 ;
      RECT 97.995 3.242 98.215 3.608 ;
      RECT 97.995 3.242 98.23 3.59 ;
      RECT 98.02 3.22 98.25 3.505 ;
      RECT 97.99 3.247 98.25 3.503 ;
      RECT 98 3.24 98.255 3.441 ;
      RECT 97.99 3.362 98.26 3.424 ;
      RECT 97.975 3.257 98.255 3.375 ;
      RECT 97.97 3.267 98.255 3.275 ;
      RECT 98.05 4.038 98.055 4.115 ;
      RECT 98.04 4.032 98.05 4.305 ;
      RECT 98.03 4.024 98.04 4.326 ;
      RECT 98.02 4.015 98.03 4.348 ;
      RECT 98.015 4.01 98.02 4.365 ;
      RECT 97.975 4.01 98.015 4.405 ;
      RECT 97.955 4.01 97.975 4.46 ;
      RECT 97.95 4.01 97.955 4.488 ;
      RECT 97.94 4.01 97.95 4.503 ;
      RECT 97.905 4.01 97.94 4.545 ;
      RECT 97.9 4.01 97.905 4.588 ;
      RECT 97.89 4.01 97.9 4.603 ;
      RECT 97.875 4.01 97.89 4.623 ;
      RECT 97.86 4.01 97.875 4.65 ;
      RECT 97.855 4.011 97.86 4.668 ;
      RECT 97.835 4.012 97.855 4.675 ;
      RECT 97.78 4.013 97.835 4.695 ;
      RECT 97.77 4.014 97.78 4.709 ;
      RECT 97.765 4.017 97.77 4.708 ;
      RECT 97.725 4.09 97.765 4.706 ;
      RECT 97.71 4.17 97.725 4.704 ;
      RECT 97.685 4.225 97.71 4.702 ;
      RECT 97.67 4.29 97.685 4.701 ;
      RECT 97.625 4.322 97.67 4.698 ;
      RECT 97.54 4.345 97.625 4.693 ;
      RECT 97.515 4.365 97.54 4.688 ;
      RECT 97.445 4.37 97.515 4.684 ;
      RECT 97.425 4.372 97.445 4.681 ;
      RECT 97.34 4.383 97.425 4.675 ;
      RECT 97.335 4.394 97.34 4.67 ;
      RECT 97.325 4.396 97.335 4.67 ;
      RECT 97.29 4.4 97.325 4.668 ;
      RECT 97.24 4.41 97.29 4.655 ;
      RECT 97.22 4.418 97.24 4.64 ;
      RECT 97.14 4.43 97.22 4.623 ;
      RECT 97.305 3.98 97.475 4.19 ;
      RECT 97.421 3.976 97.475 4.19 ;
      RECT 97.226 3.98 97.475 4.181 ;
      RECT 97.226 3.98 97.48 4.17 ;
      RECT 97.14 3.98 97.48 4.161 ;
      RECT 97.14 3.988 97.49 4.105 ;
      RECT 97.14 4 97.495 4.018 ;
      RECT 97.14 4.007 97.5 4.01 ;
      RECT 97.335 3.978 97.475 4.19 ;
      RECT 97.09 4.923 97.335 5.255 ;
      RECT 97.085 4.915 97.09 5.252 ;
      RECT 97.055 4.935 97.335 5.233 ;
      RECT 97.035 4.967 97.335 5.206 ;
      RECT 97.085 4.92 97.262 5.252 ;
      RECT 97.085 4.917 97.176 5.252 ;
      RECT 97.025 3.265 97.195 3.685 ;
      RECT 97.02 3.265 97.195 3.683 ;
      RECT 97.02 3.265 97.22 3.673 ;
      RECT 97.02 3.265 97.24 3.648 ;
      RECT 97.015 3.265 97.24 3.643 ;
      RECT 97.015 3.265 97.25 3.633 ;
      RECT 97.015 3.265 97.255 3.628 ;
      RECT 97.015 3.27 97.26 3.623 ;
      RECT 97.015 3.302 97.275 3.613 ;
      RECT 97.015 3.372 97.3 3.596 ;
      RECT 96.995 3.372 97.3 3.588 ;
      RECT 96.995 3.432 97.31 3.565 ;
      RECT 96.995 3.472 97.32 3.51 ;
      RECT 96.98 3.265 97.255 3.49 ;
      RECT 96.97 3.28 97.26 3.388 ;
      RECT 96.56 4.67 96.73 5.195 ;
      RECT 96.555 4.67 96.73 5.188 ;
      RECT 96.545 4.67 96.735 5.153 ;
      RECT 96.54 4.68 96.735 5.125 ;
      RECT 96.535 4.7 96.735 5.108 ;
      RECT 96.545 4.675 96.74 5.098 ;
      RECT 96.53 4.72 96.74 5.09 ;
      RECT 96.525 4.74 96.74 5.075 ;
      RECT 96.52 4.77 96.74 5.065 ;
      RECT 96.51 4.815 96.74 5.04 ;
      RECT 96.54 4.685 96.745 5.023 ;
      RECT 96.505 4.867 96.745 5.018 ;
      RECT 96.54 4.695 96.75 4.988 ;
      RECT 96.5 4.9 96.75 4.985 ;
      RECT 96.495 4.925 96.75 4.965 ;
      RECT 96.535 4.712 96.76 4.905 ;
      RECT 96.53 4.734 96.77 4.798 ;
      RECT 96.48 3.981 96.495 4.25 ;
      RECT 96.435 3.965 96.48 4.295 ;
      RECT 96.43 3.953 96.435 4.345 ;
      RECT 96.42 3.949 96.43 4.378 ;
      RECT 96.415 3.946 96.42 4.406 ;
      RECT 96.4 3.948 96.415 4.448 ;
      RECT 96.395 3.952 96.4 4.488 ;
      RECT 96.375 3.957 96.395 4.54 ;
      RECT 96.371 3.962 96.375 4.597 ;
      RECT 96.285 3.981 96.371 4.634 ;
      RECT 96.275 4.002 96.285 4.67 ;
      RECT 96.27 4.01 96.275 4.671 ;
      RECT 96.265 4.052 96.27 4.672 ;
      RECT 96.25 4.14 96.265 4.673 ;
      RECT 96.24 4.29 96.25 4.675 ;
      RECT 96.235 4.335 96.24 4.677 ;
      RECT 96.2 4.377 96.235 4.68 ;
      RECT 96.195 4.395 96.2 4.683 ;
      RECT 96.118 4.401 96.195 4.689 ;
      RECT 96.032 4.415 96.118 4.702 ;
      RECT 95.946 4.429 96.032 4.716 ;
      RECT 95.86 4.443 95.946 4.729 ;
      RECT 95.8 4.455 95.86 4.741 ;
      RECT 95.775 4.462 95.8 4.748 ;
      RECT 95.761 4.465 95.775 4.753 ;
      RECT 95.675 4.473 95.761 4.769 ;
      RECT 95.67 4.48 95.675 4.784 ;
      RECT 95.646 4.48 95.67 4.791 ;
      RECT 95.56 4.483 95.646 4.819 ;
      RECT 95.475 4.487 95.56 4.863 ;
      RECT 95.41 4.491 95.475 4.9 ;
      RECT 95.385 4.494 95.41 4.916 ;
      RECT 95.31 4.507 95.385 4.92 ;
      RECT 95.285 4.525 95.31 4.924 ;
      RECT 95.275 4.532 95.285 4.926 ;
      RECT 95.26 4.535 95.275 4.927 ;
      RECT 95.2 4.547 95.26 4.931 ;
      RECT 95.19 4.561 95.2 4.935 ;
      RECT 95.135 4.571 95.19 4.923 ;
      RECT 95.11 4.592 95.135 4.906 ;
      RECT 95.09 4.612 95.11 4.897 ;
      RECT 95.085 4.625 95.09 4.892 ;
      RECT 95.07 4.637 95.085 4.888 ;
      RECT 96.305 3.292 96.31 3.315 ;
      RECT 96.3 3.283 96.305 3.355 ;
      RECT 96.295 3.281 96.3 3.398 ;
      RECT 96.29 3.272 96.295 3.433 ;
      RECT 96.285 3.262 96.29 3.505 ;
      RECT 96.28 3.252 96.285 3.57 ;
      RECT 96.275 3.249 96.28 3.61 ;
      RECT 96.25 3.243 96.275 3.7 ;
      RECT 96.215 3.231 96.25 3.725 ;
      RECT 96.205 3.222 96.215 3.725 ;
      RECT 96.07 3.22 96.08 3.708 ;
      RECT 96.06 3.22 96.07 3.675 ;
      RECT 96.055 3.22 96.06 3.65 ;
      RECT 96.05 3.22 96.055 3.638 ;
      RECT 96.045 3.22 96.05 3.62 ;
      RECT 96.035 3.22 96.045 3.585 ;
      RECT 96.03 3.222 96.035 3.563 ;
      RECT 96.025 3.228 96.03 3.548 ;
      RECT 96.02 3.234 96.025 3.533 ;
      RECT 96.005 3.246 96.02 3.506 ;
      RECT 96 3.257 96.005 3.474 ;
      RECT 95.995 3.267 96 3.458 ;
      RECT 95.985 3.275 95.995 3.427 ;
      RECT 95.98 3.285 95.985 3.401 ;
      RECT 95.975 3.342 95.98 3.384 ;
      RECT 96.08 3.22 96.205 3.725 ;
      RECT 95.795 3.907 96.055 4.205 ;
      RECT 95.79 3.914 96.055 4.203 ;
      RECT 95.795 3.909 96.07 4.198 ;
      RECT 95.785 3.922 96.07 4.195 ;
      RECT 95.785 3.927 96.075 4.188 ;
      RECT 95.78 3.935 96.075 4.185 ;
      RECT 95.78 3.952 96.08 3.983 ;
      RECT 95.795 3.904 96.026 4.205 ;
      RECT 95.85 3.903 96.026 4.205 ;
      RECT 95.85 3.9 95.94 4.205 ;
      RECT 95.85 3.897 95.936 4.205 ;
      RECT 95.54 4.17 95.545 4.183 ;
      RECT 95.535 4.137 95.54 4.188 ;
      RECT 95.53 4.092 95.535 4.195 ;
      RECT 95.525 4.047 95.53 4.203 ;
      RECT 95.52 4.015 95.525 4.211 ;
      RECT 95.515 3.975 95.52 4.212 ;
      RECT 95.5 3.955 95.515 4.214 ;
      RECT 95.425 3.937 95.5 4.226 ;
      RECT 95.415 3.93 95.425 4.237 ;
      RECT 95.41 3.93 95.415 4.239 ;
      RECT 95.38 3.936 95.41 4.243 ;
      RECT 95.34 3.949 95.38 4.243 ;
      RECT 95.315 3.96 95.34 4.229 ;
      RECT 95.3 3.966 95.315 4.212 ;
      RECT 95.29 3.968 95.3 4.203 ;
      RECT 95.285 3.969 95.29 4.198 ;
      RECT 95.28 3.97 95.285 4.193 ;
      RECT 95.275 3.971 95.28 4.19 ;
      RECT 95.25 3.976 95.275 4.18 ;
      RECT 95.24 3.992 95.25 4.167 ;
      RECT 95.235 4.012 95.24 4.162 ;
      RECT 95.245 3.405 95.25 3.601 ;
      RECT 95.23 3.369 95.245 3.603 ;
      RECT 95.22 3.351 95.23 3.608 ;
      RECT 95.21 3.337 95.22 3.612 ;
      RECT 95.165 3.321 95.21 3.622 ;
      RECT 95.16 3.311 95.165 3.631 ;
      RECT 95.115 3.3 95.16 3.637 ;
      RECT 95.11 3.288 95.115 3.644 ;
      RECT 95.095 3.283 95.11 3.648 ;
      RECT 95.08 3.275 95.095 3.653 ;
      RECT 95.07 3.268 95.08 3.658 ;
      RECT 95.06 3.265 95.07 3.663 ;
      RECT 95.05 3.265 95.06 3.664 ;
      RECT 95.045 3.262 95.05 3.663 ;
      RECT 95.01 3.257 95.035 3.662 ;
      RECT 94.986 3.253 95.01 3.661 ;
      RECT 94.9 3.244 94.986 3.658 ;
      RECT 94.885 3.236 94.9 3.655 ;
      RECT 94.863 3.235 94.885 3.654 ;
      RECT 94.777 3.235 94.863 3.652 ;
      RECT 94.691 3.235 94.777 3.65 ;
      RECT 94.605 3.235 94.691 3.647 ;
      RECT 94.595 3.235 94.605 3.638 ;
      RECT 94.565 3.235 94.595 3.598 ;
      RECT 94.555 3.245 94.565 3.553 ;
      RECT 94.55 3.285 94.555 3.538 ;
      RECT 94.545 3.3 94.55 3.525 ;
      RECT 94.515 3.38 94.545 3.487 ;
      RECT 95.035 3.26 95.045 3.663 ;
      RECT 94.86 4.025 94.875 4.63 ;
      RECT 94.865 4.02 94.875 4.63 ;
      RECT 95.03 4.02 95.035 4.203 ;
      RECT 95.02 4.02 95.03 4.233 ;
      RECT 95.005 4.02 95.02 4.293 ;
      RECT 95 4.02 95.005 4.338 ;
      RECT 94.995 4.02 95 4.368 ;
      RECT 94.99 4.02 94.995 4.388 ;
      RECT 94.98 4.02 94.99 4.423 ;
      RECT 94.965 4.02 94.98 4.455 ;
      RECT 94.92 4.02 94.965 4.483 ;
      RECT 94.915 4.02 94.92 4.513 ;
      RECT 94.91 4.02 94.915 4.525 ;
      RECT 94.905 4.02 94.91 4.533 ;
      RECT 94.895 4.02 94.905 4.548 ;
      RECT 94.89 4.02 94.895 4.57 ;
      RECT 94.88 4.02 94.89 4.593 ;
      RECT 94.875 4.02 94.88 4.613 ;
      RECT 94.84 4.035 94.86 4.63 ;
      RECT 94.815 4.052 94.84 4.63 ;
      RECT 94.81 4.062 94.815 4.63 ;
      RECT 94.78 4.077 94.81 4.63 ;
      RECT 94.705 4.119 94.78 4.63 ;
      RECT 94.7 4.15 94.705 4.613 ;
      RECT 94.695 4.154 94.7 4.595 ;
      RECT 94.69 4.158 94.695 4.558 ;
      RECT 94.685 4.342 94.69 4.525 ;
      RECT 94.17 4.531 94.256 5.096 ;
      RECT 94.125 4.533 94.29 5.09 ;
      RECT 94.256 4.53 94.29 5.09 ;
      RECT 94.17 4.532 94.375 5.084 ;
      RECT 94.125 4.542 94.385 5.08 ;
      RECT 94.1 4.534 94.375 5.076 ;
      RECT 94.095 4.537 94.375 5.071 ;
      RECT 94.07 4.552 94.385 5.065 ;
      RECT 94.07 4.577 94.425 5.06 ;
      RECT 94.03 4.585 94.425 5.035 ;
      RECT 94.03 4.612 94.44 5.033 ;
      RECT 94.03 4.642 94.45 5.02 ;
      RECT 94.025 4.787 94.45 5.008 ;
      RECT 94.03 4.716 94.47 5.005 ;
      RECT 94.03 4.773 94.475 4.813 ;
      RECT 94.22 4.052 94.39 4.23 ;
      RECT 94.17 3.991 94.22 4.215 ;
      RECT 93.905 3.971 94.17 4.2 ;
      RECT 93.865 4.035 94.34 4.2 ;
      RECT 93.865 4.025 94.295 4.2 ;
      RECT 93.865 4.022 94.285 4.2 ;
      RECT 93.865 4.01 94.275 4.2 ;
      RECT 93.865 3.995 94.22 4.2 ;
      RECT 93.905 3.967 94.106 4.2 ;
      RECT 93.915 3.945 94.106 4.2 ;
      RECT 93.94 3.93 94.02 4.2 ;
      RECT 93.695 4.46 93.815 4.905 ;
      RECT 93.68 4.46 93.815 4.904 ;
      RECT 93.635 4.482 93.815 4.899 ;
      RECT 93.595 4.531 93.815 4.893 ;
      RECT 93.595 4.531 93.82 4.868 ;
      RECT 93.595 4.531 93.84 4.758 ;
      RECT 93.59 4.561 93.84 4.755 ;
      RECT 93.68 4.46 93.85 4.65 ;
      RECT 93.34 3.245 93.345 3.69 ;
      RECT 93.15 3.245 93.17 3.655 ;
      RECT 93.12 3.245 93.125 3.63 ;
      RECT 93.8 3.552 93.815 3.74 ;
      RECT 93.795 3.537 93.8 3.746 ;
      RECT 93.775 3.51 93.795 3.749 ;
      RECT 93.725 3.477 93.775 3.758 ;
      RECT 93.695 3.457 93.725 3.762 ;
      RECT 93.676 3.445 93.695 3.758 ;
      RECT 93.59 3.417 93.676 3.748 ;
      RECT 93.58 3.392 93.59 3.738 ;
      RECT 93.51 3.36 93.58 3.73 ;
      RECT 93.485 3.32 93.51 3.722 ;
      RECT 93.465 3.302 93.485 3.716 ;
      RECT 93.455 3.292 93.465 3.713 ;
      RECT 93.445 3.285 93.455 3.711 ;
      RECT 93.425 3.272 93.445 3.708 ;
      RECT 93.415 3.262 93.425 3.705 ;
      RECT 93.405 3.255 93.415 3.703 ;
      RECT 93.355 3.247 93.405 3.697 ;
      RECT 93.345 3.245 93.355 3.691 ;
      RECT 93.315 3.245 93.34 3.688 ;
      RECT 93.286 3.245 93.315 3.683 ;
      RECT 93.2 3.245 93.286 3.673 ;
      RECT 93.17 3.245 93.2 3.66 ;
      RECT 93.125 3.245 93.15 3.643 ;
      RECT 93.11 3.245 93.12 3.625 ;
      RECT 93.09 3.252 93.11 3.61 ;
      RECT 93.085 3.267 93.09 3.598 ;
      RECT 93.08 3.272 93.085 3.538 ;
      RECT 93.075 3.277 93.08 3.38 ;
      RECT 93.07 3.28 93.075 3.298 ;
      RECT 92.81 4.57 92.845 4.89 ;
      RECT 93.395 4.755 93.4 4.937 ;
      RECT 93.35 4.637 93.395 4.956 ;
      RECT 93.335 4.614 93.35 4.979 ;
      RECT 93.325 4.604 93.335 4.989 ;
      RECT 93.305 4.599 93.325 5.002 ;
      RECT 93.28 4.597 93.305 5.023 ;
      RECT 93.261 4.596 93.28 5.035 ;
      RECT 93.175 4.593 93.261 5.035 ;
      RECT 93.105 4.588 93.175 5.023 ;
      RECT 93.03 4.584 93.105 4.998 ;
      RECT 92.965 4.58 93.03 4.965 ;
      RECT 92.895 4.577 92.965 4.925 ;
      RECT 92.865 4.573 92.895 4.9 ;
      RECT 92.845 4.571 92.865 4.893 ;
      RECT 92.761 4.569 92.81 4.891 ;
      RECT 92.675 4.566 92.761 4.892 ;
      RECT 92.6 4.565 92.675 4.894 ;
      RECT 92.515 4.565 92.6 4.92 ;
      RECT 92.438 4.566 92.515 4.945 ;
      RECT 92.352 4.567 92.438 4.945 ;
      RECT 92.266 4.567 92.352 4.945 ;
      RECT 92.18 4.568 92.266 4.945 ;
      RECT 92.16 4.569 92.18 4.937 ;
      RECT 92.145 4.575 92.16 4.922 ;
      RECT 92.11 4.595 92.145 4.902 ;
      RECT 92.1 4.615 92.11 4.884 ;
      RECT 93.07 3.92 93.075 4.19 ;
      RECT 93.065 3.911 93.07 4.195 ;
      RECT 93.055 3.901 93.065 4.207 ;
      RECT 93.05 3.89 93.055 4.218 ;
      RECT 93.03 3.884 93.05 4.236 ;
      RECT 92.985 3.881 93.03 4.285 ;
      RECT 92.97 3.88 92.985 4.33 ;
      RECT 92.965 3.88 92.97 4.343 ;
      RECT 92.955 3.88 92.965 4.355 ;
      RECT 92.95 3.881 92.955 4.37 ;
      RECT 92.93 3.889 92.95 4.375 ;
      RECT 92.9 3.905 92.93 4.375 ;
      RECT 92.89 3.917 92.895 4.375 ;
      RECT 92.855 3.932 92.89 4.375 ;
      RECT 92.825 3.952 92.855 4.375 ;
      RECT 92.815 3.977 92.825 4.375 ;
      RECT 92.81 4.005 92.815 4.375 ;
      RECT 92.805 4.035 92.81 4.375 ;
      RECT 92.8 4.052 92.805 4.375 ;
      RECT 92.79 4.08 92.8 4.375 ;
      RECT 92.78 4.115 92.79 4.375 ;
      RECT 92.775 4.15 92.78 4.375 ;
      RECT 92.895 3.915 92.9 4.375 ;
      RECT 91.885 3.245 91.89 3.644 ;
      RECT 91.63 3.245 91.665 3.642 ;
      RECT 91.225 3.28 91.23 3.636 ;
      RECT 91.97 3.283 91.975 3.538 ;
      RECT 91.965 3.281 91.97 3.544 ;
      RECT 91.96 3.28 91.965 3.551 ;
      RECT 91.935 3.273 91.96 3.575 ;
      RECT 91.93 3.266 91.935 3.599 ;
      RECT 91.925 3.262 91.93 3.608 ;
      RECT 91.915 3.257 91.925 3.621 ;
      RECT 91.91 3.254 91.915 3.63 ;
      RECT 91.905 3.252 91.91 3.635 ;
      RECT 91.89 3.248 91.905 3.645 ;
      RECT 91.875 3.242 91.885 3.644 ;
      RECT 91.837 3.24 91.875 3.644 ;
      RECT 91.751 3.242 91.837 3.644 ;
      RECT 91.665 3.244 91.751 3.643 ;
      RECT 91.594 3.245 91.63 3.642 ;
      RECT 91.508 3.247 91.594 3.642 ;
      RECT 91.422 3.249 91.508 3.641 ;
      RECT 91.336 3.251 91.422 3.641 ;
      RECT 91.25 3.254 91.336 3.64 ;
      RECT 91.24 3.26 91.25 3.639 ;
      RECT 91.23 3.272 91.24 3.637 ;
      RECT 91.17 3.307 91.225 3.633 ;
      RECT 91.165 3.337 91.17 3.395 ;
      RECT 91.51 4.552 91.515 4.809 ;
      RECT 91.49 4.471 91.51 4.826 ;
      RECT 91.47 4.465 91.49 4.855 ;
      RECT 91.41 4.452 91.47 4.875 ;
      RECT 91.365 4.436 91.41 4.876 ;
      RECT 91.281 4.424 91.365 4.864 ;
      RECT 91.195 4.411 91.281 4.848 ;
      RECT 91.185 4.404 91.195 4.84 ;
      RECT 91.14 4.401 91.185 4.78 ;
      RECT 91.12 4.397 91.14 4.695 ;
      RECT 91.105 4.395 91.12 4.648 ;
      RECT 91.075 4.392 91.105 4.618 ;
      RECT 91.04 4.388 91.075 4.595 ;
      RECT 90.997 4.383 91.04 4.583 ;
      RECT 90.911 4.374 90.997 4.592 ;
      RECT 90.825 4.363 90.911 4.604 ;
      RECT 90.76 4.354 90.825 4.613 ;
      RECT 90.74 4.345 90.76 4.618 ;
      RECT 90.735 4.338 90.74 4.62 ;
      RECT 90.695 4.323 90.735 4.617 ;
      RECT 90.675 4.302 90.695 4.612 ;
      RECT 90.66 4.29 90.675 4.605 ;
      RECT 90.655 4.282 90.66 4.598 ;
      RECT 90.64 4.262 90.655 4.591 ;
      RECT 90.635 4.125 90.64 4.585 ;
      RECT 90.555 4.014 90.635 4.557 ;
      RECT 90.546 4.007 90.555 4.523 ;
      RECT 90.46 4.001 90.546 4.448 ;
      RECT 90.435 3.992 90.46 4.36 ;
      RECT 90.405 3.987 90.435 4.335 ;
      RECT 90.34 3.996 90.405 4.32 ;
      RECT 90.32 4.012 90.34 4.295 ;
      RECT 90.31 4.018 90.32 4.243 ;
      RECT 90.29 4.04 90.31 4.125 ;
      RECT 90.945 4.072 91.17 4.19 ;
      RECT 90.945 3.915 91.165 4.19 ;
      RECT 90.16 4.683 90.225 5.126 ;
      RECT 90.1 4.708 90.225 5.124 ;
      RECT 90.1 4.708 90.28 5.118 ;
      RECT 90.085 4.733 90.28 5.117 ;
      RECT 90.225 4.67 90.3 5.114 ;
      RECT 90.16 4.695 90.38 5.108 ;
      RECT 90.085 4.734 90.425 5.102 ;
      RECT 90.07 4.761 90.425 5.093 ;
      RECT 90.085 4.754 90.445 5.085 ;
      RECT 90.07 4.763 90.45 5.068 ;
      RECT 90.065 4.78 90.45 4.895 ;
      RECT 90.07 3.502 90.105 3.74 ;
      RECT 90.07 3.502 90.135 3.739 ;
      RECT 90.07 3.502 90.25 3.735 ;
      RECT 90.07 3.502 90.305 3.713 ;
      RECT 90.08 3.445 90.36 3.613 ;
      RECT 90.185 3.285 90.215 3.736 ;
      RECT 90.215 3.28 90.395 3.493 ;
      RECT 90.085 3.421 90.395 3.493 ;
      RECT 90.135 3.317 90.185 3.737 ;
      RECT 90.105 3.373 90.395 3.493 ;
      RECT 88.965 7.455 89.135 8.925 ;
      RECT 88.965 7.455 89.14 8.715 ;
      RECT 88.595 9.405 89.065 9.575 ;
      RECT 88.595 8.385 88.765 9.575 ;
      RECT 88.59 3.035 88.76 4.225 ;
      RECT 88.59 3.035 89.06 3.205 ;
      RECT 87.975 3.895 88.15 5.155 ;
      RECT 87.975 3.685 88.145 5.155 ;
      RECT 87.975 7.455 88.145 8.925 ;
      RECT 87.975 7.455 88.15 8.715 ;
      RECT 87.605 3.035 87.775 4.225 ;
      RECT 87.605 3.035 88.075 3.205 ;
      RECT 87.605 9.405 88.075 9.575 ;
      RECT 87.605 8.385 87.775 9.575 ;
      RECT 86.615 4.015 86.79 5.155 ;
      RECT 86.615 1.865 86.785 5.155 ;
      RECT 86.615 1.865 86.79 2.415 ;
      RECT 86.615 10.195 86.79 10.745 ;
      RECT 86.615 7.455 86.785 10.745 ;
      RECT 86.615 7.455 86.79 8.595 ;
      RECT 86.185 3.895 86.36 5.155 ;
      RECT 86.185 2.945 86.355 5.155 ;
      RECT 86.185 7.455 86.355 9.665 ;
      RECT 86.185 7.455 86.36 8.715 ;
      RECT 85.755 3.925 85.925 5.155 ;
      RECT 85.815 2.145 85.985 4.095 ;
      RECT 85.755 1.865 85.925 2.315 ;
      RECT 85.755 10.295 85.925 10.745 ;
      RECT 85.815 8.515 85.985 10.465 ;
      RECT 85.755 7.455 85.925 8.685 ;
      RECT 85.23 3.895 85.405 5.155 ;
      RECT 85.23 1.865 85.4 5.155 ;
      RECT 85.23 3.365 85.64 3.695 ;
      RECT 85.23 2.525 85.64 2.855 ;
      RECT 85.23 1.865 85.405 2.355 ;
      RECT 85.23 10.255 85.405 10.745 ;
      RECT 85.23 7.455 85.4 10.745 ;
      RECT 85.23 9.755 85.64 10.085 ;
      RECT 85.23 8.915 85.64 9.245 ;
      RECT 85.23 7.455 85.405 8.715 ;
      RECT 83.345 4.687 83.36 4.738 ;
      RECT 83.34 4.667 83.345 4.785 ;
      RECT 83.325 4.657 83.34 4.853 ;
      RECT 83.3 4.637 83.325 4.908 ;
      RECT 83.26 4.622 83.3 4.928 ;
      RECT 83.215 4.616 83.26 4.956 ;
      RECT 83.145 4.606 83.215 4.973 ;
      RECT 83.125 4.598 83.145 4.973 ;
      RECT 83.065 4.592 83.125 4.965 ;
      RECT 83.006 4.583 83.065 4.953 ;
      RECT 82.92 4.572 83.006 4.936 ;
      RECT 82.898 4.563 82.92 4.924 ;
      RECT 82.812 4.556 82.898 4.911 ;
      RECT 82.726 4.543 82.812 4.892 ;
      RECT 82.64 4.531 82.726 4.872 ;
      RECT 82.61 4.52 82.64 4.859 ;
      RECT 82.56 4.506 82.61 4.851 ;
      RECT 82.54 4.495 82.56 4.843 ;
      RECT 82.491 4.484 82.54 4.835 ;
      RECT 82.405 4.463 82.491 4.82 ;
      RECT 82.36 4.45 82.405 4.805 ;
      RECT 82.315 4.45 82.36 4.785 ;
      RECT 82.26 4.45 82.315 4.72 ;
      RECT 82.235 4.45 82.26 4.643 ;
      RECT 82.76 4.187 82.93 4.37 ;
      RECT 82.76 4.187 82.945 4.328 ;
      RECT 82.76 4.187 82.95 4.27 ;
      RECT 82.82 3.955 82.955 4.246 ;
      RECT 82.82 3.959 82.96 4.229 ;
      RECT 82.765 4.122 82.96 4.229 ;
      RECT 82.79 3.967 82.93 4.37 ;
      RECT 82.79 3.971 82.97 4.17 ;
      RECT 82.775 4.057 82.97 4.17 ;
      RECT 82.785 3.987 82.93 4.37 ;
      RECT 82.785 3.99 82.98 4.083 ;
      RECT 82.78 4.007 82.98 4.083 ;
      RECT 82.55 3.227 82.72 3.71 ;
      RECT 82.545 3.222 82.695 3.7 ;
      RECT 82.545 3.229 82.725 3.694 ;
      RECT 82.535 3.223 82.695 3.673 ;
      RECT 82.535 3.239 82.74 3.632 ;
      RECT 82.505 3.224 82.695 3.595 ;
      RECT 82.505 3.254 82.75 3.535 ;
      RECT 82.5 3.226 82.695 3.533 ;
      RECT 82.48 3.235 82.725 3.49 ;
      RECT 82.455 3.251 82.74 3.402 ;
      RECT 82.455 3.27 82.765 3.393 ;
      RECT 82.45 3.307 82.765 3.345 ;
      RECT 82.455 3.287 82.77 3.313 ;
      RECT 82.55 3.221 82.66 3.71 ;
      RECT 82.636 3.22 82.66 3.71 ;
      RECT 81.87 4.005 81.875 4.216 ;
      RECT 82.47 4.005 82.475 4.19 ;
      RECT 82.535 4.045 82.54 4.158 ;
      RECT 82.53 4.037 82.535 4.164 ;
      RECT 82.525 4.027 82.53 4.172 ;
      RECT 82.52 4.017 82.525 4.181 ;
      RECT 82.515 4.007 82.52 4.185 ;
      RECT 82.475 4.005 82.515 4.188 ;
      RECT 82.447 4.004 82.47 4.192 ;
      RECT 82.361 4.001 82.447 4.199 ;
      RECT 82.275 3.997 82.361 4.21 ;
      RECT 82.255 3.995 82.275 4.216 ;
      RECT 82.237 3.994 82.255 4.219 ;
      RECT 82.151 3.992 82.237 4.226 ;
      RECT 82.065 3.987 82.151 4.239 ;
      RECT 82.046 3.984 82.065 4.244 ;
      RECT 81.96 3.982 82.046 4.235 ;
      RECT 81.95 3.982 81.96 4.228 ;
      RECT 81.875 3.995 81.95 4.222 ;
      RECT 81.86 4.006 81.87 4.216 ;
      RECT 81.85 4.008 81.86 4.215 ;
      RECT 81.84 4.012 81.85 4.211 ;
      RECT 81.835 4.015 81.84 4.205 ;
      RECT 81.825 4.017 81.835 4.199 ;
      RECT 81.82 4.02 81.825 4.193 ;
      RECT 81.855 10.195 82.03 10.745 ;
      RECT 81.855 7.455 82.025 10.745 ;
      RECT 81.855 7.455 82.03 8.595 ;
      RECT 81.8 4.606 81.805 4.81 ;
      RECT 81.785 4.593 81.8 4.903 ;
      RECT 81.77 4.574 81.785 5.18 ;
      RECT 81.735 4.54 81.77 5.18 ;
      RECT 81.731 4.51 81.735 5.18 ;
      RECT 81.645 4.392 81.731 5.18 ;
      RECT 81.635 4.267 81.645 5.18 ;
      RECT 81.62 4.235 81.635 5.18 ;
      RECT 81.615 4.21 81.62 5.18 ;
      RECT 81.61 4.2 81.615 5.136 ;
      RECT 81.595 4.172 81.61 5.041 ;
      RECT 81.58 4.138 81.595 4.94 ;
      RECT 81.575 4.116 81.58 4.893 ;
      RECT 81.57 4.105 81.575 4.863 ;
      RECT 81.565 4.095 81.57 4.829 ;
      RECT 81.555 4.082 81.565 4.797 ;
      RECT 81.53 4.058 81.555 4.723 ;
      RECT 81.525 4.038 81.53 4.648 ;
      RECT 81.52 4.032 81.525 4.623 ;
      RECT 81.515 4.027 81.52 4.588 ;
      RECT 81.51 4.022 81.515 4.563 ;
      RECT 81.505 4.02 81.51 4.543 ;
      RECT 81.5 4.02 81.505 4.528 ;
      RECT 81.495 4.02 81.5 4.488 ;
      RECT 81.485 4.02 81.495 4.46 ;
      RECT 81.475 4.02 81.485 4.405 ;
      RECT 81.46 4.02 81.475 4.343 ;
      RECT 81.455 4.019 81.46 4.288 ;
      RECT 81.44 4.018 81.455 4.268 ;
      RECT 81.38 4.016 81.44 4.242 ;
      RECT 81.345 4.017 81.38 4.222 ;
      RECT 81.34 4.019 81.345 4.212 ;
      RECT 81.33 4.038 81.34 4.202 ;
      RECT 81.325 4.065 81.33 4.133 ;
      RECT 81.44 3.49 81.61 3.735 ;
      RECT 81.475 3.261 81.61 3.735 ;
      RECT 81.475 3.263 81.62 3.73 ;
      RECT 81.475 3.265 81.645 3.718 ;
      RECT 81.475 3.268 81.67 3.7 ;
      RECT 81.475 3.273 81.72 3.673 ;
      RECT 81.475 3.278 81.74 3.638 ;
      RECT 81.455 3.28 81.75 3.613 ;
      RECT 81.445 3.375 81.75 3.613 ;
      RECT 81.475 3.26 81.585 3.735 ;
      RECT 81.485 3.257 81.58 3.735 ;
      RECT 81.425 7.455 81.595 9.665 ;
      RECT 81.425 7.455 81.6 8.715 ;
      RECT 81.005 4.522 81.195 4.88 ;
      RECT 81.005 4.534 81.23 4.879 ;
      RECT 81.005 4.562 81.25 4.877 ;
      RECT 81.005 4.587 81.255 4.876 ;
      RECT 81.005 4.645 81.27 4.875 ;
      RECT 80.99 4.518 81.15 4.86 ;
      RECT 80.97 4.527 81.195 4.813 ;
      RECT 80.945 4.538 81.23 4.75 ;
      RECT 80.945 4.622 81.265 4.75 ;
      RECT 80.945 4.597 81.26 4.75 ;
      RECT 81.005 4.513 81.15 4.88 ;
      RECT 81.091 4.512 81.15 4.88 ;
      RECT 81.091 4.511 81.135 4.88 ;
      RECT 80.47 10.255 80.645 10.745 ;
      RECT 80.47 7.455 80.64 10.745 ;
      RECT 80.47 9.755 80.88 10.085 ;
      RECT 80.47 8.915 80.88 9.245 ;
      RECT 80.47 7.455 80.645 8.715 ;
      RECT 80.79 4.027 80.795 4.405 ;
      RECT 80.785 3.995 80.79 4.405 ;
      RECT 80.78 3.967 80.785 4.405 ;
      RECT 80.775 3.947 80.78 4.405 ;
      RECT 80.72 3.93 80.775 4.405 ;
      RECT 80.68 3.915 80.72 4.405 ;
      RECT 80.625 3.902 80.68 4.405 ;
      RECT 80.59 3.893 80.625 4.405 ;
      RECT 80.586 3.891 80.59 4.404 ;
      RECT 80.5 3.887 80.586 4.387 ;
      RECT 80.415 3.879 80.5 4.35 ;
      RECT 80.405 3.875 80.415 4.323 ;
      RECT 80.395 3.875 80.405 4.305 ;
      RECT 80.385 3.877 80.395 4.288 ;
      RECT 80.38 3.882 80.385 4.274 ;
      RECT 80.375 3.886 80.38 4.261 ;
      RECT 80.365 3.891 80.375 4.245 ;
      RECT 80.35 3.905 80.365 4.22 ;
      RECT 80.345 3.911 80.35 4.2 ;
      RECT 80.34 3.913 80.345 4.193 ;
      RECT 80.335 3.917 80.34 4.068 ;
      RECT 80.515 4.717 80.76 5.18 ;
      RECT 80.435 4.69 80.755 5.176 ;
      RECT 80.365 4.725 80.76 5.169 ;
      RECT 80.155 4.98 80.76 5.165 ;
      RECT 80.335 4.748 80.76 5.165 ;
      RECT 80.175 4.94 80.76 5.165 ;
      RECT 80.325 4.76 80.76 5.165 ;
      RECT 80.21 4.877 80.76 5.165 ;
      RECT 80.265 4.802 80.76 5.165 ;
      RECT 80.515 4.667 80.755 5.18 ;
      RECT 80.545 4.66 80.755 5.18 ;
      RECT 80.535 4.662 80.755 5.18 ;
      RECT 80.545 4.657 80.675 5.18 ;
      RECT 80.1 3.22 80.186 3.659 ;
      RECT 80.095 3.22 80.186 3.657 ;
      RECT 80.095 3.22 80.255 3.656 ;
      RECT 80.095 3.22 80.285 3.653 ;
      RECT 80.08 3.227 80.285 3.644 ;
      RECT 80.08 3.227 80.29 3.64 ;
      RECT 80.075 3.237 80.29 3.633 ;
      RECT 80.07 3.242 80.29 3.608 ;
      RECT 80.07 3.242 80.305 3.59 ;
      RECT 80.095 3.22 80.325 3.505 ;
      RECT 80.065 3.247 80.325 3.503 ;
      RECT 80.075 3.24 80.33 3.441 ;
      RECT 80.065 3.362 80.335 3.424 ;
      RECT 80.05 3.257 80.33 3.375 ;
      RECT 80.045 3.267 80.33 3.275 ;
      RECT 80.125 4.038 80.13 4.115 ;
      RECT 80.115 4.032 80.125 4.305 ;
      RECT 80.105 4.024 80.115 4.326 ;
      RECT 80.095 4.015 80.105 4.348 ;
      RECT 80.09 4.01 80.095 4.365 ;
      RECT 80.05 4.01 80.09 4.405 ;
      RECT 80.03 4.01 80.05 4.46 ;
      RECT 80.025 4.01 80.03 4.488 ;
      RECT 80.015 4.01 80.025 4.503 ;
      RECT 79.98 4.01 80.015 4.545 ;
      RECT 79.975 4.01 79.98 4.588 ;
      RECT 79.965 4.01 79.975 4.603 ;
      RECT 79.95 4.01 79.965 4.623 ;
      RECT 79.935 4.01 79.95 4.65 ;
      RECT 79.93 4.011 79.935 4.668 ;
      RECT 79.91 4.012 79.93 4.675 ;
      RECT 79.855 4.013 79.91 4.695 ;
      RECT 79.845 4.014 79.855 4.709 ;
      RECT 79.84 4.017 79.845 4.708 ;
      RECT 79.8 4.09 79.84 4.706 ;
      RECT 79.785 4.17 79.8 4.704 ;
      RECT 79.76 4.225 79.785 4.702 ;
      RECT 79.745 4.29 79.76 4.701 ;
      RECT 79.7 4.322 79.745 4.698 ;
      RECT 79.615 4.345 79.7 4.693 ;
      RECT 79.59 4.365 79.615 4.688 ;
      RECT 79.52 4.37 79.59 4.684 ;
      RECT 79.5 4.372 79.52 4.681 ;
      RECT 79.415 4.383 79.5 4.675 ;
      RECT 79.41 4.394 79.415 4.67 ;
      RECT 79.4 4.396 79.41 4.67 ;
      RECT 79.365 4.4 79.4 4.668 ;
      RECT 79.315 4.41 79.365 4.655 ;
      RECT 79.295 4.418 79.315 4.64 ;
      RECT 79.215 4.43 79.295 4.623 ;
      RECT 79.38 3.98 79.55 4.19 ;
      RECT 79.496 3.976 79.55 4.19 ;
      RECT 79.301 3.98 79.55 4.181 ;
      RECT 79.301 3.98 79.555 4.17 ;
      RECT 79.215 3.98 79.555 4.161 ;
      RECT 79.215 3.988 79.565 4.105 ;
      RECT 79.215 4 79.57 4.018 ;
      RECT 79.215 4.007 79.575 4.01 ;
      RECT 79.41 3.978 79.55 4.19 ;
      RECT 79.165 4.923 79.41 5.255 ;
      RECT 79.16 4.915 79.165 5.252 ;
      RECT 79.13 4.935 79.41 5.233 ;
      RECT 79.11 4.967 79.41 5.206 ;
      RECT 79.16 4.92 79.337 5.252 ;
      RECT 79.16 4.917 79.251 5.252 ;
      RECT 79.1 3.265 79.27 3.685 ;
      RECT 79.095 3.265 79.27 3.683 ;
      RECT 79.095 3.265 79.295 3.673 ;
      RECT 79.095 3.265 79.315 3.648 ;
      RECT 79.09 3.265 79.315 3.643 ;
      RECT 79.09 3.265 79.325 3.633 ;
      RECT 79.09 3.265 79.33 3.628 ;
      RECT 79.09 3.27 79.335 3.623 ;
      RECT 79.09 3.302 79.35 3.613 ;
      RECT 79.09 3.372 79.375 3.596 ;
      RECT 79.07 3.372 79.375 3.588 ;
      RECT 79.07 3.432 79.385 3.565 ;
      RECT 79.07 3.472 79.395 3.51 ;
      RECT 79.055 3.265 79.33 3.49 ;
      RECT 79.045 3.28 79.335 3.388 ;
      RECT 78.635 4.67 78.805 5.195 ;
      RECT 78.63 4.67 78.805 5.188 ;
      RECT 78.62 4.67 78.81 5.153 ;
      RECT 78.615 4.68 78.81 5.125 ;
      RECT 78.61 4.7 78.81 5.108 ;
      RECT 78.62 4.675 78.815 5.098 ;
      RECT 78.605 4.72 78.815 5.09 ;
      RECT 78.6 4.74 78.815 5.075 ;
      RECT 78.595 4.77 78.815 5.065 ;
      RECT 78.585 4.815 78.815 5.04 ;
      RECT 78.615 4.685 78.82 5.023 ;
      RECT 78.58 4.867 78.82 5.018 ;
      RECT 78.615 4.695 78.825 4.988 ;
      RECT 78.575 4.9 78.825 4.985 ;
      RECT 78.57 4.925 78.825 4.965 ;
      RECT 78.61 4.712 78.835 4.905 ;
      RECT 78.605 4.734 78.845 4.798 ;
      RECT 78.555 3.981 78.57 4.25 ;
      RECT 78.51 3.965 78.555 4.295 ;
      RECT 78.505 3.953 78.51 4.345 ;
      RECT 78.495 3.949 78.505 4.378 ;
      RECT 78.49 3.946 78.495 4.406 ;
      RECT 78.475 3.948 78.49 4.448 ;
      RECT 78.47 3.952 78.475 4.488 ;
      RECT 78.45 3.957 78.47 4.54 ;
      RECT 78.446 3.962 78.45 4.597 ;
      RECT 78.36 3.981 78.446 4.634 ;
      RECT 78.35 4.002 78.36 4.67 ;
      RECT 78.345 4.01 78.35 4.671 ;
      RECT 78.34 4.052 78.345 4.672 ;
      RECT 78.325 4.14 78.34 4.673 ;
      RECT 78.315 4.29 78.325 4.675 ;
      RECT 78.31 4.335 78.315 4.677 ;
      RECT 78.275 4.377 78.31 4.68 ;
      RECT 78.27 4.395 78.275 4.683 ;
      RECT 78.193 4.401 78.27 4.689 ;
      RECT 78.107 4.415 78.193 4.702 ;
      RECT 78.021 4.429 78.107 4.716 ;
      RECT 77.935 4.443 78.021 4.729 ;
      RECT 77.875 4.455 77.935 4.741 ;
      RECT 77.85 4.462 77.875 4.748 ;
      RECT 77.836 4.465 77.85 4.753 ;
      RECT 77.75 4.473 77.836 4.769 ;
      RECT 77.745 4.48 77.75 4.784 ;
      RECT 77.721 4.48 77.745 4.791 ;
      RECT 77.635 4.483 77.721 4.819 ;
      RECT 77.55 4.487 77.635 4.863 ;
      RECT 77.485 4.491 77.55 4.9 ;
      RECT 77.46 4.494 77.485 4.916 ;
      RECT 77.385 4.507 77.46 4.92 ;
      RECT 77.36 4.525 77.385 4.924 ;
      RECT 77.35 4.532 77.36 4.926 ;
      RECT 77.335 4.535 77.35 4.927 ;
      RECT 77.275 4.547 77.335 4.931 ;
      RECT 77.265 4.561 77.275 4.935 ;
      RECT 77.21 4.571 77.265 4.923 ;
      RECT 77.185 4.592 77.21 4.906 ;
      RECT 77.165 4.612 77.185 4.897 ;
      RECT 77.16 4.625 77.165 4.892 ;
      RECT 77.145 4.637 77.16 4.888 ;
      RECT 78.38 3.292 78.385 3.315 ;
      RECT 78.375 3.283 78.38 3.355 ;
      RECT 78.37 3.281 78.375 3.398 ;
      RECT 78.365 3.272 78.37 3.433 ;
      RECT 78.36 3.262 78.365 3.505 ;
      RECT 78.355 3.252 78.36 3.57 ;
      RECT 78.35 3.249 78.355 3.61 ;
      RECT 78.325 3.243 78.35 3.7 ;
      RECT 78.29 3.231 78.325 3.725 ;
      RECT 78.28 3.222 78.29 3.725 ;
      RECT 78.145 3.22 78.155 3.708 ;
      RECT 78.135 3.22 78.145 3.675 ;
      RECT 78.13 3.22 78.135 3.65 ;
      RECT 78.125 3.22 78.13 3.638 ;
      RECT 78.12 3.22 78.125 3.62 ;
      RECT 78.11 3.22 78.12 3.585 ;
      RECT 78.105 3.222 78.11 3.563 ;
      RECT 78.1 3.228 78.105 3.548 ;
      RECT 78.095 3.234 78.1 3.533 ;
      RECT 78.08 3.246 78.095 3.506 ;
      RECT 78.075 3.257 78.08 3.474 ;
      RECT 78.07 3.267 78.075 3.458 ;
      RECT 78.06 3.275 78.07 3.427 ;
      RECT 78.055 3.285 78.06 3.401 ;
      RECT 78.05 3.342 78.055 3.384 ;
      RECT 78.155 3.22 78.28 3.725 ;
      RECT 77.87 3.907 78.13 4.205 ;
      RECT 77.865 3.914 78.13 4.203 ;
      RECT 77.87 3.909 78.145 4.198 ;
      RECT 77.86 3.922 78.145 4.195 ;
      RECT 77.86 3.927 78.15 4.188 ;
      RECT 77.855 3.935 78.15 4.185 ;
      RECT 77.855 3.952 78.155 3.983 ;
      RECT 77.87 3.904 78.101 4.205 ;
      RECT 77.925 3.903 78.101 4.205 ;
      RECT 77.925 3.9 78.015 4.205 ;
      RECT 77.925 3.897 78.011 4.205 ;
      RECT 77.615 4.17 77.62 4.183 ;
      RECT 77.61 4.137 77.615 4.188 ;
      RECT 77.605 4.092 77.61 4.195 ;
      RECT 77.6 4.047 77.605 4.203 ;
      RECT 77.595 4.015 77.6 4.211 ;
      RECT 77.59 3.975 77.595 4.212 ;
      RECT 77.575 3.955 77.59 4.214 ;
      RECT 77.5 3.937 77.575 4.226 ;
      RECT 77.49 3.93 77.5 4.237 ;
      RECT 77.485 3.93 77.49 4.239 ;
      RECT 77.455 3.936 77.485 4.243 ;
      RECT 77.415 3.949 77.455 4.243 ;
      RECT 77.39 3.96 77.415 4.229 ;
      RECT 77.375 3.966 77.39 4.212 ;
      RECT 77.365 3.968 77.375 4.203 ;
      RECT 77.36 3.969 77.365 4.198 ;
      RECT 77.355 3.97 77.36 4.193 ;
      RECT 77.35 3.971 77.355 4.19 ;
      RECT 77.325 3.976 77.35 4.18 ;
      RECT 77.315 3.992 77.325 4.167 ;
      RECT 77.31 4.012 77.315 4.162 ;
      RECT 77.32 3.405 77.325 3.601 ;
      RECT 77.305 3.369 77.32 3.603 ;
      RECT 77.295 3.351 77.305 3.608 ;
      RECT 77.285 3.337 77.295 3.612 ;
      RECT 77.24 3.321 77.285 3.622 ;
      RECT 77.235 3.311 77.24 3.631 ;
      RECT 77.19 3.3 77.235 3.637 ;
      RECT 77.185 3.288 77.19 3.644 ;
      RECT 77.17 3.283 77.185 3.648 ;
      RECT 77.155 3.275 77.17 3.653 ;
      RECT 77.145 3.268 77.155 3.658 ;
      RECT 77.135 3.265 77.145 3.663 ;
      RECT 77.125 3.265 77.135 3.664 ;
      RECT 77.12 3.262 77.125 3.663 ;
      RECT 77.085 3.257 77.11 3.662 ;
      RECT 77.061 3.253 77.085 3.661 ;
      RECT 76.975 3.244 77.061 3.658 ;
      RECT 76.96 3.236 76.975 3.655 ;
      RECT 76.938 3.235 76.96 3.654 ;
      RECT 76.852 3.235 76.938 3.652 ;
      RECT 76.766 3.235 76.852 3.65 ;
      RECT 76.68 3.235 76.766 3.647 ;
      RECT 76.67 3.235 76.68 3.638 ;
      RECT 76.64 3.235 76.67 3.598 ;
      RECT 76.63 3.245 76.64 3.553 ;
      RECT 76.625 3.285 76.63 3.538 ;
      RECT 76.62 3.3 76.625 3.525 ;
      RECT 76.59 3.38 76.62 3.487 ;
      RECT 77.11 3.26 77.12 3.663 ;
      RECT 76.935 4.025 76.95 4.63 ;
      RECT 76.94 4.02 76.95 4.63 ;
      RECT 77.105 4.02 77.11 4.203 ;
      RECT 77.095 4.02 77.105 4.233 ;
      RECT 77.08 4.02 77.095 4.293 ;
      RECT 77.075 4.02 77.08 4.338 ;
      RECT 77.07 4.02 77.075 4.368 ;
      RECT 77.065 4.02 77.07 4.388 ;
      RECT 77.055 4.02 77.065 4.423 ;
      RECT 77.04 4.02 77.055 4.455 ;
      RECT 76.995 4.02 77.04 4.483 ;
      RECT 76.99 4.02 76.995 4.513 ;
      RECT 76.985 4.02 76.99 4.525 ;
      RECT 76.98 4.02 76.985 4.533 ;
      RECT 76.97 4.02 76.98 4.548 ;
      RECT 76.965 4.02 76.97 4.57 ;
      RECT 76.955 4.02 76.965 4.593 ;
      RECT 76.95 4.02 76.955 4.613 ;
      RECT 76.915 4.035 76.935 4.63 ;
      RECT 76.89 4.052 76.915 4.63 ;
      RECT 76.885 4.062 76.89 4.63 ;
      RECT 76.855 4.077 76.885 4.63 ;
      RECT 76.78 4.119 76.855 4.63 ;
      RECT 76.775 4.15 76.78 4.613 ;
      RECT 76.77 4.154 76.775 4.595 ;
      RECT 76.765 4.158 76.77 4.558 ;
      RECT 76.76 4.342 76.765 4.525 ;
      RECT 76.245 4.531 76.331 5.096 ;
      RECT 76.2 4.533 76.365 5.09 ;
      RECT 76.331 4.53 76.365 5.09 ;
      RECT 76.245 4.532 76.45 5.084 ;
      RECT 76.2 4.542 76.46 5.08 ;
      RECT 76.175 4.534 76.45 5.076 ;
      RECT 76.17 4.537 76.45 5.071 ;
      RECT 76.145 4.552 76.46 5.065 ;
      RECT 76.145 4.577 76.5 5.06 ;
      RECT 76.105 4.585 76.5 5.035 ;
      RECT 76.105 4.612 76.515 5.033 ;
      RECT 76.105 4.642 76.525 5.02 ;
      RECT 76.1 4.787 76.525 5.008 ;
      RECT 76.105 4.716 76.545 5.005 ;
      RECT 76.105 4.773 76.55 4.813 ;
      RECT 76.295 4.052 76.465 4.23 ;
      RECT 76.245 3.991 76.295 4.215 ;
      RECT 75.98 3.971 76.245 4.2 ;
      RECT 75.94 4.035 76.415 4.2 ;
      RECT 75.94 4.025 76.37 4.2 ;
      RECT 75.94 4.022 76.36 4.2 ;
      RECT 75.94 4.01 76.35 4.2 ;
      RECT 75.94 3.995 76.295 4.2 ;
      RECT 75.98 3.967 76.181 4.2 ;
      RECT 75.99 3.945 76.181 4.2 ;
      RECT 76.015 3.93 76.095 4.2 ;
      RECT 75.77 4.46 75.89 4.905 ;
      RECT 75.755 4.46 75.89 4.904 ;
      RECT 75.71 4.482 75.89 4.899 ;
      RECT 75.67 4.531 75.89 4.893 ;
      RECT 75.67 4.531 75.895 4.868 ;
      RECT 75.67 4.531 75.915 4.758 ;
      RECT 75.665 4.561 75.915 4.755 ;
      RECT 75.755 4.46 75.925 4.65 ;
      RECT 75.415 3.245 75.42 3.69 ;
      RECT 75.225 3.245 75.245 3.655 ;
      RECT 75.195 3.245 75.2 3.63 ;
      RECT 75.875 3.552 75.89 3.74 ;
      RECT 75.87 3.537 75.875 3.746 ;
      RECT 75.85 3.51 75.87 3.749 ;
      RECT 75.8 3.477 75.85 3.758 ;
      RECT 75.77 3.457 75.8 3.762 ;
      RECT 75.751 3.445 75.77 3.758 ;
      RECT 75.665 3.417 75.751 3.748 ;
      RECT 75.655 3.392 75.665 3.738 ;
      RECT 75.585 3.36 75.655 3.73 ;
      RECT 75.56 3.32 75.585 3.722 ;
      RECT 75.54 3.302 75.56 3.716 ;
      RECT 75.53 3.292 75.54 3.713 ;
      RECT 75.52 3.285 75.53 3.711 ;
      RECT 75.5 3.272 75.52 3.708 ;
      RECT 75.49 3.262 75.5 3.705 ;
      RECT 75.48 3.255 75.49 3.703 ;
      RECT 75.43 3.247 75.48 3.697 ;
      RECT 75.42 3.245 75.43 3.691 ;
      RECT 75.39 3.245 75.415 3.688 ;
      RECT 75.361 3.245 75.39 3.683 ;
      RECT 75.275 3.245 75.361 3.673 ;
      RECT 75.245 3.245 75.275 3.66 ;
      RECT 75.2 3.245 75.225 3.643 ;
      RECT 75.185 3.245 75.195 3.625 ;
      RECT 75.165 3.252 75.185 3.61 ;
      RECT 75.16 3.267 75.165 3.598 ;
      RECT 75.155 3.272 75.16 3.538 ;
      RECT 75.15 3.277 75.155 3.38 ;
      RECT 75.145 3.28 75.15 3.298 ;
      RECT 74.885 4.57 74.92 4.89 ;
      RECT 75.47 4.755 75.475 4.937 ;
      RECT 75.425 4.637 75.47 4.956 ;
      RECT 75.41 4.614 75.425 4.979 ;
      RECT 75.4 4.604 75.41 4.989 ;
      RECT 75.38 4.599 75.4 5.002 ;
      RECT 75.355 4.597 75.38 5.023 ;
      RECT 75.336 4.596 75.355 5.035 ;
      RECT 75.25 4.593 75.336 5.035 ;
      RECT 75.18 4.588 75.25 5.023 ;
      RECT 75.105 4.584 75.18 4.998 ;
      RECT 75.04 4.58 75.105 4.965 ;
      RECT 74.97 4.577 75.04 4.925 ;
      RECT 74.94 4.573 74.97 4.9 ;
      RECT 74.92 4.571 74.94 4.893 ;
      RECT 74.836 4.569 74.885 4.891 ;
      RECT 74.75 4.566 74.836 4.892 ;
      RECT 74.675 4.565 74.75 4.894 ;
      RECT 74.59 4.565 74.675 4.92 ;
      RECT 74.513 4.566 74.59 4.945 ;
      RECT 74.427 4.567 74.513 4.945 ;
      RECT 74.341 4.567 74.427 4.945 ;
      RECT 74.255 4.568 74.341 4.945 ;
      RECT 74.235 4.569 74.255 4.937 ;
      RECT 74.22 4.575 74.235 4.922 ;
      RECT 74.185 4.595 74.22 4.902 ;
      RECT 74.175 4.615 74.185 4.884 ;
      RECT 75.145 3.92 75.15 4.19 ;
      RECT 75.14 3.911 75.145 4.195 ;
      RECT 75.13 3.901 75.14 4.207 ;
      RECT 75.125 3.89 75.13 4.218 ;
      RECT 75.105 3.884 75.125 4.236 ;
      RECT 75.06 3.881 75.105 4.285 ;
      RECT 75.045 3.88 75.06 4.33 ;
      RECT 75.04 3.88 75.045 4.343 ;
      RECT 75.03 3.88 75.04 4.355 ;
      RECT 75.025 3.881 75.03 4.37 ;
      RECT 75.005 3.889 75.025 4.375 ;
      RECT 74.975 3.905 75.005 4.375 ;
      RECT 74.965 3.917 74.97 4.375 ;
      RECT 74.93 3.932 74.965 4.375 ;
      RECT 74.9 3.952 74.93 4.375 ;
      RECT 74.89 3.977 74.9 4.375 ;
      RECT 74.885 4.005 74.89 4.375 ;
      RECT 74.88 4.035 74.885 4.375 ;
      RECT 74.875 4.052 74.88 4.375 ;
      RECT 74.865 4.08 74.875 4.375 ;
      RECT 74.855 4.115 74.865 4.375 ;
      RECT 74.85 4.15 74.855 4.375 ;
      RECT 74.97 3.915 74.975 4.375 ;
      RECT 73.96 3.245 73.965 3.644 ;
      RECT 73.705 3.245 73.74 3.642 ;
      RECT 73.3 3.28 73.305 3.636 ;
      RECT 74.045 3.283 74.05 3.538 ;
      RECT 74.04 3.281 74.045 3.544 ;
      RECT 74.035 3.28 74.04 3.551 ;
      RECT 74.01 3.273 74.035 3.575 ;
      RECT 74.005 3.266 74.01 3.599 ;
      RECT 74 3.262 74.005 3.608 ;
      RECT 73.99 3.257 74 3.621 ;
      RECT 73.985 3.254 73.99 3.63 ;
      RECT 73.98 3.252 73.985 3.635 ;
      RECT 73.965 3.248 73.98 3.645 ;
      RECT 73.95 3.242 73.96 3.644 ;
      RECT 73.912 3.24 73.95 3.644 ;
      RECT 73.826 3.242 73.912 3.644 ;
      RECT 73.74 3.244 73.826 3.643 ;
      RECT 73.669 3.245 73.705 3.642 ;
      RECT 73.583 3.247 73.669 3.642 ;
      RECT 73.497 3.249 73.583 3.641 ;
      RECT 73.411 3.251 73.497 3.641 ;
      RECT 73.325 3.254 73.411 3.64 ;
      RECT 73.315 3.26 73.325 3.639 ;
      RECT 73.305 3.272 73.315 3.637 ;
      RECT 73.245 3.307 73.3 3.633 ;
      RECT 73.24 3.337 73.245 3.395 ;
      RECT 73.585 4.552 73.59 4.809 ;
      RECT 73.565 4.471 73.585 4.826 ;
      RECT 73.545 4.465 73.565 4.855 ;
      RECT 73.485 4.452 73.545 4.875 ;
      RECT 73.44 4.436 73.485 4.876 ;
      RECT 73.356 4.424 73.44 4.864 ;
      RECT 73.27 4.411 73.356 4.848 ;
      RECT 73.26 4.404 73.27 4.84 ;
      RECT 73.215 4.401 73.26 4.78 ;
      RECT 73.195 4.397 73.215 4.695 ;
      RECT 73.18 4.395 73.195 4.648 ;
      RECT 73.15 4.392 73.18 4.618 ;
      RECT 73.115 4.388 73.15 4.595 ;
      RECT 73.072 4.383 73.115 4.583 ;
      RECT 72.986 4.374 73.072 4.592 ;
      RECT 72.9 4.363 72.986 4.604 ;
      RECT 72.835 4.354 72.9 4.613 ;
      RECT 72.815 4.345 72.835 4.618 ;
      RECT 72.81 4.338 72.815 4.62 ;
      RECT 72.77 4.323 72.81 4.617 ;
      RECT 72.75 4.302 72.77 4.612 ;
      RECT 72.735 4.29 72.75 4.605 ;
      RECT 72.73 4.282 72.735 4.598 ;
      RECT 72.715 4.262 72.73 4.591 ;
      RECT 72.71 4.125 72.715 4.585 ;
      RECT 72.63 4.014 72.71 4.557 ;
      RECT 72.621 4.007 72.63 4.523 ;
      RECT 72.535 4.001 72.621 4.448 ;
      RECT 72.51 3.992 72.535 4.36 ;
      RECT 72.48 3.987 72.51 4.335 ;
      RECT 72.415 3.996 72.48 4.32 ;
      RECT 72.395 4.012 72.415 4.295 ;
      RECT 72.385 4.018 72.395 4.243 ;
      RECT 72.365 4.04 72.385 4.125 ;
      RECT 73.02 4.072 73.245 4.19 ;
      RECT 73.02 3.915 73.24 4.19 ;
      RECT 72.235 4.683 72.3 5.126 ;
      RECT 72.175 4.708 72.3 5.124 ;
      RECT 72.175 4.708 72.355 5.118 ;
      RECT 72.16 4.733 72.355 5.117 ;
      RECT 72.3 4.67 72.375 5.114 ;
      RECT 72.235 4.695 72.455 5.108 ;
      RECT 72.16 4.734 72.5 5.102 ;
      RECT 72.145 4.761 72.5 5.093 ;
      RECT 72.16 4.754 72.52 5.085 ;
      RECT 72.145 4.763 72.525 5.068 ;
      RECT 72.14 4.78 72.525 4.895 ;
      RECT 72.145 3.502 72.18 3.74 ;
      RECT 72.145 3.502 72.21 3.739 ;
      RECT 72.145 3.502 72.325 3.735 ;
      RECT 72.145 3.502 72.38 3.713 ;
      RECT 72.155 3.445 72.435 3.613 ;
      RECT 72.26 3.285 72.29 3.736 ;
      RECT 72.29 3.28 72.47 3.493 ;
      RECT 72.16 3.421 72.47 3.493 ;
      RECT 72.21 3.317 72.26 3.737 ;
      RECT 72.18 3.373 72.47 3.493 ;
      RECT 71.04 7.455 71.21 8.925 ;
      RECT 71.04 7.455 71.215 8.715 ;
      RECT 70.67 9.405 71.14 9.575 ;
      RECT 70.67 8.385 70.84 9.575 ;
      RECT 70.665 3.035 70.835 4.225 ;
      RECT 70.665 3.035 71.135 3.205 ;
      RECT 70.05 3.895 70.225 5.155 ;
      RECT 70.05 3.685 70.22 5.155 ;
      RECT 70.05 7.455 70.22 8.925 ;
      RECT 70.05 7.455 70.225 8.715 ;
      RECT 69.68 3.035 69.85 4.225 ;
      RECT 69.68 3.035 70.15 3.205 ;
      RECT 69.68 9.405 70.15 9.575 ;
      RECT 69.68 8.385 69.85 9.575 ;
      RECT 68.69 4.015 68.865 5.155 ;
      RECT 68.69 1.865 68.86 5.155 ;
      RECT 68.69 1.865 68.865 2.415 ;
      RECT 68.69 10.195 68.865 10.745 ;
      RECT 68.69 7.455 68.86 10.745 ;
      RECT 68.69 7.455 68.865 8.595 ;
      RECT 68.26 3.895 68.435 5.155 ;
      RECT 68.26 2.945 68.43 5.155 ;
      RECT 68.26 7.455 68.43 9.665 ;
      RECT 68.26 7.455 68.435 8.715 ;
      RECT 67.83 3.925 68 5.155 ;
      RECT 67.89 2.145 68.06 4.095 ;
      RECT 67.83 1.865 68 2.315 ;
      RECT 67.83 10.295 68 10.745 ;
      RECT 67.89 8.515 68.06 10.465 ;
      RECT 67.83 7.455 68 8.685 ;
      RECT 67.305 3.895 67.48 5.155 ;
      RECT 67.305 1.865 67.475 5.155 ;
      RECT 67.305 3.365 67.715 3.695 ;
      RECT 67.305 2.525 67.715 2.855 ;
      RECT 67.305 1.865 67.48 2.355 ;
      RECT 67.305 10.255 67.48 10.745 ;
      RECT 67.305 7.455 67.475 10.745 ;
      RECT 67.305 9.755 67.715 10.085 ;
      RECT 67.305 8.915 67.715 9.245 ;
      RECT 67.305 7.455 67.48 8.715 ;
      RECT 65.42 4.687 65.435 4.738 ;
      RECT 65.415 4.667 65.42 4.785 ;
      RECT 65.4 4.657 65.415 4.853 ;
      RECT 65.375 4.637 65.4 4.908 ;
      RECT 65.335 4.622 65.375 4.928 ;
      RECT 65.29 4.616 65.335 4.956 ;
      RECT 65.22 4.606 65.29 4.973 ;
      RECT 65.2 4.598 65.22 4.973 ;
      RECT 65.14 4.592 65.2 4.965 ;
      RECT 65.081 4.583 65.14 4.953 ;
      RECT 64.995 4.572 65.081 4.936 ;
      RECT 64.973 4.563 64.995 4.924 ;
      RECT 64.887 4.556 64.973 4.911 ;
      RECT 64.801 4.543 64.887 4.892 ;
      RECT 64.715 4.531 64.801 4.872 ;
      RECT 64.685 4.52 64.715 4.859 ;
      RECT 64.635 4.506 64.685 4.851 ;
      RECT 64.615 4.495 64.635 4.843 ;
      RECT 64.566 4.484 64.615 4.835 ;
      RECT 64.48 4.463 64.566 4.82 ;
      RECT 64.435 4.45 64.48 4.805 ;
      RECT 64.39 4.45 64.435 4.785 ;
      RECT 64.335 4.45 64.39 4.72 ;
      RECT 64.31 4.45 64.335 4.643 ;
      RECT 64.835 4.187 65.005 4.37 ;
      RECT 64.835 4.187 65.02 4.328 ;
      RECT 64.835 4.187 65.025 4.27 ;
      RECT 64.895 3.955 65.03 4.246 ;
      RECT 64.895 3.959 65.035 4.229 ;
      RECT 64.84 4.122 65.035 4.229 ;
      RECT 64.865 3.967 65.005 4.37 ;
      RECT 64.865 3.971 65.045 4.17 ;
      RECT 64.85 4.057 65.045 4.17 ;
      RECT 64.86 3.987 65.005 4.37 ;
      RECT 64.86 3.99 65.055 4.083 ;
      RECT 64.855 4.007 65.055 4.083 ;
      RECT 64.625 3.227 64.795 3.71 ;
      RECT 64.62 3.222 64.77 3.7 ;
      RECT 64.62 3.229 64.8 3.694 ;
      RECT 64.61 3.223 64.77 3.673 ;
      RECT 64.61 3.239 64.815 3.632 ;
      RECT 64.58 3.224 64.77 3.595 ;
      RECT 64.58 3.254 64.825 3.535 ;
      RECT 64.575 3.226 64.77 3.533 ;
      RECT 64.555 3.235 64.8 3.49 ;
      RECT 64.53 3.251 64.815 3.402 ;
      RECT 64.53 3.27 64.84 3.393 ;
      RECT 64.525 3.307 64.84 3.345 ;
      RECT 64.53 3.287 64.845 3.313 ;
      RECT 64.625 3.221 64.735 3.71 ;
      RECT 64.711 3.22 64.735 3.71 ;
      RECT 63.945 4.005 63.95 4.216 ;
      RECT 64.545 4.005 64.55 4.19 ;
      RECT 64.61 4.045 64.615 4.158 ;
      RECT 64.605 4.037 64.61 4.164 ;
      RECT 64.6 4.027 64.605 4.172 ;
      RECT 64.595 4.017 64.6 4.181 ;
      RECT 64.59 4.007 64.595 4.185 ;
      RECT 64.55 4.005 64.59 4.188 ;
      RECT 64.522 4.004 64.545 4.192 ;
      RECT 64.436 4.001 64.522 4.199 ;
      RECT 64.35 3.997 64.436 4.21 ;
      RECT 64.33 3.995 64.35 4.216 ;
      RECT 64.312 3.994 64.33 4.219 ;
      RECT 64.226 3.992 64.312 4.226 ;
      RECT 64.14 3.987 64.226 4.239 ;
      RECT 64.121 3.984 64.14 4.244 ;
      RECT 64.035 3.982 64.121 4.235 ;
      RECT 64.025 3.982 64.035 4.228 ;
      RECT 63.95 3.995 64.025 4.222 ;
      RECT 63.935 4.006 63.945 4.216 ;
      RECT 63.925 4.008 63.935 4.215 ;
      RECT 63.915 4.012 63.925 4.211 ;
      RECT 63.91 4.015 63.915 4.205 ;
      RECT 63.9 4.017 63.91 4.199 ;
      RECT 63.895 4.02 63.9 4.193 ;
      RECT 63.93 10.195 64.105 10.745 ;
      RECT 63.93 7.455 64.1 10.745 ;
      RECT 63.93 7.455 64.105 8.595 ;
      RECT 63.875 4.606 63.88 4.81 ;
      RECT 63.86 4.593 63.875 4.903 ;
      RECT 63.845 4.574 63.86 5.18 ;
      RECT 63.81 4.54 63.845 5.18 ;
      RECT 63.806 4.51 63.81 5.18 ;
      RECT 63.72 4.392 63.806 5.18 ;
      RECT 63.71 4.267 63.72 5.18 ;
      RECT 63.695 4.235 63.71 5.18 ;
      RECT 63.69 4.21 63.695 5.18 ;
      RECT 63.685 4.2 63.69 5.136 ;
      RECT 63.67 4.172 63.685 5.041 ;
      RECT 63.655 4.138 63.67 4.94 ;
      RECT 63.65 4.116 63.655 4.893 ;
      RECT 63.645 4.105 63.65 4.863 ;
      RECT 63.64 4.095 63.645 4.829 ;
      RECT 63.63 4.082 63.64 4.797 ;
      RECT 63.605 4.058 63.63 4.723 ;
      RECT 63.6 4.038 63.605 4.648 ;
      RECT 63.595 4.032 63.6 4.623 ;
      RECT 63.59 4.027 63.595 4.588 ;
      RECT 63.585 4.022 63.59 4.563 ;
      RECT 63.58 4.02 63.585 4.543 ;
      RECT 63.575 4.02 63.58 4.528 ;
      RECT 63.57 4.02 63.575 4.488 ;
      RECT 63.56 4.02 63.57 4.46 ;
      RECT 63.55 4.02 63.56 4.405 ;
      RECT 63.535 4.02 63.55 4.343 ;
      RECT 63.53 4.019 63.535 4.288 ;
      RECT 63.515 4.018 63.53 4.268 ;
      RECT 63.455 4.016 63.515 4.242 ;
      RECT 63.42 4.017 63.455 4.222 ;
      RECT 63.415 4.019 63.42 4.212 ;
      RECT 63.405 4.038 63.415 4.202 ;
      RECT 63.4 4.065 63.405 4.133 ;
      RECT 63.515 3.49 63.685 3.735 ;
      RECT 63.55 3.261 63.685 3.735 ;
      RECT 63.55 3.263 63.695 3.73 ;
      RECT 63.55 3.265 63.72 3.718 ;
      RECT 63.55 3.268 63.745 3.7 ;
      RECT 63.55 3.273 63.795 3.673 ;
      RECT 63.55 3.278 63.815 3.638 ;
      RECT 63.53 3.28 63.825 3.613 ;
      RECT 63.52 3.375 63.825 3.613 ;
      RECT 63.55 3.26 63.66 3.735 ;
      RECT 63.56 3.257 63.655 3.735 ;
      RECT 63.5 7.455 63.67 9.665 ;
      RECT 63.5 7.455 63.675 8.715 ;
      RECT 63.08 4.522 63.27 4.88 ;
      RECT 63.08 4.534 63.305 4.879 ;
      RECT 63.08 4.562 63.325 4.877 ;
      RECT 63.08 4.587 63.33 4.876 ;
      RECT 63.08 4.645 63.345 4.875 ;
      RECT 63.065 4.518 63.225 4.86 ;
      RECT 63.045 4.527 63.27 4.813 ;
      RECT 63.02 4.538 63.305 4.75 ;
      RECT 63.02 4.622 63.34 4.75 ;
      RECT 63.02 4.597 63.335 4.75 ;
      RECT 63.08 4.513 63.225 4.88 ;
      RECT 63.166 4.512 63.225 4.88 ;
      RECT 63.166 4.511 63.21 4.88 ;
      RECT 62.545 10.255 62.72 10.745 ;
      RECT 62.545 7.455 62.715 10.745 ;
      RECT 62.545 9.755 62.955 10.085 ;
      RECT 62.545 8.915 62.955 9.245 ;
      RECT 62.545 7.455 62.72 8.715 ;
      RECT 62.865 4.027 62.87 4.405 ;
      RECT 62.86 3.995 62.865 4.405 ;
      RECT 62.855 3.967 62.86 4.405 ;
      RECT 62.85 3.947 62.855 4.405 ;
      RECT 62.795 3.93 62.85 4.405 ;
      RECT 62.755 3.915 62.795 4.405 ;
      RECT 62.7 3.902 62.755 4.405 ;
      RECT 62.665 3.893 62.7 4.405 ;
      RECT 62.661 3.891 62.665 4.404 ;
      RECT 62.575 3.887 62.661 4.387 ;
      RECT 62.49 3.879 62.575 4.35 ;
      RECT 62.48 3.875 62.49 4.323 ;
      RECT 62.47 3.875 62.48 4.305 ;
      RECT 62.46 3.877 62.47 4.288 ;
      RECT 62.455 3.882 62.46 4.274 ;
      RECT 62.45 3.886 62.455 4.261 ;
      RECT 62.44 3.891 62.45 4.245 ;
      RECT 62.425 3.905 62.44 4.22 ;
      RECT 62.42 3.911 62.425 4.2 ;
      RECT 62.415 3.913 62.42 4.193 ;
      RECT 62.41 3.917 62.415 4.068 ;
      RECT 62.59 4.717 62.835 5.18 ;
      RECT 62.51 4.69 62.83 5.176 ;
      RECT 62.44 4.725 62.835 5.169 ;
      RECT 62.23 4.98 62.835 5.165 ;
      RECT 62.41 4.748 62.835 5.165 ;
      RECT 62.25 4.94 62.835 5.165 ;
      RECT 62.4 4.76 62.835 5.165 ;
      RECT 62.285 4.877 62.835 5.165 ;
      RECT 62.34 4.802 62.835 5.165 ;
      RECT 62.59 4.667 62.83 5.18 ;
      RECT 62.62 4.66 62.83 5.18 ;
      RECT 62.61 4.662 62.83 5.18 ;
      RECT 62.62 4.657 62.75 5.18 ;
      RECT 62.175 3.22 62.261 3.659 ;
      RECT 62.17 3.22 62.261 3.657 ;
      RECT 62.17 3.22 62.33 3.656 ;
      RECT 62.17 3.22 62.36 3.653 ;
      RECT 62.155 3.227 62.36 3.644 ;
      RECT 62.155 3.227 62.365 3.64 ;
      RECT 62.15 3.237 62.365 3.633 ;
      RECT 62.145 3.242 62.365 3.608 ;
      RECT 62.145 3.242 62.38 3.59 ;
      RECT 62.17 3.22 62.4 3.505 ;
      RECT 62.14 3.247 62.4 3.503 ;
      RECT 62.15 3.24 62.405 3.441 ;
      RECT 62.14 3.362 62.41 3.424 ;
      RECT 62.125 3.257 62.405 3.375 ;
      RECT 62.12 3.267 62.405 3.275 ;
      RECT 62.2 4.038 62.205 4.115 ;
      RECT 62.19 4.032 62.2 4.305 ;
      RECT 62.18 4.024 62.19 4.326 ;
      RECT 62.17 4.015 62.18 4.348 ;
      RECT 62.165 4.01 62.17 4.365 ;
      RECT 62.125 4.01 62.165 4.405 ;
      RECT 62.105 4.01 62.125 4.46 ;
      RECT 62.1 4.01 62.105 4.488 ;
      RECT 62.09 4.01 62.1 4.503 ;
      RECT 62.055 4.01 62.09 4.545 ;
      RECT 62.05 4.01 62.055 4.588 ;
      RECT 62.04 4.01 62.05 4.603 ;
      RECT 62.025 4.01 62.04 4.623 ;
      RECT 62.01 4.01 62.025 4.65 ;
      RECT 62.005 4.011 62.01 4.668 ;
      RECT 61.985 4.012 62.005 4.675 ;
      RECT 61.93 4.013 61.985 4.695 ;
      RECT 61.92 4.014 61.93 4.709 ;
      RECT 61.915 4.017 61.92 4.708 ;
      RECT 61.875 4.09 61.915 4.706 ;
      RECT 61.86 4.17 61.875 4.704 ;
      RECT 61.835 4.225 61.86 4.702 ;
      RECT 61.82 4.29 61.835 4.701 ;
      RECT 61.775 4.322 61.82 4.698 ;
      RECT 61.69 4.345 61.775 4.693 ;
      RECT 61.665 4.365 61.69 4.688 ;
      RECT 61.595 4.37 61.665 4.684 ;
      RECT 61.575 4.372 61.595 4.681 ;
      RECT 61.49 4.383 61.575 4.675 ;
      RECT 61.485 4.394 61.49 4.67 ;
      RECT 61.475 4.396 61.485 4.67 ;
      RECT 61.44 4.4 61.475 4.668 ;
      RECT 61.39 4.41 61.44 4.655 ;
      RECT 61.37 4.418 61.39 4.64 ;
      RECT 61.29 4.43 61.37 4.623 ;
      RECT 61.455 3.98 61.625 4.19 ;
      RECT 61.571 3.976 61.625 4.19 ;
      RECT 61.376 3.98 61.625 4.181 ;
      RECT 61.376 3.98 61.63 4.17 ;
      RECT 61.29 3.98 61.63 4.161 ;
      RECT 61.29 3.988 61.64 4.105 ;
      RECT 61.29 4 61.645 4.018 ;
      RECT 61.29 4.007 61.65 4.01 ;
      RECT 61.485 3.978 61.625 4.19 ;
      RECT 61.24 4.923 61.485 5.255 ;
      RECT 61.235 4.915 61.24 5.252 ;
      RECT 61.205 4.935 61.485 5.233 ;
      RECT 61.185 4.967 61.485 5.206 ;
      RECT 61.235 4.92 61.412 5.252 ;
      RECT 61.235 4.917 61.326 5.252 ;
      RECT 61.175 3.265 61.345 3.685 ;
      RECT 61.17 3.265 61.345 3.683 ;
      RECT 61.17 3.265 61.37 3.673 ;
      RECT 61.17 3.265 61.39 3.648 ;
      RECT 61.165 3.265 61.39 3.643 ;
      RECT 61.165 3.265 61.4 3.633 ;
      RECT 61.165 3.265 61.405 3.628 ;
      RECT 61.165 3.27 61.41 3.623 ;
      RECT 61.165 3.302 61.425 3.613 ;
      RECT 61.165 3.372 61.45 3.596 ;
      RECT 61.145 3.372 61.45 3.588 ;
      RECT 61.145 3.432 61.46 3.565 ;
      RECT 61.145 3.472 61.47 3.51 ;
      RECT 61.13 3.265 61.405 3.49 ;
      RECT 61.12 3.28 61.41 3.388 ;
      RECT 60.71 4.67 60.88 5.195 ;
      RECT 60.705 4.67 60.88 5.188 ;
      RECT 60.695 4.67 60.885 5.153 ;
      RECT 60.69 4.68 60.885 5.125 ;
      RECT 60.685 4.7 60.885 5.108 ;
      RECT 60.695 4.675 60.89 5.098 ;
      RECT 60.68 4.72 60.89 5.09 ;
      RECT 60.675 4.74 60.89 5.075 ;
      RECT 60.67 4.77 60.89 5.065 ;
      RECT 60.66 4.815 60.89 5.04 ;
      RECT 60.69 4.685 60.895 5.023 ;
      RECT 60.655 4.867 60.895 5.018 ;
      RECT 60.69 4.695 60.9 4.988 ;
      RECT 60.65 4.9 60.9 4.985 ;
      RECT 60.645 4.925 60.9 4.965 ;
      RECT 60.685 4.712 60.91 4.905 ;
      RECT 60.68 4.734 60.92 4.798 ;
      RECT 60.63 3.981 60.645 4.25 ;
      RECT 60.585 3.965 60.63 4.295 ;
      RECT 60.58 3.953 60.585 4.345 ;
      RECT 60.57 3.949 60.58 4.378 ;
      RECT 60.565 3.946 60.57 4.406 ;
      RECT 60.55 3.948 60.565 4.448 ;
      RECT 60.545 3.952 60.55 4.488 ;
      RECT 60.525 3.957 60.545 4.54 ;
      RECT 60.521 3.962 60.525 4.597 ;
      RECT 60.435 3.981 60.521 4.634 ;
      RECT 60.425 4.002 60.435 4.67 ;
      RECT 60.42 4.01 60.425 4.671 ;
      RECT 60.415 4.052 60.42 4.672 ;
      RECT 60.4 4.14 60.415 4.673 ;
      RECT 60.39 4.29 60.4 4.675 ;
      RECT 60.385 4.335 60.39 4.677 ;
      RECT 60.35 4.377 60.385 4.68 ;
      RECT 60.345 4.395 60.35 4.683 ;
      RECT 60.268 4.401 60.345 4.689 ;
      RECT 60.182 4.415 60.268 4.702 ;
      RECT 60.096 4.429 60.182 4.716 ;
      RECT 60.01 4.443 60.096 4.729 ;
      RECT 59.95 4.455 60.01 4.741 ;
      RECT 59.925 4.462 59.95 4.748 ;
      RECT 59.911 4.465 59.925 4.753 ;
      RECT 59.825 4.473 59.911 4.769 ;
      RECT 59.82 4.48 59.825 4.784 ;
      RECT 59.796 4.48 59.82 4.791 ;
      RECT 59.71 4.483 59.796 4.819 ;
      RECT 59.625 4.487 59.71 4.863 ;
      RECT 59.56 4.491 59.625 4.9 ;
      RECT 59.535 4.494 59.56 4.916 ;
      RECT 59.46 4.507 59.535 4.92 ;
      RECT 59.435 4.525 59.46 4.924 ;
      RECT 59.425 4.532 59.435 4.926 ;
      RECT 59.41 4.535 59.425 4.927 ;
      RECT 59.35 4.547 59.41 4.931 ;
      RECT 59.34 4.561 59.35 4.935 ;
      RECT 59.285 4.571 59.34 4.923 ;
      RECT 59.26 4.592 59.285 4.906 ;
      RECT 59.24 4.612 59.26 4.897 ;
      RECT 59.235 4.625 59.24 4.892 ;
      RECT 59.22 4.637 59.235 4.888 ;
      RECT 60.455 3.292 60.46 3.315 ;
      RECT 60.45 3.283 60.455 3.355 ;
      RECT 60.445 3.281 60.45 3.398 ;
      RECT 60.44 3.272 60.445 3.433 ;
      RECT 60.435 3.262 60.44 3.505 ;
      RECT 60.43 3.252 60.435 3.57 ;
      RECT 60.425 3.249 60.43 3.61 ;
      RECT 60.4 3.243 60.425 3.7 ;
      RECT 60.365 3.231 60.4 3.725 ;
      RECT 60.355 3.222 60.365 3.725 ;
      RECT 60.22 3.22 60.23 3.708 ;
      RECT 60.21 3.22 60.22 3.675 ;
      RECT 60.205 3.22 60.21 3.65 ;
      RECT 60.2 3.22 60.205 3.638 ;
      RECT 60.195 3.22 60.2 3.62 ;
      RECT 60.185 3.22 60.195 3.585 ;
      RECT 60.18 3.222 60.185 3.563 ;
      RECT 60.175 3.228 60.18 3.548 ;
      RECT 60.17 3.234 60.175 3.533 ;
      RECT 60.155 3.246 60.17 3.506 ;
      RECT 60.15 3.257 60.155 3.474 ;
      RECT 60.145 3.267 60.15 3.458 ;
      RECT 60.135 3.275 60.145 3.427 ;
      RECT 60.13 3.285 60.135 3.401 ;
      RECT 60.125 3.342 60.13 3.384 ;
      RECT 60.23 3.22 60.355 3.725 ;
      RECT 59.945 3.907 60.205 4.205 ;
      RECT 59.94 3.914 60.205 4.203 ;
      RECT 59.945 3.909 60.22 4.198 ;
      RECT 59.935 3.922 60.22 4.195 ;
      RECT 59.935 3.927 60.225 4.188 ;
      RECT 59.93 3.935 60.225 4.185 ;
      RECT 59.93 3.952 60.23 3.983 ;
      RECT 59.945 3.904 60.176 4.205 ;
      RECT 60 3.903 60.176 4.205 ;
      RECT 60 3.9 60.09 4.205 ;
      RECT 60 3.897 60.086 4.205 ;
      RECT 59.69 4.17 59.695 4.183 ;
      RECT 59.685 4.137 59.69 4.188 ;
      RECT 59.68 4.092 59.685 4.195 ;
      RECT 59.675 4.047 59.68 4.203 ;
      RECT 59.67 4.015 59.675 4.211 ;
      RECT 59.665 3.975 59.67 4.212 ;
      RECT 59.65 3.955 59.665 4.214 ;
      RECT 59.575 3.937 59.65 4.226 ;
      RECT 59.565 3.93 59.575 4.237 ;
      RECT 59.56 3.93 59.565 4.239 ;
      RECT 59.53 3.936 59.56 4.243 ;
      RECT 59.49 3.949 59.53 4.243 ;
      RECT 59.465 3.96 59.49 4.229 ;
      RECT 59.45 3.966 59.465 4.212 ;
      RECT 59.44 3.968 59.45 4.203 ;
      RECT 59.435 3.969 59.44 4.198 ;
      RECT 59.43 3.97 59.435 4.193 ;
      RECT 59.425 3.971 59.43 4.19 ;
      RECT 59.4 3.976 59.425 4.18 ;
      RECT 59.39 3.992 59.4 4.167 ;
      RECT 59.385 4.012 59.39 4.162 ;
      RECT 59.395 3.405 59.4 3.601 ;
      RECT 59.38 3.369 59.395 3.603 ;
      RECT 59.37 3.351 59.38 3.608 ;
      RECT 59.36 3.337 59.37 3.612 ;
      RECT 59.315 3.321 59.36 3.622 ;
      RECT 59.31 3.311 59.315 3.631 ;
      RECT 59.265 3.3 59.31 3.637 ;
      RECT 59.26 3.288 59.265 3.644 ;
      RECT 59.245 3.283 59.26 3.648 ;
      RECT 59.23 3.275 59.245 3.653 ;
      RECT 59.22 3.268 59.23 3.658 ;
      RECT 59.21 3.265 59.22 3.663 ;
      RECT 59.2 3.265 59.21 3.664 ;
      RECT 59.195 3.262 59.2 3.663 ;
      RECT 59.16 3.257 59.185 3.662 ;
      RECT 59.136 3.253 59.16 3.661 ;
      RECT 59.05 3.244 59.136 3.658 ;
      RECT 59.035 3.236 59.05 3.655 ;
      RECT 59.013 3.235 59.035 3.654 ;
      RECT 58.927 3.235 59.013 3.652 ;
      RECT 58.841 3.235 58.927 3.65 ;
      RECT 58.755 3.235 58.841 3.647 ;
      RECT 58.745 3.235 58.755 3.638 ;
      RECT 58.715 3.235 58.745 3.598 ;
      RECT 58.705 3.245 58.715 3.553 ;
      RECT 58.7 3.285 58.705 3.538 ;
      RECT 58.695 3.3 58.7 3.525 ;
      RECT 58.665 3.38 58.695 3.487 ;
      RECT 59.185 3.26 59.195 3.663 ;
      RECT 59.01 4.025 59.025 4.63 ;
      RECT 59.015 4.02 59.025 4.63 ;
      RECT 59.18 4.02 59.185 4.203 ;
      RECT 59.17 4.02 59.18 4.233 ;
      RECT 59.155 4.02 59.17 4.293 ;
      RECT 59.15 4.02 59.155 4.338 ;
      RECT 59.145 4.02 59.15 4.368 ;
      RECT 59.14 4.02 59.145 4.388 ;
      RECT 59.13 4.02 59.14 4.423 ;
      RECT 59.115 4.02 59.13 4.455 ;
      RECT 59.07 4.02 59.115 4.483 ;
      RECT 59.065 4.02 59.07 4.513 ;
      RECT 59.06 4.02 59.065 4.525 ;
      RECT 59.055 4.02 59.06 4.533 ;
      RECT 59.045 4.02 59.055 4.548 ;
      RECT 59.04 4.02 59.045 4.57 ;
      RECT 59.03 4.02 59.04 4.593 ;
      RECT 59.025 4.02 59.03 4.613 ;
      RECT 58.99 4.035 59.01 4.63 ;
      RECT 58.965 4.052 58.99 4.63 ;
      RECT 58.96 4.062 58.965 4.63 ;
      RECT 58.93 4.077 58.96 4.63 ;
      RECT 58.855 4.119 58.93 4.63 ;
      RECT 58.85 4.15 58.855 4.613 ;
      RECT 58.845 4.154 58.85 4.595 ;
      RECT 58.84 4.158 58.845 4.558 ;
      RECT 58.835 4.342 58.84 4.525 ;
      RECT 58.32 4.531 58.406 5.096 ;
      RECT 58.275 4.533 58.44 5.09 ;
      RECT 58.406 4.53 58.44 5.09 ;
      RECT 58.32 4.532 58.525 5.084 ;
      RECT 58.275 4.542 58.535 5.08 ;
      RECT 58.25 4.534 58.525 5.076 ;
      RECT 58.245 4.537 58.525 5.071 ;
      RECT 58.22 4.552 58.535 5.065 ;
      RECT 58.22 4.577 58.575 5.06 ;
      RECT 58.18 4.585 58.575 5.035 ;
      RECT 58.18 4.612 58.59 5.033 ;
      RECT 58.18 4.642 58.6 5.02 ;
      RECT 58.175 4.787 58.6 5.008 ;
      RECT 58.18 4.716 58.62 5.005 ;
      RECT 58.18 4.773 58.625 4.813 ;
      RECT 58.37 4.052 58.54 4.23 ;
      RECT 58.32 3.991 58.37 4.215 ;
      RECT 58.055 3.971 58.32 4.2 ;
      RECT 58.015 4.035 58.49 4.2 ;
      RECT 58.015 4.025 58.445 4.2 ;
      RECT 58.015 4.022 58.435 4.2 ;
      RECT 58.015 4.01 58.425 4.2 ;
      RECT 58.015 3.995 58.37 4.2 ;
      RECT 58.055 3.967 58.256 4.2 ;
      RECT 58.065 3.945 58.256 4.2 ;
      RECT 58.09 3.93 58.17 4.2 ;
      RECT 57.845 4.46 57.965 4.905 ;
      RECT 57.83 4.46 57.965 4.904 ;
      RECT 57.785 4.482 57.965 4.899 ;
      RECT 57.745 4.531 57.965 4.893 ;
      RECT 57.745 4.531 57.97 4.868 ;
      RECT 57.745 4.531 57.99 4.758 ;
      RECT 57.74 4.561 57.99 4.755 ;
      RECT 57.83 4.46 58 4.65 ;
      RECT 57.49 3.245 57.495 3.69 ;
      RECT 57.3 3.245 57.32 3.655 ;
      RECT 57.27 3.245 57.275 3.63 ;
      RECT 57.95 3.552 57.965 3.74 ;
      RECT 57.945 3.537 57.95 3.746 ;
      RECT 57.925 3.51 57.945 3.749 ;
      RECT 57.875 3.477 57.925 3.758 ;
      RECT 57.845 3.457 57.875 3.762 ;
      RECT 57.826 3.445 57.845 3.758 ;
      RECT 57.74 3.417 57.826 3.748 ;
      RECT 57.73 3.392 57.74 3.738 ;
      RECT 57.66 3.36 57.73 3.73 ;
      RECT 57.635 3.32 57.66 3.722 ;
      RECT 57.615 3.302 57.635 3.716 ;
      RECT 57.605 3.292 57.615 3.713 ;
      RECT 57.595 3.285 57.605 3.711 ;
      RECT 57.575 3.272 57.595 3.708 ;
      RECT 57.565 3.262 57.575 3.705 ;
      RECT 57.555 3.255 57.565 3.703 ;
      RECT 57.505 3.247 57.555 3.697 ;
      RECT 57.495 3.245 57.505 3.691 ;
      RECT 57.465 3.245 57.49 3.688 ;
      RECT 57.436 3.245 57.465 3.683 ;
      RECT 57.35 3.245 57.436 3.673 ;
      RECT 57.32 3.245 57.35 3.66 ;
      RECT 57.275 3.245 57.3 3.643 ;
      RECT 57.26 3.245 57.27 3.625 ;
      RECT 57.24 3.252 57.26 3.61 ;
      RECT 57.235 3.267 57.24 3.598 ;
      RECT 57.23 3.272 57.235 3.538 ;
      RECT 57.225 3.277 57.23 3.38 ;
      RECT 57.22 3.28 57.225 3.298 ;
      RECT 56.96 4.57 56.995 4.89 ;
      RECT 57.545 4.755 57.55 4.937 ;
      RECT 57.5 4.637 57.545 4.956 ;
      RECT 57.485 4.614 57.5 4.979 ;
      RECT 57.475 4.604 57.485 4.989 ;
      RECT 57.455 4.599 57.475 5.002 ;
      RECT 57.43 4.597 57.455 5.023 ;
      RECT 57.411 4.596 57.43 5.035 ;
      RECT 57.325 4.593 57.411 5.035 ;
      RECT 57.255 4.588 57.325 5.023 ;
      RECT 57.18 4.584 57.255 4.998 ;
      RECT 57.115 4.58 57.18 4.965 ;
      RECT 57.045 4.577 57.115 4.925 ;
      RECT 57.015 4.573 57.045 4.9 ;
      RECT 56.995 4.571 57.015 4.893 ;
      RECT 56.911 4.569 56.96 4.891 ;
      RECT 56.825 4.566 56.911 4.892 ;
      RECT 56.75 4.565 56.825 4.894 ;
      RECT 56.665 4.565 56.75 4.92 ;
      RECT 56.588 4.566 56.665 4.945 ;
      RECT 56.502 4.567 56.588 4.945 ;
      RECT 56.416 4.567 56.502 4.945 ;
      RECT 56.33 4.568 56.416 4.945 ;
      RECT 56.31 4.569 56.33 4.937 ;
      RECT 56.295 4.575 56.31 4.922 ;
      RECT 56.26 4.595 56.295 4.902 ;
      RECT 56.25 4.615 56.26 4.884 ;
      RECT 57.22 3.92 57.225 4.19 ;
      RECT 57.215 3.911 57.22 4.195 ;
      RECT 57.205 3.901 57.215 4.207 ;
      RECT 57.2 3.89 57.205 4.218 ;
      RECT 57.18 3.884 57.2 4.236 ;
      RECT 57.135 3.881 57.18 4.285 ;
      RECT 57.12 3.88 57.135 4.33 ;
      RECT 57.115 3.88 57.12 4.343 ;
      RECT 57.105 3.88 57.115 4.355 ;
      RECT 57.1 3.881 57.105 4.37 ;
      RECT 57.08 3.889 57.1 4.375 ;
      RECT 57.05 3.905 57.08 4.375 ;
      RECT 57.04 3.917 57.045 4.375 ;
      RECT 57.005 3.932 57.04 4.375 ;
      RECT 56.975 3.952 57.005 4.375 ;
      RECT 56.965 3.977 56.975 4.375 ;
      RECT 56.96 4.005 56.965 4.375 ;
      RECT 56.955 4.035 56.96 4.375 ;
      RECT 56.95 4.052 56.955 4.375 ;
      RECT 56.94 4.08 56.95 4.375 ;
      RECT 56.93 4.115 56.94 4.375 ;
      RECT 56.925 4.15 56.93 4.375 ;
      RECT 57.045 3.915 57.05 4.375 ;
      RECT 56.035 3.245 56.04 3.644 ;
      RECT 55.78 3.245 55.815 3.642 ;
      RECT 55.375 3.28 55.38 3.636 ;
      RECT 56.12 3.283 56.125 3.538 ;
      RECT 56.115 3.281 56.12 3.544 ;
      RECT 56.11 3.28 56.115 3.551 ;
      RECT 56.085 3.273 56.11 3.575 ;
      RECT 56.08 3.266 56.085 3.599 ;
      RECT 56.075 3.262 56.08 3.608 ;
      RECT 56.065 3.257 56.075 3.621 ;
      RECT 56.06 3.254 56.065 3.63 ;
      RECT 56.055 3.252 56.06 3.635 ;
      RECT 56.04 3.248 56.055 3.645 ;
      RECT 56.025 3.242 56.035 3.644 ;
      RECT 55.987 3.24 56.025 3.644 ;
      RECT 55.901 3.242 55.987 3.644 ;
      RECT 55.815 3.244 55.901 3.643 ;
      RECT 55.744 3.245 55.78 3.642 ;
      RECT 55.658 3.247 55.744 3.642 ;
      RECT 55.572 3.249 55.658 3.641 ;
      RECT 55.486 3.251 55.572 3.641 ;
      RECT 55.4 3.254 55.486 3.64 ;
      RECT 55.39 3.26 55.4 3.639 ;
      RECT 55.38 3.272 55.39 3.637 ;
      RECT 55.32 3.307 55.375 3.633 ;
      RECT 55.315 3.337 55.32 3.395 ;
      RECT 55.66 4.552 55.665 4.809 ;
      RECT 55.64 4.471 55.66 4.826 ;
      RECT 55.62 4.465 55.64 4.855 ;
      RECT 55.56 4.452 55.62 4.875 ;
      RECT 55.515 4.436 55.56 4.876 ;
      RECT 55.431 4.424 55.515 4.864 ;
      RECT 55.345 4.411 55.431 4.848 ;
      RECT 55.335 4.404 55.345 4.84 ;
      RECT 55.29 4.401 55.335 4.78 ;
      RECT 55.27 4.397 55.29 4.695 ;
      RECT 55.255 4.395 55.27 4.648 ;
      RECT 55.225 4.392 55.255 4.618 ;
      RECT 55.19 4.388 55.225 4.595 ;
      RECT 55.147 4.383 55.19 4.583 ;
      RECT 55.061 4.374 55.147 4.592 ;
      RECT 54.975 4.363 55.061 4.604 ;
      RECT 54.91 4.354 54.975 4.613 ;
      RECT 54.89 4.345 54.91 4.618 ;
      RECT 54.885 4.338 54.89 4.62 ;
      RECT 54.845 4.323 54.885 4.617 ;
      RECT 54.825 4.302 54.845 4.612 ;
      RECT 54.81 4.29 54.825 4.605 ;
      RECT 54.805 4.282 54.81 4.598 ;
      RECT 54.79 4.262 54.805 4.591 ;
      RECT 54.785 4.125 54.79 4.585 ;
      RECT 54.705 4.014 54.785 4.557 ;
      RECT 54.696 4.007 54.705 4.523 ;
      RECT 54.61 4.001 54.696 4.448 ;
      RECT 54.585 3.992 54.61 4.36 ;
      RECT 54.555 3.987 54.585 4.335 ;
      RECT 54.49 3.996 54.555 4.32 ;
      RECT 54.47 4.012 54.49 4.295 ;
      RECT 54.46 4.018 54.47 4.243 ;
      RECT 54.44 4.04 54.46 4.125 ;
      RECT 55.095 4.072 55.32 4.19 ;
      RECT 55.095 3.915 55.315 4.19 ;
      RECT 54.31 4.683 54.375 5.126 ;
      RECT 54.25 4.708 54.375 5.124 ;
      RECT 54.25 4.708 54.43 5.118 ;
      RECT 54.235 4.733 54.43 5.117 ;
      RECT 54.375 4.67 54.45 5.114 ;
      RECT 54.31 4.695 54.53 5.108 ;
      RECT 54.235 4.734 54.575 5.102 ;
      RECT 54.22 4.761 54.575 5.093 ;
      RECT 54.235 4.754 54.595 5.085 ;
      RECT 54.22 4.763 54.6 5.068 ;
      RECT 54.215 4.78 54.6 4.895 ;
      RECT 54.22 3.502 54.255 3.74 ;
      RECT 54.22 3.502 54.285 3.739 ;
      RECT 54.22 3.502 54.4 3.735 ;
      RECT 54.22 3.502 54.455 3.713 ;
      RECT 54.23 3.445 54.51 3.613 ;
      RECT 54.335 3.285 54.365 3.736 ;
      RECT 54.365 3.28 54.545 3.493 ;
      RECT 54.235 3.421 54.545 3.493 ;
      RECT 54.285 3.317 54.335 3.737 ;
      RECT 54.255 3.373 54.545 3.493 ;
      RECT 53.115 7.455 53.285 8.925 ;
      RECT 53.115 7.455 53.29 8.715 ;
      RECT 52.745 9.405 53.215 9.575 ;
      RECT 52.745 8.385 52.915 9.575 ;
      RECT 52.74 3.035 52.91 4.225 ;
      RECT 52.74 3.035 53.21 3.205 ;
      RECT 52.125 3.895 52.3 5.155 ;
      RECT 52.125 3.685 52.295 5.155 ;
      RECT 52.125 7.455 52.295 8.925 ;
      RECT 52.125 7.455 52.3 8.715 ;
      RECT 51.755 3.035 51.925 4.225 ;
      RECT 51.755 3.035 52.225 3.205 ;
      RECT 51.755 9.405 52.225 9.575 ;
      RECT 51.755 8.385 51.925 9.575 ;
      RECT 50.765 4.015 50.94 5.155 ;
      RECT 50.765 1.865 50.935 5.155 ;
      RECT 50.765 1.865 50.94 2.415 ;
      RECT 50.765 10.195 50.94 10.745 ;
      RECT 50.765 7.455 50.935 10.745 ;
      RECT 50.765 7.455 50.94 8.595 ;
      RECT 50.335 3.895 50.51 5.155 ;
      RECT 50.335 2.945 50.505 5.155 ;
      RECT 50.335 7.455 50.505 9.665 ;
      RECT 50.335 7.455 50.51 8.715 ;
      RECT 49.905 3.925 50.075 5.155 ;
      RECT 49.965 2.145 50.135 4.095 ;
      RECT 49.905 1.865 50.075 2.315 ;
      RECT 49.905 10.295 50.075 10.745 ;
      RECT 49.965 8.515 50.135 10.465 ;
      RECT 49.905 7.455 50.075 8.685 ;
      RECT 49.38 3.895 49.555 5.155 ;
      RECT 49.38 1.865 49.55 5.155 ;
      RECT 49.38 3.365 49.79 3.695 ;
      RECT 49.38 2.525 49.79 2.855 ;
      RECT 49.38 1.865 49.555 2.355 ;
      RECT 49.38 10.255 49.555 10.745 ;
      RECT 49.38 7.455 49.55 10.745 ;
      RECT 49.38 9.755 49.79 10.085 ;
      RECT 49.38 8.915 49.79 9.245 ;
      RECT 49.38 7.455 49.555 8.715 ;
      RECT 47.495 4.687 47.51 4.738 ;
      RECT 47.49 4.667 47.495 4.785 ;
      RECT 47.475 4.657 47.49 4.853 ;
      RECT 47.45 4.637 47.475 4.908 ;
      RECT 47.41 4.622 47.45 4.928 ;
      RECT 47.365 4.616 47.41 4.956 ;
      RECT 47.295 4.606 47.365 4.973 ;
      RECT 47.275 4.598 47.295 4.973 ;
      RECT 47.215 4.592 47.275 4.965 ;
      RECT 47.156 4.583 47.215 4.953 ;
      RECT 47.07 4.572 47.156 4.936 ;
      RECT 47.048 4.563 47.07 4.924 ;
      RECT 46.962 4.556 47.048 4.911 ;
      RECT 46.876 4.543 46.962 4.892 ;
      RECT 46.79 4.531 46.876 4.872 ;
      RECT 46.76 4.52 46.79 4.859 ;
      RECT 46.71 4.506 46.76 4.851 ;
      RECT 46.69 4.495 46.71 4.843 ;
      RECT 46.641 4.484 46.69 4.835 ;
      RECT 46.555 4.463 46.641 4.82 ;
      RECT 46.51 4.45 46.555 4.805 ;
      RECT 46.465 4.45 46.51 4.785 ;
      RECT 46.41 4.45 46.465 4.72 ;
      RECT 46.385 4.45 46.41 4.643 ;
      RECT 46.91 4.187 47.08 4.37 ;
      RECT 46.91 4.187 47.095 4.328 ;
      RECT 46.91 4.187 47.1 4.27 ;
      RECT 46.97 3.955 47.105 4.246 ;
      RECT 46.97 3.959 47.11 4.229 ;
      RECT 46.915 4.122 47.11 4.229 ;
      RECT 46.94 3.967 47.08 4.37 ;
      RECT 46.94 3.971 47.12 4.17 ;
      RECT 46.925 4.057 47.12 4.17 ;
      RECT 46.935 3.987 47.08 4.37 ;
      RECT 46.935 3.99 47.13 4.083 ;
      RECT 46.93 4.007 47.13 4.083 ;
      RECT 46.7 3.227 46.87 3.71 ;
      RECT 46.695 3.222 46.845 3.7 ;
      RECT 46.695 3.229 46.875 3.694 ;
      RECT 46.685 3.223 46.845 3.673 ;
      RECT 46.685 3.239 46.89 3.632 ;
      RECT 46.655 3.224 46.845 3.595 ;
      RECT 46.655 3.254 46.9 3.535 ;
      RECT 46.65 3.226 46.845 3.533 ;
      RECT 46.63 3.235 46.875 3.49 ;
      RECT 46.605 3.251 46.89 3.402 ;
      RECT 46.605 3.27 46.915 3.393 ;
      RECT 46.6 3.307 46.915 3.345 ;
      RECT 46.605 3.287 46.92 3.313 ;
      RECT 46.7 3.221 46.81 3.71 ;
      RECT 46.786 3.22 46.81 3.71 ;
      RECT 46.02 4.005 46.025 4.216 ;
      RECT 46.62 4.005 46.625 4.19 ;
      RECT 46.685 4.045 46.69 4.158 ;
      RECT 46.68 4.037 46.685 4.164 ;
      RECT 46.675 4.027 46.68 4.172 ;
      RECT 46.67 4.017 46.675 4.181 ;
      RECT 46.665 4.007 46.67 4.185 ;
      RECT 46.625 4.005 46.665 4.188 ;
      RECT 46.597 4.004 46.62 4.192 ;
      RECT 46.511 4.001 46.597 4.199 ;
      RECT 46.425 3.997 46.511 4.21 ;
      RECT 46.405 3.995 46.425 4.216 ;
      RECT 46.387 3.994 46.405 4.219 ;
      RECT 46.301 3.992 46.387 4.226 ;
      RECT 46.215 3.987 46.301 4.239 ;
      RECT 46.196 3.984 46.215 4.244 ;
      RECT 46.11 3.982 46.196 4.235 ;
      RECT 46.1 3.982 46.11 4.228 ;
      RECT 46.025 3.995 46.1 4.222 ;
      RECT 46.01 4.006 46.02 4.216 ;
      RECT 46 4.008 46.01 4.215 ;
      RECT 45.99 4.012 46 4.211 ;
      RECT 45.985 4.015 45.99 4.205 ;
      RECT 45.975 4.017 45.985 4.199 ;
      RECT 45.97 4.02 45.975 4.193 ;
      RECT 46.005 10.195 46.18 10.745 ;
      RECT 46.005 7.455 46.175 10.745 ;
      RECT 46.005 7.455 46.18 8.595 ;
      RECT 45.95 4.606 45.955 4.81 ;
      RECT 45.935 4.593 45.95 4.903 ;
      RECT 45.92 4.574 45.935 5.18 ;
      RECT 45.885 4.54 45.92 5.18 ;
      RECT 45.881 4.51 45.885 5.18 ;
      RECT 45.795 4.392 45.881 5.18 ;
      RECT 45.785 4.267 45.795 5.18 ;
      RECT 45.77 4.235 45.785 5.18 ;
      RECT 45.765 4.21 45.77 5.18 ;
      RECT 45.76 4.2 45.765 5.136 ;
      RECT 45.745 4.172 45.76 5.041 ;
      RECT 45.73 4.138 45.745 4.94 ;
      RECT 45.725 4.116 45.73 4.893 ;
      RECT 45.72 4.105 45.725 4.863 ;
      RECT 45.715 4.095 45.72 4.829 ;
      RECT 45.705 4.082 45.715 4.797 ;
      RECT 45.68 4.058 45.705 4.723 ;
      RECT 45.675 4.038 45.68 4.648 ;
      RECT 45.67 4.032 45.675 4.623 ;
      RECT 45.665 4.027 45.67 4.588 ;
      RECT 45.66 4.022 45.665 4.563 ;
      RECT 45.655 4.02 45.66 4.543 ;
      RECT 45.65 4.02 45.655 4.528 ;
      RECT 45.645 4.02 45.65 4.488 ;
      RECT 45.635 4.02 45.645 4.46 ;
      RECT 45.625 4.02 45.635 4.405 ;
      RECT 45.61 4.02 45.625 4.343 ;
      RECT 45.605 4.019 45.61 4.288 ;
      RECT 45.59 4.018 45.605 4.268 ;
      RECT 45.53 4.016 45.59 4.242 ;
      RECT 45.495 4.017 45.53 4.222 ;
      RECT 45.49 4.019 45.495 4.212 ;
      RECT 45.48 4.038 45.49 4.202 ;
      RECT 45.475 4.065 45.48 4.133 ;
      RECT 45.59 3.49 45.76 3.735 ;
      RECT 45.625 3.261 45.76 3.735 ;
      RECT 45.625 3.263 45.77 3.73 ;
      RECT 45.625 3.265 45.795 3.718 ;
      RECT 45.625 3.268 45.82 3.7 ;
      RECT 45.625 3.273 45.87 3.673 ;
      RECT 45.625 3.278 45.89 3.638 ;
      RECT 45.605 3.28 45.9 3.613 ;
      RECT 45.595 3.375 45.9 3.613 ;
      RECT 45.625 3.26 45.735 3.735 ;
      RECT 45.635 3.257 45.73 3.735 ;
      RECT 45.575 7.455 45.745 9.665 ;
      RECT 45.575 7.455 45.75 8.715 ;
      RECT 45.155 4.522 45.345 4.88 ;
      RECT 45.155 4.534 45.38 4.879 ;
      RECT 45.155 4.562 45.4 4.877 ;
      RECT 45.155 4.587 45.405 4.876 ;
      RECT 45.155 4.645 45.42 4.875 ;
      RECT 45.14 4.518 45.3 4.86 ;
      RECT 45.12 4.527 45.345 4.813 ;
      RECT 45.095 4.538 45.38 4.75 ;
      RECT 45.095 4.622 45.415 4.75 ;
      RECT 45.095 4.597 45.41 4.75 ;
      RECT 45.155 4.513 45.3 4.88 ;
      RECT 45.241 4.512 45.3 4.88 ;
      RECT 45.241 4.511 45.285 4.88 ;
      RECT 44.62 10.255 44.795 10.745 ;
      RECT 44.62 7.455 44.79 10.745 ;
      RECT 44.62 9.755 45.03 10.085 ;
      RECT 44.62 8.915 45.03 9.245 ;
      RECT 44.62 7.455 44.795 8.715 ;
      RECT 44.94 4.027 44.945 4.405 ;
      RECT 44.935 3.995 44.94 4.405 ;
      RECT 44.93 3.967 44.935 4.405 ;
      RECT 44.925 3.947 44.93 4.405 ;
      RECT 44.87 3.93 44.925 4.405 ;
      RECT 44.83 3.915 44.87 4.405 ;
      RECT 44.775 3.902 44.83 4.405 ;
      RECT 44.74 3.893 44.775 4.405 ;
      RECT 44.736 3.891 44.74 4.404 ;
      RECT 44.65 3.887 44.736 4.387 ;
      RECT 44.565 3.879 44.65 4.35 ;
      RECT 44.555 3.875 44.565 4.323 ;
      RECT 44.545 3.875 44.555 4.305 ;
      RECT 44.535 3.877 44.545 4.288 ;
      RECT 44.53 3.882 44.535 4.274 ;
      RECT 44.525 3.886 44.53 4.261 ;
      RECT 44.515 3.891 44.525 4.245 ;
      RECT 44.5 3.905 44.515 4.22 ;
      RECT 44.495 3.911 44.5 4.2 ;
      RECT 44.49 3.913 44.495 4.193 ;
      RECT 44.485 3.917 44.49 4.068 ;
      RECT 44.665 4.717 44.91 5.18 ;
      RECT 44.585 4.69 44.905 5.176 ;
      RECT 44.515 4.725 44.91 5.169 ;
      RECT 44.305 4.98 44.91 5.165 ;
      RECT 44.485 4.748 44.91 5.165 ;
      RECT 44.325 4.94 44.91 5.165 ;
      RECT 44.475 4.76 44.91 5.165 ;
      RECT 44.36 4.877 44.91 5.165 ;
      RECT 44.415 4.802 44.91 5.165 ;
      RECT 44.665 4.667 44.905 5.18 ;
      RECT 44.695 4.66 44.905 5.18 ;
      RECT 44.685 4.662 44.905 5.18 ;
      RECT 44.695 4.657 44.825 5.18 ;
      RECT 44.25 3.22 44.336 3.659 ;
      RECT 44.245 3.22 44.336 3.657 ;
      RECT 44.245 3.22 44.405 3.656 ;
      RECT 44.245 3.22 44.435 3.653 ;
      RECT 44.23 3.227 44.435 3.644 ;
      RECT 44.23 3.227 44.44 3.64 ;
      RECT 44.225 3.237 44.44 3.633 ;
      RECT 44.22 3.242 44.44 3.608 ;
      RECT 44.22 3.242 44.455 3.59 ;
      RECT 44.245 3.22 44.475 3.505 ;
      RECT 44.215 3.247 44.475 3.503 ;
      RECT 44.225 3.24 44.48 3.441 ;
      RECT 44.215 3.362 44.485 3.424 ;
      RECT 44.2 3.257 44.48 3.375 ;
      RECT 44.195 3.267 44.48 3.275 ;
      RECT 44.275 4.038 44.28 4.115 ;
      RECT 44.265 4.032 44.275 4.305 ;
      RECT 44.255 4.024 44.265 4.326 ;
      RECT 44.245 4.015 44.255 4.348 ;
      RECT 44.24 4.01 44.245 4.365 ;
      RECT 44.2 4.01 44.24 4.405 ;
      RECT 44.18 4.01 44.2 4.46 ;
      RECT 44.175 4.01 44.18 4.488 ;
      RECT 44.165 4.01 44.175 4.503 ;
      RECT 44.13 4.01 44.165 4.545 ;
      RECT 44.125 4.01 44.13 4.588 ;
      RECT 44.115 4.01 44.125 4.603 ;
      RECT 44.1 4.01 44.115 4.623 ;
      RECT 44.085 4.01 44.1 4.65 ;
      RECT 44.08 4.011 44.085 4.668 ;
      RECT 44.06 4.012 44.08 4.675 ;
      RECT 44.005 4.013 44.06 4.695 ;
      RECT 43.995 4.014 44.005 4.709 ;
      RECT 43.99 4.017 43.995 4.708 ;
      RECT 43.95 4.09 43.99 4.706 ;
      RECT 43.935 4.17 43.95 4.704 ;
      RECT 43.91 4.225 43.935 4.702 ;
      RECT 43.895 4.29 43.91 4.701 ;
      RECT 43.85 4.322 43.895 4.698 ;
      RECT 43.765 4.345 43.85 4.693 ;
      RECT 43.74 4.365 43.765 4.688 ;
      RECT 43.67 4.37 43.74 4.684 ;
      RECT 43.65 4.372 43.67 4.681 ;
      RECT 43.565 4.383 43.65 4.675 ;
      RECT 43.56 4.394 43.565 4.67 ;
      RECT 43.55 4.396 43.56 4.67 ;
      RECT 43.515 4.4 43.55 4.668 ;
      RECT 43.465 4.41 43.515 4.655 ;
      RECT 43.445 4.418 43.465 4.64 ;
      RECT 43.365 4.43 43.445 4.623 ;
      RECT 43.53 3.98 43.7 4.19 ;
      RECT 43.646 3.976 43.7 4.19 ;
      RECT 43.451 3.98 43.7 4.181 ;
      RECT 43.451 3.98 43.705 4.17 ;
      RECT 43.365 3.98 43.705 4.161 ;
      RECT 43.365 3.988 43.715 4.105 ;
      RECT 43.365 4 43.72 4.018 ;
      RECT 43.365 4.007 43.725 4.01 ;
      RECT 43.56 3.978 43.7 4.19 ;
      RECT 43.315 4.923 43.56 5.255 ;
      RECT 43.31 4.915 43.315 5.252 ;
      RECT 43.28 4.935 43.56 5.233 ;
      RECT 43.26 4.967 43.56 5.206 ;
      RECT 43.31 4.92 43.487 5.252 ;
      RECT 43.31 4.917 43.401 5.252 ;
      RECT 43.25 3.265 43.42 3.685 ;
      RECT 43.245 3.265 43.42 3.683 ;
      RECT 43.245 3.265 43.445 3.673 ;
      RECT 43.245 3.265 43.465 3.648 ;
      RECT 43.24 3.265 43.465 3.643 ;
      RECT 43.24 3.265 43.475 3.633 ;
      RECT 43.24 3.265 43.48 3.628 ;
      RECT 43.24 3.27 43.485 3.623 ;
      RECT 43.24 3.302 43.5 3.613 ;
      RECT 43.24 3.372 43.525 3.596 ;
      RECT 43.22 3.372 43.525 3.588 ;
      RECT 43.22 3.432 43.535 3.565 ;
      RECT 43.22 3.472 43.545 3.51 ;
      RECT 43.205 3.265 43.48 3.49 ;
      RECT 43.195 3.28 43.485 3.388 ;
      RECT 42.785 4.67 42.955 5.195 ;
      RECT 42.78 4.67 42.955 5.188 ;
      RECT 42.77 4.67 42.96 5.153 ;
      RECT 42.765 4.68 42.96 5.125 ;
      RECT 42.76 4.7 42.96 5.108 ;
      RECT 42.77 4.675 42.965 5.098 ;
      RECT 42.755 4.72 42.965 5.09 ;
      RECT 42.75 4.74 42.965 5.075 ;
      RECT 42.745 4.77 42.965 5.065 ;
      RECT 42.735 4.815 42.965 5.04 ;
      RECT 42.765 4.685 42.97 5.023 ;
      RECT 42.73 4.867 42.97 5.018 ;
      RECT 42.765 4.695 42.975 4.988 ;
      RECT 42.725 4.9 42.975 4.985 ;
      RECT 42.72 4.925 42.975 4.965 ;
      RECT 42.76 4.712 42.985 4.905 ;
      RECT 42.755 4.734 42.995 4.798 ;
      RECT 42.705 3.981 42.72 4.25 ;
      RECT 42.66 3.965 42.705 4.295 ;
      RECT 42.655 3.953 42.66 4.345 ;
      RECT 42.645 3.949 42.655 4.378 ;
      RECT 42.64 3.946 42.645 4.406 ;
      RECT 42.625 3.948 42.64 4.448 ;
      RECT 42.62 3.952 42.625 4.488 ;
      RECT 42.6 3.957 42.62 4.54 ;
      RECT 42.596 3.962 42.6 4.597 ;
      RECT 42.51 3.981 42.596 4.634 ;
      RECT 42.5 4.002 42.51 4.67 ;
      RECT 42.495 4.01 42.5 4.671 ;
      RECT 42.49 4.052 42.495 4.672 ;
      RECT 42.475 4.14 42.49 4.673 ;
      RECT 42.465 4.29 42.475 4.675 ;
      RECT 42.46 4.335 42.465 4.677 ;
      RECT 42.425 4.377 42.46 4.68 ;
      RECT 42.42 4.395 42.425 4.683 ;
      RECT 42.343 4.401 42.42 4.689 ;
      RECT 42.257 4.415 42.343 4.702 ;
      RECT 42.171 4.429 42.257 4.716 ;
      RECT 42.085 4.443 42.171 4.729 ;
      RECT 42.025 4.455 42.085 4.741 ;
      RECT 42 4.462 42.025 4.748 ;
      RECT 41.986 4.465 42 4.753 ;
      RECT 41.9 4.473 41.986 4.769 ;
      RECT 41.895 4.48 41.9 4.784 ;
      RECT 41.871 4.48 41.895 4.791 ;
      RECT 41.785 4.483 41.871 4.819 ;
      RECT 41.7 4.487 41.785 4.863 ;
      RECT 41.635 4.491 41.7 4.9 ;
      RECT 41.61 4.494 41.635 4.916 ;
      RECT 41.535 4.507 41.61 4.92 ;
      RECT 41.51 4.525 41.535 4.924 ;
      RECT 41.5 4.532 41.51 4.926 ;
      RECT 41.485 4.535 41.5 4.927 ;
      RECT 41.425 4.547 41.485 4.931 ;
      RECT 41.415 4.561 41.425 4.935 ;
      RECT 41.36 4.571 41.415 4.923 ;
      RECT 41.335 4.592 41.36 4.906 ;
      RECT 41.315 4.612 41.335 4.897 ;
      RECT 41.31 4.625 41.315 4.892 ;
      RECT 41.295 4.637 41.31 4.888 ;
      RECT 42.53 3.292 42.535 3.315 ;
      RECT 42.525 3.283 42.53 3.355 ;
      RECT 42.52 3.281 42.525 3.398 ;
      RECT 42.515 3.272 42.52 3.433 ;
      RECT 42.51 3.262 42.515 3.505 ;
      RECT 42.505 3.252 42.51 3.57 ;
      RECT 42.5 3.249 42.505 3.61 ;
      RECT 42.475 3.243 42.5 3.7 ;
      RECT 42.44 3.231 42.475 3.725 ;
      RECT 42.43 3.222 42.44 3.725 ;
      RECT 42.295 3.22 42.305 3.708 ;
      RECT 42.285 3.22 42.295 3.675 ;
      RECT 42.28 3.22 42.285 3.65 ;
      RECT 42.275 3.22 42.28 3.638 ;
      RECT 42.27 3.22 42.275 3.62 ;
      RECT 42.26 3.22 42.27 3.585 ;
      RECT 42.255 3.222 42.26 3.563 ;
      RECT 42.25 3.228 42.255 3.548 ;
      RECT 42.245 3.234 42.25 3.533 ;
      RECT 42.23 3.246 42.245 3.506 ;
      RECT 42.225 3.257 42.23 3.474 ;
      RECT 42.22 3.267 42.225 3.458 ;
      RECT 42.21 3.275 42.22 3.427 ;
      RECT 42.205 3.285 42.21 3.401 ;
      RECT 42.2 3.342 42.205 3.384 ;
      RECT 42.305 3.22 42.43 3.725 ;
      RECT 42.02 3.907 42.28 4.205 ;
      RECT 42.015 3.914 42.28 4.203 ;
      RECT 42.02 3.909 42.295 4.198 ;
      RECT 42.01 3.922 42.295 4.195 ;
      RECT 42.01 3.927 42.3 4.188 ;
      RECT 42.005 3.935 42.3 4.185 ;
      RECT 42.005 3.952 42.305 3.983 ;
      RECT 42.02 3.904 42.251 4.205 ;
      RECT 42.075 3.903 42.251 4.205 ;
      RECT 42.075 3.9 42.165 4.205 ;
      RECT 42.075 3.897 42.161 4.205 ;
      RECT 41.765 4.17 41.77 4.183 ;
      RECT 41.76 4.137 41.765 4.188 ;
      RECT 41.755 4.092 41.76 4.195 ;
      RECT 41.75 4.047 41.755 4.203 ;
      RECT 41.745 4.015 41.75 4.211 ;
      RECT 41.74 3.975 41.745 4.212 ;
      RECT 41.725 3.955 41.74 4.214 ;
      RECT 41.65 3.937 41.725 4.226 ;
      RECT 41.64 3.93 41.65 4.237 ;
      RECT 41.635 3.93 41.64 4.239 ;
      RECT 41.605 3.936 41.635 4.243 ;
      RECT 41.565 3.949 41.605 4.243 ;
      RECT 41.54 3.96 41.565 4.229 ;
      RECT 41.525 3.966 41.54 4.212 ;
      RECT 41.515 3.968 41.525 4.203 ;
      RECT 41.51 3.969 41.515 4.198 ;
      RECT 41.505 3.97 41.51 4.193 ;
      RECT 41.5 3.971 41.505 4.19 ;
      RECT 41.475 3.976 41.5 4.18 ;
      RECT 41.465 3.992 41.475 4.167 ;
      RECT 41.46 4.012 41.465 4.162 ;
      RECT 41.47 3.405 41.475 3.601 ;
      RECT 41.455 3.369 41.47 3.603 ;
      RECT 41.445 3.351 41.455 3.608 ;
      RECT 41.435 3.337 41.445 3.612 ;
      RECT 41.39 3.321 41.435 3.622 ;
      RECT 41.385 3.311 41.39 3.631 ;
      RECT 41.34 3.3 41.385 3.637 ;
      RECT 41.335 3.288 41.34 3.644 ;
      RECT 41.32 3.283 41.335 3.648 ;
      RECT 41.305 3.275 41.32 3.653 ;
      RECT 41.295 3.268 41.305 3.658 ;
      RECT 41.285 3.265 41.295 3.663 ;
      RECT 41.275 3.265 41.285 3.664 ;
      RECT 41.27 3.262 41.275 3.663 ;
      RECT 41.235 3.257 41.26 3.662 ;
      RECT 41.211 3.253 41.235 3.661 ;
      RECT 41.125 3.244 41.211 3.658 ;
      RECT 41.11 3.236 41.125 3.655 ;
      RECT 41.088 3.235 41.11 3.654 ;
      RECT 41.002 3.235 41.088 3.652 ;
      RECT 40.916 3.235 41.002 3.65 ;
      RECT 40.83 3.235 40.916 3.647 ;
      RECT 40.82 3.235 40.83 3.638 ;
      RECT 40.79 3.235 40.82 3.598 ;
      RECT 40.78 3.245 40.79 3.553 ;
      RECT 40.775 3.285 40.78 3.538 ;
      RECT 40.77 3.3 40.775 3.525 ;
      RECT 40.74 3.38 40.77 3.487 ;
      RECT 41.26 3.26 41.27 3.663 ;
      RECT 41.085 4.025 41.1 4.63 ;
      RECT 41.09 4.02 41.1 4.63 ;
      RECT 41.255 4.02 41.26 4.203 ;
      RECT 41.245 4.02 41.255 4.233 ;
      RECT 41.23 4.02 41.245 4.293 ;
      RECT 41.225 4.02 41.23 4.338 ;
      RECT 41.22 4.02 41.225 4.368 ;
      RECT 41.215 4.02 41.22 4.388 ;
      RECT 41.205 4.02 41.215 4.423 ;
      RECT 41.19 4.02 41.205 4.455 ;
      RECT 41.145 4.02 41.19 4.483 ;
      RECT 41.14 4.02 41.145 4.513 ;
      RECT 41.135 4.02 41.14 4.525 ;
      RECT 41.13 4.02 41.135 4.533 ;
      RECT 41.12 4.02 41.13 4.548 ;
      RECT 41.115 4.02 41.12 4.57 ;
      RECT 41.105 4.02 41.115 4.593 ;
      RECT 41.1 4.02 41.105 4.613 ;
      RECT 41.065 4.035 41.085 4.63 ;
      RECT 41.04 4.052 41.065 4.63 ;
      RECT 41.035 4.062 41.04 4.63 ;
      RECT 41.005 4.077 41.035 4.63 ;
      RECT 40.93 4.119 41.005 4.63 ;
      RECT 40.925 4.15 40.93 4.613 ;
      RECT 40.92 4.154 40.925 4.595 ;
      RECT 40.915 4.158 40.92 4.558 ;
      RECT 40.91 4.342 40.915 4.525 ;
      RECT 40.395 4.531 40.481 5.096 ;
      RECT 40.35 4.533 40.515 5.09 ;
      RECT 40.481 4.53 40.515 5.09 ;
      RECT 40.395 4.532 40.6 5.084 ;
      RECT 40.35 4.542 40.61 5.08 ;
      RECT 40.325 4.534 40.6 5.076 ;
      RECT 40.32 4.537 40.6 5.071 ;
      RECT 40.295 4.552 40.61 5.065 ;
      RECT 40.295 4.577 40.65 5.06 ;
      RECT 40.255 4.585 40.65 5.035 ;
      RECT 40.255 4.612 40.665 5.033 ;
      RECT 40.255 4.642 40.675 5.02 ;
      RECT 40.25 4.787 40.675 5.008 ;
      RECT 40.255 4.716 40.695 5.005 ;
      RECT 40.255 4.773 40.7 4.813 ;
      RECT 40.445 4.052 40.615 4.23 ;
      RECT 40.395 3.991 40.445 4.215 ;
      RECT 40.13 3.971 40.395 4.2 ;
      RECT 40.09 4.035 40.565 4.2 ;
      RECT 40.09 4.025 40.52 4.2 ;
      RECT 40.09 4.022 40.51 4.2 ;
      RECT 40.09 4.01 40.5 4.2 ;
      RECT 40.09 3.995 40.445 4.2 ;
      RECT 40.13 3.967 40.331 4.2 ;
      RECT 40.14 3.945 40.331 4.2 ;
      RECT 40.165 3.93 40.245 4.2 ;
      RECT 39.92 4.46 40.04 4.905 ;
      RECT 39.905 4.46 40.04 4.904 ;
      RECT 39.86 4.482 40.04 4.899 ;
      RECT 39.82 4.531 40.04 4.893 ;
      RECT 39.82 4.531 40.045 4.868 ;
      RECT 39.82 4.531 40.065 4.758 ;
      RECT 39.815 4.561 40.065 4.755 ;
      RECT 39.905 4.46 40.075 4.65 ;
      RECT 39.565 3.245 39.57 3.69 ;
      RECT 39.375 3.245 39.395 3.655 ;
      RECT 39.345 3.245 39.35 3.63 ;
      RECT 40.025 3.552 40.04 3.74 ;
      RECT 40.02 3.537 40.025 3.746 ;
      RECT 40 3.51 40.02 3.749 ;
      RECT 39.95 3.477 40 3.758 ;
      RECT 39.92 3.457 39.95 3.762 ;
      RECT 39.901 3.445 39.92 3.758 ;
      RECT 39.815 3.417 39.901 3.748 ;
      RECT 39.805 3.392 39.815 3.738 ;
      RECT 39.735 3.36 39.805 3.73 ;
      RECT 39.71 3.32 39.735 3.722 ;
      RECT 39.69 3.302 39.71 3.716 ;
      RECT 39.68 3.292 39.69 3.713 ;
      RECT 39.67 3.285 39.68 3.711 ;
      RECT 39.65 3.272 39.67 3.708 ;
      RECT 39.64 3.262 39.65 3.705 ;
      RECT 39.63 3.255 39.64 3.703 ;
      RECT 39.58 3.247 39.63 3.697 ;
      RECT 39.57 3.245 39.58 3.691 ;
      RECT 39.54 3.245 39.565 3.688 ;
      RECT 39.511 3.245 39.54 3.683 ;
      RECT 39.425 3.245 39.511 3.673 ;
      RECT 39.395 3.245 39.425 3.66 ;
      RECT 39.35 3.245 39.375 3.643 ;
      RECT 39.335 3.245 39.345 3.625 ;
      RECT 39.315 3.252 39.335 3.61 ;
      RECT 39.31 3.267 39.315 3.598 ;
      RECT 39.305 3.272 39.31 3.538 ;
      RECT 39.3 3.277 39.305 3.38 ;
      RECT 39.295 3.28 39.3 3.298 ;
      RECT 39.035 4.57 39.07 4.89 ;
      RECT 39.62 4.755 39.625 4.937 ;
      RECT 39.575 4.637 39.62 4.956 ;
      RECT 39.56 4.614 39.575 4.979 ;
      RECT 39.55 4.604 39.56 4.989 ;
      RECT 39.53 4.599 39.55 5.002 ;
      RECT 39.505 4.597 39.53 5.023 ;
      RECT 39.486 4.596 39.505 5.035 ;
      RECT 39.4 4.593 39.486 5.035 ;
      RECT 39.33 4.588 39.4 5.023 ;
      RECT 39.255 4.584 39.33 4.998 ;
      RECT 39.19 4.58 39.255 4.965 ;
      RECT 39.12 4.577 39.19 4.925 ;
      RECT 39.09 4.573 39.12 4.9 ;
      RECT 39.07 4.571 39.09 4.893 ;
      RECT 38.986 4.569 39.035 4.891 ;
      RECT 38.9 4.566 38.986 4.892 ;
      RECT 38.825 4.565 38.9 4.894 ;
      RECT 38.74 4.565 38.825 4.92 ;
      RECT 38.663 4.566 38.74 4.945 ;
      RECT 38.577 4.567 38.663 4.945 ;
      RECT 38.491 4.567 38.577 4.945 ;
      RECT 38.405 4.568 38.491 4.945 ;
      RECT 38.385 4.569 38.405 4.937 ;
      RECT 38.37 4.575 38.385 4.922 ;
      RECT 38.335 4.595 38.37 4.902 ;
      RECT 38.325 4.615 38.335 4.884 ;
      RECT 39.295 3.92 39.3 4.19 ;
      RECT 39.29 3.911 39.295 4.195 ;
      RECT 39.28 3.901 39.29 4.207 ;
      RECT 39.275 3.89 39.28 4.218 ;
      RECT 39.255 3.884 39.275 4.236 ;
      RECT 39.21 3.881 39.255 4.285 ;
      RECT 39.195 3.88 39.21 4.33 ;
      RECT 39.19 3.88 39.195 4.343 ;
      RECT 39.18 3.88 39.19 4.355 ;
      RECT 39.175 3.881 39.18 4.37 ;
      RECT 39.155 3.889 39.175 4.375 ;
      RECT 39.125 3.905 39.155 4.375 ;
      RECT 39.115 3.917 39.12 4.375 ;
      RECT 39.08 3.932 39.115 4.375 ;
      RECT 39.05 3.952 39.08 4.375 ;
      RECT 39.04 3.977 39.05 4.375 ;
      RECT 39.035 4.005 39.04 4.375 ;
      RECT 39.03 4.035 39.035 4.375 ;
      RECT 39.025 4.052 39.03 4.375 ;
      RECT 39.015 4.08 39.025 4.375 ;
      RECT 39.005 4.115 39.015 4.375 ;
      RECT 39 4.15 39.005 4.375 ;
      RECT 39.12 3.915 39.125 4.375 ;
      RECT 38.11 3.245 38.115 3.644 ;
      RECT 37.855 3.245 37.89 3.642 ;
      RECT 37.45 3.28 37.455 3.636 ;
      RECT 38.195 3.283 38.2 3.538 ;
      RECT 38.19 3.281 38.195 3.544 ;
      RECT 38.185 3.28 38.19 3.551 ;
      RECT 38.16 3.273 38.185 3.575 ;
      RECT 38.155 3.266 38.16 3.599 ;
      RECT 38.15 3.262 38.155 3.608 ;
      RECT 38.14 3.257 38.15 3.621 ;
      RECT 38.135 3.254 38.14 3.63 ;
      RECT 38.13 3.252 38.135 3.635 ;
      RECT 38.115 3.248 38.13 3.645 ;
      RECT 38.1 3.242 38.11 3.644 ;
      RECT 38.062 3.24 38.1 3.644 ;
      RECT 37.976 3.242 38.062 3.644 ;
      RECT 37.89 3.244 37.976 3.643 ;
      RECT 37.819 3.245 37.855 3.642 ;
      RECT 37.733 3.247 37.819 3.642 ;
      RECT 37.647 3.249 37.733 3.641 ;
      RECT 37.561 3.251 37.647 3.641 ;
      RECT 37.475 3.254 37.561 3.64 ;
      RECT 37.465 3.26 37.475 3.639 ;
      RECT 37.455 3.272 37.465 3.637 ;
      RECT 37.395 3.307 37.45 3.633 ;
      RECT 37.39 3.337 37.395 3.395 ;
      RECT 37.735 4.552 37.74 4.809 ;
      RECT 37.715 4.471 37.735 4.826 ;
      RECT 37.695 4.465 37.715 4.855 ;
      RECT 37.635 4.452 37.695 4.875 ;
      RECT 37.59 4.436 37.635 4.876 ;
      RECT 37.506 4.424 37.59 4.864 ;
      RECT 37.42 4.411 37.506 4.848 ;
      RECT 37.41 4.404 37.42 4.84 ;
      RECT 37.365 4.401 37.41 4.78 ;
      RECT 37.345 4.397 37.365 4.695 ;
      RECT 37.33 4.395 37.345 4.648 ;
      RECT 37.3 4.392 37.33 4.618 ;
      RECT 37.265 4.388 37.3 4.595 ;
      RECT 37.222 4.383 37.265 4.583 ;
      RECT 37.136 4.374 37.222 4.592 ;
      RECT 37.05 4.363 37.136 4.604 ;
      RECT 36.985 4.354 37.05 4.613 ;
      RECT 36.965 4.345 36.985 4.618 ;
      RECT 36.96 4.338 36.965 4.62 ;
      RECT 36.92 4.323 36.96 4.617 ;
      RECT 36.9 4.302 36.92 4.612 ;
      RECT 36.885 4.29 36.9 4.605 ;
      RECT 36.88 4.282 36.885 4.598 ;
      RECT 36.865 4.262 36.88 4.591 ;
      RECT 36.86 4.125 36.865 4.585 ;
      RECT 36.78 4.014 36.86 4.557 ;
      RECT 36.771 4.007 36.78 4.523 ;
      RECT 36.685 4.001 36.771 4.448 ;
      RECT 36.66 3.992 36.685 4.36 ;
      RECT 36.63 3.987 36.66 4.335 ;
      RECT 36.565 3.996 36.63 4.32 ;
      RECT 36.545 4.012 36.565 4.295 ;
      RECT 36.535 4.018 36.545 4.243 ;
      RECT 36.515 4.04 36.535 4.125 ;
      RECT 37.17 4.072 37.395 4.19 ;
      RECT 37.17 3.915 37.39 4.19 ;
      RECT 36.385 4.683 36.45 5.126 ;
      RECT 36.325 4.708 36.45 5.124 ;
      RECT 36.325 4.708 36.505 5.118 ;
      RECT 36.31 4.733 36.505 5.117 ;
      RECT 36.45 4.67 36.525 5.114 ;
      RECT 36.385 4.695 36.605 5.108 ;
      RECT 36.31 4.734 36.65 5.102 ;
      RECT 36.295 4.761 36.65 5.093 ;
      RECT 36.31 4.754 36.67 5.085 ;
      RECT 36.295 4.763 36.675 5.068 ;
      RECT 36.29 4.78 36.675 4.895 ;
      RECT 36.295 3.502 36.33 3.74 ;
      RECT 36.295 3.502 36.36 3.739 ;
      RECT 36.295 3.502 36.475 3.735 ;
      RECT 36.295 3.502 36.53 3.713 ;
      RECT 36.305 3.445 36.585 3.613 ;
      RECT 36.41 3.285 36.44 3.736 ;
      RECT 36.44 3.28 36.62 3.493 ;
      RECT 36.31 3.421 36.62 3.493 ;
      RECT 36.36 3.317 36.41 3.737 ;
      RECT 36.33 3.373 36.62 3.493 ;
      RECT 35.19 7.455 35.36 8.925 ;
      RECT 35.19 7.455 35.365 8.715 ;
      RECT 34.82 9.405 35.29 9.575 ;
      RECT 34.82 8.385 34.99 9.575 ;
      RECT 34.815 3.035 34.985 4.225 ;
      RECT 34.815 3.035 35.285 3.205 ;
      RECT 34.2 3.895 34.375 5.155 ;
      RECT 34.2 3.685 34.37 5.155 ;
      RECT 34.2 7.455 34.37 8.925 ;
      RECT 34.2 7.455 34.375 8.715 ;
      RECT 33.83 3.035 34 4.225 ;
      RECT 33.83 3.035 34.3 3.205 ;
      RECT 33.83 9.405 34.3 9.575 ;
      RECT 33.83 8.385 34 9.575 ;
      RECT 32.84 4.015 33.015 5.155 ;
      RECT 32.84 1.865 33.01 5.155 ;
      RECT 32.84 1.865 33.015 2.415 ;
      RECT 32.84 10.195 33.015 10.745 ;
      RECT 32.84 7.455 33.01 10.745 ;
      RECT 32.84 7.455 33.015 8.595 ;
      RECT 32.41 3.895 32.585 5.155 ;
      RECT 32.41 2.945 32.58 5.155 ;
      RECT 32.41 7.455 32.58 9.665 ;
      RECT 32.41 7.455 32.585 8.715 ;
      RECT 31.98 3.925 32.15 5.155 ;
      RECT 32.04 2.145 32.21 4.095 ;
      RECT 31.98 1.865 32.15 2.315 ;
      RECT 31.98 10.295 32.15 10.745 ;
      RECT 32.04 8.515 32.21 10.465 ;
      RECT 31.98 7.455 32.15 8.685 ;
      RECT 31.455 3.895 31.63 5.155 ;
      RECT 31.455 1.865 31.625 5.155 ;
      RECT 31.455 3.365 31.865 3.695 ;
      RECT 31.455 2.525 31.865 2.855 ;
      RECT 31.455 1.865 31.63 2.355 ;
      RECT 31.455 10.255 31.63 10.745 ;
      RECT 31.455 7.455 31.625 10.745 ;
      RECT 31.455 9.755 31.865 10.085 ;
      RECT 31.455 8.915 31.865 9.245 ;
      RECT 31.455 7.455 31.63 8.715 ;
      RECT 29.57 4.687 29.585 4.738 ;
      RECT 29.565 4.667 29.57 4.785 ;
      RECT 29.55 4.657 29.565 4.853 ;
      RECT 29.525 4.637 29.55 4.908 ;
      RECT 29.485 4.622 29.525 4.928 ;
      RECT 29.44 4.616 29.485 4.956 ;
      RECT 29.37 4.606 29.44 4.973 ;
      RECT 29.35 4.598 29.37 4.973 ;
      RECT 29.29 4.592 29.35 4.965 ;
      RECT 29.231 4.583 29.29 4.953 ;
      RECT 29.145 4.572 29.231 4.936 ;
      RECT 29.123 4.563 29.145 4.924 ;
      RECT 29.037 4.556 29.123 4.911 ;
      RECT 28.951 4.543 29.037 4.892 ;
      RECT 28.865 4.531 28.951 4.872 ;
      RECT 28.835 4.52 28.865 4.859 ;
      RECT 28.785 4.506 28.835 4.851 ;
      RECT 28.765 4.495 28.785 4.843 ;
      RECT 28.716 4.484 28.765 4.835 ;
      RECT 28.63 4.463 28.716 4.82 ;
      RECT 28.585 4.45 28.63 4.805 ;
      RECT 28.54 4.45 28.585 4.785 ;
      RECT 28.485 4.45 28.54 4.72 ;
      RECT 28.46 4.45 28.485 4.643 ;
      RECT 28.985 4.187 29.155 4.37 ;
      RECT 28.985 4.187 29.17 4.328 ;
      RECT 28.985 4.187 29.175 4.27 ;
      RECT 29.045 3.955 29.18 4.246 ;
      RECT 29.045 3.959 29.185 4.229 ;
      RECT 28.99 4.122 29.185 4.229 ;
      RECT 29.015 3.967 29.155 4.37 ;
      RECT 29.015 3.971 29.195 4.17 ;
      RECT 29 4.057 29.195 4.17 ;
      RECT 29.01 3.987 29.155 4.37 ;
      RECT 29.01 3.99 29.205 4.083 ;
      RECT 29.005 4.007 29.205 4.083 ;
      RECT 28.775 3.227 28.945 3.71 ;
      RECT 28.77 3.222 28.92 3.7 ;
      RECT 28.77 3.229 28.95 3.694 ;
      RECT 28.76 3.223 28.92 3.673 ;
      RECT 28.76 3.239 28.965 3.632 ;
      RECT 28.73 3.224 28.92 3.595 ;
      RECT 28.73 3.254 28.975 3.535 ;
      RECT 28.725 3.226 28.92 3.533 ;
      RECT 28.705 3.235 28.95 3.49 ;
      RECT 28.68 3.251 28.965 3.402 ;
      RECT 28.68 3.27 28.99 3.393 ;
      RECT 28.675 3.307 28.99 3.345 ;
      RECT 28.68 3.287 28.995 3.313 ;
      RECT 28.775 3.221 28.885 3.71 ;
      RECT 28.861 3.22 28.885 3.71 ;
      RECT 28.095 4.005 28.1 4.216 ;
      RECT 28.695 4.005 28.7 4.19 ;
      RECT 28.76 4.045 28.765 4.158 ;
      RECT 28.755 4.037 28.76 4.164 ;
      RECT 28.75 4.027 28.755 4.172 ;
      RECT 28.745 4.017 28.75 4.181 ;
      RECT 28.74 4.007 28.745 4.185 ;
      RECT 28.7 4.005 28.74 4.188 ;
      RECT 28.672 4.004 28.695 4.192 ;
      RECT 28.586 4.001 28.672 4.199 ;
      RECT 28.5 3.997 28.586 4.21 ;
      RECT 28.48 3.995 28.5 4.216 ;
      RECT 28.462 3.994 28.48 4.219 ;
      RECT 28.376 3.992 28.462 4.226 ;
      RECT 28.29 3.987 28.376 4.239 ;
      RECT 28.271 3.984 28.29 4.244 ;
      RECT 28.185 3.982 28.271 4.235 ;
      RECT 28.175 3.982 28.185 4.228 ;
      RECT 28.1 3.995 28.175 4.222 ;
      RECT 28.085 4.006 28.095 4.216 ;
      RECT 28.075 4.008 28.085 4.215 ;
      RECT 28.065 4.012 28.075 4.211 ;
      RECT 28.06 4.015 28.065 4.205 ;
      RECT 28.05 4.017 28.06 4.199 ;
      RECT 28.045 4.02 28.05 4.193 ;
      RECT 28.08 10.195 28.255 10.745 ;
      RECT 28.08 7.455 28.25 10.745 ;
      RECT 28.08 7.455 28.255 8.595 ;
      RECT 28.025 4.606 28.03 4.81 ;
      RECT 28.01 4.593 28.025 4.903 ;
      RECT 27.995 4.574 28.01 5.18 ;
      RECT 27.96 4.54 27.995 5.18 ;
      RECT 27.956 4.51 27.96 5.18 ;
      RECT 27.87 4.392 27.956 5.18 ;
      RECT 27.86 4.267 27.87 5.18 ;
      RECT 27.845 4.235 27.86 5.18 ;
      RECT 27.84 4.21 27.845 5.18 ;
      RECT 27.835 4.2 27.84 5.136 ;
      RECT 27.82 4.172 27.835 5.041 ;
      RECT 27.805 4.138 27.82 4.94 ;
      RECT 27.8 4.116 27.805 4.893 ;
      RECT 27.795 4.105 27.8 4.863 ;
      RECT 27.79 4.095 27.795 4.829 ;
      RECT 27.78 4.082 27.79 4.797 ;
      RECT 27.755 4.058 27.78 4.723 ;
      RECT 27.75 4.038 27.755 4.648 ;
      RECT 27.745 4.032 27.75 4.623 ;
      RECT 27.74 4.027 27.745 4.588 ;
      RECT 27.735 4.022 27.74 4.563 ;
      RECT 27.73 4.02 27.735 4.543 ;
      RECT 27.725 4.02 27.73 4.528 ;
      RECT 27.72 4.02 27.725 4.488 ;
      RECT 27.71 4.02 27.72 4.46 ;
      RECT 27.7 4.02 27.71 4.405 ;
      RECT 27.685 4.02 27.7 4.343 ;
      RECT 27.68 4.019 27.685 4.288 ;
      RECT 27.665 4.018 27.68 4.268 ;
      RECT 27.605 4.016 27.665 4.242 ;
      RECT 27.57 4.017 27.605 4.222 ;
      RECT 27.565 4.019 27.57 4.212 ;
      RECT 27.555 4.038 27.565 4.202 ;
      RECT 27.55 4.065 27.555 4.133 ;
      RECT 27.665 3.49 27.835 3.735 ;
      RECT 27.7 3.261 27.835 3.735 ;
      RECT 27.7 3.263 27.845 3.73 ;
      RECT 27.7 3.265 27.87 3.718 ;
      RECT 27.7 3.268 27.895 3.7 ;
      RECT 27.7 3.273 27.945 3.673 ;
      RECT 27.7 3.278 27.965 3.638 ;
      RECT 27.68 3.28 27.975 3.613 ;
      RECT 27.67 3.375 27.975 3.613 ;
      RECT 27.7 3.26 27.81 3.735 ;
      RECT 27.71 3.257 27.805 3.735 ;
      RECT 27.65 7.455 27.82 9.665 ;
      RECT 27.65 7.455 27.825 8.715 ;
      RECT 27.23 4.522 27.42 4.88 ;
      RECT 27.23 4.534 27.455 4.879 ;
      RECT 27.23 4.562 27.475 4.877 ;
      RECT 27.23 4.587 27.48 4.876 ;
      RECT 27.23 4.645 27.495 4.875 ;
      RECT 27.215 4.518 27.375 4.86 ;
      RECT 27.195 4.527 27.42 4.813 ;
      RECT 27.17 4.538 27.455 4.75 ;
      RECT 27.17 4.622 27.49 4.75 ;
      RECT 27.17 4.597 27.485 4.75 ;
      RECT 27.23 4.513 27.375 4.88 ;
      RECT 27.316 4.512 27.375 4.88 ;
      RECT 27.316 4.511 27.36 4.88 ;
      RECT 26.695 10.255 26.87 10.745 ;
      RECT 26.695 7.455 26.865 10.745 ;
      RECT 26.695 9.755 27.105 10.085 ;
      RECT 26.695 8.915 27.105 9.245 ;
      RECT 26.695 7.455 26.87 8.715 ;
      RECT 27.015 4.027 27.02 4.405 ;
      RECT 27.01 3.995 27.015 4.405 ;
      RECT 27.005 3.967 27.01 4.405 ;
      RECT 27 3.947 27.005 4.405 ;
      RECT 26.945 3.93 27 4.405 ;
      RECT 26.905 3.915 26.945 4.405 ;
      RECT 26.85 3.902 26.905 4.405 ;
      RECT 26.815 3.893 26.85 4.405 ;
      RECT 26.811 3.891 26.815 4.404 ;
      RECT 26.725 3.887 26.811 4.387 ;
      RECT 26.64 3.879 26.725 4.35 ;
      RECT 26.63 3.875 26.64 4.323 ;
      RECT 26.62 3.875 26.63 4.305 ;
      RECT 26.61 3.877 26.62 4.288 ;
      RECT 26.605 3.882 26.61 4.274 ;
      RECT 26.6 3.886 26.605 4.261 ;
      RECT 26.59 3.891 26.6 4.245 ;
      RECT 26.575 3.905 26.59 4.22 ;
      RECT 26.57 3.911 26.575 4.2 ;
      RECT 26.565 3.913 26.57 4.193 ;
      RECT 26.56 3.917 26.565 4.068 ;
      RECT 26.74 4.717 26.985 5.18 ;
      RECT 26.66 4.69 26.98 5.176 ;
      RECT 26.59 4.725 26.985 5.169 ;
      RECT 26.38 4.98 26.985 5.165 ;
      RECT 26.56 4.748 26.985 5.165 ;
      RECT 26.4 4.94 26.985 5.165 ;
      RECT 26.55 4.76 26.985 5.165 ;
      RECT 26.435 4.877 26.985 5.165 ;
      RECT 26.49 4.802 26.985 5.165 ;
      RECT 26.74 4.667 26.98 5.18 ;
      RECT 26.77 4.66 26.98 5.18 ;
      RECT 26.76 4.662 26.98 5.18 ;
      RECT 26.77 4.657 26.9 5.18 ;
      RECT 26.325 3.22 26.411 3.659 ;
      RECT 26.32 3.22 26.411 3.657 ;
      RECT 26.32 3.22 26.48 3.656 ;
      RECT 26.32 3.22 26.51 3.653 ;
      RECT 26.305 3.227 26.51 3.644 ;
      RECT 26.305 3.227 26.515 3.64 ;
      RECT 26.3 3.237 26.515 3.633 ;
      RECT 26.295 3.242 26.515 3.608 ;
      RECT 26.295 3.242 26.53 3.59 ;
      RECT 26.32 3.22 26.55 3.505 ;
      RECT 26.29 3.247 26.55 3.503 ;
      RECT 26.3 3.24 26.555 3.441 ;
      RECT 26.29 3.362 26.56 3.424 ;
      RECT 26.275 3.257 26.555 3.375 ;
      RECT 26.27 3.267 26.555 3.275 ;
      RECT 26.35 4.038 26.355 4.115 ;
      RECT 26.34 4.032 26.35 4.305 ;
      RECT 26.33 4.024 26.34 4.326 ;
      RECT 26.32 4.015 26.33 4.348 ;
      RECT 26.315 4.01 26.32 4.365 ;
      RECT 26.275 4.01 26.315 4.405 ;
      RECT 26.255 4.01 26.275 4.46 ;
      RECT 26.25 4.01 26.255 4.488 ;
      RECT 26.24 4.01 26.25 4.503 ;
      RECT 26.205 4.01 26.24 4.545 ;
      RECT 26.2 4.01 26.205 4.588 ;
      RECT 26.19 4.01 26.2 4.603 ;
      RECT 26.175 4.01 26.19 4.623 ;
      RECT 26.16 4.01 26.175 4.65 ;
      RECT 26.155 4.011 26.16 4.668 ;
      RECT 26.135 4.012 26.155 4.675 ;
      RECT 26.08 4.013 26.135 4.695 ;
      RECT 26.07 4.014 26.08 4.709 ;
      RECT 26.065 4.017 26.07 4.708 ;
      RECT 26.025 4.09 26.065 4.706 ;
      RECT 26.01 4.17 26.025 4.704 ;
      RECT 25.985 4.225 26.01 4.702 ;
      RECT 25.97 4.29 25.985 4.701 ;
      RECT 25.925 4.322 25.97 4.698 ;
      RECT 25.84 4.345 25.925 4.693 ;
      RECT 25.815 4.365 25.84 4.688 ;
      RECT 25.745 4.37 25.815 4.684 ;
      RECT 25.725 4.372 25.745 4.681 ;
      RECT 25.64 4.383 25.725 4.675 ;
      RECT 25.635 4.394 25.64 4.67 ;
      RECT 25.625 4.396 25.635 4.67 ;
      RECT 25.59 4.4 25.625 4.668 ;
      RECT 25.54 4.41 25.59 4.655 ;
      RECT 25.52 4.418 25.54 4.64 ;
      RECT 25.44 4.43 25.52 4.623 ;
      RECT 25.605 3.98 25.775 4.19 ;
      RECT 25.721 3.976 25.775 4.19 ;
      RECT 25.526 3.98 25.775 4.181 ;
      RECT 25.526 3.98 25.78 4.17 ;
      RECT 25.44 3.98 25.78 4.161 ;
      RECT 25.44 3.988 25.79 4.105 ;
      RECT 25.44 4 25.795 4.018 ;
      RECT 25.44 4.007 25.8 4.01 ;
      RECT 25.635 3.978 25.775 4.19 ;
      RECT 25.39 4.923 25.635 5.255 ;
      RECT 25.385 4.915 25.39 5.252 ;
      RECT 25.355 4.935 25.635 5.233 ;
      RECT 25.335 4.967 25.635 5.206 ;
      RECT 25.385 4.92 25.562 5.252 ;
      RECT 25.385 4.917 25.476 5.252 ;
      RECT 25.325 3.265 25.495 3.685 ;
      RECT 25.32 3.265 25.495 3.683 ;
      RECT 25.32 3.265 25.52 3.673 ;
      RECT 25.32 3.265 25.54 3.648 ;
      RECT 25.315 3.265 25.54 3.643 ;
      RECT 25.315 3.265 25.55 3.633 ;
      RECT 25.315 3.265 25.555 3.628 ;
      RECT 25.315 3.27 25.56 3.623 ;
      RECT 25.315 3.302 25.575 3.613 ;
      RECT 25.315 3.372 25.6 3.596 ;
      RECT 25.295 3.372 25.6 3.588 ;
      RECT 25.295 3.432 25.61 3.565 ;
      RECT 25.295 3.472 25.62 3.51 ;
      RECT 25.28 3.265 25.555 3.49 ;
      RECT 25.27 3.28 25.56 3.388 ;
      RECT 24.86 4.67 25.03 5.195 ;
      RECT 24.855 4.67 25.03 5.188 ;
      RECT 24.845 4.67 25.035 5.153 ;
      RECT 24.84 4.68 25.035 5.125 ;
      RECT 24.835 4.7 25.035 5.108 ;
      RECT 24.845 4.675 25.04 5.098 ;
      RECT 24.83 4.72 25.04 5.09 ;
      RECT 24.825 4.74 25.04 5.075 ;
      RECT 24.82 4.77 25.04 5.065 ;
      RECT 24.81 4.815 25.04 5.04 ;
      RECT 24.84 4.685 25.045 5.023 ;
      RECT 24.805 4.867 25.045 5.018 ;
      RECT 24.84 4.695 25.05 4.988 ;
      RECT 24.8 4.9 25.05 4.985 ;
      RECT 24.795 4.925 25.05 4.965 ;
      RECT 24.835 4.712 25.06 4.905 ;
      RECT 24.83 4.734 25.07 4.798 ;
      RECT 24.78 3.981 24.795 4.25 ;
      RECT 24.735 3.965 24.78 4.295 ;
      RECT 24.73 3.953 24.735 4.345 ;
      RECT 24.72 3.949 24.73 4.378 ;
      RECT 24.715 3.946 24.72 4.406 ;
      RECT 24.7 3.948 24.715 4.448 ;
      RECT 24.695 3.952 24.7 4.488 ;
      RECT 24.675 3.957 24.695 4.54 ;
      RECT 24.671 3.962 24.675 4.597 ;
      RECT 24.585 3.981 24.671 4.634 ;
      RECT 24.575 4.002 24.585 4.67 ;
      RECT 24.57 4.01 24.575 4.671 ;
      RECT 24.565 4.052 24.57 4.672 ;
      RECT 24.55 4.14 24.565 4.673 ;
      RECT 24.54 4.29 24.55 4.675 ;
      RECT 24.535 4.335 24.54 4.677 ;
      RECT 24.5 4.377 24.535 4.68 ;
      RECT 24.495 4.395 24.5 4.683 ;
      RECT 24.418 4.401 24.495 4.689 ;
      RECT 24.332 4.415 24.418 4.702 ;
      RECT 24.246 4.429 24.332 4.716 ;
      RECT 24.16 4.443 24.246 4.729 ;
      RECT 24.1 4.455 24.16 4.741 ;
      RECT 24.075 4.462 24.1 4.748 ;
      RECT 24.061 4.465 24.075 4.753 ;
      RECT 23.975 4.473 24.061 4.769 ;
      RECT 23.97 4.48 23.975 4.784 ;
      RECT 23.946 4.48 23.97 4.791 ;
      RECT 23.86 4.483 23.946 4.819 ;
      RECT 23.775 4.487 23.86 4.863 ;
      RECT 23.71 4.491 23.775 4.9 ;
      RECT 23.685 4.494 23.71 4.916 ;
      RECT 23.61 4.507 23.685 4.92 ;
      RECT 23.585 4.525 23.61 4.924 ;
      RECT 23.575 4.532 23.585 4.926 ;
      RECT 23.56 4.535 23.575 4.927 ;
      RECT 23.5 4.547 23.56 4.931 ;
      RECT 23.49 4.561 23.5 4.935 ;
      RECT 23.435 4.571 23.49 4.923 ;
      RECT 23.41 4.592 23.435 4.906 ;
      RECT 23.39 4.612 23.41 4.897 ;
      RECT 23.385 4.625 23.39 4.892 ;
      RECT 23.37 4.637 23.385 4.888 ;
      RECT 24.605 3.292 24.61 3.315 ;
      RECT 24.6 3.283 24.605 3.355 ;
      RECT 24.595 3.281 24.6 3.398 ;
      RECT 24.59 3.272 24.595 3.433 ;
      RECT 24.585 3.262 24.59 3.505 ;
      RECT 24.58 3.252 24.585 3.57 ;
      RECT 24.575 3.249 24.58 3.61 ;
      RECT 24.55 3.243 24.575 3.7 ;
      RECT 24.515 3.231 24.55 3.725 ;
      RECT 24.505 3.222 24.515 3.725 ;
      RECT 24.37 3.22 24.38 3.708 ;
      RECT 24.36 3.22 24.37 3.675 ;
      RECT 24.355 3.22 24.36 3.65 ;
      RECT 24.35 3.22 24.355 3.638 ;
      RECT 24.345 3.22 24.35 3.62 ;
      RECT 24.335 3.22 24.345 3.585 ;
      RECT 24.33 3.222 24.335 3.563 ;
      RECT 24.325 3.228 24.33 3.548 ;
      RECT 24.32 3.234 24.325 3.533 ;
      RECT 24.305 3.246 24.32 3.506 ;
      RECT 24.3 3.257 24.305 3.474 ;
      RECT 24.295 3.267 24.3 3.458 ;
      RECT 24.285 3.275 24.295 3.427 ;
      RECT 24.28 3.285 24.285 3.401 ;
      RECT 24.275 3.342 24.28 3.384 ;
      RECT 24.38 3.22 24.505 3.725 ;
      RECT 24.095 3.907 24.355 4.205 ;
      RECT 24.09 3.914 24.355 4.203 ;
      RECT 24.095 3.909 24.37 4.198 ;
      RECT 24.085 3.922 24.37 4.195 ;
      RECT 24.085 3.927 24.375 4.188 ;
      RECT 24.08 3.935 24.375 4.185 ;
      RECT 24.08 3.952 24.38 3.983 ;
      RECT 24.095 3.904 24.326 4.205 ;
      RECT 24.15 3.903 24.326 4.205 ;
      RECT 24.15 3.9 24.24 4.205 ;
      RECT 24.15 3.897 24.236 4.205 ;
      RECT 23.84 4.17 23.845 4.183 ;
      RECT 23.835 4.137 23.84 4.188 ;
      RECT 23.83 4.092 23.835 4.195 ;
      RECT 23.825 4.047 23.83 4.203 ;
      RECT 23.82 4.015 23.825 4.211 ;
      RECT 23.815 3.975 23.82 4.212 ;
      RECT 23.8 3.955 23.815 4.214 ;
      RECT 23.725 3.937 23.8 4.226 ;
      RECT 23.715 3.93 23.725 4.237 ;
      RECT 23.71 3.93 23.715 4.239 ;
      RECT 23.68 3.936 23.71 4.243 ;
      RECT 23.64 3.949 23.68 4.243 ;
      RECT 23.615 3.96 23.64 4.229 ;
      RECT 23.6 3.966 23.615 4.212 ;
      RECT 23.59 3.968 23.6 4.203 ;
      RECT 23.585 3.969 23.59 4.198 ;
      RECT 23.58 3.97 23.585 4.193 ;
      RECT 23.575 3.971 23.58 4.19 ;
      RECT 23.55 3.976 23.575 4.18 ;
      RECT 23.54 3.992 23.55 4.167 ;
      RECT 23.535 4.012 23.54 4.162 ;
      RECT 23.545 3.405 23.55 3.601 ;
      RECT 23.53 3.369 23.545 3.603 ;
      RECT 23.52 3.351 23.53 3.608 ;
      RECT 23.51 3.337 23.52 3.612 ;
      RECT 23.465 3.321 23.51 3.622 ;
      RECT 23.46 3.311 23.465 3.631 ;
      RECT 23.415 3.3 23.46 3.637 ;
      RECT 23.41 3.288 23.415 3.644 ;
      RECT 23.395 3.283 23.41 3.648 ;
      RECT 23.38 3.275 23.395 3.653 ;
      RECT 23.37 3.268 23.38 3.658 ;
      RECT 23.36 3.265 23.37 3.663 ;
      RECT 23.35 3.265 23.36 3.664 ;
      RECT 23.345 3.262 23.35 3.663 ;
      RECT 23.31 3.257 23.335 3.662 ;
      RECT 23.286 3.253 23.31 3.661 ;
      RECT 23.2 3.244 23.286 3.658 ;
      RECT 23.185 3.236 23.2 3.655 ;
      RECT 23.163 3.235 23.185 3.654 ;
      RECT 23.077 3.235 23.163 3.652 ;
      RECT 22.991 3.235 23.077 3.65 ;
      RECT 22.905 3.235 22.991 3.647 ;
      RECT 22.895 3.235 22.905 3.638 ;
      RECT 22.865 3.235 22.895 3.598 ;
      RECT 22.855 3.245 22.865 3.553 ;
      RECT 22.85 3.285 22.855 3.538 ;
      RECT 22.845 3.3 22.85 3.525 ;
      RECT 22.815 3.38 22.845 3.487 ;
      RECT 23.335 3.26 23.345 3.663 ;
      RECT 23.16 4.025 23.175 4.63 ;
      RECT 23.165 4.02 23.175 4.63 ;
      RECT 23.33 4.02 23.335 4.203 ;
      RECT 23.32 4.02 23.33 4.233 ;
      RECT 23.305 4.02 23.32 4.293 ;
      RECT 23.3 4.02 23.305 4.338 ;
      RECT 23.295 4.02 23.3 4.368 ;
      RECT 23.29 4.02 23.295 4.388 ;
      RECT 23.28 4.02 23.29 4.423 ;
      RECT 23.265 4.02 23.28 4.455 ;
      RECT 23.22 4.02 23.265 4.483 ;
      RECT 23.215 4.02 23.22 4.513 ;
      RECT 23.21 4.02 23.215 4.525 ;
      RECT 23.205 4.02 23.21 4.533 ;
      RECT 23.195 4.02 23.205 4.548 ;
      RECT 23.19 4.02 23.195 4.57 ;
      RECT 23.18 4.02 23.19 4.593 ;
      RECT 23.175 4.02 23.18 4.613 ;
      RECT 23.14 4.035 23.16 4.63 ;
      RECT 23.115 4.052 23.14 4.63 ;
      RECT 23.11 4.062 23.115 4.63 ;
      RECT 23.08 4.077 23.11 4.63 ;
      RECT 23.005 4.119 23.08 4.63 ;
      RECT 23 4.15 23.005 4.613 ;
      RECT 22.995 4.154 23 4.595 ;
      RECT 22.99 4.158 22.995 4.558 ;
      RECT 22.985 4.342 22.99 4.525 ;
      RECT 22.47 4.531 22.556 5.096 ;
      RECT 22.425 4.533 22.59 5.09 ;
      RECT 22.556 4.53 22.59 5.09 ;
      RECT 22.47 4.532 22.675 5.084 ;
      RECT 22.425 4.542 22.685 5.08 ;
      RECT 22.4 4.534 22.675 5.076 ;
      RECT 22.395 4.537 22.675 5.071 ;
      RECT 22.37 4.552 22.685 5.065 ;
      RECT 22.37 4.577 22.725 5.06 ;
      RECT 22.33 4.585 22.725 5.035 ;
      RECT 22.33 4.612 22.74 5.033 ;
      RECT 22.33 4.642 22.75 5.02 ;
      RECT 22.325 4.787 22.75 5.008 ;
      RECT 22.33 4.716 22.77 5.005 ;
      RECT 22.33 4.773 22.775 4.813 ;
      RECT 22.52 4.052 22.69 4.23 ;
      RECT 22.47 3.991 22.52 4.215 ;
      RECT 22.205 3.971 22.47 4.2 ;
      RECT 22.165 4.035 22.64 4.2 ;
      RECT 22.165 4.025 22.595 4.2 ;
      RECT 22.165 4.022 22.585 4.2 ;
      RECT 22.165 4.01 22.575 4.2 ;
      RECT 22.165 3.995 22.52 4.2 ;
      RECT 22.205 3.967 22.406 4.2 ;
      RECT 22.215 3.945 22.406 4.2 ;
      RECT 22.24 3.93 22.32 4.2 ;
      RECT 21.995 4.46 22.115 4.905 ;
      RECT 21.98 4.46 22.115 4.904 ;
      RECT 21.935 4.482 22.115 4.899 ;
      RECT 21.895 4.531 22.115 4.893 ;
      RECT 21.895 4.531 22.12 4.868 ;
      RECT 21.895 4.531 22.14 4.758 ;
      RECT 21.89 4.561 22.14 4.755 ;
      RECT 21.98 4.46 22.15 4.65 ;
      RECT 21.64 3.245 21.645 3.69 ;
      RECT 21.45 3.245 21.47 3.655 ;
      RECT 21.42 3.245 21.425 3.63 ;
      RECT 22.1 3.552 22.115 3.74 ;
      RECT 22.095 3.537 22.1 3.746 ;
      RECT 22.075 3.51 22.095 3.749 ;
      RECT 22.025 3.477 22.075 3.758 ;
      RECT 21.995 3.457 22.025 3.762 ;
      RECT 21.976 3.445 21.995 3.758 ;
      RECT 21.89 3.417 21.976 3.748 ;
      RECT 21.88 3.392 21.89 3.738 ;
      RECT 21.81 3.36 21.88 3.73 ;
      RECT 21.785 3.32 21.81 3.722 ;
      RECT 21.765 3.302 21.785 3.716 ;
      RECT 21.755 3.292 21.765 3.713 ;
      RECT 21.745 3.285 21.755 3.711 ;
      RECT 21.725 3.272 21.745 3.708 ;
      RECT 21.715 3.262 21.725 3.705 ;
      RECT 21.705 3.255 21.715 3.703 ;
      RECT 21.655 3.247 21.705 3.697 ;
      RECT 21.645 3.245 21.655 3.691 ;
      RECT 21.615 3.245 21.64 3.688 ;
      RECT 21.586 3.245 21.615 3.683 ;
      RECT 21.5 3.245 21.586 3.673 ;
      RECT 21.47 3.245 21.5 3.66 ;
      RECT 21.425 3.245 21.45 3.643 ;
      RECT 21.41 3.245 21.42 3.625 ;
      RECT 21.39 3.252 21.41 3.61 ;
      RECT 21.385 3.267 21.39 3.598 ;
      RECT 21.38 3.272 21.385 3.538 ;
      RECT 21.375 3.277 21.38 3.38 ;
      RECT 21.37 3.28 21.375 3.298 ;
      RECT 21.11 4.57 21.145 4.89 ;
      RECT 21.695 4.755 21.7 4.937 ;
      RECT 21.65 4.637 21.695 4.956 ;
      RECT 21.635 4.614 21.65 4.979 ;
      RECT 21.625 4.604 21.635 4.989 ;
      RECT 21.605 4.599 21.625 5.002 ;
      RECT 21.58 4.597 21.605 5.023 ;
      RECT 21.561 4.596 21.58 5.035 ;
      RECT 21.475 4.593 21.561 5.035 ;
      RECT 21.405 4.588 21.475 5.023 ;
      RECT 21.33 4.584 21.405 4.998 ;
      RECT 21.265 4.58 21.33 4.965 ;
      RECT 21.195 4.577 21.265 4.925 ;
      RECT 21.165 4.573 21.195 4.9 ;
      RECT 21.145 4.571 21.165 4.893 ;
      RECT 21.061 4.569 21.11 4.891 ;
      RECT 20.975 4.566 21.061 4.892 ;
      RECT 20.9 4.565 20.975 4.894 ;
      RECT 20.815 4.565 20.9 4.92 ;
      RECT 20.738 4.566 20.815 4.945 ;
      RECT 20.652 4.567 20.738 4.945 ;
      RECT 20.566 4.567 20.652 4.945 ;
      RECT 20.48 4.568 20.566 4.945 ;
      RECT 20.46 4.569 20.48 4.937 ;
      RECT 20.445 4.575 20.46 4.922 ;
      RECT 20.41 4.595 20.445 4.902 ;
      RECT 20.4 4.615 20.41 4.884 ;
      RECT 21.37 3.92 21.375 4.19 ;
      RECT 21.365 3.911 21.37 4.195 ;
      RECT 21.355 3.901 21.365 4.207 ;
      RECT 21.35 3.89 21.355 4.218 ;
      RECT 21.33 3.884 21.35 4.236 ;
      RECT 21.285 3.881 21.33 4.285 ;
      RECT 21.27 3.88 21.285 4.33 ;
      RECT 21.265 3.88 21.27 4.343 ;
      RECT 21.255 3.88 21.265 4.355 ;
      RECT 21.25 3.881 21.255 4.37 ;
      RECT 21.23 3.889 21.25 4.375 ;
      RECT 21.2 3.905 21.23 4.375 ;
      RECT 21.19 3.917 21.195 4.375 ;
      RECT 21.155 3.932 21.19 4.375 ;
      RECT 21.125 3.952 21.155 4.375 ;
      RECT 21.115 3.977 21.125 4.375 ;
      RECT 21.11 4.005 21.115 4.375 ;
      RECT 21.105 4.035 21.11 4.375 ;
      RECT 21.1 4.052 21.105 4.375 ;
      RECT 21.09 4.08 21.1 4.375 ;
      RECT 21.08 4.115 21.09 4.375 ;
      RECT 21.075 4.15 21.08 4.375 ;
      RECT 21.195 3.915 21.2 4.375 ;
      RECT 20.185 3.245 20.19 3.644 ;
      RECT 19.93 3.245 19.965 3.642 ;
      RECT 19.525 3.28 19.53 3.636 ;
      RECT 20.27 3.283 20.275 3.538 ;
      RECT 20.265 3.281 20.27 3.544 ;
      RECT 20.26 3.28 20.265 3.551 ;
      RECT 20.235 3.273 20.26 3.575 ;
      RECT 20.23 3.266 20.235 3.599 ;
      RECT 20.225 3.262 20.23 3.608 ;
      RECT 20.215 3.257 20.225 3.621 ;
      RECT 20.21 3.254 20.215 3.63 ;
      RECT 20.205 3.252 20.21 3.635 ;
      RECT 20.19 3.248 20.205 3.645 ;
      RECT 20.175 3.242 20.185 3.644 ;
      RECT 20.137 3.24 20.175 3.644 ;
      RECT 20.051 3.242 20.137 3.644 ;
      RECT 19.965 3.244 20.051 3.643 ;
      RECT 19.894 3.245 19.93 3.642 ;
      RECT 19.808 3.247 19.894 3.642 ;
      RECT 19.722 3.249 19.808 3.641 ;
      RECT 19.636 3.251 19.722 3.641 ;
      RECT 19.55 3.254 19.636 3.64 ;
      RECT 19.54 3.26 19.55 3.639 ;
      RECT 19.53 3.272 19.54 3.637 ;
      RECT 19.47 3.307 19.525 3.633 ;
      RECT 19.465 3.337 19.47 3.395 ;
      RECT 19.81 4.552 19.815 4.809 ;
      RECT 19.79 4.471 19.81 4.826 ;
      RECT 19.77 4.465 19.79 4.855 ;
      RECT 19.71 4.452 19.77 4.875 ;
      RECT 19.665 4.436 19.71 4.876 ;
      RECT 19.581 4.424 19.665 4.864 ;
      RECT 19.495 4.411 19.581 4.848 ;
      RECT 19.485 4.404 19.495 4.84 ;
      RECT 19.44 4.401 19.485 4.78 ;
      RECT 19.42 4.397 19.44 4.695 ;
      RECT 19.405 4.395 19.42 4.648 ;
      RECT 19.375 4.392 19.405 4.618 ;
      RECT 19.34 4.388 19.375 4.595 ;
      RECT 19.297 4.383 19.34 4.583 ;
      RECT 19.211 4.374 19.297 4.592 ;
      RECT 19.125 4.363 19.211 4.604 ;
      RECT 19.06 4.354 19.125 4.613 ;
      RECT 19.04 4.345 19.06 4.618 ;
      RECT 19.035 4.338 19.04 4.62 ;
      RECT 18.995 4.323 19.035 4.617 ;
      RECT 18.975 4.302 18.995 4.612 ;
      RECT 18.96 4.29 18.975 4.605 ;
      RECT 18.955 4.282 18.96 4.598 ;
      RECT 18.94 4.262 18.955 4.591 ;
      RECT 18.935 4.125 18.94 4.585 ;
      RECT 18.855 4.014 18.935 4.557 ;
      RECT 18.846 4.007 18.855 4.523 ;
      RECT 18.76 4.001 18.846 4.448 ;
      RECT 18.735 3.992 18.76 4.36 ;
      RECT 18.705 3.987 18.735 4.335 ;
      RECT 18.64 3.996 18.705 4.32 ;
      RECT 18.62 4.012 18.64 4.295 ;
      RECT 18.61 4.018 18.62 4.243 ;
      RECT 18.59 4.04 18.61 4.125 ;
      RECT 19.245 4.072 19.47 4.19 ;
      RECT 19.245 3.915 19.465 4.19 ;
      RECT 18.46 4.683 18.525 5.126 ;
      RECT 18.4 4.708 18.525 5.124 ;
      RECT 18.4 4.708 18.58 5.118 ;
      RECT 18.385 4.733 18.58 5.117 ;
      RECT 18.525 4.67 18.6 5.114 ;
      RECT 18.46 4.695 18.68 5.108 ;
      RECT 18.385 4.734 18.725 5.102 ;
      RECT 18.37 4.761 18.725 5.093 ;
      RECT 18.385 4.754 18.745 5.085 ;
      RECT 18.37 4.763 18.75 5.068 ;
      RECT 18.365 4.78 18.75 4.895 ;
      RECT 18.37 3.502 18.405 3.74 ;
      RECT 18.37 3.502 18.435 3.739 ;
      RECT 18.37 3.502 18.55 3.735 ;
      RECT 18.37 3.502 18.605 3.713 ;
      RECT 18.38 3.445 18.66 3.613 ;
      RECT 18.485 3.285 18.515 3.736 ;
      RECT 18.515 3.28 18.695 3.493 ;
      RECT 18.385 3.421 18.695 3.493 ;
      RECT 18.435 3.317 18.485 3.737 ;
      RECT 18.405 3.373 18.695 3.493 ;
      RECT 16.62 7.455 16.79 9.665 ;
      RECT 16.62 7.455 16.795 8.715 ;
      RECT 16.19 10.295 16.36 10.745 ;
      RECT 16.25 8.515 16.42 10.465 ;
      RECT 16.19 7.455 16.36 8.685 ;
      RECT 15.665 10.255 15.84 10.745 ;
      RECT 15.665 7.455 15.835 10.745 ;
      RECT 15.665 9.755 16.075 10.085 ;
      RECT 15.665 8.915 16.075 9.245 ;
      RECT 15.665 7.455 15.84 8.715 ;
      RECT 106.89 10.235 107.065 10.745 ;
      RECT 105.9 1.865 106.075 2.375 ;
      RECT 105.9 10.235 106.075 10.745 ;
      RECT 104.11 1.865 104.285 2.375 ;
      RECT 104.11 10.235 104.285 10.745 ;
      RECT 99.35 10.235 99.525 10.745 ;
      RECT 92.07 3.915 92.595 4.19 ;
      RECT 88.965 10.235 89.14 10.745 ;
      RECT 87.975 1.865 88.15 2.375 ;
      RECT 87.975 10.235 88.15 10.745 ;
      RECT 86.185 1.865 86.36 2.375 ;
      RECT 86.185 10.235 86.36 10.745 ;
      RECT 81.425 10.235 81.6 10.745 ;
      RECT 74.145 3.915 74.67 4.19 ;
      RECT 71.04 10.235 71.215 10.745 ;
      RECT 70.05 1.865 70.225 2.375 ;
      RECT 70.05 10.235 70.225 10.745 ;
      RECT 68.26 1.865 68.435 2.375 ;
      RECT 68.26 10.235 68.435 10.745 ;
      RECT 63.5 10.235 63.675 10.745 ;
      RECT 56.22 3.915 56.745 4.19 ;
      RECT 53.115 10.235 53.29 10.745 ;
      RECT 52.125 1.865 52.3 2.375 ;
      RECT 52.125 10.235 52.3 10.745 ;
      RECT 50.335 1.865 50.51 2.375 ;
      RECT 50.335 10.235 50.51 10.745 ;
      RECT 45.575 10.235 45.75 10.745 ;
      RECT 38.295 3.915 38.82 4.19 ;
      RECT 35.19 10.235 35.365 10.745 ;
      RECT 34.2 1.865 34.375 2.375 ;
      RECT 34.2 10.235 34.375 10.745 ;
      RECT 32.41 1.865 32.585 2.375 ;
      RECT 32.41 10.235 32.585 10.745 ;
      RECT 27.65 10.235 27.825 10.745 ;
      RECT 20.37 3.915 20.895 4.19 ;
      RECT 16.62 10.235 16.795 10.745 ;
  END
END sky130_osu_ring_oscillator_mpr2at_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2at_8_b0r2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2at_8_b0r2 ;
  SIZE 107.585 BY 12.61 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 35.23 0 35.61 5.265 ;
      LAYER met2 ;
        RECT 35.23 4.885 35.61 5.265 ;
      LAYER li1 ;
        RECT 35.33 1.865 35.505 2.375 ;
        RECT 35.33 3.895 35.505 5.155 ;
        RECT 35.33 3.685 35.5 5.155 ;
      LAYER met1 ;
        RECT 35.23 4.885 35.61 5.265 ;
        RECT 35.27 2.175 35.565 2.405 ;
        RECT 35.27 3.655 35.56 3.885 ;
        RECT 35.33 2.175 35.5 3.885 ;
      LAYER via1 ;
        RECT 35.345 5 35.495 5.15 ;
      LAYER via2 ;
        RECT 35.32 4.975 35.52 5.175 ;
      LAYER mcon ;
        RECT 35.33 3.685 35.5 3.855 ;
        RECT 35.335 4.985 35.505 5.155 ;
        RECT 35.33 2.205 35.505 2.375 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 53.155 0 53.535 5.265 ;
      LAYER met2 ;
        RECT 53.155 4.885 53.535 5.265 ;
      LAYER li1 ;
        RECT 53.255 1.865 53.43 2.375 ;
        RECT 53.255 3.895 53.43 5.155 ;
        RECT 53.255 3.685 53.425 5.155 ;
      LAYER met1 ;
        RECT 53.155 4.885 53.535 5.265 ;
        RECT 53.195 2.175 53.49 2.405 ;
        RECT 53.195 3.655 53.485 3.885 ;
        RECT 53.255 2.175 53.425 3.885 ;
      LAYER via1 ;
        RECT 53.27 5 53.42 5.15 ;
      LAYER via2 ;
        RECT 53.245 4.975 53.445 5.175 ;
      LAYER mcon ;
        RECT 53.255 3.685 53.425 3.855 ;
        RECT 53.26 4.985 53.43 5.155 ;
        RECT 53.255 2.205 53.43 2.375 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 71.08 0 71.46 5.265 ;
      LAYER met2 ;
        RECT 71.08 4.885 71.46 5.265 ;
      LAYER li1 ;
        RECT 71.18 1.865 71.355 2.375 ;
        RECT 71.18 3.895 71.355 5.155 ;
        RECT 71.18 3.685 71.35 5.155 ;
      LAYER met1 ;
        RECT 71.08 4.885 71.46 5.265 ;
        RECT 71.12 2.175 71.415 2.405 ;
        RECT 71.12 3.655 71.41 3.885 ;
        RECT 71.18 2.175 71.35 3.885 ;
      LAYER via1 ;
        RECT 71.195 5 71.345 5.15 ;
      LAYER via2 ;
        RECT 71.17 4.975 71.37 5.175 ;
      LAYER mcon ;
        RECT 71.18 3.685 71.35 3.855 ;
        RECT 71.185 4.985 71.355 5.155 ;
        RECT 71.18 2.205 71.355 2.375 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 89.005 0 89.385 5.265 ;
      LAYER met2 ;
        RECT 89.005 4.885 89.385 5.265 ;
      LAYER li1 ;
        RECT 89.105 1.865 89.28 2.375 ;
        RECT 89.105 3.895 89.28 5.155 ;
        RECT 89.105 3.685 89.275 5.155 ;
      LAYER met1 ;
        RECT 89.005 4.885 89.385 5.265 ;
        RECT 89.045 2.175 89.34 2.405 ;
        RECT 89.045 3.655 89.335 3.885 ;
        RECT 89.105 2.175 89.275 3.885 ;
      LAYER via1 ;
        RECT 89.12 5 89.27 5.15 ;
      LAYER via2 ;
        RECT 89.095 4.975 89.295 5.175 ;
      LAYER mcon ;
        RECT 89.105 3.685 89.275 3.855 ;
        RECT 89.11 4.985 89.28 5.155 ;
        RECT 89.105 2.205 89.28 2.375 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 106.93 0 107.31 5.265 ;
      LAYER met2 ;
        RECT 106.93 4.885 107.31 5.265 ;
      LAYER li1 ;
        RECT 107.03 1.865 107.205 2.375 ;
        RECT 107.03 3.895 107.205 5.155 ;
        RECT 107.03 3.685 107.2 5.155 ;
      LAYER met1 ;
        RECT 106.93 4.885 107.31 5.265 ;
        RECT 106.97 2.175 107.265 2.405 ;
        RECT 106.97 3.655 107.26 3.885 ;
        RECT 107.03 2.175 107.2 3.885 ;
      LAYER via1 ;
        RECT 107.045 5 107.195 5.15 ;
      LAYER via2 ;
        RECT 107.02 4.975 107.22 5.175 ;
      LAYER mcon ;
        RECT 107.03 3.685 107.2 3.855 ;
        RECT 107.035 4.985 107.205 5.155 ;
        RECT 107.03 2.205 107.205 2.375 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 31.105 4 31.455 4.35 ;
        RECT 31.095 8.275 31.445 8.625 ;
        RECT 31.17 4 31.345 8.625 ;
      LAYER li1 ;
        RECT 31.18 2.955 31.35 4.225 ;
        RECT 31.18 8.385 31.35 9.655 ;
        RECT 26.42 8.385 26.59 9.655 ;
      LAYER met1 ;
        RECT 31.105 4.055 31.58 4.225 ;
        RECT 31.105 4 31.455 4.35 ;
        RECT 31.095 8.385 31.58 8.555 ;
        RECT 31.095 8.275 31.445 8.625 ;
        RECT 26.67 8.38 31.445 8.55 ;
        RECT 26.36 8.385 26.82 8.555 ;
        RECT 26.36 8.355 26.65 8.585 ;
      LAYER via1 ;
        RECT 31.195 8.375 31.345 8.525 ;
        RECT 31.205 4.1 31.355 4.25 ;
      LAYER mcon ;
        RECT 26.42 8.385 26.59 8.555 ;
        RECT 31.18 8.385 31.35 8.555 ;
        RECT 31.18 4.055 31.35 4.225 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 49.03 4 49.38 4.35 ;
        RECT 49.02 8.275 49.37 8.625 ;
        RECT 49.095 4 49.27 8.625 ;
      LAYER li1 ;
        RECT 49.105 2.955 49.275 4.225 ;
        RECT 49.105 8.385 49.275 9.655 ;
        RECT 44.345 8.385 44.515 9.655 ;
      LAYER met1 ;
        RECT 49.03 4.055 49.505 4.225 ;
        RECT 49.03 4 49.38 4.35 ;
        RECT 49.02 8.385 49.505 8.555 ;
        RECT 49.02 8.275 49.37 8.625 ;
        RECT 44.595 8.38 49.37 8.55 ;
        RECT 44.285 8.385 44.745 8.555 ;
        RECT 44.285 8.355 44.575 8.585 ;
      LAYER via1 ;
        RECT 49.12 8.375 49.27 8.525 ;
        RECT 49.13 4.1 49.28 4.25 ;
      LAYER mcon ;
        RECT 44.345 8.385 44.515 8.555 ;
        RECT 49.105 8.385 49.275 8.555 ;
        RECT 49.105 4.055 49.275 4.225 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 66.955 4 67.305 4.35 ;
        RECT 66.945 8.275 67.295 8.625 ;
        RECT 67.02 4 67.195 8.625 ;
      LAYER li1 ;
        RECT 67.03 2.955 67.2 4.225 ;
        RECT 67.03 8.385 67.2 9.655 ;
        RECT 62.27 8.385 62.44 9.655 ;
      LAYER met1 ;
        RECT 66.955 4.055 67.43 4.225 ;
        RECT 66.955 4 67.305 4.35 ;
        RECT 66.945 8.385 67.43 8.555 ;
        RECT 66.945 8.275 67.295 8.625 ;
        RECT 62.52 8.38 67.295 8.55 ;
        RECT 62.21 8.385 62.67 8.555 ;
        RECT 62.21 8.355 62.5 8.585 ;
      LAYER via1 ;
        RECT 67.045 8.375 67.195 8.525 ;
        RECT 67.055 4.1 67.205 4.25 ;
      LAYER mcon ;
        RECT 62.27 8.385 62.44 8.555 ;
        RECT 67.03 8.385 67.2 8.555 ;
        RECT 67.03 4.055 67.2 4.225 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 84.88 4 85.23 4.35 ;
        RECT 84.87 8.275 85.22 8.625 ;
        RECT 84.945 4 85.12 8.625 ;
      LAYER li1 ;
        RECT 84.955 2.955 85.125 4.225 ;
        RECT 84.955 8.385 85.125 9.655 ;
        RECT 80.195 8.385 80.365 9.655 ;
      LAYER met1 ;
        RECT 84.88 4.055 85.355 4.225 ;
        RECT 84.88 4 85.23 4.35 ;
        RECT 84.87 8.385 85.355 8.555 ;
        RECT 84.87 8.275 85.22 8.625 ;
        RECT 80.445 8.38 85.22 8.55 ;
        RECT 80.135 8.385 80.595 8.555 ;
        RECT 80.135 8.355 80.425 8.585 ;
      LAYER via1 ;
        RECT 84.97 8.375 85.12 8.525 ;
        RECT 84.98 4.1 85.13 4.25 ;
      LAYER mcon ;
        RECT 80.195 8.385 80.365 8.555 ;
        RECT 84.955 8.385 85.125 8.555 ;
        RECT 84.955 4.055 85.125 4.225 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 102.805 4 103.155 4.35 ;
        RECT 102.795 8.275 103.145 8.625 ;
        RECT 102.87 4 103.045 8.625 ;
      LAYER li1 ;
        RECT 102.88 2.955 103.05 4.225 ;
        RECT 102.88 8.385 103.05 9.655 ;
        RECT 98.12 8.385 98.29 9.655 ;
      LAYER met1 ;
        RECT 102.805 4.055 103.28 4.225 ;
        RECT 102.805 4 103.155 4.35 ;
        RECT 102.795 8.385 103.28 8.555 ;
        RECT 102.795 8.275 103.145 8.625 ;
        RECT 98.37 8.38 103.145 8.55 ;
        RECT 98.06 8.385 98.52 8.555 ;
        RECT 98.06 8.355 98.35 8.585 ;
      LAYER via1 ;
        RECT 102.895 8.375 103.045 8.525 ;
        RECT 102.905 4.1 103.055 4.25 ;
      LAYER mcon ;
        RECT 98.12 8.385 98.29 8.555 ;
        RECT 102.88 8.385 103.05 8.555 ;
        RECT 102.88 4.055 103.05 4.225 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 15.39 8.385 15.56 9.655 ;
      LAYER met1 ;
        RECT 15.33 8.385 15.79 8.555 ;
        RECT 15.335 8.35 15.625 8.58 ;
        RECT 15.33 8.355 15.62 8.585 ;
      LAYER mcon ;
        RECT 15.39 8.385 15.56 8.555 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.005 5.58 107.58 7.18 ;
        RECT 101.62 5.43 107.58 7.18 ;
        RECT 102.7 5.43 107.425 7.185 ;
        RECT 102.7 5.425 107.42 7.185 ;
        RECT 106.605 5.425 106.775 7.915 ;
        RECT 106.6 4.695 106.77 7.185 ;
        RECT 105.615 4.695 105.785 7.915 ;
        RECT 102.87 4.695 103.04 7.915 ;
        RECT 97.94 5.58 100.69 7.185 ;
        RECT 100.13 5.08 100.3 7.185 ;
        RECT 98.11 5.58 98.28 7.915 ;
        RECT 97.69 5.08 97.86 7.18 ;
        RECT 95.73 5.08 95.9 7.18 ;
        RECT 94.77 5.08 94.94 7.18 ;
        RECT 92.81 5.08 92.98 7.18 ;
        RECT 91.81 5.08 91.98 7.18 ;
        RECT 90.85 5.08 91.02 7.18 ;
        RECT 83.695 5.43 89.655 7.18 ;
        RECT 84.775 5.43 89.5 7.185 ;
        RECT 84.775 5.425 89.495 7.185 ;
        RECT 88.68 5.425 88.85 7.915 ;
        RECT 88.675 4.695 88.845 7.185 ;
        RECT 87.69 4.695 87.86 7.915 ;
        RECT 84.945 4.695 85.115 7.915 ;
        RECT 80.015 5.58 82.765 7.185 ;
        RECT 82.205 5.08 82.375 7.185 ;
        RECT 80.185 5.58 80.355 7.915 ;
        RECT 79.765 5.08 79.935 7.18 ;
        RECT 77.805 5.08 77.975 7.18 ;
        RECT 76.845 5.08 77.015 7.18 ;
        RECT 74.885 5.08 75.055 7.18 ;
        RECT 73.885 5.08 74.055 7.18 ;
        RECT 72.925 5.08 73.095 7.18 ;
        RECT 65.77 5.43 71.73 7.18 ;
        RECT 66.85 5.43 71.575 7.185 ;
        RECT 66.85 5.425 71.57 7.185 ;
        RECT 70.755 5.425 70.925 7.915 ;
        RECT 70.75 4.695 70.92 7.185 ;
        RECT 69.765 4.695 69.935 7.915 ;
        RECT 67.02 4.695 67.19 7.915 ;
        RECT 62.09 5.58 64.84 7.185 ;
        RECT 64.28 5.08 64.45 7.185 ;
        RECT 62.26 5.58 62.43 7.915 ;
        RECT 61.84 5.08 62.01 7.18 ;
        RECT 59.88 5.08 60.05 7.18 ;
        RECT 58.92 5.08 59.09 7.18 ;
        RECT 56.96 5.08 57.13 7.18 ;
        RECT 55.96 5.08 56.13 7.18 ;
        RECT 55 5.08 55.17 7.18 ;
        RECT 47.845 5.43 53.805 7.18 ;
        RECT 48.925 5.43 53.65 7.185 ;
        RECT 48.925 5.425 53.645 7.185 ;
        RECT 52.83 5.425 53 7.915 ;
        RECT 52.825 4.695 52.995 7.185 ;
        RECT 51.84 4.695 52.01 7.915 ;
        RECT 49.095 4.695 49.265 7.915 ;
        RECT 44.165 5.58 46.915 7.185 ;
        RECT 46.355 5.08 46.525 7.185 ;
        RECT 44.335 5.58 44.505 7.915 ;
        RECT 43.915 5.08 44.085 7.18 ;
        RECT 41.955 5.08 42.125 7.18 ;
        RECT 40.995 5.08 41.165 7.18 ;
        RECT 39.035 5.08 39.205 7.18 ;
        RECT 38.035 5.08 38.205 7.18 ;
        RECT 37.075 5.08 37.245 7.18 ;
        RECT 29.92 5.43 35.88 7.18 ;
        RECT 31 5.43 35.725 7.185 ;
        RECT 31 5.425 35.72 7.185 ;
        RECT 34.905 5.425 35.075 7.915 ;
        RECT 34.9 4.695 35.07 7.185 ;
        RECT 33.915 4.695 34.085 7.915 ;
        RECT 31.17 4.695 31.34 7.915 ;
        RECT 26.24 5.58 28.99 7.185 ;
        RECT 28.43 5.08 28.6 7.185 ;
        RECT 26.41 5.58 26.58 7.915 ;
        RECT 25.99 5.08 26.16 7.18 ;
        RECT 24.03 5.08 24.2 7.18 ;
        RECT 23.07 5.08 23.24 7.18 ;
        RECT 21.11 5.08 21.28 7.18 ;
        RECT 20.11 5.08 20.28 7.18 ;
        RECT 19.15 5.08 19.32 7.18 ;
        RECT 15.21 5.58 17.96 7.185 ;
        RECT 17.195 10.195 17.37 10.745 ;
        RECT 17.195 7.455 17.37 8.595 ;
        RECT 17.195 5.58 17.365 10.745 ;
        RECT 15.38 5.58 15.55 7.915 ;
      LAYER met1 ;
        RECT 0.005 5.58 107.58 7.18 ;
        RECT 90.04 5.43 107.58 7.18 ;
        RECT 102.7 5.43 107.425 7.185 ;
        RECT 102.7 5.425 107.42 7.185 ;
        RECT 90.04 5.425 102 7.18 ;
        RECT 97.94 5.425 100.69 7.185 ;
        RECT 72.115 5.43 89.655 7.18 ;
        RECT 84.775 5.43 89.5 7.185 ;
        RECT 84.775 5.425 89.495 7.185 ;
        RECT 72.115 5.425 84.075 7.18 ;
        RECT 80.015 5.425 82.765 7.185 ;
        RECT 54.19 5.43 71.73 7.18 ;
        RECT 66.85 5.43 71.575 7.185 ;
        RECT 66.85 5.425 71.57 7.185 ;
        RECT 54.19 5.425 66.15 7.18 ;
        RECT 62.09 5.425 64.84 7.185 ;
        RECT 36.265 5.43 53.805 7.18 ;
        RECT 48.925 5.43 53.65 7.185 ;
        RECT 48.925 5.425 53.645 7.185 ;
        RECT 36.265 5.425 48.225 7.18 ;
        RECT 44.165 5.425 46.915 7.185 ;
        RECT 18.34 5.43 35.88 7.18 ;
        RECT 31 5.43 35.725 7.185 ;
        RECT 31 5.425 35.72 7.185 ;
        RECT 18.34 5.425 30.3 7.18 ;
        RECT 26.24 5.425 28.99 7.185 ;
        RECT 15.21 5.58 17.96 7.185 ;
        RECT 17.135 9.095 17.425 9.325 ;
        RECT 16.965 9.125 17.425 9.295 ;
      LAYER mcon ;
        RECT 17.195 9.125 17.365 9.295 ;
        RECT 17.5 6.985 17.67 7.155 ;
        RECT 18.485 5.58 18.655 5.75 ;
        RECT 18.945 5.58 19.115 5.75 ;
        RECT 19.405 5.58 19.575 5.75 ;
        RECT 19.865 5.58 20.035 5.75 ;
        RECT 20.325 5.58 20.495 5.75 ;
        RECT 20.785 5.58 20.955 5.75 ;
        RECT 21.245 5.58 21.415 5.75 ;
        RECT 21.705 5.58 21.875 5.75 ;
        RECT 22.165 5.58 22.335 5.75 ;
        RECT 22.625 5.58 22.795 5.75 ;
        RECT 23.085 5.58 23.255 5.75 ;
        RECT 23.545 5.58 23.715 5.75 ;
        RECT 24.005 5.58 24.175 5.75 ;
        RECT 24.465 5.58 24.635 5.75 ;
        RECT 24.925 5.58 25.095 5.75 ;
        RECT 25.385 5.58 25.555 5.75 ;
        RECT 25.845 5.58 26.015 5.75 ;
        RECT 26.305 5.58 26.475 5.75 ;
        RECT 26.765 5.58 26.935 5.75 ;
        RECT 27.225 5.58 27.395 5.75 ;
        RECT 27.685 5.58 27.855 5.75 ;
        RECT 28.145 5.58 28.315 5.75 ;
        RECT 28.53 6.985 28.7 7.155 ;
        RECT 28.605 5.58 28.775 5.75 ;
        RECT 29.065 5.58 29.235 5.75 ;
        RECT 29.525 5.58 29.695 5.75 ;
        RECT 29.985 5.58 30.155 5.75 ;
        RECT 33.29 6.985 33.46 7.155 ;
        RECT 33.29 5.455 33.46 5.625 ;
        RECT 33.995 6.985 34.165 7.155 ;
        RECT 33.995 5.455 34.165 5.625 ;
        RECT 34.98 5.455 35.15 5.625 ;
        RECT 34.985 6.985 35.155 7.155 ;
        RECT 36.41 5.58 36.58 5.75 ;
        RECT 36.87 5.58 37.04 5.75 ;
        RECT 37.33 5.58 37.5 5.75 ;
        RECT 37.79 5.58 37.96 5.75 ;
        RECT 38.25 5.58 38.42 5.75 ;
        RECT 38.71 5.58 38.88 5.75 ;
        RECT 39.17 5.58 39.34 5.75 ;
        RECT 39.63 5.58 39.8 5.75 ;
        RECT 40.09 5.58 40.26 5.75 ;
        RECT 40.55 5.58 40.72 5.75 ;
        RECT 41.01 5.58 41.18 5.75 ;
        RECT 41.47 5.58 41.64 5.75 ;
        RECT 41.93 5.58 42.1 5.75 ;
        RECT 42.39 5.58 42.56 5.75 ;
        RECT 42.85 5.58 43.02 5.75 ;
        RECT 43.31 5.58 43.48 5.75 ;
        RECT 43.77 5.58 43.94 5.75 ;
        RECT 44.23 5.58 44.4 5.75 ;
        RECT 44.69 5.58 44.86 5.75 ;
        RECT 45.15 5.58 45.32 5.75 ;
        RECT 45.61 5.58 45.78 5.75 ;
        RECT 46.07 5.58 46.24 5.75 ;
        RECT 46.455 6.985 46.625 7.155 ;
        RECT 46.53 5.58 46.7 5.75 ;
        RECT 46.99 5.58 47.16 5.75 ;
        RECT 47.45 5.58 47.62 5.75 ;
        RECT 47.91 5.58 48.08 5.75 ;
        RECT 51.215 6.985 51.385 7.155 ;
        RECT 51.215 5.455 51.385 5.625 ;
        RECT 51.92 6.985 52.09 7.155 ;
        RECT 51.92 5.455 52.09 5.625 ;
        RECT 52.905 5.455 53.075 5.625 ;
        RECT 52.91 6.985 53.08 7.155 ;
        RECT 54.335 5.58 54.505 5.75 ;
        RECT 54.795 5.58 54.965 5.75 ;
        RECT 55.255 5.58 55.425 5.75 ;
        RECT 55.715 5.58 55.885 5.75 ;
        RECT 56.175 5.58 56.345 5.75 ;
        RECT 56.635 5.58 56.805 5.75 ;
        RECT 57.095 5.58 57.265 5.75 ;
        RECT 57.555 5.58 57.725 5.75 ;
        RECT 58.015 5.58 58.185 5.75 ;
        RECT 58.475 5.58 58.645 5.75 ;
        RECT 58.935 5.58 59.105 5.75 ;
        RECT 59.395 5.58 59.565 5.75 ;
        RECT 59.855 5.58 60.025 5.75 ;
        RECT 60.315 5.58 60.485 5.75 ;
        RECT 60.775 5.58 60.945 5.75 ;
        RECT 61.235 5.58 61.405 5.75 ;
        RECT 61.695 5.58 61.865 5.75 ;
        RECT 62.155 5.58 62.325 5.75 ;
        RECT 62.615 5.58 62.785 5.75 ;
        RECT 63.075 5.58 63.245 5.75 ;
        RECT 63.535 5.58 63.705 5.75 ;
        RECT 63.995 5.58 64.165 5.75 ;
        RECT 64.38 6.985 64.55 7.155 ;
        RECT 64.455 5.58 64.625 5.75 ;
        RECT 64.915 5.58 65.085 5.75 ;
        RECT 65.375 5.58 65.545 5.75 ;
        RECT 65.835 5.58 66.005 5.75 ;
        RECT 69.14 6.985 69.31 7.155 ;
        RECT 69.14 5.455 69.31 5.625 ;
        RECT 69.845 6.985 70.015 7.155 ;
        RECT 69.845 5.455 70.015 5.625 ;
        RECT 70.83 5.455 71 5.625 ;
        RECT 70.835 6.985 71.005 7.155 ;
        RECT 72.26 5.58 72.43 5.75 ;
        RECT 72.72 5.58 72.89 5.75 ;
        RECT 73.18 5.58 73.35 5.75 ;
        RECT 73.64 5.58 73.81 5.75 ;
        RECT 74.1 5.58 74.27 5.75 ;
        RECT 74.56 5.58 74.73 5.75 ;
        RECT 75.02 5.58 75.19 5.75 ;
        RECT 75.48 5.58 75.65 5.75 ;
        RECT 75.94 5.58 76.11 5.75 ;
        RECT 76.4 5.58 76.57 5.75 ;
        RECT 76.86 5.58 77.03 5.75 ;
        RECT 77.32 5.58 77.49 5.75 ;
        RECT 77.78 5.58 77.95 5.75 ;
        RECT 78.24 5.58 78.41 5.75 ;
        RECT 78.7 5.58 78.87 5.75 ;
        RECT 79.16 5.58 79.33 5.75 ;
        RECT 79.62 5.58 79.79 5.75 ;
        RECT 80.08 5.58 80.25 5.75 ;
        RECT 80.54 5.58 80.71 5.75 ;
        RECT 81 5.58 81.17 5.75 ;
        RECT 81.46 5.58 81.63 5.75 ;
        RECT 81.92 5.58 82.09 5.75 ;
        RECT 82.305 6.985 82.475 7.155 ;
        RECT 82.38 5.58 82.55 5.75 ;
        RECT 82.84 5.58 83.01 5.75 ;
        RECT 83.3 5.58 83.47 5.75 ;
        RECT 83.76 5.58 83.93 5.75 ;
        RECT 87.065 6.985 87.235 7.155 ;
        RECT 87.065 5.455 87.235 5.625 ;
        RECT 87.77 6.985 87.94 7.155 ;
        RECT 87.77 5.455 87.94 5.625 ;
        RECT 88.755 5.455 88.925 5.625 ;
        RECT 88.76 6.985 88.93 7.155 ;
        RECT 90.185 5.58 90.355 5.75 ;
        RECT 90.645 5.58 90.815 5.75 ;
        RECT 91.105 5.58 91.275 5.75 ;
        RECT 91.565 5.58 91.735 5.75 ;
        RECT 92.025 5.58 92.195 5.75 ;
        RECT 92.485 5.58 92.655 5.75 ;
        RECT 92.945 5.58 93.115 5.75 ;
        RECT 93.405 5.58 93.575 5.75 ;
        RECT 93.865 5.58 94.035 5.75 ;
        RECT 94.325 5.58 94.495 5.75 ;
        RECT 94.785 5.58 94.955 5.75 ;
        RECT 95.245 5.58 95.415 5.75 ;
        RECT 95.705 5.58 95.875 5.75 ;
        RECT 96.165 5.58 96.335 5.75 ;
        RECT 96.625 5.58 96.795 5.75 ;
        RECT 97.085 5.58 97.255 5.75 ;
        RECT 97.545 5.58 97.715 5.75 ;
        RECT 98.005 5.58 98.175 5.75 ;
        RECT 98.465 5.58 98.635 5.75 ;
        RECT 98.925 5.58 99.095 5.75 ;
        RECT 99.385 5.58 99.555 5.75 ;
        RECT 99.845 5.58 100.015 5.75 ;
        RECT 100.23 6.985 100.4 7.155 ;
        RECT 100.305 5.58 100.475 5.75 ;
        RECT 100.765 5.58 100.935 5.75 ;
        RECT 101.225 5.58 101.395 5.75 ;
        RECT 101.685 5.58 101.855 5.75 ;
        RECT 104.99 6.985 105.16 7.155 ;
        RECT 104.99 5.455 105.16 5.625 ;
        RECT 105.695 6.985 105.865 7.155 ;
        RECT 105.695 5.455 105.865 5.625 ;
        RECT 106.68 5.455 106.85 5.625 ;
        RECT 106.685 6.985 106.855 7.155 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 91.655 3.86 92.385 4.19 ;
        RECT 73.73 3.86 74.46 4.19 ;
        RECT 55.805 3.86 56.535 4.19 ;
        RECT 37.88 3.86 38.61 4.19 ;
        RECT 19.955 3.86 20.685 4.19 ;
      LAYER met2 ;
        RECT 93.33 3.93 93.59 4.19 ;
        RECT 91.96 3.91 93.37 4.125 ;
        RECT 91.96 3.885 92.45 4.165 ;
        RECT 91.99 3.885 92.415 4.205 ;
        RECT 91.99 3.885 92.395 4.225 ;
        RECT 91.99 3.885 92.37 4.235 ;
        RECT 92 2.5 92.345 2.845 ;
        RECT 91.99 3.885 92.295 4.255 ;
        RECT 91.99 3.885 92.27 4.335 ;
        RECT 92.095 2.5 92.265 4.335 ;
        RECT 91.99 3.885 92.245 4.35 ;
        RECT 91.96 4.41 92.22 4.67 ;
        RECT 91.99 3.885 92.24 4.415 ;
        RECT 75.405 3.93 75.665 4.19 ;
        RECT 74.035 3.91 75.445 4.125 ;
        RECT 74.035 3.885 74.525 4.165 ;
        RECT 74.065 3.885 74.49 4.205 ;
        RECT 74.065 3.885 74.47 4.225 ;
        RECT 74.065 3.885 74.445 4.235 ;
        RECT 74.075 2.5 74.42 2.845 ;
        RECT 74.065 3.885 74.37 4.255 ;
        RECT 74.065 3.885 74.345 4.335 ;
        RECT 74.17 2.5 74.34 4.335 ;
        RECT 74.065 3.885 74.32 4.35 ;
        RECT 74.035 4.41 74.295 4.67 ;
        RECT 74.065 3.885 74.315 4.415 ;
        RECT 57.48 3.93 57.74 4.19 ;
        RECT 56.11 3.91 57.52 4.125 ;
        RECT 56.11 3.885 56.6 4.165 ;
        RECT 56.14 3.885 56.565 4.205 ;
        RECT 56.14 3.885 56.545 4.225 ;
        RECT 56.14 3.885 56.52 4.235 ;
        RECT 56.15 2.5 56.495 2.845 ;
        RECT 56.14 3.885 56.445 4.255 ;
        RECT 56.14 3.885 56.42 4.335 ;
        RECT 56.245 2.5 56.415 4.335 ;
        RECT 56.14 3.885 56.395 4.35 ;
        RECT 56.11 4.41 56.37 4.67 ;
        RECT 56.14 3.885 56.39 4.415 ;
        RECT 39.555 3.93 39.815 4.19 ;
        RECT 38.185 3.91 39.595 4.125 ;
        RECT 38.185 3.885 38.675 4.165 ;
        RECT 38.215 3.885 38.64 4.205 ;
        RECT 38.215 3.885 38.62 4.225 ;
        RECT 38.215 3.885 38.595 4.235 ;
        RECT 38.225 2.5 38.57 2.845 ;
        RECT 38.215 3.885 38.52 4.255 ;
        RECT 38.215 3.885 38.495 4.335 ;
        RECT 38.32 2.5 38.49 4.335 ;
        RECT 38.215 3.885 38.47 4.35 ;
        RECT 38.185 4.41 38.445 4.67 ;
        RECT 38.215 3.885 38.465 4.415 ;
        RECT 21.63 3.93 21.89 4.19 ;
        RECT 20.26 3.91 21.67 4.125 ;
        RECT 20.26 3.885 20.75 4.165 ;
        RECT 20.29 3.885 20.715 4.205 ;
        RECT 20.29 3.885 20.695 4.225 ;
        RECT 20.29 3.885 20.67 4.235 ;
        RECT 20.3 2.5 20.645 2.845 ;
        RECT 20.29 3.885 20.595 4.255 ;
        RECT 20.29 3.885 20.57 4.335 ;
        RECT 20.395 2.5 20.565 4.335 ;
        RECT 20.29 3.885 20.545 4.35 ;
        RECT 20.26 4.41 20.52 4.67 ;
        RECT 20.29 3.885 20.54 4.415 ;
      LAYER li1 ;
        RECT 0.03 11.445 107.585 12.61 ;
        RECT 0.035 11.01 107.585 12.61 ;
        RECT 106.605 10.385 106.775 12.61 ;
        RECT 105.615 10.385 105.785 12.61 ;
        RECT 102.87 10.385 103.04 12.61 ;
        RECT 98.11 10.385 98.28 12.61 ;
        RECT 88.68 10.385 88.85 12.61 ;
        RECT 87.69 10.385 87.86 12.61 ;
        RECT 84.945 10.385 85.115 12.61 ;
        RECT 80.185 10.385 80.355 12.61 ;
        RECT 70.755 10.385 70.925 12.61 ;
        RECT 69.765 10.385 69.935 12.61 ;
        RECT 67.02 10.385 67.19 12.61 ;
        RECT 62.26 10.385 62.43 12.61 ;
        RECT 52.83 10.385 53 12.61 ;
        RECT 51.84 10.385 52.01 12.61 ;
        RECT 49.095 10.385 49.265 12.61 ;
        RECT 44.335 10.385 44.505 12.61 ;
        RECT 34.905 10.385 35.075 12.61 ;
        RECT 33.915 10.385 34.085 12.61 ;
        RECT 31.17 10.385 31.34 12.61 ;
        RECT 26.41 10.385 26.58 12.61 ;
        RECT 15.38 10.385 15.55 12.61 ;
        RECT 0 0 107.58 1.6 ;
        RECT 106.6 0 106.77 2.225 ;
        RECT 105.615 0 105.785 2.225 ;
        RECT 102.87 0 103.04 2.225 ;
        RECT 90.04 2.86 102 3.03 ;
        RECT 90.025 0 101.935 2.975 ;
        RECT 101.09 0 101.26 3.53 ;
        RECT 100.13 0 100.3 3.53 ;
        RECT 99.17 0 99.34 3.53 ;
        RECT 98.65 0 98.82 3.53 ;
        RECT 97.69 0 97.86 3.53 ;
        RECT 96.69 0 96.86 3.53 ;
        RECT 95.73 0 95.9 3.53 ;
        RECT 94.25 0 94.42 3.53 ;
        RECT 92.33 0 92.5 3.53 ;
        RECT 90.85 0 91.02 3.53 ;
        RECT 88.675 0 88.845 2.225 ;
        RECT 87.69 0 87.86 2.225 ;
        RECT 84.945 0 85.115 2.225 ;
        RECT 72.115 2.86 84.075 3.03 ;
        RECT 72.1 0 84.01 2.975 ;
        RECT 83.165 0 83.335 3.53 ;
        RECT 82.205 0 82.375 3.53 ;
        RECT 81.245 0 81.415 3.53 ;
        RECT 80.725 0 80.895 3.53 ;
        RECT 79.765 0 79.935 3.53 ;
        RECT 78.765 0 78.935 3.53 ;
        RECT 77.805 0 77.975 3.53 ;
        RECT 76.325 0 76.495 3.53 ;
        RECT 74.405 0 74.575 3.53 ;
        RECT 72.925 0 73.095 3.53 ;
        RECT 70.75 0 70.92 2.225 ;
        RECT 69.765 0 69.935 2.225 ;
        RECT 67.02 0 67.19 2.225 ;
        RECT 54.19 2.86 66.15 3.03 ;
        RECT 54.175 0 66.085 2.975 ;
        RECT 65.24 0 65.41 3.53 ;
        RECT 64.28 0 64.45 3.53 ;
        RECT 63.32 0 63.49 3.53 ;
        RECT 62.8 0 62.97 3.53 ;
        RECT 61.84 0 62.01 3.53 ;
        RECT 60.84 0 61.01 3.53 ;
        RECT 59.88 0 60.05 3.53 ;
        RECT 58.4 0 58.57 3.53 ;
        RECT 56.48 0 56.65 3.53 ;
        RECT 55 0 55.17 3.53 ;
        RECT 52.825 0 52.995 2.225 ;
        RECT 51.84 0 52.01 2.225 ;
        RECT 49.095 0 49.265 2.225 ;
        RECT 36.265 2.86 48.225 3.03 ;
        RECT 36.25 0 48.16 2.975 ;
        RECT 47.315 0 47.485 3.53 ;
        RECT 46.355 0 46.525 3.53 ;
        RECT 45.395 0 45.565 3.53 ;
        RECT 44.875 0 45.045 3.53 ;
        RECT 43.915 0 44.085 3.53 ;
        RECT 42.915 0 43.085 3.53 ;
        RECT 41.955 0 42.125 3.53 ;
        RECT 40.475 0 40.645 3.53 ;
        RECT 38.555 0 38.725 3.53 ;
        RECT 37.075 0 37.245 3.53 ;
        RECT 34.9 0 35.07 2.225 ;
        RECT 33.915 0 34.085 2.225 ;
        RECT 31.17 0 31.34 2.225 ;
        RECT 18.34 2.86 30.3 3.03 ;
        RECT 18.325 0 30.235 2.975 ;
        RECT 29.39 0 29.56 3.53 ;
        RECT 28.43 0 28.6 3.53 ;
        RECT 27.47 0 27.64 3.53 ;
        RECT 26.95 0 27.12 3.53 ;
        RECT 25.99 0 26.16 3.53 ;
        RECT 24.99 0 25.16 3.53 ;
        RECT 24.03 0 24.2 3.53 ;
        RECT 22.55 0 22.72 3.53 ;
        RECT 20.63 0 20.8 3.53 ;
        RECT 19.15 0 19.32 3.53 ;
        RECT 99.125 8.515 99.295 10.465 ;
        RECT 99.065 10.295 99.235 10.745 ;
        RECT 99.065 7.455 99.235 8.685 ;
        RECT 93.43 3.96 93.74 4.265 ;
        RECT 93.43 3.96 93.72 4.29 ;
        RECT 91.87 4.21 92.07 4.61 ;
        RECT 91.555 3.995 92.025 4.245 ;
        RECT 91.865 4.21 92.07 4.43 ;
        RECT 91.86 4.21 92.07 4.395 ;
        RECT 91.84 4.21 92.07 4.375 ;
        RECT 91.835 4.21 92.07 4.35 ;
        RECT 91.81 4.21 92.07 4.345 ;
        RECT 91.74 4.21 92.07 4.34 ;
        RECT 91.725 4.21 92.07 4.32 ;
        RECT 91.695 4.21 92.07 4.31 ;
        RECT 91.69 4.21 92.07 4.285 ;
        RECT 91.64 4.21 92.07 4.28 ;
        RECT 81.2 8.515 81.37 10.465 ;
        RECT 81.14 10.295 81.31 10.745 ;
        RECT 81.14 7.455 81.31 8.685 ;
        RECT 75.505 3.96 75.815 4.265 ;
        RECT 75.505 3.96 75.795 4.29 ;
        RECT 73.945 4.21 74.145 4.61 ;
        RECT 73.63 3.995 74.1 4.245 ;
        RECT 73.94 4.21 74.145 4.43 ;
        RECT 73.935 4.21 74.145 4.395 ;
        RECT 73.915 4.21 74.145 4.375 ;
        RECT 73.91 4.21 74.145 4.35 ;
        RECT 73.885 4.21 74.145 4.345 ;
        RECT 73.815 4.21 74.145 4.34 ;
        RECT 73.8 4.21 74.145 4.32 ;
        RECT 73.77 4.21 74.145 4.31 ;
        RECT 73.765 4.21 74.145 4.285 ;
        RECT 73.715 4.21 74.145 4.28 ;
        RECT 63.275 8.515 63.445 10.465 ;
        RECT 63.215 10.295 63.385 10.745 ;
        RECT 63.215 7.455 63.385 8.685 ;
        RECT 57.58 3.96 57.89 4.265 ;
        RECT 57.58 3.96 57.87 4.29 ;
        RECT 56.02 4.21 56.22 4.61 ;
        RECT 55.705 3.995 56.175 4.245 ;
        RECT 56.015 4.21 56.22 4.43 ;
        RECT 56.01 4.21 56.22 4.395 ;
        RECT 55.99 4.21 56.22 4.375 ;
        RECT 55.985 4.21 56.22 4.35 ;
        RECT 55.96 4.21 56.22 4.345 ;
        RECT 55.89 4.21 56.22 4.34 ;
        RECT 55.875 4.21 56.22 4.32 ;
        RECT 55.845 4.21 56.22 4.31 ;
        RECT 55.84 4.21 56.22 4.285 ;
        RECT 55.79 4.21 56.22 4.28 ;
        RECT 45.35 8.515 45.52 10.465 ;
        RECT 45.29 10.295 45.46 10.745 ;
        RECT 45.29 7.455 45.46 8.685 ;
        RECT 39.655 3.96 39.965 4.265 ;
        RECT 39.655 3.96 39.945 4.29 ;
        RECT 38.095 4.21 38.295 4.61 ;
        RECT 37.78 3.995 38.25 4.245 ;
        RECT 38.09 4.21 38.295 4.43 ;
        RECT 38.085 4.21 38.295 4.395 ;
        RECT 38.065 4.21 38.295 4.375 ;
        RECT 38.06 4.21 38.295 4.35 ;
        RECT 38.035 4.21 38.295 4.345 ;
        RECT 37.965 4.21 38.295 4.34 ;
        RECT 37.95 4.21 38.295 4.32 ;
        RECT 37.92 4.21 38.295 4.31 ;
        RECT 37.915 4.21 38.295 4.285 ;
        RECT 37.865 4.21 38.295 4.28 ;
        RECT 27.425 8.515 27.595 10.465 ;
        RECT 27.365 10.295 27.535 10.745 ;
        RECT 27.365 7.455 27.535 8.685 ;
        RECT 21.73 3.96 22.04 4.265 ;
        RECT 21.73 3.96 22.02 4.29 ;
        RECT 20.17 4.21 20.37 4.61 ;
        RECT 19.855 3.995 20.325 4.245 ;
        RECT 20.165 4.21 20.37 4.43 ;
        RECT 20.16 4.21 20.37 4.395 ;
        RECT 20.14 4.21 20.37 4.375 ;
        RECT 20.135 4.21 20.37 4.35 ;
        RECT 20.11 4.21 20.37 4.345 ;
        RECT 20.04 4.21 20.37 4.34 ;
        RECT 20.025 4.21 20.37 4.32 ;
        RECT 19.995 4.21 20.37 4.31 ;
        RECT 19.99 4.21 20.37 4.285 ;
        RECT 19.94 4.21 20.37 4.28 ;
      LAYER met1 ;
        RECT 0.035 11.01 107.585 12.61 ;
        RECT 99.065 8.725 99.355 8.955 ;
        RECT 98.725 8.75 99.355 8.925 ;
        RECT 98.725 8.75 98.895 12.61 ;
        RECT 81.14 8.725 81.43 8.955 ;
        RECT 80.8 8.75 81.43 8.925 ;
        RECT 80.8 8.75 80.97 12.61 ;
        RECT 63.215 8.725 63.505 8.955 ;
        RECT 62.875 8.75 63.505 8.925 ;
        RECT 62.875 8.75 63.045 12.61 ;
        RECT 45.29 8.725 45.58 8.955 ;
        RECT 44.95 8.75 45.58 8.925 ;
        RECT 44.95 8.75 45.12 12.61 ;
        RECT 27.365 8.725 27.655 8.955 ;
        RECT 27.025 8.75 27.655 8.925 ;
        RECT 27.025 8.75 27.195 12.61 ;
        RECT 0 0 107.58 1.6 ;
        RECT 90.04 2.705 102 3.185 ;
        RECT 90.025 2.58 101.935 2.975 ;
        RECT 94.455 0 101.935 3.185 ;
        RECT 91.05 0 101.935 2.3 ;
        RECT 93.02 0 94.175 3.185 ;
        RECT 90.025 2.55 92.74 2.975 ;
        RECT 91.05 0 92.74 3.185 ;
        RECT 90.025 0 101.935 2.27 ;
        RECT 90.025 0 90.77 2.975 ;
        RECT 72.115 2.705 84.075 3.185 ;
        RECT 72.1 2.58 84.01 2.975 ;
        RECT 76.53 0 84.01 3.185 ;
        RECT 73.125 0 84.01 2.3 ;
        RECT 75.095 0 76.25 3.185 ;
        RECT 72.1 2.55 74.815 2.975 ;
        RECT 73.125 0 74.815 3.185 ;
        RECT 72.1 0 84.01 2.27 ;
        RECT 72.1 0 72.845 2.975 ;
        RECT 54.19 2.705 66.15 3.185 ;
        RECT 54.175 2.58 66.085 2.975 ;
        RECT 58.605 0 66.085 3.185 ;
        RECT 55.2 0 66.085 2.3 ;
        RECT 57.17 0 58.325 3.185 ;
        RECT 54.175 2.55 56.89 2.975 ;
        RECT 55.2 0 56.89 3.185 ;
        RECT 54.175 0 66.085 2.27 ;
        RECT 54.175 0 54.92 2.975 ;
        RECT 36.265 2.705 48.225 3.185 ;
        RECT 36.25 2.58 48.16 2.975 ;
        RECT 40.68 0 48.16 3.185 ;
        RECT 37.275 0 48.16 2.3 ;
        RECT 39.245 0 40.4 3.185 ;
        RECT 36.25 2.55 38.965 2.975 ;
        RECT 37.275 0 38.965 3.185 ;
        RECT 36.25 0 48.16 2.27 ;
        RECT 36.25 0 36.995 2.975 ;
        RECT 18.34 2.705 30.3 3.185 ;
        RECT 18.325 2.46 30.235 2.975 ;
        RECT 22.755 0 30.235 3.185 ;
        RECT 19.35 0 30.235 2.3 ;
        RECT 21.32 0 22.475 3.185 ;
        RECT 19.35 0 21.04 3.185 ;
        RECT 18.325 0 30.235 2.27 ;
        RECT 18.325 0 19.07 2.975 ;
        RECT 93.33 3.94 93.62 4.155 ;
        RECT 93.33 3.93 93.59 4.19 ;
        RECT 91.96 4.41 92.22 4.67 ;
        RECT 91.88 4.42 92.22 4.63 ;
        RECT 75.405 3.94 75.695 4.155 ;
        RECT 75.405 3.93 75.665 4.19 ;
        RECT 74.035 4.41 74.295 4.67 ;
        RECT 73.955 4.42 74.295 4.63 ;
        RECT 57.48 3.94 57.77 4.155 ;
        RECT 57.48 3.93 57.74 4.19 ;
        RECT 56.11 4.41 56.37 4.67 ;
        RECT 56.03 4.42 56.37 4.63 ;
        RECT 39.555 3.94 39.845 4.155 ;
        RECT 39.555 3.93 39.815 4.19 ;
        RECT 38.185 4.41 38.445 4.67 ;
        RECT 38.105 4.42 38.445 4.63 ;
        RECT 21.63 3.94 21.92 4.155 ;
        RECT 21.63 3.93 21.89 4.19 ;
        RECT 20.26 4.41 20.52 4.67 ;
        RECT 20.18 4.42 20.52 4.63 ;
      LAYER via1 ;
        RECT 20.315 4.465 20.465 4.615 ;
        RECT 20.395 2.595 20.545 2.745 ;
        RECT 21.685 3.985 21.835 4.135 ;
        RECT 38.24 4.465 38.39 4.615 ;
        RECT 38.32 2.595 38.47 2.745 ;
        RECT 39.61 3.985 39.76 4.135 ;
        RECT 56.165 4.465 56.315 4.615 ;
        RECT 56.245 2.595 56.395 2.745 ;
        RECT 57.535 3.985 57.685 4.135 ;
        RECT 74.09 4.465 74.24 4.615 ;
        RECT 74.17 2.595 74.32 2.745 ;
        RECT 75.46 3.985 75.61 4.135 ;
        RECT 92.015 4.465 92.165 4.615 ;
        RECT 92.095 2.595 92.245 2.745 ;
        RECT 93.385 3.985 93.535 4.135 ;
      LAYER via2 ;
        RECT 20.345 3.925 20.555 4.125 ;
        RECT 38.27 3.925 38.48 4.125 ;
        RECT 56.195 3.925 56.405 4.125 ;
        RECT 74.12 3.925 74.33 4.125 ;
        RECT 92.045 3.925 92.255 4.125 ;
      LAYER mcon ;
        RECT 15.46 11.045 15.63 11.215 ;
        RECT 16.14 11.045 16.31 11.215 ;
        RECT 16.82 11.045 16.99 11.215 ;
        RECT 17.5 11.045 17.67 11.215 ;
        RECT 18.485 2.86 18.655 3.03 ;
        RECT 18.945 2.86 19.115 3.03 ;
        RECT 19.405 2.86 19.575 3.03 ;
        RECT 19.865 2.86 20.035 3.03 ;
        RECT 20.2 4.44 20.37 4.61 ;
        RECT 20.325 2.86 20.495 3.03 ;
        RECT 20.785 2.86 20.955 3.03 ;
        RECT 21.245 2.86 21.415 3.03 ;
        RECT 21.705 2.86 21.875 3.03 ;
        RECT 21.73 3.965 21.9 4.135 ;
        RECT 22.165 2.86 22.335 3.03 ;
        RECT 22.625 2.86 22.795 3.03 ;
        RECT 23.085 2.86 23.255 3.03 ;
        RECT 23.545 2.86 23.715 3.03 ;
        RECT 24.005 2.86 24.175 3.03 ;
        RECT 24.465 2.86 24.635 3.03 ;
        RECT 24.925 2.86 25.095 3.03 ;
        RECT 25.385 2.86 25.555 3.03 ;
        RECT 25.845 2.86 26.015 3.03 ;
        RECT 26.305 2.86 26.475 3.03 ;
        RECT 26.49 11.045 26.66 11.215 ;
        RECT 26.765 2.86 26.935 3.03 ;
        RECT 27.17 11.045 27.34 11.215 ;
        RECT 27.225 2.86 27.395 3.03 ;
        RECT 27.425 8.755 27.595 8.925 ;
        RECT 27.685 2.86 27.855 3.03 ;
        RECT 27.85 11.045 28.02 11.215 ;
        RECT 28.145 2.86 28.315 3.03 ;
        RECT 28.53 11.045 28.7 11.215 ;
        RECT 28.605 2.86 28.775 3.03 ;
        RECT 29.065 2.86 29.235 3.03 ;
        RECT 29.525 2.86 29.695 3.03 ;
        RECT 29.985 2.86 30.155 3.03 ;
        RECT 31.25 11.045 31.42 11.215 ;
        RECT 31.25 1.395 31.42 1.565 ;
        RECT 31.93 11.045 32.1 11.215 ;
        RECT 31.93 1.395 32.1 1.565 ;
        RECT 32.61 11.045 32.78 11.215 ;
        RECT 32.61 1.395 32.78 1.565 ;
        RECT 33.29 11.045 33.46 11.215 ;
        RECT 33.29 1.395 33.46 1.565 ;
        RECT 33.995 11.045 34.165 11.215 ;
        RECT 33.995 1.395 34.165 1.565 ;
        RECT 34.98 1.395 35.15 1.565 ;
        RECT 34.985 11.045 35.155 11.215 ;
        RECT 36.41 2.86 36.58 3.03 ;
        RECT 36.87 2.86 37.04 3.03 ;
        RECT 37.33 2.86 37.5 3.03 ;
        RECT 37.79 2.86 37.96 3.03 ;
        RECT 38.125 4.44 38.295 4.61 ;
        RECT 38.25 2.86 38.42 3.03 ;
        RECT 38.71 2.86 38.88 3.03 ;
        RECT 39.17 2.86 39.34 3.03 ;
        RECT 39.63 2.86 39.8 3.03 ;
        RECT 39.655 3.965 39.825 4.135 ;
        RECT 40.09 2.86 40.26 3.03 ;
        RECT 40.55 2.86 40.72 3.03 ;
        RECT 41.01 2.86 41.18 3.03 ;
        RECT 41.47 2.86 41.64 3.03 ;
        RECT 41.93 2.86 42.1 3.03 ;
        RECT 42.39 2.86 42.56 3.03 ;
        RECT 42.85 2.86 43.02 3.03 ;
        RECT 43.31 2.86 43.48 3.03 ;
        RECT 43.77 2.86 43.94 3.03 ;
        RECT 44.23 2.86 44.4 3.03 ;
        RECT 44.415 11.045 44.585 11.215 ;
        RECT 44.69 2.86 44.86 3.03 ;
        RECT 45.095 11.045 45.265 11.215 ;
        RECT 45.15 2.86 45.32 3.03 ;
        RECT 45.35 8.755 45.52 8.925 ;
        RECT 45.61 2.86 45.78 3.03 ;
        RECT 45.775 11.045 45.945 11.215 ;
        RECT 46.07 2.86 46.24 3.03 ;
        RECT 46.455 11.045 46.625 11.215 ;
        RECT 46.53 2.86 46.7 3.03 ;
        RECT 46.99 2.86 47.16 3.03 ;
        RECT 47.45 2.86 47.62 3.03 ;
        RECT 47.91 2.86 48.08 3.03 ;
        RECT 49.175 11.045 49.345 11.215 ;
        RECT 49.175 1.395 49.345 1.565 ;
        RECT 49.855 11.045 50.025 11.215 ;
        RECT 49.855 1.395 50.025 1.565 ;
        RECT 50.535 11.045 50.705 11.215 ;
        RECT 50.535 1.395 50.705 1.565 ;
        RECT 51.215 11.045 51.385 11.215 ;
        RECT 51.215 1.395 51.385 1.565 ;
        RECT 51.92 11.045 52.09 11.215 ;
        RECT 51.92 1.395 52.09 1.565 ;
        RECT 52.905 1.395 53.075 1.565 ;
        RECT 52.91 11.045 53.08 11.215 ;
        RECT 54.335 2.86 54.505 3.03 ;
        RECT 54.795 2.86 54.965 3.03 ;
        RECT 55.255 2.86 55.425 3.03 ;
        RECT 55.715 2.86 55.885 3.03 ;
        RECT 56.05 4.44 56.22 4.61 ;
        RECT 56.175 2.86 56.345 3.03 ;
        RECT 56.635 2.86 56.805 3.03 ;
        RECT 57.095 2.86 57.265 3.03 ;
        RECT 57.555 2.86 57.725 3.03 ;
        RECT 57.58 3.965 57.75 4.135 ;
        RECT 58.015 2.86 58.185 3.03 ;
        RECT 58.475 2.86 58.645 3.03 ;
        RECT 58.935 2.86 59.105 3.03 ;
        RECT 59.395 2.86 59.565 3.03 ;
        RECT 59.855 2.86 60.025 3.03 ;
        RECT 60.315 2.86 60.485 3.03 ;
        RECT 60.775 2.86 60.945 3.03 ;
        RECT 61.235 2.86 61.405 3.03 ;
        RECT 61.695 2.86 61.865 3.03 ;
        RECT 62.155 2.86 62.325 3.03 ;
        RECT 62.34 11.045 62.51 11.215 ;
        RECT 62.615 2.86 62.785 3.03 ;
        RECT 63.02 11.045 63.19 11.215 ;
        RECT 63.075 2.86 63.245 3.03 ;
        RECT 63.275 8.755 63.445 8.925 ;
        RECT 63.535 2.86 63.705 3.03 ;
        RECT 63.7 11.045 63.87 11.215 ;
        RECT 63.995 2.86 64.165 3.03 ;
        RECT 64.38 11.045 64.55 11.215 ;
        RECT 64.455 2.86 64.625 3.03 ;
        RECT 64.915 2.86 65.085 3.03 ;
        RECT 65.375 2.86 65.545 3.03 ;
        RECT 65.835 2.86 66.005 3.03 ;
        RECT 67.1 11.045 67.27 11.215 ;
        RECT 67.1 1.395 67.27 1.565 ;
        RECT 67.78 11.045 67.95 11.215 ;
        RECT 67.78 1.395 67.95 1.565 ;
        RECT 68.46 11.045 68.63 11.215 ;
        RECT 68.46 1.395 68.63 1.565 ;
        RECT 69.14 11.045 69.31 11.215 ;
        RECT 69.14 1.395 69.31 1.565 ;
        RECT 69.845 11.045 70.015 11.215 ;
        RECT 69.845 1.395 70.015 1.565 ;
        RECT 70.83 1.395 71 1.565 ;
        RECT 70.835 11.045 71.005 11.215 ;
        RECT 72.26 2.86 72.43 3.03 ;
        RECT 72.72 2.86 72.89 3.03 ;
        RECT 73.18 2.86 73.35 3.03 ;
        RECT 73.64 2.86 73.81 3.03 ;
        RECT 73.975 4.44 74.145 4.61 ;
        RECT 74.1 2.86 74.27 3.03 ;
        RECT 74.56 2.86 74.73 3.03 ;
        RECT 75.02 2.86 75.19 3.03 ;
        RECT 75.48 2.86 75.65 3.03 ;
        RECT 75.505 3.965 75.675 4.135 ;
        RECT 75.94 2.86 76.11 3.03 ;
        RECT 76.4 2.86 76.57 3.03 ;
        RECT 76.86 2.86 77.03 3.03 ;
        RECT 77.32 2.86 77.49 3.03 ;
        RECT 77.78 2.86 77.95 3.03 ;
        RECT 78.24 2.86 78.41 3.03 ;
        RECT 78.7 2.86 78.87 3.03 ;
        RECT 79.16 2.86 79.33 3.03 ;
        RECT 79.62 2.86 79.79 3.03 ;
        RECT 80.08 2.86 80.25 3.03 ;
        RECT 80.265 11.045 80.435 11.215 ;
        RECT 80.54 2.86 80.71 3.03 ;
        RECT 80.945 11.045 81.115 11.215 ;
        RECT 81 2.86 81.17 3.03 ;
        RECT 81.2 8.755 81.37 8.925 ;
        RECT 81.46 2.86 81.63 3.03 ;
        RECT 81.625 11.045 81.795 11.215 ;
        RECT 81.92 2.86 82.09 3.03 ;
        RECT 82.305 11.045 82.475 11.215 ;
        RECT 82.38 2.86 82.55 3.03 ;
        RECT 82.84 2.86 83.01 3.03 ;
        RECT 83.3 2.86 83.47 3.03 ;
        RECT 83.76 2.86 83.93 3.03 ;
        RECT 85.025 11.045 85.195 11.215 ;
        RECT 85.025 1.395 85.195 1.565 ;
        RECT 85.705 11.045 85.875 11.215 ;
        RECT 85.705 1.395 85.875 1.565 ;
        RECT 86.385 11.045 86.555 11.215 ;
        RECT 86.385 1.395 86.555 1.565 ;
        RECT 87.065 11.045 87.235 11.215 ;
        RECT 87.065 1.395 87.235 1.565 ;
        RECT 87.77 11.045 87.94 11.215 ;
        RECT 87.77 1.395 87.94 1.565 ;
        RECT 88.755 1.395 88.925 1.565 ;
        RECT 88.76 11.045 88.93 11.215 ;
        RECT 90.185 2.86 90.355 3.03 ;
        RECT 90.645 2.86 90.815 3.03 ;
        RECT 91.105 2.86 91.275 3.03 ;
        RECT 91.565 2.86 91.735 3.03 ;
        RECT 91.9 4.44 92.07 4.61 ;
        RECT 92.025 2.86 92.195 3.03 ;
        RECT 92.485 2.86 92.655 3.03 ;
        RECT 92.945 2.86 93.115 3.03 ;
        RECT 93.405 2.86 93.575 3.03 ;
        RECT 93.43 3.965 93.6 4.135 ;
        RECT 93.865 2.86 94.035 3.03 ;
        RECT 94.325 2.86 94.495 3.03 ;
        RECT 94.785 2.86 94.955 3.03 ;
        RECT 95.245 2.86 95.415 3.03 ;
        RECT 95.705 2.86 95.875 3.03 ;
        RECT 96.165 2.86 96.335 3.03 ;
        RECT 96.625 2.86 96.795 3.03 ;
        RECT 97.085 2.86 97.255 3.03 ;
        RECT 97.545 2.86 97.715 3.03 ;
        RECT 98.005 2.86 98.175 3.03 ;
        RECT 98.19 11.045 98.36 11.215 ;
        RECT 98.465 2.86 98.635 3.03 ;
        RECT 98.87 11.045 99.04 11.215 ;
        RECT 98.925 2.86 99.095 3.03 ;
        RECT 99.125 8.755 99.295 8.925 ;
        RECT 99.385 2.86 99.555 3.03 ;
        RECT 99.55 11.045 99.72 11.215 ;
        RECT 99.845 2.86 100.015 3.03 ;
        RECT 100.23 11.045 100.4 11.215 ;
        RECT 100.305 2.86 100.475 3.03 ;
        RECT 100.765 2.86 100.935 3.03 ;
        RECT 101.225 2.86 101.395 3.03 ;
        RECT 101.685 2.86 101.855 3.03 ;
        RECT 102.95 11.045 103.12 11.215 ;
        RECT 102.95 1.395 103.12 1.565 ;
        RECT 103.63 11.045 103.8 11.215 ;
        RECT 103.63 1.395 103.8 1.565 ;
        RECT 104.31 11.045 104.48 11.215 ;
        RECT 104.31 1.395 104.48 1.565 ;
        RECT 104.99 11.045 105.16 11.215 ;
        RECT 104.99 1.395 105.16 1.565 ;
        RECT 105.695 11.045 105.865 11.215 ;
        RECT 105.695 1.395 105.865 1.565 ;
        RECT 106.68 1.395 106.85 1.565 ;
        RECT 106.685 11.045 106.855 11.215 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 99.385 9.49 99.76 9.86 ;
      RECT 99.42 7.36 99.73 9.86 ;
      RECT 99.42 7.36 102.515 7.67 ;
      RECT 102.205 2.805 102.515 7.67 ;
      RECT 102.215 2.435 102.59 2.805 ;
      RECT 102.215 2.42 102.525 2.805 ;
      RECT 99.345 4.98 99.9 5.31 ;
      RECT 99.345 3.315 99.645 5.31 ;
      RECT 95.41 4.42 95.965 4.75 ;
      RECT 95.665 3.315 95.965 4.75 ;
      RECT 96.46 3.18 96.61 3.83 ;
      RECT 95.665 3.315 99.645 3.615 ;
      RECT 94.17 2.255 94.47 5.205 ;
      RECT 94.17 3.86 94.9 4.19 ;
      RECT 94.125 2.255 94.5 2.625 ;
      RECT 92.73 4.42 93.46 4.75 ;
      RECT 92.735 2.255 93.035 4.75 ;
      RECT 90.62 3.86 91.35 4.19 ;
      RECT 90.765 2.225 91.065 4.19 ;
      RECT 92.69 2.255 93.065 2.625 ;
      RECT 90.72 2.225 91.095 2.595 ;
      RECT 90.72 2.265 93.065 2.565 ;
      RECT 81.46 9.49 81.835 9.86 ;
      RECT 81.495 7.36 81.805 9.86 ;
      RECT 81.495 7.36 84.59 7.67 ;
      RECT 84.28 2.805 84.59 7.67 ;
      RECT 84.29 2.435 84.665 2.805 ;
      RECT 84.29 2.42 84.6 2.805 ;
      RECT 81.42 4.98 81.975 5.31 ;
      RECT 81.42 3.315 81.72 5.31 ;
      RECT 77.485 4.42 78.04 4.75 ;
      RECT 77.74 3.315 78.04 4.75 ;
      RECT 78.535 3.18 78.685 3.83 ;
      RECT 77.74 3.315 81.72 3.615 ;
      RECT 76.245 2.255 76.545 5.205 ;
      RECT 76.245 3.86 76.975 4.19 ;
      RECT 76.2 2.255 76.575 2.625 ;
      RECT 74.805 4.42 75.535 4.75 ;
      RECT 74.81 2.255 75.11 4.75 ;
      RECT 72.695 3.86 73.425 4.19 ;
      RECT 72.84 2.225 73.14 4.19 ;
      RECT 74.765 2.255 75.14 2.625 ;
      RECT 72.795 2.225 73.17 2.595 ;
      RECT 72.795 2.265 75.14 2.565 ;
      RECT 63.535 9.49 63.91 9.86 ;
      RECT 63.57 7.36 63.88 9.86 ;
      RECT 63.57 7.36 66.665 7.67 ;
      RECT 66.355 2.805 66.665 7.67 ;
      RECT 66.365 2.435 66.74 2.805 ;
      RECT 66.365 2.42 66.675 2.805 ;
      RECT 63.495 4.98 64.05 5.31 ;
      RECT 63.495 3.315 63.795 5.31 ;
      RECT 59.56 4.42 60.115 4.75 ;
      RECT 59.815 3.315 60.115 4.75 ;
      RECT 60.61 3.18 60.76 3.83 ;
      RECT 59.815 3.315 63.795 3.615 ;
      RECT 58.32 2.255 58.62 5.205 ;
      RECT 58.32 3.86 59.05 4.19 ;
      RECT 58.275 2.255 58.65 2.625 ;
      RECT 56.88 4.42 57.61 4.75 ;
      RECT 56.885 2.255 57.185 4.75 ;
      RECT 54.77 3.86 55.5 4.19 ;
      RECT 54.915 2.225 55.215 4.19 ;
      RECT 56.84 2.255 57.215 2.625 ;
      RECT 54.87 2.225 55.245 2.595 ;
      RECT 54.87 2.265 57.215 2.565 ;
      RECT 45.61 9.49 45.985 9.86 ;
      RECT 45.645 7.36 45.955 9.86 ;
      RECT 45.645 7.36 48.74 7.67 ;
      RECT 48.43 2.805 48.74 7.67 ;
      RECT 48.44 2.435 48.815 2.805 ;
      RECT 48.44 2.42 48.75 2.805 ;
      RECT 45.57 4.98 46.125 5.31 ;
      RECT 45.57 3.315 45.87 5.31 ;
      RECT 41.635 4.42 42.19 4.75 ;
      RECT 41.89 3.315 42.19 4.75 ;
      RECT 42.685 3.18 42.835 3.83 ;
      RECT 41.89 3.315 45.87 3.615 ;
      RECT 40.395 2.255 40.695 5.205 ;
      RECT 40.395 3.86 41.125 4.19 ;
      RECT 40.35 2.255 40.725 2.625 ;
      RECT 38.955 4.42 39.685 4.75 ;
      RECT 38.96 2.255 39.26 4.75 ;
      RECT 36.845 3.86 37.575 4.19 ;
      RECT 36.99 2.225 37.29 4.19 ;
      RECT 38.915 2.255 39.29 2.625 ;
      RECT 36.945 2.225 37.32 2.595 ;
      RECT 36.945 2.265 39.29 2.565 ;
      RECT 27.685 9.49 28.06 9.86 ;
      RECT 27.72 7.36 28.03 9.86 ;
      RECT 27.72 7.36 30.815 7.67 ;
      RECT 30.505 2.805 30.815 7.67 ;
      RECT 30.515 2.435 30.89 2.805 ;
      RECT 30.515 2.42 30.825 2.805 ;
      RECT 27.645 4.98 28.2 5.31 ;
      RECT 27.645 3.315 27.945 5.31 ;
      RECT 23.71 4.42 24.265 4.75 ;
      RECT 23.965 3.315 24.265 4.75 ;
      RECT 24.76 3.18 24.91 3.83 ;
      RECT 23.965 3.315 27.945 3.615 ;
      RECT 22.47 2.255 22.77 5.205 ;
      RECT 22.47 3.86 23.2 4.19 ;
      RECT 22.425 2.255 22.8 2.625 ;
      RECT 21.03 4.42 21.76 4.75 ;
      RECT 21.035 2.255 21.335 4.75 ;
      RECT 18.92 3.86 19.65 4.19 ;
      RECT 19.065 2.225 19.365 4.19 ;
      RECT 20.99 2.255 21.365 2.625 ;
      RECT 19.02 2.225 19.395 2.595 ;
      RECT 19.02 2.265 21.365 2.565 ;
      RECT 106.94 7.35 107.315 12.61 ;
      RECT 100.53 3.3 101.26 3.63 ;
      RECT 98.31 4.98 99.04 5.31 ;
      RECT 96.61 4.98 97.34 5.31 ;
      RECT 90.29 4.98 91.02 5.31 ;
      RECT 89.015 7.35 89.39 12.61 ;
      RECT 82.605 3.3 83.335 3.63 ;
      RECT 80.385 4.98 81.115 5.31 ;
      RECT 78.685 4.98 79.415 5.31 ;
      RECT 72.365 4.98 73.095 5.31 ;
      RECT 71.09 7.35 71.465 12.61 ;
      RECT 64.68 3.3 65.41 3.63 ;
      RECT 62.46 4.98 63.19 5.31 ;
      RECT 60.76 4.98 61.49 5.31 ;
      RECT 54.44 4.98 55.17 5.31 ;
      RECT 53.165 7.35 53.54 12.61 ;
      RECT 46.755 3.3 47.485 3.63 ;
      RECT 44.535 4.98 45.265 5.31 ;
      RECT 42.835 4.98 43.565 5.31 ;
      RECT 36.515 4.98 37.245 5.31 ;
      RECT 35.24 7.35 35.615 12.61 ;
      RECT 28.83 3.3 29.56 3.63 ;
      RECT 26.61 4.98 27.34 5.31 ;
      RECT 24.91 4.98 25.64 5.31 ;
      RECT 18.59 4.98 19.32 5.31 ;
    LAYER via2 ;
      RECT 107.025 7.44 107.225 7.64 ;
      RECT 102.305 2.52 102.505 2.72 ;
      RECT 100.595 3.365 100.795 3.565 ;
      RECT 99.635 5.045 99.835 5.245 ;
      RECT 99.475 9.575 99.675 9.775 ;
      RECT 98.635 5.045 98.835 5.245 ;
      RECT 96.675 5.045 96.875 5.245 ;
      RECT 95.475 4.485 95.675 4.685 ;
      RECT 94.235 3.925 94.435 4.125 ;
      RECT 94.215 2.34 94.415 2.54 ;
      RECT 92.795 4.485 92.995 4.685 ;
      RECT 92.78 2.335 92.98 2.535 ;
      RECT 90.835 3.925 91.035 4.125 ;
      RECT 90.81 2.31 91.01 2.51 ;
      RECT 90.355 5.045 90.555 5.245 ;
      RECT 89.1 7.44 89.3 7.64 ;
      RECT 84.38 2.52 84.58 2.72 ;
      RECT 82.67 3.365 82.87 3.565 ;
      RECT 81.71 5.045 81.91 5.245 ;
      RECT 81.55 9.575 81.75 9.775 ;
      RECT 80.71 5.045 80.91 5.245 ;
      RECT 78.75 5.045 78.95 5.245 ;
      RECT 77.55 4.485 77.75 4.685 ;
      RECT 76.31 3.925 76.51 4.125 ;
      RECT 76.29 2.34 76.49 2.54 ;
      RECT 74.87 4.485 75.07 4.685 ;
      RECT 74.855 2.335 75.055 2.535 ;
      RECT 72.91 3.925 73.11 4.125 ;
      RECT 72.885 2.31 73.085 2.51 ;
      RECT 72.43 5.045 72.63 5.245 ;
      RECT 71.175 7.44 71.375 7.64 ;
      RECT 66.455 2.52 66.655 2.72 ;
      RECT 64.745 3.365 64.945 3.565 ;
      RECT 63.785 5.045 63.985 5.245 ;
      RECT 63.625 9.575 63.825 9.775 ;
      RECT 62.785 5.045 62.985 5.245 ;
      RECT 60.825 5.045 61.025 5.245 ;
      RECT 59.625 4.485 59.825 4.685 ;
      RECT 58.385 3.925 58.585 4.125 ;
      RECT 58.365 2.34 58.565 2.54 ;
      RECT 56.945 4.485 57.145 4.685 ;
      RECT 56.93 2.335 57.13 2.535 ;
      RECT 54.985 3.925 55.185 4.125 ;
      RECT 54.96 2.31 55.16 2.51 ;
      RECT 54.505 5.045 54.705 5.245 ;
      RECT 53.25 7.44 53.45 7.64 ;
      RECT 48.53 2.52 48.73 2.72 ;
      RECT 46.82 3.365 47.02 3.565 ;
      RECT 45.86 5.045 46.06 5.245 ;
      RECT 45.7 9.575 45.9 9.775 ;
      RECT 44.86 5.045 45.06 5.245 ;
      RECT 42.9 5.045 43.1 5.245 ;
      RECT 41.7 4.485 41.9 4.685 ;
      RECT 40.46 3.925 40.66 4.125 ;
      RECT 40.44 2.34 40.64 2.54 ;
      RECT 39.02 4.485 39.22 4.685 ;
      RECT 39.005 2.335 39.205 2.535 ;
      RECT 37.06 3.925 37.26 4.125 ;
      RECT 37.035 2.31 37.235 2.51 ;
      RECT 36.58 5.045 36.78 5.245 ;
      RECT 35.325 7.44 35.525 7.64 ;
      RECT 30.605 2.52 30.805 2.72 ;
      RECT 28.895 3.365 29.095 3.565 ;
      RECT 27.935 5.045 28.135 5.245 ;
      RECT 27.775 9.575 27.975 9.775 ;
      RECT 26.935 5.045 27.135 5.245 ;
      RECT 24.975 5.045 25.175 5.245 ;
      RECT 23.775 4.485 23.975 4.685 ;
      RECT 22.535 3.925 22.735 4.125 ;
      RECT 22.515 2.34 22.715 2.54 ;
      RECT 21.095 4.485 21.295 4.685 ;
      RECT 21.08 2.335 21.28 2.535 ;
      RECT 19.135 3.925 19.335 4.125 ;
      RECT 19.11 2.31 19.31 2.51 ;
      RECT 18.655 5.045 18.855 5.245 ;
    LAYER met2 ;
      RECT 16.39 10.835 107.205 11.005 ;
      RECT 107.035 9.71 107.205 11.005 ;
      RECT 16.39 8.69 16.56 11.005 ;
      RECT 107.005 9.71 107.355 10.06 ;
      RECT 16.33 8.69 16.62 9.04 ;
      RECT 103.85 8.66 104.17 8.98 ;
      RECT 103.88 8.13 104.05 8.98 ;
      RECT 103.88 8.13 104.055 8.48 ;
      RECT 103.88 8.13 104.855 8.305 ;
      RECT 104.68 3.26 104.855 8.305 ;
      RECT 104.625 3.26 104.975 3.61 ;
      RECT 104.65 9.09 104.975 9.415 ;
      RECT 103.535 9.18 104.975 9.35 ;
      RECT 103.535 3.69 103.695 9.35 ;
      RECT 103.85 3.66 104.17 3.98 ;
      RECT 103.535 3.69 104.17 3.86 ;
      RECT 102.215 2.435 102.59 2.805 ;
      RECT 94.125 2.255 94.5 2.625 ;
      RECT 92.69 2.255 93.065 2.625 ;
      RECT 92.69 2.375 102.52 2.545 ;
      RECT 96.81 5.655 102.49 5.825 ;
      RECT 102.32 4.72 102.49 5.825 ;
      RECT 96.62 4.895 96.655 5.825 ;
      RECT 96.885 5.005 96.915 5.285 ;
      RECT 96.59 4.895 96.655 5.155 ;
      RECT 102.23 4.725 102.58 5.075 ;
      RECT 96.42 3.52 96.455 3.78 ;
      RECT 96.195 3.52 96.255 3.78 ;
      RECT 96.875 4.985 96.885 5.285 ;
      RECT 96.87 4.945 96.875 5.285 ;
      RECT 96.855 4.9 96.87 5.285 ;
      RECT 96.85 4.865 96.855 5.285 ;
      RECT 96.845 4.845 96.85 5.285 ;
      RECT 96.815 4.772 96.845 5.285 ;
      RECT 96.81 4.7 96.815 5.285 ;
      RECT 96.795 4.66 96.81 5.825 ;
      RECT 96.785 4.6 96.795 5.825 ;
      RECT 96.74 4.54 96.785 5.825 ;
      RECT 96.655 4.501 96.74 5.825 ;
      RECT 96.65 4.492 96.655 4.865 ;
      RECT 96.64 4.491 96.65 4.848 ;
      RECT 96.615 4.472 96.64 4.818 ;
      RECT 96.61 4.447 96.615 4.797 ;
      RECT 96.6 4.425 96.61 4.788 ;
      RECT 96.595 4.396 96.6 4.778 ;
      RECT 96.555 4.322 96.595 4.75 ;
      RECT 96.535 4.223 96.555 4.715 ;
      RECT 96.52 4.159 96.535 4.698 ;
      RECT 96.49 4.083 96.52 4.67 ;
      RECT 96.47 3.998 96.49 4.643 ;
      RECT 96.43 3.894 96.47 4.55 ;
      RECT 96.425 3.815 96.43 4.458 ;
      RECT 96.42 3.798 96.425 4.435 ;
      RECT 96.415 3.52 96.42 4.415 ;
      RECT 96.385 3.52 96.415 4.353 ;
      RECT 96.38 3.52 96.385 4.285 ;
      RECT 96.37 3.52 96.38 4.25 ;
      RECT 96.36 3.52 96.37 4.215 ;
      RECT 96.295 3.52 96.36 4.07 ;
      RECT 96.29 3.52 96.295 3.94 ;
      RECT 96.26 3.52 96.29 3.873 ;
      RECT 96.255 3.52 96.26 3.798 ;
      RECT 100.59 3.455 100.85 3.715 ;
      RECT 100.585 3.455 100.85 3.663 ;
      RECT 100.58 3.455 100.85 3.633 ;
      RECT 100.555 3.325 100.835 3.605 ;
      RECT 89.06 9.095 89.41 9.445 ;
      RECT 100.305 9.05 100.655 9.4 ;
      RECT 89.06 9.125 100.655 9.325 ;
      RECT 99.595 5.005 99.875 5.285 ;
      RECT 99.635 4.96 99.9 5.22 ;
      RECT 99.625 4.995 99.9 5.22 ;
      RECT 99.63 4.98 99.875 5.285 ;
      RECT 99.635 4.957 99.845 5.285 ;
      RECT 99.635 4.955 99.83 5.285 ;
      RECT 99.675 4.945 99.83 5.285 ;
      RECT 99.645 4.95 99.83 5.285 ;
      RECT 99.675 4.942 99.775 5.285 ;
      RECT 99.7 4.935 99.775 5.285 ;
      RECT 99.68 4.937 99.775 5.285 ;
      RECT 99.01 4.45 99.27 4.71 ;
      RECT 99.06 4.442 99.25 4.71 ;
      RECT 99.065 4.362 99.25 4.71 ;
      RECT 99.185 3.75 99.25 4.71 ;
      RECT 99.09 4.147 99.25 4.71 ;
      RECT 99.165 3.835 99.25 4.71 ;
      RECT 99.2 3.46 99.336 4.188 ;
      RECT 99.145 3.957 99.336 4.188 ;
      RECT 99.16 3.897 99.25 4.71 ;
      RECT 99.2 3.46 99.36 3.853 ;
      RECT 99.2 3.46 99.37 3.75 ;
      RECT 99.19 3.46 99.45 3.72 ;
      RECT 98.595 5.005 98.875 5.285 ;
      RECT 98.615 4.965 98.875 5.285 ;
      RECT 98.255 4.92 98.36 5.18 ;
      RECT 98.11 3.41 98.2 3.67 ;
      RECT 98.65 4.475 98.655 4.515 ;
      RECT 98.645 4.465 98.65 4.6 ;
      RECT 98.64 4.455 98.645 4.693 ;
      RECT 98.63 4.435 98.64 4.749 ;
      RECT 98.55 4.363 98.63 4.829 ;
      RECT 98.585 5.007 98.595 5.232 ;
      RECT 98.58 5.004 98.585 5.227 ;
      RECT 98.565 5.001 98.58 5.22 ;
      RECT 98.53 4.995 98.565 5.202 ;
      RECT 98.545 4.298 98.55 4.903 ;
      RECT 98.525 4.249 98.545 4.918 ;
      RECT 98.515 4.982 98.53 5.185 ;
      RECT 98.52 4.191 98.525 4.933 ;
      RECT 98.515 4.169 98.52 4.943 ;
      RECT 98.48 4.079 98.515 5.18 ;
      RECT 98.465 3.957 98.48 5.18 ;
      RECT 98.46 3.91 98.465 5.18 ;
      RECT 98.435 3.835 98.46 5.18 ;
      RECT 98.42 3.75 98.435 5.18 ;
      RECT 98.415 3.697 98.42 5.18 ;
      RECT 98.41 3.677 98.415 5.18 ;
      RECT 98.405 3.652 98.41 4.414 ;
      RECT 98.39 4.612 98.41 5.18 ;
      RECT 98.4 3.63 98.405 4.391 ;
      RECT 98.39 3.582 98.4 4.356 ;
      RECT 98.385 3.545 98.39 4.322 ;
      RECT 98.385 4.692 98.39 5.18 ;
      RECT 98.37 3.522 98.385 4.277 ;
      RECT 98.365 4.79 98.385 5.18 ;
      RECT 98.315 3.41 98.37 4.119 ;
      RECT 98.36 4.912 98.365 5.18 ;
      RECT 98.3 3.41 98.315 3.958 ;
      RECT 98.295 3.41 98.3 3.91 ;
      RECT 98.29 3.41 98.295 3.898 ;
      RECT 98.245 3.41 98.29 3.835 ;
      RECT 98.22 3.41 98.245 3.753 ;
      RECT 98.205 3.41 98.22 3.705 ;
      RECT 98.2 3.41 98.205 3.675 ;
      RECT 97.525 4.86 97.57 5.12 ;
      RECT 97.43 3.395 97.575 3.655 ;
      RECT 97.935 4.017 97.945 4.108 ;
      RECT 97.92 3.955 97.935 4.164 ;
      RECT 97.915 3.902 97.92 4.21 ;
      RECT 97.865 3.849 97.915 4.336 ;
      RECT 97.86 3.804 97.865 4.483 ;
      RECT 97.85 3.792 97.86 4.525 ;
      RECT 97.815 3.756 97.85 4.63 ;
      RECT 97.81 3.724 97.815 4.736 ;
      RECT 97.795 3.706 97.81 4.781 ;
      RECT 97.79 3.689 97.795 4.015 ;
      RECT 97.785 4.07 97.795 4.838 ;
      RECT 97.78 3.675 97.79 3.988 ;
      RECT 97.775 4.125 97.785 5.12 ;
      RECT 97.77 3.661 97.78 3.973 ;
      RECT 97.77 4.175 97.775 5.12 ;
      RECT 97.755 3.638 97.77 3.953 ;
      RECT 97.735 4.297 97.77 5.12 ;
      RECT 97.75 3.62 97.755 3.935 ;
      RECT 97.745 3.612 97.75 3.925 ;
      RECT 97.715 3.58 97.745 3.889 ;
      RECT 97.725 4.425 97.735 5.12 ;
      RECT 97.72 4.452 97.725 5.12 ;
      RECT 97.715 4.502 97.72 5.12 ;
      RECT 97.705 3.546 97.715 3.854 ;
      RECT 97.665 4.57 97.715 5.12 ;
      RECT 97.69 3.523 97.705 3.83 ;
      RECT 97.665 3.395 97.69 3.793 ;
      RECT 97.66 3.395 97.665 3.765 ;
      RECT 97.63 4.67 97.665 5.12 ;
      RECT 97.655 3.395 97.66 3.758 ;
      RECT 97.65 3.395 97.655 3.748 ;
      RECT 97.635 3.395 97.65 3.733 ;
      RECT 97.62 3.395 97.635 3.705 ;
      RECT 97.585 4.775 97.63 5.12 ;
      RECT 97.605 3.395 97.62 3.678 ;
      RECT 97.575 3.395 97.605 3.663 ;
      RECT 97.57 4.847 97.585 5.12 ;
      RECT 97.495 3.93 97.535 4.19 ;
      RECT 97.27 3.877 97.275 4.135 ;
      RECT 93.225 3.355 93.485 3.615 ;
      RECT 93.225 3.38 93.5 3.595 ;
      RECT 95.615 3.205 95.62 3.35 ;
      RECT 97.485 3.925 97.495 4.19 ;
      RECT 97.465 3.917 97.485 4.19 ;
      RECT 97.447 3.913 97.465 4.19 ;
      RECT 97.361 3.902 97.447 4.19 ;
      RECT 97.275 3.885 97.361 4.19 ;
      RECT 97.22 3.872 97.27 4.12 ;
      RECT 97.186 3.864 97.22 4.095 ;
      RECT 97.1 3.853 97.186 4.06 ;
      RECT 97.065 3.83 97.1 4.025 ;
      RECT 97.055 3.792 97.065 4.011 ;
      RECT 97.05 3.765 97.055 4.007 ;
      RECT 97.045 3.752 97.05 4.004 ;
      RECT 97.035 3.732 97.045 4 ;
      RECT 97.03 3.707 97.035 3.996 ;
      RECT 97.005 3.662 97.03 3.99 ;
      RECT 96.995 3.603 97.005 3.982 ;
      RECT 96.985 3.571 96.995 3.973 ;
      RECT 96.965 3.523 96.985 3.953 ;
      RECT 96.96 3.483 96.965 3.923 ;
      RECT 96.945 3.457 96.96 3.897 ;
      RECT 96.94 3.435 96.945 3.873 ;
      RECT 96.925 3.407 96.94 3.849 ;
      RECT 96.91 3.38 96.925 3.813 ;
      RECT 96.895 3.357 96.91 3.775 ;
      RECT 96.89 3.347 96.895 3.75 ;
      RECT 96.88 3.34 96.89 3.733 ;
      RECT 96.865 3.327 96.88 3.703 ;
      RECT 96.86 3.317 96.865 3.678 ;
      RECT 96.855 3.312 96.86 3.665 ;
      RECT 96.845 3.305 96.855 3.645 ;
      RECT 96.84 3.298 96.845 3.63 ;
      RECT 96.815 3.291 96.84 3.588 ;
      RECT 96.8 3.281 96.815 3.538 ;
      RECT 96.79 3.276 96.8 3.508 ;
      RECT 96.78 3.272 96.79 3.483 ;
      RECT 96.765 3.269 96.78 3.473 ;
      RECT 96.715 3.266 96.765 3.458 ;
      RECT 96.695 3.264 96.715 3.443 ;
      RECT 96.646 3.262 96.695 3.438 ;
      RECT 96.56 3.258 96.646 3.433 ;
      RECT 96.521 3.255 96.56 3.429 ;
      RECT 96.435 3.251 96.521 3.424 ;
      RECT 96.385 3.248 96.435 3.418 ;
      RECT 96.336 3.245 96.385 3.413 ;
      RECT 96.25 3.242 96.336 3.408 ;
      RECT 96.246 3.24 96.25 3.405 ;
      RECT 96.16 3.237 96.246 3.4 ;
      RECT 96.111 3.233 96.16 3.393 ;
      RECT 96.025 3.23 96.111 3.388 ;
      RECT 96.001 3.227 96.025 3.384 ;
      RECT 95.915 3.225 96.001 3.379 ;
      RECT 95.85 3.221 95.915 3.372 ;
      RECT 95.847 3.22 95.85 3.369 ;
      RECT 95.761 3.217 95.847 3.366 ;
      RECT 95.675 3.211 95.761 3.359 ;
      RECT 95.645 3.207 95.675 3.355 ;
      RECT 95.62 3.205 95.645 3.353 ;
      RECT 95.565 3.202 95.615 3.35 ;
      RECT 95.485 3.201 95.565 3.35 ;
      RECT 95.43 3.203 95.485 3.353 ;
      RECT 95.415 3.204 95.43 3.357 ;
      RECT 95.36 3.212 95.415 3.367 ;
      RECT 95.33 3.22 95.36 3.38 ;
      RECT 95.311 3.221 95.33 3.386 ;
      RECT 95.225 3.224 95.311 3.391 ;
      RECT 95.155 3.229 95.225 3.4 ;
      RECT 95.136 3.232 95.155 3.406 ;
      RECT 95.05 3.236 95.136 3.411 ;
      RECT 95.01 3.24 95.05 3.418 ;
      RECT 95.001 3.242 95.01 3.421 ;
      RECT 94.915 3.246 95.001 3.426 ;
      RECT 94.912 3.249 94.915 3.43 ;
      RECT 94.826 3.252 94.912 3.434 ;
      RECT 94.74 3.258 94.826 3.442 ;
      RECT 94.716 3.262 94.74 3.446 ;
      RECT 94.63 3.266 94.716 3.451 ;
      RECT 94.585 3.271 94.63 3.458 ;
      RECT 94.505 3.276 94.585 3.465 ;
      RECT 94.425 3.282 94.505 3.48 ;
      RECT 94.4 3.286 94.425 3.493 ;
      RECT 94.335 3.289 94.4 3.505 ;
      RECT 94.28 3.294 94.335 3.52 ;
      RECT 94.25 3.297 94.28 3.538 ;
      RECT 94.24 3.299 94.25 3.551 ;
      RECT 94.18 3.314 94.24 3.561 ;
      RECT 94.165 3.331 94.18 3.57 ;
      RECT 94.16 3.34 94.165 3.57 ;
      RECT 94.15 3.35 94.16 3.57 ;
      RECT 94.14 3.367 94.15 3.57 ;
      RECT 94.12 3.377 94.14 3.571 ;
      RECT 94.075 3.387 94.12 3.572 ;
      RECT 94.04 3.396 94.075 3.574 ;
      RECT 93.975 3.401 94.04 3.576 ;
      RECT 93.895 3.402 93.975 3.579 ;
      RECT 93.891 3.4 93.895 3.58 ;
      RECT 93.805 3.397 93.891 3.582 ;
      RECT 93.758 3.394 93.805 3.584 ;
      RECT 93.672 3.39 93.758 3.587 ;
      RECT 93.586 3.386 93.672 3.59 ;
      RECT 93.5 3.382 93.586 3.594 ;
      RECT 95.435 4.445 95.715 4.725 ;
      RECT 95.475 4.425 95.735 4.685 ;
      RECT 95.465 4.435 95.735 4.685 ;
      RECT 95.475 4.362 95.69 4.725 ;
      RECT 95.53 4.285 95.685 4.725 ;
      RECT 95.535 4.07 95.685 4.725 ;
      RECT 95.525 3.872 95.675 4.123 ;
      RECT 95.515 3.872 95.675 3.99 ;
      RECT 95.51 3.75 95.67 3.893 ;
      RECT 95.495 3.75 95.67 3.798 ;
      RECT 95.49 3.46 95.665 3.775 ;
      RECT 95.475 3.46 95.665 3.745 ;
      RECT 95.435 3.46 95.695 3.72 ;
      RECT 95.345 4.93 95.425 5.19 ;
      RECT 94.75 3.65 94.755 3.915 ;
      RECT 94.63 3.65 94.755 3.91 ;
      RECT 95.305 4.895 95.345 5.19 ;
      RECT 95.26 4.817 95.305 5.19 ;
      RECT 95.24 4.745 95.26 5.19 ;
      RECT 95.23 4.697 95.24 5.19 ;
      RECT 95.195 4.63 95.23 5.19 ;
      RECT 95.165 4.53 95.195 5.19 ;
      RECT 95.145 4.455 95.165 4.99 ;
      RECT 95.135 4.405 95.145 4.945 ;
      RECT 95.13 4.382 95.135 4.918 ;
      RECT 95.125 4.367 95.13 4.905 ;
      RECT 95.12 4.352 95.125 4.883 ;
      RECT 95.115 4.337 95.12 4.865 ;
      RECT 95.09 4.292 95.115 4.82 ;
      RECT 95.08 4.24 95.09 4.763 ;
      RECT 95.07 4.21 95.08 4.73 ;
      RECT 95.06 4.175 95.07 4.698 ;
      RECT 95.025 4.107 95.06 4.63 ;
      RECT 95.02 4.046 95.025 4.565 ;
      RECT 95.01 4.034 95.02 4.545 ;
      RECT 95.005 4.022 95.01 4.525 ;
      RECT 95 4.014 95.005 4.513 ;
      RECT 94.995 4.006 95 4.493 ;
      RECT 94.985 3.994 94.995 4.465 ;
      RECT 94.975 3.978 94.985 4.435 ;
      RECT 94.95 3.95 94.975 4.373 ;
      RECT 94.94 3.921 94.95 4.318 ;
      RECT 94.925 3.9 94.94 4.278 ;
      RECT 94.92 3.884 94.925 4.25 ;
      RECT 94.915 3.872 94.92 4.24 ;
      RECT 94.91 3.867 94.915 4.213 ;
      RECT 94.905 3.86 94.91 4.2 ;
      RECT 94.89 3.843 94.905 4.173 ;
      RECT 94.88 3.65 94.89 4.133 ;
      RECT 94.87 3.65 94.88 4.1 ;
      RECT 94.86 3.65 94.87 4.075 ;
      RECT 94.79 3.65 94.86 4.01 ;
      RECT 94.78 3.65 94.79 3.958 ;
      RECT 94.765 3.65 94.78 3.94 ;
      RECT 94.755 3.65 94.765 3.925 ;
      RECT 94.585 4.52 94.845 4.78 ;
      RECT 93.12 4.555 93.125 4.762 ;
      RECT 92.755 4.445 92.83 4.76 ;
      RECT 92.57 4.5 92.725 4.76 ;
      RECT 92.755 4.445 92.86 4.725 ;
      RECT 94.57 4.617 94.585 4.778 ;
      RECT 94.545 4.625 94.57 4.783 ;
      RECT 94.52 4.632 94.545 4.788 ;
      RECT 94.457 4.643 94.52 4.797 ;
      RECT 94.371 4.662 94.457 4.814 ;
      RECT 94.285 4.684 94.371 4.833 ;
      RECT 94.27 4.697 94.285 4.844 ;
      RECT 94.23 4.705 94.27 4.851 ;
      RECT 94.21 4.71 94.23 4.858 ;
      RECT 94.172 4.711 94.21 4.861 ;
      RECT 94.086 4.714 94.172 4.862 ;
      RECT 94 4.718 94.086 4.863 ;
      RECT 93.951 4.72 94 4.865 ;
      RECT 93.865 4.72 93.951 4.867 ;
      RECT 93.825 4.715 93.865 4.869 ;
      RECT 93.815 4.709 93.825 4.87 ;
      RECT 93.775 4.704 93.815 4.867 ;
      RECT 93.765 4.697 93.775 4.863 ;
      RECT 93.75 4.693 93.765 4.861 ;
      RECT 93.733 4.689 93.75 4.859 ;
      RECT 93.647 4.679 93.733 4.851 ;
      RECT 93.561 4.661 93.647 4.837 ;
      RECT 93.475 4.644 93.561 4.823 ;
      RECT 93.45 4.632 93.475 4.814 ;
      RECT 93.38 4.622 93.45 4.807 ;
      RECT 93.335 4.61 93.38 4.798 ;
      RECT 93.275 4.597 93.335 4.79 ;
      RECT 93.27 4.589 93.275 4.785 ;
      RECT 93.235 4.584 93.27 4.783 ;
      RECT 93.18 4.575 93.235 4.776 ;
      RECT 93.14 4.564 93.18 4.768 ;
      RECT 93.125 4.557 93.14 4.764 ;
      RECT 93.105 4.55 93.12 4.761 ;
      RECT 93.09 4.54 93.105 4.759 ;
      RECT 93.075 4.527 93.09 4.756 ;
      RECT 93.05 4.51 93.075 4.752 ;
      RECT 93.035 4.492 93.05 4.749 ;
      RECT 93.01 4.445 93.035 4.747 ;
      RECT 92.986 4.445 93.01 4.744 ;
      RECT 92.9 4.445 92.986 4.736 ;
      RECT 92.86 4.445 92.9 4.728 ;
      RECT 92.725 4.492 92.755 4.76 ;
      RECT 94.405 4.075 94.665 4.335 ;
      RECT 94.365 4.075 94.665 4.213 ;
      RECT 94.33 4.075 94.665 4.198 ;
      RECT 94.275 4.075 94.665 4.178 ;
      RECT 94.195 3.885 94.475 4.165 ;
      RECT 94.195 4.067 94.545 4.165 ;
      RECT 94.195 4.01 94.53 4.165 ;
      RECT 94.195 3.957 94.48 4.165 ;
      RECT 91.355 4.244 91.37 4.7 ;
      RECT 91.35 4.316 91.456 4.698 ;
      RECT 91.37 3.41 91.505 4.696 ;
      RECT 91.355 4.26 91.51 4.695 ;
      RECT 91.355 4.31 91.515 4.693 ;
      RECT 91.34 4.375 91.515 4.692 ;
      RECT 91.35 4.367 91.52 4.689 ;
      RECT 91.33 4.415 91.52 4.684 ;
      RECT 91.33 4.415 91.535 4.681 ;
      RECT 91.325 4.415 91.535 4.678 ;
      RECT 91.3 4.415 91.56 4.675 ;
      RECT 91.37 3.41 91.53 4.063 ;
      RECT 91.365 3.41 91.53 4.035 ;
      RECT 91.36 3.41 91.53 3.863 ;
      RECT 91.36 3.41 91.55 3.803 ;
      RECT 91.315 3.41 91.575 3.67 ;
      RECT 90.795 3.885 91.075 4.165 ;
      RECT 90.785 3.9 91.075 4.16 ;
      RECT 90.74 3.962 91.075 4.158 ;
      RECT 90.815 3.877 90.98 4.165 ;
      RECT 90.815 3.862 90.936 4.165 ;
      RECT 90.85 3.855 90.936 4.165 ;
      RECT 90.315 5.005 90.595 5.285 ;
      RECT 90.275 4.967 90.57 5.078 ;
      RECT 90.26 4.917 90.55 4.973 ;
      RECT 90.205 4.68 90.465 4.94 ;
      RECT 90.205 4.882 90.545 4.94 ;
      RECT 90.205 4.822 90.54 4.94 ;
      RECT 90.205 4.772 90.52 4.94 ;
      RECT 90.205 4.752 90.515 4.94 ;
      RECT 90.205 4.73 90.51 4.94 ;
      RECT 90.205 4.715 90.48 4.94 ;
      RECT 85.925 8.66 86.245 8.98 ;
      RECT 85.955 8.13 86.125 8.98 ;
      RECT 85.955 8.13 86.13 8.48 ;
      RECT 85.955 8.13 86.93 8.305 ;
      RECT 86.755 3.26 86.93 8.305 ;
      RECT 86.7 3.26 87.05 3.61 ;
      RECT 86.725 9.09 87.05 9.415 ;
      RECT 85.61 9.18 87.05 9.35 ;
      RECT 85.61 3.69 85.77 9.35 ;
      RECT 85.925 3.66 86.245 3.98 ;
      RECT 85.61 3.69 86.245 3.86 ;
      RECT 84.29 2.435 84.665 2.805 ;
      RECT 76.2 2.255 76.575 2.625 ;
      RECT 74.765 2.255 75.14 2.625 ;
      RECT 74.765 2.375 84.595 2.545 ;
      RECT 78.885 5.655 84.565 5.825 ;
      RECT 84.395 4.72 84.565 5.825 ;
      RECT 78.695 4.895 78.73 5.825 ;
      RECT 78.96 5.005 78.99 5.285 ;
      RECT 78.665 4.895 78.73 5.155 ;
      RECT 84.305 4.725 84.655 5.075 ;
      RECT 78.495 3.52 78.53 3.78 ;
      RECT 78.27 3.52 78.33 3.78 ;
      RECT 78.95 4.985 78.96 5.285 ;
      RECT 78.945 4.945 78.95 5.285 ;
      RECT 78.93 4.9 78.945 5.285 ;
      RECT 78.925 4.865 78.93 5.285 ;
      RECT 78.92 4.845 78.925 5.285 ;
      RECT 78.89 4.772 78.92 5.285 ;
      RECT 78.885 4.7 78.89 5.285 ;
      RECT 78.87 4.66 78.885 5.825 ;
      RECT 78.86 4.6 78.87 5.825 ;
      RECT 78.815 4.54 78.86 5.825 ;
      RECT 78.73 4.501 78.815 5.825 ;
      RECT 78.725 4.492 78.73 4.865 ;
      RECT 78.715 4.491 78.725 4.848 ;
      RECT 78.69 4.472 78.715 4.818 ;
      RECT 78.685 4.447 78.69 4.797 ;
      RECT 78.675 4.425 78.685 4.788 ;
      RECT 78.67 4.396 78.675 4.778 ;
      RECT 78.63 4.322 78.67 4.75 ;
      RECT 78.61 4.223 78.63 4.715 ;
      RECT 78.595 4.159 78.61 4.698 ;
      RECT 78.565 4.083 78.595 4.67 ;
      RECT 78.545 3.998 78.565 4.643 ;
      RECT 78.505 3.894 78.545 4.55 ;
      RECT 78.5 3.815 78.505 4.458 ;
      RECT 78.495 3.798 78.5 4.435 ;
      RECT 78.49 3.52 78.495 4.415 ;
      RECT 78.46 3.52 78.49 4.353 ;
      RECT 78.455 3.52 78.46 4.285 ;
      RECT 78.445 3.52 78.455 4.25 ;
      RECT 78.435 3.52 78.445 4.215 ;
      RECT 78.37 3.52 78.435 4.07 ;
      RECT 78.365 3.52 78.37 3.94 ;
      RECT 78.335 3.52 78.365 3.873 ;
      RECT 78.33 3.52 78.335 3.798 ;
      RECT 82.665 3.455 82.925 3.715 ;
      RECT 82.66 3.455 82.925 3.663 ;
      RECT 82.655 3.455 82.925 3.633 ;
      RECT 82.63 3.325 82.91 3.605 ;
      RECT 71.135 9.095 71.485 9.445 ;
      RECT 82.1 9.05 82.45 9.4 ;
      RECT 71.135 9.125 82.45 9.325 ;
      RECT 81.67 5.005 81.95 5.285 ;
      RECT 81.71 4.96 81.975 5.22 ;
      RECT 81.7 4.995 81.975 5.22 ;
      RECT 81.705 4.98 81.95 5.285 ;
      RECT 81.71 4.957 81.92 5.285 ;
      RECT 81.71 4.955 81.905 5.285 ;
      RECT 81.75 4.945 81.905 5.285 ;
      RECT 81.72 4.95 81.905 5.285 ;
      RECT 81.75 4.942 81.85 5.285 ;
      RECT 81.775 4.935 81.85 5.285 ;
      RECT 81.755 4.937 81.85 5.285 ;
      RECT 81.085 4.45 81.345 4.71 ;
      RECT 81.135 4.442 81.325 4.71 ;
      RECT 81.14 4.362 81.325 4.71 ;
      RECT 81.26 3.75 81.325 4.71 ;
      RECT 81.165 4.147 81.325 4.71 ;
      RECT 81.24 3.835 81.325 4.71 ;
      RECT 81.275 3.46 81.411 4.188 ;
      RECT 81.22 3.957 81.411 4.188 ;
      RECT 81.235 3.897 81.325 4.71 ;
      RECT 81.275 3.46 81.435 3.853 ;
      RECT 81.275 3.46 81.445 3.75 ;
      RECT 81.265 3.46 81.525 3.72 ;
      RECT 80.67 5.005 80.95 5.285 ;
      RECT 80.69 4.965 80.95 5.285 ;
      RECT 80.33 4.92 80.435 5.18 ;
      RECT 80.185 3.41 80.275 3.67 ;
      RECT 80.725 4.475 80.73 4.515 ;
      RECT 80.72 4.465 80.725 4.6 ;
      RECT 80.715 4.455 80.72 4.693 ;
      RECT 80.705 4.435 80.715 4.749 ;
      RECT 80.625 4.363 80.705 4.829 ;
      RECT 80.66 5.007 80.67 5.232 ;
      RECT 80.655 5.004 80.66 5.227 ;
      RECT 80.64 5.001 80.655 5.22 ;
      RECT 80.605 4.995 80.64 5.202 ;
      RECT 80.62 4.298 80.625 4.903 ;
      RECT 80.6 4.249 80.62 4.918 ;
      RECT 80.59 4.982 80.605 5.185 ;
      RECT 80.595 4.191 80.6 4.933 ;
      RECT 80.59 4.169 80.595 4.943 ;
      RECT 80.555 4.079 80.59 5.18 ;
      RECT 80.54 3.957 80.555 5.18 ;
      RECT 80.535 3.91 80.54 5.18 ;
      RECT 80.51 3.835 80.535 5.18 ;
      RECT 80.495 3.75 80.51 5.18 ;
      RECT 80.49 3.697 80.495 5.18 ;
      RECT 80.485 3.677 80.49 5.18 ;
      RECT 80.48 3.652 80.485 4.414 ;
      RECT 80.465 4.612 80.485 5.18 ;
      RECT 80.475 3.63 80.48 4.391 ;
      RECT 80.465 3.582 80.475 4.356 ;
      RECT 80.46 3.545 80.465 4.322 ;
      RECT 80.46 4.692 80.465 5.18 ;
      RECT 80.445 3.522 80.46 4.277 ;
      RECT 80.44 4.79 80.46 5.18 ;
      RECT 80.39 3.41 80.445 4.119 ;
      RECT 80.435 4.912 80.44 5.18 ;
      RECT 80.375 3.41 80.39 3.958 ;
      RECT 80.37 3.41 80.375 3.91 ;
      RECT 80.365 3.41 80.37 3.898 ;
      RECT 80.32 3.41 80.365 3.835 ;
      RECT 80.295 3.41 80.32 3.753 ;
      RECT 80.28 3.41 80.295 3.705 ;
      RECT 80.275 3.41 80.28 3.675 ;
      RECT 79.6 4.86 79.645 5.12 ;
      RECT 79.505 3.395 79.65 3.655 ;
      RECT 80.01 4.017 80.02 4.108 ;
      RECT 79.995 3.955 80.01 4.164 ;
      RECT 79.99 3.902 79.995 4.21 ;
      RECT 79.94 3.849 79.99 4.336 ;
      RECT 79.935 3.804 79.94 4.483 ;
      RECT 79.925 3.792 79.935 4.525 ;
      RECT 79.89 3.756 79.925 4.63 ;
      RECT 79.885 3.724 79.89 4.736 ;
      RECT 79.87 3.706 79.885 4.781 ;
      RECT 79.865 3.689 79.87 4.015 ;
      RECT 79.86 4.07 79.87 4.838 ;
      RECT 79.855 3.675 79.865 3.988 ;
      RECT 79.85 4.125 79.86 5.12 ;
      RECT 79.845 3.661 79.855 3.973 ;
      RECT 79.845 4.175 79.85 5.12 ;
      RECT 79.83 3.638 79.845 3.953 ;
      RECT 79.81 4.297 79.845 5.12 ;
      RECT 79.825 3.62 79.83 3.935 ;
      RECT 79.82 3.612 79.825 3.925 ;
      RECT 79.79 3.58 79.82 3.889 ;
      RECT 79.8 4.425 79.81 5.12 ;
      RECT 79.795 4.452 79.8 5.12 ;
      RECT 79.79 4.502 79.795 5.12 ;
      RECT 79.78 3.546 79.79 3.854 ;
      RECT 79.74 4.57 79.79 5.12 ;
      RECT 79.765 3.523 79.78 3.83 ;
      RECT 79.74 3.395 79.765 3.793 ;
      RECT 79.735 3.395 79.74 3.765 ;
      RECT 79.705 4.67 79.74 5.12 ;
      RECT 79.73 3.395 79.735 3.758 ;
      RECT 79.725 3.395 79.73 3.748 ;
      RECT 79.71 3.395 79.725 3.733 ;
      RECT 79.695 3.395 79.71 3.705 ;
      RECT 79.66 4.775 79.705 5.12 ;
      RECT 79.68 3.395 79.695 3.678 ;
      RECT 79.65 3.395 79.68 3.663 ;
      RECT 79.645 4.847 79.66 5.12 ;
      RECT 79.57 3.93 79.61 4.19 ;
      RECT 79.345 3.877 79.35 4.135 ;
      RECT 75.3 3.355 75.56 3.615 ;
      RECT 75.3 3.38 75.575 3.595 ;
      RECT 77.69 3.205 77.695 3.35 ;
      RECT 79.56 3.925 79.57 4.19 ;
      RECT 79.54 3.917 79.56 4.19 ;
      RECT 79.522 3.913 79.54 4.19 ;
      RECT 79.436 3.902 79.522 4.19 ;
      RECT 79.35 3.885 79.436 4.19 ;
      RECT 79.295 3.872 79.345 4.12 ;
      RECT 79.261 3.864 79.295 4.095 ;
      RECT 79.175 3.853 79.261 4.06 ;
      RECT 79.14 3.83 79.175 4.025 ;
      RECT 79.13 3.792 79.14 4.011 ;
      RECT 79.125 3.765 79.13 4.007 ;
      RECT 79.12 3.752 79.125 4.004 ;
      RECT 79.11 3.732 79.12 4 ;
      RECT 79.105 3.707 79.11 3.996 ;
      RECT 79.08 3.662 79.105 3.99 ;
      RECT 79.07 3.603 79.08 3.982 ;
      RECT 79.06 3.571 79.07 3.973 ;
      RECT 79.04 3.523 79.06 3.953 ;
      RECT 79.035 3.483 79.04 3.923 ;
      RECT 79.02 3.457 79.035 3.897 ;
      RECT 79.015 3.435 79.02 3.873 ;
      RECT 79 3.407 79.015 3.849 ;
      RECT 78.985 3.38 79 3.813 ;
      RECT 78.97 3.357 78.985 3.775 ;
      RECT 78.965 3.347 78.97 3.75 ;
      RECT 78.955 3.34 78.965 3.733 ;
      RECT 78.94 3.327 78.955 3.703 ;
      RECT 78.935 3.317 78.94 3.678 ;
      RECT 78.93 3.312 78.935 3.665 ;
      RECT 78.92 3.305 78.93 3.645 ;
      RECT 78.915 3.298 78.92 3.63 ;
      RECT 78.89 3.291 78.915 3.588 ;
      RECT 78.875 3.281 78.89 3.538 ;
      RECT 78.865 3.276 78.875 3.508 ;
      RECT 78.855 3.272 78.865 3.483 ;
      RECT 78.84 3.269 78.855 3.473 ;
      RECT 78.79 3.266 78.84 3.458 ;
      RECT 78.77 3.264 78.79 3.443 ;
      RECT 78.721 3.262 78.77 3.438 ;
      RECT 78.635 3.258 78.721 3.433 ;
      RECT 78.596 3.255 78.635 3.429 ;
      RECT 78.51 3.251 78.596 3.424 ;
      RECT 78.46 3.248 78.51 3.418 ;
      RECT 78.411 3.245 78.46 3.413 ;
      RECT 78.325 3.242 78.411 3.408 ;
      RECT 78.321 3.24 78.325 3.405 ;
      RECT 78.235 3.237 78.321 3.4 ;
      RECT 78.186 3.233 78.235 3.393 ;
      RECT 78.1 3.23 78.186 3.388 ;
      RECT 78.076 3.227 78.1 3.384 ;
      RECT 77.99 3.225 78.076 3.379 ;
      RECT 77.925 3.221 77.99 3.372 ;
      RECT 77.922 3.22 77.925 3.369 ;
      RECT 77.836 3.217 77.922 3.366 ;
      RECT 77.75 3.211 77.836 3.359 ;
      RECT 77.72 3.207 77.75 3.355 ;
      RECT 77.695 3.205 77.72 3.353 ;
      RECT 77.64 3.202 77.69 3.35 ;
      RECT 77.56 3.201 77.64 3.35 ;
      RECT 77.505 3.203 77.56 3.353 ;
      RECT 77.49 3.204 77.505 3.357 ;
      RECT 77.435 3.212 77.49 3.367 ;
      RECT 77.405 3.22 77.435 3.38 ;
      RECT 77.386 3.221 77.405 3.386 ;
      RECT 77.3 3.224 77.386 3.391 ;
      RECT 77.23 3.229 77.3 3.4 ;
      RECT 77.211 3.232 77.23 3.406 ;
      RECT 77.125 3.236 77.211 3.411 ;
      RECT 77.085 3.24 77.125 3.418 ;
      RECT 77.076 3.242 77.085 3.421 ;
      RECT 76.99 3.246 77.076 3.426 ;
      RECT 76.987 3.249 76.99 3.43 ;
      RECT 76.901 3.252 76.987 3.434 ;
      RECT 76.815 3.258 76.901 3.442 ;
      RECT 76.791 3.262 76.815 3.446 ;
      RECT 76.705 3.266 76.791 3.451 ;
      RECT 76.66 3.271 76.705 3.458 ;
      RECT 76.58 3.276 76.66 3.465 ;
      RECT 76.5 3.282 76.58 3.48 ;
      RECT 76.475 3.286 76.5 3.493 ;
      RECT 76.41 3.289 76.475 3.505 ;
      RECT 76.355 3.294 76.41 3.52 ;
      RECT 76.325 3.297 76.355 3.538 ;
      RECT 76.315 3.299 76.325 3.551 ;
      RECT 76.255 3.314 76.315 3.561 ;
      RECT 76.24 3.331 76.255 3.57 ;
      RECT 76.235 3.34 76.24 3.57 ;
      RECT 76.225 3.35 76.235 3.57 ;
      RECT 76.215 3.367 76.225 3.57 ;
      RECT 76.195 3.377 76.215 3.571 ;
      RECT 76.15 3.387 76.195 3.572 ;
      RECT 76.115 3.396 76.15 3.574 ;
      RECT 76.05 3.401 76.115 3.576 ;
      RECT 75.97 3.402 76.05 3.579 ;
      RECT 75.966 3.4 75.97 3.58 ;
      RECT 75.88 3.397 75.966 3.582 ;
      RECT 75.833 3.394 75.88 3.584 ;
      RECT 75.747 3.39 75.833 3.587 ;
      RECT 75.661 3.386 75.747 3.59 ;
      RECT 75.575 3.382 75.661 3.594 ;
      RECT 77.51 4.445 77.79 4.725 ;
      RECT 77.55 4.425 77.81 4.685 ;
      RECT 77.54 4.435 77.81 4.685 ;
      RECT 77.55 4.362 77.765 4.725 ;
      RECT 77.605 4.285 77.76 4.725 ;
      RECT 77.61 4.07 77.76 4.725 ;
      RECT 77.6 3.872 77.75 4.123 ;
      RECT 77.59 3.872 77.75 3.99 ;
      RECT 77.585 3.75 77.745 3.893 ;
      RECT 77.57 3.75 77.745 3.798 ;
      RECT 77.565 3.46 77.74 3.775 ;
      RECT 77.55 3.46 77.74 3.745 ;
      RECT 77.51 3.46 77.77 3.72 ;
      RECT 77.42 4.93 77.5 5.19 ;
      RECT 76.825 3.65 76.83 3.915 ;
      RECT 76.705 3.65 76.83 3.91 ;
      RECT 77.38 4.895 77.42 5.19 ;
      RECT 77.335 4.817 77.38 5.19 ;
      RECT 77.315 4.745 77.335 5.19 ;
      RECT 77.305 4.697 77.315 5.19 ;
      RECT 77.27 4.63 77.305 5.19 ;
      RECT 77.24 4.53 77.27 5.19 ;
      RECT 77.22 4.455 77.24 4.99 ;
      RECT 77.21 4.405 77.22 4.945 ;
      RECT 77.205 4.382 77.21 4.918 ;
      RECT 77.2 4.367 77.205 4.905 ;
      RECT 77.195 4.352 77.2 4.883 ;
      RECT 77.19 4.337 77.195 4.865 ;
      RECT 77.165 4.292 77.19 4.82 ;
      RECT 77.155 4.24 77.165 4.763 ;
      RECT 77.145 4.21 77.155 4.73 ;
      RECT 77.135 4.175 77.145 4.698 ;
      RECT 77.1 4.107 77.135 4.63 ;
      RECT 77.095 4.046 77.1 4.565 ;
      RECT 77.085 4.034 77.095 4.545 ;
      RECT 77.08 4.022 77.085 4.525 ;
      RECT 77.075 4.014 77.08 4.513 ;
      RECT 77.07 4.006 77.075 4.493 ;
      RECT 77.06 3.994 77.07 4.465 ;
      RECT 77.05 3.978 77.06 4.435 ;
      RECT 77.025 3.95 77.05 4.373 ;
      RECT 77.015 3.921 77.025 4.318 ;
      RECT 77 3.9 77.015 4.278 ;
      RECT 76.995 3.884 77 4.25 ;
      RECT 76.99 3.872 76.995 4.24 ;
      RECT 76.985 3.867 76.99 4.213 ;
      RECT 76.98 3.86 76.985 4.2 ;
      RECT 76.965 3.843 76.98 4.173 ;
      RECT 76.955 3.65 76.965 4.133 ;
      RECT 76.945 3.65 76.955 4.1 ;
      RECT 76.935 3.65 76.945 4.075 ;
      RECT 76.865 3.65 76.935 4.01 ;
      RECT 76.855 3.65 76.865 3.958 ;
      RECT 76.84 3.65 76.855 3.94 ;
      RECT 76.83 3.65 76.84 3.925 ;
      RECT 76.66 4.52 76.92 4.78 ;
      RECT 75.195 4.555 75.2 4.762 ;
      RECT 74.83 4.445 74.905 4.76 ;
      RECT 74.645 4.5 74.8 4.76 ;
      RECT 74.83 4.445 74.935 4.725 ;
      RECT 76.645 4.617 76.66 4.778 ;
      RECT 76.62 4.625 76.645 4.783 ;
      RECT 76.595 4.632 76.62 4.788 ;
      RECT 76.532 4.643 76.595 4.797 ;
      RECT 76.446 4.662 76.532 4.814 ;
      RECT 76.36 4.684 76.446 4.833 ;
      RECT 76.345 4.697 76.36 4.844 ;
      RECT 76.305 4.705 76.345 4.851 ;
      RECT 76.285 4.71 76.305 4.858 ;
      RECT 76.247 4.711 76.285 4.861 ;
      RECT 76.161 4.714 76.247 4.862 ;
      RECT 76.075 4.718 76.161 4.863 ;
      RECT 76.026 4.72 76.075 4.865 ;
      RECT 75.94 4.72 76.026 4.867 ;
      RECT 75.9 4.715 75.94 4.869 ;
      RECT 75.89 4.709 75.9 4.87 ;
      RECT 75.85 4.704 75.89 4.867 ;
      RECT 75.84 4.697 75.85 4.863 ;
      RECT 75.825 4.693 75.84 4.861 ;
      RECT 75.808 4.689 75.825 4.859 ;
      RECT 75.722 4.679 75.808 4.851 ;
      RECT 75.636 4.661 75.722 4.837 ;
      RECT 75.55 4.644 75.636 4.823 ;
      RECT 75.525 4.632 75.55 4.814 ;
      RECT 75.455 4.622 75.525 4.807 ;
      RECT 75.41 4.61 75.455 4.798 ;
      RECT 75.35 4.597 75.41 4.79 ;
      RECT 75.345 4.589 75.35 4.785 ;
      RECT 75.31 4.584 75.345 4.783 ;
      RECT 75.255 4.575 75.31 4.776 ;
      RECT 75.215 4.564 75.255 4.768 ;
      RECT 75.2 4.557 75.215 4.764 ;
      RECT 75.18 4.55 75.195 4.761 ;
      RECT 75.165 4.54 75.18 4.759 ;
      RECT 75.15 4.527 75.165 4.756 ;
      RECT 75.125 4.51 75.15 4.752 ;
      RECT 75.11 4.492 75.125 4.749 ;
      RECT 75.085 4.445 75.11 4.747 ;
      RECT 75.061 4.445 75.085 4.744 ;
      RECT 74.975 4.445 75.061 4.736 ;
      RECT 74.935 4.445 74.975 4.728 ;
      RECT 74.8 4.492 74.83 4.76 ;
      RECT 76.48 4.075 76.74 4.335 ;
      RECT 76.44 4.075 76.74 4.213 ;
      RECT 76.405 4.075 76.74 4.198 ;
      RECT 76.35 4.075 76.74 4.178 ;
      RECT 76.27 3.885 76.55 4.165 ;
      RECT 76.27 4.067 76.62 4.165 ;
      RECT 76.27 4.01 76.605 4.165 ;
      RECT 76.27 3.957 76.555 4.165 ;
      RECT 73.43 4.244 73.445 4.7 ;
      RECT 73.425 4.316 73.531 4.698 ;
      RECT 73.445 3.41 73.58 4.696 ;
      RECT 73.43 4.26 73.585 4.695 ;
      RECT 73.43 4.31 73.59 4.693 ;
      RECT 73.415 4.375 73.59 4.692 ;
      RECT 73.425 4.367 73.595 4.689 ;
      RECT 73.405 4.415 73.595 4.684 ;
      RECT 73.405 4.415 73.61 4.681 ;
      RECT 73.4 4.415 73.61 4.678 ;
      RECT 73.375 4.415 73.635 4.675 ;
      RECT 73.445 3.41 73.605 4.063 ;
      RECT 73.44 3.41 73.605 4.035 ;
      RECT 73.435 3.41 73.605 3.863 ;
      RECT 73.435 3.41 73.625 3.803 ;
      RECT 73.39 3.41 73.65 3.67 ;
      RECT 72.87 3.885 73.15 4.165 ;
      RECT 72.86 3.9 73.15 4.16 ;
      RECT 72.815 3.962 73.15 4.158 ;
      RECT 72.89 3.877 73.055 4.165 ;
      RECT 72.89 3.862 73.011 4.165 ;
      RECT 72.925 3.855 73.011 4.165 ;
      RECT 72.39 5.005 72.67 5.285 ;
      RECT 72.35 4.967 72.645 5.078 ;
      RECT 72.335 4.917 72.625 4.973 ;
      RECT 72.28 4.68 72.54 4.94 ;
      RECT 72.28 4.882 72.62 4.94 ;
      RECT 72.28 4.822 72.615 4.94 ;
      RECT 72.28 4.772 72.595 4.94 ;
      RECT 72.28 4.752 72.59 4.94 ;
      RECT 72.28 4.73 72.585 4.94 ;
      RECT 72.28 4.715 72.555 4.94 ;
      RECT 68 8.66 68.32 8.98 ;
      RECT 68.03 8.13 68.2 8.98 ;
      RECT 68.03 8.13 68.205 8.48 ;
      RECT 68.03 8.13 69.005 8.305 ;
      RECT 68.83 3.26 69.005 8.305 ;
      RECT 68.775 3.26 69.125 3.61 ;
      RECT 68.8 9.09 69.125 9.415 ;
      RECT 67.685 9.18 69.125 9.35 ;
      RECT 67.685 3.69 67.845 9.35 ;
      RECT 68 3.66 68.32 3.98 ;
      RECT 67.685 3.69 68.32 3.86 ;
      RECT 66.365 2.435 66.74 2.805 ;
      RECT 58.275 2.255 58.65 2.625 ;
      RECT 56.84 2.255 57.215 2.625 ;
      RECT 56.84 2.375 66.67 2.545 ;
      RECT 60.96 5.655 66.64 5.825 ;
      RECT 66.47 4.72 66.64 5.825 ;
      RECT 60.77 4.895 60.805 5.825 ;
      RECT 61.035 5.005 61.065 5.285 ;
      RECT 60.74 4.895 60.805 5.155 ;
      RECT 66.38 4.725 66.73 5.075 ;
      RECT 60.57 3.52 60.605 3.78 ;
      RECT 60.345 3.52 60.405 3.78 ;
      RECT 61.025 4.985 61.035 5.285 ;
      RECT 61.02 4.945 61.025 5.285 ;
      RECT 61.005 4.9 61.02 5.285 ;
      RECT 61 4.865 61.005 5.285 ;
      RECT 60.995 4.845 61 5.285 ;
      RECT 60.965 4.772 60.995 5.285 ;
      RECT 60.96 4.7 60.965 5.285 ;
      RECT 60.945 4.66 60.96 5.825 ;
      RECT 60.935 4.6 60.945 5.825 ;
      RECT 60.89 4.54 60.935 5.825 ;
      RECT 60.805 4.501 60.89 5.825 ;
      RECT 60.8 4.492 60.805 4.865 ;
      RECT 60.79 4.491 60.8 4.848 ;
      RECT 60.765 4.472 60.79 4.818 ;
      RECT 60.76 4.447 60.765 4.797 ;
      RECT 60.75 4.425 60.76 4.788 ;
      RECT 60.745 4.396 60.75 4.778 ;
      RECT 60.705 4.322 60.745 4.75 ;
      RECT 60.685 4.223 60.705 4.715 ;
      RECT 60.67 4.159 60.685 4.698 ;
      RECT 60.64 4.083 60.67 4.67 ;
      RECT 60.62 3.998 60.64 4.643 ;
      RECT 60.58 3.894 60.62 4.55 ;
      RECT 60.575 3.815 60.58 4.458 ;
      RECT 60.57 3.798 60.575 4.435 ;
      RECT 60.565 3.52 60.57 4.415 ;
      RECT 60.535 3.52 60.565 4.353 ;
      RECT 60.53 3.52 60.535 4.285 ;
      RECT 60.52 3.52 60.53 4.25 ;
      RECT 60.51 3.52 60.52 4.215 ;
      RECT 60.445 3.52 60.51 4.07 ;
      RECT 60.44 3.52 60.445 3.94 ;
      RECT 60.41 3.52 60.44 3.873 ;
      RECT 60.405 3.52 60.41 3.798 ;
      RECT 64.74 3.455 65 3.715 ;
      RECT 64.735 3.455 65 3.663 ;
      RECT 64.73 3.455 65 3.633 ;
      RECT 64.705 3.325 64.985 3.605 ;
      RECT 53.255 9.095 53.605 9.445 ;
      RECT 64.23 9.05 64.58 9.4 ;
      RECT 53.255 9.125 64.58 9.325 ;
      RECT 63.745 5.005 64.025 5.285 ;
      RECT 63.785 4.96 64.05 5.22 ;
      RECT 63.775 4.995 64.05 5.22 ;
      RECT 63.78 4.98 64.025 5.285 ;
      RECT 63.785 4.957 63.995 5.285 ;
      RECT 63.785 4.955 63.98 5.285 ;
      RECT 63.825 4.945 63.98 5.285 ;
      RECT 63.795 4.95 63.98 5.285 ;
      RECT 63.825 4.942 63.925 5.285 ;
      RECT 63.85 4.935 63.925 5.285 ;
      RECT 63.83 4.937 63.925 5.285 ;
      RECT 63.16 4.45 63.42 4.71 ;
      RECT 63.21 4.442 63.4 4.71 ;
      RECT 63.215 4.362 63.4 4.71 ;
      RECT 63.335 3.75 63.4 4.71 ;
      RECT 63.24 4.147 63.4 4.71 ;
      RECT 63.315 3.835 63.4 4.71 ;
      RECT 63.35 3.46 63.486 4.188 ;
      RECT 63.295 3.957 63.486 4.188 ;
      RECT 63.31 3.897 63.4 4.71 ;
      RECT 63.35 3.46 63.51 3.853 ;
      RECT 63.35 3.46 63.52 3.75 ;
      RECT 63.34 3.46 63.6 3.72 ;
      RECT 62.745 5.005 63.025 5.285 ;
      RECT 62.765 4.965 63.025 5.285 ;
      RECT 62.405 4.92 62.51 5.18 ;
      RECT 62.26 3.41 62.35 3.67 ;
      RECT 62.8 4.475 62.805 4.515 ;
      RECT 62.795 4.465 62.8 4.6 ;
      RECT 62.79 4.455 62.795 4.693 ;
      RECT 62.78 4.435 62.79 4.749 ;
      RECT 62.7 4.363 62.78 4.829 ;
      RECT 62.735 5.007 62.745 5.232 ;
      RECT 62.73 5.004 62.735 5.227 ;
      RECT 62.715 5.001 62.73 5.22 ;
      RECT 62.68 4.995 62.715 5.202 ;
      RECT 62.695 4.298 62.7 4.903 ;
      RECT 62.675 4.249 62.695 4.918 ;
      RECT 62.665 4.982 62.68 5.185 ;
      RECT 62.67 4.191 62.675 4.933 ;
      RECT 62.665 4.169 62.67 4.943 ;
      RECT 62.63 4.079 62.665 5.18 ;
      RECT 62.615 3.957 62.63 5.18 ;
      RECT 62.61 3.91 62.615 5.18 ;
      RECT 62.585 3.835 62.61 5.18 ;
      RECT 62.57 3.75 62.585 5.18 ;
      RECT 62.565 3.697 62.57 5.18 ;
      RECT 62.56 3.677 62.565 5.18 ;
      RECT 62.555 3.652 62.56 4.414 ;
      RECT 62.54 4.612 62.56 5.18 ;
      RECT 62.55 3.63 62.555 4.391 ;
      RECT 62.54 3.582 62.55 4.356 ;
      RECT 62.535 3.545 62.54 4.322 ;
      RECT 62.535 4.692 62.54 5.18 ;
      RECT 62.52 3.522 62.535 4.277 ;
      RECT 62.515 4.79 62.535 5.18 ;
      RECT 62.465 3.41 62.52 4.119 ;
      RECT 62.51 4.912 62.515 5.18 ;
      RECT 62.45 3.41 62.465 3.958 ;
      RECT 62.445 3.41 62.45 3.91 ;
      RECT 62.44 3.41 62.445 3.898 ;
      RECT 62.395 3.41 62.44 3.835 ;
      RECT 62.37 3.41 62.395 3.753 ;
      RECT 62.355 3.41 62.37 3.705 ;
      RECT 62.35 3.41 62.355 3.675 ;
      RECT 61.675 4.86 61.72 5.12 ;
      RECT 61.58 3.395 61.725 3.655 ;
      RECT 62.085 4.017 62.095 4.108 ;
      RECT 62.07 3.955 62.085 4.164 ;
      RECT 62.065 3.902 62.07 4.21 ;
      RECT 62.015 3.849 62.065 4.336 ;
      RECT 62.01 3.804 62.015 4.483 ;
      RECT 62 3.792 62.01 4.525 ;
      RECT 61.965 3.756 62 4.63 ;
      RECT 61.96 3.724 61.965 4.736 ;
      RECT 61.945 3.706 61.96 4.781 ;
      RECT 61.94 3.689 61.945 4.015 ;
      RECT 61.935 4.07 61.945 4.838 ;
      RECT 61.93 3.675 61.94 3.988 ;
      RECT 61.925 4.125 61.935 5.12 ;
      RECT 61.92 3.661 61.93 3.973 ;
      RECT 61.92 4.175 61.925 5.12 ;
      RECT 61.905 3.638 61.92 3.953 ;
      RECT 61.885 4.297 61.92 5.12 ;
      RECT 61.9 3.62 61.905 3.935 ;
      RECT 61.895 3.612 61.9 3.925 ;
      RECT 61.865 3.58 61.895 3.889 ;
      RECT 61.875 4.425 61.885 5.12 ;
      RECT 61.87 4.452 61.875 5.12 ;
      RECT 61.865 4.502 61.87 5.12 ;
      RECT 61.855 3.546 61.865 3.854 ;
      RECT 61.815 4.57 61.865 5.12 ;
      RECT 61.84 3.523 61.855 3.83 ;
      RECT 61.815 3.395 61.84 3.793 ;
      RECT 61.81 3.395 61.815 3.765 ;
      RECT 61.78 4.67 61.815 5.12 ;
      RECT 61.805 3.395 61.81 3.758 ;
      RECT 61.8 3.395 61.805 3.748 ;
      RECT 61.785 3.395 61.8 3.733 ;
      RECT 61.77 3.395 61.785 3.705 ;
      RECT 61.735 4.775 61.78 5.12 ;
      RECT 61.755 3.395 61.77 3.678 ;
      RECT 61.725 3.395 61.755 3.663 ;
      RECT 61.72 4.847 61.735 5.12 ;
      RECT 61.645 3.93 61.685 4.19 ;
      RECT 61.42 3.877 61.425 4.135 ;
      RECT 57.375 3.355 57.635 3.615 ;
      RECT 57.375 3.38 57.65 3.595 ;
      RECT 59.765 3.205 59.77 3.35 ;
      RECT 61.635 3.925 61.645 4.19 ;
      RECT 61.615 3.917 61.635 4.19 ;
      RECT 61.597 3.913 61.615 4.19 ;
      RECT 61.511 3.902 61.597 4.19 ;
      RECT 61.425 3.885 61.511 4.19 ;
      RECT 61.37 3.872 61.42 4.12 ;
      RECT 61.336 3.864 61.37 4.095 ;
      RECT 61.25 3.853 61.336 4.06 ;
      RECT 61.215 3.83 61.25 4.025 ;
      RECT 61.205 3.792 61.215 4.011 ;
      RECT 61.2 3.765 61.205 4.007 ;
      RECT 61.195 3.752 61.2 4.004 ;
      RECT 61.185 3.732 61.195 4 ;
      RECT 61.18 3.707 61.185 3.996 ;
      RECT 61.155 3.662 61.18 3.99 ;
      RECT 61.145 3.603 61.155 3.982 ;
      RECT 61.135 3.571 61.145 3.973 ;
      RECT 61.115 3.523 61.135 3.953 ;
      RECT 61.11 3.483 61.115 3.923 ;
      RECT 61.095 3.457 61.11 3.897 ;
      RECT 61.09 3.435 61.095 3.873 ;
      RECT 61.075 3.407 61.09 3.849 ;
      RECT 61.06 3.38 61.075 3.813 ;
      RECT 61.045 3.357 61.06 3.775 ;
      RECT 61.04 3.347 61.045 3.75 ;
      RECT 61.03 3.34 61.04 3.733 ;
      RECT 61.015 3.327 61.03 3.703 ;
      RECT 61.01 3.317 61.015 3.678 ;
      RECT 61.005 3.312 61.01 3.665 ;
      RECT 60.995 3.305 61.005 3.645 ;
      RECT 60.99 3.298 60.995 3.63 ;
      RECT 60.965 3.291 60.99 3.588 ;
      RECT 60.95 3.281 60.965 3.538 ;
      RECT 60.94 3.276 60.95 3.508 ;
      RECT 60.93 3.272 60.94 3.483 ;
      RECT 60.915 3.269 60.93 3.473 ;
      RECT 60.865 3.266 60.915 3.458 ;
      RECT 60.845 3.264 60.865 3.443 ;
      RECT 60.796 3.262 60.845 3.438 ;
      RECT 60.71 3.258 60.796 3.433 ;
      RECT 60.671 3.255 60.71 3.429 ;
      RECT 60.585 3.251 60.671 3.424 ;
      RECT 60.535 3.248 60.585 3.418 ;
      RECT 60.486 3.245 60.535 3.413 ;
      RECT 60.4 3.242 60.486 3.408 ;
      RECT 60.396 3.24 60.4 3.405 ;
      RECT 60.31 3.237 60.396 3.4 ;
      RECT 60.261 3.233 60.31 3.393 ;
      RECT 60.175 3.23 60.261 3.388 ;
      RECT 60.151 3.227 60.175 3.384 ;
      RECT 60.065 3.225 60.151 3.379 ;
      RECT 60 3.221 60.065 3.372 ;
      RECT 59.997 3.22 60 3.369 ;
      RECT 59.911 3.217 59.997 3.366 ;
      RECT 59.825 3.211 59.911 3.359 ;
      RECT 59.795 3.207 59.825 3.355 ;
      RECT 59.77 3.205 59.795 3.353 ;
      RECT 59.715 3.202 59.765 3.35 ;
      RECT 59.635 3.201 59.715 3.35 ;
      RECT 59.58 3.203 59.635 3.353 ;
      RECT 59.565 3.204 59.58 3.357 ;
      RECT 59.51 3.212 59.565 3.367 ;
      RECT 59.48 3.22 59.51 3.38 ;
      RECT 59.461 3.221 59.48 3.386 ;
      RECT 59.375 3.224 59.461 3.391 ;
      RECT 59.305 3.229 59.375 3.4 ;
      RECT 59.286 3.232 59.305 3.406 ;
      RECT 59.2 3.236 59.286 3.411 ;
      RECT 59.16 3.24 59.2 3.418 ;
      RECT 59.151 3.242 59.16 3.421 ;
      RECT 59.065 3.246 59.151 3.426 ;
      RECT 59.062 3.249 59.065 3.43 ;
      RECT 58.976 3.252 59.062 3.434 ;
      RECT 58.89 3.258 58.976 3.442 ;
      RECT 58.866 3.262 58.89 3.446 ;
      RECT 58.78 3.266 58.866 3.451 ;
      RECT 58.735 3.271 58.78 3.458 ;
      RECT 58.655 3.276 58.735 3.465 ;
      RECT 58.575 3.282 58.655 3.48 ;
      RECT 58.55 3.286 58.575 3.493 ;
      RECT 58.485 3.289 58.55 3.505 ;
      RECT 58.43 3.294 58.485 3.52 ;
      RECT 58.4 3.297 58.43 3.538 ;
      RECT 58.39 3.299 58.4 3.551 ;
      RECT 58.33 3.314 58.39 3.561 ;
      RECT 58.315 3.331 58.33 3.57 ;
      RECT 58.31 3.34 58.315 3.57 ;
      RECT 58.3 3.35 58.31 3.57 ;
      RECT 58.29 3.367 58.3 3.57 ;
      RECT 58.27 3.377 58.29 3.571 ;
      RECT 58.225 3.387 58.27 3.572 ;
      RECT 58.19 3.396 58.225 3.574 ;
      RECT 58.125 3.401 58.19 3.576 ;
      RECT 58.045 3.402 58.125 3.579 ;
      RECT 58.041 3.4 58.045 3.58 ;
      RECT 57.955 3.397 58.041 3.582 ;
      RECT 57.908 3.394 57.955 3.584 ;
      RECT 57.822 3.39 57.908 3.587 ;
      RECT 57.736 3.386 57.822 3.59 ;
      RECT 57.65 3.382 57.736 3.594 ;
      RECT 59.585 4.445 59.865 4.725 ;
      RECT 59.625 4.425 59.885 4.685 ;
      RECT 59.615 4.435 59.885 4.685 ;
      RECT 59.625 4.362 59.84 4.725 ;
      RECT 59.68 4.285 59.835 4.725 ;
      RECT 59.685 4.07 59.835 4.725 ;
      RECT 59.675 3.872 59.825 4.123 ;
      RECT 59.665 3.872 59.825 3.99 ;
      RECT 59.66 3.75 59.82 3.893 ;
      RECT 59.645 3.75 59.82 3.798 ;
      RECT 59.64 3.46 59.815 3.775 ;
      RECT 59.625 3.46 59.815 3.745 ;
      RECT 59.585 3.46 59.845 3.72 ;
      RECT 59.495 4.93 59.575 5.19 ;
      RECT 58.9 3.65 58.905 3.915 ;
      RECT 58.78 3.65 58.905 3.91 ;
      RECT 59.455 4.895 59.495 5.19 ;
      RECT 59.41 4.817 59.455 5.19 ;
      RECT 59.39 4.745 59.41 5.19 ;
      RECT 59.38 4.697 59.39 5.19 ;
      RECT 59.345 4.63 59.38 5.19 ;
      RECT 59.315 4.53 59.345 5.19 ;
      RECT 59.295 4.455 59.315 4.99 ;
      RECT 59.285 4.405 59.295 4.945 ;
      RECT 59.28 4.382 59.285 4.918 ;
      RECT 59.275 4.367 59.28 4.905 ;
      RECT 59.27 4.352 59.275 4.883 ;
      RECT 59.265 4.337 59.27 4.865 ;
      RECT 59.24 4.292 59.265 4.82 ;
      RECT 59.23 4.24 59.24 4.763 ;
      RECT 59.22 4.21 59.23 4.73 ;
      RECT 59.21 4.175 59.22 4.698 ;
      RECT 59.175 4.107 59.21 4.63 ;
      RECT 59.17 4.046 59.175 4.565 ;
      RECT 59.16 4.034 59.17 4.545 ;
      RECT 59.155 4.022 59.16 4.525 ;
      RECT 59.15 4.014 59.155 4.513 ;
      RECT 59.145 4.006 59.15 4.493 ;
      RECT 59.135 3.994 59.145 4.465 ;
      RECT 59.125 3.978 59.135 4.435 ;
      RECT 59.1 3.95 59.125 4.373 ;
      RECT 59.09 3.921 59.1 4.318 ;
      RECT 59.075 3.9 59.09 4.278 ;
      RECT 59.07 3.884 59.075 4.25 ;
      RECT 59.065 3.872 59.07 4.24 ;
      RECT 59.06 3.867 59.065 4.213 ;
      RECT 59.055 3.86 59.06 4.2 ;
      RECT 59.04 3.843 59.055 4.173 ;
      RECT 59.03 3.65 59.04 4.133 ;
      RECT 59.02 3.65 59.03 4.1 ;
      RECT 59.01 3.65 59.02 4.075 ;
      RECT 58.94 3.65 59.01 4.01 ;
      RECT 58.93 3.65 58.94 3.958 ;
      RECT 58.915 3.65 58.93 3.94 ;
      RECT 58.905 3.65 58.915 3.925 ;
      RECT 58.735 4.52 58.995 4.78 ;
      RECT 57.27 4.555 57.275 4.762 ;
      RECT 56.905 4.445 56.98 4.76 ;
      RECT 56.72 4.5 56.875 4.76 ;
      RECT 56.905 4.445 57.01 4.725 ;
      RECT 58.72 4.617 58.735 4.778 ;
      RECT 58.695 4.625 58.72 4.783 ;
      RECT 58.67 4.632 58.695 4.788 ;
      RECT 58.607 4.643 58.67 4.797 ;
      RECT 58.521 4.662 58.607 4.814 ;
      RECT 58.435 4.684 58.521 4.833 ;
      RECT 58.42 4.697 58.435 4.844 ;
      RECT 58.38 4.705 58.42 4.851 ;
      RECT 58.36 4.71 58.38 4.858 ;
      RECT 58.322 4.711 58.36 4.861 ;
      RECT 58.236 4.714 58.322 4.862 ;
      RECT 58.15 4.718 58.236 4.863 ;
      RECT 58.101 4.72 58.15 4.865 ;
      RECT 58.015 4.72 58.101 4.867 ;
      RECT 57.975 4.715 58.015 4.869 ;
      RECT 57.965 4.709 57.975 4.87 ;
      RECT 57.925 4.704 57.965 4.867 ;
      RECT 57.915 4.697 57.925 4.863 ;
      RECT 57.9 4.693 57.915 4.861 ;
      RECT 57.883 4.689 57.9 4.859 ;
      RECT 57.797 4.679 57.883 4.851 ;
      RECT 57.711 4.661 57.797 4.837 ;
      RECT 57.625 4.644 57.711 4.823 ;
      RECT 57.6 4.632 57.625 4.814 ;
      RECT 57.53 4.622 57.6 4.807 ;
      RECT 57.485 4.61 57.53 4.798 ;
      RECT 57.425 4.597 57.485 4.79 ;
      RECT 57.42 4.589 57.425 4.785 ;
      RECT 57.385 4.584 57.42 4.783 ;
      RECT 57.33 4.575 57.385 4.776 ;
      RECT 57.29 4.564 57.33 4.768 ;
      RECT 57.275 4.557 57.29 4.764 ;
      RECT 57.255 4.55 57.27 4.761 ;
      RECT 57.24 4.54 57.255 4.759 ;
      RECT 57.225 4.527 57.24 4.756 ;
      RECT 57.2 4.51 57.225 4.752 ;
      RECT 57.185 4.492 57.2 4.749 ;
      RECT 57.16 4.445 57.185 4.747 ;
      RECT 57.136 4.445 57.16 4.744 ;
      RECT 57.05 4.445 57.136 4.736 ;
      RECT 57.01 4.445 57.05 4.728 ;
      RECT 56.875 4.492 56.905 4.76 ;
      RECT 58.555 4.075 58.815 4.335 ;
      RECT 58.515 4.075 58.815 4.213 ;
      RECT 58.48 4.075 58.815 4.198 ;
      RECT 58.425 4.075 58.815 4.178 ;
      RECT 58.345 3.885 58.625 4.165 ;
      RECT 58.345 4.067 58.695 4.165 ;
      RECT 58.345 4.01 58.68 4.165 ;
      RECT 58.345 3.957 58.63 4.165 ;
      RECT 55.505 4.244 55.52 4.7 ;
      RECT 55.5 4.316 55.606 4.698 ;
      RECT 55.52 3.41 55.655 4.696 ;
      RECT 55.505 4.26 55.66 4.695 ;
      RECT 55.505 4.31 55.665 4.693 ;
      RECT 55.49 4.375 55.665 4.692 ;
      RECT 55.5 4.367 55.67 4.689 ;
      RECT 55.48 4.415 55.67 4.684 ;
      RECT 55.48 4.415 55.685 4.681 ;
      RECT 55.475 4.415 55.685 4.678 ;
      RECT 55.45 4.415 55.71 4.675 ;
      RECT 55.52 3.41 55.68 4.063 ;
      RECT 55.515 3.41 55.68 4.035 ;
      RECT 55.51 3.41 55.68 3.863 ;
      RECT 55.51 3.41 55.7 3.803 ;
      RECT 55.465 3.41 55.725 3.67 ;
      RECT 54.945 3.885 55.225 4.165 ;
      RECT 54.935 3.9 55.225 4.16 ;
      RECT 54.89 3.962 55.225 4.158 ;
      RECT 54.965 3.877 55.13 4.165 ;
      RECT 54.965 3.862 55.086 4.165 ;
      RECT 55 3.855 55.086 4.165 ;
      RECT 54.465 5.005 54.745 5.285 ;
      RECT 54.425 4.967 54.72 5.078 ;
      RECT 54.41 4.917 54.7 4.973 ;
      RECT 54.355 4.68 54.615 4.94 ;
      RECT 54.355 4.882 54.695 4.94 ;
      RECT 54.355 4.822 54.69 4.94 ;
      RECT 54.355 4.772 54.67 4.94 ;
      RECT 54.355 4.752 54.665 4.94 ;
      RECT 54.355 4.73 54.66 4.94 ;
      RECT 54.355 4.715 54.63 4.94 ;
      RECT 50.075 8.66 50.395 8.98 ;
      RECT 50.105 8.13 50.275 8.98 ;
      RECT 50.105 8.13 50.28 8.48 ;
      RECT 50.105 8.13 51.08 8.305 ;
      RECT 50.905 3.26 51.08 8.305 ;
      RECT 50.85 3.26 51.2 3.61 ;
      RECT 50.875 9.09 51.2 9.415 ;
      RECT 49.76 9.18 51.2 9.35 ;
      RECT 49.76 3.69 49.92 9.35 ;
      RECT 50.075 3.66 50.395 3.98 ;
      RECT 49.76 3.69 50.395 3.86 ;
      RECT 48.44 2.435 48.815 2.805 ;
      RECT 40.35 2.255 40.725 2.625 ;
      RECT 38.915 2.255 39.29 2.625 ;
      RECT 38.915 2.375 48.745 2.545 ;
      RECT 43.035 5.655 48.715 5.825 ;
      RECT 48.545 4.72 48.715 5.825 ;
      RECT 42.845 4.895 42.88 5.825 ;
      RECT 43.11 5.005 43.14 5.285 ;
      RECT 42.815 4.895 42.88 5.155 ;
      RECT 48.455 4.725 48.805 5.075 ;
      RECT 42.645 3.52 42.68 3.78 ;
      RECT 42.42 3.52 42.48 3.78 ;
      RECT 43.1 4.985 43.11 5.285 ;
      RECT 43.095 4.945 43.1 5.285 ;
      RECT 43.08 4.9 43.095 5.285 ;
      RECT 43.075 4.865 43.08 5.285 ;
      RECT 43.07 4.845 43.075 5.285 ;
      RECT 43.04 4.772 43.07 5.285 ;
      RECT 43.035 4.7 43.04 5.285 ;
      RECT 43.02 4.66 43.035 5.825 ;
      RECT 43.01 4.6 43.02 5.825 ;
      RECT 42.965 4.54 43.01 5.825 ;
      RECT 42.88 4.501 42.965 5.825 ;
      RECT 42.875 4.492 42.88 4.865 ;
      RECT 42.865 4.491 42.875 4.848 ;
      RECT 42.84 4.472 42.865 4.818 ;
      RECT 42.835 4.447 42.84 4.797 ;
      RECT 42.825 4.425 42.835 4.788 ;
      RECT 42.82 4.396 42.825 4.778 ;
      RECT 42.78 4.322 42.82 4.75 ;
      RECT 42.76 4.223 42.78 4.715 ;
      RECT 42.745 4.159 42.76 4.698 ;
      RECT 42.715 4.083 42.745 4.67 ;
      RECT 42.695 3.998 42.715 4.643 ;
      RECT 42.655 3.894 42.695 4.55 ;
      RECT 42.65 3.815 42.655 4.458 ;
      RECT 42.645 3.798 42.65 4.435 ;
      RECT 42.64 3.52 42.645 4.415 ;
      RECT 42.61 3.52 42.64 4.353 ;
      RECT 42.605 3.52 42.61 4.285 ;
      RECT 42.595 3.52 42.605 4.25 ;
      RECT 42.585 3.52 42.595 4.215 ;
      RECT 42.52 3.52 42.585 4.07 ;
      RECT 42.515 3.52 42.52 3.94 ;
      RECT 42.485 3.52 42.515 3.873 ;
      RECT 42.48 3.52 42.485 3.798 ;
      RECT 46.815 3.455 47.075 3.715 ;
      RECT 46.81 3.455 47.075 3.663 ;
      RECT 46.805 3.455 47.075 3.633 ;
      RECT 46.78 3.325 47.06 3.605 ;
      RECT 35.33 9.095 35.68 9.445 ;
      RECT 46.3 9.05 46.65 9.4 ;
      RECT 35.33 9.125 46.65 9.325 ;
      RECT 45.82 5.005 46.1 5.285 ;
      RECT 45.86 4.96 46.125 5.22 ;
      RECT 45.85 4.995 46.125 5.22 ;
      RECT 45.855 4.98 46.1 5.285 ;
      RECT 45.86 4.957 46.07 5.285 ;
      RECT 45.86 4.955 46.055 5.285 ;
      RECT 45.9 4.945 46.055 5.285 ;
      RECT 45.87 4.95 46.055 5.285 ;
      RECT 45.9 4.942 46 5.285 ;
      RECT 45.925 4.935 46 5.285 ;
      RECT 45.905 4.937 46 5.285 ;
      RECT 45.235 4.45 45.495 4.71 ;
      RECT 45.285 4.442 45.475 4.71 ;
      RECT 45.29 4.362 45.475 4.71 ;
      RECT 45.41 3.75 45.475 4.71 ;
      RECT 45.315 4.147 45.475 4.71 ;
      RECT 45.39 3.835 45.475 4.71 ;
      RECT 45.425 3.46 45.561 4.188 ;
      RECT 45.37 3.957 45.561 4.188 ;
      RECT 45.385 3.897 45.475 4.71 ;
      RECT 45.425 3.46 45.585 3.853 ;
      RECT 45.425 3.46 45.595 3.75 ;
      RECT 45.415 3.46 45.675 3.72 ;
      RECT 44.82 5.005 45.1 5.285 ;
      RECT 44.84 4.965 45.1 5.285 ;
      RECT 44.48 4.92 44.585 5.18 ;
      RECT 44.335 3.41 44.425 3.67 ;
      RECT 44.875 4.475 44.88 4.515 ;
      RECT 44.87 4.465 44.875 4.6 ;
      RECT 44.865 4.455 44.87 4.693 ;
      RECT 44.855 4.435 44.865 4.749 ;
      RECT 44.775 4.363 44.855 4.829 ;
      RECT 44.81 5.007 44.82 5.232 ;
      RECT 44.805 5.004 44.81 5.227 ;
      RECT 44.79 5.001 44.805 5.22 ;
      RECT 44.755 4.995 44.79 5.202 ;
      RECT 44.77 4.298 44.775 4.903 ;
      RECT 44.75 4.249 44.77 4.918 ;
      RECT 44.74 4.982 44.755 5.185 ;
      RECT 44.745 4.191 44.75 4.933 ;
      RECT 44.74 4.169 44.745 4.943 ;
      RECT 44.705 4.079 44.74 5.18 ;
      RECT 44.69 3.957 44.705 5.18 ;
      RECT 44.685 3.91 44.69 5.18 ;
      RECT 44.66 3.835 44.685 5.18 ;
      RECT 44.645 3.75 44.66 5.18 ;
      RECT 44.64 3.697 44.645 5.18 ;
      RECT 44.635 3.677 44.64 5.18 ;
      RECT 44.63 3.652 44.635 4.414 ;
      RECT 44.615 4.612 44.635 5.18 ;
      RECT 44.625 3.63 44.63 4.391 ;
      RECT 44.615 3.582 44.625 4.356 ;
      RECT 44.61 3.545 44.615 4.322 ;
      RECT 44.61 4.692 44.615 5.18 ;
      RECT 44.595 3.522 44.61 4.277 ;
      RECT 44.59 4.79 44.61 5.18 ;
      RECT 44.54 3.41 44.595 4.119 ;
      RECT 44.585 4.912 44.59 5.18 ;
      RECT 44.525 3.41 44.54 3.958 ;
      RECT 44.52 3.41 44.525 3.91 ;
      RECT 44.515 3.41 44.52 3.898 ;
      RECT 44.47 3.41 44.515 3.835 ;
      RECT 44.445 3.41 44.47 3.753 ;
      RECT 44.43 3.41 44.445 3.705 ;
      RECT 44.425 3.41 44.43 3.675 ;
      RECT 43.75 4.86 43.795 5.12 ;
      RECT 43.655 3.395 43.8 3.655 ;
      RECT 44.16 4.017 44.17 4.108 ;
      RECT 44.145 3.955 44.16 4.164 ;
      RECT 44.14 3.902 44.145 4.21 ;
      RECT 44.09 3.849 44.14 4.336 ;
      RECT 44.085 3.804 44.09 4.483 ;
      RECT 44.075 3.792 44.085 4.525 ;
      RECT 44.04 3.756 44.075 4.63 ;
      RECT 44.035 3.724 44.04 4.736 ;
      RECT 44.02 3.706 44.035 4.781 ;
      RECT 44.015 3.689 44.02 4.015 ;
      RECT 44.01 4.07 44.02 4.838 ;
      RECT 44.005 3.675 44.015 3.988 ;
      RECT 44 4.125 44.01 5.12 ;
      RECT 43.995 3.661 44.005 3.973 ;
      RECT 43.995 4.175 44 5.12 ;
      RECT 43.98 3.638 43.995 3.953 ;
      RECT 43.96 4.297 43.995 5.12 ;
      RECT 43.975 3.62 43.98 3.935 ;
      RECT 43.97 3.612 43.975 3.925 ;
      RECT 43.94 3.58 43.97 3.889 ;
      RECT 43.95 4.425 43.96 5.12 ;
      RECT 43.945 4.452 43.95 5.12 ;
      RECT 43.94 4.502 43.945 5.12 ;
      RECT 43.93 3.546 43.94 3.854 ;
      RECT 43.89 4.57 43.94 5.12 ;
      RECT 43.915 3.523 43.93 3.83 ;
      RECT 43.89 3.395 43.915 3.793 ;
      RECT 43.885 3.395 43.89 3.765 ;
      RECT 43.855 4.67 43.89 5.12 ;
      RECT 43.88 3.395 43.885 3.758 ;
      RECT 43.875 3.395 43.88 3.748 ;
      RECT 43.86 3.395 43.875 3.733 ;
      RECT 43.845 3.395 43.86 3.705 ;
      RECT 43.81 4.775 43.855 5.12 ;
      RECT 43.83 3.395 43.845 3.678 ;
      RECT 43.8 3.395 43.83 3.663 ;
      RECT 43.795 4.847 43.81 5.12 ;
      RECT 43.72 3.93 43.76 4.19 ;
      RECT 43.495 3.877 43.5 4.135 ;
      RECT 39.45 3.355 39.71 3.615 ;
      RECT 39.45 3.38 39.725 3.595 ;
      RECT 41.84 3.205 41.845 3.35 ;
      RECT 43.71 3.925 43.72 4.19 ;
      RECT 43.69 3.917 43.71 4.19 ;
      RECT 43.672 3.913 43.69 4.19 ;
      RECT 43.586 3.902 43.672 4.19 ;
      RECT 43.5 3.885 43.586 4.19 ;
      RECT 43.445 3.872 43.495 4.12 ;
      RECT 43.411 3.864 43.445 4.095 ;
      RECT 43.325 3.853 43.411 4.06 ;
      RECT 43.29 3.83 43.325 4.025 ;
      RECT 43.28 3.792 43.29 4.011 ;
      RECT 43.275 3.765 43.28 4.007 ;
      RECT 43.27 3.752 43.275 4.004 ;
      RECT 43.26 3.732 43.27 4 ;
      RECT 43.255 3.707 43.26 3.996 ;
      RECT 43.23 3.662 43.255 3.99 ;
      RECT 43.22 3.603 43.23 3.982 ;
      RECT 43.21 3.571 43.22 3.973 ;
      RECT 43.19 3.523 43.21 3.953 ;
      RECT 43.185 3.483 43.19 3.923 ;
      RECT 43.17 3.457 43.185 3.897 ;
      RECT 43.165 3.435 43.17 3.873 ;
      RECT 43.15 3.407 43.165 3.849 ;
      RECT 43.135 3.38 43.15 3.813 ;
      RECT 43.12 3.357 43.135 3.775 ;
      RECT 43.115 3.347 43.12 3.75 ;
      RECT 43.105 3.34 43.115 3.733 ;
      RECT 43.09 3.327 43.105 3.703 ;
      RECT 43.085 3.317 43.09 3.678 ;
      RECT 43.08 3.312 43.085 3.665 ;
      RECT 43.07 3.305 43.08 3.645 ;
      RECT 43.065 3.298 43.07 3.63 ;
      RECT 43.04 3.291 43.065 3.588 ;
      RECT 43.025 3.281 43.04 3.538 ;
      RECT 43.015 3.276 43.025 3.508 ;
      RECT 43.005 3.272 43.015 3.483 ;
      RECT 42.99 3.269 43.005 3.473 ;
      RECT 42.94 3.266 42.99 3.458 ;
      RECT 42.92 3.264 42.94 3.443 ;
      RECT 42.871 3.262 42.92 3.438 ;
      RECT 42.785 3.258 42.871 3.433 ;
      RECT 42.746 3.255 42.785 3.429 ;
      RECT 42.66 3.251 42.746 3.424 ;
      RECT 42.61 3.248 42.66 3.418 ;
      RECT 42.561 3.245 42.61 3.413 ;
      RECT 42.475 3.242 42.561 3.408 ;
      RECT 42.471 3.24 42.475 3.405 ;
      RECT 42.385 3.237 42.471 3.4 ;
      RECT 42.336 3.233 42.385 3.393 ;
      RECT 42.25 3.23 42.336 3.388 ;
      RECT 42.226 3.227 42.25 3.384 ;
      RECT 42.14 3.225 42.226 3.379 ;
      RECT 42.075 3.221 42.14 3.372 ;
      RECT 42.072 3.22 42.075 3.369 ;
      RECT 41.986 3.217 42.072 3.366 ;
      RECT 41.9 3.211 41.986 3.359 ;
      RECT 41.87 3.207 41.9 3.355 ;
      RECT 41.845 3.205 41.87 3.353 ;
      RECT 41.79 3.202 41.84 3.35 ;
      RECT 41.71 3.201 41.79 3.35 ;
      RECT 41.655 3.203 41.71 3.353 ;
      RECT 41.64 3.204 41.655 3.357 ;
      RECT 41.585 3.212 41.64 3.367 ;
      RECT 41.555 3.22 41.585 3.38 ;
      RECT 41.536 3.221 41.555 3.386 ;
      RECT 41.45 3.224 41.536 3.391 ;
      RECT 41.38 3.229 41.45 3.4 ;
      RECT 41.361 3.232 41.38 3.406 ;
      RECT 41.275 3.236 41.361 3.411 ;
      RECT 41.235 3.24 41.275 3.418 ;
      RECT 41.226 3.242 41.235 3.421 ;
      RECT 41.14 3.246 41.226 3.426 ;
      RECT 41.137 3.249 41.14 3.43 ;
      RECT 41.051 3.252 41.137 3.434 ;
      RECT 40.965 3.258 41.051 3.442 ;
      RECT 40.941 3.262 40.965 3.446 ;
      RECT 40.855 3.266 40.941 3.451 ;
      RECT 40.81 3.271 40.855 3.458 ;
      RECT 40.73 3.276 40.81 3.465 ;
      RECT 40.65 3.282 40.73 3.48 ;
      RECT 40.625 3.286 40.65 3.493 ;
      RECT 40.56 3.289 40.625 3.505 ;
      RECT 40.505 3.294 40.56 3.52 ;
      RECT 40.475 3.297 40.505 3.538 ;
      RECT 40.465 3.299 40.475 3.551 ;
      RECT 40.405 3.314 40.465 3.561 ;
      RECT 40.39 3.331 40.405 3.57 ;
      RECT 40.385 3.34 40.39 3.57 ;
      RECT 40.375 3.35 40.385 3.57 ;
      RECT 40.365 3.367 40.375 3.57 ;
      RECT 40.345 3.377 40.365 3.571 ;
      RECT 40.3 3.387 40.345 3.572 ;
      RECT 40.265 3.396 40.3 3.574 ;
      RECT 40.2 3.401 40.265 3.576 ;
      RECT 40.12 3.402 40.2 3.579 ;
      RECT 40.116 3.4 40.12 3.58 ;
      RECT 40.03 3.397 40.116 3.582 ;
      RECT 39.983 3.394 40.03 3.584 ;
      RECT 39.897 3.39 39.983 3.587 ;
      RECT 39.811 3.386 39.897 3.59 ;
      RECT 39.725 3.382 39.811 3.594 ;
      RECT 41.66 4.445 41.94 4.725 ;
      RECT 41.7 4.425 41.96 4.685 ;
      RECT 41.69 4.435 41.96 4.685 ;
      RECT 41.7 4.362 41.915 4.725 ;
      RECT 41.755 4.285 41.91 4.725 ;
      RECT 41.76 4.07 41.91 4.725 ;
      RECT 41.75 3.872 41.9 4.123 ;
      RECT 41.74 3.872 41.9 3.99 ;
      RECT 41.735 3.75 41.895 3.893 ;
      RECT 41.72 3.75 41.895 3.798 ;
      RECT 41.715 3.46 41.89 3.775 ;
      RECT 41.7 3.46 41.89 3.745 ;
      RECT 41.66 3.46 41.92 3.72 ;
      RECT 41.57 4.93 41.65 5.19 ;
      RECT 40.975 3.65 40.98 3.915 ;
      RECT 40.855 3.65 40.98 3.91 ;
      RECT 41.53 4.895 41.57 5.19 ;
      RECT 41.485 4.817 41.53 5.19 ;
      RECT 41.465 4.745 41.485 5.19 ;
      RECT 41.455 4.697 41.465 5.19 ;
      RECT 41.42 4.63 41.455 5.19 ;
      RECT 41.39 4.53 41.42 5.19 ;
      RECT 41.37 4.455 41.39 4.99 ;
      RECT 41.36 4.405 41.37 4.945 ;
      RECT 41.355 4.382 41.36 4.918 ;
      RECT 41.35 4.367 41.355 4.905 ;
      RECT 41.345 4.352 41.35 4.883 ;
      RECT 41.34 4.337 41.345 4.865 ;
      RECT 41.315 4.292 41.34 4.82 ;
      RECT 41.305 4.24 41.315 4.763 ;
      RECT 41.295 4.21 41.305 4.73 ;
      RECT 41.285 4.175 41.295 4.698 ;
      RECT 41.25 4.107 41.285 4.63 ;
      RECT 41.245 4.046 41.25 4.565 ;
      RECT 41.235 4.034 41.245 4.545 ;
      RECT 41.23 4.022 41.235 4.525 ;
      RECT 41.225 4.014 41.23 4.513 ;
      RECT 41.22 4.006 41.225 4.493 ;
      RECT 41.21 3.994 41.22 4.465 ;
      RECT 41.2 3.978 41.21 4.435 ;
      RECT 41.175 3.95 41.2 4.373 ;
      RECT 41.165 3.921 41.175 4.318 ;
      RECT 41.15 3.9 41.165 4.278 ;
      RECT 41.145 3.884 41.15 4.25 ;
      RECT 41.14 3.872 41.145 4.24 ;
      RECT 41.135 3.867 41.14 4.213 ;
      RECT 41.13 3.86 41.135 4.2 ;
      RECT 41.115 3.843 41.13 4.173 ;
      RECT 41.105 3.65 41.115 4.133 ;
      RECT 41.095 3.65 41.105 4.1 ;
      RECT 41.085 3.65 41.095 4.075 ;
      RECT 41.015 3.65 41.085 4.01 ;
      RECT 41.005 3.65 41.015 3.958 ;
      RECT 40.99 3.65 41.005 3.94 ;
      RECT 40.98 3.65 40.99 3.925 ;
      RECT 40.81 4.52 41.07 4.78 ;
      RECT 39.345 4.555 39.35 4.762 ;
      RECT 38.98 4.445 39.055 4.76 ;
      RECT 38.795 4.5 38.95 4.76 ;
      RECT 38.98 4.445 39.085 4.725 ;
      RECT 40.795 4.617 40.81 4.778 ;
      RECT 40.77 4.625 40.795 4.783 ;
      RECT 40.745 4.632 40.77 4.788 ;
      RECT 40.682 4.643 40.745 4.797 ;
      RECT 40.596 4.662 40.682 4.814 ;
      RECT 40.51 4.684 40.596 4.833 ;
      RECT 40.495 4.697 40.51 4.844 ;
      RECT 40.455 4.705 40.495 4.851 ;
      RECT 40.435 4.71 40.455 4.858 ;
      RECT 40.397 4.711 40.435 4.861 ;
      RECT 40.311 4.714 40.397 4.862 ;
      RECT 40.225 4.718 40.311 4.863 ;
      RECT 40.176 4.72 40.225 4.865 ;
      RECT 40.09 4.72 40.176 4.867 ;
      RECT 40.05 4.715 40.09 4.869 ;
      RECT 40.04 4.709 40.05 4.87 ;
      RECT 40 4.704 40.04 4.867 ;
      RECT 39.99 4.697 40 4.863 ;
      RECT 39.975 4.693 39.99 4.861 ;
      RECT 39.958 4.689 39.975 4.859 ;
      RECT 39.872 4.679 39.958 4.851 ;
      RECT 39.786 4.661 39.872 4.837 ;
      RECT 39.7 4.644 39.786 4.823 ;
      RECT 39.675 4.632 39.7 4.814 ;
      RECT 39.605 4.622 39.675 4.807 ;
      RECT 39.56 4.61 39.605 4.798 ;
      RECT 39.5 4.597 39.56 4.79 ;
      RECT 39.495 4.589 39.5 4.785 ;
      RECT 39.46 4.584 39.495 4.783 ;
      RECT 39.405 4.575 39.46 4.776 ;
      RECT 39.365 4.564 39.405 4.768 ;
      RECT 39.35 4.557 39.365 4.764 ;
      RECT 39.33 4.55 39.345 4.761 ;
      RECT 39.315 4.54 39.33 4.759 ;
      RECT 39.3 4.527 39.315 4.756 ;
      RECT 39.275 4.51 39.3 4.752 ;
      RECT 39.26 4.492 39.275 4.749 ;
      RECT 39.235 4.445 39.26 4.747 ;
      RECT 39.211 4.445 39.235 4.744 ;
      RECT 39.125 4.445 39.211 4.736 ;
      RECT 39.085 4.445 39.125 4.728 ;
      RECT 38.95 4.492 38.98 4.76 ;
      RECT 40.63 4.075 40.89 4.335 ;
      RECT 40.59 4.075 40.89 4.213 ;
      RECT 40.555 4.075 40.89 4.198 ;
      RECT 40.5 4.075 40.89 4.178 ;
      RECT 40.42 3.885 40.7 4.165 ;
      RECT 40.42 4.067 40.77 4.165 ;
      RECT 40.42 4.01 40.755 4.165 ;
      RECT 40.42 3.957 40.705 4.165 ;
      RECT 37.58 4.244 37.595 4.7 ;
      RECT 37.575 4.316 37.681 4.698 ;
      RECT 37.595 3.41 37.73 4.696 ;
      RECT 37.58 4.26 37.735 4.695 ;
      RECT 37.58 4.31 37.74 4.693 ;
      RECT 37.565 4.375 37.74 4.692 ;
      RECT 37.575 4.367 37.745 4.689 ;
      RECT 37.555 4.415 37.745 4.684 ;
      RECT 37.555 4.415 37.76 4.681 ;
      RECT 37.55 4.415 37.76 4.678 ;
      RECT 37.525 4.415 37.785 4.675 ;
      RECT 37.595 3.41 37.755 4.063 ;
      RECT 37.59 3.41 37.755 4.035 ;
      RECT 37.585 3.41 37.755 3.863 ;
      RECT 37.585 3.41 37.775 3.803 ;
      RECT 37.54 3.41 37.8 3.67 ;
      RECT 37.02 3.885 37.3 4.165 ;
      RECT 37.01 3.9 37.3 4.16 ;
      RECT 36.965 3.962 37.3 4.158 ;
      RECT 37.04 3.877 37.205 4.165 ;
      RECT 37.04 3.862 37.161 4.165 ;
      RECT 37.075 3.855 37.161 4.165 ;
      RECT 36.54 5.005 36.82 5.285 ;
      RECT 36.5 4.967 36.795 5.078 ;
      RECT 36.485 4.917 36.775 4.973 ;
      RECT 36.43 4.68 36.69 4.94 ;
      RECT 36.43 4.882 36.77 4.94 ;
      RECT 36.43 4.822 36.765 4.94 ;
      RECT 36.43 4.772 36.745 4.94 ;
      RECT 36.43 4.752 36.74 4.94 ;
      RECT 36.43 4.73 36.735 4.94 ;
      RECT 36.43 4.715 36.705 4.94 ;
      RECT 32.15 8.66 32.47 8.98 ;
      RECT 32.18 8.13 32.35 8.98 ;
      RECT 32.18 8.13 32.355 8.48 ;
      RECT 32.18 8.13 33.155 8.305 ;
      RECT 32.98 3.26 33.155 8.305 ;
      RECT 32.925 3.26 33.275 3.61 ;
      RECT 32.95 9.09 33.275 9.415 ;
      RECT 31.835 9.18 33.275 9.35 ;
      RECT 31.835 3.69 31.995 9.35 ;
      RECT 32.15 3.66 32.47 3.98 ;
      RECT 31.835 3.69 32.47 3.86 ;
      RECT 30.515 2.435 30.89 2.805 ;
      RECT 22.425 2.255 22.8 2.625 ;
      RECT 20.99 2.255 21.365 2.625 ;
      RECT 20.99 2.375 30.82 2.545 ;
      RECT 25.11 5.655 30.79 5.825 ;
      RECT 30.62 4.72 30.79 5.825 ;
      RECT 24.92 4.895 24.955 5.825 ;
      RECT 25.185 5.005 25.215 5.285 ;
      RECT 24.89 4.895 24.955 5.155 ;
      RECT 30.53 4.725 30.88 5.075 ;
      RECT 24.72 3.52 24.755 3.78 ;
      RECT 24.495 3.52 24.555 3.78 ;
      RECT 25.175 4.985 25.185 5.285 ;
      RECT 25.17 4.945 25.175 5.285 ;
      RECT 25.155 4.9 25.17 5.285 ;
      RECT 25.15 4.865 25.155 5.285 ;
      RECT 25.145 4.845 25.15 5.285 ;
      RECT 25.115 4.772 25.145 5.285 ;
      RECT 25.11 4.7 25.115 5.285 ;
      RECT 25.095 4.66 25.11 5.825 ;
      RECT 25.085 4.6 25.095 5.825 ;
      RECT 25.04 4.54 25.085 5.825 ;
      RECT 24.955 4.501 25.04 5.825 ;
      RECT 24.95 4.492 24.955 4.865 ;
      RECT 24.94 4.491 24.95 4.848 ;
      RECT 24.915 4.472 24.94 4.818 ;
      RECT 24.91 4.447 24.915 4.797 ;
      RECT 24.9 4.425 24.91 4.788 ;
      RECT 24.895 4.396 24.9 4.778 ;
      RECT 24.855 4.322 24.895 4.75 ;
      RECT 24.835 4.223 24.855 4.715 ;
      RECT 24.82 4.159 24.835 4.698 ;
      RECT 24.79 4.083 24.82 4.67 ;
      RECT 24.77 3.998 24.79 4.643 ;
      RECT 24.73 3.894 24.77 4.55 ;
      RECT 24.725 3.815 24.73 4.458 ;
      RECT 24.72 3.798 24.725 4.435 ;
      RECT 24.715 3.52 24.72 4.415 ;
      RECT 24.685 3.52 24.715 4.353 ;
      RECT 24.68 3.52 24.685 4.285 ;
      RECT 24.67 3.52 24.68 4.25 ;
      RECT 24.66 3.52 24.67 4.215 ;
      RECT 24.595 3.52 24.66 4.07 ;
      RECT 24.59 3.52 24.595 3.94 ;
      RECT 24.56 3.52 24.59 3.873 ;
      RECT 24.555 3.52 24.56 3.798 ;
      RECT 28.89 3.455 29.15 3.715 ;
      RECT 28.885 3.455 29.15 3.663 ;
      RECT 28.88 3.455 29.15 3.633 ;
      RECT 28.855 3.325 29.135 3.605 ;
      RECT 16.705 9.43 16.995 9.78 ;
      RECT 16.705 9.49 18.015 9.66 ;
      RECT 17.845 9.12 18.015 9.66 ;
      RECT 28.345 9.04 28.695 9.39 ;
      RECT 17.845 9.12 28.695 9.29 ;
      RECT 27.895 5.005 28.175 5.285 ;
      RECT 27.935 4.96 28.2 5.22 ;
      RECT 27.925 4.995 28.2 5.22 ;
      RECT 27.93 4.98 28.175 5.285 ;
      RECT 27.935 4.957 28.145 5.285 ;
      RECT 27.935 4.955 28.13 5.285 ;
      RECT 27.975 4.945 28.13 5.285 ;
      RECT 27.945 4.95 28.13 5.285 ;
      RECT 27.975 4.942 28.075 5.285 ;
      RECT 28 4.935 28.075 5.285 ;
      RECT 27.98 4.937 28.075 5.285 ;
      RECT 27.31 4.45 27.57 4.71 ;
      RECT 27.36 4.442 27.55 4.71 ;
      RECT 27.365 4.362 27.55 4.71 ;
      RECT 27.485 3.75 27.55 4.71 ;
      RECT 27.39 4.147 27.55 4.71 ;
      RECT 27.465 3.835 27.55 4.71 ;
      RECT 27.5 3.46 27.636 4.188 ;
      RECT 27.445 3.957 27.636 4.188 ;
      RECT 27.46 3.897 27.55 4.71 ;
      RECT 27.5 3.46 27.66 3.853 ;
      RECT 27.5 3.46 27.67 3.75 ;
      RECT 27.49 3.46 27.75 3.72 ;
      RECT 26.895 5.005 27.175 5.285 ;
      RECT 26.915 4.965 27.175 5.285 ;
      RECT 26.555 4.92 26.66 5.18 ;
      RECT 26.41 3.41 26.5 3.67 ;
      RECT 26.95 4.475 26.955 4.515 ;
      RECT 26.945 4.465 26.95 4.6 ;
      RECT 26.94 4.455 26.945 4.693 ;
      RECT 26.93 4.435 26.94 4.749 ;
      RECT 26.85 4.363 26.93 4.829 ;
      RECT 26.885 5.007 26.895 5.232 ;
      RECT 26.88 5.004 26.885 5.227 ;
      RECT 26.865 5.001 26.88 5.22 ;
      RECT 26.83 4.995 26.865 5.202 ;
      RECT 26.845 4.298 26.85 4.903 ;
      RECT 26.825 4.249 26.845 4.918 ;
      RECT 26.815 4.982 26.83 5.185 ;
      RECT 26.82 4.191 26.825 4.933 ;
      RECT 26.815 4.169 26.82 4.943 ;
      RECT 26.78 4.079 26.815 5.18 ;
      RECT 26.765 3.957 26.78 5.18 ;
      RECT 26.76 3.91 26.765 5.18 ;
      RECT 26.735 3.835 26.76 5.18 ;
      RECT 26.72 3.75 26.735 5.18 ;
      RECT 26.715 3.697 26.72 5.18 ;
      RECT 26.71 3.677 26.715 5.18 ;
      RECT 26.705 3.652 26.71 4.414 ;
      RECT 26.69 4.612 26.71 5.18 ;
      RECT 26.7 3.63 26.705 4.391 ;
      RECT 26.69 3.582 26.7 4.356 ;
      RECT 26.685 3.545 26.69 4.322 ;
      RECT 26.685 4.692 26.69 5.18 ;
      RECT 26.67 3.522 26.685 4.277 ;
      RECT 26.665 4.79 26.685 5.18 ;
      RECT 26.615 3.41 26.67 4.119 ;
      RECT 26.66 4.912 26.665 5.18 ;
      RECT 26.6 3.41 26.615 3.958 ;
      RECT 26.595 3.41 26.6 3.91 ;
      RECT 26.59 3.41 26.595 3.898 ;
      RECT 26.545 3.41 26.59 3.835 ;
      RECT 26.52 3.41 26.545 3.753 ;
      RECT 26.505 3.41 26.52 3.705 ;
      RECT 26.5 3.41 26.505 3.675 ;
      RECT 25.825 4.86 25.87 5.12 ;
      RECT 25.73 3.395 25.875 3.655 ;
      RECT 26.235 4.017 26.245 4.108 ;
      RECT 26.22 3.955 26.235 4.164 ;
      RECT 26.215 3.902 26.22 4.21 ;
      RECT 26.165 3.849 26.215 4.336 ;
      RECT 26.16 3.804 26.165 4.483 ;
      RECT 26.15 3.792 26.16 4.525 ;
      RECT 26.115 3.756 26.15 4.63 ;
      RECT 26.11 3.724 26.115 4.736 ;
      RECT 26.095 3.706 26.11 4.781 ;
      RECT 26.09 3.689 26.095 4.015 ;
      RECT 26.085 4.07 26.095 4.838 ;
      RECT 26.08 3.675 26.09 3.988 ;
      RECT 26.075 4.125 26.085 5.12 ;
      RECT 26.07 3.661 26.08 3.973 ;
      RECT 26.07 4.175 26.075 5.12 ;
      RECT 26.055 3.638 26.07 3.953 ;
      RECT 26.035 4.297 26.07 5.12 ;
      RECT 26.05 3.62 26.055 3.935 ;
      RECT 26.045 3.612 26.05 3.925 ;
      RECT 26.015 3.58 26.045 3.889 ;
      RECT 26.025 4.425 26.035 5.12 ;
      RECT 26.02 4.452 26.025 5.12 ;
      RECT 26.015 4.502 26.02 5.12 ;
      RECT 26.005 3.546 26.015 3.854 ;
      RECT 25.965 4.57 26.015 5.12 ;
      RECT 25.99 3.523 26.005 3.83 ;
      RECT 25.965 3.395 25.99 3.793 ;
      RECT 25.96 3.395 25.965 3.765 ;
      RECT 25.93 4.67 25.965 5.12 ;
      RECT 25.955 3.395 25.96 3.758 ;
      RECT 25.95 3.395 25.955 3.748 ;
      RECT 25.935 3.395 25.95 3.733 ;
      RECT 25.92 3.395 25.935 3.705 ;
      RECT 25.885 4.775 25.93 5.12 ;
      RECT 25.905 3.395 25.92 3.678 ;
      RECT 25.875 3.395 25.905 3.663 ;
      RECT 25.87 4.847 25.885 5.12 ;
      RECT 25.795 3.93 25.835 4.19 ;
      RECT 25.57 3.877 25.575 4.135 ;
      RECT 21.525 3.355 21.785 3.615 ;
      RECT 21.525 3.38 21.8 3.595 ;
      RECT 23.915 3.205 23.92 3.35 ;
      RECT 25.785 3.925 25.795 4.19 ;
      RECT 25.765 3.917 25.785 4.19 ;
      RECT 25.747 3.913 25.765 4.19 ;
      RECT 25.661 3.902 25.747 4.19 ;
      RECT 25.575 3.885 25.661 4.19 ;
      RECT 25.52 3.872 25.57 4.12 ;
      RECT 25.486 3.864 25.52 4.095 ;
      RECT 25.4 3.853 25.486 4.06 ;
      RECT 25.365 3.83 25.4 4.025 ;
      RECT 25.355 3.792 25.365 4.011 ;
      RECT 25.35 3.765 25.355 4.007 ;
      RECT 25.345 3.752 25.35 4.004 ;
      RECT 25.335 3.732 25.345 4 ;
      RECT 25.33 3.707 25.335 3.996 ;
      RECT 25.305 3.662 25.33 3.99 ;
      RECT 25.295 3.603 25.305 3.982 ;
      RECT 25.285 3.571 25.295 3.973 ;
      RECT 25.265 3.523 25.285 3.953 ;
      RECT 25.26 3.483 25.265 3.923 ;
      RECT 25.245 3.457 25.26 3.897 ;
      RECT 25.24 3.435 25.245 3.873 ;
      RECT 25.225 3.407 25.24 3.849 ;
      RECT 25.21 3.38 25.225 3.813 ;
      RECT 25.195 3.357 25.21 3.775 ;
      RECT 25.19 3.347 25.195 3.75 ;
      RECT 25.18 3.34 25.19 3.733 ;
      RECT 25.165 3.327 25.18 3.703 ;
      RECT 25.16 3.317 25.165 3.678 ;
      RECT 25.155 3.312 25.16 3.665 ;
      RECT 25.145 3.305 25.155 3.645 ;
      RECT 25.14 3.298 25.145 3.63 ;
      RECT 25.115 3.291 25.14 3.588 ;
      RECT 25.1 3.281 25.115 3.538 ;
      RECT 25.09 3.276 25.1 3.508 ;
      RECT 25.08 3.272 25.09 3.483 ;
      RECT 25.065 3.269 25.08 3.473 ;
      RECT 25.015 3.266 25.065 3.458 ;
      RECT 24.995 3.264 25.015 3.443 ;
      RECT 24.946 3.262 24.995 3.438 ;
      RECT 24.86 3.258 24.946 3.433 ;
      RECT 24.821 3.255 24.86 3.429 ;
      RECT 24.735 3.251 24.821 3.424 ;
      RECT 24.685 3.248 24.735 3.418 ;
      RECT 24.636 3.245 24.685 3.413 ;
      RECT 24.55 3.242 24.636 3.408 ;
      RECT 24.546 3.24 24.55 3.405 ;
      RECT 24.46 3.237 24.546 3.4 ;
      RECT 24.411 3.233 24.46 3.393 ;
      RECT 24.325 3.23 24.411 3.388 ;
      RECT 24.301 3.227 24.325 3.384 ;
      RECT 24.215 3.225 24.301 3.379 ;
      RECT 24.15 3.221 24.215 3.372 ;
      RECT 24.147 3.22 24.15 3.369 ;
      RECT 24.061 3.217 24.147 3.366 ;
      RECT 23.975 3.211 24.061 3.359 ;
      RECT 23.945 3.207 23.975 3.355 ;
      RECT 23.92 3.205 23.945 3.353 ;
      RECT 23.865 3.202 23.915 3.35 ;
      RECT 23.785 3.201 23.865 3.35 ;
      RECT 23.73 3.203 23.785 3.353 ;
      RECT 23.715 3.204 23.73 3.357 ;
      RECT 23.66 3.212 23.715 3.367 ;
      RECT 23.63 3.22 23.66 3.38 ;
      RECT 23.611 3.221 23.63 3.386 ;
      RECT 23.525 3.224 23.611 3.391 ;
      RECT 23.455 3.229 23.525 3.4 ;
      RECT 23.436 3.232 23.455 3.406 ;
      RECT 23.35 3.236 23.436 3.411 ;
      RECT 23.31 3.24 23.35 3.418 ;
      RECT 23.301 3.242 23.31 3.421 ;
      RECT 23.215 3.246 23.301 3.426 ;
      RECT 23.212 3.249 23.215 3.43 ;
      RECT 23.126 3.252 23.212 3.434 ;
      RECT 23.04 3.258 23.126 3.442 ;
      RECT 23.016 3.262 23.04 3.446 ;
      RECT 22.93 3.266 23.016 3.451 ;
      RECT 22.885 3.271 22.93 3.458 ;
      RECT 22.805 3.276 22.885 3.465 ;
      RECT 22.725 3.282 22.805 3.48 ;
      RECT 22.7 3.286 22.725 3.493 ;
      RECT 22.635 3.289 22.7 3.505 ;
      RECT 22.58 3.294 22.635 3.52 ;
      RECT 22.55 3.297 22.58 3.538 ;
      RECT 22.54 3.299 22.55 3.551 ;
      RECT 22.48 3.314 22.54 3.561 ;
      RECT 22.465 3.331 22.48 3.57 ;
      RECT 22.46 3.34 22.465 3.57 ;
      RECT 22.45 3.35 22.46 3.57 ;
      RECT 22.44 3.367 22.45 3.57 ;
      RECT 22.42 3.377 22.44 3.571 ;
      RECT 22.375 3.387 22.42 3.572 ;
      RECT 22.34 3.396 22.375 3.574 ;
      RECT 22.275 3.401 22.34 3.576 ;
      RECT 22.195 3.402 22.275 3.579 ;
      RECT 22.191 3.4 22.195 3.58 ;
      RECT 22.105 3.397 22.191 3.582 ;
      RECT 22.058 3.394 22.105 3.584 ;
      RECT 21.972 3.39 22.058 3.587 ;
      RECT 21.886 3.386 21.972 3.59 ;
      RECT 21.8 3.382 21.886 3.594 ;
      RECT 23.735 4.445 24.015 4.725 ;
      RECT 23.775 4.425 24.035 4.685 ;
      RECT 23.765 4.435 24.035 4.685 ;
      RECT 23.775 4.362 23.99 4.725 ;
      RECT 23.83 4.285 23.985 4.725 ;
      RECT 23.835 4.07 23.985 4.725 ;
      RECT 23.825 3.872 23.975 4.123 ;
      RECT 23.815 3.872 23.975 3.99 ;
      RECT 23.81 3.75 23.97 3.893 ;
      RECT 23.795 3.75 23.97 3.798 ;
      RECT 23.79 3.46 23.965 3.775 ;
      RECT 23.775 3.46 23.965 3.745 ;
      RECT 23.735 3.46 23.995 3.72 ;
      RECT 23.645 4.93 23.725 5.19 ;
      RECT 23.05 3.65 23.055 3.915 ;
      RECT 22.93 3.65 23.055 3.91 ;
      RECT 23.605 4.895 23.645 5.19 ;
      RECT 23.56 4.817 23.605 5.19 ;
      RECT 23.54 4.745 23.56 5.19 ;
      RECT 23.53 4.697 23.54 5.19 ;
      RECT 23.495 4.63 23.53 5.19 ;
      RECT 23.465 4.53 23.495 5.19 ;
      RECT 23.445 4.455 23.465 4.99 ;
      RECT 23.435 4.405 23.445 4.945 ;
      RECT 23.43 4.382 23.435 4.918 ;
      RECT 23.425 4.367 23.43 4.905 ;
      RECT 23.42 4.352 23.425 4.883 ;
      RECT 23.415 4.337 23.42 4.865 ;
      RECT 23.39 4.292 23.415 4.82 ;
      RECT 23.38 4.24 23.39 4.763 ;
      RECT 23.37 4.21 23.38 4.73 ;
      RECT 23.36 4.175 23.37 4.698 ;
      RECT 23.325 4.107 23.36 4.63 ;
      RECT 23.32 4.046 23.325 4.565 ;
      RECT 23.31 4.034 23.32 4.545 ;
      RECT 23.305 4.022 23.31 4.525 ;
      RECT 23.3 4.014 23.305 4.513 ;
      RECT 23.295 4.006 23.3 4.493 ;
      RECT 23.285 3.994 23.295 4.465 ;
      RECT 23.275 3.978 23.285 4.435 ;
      RECT 23.25 3.95 23.275 4.373 ;
      RECT 23.24 3.921 23.25 4.318 ;
      RECT 23.225 3.9 23.24 4.278 ;
      RECT 23.22 3.884 23.225 4.25 ;
      RECT 23.215 3.872 23.22 4.24 ;
      RECT 23.21 3.867 23.215 4.213 ;
      RECT 23.205 3.86 23.21 4.2 ;
      RECT 23.19 3.843 23.205 4.173 ;
      RECT 23.18 3.65 23.19 4.133 ;
      RECT 23.17 3.65 23.18 4.1 ;
      RECT 23.16 3.65 23.17 4.075 ;
      RECT 23.09 3.65 23.16 4.01 ;
      RECT 23.08 3.65 23.09 3.958 ;
      RECT 23.065 3.65 23.08 3.94 ;
      RECT 23.055 3.65 23.065 3.925 ;
      RECT 22.885 4.52 23.145 4.78 ;
      RECT 21.42 4.555 21.425 4.762 ;
      RECT 21.055 4.445 21.13 4.76 ;
      RECT 20.87 4.5 21.025 4.76 ;
      RECT 21.055 4.445 21.16 4.725 ;
      RECT 22.87 4.617 22.885 4.778 ;
      RECT 22.845 4.625 22.87 4.783 ;
      RECT 22.82 4.632 22.845 4.788 ;
      RECT 22.757 4.643 22.82 4.797 ;
      RECT 22.671 4.662 22.757 4.814 ;
      RECT 22.585 4.684 22.671 4.833 ;
      RECT 22.57 4.697 22.585 4.844 ;
      RECT 22.53 4.705 22.57 4.851 ;
      RECT 22.51 4.71 22.53 4.858 ;
      RECT 22.472 4.711 22.51 4.861 ;
      RECT 22.386 4.714 22.472 4.862 ;
      RECT 22.3 4.718 22.386 4.863 ;
      RECT 22.251 4.72 22.3 4.865 ;
      RECT 22.165 4.72 22.251 4.867 ;
      RECT 22.125 4.715 22.165 4.869 ;
      RECT 22.115 4.709 22.125 4.87 ;
      RECT 22.075 4.704 22.115 4.867 ;
      RECT 22.065 4.697 22.075 4.863 ;
      RECT 22.05 4.693 22.065 4.861 ;
      RECT 22.033 4.689 22.05 4.859 ;
      RECT 21.947 4.679 22.033 4.851 ;
      RECT 21.861 4.661 21.947 4.837 ;
      RECT 21.775 4.644 21.861 4.823 ;
      RECT 21.75 4.632 21.775 4.814 ;
      RECT 21.68 4.622 21.75 4.807 ;
      RECT 21.635 4.61 21.68 4.798 ;
      RECT 21.575 4.597 21.635 4.79 ;
      RECT 21.57 4.589 21.575 4.785 ;
      RECT 21.535 4.584 21.57 4.783 ;
      RECT 21.48 4.575 21.535 4.776 ;
      RECT 21.44 4.564 21.48 4.768 ;
      RECT 21.425 4.557 21.44 4.764 ;
      RECT 21.405 4.55 21.42 4.761 ;
      RECT 21.39 4.54 21.405 4.759 ;
      RECT 21.375 4.527 21.39 4.756 ;
      RECT 21.35 4.51 21.375 4.752 ;
      RECT 21.335 4.492 21.35 4.749 ;
      RECT 21.31 4.445 21.335 4.747 ;
      RECT 21.286 4.445 21.31 4.744 ;
      RECT 21.2 4.445 21.286 4.736 ;
      RECT 21.16 4.445 21.2 4.728 ;
      RECT 21.025 4.492 21.055 4.76 ;
      RECT 22.705 4.075 22.965 4.335 ;
      RECT 22.665 4.075 22.965 4.213 ;
      RECT 22.63 4.075 22.965 4.198 ;
      RECT 22.575 4.075 22.965 4.178 ;
      RECT 22.495 3.885 22.775 4.165 ;
      RECT 22.495 4.067 22.845 4.165 ;
      RECT 22.495 4.01 22.83 4.165 ;
      RECT 22.495 3.957 22.78 4.165 ;
      RECT 19.655 4.244 19.67 4.7 ;
      RECT 19.65 4.316 19.756 4.698 ;
      RECT 19.67 3.41 19.805 4.696 ;
      RECT 19.655 4.26 19.81 4.695 ;
      RECT 19.655 4.31 19.815 4.693 ;
      RECT 19.64 4.375 19.815 4.692 ;
      RECT 19.65 4.367 19.82 4.689 ;
      RECT 19.63 4.415 19.82 4.684 ;
      RECT 19.63 4.415 19.835 4.681 ;
      RECT 19.625 4.415 19.835 4.678 ;
      RECT 19.6 4.415 19.86 4.675 ;
      RECT 19.67 3.41 19.83 4.063 ;
      RECT 19.665 3.41 19.83 4.035 ;
      RECT 19.66 3.41 19.83 3.863 ;
      RECT 19.66 3.41 19.85 3.803 ;
      RECT 19.615 3.41 19.875 3.67 ;
      RECT 19.095 3.885 19.375 4.165 ;
      RECT 19.085 3.9 19.375 4.16 ;
      RECT 19.04 3.962 19.375 4.158 ;
      RECT 19.115 3.877 19.28 4.165 ;
      RECT 19.115 3.862 19.236 4.165 ;
      RECT 19.15 3.855 19.236 4.165 ;
      RECT 18.615 5.005 18.895 5.285 ;
      RECT 18.575 4.967 18.87 5.078 ;
      RECT 18.56 4.917 18.85 4.973 ;
      RECT 18.505 4.68 18.765 4.94 ;
      RECT 18.505 4.882 18.845 4.94 ;
      RECT 18.505 4.822 18.84 4.94 ;
      RECT 18.505 4.772 18.82 4.94 ;
      RECT 18.505 4.752 18.815 4.94 ;
      RECT 18.505 4.73 18.81 4.94 ;
      RECT 18.505 4.715 18.78 4.94 ;
      RECT 106.94 7.35 107.315 7.73 ;
      RECT 99.385 9.49 99.76 9.86 ;
      RECT 90.72 2.225 91.095 2.595 ;
      RECT 89.015 7.35 89.39 7.73 ;
      RECT 81.46 9.49 81.835 9.86 ;
      RECT 72.795 2.225 73.17 2.595 ;
      RECT 71.09 7.35 71.465 7.73 ;
      RECT 63.535 9.49 63.91 9.86 ;
      RECT 54.87 2.225 55.245 2.595 ;
      RECT 53.165 7.35 53.54 7.73 ;
      RECT 45.61 9.49 45.985 9.86 ;
      RECT 36.945 2.225 37.32 2.595 ;
      RECT 35.24 7.35 35.615 7.73 ;
      RECT 27.685 9.49 28.06 9.86 ;
      RECT 19.02 2.225 19.395 2.595 ;
    LAYER via1 ;
      RECT 107.105 9.81 107.255 9.96 ;
      RECT 107.05 7.465 107.2 7.615 ;
      RECT 104.74 9.175 104.89 9.325 ;
      RECT 104.725 3.36 104.875 3.51 ;
      RECT 103.935 3.745 104.085 3.895 ;
      RECT 103.935 8.76 104.085 8.91 ;
      RECT 102.33 2.545 102.48 2.695 ;
      RECT 102.33 4.825 102.48 4.975 ;
      RECT 100.645 3.51 100.795 3.66 ;
      RECT 100.405 9.15 100.555 9.3 ;
      RECT 99.695 5.015 99.845 5.165 ;
      RECT 99.5 9.6 99.65 9.75 ;
      RECT 99.245 3.515 99.395 3.665 ;
      RECT 99.065 4.505 99.215 4.655 ;
      RECT 98.67 5.02 98.82 5.17 ;
      RECT 98.31 4.975 98.46 5.125 ;
      RECT 98.165 3.465 98.315 3.615 ;
      RECT 97.58 4.915 97.73 5.065 ;
      RECT 97.485 3.45 97.635 3.6 ;
      RECT 97.33 3.985 97.48 4.135 ;
      RECT 96.645 4.95 96.795 5.1 ;
      RECT 96.25 3.575 96.4 3.725 ;
      RECT 95.53 4.48 95.68 4.63 ;
      RECT 95.49 3.515 95.64 3.665 ;
      RECT 95.22 4.985 95.37 5.135 ;
      RECT 94.685 3.705 94.835 3.855 ;
      RECT 94.64 4.575 94.79 4.725 ;
      RECT 94.46 4.13 94.61 4.28 ;
      RECT 93.28 3.41 93.43 3.56 ;
      RECT 92.625 4.555 92.775 4.705 ;
      RECT 91.37 3.465 91.52 3.615 ;
      RECT 91.355 4.47 91.505 4.62 ;
      RECT 90.84 3.955 90.99 4.105 ;
      RECT 90.26 4.735 90.41 4.885 ;
      RECT 89.16 9.195 89.31 9.345 ;
      RECT 89.125 7.465 89.275 7.615 ;
      RECT 86.815 9.175 86.965 9.325 ;
      RECT 86.8 3.36 86.95 3.51 ;
      RECT 86.01 3.745 86.16 3.895 ;
      RECT 86.01 8.76 86.16 8.91 ;
      RECT 84.405 2.545 84.555 2.695 ;
      RECT 84.405 4.825 84.555 4.975 ;
      RECT 82.72 3.51 82.87 3.66 ;
      RECT 82.2 9.15 82.35 9.3 ;
      RECT 81.77 5.015 81.92 5.165 ;
      RECT 81.575 9.6 81.725 9.75 ;
      RECT 81.32 3.515 81.47 3.665 ;
      RECT 81.14 4.505 81.29 4.655 ;
      RECT 80.745 5.02 80.895 5.17 ;
      RECT 80.385 4.975 80.535 5.125 ;
      RECT 80.24 3.465 80.39 3.615 ;
      RECT 79.655 4.915 79.805 5.065 ;
      RECT 79.56 3.45 79.71 3.6 ;
      RECT 79.405 3.985 79.555 4.135 ;
      RECT 78.72 4.95 78.87 5.1 ;
      RECT 78.325 3.575 78.475 3.725 ;
      RECT 77.605 4.48 77.755 4.63 ;
      RECT 77.565 3.515 77.715 3.665 ;
      RECT 77.295 4.985 77.445 5.135 ;
      RECT 76.76 3.705 76.91 3.855 ;
      RECT 76.715 4.575 76.865 4.725 ;
      RECT 76.535 4.13 76.685 4.28 ;
      RECT 75.355 3.41 75.505 3.56 ;
      RECT 74.7 4.555 74.85 4.705 ;
      RECT 73.445 3.465 73.595 3.615 ;
      RECT 73.43 4.47 73.58 4.62 ;
      RECT 72.915 3.955 73.065 4.105 ;
      RECT 72.335 4.735 72.485 4.885 ;
      RECT 71.235 9.195 71.385 9.345 ;
      RECT 71.2 7.465 71.35 7.615 ;
      RECT 68.89 9.175 69.04 9.325 ;
      RECT 68.875 3.36 69.025 3.51 ;
      RECT 68.085 3.745 68.235 3.895 ;
      RECT 68.085 8.76 68.235 8.91 ;
      RECT 66.48 2.545 66.63 2.695 ;
      RECT 66.48 4.825 66.63 4.975 ;
      RECT 64.795 3.51 64.945 3.66 ;
      RECT 64.33 9.15 64.48 9.3 ;
      RECT 63.845 5.015 63.995 5.165 ;
      RECT 63.65 9.6 63.8 9.75 ;
      RECT 63.395 3.515 63.545 3.665 ;
      RECT 63.215 4.505 63.365 4.655 ;
      RECT 62.82 5.02 62.97 5.17 ;
      RECT 62.46 4.975 62.61 5.125 ;
      RECT 62.315 3.465 62.465 3.615 ;
      RECT 61.73 4.915 61.88 5.065 ;
      RECT 61.635 3.45 61.785 3.6 ;
      RECT 61.48 3.985 61.63 4.135 ;
      RECT 60.795 4.95 60.945 5.1 ;
      RECT 60.4 3.575 60.55 3.725 ;
      RECT 59.68 4.48 59.83 4.63 ;
      RECT 59.64 3.515 59.79 3.665 ;
      RECT 59.37 4.985 59.52 5.135 ;
      RECT 58.835 3.705 58.985 3.855 ;
      RECT 58.79 4.575 58.94 4.725 ;
      RECT 58.61 4.13 58.76 4.28 ;
      RECT 57.43 3.41 57.58 3.56 ;
      RECT 56.775 4.555 56.925 4.705 ;
      RECT 55.52 3.465 55.67 3.615 ;
      RECT 55.505 4.47 55.655 4.62 ;
      RECT 54.99 3.955 55.14 4.105 ;
      RECT 54.41 4.735 54.56 4.885 ;
      RECT 53.355 9.195 53.505 9.345 ;
      RECT 53.275 7.465 53.425 7.615 ;
      RECT 50.965 9.175 51.115 9.325 ;
      RECT 50.95 3.36 51.1 3.51 ;
      RECT 50.16 3.745 50.31 3.895 ;
      RECT 50.16 8.76 50.31 8.91 ;
      RECT 48.555 2.545 48.705 2.695 ;
      RECT 48.555 4.825 48.705 4.975 ;
      RECT 46.87 3.51 47.02 3.66 ;
      RECT 46.4 9.15 46.55 9.3 ;
      RECT 45.92 5.015 46.07 5.165 ;
      RECT 45.725 9.6 45.875 9.75 ;
      RECT 45.47 3.515 45.62 3.665 ;
      RECT 45.29 4.505 45.44 4.655 ;
      RECT 44.895 5.02 45.045 5.17 ;
      RECT 44.535 4.975 44.685 5.125 ;
      RECT 44.39 3.465 44.54 3.615 ;
      RECT 43.805 4.915 43.955 5.065 ;
      RECT 43.71 3.45 43.86 3.6 ;
      RECT 43.555 3.985 43.705 4.135 ;
      RECT 42.87 4.95 43.02 5.1 ;
      RECT 42.475 3.575 42.625 3.725 ;
      RECT 41.755 4.48 41.905 4.63 ;
      RECT 41.715 3.515 41.865 3.665 ;
      RECT 41.445 4.985 41.595 5.135 ;
      RECT 40.91 3.705 41.06 3.855 ;
      RECT 40.865 4.575 41.015 4.725 ;
      RECT 40.685 4.13 40.835 4.28 ;
      RECT 39.505 3.41 39.655 3.56 ;
      RECT 38.85 4.555 39 4.705 ;
      RECT 37.595 3.465 37.745 3.615 ;
      RECT 37.58 4.47 37.73 4.62 ;
      RECT 37.065 3.955 37.215 4.105 ;
      RECT 36.485 4.735 36.635 4.885 ;
      RECT 35.43 9.195 35.58 9.345 ;
      RECT 35.35 7.465 35.5 7.615 ;
      RECT 33.04 9.175 33.19 9.325 ;
      RECT 33.025 3.36 33.175 3.51 ;
      RECT 32.235 3.745 32.385 3.895 ;
      RECT 32.235 8.76 32.385 8.91 ;
      RECT 30.63 2.545 30.78 2.695 ;
      RECT 30.63 4.825 30.78 4.975 ;
      RECT 28.945 3.51 29.095 3.66 ;
      RECT 28.445 9.14 28.595 9.29 ;
      RECT 27.995 5.015 28.145 5.165 ;
      RECT 27.8 9.6 27.95 9.75 ;
      RECT 27.545 3.515 27.695 3.665 ;
      RECT 27.365 4.505 27.515 4.655 ;
      RECT 26.97 5.02 27.12 5.17 ;
      RECT 26.61 4.975 26.76 5.125 ;
      RECT 26.465 3.465 26.615 3.615 ;
      RECT 25.88 4.915 26.03 5.065 ;
      RECT 25.785 3.45 25.935 3.6 ;
      RECT 25.63 3.985 25.78 4.135 ;
      RECT 24.945 4.95 25.095 5.1 ;
      RECT 24.55 3.575 24.7 3.725 ;
      RECT 23.83 4.48 23.98 4.63 ;
      RECT 23.79 3.515 23.94 3.665 ;
      RECT 23.52 4.985 23.67 5.135 ;
      RECT 22.985 3.705 23.135 3.855 ;
      RECT 22.94 4.575 23.09 4.725 ;
      RECT 22.76 4.13 22.91 4.28 ;
      RECT 21.58 3.41 21.73 3.56 ;
      RECT 20.925 4.555 21.075 4.705 ;
      RECT 19.67 3.465 19.82 3.615 ;
      RECT 19.655 4.47 19.805 4.62 ;
      RECT 19.14 3.955 19.29 4.105 ;
      RECT 18.56 4.735 18.71 4.885 ;
      RECT 16.775 9.53 16.925 9.68 ;
      RECT 16.4 8.79 16.55 8.94 ;
    LAYER met1 ;
      RECT 106.975 10.205 107.27 10.435 ;
      RECT 107.035 9.71 107.21 10.435 ;
      RECT 107.005 9.71 107.355 10.06 ;
      RECT 107.035 8.725 107.205 10.435 ;
      RECT 106.975 8.725 107.265 8.955 ;
      RECT 105.985 10.205 106.28 10.435 ;
      RECT 106.045 8.725 106.215 10.435 ;
      RECT 105.985 8.725 106.275 8.955 ;
      RECT 105.985 8.76 106.835 8.92 ;
      RECT 106.67 8.355 106.835 8.92 ;
      RECT 105.985 8.755 106.38 8.92 ;
      RECT 106.605 8.355 106.895 8.585 ;
      RECT 106.605 8.385 107.065 8.555 ;
      RECT 106.57 4.025 106.895 4.26 ;
      RECT 106.57 4.055 107.06 4.225 ;
      RECT 106.57 3.69 106.76 4.26 ;
      RECT 105.985 3.655 106.275 3.885 ;
      RECT 105.985 3.69 106.76 3.86 ;
      RECT 106.045 2.175 106.215 3.885 ;
      RECT 105.985 2.175 106.28 2.405 ;
      RECT 105.615 4.025 105.905 4.255 ;
      RECT 105.615 4.055 106.075 4.225 ;
      RECT 105.68 2.95 105.845 4.255 ;
      RECT 104.195 2.915 104.485 3.145 ;
      RECT 104.195 2.95 105.845 3.12 ;
      RECT 104.255 2.175 104.425 3.145 ;
      RECT 104.195 2.175 104.485 2.405 ;
      RECT 104.195 10.205 104.485 10.435 ;
      RECT 104.255 9.465 104.425 10.435 ;
      RECT 104.255 9.555 105.845 9.725 ;
      RECT 105.675 8.355 105.845 9.725 ;
      RECT 104.195 9.465 104.485 9.695 ;
      RECT 105.615 8.355 105.905 8.585 ;
      RECT 105.615 8.385 106.075 8.555 ;
      RECT 102.23 4.725 102.58 5.075 ;
      RECT 102.32 3.32 102.49 5.075 ;
      RECT 104.625 3.26 104.975 3.61 ;
      RECT 102.32 3.32 103.94 3.495 ;
      RECT 102.32 3.32 104.595 3.49 ;
      RECT 104.455 3.315 104.975 3.485 ;
      RECT 104.65 9.09 104.975 9.415 ;
      RECT 100.305 9.05 100.655 9.4 ;
      RECT 104.625 9.095 104.975 9.325 ;
      RECT 99.865 9.095 100.155 9.325 ;
      RECT 104.455 9.12 104.975 9.295 ;
      RECT 99.695 9.125 100.155 9.295 ;
      RECT 99.865 9.12 104.975 9.29 ;
      RECT 103.85 3.66 104.17 3.98 ;
      RECT 103.825 3.655 104.115 3.885 ;
      RECT 103.78 3.685 104.17 3.86 ;
      RECT 103.65 3.685 104.17 3.855 ;
      RECT 103.85 8.66 104.17 8.98 ;
      RECT 103.825 8.725 104.17 8.955 ;
      RECT 103.65 8.755 104.17 8.925 ;
      RECT 99.64 4.96 99.68 5.22 ;
      RECT 99.68 4.94 99.685 4.95 ;
      RECT 101.01 4.185 101.02 4.406 ;
      RECT 100.94 4.18 101.01 4.531 ;
      RECT 100.93 4.18 100.94 4.658 ;
      RECT 100.905 4.18 100.93 4.705 ;
      RECT 100.88 4.18 100.905 4.783 ;
      RECT 100.86 4.18 100.88 4.853 ;
      RECT 100.835 4.18 100.86 4.893 ;
      RECT 100.825 4.18 100.835 4.913 ;
      RECT 100.815 4.182 100.825 4.921 ;
      RECT 100.81 4.187 100.815 4.378 ;
      RECT 100.81 4.387 100.815 4.922 ;
      RECT 100.805 4.432 100.81 4.923 ;
      RECT 100.795 4.497 100.805 4.924 ;
      RECT 100.785 4.592 100.795 4.926 ;
      RECT 100.78 4.645 100.785 4.928 ;
      RECT 100.775 4.665 100.78 4.929 ;
      RECT 100.72 4.69 100.775 4.935 ;
      RECT 100.68 4.725 100.72 4.944 ;
      RECT 100.67 4.742 100.68 4.949 ;
      RECT 100.661 4.748 100.67 4.951 ;
      RECT 100.575 4.786 100.661 4.962 ;
      RECT 100.57 4.825 100.575 4.972 ;
      RECT 100.495 4.832 100.57 4.982 ;
      RECT 100.475 4.842 100.495 4.993 ;
      RECT 100.445 4.849 100.475 5.001 ;
      RECT 100.42 4.856 100.445 5.008 ;
      RECT 100.396 4.862 100.42 5.013 ;
      RECT 100.31 4.875 100.396 5.025 ;
      RECT 100.232 4.882 100.31 5.043 ;
      RECT 100.146 4.877 100.232 5.061 ;
      RECT 100.06 4.872 100.146 5.081 ;
      RECT 99.98 4.866 100.06 5.098 ;
      RECT 99.915 4.862 99.98 5.127 ;
      RECT 99.91 4.576 99.915 4.6 ;
      RECT 99.9 4.852 99.915 5.155 ;
      RECT 99.905 4.57 99.91 4.64 ;
      RECT 99.9 4.564 99.905 4.71 ;
      RECT 99.895 4.558 99.9 4.788 ;
      RECT 99.895 4.835 99.9 5.22 ;
      RECT 99.887 4.555 99.895 5.22 ;
      RECT 99.801 4.553 99.887 5.22 ;
      RECT 99.715 4.551 99.801 5.22 ;
      RECT 99.705 4.552 99.715 5.22 ;
      RECT 99.7 4.557 99.705 5.22 ;
      RECT 99.69 4.57 99.7 5.22 ;
      RECT 99.685 4.592 99.69 5.22 ;
      RECT 99.68 4.952 99.685 5.22 ;
      RECT 100.31 4.42 100.315 4.64 ;
      RECT 100.815 3.455 100.85 3.715 ;
      RECT 100.8 3.455 100.815 3.723 ;
      RECT 100.771 3.455 100.8 3.745 ;
      RECT 100.685 3.455 100.771 3.805 ;
      RECT 100.665 3.455 100.685 3.87 ;
      RECT 100.605 3.455 100.665 4.035 ;
      RECT 100.6 3.455 100.605 4.183 ;
      RECT 100.595 3.455 100.6 4.195 ;
      RECT 100.59 3.455 100.595 4.221 ;
      RECT 100.56 3.641 100.59 4.301 ;
      RECT 100.555 3.689 100.56 4.39 ;
      RECT 100.55 3.703 100.555 4.405 ;
      RECT 100.545 3.722 100.55 4.435 ;
      RECT 100.54 3.737 100.545 4.451 ;
      RECT 100.535 3.752 100.54 4.473 ;
      RECT 100.53 3.772 100.535 4.495 ;
      RECT 100.52 3.792 100.53 4.528 ;
      RECT 100.505 3.834 100.52 4.59 ;
      RECT 100.5 3.865 100.505 4.63 ;
      RECT 100.495 3.877 100.5 4.635 ;
      RECT 100.49 3.889 100.495 4.64 ;
      RECT 100.485 3.902 100.49 4.64 ;
      RECT 100.48 3.92 100.485 4.64 ;
      RECT 100.475 3.94 100.48 4.64 ;
      RECT 100.47 3.952 100.475 4.64 ;
      RECT 100.465 3.965 100.47 4.64 ;
      RECT 100.445 4 100.465 4.64 ;
      RECT 100.395 4.102 100.445 4.64 ;
      RECT 100.39 4.187 100.395 4.64 ;
      RECT 100.385 4.195 100.39 4.64 ;
      RECT 100.38 4.212 100.385 4.64 ;
      RECT 100.375 4.227 100.38 4.64 ;
      RECT 100.34 4.292 100.375 4.64 ;
      RECT 100.325 4.357 100.34 4.64 ;
      RECT 100.32 4.387 100.325 4.64 ;
      RECT 100.315 4.412 100.32 4.64 ;
      RECT 100.3 4.422 100.31 4.64 ;
      RECT 100.285 4.435 100.3 4.633 ;
      RECT 100.03 4.025 100.1 4.235 ;
      RECT 99.82 4.002 99.825 4.195 ;
      RECT 97.275 3.93 97.535 4.19 ;
      RECT 100.11 4.212 100.115 4.215 ;
      RECT 100.1 4.03 100.11 4.23 ;
      RECT 100.001 4.023 100.03 4.235 ;
      RECT 99.915 4.015 100.001 4.235 ;
      RECT 99.9 4.009 99.915 4.233 ;
      RECT 99.88 4.008 99.9 4.22 ;
      RECT 99.875 4.007 99.88 4.203 ;
      RECT 99.825 4.004 99.875 4.198 ;
      RECT 99.795 4.001 99.82 4.193 ;
      RECT 99.775 3.999 99.795 4.188 ;
      RECT 99.76 3.997 99.775 4.185 ;
      RECT 99.73 3.995 99.76 4.183 ;
      RECT 99.665 3.991 99.73 4.175 ;
      RECT 99.635 3.986 99.665 4.17 ;
      RECT 99.615 3.984 99.635 4.168 ;
      RECT 99.585 3.981 99.615 4.163 ;
      RECT 99.525 3.977 99.585 4.155 ;
      RECT 99.52 3.974 99.525 4.15 ;
      RECT 99.45 3.972 99.52 4.145 ;
      RECT 99.421 3.968 99.45 4.138 ;
      RECT 99.335 3.963 99.421 4.13 ;
      RECT 99.301 3.958 99.335 4.122 ;
      RECT 99.215 3.95 99.301 4.114 ;
      RECT 99.176 3.943 99.215 4.106 ;
      RECT 99.09 3.938 99.176 4.098 ;
      RECT 99.025 3.932 99.09 4.088 ;
      RECT 99.005 3.927 99.025 4.083 ;
      RECT 98.996 3.924 99.005 4.082 ;
      RECT 98.91 3.92 98.996 4.076 ;
      RECT 98.87 3.916 98.91 4.068 ;
      RECT 98.85 3.912 98.87 4.066 ;
      RECT 98.79 3.912 98.85 4.063 ;
      RECT 98.77 3.915 98.79 4.061 ;
      RECT 98.749 3.915 98.77 4.061 ;
      RECT 98.663 3.917 98.749 4.065 ;
      RECT 98.577 3.919 98.663 4.071 ;
      RECT 98.491 3.921 98.577 4.078 ;
      RECT 98.405 3.924 98.491 4.084 ;
      RECT 98.371 3.925 98.405 4.089 ;
      RECT 98.285 3.928 98.371 4.094 ;
      RECT 98.256 3.935 98.285 4.099 ;
      RECT 98.17 3.935 98.256 4.104 ;
      RECT 98.137 3.935 98.17 4.109 ;
      RECT 98.051 3.937 98.137 4.114 ;
      RECT 97.965 3.939 98.051 4.121 ;
      RECT 97.901 3.941 97.965 4.127 ;
      RECT 97.815 3.943 97.901 4.133 ;
      RECT 97.812 3.945 97.815 4.136 ;
      RECT 97.726 3.946 97.812 4.14 ;
      RECT 97.64 3.949 97.726 4.147 ;
      RECT 97.621 3.951 97.64 4.151 ;
      RECT 97.535 3.953 97.621 4.156 ;
      RECT 97.265 3.965 97.275 4.16 ;
      RECT 99.435 10.205 99.725 10.435 ;
      RECT 99.495 9.465 99.665 10.435 ;
      RECT 99.385 9.49 99.76 9.86 ;
      RECT 99.435 9.465 99.725 9.86 ;
      RECT 99.5 3.545 99.685 3.755 ;
      RECT 99.495 3.546 99.69 3.753 ;
      RECT 99.49 3.551 99.7 3.748 ;
      RECT 99.485 3.527 99.49 3.745 ;
      RECT 99.455 3.524 99.485 3.738 ;
      RECT 99.45 3.52 99.455 3.729 ;
      RECT 99.415 3.551 99.7 3.724 ;
      RECT 99.19 3.46 99.45 3.72 ;
      RECT 99.49 3.529 99.495 3.748 ;
      RECT 99.495 3.53 99.5 3.753 ;
      RECT 99.19 3.542 99.57 3.72 ;
      RECT 99.19 3.54 99.555 3.72 ;
      RECT 99.19 3.535 99.545 3.72 ;
      RECT 99.145 4.45 99.195 4.735 ;
      RECT 99.09 4.42 99.095 4.735 ;
      RECT 99.06 4.4 99.065 4.735 ;
      RECT 99.21 4.45 99.27 4.71 ;
      RECT 99.205 4.45 99.21 4.718 ;
      RECT 99.195 4.45 99.205 4.73 ;
      RECT 99.11 4.44 99.145 4.735 ;
      RECT 99.105 4.427 99.11 4.735 ;
      RECT 99.095 4.422 99.105 4.735 ;
      RECT 99.075 4.412 99.09 4.735 ;
      RECT 99.065 4.405 99.075 4.735 ;
      RECT 99.055 4.397 99.06 4.735 ;
      RECT 99.025 4.387 99.055 4.735 ;
      RECT 99.01 4.375 99.025 4.735 ;
      RECT 98.995 4.365 99.01 4.73 ;
      RECT 98.975 4.355 98.995 4.705 ;
      RECT 98.965 4.347 98.975 4.682 ;
      RECT 98.935 4.33 98.965 4.672 ;
      RECT 98.93 4.307 98.935 4.663 ;
      RECT 98.925 4.294 98.93 4.661 ;
      RECT 98.91 4.27 98.925 4.655 ;
      RECT 98.905 4.246 98.91 4.649 ;
      RECT 98.895 4.235 98.905 4.644 ;
      RECT 98.89 4.225 98.895 4.64 ;
      RECT 98.885 4.217 98.89 4.637 ;
      RECT 98.875 4.212 98.885 4.633 ;
      RECT 98.87 4.207 98.875 4.629 ;
      RECT 98.785 4.205 98.87 4.604 ;
      RECT 98.755 4.205 98.785 4.57 ;
      RECT 98.74 4.205 98.755 4.553 ;
      RECT 98.685 4.205 98.74 4.498 ;
      RECT 98.68 4.21 98.685 4.447 ;
      RECT 98.67 4.215 98.68 4.437 ;
      RECT 98.665 4.225 98.67 4.423 ;
      RECT 98.615 4.965 98.875 5.225 ;
      RECT 98.535 4.98 98.875 5.201 ;
      RECT 98.515 4.98 98.875 5.196 ;
      RECT 98.491 4.98 98.875 5.194 ;
      RECT 98.405 4.98 98.875 5.189 ;
      RECT 98.255 4.92 98.515 5.185 ;
      RECT 98.21 4.98 98.875 5.18 ;
      RECT 98.205 4.987 98.875 5.175 ;
      RECT 98.22 4.975 98.535 5.185 ;
      RECT 98.11 3.41 98.37 3.67 ;
      RECT 98.11 3.467 98.375 3.663 ;
      RECT 98.11 3.497 98.38 3.595 ;
      RECT 98.17 3.928 98.285 3.93 ;
      RECT 98.256 3.925 98.285 3.93 ;
      RECT 97.28 4.929 97.305 5.169 ;
      RECT 97.265 4.932 97.355 5.163 ;
      RECT 97.26 4.937 97.441 5.158 ;
      RECT 97.255 4.945 97.505 5.156 ;
      RECT 97.255 4.945 97.515 5.155 ;
      RECT 97.25 4.952 97.525 5.148 ;
      RECT 97.25 4.952 97.611 5.137 ;
      RECT 97.245 4.987 97.611 5.133 ;
      RECT 97.245 4.987 97.62 5.122 ;
      RECT 97.525 4.86 97.785 5.12 ;
      RECT 97.235 5.037 97.785 5.118 ;
      RECT 97.505 4.905 97.525 5.153 ;
      RECT 97.441 4.908 97.505 5.157 ;
      RECT 97.355 4.913 97.441 5.162 ;
      RECT 97.285 4.924 97.785 5.12 ;
      RECT 97.305 4.918 97.355 5.167 ;
      RECT 97.43 3.395 97.44 3.657 ;
      RECT 97.42 3.452 97.43 3.66 ;
      RECT 97.395 3.457 97.42 3.666 ;
      RECT 97.37 3.461 97.395 3.678 ;
      RECT 97.36 3.464 97.37 3.688 ;
      RECT 97.355 3.465 97.36 3.693 ;
      RECT 97.35 3.466 97.355 3.698 ;
      RECT 97.345 3.467 97.35 3.7 ;
      RECT 97.32 3.47 97.345 3.703 ;
      RECT 97.29 3.476 97.32 3.706 ;
      RECT 97.225 3.487 97.29 3.709 ;
      RECT 97.18 3.495 97.225 3.713 ;
      RECT 97.165 3.495 97.18 3.721 ;
      RECT 97.16 3.496 97.165 3.728 ;
      RECT 97.155 3.498 97.16 3.731 ;
      RECT 97.15 3.502 97.155 3.734 ;
      RECT 97.14 3.51 97.15 3.738 ;
      RECT 97.135 3.523 97.14 3.743 ;
      RECT 97.13 3.531 97.135 3.745 ;
      RECT 97.125 3.537 97.13 3.745 ;
      RECT 97.12 3.541 97.125 3.748 ;
      RECT 97.115 3.543 97.12 3.751 ;
      RECT 97.11 3.546 97.115 3.754 ;
      RECT 97.1 3.551 97.11 3.758 ;
      RECT 97.095 3.557 97.1 3.763 ;
      RECT 97.085 3.563 97.095 3.767 ;
      RECT 97.07 3.57 97.085 3.773 ;
      RECT 97.041 3.584 97.07 3.783 ;
      RECT 96.955 3.619 97.041 3.815 ;
      RECT 96.935 3.652 96.955 3.844 ;
      RECT 96.915 3.665 96.935 3.855 ;
      RECT 96.895 3.677 96.915 3.866 ;
      RECT 96.845 3.699 96.895 3.886 ;
      RECT 96.83 3.717 96.845 3.903 ;
      RECT 96.825 3.723 96.83 3.906 ;
      RECT 96.82 3.727 96.825 3.909 ;
      RECT 96.815 3.731 96.82 3.913 ;
      RECT 96.81 3.733 96.815 3.916 ;
      RECT 96.8 3.74 96.81 3.919 ;
      RECT 96.795 3.745 96.8 3.923 ;
      RECT 96.79 3.747 96.795 3.926 ;
      RECT 96.785 3.751 96.79 3.929 ;
      RECT 96.78 3.753 96.785 3.933 ;
      RECT 96.765 3.758 96.78 3.938 ;
      RECT 96.76 3.763 96.765 3.941 ;
      RECT 96.755 3.771 96.76 3.944 ;
      RECT 96.75 3.773 96.755 3.947 ;
      RECT 96.745 3.775 96.75 3.95 ;
      RECT 96.735 3.777 96.745 3.956 ;
      RECT 96.7 3.791 96.735 3.968 ;
      RECT 96.69 3.806 96.7 3.978 ;
      RECT 96.615 3.835 96.69 4.002 ;
      RECT 96.61 3.86 96.615 4.025 ;
      RECT 96.595 3.864 96.61 4.031 ;
      RECT 96.585 3.872 96.595 4.036 ;
      RECT 96.555 3.885 96.585 4.04 ;
      RECT 96.545 3.9 96.555 4.045 ;
      RECT 96.535 3.905 96.545 4.048 ;
      RECT 96.53 3.907 96.535 4.05 ;
      RECT 96.515 3.91 96.53 4.053 ;
      RECT 96.51 3.912 96.515 4.056 ;
      RECT 96.49 3.917 96.51 4.06 ;
      RECT 96.46 3.922 96.49 4.068 ;
      RECT 96.435 3.929 96.46 4.076 ;
      RECT 96.43 3.934 96.435 4.081 ;
      RECT 96.4 3.937 96.43 4.085 ;
      RECT 96.36 3.94 96.4 4.095 ;
      RECT 96.325 3.937 96.36 4.107 ;
      RECT 96.315 3.933 96.325 4.114 ;
      RECT 96.29 3.929 96.315 4.12 ;
      RECT 96.285 3.925 96.29 4.125 ;
      RECT 96.245 3.922 96.285 4.125 ;
      RECT 96.23 3.907 96.245 4.126 ;
      RECT 96.207 3.895 96.23 4.126 ;
      RECT 96.121 3.895 96.207 4.127 ;
      RECT 96.035 3.895 96.121 4.129 ;
      RECT 96.015 3.895 96.035 4.126 ;
      RECT 96.01 3.9 96.015 4.121 ;
      RECT 96.005 3.905 96.01 4.119 ;
      RECT 95.995 3.915 96.005 4.117 ;
      RECT 95.99 3.921 95.995 4.11 ;
      RECT 95.985 3.923 95.99 4.095 ;
      RECT 95.98 3.927 95.985 4.085 ;
      RECT 97.44 3.395 97.69 3.655 ;
      RECT 95.165 4.93 95.425 5.19 ;
      RECT 97.46 4.42 97.465 4.63 ;
      RECT 97.465 4.425 97.475 4.625 ;
      RECT 97.415 4.42 97.46 4.645 ;
      RECT 97.405 4.42 97.415 4.665 ;
      RECT 97.386 4.42 97.405 4.67 ;
      RECT 97.3 4.42 97.386 4.667 ;
      RECT 97.27 4.422 97.3 4.665 ;
      RECT 97.215 4.432 97.27 4.663 ;
      RECT 97.15 4.446 97.215 4.661 ;
      RECT 97.145 4.454 97.15 4.66 ;
      RECT 97.13 4.457 97.145 4.658 ;
      RECT 97.065 4.467 97.13 4.654 ;
      RECT 97.017 4.481 97.065 4.655 ;
      RECT 96.931 4.498 97.017 4.669 ;
      RECT 96.845 4.519 96.931 4.686 ;
      RECT 96.825 4.532 96.845 4.696 ;
      RECT 96.78 4.54 96.825 4.703 ;
      RECT 96.745 4.548 96.78 4.711 ;
      RECT 96.711 4.556 96.745 4.719 ;
      RECT 96.625 4.57 96.711 4.731 ;
      RECT 96.59 4.587 96.625 4.743 ;
      RECT 96.581 4.596 96.59 4.747 ;
      RECT 96.495 4.614 96.581 4.764 ;
      RECT 96.436 4.641 96.495 4.791 ;
      RECT 96.35 4.668 96.436 4.819 ;
      RECT 96.33 4.69 96.35 4.839 ;
      RECT 96.27 4.705 96.33 4.855 ;
      RECT 96.26 4.717 96.27 4.868 ;
      RECT 96.255 4.722 96.26 4.871 ;
      RECT 96.245 4.725 96.255 4.874 ;
      RECT 96.24 4.727 96.245 4.877 ;
      RECT 96.21 4.735 96.24 4.884 ;
      RECT 96.195 4.742 96.21 4.892 ;
      RECT 96.185 4.747 96.195 4.896 ;
      RECT 96.18 4.75 96.185 4.899 ;
      RECT 96.17 4.752 96.18 4.902 ;
      RECT 96.135 4.762 96.17 4.911 ;
      RECT 96.06 4.785 96.135 4.933 ;
      RECT 96.04 4.803 96.06 4.951 ;
      RECT 96.01 4.81 96.04 4.961 ;
      RECT 95.99 4.818 96.01 4.971 ;
      RECT 95.98 4.824 95.99 4.978 ;
      RECT 95.961 4.829 95.98 4.984 ;
      RECT 95.875 4.849 95.961 5.004 ;
      RECT 95.86 4.869 95.875 5.023 ;
      RECT 95.815 4.881 95.86 5.034 ;
      RECT 95.75 4.902 95.815 5.057 ;
      RECT 95.71 4.922 95.75 5.078 ;
      RECT 95.7 4.932 95.71 5.088 ;
      RECT 95.65 4.944 95.7 5.099 ;
      RECT 95.63 4.96 95.65 5.111 ;
      RECT 95.6 4.97 95.63 5.117 ;
      RECT 95.59 4.975 95.6 5.119 ;
      RECT 95.521 4.976 95.59 5.125 ;
      RECT 95.435 4.978 95.521 5.135 ;
      RECT 95.425 4.979 95.435 5.14 ;
      RECT 96.695 5.005 96.885 5.215 ;
      RECT 96.685 5.01 96.895 5.208 ;
      RECT 96.67 5.01 96.895 5.173 ;
      RECT 96.59 4.895 96.85 5.155 ;
      RECT 95.505 4.425 95.69 4.72 ;
      RECT 95.495 4.425 95.69 4.718 ;
      RECT 95.48 4.425 95.695 4.713 ;
      RECT 95.48 4.425 95.7 4.71 ;
      RECT 95.475 4.425 95.7 4.708 ;
      RECT 95.47 4.68 95.7 4.698 ;
      RECT 95.475 4.425 95.735 4.685 ;
      RECT 95.435 3.46 95.695 3.72 ;
      RECT 95.245 3.385 95.331 3.718 ;
      RECT 95.22 3.389 95.375 3.714 ;
      RECT 95.331 3.381 95.375 3.714 ;
      RECT 95.331 3.382 95.38 3.713 ;
      RECT 95.245 3.387 95.395 3.712 ;
      RECT 95.22 3.395 95.435 3.711 ;
      RECT 95.215 3.39 95.395 3.706 ;
      RECT 95.205 3.405 95.435 3.613 ;
      RECT 95.205 3.457 95.635 3.613 ;
      RECT 95.205 3.45 95.615 3.613 ;
      RECT 95.205 3.437 95.585 3.613 ;
      RECT 95.205 3.425 95.525 3.613 ;
      RECT 95.205 3.41 95.5 3.613 ;
      RECT 94.405 4.04 94.54 4.335 ;
      RECT 94.665 4.063 94.67 4.25 ;
      RECT 95.385 3.96 95.53 4.195 ;
      RECT 95.545 3.96 95.55 4.185 ;
      RECT 95.58 3.971 95.585 4.165 ;
      RECT 95.575 3.963 95.58 4.17 ;
      RECT 95.555 3.96 95.575 4.175 ;
      RECT 95.55 3.96 95.555 4.183 ;
      RECT 95.54 3.96 95.545 4.188 ;
      RECT 95.53 3.96 95.54 4.193 ;
      RECT 95.36 3.962 95.385 4.195 ;
      RECT 95.31 3.969 95.36 4.195 ;
      RECT 95.305 3.974 95.31 4.195 ;
      RECT 95.266 3.979 95.305 4.196 ;
      RECT 95.18 3.991 95.266 4.197 ;
      RECT 95.171 4.001 95.18 4.197 ;
      RECT 95.085 4.01 95.171 4.199 ;
      RECT 95.061 4.02 95.085 4.201 ;
      RECT 94.975 4.031 95.061 4.202 ;
      RECT 94.945 4.042 94.975 4.204 ;
      RECT 94.915 4.047 94.945 4.206 ;
      RECT 94.89 4.053 94.915 4.209 ;
      RECT 94.875 4.058 94.89 4.21 ;
      RECT 94.83 4.064 94.875 4.21 ;
      RECT 94.825 4.069 94.83 4.211 ;
      RECT 94.805 4.069 94.825 4.213 ;
      RECT 94.785 4.067 94.805 4.218 ;
      RECT 94.75 4.066 94.785 4.225 ;
      RECT 94.72 4.065 94.75 4.235 ;
      RECT 94.67 4.064 94.72 4.245 ;
      RECT 94.58 4.061 94.665 4.335 ;
      RECT 94.555 4.055 94.58 4.335 ;
      RECT 94.54 4.045 94.555 4.335 ;
      RECT 94.355 4.04 94.405 4.255 ;
      RECT 94.345 4.045 94.355 4.245 ;
      RECT 94.585 4.52 94.845 4.78 ;
      RECT 94.585 4.52 94.875 4.673 ;
      RECT 94.585 4.52 94.91 4.658 ;
      RECT 94.84 4.44 95.03 4.65 ;
      RECT 94.83 4.445 95.04 4.643 ;
      RECT 94.795 4.515 95.04 4.643 ;
      RECT 94.825 4.457 94.845 4.78 ;
      RECT 94.81 4.505 95.04 4.643 ;
      RECT 94.815 4.477 94.845 4.78 ;
      RECT 93.895 3.545 93.965 4.65 ;
      RECT 94.63 3.65 94.89 3.91 ;
      RECT 94.21 3.696 94.225 3.905 ;
      RECT 94.546 3.709 94.63 3.86 ;
      RECT 94.46 3.706 94.546 3.86 ;
      RECT 94.421 3.704 94.46 3.86 ;
      RECT 94.335 3.702 94.421 3.86 ;
      RECT 94.275 3.7 94.335 3.871 ;
      RECT 94.24 3.698 94.275 3.889 ;
      RECT 94.225 3.696 94.24 3.9 ;
      RECT 94.195 3.696 94.21 3.913 ;
      RECT 94.185 3.696 94.195 3.918 ;
      RECT 94.16 3.695 94.185 3.923 ;
      RECT 94.145 3.69 94.16 3.929 ;
      RECT 94.14 3.683 94.145 3.934 ;
      RECT 94.115 3.674 94.14 3.94 ;
      RECT 94.07 3.653 94.115 3.953 ;
      RECT 94.06 3.637 94.07 3.963 ;
      RECT 94.045 3.63 94.06 3.973 ;
      RECT 94.035 3.623 94.045 3.99 ;
      RECT 94.03 3.62 94.035 4.02 ;
      RECT 94.025 3.618 94.03 4.05 ;
      RECT 94.02 3.616 94.025 4.087 ;
      RECT 94.005 3.612 94.02 4.154 ;
      RECT 94.005 4.445 94.015 4.645 ;
      RECT 94 3.608 94.005 4.28 ;
      RECT 94 4.432 94.005 4.65 ;
      RECT 93.995 3.606 94 4.365 ;
      RECT 93.995 4.422 94 4.65 ;
      RECT 93.98 3.577 93.995 4.65 ;
      RECT 93.965 3.55 93.98 4.65 ;
      RECT 93.89 3.545 93.895 3.9 ;
      RECT 93.89 3.955 93.895 4.65 ;
      RECT 93.875 3.545 93.89 3.878 ;
      RECT 93.885 3.977 93.89 4.65 ;
      RECT 93.875 4.017 93.885 4.65 ;
      RECT 93.84 3.545 93.875 3.82 ;
      RECT 93.87 4.052 93.875 4.65 ;
      RECT 93.855 4.107 93.87 4.65 ;
      RECT 93.85 4.172 93.855 4.65 ;
      RECT 93.835 4.22 93.85 4.65 ;
      RECT 93.81 3.545 93.84 3.775 ;
      RECT 93.83 4.275 93.835 4.65 ;
      RECT 93.815 4.335 93.83 4.65 ;
      RECT 93.81 4.383 93.815 4.648 ;
      RECT 93.805 3.545 93.81 3.768 ;
      RECT 93.805 4.415 93.81 4.643 ;
      RECT 93.78 3.545 93.805 3.76 ;
      RECT 93.77 3.55 93.78 3.75 ;
      RECT 93.985 4.825 94.005 5.065 ;
      RECT 93.215 4.755 93.22 4.965 ;
      RECT 94.495 4.828 94.505 5.023 ;
      RECT 94.49 4.818 94.495 5.026 ;
      RECT 94.41 4.815 94.49 5.049 ;
      RECT 94.406 4.815 94.41 5.071 ;
      RECT 94.32 4.815 94.406 5.081 ;
      RECT 94.305 4.815 94.32 5.089 ;
      RECT 94.276 4.816 94.305 5.087 ;
      RECT 94.19 4.821 94.276 5.083 ;
      RECT 94.177 4.825 94.19 5.079 ;
      RECT 94.091 4.825 94.177 5.075 ;
      RECT 94.005 4.825 94.091 5.069 ;
      RECT 93.921 4.825 93.985 5.063 ;
      RECT 93.835 4.825 93.921 5.058 ;
      RECT 93.815 4.825 93.835 5.054 ;
      RECT 93.755 4.82 93.815 5.051 ;
      RECT 93.727 4.814 93.755 5.048 ;
      RECT 93.641 4.809 93.727 5.044 ;
      RECT 93.555 4.803 93.641 5.038 ;
      RECT 93.48 4.785 93.555 5.033 ;
      RECT 93.445 4.762 93.48 5.029 ;
      RECT 93.435 4.752 93.445 5.028 ;
      RECT 93.38 4.75 93.435 5.027 ;
      RECT 93.305 4.75 93.38 5.023 ;
      RECT 93.295 4.75 93.305 5.018 ;
      RECT 93.28 4.75 93.295 5.01 ;
      RECT 93.23 4.752 93.28 4.988 ;
      RECT 93.22 4.755 93.23 4.968 ;
      RECT 93.21 4.76 93.215 4.963 ;
      RECT 93.205 4.765 93.21 4.958 ;
      RECT 91.315 3.41 91.575 3.67 ;
      RECT 91.305 3.44 91.575 3.65 ;
      RECT 93.225 3.355 93.485 3.615 ;
      RECT 93.22 3.43 93.225 3.616 ;
      RECT 93.195 3.435 93.22 3.618 ;
      RECT 93.18 3.442 93.195 3.621 ;
      RECT 93.12 3.46 93.18 3.626 ;
      RECT 93.09 3.48 93.12 3.633 ;
      RECT 93.065 3.488 93.09 3.638 ;
      RECT 93.04 3.496 93.065 3.64 ;
      RECT 93.022 3.5 93.04 3.639 ;
      RECT 92.936 3.498 93.022 3.639 ;
      RECT 92.85 3.496 92.936 3.639 ;
      RECT 92.764 3.494 92.85 3.638 ;
      RECT 92.678 3.492 92.764 3.638 ;
      RECT 92.592 3.49 92.678 3.638 ;
      RECT 92.506 3.488 92.592 3.638 ;
      RECT 92.42 3.486 92.506 3.637 ;
      RECT 92.402 3.485 92.42 3.637 ;
      RECT 92.316 3.484 92.402 3.637 ;
      RECT 92.23 3.482 92.316 3.637 ;
      RECT 92.144 3.481 92.23 3.636 ;
      RECT 92.058 3.48 92.144 3.636 ;
      RECT 91.972 3.478 92.058 3.636 ;
      RECT 91.886 3.477 91.972 3.636 ;
      RECT 91.8 3.475 91.886 3.635 ;
      RECT 91.776 3.473 91.8 3.635 ;
      RECT 91.69 3.466 91.776 3.635 ;
      RECT 91.661 3.458 91.69 3.635 ;
      RECT 91.575 3.45 91.661 3.635 ;
      RECT 91.295 3.447 91.305 3.645 ;
      RECT 92.8 4.41 92.805 4.76 ;
      RECT 92.57 4.5 92.71 4.76 ;
      RECT 93.045 4.185 93.09 4.395 ;
      RECT 93.1 4.196 93.11 4.39 ;
      RECT 93.09 4.188 93.1 4.395 ;
      RECT 93.025 4.185 93.045 4.4 ;
      RECT 92.995 4.185 93.025 4.423 ;
      RECT 92.985 4.185 92.995 4.448 ;
      RECT 92.98 4.185 92.985 4.458 ;
      RECT 92.925 4.185 92.98 4.498 ;
      RECT 92.92 4.185 92.925 4.538 ;
      RECT 92.915 4.187 92.92 4.543 ;
      RECT 92.9 4.197 92.915 4.554 ;
      RECT 92.855 4.255 92.9 4.59 ;
      RECT 92.845 4.31 92.855 4.624 ;
      RECT 92.83 4.337 92.845 4.64 ;
      RECT 92.82 4.364 92.83 4.76 ;
      RECT 92.805 4.387 92.82 4.76 ;
      RECT 92.795 4.427 92.8 4.76 ;
      RECT 92.79 4.437 92.795 4.76 ;
      RECT 92.785 4.452 92.79 4.76 ;
      RECT 92.775 4.457 92.785 4.76 ;
      RECT 92.71 4.48 92.775 4.76 ;
      RECT 92.18 3.875 92.41 4.185 ;
      RECT 92.08 3.875 92.41 4.165 ;
      RECT 90.785 3.9 91.045 4.16 ;
      RECT 91.91 3.875 92.41 4.155 ;
      RECT 91.725 3.875 92.41 4.145 ;
      RECT 91.54 3.925 92.41 4.135 ;
      RECT 91.42 3.925 92.41 4.125 ;
      RECT 91.09 3.925 92.41 4.115 ;
      RECT 91.085 3.925 92.41 4.101 ;
      RECT 90.785 3.915 91.37 4.098 ;
      RECT 91.655 3.875 92.47 4.015 ;
      RECT 91.09 3.91 91.36 4.115 ;
      RECT 91.09 3.895 91.35 4.115 ;
      RECT 91.3 4.415 91.56 4.675 ;
      RECT 91.3 4.455 91.665 4.665 ;
      RECT 91.3 4.457 91.67 4.664 ;
      RECT 91.3 4.465 91.675 4.661 ;
      RECT 90.225 3.54 90.325 5.065 ;
      RECT 90.415 4.68 90.465 4.94 ;
      RECT 90.41 3.553 90.415 3.74 ;
      RECT 90.405 4.661 90.415 4.94 ;
      RECT 90.405 3.55 90.41 3.748 ;
      RECT 90.39 3.544 90.405 3.755 ;
      RECT 90.4 4.649 90.405 5.023 ;
      RECT 90.39 4.637 90.4 5.06 ;
      RECT 90.38 3.54 90.39 3.762 ;
      RECT 90.38 4.622 90.39 5.065 ;
      RECT 90.375 3.54 90.38 3.77 ;
      RECT 90.355 4.592 90.38 5.065 ;
      RECT 90.335 3.54 90.375 3.818 ;
      RECT 90.345 4.552 90.355 5.065 ;
      RECT 90.335 4.507 90.345 5.065 ;
      RECT 90.33 3.54 90.335 3.888 ;
      RECT 90.33 4.465 90.335 5.065 ;
      RECT 90.325 3.54 90.33 4.365 ;
      RECT 90.325 4.447 90.33 5.065 ;
      RECT 90.215 3.543 90.225 5.065 ;
      RECT 90.2 3.55 90.215 5.061 ;
      RECT 90.195 3.56 90.2 5.056 ;
      RECT 90.19 3.76 90.195 4.948 ;
      RECT 90.185 3.845 90.19 4.5 ;
      RECT 89.05 10.205 89.345 10.435 ;
      RECT 89.11 8.725 89.28 10.435 ;
      RECT 89.06 9.095 89.41 9.445 ;
      RECT 89.05 8.725 89.34 8.955 ;
      RECT 88.06 10.205 88.355 10.435 ;
      RECT 88.12 8.725 88.29 10.435 ;
      RECT 88.06 8.725 88.35 8.955 ;
      RECT 88.06 8.76 88.91 8.92 ;
      RECT 88.745 8.355 88.91 8.92 ;
      RECT 88.06 8.755 88.455 8.92 ;
      RECT 88.68 8.355 88.97 8.585 ;
      RECT 88.68 8.385 89.14 8.555 ;
      RECT 88.645 4.025 88.97 4.26 ;
      RECT 88.645 4.055 89.135 4.225 ;
      RECT 88.645 3.69 88.835 4.26 ;
      RECT 88.06 3.655 88.35 3.885 ;
      RECT 88.06 3.69 88.835 3.86 ;
      RECT 88.12 2.175 88.29 3.885 ;
      RECT 88.06 2.175 88.355 2.405 ;
      RECT 87.69 4.025 87.98 4.255 ;
      RECT 87.69 4.055 88.15 4.225 ;
      RECT 87.755 2.95 87.92 4.255 ;
      RECT 86.27 2.915 86.56 3.145 ;
      RECT 86.27 2.95 87.92 3.12 ;
      RECT 86.33 2.175 86.5 3.145 ;
      RECT 86.27 2.175 86.56 2.405 ;
      RECT 86.27 10.205 86.56 10.435 ;
      RECT 86.33 9.465 86.5 10.435 ;
      RECT 86.33 9.555 87.92 9.725 ;
      RECT 87.75 8.355 87.92 9.725 ;
      RECT 86.27 9.465 86.56 9.695 ;
      RECT 87.69 8.355 87.98 8.585 ;
      RECT 87.69 8.385 88.15 8.555 ;
      RECT 84.305 4.725 84.655 5.075 ;
      RECT 84.395 3.32 84.565 5.075 ;
      RECT 86.7 3.26 87.05 3.61 ;
      RECT 84.395 3.32 86.015 3.495 ;
      RECT 84.395 3.32 86.67 3.49 ;
      RECT 86.53 3.315 87.05 3.485 ;
      RECT 86.725 9.09 87.05 9.415 ;
      RECT 82.1 9.05 82.45 9.4 ;
      RECT 86.7 9.095 87.05 9.325 ;
      RECT 81.94 9.095 82.45 9.325 ;
      RECT 86.53 9.12 87.05 9.295 ;
      RECT 81.77 9.125 82.45 9.295 ;
      RECT 81.94 9.12 87.05 9.29 ;
      RECT 85.925 3.66 86.245 3.98 ;
      RECT 85.9 3.655 86.19 3.885 ;
      RECT 85.855 3.685 86.245 3.86 ;
      RECT 85.725 3.685 86.245 3.855 ;
      RECT 85.925 8.66 86.245 8.98 ;
      RECT 85.9 8.725 86.245 8.955 ;
      RECT 85.725 8.755 86.245 8.925 ;
      RECT 81.715 4.96 81.755 5.22 ;
      RECT 81.755 4.94 81.76 4.95 ;
      RECT 83.085 4.185 83.095 4.406 ;
      RECT 83.015 4.18 83.085 4.531 ;
      RECT 83.005 4.18 83.015 4.658 ;
      RECT 82.98 4.18 83.005 4.705 ;
      RECT 82.955 4.18 82.98 4.783 ;
      RECT 82.935 4.18 82.955 4.853 ;
      RECT 82.91 4.18 82.935 4.893 ;
      RECT 82.9 4.18 82.91 4.913 ;
      RECT 82.89 4.182 82.9 4.921 ;
      RECT 82.885 4.187 82.89 4.378 ;
      RECT 82.885 4.387 82.89 4.922 ;
      RECT 82.88 4.432 82.885 4.923 ;
      RECT 82.87 4.497 82.88 4.924 ;
      RECT 82.86 4.592 82.87 4.926 ;
      RECT 82.855 4.645 82.86 4.928 ;
      RECT 82.85 4.665 82.855 4.929 ;
      RECT 82.795 4.69 82.85 4.935 ;
      RECT 82.755 4.725 82.795 4.944 ;
      RECT 82.745 4.742 82.755 4.949 ;
      RECT 82.736 4.748 82.745 4.951 ;
      RECT 82.65 4.786 82.736 4.962 ;
      RECT 82.645 4.825 82.65 4.972 ;
      RECT 82.57 4.832 82.645 4.982 ;
      RECT 82.55 4.842 82.57 4.993 ;
      RECT 82.52 4.849 82.55 5.001 ;
      RECT 82.495 4.856 82.52 5.008 ;
      RECT 82.471 4.862 82.495 5.013 ;
      RECT 82.385 4.875 82.471 5.025 ;
      RECT 82.307 4.882 82.385 5.043 ;
      RECT 82.221 4.877 82.307 5.061 ;
      RECT 82.135 4.872 82.221 5.081 ;
      RECT 82.055 4.866 82.135 5.098 ;
      RECT 81.99 4.862 82.055 5.127 ;
      RECT 81.985 4.576 81.99 4.6 ;
      RECT 81.975 4.852 81.99 5.155 ;
      RECT 81.98 4.57 81.985 4.64 ;
      RECT 81.975 4.564 81.98 4.71 ;
      RECT 81.97 4.558 81.975 4.788 ;
      RECT 81.97 4.835 81.975 5.22 ;
      RECT 81.962 4.555 81.97 5.22 ;
      RECT 81.876 4.553 81.962 5.22 ;
      RECT 81.79 4.551 81.876 5.22 ;
      RECT 81.78 4.552 81.79 5.22 ;
      RECT 81.775 4.557 81.78 5.22 ;
      RECT 81.765 4.57 81.775 5.22 ;
      RECT 81.76 4.592 81.765 5.22 ;
      RECT 81.755 4.952 81.76 5.22 ;
      RECT 82.385 4.42 82.39 4.64 ;
      RECT 82.89 3.455 82.925 3.715 ;
      RECT 82.875 3.455 82.89 3.723 ;
      RECT 82.846 3.455 82.875 3.745 ;
      RECT 82.76 3.455 82.846 3.805 ;
      RECT 82.74 3.455 82.76 3.87 ;
      RECT 82.68 3.455 82.74 4.035 ;
      RECT 82.675 3.455 82.68 4.183 ;
      RECT 82.67 3.455 82.675 4.195 ;
      RECT 82.665 3.455 82.67 4.221 ;
      RECT 82.635 3.641 82.665 4.301 ;
      RECT 82.63 3.689 82.635 4.39 ;
      RECT 82.625 3.703 82.63 4.405 ;
      RECT 82.62 3.722 82.625 4.435 ;
      RECT 82.615 3.737 82.62 4.451 ;
      RECT 82.61 3.752 82.615 4.473 ;
      RECT 82.605 3.772 82.61 4.495 ;
      RECT 82.595 3.792 82.605 4.528 ;
      RECT 82.58 3.834 82.595 4.59 ;
      RECT 82.575 3.865 82.58 4.63 ;
      RECT 82.57 3.877 82.575 4.635 ;
      RECT 82.565 3.889 82.57 4.64 ;
      RECT 82.56 3.902 82.565 4.64 ;
      RECT 82.555 3.92 82.56 4.64 ;
      RECT 82.55 3.94 82.555 4.64 ;
      RECT 82.545 3.952 82.55 4.64 ;
      RECT 82.54 3.965 82.545 4.64 ;
      RECT 82.52 4 82.54 4.64 ;
      RECT 82.47 4.102 82.52 4.64 ;
      RECT 82.465 4.187 82.47 4.64 ;
      RECT 82.46 4.195 82.465 4.64 ;
      RECT 82.455 4.212 82.46 4.64 ;
      RECT 82.45 4.227 82.455 4.64 ;
      RECT 82.415 4.292 82.45 4.64 ;
      RECT 82.4 4.357 82.415 4.64 ;
      RECT 82.395 4.387 82.4 4.64 ;
      RECT 82.39 4.412 82.395 4.64 ;
      RECT 82.375 4.422 82.385 4.64 ;
      RECT 82.36 4.435 82.375 4.633 ;
      RECT 82.105 4.025 82.175 4.235 ;
      RECT 81.895 4.002 81.9 4.195 ;
      RECT 79.35 3.93 79.61 4.19 ;
      RECT 82.185 4.212 82.19 4.215 ;
      RECT 82.175 4.03 82.185 4.23 ;
      RECT 82.076 4.023 82.105 4.235 ;
      RECT 81.99 4.015 82.076 4.235 ;
      RECT 81.975 4.009 81.99 4.233 ;
      RECT 81.955 4.008 81.975 4.22 ;
      RECT 81.95 4.007 81.955 4.203 ;
      RECT 81.9 4.004 81.95 4.198 ;
      RECT 81.87 4.001 81.895 4.193 ;
      RECT 81.85 3.999 81.87 4.188 ;
      RECT 81.835 3.997 81.85 4.185 ;
      RECT 81.805 3.995 81.835 4.183 ;
      RECT 81.74 3.991 81.805 4.175 ;
      RECT 81.71 3.986 81.74 4.17 ;
      RECT 81.69 3.984 81.71 4.168 ;
      RECT 81.66 3.981 81.69 4.163 ;
      RECT 81.6 3.977 81.66 4.155 ;
      RECT 81.595 3.974 81.6 4.15 ;
      RECT 81.525 3.972 81.595 4.145 ;
      RECT 81.496 3.968 81.525 4.138 ;
      RECT 81.41 3.963 81.496 4.13 ;
      RECT 81.376 3.958 81.41 4.122 ;
      RECT 81.29 3.95 81.376 4.114 ;
      RECT 81.251 3.943 81.29 4.106 ;
      RECT 81.165 3.938 81.251 4.098 ;
      RECT 81.1 3.932 81.165 4.088 ;
      RECT 81.08 3.927 81.1 4.083 ;
      RECT 81.071 3.924 81.08 4.082 ;
      RECT 80.985 3.92 81.071 4.076 ;
      RECT 80.945 3.916 80.985 4.068 ;
      RECT 80.925 3.912 80.945 4.066 ;
      RECT 80.865 3.912 80.925 4.063 ;
      RECT 80.845 3.915 80.865 4.061 ;
      RECT 80.824 3.915 80.845 4.061 ;
      RECT 80.738 3.917 80.824 4.065 ;
      RECT 80.652 3.919 80.738 4.071 ;
      RECT 80.566 3.921 80.652 4.078 ;
      RECT 80.48 3.924 80.566 4.084 ;
      RECT 80.446 3.925 80.48 4.089 ;
      RECT 80.36 3.928 80.446 4.094 ;
      RECT 80.331 3.935 80.36 4.099 ;
      RECT 80.245 3.935 80.331 4.104 ;
      RECT 80.212 3.935 80.245 4.109 ;
      RECT 80.126 3.937 80.212 4.114 ;
      RECT 80.04 3.939 80.126 4.121 ;
      RECT 79.976 3.941 80.04 4.127 ;
      RECT 79.89 3.943 79.976 4.133 ;
      RECT 79.887 3.945 79.89 4.136 ;
      RECT 79.801 3.946 79.887 4.14 ;
      RECT 79.715 3.949 79.801 4.147 ;
      RECT 79.696 3.951 79.715 4.151 ;
      RECT 79.61 3.953 79.696 4.156 ;
      RECT 79.34 3.965 79.35 4.16 ;
      RECT 81.51 10.205 81.8 10.435 ;
      RECT 81.57 9.465 81.74 10.435 ;
      RECT 81.46 9.49 81.835 9.86 ;
      RECT 81.51 9.465 81.8 9.86 ;
      RECT 81.575 3.545 81.76 3.755 ;
      RECT 81.57 3.546 81.765 3.753 ;
      RECT 81.565 3.551 81.775 3.748 ;
      RECT 81.56 3.527 81.565 3.745 ;
      RECT 81.53 3.524 81.56 3.738 ;
      RECT 81.525 3.52 81.53 3.729 ;
      RECT 81.49 3.551 81.775 3.724 ;
      RECT 81.265 3.46 81.525 3.72 ;
      RECT 81.565 3.529 81.57 3.748 ;
      RECT 81.57 3.53 81.575 3.753 ;
      RECT 81.265 3.542 81.645 3.72 ;
      RECT 81.265 3.54 81.63 3.72 ;
      RECT 81.265 3.535 81.62 3.72 ;
      RECT 81.22 4.45 81.27 4.735 ;
      RECT 81.165 4.42 81.17 4.735 ;
      RECT 81.135 4.4 81.14 4.735 ;
      RECT 81.285 4.45 81.345 4.71 ;
      RECT 81.28 4.45 81.285 4.718 ;
      RECT 81.27 4.45 81.28 4.73 ;
      RECT 81.185 4.44 81.22 4.735 ;
      RECT 81.18 4.427 81.185 4.735 ;
      RECT 81.17 4.422 81.18 4.735 ;
      RECT 81.15 4.412 81.165 4.735 ;
      RECT 81.14 4.405 81.15 4.735 ;
      RECT 81.13 4.397 81.135 4.735 ;
      RECT 81.1 4.387 81.13 4.735 ;
      RECT 81.085 4.375 81.1 4.735 ;
      RECT 81.07 4.365 81.085 4.73 ;
      RECT 81.05 4.355 81.07 4.705 ;
      RECT 81.04 4.347 81.05 4.682 ;
      RECT 81.01 4.33 81.04 4.672 ;
      RECT 81.005 4.307 81.01 4.663 ;
      RECT 81 4.294 81.005 4.661 ;
      RECT 80.985 4.27 81 4.655 ;
      RECT 80.98 4.246 80.985 4.649 ;
      RECT 80.97 4.235 80.98 4.644 ;
      RECT 80.965 4.225 80.97 4.64 ;
      RECT 80.96 4.217 80.965 4.637 ;
      RECT 80.95 4.212 80.96 4.633 ;
      RECT 80.945 4.207 80.95 4.629 ;
      RECT 80.86 4.205 80.945 4.604 ;
      RECT 80.83 4.205 80.86 4.57 ;
      RECT 80.815 4.205 80.83 4.553 ;
      RECT 80.76 4.205 80.815 4.498 ;
      RECT 80.755 4.21 80.76 4.447 ;
      RECT 80.745 4.215 80.755 4.437 ;
      RECT 80.74 4.225 80.745 4.423 ;
      RECT 80.69 4.965 80.95 5.225 ;
      RECT 80.61 4.98 80.95 5.201 ;
      RECT 80.59 4.98 80.95 5.196 ;
      RECT 80.566 4.98 80.95 5.194 ;
      RECT 80.48 4.98 80.95 5.189 ;
      RECT 80.33 4.92 80.59 5.185 ;
      RECT 80.285 4.98 80.95 5.18 ;
      RECT 80.28 4.987 80.95 5.175 ;
      RECT 80.295 4.975 80.61 5.185 ;
      RECT 80.185 3.41 80.445 3.67 ;
      RECT 80.185 3.467 80.45 3.663 ;
      RECT 80.185 3.497 80.455 3.595 ;
      RECT 80.245 3.928 80.36 3.93 ;
      RECT 80.331 3.925 80.36 3.93 ;
      RECT 79.355 4.929 79.38 5.169 ;
      RECT 79.34 4.932 79.43 5.163 ;
      RECT 79.335 4.937 79.516 5.158 ;
      RECT 79.33 4.945 79.58 5.156 ;
      RECT 79.33 4.945 79.59 5.155 ;
      RECT 79.325 4.952 79.6 5.148 ;
      RECT 79.325 4.952 79.686 5.137 ;
      RECT 79.32 4.987 79.686 5.133 ;
      RECT 79.32 4.987 79.695 5.122 ;
      RECT 79.6 4.86 79.86 5.12 ;
      RECT 79.31 5.037 79.86 5.118 ;
      RECT 79.58 4.905 79.6 5.153 ;
      RECT 79.516 4.908 79.58 5.157 ;
      RECT 79.43 4.913 79.516 5.162 ;
      RECT 79.36 4.924 79.86 5.12 ;
      RECT 79.38 4.918 79.43 5.167 ;
      RECT 79.505 3.395 79.515 3.657 ;
      RECT 79.495 3.452 79.505 3.66 ;
      RECT 79.47 3.457 79.495 3.666 ;
      RECT 79.445 3.461 79.47 3.678 ;
      RECT 79.435 3.464 79.445 3.688 ;
      RECT 79.43 3.465 79.435 3.693 ;
      RECT 79.425 3.466 79.43 3.698 ;
      RECT 79.42 3.467 79.425 3.7 ;
      RECT 79.395 3.47 79.42 3.703 ;
      RECT 79.365 3.476 79.395 3.706 ;
      RECT 79.3 3.487 79.365 3.709 ;
      RECT 79.255 3.495 79.3 3.713 ;
      RECT 79.24 3.495 79.255 3.721 ;
      RECT 79.235 3.496 79.24 3.728 ;
      RECT 79.23 3.498 79.235 3.731 ;
      RECT 79.225 3.502 79.23 3.734 ;
      RECT 79.215 3.51 79.225 3.738 ;
      RECT 79.21 3.523 79.215 3.743 ;
      RECT 79.205 3.531 79.21 3.745 ;
      RECT 79.2 3.537 79.205 3.745 ;
      RECT 79.195 3.541 79.2 3.748 ;
      RECT 79.19 3.543 79.195 3.751 ;
      RECT 79.185 3.546 79.19 3.754 ;
      RECT 79.175 3.551 79.185 3.758 ;
      RECT 79.17 3.557 79.175 3.763 ;
      RECT 79.16 3.563 79.17 3.767 ;
      RECT 79.145 3.57 79.16 3.773 ;
      RECT 79.116 3.584 79.145 3.783 ;
      RECT 79.03 3.619 79.116 3.815 ;
      RECT 79.01 3.652 79.03 3.844 ;
      RECT 78.99 3.665 79.01 3.855 ;
      RECT 78.97 3.677 78.99 3.866 ;
      RECT 78.92 3.699 78.97 3.886 ;
      RECT 78.905 3.717 78.92 3.903 ;
      RECT 78.9 3.723 78.905 3.906 ;
      RECT 78.895 3.727 78.9 3.909 ;
      RECT 78.89 3.731 78.895 3.913 ;
      RECT 78.885 3.733 78.89 3.916 ;
      RECT 78.875 3.74 78.885 3.919 ;
      RECT 78.87 3.745 78.875 3.923 ;
      RECT 78.865 3.747 78.87 3.926 ;
      RECT 78.86 3.751 78.865 3.929 ;
      RECT 78.855 3.753 78.86 3.933 ;
      RECT 78.84 3.758 78.855 3.938 ;
      RECT 78.835 3.763 78.84 3.941 ;
      RECT 78.83 3.771 78.835 3.944 ;
      RECT 78.825 3.773 78.83 3.947 ;
      RECT 78.82 3.775 78.825 3.95 ;
      RECT 78.81 3.777 78.82 3.956 ;
      RECT 78.775 3.791 78.81 3.968 ;
      RECT 78.765 3.806 78.775 3.978 ;
      RECT 78.69 3.835 78.765 4.002 ;
      RECT 78.685 3.86 78.69 4.025 ;
      RECT 78.67 3.864 78.685 4.031 ;
      RECT 78.66 3.872 78.67 4.036 ;
      RECT 78.63 3.885 78.66 4.04 ;
      RECT 78.62 3.9 78.63 4.045 ;
      RECT 78.61 3.905 78.62 4.048 ;
      RECT 78.605 3.907 78.61 4.05 ;
      RECT 78.59 3.91 78.605 4.053 ;
      RECT 78.585 3.912 78.59 4.056 ;
      RECT 78.565 3.917 78.585 4.06 ;
      RECT 78.535 3.922 78.565 4.068 ;
      RECT 78.51 3.929 78.535 4.076 ;
      RECT 78.505 3.934 78.51 4.081 ;
      RECT 78.475 3.937 78.505 4.085 ;
      RECT 78.435 3.94 78.475 4.095 ;
      RECT 78.4 3.937 78.435 4.107 ;
      RECT 78.39 3.933 78.4 4.114 ;
      RECT 78.365 3.929 78.39 4.12 ;
      RECT 78.36 3.925 78.365 4.125 ;
      RECT 78.32 3.922 78.36 4.125 ;
      RECT 78.305 3.907 78.32 4.126 ;
      RECT 78.282 3.895 78.305 4.126 ;
      RECT 78.196 3.895 78.282 4.127 ;
      RECT 78.11 3.895 78.196 4.129 ;
      RECT 78.09 3.895 78.11 4.126 ;
      RECT 78.085 3.9 78.09 4.121 ;
      RECT 78.08 3.905 78.085 4.119 ;
      RECT 78.07 3.915 78.08 4.117 ;
      RECT 78.065 3.921 78.07 4.11 ;
      RECT 78.06 3.923 78.065 4.095 ;
      RECT 78.055 3.927 78.06 4.085 ;
      RECT 79.515 3.395 79.765 3.655 ;
      RECT 77.24 4.93 77.5 5.19 ;
      RECT 79.535 4.42 79.54 4.63 ;
      RECT 79.54 4.425 79.55 4.625 ;
      RECT 79.49 4.42 79.535 4.645 ;
      RECT 79.48 4.42 79.49 4.665 ;
      RECT 79.461 4.42 79.48 4.67 ;
      RECT 79.375 4.42 79.461 4.667 ;
      RECT 79.345 4.422 79.375 4.665 ;
      RECT 79.29 4.432 79.345 4.663 ;
      RECT 79.225 4.446 79.29 4.661 ;
      RECT 79.22 4.454 79.225 4.66 ;
      RECT 79.205 4.457 79.22 4.658 ;
      RECT 79.14 4.467 79.205 4.654 ;
      RECT 79.092 4.481 79.14 4.655 ;
      RECT 79.006 4.498 79.092 4.669 ;
      RECT 78.92 4.519 79.006 4.686 ;
      RECT 78.9 4.532 78.92 4.696 ;
      RECT 78.855 4.54 78.9 4.703 ;
      RECT 78.82 4.548 78.855 4.711 ;
      RECT 78.786 4.556 78.82 4.719 ;
      RECT 78.7 4.57 78.786 4.731 ;
      RECT 78.665 4.587 78.7 4.743 ;
      RECT 78.656 4.596 78.665 4.747 ;
      RECT 78.57 4.614 78.656 4.764 ;
      RECT 78.511 4.641 78.57 4.791 ;
      RECT 78.425 4.668 78.511 4.819 ;
      RECT 78.405 4.69 78.425 4.839 ;
      RECT 78.345 4.705 78.405 4.855 ;
      RECT 78.335 4.717 78.345 4.868 ;
      RECT 78.33 4.722 78.335 4.871 ;
      RECT 78.32 4.725 78.33 4.874 ;
      RECT 78.315 4.727 78.32 4.877 ;
      RECT 78.285 4.735 78.315 4.884 ;
      RECT 78.27 4.742 78.285 4.892 ;
      RECT 78.26 4.747 78.27 4.896 ;
      RECT 78.255 4.75 78.26 4.899 ;
      RECT 78.245 4.752 78.255 4.902 ;
      RECT 78.21 4.762 78.245 4.911 ;
      RECT 78.135 4.785 78.21 4.933 ;
      RECT 78.115 4.803 78.135 4.951 ;
      RECT 78.085 4.81 78.115 4.961 ;
      RECT 78.065 4.818 78.085 4.971 ;
      RECT 78.055 4.824 78.065 4.978 ;
      RECT 78.036 4.829 78.055 4.984 ;
      RECT 77.95 4.849 78.036 5.004 ;
      RECT 77.935 4.869 77.95 5.023 ;
      RECT 77.89 4.881 77.935 5.034 ;
      RECT 77.825 4.902 77.89 5.057 ;
      RECT 77.785 4.922 77.825 5.078 ;
      RECT 77.775 4.932 77.785 5.088 ;
      RECT 77.725 4.944 77.775 5.099 ;
      RECT 77.705 4.96 77.725 5.111 ;
      RECT 77.675 4.97 77.705 5.117 ;
      RECT 77.665 4.975 77.675 5.119 ;
      RECT 77.596 4.976 77.665 5.125 ;
      RECT 77.51 4.978 77.596 5.135 ;
      RECT 77.5 4.979 77.51 5.14 ;
      RECT 78.77 5.005 78.96 5.215 ;
      RECT 78.76 5.01 78.97 5.208 ;
      RECT 78.745 5.01 78.97 5.173 ;
      RECT 78.665 4.895 78.925 5.155 ;
      RECT 77.58 4.425 77.765 4.72 ;
      RECT 77.57 4.425 77.765 4.718 ;
      RECT 77.555 4.425 77.77 4.713 ;
      RECT 77.555 4.425 77.775 4.71 ;
      RECT 77.55 4.425 77.775 4.708 ;
      RECT 77.545 4.68 77.775 4.698 ;
      RECT 77.55 4.425 77.81 4.685 ;
      RECT 77.51 3.46 77.77 3.72 ;
      RECT 77.32 3.385 77.406 3.718 ;
      RECT 77.295 3.389 77.45 3.714 ;
      RECT 77.406 3.381 77.45 3.714 ;
      RECT 77.406 3.382 77.455 3.713 ;
      RECT 77.32 3.387 77.47 3.712 ;
      RECT 77.295 3.395 77.51 3.711 ;
      RECT 77.29 3.39 77.47 3.706 ;
      RECT 77.28 3.405 77.51 3.613 ;
      RECT 77.28 3.457 77.71 3.613 ;
      RECT 77.28 3.45 77.69 3.613 ;
      RECT 77.28 3.437 77.66 3.613 ;
      RECT 77.28 3.425 77.6 3.613 ;
      RECT 77.28 3.41 77.575 3.613 ;
      RECT 76.48 4.04 76.615 4.335 ;
      RECT 76.74 4.063 76.745 4.25 ;
      RECT 77.46 3.96 77.605 4.195 ;
      RECT 77.62 3.96 77.625 4.185 ;
      RECT 77.655 3.971 77.66 4.165 ;
      RECT 77.65 3.963 77.655 4.17 ;
      RECT 77.63 3.96 77.65 4.175 ;
      RECT 77.625 3.96 77.63 4.183 ;
      RECT 77.615 3.96 77.62 4.188 ;
      RECT 77.605 3.96 77.615 4.193 ;
      RECT 77.435 3.962 77.46 4.195 ;
      RECT 77.385 3.969 77.435 4.195 ;
      RECT 77.38 3.974 77.385 4.195 ;
      RECT 77.341 3.979 77.38 4.196 ;
      RECT 77.255 3.991 77.341 4.197 ;
      RECT 77.246 4.001 77.255 4.197 ;
      RECT 77.16 4.01 77.246 4.199 ;
      RECT 77.136 4.02 77.16 4.201 ;
      RECT 77.05 4.031 77.136 4.202 ;
      RECT 77.02 4.042 77.05 4.204 ;
      RECT 76.99 4.047 77.02 4.206 ;
      RECT 76.965 4.053 76.99 4.209 ;
      RECT 76.95 4.058 76.965 4.21 ;
      RECT 76.905 4.064 76.95 4.21 ;
      RECT 76.9 4.069 76.905 4.211 ;
      RECT 76.88 4.069 76.9 4.213 ;
      RECT 76.86 4.067 76.88 4.218 ;
      RECT 76.825 4.066 76.86 4.225 ;
      RECT 76.795 4.065 76.825 4.235 ;
      RECT 76.745 4.064 76.795 4.245 ;
      RECT 76.655 4.061 76.74 4.335 ;
      RECT 76.63 4.055 76.655 4.335 ;
      RECT 76.615 4.045 76.63 4.335 ;
      RECT 76.43 4.04 76.48 4.255 ;
      RECT 76.42 4.045 76.43 4.245 ;
      RECT 76.66 4.52 76.92 4.78 ;
      RECT 76.66 4.52 76.95 4.673 ;
      RECT 76.66 4.52 76.985 4.658 ;
      RECT 76.915 4.44 77.105 4.65 ;
      RECT 76.905 4.445 77.115 4.643 ;
      RECT 76.87 4.515 77.115 4.643 ;
      RECT 76.9 4.457 76.92 4.78 ;
      RECT 76.885 4.505 77.115 4.643 ;
      RECT 76.89 4.477 76.92 4.78 ;
      RECT 75.97 3.545 76.04 4.65 ;
      RECT 76.705 3.65 76.965 3.91 ;
      RECT 76.285 3.696 76.3 3.905 ;
      RECT 76.621 3.709 76.705 3.86 ;
      RECT 76.535 3.706 76.621 3.86 ;
      RECT 76.496 3.704 76.535 3.86 ;
      RECT 76.41 3.702 76.496 3.86 ;
      RECT 76.35 3.7 76.41 3.871 ;
      RECT 76.315 3.698 76.35 3.889 ;
      RECT 76.3 3.696 76.315 3.9 ;
      RECT 76.27 3.696 76.285 3.913 ;
      RECT 76.26 3.696 76.27 3.918 ;
      RECT 76.235 3.695 76.26 3.923 ;
      RECT 76.22 3.69 76.235 3.929 ;
      RECT 76.215 3.683 76.22 3.934 ;
      RECT 76.19 3.674 76.215 3.94 ;
      RECT 76.145 3.653 76.19 3.953 ;
      RECT 76.135 3.637 76.145 3.963 ;
      RECT 76.12 3.63 76.135 3.973 ;
      RECT 76.11 3.623 76.12 3.99 ;
      RECT 76.105 3.62 76.11 4.02 ;
      RECT 76.1 3.618 76.105 4.05 ;
      RECT 76.095 3.616 76.1 4.087 ;
      RECT 76.08 3.612 76.095 4.154 ;
      RECT 76.08 4.445 76.09 4.645 ;
      RECT 76.075 3.608 76.08 4.28 ;
      RECT 76.075 4.432 76.08 4.65 ;
      RECT 76.07 3.606 76.075 4.365 ;
      RECT 76.07 4.422 76.075 4.65 ;
      RECT 76.055 3.577 76.07 4.65 ;
      RECT 76.04 3.55 76.055 4.65 ;
      RECT 75.965 3.545 75.97 3.9 ;
      RECT 75.965 3.955 75.97 4.65 ;
      RECT 75.95 3.545 75.965 3.878 ;
      RECT 75.96 3.977 75.965 4.65 ;
      RECT 75.95 4.017 75.96 4.65 ;
      RECT 75.915 3.545 75.95 3.82 ;
      RECT 75.945 4.052 75.95 4.65 ;
      RECT 75.93 4.107 75.945 4.65 ;
      RECT 75.925 4.172 75.93 4.65 ;
      RECT 75.91 4.22 75.925 4.65 ;
      RECT 75.885 3.545 75.915 3.775 ;
      RECT 75.905 4.275 75.91 4.65 ;
      RECT 75.89 4.335 75.905 4.65 ;
      RECT 75.885 4.383 75.89 4.648 ;
      RECT 75.88 3.545 75.885 3.768 ;
      RECT 75.88 4.415 75.885 4.643 ;
      RECT 75.855 3.545 75.88 3.76 ;
      RECT 75.845 3.55 75.855 3.75 ;
      RECT 76.06 4.825 76.08 5.065 ;
      RECT 75.29 4.755 75.295 4.965 ;
      RECT 76.57 4.828 76.58 5.023 ;
      RECT 76.565 4.818 76.57 5.026 ;
      RECT 76.485 4.815 76.565 5.049 ;
      RECT 76.481 4.815 76.485 5.071 ;
      RECT 76.395 4.815 76.481 5.081 ;
      RECT 76.38 4.815 76.395 5.089 ;
      RECT 76.351 4.816 76.38 5.087 ;
      RECT 76.265 4.821 76.351 5.083 ;
      RECT 76.252 4.825 76.265 5.079 ;
      RECT 76.166 4.825 76.252 5.075 ;
      RECT 76.08 4.825 76.166 5.069 ;
      RECT 75.996 4.825 76.06 5.063 ;
      RECT 75.91 4.825 75.996 5.058 ;
      RECT 75.89 4.825 75.91 5.054 ;
      RECT 75.83 4.82 75.89 5.051 ;
      RECT 75.802 4.814 75.83 5.048 ;
      RECT 75.716 4.809 75.802 5.044 ;
      RECT 75.63 4.803 75.716 5.038 ;
      RECT 75.555 4.785 75.63 5.033 ;
      RECT 75.52 4.762 75.555 5.029 ;
      RECT 75.51 4.752 75.52 5.028 ;
      RECT 75.455 4.75 75.51 5.027 ;
      RECT 75.38 4.75 75.455 5.023 ;
      RECT 75.37 4.75 75.38 5.018 ;
      RECT 75.355 4.75 75.37 5.01 ;
      RECT 75.305 4.752 75.355 4.988 ;
      RECT 75.295 4.755 75.305 4.968 ;
      RECT 75.285 4.76 75.29 4.963 ;
      RECT 75.28 4.765 75.285 4.958 ;
      RECT 73.39 3.41 73.65 3.67 ;
      RECT 73.38 3.44 73.65 3.65 ;
      RECT 75.3 3.355 75.56 3.615 ;
      RECT 75.295 3.43 75.3 3.616 ;
      RECT 75.27 3.435 75.295 3.618 ;
      RECT 75.255 3.442 75.27 3.621 ;
      RECT 75.195 3.46 75.255 3.626 ;
      RECT 75.165 3.48 75.195 3.633 ;
      RECT 75.14 3.488 75.165 3.638 ;
      RECT 75.115 3.496 75.14 3.64 ;
      RECT 75.097 3.5 75.115 3.639 ;
      RECT 75.011 3.498 75.097 3.639 ;
      RECT 74.925 3.496 75.011 3.639 ;
      RECT 74.839 3.494 74.925 3.638 ;
      RECT 74.753 3.492 74.839 3.638 ;
      RECT 74.667 3.49 74.753 3.638 ;
      RECT 74.581 3.488 74.667 3.638 ;
      RECT 74.495 3.486 74.581 3.637 ;
      RECT 74.477 3.485 74.495 3.637 ;
      RECT 74.391 3.484 74.477 3.637 ;
      RECT 74.305 3.482 74.391 3.637 ;
      RECT 74.219 3.481 74.305 3.636 ;
      RECT 74.133 3.48 74.219 3.636 ;
      RECT 74.047 3.478 74.133 3.636 ;
      RECT 73.961 3.477 74.047 3.636 ;
      RECT 73.875 3.475 73.961 3.635 ;
      RECT 73.851 3.473 73.875 3.635 ;
      RECT 73.765 3.466 73.851 3.635 ;
      RECT 73.736 3.458 73.765 3.635 ;
      RECT 73.65 3.45 73.736 3.635 ;
      RECT 73.37 3.447 73.38 3.645 ;
      RECT 74.875 4.41 74.88 4.76 ;
      RECT 74.645 4.5 74.785 4.76 ;
      RECT 75.12 4.185 75.165 4.395 ;
      RECT 75.175 4.196 75.185 4.39 ;
      RECT 75.165 4.188 75.175 4.395 ;
      RECT 75.1 4.185 75.12 4.4 ;
      RECT 75.07 4.185 75.1 4.423 ;
      RECT 75.06 4.185 75.07 4.448 ;
      RECT 75.055 4.185 75.06 4.458 ;
      RECT 75 4.185 75.055 4.498 ;
      RECT 74.995 4.185 75 4.538 ;
      RECT 74.99 4.187 74.995 4.543 ;
      RECT 74.975 4.197 74.99 4.554 ;
      RECT 74.93 4.255 74.975 4.59 ;
      RECT 74.92 4.31 74.93 4.624 ;
      RECT 74.905 4.337 74.92 4.64 ;
      RECT 74.895 4.364 74.905 4.76 ;
      RECT 74.88 4.387 74.895 4.76 ;
      RECT 74.87 4.427 74.875 4.76 ;
      RECT 74.865 4.437 74.87 4.76 ;
      RECT 74.86 4.452 74.865 4.76 ;
      RECT 74.85 4.457 74.86 4.76 ;
      RECT 74.785 4.48 74.85 4.76 ;
      RECT 74.255 3.875 74.485 4.185 ;
      RECT 74.155 3.875 74.485 4.165 ;
      RECT 72.86 3.9 73.12 4.16 ;
      RECT 73.985 3.875 74.485 4.155 ;
      RECT 73.8 3.875 74.485 4.145 ;
      RECT 73.615 3.925 74.485 4.135 ;
      RECT 73.495 3.925 74.485 4.125 ;
      RECT 73.165 3.925 74.485 4.115 ;
      RECT 73.16 3.925 74.485 4.101 ;
      RECT 72.86 3.915 73.445 4.098 ;
      RECT 73.73 3.875 74.545 4.015 ;
      RECT 73.165 3.91 73.435 4.115 ;
      RECT 73.165 3.895 73.425 4.115 ;
      RECT 73.375 4.415 73.635 4.675 ;
      RECT 73.375 4.455 73.74 4.665 ;
      RECT 73.375 4.457 73.745 4.664 ;
      RECT 73.375 4.465 73.75 4.661 ;
      RECT 72.3 3.54 72.4 5.065 ;
      RECT 72.49 4.68 72.54 4.94 ;
      RECT 72.485 3.553 72.49 3.74 ;
      RECT 72.48 4.661 72.49 4.94 ;
      RECT 72.48 3.55 72.485 3.748 ;
      RECT 72.465 3.544 72.48 3.755 ;
      RECT 72.475 4.649 72.48 5.023 ;
      RECT 72.465 4.637 72.475 5.06 ;
      RECT 72.455 3.54 72.465 3.762 ;
      RECT 72.455 4.622 72.465 5.065 ;
      RECT 72.45 3.54 72.455 3.77 ;
      RECT 72.43 4.592 72.455 5.065 ;
      RECT 72.41 3.54 72.45 3.818 ;
      RECT 72.42 4.552 72.43 5.065 ;
      RECT 72.41 4.507 72.42 5.065 ;
      RECT 72.405 3.54 72.41 3.888 ;
      RECT 72.405 4.465 72.41 5.065 ;
      RECT 72.4 3.54 72.405 4.365 ;
      RECT 72.4 4.447 72.405 5.065 ;
      RECT 72.29 3.543 72.3 5.065 ;
      RECT 72.275 3.55 72.29 5.061 ;
      RECT 72.27 3.56 72.275 5.056 ;
      RECT 72.265 3.76 72.27 4.948 ;
      RECT 72.26 3.845 72.265 4.5 ;
      RECT 71.125 10.205 71.42 10.435 ;
      RECT 71.185 8.725 71.355 10.435 ;
      RECT 71.135 9.095 71.485 9.445 ;
      RECT 71.125 8.725 71.415 8.955 ;
      RECT 70.135 10.205 70.43 10.435 ;
      RECT 70.195 8.725 70.365 10.435 ;
      RECT 70.135 8.725 70.425 8.955 ;
      RECT 70.135 8.76 70.985 8.92 ;
      RECT 70.82 8.355 70.985 8.92 ;
      RECT 70.135 8.755 70.53 8.92 ;
      RECT 70.755 8.355 71.045 8.585 ;
      RECT 70.755 8.385 71.215 8.555 ;
      RECT 70.72 4.025 71.045 4.26 ;
      RECT 70.72 4.055 71.21 4.225 ;
      RECT 70.72 3.69 70.91 4.26 ;
      RECT 70.135 3.655 70.425 3.885 ;
      RECT 70.135 3.69 70.91 3.86 ;
      RECT 70.195 2.175 70.365 3.885 ;
      RECT 70.135 2.175 70.43 2.405 ;
      RECT 69.765 4.025 70.055 4.255 ;
      RECT 69.765 4.055 70.225 4.225 ;
      RECT 69.83 2.95 69.995 4.255 ;
      RECT 68.345 2.915 68.635 3.145 ;
      RECT 68.345 2.95 69.995 3.12 ;
      RECT 68.405 2.175 68.575 3.145 ;
      RECT 68.345 2.175 68.635 2.405 ;
      RECT 68.345 10.205 68.635 10.435 ;
      RECT 68.405 9.465 68.575 10.435 ;
      RECT 68.405 9.555 69.995 9.725 ;
      RECT 69.825 8.355 69.995 9.725 ;
      RECT 68.345 9.465 68.635 9.695 ;
      RECT 69.765 8.355 70.055 8.585 ;
      RECT 69.765 8.385 70.225 8.555 ;
      RECT 66.38 4.725 66.73 5.075 ;
      RECT 66.47 3.32 66.64 5.075 ;
      RECT 68.775 3.26 69.125 3.61 ;
      RECT 66.47 3.32 68.09 3.495 ;
      RECT 66.47 3.32 68.745 3.49 ;
      RECT 68.605 3.315 69.125 3.485 ;
      RECT 68.8 9.09 69.125 9.415 ;
      RECT 64.23 9.05 64.58 9.4 ;
      RECT 68.775 9.095 69.125 9.325 ;
      RECT 64.015 9.095 64.58 9.325 ;
      RECT 68.605 9.12 69.125 9.295 ;
      RECT 63.845 9.125 64.58 9.295 ;
      RECT 64.015 9.12 69.125 9.29 ;
      RECT 68 3.66 68.32 3.98 ;
      RECT 67.975 3.655 68.265 3.885 ;
      RECT 67.93 3.685 68.32 3.86 ;
      RECT 67.8 3.685 68.32 3.855 ;
      RECT 68 8.66 68.32 8.98 ;
      RECT 67.975 8.725 68.32 8.955 ;
      RECT 67.8 8.755 68.32 8.925 ;
      RECT 63.79 4.96 63.83 5.22 ;
      RECT 63.83 4.94 63.835 4.95 ;
      RECT 65.16 4.185 65.17 4.406 ;
      RECT 65.09 4.18 65.16 4.531 ;
      RECT 65.08 4.18 65.09 4.658 ;
      RECT 65.055 4.18 65.08 4.705 ;
      RECT 65.03 4.18 65.055 4.783 ;
      RECT 65.01 4.18 65.03 4.853 ;
      RECT 64.985 4.18 65.01 4.893 ;
      RECT 64.975 4.18 64.985 4.913 ;
      RECT 64.965 4.182 64.975 4.921 ;
      RECT 64.96 4.187 64.965 4.378 ;
      RECT 64.96 4.387 64.965 4.922 ;
      RECT 64.955 4.432 64.96 4.923 ;
      RECT 64.945 4.497 64.955 4.924 ;
      RECT 64.935 4.592 64.945 4.926 ;
      RECT 64.93 4.645 64.935 4.928 ;
      RECT 64.925 4.665 64.93 4.929 ;
      RECT 64.87 4.69 64.925 4.935 ;
      RECT 64.83 4.725 64.87 4.944 ;
      RECT 64.82 4.742 64.83 4.949 ;
      RECT 64.811 4.748 64.82 4.951 ;
      RECT 64.725 4.786 64.811 4.962 ;
      RECT 64.72 4.825 64.725 4.972 ;
      RECT 64.645 4.832 64.72 4.982 ;
      RECT 64.625 4.842 64.645 4.993 ;
      RECT 64.595 4.849 64.625 5.001 ;
      RECT 64.57 4.856 64.595 5.008 ;
      RECT 64.546 4.862 64.57 5.013 ;
      RECT 64.46 4.875 64.546 5.025 ;
      RECT 64.382 4.882 64.46 5.043 ;
      RECT 64.296 4.877 64.382 5.061 ;
      RECT 64.21 4.872 64.296 5.081 ;
      RECT 64.13 4.866 64.21 5.098 ;
      RECT 64.065 4.862 64.13 5.127 ;
      RECT 64.06 4.576 64.065 4.6 ;
      RECT 64.05 4.852 64.065 5.155 ;
      RECT 64.055 4.57 64.06 4.64 ;
      RECT 64.05 4.564 64.055 4.71 ;
      RECT 64.045 4.558 64.05 4.788 ;
      RECT 64.045 4.835 64.05 5.22 ;
      RECT 64.037 4.555 64.045 5.22 ;
      RECT 63.951 4.553 64.037 5.22 ;
      RECT 63.865 4.551 63.951 5.22 ;
      RECT 63.855 4.552 63.865 5.22 ;
      RECT 63.85 4.557 63.855 5.22 ;
      RECT 63.84 4.57 63.85 5.22 ;
      RECT 63.835 4.592 63.84 5.22 ;
      RECT 63.83 4.952 63.835 5.22 ;
      RECT 64.46 4.42 64.465 4.64 ;
      RECT 64.965 3.455 65 3.715 ;
      RECT 64.95 3.455 64.965 3.723 ;
      RECT 64.921 3.455 64.95 3.745 ;
      RECT 64.835 3.455 64.921 3.805 ;
      RECT 64.815 3.455 64.835 3.87 ;
      RECT 64.755 3.455 64.815 4.035 ;
      RECT 64.75 3.455 64.755 4.183 ;
      RECT 64.745 3.455 64.75 4.195 ;
      RECT 64.74 3.455 64.745 4.221 ;
      RECT 64.71 3.641 64.74 4.301 ;
      RECT 64.705 3.689 64.71 4.39 ;
      RECT 64.7 3.703 64.705 4.405 ;
      RECT 64.695 3.722 64.7 4.435 ;
      RECT 64.69 3.737 64.695 4.451 ;
      RECT 64.685 3.752 64.69 4.473 ;
      RECT 64.68 3.772 64.685 4.495 ;
      RECT 64.67 3.792 64.68 4.528 ;
      RECT 64.655 3.834 64.67 4.59 ;
      RECT 64.65 3.865 64.655 4.63 ;
      RECT 64.645 3.877 64.65 4.635 ;
      RECT 64.64 3.889 64.645 4.64 ;
      RECT 64.635 3.902 64.64 4.64 ;
      RECT 64.63 3.92 64.635 4.64 ;
      RECT 64.625 3.94 64.63 4.64 ;
      RECT 64.62 3.952 64.625 4.64 ;
      RECT 64.615 3.965 64.62 4.64 ;
      RECT 64.595 4 64.615 4.64 ;
      RECT 64.545 4.102 64.595 4.64 ;
      RECT 64.54 4.187 64.545 4.64 ;
      RECT 64.535 4.195 64.54 4.64 ;
      RECT 64.53 4.212 64.535 4.64 ;
      RECT 64.525 4.227 64.53 4.64 ;
      RECT 64.49 4.292 64.525 4.64 ;
      RECT 64.475 4.357 64.49 4.64 ;
      RECT 64.47 4.387 64.475 4.64 ;
      RECT 64.465 4.412 64.47 4.64 ;
      RECT 64.45 4.422 64.46 4.64 ;
      RECT 64.435 4.435 64.45 4.633 ;
      RECT 64.18 4.025 64.25 4.235 ;
      RECT 63.97 4.002 63.975 4.195 ;
      RECT 61.425 3.93 61.685 4.19 ;
      RECT 64.26 4.212 64.265 4.215 ;
      RECT 64.25 4.03 64.26 4.23 ;
      RECT 64.151 4.023 64.18 4.235 ;
      RECT 64.065 4.015 64.151 4.235 ;
      RECT 64.05 4.009 64.065 4.233 ;
      RECT 64.03 4.008 64.05 4.22 ;
      RECT 64.025 4.007 64.03 4.203 ;
      RECT 63.975 4.004 64.025 4.198 ;
      RECT 63.945 4.001 63.97 4.193 ;
      RECT 63.925 3.999 63.945 4.188 ;
      RECT 63.91 3.997 63.925 4.185 ;
      RECT 63.88 3.995 63.91 4.183 ;
      RECT 63.815 3.991 63.88 4.175 ;
      RECT 63.785 3.986 63.815 4.17 ;
      RECT 63.765 3.984 63.785 4.168 ;
      RECT 63.735 3.981 63.765 4.163 ;
      RECT 63.675 3.977 63.735 4.155 ;
      RECT 63.67 3.974 63.675 4.15 ;
      RECT 63.6 3.972 63.67 4.145 ;
      RECT 63.571 3.968 63.6 4.138 ;
      RECT 63.485 3.963 63.571 4.13 ;
      RECT 63.451 3.958 63.485 4.122 ;
      RECT 63.365 3.95 63.451 4.114 ;
      RECT 63.326 3.943 63.365 4.106 ;
      RECT 63.24 3.938 63.326 4.098 ;
      RECT 63.175 3.932 63.24 4.088 ;
      RECT 63.155 3.927 63.175 4.083 ;
      RECT 63.146 3.924 63.155 4.082 ;
      RECT 63.06 3.92 63.146 4.076 ;
      RECT 63.02 3.916 63.06 4.068 ;
      RECT 63 3.912 63.02 4.066 ;
      RECT 62.94 3.912 63 4.063 ;
      RECT 62.92 3.915 62.94 4.061 ;
      RECT 62.899 3.915 62.92 4.061 ;
      RECT 62.813 3.917 62.899 4.065 ;
      RECT 62.727 3.919 62.813 4.071 ;
      RECT 62.641 3.921 62.727 4.078 ;
      RECT 62.555 3.924 62.641 4.084 ;
      RECT 62.521 3.925 62.555 4.089 ;
      RECT 62.435 3.928 62.521 4.094 ;
      RECT 62.406 3.935 62.435 4.099 ;
      RECT 62.32 3.935 62.406 4.104 ;
      RECT 62.287 3.935 62.32 4.109 ;
      RECT 62.201 3.937 62.287 4.114 ;
      RECT 62.115 3.939 62.201 4.121 ;
      RECT 62.051 3.941 62.115 4.127 ;
      RECT 61.965 3.943 62.051 4.133 ;
      RECT 61.962 3.945 61.965 4.136 ;
      RECT 61.876 3.946 61.962 4.14 ;
      RECT 61.79 3.949 61.876 4.147 ;
      RECT 61.771 3.951 61.79 4.151 ;
      RECT 61.685 3.953 61.771 4.156 ;
      RECT 61.415 3.965 61.425 4.16 ;
      RECT 63.585 10.205 63.875 10.435 ;
      RECT 63.645 9.465 63.815 10.435 ;
      RECT 63.535 9.49 63.91 9.86 ;
      RECT 63.585 9.465 63.875 9.86 ;
      RECT 63.65 3.545 63.835 3.755 ;
      RECT 63.645 3.546 63.84 3.753 ;
      RECT 63.64 3.551 63.85 3.748 ;
      RECT 63.635 3.527 63.64 3.745 ;
      RECT 63.605 3.524 63.635 3.738 ;
      RECT 63.6 3.52 63.605 3.729 ;
      RECT 63.565 3.551 63.85 3.724 ;
      RECT 63.34 3.46 63.6 3.72 ;
      RECT 63.64 3.529 63.645 3.748 ;
      RECT 63.645 3.53 63.65 3.753 ;
      RECT 63.34 3.542 63.72 3.72 ;
      RECT 63.34 3.54 63.705 3.72 ;
      RECT 63.34 3.535 63.695 3.72 ;
      RECT 63.295 4.45 63.345 4.735 ;
      RECT 63.24 4.42 63.245 4.735 ;
      RECT 63.21 4.4 63.215 4.735 ;
      RECT 63.36 4.45 63.42 4.71 ;
      RECT 63.355 4.45 63.36 4.718 ;
      RECT 63.345 4.45 63.355 4.73 ;
      RECT 63.26 4.44 63.295 4.735 ;
      RECT 63.255 4.427 63.26 4.735 ;
      RECT 63.245 4.422 63.255 4.735 ;
      RECT 63.225 4.412 63.24 4.735 ;
      RECT 63.215 4.405 63.225 4.735 ;
      RECT 63.205 4.397 63.21 4.735 ;
      RECT 63.175 4.387 63.205 4.735 ;
      RECT 63.16 4.375 63.175 4.735 ;
      RECT 63.145 4.365 63.16 4.73 ;
      RECT 63.125 4.355 63.145 4.705 ;
      RECT 63.115 4.347 63.125 4.682 ;
      RECT 63.085 4.33 63.115 4.672 ;
      RECT 63.08 4.307 63.085 4.663 ;
      RECT 63.075 4.294 63.08 4.661 ;
      RECT 63.06 4.27 63.075 4.655 ;
      RECT 63.055 4.246 63.06 4.649 ;
      RECT 63.045 4.235 63.055 4.644 ;
      RECT 63.04 4.225 63.045 4.64 ;
      RECT 63.035 4.217 63.04 4.637 ;
      RECT 63.025 4.212 63.035 4.633 ;
      RECT 63.02 4.207 63.025 4.629 ;
      RECT 62.935 4.205 63.02 4.604 ;
      RECT 62.905 4.205 62.935 4.57 ;
      RECT 62.89 4.205 62.905 4.553 ;
      RECT 62.835 4.205 62.89 4.498 ;
      RECT 62.83 4.21 62.835 4.447 ;
      RECT 62.82 4.215 62.83 4.437 ;
      RECT 62.815 4.225 62.82 4.423 ;
      RECT 62.765 4.965 63.025 5.225 ;
      RECT 62.685 4.98 63.025 5.201 ;
      RECT 62.665 4.98 63.025 5.196 ;
      RECT 62.641 4.98 63.025 5.194 ;
      RECT 62.555 4.98 63.025 5.189 ;
      RECT 62.405 4.92 62.665 5.185 ;
      RECT 62.36 4.98 63.025 5.18 ;
      RECT 62.355 4.987 63.025 5.175 ;
      RECT 62.37 4.975 62.685 5.185 ;
      RECT 62.26 3.41 62.52 3.67 ;
      RECT 62.26 3.467 62.525 3.663 ;
      RECT 62.26 3.497 62.53 3.595 ;
      RECT 62.32 3.928 62.435 3.93 ;
      RECT 62.406 3.925 62.435 3.93 ;
      RECT 61.43 4.929 61.455 5.169 ;
      RECT 61.415 4.932 61.505 5.163 ;
      RECT 61.41 4.937 61.591 5.158 ;
      RECT 61.405 4.945 61.655 5.156 ;
      RECT 61.405 4.945 61.665 5.155 ;
      RECT 61.4 4.952 61.675 5.148 ;
      RECT 61.4 4.952 61.761 5.137 ;
      RECT 61.395 4.987 61.761 5.133 ;
      RECT 61.395 4.987 61.77 5.122 ;
      RECT 61.675 4.86 61.935 5.12 ;
      RECT 61.385 5.037 61.935 5.118 ;
      RECT 61.655 4.905 61.675 5.153 ;
      RECT 61.591 4.908 61.655 5.157 ;
      RECT 61.505 4.913 61.591 5.162 ;
      RECT 61.435 4.924 61.935 5.12 ;
      RECT 61.455 4.918 61.505 5.167 ;
      RECT 61.58 3.395 61.59 3.657 ;
      RECT 61.57 3.452 61.58 3.66 ;
      RECT 61.545 3.457 61.57 3.666 ;
      RECT 61.52 3.461 61.545 3.678 ;
      RECT 61.51 3.464 61.52 3.688 ;
      RECT 61.505 3.465 61.51 3.693 ;
      RECT 61.5 3.466 61.505 3.698 ;
      RECT 61.495 3.467 61.5 3.7 ;
      RECT 61.47 3.47 61.495 3.703 ;
      RECT 61.44 3.476 61.47 3.706 ;
      RECT 61.375 3.487 61.44 3.709 ;
      RECT 61.33 3.495 61.375 3.713 ;
      RECT 61.315 3.495 61.33 3.721 ;
      RECT 61.31 3.496 61.315 3.728 ;
      RECT 61.305 3.498 61.31 3.731 ;
      RECT 61.3 3.502 61.305 3.734 ;
      RECT 61.29 3.51 61.3 3.738 ;
      RECT 61.285 3.523 61.29 3.743 ;
      RECT 61.28 3.531 61.285 3.745 ;
      RECT 61.275 3.537 61.28 3.745 ;
      RECT 61.27 3.541 61.275 3.748 ;
      RECT 61.265 3.543 61.27 3.751 ;
      RECT 61.26 3.546 61.265 3.754 ;
      RECT 61.25 3.551 61.26 3.758 ;
      RECT 61.245 3.557 61.25 3.763 ;
      RECT 61.235 3.563 61.245 3.767 ;
      RECT 61.22 3.57 61.235 3.773 ;
      RECT 61.191 3.584 61.22 3.783 ;
      RECT 61.105 3.619 61.191 3.815 ;
      RECT 61.085 3.652 61.105 3.844 ;
      RECT 61.065 3.665 61.085 3.855 ;
      RECT 61.045 3.677 61.065 3.866 ;
      RECT 60.995 3.699 61.045 3.886 ;
      RECT 60.98 3.717 60.995 3.903 ;
      RECT 60.975 3.723 60.98 3.906 ;
      RECT 60.97 3.727 60.975 3.909 ;
      RECT 60.965 3.731 60.97 3.913 ;
      RECT 60.96 3.733 60.965 3.916 ;
      RECT 60.95 3.74 60.96 3.919 ;
      RECT 60.945 3.745 60.95 3.923 ;
      RECT 60.94 3.747 60.945 3.926 ;
      RECT 60.935 3.751 60.94 3.929 ;
      RECT 60.93 3.753 60.935 3.933 ;
      RECT 60.915 3.758 60.93 3.938 ;
      RECT 60.91 3.763 60.915 3.941 ;
      RECT 60.905 3.771 60.91 3.944 ;
      RECT 60.9 3.773 60.905 3.947 ;
      RECT 60.895 3.775 60.9 3.95 ;
      RECT 60.885 3.777 60.895 3.956 ;
      RECT 60.85 3.791 60.885 3.968 ;
      RECT 60.84 3.806 60.85 3.978 ;
      RECT 60.765 3.835 60.84 4.002 ;
      RECT 60.76 3.86 60.765 4.025 ;
      RECT 60.745 3.864 60.76 4.031 ;
      RECT 60.735 3.872 60.745 4.036 ;
      RECT 60.705 3.885 60.735 4.04 ;
      RECT 60.695 3.9 60.705 4.045 ;
      RECT 60.685 3.905 60.695 4.048 ;
      RECT 60.68 3.907 60.685 4.05 ;
      RECT 60.665 3.91 60.68 4.053 ;
      RECT 60.66 3.912 60.665 4.056 ;
      RECT 60.64 3.917 60.66 4.06 ;
      RECT 60.61 3.922 60.64 4.068 ;
      RECT 60.585 3.929 60.61 4.076 ;
      RECT 60.58 3.934 60.585 4.081 ;
      RECT 60.55 3.937 60.58 4.085 ;
      RECT 60.51 3.94 60.55 4.095 ;
      RECT 60.475 3.937 60.51 4.107 ;
      RECT 60.465 3.933 60.475 4.114 ;
      RECT 60.44 3.929 60.465 4.12 ;
      RECT 60.435 3.925 60.44 4.125 ;
      RECT 60.395 3.922 60.435 4.125 ;
      RECT 60.38 3.907 60.395 4.126 ;
      RECT 60.357 3.895 60.38 4.126 ;
      RECT 60.271 3.895 60.357 4.127 ;
      RECT 60.185 3.895 60.271 4.129 ;
      RECT 60.165 3.895 60.185 4.126 ;
      RECT 60.16 3.9 60.165 4.121 ;
      RECT 60.155 3.905 60.16 4.119 ;
      RECT 60.145 3.915 60.155 4.117 ;
      RECT 60.14 3.921 60.145 4.11 ;
      RECT 60.135 3.923 60.14 4.095 ;
      RECT 60.13 3.927 60.135 4.085 ;
      RECT 61.59 3.395 61.84 3.655 ;
      RECT 59.315 4.93 59.575 5.19 ;
      RECT 61.61 4.42 61.615 4.63 ;
      RECT 61.615 4.425 61.625 4.625 ;
      RECT 61.565 4.42 61.61 4.645 ;
      RECT 61.555 4.42 61.565 4.665 ;
      RECT 61.536 4.42 61.555 4.67 ;
      RECT 61.45 4.42 61.536 4.667 ;
      RECT 61.42 4.422 61.45 4.665 ;
      RECT 61.365 4.432 61.42 4.663 ;
      RECT 61.3 4.446 61.365 4.661 ;
      RECT 61.295 4.454 61.3 4.66 ;
      RECT 61.28 4.457 61.295 4.658 ;
      RECT 61.215 4.467 61.28 4.654 ;
      RECT 61.167 4.481 61.215 4.655 ;
      RECT 61.081 4.498 61.167 4.669 ;
      RECT 60.995 4.519 61.081 4.686 ;
      RECT 60.975 4.532 60.995 4.696 ;
      RECT 60.93 4.54 60.975 4.703 ;
      RECT 60.895 4.548 60.93 4.711 ;
      RECT 60.861 4.556 60.895 4.719 ;
      RECT 60.775 4.57 60.861 4.731 ;
      RECT 60.74 4.587 60.775 4.743 ;
      RECT 60.731 4.596 60.74 4.747 ;
      RECT 60.645 4.614 60.731 4.764 ;
      RECT 60.586 4.641 60.645 4.791 ;
      RECT 60.5 4.668 60.586 4.819 ;
      RECT 60.48 4.69 60.5 4.839 ;
      RECT 60.42 4.705 60.48 4.855 ;
      RECT 60.41 4.717 60.42 4.868 ;
      RECT 60.405 4.722 60.41 4.871 ;
      RECT 60.395 4.725 60.405 4.874 ;
      RECT 60.39 4.727 60.395 4.877 ;
      RECT 60.36 4.735 60.39 4.884 ;
      RECT 60.345 4.742 60.36 4.892 ;
      RECT 60.335 4.747 60.345 4.896 ;
      RECT 60.33 4.75 60.335 4.899 ;
      RECT 60.32 4.752 60.33 4.902 ;
      RECT 60.285 4.762 60.32 4.911 ;
      RECT 60.21 4.785 60.285 4.933 ;
      RECT 60.19 4.803 60.21 4.951 ;
      RECT 60.16 4.81 60.19 4.961 ;
      RECT 60.14 4.818 60.16 4.971 ;
      RECT 60.13 4.824 60.14 4.978 ;
      RECT 60.111 4.829 60.13 4.984 ;
      RECT 60.025 4.849 60.111 5.004 ;
      RECT 60.01 4.869 60.025 5.023 ;
      RECT 59.965 4.881 60.01 5.034 ;
      RECT 59.9 4.902 59.965 5.057 ;
      RECT 59.86 4.922 59.9 5.078 ;
      RECT 59.85 4.932 59.86 5.088 ;
      RECT 59.8 4.944 59.85 5.099 ;
      RECT 59.78 4.96 59.8 5.111 ;
      RECT 59.75 4.97 59.78 5.117 ;
      RECT 59.74 4.975 59.75 5.119 ;
      RECT 59.671 4.976 59.74 5.125 ;
      RECT 59.585 4.978 59.671 5.135 ;
      RECT 59.575 4.979 59.585 5.14 ;
      RECT 60.845 5.005 61.035 5.215 ;
      RECT 60.835 5.01 61.045 5.208 ;
      RECT 60.82 5.01 61.045 5.173 ;
      RECT 60.74 4.895 61 5.155 ;
      RECT 59.655 4.425 59.84 4.72 ;
      RECT 59.645 4.425 59.84 4.718 ;
      RECT 59.63 4.425 59.845 4.713 ;
      RECT 59.63 4.425 59.85 4.71 ;
      RECT 59.625 4.425 59.85 4.708 ;
      RECT 59.62 4.68 59.85 4.698 ;
      RECT 59.625 4.425 59.885 4.685 ;
      RECT 59.585 3.46 59.845 3.72 ;
      RECT 59.395 3.385 59.481 3.718 ;
      RECT 59.37 3.389 59.525 3.714 ;
      RECT 59.481 3.381 59.525 3.714 ;
      RECT 59.481 3.382 59.53 3.713 ;
      RECT 59.395 3.387 59.545 3.712 ;
      RECT 59.37 3.395 59.585 3.711 ;
      RECT 59.365 3.39 59.545 3.706 ;
      RECT 59.355 3.405 59.585 3.613 ;
      RECT 59.355 3.457 59.785 3.613 ;
      RECT 59.355 3.45 59.765 3.613 ;
      RECT 59.355 3.437 59.735 3.613 ;
      RECT 59.355 3.425 59.675 3.613 ;
      RECT 59.355 3.41 59.65 3.613 ;
      RECT 58.555 4.04 58.69 4.335 ;
      RECT 58.815 4.063 58.82 4.25 ;
      RECT 59.535 3.96 59.68 4.195 ;
      RECT 59.695 3.96 59.7 4.185 ;
      RECT 59.73 3.971 59.735 4.165 ;
      RECT 59.725 3.963 59.73 4.17 ;
      RECT 59.705 3.96 59.725 4.175 ;
      RECT 59.7 3.96 59.705 4.183 ;
      RECT 59.69 3.96 59.695 4.188 ;
      RECT 59.68 3.96 59.69 4.193 ;
      RECT 59.51 3.962 59.535 4.195 ;
      RECT 59.46 3.969 59.51 4.195 ;
      RECT 59.455 3.974 59.46 4.195 ;
      RECT 59.416 3.979 59.455 4.196 ;
      RECT 59.33 3.991 59.416 4.197 ;
      RECT 59.321 4.001 59.33 4.197 ;
      RECT 59.235 4.01 59.321 4.199 ;
      RECT 59.211 4.02 59.235 4.201 ;
      RECT 59.125 4.031 59.211 4.202 ;
      RECT 59.095 4.042 59.125 4.204 ;
      RECT 59.065 4.047 59.095 4.206 ;
      RECT 59.04 4.053 59.065 4.209 ;
      RECT 59.025 4.058 59.04 4.21 ;
      RECT 58.98 4.064 59.025 4.21 ;
      RECT 58.975 4.069 58.98 4.211 ;
      RECT 58.955 4.069 58.975 4.213 ;
      RECT 58.935 4.067 58.955 4.218 ;
      RECT 58.9 4.066 58.935 4.225 ;
      RECT 58.87 4.065 58.9 4.235 ;
      RECT 58.82 4.064 58.87 4.245 ;
      RECT 58.73 4.061 58.815 4.335 ;
      RECT 58.705 4.055 58.73 4.335 ;
      RECT 58.69 4.045 58.705 4.335 ;
      RECT 58.505 4.04 58.555 4.255 ;
      RECT 58.495 4.045 58.505 4.245 ;
      RECT 58.735 4.52 58.995 4.78 ;
      RECT 58.735 4.52 59.025 4.673 ;
      RECT 58.735 4.52 59.06 4.658 ;
      RECT 58.99 4.44 59.18 4.65 ;
      RECT 58.98 4.445 59.19 4.643 ;
      RECT 58.945 4.515 59.19 4.643 ;
      RECT 58.975 4.457 58.995 4.78 ;
      RECT 58.96 4.505 59.19 4.643 ;
      RECT 58.965 4.477 58.995 4.78 ;
      RECT 58.045 3.545 58.115 4.65 ;
      RECT 58.78 3.65 59.04 3.91 ;
      RECT 58.36 3.696 58.375 3.905 ;
      RECT 58.696 3.709 58.78 3.86 ;
      RECT 58.61 3.706 58.696 3.86 ;
      RECT 58.571 3.704 58.61 3.86 ;
      RECT 58.485 3.702 58.571 3.86 ;
      RECT 58.425 3.7 58.485 3.871 ;
      RECT 58.39 3.698 58.425 3.889 ;
      RECT 58.375 3.696 58.39 3.9 ;
      RECT 58.345 3.696 58.36 3.913 ;
      RECT 58.335 3.696 58.345 3.918 ;
      RECT 58.31 3.695 58.335 3.923 ;
      RECT 58.295 3.69 58.31 3.929 ;
      RECT 58.29 3.683 58.295 3.934 ;
      RECT 58.265 3.674 58.29 3.94 ;
      RECT 58.22 3.653 58.265 3.953 ;
      RECT 58.21 3.637 58.22 3.963 ;
      RECT 58.195 3.63 58.21 3.973 ;
      RECT 58.185 3.623 58.195 3.99 ;
      RECT 58.18 3.62 58.185 4.02 ;
      RECT 58.175 3.618 58.18 4.05 ;
      RECT 58.17 3.616 58.175 4.087 ;
      RECT 58.155 3.612 58.17 4.154 ;
      RECT 58.155 4.445 58.165 4.645 ;
      RECT 58.15 3.608 58.155 4.28 ;
      RECT 58.15 4.432 58.155 4.65 ;
      RECT 58.145 3.606 58.15 4.365 ;
      RECT 58.145 4.422 58.15 4.65 ;
      RECT 58.13 3.577 58.145 4.65 ;
      RECT 58.115 3.55 58.13 4.65 ;
      RECT 58.04 3.545 58.045 3.9 ;
      RECT 58.04 3.955 58.045 4.65 ;
      RECT 58.025 3.545 58.04 3.878 ;
      RECT 58.035 3.977 58.04 4.65 ;
      RECT 58.025 4.017 58.035 4.65 ;
      RECT 57.99 3.545 58.025 3.82 ;
      RECT 58.02 4.052 58.025 4.65 ;
      RECT 58.005 4.107 58.02 4.65 ;
      RECT 58 4.172 58.005 4.65 ;
      RECT 57.985 4.22 58 4.65 ;
      RECT 57.96 3.545 57.99 3.775 ;
      RECT 57.98 4.275 57.985 4.65 ;
      RECT 57.965 4.335 57.98 4.65 ;
      RECT 57.96 4.383 57.965 4.648 ;
      RECT 57.955 3.545 57.96 3.768 ;
      RECT 57.955 4.415 57.96 4.643 ;
      RECT 57.93 3.545 57.955 3.76 ;
      RECT 57.92 3.55 57.93 3.75 ;
      RECT 58.135 4.825 58.155 5.065 ;
      RECT 57.365 4.755 57.37 4.965 ;
      RECT 58.645 4.828 58.655 5.023 ;
      RECT 58.64 4.818 58.645 5.026 ;
      RECT 58.56 4.815 58.64 5.049 ;
      RECT 58.556 4.815 58.56 5.071 ;
      RECT 58.47 4.815 58.556 5.081 ;
      RECT 58.455 4.815 58.47 5.089 ;
      RECT 58.426 4.816 58.455 5.087 ;
      RECT 58.34 4.821 58.426 5.083 ;
      RECT 58.327 4.825 58.34 5.079 ;
      RECT 58.241 4.825 58.327 5.075 ;
      RECT 58.155 4.825 58.241 5.069 ;
      RECT 58.071 4.825 58.135 5.063 ;
      RECT 57.985 4.825 58.071 5.058 ;
      RECT 57.965 4.825 57.985 5.054 ;
      RECT 57.905 4.82 57.965 5.051 ;
      RECT 57.877 4.814 57.905 5.048 ;
      RECT 57.791 4.809 57.877 5.044 ;
      RECT 57.705 4.803 57.791 5.038 ;
      RECT 57.63 4.785 57.705 5.033 ;
      RECT 57.595 4.762 57.63 5.029 ;
      RECT 57.585 4.752 57.595 5.028 ;
      RECT 57.53 4.75 57.585 5.027 ;
      RECT 57.455 4.75 57.53 5.023 ;
      RECT 57.445 4.75 57.455 5.018 ;
      RECT 57.43 4.75 57.445 5.01 ;
      RECT 57.38 4.752 57.43 4.988 ;
      RECT 57.37 4.755 57.38 4.968 ;
      RECT 57.36 4.76 57.365 4.963 ;
      RECT 57.355 4.765 57.36 4.958 ;
      RECT 55.465 3.41 55.725 3.67 ;
      RECT 55.455 3.44 55.725 3.65 ;
      RECT 57.375 3.355 57.635 3.615 ;
      RECT 57.37 3.43 57.375 3.616 ;
      RECT 57.345 3.435 57.37 3.618 ;
      RECT 57.33 3.442 57.345 3.621 ;
      RECT 57.27 3.46 57.33 3.626 ;
      RECT 57.24 3.48 57.27 3.633 ;
      RECT 57.215 3.488 57.24 3.638 ;
      RECT 57.19 3.496 57.215 3.64 ;
      RECT 57.172 3.5 57.19 3.639 ;
      RECT 57.086 3.498 57.172 3.639 ;
      RECT 57 3.496 57.086 3.639 ;
      RECT 56.914 3.494 57 3.638 ;
      RECT 56.828 3.492 56.914 3.638 ;
      RECT 56.742 3.49 56.828 3.638 ;
      RECT 56.656 3.488 56.742 3.638 ;
      RECT 56.57 3.486 56.656 3.637 ;
      RECT 56.552 3.485 56.57 3.637 ;
      RECT 56.466 3.484 56.552 3.637 ;
      RECT 56.38 3.482 56.466 3.637 ;
      RECT 56.294 3.481 56.38 3.636 ;
      RECT 56.208 3.48 56.294 3.636 ;
      RECT 56.122 3.478 56.208 3.636 ;
      RECT 56.036 3.477 56.122 3.636 ;
      RECT 55.95 3.475 56.036 3.635 ;
      RECT 55.926 3.473 55.95 3.635 ;
      RECT 55.84 3.466 55.926 3.635 ;
      RECT 55.811 3.458 55.84 3.635 ;
      RECT 55.725 3.45 55.811 3.635 ;
      RECT 55.445 3.447 55.455 3.645 ;
      RECT 56.95 4.41 56.955 4.76 ;
      RECT 56.72 4.5 56.86 4.76 ;
      RECT 57.195 4.185 57.24 4.395 ;
      RECT 57.25 4.196 57.26 4.39 ;
      RECT 57.24 4.188 57.25 4.395 ;
      RECT 57.175 4.185 57.195 4.4 ;
      RECT 57.145 4.185 57.175 4.423 ;
      RECT 57.135 4.185 57.145 4.448 ;
      RECT 57.13 4.185 57.135 4.458 ;
      RECT 57.075 4.185 57.13 4.498 ;
      RECT 57.07 4.185 57.075 4.538 ;
      RECT 57.065 4.187 57.07 4.543 ;
      RECT 57.05 4.197 57.065 4.554 ;
      RECT 57.005 4.255 57.05 4.59 ;
      RECT 56.995 4.31 57.005 4.624 ;
      RECT 56.98 4.337 56.995 4.64 ;
      RECT 56.97 4.364 56.98 4.76 ;
      RECT 56.955 4.387 56.97 4.76 ;
      RECT 56.945 4.427 56.95 4.76 ;
      RECT 56.94 4.437 56.945 4.76 ;
      RECT 56.935 4.452 56.94 4.76 ;
      RECT 56.925 4.457 56.935 4.76 ;
      RECT 56.86 4.48 56.925 4.76 ;
      RECT 56.33 3.875 56.56 4.185 ;
      RECT 56.23 3.875 56.56 4.165 ;
      RECT 54.935 3.9 55.195 4.16 ;
      RECT 56.06 3.875 56.56 4.155 ;
      RECT 55.875 3.875 56.56 4.145 ;
      RECT 55.69 3.925 56.56 4.135 ;
      RECT 55.57 3.925 56.56 4.125 ;
      RECT 55.24 3.925 56.56 4.115 ;
      RECT 55.235 3.925 56.56 4.101 ;
      RECT 54.935 3.915 55.52 4.098 ;
      RECT 55.805 3.875 56.62 4.015 ;
      RECT 55.24 3.91 55.51 4.115 ;
      RECT 55.24 3.895 55.5 4.115 ;
      RECT 55.45 4.415 55.71 4.675 ;
      RECT 55.45 4.455 55.815 4.665 ;
      RECT 55.45 4.457 55.82 4.664 ;
      RECT 55.45 4.465 55.825 4.661 ;
      RECT 54.375 3.54 54.475 5.065 ;
      RECT 54.565 4.68 54.615 4.94 ;
      RECT 54.56 3.553 54.565 3.74 ;
      RECT 54.555 4.661 54.565 4.94 ;
      RECT 54.555 3.55 54.56 3.748 ;
      RECT 54.54 3.544 54.555 3.755 ;
      RECT 54.55 4.649 54.555 5.023 ;
      RECT 54.54 4.637 54.55 5.06 ;
      RECT 54.53 3.54 54.54 3.762 ;
      RECT 54.53 4.622 54.54 5.065 ;
      RECT 54.525 3.54 54.53 3.77 ;
      RECT 54.505 4.592 54.53 5.065 ;
      RECT 54.485 3.54 54.525 3.818 ;
      RECT 54.495 4.552 54.505 5.065 ;
      RECT 54.485 4.507 54.495 5.065 ;
      RECT 54.48 3.54 54.485 3.888 ;
      RECT 54.48 4.465 54.485 5.065 ;
      RECT 54.475 3.54 54.48 4.365 ;
      RECT 54.475 4.447 54.48 5.065 ;
      RECT 54.365 3.543 54.375 5.065 ;
      RECT 54.35 3.55 54.365 5.061 ;
      RECT 54.345 3.56 54.35 5.056 ;
      RECT 54.34 3.76 54.345 4.948 ;
      RECT 54.335 3.845 54.34 4.5 ;
      RECT 53.2 10.205 53.495 10.435 ;
      RECT 53.26 8.725 53.43 10.435 ;
      RECT 53.25 9.095 53.605 9.45 ;
      RECT 53.2 8.725 53.49 8.955 ;
      RECT 52.21 10.205 52.505 10.435 ;
      RECT 52.27 8.725 52.44 10.435 ;
      RECT 52.21 8.725 52.5 8.955 ;
      RECT 52.21 8.76 53.06 8.92 ;
      RECT 52.895 8.355 53.06 8.92 ;
      RECT 52.21 8.755 52.605 8.92 ;
      RECT 52.83 8.355 53.12 8.585 ;
      RECT 52.83 8.385 53.29 8.555 ;
      RECT 52.795 4.025 53.12 4.26 ;
      RECT 52.795 4.055 53.285 4.225 ;
      RECT 52.795 3.69 52.985 4.26 ;
      RECT 52.21 3.655 52.5 3.885 ;
      RECT 52.21 3.69 52.985 3.86 ;
      RECT 52.27 2.175 52.44 3.885 ;
      RECT 52.21 2.175 52.505 2.405 ;
      RECT 51.84 4.025 52.13 4.255 ;
      RECT 51.84 4.055 52.3 4.225 ;
      RECT 51.905 2.95 52.07 4.255 ;
      RECT 50.42 2.915 50.71 3.145 ;
      RECT 50.42 2.95 52.07 3.12 ;
      RECT 50.48 2.175 50.65 3.145 ;
      RECT 50.42 2.175 50.71 2.405 ;
      RECT 50.42 10.205 50.71 10.435 ;
      RECT 50.48 9.465 50.65 10.435 ;
      RECT 50.48 9.555 52.07 9.725 ;
      RECT 51.9 8.355 52.07 9.725 ;
      RECT 50.42 9.465 50.71 9.695 ;
      RECT 51.84 8.355 52.13 8.585 ;
      RECT 51.84 8.385 52.3 8.555 ;
      RECT 48.455 4.725 48.805 5.075 ;
      RECT 48.545 3.32 48.715 5.075 ;
      RECT 50.85 3.26 51.2 3.61 ;
      RECT 48.545 3.32 50.165 3.495 ;
      RECT 48.545 3.32 50.82 3.49 ;
      RECT 50.68 3.315 51.2 3.485 ;
      RECT 50.875 9.09 51.2 9.415 ;
      RECT 46.3 9.05 46.65 9.4 ;
      RECT 50.85 9.095 51.2 9.325 ;
      RECT 46.09 9.095 46.65 9.325 ;
      RECT 50.68 9.12 51.2 9.295 ;
      RECT 45.92 9.125 46.65 9.295 ;
      RECT 46.09 9.12 51.2 9.29 ;
      RECT 50.075 3.66 50.395 3.98 ;
      RECT 50.05 3.655 50.34 3.885 ;
      RECT 50.005 3.685 50.395 3.86 ;
      RECT 49.875 3.685 50.395 3.855 ;
      RECT 50.075 8.66 50.395 8.98 ;
      RECT 50.05 8.725 50.395 8.955 ;
      RECT 49.875 8.755 50.395 8.925 ;
      RECT 45.865 4.96 45.905 5.22 ;
      RECT 45.905 4.94 45.91 4.95 ;
      RECT 47.235 4.185 47.245 4.406 ;
      RECT 47.165 4.18 47.235 4.531 ;
      RECT 47.155 4.18 47.165 4.658 ;
      RECT 47.13 4.18 47.155 4.705 ;
      RECT 47.105 4.18 47.13 4.783 ;
      RECT 47.085 4.18 47.105 4.853 ;
      RECT 47.06 4.18 47.085 4.893 ;
      RECT 47.05 4.18 47.06 4.913 ;
      RECT 47.04 4.182 47.05 4.921 ;
      RECT 47.035 4.187 47.04 4.378 ;
      RECT 47.035 4.387 47.04 4.922 ;
      RECT 47.03 4.432 47.035 4.923 ;
      RECT 47.02 4.497 47.03 4.924 ;
      RECT 47.01 4.592 47.02 4.926 ;
      RECT 47.005 4.645 47.01 4.928 ;
      RECT 47 4.665 47.005 4.929 ;
      RECT 46.945 4.69 47 4.935 ;
      RECT 46.905 4.725 46.945 4.944 ;
      RECT 46.895 4.742 46.905 4.949 ;
      RECT 46.886 4.748 46.895 4.951 ;
      RECT 46.8 4.786 46.886 4.962 ;
      RECT 46.795 4.825 46.8 4.972 ;
      RECT 46.72 4.832 46.795 4.982 ;
      RECT 46.7 4.842 46.72 4.993 ;
      RECT 46.67 4.849 46.7 5.001 ;
      RECT 46.645 4.856 46.67 5.008 ;
      RECT 46.621 4.862 46.645 5.013 ;
      RECT 46.535 4.875 46.621 5.025 ;
      RECT 46.457 4.882 46.535 5.043 ;
      RECT 46.371 4.877 46.457 5.061 ;
      RECT 46.285 4.872 46.371 5.081 ;
      RECT 46.205 4.866 46.285 5.098 ;
      RECT 46.14 4.862 46.205 5.127 ;
      RECT 46.135 4.576 46.14 4.6 ;
      RECT 46.125 4.852 46.14 5.155 ;
      RECT 46.13 4.57 46.135 4.64 ;
      RECT 46.125 4.564 46.13 4.71 ;
      RECT 46.12 4.558 46.125 4.788 ;
      RECT 46.12 4.835 46.125 5.22 ;
      RECT 46.112 4.555 46.12 5.22 ;
      RECT 46.026 4.553 46.112 5.22 ;
      RECT 45.94 4.551 46.026 5.22 ;
      RECT 45.93 4.552 45.94 5.22 ;
      RECT 45.925 4.557 45.93 5.22 ;
      RECT 45.915 4.57 45.925 5.22 ;
      RECT 45.91 4.592 45.915 5.22 ;
      RECT 45.905 4.952 45.91 5.22 ;
      RECT 46.535 4.42 46.54 4.64 ;
      RECT 47.04 3.455 47.075 3.715 ;
      RECT 47.025 3.455 47.04 3.723 ;
      RECT 46.996 3.455 47.025 3.745 ;
      RECT 46.91 3.455 46.996 3.805 ;
      RECT 46.89 3.455 46.91 3.87 ;
      RECT 46.83 3.455 46.89 4.035 ;
      RECT 46.825 3.455 46.83 4.183 ;
      RECT 46.82 3.455 46.825 4.195 ;
      RECT 46.815 3.455 46.82 4.221 ;
      RECT 46.785 3.641 46.815 4.301 ;
      RECT 46.78 3.689 46.785 4.39 ;
      RECT 46.775 3.703 46.78 4.405 ;
      RECT 46.77 3.722 46.775 4.435 ;
      RECT 46.765 3.737 46.77 4.451 ;
      RECT 46.76 3.752 46.765 4.473 ;
      RECT 46.755 3.772 46.76 4.495 ;
      RECT 46.745 3.792 46.755 4.528 ;
      RECT 46.73 3.834 46.745 4.59 ;
      RECT 46.725 3.865 46.73 4.63 ;
      RECT 46.72 3.877 46.725 4.635 ;
      RECT 46.715 3.889 46.72 4.64 ;
      RECT 46.71 3.902 46.715 4.64 ;
      RECT 46.705 3.92 46.71 4.64 ;
      RECT 46.7 3.94 46.705 4.64 ;
      RECT 46.695 3.952 46.7 4.64 ;
      RECT 46.69 3.965 46.695 4.64 ;
      RECT 46.67 4 46.69 4.64 ;
      RECT 46.62 4.102 46.67 4.64 ;
      RECT 46.615 4.187 46.62 4.64 ;
      RECT 46.61 4.195 46.615 4.64 ;
      RECT 46.605 4.212 46.61 4.64 ;
      RECT 46.6 4.227 46.605 4.64 ;
      RECT 46.565 4.292 46.6 4.64 ;
      RECT 46.55 4.357 46.565 4.64 ;
      RECT 46.545 4.387 46.55 4.64 ;
      RECT 46.54 4.412 46.545 4.64 ;
      RECT 46.525 4.422 46.535 4.64 ;
      RECT 46.51 4.435 46.525 4.633 ;
      RECT 46.255 4.025 46.325 4.235 ;
      RECT 46.045 4.002 46.05 4.195 ;
      RECT 43.5 3.93 43.76 4.19 ;
      RECT 46.335 4.212 46.34 4.215 ;
      RECT 46.325 4.03 46.335 4.23 ;
      RECT 46.226 4.023 46.255 4.235 ;
      RECT 46.14 4.015 46.226 4.235 ;
      RECT 46.125 4.009 46.14 4.233 ;
      RECT 46.105 4.008 46.125 4.22 ;
      RECT 46.1 4.007 46.105 4.203 ;
      RECT 46.05 4.004 46.1 4.198 ;
      RECT 46.02 4.001 46.045 4.193 ;
      RECT 46 3.999 46.02 4.188 ;
      RECT 45.985 3.997 46 4.185 ;
      RECT 45.955 3.995 45.985 4.183 ;
      RECT 45.89 3.991 45.955 4.175 ;
      RECT 45.86 3.986 45.89 4.17 ;
      RECT 45.84 3.984 45.86 4.168 ;
      RECT 45.81 3.981 45.84 4.163 ;
      RECT 45.75 3.977 45.81 4.155 ;
      RECT 45.745 3.974 45.75 4.15 ;
      RECT 45.675 3.972 45.745 4.145 ;
      RECT 45.646 3.968 45.675 4.138 ;
      RECT 45.56 3.963 45.646 4.13 ;
      RECT 45.526 3.958 45.56 4.122 ;
      RECT 45.44 3.95 45.526 4.114 ;
      RECT 45.401 3.943 45.44 4.106 ;
      RECT 45.315 3.938 45.401 4.098 ;
      RECT 45.25 3.932 45.315 4.088 ;
      RECT 45.23 3.927 45.25 4.083 ;
      RECT 45.221 3.924 45.23 4.082 ;
      RECT 45.135 3.92 45.221 4.076 ;
      RECT 45.095 3.916 45.135 4.068 ;
      RECT 45.075 3.912 45.095 4.066 ;
      RECT 45.015 3.912 45.075 4.063 ;
      RECT 44.995 3.915 45.015 4.061 ;
      RECT 44.974 3.915 44.995 4.061 ;
      RECT 44.888 3.917 44.974 4.065 ;
      RECT 44.802 3.919 44.888 4.071 ;
      RECT 44.716 3.921 44.802 4.078 ;
      RECT 44.63 3.924 44.716 4.084 ;
      RECT 44.596 3.925 44.63 4.089 ;
      RECT 44.51 3.928 44.596 4.094 ;
      RECT 44.481 3.935 44.51 4.099 ;
      RECT 44.395 3.935 44.481 4.104 ;
      RECT 44.362 3.935 44.395 4.109 ;
      RECT 44.276 3.937 44.362 4.114 ;
      RECT 44.19 3.939 44.276 4.121 ;
      RECT 44.126 3.941 44.19 4.127 ;
      RECT 44.04 3.943 44.126 4.133 ;
      RECT 44.037 3.945 44.04 4.136 ;
      RECT 43.951 3.946 44.037 4.14 ;
      RECT 43.865 3.949 43.951 4.147 ;
      RECT 43.846 3.951 43.865 4.151 ;
      RECT 43.76 3.953 43.846 4.156 ;
      RECT 43.49 3.965 43.5 4.16 ;
      RECT 45.66 10.205 45.95 10.435 ;
      RECT 45.72 9.465 45.89 10.435 ;
      RECT 45.61 9.49 45.985 9.86 ;
      RECT 45.66 9.465 45.95 9.86 ;
      RECT 45.725 3.545 45.91 3.755 ;
      RECT 45.72 3.546 45.915 3.753 ;
      RECT 45.715 3.551 45.925 3.748 ;
      RECT 45.71 3.527 45.715 3.745 ;
      RECT 45.68 3.524 45.71 3.738 ;
      RECT 45.675 3.52 45.68 3.729 ;
      RECT 45.64 3.551 45.925 3.724 ;
      RECT 45.415 3.46 45.675 3.72 ;
      RECT 45.715 3.529 45.72 3.748 ;
      RECT 45.72 3.53 45.725 3.753 ;
      RECT 45.415 3.542 45.795 3.72 ;
      RECT 45.415 3.54 45.78 3.72 ;
      RECT 45.415 3.535 45.77 3.72 ;
      RECT 45.37 4.45 45.42 4.735 ;
      RECT 45.315 4.42 45.32 4.735 ;
      RECT 45.285 4.4 45.29 4.735 ;
      RECT 45.435 4.45 45.495 4.71 ;
      RECT 45.43 4.45 45.435 4.718 ;
      RECT 45.42 4.45 45.43 4.73 ;
      RECT 45.335 4.44 45.37 4.735 ;
      RECT 45.33 4.427 45.335 4.735 ;
      RECT 45.32 4.422 45.33 4.735 ;
      RECT 45.3 4.412 45.315 4.735 ;
      RECT 45.29 4.405 45.3 4.735 ;
      RECT 45.28 4.397 45.285 4.735 ;
      RECT 45.25 4.387 45.28 4.735 ;
      RECT 45.235 4.375 45.25 4.735 ;
      RECT 45.22 4.365 45.235 4.73 ;
      RECT 45.2 4.355 45.22 4.705 ;
      RECT 45.19 4.347 45.2 4.682 ;
      RECT 45.16 4.33 45.19 4.672 ;
      RECT 45.155 4.307 45.16 4.663 ;
      RECT 45.15 4.294 45.155 4.661 ;
      RECT 45.135 4.27 45.15 4.655 ;
      RECT 45.13 4.246 45.135 4.649 ;
      RECT 45.12 4.235 45.13 4.644 ;
      RECT 45.115 4.225 45.12 4.64 ;
      RECT 45.11 4.217 45.115 4.637 ;
      RECT 45.1 4.212 45.11 4.633 ;
      RECT 45.095 4.207 45.1 4.629 ;
      RECT 45.01 4.205 45.095 4.604 ;
      RECT 44.98 4.205 45.01 4.57 ;
      RECT 44.965 4.205 44.98 4.553 ;
      RECT 44.91 4.205 44.965 4.498 ;
      RECT 44.905 4.21 44.91 4.447 ;
      RECT 44.895 4.215 44.905 4.437 ;
      RECT 44.89 4.225 44.895 4.423 ;
      RECT 44.84 4.965 45.1 5.225 ;
      RECT 44.76 4.98 45.1 5.201 ;
      RECT 44.74 4.98 45.1 5.196 ;
      RECT 44.716 4.98 45.1 5.194 ;
      RECT 44.63 4.98 45.1 5.189 ;
      RECT 44.48 4.92 44.74 5.185 ;
      RECT 44.435 4.98 45.1 5.18 ;
      RECT 44.43 4.987 45.1 5.175 ;
      RECT 44.445 4.975 44.76 5.185 ;
      RECT 44.335 3.41 44.595 3.67 ;
      RECT 44.335 3.467 44.6 3.663 ;
      RECT 44.335 3.497 44.605 3.595 ;
      RECT 44.395 3.928 44.51 3.93 ;
      RECT 44.481 3.925 44.51 3.93 ;
      RECT 43.505 4.929 43.53 5.169 ;
      RECT 43.49 4.932 43.58 5.163 ;
      RECT 43.485 4.937 43.666 5.158 ;
      RECT 43.48 4.945 43.73 5.156 ;
      RECT 43.48 4.945 43.74 5.155 ;
      RECT 43.475 4.952 43.75 5.148 ;
      RECT 43.475 4.952 43.836 5.137 ;
      RECT 43.47 4.987 43.836 5.133 ;
      RECT 43.47 4.987 43.845 5.122 ;
      RECT 43.75 4.86 44.01 5.12 ;
      RECT 43.46 5.037 44.01 5.118 ;
      RECT 43.73 4.905 43.75 5.153 ;
      RECT 43.666 4.908 43.73 5.157 ;
      RECT 43.58 4.913 43.666 5.162 ;
      RECT 43.51 4.924 44.01 5.12 ;
      RECT 43.53 4.918 43.58 5.167 ;
      RECT 43.655 3.395 43.665 3.657 ;
      RECT 43.645 3.452 43.655 3.66 ;
      RECT 43.62 3.457 43.645 3.666 ;
      RECT 43.595 3.461 43.62 3.678 ;
      RECT 43.585 3.464 43.595 3.688 ;
      RECT 43.58 3.465 43.585 3.693 ;
      RECT 43.575 3.466 43.58 3.698 ;
      RECT 43.57 3.467 43.575 3.7 ;
      RECT 43.545 3.47 43.57 3.703 ;
      RECT 43.515 3.476 43.545 3.706 ;
      RECT 43.45 3.487 43.515 3.709 ;
      RECT 43.405 3.495 43.45 3.713 ;
      RECT 43.39 3.495 43.405 3.721 ;
      RECT 43.385 3.496 43.39 3.728 ;
      RECT 43.38 3.498 43.385 3.731 ;
      RECT 43.375 3.502 43.38 3.734 ;
      RECT 43.365 3.51 43.375 3.738 ;
      RECT 43.36 3.523 43.365 3.743 ;
      RECT 43.355 3.531 43.36 3.745 ;
      RECT 43.35 3.537 43.355 3.745 ;
      RECT 43.345 3.541 43.35 3.748 ;
      RECT 43.34 3.543 43.345 3.751 ;
      RECT 43.335 3.546 43.34 3.754 ;
      RECT 43.325 3.551 43.335 3.758 ;
      RECT 43.32 3.557 43.325 3.763 ;
      RECT 43.31 3.563 43.32 3.767 ;
      RECT 43.295 3.57 43.31 3.773 ;
      RECT 43.266 3.584 43.295 3.783 ;
      RECT 43.18 3.619 43.266 3.815 ;
      RECT 43.16 3.652 43.18 3.844 ;
      RECT 43.14 3.665 43.16 3.855 ;
      RECT 43.12 3.677 43.14 3.866 ;
      RECT 43.07 3.699 43.12 3.886 ;
      RECT 43.055 3.717 43.07 3.903 ;
      RECT 43.05 3.723 43.055 3.906 ;
      RECT 43.045 3.727 43.05 3.909 ;
      RECT 43.04 3.731 43.045 3.913 ;
      RECT 43.035 3.733 43.04 3.916 ;
      RECT 43.025 3.74 43.035 3.919 ;
      RECT 43.02 3.745 43.025 3.923 ;
      RECT 43.015 3.747 43.02 3.926 ;
      RECT 43.01 3.751 43.015 3.929 ;
      RECT 43.005 3.753 43.01 3.933 ;
      RECT 42.99 3.758 43.005 3.938 ;
      RECT 42.985 3.763 42.99 3.941 ;
      RECT 42.98 3.771 42.985 3.944 ;
      RECT 42.975 3.773 42.98 3.947 ;
      RECT 42.97 3.775 42.975 3.95 ;
      RECT 42.96 3.777 42.97 3.956 ;
      RECT 42.925 3.791 42.96 3.968 ;
      RECT 42.915 3.806 42.925 3.978 ;
      RECT 42.84 3.835 42.915 4.002 ;
      RECT 42.835 3.86 42.84 4.025 ;
      RECT 42.82 3.864 42.835 4.031 ;
      RECT 42.81 3.872 42.82 4.036 ;
      RECT 42.78 3.885 42.81 4.04 ;
      RECT 42.77 3.9 42.78 4.045 ;
      RECT 42.76 3.905 42.77 4.048 ;
      RECT 42.755 3.907 42.76 4.05 ;
      RECT 42.74 3.91 42.755 4.053 ;
      RECT 42.735 3.912 42.74 4.056 ;
      RECT 42.715 3.917 42.735 4.06 ;
      RECT 42.685 3.922 42.715 4.068 ;
      RECT 42.66 3.929 42.685 4.076 ;
      RECT 42.655 3.934 42.66 4.081 ;
      RECT 42.625 3.937 42.655 4.085 ;
      RECT 42.585 3.94 42.625 4.095 ;
      RECT 42.55 3.937 42.585 4.107 ;
      RECT 42.54 3.933 42.55 4.114 ;
      RECT 42.515 3.929 42.54 4.12 ;
      RECT 42.51 3.925 42.515 4.125 ;
      RECT 42.47 3.922 42.51 4.125 ;
      RECT 42.455 3.907 42.47 4.126 ;
      RECT 42.432 3.895 42.455 4.126 ;
      RECT 42.346 3.895 42.432 4.127 ;
      RECT 42.26 3.895 42.346 4.129 ;
      RECT 42.24 3.895 42.26 4.126 ;
      RECT 42.235 3.9 42.24 4.121 ;
      RECT 42.23 3.905 42.235 4.119 ;
      RECT 42.22 3.915 42.23 4.117 ;
      RECT 42.215 3.921 42.22 4.11 ;
      RECT 42.21 3.923 42.215 4.095 ;
      RECT 42.205 3.927 42.21 4.085 ;
      RECT 43.665 3.395 43.915 3.655 ;
      RECT 41.39 4.93 41.65 5.19 ;
      RECT 43.685 4.42 43.69 4.63 ;
      RECT 43.69 4.425 43.7 4.625 ;
      RECT 43.64 4.42 43.685 4.645 ;
      RECT 43.63 4.42 43.64 4.665 ;
      RECT 43.611 4.42 43.63 4.67 ;
      RECT 43.525 4.42 43.611 4.667 ;
      RECT 43.495 4.422 43.525 4.665 ;
      RECT 43.44 4.432 43.495 4.663 ;
      RECT 43.375 4.446 43.44 4.661 ;
      RECT 43.37 4.454 43.375 4.66 ;
      RECT 43.355 4.457 43.37 4.658 ;
      RECT 43.29 4.467 43.355 4.654 ;
      RECT 43.242 4.481 43.29 4.655 ;
      RECT 43.156 4.498 43.242 4.669 ;
      RECT 43.07 4.519 43.156 4.686 ;
      RECT 43.05 4.532 43.07 4.696 ;
      RECT 43.005 4.54 43.05 4.703 ;
      RECT 42.97 4.548 43.005 4.711 ;
      RECT 42.936 4.556 42.97 4.719 ;
      RECT 42.85 4.57 42.936 4.731 ;
      RECT 42.815 4.587 42.85 4.743 ;
      RECT 42.806 4.596 42.815 4.747 ;
      RECT 42.72 4.614 42.806 4.764 ;
      RECT 42.661 4.641 42.72 4.791 ;
      RECT 42.575 4.668 42.661 4.819 ;
      RECT 42.555 4.69 42.575 4.839 ;
      RECT 42.495 4.705 42.555 4.855 ;
      RECT 42.485 4.717 42.495 4.868 ;
      RECT 42.48 4.722 42.485 4.871 ;
      RECT 42.47 4.725 42.48 4.874 ;
      RECT 42.465 4.727 42.47 4.877 ;
      RECT 42.435 4.735 42.465 4.884 ;
      RECT 42.42 4.742 42.435 4.892 ;
      RECT 42.41 4.747 42.42 4.896 ;
      RECT 42.405 4.75 42.41 4.899 ;
      RECT 42.395 4.752 42.405 4.902 ;
      RECT 42.36 4.762 42.395 4.911 ;
      RECT 42.285 4.785 42.36 4.933 ;
      RECT 42.265 4.803 42.285 4.951 ;
      RECT 42.235 4.81 42.265 4.961 ;
      RECT 42.215 4.818 42.235 4.971 ;
      RECT 42.205 4.824 42.215 4.978 ;
      RECT 42.186 4.829 42.205 4.984 ;
      RECT 42.1 4.849 42.186 5.004 ;
      RECT 42.085 4.869 42.1 5.023 ;
      RECT 42.04 4.881 42.085 5.034 ;
      RECT 41.975 4.902 42.04 5.057 ;
      RECT 41.935 4.922 41.975 5.078 ;
      RECT 41.925 4.932 41.935 5.088 ;
      RECT 41.875 4.944 41.925 5.099 ;
      RECT 41.855 4.96 41.875 5.111 ;
      RECT 41.825 4.97 41.855 5.117 ;
      RECT 41.815 4.975 41.825 5.119 ;
      RECT 41.746 4.976 41.815 5.125 ;
      RECT 41.66 4.978 41.746 5.135 ;
      RECT 41.65 4.979 41.66 5.14 ;
      RECT 42.92 5.005 43.11 5.215 ;
      RECT 42.91 5.01 43.12 5.208 ;
      RECT 42.895 5.01 43.12 5.173 ;
      RECT 42.815 4.895 43.075 5.155 ;
      RECT 41.73 4.425 41.915 4.72 ;
      RECT 41.72 4.425 41.915 4.718 ;
      RECT 41.705 4.425 41.92 4.713 ;
      RECT 41.705 4.425 41.925 4.71 ;
      RECT 41.7 4.425 41.925 4.708 ;
      RECT 41.695 4.68 41.925 4.698 ;
      RECT 41.7 4.425 41.96 4.685 ;
      RECT 41.66 3.46 41.92 3.72 ;
      RECT 41.47 3.385 41.556 3.718 ;
      RECT 41.445 3.389 41.6 3.714 ;
      RECT 41.556 3.381 41.6 3.714 ;
      RECT 41.556 3.382 41.605 3.713 ;
      RECT 41.47 3.387 41.62 3.712 ;
      RECT 41.445 3.395 41.66 3.711 ;
      RECT 41.44 3.39 41.62 3.706 ;
      RECT 41.43 3.405 41.66 3.613 ;
      RECT 41.43 3.457 41.86 3.613 ;
      RECT 41.43 3.45 41.84 3.613 ;
      RECT 41.43 3.437 41.81 3.613 ;
      RECT 41.43 3.425 41.75 3.613 ;
      RECT 41.43 3.41 41.725 3.613 ;
      RECT 40.63 4.04 40.765 4.335 ;
      RECT 40.89 4.063 40.895 4.25 ;
      RECT 41.61 3.96 41.755 4.195 ;
      RECT 41.77 3.96 41.775 4.185 ;
      RECT 41.805 3.971 41.81 4.165 ;
      RECT 41.8 3.963 41.805 4.17 ;
      RECT 41.78 3.96 41.8 4.175 ;
      RECT 41.775 3.96 41.78 4.183 ;
      RECT 41.765 3.96 41.77 4.188 ;
      RECT 41.755 3.96 41.765 4.193 ;
      RECT 41.585 3.962 41.61 4.195 ;
      RECT 41.535 3.969 41.585 4.195 ;
      RECT 41.53 3.974 41.535 4.195 ;
      RECT 41.491 3.979 41.53 4.196 ;
      RECT 41.405 3.991 41.491 4.197 ;
      RECT 41.396 4.001 41.405 4.197 ;
      RECT 41.31 4.01 41.396 4.199 ;
      RECT 41.286 4.02 41.31 4.201 ;
      RECT 41.2 4.031 41.286 4.202 ;
      RECT 41.17 4.042 41.2 4.204 ;
      RECT 41.14 4.047 41.17 4.206 ;
      RECT 41.115 4.053 41.14 4.209 ;
      RECT 41.1 4.058 41.115 4.21 ;
      RECT 41.055 4.064 41.1 4.21 ;
      RECT 41.05 4.069 41.055 4.211 ;
      RECT 41.03 4.069 41.05 4.213 ;
      RECT 41.01 4.067 41.03 4.218 ;
      RECT 40.975 4.066 41.01 4.225 ;
      RECT 40.945 4.065 40.975 4.235 ;
      RECT 40.895 4.064 40.945 4.245 ;
      RECT 40.805 4.061 40.89 4.335 ;
      RECT 40.78 4.055 40.805 4.335 ;
      RECT 40.765 4.045 40.78 4.335 ;
      RECT 40.58 4.04 40.63 4.255 ;
      RECT 40.57 4.045 40.58 4.245 ;
      RECT 40.81 4.52 41.07 4.78 ;
      RECT 40.81 4.52 41.1 4.673 ;
      RECT 40.81 4.52 41.135 4.658 ;
      RECT 41.065 4.44 41.255 4.65 ;
      RECT 41.055 4.445 41.265 4.643 ;
      RECT 41.02 4.515 41.265 4.643 ;
      RECT 41.05 4.457 41.07 4.78 ;
      RECT 41.035 4.505 41.265 4.643 ;
      RECT 41.04 4.477 41.07 4.78 ;
      RECT 40.12 3.545 40.19 4.65 ;
      RECT 40.855 3.65 41.115 3.91 ;
      RECT 40.435 3.696 40.45 3.905 ;
      RECT 40.771 3.709 40.855 3.86 ;
      RECT 40.685 3.706 40.771 3.86 ;
      RECT 40.646 3.704 40.685 3.86 ;
      RECT 40.56 3.702 40.646 3.86 ;
      RECT 40.5 3.7 40.56 3.871 ;
      RECT 40.465 3.698 40.5 3.889 ;
      RECT 40.45 3.696 40.465 3.9 ;
      RECT 40.42 3.696 40.435 3.913 ;
      RECT 40.41 3.696 40.42 3.918 ;
      RECT 40.385 3.695 40.41 3.923 ;
      RECT 40.37 3.69 40.385 3.929 ;
      RECT 40.365 3.683 40.37 3.934 ;
      RECT 40.34 3.674 40.365 3.94 ;
      RECT 40.295 3.653 40.34 3.953 ;
      RECT 40.285 3.637 40.295 3.963 ;
      RECT 40.27 3.63 40.285 3.973 ;
      RECT 40.26 3.623 40.27 3.99 ;
      RECT 40.255 3.62 40.26 4.02 ;
      RECT 40.25 3.618 40.255 4.05 ;
      RECT 40.245 3.616 40.25 4.087 ;
      RECT 40.23 3.612 40.245 4.154 ;
      RECT 40.23 4.445 40.24 4.645 ;
      RECT 40.225 3.608 40.23 4.28 ;
      RECT 40.225 4.432 40.23 4.65 ;
      RECT 40.22 3.606 40.225 4.365 ;
      RECT 40.22 4.422 40.225 4.65 ;
      RECT 40.205 3.577 40.22 4.65 ;
      RECT 40.19 3.55 40.205 4.65 ;
      RECT 40.115 3.545 40.12 3.9 ;
      RECT 40.115 3.955 40.12 4.65 ;
      RECT 40.1 3.545 40.115 3.878 ;
      RECT 40.11 3.977 40.115 4.65 ;
      RECT 40.1 4.017 40.11 4.65 ;
      RECT 40.065 3.545 40.1 3.82 ;
      RECT 40.095 4.052 40.1 4.65 ;
      RECT 40.08 4.107 40.095 4.65 ;
      RECT 40.075 4.172 40.08 4.65 ;
      RECT 40.06 4.22 40.075 4.65 ;
      RECT 40.035 3.545 40.065 3.775 ;
      RECT 40.055 4.275 40.06 4.65 ;
      RECT 40.04 4.335 40.055 4.65 ;
      RECT 40.035 4.383 40.04 4.648 ;
      RECT 40.03 3.545 40.035 3.768 ;
      RECT 40.03 4.415 40.035 4.643 ;
      RECT 40.005 3.545 40.03 3.76 ;
      RECT 39.995 3.55 40.005 3.75 ;
      RECT 40.21 4.825 40.23 5.065 ;
      RECT 39.44 4.755 39.445 4.965 ;
      RECT 40.72 4.828 40.73 5.023 ;
      RECT 40.715 4.818 40.72 5.026 ;
      RECT 40.635 4.815 40.715 5.049 ;
      RECT 40.631 4.815 40.635 5.071 ;
      RECT 40.545 4.815 40.631 5.081 ;
      RECT 40.53 4.815 40.545 5.089 ;
      RECT 40.501 4.816 40.53 5.087 ;
      RECT 40.415 4.821 40.501 5.083 ;
      RECT 40.402 4.825 40.415 5.079 ;
      RECT 40.316 4.825 40.402 5.075 ;
      RECT 40.23 4.825 40.316 5.069 ;
      RECT 40.146 4.825 40.21 5.063 ;
      RECT 40.06 4.825 40.146 5.058 ;
      RECT 40.04 4.825 40.06 5.054 ;
      RECT 39.98 4.82 40.04 5.051 ;
      RECT 39.952 4.814 39.98 5.048 ;
      RECT 39.866 4.809 39.952 5.044 ;
      RECT 39.78 4.803 39.866 5.038 ;
      RECT 39.705 4.785 39.78 5.033 ;
      RECT 39.67 4.762 39.705 5.029 ;
      RECT 39.66 4.752 39.67 5.028 ;
      RECT 39.605 4.75 39.66 5.027 ;
      RECT 39.53 4.75 39.605 5.023 ;
      RECT 39.52 4.75 39.53 5.018 ;
      RECT 39.505 4.75 39.52 5.01 ;
      RECT 39.455 4.752 39.505 4.988 ;
      RECT 39.445 4.755 39.455 4.968 ;
      RECT 39.435 4.76 39.44 4.963 ;
      RECT 39.43 4.765 39.435 4.958 ;
      RECT 37.54 3.41 37.8 3.67 ;
      RECT 37.53 3.44 37.8 3.65 ;
      RECT 39.45 3.355 39.71 3.615 ;
      RECT 39.445 3.43 39.45 3.616 ;
      RECT 39.42 3.435 39.445 3.618 ;
      RECT 39.405 3.442 39.42 3.621 ;
      RECT 39.345 3.46 39.405 3.626 ;
      RECT 39.315 3.48 39.345 3.633 ;
      RECT 39.29 3.488 39.315 3.638 ;
      RECT 39.265 3.496 39.29 3.64 ;
      RECT 39.247 3.5 39.265 3.639 ;
      RECT 39.161 3.498 39.247 3.639 ;
      RECT 39.075 3.496 39.161 3.639 ;
      RECT 38.989 3.494 39.075 3.638 ;
      RECT 38.903 3.492 38.989 3.638 ;
      RECT 38.817 3.49 38.903 3.638 ;
      RECT 38.731 3.488 38.817 3.638 ;
      RECT 38.645 3.486 38.731 3.637 ;
      RECT 38.627 3.485 38.645 3.637 ;
      RECT 38.541 3.484 38.627 3.637 ;
      RECT 38.455 3.482 38.541 3.637 ;
      RECT 38.369 3.481 38.455 3.636 ;
      RECT 38.283 3.48 38.369 3.636 ;
      RECT 38.197 3.478 38.283 3.636 ;
      RECT 38.111 3.477 38.197 3.636 ;
      RECT 38.025 3.475 38.111 3.635 ;
      RECT 38.001 3.473 38.025 3.635 ;
      RECT 37.915 3.466 38.001 3.635 ;
      RECT 37.886 3.458 37.915 3.635 ;
      RECT 37.8 3.45 37.886 3.635 ;
      RECT 37.52 3.447 37.53 3.645 ;
      RECT 39.025 4.41 39.03 4.76 ;
      RECT 38.795 4.5 38.935 4.76 ;
      RECT 39.27 4.185 39.315 4.395 ;
      RECT 39.325 4.196 39.335 4.39 ;
      RECT 39.315 4.188 39.325 4.395 ;
      RECT 39.25 4.185 39.27 4.4 ;
      RECT 39.22 4.185 39.25 4.423 ;
      RECT 39.21 4.185 39.22 4.448 ;
      RECT 39.205 4.185 39.21 4.458 ;
      RECT 39.15 4.185 39.205 4.498 ;
      RECT 39.145 4.185 39.15 4.538 ;
      RECT 39.14 4.187 39.145 4.543 ;
      RECT 39.125 4.197 39.14 4.554 ;
      RECT 39.08 4.255 39.125 4.59 ;
      RECT 39.07 4.31 39.08 4.624 ;
      RECT 39.055 4.337 39.07 4.64 ;
      RECT 39.045 4.364 39.055 4.76 ;
      RECT 39.03 4.387 39.045 4.76 ;
      RECT 39.02 4.427 39.025 4.76 ;
      RECT 39.015 4.437 39.02 4.76 ;
      RECT 39.01 4.452 39.015 4.76 ;
      RECT 39 4.457 39.01 4.76 ;
      RECT 38.935 4.48 39 4.76 ;
      RECT 38.405 3.875 38.635 4.185 ;
      RECT 38.305 3.875 38.635 4.165 ;
      RECT 37.01 3.9 37.27 4.16 ;
      RECT 38.135 3.875 38.635 4.155 ;
      RECT 37.95 3.875 38.635 4.145 ;
      RECT 37.765 3.925 38.635 4.135 ;
      RECT 37.645 3.925 38.635 4.125 ;
      RECT 37.315 3.925 38.635 4.115 ;
      RECT 37.31 3.925 38.635 4.101 ;
      RECT 37.01 3.915 37.595 4.098 ;
      RECT 37.88 3.875 38.695 4.015 ;
      RECT 37.315 3.91 37.585 4.115 ;
      RECT 37.315 3.895 37.575 4.115 ;
      RECT 37.525 4.415 37.785 4.675 ;
      RECT 37.525 4.455 37.89 4.665 ;
      RECT 37.525 4.457 37.895 4.664 ;
      RECT 37.525 4.465 37.9 4.661 ;
      RECT 36.45 3.54 36.55 5.065 ;
      RECT 36.64 4.68 36.69 4.94 ;
      RECT 36.635 3.553 36.64 3.74 ;
      RECT 36.63 4.661 36.64 4.94 ;
      RECT 36.63 3.55 36.635 3.748 ;
      RECT 36.615 3.544 36.63 3.755 ;
      RECT 36.625 4.649 36.63 5.023 ;
      RECT 36.615 4.637 36.625 5.06 ;
      RECT 36.605 3.54 36.615 3.762 ;
      RECT 36.605 4.622 36.615 5.065 ;
      RECT 36.6 3.54 36.605 3.77 ;
      RECT 36.58 4.592 36.605 5.065 ;
      RECT 36.56 3.54 36.6 3.818 ;
      RECT 36.57 4.552 36.58 5.065 ;
      RECT 36.56 4.507 36.57 5.065 ;
      RECT 36.555 3.54 36.56 3.888 ;
      RECT 36.555 4.465 36.56 5.065 ;
      RECT 36.55 3.54 36.555 4.365 ;
      RECT 36.55 4.447 36.555 5.065 ;
      RECT 36.44 3.543 36.45 5.065 ;
      RECT 36.425 3.55 36.44 5.061 ;
      RECT 36.42 3.56 36.425 5.056 ;
      RECT 36.415 3.76 36.42 4.948 ;
      RECT 36.41 3.845 36.415 4.5 ;
      RECT 35.275 10.205 35.57 10.435 ;
      RECT 35.335 8.725 35.505 10.435 ;
      RECT 35.33 9.095 35.68 9.445 ;
      RECT 35.275 8.725 35.565 8.955 ;
      RECT 34.285 10.205 34.58 10.435 ;
      RECT 34.345 8.725 34.515 10.435 ;
      RECT 34.285 8.725 34.575 8.955 ;
      RECT 34.285 8.76 35.135 8.92 ;
      RECT 34.97 8.355 35.135 8.92 ;
      RECT 34.285 8.755 34.68 8.92 ;
      RECT 34.905 8.355 35.195 8.585 ;
      RECT 34.905 8.385 35.365 8.555 ;
      RECT 34.87 4.025 35.195 4.26 ;
      RECT 34.87 4.055 35.36 4.225 ;
      RECT 34.87 3.69 35.06 4.26 ;
      RECT 34.285 3.655 34.575 3.885 ;
      RECT 34.285 3.69 35.06 3.86 ;
      RECT 34.345 2.175 34.515 3.885 ;
      RECT 34.285 2.175 34.58 2.405 ;
      RECT 33.915 4.025 34.205 4.255 ;
      RECT 33.915 4.055 34.375 4.225 ;
      RECT 33.98 2.95 34.145 4.255 ;
      RECT 32.495 2.915 32.785 3.145 ;
      RECT 32.495 2.95 34.145 3.12 ;
      RECT 32.555 2.175 32.725 3.145 ;
      RECT 32.495 2.175 32.785 2.405 ;
      RECT 32.495 10.205 32.785 10.435 ;
      RECT 32.555 9.465 32.725 10.435 ;
      RECT 32.555 9.555 34.145 9.725 ;
      RECT 33.975 8.355 34.145 9.725 ;
      RECT 32.495 9.465 32.785 9.695 ;
      RECT 33.915 8.355 34.205 8.585 ;
      RECT 33.915 8.385 34.375 8.555 ;
      RECT 30.53 4.725 30.88 5.075 ;
      RECT 30.62 3.32 30.79 5.075 ;
      RECT 32.925 3.26 33.275 3.61 ;
      RECT 30.62 3.32 32.24 3.495 ;
      RECT 30.62 3.32 32.895 3.49 ;
      RECT 32.755 3.315 33.275 3.485 ;
      RECT 32.95 9.09 33.275 9.415 ;
      RECT 28.345 9.04 28.695 9.39 ;
      RECT 32.925 9.095 33.275 9.325 ;
      RECT 28.165 9.095 28.695 9.325 ;
      RECT 32.755 9.12 33.275 9.295 ;
      RECT 27.995 9.125 28.695 9.295 ;
      RECT 28.165 9.12 33.275 9.29 ;
      RECT 32.15 3.66 32.47 3.98 ;
      RECT 32.125 3.655 32.415 3.885 ;
      RECT 32.08 3.685 32.47 3.86 ;
      RECT 31.95 3.685 32.47 3.855 ;
      RECT 32.15 8.66 32.47 8.98 ;
      RECT 32.125 8.725 32.47 8.955 ;
      RECT 31.95 8.755 32.47 8.925 ;
      RECT 27.94 4.96 27.98 5.22 ;
      RECT 27.98 4.94 27.985 4.95 ;
      RECT 29.31 4.185 29.32 4.406 ;
      RECT 29.24 4.18 29.31 4.531 ;
      RECT 29.23 4.18 29.24 4.658 ;
      RECT 29.205 4.18 29.23 4.705 ;
      RECT 29.18 4.18 29.205 4.783 ;
      RECT 29.16 4.18 29.18 4.853 ;
      RECT 29.135 4.18 29.16 4.893 ;
      RECT 29.125 4.18 29.135 4.913 ;
      RECT 29.115 4.182 29.125 4.921 ;
      RECT 29.11 4.187 29.115 4.378 ;
      RECT 29.11 4.387 29.115 4.922 ;
      RECT 29.105 4.432 29.11 4.923 ;
      RECT 29.095 4.497 29.105 4.924 ;
      RECT 29.085 4.592 29.095 4.926 ;
      RECT 29.08 4.645 29.085 4.928 ;
      RECT 29.075 4.665 29.08 4.929 ;
      RECT 29.02 4.69 29.075 4.935 ;
      RECT 28.98 4.725 29.02 4.944 ;
      RECT 28.97 4.742 28.98 4.949 ;
      RECT 28.961 4.748 28.97 4.951 ;
      RECT 28.875 4.786 28.961 4.962 ;
      RECT 28.87 4.825 28.875 4.972 ;
      RECT 28.795 4.832 28.87 4.982 ;
      RECT 28.775 4.842 28.795 4.993 ;
      RECT 28.745 4.849 28.775 5.001 ;
      RECT 28.72 4.856 28.745 5.008 ;
      RECT 28.696 4.862 28.72 5.013 ;
      RECT 28.61 4.875 28.696 5.025 ;
      RECT 28.532 4.882 28.61 5.043 ;
      RECT 28.446 4.877 28.532 5.061 ;
      RECT 28.36 4.872 28.446 5.081 ;
      RECT 28.28 4.866 28.36 5.098 ;
      RECT 28.215 4.862 28.28 5.127 ;
      RECT 28.21 4.576 28.215 4.6 ;
      RECT 28.2 4.852 28.215 5.155 ;
      RECT 28.205 4.57 28.21 4.64 ;
      RECT 28.2 4.564 28.205 4.71 ;
      RECT 28.195 4.558 28.2 4.788 ;
      RECT 28.195 4.835 28.2 5.22 ;
      RECT 28.187 4.555 28.195 5.22 ;
      RECT 28.101 4.553 28.187 5.22 ;
      RECT 28.015 4.551 28.101 5.22 ;
      RECT 28.005 4.552 28.015 5.22 ;
      RECT 28 4.557 28.005 5.22 ;
      RECT 27.99 4.57 28 5.22 ;
      RECT 27.985 4.592 27.99 5.22 ;
      RECT 27.98 4.952 27.985 5.22 ;
      RECT 28.61 4.42 28.615 4.64 ;
      RECT 29.115 3.455 29.15 3.715 ;
      RECT 29.1 3.455 29.115 3.723 ;
      RECT 29.071 3.455 29.1 3.745 ;
      RECT 28.985 3.455 29.071 3.805 ;
      RECT 28.965 3.455 28.985 3.87 ;
      RECT 28.905 3.455 28.965 4.035 ;
      RECT 28.9 3.455 28.905 4.183 ;
      RECT 28.895 3.455 28.9 4.195 ;
      RECT 28.89 3.455 28.895 4.221 ;
      RECT 28.86 3.641 28.89 4.301 ;
      RECT 28.855 3.689 28.86 4.39 ;
      RECT 28.85 3.703 28.855 4.405 ;
      RECT 28.845 3.722 28.85 4.435 ;
      RECT 28.84 3.737 28.845 4.451 ;
      RECT 28.835 3.752 28.84 4.473 ;
      RECT 28.83 3.772 28.835 4.495 ;
      RECT 28.82 3.792 28.83 4.528 ;
      RECT 28.805 3.834 28.82 4.59 ;
      RECT 28.8 3.865 28.805 4.63 ;
      RECT 28.795 3.877 28.8 4.635 ;
      RECT 28.79 3.889 28.795 4.64 ;
      RECT 28.785 3.902 28.79 4.64 ;
      RECT 28.78 3.92 28.785 4.64 ;
      RECT 28.775 3.94 28.78 4.64 ;
      RECT 28.77 3.952 28.775 4.64 ;
      RECT 28.765 3.965 28.77 4.64 ;
      RECT 28.745 4 28.765 4.64 ;
      RECT 28.695 4.102 28.745 4.64 ;
      RECT 28.69 4.187 28.695 4.64 ;
      RECT 28.685 4.195 28.69 4.64 ;
      RECT 28.68 4.212 28.685 4.64 ;
      RECT 28.675 4.227 28.68 4.64 ;
      RECT 28.64 4.292 28.675 4.64 ;
      RECT 28.625 4.357 28.64 4.64 ;
      RECT 28.62 4.387 28.625 4.64 ;
      RECT 28.615 4.412 28.62 4.64 ;
      RECT 28.6 4.422 28.61 4.64 ;
      RECT 28.585 4.435 28.6 4.633 ;
      RECT 28.33 4.025 28.4 4.235 ;
      RECT 28.12 4.002 28.125 4.195 ;
      RECT 25.575 3.93 25.835 4.19 ;
      RECT 28.41 4.212 28.415 4.215 ;
      RECT 28.4 4.03 28.41 4.23 ;
      RECT 28.301 4.023 28.33 4.235 ;
      RECT 28.215 4.015 28.301 4.235 ;
      RECT 28.2 4.009 28.215 4.233 ;
      RECT 28.18 4.008 28.2 4.22 ;
      RECT 28.175 4.007 28.18 4.203 ;
      RECT 28.125 4.004 28.175 4.198 ;
      RECT 28.095 4.001 28.12 4.193 ;
      RECT 28.075 3.999 28.095 4.188 ;
      RECT 28.06 3.997 28.075 4.185 ;
      RECT 28.03 3.995 28.06 4.183 ;
      RECT 27.965 3.991 28.03 4.175 ;
      RECT 27.935 3.986 27.965 4.17 ;
      RECT 27.915 3.984 27.935 4.168 ;
      RECT 27.885 3.981 27.915 4.163 ;
      RECT 27.825 3.977 27.885 4.155 ;
      RECT 27.82 3.974 27.825 4.15 ;
      RECT 27.75 3.972 27.82 4.145 ;
      RECT 27.721 3.968 27.75 4.138 ;
      RECT 27.635 3.963 27.721 4.13 ;
      RECT 27.601 3.958 27.635 4.122 ;
      RECT 27.515 3.95 27.601 4.114 ;
      RECT 27.476 3.943 27.515 4.106 ;
      RECT 27.39 3.938 27.476 4.098 ;
      RECT 27.325 3.932 27.39 4.088 ;
      RECT 27.305 3.927 27.325 4.083 ;
      RECT 27.296 3.924 27.305 4.082 ;
      RECT 27.21 3.92 27.296 4.076 ;
      RECT 27.17 3.916 27.21 4.068 ;
      RECT 27.15 3.912 27.17 4.066 ;
      RECT 27.09 3.912 27.15 4.063 ;
      RECT 27.07 3.915 27.09 4.061 ;
      RECT 27.049 3.915 27.07 4.061 ;
      RECT 26.963 3.917 27.049 4.065 ;
      RECT 26.877 3.919 26.963 4.071 ;
      RECT 26.791 3.921 26.877 4.078 ;
      RECT 26.705 3.924 26.791 4.084 ;
      RECT 26.671 3.925 26.705 4.089 ;
      RECT 26.585 3.928 26.671 4.094 ;
      RECT 26.556 3.935 26.585 4.099 ;
      RECT 26.47 3.935 26.556 4.104 ;
      RECT 26.437 3.935 26.47 4.109 ;
      RECT 26.351 3.937 26.437 4.114 ;
      RECT 26.265 3.939 26.351 4.121 ;
      RECT 26.201 3.941 26.265 4.127 ;
      RECT 26.115 3.943 26.201 4.133 ;
      RECT 26.112 3.945 26.115 4.136 ;
      RECT 26.026 3.946 26.112 4.14 ;
      RECT 25.94 3.949 26.026 4.147 ;
      RECT 25.921 3.951 25.94 4.151 ;
      RECT 25.835 3.953 25.921 4.156 ;
      RECT 25.565 3.965 25.575 4.16 ;
      RECT 27.735 10.205 28.025 10.435 ;
      RECT 27.795 9.465 27.965 10.435 ;
      RECT 27.685 9.49 28.06 9.86 ;
      RECT 27.735 9.465 28.025 9.86 ;
      RECT 27.8 3.545 27.985 3.755 ;
      RECT 27.795 3.546 27.99 3.753 ;
      RECT 27.79 3.551 28 3.748 ;
      RECT 27.785 3.527 27.79 3.745 ;
      RECT 27.755 3.524 27.785 3.738 ;
      RECT 27.75 3.52 27.755 3.729 ;
      RECT 27.715 3.551 28 3.724 ;
      RECT 27.49 3.46 27.75 3.72 ;
      RECT 27.79 3.529 27.795 3.748 ;
      RECT 27.795 3.53 27.8 3.753 ;
      RECT 27.49 3.542 27.87 3.72 ;
      RECT 27.49 3.54 27.855 3.72 ;
      RECT 27.49 3.535 27.845 3.72 ;
      RECT 27.445 4.45 27.495 4.735 ;
      RECT 27.39 4.42 27.395 4.735 ;
      RECT 27.36 4.4 27.365 4.735 ;
      RECT 27.51 4.45 27.57 4.71 ;
      RECT 27.505 4.45 27.51 4.718 ;
      RECT 27.495 4.45 27.505 4.73 ;
      RECT 27.41 4.44 27.445 4.735 ;
      RECT 27.405 4.427 27.41 4.735 ;
      RECT 27.395 4.422 27.405 4.735 ;
      RECT 27.375 4.412 27.39 4.735 ;
      RECT 27.365 4.405 27.375 4.735 ;
      RECT 27.355 4.397 27.36 4.735 ;
      RECT 27.325 4.387 27.355 4.735 ;
      RECT 27.31 4.375 27.325 4.735 ;
      RECT 27.295 4.365 27.31 4.73 ;
      RECT 27.275 4.355 27.295 4.705 ;
      RECT 27.265 4.347 27.275 4.682 ;
      RECT 27.235 4.33 27.265 4.672 ;
      RECT 27.23 4.307 27.235 4.663 ;
      RECT 27.225 4.294 27.23 4.661 ;
      RECT 27.21 4.27 27.225 4.655 ;
      RECT 27.205 4.246 27.21 4.649 ;
      RECT 27.195 4.235 27.205 4.644 ;
      RECT 27.19 4.225 27.195 4.64 ;
      RECT 27.185 4.217 27.19 4.637 ;
      RECT 27.175 4.212 27.185 4.633 ;
      RECT 27.17 4.207 27.175 4.629 ;
      RECT 27.085 4.205 27.17 4.604 ;
      RECT 27.055 4.205 27.085 4.57 ;
      RECT 27.04 4.205 27.055 4.553 ;
      RECT 26.985 4.205 27.04 4.498 ;
      RECT 26.98 4.21 26.985 4.447 ;
      RECT 26.97 4.215 26.98 4.437 ;
      RECT 26.965 4.225 26.97 4.423 ;
      RECT 26.915 4.965 27.175 5.225 ;
      RECT 26.835 4.98 27.175 5.201 ;
      RECT 26.815 4.98 27.175 5.196 ;
      RECT 26.791 4.98 27.175 5.194 ;
      RECT 26.705 4.98 27.175 5.189 ;
      RECT 26.555 4.92 26.815 5.185 ;
      RECT 26.51 4.98 27.175 5.18 ;
      RECT 26.505 4.987 27.175 5.175 ;
      RECT 26.52 4.975 26.835 5.185 ;
      RECT 26.41 3.41 26.67 3.67 ;
      RECT 26.41 3.467 26.675 3.663 ;
      RECT 26.41 3.497 26.68 3.595 ;
      RECT 26.47 3.928 26.585 3.93 ;
      RECT 26.556 3.925 26.585 3.93 ;
      RECT 25.58 4.929 25.605 5.169 ;
      RECT 25.565 4.932 25.655 5.163 ;
      RECT 25.56 4.937 25.741 5.158 ;
      RECT 25.555 4.945 25.805 5.156 ;
      RECT 25.555 4.945 25.815 5.155 ;
      RECT 25.55 4.952 25.825 5.148 ;
      RECT 25.55 4.952 25.911 5.137 ;
      RECT 25.545 4.987 25.911 5.133 ;
      RECT 25.545 4.987 25.92 5.122 ;
      RECT 25.825 4.86 26.085 5.12 ;
      RECT 25.535 5.037 26.085 5.118 ;
      RECT 25.805 4.905 25.825 5.153 ;
      RECT 25.741 4.908 25.805 5.157 ;
      RECT 25.655 4.913 25.741 5.162 ;
      RECT 25.585 4.924 26.085 5.12 ;
      RECT 25.605 4.918 25.655 5.167 ;
      RECT 25.73 3.395 25.74 3.657 ;
      RECT 25.72 3.452 25.73 3.66 ;
      RECT 25.695 3.457 25.72 3.666 ;
      RECT 25.67 3.461 25.695 3.678 ;
      RECT 25.66 3.464 25.67 3.688 ;
      RECT 25.655 3.465 25.66 3.693 ;
      RECT 25.65 3.466 25.655 3.698 ;
      RECT 25.645 3.467 25.65 3.7 ;
      RECT 25.62 3.47 25.645 3.703 ;
      RECT 25.59 3.476 25.62 3.706 ;
      RECT 25.525 3.487 25.59 3.709 ;
      RECT 25.48 3.495 25.525 3.713 ;
      RECT 25.465 3.495 25.48 3.721 ;
      RECT 25.46 3.496 25.465 3.728 ;
      RECT 25.455 3.498 25.46 3.731 ;
      RECT 25.45 3.502 25.455 3.734 ;
      RECT 25.44 3.51 25.45 3.738 ;
      RECT 25.435 3.523 25.44 3.743 ;
      RECT 25.43 3.531 25.435 3.745 ;
      RECT 25.425 3.537 25.43 3.745 ;
      RECT 25.42 3.541 25.425 3.748 ;
      RECT 25.415 3.543 25.42 3.751 ;
      RECT 25.41 3.546 25.415 3.754 ;
      RECT 25.4 3.551 25.41 3.758 ;
      RECT 25.395 3.557 25.4 3.763 ;
      RECT 25.385 3.563 25.395 3.767 ;
      RECT 25.37 3.57 25.385 3.773 ;
      RECT 25.341 3.584 25.37 3.783 ;
      RECT 25.255 3.619 25.341 3.815 ;
      RECT 25.235 3.652 25.255 3.844 ;
      RECT 25.215 3.665 25.235 3.855 ;
      RECT 25.195 3.677 25.215 3.866 ;
      RECT 25.145 3.699 25.195 3.886 ;
      RECT 25.13 3.717 25.145 3.903 ;
      RECT 25.125 3.723 25.13 3.906 ;
      RECT 25.12 3.727 25.125 3.909 ;
      RECT 25.115 3.731 25.12 3.913 ;
      RECT 25.11 3.733 25.115 3.916 ;
      RECT 25.1 3.74 25.11 3.919 ;
      RECT 25.095 3.745 25.1 3.923 ;
      RECT 25.09 3.747 25.095 3.926 ;
      RECT 25.085 3.751 25.09 3.929 ;
      RECT 25.08 3.753 25.085 3.933 ;
      RECT 25.065 3.758 25.08 3.938 ;
      RECT 25.06 3.763 25.065 3.941 ;
      RECT 25.055 3.771 25.06 3.944 ;
      RECT 25.05 3.773 25.055 3.947 ;
      RECT 25.045 3.775 25.05 3.95 ;
      RECT 25.035 3.777 25.045 3.956 ;
      RECT 25 3.791 25.035 3.968 ;
      RECT 24.99 3.806 25 3.978 ;
      RECT 24.915 3.835 24.99 4.002 ;
      RECT 24.91 3.86 24.915 4.025 ;
      RECT 24.895 3.864 24.91 4.031 ;
      RECT 24.885 3.872 24.895 4.036 ;
      RECT 24.855 3.885 24.885 4.04 ;
      RECT 24.845 3.9 24.855 4.045 ;
      RECT 24.835 3.905 24.845 4.048 ;
      RECT 24.83 3.907 24.835 4.05 ;
      RECT 24.815 3.91 24.83 4.053 ;
      RECT 24.81 3.912 24.815 4.056 ;
      RECT 24.79 3.917 24.81 4.06 ;
      RECT 24.76 3.922 24.79 4.068 ;
      RECT 24.735 3.929 24.76 4.076 ;
      RECT 24.73 3.934 24.735 4.081 ;
      RECT 24.7 3.937 24.73 4.085 ;
      RECT 24.66 3.94 24.7 4.095 ;
      RECT 24.625 3.937 24.66 4.107 ;
      RECT 24.615 3.933 24.625 4.114 ;
      RECT 24.59 3.929 24.615 4.12 ;
      RECT 24.585 3.925 24.59 4.125 ;
      RECT 24.545 3.922 24.585 4.125 ;
      RECT 24.53 3.907 24.545 4.126 ;
      RECT 24.507 3.895 24.53 4.126 ;
      RECT 24.421 3.895 24.507 4.127 ;
      RECT 24.335 3.895 24.421 4.129 ;
      RECT 24.315 3.895 24.335 4.126 ;
      RECT 24.31 3.9 24.315 4.121 ;
      RECT 24.305 3.905 24.31 4.119 ;
      RECT 24.295 3.915 24.305 4.117 ;
      RECT 24.29 3.921 24.295 4.11 ;
      RECT 24.285 3.923 24.29 4.095 ;
      RECT 24.28 3.927 24.285 4.085 ;
      RECT 25.74 3.395 25.99 3.655 ;
      RECT 23.465 4.93 23.725 5.19 ;
      RECT 25.76 4.42 25.765 4.63 ;
      RECT 25.765 4.425 25.775 4.625 ;
      RECT 25.715 4.42 25.76 4.645 ;
      RECT 25.705 4.42 25.715 4.665 ;
      RECT 25.686 4.42 25.705 4.67 ;
      RECT 25.6 4.42 25.686 4.667 ;
      RECT 25.57 4.422 25.6 4.665 ;
      RECT 25.515 4.432 25.57 4.663 ;
      RECT 25.45 4.446 25.515 4.661 ;
      RECT 25.445 4.454 25.45 4.66 ;
      RECT 25.43 4.457 25.445 4.658 ;
      RECT 25.365 4.467 25.43 4.654 ;
      RECT 25.317 4.481 25.365 4.655 ;
      RECT 25.231 4.498 25.317 4.669 ;
      RECT 25.145 4.519 25.231 4.686 ;
      RECT 25.125 4.532 25.145 4.696 ;
      RECT 25.08 4.54 25.125 4.703 ;
      RECT 25.045 4.548 25.08 4.711 ;
      RECT 25.011 4.556 25.045 4.719 ;
      RECT 24.925 4.57 25.011 4.731 ;
      RECT 24.89 4.587 24.925 4.743 ;
      RECT 24.881 4.596 24.89 4.747 ;
      RECT 24.795 4.614 24.881 4.764 ;
      RECT 24.736 4.641 24.795 4.791 ;
      RECT 24.65 4.668 24.736 4.819 ;
      RECT 24.63 4.69 24.65 4.839 ;
      RECT 24.57 4.705 24.63 4.855 ;
      RECT 24.56 4.717 24.57 4.868 ;
      RECT 24.555 4.722 24.56 4.871 ;
      RECT 24.545 4.725 24.555 4.874 ;
      RECT 24.54 4.727 24.545 4.877 ;
      RECT 24.51 4.735 24.54 4.884 ;
      RECT 24.495 4.742 24.51 4.892 ;
      RECT 24.485 4.747 24.495 4.896 ;
      RECT 24.48 4.75 24.485 4.899 ;
      RECT 24.47 4.752 24.48 4.902 ;
      RECT 24.435 4.762 24.47 4.911 ;
      RECT 24.36 4.785 24.435 4.933 ;
      RECT 24.34 4.803 24.36 4.951 ;
      RECT 24.31 4.81 24.34 4.961 ;
      RECT 24.29 4.818 24.31 4.971 ;
      RECT 24.28 4.824 24.29 4.978 ;
      RECT 24.261 4.829 24.28 4.984 ;
      RECT 24.175 4.849 24.261 5.004 ;
      RECT 24.16 4.869 24.175 5.023 ;
      RECT 24.115 4.881 24.16 5.034 ;
      RECT 24.05 4.902 24.115 5.057 ;
      RECT 24.01 4.922 24.05 5.078 ;
      RECT 24 4.932 24.01 5.088 ;
      RECT 23.95 4.944 24 5.099 ;
      RECT 23.93 4.96 23.95 5.111 ;
      RECT 23.9 4.97 23.93 5.117 ;
      RECT 23.89 4.975 23.9 5.119 ;
      RECT 23.821 4.976 23.89 5.125 ;
      RECT 23.735 4.978 23.821 5.135 ;
      RECT 23.725 4.979 23.735 5.14 ;
      RECT 24.995 5.005 25.185 5.215 ;
      RECT 24.985 5.01 25.195 5.208 ;
      RECT 24.97 5.01 25.195 5.173 ;
      RECT 24.89 4.895 25.15 5.155 ;
      RECT 23.805 4.425 23.99 4.72 ;
      RECT 23.795 4.425 23.99 4.718 ;
      RECT 23.78 4.425 23.995 4.713 ;
      RECT 23.78 4.425 24 4.71 ;
      RECT 23.775 4.425 24 4.708 ;
      RECT 23.77 4.68 24 4.698 ;
      RECT 23.775 4.425 24.035 4.685 ;
      RECT 23.735 3.46 23.995 3.72 ;
      RECT 23.545 3.385 23.631 3.718 ;
      RECT 23.52 3.389 23.675 3.714 ;
      RECT 23.631 3.381 23.675 3.714 ;
      RECT 23.631 3.382 23.68 3.713 ;
      RECT 23.545 3.387 23.695 3.712 ;
      RECT 23.52 3.395 23.735 3.711 ;
      RECT 23.515 3.39 23.695 3.706 ;
      RECT 23.505 3.405 23.735 3.613 ;
      RECT 23.505 3.457 23.935 3.613 ;
      RECT 23.505 3.45 23.915 3.613 ;
      RECT 23.505 3.437 23.885 3.613 ;
      RECT 23.505 3.425 23.825 3.613 ;
      RECT 23.505 3.41 23.8 3.613 ;
      RECT 22.705 4.04 22.84 4.335 ;
      RECT 22.965 4.063 22.97 4.25 ;
      RECT 23.685 3.96 23.83 4.195 ;
      RECT 23.845 3.96 23.85 4.185 ;
      RECT 23.88 3.971 23.885 4.165 ;
      RECT 23.875 3.963 23.88 4.17 ;
      RECT 23.855 3.96 23.875 4.175 ;
      RECT 23.85 3.96 23.855 4.183 ;
      RECT 23.84 3.96 23.845 4.188 ;
      RECT 23.83 3.96 23.84 4.193 ;
      RECT 23.66 3.962 23.685 4.195 ;
      RECT 23.61 3.969 23.66 4.195 ;
      RECT 23.605 3.974 23.61 4.195 ;
      RECT 23.566 3.979 23.605 4.196 ;
      RECT 23.48 3.991 23.566 4.197 ;
      RECT 23.471 4.001 23.48 4.197 ;
      RECT 23.385 4.01 23.471 4.199 ;
      RECT 23.361 4.02 23.385 4.201 ;
      RECT 23.275 4.031 23.361 4.202 ;
      RECT 23.245 4.042 23.275 4.204 ;
      RECT 23.215 4.047 23.245 4.206 ;
      RECT 23.19 4.053 23.215 4.209 ;
      RECT 23.175 4.058 23.19 4.21 ;
      RECT 23.13 4.064 23.175 4.21 ;
      RECT 23.125 4.069 23.13 4.211 ;
      RECT 23.105 4.069 23.125 4.213 ;
      RECT 23.085 4.067 23.105 4.218 ;
      RECT 23.05 4.066 23.085 4.225 ;
      RECT 23.02 4.065 23.05 4.235 ;
      RECT 22.97 4.064 23.02 4.245 ;
      RECT 22.88 4.061 22.965 4.335 ;
      RECT 22.855 4.055 22.88 4.335 ;
      RECT 22.84 4.045 22.855 4.335 ;
      RECT 22.655 4.04 22.705 4.255 ;
      RECT 22.645 4.045 22.655 4.245 ;
      RECT 22.885 4.52 23.145 4.78 ;
      RECT 22.885 4.52 23.175 4.673 ;
      RECT 22.885 4.52 23.21 4.658 ;
      RECT 23.14 4.44 23.33 4.65 ;
      RECT 23.13 4.445 23.34 4.643 ;
      RECT 23.095 4.515 23.34 4.643 ;
      RECT 23.125 4.457 23.145 4.78 ;
      RECT 23.11 4.505 23.34 4.643 ;
      RECT 23.115 4.477 23.145 4.78 ;
      RECT 22.195 3.545 22.265 4.65 ;
      RECT 22.93 3.65 23.19 3.91 ;
      RECT 22.51 3.696 22.525 3.905 ;
      RECT 22.846 3.709 22.93 3.86 ;
      RECT 22.76 3.706 22.846 3.86 ;
      RECT 22.721 3.704 22.76 3.86 ;
      RECT 22.635 3.702 22.721 3.86 ;
      RECT 22.575 3.7 22.635 3.871 ;
      RECT 22.54 3.698 22.575 3.889 ;
      RECT 22.525 3.696 22.54 3.9 ;
      RECT 22.495 3.696 22.51 3.913 ;
      RECT 22.485 3.696 22.495 3.918 ;
      RECT 22.46 3.695 22.485 3.923 ;
      RECT 22.445 3.69 22.46 3.929 ;
      RECT 22.44 3.683 22.445 3.934 ;
      RECT 22.415 3.674 22.44 3.94 ;
      RECT 22.37 3.653 22.415 3.953 ;
      RECT 22.36 3.637 22.37 3.963 ;
      RECT 22.345 3.63 22.36 3.973 ;
      RECT 22.335 3.623 22.345 3.99 ;
      RECT 22.33 3.62 22.335 4.02 ;
      RECT 22.325 3.618 22.33 4.05 ;
      RECT 22.32 3.616 22.325 4.087 ;
      RECT 22.305 3.612 22.32 4.154 ;
      RECT 22.305 4.445 22.315 4.645 ;
      RECT 22.3 3.608 22.305 4.28 ;
      RECT 22.3 4.432 22.305 4.65 ;
      RECT 22.295 3.606 22.3 4.365 ;
      RECT 22.295 4.422 22.3 4.65 ;
      RECT 22.28 3.577 22.295 4.65 ;
      RECT 22.265 3.55 22.28 4.65 ;
      RECT 22.19 3.545 22.195 3.9 ;
      RECT 22.19 3.955 22.195 4.65 ;
      RECT 22.175 3.545 22.19 3.878 ;
      RECT 22.185 3.977 22.19 4.65 ;
      RECT 22.175 4.017 22.185 4.65 ;
      RECT 22.14 3.545 22.175 3.82 ;
      RECT 22.17 4.052 22.175 4.65 ;
      RECT 22.155 4.107 22.17 4.65 ;
      RECT 22.15 4.172 22.155 4.65 ;
      RECT 22.135 4.22 22.15 4.65 ;
      RECT 22.11 3.545 22.14 3.775 ;
      RECT 22.13 4.275 22.135 4.65 ;
      RECT 22.115 4.335 22.13 4.65 ;
      RECT 22.11 4.383 22.115 4.648 ;
      RECT 22.105 3.545 22.11 3.768 ;
      RECT 22.105 4.415 22.11 4.643 ;
      RECT 22.08 3.545 22.105 3.76 ;
      RECT 22.07 3.55 22.08 3.75 ;
      RECT 22.285 4.825 22.305 5.065 ;
      RECT 21.515 4.755 21.52 4.965 ;
      RECT 22.795 4.828 22.805 5.023 ;
      RECT 22.79 4.818 22.795 5.026 ;
      RECT 22.71 4.815 22.79 5.049 ;
      RECT 22.706 4.815 22.71 5.071 ;
      RECT 22.62 4.815 22.706 5.081 ;
      RECT 22.605 4.815 22.62 5.089 ;
      RECT 22.576 4.816 22.605 5.087 ;
      RECT 22.49 4.821 22.576 5.083 ;
      RECT 22.477 4.825 22.49 5.079 ;
      RECT 22.391 4.825 22.477 5.075 ;
      RECT 22.305 4.825 22.391 5.069 ;
      RECT 22.221 4.825 22.285 5.063 ;
      RECT 22.135 4.825 22.221 5.058 ;
      RECT 22.115 4.825 22.135 5.054 ;
      RECT 22.055 4.82 22.115 5.051 ;
      RECT 22.027 4.814 22.055 5.048 ;
      RECT 21.941 4.809 22.027 5.044 ;
      RECT 21.855 4.803 21.941 5.038 ;
      RECT 21.78 4.785 21.855 5.033 ;
      RECT 21.745 4.762 21.78 5.029 ;
      RECT 21.735 4.752 21.745 5.028 ;
      RECT 21.68 4.75 21.735 5.027 ;
      RECT 21.605 4.75 21.68 5.023 ;
      RECT 21.595 4.75 21.605 5.018 ;
      RECT 21.58 4.75 21.595 5.01 ;
      RECT 21.53 4.752 21.58 4.988 ;
      RECT 21.52 4.755 21.53 4.968 ;
      RECT 21.51 4.76 21.515 4.963 ;
      RECT 21.505 4.765 21.51 4.958 ;
      RECT 19.615 3.41 19.875 3.67 ;
      RECT 19.605 3.44 19.875 3.65 ;
      RECT 21.525 3.355 21.785 3.615 ;
      RECT 21.52 3.43 21.525 3.616 ;
      RECT 21.495 3.435 21.52 3.618 ;
      RECT 21.48 3.442 21.495 3.621 ;
      RECT 21.42 3.46 21.48 3.626 ;
      RECT 21.39 3.48 21.42 3.633 ;
      RECT 21.365 3.488 21.39 3.638 ;
      RECT 21.34 3.496 21.365 3.64 ;
      RECT 21.322 3.5 21.34 3.639 ;
      RECT 21.236 3.498 21.322 3.639 ;
      RECT 21.15 3.496 21.236 3.639 ;
      RECT 21.064 3.494 21.15 3.638 ;
      RECT 20.978 3.492 21.064 3.638 ;
      RECT 20.892 3.49 20.978 3.638 ;
      RECT 20.806 3.488 20.892 3.638 ;
      RECT 20.72 3.486 20.806 3.637 ;
      RECT 20.702 3.485 20.72 3.637 ;
      RECT 20.616 3.484 20.702 3.637 ;
      RECT 20.53 3.482 20.616 3.637 ;
      RECT 20.444 3.481 20.53 3.636 ;
      RECT 20.358 3.48 20.444 3.636 ;
      RECT 20.272 3.478 20.358 3.636 ;
      RECT 20.186 3.477 20.272 3.636 ;
      RECT 20.1 3.475 20.186 3.635 ;
      RECT 20.076 3.473 20.1 3.635 ;
      RECT 19.99 3.466 20.076 3.635 ;
      RECT 19.961 3.458 19.99 3.635 ;
      RECT 19.875 3.45 19.961 3.635 ;
      RECT 19.595 3.447 19.605 3.645 ;
      RECT 21.1 4.41 21.105 4.76 ;
      RECT 20.87 4.5 21.01 4.76 ;
      RECT 21.345 4.185 21.39 4.395 ;
      RECT 21.4 4.196 21.41 4.39 ;
      RECT 21.39 4.188 21.4 4.395 ;
      RECT 21.325 4.185 21.345 4.4 ;
      RECT 21.295 4.185 21.325 4.423 ;
      RECT 21.285 4.185 21.295 4.448 ;
      RECT 21.28 4.185 21.285 4.458 ;
      RECT 21.225 4.185 21.28 4.498 ;
      RECT 21.22 4.185 21.225 4.538 ;
      RECT 21.215 4.187 21.22 4.543 ;
      RECT 21.2 4.197 21.215 4.554 ;
      RECT 21.155 4.255 21.2 4.59 ;
      RECT 21.145 4.31 21.155 4.624 ;
      RECT 21.13 4.337 21.145 4.64 ;
      RECT 21.12 4.364 21.13 4.76 ;
      RECT 21.105 4.387 21.12 4.76 ;
      RECT 21.095 4.427 21.1 4.76 ;
      RECT 21.09 4.437 21.095 4.76 ;
      RECT 21.085 4.452 21.09 4.76 ;
      RECT 21.075 4.457 21.085 4.76 ;
      RECT 21.01 4.48 21.075 4.76 ;
      RECT 20.48 3.875 20.71 4.185 ;
      RECT 20.38 3.875 20.71 4.165 ;
      RECT 19.085 3.9 19.345 4.16 ;
      RECT 20.21 3.875 20.71 4.155 ;
      RECT 20.025 3.875 20.71 4.145 ;
      RECT 19.84 3.925 20.71 4.135 ;
      RECT 19.72 3.925 20.71 4.125 ;
      RECT 19.39 3.925 20.71 4.115 ;
      RECT 19.385 3.925 20.71 4.101 ;
      RECT 19.085 3.915 19.67 4.098 ;
      RECT 19.955 3.875 20.77 4.015 ;
      RECT 19.39 3.91 19.66 4.115 ;
      RECT 19.39 3.895 19.65 4.115 ;
      RECT 19.6 4.415 19.86 4.675 ;
      RECT 19.6 4.455 19.965 4.665 ;
      RECT 19.6 4.457 19.97 4.664 ;
      RECT 19.6 4.465 19.975 4.661 ;
      RECT 18.525 3.54 18.625 5.065 ;
      RECT 18.715 4.68 18.765 4.94 ;
      RECT 18.71 3.553 18.715 3.74 ;
      RECT 18.705 4.661 18.715 4.94 ;
      RECT 18.705 3.55 18.71 3.748 ;
      RECT 18.69 3.544 18.705 3.755 ;
      RECT 18.7 4.649 18.705 5.023 ;
      RECT 18.69 4.637 18.7 5.06 ;
      RECT 18.68 3.54 18.69 3.762 ;
      RECT 18.68 4.622 18.69 5.065 ;
      RECT 18.675 3.54 18.68 3.77 ;
      RECT 18.655 4.592 18.68 5.065 ;
      RECT 18.635 3.54 18.675 3.818 ;
      RECT 18.645 4.552 18.655 5.065 ;
      RECT 18.635 4.507 18.645 5.065 ;
      RECT 18.63 3.54 18.635 3.888 ;
      RECT 18.63 4.465 18.635 5.065 ;
      RECT 18.625 3.54 18.63 4.365 ;
      RECT 18.625 4.447 18.63 5.065 ;
      RECT 18.515 3.543 18.525 5.065 ;
      RECT 18.5 3.55 18.515 5.061 ;
      RECT 18.495 3.56 18.5 5.056 ;
      RECT 18.49 3.76 18.495 4.948 ;
      RECT 18.485 3.845 18.49 4.5 ;
      RECT 16.705 10.205 16.995 10.435 ;
      RECT 16.765 9.46 16.935 10.435 ;
      RECT 16.675 9.46 17.025 9.75 ;
      RECT 16.3 8.72 16.65 9.01 ;
      RECT 16.16 8.755 16.65 8.925 ;
      RECT 106.94 7.35 107.315 7.73 ;
      RECT 102.215 2.435 102.59 2.805 ;
      RECT 96.195 3.52 96.455 3.78 ;
      RECT 89.015 7.35 89.39 7.73 ;
      RECT 84.29 2.435 84.665 2.805 ;
      RECT 78.27 3.52 78.53 3.78 ;
      RECT 71.09 7.35 71.465 7.73 ;
      RECT 66.365 2.435 66.74 2.805 ;
      RECT 60.345 3.52 60.605 3.78 ;
      RECT 53.165 7.35 53.54 7.73 ;
      RECT 48.44 2.435 48.815 2.805 ;
      RECT 42.42 3.52 42.68 3.78 ;
      RECT 35.24 7.35 35.615 7.73 ;
      RECT 30.515 2.435 30.89 2.805 ;
      RECT 24.495 3.52 24.755 3.78 ;
    LAYER mcon ;
      RECT 107.04 7.455 107.21 7.625 ;
      RECT 107.035 8.755 107.205 8.925 ;
      RECT 107.035 10.235 107.205 10.405 ;
      RECT 106.665 8.385 106.835 8.555 ;
      RECT 106.66 4.055 106.83 4.225 ;
      RECT 106.045 2.205 106.215 2.375 ;
      RECT 106.045 3.685 106.215 3.855 ;
      RECT 106.045 8.755 106.215 8.925 ;
      RECT 106.045 10.235 106.215 10.405 ;
      RECT 105.675 4.055 105.845 4.225 ;
      RECT 105.675 8.385 105.845 8.555 ;
      RECT 104.685 3.315 104.855 3.485 ;
      RECT 104.685 9.125 104.855 9.295 ;
      RECT 104.255 2.205 104.425 2.375 ;
      RECT 104.255 2.945 104.425 3.115 ;
      RECT 104.255 9.495 104.425 9.665 ;
      RECT 104.255 10.235 104.425 10.405 ;
      RECT 103.885 3.685 104.055 3.855 ;
      RECT 103.885 8.755 104.055 8.925 ;
      RECT 100.83 4.2 101 4.37 ;
      RECT 100.62 3.54 100.79 3.71 ;
      RECT 100.305 4.45 100.475 4.62 ;
      RECT 99.925 9.125 100.095 9.295 ;
      RECT 99.92 4.045 100.09 4.215 ;
      RECT 99.705 4.61 99.875 4.78 ;
      RECT 99.685 5.01 99.855 5.18 ;
      RECT 99.51 3.565 99.68 3.735 ;
      RECT 99.495 9.495 99.665 9.665 ;
      RECT 99.495 10.235 99.665 10.405 ;
      RECT 99.015 4.545 99.185 4.715 ;
      RECT 98.69 4.23 98.86 4.4 ;
      RECT 98.625 5.01 98.795 5.18 ;
      RECT 98.225 4.995 98.395 5.165 ;
      RECT 98.185 3.48 98.355 3.65 ;
      RECT 97.285 3.98 97.455 4.15 ;
      RECT 97.285 4.44 97.455 4.61 ;
      RECT 97.285 4.955 97.455 5.125 ;
      RECT 97.17 3.515 97.34 3.685 ;
      RECT 96.705 5.025 96.875 5.195 ;
      RECT 96.225 3.555 96.395 3.725 ;
      RECT 96.01 3.93 96.18 4.1 ;
      RECT 95.51 4.53 95.68 4.7 ;
      RECT 95.395 3.98 95.565 4.15 ;
      RECT 95.225 3.43 95.395 3.6 ;
      RECT 94.85 4.46 95.02 4.63 ;
      RECT 94.365 4.06 94.535 4.23 ;
      RECT 94.315 4.835 94.485 5.005 ;
      RECT 93.825 4.46 93.995 4.63 ;
      RECT 93.79 3.565 93.96 3.735 ;
      RECT 93.225 4.775 93.395 4.945 ;
      RECT 92.92 4.205 93.09 4.375 ;
      RECT 92.22 3.995 92.39 4.165 ;
      RECT 91.485 4.475 91.655 4.645 ;
      RECT 91.315 3.46 91.485 3.63 ;
      RECT 91.14 3.915 91.31 4.085 ;
      RECT 90.22 3.565 90.39 3.735 ;
      RECT 90.215 4.88 90.385 5.05 ;
      RECT 89.115 7.455 89.285 7.625 ;
      RECT 89.11 8.755 89.28 8.925 ;
      RECT 89.11 10.235 89.28 10.405 ;
      RECT 88.74 8.385 88.91 8.555 ;
      RECT 88.735 4.055 88.905 4.225 ;
      RECT 88.12 2.205 88.29 2.375 ;
      RECT 88.12 3.685 88.29 3.855 ;
      RECT 88.12 8.755 88.29 8.925 ;
      RECT 88.12 10.235 88.29 10.405 ;
      RECT 87.75 4.055 87.92 4.225 ;
      RECT 87.75 8.385 87.92 8.555 ;
      RECT 86.76 3.315 86.93 3.485 ;
      RECT 86.76 9.125 86.93 9.295 ;
      RECT 86.33 2.205 86.5 2.375 ;
      RECT 86.33 2.945 86.5 3.115 ;
      RECT 86.33 9.495 86.5 9.665 ;
      RECT 86.33 10.235 86.5 10.405 ;
      RECT 85.96 3.685 86.13 3.855 ;
      RECT 85.96 8.755 86.13 8.925 ;
      RECT 82.905 4.2 83.075 4.37 ;
      RECT 82.695 3.54 82.865 3.71 ;
      RECT 82.38 4.45 82.55 4.62 ;
      RECT 82 9.125 82.17 9.295 ;
      RECT 81.995 4.045 82.165 4.215 ;
      RECT 81.78 4.61 81.95 4.78 ;
      RECT 81.76 5.01 81.93 5.18 ;
      RECT 81.585 3.565 81.755 3.735 ;
      RECT 81.57 9.495 81.74 9.665 ;
      RECT 81.57 10.235 81.74 10.405 ;
      RECT 81.09 4.545 81.26 4.715 ;
      RECT 80.765 4.23 80.935 4.4 ;
      RECT 80.7 5.01 80.87 5.18 ;
      RECT 80.3 4.995 80.47 5.165 ;
      RECT 80.26 3.48 80.43 3.65 ;
      RECT 79.36 3.98 79.53 4.15 ;
      RECT 79.36 4.44 79.53 4.61 ;
      RECT 79.36 4.955 79.53 5.125 ;
      RECT 79.245 3.515 79.415 3.685 ;
      RECT 78.78 5.025 78.95 5.195 ;
      RECT 78.3 3.555 78.47 3.725 ;
      RECT 78.085 3.93 78.255 4.1 ;
      RECT 77.585 4.53 77.755 4.7 ;
      RECT 77.47 3.98 77.64 4.15 ;
      RECT 77.3 3.43 77.47 3.6 ;
      RECT 76.925 4.46 77.095 4.63 ;
      RECT 76.44 4.06 76.61 4.23 ;
      RECT 76.39 4.835 76.56 5.005 ;
      RECT 75.9 4.46 76.07 4.63 ;
      RECT 75.865 3.565 76.035 3.735 ;
      RECT 75.3 4.775 75.47 4.945 ;
      RECT 74.995 4.205 75.165 4.375 ;
      RECT 74.295 3.995 74.465 4.165 ;
      RECT 73.56 4.475 73.73 4.645 ;
      RECT 73.39 3.46 73.56 3.63 ;
      RECT 73.215 3.915 73.385 4.085 ;
      RECT 72.295 3.565 72.465 3.735 ;
      RECT 72.29 4.88 72.46 5.05 ;
      RECT 71.19 7.455 71.36 7.625 ;
      RECT 71.185 8.755 71.355 8.925 ;
      RECT 71.185 10.235 71.355 10.405 ;
      RECT 70.815 8.385 70.985 8.555 ;
      RECT 70.81 4.055 70.98 4.225 ;
      RECT 70.195 2.205 70.365 2.375 ;
      RECT 70.195 3.685 70.365 3.855 ;
      RECT 70.195 8.755 70.365 8.925 ;
      RECT 70.195 10.235 70.365 10.405 ;
      RECT 69.825 4.055 69.995 4.225 ;
      RECT 69.825 8.385 69.995 8.555 ;
      RECT 68.835 3.315 69.005 3.485 ;
      RECT 68.835 9.125 69.005 9.295 ;
      RECT 68.405 2.205 68.575 2.375 ;
      RECT 68.405 2.945 68.575 3.115 ;
      RECT 68.405 9.495 68.575 9.665 ;
      RECT 68.405 10.235 68.575 10.405 ;
      RECT 68.035 3.685 68.205 3.855 ;
      RECT 68.035 8.755 68.205 8.925 ;
      RECT 64.98 4.2 65.15 4.37 ;
      RECT 64.77 3.54 64.94 3.71 ;
      RECT 64.455 4.45 64.625 4.62 ;
      RECT 64.075 9.125 64.245 9.295 ;
      RECT 64.07 4.045 64.24 4.215 ;
      RECT 63.855 4.61 64.025 4.78 ;
      RECT 63.835 5.01 64.005 5.18 ;
      RECT 63.66 3.565 63.83 3.735 ;
      RECT 63.645 9.495 63.815 9.665 ;
      RECT 63.645 10.235 63.815 10.405 ;
      RECT 63.165 4.545 63.335 4.715 ;
      RECT 62.84 4.23 63.01 4.4 ;
      RECT 62.775 5.01 62.945 5.18 ;
      RECT 62.375 4.995 62.545 5.165 ;
      RECT 62.335 3.48 62.505 3.65 ;
      RECT 61.435 3.98 61.605 4.15 ;
      RECT 61.435 4.44 61.605 4.61 ;
      RECT 61.435 4.955 61.605 5.125 ;
      RECT 61.32 3.515 61.49 3.685 ;
      RECT 60.855 5.025 61.025 5.195 ;
      RECT 60.375 3.555 60.545 3.725 ;
      RECT 60.16 3.93 60.33 4.1 ;
      RECT 59.66 4.53 59.83 4.7 ;
      RECT 59.545 3.98 59.715 4.15 ;
      RECT 59.375 3.43 59.545 3.6 ;
      RECT 59 4.46 59.17 4.63 ;
      RECT 58.515 4.06 58.685 4.23 ;
      RECT 58.465 4.835 58.635 5.005 ;
      RECT 57.975 4.46 58.145 4.63 ;
      RECT 57.94 3.565 58.11 3.735 ;
      RECT 57.375 4.775 57.545 4.945 ;
      RECT 57.07 4.205 57.24 4.375 ;
      RECT 56.37 3.995 56.54 4.165 ;
      RECT 55.635 4.475 55.805 4.645 ;
      RECT 55.465 3.46 55.635 3.63 ;
      RECT 55.29 3.915 55.46 4.085 ;
      RECT 54.37 3.565 54.54 3.735 ;
      RECT 54.365 4.88 54.535 5.05 ;
      RECT 53.265 7.455 53.435 7.625 ;
      RECT 53.26 8.755 53.43 8.925 ;
      RECT 53.26 10.235 53.43 10.405 ;
      RECT 52.89 8.385 53.06 8.555 ;
      RECT 52.885 4.055 53.055 4.225 ;
      RECT 52.27 2.205 52.44 2.375 ;
      RECT 52.27 3.685 52.44 3.855 ;
      RECT 52.27 8.755 52.44 8.925 ;
      RECT 52.27 10.235 52.44 10.405 ;
      RECT 51.9 4.055 52.07 4.225 ;
      RECT 51.9 8.385 52.07 8.555 ;
      RECT 50.91 3.315 51.08 3.485 ;
      RECT 50.91 9.125 51.08 9.295 ;
      RECT 50.48 2.205 50.65 2.375 ;
      RECT 50.48 2.945 50.65 3.115 ;
      RECT 50.48 9.495 50.65 9.665 ;
      RECT 50.48 10.235 50.65 10.405 ;
      RECT 50.11 3.685 50.28 3.855 ;
      RECT 50.11 8.755 50.28 8.925 ;
      RECT 47.055 4.2 47.225 4.37 ;
      RECT 46.845 3.54 47.015 3.71 ;
      RECT 46.53 4.45 46.7 4.62 ;
      RECT 46.15 9.125 46.32 9.295 ;
      RECT 46.145 4.045 46.315 4.215 ;
      RECT 45.93 4.61 46.1 4.78 ;
      RECT 45.91 5.01 46.08 5.18 ;
      RECT 45.735 3.565 45.905 3.735 ;
      RECT 45.72 9.495 45.89 9.665 ;
      RECT 45.72 10.235 45.89 10.405 ;
      RECT 45.24 4.545 45.41 4.715 ;
      RECT 44.915 4.23 45.085 4.4 ;
      RECT 44.85 5.01 45.02 5.18 ;
      RECT 44.45 4.995 44.62 5.165 ;
      RECT 44.41 3.48 44.58 3.65 ;
      RECT 43.51 3.98 43.68 4.15 ;
      RECT 43.51 4.44 43.68 4.61 ;
      RECT 43.51 4.955 43.68 5.125 ;
      RECT 43.395 3.515 43.565 3.685 ;
      RECT 42.93 5.025 43.1 5.195 ;
      RECT 42.45 3.555 42.62 3.725 ;
      RECT 42.235 3.93 42.405 4.1 ;
      RECT 41.735 4.53 41.905 4.7 ;
      RECT 41.62 3.98 41.79 4.15 ;
      RECT 41.45 3.43 41.62 3.6 ;
      RECT 41.075 4.46 41.245 4.63 ;
      RECT 40.59 4.06 40.76 4.23 ;
      RECT 40.54 4.835 40.71 5.005 ;
      RECT 40.05 4.46 40.22 4.63 ;
      RECT 40.015 3.565 40.185 3.735 ;
      RECT 39.45 4.775 39.62 4.945 ;
      RECT 39.145 4.205 39.315 4.375 ;
      RECT 38.445 3.995 38.615 4.165 ;
      RECT 37.71 4.475 37.88 4.645 ;
      RECT 37.54 3.46 37.71 3.63 ;
      RECT 37.365 3.915 37.535 4.085 ;
      RECT 36.445 3.565 36.615 3.735 ;
      RECT 36.44 4.88 36.61 5.05 ;
      RECT 35.34 7.455 35.51 7.625 ;
      RECT 35.335 8.755 35.505 8.925 ;
      RECT 35.335 10.235 35.505 10.405 ;
      RECT 34.965 8.385 35.135 8.555 ;
      RECT 34.96 4.055 35.13 4.225 ;
      RECT 34.345 2.205 34.515 2.375 ;
      RECT 34.345 3.685 34.515 3.855 ;
      RECT 34.345 8.755 34.515 8.925 ;
      RECT 34.345 10.235 34.515 10.405 ;
      RECT 33.975 4.055 34.145 4.225 ;
      RECT 33.975 8.385 34.145 8.555 ;
      RECT 32.985 3.315 33.155 3.485 ;
      RECT 32.985 9.125 33.155 9.295 ;
      RECT 32.555 2.205 32.725 2.375 ;
      RECT 32.555 2.945 32.725 3.115 ;
      RECT 32.555 9.495 32.725 9.665 ;
      RECT 32.555 10.235 32.725 10.405 ;
      RECT 32.185 3.685 32.355 3.855 ;
      RECT 32.185 8.755 32.355 8.925 ;
      RECT 29.13 4.2 29.3 4.37 ;
      RECT 28.92 3.54 29.09 3.71 ;
      RECT 28.605 4.45 28.775 4.62 ;
      RECT 28.225 9.125 28.395 9.295 ;
      RECT 28.22 4.045 28.39 4.215 ;
      RECT 28.005 4.61 28.175 4.78 ;
      RECT 27.985 5.01 28.155 5.18 ;
      RECT 27.81 3.565 27.98 3.735 ;
      RECT 27.795 9.495 27.965 9.665 ;
      RECT 27.795 10.235 27.965 10.405 ;
      RECT 27.315 4.545 27.485 4.715 ;
      RECT 26.99 4.23 27.16 4.4 ;
      RECT 26.925 5.01 27.095 5.18 ;
      RECT 26.525 4.995 26.695 5.165 ;
      RECT 26.485 3.48 26.655 3.65 ;
      RECT 25.585 3.98 25.755 4.15 ;
      RECT 25.585 4.44 25.755 4.61 ;
      RECT 25.585 4.955 25.755 5.125 ;
      RECT 25.47 3.515 25.64 3.685 ;
      RECT 25.005 5.025 25.175 5.195 ;
      RECT 24.525 3.555 24.695 3.725 ;
      RECT 24.31 3.93 24.48 4.1 ;
      RECT 23.81 4.53 23.98 4.7 ;
      RECT 23.695 3.98 23.865 4.15 ;
      RECT 23.525 3.43 23.695 3.6 ;
      RECT 23.15 4.46 23.32 4.63 ;
      RECT 22.665 4.06 22.835 4.23 ;
      RECT 22.615 4.835 22.785 5.005 ;
      RECT 22.125 4.46 22.295 4.63 ;
      RECT 22.09 3.565 22.26 3.735 ;
      RECT 21.525 4.775 21.695 4.945 ;
      RECT 21.22 4.205 21.39 4.375 ;
      RECT 20.52 3.995 20.69 4.165 ;
      RECT 19.785 4.475 19.955 4.645 ;
      RECT 19.615 3.46 19.785 3.63 ;
      RECT 19.44 3.915 19.61 4.085 ;
      RECT 18.52 3.565 18.69 3.735 ;
      RECT 18.515 4.88 18.685 5.05 ;
      RECT 16.765 9.495 16.935 9.665 ;
      RECT 16.765 10.235 16.935 10.405 ;
      RECT 16.395 8.755 16.565 8.925 ;
    LAYER li1 ;
      RECT 107.035 7.455 107.205 8.925 ;
      RECT 107.035 7.455 107.21 8.715 ;
      RECT 106.665 9.405 107.135 9.575 ;
      RECT 106.665 8.385 106.835 9.575 ;
      RECT 106.66 3.035 106.83 4.225 ;
      RECT 106.66 3.035 107.13 3.205 ;
      RECT 106.045 3.895 106.22 5.155 ;
      RECT 106.045 3.685 106.215 5.155 ;
      RECT 106.045 7.455 106.215 8.925 ;
      RECT 106.045 7.455 106.22 8.715 ;
      RECT 105.675 3.035 105.845 4.225 ;
      RECT 105.675 3.035 106.145 3.205 ;
      RECT 105.675 9.405 106.145 9.575 ;
      RECT 105.675 8.385 105.845 9.575 ;
      RECT 104.685 4.015 104.86 5.155 ;
      RECT 104.685 1.865 104.855 5.155 ;
      RECT 104.685 1.865 104.86 2.415 ;
      RECT 104.685 10.195 104.86 10.745 ;
      RECT 104.685 7.455 104.855 10.745 ;
      RECT 104.685 7.455 104.86 8.595 ;
      RECT 104.255 3.895 104.43 5.155 ;
      RECT 104.255 2.945 104.425 5.155 ;
      RECT 104.255 7.455 104.425 9.665 ;
      RECT 104.255 7.455 104.43 8.715 ;
      RECT 103.825 3.925 103.995 5.155 ;
      RECT 103.885 2.145 104.055 4.095 ;
      RECT 103.825 1.865 103.995 2.315 ;
      RECT 103.825 10.295 103.995 10.745 ;
      RECT 103.885 8.515 104.055 10.465 ;
      RECT 103.825 7.455 103.995 8.685 ;
      RECT 103.3 3.895 103.475 5.155 ;
      RECT 103.3 1.865 103.47 5.155 ;
      RECT 103.3 3.365 103.71 3.695 ;
      RECT 103.3 2.525 103.71 2.855 ;
      RECT 103.3 1.865 103.475 2.355 ;
      RECT 103.3 10.255 103.475 10.745 ;
      RECT 103.3 7.455 103.47 10.745 ;
      RECT 103.3 9.755 103.71 10.085 ;
      RECT 103.3 8.915 103.71 9.245 ;
      RECT 103.3 7.455 103.475 8.715 ;
      RECT 101.415 4.687 101.43 4.738 ;
      RECT 101.41 4.667 101.415 4.785 ;
      RECT 101.395 4.657 101.41 4.853 ;
      RECT 101.37 4.637 101.395 4.908 ;
      RECT 101.33 4.622 101.37 4.928 ;
      RECT 101.285 4.616 101.33 4.956 ;
      RECT 101.215 4.606 101.285 4.973 ;
      RECT 101.195 4.598 101.215 4.973 ;
      RECT 101.135 4.592 101.195 4.965 ;
      RECT 101.076 4.583 101.135 4.953 ;
      RECT 100.99 4.572 101.076 4.936 ;
      RECT 100.968 4.563 100.99 4.924 ;
      RECT 100.882 4.556 100.968 4.911 ;
      RECT 100.796 4.543 100.882 4.892 ;
      RECT 100.71 4.531 100.796 4.872 ;
      RECT 100.68 4.52 100.71 4.859 ;
      RECT 100.63 4.506 100.68 4.851 ;
      RECT 100.61 4.495 100.63 4.843 ;
      RECT 100.561 4.484 100.61 4.835 ;
      RECT 100.475 4.463 100.561 4.82 ;
      RECT 100.43 4.45 100.475 4.805 ;
      RECT 100.385 4.45 100.43 4.785 ;
      RECT 100.33 4.45 100.385 4.72 ;
      RECT 100.305 4.45 100.33 4.643 ;
      RECT 100.83 4.187 101 4.37 ;
      RECT 100.83 4.187 101.015 4.328 ;
      RECT 100.83 4.187 101.02 4.27 ;
      RECT 100.89 3.955 101.025 4.246 ;
      RECT 100.89 3.959 101.03 4.229 ;
      RECT 100.835 4.122 101.03 4.229 ;
      RECT 100.86 3.967 101 4.37 ;
      RECT 100.86 3.971 101.04 4.17 ;
      RECT 100.845 4.057 101.04 4.17 ;
      RECT 100.855 3.987 101 4.37 ;
      RECT 100.855 3.99 101.05 4.083 ;
      RECT 100.85 4.007 101.05 4.083 ;
      RECT 100.62 3.227 100.79 3.71 ;
      RECT 100.615 3.222 100.765 3.7 ;
      RECT 100.615 3.229 100.795 3.694 ;
      RECT 100.605 3.223 100.765 3.673 ;
      RECT 100.605 3.239 100.81 3.632 ;
      RECT 100.575 3.224 100.765 3.595 ;
      RECT 100.575 3.254 100.82 3.535 ;
      RECT 100.57 3.226 100.765 3.533 ;
      RECT 100.55 3.235 100.795 3.49 ;
      RECT 100.525 3.251 100.81 3.402 ;
      RECT 100.525 3.27 100.835 3.393 ;
      RECT 100.52 3.307 100.835 3.345 ;
      RECT 100.525 3.287 100.84 3.313 ;
      RECT 100.62 3.221 100.73 3.71 ;
      RECT 100.706 3.22 100.73 3.71 ;
      RECT 99.94 4.005 99.945 4.216 ;
      RECT 100.54 4.005 100.545 4.19 ;
      RECT 100.605 4.045 100.61 4.158 ;
      RECT 100.6 4.037 100.605 4.164 ;
      RECT 100.595 4.027 100.6 4.172 ;
      RECT 100.59 4.017 100.595 4.181 ;
      RECT 100.585 4.007 100.59 4.185 ;
      RECT 100.545 4.005 100.585 4.188 ;
      RECT 100.517 4.004 100.54 4.192 ;
      RECT 100.431 4.001 100.517 4.199 ;
      RECT 100.345 3.997 100.431 4.21 ;
      RECT 100.325 3.995 100.345 4.216 ;
      RECT 100.307 3.994 100.325 4.219 ;
      RECT 100.221 3.992 100.307 4.226 ;
      RECT 100.135 3.987 100.221 4.239 ;
      RECT 100.116 3.984 100.135 4.244 ;
      RECT 100.03 3.982 100.116 4.235 ;
      RECT 100.02 3.982 100.03 4.228 ;
      RECT 99.945 3.995 100.02 4.222 ;
      RECT 99.93 4.006 99.94 4.216 ;
      RECT 99.92 4.008 99.93 4.215 ;
      RECT 99.91 4.012 99.92 4.211 ;
      RECT 99.905 4.015 99.91 4.205 ;
      RECT 99.895 4.017 99.905 4.199 ;
      RECT 99.89 4.02 99.895 4.193 ;
      RECT 99.925 10.195 100.1 10.745 ;
      RECT 99.925 7.455 100.095 10.745 ;
      RECT 99.925 7.455 100.1 8.595 ;
      RECT 99.87 4.606 99.875 4.81 ;
      RECT 99.855 4.593 99.87 4.903 ;
      RECT 99.84 4.574 99.855 5.18 ;
      RECT 99.805 4.54 99.84 5.18 ;
      RECT 99.801 4.51 99.805 5.18 ;
      RECT 99.715 4.392 99.801 5.18 ;
      RECT 99.705 4.267 99.715 5.18 ;
      RECT 99.69 4.235 99.705 5.18 ;
      RECT 99.685 4.21 99.69 5.18 ;
      RECT 99.68 4.2 99.685 5.136 ;
      RECT 99.665 4.172 99.68 5.041 ;
      RECT 99.65 4.138 99.665 4.94 ;
      RECT 99.645 4.116 99.65 4.893 ;
      RECT 99.64 4.105 99.645 4.863 ;
      RECT 99.635 4.095 99.64 4.829 ;
      RECT 99.625 4.082 99.635 4.797 ;
      RECT 99.6 4.058 99.625 4.723 ;
      RECT 99.595 4.038 99.6 4.648 ;
      RECT 99.59 4.032 99.595 4.623 ;
      RECT 99.585 4.027 99.59 4.588 ;
      RECT 99.58 4.022 99.585 4.563 ;
      RECT 99.575 4.02 99.58 4.543 ;
      RECT 99.57 4.02 99.575 4.528 ;
      RECT 99.565 4.02 99.57 4.488 ;
      RECT 99.555 4.02 99.565 4.46 ;
      RECT 99.545 4.02 99.555 4.405 ;
      RECT 99.53 4.02 99.545 4.343 ;
      RECT 99.525 4.019 99.53 4.288 ;
      RECT 99.51 4.018 99.525 4.268 ;
      RECT 99.45 4.016 99.51 4.242 ;
      RECT 99.415 4.017 99.45 4.222 ;
      RECT 99.41 4.019 99.415 4.212 ;
      RECT 99.4 4.038 99.41 4.202 ;
      RECT 99.395 4.065 99.4 4.133 ;
      RECT 99.51 3.49 99.68 3.735 ;
      RECT 99.545 3.261 99.68 3.735 ;
      RECT 99.545 3.263 99.69 3.73 ;
      RECT 99.545 3.265 99.715 3.718 ;
      RECT 99.545 3.268 99.74 3.7 ;
      RECT 99.545 3.273 99.79 3.673 ;
      RECT 99.545 3.278 99.81 3.638 ;
      RECT 99.525 3.28 99.82 3.613 ;
      RECT 99.515 3.375 99.82 3.613 ;
      RECT 99.545 3.26 99.655 3.735 ;
      RECT 99.555 3.257 99.65 3.735 ;
      RECT 99.495 7.455 99.665 9.665 ;
      RECT 99.495 7.455 99.67 8.715 ;
      RECT 99.075 4.522 99.265 4.88 ;
      RECT 99.075 4.534 99.3 4.879 ;
      RECT 99.075 4.562 99.32 4.877 ;
      RECT 99.075 4.587 99.325 4.876 ;
      RECT 99.075 4.645 99.34 4.875 ;
      RECT 99.06 4.518 99.22 4.86 ;
      RECT 99.04 4.527 99.265 4.813 ;
      RECT 99.015 4.538 99.3 4.75 ;
      RECT 99.015 4.622 99.335 4.75 ;
      RECT 99.015 4.597 99.33 4.75 ;
      RECT 99.075 4.513 99.22 4.88 ;
      RECT 99.161 4.512 99.22 4.88 ;
      RECT 99.161 4.511 99.205 4.88 ;
      RECT 98.54 10.255 98.715 10.745 ;
      RECT 98.54 7.455 98.71 10.745 ;
      RECT 98.54 9.755 98.95 10.085 ;
      RECT 98.54 8.915 98.95 9.245 ;
      RECT 98.54 7.455 98.715 8.715 ;
      RECT 98.86 4.027 98.865 4.405 ;
      RECT 98.855 3.995 98.86 4.405 ;
      RECT 98.85 3.967 98.855 4.405 ;
      RECT 98.845 3.947 98.85 4.405 ;
      RECT 98.79 3.93 98.845 4.405 ;
      RECT 98.75 3.915 98.79 4.405 ;
      RECT 98.695 3.902 98.75 4.405 ;
      RECT 98.66 3.893 98.695 4.405 ;
      RECT 98.656 3.891 98.66 4.404 ;
      RECT 98.57 3.887 98.656 4.387 ;
      RECT 98.485 3.879 98.57 4.35 ;
      RECT 98.475 3.875 98.485 4.323 ;
      RECT 98.465 3.875 98.475 4.305 ;
      RECT 98.455 3.877 98.465 4.288 ;
      RECT 98.45 3.882 98.455 4.274 ;
      RECT 98.445 3.886 98.45 4.261 ;
      RECT 98.435 3.891 98.445 4.245 ;
      RECT 98.42 3.905 98.435 4.22 ;
      RECT 98.415 3.911 98.42 4.2 ;
      RECT 98.41 3.913 98.415 4.193 ;
      RECT 98.405 3.917 98.41 4.068 ;
      RECT 98.585 4.717 98.83 5.18 ;
      RECT 98.505 4.69 98.825 5.176 ;
      RECT 98.435 4.725 98.83 5.169 ;
      RECT 98.225 4.98 98.83 5.165 ;
      RECT 98.405 4.748 98.83 5.165 ;
      RECT 98.245 4.94 98.83 5.165 ;
      RECT 98.395 4.76 98.83 5.165 ;
      RECT 98.28 4.877 98.83 5.165 ;
      RECT 98.335 4.802 98.83 5.165 ;
      RECT 98.585 4.667 98.825 5.18 ;
      RECT 98.615 4.66 98.825 5.18 ;
      RECT 98.605 4.662 98.825 5.18 ;
      RECT 98.615 4.657 98.745 5.18 ;
      RECT 98.17 3.22 98.256 3.659 ;
      RECT 98.165 3.22 98.256 3.657 ;
      RECT 98.165 3.22 98.325 3.656 ;
      RECT 98.165 3.22 98.355 3.653 ;
      RECT 98.15 3.227 98.355 3.644 ;
      RECT 98.15 3.227 98.36 3.64 ;
      RECT 98.145 3.237 98.36 3.633 ;
      RECT 98.14 3.242 98.36 3.608 ;
      RECT 98.14 3.242 98.375 3.59 ;
      RECT 98.165 3.22 98.395 3.505 ;
      RECT 98.135 3.247 98.395 3.503 ;
      RECT 98.145 3.24 98.4 3.441 ;
      RECT 98.135 3.362 98.405 3.424 ;
      RECT 98.12 3.257 98.4 3.375 ;
      RECT 98.115 3.267 98.4 3.275 ;
      RECT 98.195 4.038 98.2 4.115 ;
      RECT 98.185 4.032 98.195 4.305 ;
      RECT 98.175 4.024 98.185 4.326 ;
      RECT 98.165 4.015 98.175 4.348 ;
      RECT 98.16 4.01 98.165 4.365 ;
      RECT 98.12 4.01 98.16 4.405 ;
      RECT 98.1 4.01 98.12 4.46 ;
      RECT 98.095 4.01 98.1 4.488 ;
      RECT 98.085 4.01 98.095 4.503 ;
      RECT 98.05 4.01 98.085 4.545 ;
      RECT 98.045 4.01 98.05 4.588 ;
      RECT 98.035 4.01 98.045 4.603 ;
      RECT 98.02 4.01 98.035 4.623 ;
      RECT 98.005 4.01 98.02 4.65 ;
      RECT 98 4.011 98.005 4.668 ;
      RECT 97.98 4.012 98 4.675 ;
      RECT 97.925 4.013 97.98 4.695 ;
      RECT 97.915 4.014 97.925 4.709 ;
      RECT 97.91 4.017 97.915 4.708 ;
      RECT 97.87 4.09 97.91 4.706 ;
      RECT 97.855 4.17 97.87 4.704 ;
      RECT 97.83 4.225 97.855 4.702 ;
      RECT 97.815 4.29 97.83 4.701 ;
      RECT 97.77 4.322 97.815 4.698 ;
      RECT 97.685 4.345 97.77 4.693 ;
      RECT 97.66 4.365 97.685 4.688 ;
      RECT 97.59 4.37 97.66 4.684 ;
      RECT 97.57 4.372 97.59 4.681 ;
      RECT 97.485 4.383 97.57 4.675 ;
      RECT 97.48 4.394 97.485 4.67 ;
      RECT 97.47 4.396 97.48 4.67 ;
      RECT 97.435 4.4 97.47 4.668 ;
      RECT 97.385 4.41 97.435 4.655 ;
      RECT 97.365 4.418 97.385 4.64 ;
      RECT 97.285 4.43 97.365 4.623 ;
      RECT 97.45 3.98 97.62 4.19 ;
      RECT 97.566 3.976 97.62 4.19 ;
      RECT 97.371 3.98 97.62 4.181 ;
      RECT 97.371 3.98 97.625 4.17 ;
      RECT 97.285 3.98 97.625 4.161 ;
      RECT 97.285 3.988 97.635 4.105 ;
      RECT 97.285 4 97.64 4.018 ;
      RECT 97.285 4.007 97.645 4.01 ;
      RECT 97.48 3.978 97.62 4.19 ;
      RECT 97.235 4.923 97.48 5.255 ;
      RECT 97.23 4.915 97.235 5.252 ;
      RECT 97.2 4.935 97.48 5.233 ;
      RECT 97.18 4.967 97.48 5.206 ;
      RECT 97.23 4.92 97.407 5.252 ;
      RECT 97.23 4.917 97.321 5.252 ;
      RECT 97.17 3.265 97.34 3.685 ;
      RECT 97.165 3.265 97.34 3.683 ;
      RECT 97.165 3.265 97.365 3.673 ;
      RECT 97.165 3.265 97.385 3.648 ;
      RECT 97.16 3.265 97.385 3.643 ;
      RECT 97.16 3.265 97.395 3.633 ;
      RECT 97.16 3.265 97.4 3.628 ;
      RECT 97.16 3.27 97.405 3.623 ;
      RECT 97.16 3.302 97.42 3.613 ;
      RECT 97.16 3.372 97.445 3.596 ;
      RECT 97.14 3.372 97.445 3.588 ;
      RECT 97.14 3.432 97.455 3.565 ;
      RECT 97.14 3.472 97.465 3.51 ;
      RECT 97.125 3.265 97.4 3.49 ;
      RECT 97.115 3.28 97.405 3.388 ;
      RECT 96.705 4.67 96.875 5.195 ;
      RECT 96.7 4.67 96.875 5.188 ;
      RECT 96.69 4.67 96.88 5.153 ;
      RECT 96.685 4.68 96.88 5.125 ;
      RECT 96.68 4.7 96.88 5.108 ;
      RECT 96.69 4.675 96.885 5.098 ;
      RECT 96.675 4.72 96.885 5.09 ;
      RECT 96.67 4.74 96.885 5.075 ;
      RECT 96.665 4.77 96.885 5.065 ;
      RECT 96.655 4.815 96.885 5.04 ;
      RECT 96.685 4.685 96.89 5.023 ;
      RECT 96.65 4.867 96.89 5.018 ;
      RECT 96.685 4.695 96.895 4.988 ;
      RECT 96.645 4.9 96.895 4.985 ;
      RECT 96.64 4.925 96.895 4.965 ;
      RECT 96.68 4.712 96.905 4.905 ;
      RECT 96.675 4.734 96.915 4.798 ;
      RECT 96.625 3.981 96.64 4.25 ;
      RECT 96.58 3.965 96.625 4.295 ;
      RECT 96.575 3.953 96.58 4.345 ;
      RECT 96.565 3.949 96.575 4.378 ;
      RECT 96.56 3.946 96.565 4.406 ;
      RECT 96.545 3.948 96.56 4.448 ;
      RECT 96.54 3.952 96.545 4.488 ;
      RECT 96.52 3.957 96.54 4.54 ;
      RECT 96.516 3.962 96.52 4.597 ;
      RECT 96.43 3.981 96.516 4.634 ;
      RECT 96.42 4.002 96.43 4.67 ;
      RECT 96.415 4.01 96.42 4.671 ;
      RECT 96.41 4.052 96.415 4.672 ;
      RECT 96.395 4.14 96.41 4.673 ;
      RECT 96.385 4.29 96.395 4.675 ;
      RECT 96.38 4.335 96.385 4.677 ;
      RECT 96.345 4.377 96.38 4.68 ;
      RECT 96.34 4.395 96.345 4.683 ;
      RECT 96.263 4.401 96.34 4.689 ;
      RECT 96.177 4.415 96.263 4.702 ;
      RECT 96.091 4.429 96.177 4.716 ;
      RECT 96.005 4.443 96.091 4.729 ;
      RECT 95.945 4.455 96.005 4.741 ;
      RECT 95.92 4.462 95.945 4.748 ;
      RECT 95.906 4.465 95.92 4.753 ;
      RECT 95.82 4.473 95.906 4.769 ;
      RECT 95.815 4.48 95.82 4.784 ;
      RECT 95.791 4.48 95.815 4.791 ;
      RECT 95.705 4.483 95.791 4.819 ;
      RECT 95.62 4.487 95.705 4.863 ;
      RECT 95.555 4.491 95.62 4.9 ;
      RECT 95.53 4.494 95.555 4.916 ;
      RECT 95.455 4.507 95.53 4.92 ;
      RECT 95.43 4.525 95.455 4.924 ;
      RECT 95.42 4.532 95.43 4.926 ;
      RECT 95.405 4.535 95.42 4.927 ;
      RECT 95.345 4.547 95.405 4.931 ;
      RECT 95.335 4.561 95.345 4.935 ;
      RECT 95.28 4.571 95.335 4.923 ;
      RECT 95.255 4.592 95.28 4.906 ;
      RECT 95.235 4.612 95.255 4.897 ;
      RECT 95.23 4.625 95.235 4.892 ;
      RECT 95.215 4.637 95.23 4.888 ;
      RECT 96.45 3.292 96.455 3.315 ;
      RECT 96.445 3.283 96.45 3.355 ;
      RECT 96.44 3.281 96.445 3.398 ;
      RECT 96.435 3.272 96.44 3.433 ;
      RECT 96.43 3.262 96.435 3.505 ;
      RECT 96.425 3.252 96.43 3.57 ;
      RECT 96.42 3.249 96.425 3.61 ;
      RECT 96.395 3.243 96.42 3.7 ;
      RECT 96.36 3.231 96.395 3.725 ;
      RECT 96.35 3.222 96.36 3.725 ;
      RECT 96.215 3.22 96.225 3.708 ;
      RECT 96.205 3.22 96.215 3.675 ;
      RECT 96.2 3.22 96.205 3.65 ;
      RECT 96.195 3.22 96.2 3.638 ;
      RECT 96.19 3.22 96.195 3.62 ;
      RECT 96.18 3.22 96.19 3.585 ;
      RECT 96.175 3.222 96.18 3.563 ;
      RECT 96.17 3.228 96.175 3.548 ;
      RECT 96.165 3.234 96.17 3.533 ;
      RECT 96.15 3.246 96.165 3.506 ;
      RECT 96.145 3.257 96.15 3.474 ;
      RECT 96.14 3.267 96.145 3.458 ;
      RECT 96.13 3.275 96.14 3.427 ;
      RECT 96.125 3.285 96.13 3.401 ;
      RECT 96.12 3.342 96.125 3.384 ;
      RECT 96.225 3.22 96.35 3.725 ;
      RECT 95.94 3.907 96.2 4.205 ;
      RECT 95.935 3.914 96.2 4.203 ;
      RECT 95.94 3.909 96.215 4.198 ;
      RECT 95.93 3.922 96.215 4.195 ;
      RECT 95.93 3.927 96.22 4.188 ;
      RECT 95.925 3.935 96.22 4.185 ;
      RECT 95.925 3.952 96.225 3.983 ;
      RECT 95.94 3.904 96.171 4.205 ;
      RECT 95.995 3.903 96.171 4.205 ;
      RECT 95.995 3.9 96.085 4.205 ;
      RECT 95.995 3.897 96.081 4.205 ;
      RECT 95.685 4.17 95.69 4.183 ;
      RECT 95.68 4.137 95.685 4.188 ;
      RECT 95.675 4.092 95.68 4.195 ;
      RECT 95.67 4.047 95.675 4.203 ;
      RECT 95.665 4.015 95.67 4.211 ;
      RECT 95.66 3.975 95.665 4.212 ;
      RECT 95.645 3.955 95.66 4.214 ;
      RECT 95.57 3.937 95.645 4.226 ;
      RECT 95.56 3.93 95.57 4.237 ;
      RECT 95.555 3.93 95.56 4.239 ;
      RECT 95.525 3.936 95.555 4.243 ;
      RECT 95.485 3.949 95.525 4.243 ;
      RECT 95.46 3.96 95.485 4.229 ;
      RECT 95.445 3.966 95.46 4.212 ;
      RECT 95.435 3.968 95.445 4.203 ;
      RECT 95.43 3.969 95.435 4.198 ;
      RECT 95.425 3.97 95.43 4.193 ;
      RECT 95.42 3.971 95.425 4.19 ;
      RECT 95.395 3.976 95.42 4.18 ;
      RECT 95.385 3.992 95.395 4.167 ;
      RECT 95.38 4.012 95.385 4.162 ;
      RECT 95.39 3.405 95.395 3.601 ;
      RECT 95.375 3.369 95.39 3.603 ;
      RECT 95.365 3.351 95.375 3.608 ;
      RECT 95.355 3.337 95.365 3.612 ;
      RECT 95.31 3.321 95.355 3.622 ;
      RECT 95.305 3.311 95.31 3.631 ;
      RECT 95.26 3.3 95.305 3.637 ;
      RECT 95.255 3.288 95.26 3.644 ;
      RECT 95.24 3.283 95.255 3.648 ;
      RECT 95.225 3.275 95.24 3.653 ;
      RECT 95.215 3.268 95.225 3.658 ;
      RECT 95.205 3.265 95.215 3.663 ;
      RECT 95.195 3.265 95.205 3.664 ;
      RECT 95.19 3.262 95.195 3.663 ;
      RECT 95.155 3.257 95.18 3.662 ;
      RECT 95.131 3.253 95.155 3.661 ;
      RECT 95.045 3.244 95.131 3.658 ;
      RECT 95.03 3.236 95.045 3.655 ;
      RECT 95.008 3.235 95.03 3.654 ;
      RECT 94.922 3.235 95.008 3.652 ;
      RECT 94.836 3.235 94.922 3.65 ;
      RECT 94.75 3.235 94.836 3.647 ;
      RECT 94.74 3.235 94.75 3.638 ;
      RECT 94.71 3.235 94.74 3.598 ;
      RECT 94.7 3.245 94.71 3.553 ;
      RECT 94.695 3.285 94.7 3.538 ;
      RECT 94.69 3.3 94.695 3.525 ;
      RECT 94.66 3.38 94.69 3.487 ;
      RECT 95.18 3.26 95.19 3.663 ;
      RECT 95.005 4.025 95.02 4.63 ;
      RECT 95.01 4.02 95.02 4.63 ;
      RECT 95.175 4.02 95.18 4.203 ;
      RECT 95.165 4.02 95.175 4.233 ;
      RECT 95.15 4.02 95.165 4.293 ;
      RECT 95.145 4.02 95.15 4.338 ;
      RECT 95.14 4.02 95.145 4.368 ;
      RECT 95.135 4.02 95.14 4.388 ;
      RECT 95.125 4.02 95.135 4.423 ;
      RECT 95.11 4.02 95.125 4.455 ;
      RECT 95.065 4.02 95.11 4.483 ;
      RECT 95.06 4.02 95.065 4.513 ;
      RECT 95.055 4.02 95.06 4.525 ;
      RECT 95.05 4.02 95.055 4.533 ;
      RECT 95.04 4.02 95.05 4.548 ;
      RECT 95.035 4.02 95.04 4.57 ;
      RECT 95.025 4.02 95.035 4.593 ;
      RECT 95.02 4.02 95.025 4.613 ;
      RECT 94.985 4.035 95.005 4.63 ;
      RECT 94.96 4.052 94.985 4.63 ;
      RECT 94.955 4.062 94.96 4.63 ;
      RECT 94.925 4.077 94.955 4.63 ;
      RECT 94.85 4.119 94.925 4.63 ;
      RECT 94.845 4.15 94.85 4.613 ;
      RECT 94.84 4.154 94.845 4.595 ;
      RECT 94.835 4.158 94.84 4.558 ;
      RECT 94.83 4.342 94.835 4.525 ;
      RECT 94.315 4.531 94.401 5.096 ;
      RECT 94.27 4.533 94.435 5.09 ;
      RECT 94.401 4.53 94.435 5.09 ;
      RECT 94.315 4.532 94.52 5.084 ;
      RECT 94.27 4.542 94.53 5.08 ;
      RECT 94.245 4.534 94.52 5.076 ;
      RECT 94.24 4.537 94.52 5.071 ;
      RECT 94.215 4.552 94.53 5.065 ;
      RECT 94.215 4.577 94.57 5.06 ;
      RECT 94.175 4.585 94.57 5.035 ;
      RECT 94.175 4.612 94.585 5.033 ;
      RECT 94.175 4.642 94.595 5.02 ;
      RECT 94.17 4.787 94.595 5.008 ;
      RECT 94.175 4.716 94.615 5.005 ;
      RECT 94.175 4.773 94.62 4.813 ;
      RECT 94.365 4.052 94.535 4.23 ;
      RECT 94.315 3.991 94.365 4.215 ;
      RECT 94.05 3.971 94.315 4.2 ;
      RECT 94.01 4.035 94.485 4.2 ;
      RECT 94.01 4.025 94.44 4.2 ;
      RECT 94.01 4.022 94.43 4.2 ;
      RECT 94.01 4.01 94.42 4.2 ;
      RECT 94.01 3.995 94.365 4.2 ;
      RECT 94.05 3.967 94.251 4.2 ;
      RECT 94.06 3.945 94.251 4.2 ;
      RECT 94.085 3.93 94.165 4.2 ;
      RECT 93.84 4.46 93.96 4.905 ;
      RECT 93.825 4.46 93.96 4.904 ;
      RECT 93.78 4.482 93.96 4.899 ;
      RECT 93.74 4.531 93.96 4.893 ;
      RECT 93.74 4.531 93.965 4.868 ;
      RECT 93.74 4.531 93.985 4.758 ;
      RECT 93.735 4.561 93.985 4.755 ;
      RECT 93.825 4.46 93.995 4.65 ;
      RECT 93.485 3.245 93.49 3.69 ;
      RECT 93.295 3.245 93.315 3.655 ;
      RECT 93.265 3.245 93.27 3.63 ;
      RECT 93.945 3.552 93.96 3.74 ;
      RECT 93.94 3.537 93.945 3.746 ;
      RECT 93.92 3.51 93.94 3.749 ;
      RECT 93.87 3.477 93.92 3.758 ;
      RECT 93.84 3.457 93.87 3.762 ;
      RECT 93.821 3.445 93.84 3.758 ;
      RECT 93.735 3.417 93.821 3.748 ;
      RECT 93.725 3.392 93.735 3.738 ;
      RECT 93.655 3.36 93.725 3.73 ;
      RECT 93.63 3.32 93.655 3.722 ;
      RECT 93.61 3.302 93.63 3.716 ;
      RECT 93.6 3.292 93.61 3.713 ;
      RECT 93.59 3.285 93.6 3.711 ;
      RECT 93.57 3.272 93.59 3.708 ;
      RECT 93.56 3.262 93.57 3.705 ;
      RECT 93.55 3.255 93.56 3.703 ;
      RECT 93.5 3.247 93.55 3.697 ;
      RECT 93.49 3.245 93.5 3.691 ;
      RECT 93.46 3.245 93.485 3.688 ;
      RECT 93.431 3.245 93.46 3.683 ;
      RECT 93.345 3.245 93.431 3.673 ;
      RECT 93.315 3.245 93.345 3.66 ;
      RECT 93.27 3.245 93.295 3.643 ;
      RECT 93.255 3.245 93.265 3.625 ;
      RECT 93.235 3.252 93.255 3.61 ;
      RECT 93.23 3.267 93.235 3.598 ;
      RECT 93.225 3.272 93.23 3.538 ;
      RECT 93.22 3.277 93.225 3.38 ;
      RECT 93.215 3.28 93.22 3.298 ;
      RECT 92.955 4.57 92.99 4.89 ;
      RECT 93.54 4.755 93.545 4.937 ;
      RECT 93.495 4.637 93.54 4.956 ;
      RECT 93.48 4.614 93.495 4.979 ;
      RECT 93.47 4.604 93.48 4.989 ;
      RECT 93.45 4.599 93.47 5.002 ;
      RECT 93.425 4.597 93.45 5.023 ;
      RECT 93.406 4.596 93.425 5.035 ;
      RECT 93.32 4.593 93.406 5.035 ;
      RECT 93.25 4.588 93.32 5.023 ;
      RECT 93.175 4.584 93.25 4.998 ;
      RECT 93.11 4.58 93.175 4.965 ;
      RECT 93.04 4.577 93.11 4.925 ;
      RECT 93.01 4.573 93.04 4.9 ;
      RECT 92.99 4.571 93.01 4.893 ;
      RECT 92.906 4.569 92.955 4.891 ;
      RECT 92.82 4.566 92.906 4.892 ;
      RECT 92.745 4.565 92.82 4.894 ;
      RECT 92.66 4.565 92.745 4.92 ;
      RECT 92.583 4.566 92.66 4.945 ;
      RECT 92.497 4.567 92.583 4.945 ;
      RECT 92.411 4.567 92.497 4.945 ;
      RECT 92.325 4.568 92.411 4.945 ;
      RECT 92.305 4.569 92.325 4.937 ;
      RECT 92.29 4.575 92.305 4.922 ;
      RECT 92.255 4.595 92.29 4.902 ;
      RECT 92.245 4.615 92.255 4.884 ;
      RECT 93.215 3.92 93.22 4.19 ;
      RECT 93.21 3.911 93.215 4.195 ;
      RECT 93.2 3.901 93.21 4.207 ;
      RECT 93.195 3.89 93.2 4.218 ;
      RECT 93.175 3.884 93.195 4.236 ;
      RECT 93.13 3.881 93.175 4.285 ;
      RECT 93.115 3.88 93.13 4.33 ;
      RECT 93.11 3.88 93.115 4.343 ;
      RECT 93.1 3.88 93.11 4.355 ;
      RECT 93.095 3.881 93.1 4.37 ;
      RECT 93.075 3.889 93.095 4.375 ;
      RECT 93.045 3.905 93.075 4.375 ;
      RECT 93.035 3.917 93.04 4.375 ;
      RECT 93 3.932 93.035 4.375 ;
      RECT 92.97 3.952 93 4.375 ;
      RECT 92.96 3.977 92.97 4.375 ;
      RECT 92.955 4.005 92.96 4.375 ;
      RECT 92.95 4.035 92.955 4.375 ;
      RECT 92.945 4.052 92.95 4.375 ;
      RECT 92.935 4.08 92.945 4.375 ;
      RECT 92.925 4.115 92.935 4.375 ;
      RECT 92.92 4.15 92.925 4.375 ;
      RECT 93.04 3.915 93.045 4.375 ;
      RECT 92.22 3.975 92.74 4.19 ;
      RECT 92.3 3.915 92.74 4.19 ;
      RECT 92.03 3.245 92.035 3.644 ;
      RECT 91.775 3.245 91.81 3.642 ;
      RECT 91.37 3.28 91.375 3.636 ;
      RECT 92.115 3.283 92.12 3.538 ;
      RECT 92.11 3.281 92.115 3.544 ;
      RECT 92.105 3.28 92.11 3.551 ;
      RECT 92.08 3.273 92.105 3.575 ;
      RECT 92.075 3.266 92.08 3.599 ;
      RECT 92.07 3.262 92.075 3.608 ;
      RECT 92.06 3.257 92.07 3.621 ;
      RECT 92.055 3.254 92.06 3.63 ;
      RECT 92.05 3.252 92.055 3.635 ;
      RECT 92.035 3.248 92.05 3.645 ;
      RECT 92.02 3.242 92.03 3.644 ;
      RECT 91.982 3.24 92.02 3.644 ;
      RECT 91.896 3.242 91.982 3.644 ;
      RECT 91.81 3.244 91.896 3.643 ;
      RECT 91.739 3.245 91.775 3.642 ;
      RECT 91.653 3.247 91.739 3.642 ;
      RECT 91.567 3.249 91.653 3.641 ;
      RECT 91.481 3.251 91.567 3.641 ;
      RECT 91.395 3.254 91.481 3.64 ;
      RECT 91.385 3.26 91.395 3.639 ;
      RECT 91.375 3.272 91.385 3.637 ;
      RECT 91.315 3.307 91.37 3.633 ;
      RECT 91.31 3.337 91.315 3.395 ;
      RECT 91.655 4.552 91.66 4.809 ;
      RECT 91.635 4.471 91.655 4.826 ;
      RECT 91.615 4.465 91.635 4.855 ;
      RECT 91.555 4.452 91.615 4.875 ;
      RECT 91.51 4.436 91.555 4.876 ;
      RECT 91.426 4.424 91.51 4.864 ;
      RECT 91.34 4.411 91.426 4.848 ;
      RECT 91.33 4.404 91.34 4.84 ;
      RECT 91.285 4.401 91.33 4.78 ;
      RECT 91.265 4.397 91.285 4.695 ;
      RECT 91.25 4.395 91.265 4.648 ;
      RECT 91.22 4.392 91.25 4.618 ;
      RECT 91.185 4.388 91.22 4.595 ;
      RECT 91.142 4.383 91.185 4.583 ;
      RECT 91.056 4.374 91.142 4.592 ;
      RECT 90.97 4.363 91.056 4.604 ;
      RECT 90.905 4.354 90.97 4.613 ;
      RECT 90.885 4.345 90.905 4.618 ;
      RECT 90.88 4.338 90.885 4.62 ;
      RECT 90.84 4.323 90.88 4.617 ;
      RECT 90.82 4.302 90.84 4.612 ;
      RECT 90.805 4.29 90.82 4.605 ;
      RECT 90.8 4.282 90.805 4.598 ;
      RECT 90.785 4.262 90.8 4.591 ;
      RECT 90.78 4.125 90.785 4.585 ;
      RECT 90.7 4.014 90.78 4.557 ;
      RECT 90.691 4.007 90.7 4.523 ;
      RECT 90.605 4.001 90.691 4.448 ;
      RECT 90.58 3.992 90.605 4.36 ;
      RECT 90.55 3.987 90.58 4.335 ;
      RECT 90.485 3.996 90.55 4.32 ;
      RECT 90.465 4.012 90.485 4.295 ;
      RECT 90.455 4.018 90.465 4.243 ;
      RECT 90.435 4.04 90.455 4.125 ;
      RECT 91.09 4.005 91.26 4.19 ;
      RECT 91.09 4.005 91.295 4.188 ;
      RECT 91.14 3.915 91.31 4.179 ;
      RECT 91.09 4.072 91.315 4.172 ;
      RECT 91.105 3.95 91.31 4.179 ;
      RECT 90.305 4.683 90.37 5.126 ;
      RECT 90.245 4.708 90.37 5.124 ;
      RECT 90.245 4.708 90.425 5.118 ;
      RECT 90.23 4.733 90.425 5.117 ;
      RECT 90.37 4.67 90.445 5.114 ;
      RECT 90.305 4.695 90.525 5.108 ;
      RECT 90.23 4.734 90.57 5.102 ;
      RECT 90.215 4.761 90.57 5.093 ;
      RECT 90.23 4.754 90.59 5.085 ;
      RECT 90.215 4.763 90.595 5.068 ;
      RECT 90.21 4.78 90.595 4.895 ;
      RECT 90.215 3.502 90.25 3.74 ;
      RECT 90.215 3.502 90.28 3.739 ;
      RECT 90.215 3.502 90.395 3.735 ;
      RECT 90.215 3.502 90.45 3.713 ;
      RECT 90.225 3.445 90.505 3.613 ;
      RECT 90.33 3.285 90.36 3.736 ;
      RECT 90.36 3.28 90.54 3.493 ;
      RECT 90.23 3.421 90.54 3.493 ;
      RECT 90.28 3.317 90.33 3.737 ;
      RECT 90.25 3.373 90.54 3.493 ;
      RECT 89.11 7.455 89.28 8.925 ;
      RECT 89.11 7.455 89.285 8.715 ;
      RECT 88.74 9.405 89.21 9.575 ;
      RECT 88.74 8.385 88.91 9.575 ;
      RECT 88.735 3.035 88.905 4.225 ;
      RECT 88.735 3.035 89.205 3.205 ;
      RECT 88.12 3.895 88.295 5.155 ;
      RECT 88.12 3.685 88.29 5.155 ;
      RECT 88.12 7.455 88.29 8.925 ;
      RECT 88.12 7.455 88.295 8.715 ;
      RECT 87.75 3.035 87.92 4.225 ;
      RECT 87.75 3.035 88.22 3.205 ;
      RECT 87.75 9.405 88.22 9.575 ;
      RECT 87.75 8.385 87.92 9.575 ;
      RECT 86.76 4.015 86.935 5.155 ;
      RECT 86.76 1.865 86.93 5.155 ;
      RECT 86.76 1.865 86.935 2.415 ;
      RECT 86.76 10.195 86.935 10.745 ;
      RECT 86.76 7.455 86.93 10.745 ;
      RECT 86.76 7.455 86.935 8.595 ;
      RECT 86.33 3.895 86.505 5.155 ;
      RECT 86.33 2.945 86.5 5.155 ;
      RECT 86.33 7.455 86.5 9.665 ;
      RECT 86.33 7.455 86.505 8.715 ;
      RECT 85.9 3.925 86.07 5.155 ;
      RECT 85.96 2.145 86.13 4.095 ;
      RECT 85.9 1.865 86.07 2.315 ;
      RECT 85.9 10.295 86.07 10.745 ;
      RECT 85.96 8.515 86.13 10.465 ;
      RECT 85.9 7.455 86.07 8.685 ;
      RECT 85.375 3.895 85.55 5.155 ;
      RECT 85.375 1.865 85.545 5.155 ;
      RECT 85.375 3.365 85.785 3.695 ;
      RECT 85.375 2.525 85.785 2.855 ;
      RECT 85.375 1.865 85.55 2.355 ;
      RECT 85.375 10.255 85.55 10.745 ;
      RECT 85.375 7.455 85.545 10.745 ;
      RECT 85.375 9.755 85.785 10.085 ;
      RECT 85.375 8.915 85.785 9.245 ;
      RECT 85.375 7.455 85.55 8.715 ;
      RECT 83.49 4.687 83.505 4.738 ;
      RECT 83.485 4.667 83.49 4.785 ;
      RECT 83.47 4.657 83.485 4.853 ;
      RECT 83.445 4.637 83.47 4.908 ;
      RECT 83.405 4.622 83.445 4.928 ;
      RECT 83.36 4.616 83.405 4.956 ;
      RECT 83.29 4.606 83.36 4.973 ;
      RECT 83.27 4.598 83.29 4.973 ;
      RECT 83.21 4.592 83.27 4.965 ;
      RECT 83.151 4.583 83.21 4.953 ;
      RECT 83.065 4.572 83.151 4.936 ;
      RECT 83.043 4.563 83.065 4.924 ;
      RECT 82.957 4.556 83.043 4.911 ;
      RECT 82.871 4.543 82.957 4.892 ;
      RECT 82.785 4.531 82.871 4.872 ;
      RECT 82.755 4.52 82.785 4.859 ;
      RECT 82.705 4.506 82.755 4.851 ;
      RECT 82.685 4.495 82.705 4.843 ;
      RECT 82.636 4.484 82.685 4.835 ;
      RECT 82.55 4.463 82.636 4.82 ;
      RECT 82.505 4.45 82.55 4.805 ;
      RECT 82.46 4.45 82.505 4.785 ;
      RECT 82.405 4.45 82.46 4.72 ;
      RECT 82.38 4.45 82.405 4.643 ;
      RECT 82.905 4.187 83.075 4.37 ;
      RECT 82.905 4.187 83.09 4.328 ;
      RECT 82.905 4.187 83.095 4.27 ;
      RECT 82.965 3.955 83.1 4.246 ;
      RECT 82.965 3.959 83.105 4.229 ;
      RECT 82.91 4.122 83.105 4.229 ;
      RECT 82.935 3.967 83.075 4.37 ;
      RECT 82.935 3.971 83.115 4.17 ;
      RECT 82.92 4.057 83.115 4.17 ;
      RECT 82.93 3.987 83.075 4.37 ;
      RECT 82.93 3.99 83.125 4.083 ;
      RECT 82.925 4.007 83.125 4.083 ;
      RECT 82.695 3.227 82.865 3.71 ;
      RECT 82.69 3.222 82.84 3.7 ;
      RECT 82.69 3.229 82.87 3.694 ;
      RECT 82.68 3.223 82.84 3.673 ;
      RECT 82.68 3.239 82.885 3.632 ;
      RECT 82.65 3.224 82.84 3.595 ;
      RECT 82.65 3.254 82.895 3.535 ;
      RECT 82.645 3.226 82.84 3.533 ;
      RECT 82.625 3.235 82.87 3.49 ;
      RECT 82.6 3.251 82.885 3.402 ;
      RECT 82.6 3.27 82.91 3.393 ;
      RECT 82.595 3.307 82.91 3.345 ;
      RECT 82.6 3.287 82.915 3.313 ;
      RECT 82.695 3.221 82.805 3.71 ;
      RECT 82.781 3.22 82.805 3.71 ;
      RECT 82.015 4.005 82.02 4.216 ;
      RECT 82.615 4.005 82.62 4.19 ;
      RECT 82.68 4.045 82.685 4.158 ;
      RECT 82.675 4.037 82.68 4.164 ;
      RECT 82.67 4.027 82.675 4.172 ;
      RECT 82.665 4.017 82.67 4.181 ;
      RECT 82.66 4.007 82.665 4.185 ;
      RECT 82.62 4.005 82.66 4.188 ;
      RECT 82.592 4.004 82.615 4.192 ;
      RECT 82.506 4.001 82.592 4.199 ;
      RECT 82.42 3.997 82.506 4.21 ;
      RECT 82.4 3.995 82.42 4.216 ;
      RECT 82.382 3.994 82.4 4.219 ;
      RECT 82.296 3.992 82.382 4.226 ;
      RECT 82.21 3.987 82.296 4.239 ;
      RECT 82.191 3.984 82.21 4.244 ;
      RECT 82.105 3.982 82.191 4.235 ;
      RECT 82.095 3.982 82.105 4.228 ;
      RECT 82.02 3.995 82.095 4.222 ;
      RECT 82.005 4.006 82.015 4.216 ;
      RECT 81.995 4.008 82.005 4.215 ;
      RECT 81.985 4.012 81.995 4.211 ;
      RECT 81.98 4.015 81.985 4.205 ;
      RECT 81.97 4.017 81.98 4.199 ;
      RECT 81.965 4.02 81.97 4.193 ;
      RECT 82 10.195 82.175 10.745 ;
      RECT 82 7.455 82.17 10.745 ;
      RECT 82 7.455 82.175 8.595 ;
      RECT 81.945 4.606 81.95 4.81 ;
      RECT 81.93 4.593 81.945 4.903 ;
      RECT 81.915 4.574 81.93 5.18 ;
      RECT 81.88 4.54 81.915 5.18 ;
      RECT 81.876 4.51 81.88 5.18 ;
      RECT 81.79 4.392 81.876 5.18 ;
      RECT 81.78 4.267 81.79 5.18 ;
      RECT 81.765 4.235 81.78 5.18 ;
      RECT 81.76 4.21 81.765 5.18 ;
      RECT 81.755 4.2 81.76 5.136 ;
      RECT 81.74 4.172 81.755 5.041 ;
      RECT 81.725 4.138 81.74 4.94 ;
      RECT 81.72 4.116 81.725 4.893 ;
      RECT 81.715 4.105 81.72 4.863 ;
      RECT 81.71 4.095 81.715 4.829 ;
      RECT 81.7 4.082 81.71 4.797 ;
      RECT 81.675 4.058 81.7 4.723 ;
      RECT 81.67 4.038 81.675 4.648 ;
      RECT 81.665 4.032 81.67 4.623 ;
      RECT 81.66 4.027 81.665 4.588 ;
      RECT 81.655 4.022 81.66 4.563 ;
      RECT 81.65 4.02 81.655 4.543 ;
      RECT 81.645 4.02 81.65 4.528 ;
      RECT 81.64 4.02 81.645 4.488 ;
      RECT 81.63 4.02 81.64 4.46 ;
      RECT 81.62 4.02 81.63 4.405 ;
      RECT 81.605 4.02 81.62 4.343 ;
      RECT 81.6 4.019 81.605 4.288 ;
      RECT 81.585 4.018 81.6 4.268 ;
      RECT 81.525 4.016 81.585 4.242 ;
      RECT 81.49 4.017 81.525 4.222 ;
      RECT 81.485 4.019 81.49 4.212 ;
      RECT 81.475 4.038 81.485 4.202 ;
      RECT 81.47 4.065 81.475 4.133 ;
      RECT 81.585 3.49 81.755 3.735 ;
      RECT 81.62 3.261 81.755 3.735 ;
      RECT 81.62 3.263 81.765 3.73 ;
      RECT 81.62 3.265 81.79 3.718 ;
      RECT 81.62 3.268 81.815 3.7 ;
      RECT 81.62 3.273 81.865 3.673 ;
      RECT 81.62 3.278 81.885 3.638 ;
      RECT 81.6 3.28 81.895 3.613 ;
      RECT 81.59 3.375 81.895 3.613 ;
      RECT 81.62 3.26 81.73 3.735 ;
      RECT 81.63 3.257 81.725 3.735 ;
      RECT 81.57 7.455 81.74 9.665 ;
      RECT 81.57 7.455 81.745 8.715 ;
      RECT 81.15 4.522 81.34 4.88 ;
      RECT 81.15 4.534 81.375 4.879 ;
      RECT 81.15 4.562 81.395 4.877 ;
      RECT 81.15 4.587 81.4 4.876 ;
      RECT 81.15 4.645 81.415 4.875 ;
      RECT 81.135 4.518 81.295 4.86 ;
      RECT 81.115 4.527 81.34 4.813 ;
      RECT 81.09 4.538 81.375 4.75 ;
      RECT 81.09 4.622 81.41 4.75 ;
      RECT 81.09 4.597 81.405 4.75 ;
      RECT 81.15 4.513 81.295 4.88 ;
      RECT 81.236 4.512 81.295 4.88 ;
      RECT 81.236 4.511 81.28 4.88 ;
      RECT 80.615 10.255 80.79 10.745 ;
      RECT 80.615 7.455 80.785 10.745 ;
      RECT 80.615 9.755 81.025 10.085 ;
      RECT 80.615 8.915 81.025 9.245 ;
      RECT 80.615 7.455 80.79 8.715 ;
      RECT 80.935 4.027 80.94 4.405 ;
      RECT 80.93 3.995 80.935 4.405 ;
      RECT 80.925 3.967 80.93 4.405 ;
      RECT 80.92 3.947 80.925 4.405 ;
      RECT 80.865 3.93 80.92 4.405 ;
      RECT 80.825 3.915 80.865 4.405 ;
      RECT 80.77 3.902 80.825 4.405 ;
      RECT 80.735 3.893 80.77 4.405 ;
      RECT 80.731 3.891 80.735 4.404 ;
      RECT 80.645 3.887 80.731 4.387 ;
      RECT 80.56 3.879 80.645 4.35 ;
      RECT 80.55 3.875 80.56 4.323 ;
      RECT 80.54 3.875 80.55 4.305 ;
      RECT 80.53 3.877 80.54 4.288 ;
      RECT 80.525 3.882 80.53 4.274 ;
      RECT 80.52 3.886 80.525 4.261 ;
      RECT 80.51 3.891 80.52 4.245 ;
      RECT 80.495 3.905 80.51 4.22 ;
      RECT 80.49 3.911 80.495 4.2 ;
      RECT 80.485 3.913 80.49 4.193 ;
      RECT 80.48 3.917 80.485 4.068 ;
      RECT 80.66 4.717 80.905 5.18 ;
      RECT 80.58 4.69 80.9 5.176 ;
      RECT 80.51 4.725 80.905 5.169 ;
      RECT 80.3 4.98 80.905 5.165 ;
      RECT 80.48 4.748 80.905 5.165 ;
      RECT 80.32 4.94 80.905 5.165 ;
      RECT 80.47 4.76 80.905 5.165 ;
      RECT 80.355 4.877 80.905 5.165 ;
      RECT 80.41 4.802 80.905 5.165 ;
      RECT 80.66 4.667 80.9 5.18 ;
      RECT 80.69 4.66 80.9 5.18 ;
      RECT 80.68 4.662 80.9 5.18 ;
      RECT 80.69 4.657 80.82 5.18 ;
      RECT 80.245 3.22 80.331 3.659 ;
      RECT 80.24 3.22 80.331 3.657 ;
      RECT 80.24 3.22 80.4 3.656 ;
      RECT 80.24 3.22 80.43 3.653 ;
      RECT 80.225 3.227 80.43 3.644 ;
      RECT 80.225 3.227 80.435 3.64 ;
      RECT 80.22 3.237 80.435 3.633 ;
      RECT 80.215 3.242 80.435 3.608 ;
      RECT 80.215 3.242 80.45 3.59 ;
      RECT 80.24 3.22 80.47 3.505 ;
      RECT 80.21 3.247 80.47 3.503 ;
      RECT 80.22 3.24 80.475 3.441 ;
      RECT 80.21 3.362 80.48 3.424 ;
      RECT 80.195 3.257 80.475 3.375 ;
      RECT 80.19 3.267 80.475 3.275 ;
      RECT 80.27 4.038 80.275 4.115 ;
      RECT 80.26 4.032 80.27 4.305 ;
      RECT 80.25 4.024 80.26 4.326 ;
      RECT 80.24 4.015 80.25 4.348 ;
      RECT 80.235 4.01 80.24 4.365 ;
      RECT 80.195 4.01 80.235 4.405 ;
      RECT 80.175 4.01 80.195 4.46 ;
      RECT 80.17 4.01 80.175 4.488 ;
      RECT 80.16 4.01 80.17 4.503 ;
      RECT 80.125 4.01 80.16 4.545 ;
      RECT 80.12 4.01 80.125 4.588 ;
      RECT 80.11 4.01 80.12 4.603 ;
      RECT 80.095 4.01 80.11 4.623 ;
      RECT 80.08 4.01 80.095 4.65 ;
      RECT 80.075 4.011 80.08 4.668 ;
      RECT 80.055 4.012 80.075 4.675 ;
      RECT 80 4.013 80.055 4.695 ;
      RECT 79.99 4.014 80 4.709 ;
      RECT 79.985 4.017 79.99 4.708 ;
      RECT 79.945 4.09 79.985 4.706 ;
      RECT 79.93 4.17 79.945 4.704 ;
      RECT 79.905 4.225 79.93 4.702 ;
      RECT 79.89 4.29 79.905 4.701 ;
      RECT 79.845 4.322 79.89 4.698 ;
      RECT 79.76 4.345 79.845 4.693 ;
      RECT 79.735 4.365 79.76 4.688 ;
      RECT 79.665 4.37 79.735 4.684 ;
      RECT 79.645 4.372 79.665 4.681 ;
      RECT 79.56 4.383 79.645 4.675 ;
      RECT 79.555 4.394 79.56 4.67 ;
      RECT 79.545 4.396 79.555 4.67 ;
      RECT 79.51 4.4 79.545 4.668 ;
      RECT 79.46 4.41 79.51 4.655 ;
      RECT 79.44 4.418 79.46 4.64 ;
      RECT 79.36 4.43 79.44 4.623 ;
      RECT 79.525 3.98 79.695 4.19 ;
      RECT 79.641 3.976 79.695 4.19 ;
      RECT 79.446 3.98 79.695 4.181 ;
      RECT 79.446 3.98 79.7 4.17 ;
      RECT 79.36 3.98 79.7 4.161 ;
      RECT 79.36 3.988 79.71 4.105 ;
      RECT 79.36 4 79.715 4.018 ;
      RECT 79.36 4.007 79.72 4.01 ;
      RECT 79.555 3.978 79.695 4.19 ;
      RECT 79.31 4.923 79.555 5.255 ;
      RECT 79.305 4.915 79.31 5.252 ;
      RECT 79.275 4.935 79.555 5.233 ;
      RECT 79.255 4.967 79.555 5.206 ;
      RECT 79.305 4.92 79.482 5.252 ;
      RECT 79.305 4.917 79.396 5.252 ;
      RECT 79.245 3.265 79.415 3.685 ;
      RECT 79.24 3.265 79.415 3.683 ;
      RECT 79.24 3.265 79.44 3.673 ;
      RECT 79.24 3.265 79.46 3.648 ;
      RECT 79.235 3.265 79.46 3.643 ;
      RECT 79.235 3.265 79.47 3.633 ;
      RECT 79.235 3.265 79.475 3.628 ;
      RECT 79.235 3.27 79.48 3.623 ;
      RECT 79.235 3.302 79.495 3.613 ;
      RECT 79.235 3.372 79.52 3.596 ;
      RECT 79.215 3.372 79.52 3.588 ;
      RECT 79.215 3.432 79.53 3.565 ;
      RECT 79.215 3.472 79.54 3.51 ;
      RECT 79.2 3.265 79.475 3.49 ;
      RECT 79.19 3.28 79.48 3.388 ;
      RECT 78.78 4.67 78.95 5.195 ;
      RECT 78.775 4.67 78.95 5.188 ;
      RECT 78.765 4.67 78.955 5.153 ;
      RECT 78.76 4.68 78.955 5.125 ;
      RECT 78.755 4.7 78.955 5.108 ;
      RECT 78.765 4.675 78.96 5.098 ;
      RECT 78.75 4.72 78.96 5.09 ;
      RECT 78.745 4.74 78.96 5.075 ;
      RECT 78.74 4.77 78.96 5.065 ;
      RECT 78.73 4.815 78.96 5.04 ;
      RECT 78.76 4.685 78.965 5.023 ;
      RECT 78.725 4.867 78.965 5.018 ;
      RECT 78.76 4.695 78.97 4.988 ;
      RECT 78.72 4.9 78.97 4.985 ;
      RECT 78.715 4.925 78.97 4.965 ;
      RECT 78.755 4.712 78.98 4.905 ;
      RECT 78.75 4.734 78.99 4.798 ;
      RECT 78.7 3.981 78.715 4.25 ;
      RECT 78.655 3.965 78.7 4.295 ;
      RECT 78.65 3.953 78.655 4.345 ;
      RECT 78.64 3.949 78.65 4.378 ;
      RECT 78.635 3.946 78.64 4.406 ;
      RECT 78.62 3.948 78.635 4.448 ;
      RECT 78.615 3.952 78.62 4.488 ;
      RECT 78.595 3.957 78.615 4.54 ;
      RECT 78.591 3.962 78.595 4.597 ;
      RECT 78.505 3.981 78.591 4.634 ;
      RECT 78.495 4.002 78.505 4.67 ;
      RECT 78.49 4.01 78.495 4.671 ;
      RECT 78.485 4.052 78.49 4.672 ;
      RECT 78.47 4.14 78.485 4.673 ;
      RECT 78.46 4.29 78.47 4.675 ;
      RECT 78.455 4.335 78.46 4.677 ;
      RECT 78.42 4.377 78.455 4.68 ;
      RECT 78.415 4.395 78.42 4.683 ;
      RECT 78.338 4.401 78.415 4.689 ;
      RECT 78.252 4.415 78.338 4.702 ;
      RECT 78.166 4.429 78.252 4.716 ;
      RECT 78.08 4.443 78.166 4.729 ;
      RECT 78.02 4.455 78.08 4.741 ;
      RECT 77.995 4.462 78.02 4.748 ;
      RECT 77.981 4.465 77.995 4.753 ;
      RECT 77.895 4.473 77.981 4.769 ;
      RECT 77.89 4.48 77.895 4.784 ;
      RECT 77.866 4.48 77.89 4.791 ;
      RECT 77.78 4.483 77.866 4.819 ;
      RECT 77.695 4.487 77.78 4.863 ;
      RECT 77.63 4.491 77.695 4.9 ;
      RECT 77.605 4.494 77.63 4.916 ;
      RECT 77.53 4.507 77.605 4.92 ;
      RECT 77.505 4.525 77.53 4.924 ;
      RECT 77.495 4.532 77.505 4.926 ;
      RECT 77.48 4.535 77.495 4.927 ;
      RECT 77.42 4.547 77.48 4.931 ;
      RECT 77.41 4.561 77.42 4.935 ;
      RECT 77.355 4.571 77.41 4.923 ;
      RECT 77.33 4.592 77.355 4.906 ;
      RECT 77.31 4.612 77.33 4.897 ;
      RECT 77.305 4.625 77.31 4.892 ;
      RECT 77.29 4.637 77.305 4.888 ;
      RECT 78.525 3.292 78.53 3.315 ;
      RECT 78.52 3.283 78.525 3.355 ;
      RECT 78.515 3.281 78.52 3.398 ;
      RECT 78.51 3.272 78.515 3.433 ;
      RECT 78.505 3.262 78.51 3.505 ;
      RECT 78.5 3.252 78.505 3.57 ;
      RECT 78.495 3.249 78.5 3.61 ;
      RECT 78.47 3.243 78.495 3.7 ;
      RECT 78.435 3.231 78.47 3.725 ;
      RECT 78.425 3.222 78.435 3.725 ;
      RECT 78.29 3.22 78.3 3.708 ;
      RECT 78.28 3.22 78.29 3.675 ;
      RECT 78.275 3.22 78.28 3.65 ;
      RECT 78.27 3.22 78.275 3.638 ;
      RECT 78.265 3.22 78.27 3.62 ;
      RECT 78.255 3.22 78.265 3.585 ;
      RECT 78.25 3.222 78.255 3.563 ;
      RECT 78.245 3.228 78.25 3.548 ;
      RECT 78.24 3.234 78.245 3.533 ;
      RECT 78.225 3.246 78.24 3.506 ;
      RECT 78.22 3.257 78.225 3.474 ;
      RECT 78.215 3.267 78.22 3.458 ;
      RECT 78.205 3.275 78.215 3.427 ;
      RECT 78.2 3.285 78.205 3.401 ;
      RECT 78.195 3.342 78.2 3.384 ;
      RECT 78.3 3.22 78.425 3.725 ;
      RECT 78.015 3.907 78.275 4.205 ;
      RECT 78.01 3.914 78.275 4.203 ;
      RECT 78.015 3.909 78.29 4.198 ;
      RECT 78.005 3.922 78.29 4.195 ;
      RECT 78.005 3.927 78.295 4.188 ;
      RECT 78 3.935 78.295 4.185 ;
      RECT 78 3.952 78.3 3.983 ;
      RECT 78.015 3.904 78.246 4.205 ;
      RECT 78.07 3.903 78.246 4.205 ;
      RECT 78.07 3.9 78.16 4.205 ;
      RECT 78.07 3.897 78.156 4.205 ;
      RECT 77.76 4.17 77.765 4.183 ;
      RECT 77.755 4.137 77.76 4.188 ;
      RECT 77.75 4.092 77.755 4.195 ;
      RECT 77.745 4.047 77.75 4.203 ;
      RECT 77.74 4.015 77.745 4.211 ;
      RECT 77.735 3.975 77.74 4.212 ;
      RECT 77.72 3.955 77.735 4.214 ;
      RECT 77.645 3.937 77.72 4.226 ;
      RECT 77.635 3.93 77.645 4.237 ;
      RECT 77.63 3.93 77.635 4.239 ;
      RECT 77.6 3.936 77.63 4.243 ;
      RECT 77.56 3.949 77.6 4.243 ;
      RECT 77.535 3.96 77.56 4.229 ;
      RECT 77.52 3.966 77.535 4.212 ;
      RECT 77.51 3.968 77.52 4.203 ;
      RECT 77.505 3.969 77.51 4.198 ;
      RECT 77.5 3.97 77.505 4.193 ;
      RECT 77.495 3.971 77.5 4.19 ;
      RECT 77.47 3.976 77.495 4.18 ;
      RECT 77.46 3.992 77.47 4.167 ;
      RECT 77.455 4.012 77.46 4.162 ;
      RECT 77.465 3.405 77.47 3.601 ;
      RECT 77.45 3.369 77.465 3.603 ;
      RECT 77.44 3.351 77.45 3.608 ;
      RECT 77.43 3.337 77.44 3.612 ;
      RECT 77.385 3.321 77.43 3.622 ;
      RECT 77.38 3.311 77.385 3.631 ;
      RECT 77.335 3.3 77.38 3.637 ;
      RECT 77.33 3.288 77.335 3.644 ;
      RECT 77.315 3.283 77.33 3.648 ;
      RECT 77.3 3.275 77.315 3.653 ;
      RECT 77.29 3.268 77.3 3.658 ;
      RECT 77.28 3.265 77.29 3.663 ;
      RECT 77.27 3.265 77.28 3.664 ;
      RECT 77.265 3.262 77.27 3.663 ;
      RECT 77.23 3.257 77.255 3.662 ;
      RECT 77.206 3.253 77.23 3.661 ;
      RECT 77.12 3.244 77.206 3.658 ;
      RECT 77.105 3.236 77.12 3.655 ;
      RECT 77.083 3.235 77.105 3.654 ;
      RECT 76.997 3.235 77.083 3.652 ;
      RECT 76.911 3.235 76.997 3.65 ;
      RECT 76.825 3.235 76.911 3.647 ;
      RECT 76.815 3.235 76.825 3.638 ;
      RECT 76.785 3.235 76.815 3.598 ;
      RECT 76.775 3.245 76.785 3.553 ;
      RECT 76.77 3.285 76.775 3.538 ;
      RECT 76.765 3.3 76.77 3.525 ;
      RECT 76.735 3.38 76.765 3.487 ;
      RECT 77.255 3.26 77.265 3.663 ;
      RECT 77.08 4.025 77.095 4.63 ;
      RECT 77.085 4.02 77.095 4.63 ;
      RECT 77.25 4.02 77.255 4.203 ;
      RECT 77.24 4.02 77.25 4.233 ;
      RECT 77.225 4.02 77.24 4.293 ;
      RECT 77.22 4.02 77.225 4.338 ;
      RECT 77.215 4.02 77.22 4.368 ;
      RECT 77.21 4.02 77.215 4.388 ;
      RECT 77.2 4.02 77.21 4.423 ;
      RECT 77.185 4.02 77.2 4.455 ;
      RECT 77.14 4.02 77.185 4.483 ;
      RECT 77.135 4.02 77.14 4.513 ;
      RECT 77.13 4.02 77.135 4.525 ;
      RECT 77.125 4.02 77.13 4.533 ;
      RECT 77.115 4.02 77.125 4.548 ;
      RECT 77.11 4.02 77.115 4.57 ;
      RECT 77.1 4.02 77.11 4.593 ;
      RECT 77.095 4.02 77.1 4.613 ;
      RECT 77.06 4.035 77.08 4.63 ;
      RECT 77.035 4.052 77.06 4.63 ;
      RECT 77.03 4.062 77.035 4.63 ;
      RECT 77 4.077 77.03 4.63 ;
      RECT 76.925 4.119 77 4.63 ;
      RECT 76.92 4.15 76.925 4.613 ;
      RECT 76.915 4.154 76.92 4.595 ;
      RECT 76.91 4.158 76.915 4.558 ;
      RECT 76.905 4.342 76.91 4.525 ;
      RECT 76.39 4.531 76.476 5.096 ;
      RECT 76.345 4.533 76.51 5.09 ;
      RECT 76.476 4.53 76.51 5.09 ;
      RECT 76.39 4.532 76.595 5.084 ;
      RECT 76.345 4.542 76.605 5.08 ;
      RECT 76.32 4.534 76.595 5.076 ;
      RECT 76.315 4.537 76.595 5.071 ;
      RECT 76.29 4.552 76.605 5.065 ;
      RECT 76.29 4.577 76.645 5.06 ;
      RECT 76.25 4.585 76.645 5.035 ;
      RECT 76.25 4.612 76.66 5.033 ;
      RECT 76.25 4.642 76.67 5.02 ;
      RECT 76.245 4.787 76.67 5.008 ;
      RECT 76.25 4.716 76.69 5.005 ;
      RECT 76.25 4.773 76.695 4.813 ;
      RECT 76.44 4.052 76.61 4.23 ;
      RECT 76.39 3.991 76.44 4.215 ;
      RECT 76.125 3.971 76.39 4.2 ;
      RECT 76.085 4.035 76.56 4.2 ;
      RECT 76.085 4.025 76.515 4.2 ;
      RECT 76.085 4.022 76.505 4.2 ;
      RECT 76.085 4.01 76.495 4.2 ;
      RECT 76.085 3.995 76.44 4.2 ;
      RECT 76.125 3.967 76.326 4.2 ;
      RECT 76.135 3.945 76.326 4.2 ;
      RECT 76.16 3.93 76.24 4.2 ;
      RECT 75.915 4.46 76.035 4.905 ;
      RECT 75.9 4.46 76.035 4.904 ;
      RECT 75.855 4.482 76.035 4.899 ;
      RECT 75.815 4.531 76.035 4.893 ;
      RECT 75.815 4.531 76.04 4.868 ;
      RECT 75.815 4.531 76.06 4.758 ;
      RECT 75.81 4.561 76.06 4.755 ;
      RECT 75.9 4.46 76.07 4.65 ;
      RECT 75.56 3.245 75.565 3.69 ;
      RECT 75.37 3.245 75.39 3.655 ;
      RECT 75.34 3.245 75.345 3.63 ;
      RECT 76.02 3.552 76.035 3.74 ;
      RECT 76.015 3.537 76.02 3.746 ;
      RECT 75.995 3.51 76.015 3.749 ;
      RECT 75.945 3.477 75.995 3.758 ;
      RECT 75.915 3.457 75.945 3.762 ;
      RECT 75.896 3.445 75.915 3.758 ;
      RECT 75.81 3.417 75.896 3.748 ;
      RECT 75.8 3.392 75.81 3.738 ;
      RECT 75.73 3.36 75.8 3.73 ;
      RECT 75.705 3.32 75.73 3.722 ;
      RECT 75.685 3.302 75.705 3.716 ;
      RECT 75.675 3.292 75.685 3.713 ;
      RECT 75.665 3.285 75.675 3.711 ;
      RECT 75.645 3.272 75.665 3.708 ;
      RECT 75.635 3.262 75.645 3.705 ;
      RECT 75.625 3.255 75.635 3.703 ;
      RECT 75.575 3.247 75.625 3.697 ;
      RECT 75.565 3.245 75.575 3.691 ;
      RECT 75.535 3.245 75.56 3.688 ;
      RECT 75.506 3.245 75.535 3.683 ;
      RECT 75.42 3.245 75.506 3.673 ;
      RECT 75.39 3.245 75.42 3.66 ;
      RECT 75.345 3.245 75.37 3.643 ;
      RECT 75.33 3.245 75.34 3.625 ;
      RECT 75.31 3.252 75.33 3.61 ;
      RECT 75.305 3.267 75.31 3.598 ;
      RECT 75.3 3.272 75.305 3.538 ;
      RECT 75.295 3.277 75.3 3.38 ;
      RECT 75.29 3.28 75.295 3.298 ;
      RECT 75.03 4.57 75.065 4.89 ;
      RECT 75.615 4.755 75.62 4.937 ;
      RECT 75.57 4.637 75.615 4.956 ;
      RECT 75.555 4.614 75.57 4.979 ;
      RECT 75.545 4.604 75.555 4.989 ;
      RECT 75.525 4.599 75.545 5.002 ;
      RECT 75.5 4.597 75.525 5.023 ;
      RECT 75.481 4.596 75.5 5.035 ;
      RECT 75.395 4.593 75.481 5.035 ;
      RECT 75.325 4.588 75.395 5.023 ;
      RECT 75.25 4.584 75.325 4.998 ;
      RECT 75.185 4.58 75.25 4.965 ;
      RECT 75.115 4.577 75.185 4.925 ;
      RECT 75.085 4.573 75.115 4.9 ;
      RECT 75.065 4.571 75.085 4.893 ;
      RECT 74.981 4.569 75.03 4.891 ;
      RECT 74.895 4.566 74.981 4.892 ;
      RECT 74.82 4.565 74.895 4.894 ;
      RECT 74.735 4.565 74.82 4.92 ;
      RECT 74.658 4.566 74.735 4.945 ;
      RECT 74.572 4.567 74.658 4.945 ;
      RECT 74.486 4.567 74.572 4.945 ;
      RECT 74.4 4.568 74.486 4.945 ;
      RECT 74.38 4.569 74.4 4.937 ;
      RECT 74.365 4.575 74.38 4.922 ;
      RECT 74.33 4.595 74.365 4.902 ;
      RECT 74.32 4.615 74.33 4.884 ;
      RECT 75.29 3.92 75.295 4.19 ;
      RECT 75.285 3.911 75.29 4.195 ;
      RECT 75.275 3.901 75.285 4.207 ;
      RECT 75.27 3.89 75.275 4.218 ;
      RECT 75.25 3.884 75.27 4.236 ;
      RECT 75.205 3.881 75.25 4.285 ;
      RECT 75.19 3.88 75.205 4.33 ;
      RECT 75.185 3.88 75.19 4.343 ;
      RECT 75.175 3.88 75.185 4.355 ;
      RECT 75.17 3.881 75.175 4.37 ;
      RECT 75.15 3.889 75.17 4.375 ;
      RECT 75.12 3.905 75.15 4.375 ;
      RECT 75.11 3.917 75.115 4.375 ;
      RECT 75.075 3.932 75.11 4.375 ;
      RECT 75.045 3.952 75.075 4.375 ;
      RECT 75.035 3.977 75.045 4.375 ;
      RECT 75.03 4.005 75.035 4.375 ;
      RECT 75.025 4.035 75.03 4.375 ;
      RECT 75.02 4.052 75.025 4.375 ;
      RECT 75.01 4.08 75.02 4.375 ;
      RECT 75 4.115 75.01 4.375 ;
      RECT 74.995 4.15 75 4.375 ;
      RECT 75.115 3.915 75.12 4.375 ;
      RECT 74.295 3.975 74.815 4.19 ;
      RECT 74.375 3.915 74.815 4.19 ;
      RECT 74.105 3.245 74.11 3.644 ;
      RECT 73.85 3.245 73.885 3.642 ;
      RECT 73.445 3.28 73.45 3.636 ;
      RECT 74.19 3.283 74.195 3.538 ;
      RECT 74.185 3.281 74.19 3.544 ;
      RECT 74.18 3.28 74.185 3.551 ;
      RECT 74.155 3.273 74.18 3.575 ;
      RECT 74.15 3.266 74.155 3.599 ;
      RECT 74.145 3.262 74.15 3.608 ;
      RECT 74.135 3.257 74.145 3.621 ;
      RECT 74.13 3.254 74.135 3.63 ;
      RECT 74.125 3.252 74.13 3.635 ;
      RECT 74.11 3.248 74.125 3.645 ;
      RECT 74.095 3.242 74.105 3.644 ;
      RECT 74.057 3.24 74.095 3.644 ;
      RECT 73.971 3.242 74.057 3.644 ;
      RECT 73.885 3.244 73.971 3.643 ;
      RECT 73.814 3.245 73.85 3.642 ;
      RECT 73.728 3.247 73.814 3.642 ;
      RECT 73.642 3.249 73.728 3.641 ;
      RECT 73.556 3.251 73.642 3.641 ;
      RECT 73.47 3.254 73.556 3.64 ;
      RECT 73.46 3.26 73.47 3.639 ;
      RECT 73.45 3.272 73.46 3.637 ;
      RECT 73.39 3.307 73.445 3.633 ;
      RECT 73.385 3.337 73.39 3.395 ;
      RECT 73.73 4.552 73.735 4.809 ;
      RECT 73.71 4.471 73.73 4.826 ;
      RECT 73.69 4.465 73.71 4.855 ;
      RECT 73.63 4.452 73.69 4.875 ;
      RECT 73.585 4.436 73.63 4.876 ;
      RECT 73.501 4.424 73.585 4.864 ;
      RECT 73.415 4.411 73.501 4.848 ;
      RECT 73.405 4.404 73.415 4.84 ;
      RECT 73.36 4.401 73.405 4.78 ;
      RECT 73.34 4.397 73.36 4.695 ;
      RECT 73.325 4.395 73.34 4.648 ;
      RECT 73.295 4.392 73.325 4.618 ;
      RECT 73.26 4.388 73.295 4.595 ;
      RECT 73.217 4.383 73.26 4.583 ;
      RECT 73.131 4.374 73.217 4.592 ;
      RECT 73.045 4.363 73.131 4.604 ;
      RECT 72.98 4.354 73.045 4.613 ;
      RECT 72.96 4.345 72.98 4.618 ;
      RECT 72.955 4.338 72.96 4.62 ;
      RECT 72.915 4.323 72.955 4.617 ;
      RECT 72.895 4.302 72.915 4.612 ;
      RECT 72.88 4.29 72.895 4.605 ;
      RECT 72.875 4.282 72.88 4.598 ;
      RECT 72.86 4.262 72.875 4.591 ;
      RECT 72.855 4.125 72.86 4.585 ;
      RECT 72.775 4.014 72.855 4.557 ;
      RECT 72.766 4.007 72.775 4.523 ;
      RECT 72.68 4.001 72.766 4.448 ;
      RECT 72.655 3.992 72.68 4.36 ;
      RECT 72.625 3.987 72.655 4.335 ;
      RECT 72.56 3.996 72.625 4.32 ;
      RECT 72.54 4.012 72.56 4.295 ;
      RECT 72.53 4.018 72.54 4.243 ;
      RECT 72.51 4.04 72.53 4.125 ;
      RECT 73.165 4.005 73.335 4.19 ;
      RECT 73.165 4.005 73.37 4.188 ;
      RECT 73.215 3.915 73.385 4.179 ;
      RECT 73.165 4.072 73.39 4.172 ;
      RECT 73.18 3.95 73.385 4.179 ;
      RECT 72.38 4.683 72.445 5.126 ;
      RECT 72.32 4.708 72.445 5.124 ;
      RECT 72.32 4.708 72.5 5.118 ;
      RECT 72.305 4.733 72.5 5.117 ;
      RECT 72.445 4.67 72.52 5.114 ;
      RECT 72.38 4.695 72.6 5.108 ;
      RECT 72.305 4.734 72.645 5.102 ;
      RECT 72.29 4.761 72.645 5.093 ;
      RECT 72.305 4.754 72.665 5.085 ;
      RECT 72.29 4.763 72.67 5.068 ;
      RECT 72.285 4.78 72.67 4.895 ;
      RECT 72.29 3.502 72.325 3.74 ;
      RECT 72.29 3.502 72.355 3.739 ;
      RECT 72.29 3.502 72.47 3.735 ;
      RECT 72.29 3.502 72.525 3.713 ;
      RECT 72.3 3.445 72.58 3.613 ;
      RECT 72.405 3.285 72.435 3.736 ;
      RECT 72.435 3.28 72.615 3.493 ;
      RECT 72.305 3.421 72.615 3.493 ;
      RECT 72.355 3.317 72.405 3.737 ;
      RECT 72.325 3.373 72.615 3.493 ;
      RECT 71.185 7.455 71.355 8.925 ;
      RECT 71.185 7.455 71.36 8.715 ;
      RECT 70.815 9.405 71.285 9.575 ;
      RECT 70.815 8.385 70.985 9.575 ;
      RECT 70.81 3.035 70.98 4.225 ;
      RECT 70.81 3.035 71.28 3.205 ;
      RECT 70.195 3.895 70.37 5.155 ;
      RECT 70.195 3.685 70.365 5.155 ;
      RECT 70.195 7.455 70.365 8.925 ;
      RECT 70.195 7.455 70.37 8.715 ;
      RECT 69.825 3.035 69.995 4.225 ;
      RECT 69.825 3.035 70.295 3.205 ;
      RECT 69.825 9.405 70.295 9.575 ;
      RECT 69.825 8.385 69.995 9.575 ;
      RECT 68.835 4.015 69.01 5.155 ;
      RECT 68.835 1.865 69.005 5.155 ;
      RECT 68.835 1.865 69.01 2.415 ;
      RECT 68.835 10.195 69.01 10.745 ;
      RECT 68.835 7.455 69.005 10.745 ;
      RECT 68.835 7.455 69.01 8.595 ;
      RECT 68.405 3.895 68.58 5.155 ;
      RECT 68.405 2.945 68.575 5.155 ;
      RECT 68.405 7.455 68.575 9.665 ;
      RECT 68.405 7.455 68.58 8.715 ;
      RECT 67.975 3.925 68.145 5.155 ;
      RECT 68.035 2.145 68.205 4.095 ;
      RECT 67.975 1.865 68.145 2.315 ;
      RECT 67.975 10.295 68.145 10.745 ;
      RECT 68.035 8.515 68.205 10.465 ;
      RECT 67.975 7.455 68.145 8.685 ;
      RECT 67.45 3.895 67.625 5.155 ;
      RECT 67.45 1.865 67.62 5.155 ;
      RECT 67.45 3.365 67.86 3.695 ;
      RECT 67.45 2.525 67.86 2.855 ;
      RECT 67.45 1.865 67.625 2.355 ;
      RECT 67.45 10.255 67.625 10.745 ;
      RECT 67.45 7.455 67.62 10.745 ;
      RECT 67.45 9.755 67.86 10.085 ;
      RECT 67.45 8.915 67.86 9.245 ;
      RECT 67.45 7.455 67.625 8.715 ;
      RECT 65.565 4.687 65.58 4.738 ;
      RECT 65.56 4.667 65.565 4.785 ;
      RECT 65.545 4.657 65.56 4.853 ;
      RECT 65.52 4.637 65.545 4.908 ;
      RECT 65.48 4.622 65.52 4.928 ;
      RECT 65.435 4.616 65.48 4.956 ;
      RECT 65.365 4.606 65.435 4.973 ;
      RECT 65.345 4.598 65.365 4.973 ;
      RECT 65.285 4.592 65.345 4.965 ;
      RECT 65.226 4.583 65.285 4.953 ;
      RECT 65.14 4.572 65.226 4.936 ;
      RECT 65.118 4.563 65.14 4.924 ;
      RECT 65.032 4.556 65.118 4.911 ;
      RECT 64.946 4.543 65.032 4.892 ;
      RECT 64.86 4.531 64.946 4.872 ;
      RECT 64.83 4.52 64.86 4.859 ;
      RECT 64.78 4.506 64.83 4.851 ;
      RECT 64.76 4.495 64.78 4.843 ;
      RECT 64.711 4.484 64.76 4.835 ;
      RECT 64.625 4.463 64.711 4.82 ;
      RECT 64.58 4.45 64.625 4.805 ;
      RECT 64.535 4.45 64.58 4.785 ;
      RECT 64.48 4.45 64.535 4.72 ;
      RECT 64.455 4.45 64.48 4.643 ;
      RECT 64.98 4.187 65.15 4.37 ;
      RECT 64.98 4.187 65.165 4.328 ;
      RECT 64.98 4.187 65.17 4.27 ;
      RECT 65.04 3.955 65.175 4.246 ;
      RECT 65.04 3.959 65.18 4.229 ;
      RECT 64.985 4.122 65.18 4.229 ;
      RECT 65.01 3.967 65.15 4.37 ;
      RECT 65.01 3.971 65.19 4.17 ;
      RECT 64.995 4.057 65.19 4.17 ;
      RECT 65.005 3.987 65.15 4.37 ;
      RECT 65.005 3.99 65.2 4.083 ;
      RECT 65 4.007 65.2 4.083 ;
      RECT 64.77 3.227 64.94 3.71 ;
      RECT 64.765 3.222 64.915 3.7 ;
      RECT 64.765 3.229 64.945 3.694 ;
      RECT 64.755 3.223 64.915 3.673 ;
      RECT 64.755 3.239 64.96 3.632 ;
      RECT 64.725 3.224 64.915 3.595 ;
      RECT 64.725 3.254 64.97 3.535 ;
      RECT 64.72 3.226 64.915 3.533 ;
      RECT 64.7 3.235 64.945 3.49 ;
      RECT 64.675 3.251 64.96 3.402 ;
      RECT 64.675 3.27 64.985 3.393 ;
      RECT 64.67 3.307 64.985 3.345 ;
      RECT 64.675 3.287 64.99 3.313 ;
      RECT 64.77 3.221 64.88 3.71 ;
      RECT 64.856 3.22 64.88 3.71 ;
      RECT 64.09 4.005 64.095 4.216 ;
      RECT 64.69 4.005 64.695 4.19 ;
      RECT 64.755 4.045 64.76 4.158 ;
      RECT 64.75 4.037 64.755 4.164 ;
      RECT 64.745 4.027 64.75 4.172 ;
      RECT 64.74 4.017 64.745 4.181 ;
      RECT 64.735 4.007 64.74 4.185 ;
      RECT 64.695 4.005 64.735 4.188 ;
      RECT 64.667 4.004 64.69 4.192 ;
      RECT 64.581 4.001 64.667 4.199 ;
      RECT 64.495 3.997 64.581 4.21 ;
      RECT 64.475 3.995 64.495 4.216 ;
      RECT 64.457 3.994 64.475 4.219 ;
      RECT 64.371 3.992 64.457 4.226 ;
      RECT 64.285 3.987 64.371 4.239 ;
      RECT 64.266 3.984 64.285 4.244 ;
      RECT 64.18 3.982 64.266 4.235 ;
      RECT 64.17 3.982 64.18 4.228 ;
      RECT 64.095 3.995 64.17 4.222 ;
      RECT 64.08 4.006 64.09 4.216 ;
      RECT 64.07 4.008 64.08 4.215 ;
      RECT 64.06 4.012 64.07 4.211 ;
      RECT 64.055 4.015 64.06 4.205 ;
      RECT 64.045 4.017 64.055 4.199 ;
      RECT 64.04 4.02 64.045 4.193 ;
      RECT 64.075 10.195 64.25 10.745 ;
      RECT 64.075 7.455 64.245 10.745 ;
      RECT 64.075 7.455 64.25 8.595 ;
      RECT 64.02 4.606 64.025 4.81 ;
      RECT 64.005 4.593 64.02 4.903 ;
      RECT 63.99 4.574 64.005 5.18 ;
      RECT 63.955 4.54 63.99 5.18 ;
      RECT 63.951 4.51 63.955 5.18 ;
      RECT 63.865 4.392 63.951 5.18 ;
      RECT 63.855 4.267 63.865 5.18 ;
      RECT 63.84 4.235 63.855 5.18 ;
      RECT 63.835 4.21 63.84 5.18 ;
      RECT 63.83 4.2 63.835 5.136 ;
      RECT 63.815 4.172 63.83 5.041 ;
      RECT 63.8 4.138 63.815 4.94 ;
      RECT 63.795 4.116 63.8 4.893 ;
      RECT 63.79 4.105 63.795 4.863 ;
      RECT 63.785 4.095 63.79 4.829 ;
      RECT 63.775 4.082 63.785 4.797 ;
      RECT 63.75 4.058 63.775 4.723 ;
      RECT 63.745 4.038 63.75 4.648 ;
      RECT 63.74 4.032 63.745 4.623 ;
      RECT 63.735 4.027 63.74 4.588 ;
      RECT 63.73 4.022 63.735 4.563 ;
      RECT 63.725 4.02 63.73 4.543 ;
      RECT 63.72 4.02 63.725 4.528 ;
      RECT 63.715 4.02 63.72 4.488 ;
      RECT 63.705 4.02 63.715 4.46 ;
      RECT 63.695 4.02 63.705 4.405 ;
      RECT 63.68 4.02 63.695 4.343 ;
      RECT 63.675 4.019 63.68 4.288 ;
      RECT 63.66 4.018 63.675 4.268 ;
      RECT 63.6 4.016 63.66 4.242 ;
      RECT 63.565 4.017 63.6 4.222 ;
      RECT 63.56 4.019 63.565 4.212 ;
      RECT 63.55 4.038 63.56 4.202 ;
      RECT 63.545 4.065 63.55 4.133 ;
      RECT 63.66 3.49 63.83 3.735 ;
      RECT 63.695 3.261 63.83 3.735 ;
      RECT 63.695 3.263 63.84 3.73 ;
      RECT 63.695 3.265 63.865 3.718 ;
      RECT 63.695 3.268 63.89 3.7 ;
      RECT 63.695 3.273 63.94 3.673 ;
      RECT 63.695 3.278 63.96 3.638 ;
      RECT 63.675 3.28 63.97 3.613 ;
      RECT 63.665 3.375 63.97 3.613 ;
      RECT 63.695 3.26 63.805 3.735 ;
      RECT 63.705 3.257 63.8 3.735 ;
      RECT 63.645 7.455 63.815 9.665 ;
      RECT 63.645 7.455 63.82 8.715 ;
      RECT 63.225 4.522 63.415 4.88 ;
      RECT 63.225 4.534 63.45 4.879 ;
      RECT 63.225 4.562 63.47 4.877 ;
      RECT 63.225 4.587 63.475 4.876 ;
      RECT 63.225 4.645 63.49 4.875 ;
      RECT 63.21 4.518 63.37 4.86 ;
      RECT 63.19 4.527 63.415 4.813 ;
      RECT 63.165 4.538 63.45 4.75 ;
      RECT 63.165 4.622 63.485 4.75 ;
      RECT 63.165 4.597 63.48 4.75 ;
      RECT 63.225 4.513 63.37 4.88 ;
      RECT 63.311 4.512 63.37 4.88 ;
      RECT 63.311 4.511 63.355 4.88 ;
      RECT 62.69 10.255 62.865 10.745 ;
      RECT 62.69 7.455 62.86 10.745 ;
      RECT 62.69 9.755 63.1 10.085 ;
      RECT 62.69 8.915 63.1 9.245 ;
      RECT 62.69 7.455 62.865 8.715 ;
      RECT 63.01 4.027 63.015 4.405 ;
      RECT 63.005 3.995 63.01 4.405 ;
      RECT 63 3.967 63.005 4.405 ;
      RECT 62.995 3.947 63 4.405 ;
      RECT 62.94 3.93 62.995 4.405 ;
      RECT 62.9 3.915 62.94 4.405 ;
      RECT 62.845 3.902 62.9 4.405 ;
      RECT 62.81 3.893 62.845 4.405 ;
      RECT 62.806 3.891 62.81 4.404 ;
      RECT 62.72 3.887 62.806 4.387 ;
      RECT 62.635 3.879 62.72 4.35 ;
      RECT 62.625 3.875 62.635 4.323 ;
      RECT 62.615 3.875 62.625 4.305 ;
      RECT 62.605 3.877 62.615 4.288 ;
      RECT 62.6 3.882 62.605 4.274 ;
      RECT 62.595 3.886 62.6 4.261 ;
      RECT 62.585 3.891 62.595 4.245 ;
      RECT 62.57 3.905 62.585 4.22 ;
      RECT 62.565 3.911 62.57 4.2 ;
      RECT 62.56 3.913 62.565 4.193 ;
      RECT 62.555 3.917 62.56 4.068 ;
      RECT 62.735 4.717 62.98 5.18 ;
      RECT 62.655 4.69 62.975 5.176 ;
      RECT 62.585 4.725 62.98 5.169 ;
      RECT 62.375 4.98 62.98 5.165 ;
      RECT 62.555 4.748 62.98 5.165 ;
      RECT 62.395 4.94 62.98 5.165 ;
      RECT 62.545 4.76 62.98 5.165 ;
      RECT 62.43 4.877 62.98 5.165 ;
      RECT 62.485 4.802 62.98 5.165 ;
      RECT 62.735 4.667 62.975 5.18 ;
      RECT 62.765 4.66 62.975 5.18 ;
      RECT 62.755 4.662 62.975 5.18 ;
      RECT 62.765 4.657 62.895 5.18 ;
      RECT 62.32 3.22 62.406 3.659 ;
      RECT 62.315 3.22 62.406 3.657 ;
      RECT 62.315 3.22 62.475 3.656 ;
      RECT 62.315 3.22 62.505 3.653 ;
      RECT 62.3 3.227 62.505 3.644 ;
      RECT 62.3 3.227 62.51 3.64 ;
      RECT 62.295 3.237 62.51 3.633 ;
      RECT 62.29 3.242 62.51 3.608 ;
      RECT 62.29 3.242 62.525 3.59 ;
      RECT 62.315 3.22 62.545 3.505 ;
      RECT 62.285 3.247 62.545 3.503 ;
      RECT 62.295 3.24 62.55 3.441 ;
      RECT 62.285 3.362 62.555 3.424 ;
      RECT 62.27 3.257 62.55 3.375 ;
      RECT 62.265 3.267 62.55 3.275 ;
      RECT 62.345 4.038 62.35 4.115 ;
      RECT 62.335 4.032 62.345 4.305 ;
      RECT 62.325 4.024 62.335 4.326 ;
      RECT 62.315 4.015 62.325 4.348 ;
      RECT 62.31 4.01 62.315 4.365 ;
      RECT 62.27 4.01 62.31 4.405 ;
      RECT 62.25 4.01 62.27 4.46 ;
      RECT 62.245 4.01 62.25 4.488 ;
      RECT 62.235 4.01 62.245 4.503 ;
      RECT 62.2 4.01 62.235 4.545 ;
      RECT 62.195 4.01 62.2 4.588 ;
      RECT 62.185 4.01 62.195 4.603 ;
      RECT 62.17 4.01 62.185 4.623 ;
      RECT 62.155 4.01 62.17 4.65 ;
      RECT 62.15 4.011 62.155 4.668 ;
      RECT 62.13 4.012 62.15 4.675 ;
      RECT 62.075 4.013 62.13 4.695 ;
      RECT 62.065 4.014 62.075 4.709 ;
      RECT 62.06 4.017 62.065 4.708 ;
      RECT 62.02 4.09 62.06 4.706 ;
      RECT 62.005 4.17 62.02 4.704 ;
      RECT 61.98 4.225 62.005 4.702 ;
      RECT 61.965 4.29 61.98 4.701 ;
      RECT 61.92 4.322 61.965 4.698 ;
      RECT 61.835 4.345 61.92 4.693 ;
      RECT 61.81 4.365 61.835 4.688 ;
      RECT 61.74 4.37 61.81 4.684 ;
      RECT 61.72 4.372 61.74 4.681 ;
      RECT 61.635 4.383 61.72 4.675 ;
      RECT 61.63 4.394 61.635 4.67 ;
      RECT 61.62 4.396 61.63 4.67 ;
      RECT 61.585 4.4 61.62 4.668 ;
      RECT 61.535 4.41 61.585 4.655 ;
      RECT 61.515 4.418 61.535 4.64 ;
      RECT 61.435 4.43 61.515 4.623 ;
      RECT 61.6 3.98 61.77 4.19 ;
      RECT 61.716 3.976 61.77 4.19 ;
      RECT 61.521 3.98 61.77 4.181 ;
      RECT 61.521 3.98 61.775 4.17 ;
      RECT 61.435 3.98 61.775 4.161 ;
      RECT 61.435 3.988 61.785 4.105 ;
      RECT 61.435 4 61.79 4.018 ;
      RECT 61.435 4.007 61.795 4.01 ;
      RECT 61.63 3.978 61.77 4.19 ;
      RECT 61.385 4.923 61.63 5.255 ;
      RECT 61.38 4.915 61.385 5.252 ;
      RECT 61.35 4.935 61.63 5.233 ;
      RECT 61.33 4.967 61.63 5.206 ;
      RECT 61.38 4.92 61.557 5.252 ;
      RECT 61.38 4.917 61.471 5.252 ;
      RECT 61.32 3.265 61.49 3.685 ;
      RECT 61.315 3.265 61.49 3.683 ;
      RECT 61.315 3.265 61.515 3.673 ;
      RECT 61.315 3.265 61.535 3.648 ;
      RECT 61.31 3.265 61.535 3.643 ;
      RECT 61.31 3.265 61.545 3.633 ;
      RECT 61.31 3.265 61.55 3.628 ;
      RECT 61.31 3.27 61.555 3.623 ;
      RECT 61.31 3.302 61.57 3.613 ;
      RECT 61.31 3.372 61.595 3.596 ;
      RECT 61.29 3.372 61.595 3.588 ;
      RECT 61.29 3.432 61.605 3.565 ;
      RECT 61.29 3.472 61.615 3.51 ;
      RECT 61.275 3.265 61.55 3.49 ;
      RECT 61.265 3.28 61.555 3.388 ;
      RECT 60.855 4.67 61.025 5.195 ;
      RECT 60.85 4.67 61.025 5.188 ;
      RECT 60.84 4.67 61.03 5.153 ;
      RECT 60.835 4.68 61.03 5.125 ;
      RECT 60.83 4.7 61.03 5.108 ;
      RECT 60.84 4.675 61.035 5.098 ;
      RECT 60.825 4.72 61.035 5.09 ;
      RECT 60.82 4.74 61.035 5.075 ;
      RECT 60.815 4.77 61.035 5.065 ;
      RECT 60.805 4.815 61.035 5.04 ;
      RECT 60.835 4.685 61.04 5.023 ;
      RECT 60.8 4.867 61.04 5.018 ;
      RECT 60.835 4.695 61.045 4.988 ;
      RECT 60.795 4.9 61.045 4.985 ;
      RECT 60.79 4.925 61.045 4.965 ;
      RECT 60.83 4.712 61.055 4.905 ;
      RECT 60.825 4.734 61.065 4.798 ;
      RECT 60.775 3.981 60.79 4.25 ;
      RECT 60.73 3.965 60.775 4.295 ;
      RECT 60.725 3.953 60.73 4.345 ;
      RECT 60.715 3.949 60.725 4.378 ;
      RECT 60.71 3.946 60.715 4.406 ;
      RECT 60.695 3.948 60.71 4.448 ;
      RECT 60.69 3.952 60.695 4.488 ;
      RECT 60.67 3.957 60.69 4.54 ;
      RECT 60.666 3.962 60.67 4.597 ;
      RECT 60.58 3.981 60.666 4.634 ;
      RECT 60.57 4.002 60.58 4.67 ;
      RECT 60.565 4.01 60.57 4.671 ;
      RECT 60.56 4.052 60.565 4.672 ;
      RECT 60.545 4.14 60.56 4.673 ;
      RECT 60.535 4.29 60.545 4.675 ;
      RECT 60.53 4.335 60.535 4.677 ;
      RECT 60.495 4.377 60.53 4.68 ;
      RECT 60.49 4.395 60.495 4.683 ;
      RECT 60.413 4.401 60.49 4.689 ;
      RECT 60.327 4.415 60.413 4.702 ;
      RECT 60.241 4.429 60.327 4.716 ;
      RECT 60.155 4.443 60.241 4.729 ;
      RECT 60.095 4.455 60.155 4.741 ;
      RECT 60.07 4.462 60.095 4.748 ;
      RECT 60.056 4.465 60.07 4.753 ;
      RECT 59.97 4.473 60.056 4.769 ;
      RECT 59.965 4.48 59.97 4.784 ;
      RECT 59.941 4.48 59.965 4.791 ;
      RECT 59.855 4.483 59.941 4.819 ;
      RECT 59.77 4.487 59.855 4.863 ;
      RECT 59.705 4.491 59.77 4.9 ;
      RECT 59.68 4.494 59.705 4.916 ;
      RECT 59.605 4.507 59.68 4.92 ;
      RECT 59.58 4.525 59.605 4.924 ;
      RECT 59.57 4.532 59.58 4.926 ;
      RECT 59.555 4.535 59.57 4.927 ;
      RECT 59.495 4.547 59.555 4.931 ;
      RECT 59.485 4.561 59.495 4.935 ;
      RECT 59.43 4.571 59.485 4.923 ;
      RECT 59.405 4.592 59.43 4.906 ;
      RECT 59.385 4.612 59.405 4.897 ;
      RECT 59.38 4.625 59.385 4.892 ;
      RECT 59.365 4.637 59.38 4.888 ;
      RECT 60.6 3.292 60.605 3.315 ;
      RECT 60.595 3.283 60.6 3.355 ;
      RECT 60.59 3.281 60.595 3.398 ;
      RECT 60.585 3.272 60.59 3.433 ;
      RECT 60.58 3.262 60.585 3.505 ;
      RECT 60.575 3.252 60.58 3.57 ;
      RECT 60.57 3.249 60.575 3.61 ;
      RECT 60.545 3.243 60.57 3.7 ;
      RECT 60.51 3.231 60.545 3.725 ;
      RECT 60.5 3.222 60.51 3.725 ;
      RECT 60.365 3.22 60.375 3.708 ;
      RECT 60.355 3.22 60.365 3.675 ;
      RECT 60.35 3.22 60.355 3.65 ;
      RECT 60.345 3.22 60.35 3.638 ;
      RECT 60.34 3.22 60.345 3.62 ;
      RECT 60.33 3.22 60.34 3.585 ;
      RECT 60.325 3.222 60.33 3.563 ;
      RECT 60.32 3.228 60.325 3.548 ;
      RECT 60.315 3.234 60.32 3.533 ;
      RECT 60.3 3.246 60.315 3.506 ;
      RECT 60.295 3.257 60.3 3.474 ;
      RECT 60.29 3.267 60.295 3.458 ;
      RECT 60.28 3.275 60.29 3.427 ;
      RECT 60.275 3.285 60.28 3.401 ;
      RECT 60.27 3.342 60.275 3.384 ;
      RECT 60.375 3.22 60.5 3.725 ;
      RECT 60.09 3.907 60.35 4.205 ;
      RECT 60.085 3.914 60.35 4.203 ;
      RECT 60.09 3.909 60.365 4.198 ;
      RECT 60.08 3.922 60.365 4.195 ;
      RECT 60.08 3.927 60.37 4.188 ;
      RECT 60.075 3.935 60.37 4.185 ;
      RECT 60.075 3.952 60.375 3.983 ;
      RECT 60.09 3.904 60.321 4.205 ;
      RECT 60.145 3.903 60.321 4.205 ;
      RECT 60.145 3.9 60.235 4.205 ;
      RECT 60.145 3.897 60.231 4.205 ;
      RECT 59.835 4.17 59.84 4.183 ;
      RECT 59.83 4.137 59.835 4.188 ;
      RECT 59.825 4.092 59.83 4.195 ;
      RECT 59.82 4.047 59.825 4.203 ;
      RECT 59.815 4.015 59.82 4.211 ;
      RECT 59.81 3.975 59.815 4.212 ;
      RECT 59.795 3.955 59.81 4.214 ;
      RECT 59.72 3.937 59.795 4.226 ;
      RECT 59.71 3.93 59.72 4.237 ;
      RECT 59.705 3.93 59.71 4.239 ;
      RECT 59.675 3.936 59.705 4.243 ;
      RECT 59.635 3.949 59.675 4.243 ;
      RECT 59.61 3.96 59.635 4.229 ;
      RECT 59.595 3.966 59.61 4.212 ;
      RECT 59.585 3.968 59.595 4.203 ;
      RECT 59.58 3.969 59.585 4.198 ;
      RECT 59.575 3.97 59.58 4.193 ;
      RECT 59.57 3.971 59.575 4.19 ;
      RECT 59.545 3.976 59.57 4.18 ;
      RECT 59.535 3.992 59.545 4.167 ;
      RECT 59.53 4.012 59.535 4.162 ;
      RECT 59.54 3.405 59.545 3.601 ;
      RECT 59.525 3.369 59.54 3.603 ;
      RECT 59.515 3.351 59.525 3.608 ;
      RECT 59.505 3.337 59.515 3.612 ;
      RECT 59.46 3.321 59.505 3.622 ;
      RECT 59.455 3.311 59.46 3.631 ;
      RECT 59.41 3.3 59.455 3.637 ;
      RECT 59.405 3.288 59.41 3.644 ;
      RECT 59.39 3.283 59.405 3.648 ;
      RECT 59.375 3.275 59.39 3.653 ;
      RECT 59.365 3.268 59.375 3.658 ;
      RECT 59.355 3.265 59.365 3.663 ;
      RECT 59.345 3.265 59.355 3.664 ;
      RECT 59.34 3.262 59.345 3.663 ;
      RECT 59.305 3.257 59.33 3.662 ;
      RECT 59.281 3.253 59.305 3.661 ;
      RECT 59.195 3.244 59.281 3.658 ;
      RECT 59.18 3.236 59.195 3.655 ;
      RECT 59.158 3.235 59.18 3.654 ;
      RECT 59.072 3.235 59.158 3.652 ;
      RECT 58.986 3.235 59.072 3.65 ;
      RECT 58.9 3.235 58.986 3.647 ;
      RECT 58.89 3.235 58.9 3.638 ;
      RECT 58.86 3.235 58.89 3.598 ;
      RECT 58.85 3.245 58.86 3.553 ;
      RECT 58.845 3.285 58.85 3.538 ;
      RECT 58.84 3.3 58.845 3.525 ;
      RECT 58.81 3.38 58.84 3.487 ;
      RECT 59.33 3.26 59.34 3.663 ;
      RECT 59.155 4.025 59.17 4.63 ;
      RECT 59.16 4.02 59.17 4.63 ;
      RECT 59.325 4.02 59.33 4.203 ;
      RECT 59.315 4.02 59.325 4.233 ;
      RECT 59.3 4.02 59.315 4.293 ;
      RECT 59.295 4.02 59.3 4.338 ;
      RECT 59.29 4.02 59.295 4.368 ;
      RECT 59.285 4.02 59.29 4.388 ;
      RECT 59.275 4.02 59.285 4.423 ;
      RECT 59.26 4.02 59.275 4.455 ;
      RECT 59.215 4.02 59.26 4.483 ;
      RECT 59.21 4.02 59.215 4.513 ;
      RECT 59.205 4.02 59.21 4.525 ;
      RECT 59.2 4.02 59.205 4.533 ;
      RECT 59.19 4.02 59.2 4.548 ;
      RECT 59.185 4.02 59.19 4.57 ;
      RECT 59.175 4.02 59.185 4.593 ;
      RECT 59.17 4.02 59.175 4.613 ;
      RECT 59.135 4.035 59.155 4.63 ;
      RECT 59.11 4.052 59.135 4.63 ;
      RECT 59.105 4.062 59.11 4.63 ;
      RECT 59.075 4.077 59.105 4.63 ;
      RECT 59 4.119 59.075 4.63 ;
      RECT 58.995 4.15 59 4.613 ;
      RECT 58.99 4.154 58.995 4.595 ;
      RECT 58.985 4.158 58.99 4.558 ;
      RECT 58.98 4.342 58.985 4.525 ;
      RECT 58.465 4.531 58.551 5.096 ;
      RECT 58.42 4.533 58.585 5.09 ;
      RECT 58.551 4.53 58.585 5.09 ;
      RECT 58.465 4.532 58.67 5.084 ;
      RECT 58.42 4.542 58.68 5.08 ;
      RECT 58.395 4.534 58.67 5.076 ;
      RECT 58.39 4.537 58.67 5.071 ;
      RECT 58.365 4.552 58.68 5.065 ;
      RECT 58.365 4.577 58.72 5.06 ;
      RECT 58.325 4.585 58.72 5.035 ;
      RECT 58.325 4.612 58.735 5.033 ;
      RECT 58.325 4.642 58.745 5.02 ;
      RECT 58.32 4.787 58.745 5.008 ;
      RECT 58.325 4.716 58.765 5.005 ;
      RECT 58.325 4.773 58.77 4.813 ;
      RECT 58.515 4.052 58.685 4.23 ;
      RECT 58.465 3.991 58.515 4.215 ;
      RECT 58.2 3.971 58.465 4.2 ;
      RECT 58.16 4.035 58.635 4.2 ;
      RECT 58.16 4.025 58.59 4.2 ;
      RECT 58.16 4.022 58.58 4.2 ;
      RECT 58.16 4.01 58.57 4.2 ;
      RECT 58.16 3.995 58.515 4.2 ;
      RECT 58.2 3.967 58.401 4.2 ;
      RECT 58.21 3.945 58.401 4.2 ;
      RECT 58.235 3.93 58.315 4.2 ;
      RECT 57.99 4.46 58.11 4.905 ;
      RECT 57.975 4.46 58.11 4.904 ;
      RECT 57.93 4.482 58.11 4.899 ;
      RECT 57.89 4.531 58.11 4.893 ;
      RECT 57.89 4.531 58.115 4.868 ;
      RECT 57.89 4.531 58.135 4.758 ;
      RECT 57.885 4.561 58.135 4.755 ;
      RECT 57.975 4.46 58.145 4.65 ;
      RECT 57.635 3.245 57.64 3.69 ;
      RECT 57.445 3.245 57.465 3.655 ;
      RECT 57.415 3.245 57.42 3.63 ;
      RECT 58.095 3.552 58.11 3.74 ;
      RECT 58.09 3.537 58.095 3.746 ;
      RECT 58.07 3.51 58.09 3.749 ;
      RECT 58.02 3.477 58.07 3.758 ;
      RECT 57.99 3.457 58.02 3.762 ;
      RECT 57.971 3.445 57.99 3.758 ;
      RECT 57.885 3.417 57.971 3.748 ;
      RECT 57.875 3.392 57.885 3.738 ;
      RECT 57.805 3.36 57.875 3.73 ;
      RECT 57.78 3.32 57.805 3.722 ;
      RECT 57.76 3.302 57.78 3.716 ;
      RECT 57.75 3.292 57.76 3.713 ;
      RECT 57.74 3.285 57.75 3.711 ;
      RECT 57.72 3.272 57.74 3.708 ;
      RECT 57.71 3.262 57.72 3.705 ;
      RECT 57.7 3.255 57.71 3.703 ;
      RECT 57.65 3.247 57.7 3.697 ;
      RECT 57.64 3.245 57.65 3.691 ;
      RECT 57.61 3.245 57.635 3.688 ;
      RECT 57.581 3.245 57.61 3.683 ;
      RECT 57.495 3.245 57.581 3.673 ;
      RECT 57.465 3.245 57.495 3.66 ;
      RECT 57.42 3.245 57.445 3.643 ;
      RECT 57.405 3.245 57.415 3.625 ;
      RECT 57.385 3.252 57.405 3.61 ;
      RECT 57.38 3.267 57.385 3.598 ;
      RECT 57.375 3.272 57.38 3.538 ;
      RECT 57.37 3.277 57.375 3.38 ;
      RECT 57.365 3.28 57.37 3.298 ;
      RECT 57.105 4.57 57.14 4.89 ;
      RECT 57.69 4.755 57.695 4.937 ;
      RECT 57.645 4.637 57.69 4.956 ;
      RECT 57.63 4.614 57.645 4.979 ;
      RECT 57.62 4.604 57.63 4.989 ;
      RECT 57.6 4.599 57.62 5.002 ;
      RECT 57.575 4.597 57.6 5.023 ;
      RECT 57.556 4.596 57.575 5.035 ;
      RECT 57.47 4.593 57.556 5.035 ;
      RECT 57.4 4.588 57.47 5.023 ;
      RECT 57.325 4.584 57.4 4.998 ;
      RECT 57.26 4.58 57.325 4.965 ;
      RECT 57.19 4.577 57.26 4.925 ;
      RECT 57.16 4.573 57.19 4.9 ;
      RECT 57.14 4.571 57.16 4.893 ;
      RECT 57.056 4.569 57.105 4.891 ;
      RECT 56.97 4.566 57.056 4.892 ;
      RECT 56.895 4.565 56.97 4.894 ;
      RECT 56.81 4.565 56.895 4.92 ;
      RECT 56.733 4.566 56.81 4.945 ;
      RECT 56.647 4.567 56.733 4.945 ;
      RECT 56.561 4.567 56.647 4.945 ;
      RECT 56.475 4.568 56.561 4.945 ;
      RECT 56.455 4.569 56.475 4.937 ;
      RECT 56.44 4.575 56.455 4.922 ;
      RECT 56.405 4.595 56.44 4.902 ;
      RECT 56.395 4.615 56.405 4.884 ;
      RECT 57.365 3.92 57.37 4.19 ;
      RECT 57.36 3.911 57.365 4.195 ;
      RECT 57.35 3.901 57.36 4.207 ;
      RECT 57.345 3.89 57.35 4.218 ;
      RECT 57.325 3.884 57.345 4.236 ;
      RECT 57.28 3.881 57.325 4.285 ;
      RECT 57.265 3.88 57.28 4.33 ;
      RECT 57.26 3.88 57.265 4.343 ;
      RECT 57.25 3.88 57.26 4.355 ;
      RECT 57.245 3.881 57.25 4.37 ;
      RECT 57.225 3.889 57.245 4.375 ;
      RECT 57.195 3.905 57.225 4.375 ;
      RECT 57.185 3.917 57.19 4.375 ;
      RECT 57.15 3.932 57.185 4.375 ;
      RECT 57.12 3.952 57.15 4.375 ;
      RECT 57.11 3.977 57.12 4.375 ;
      RECT 57.105 4.005 57.11 4.375 ;
      RECT 57.1 4.035 57.105 4.375 ;
      RECT 57.095 4.052 57.1 4.375 ;
      RECT 57.085 4.08 57.095 4.375 ;
      RECT 57.075 4.115 57.085 4.375 ;
      RECT 57.07 4.15 57.075 4.375 ;
      RECT 57.19 3.915 57.195 4.375 ;
      RECT 56.37 3.975 56.89 4.19 ;
      RECT 56.45 3.915 56.89 4.19 ;
      RECT 56.18 3.245 56.185 3.644 ;
      RECT 55.925 3.245 55.96 3.642 ;
      RECT 55.52 3.28 55.525 3.636 ;
      RECT 56.265 3.283 56.27 3.538 ;
      RECT 56.26 3.281 56.265 3.544 ;
      RECT 56.255 3.28 56.26 3.551 ;
      RECT 56.23 3.273 56.255 3.575 ;
      RECT 56.225 3.266 56.23 3.599 ;
      RECT 56.22 3.262 56.225 3.608 ;
      RECT 56.21 3.257 56.22 3.621 ;
      RECT 56.205 3.254 56.21 3.63 ;
      RECT 56.2 3.252 56.205 3.635 ;
      RECT 56.185 3.248 56.2 3.645 ;
      RECT 56.17 3.242 56.18 3.644 ;
      RECT 56.132 3.24 56.17 3.644 ;
      RECT 56.046 3.242 56.132 3.644 ;
      RECT 55.96 3.244 56.046 3.643 ;
      RECT 55.889 3.245 55.925 3.642 ;
      RECT 55.803 3.247 55.889 3.642 ;
      RECT 55.717 3.249 55.803 3.641 ;
      RECT 55.631 3.251 55.717 3.641 ;
      RECT 55.545 3.254 55.631 3.64 ;
      RECT 55.535 3.26 55.545 3.639 ;
      RECT 55.525 3.272 55.535 3.637 ;
      RECT 55.465 3.307 55.52 3.633 ;
      RECT 55.46 3.337 55.465 3.395 ;
      RECT 55.805 4.552 55.81 4.809 ;
      RECT 55.785 4.471 55.805 4.826 ;
      RECT 55.765 4.465 55.785 4.855 ;
      RECT 55.705 4.452 55.765 4.875 ;
      RECT 55.66 4.436 55.705 4.876 ;
      RECT 55.576 4.424 55.66 4.864 ;
      RECT 55.49 4.411 55.576 4.848 ;
      RECT 55.48 4.404 55.49 4.84 ;
      RECT 55.435 4.401 55.48 4.78 ;
      RECT 55.415 4.397 55.435 4.695 ;
      RECT 55.4 4.395 55.415 4.648 ;
      RECT 55.37 4.392 55.4 4.618 ;
      RECT 55.335 4.388 55.37 4.595 ;
      RECT 55.292 4.383 55.335 4.583 ;
      RECT 55.206 4.374 55.292 4.592 ;
      RECT 55.12 4.363 55.206 4.604 ;
      RECT 55.055 4.354 55.12 4.613 ;
      RECT 55.035 4.345 55.055 4.618 ;
      RECT 55.03 4.338 55.035 4.62 ;
      RECT 54.99 4.323 55.03 4.617 ;
      RECT 54.97 4.302 54.99 4.612 ;
      RECT 54.955 4.29 54.97 4.605 ;
      RECT 54.95 4.282 54.955 4.598 ;
      RECT 54.935 4.262 54.95 4.591 ;
      RECT 54.93 4.125 54.935 4.585 ;
      RECT 54.85 4.014 54.93 4.557 ;
      RECT 54.841 4.007 54.85 4.523 ;
      RECT 54.755 4.001 54.841 4.448 ;
      RECT 54.73 3.992 54.755 4.36 ;
      RECT 54.7 3.987 54.73 4.335 ;
      RECT 54.635 3.996 54.7 4.32 ;
      RECT 54.615 4.012 54.635 4.295 ;
      RECT 54.605 4.018 54.615 4.243 ;
      RECT 54.585 4.04 54.605 4.125 ;
      RECT 55.24 4.005 55.41 4.19 ;
      RECT 55.24 4.005 55.445 4.188 ;
      RECT 55.29 3.915 55.46 4.179 ;
      RECT 55.24 4.072 55.465 4.172 ;
      RECT 55.255 3.95 55.46 4.179 ;
      RECT 54.455 4.683 54.52 5.126 ;
      RECT 54.395 4.708 54.52 5.124 ;
      RECT 54.395 4.708 54.575 5.118 ;
      RECT 54.38 4.733 54.575 5.117 ;
      RECT 54.52 4.67 54.595 5.114 ;
      RECT 54.455 4.695 54.675 5.108 ;
      RECT 54.38 4.734 54.72 5.102 ;
      RECT 54.365 4.761 54.72 5.093 ;
      RECT 54.38 4.754 54.74 5.085 ;
      RECT 54.365 4.763 54.745 5.068 ;
      RECT 54.36 4.78 54.745 4.895 ;
      RECT 54.365 3.502 54.4 3.74 ;
      RECT 54.365 3.502 54.43 3.739 ;
      RECT 54.365 3.502 54.545 3.735 ;
      RECT 54.365 3.502 54.6 3.713 ;
      RECT 54.375 3.445 54.655 3.613 ;
      RECT 54.48 3.285 54.51 3.736 ;
      RECT 54.51 3.28 54.69 3.493 ;
      RECT 54.38 3.421 54.69 3.493 ;
      RECT 54.43 3.317 54.48 3.737 ;
      RECT 54.4 3.373 54.69 3.493 ;
      RECT 53.26 7.455 53.43 8.925 ;
      RECT 53.26 7.455 53.435 8.715 ;
      RECT 52.89 9.405 53.36 9.575 ;
      RECT 52.89 8.385 53.06 9.575 ;
      RECT 52.885 3.035 53.055 4.225 ;
      RECT 52.885 3.035 53.355 3.205 ;
      RECT 52.27 3.895 52.445 5.155 ;
      RECT 52.27 3.685 52.44 5.155 ;
      RECT 52.27 7.455 52.44 8.925 ;
      RECT 52.27 7.455 52.445 8.715 ;
      RECT 51.9 3.035 52.07 4.225 ;
      RECT 51.9 3.035 52.37 3.205 ;
      RECT 51.9 9.405 52.37 9.575 ;
      RECT 51.9 8.385 52.07 9.575 ;
      RECT 50.91 4.015 51.085 5.155 ;
      RECT 50.91 1.865 51.08 5.155 ;
      RECT 50.91 1.865 51.085 2.415 ;
      RECT 50.91 10.195 51.085 10.745 ;
      RECT 50.91 7.455 51.08 10.745 ;
      RECT 50.91 7.455 51.085 8.595 ;
      RECT 50.48 3.895 50.655 5.155 ;
      RECT 50.48 2.945 50.65 5.155 ;
      RECT 50.48 7.455 50.65 9.665 ;
      RECT 50.48 7.455 50.655 8.715 ;
      RECT 50.05 3.925 50.22 5.155 ;
      RECT 50.11 2.145 50.28 4.095 ;
      RECT 50.05 1.865 50.22 2.315 ;
      RECT 50.05 10.295 50.22 10.745 ;
      RECT 50.11 8.515 50.28 10.465 ;
      RECT 50.05 7.455 50.22 8.685 ;
      RECT 49.525 3.895 49.7 5.155 ;
      RECT 49.525 1.865 49.695 5.155 ;
      RECT 49.525 3.365 49.935 3.695 ;
      RECT 49.525 2.525 49.935 2.855 ;
      RECT 49.525 1.865 49.7 2.355 ;
      RECT 49.525 10.255 49.7 10.745 ;
      RECT 49.525 7.455 49.695 10.745 ;
      RECT 49.525 9.755 49.935 10.085 ;
      RECT 49.525 8.915 49.935 9.245 ;
      RECT 49.525 7.455 49.7 8.715 ;
      RECT 47.64 4.687 47.655 4.738 ;
      RECT 47.635 4.667 47.64 4.785 ;
      RECT 47.62 4.657 47.635 4.853 ;
      RECT 47.595 4.637 47.62 4.908 ;
      RECT 47.555 4.622 47.595 4.928 ;
      RECT 47.51 4.616 47.555 4.956 ;
      RECT 47.44 4.606 47.51 4.973 ;
      RECT 47.42 4.598 47.44 4.973 ;
      RECT 47.36 4.592 47.42 4.965 ;
      RECT 47.301 4.583 47.36 4.953 ;
      RECT 47.215 4.572 47.301 4.936 ;
      RECT 47.193 4.563 47.215 4.924 ;
      RECT 47.107 4.556 47.193 4.911 ;
      RECT 47.021 4.543 47.107 4.892 ;
      RECT 46.935 4.531 47.021 4.872 ;
      RECT 46.905 4.52 46.935 4.859 ;
      RECT 46.855 4.506 46.905 4.851 ;
      RECT 46.835 4.495 46.855 4.843 ;
      RECT 46.786 4.484 46.835 4.835 ;
      RECT 46.7 4.463 46.786 4.82 ;
      RECT 46.655 4.45 46.7 4.805 ;
      RECT 46.61 4.45 46.655 4.785 ;
      RECT 46.555 4.45 46.61 4.72 ;
      RECT 46.53 4.45 46.555 4.643 ;
      RECT 47.055 4.187 47.225 4.37 ;
      RECT 47.055 4.187 47.24 4.328 ;
      RECT 47.055 4.187 47.245 4.27 ;
      RECT 47.115 3.955 47.25 4.246 ;
      RECT 47.115 3.959 47.255 4.229 ;
      RECT 47.06 4.122 47.255 4.229 ;
      RECT 47.085 3.967 47.225 4.37 ;
      RECT 47.085 3.971 47.265 4.17 ;
      RECT 47.07 4.057 47.265 4.17 ;
      RECT 47.08 3.987 47.225 4.37 ;
      RECT 47.08 3.99 47.275 4.083 ;
      RECT 47.075 4.007 47.275 4.083 ;
      RECT 46.845 3.227 47.015 3.71 ;
      RECT 46.84 3.222 46.99 3.7 ;
      RECT 46.84 3.229 47.02 3.694 ;
      RECT 46.83 3.223 46.99 3.673 ;
      RECT 46.83 3.239 47.035 3.632 ;
      RECT 46.8 3.224 46.99 3.595 ;
      RECT 46.8 3.254 47.045 3.535 ;
      RECT 46.795 3.226 46.99 3.533 ;
      RECT 46.775 3.235 47.02 3.49 ;
      RECT 46.75 3.251 47.035 3.402 ;
      RECT 46.75 3.27 47.06 3.393 ;
      RECT 46.745 3.307 47.06 3.345 ;
      RECT 46.75 3.287 47.065 3.313 ;
      RECT 46.845 3.221 46.955 3.71 ;
      RECT 46.931 3.22 46.955 3.71 ;
      RECT 46.165 4.005 46.17 4.216 ;
      RECT 46.765 4.005 46.77 4.19 ;
      RECT 46.83 4.045 46.835 4.158 ;
      RECT 46.825 4.037 46.83 4.164 ;
      RECT 46.82 4.027 46.825 4.172 ;
      RECT 46.815 4.017 46.82 4.181 ;
      RECT 46.81 4.007 46.815 4.185 ;
      RECT 46.77 4.005 46.81 4.188 ;
      RECT 46.742 4.004 46.765 4.192 ;
      RECT 46.656 4.001 46.742 4.199 ;
      RECT 46.57 3.997 46.656 4.21 ;
      RECT 46.55 3.995 46.57 4.216 ;
      RECT 46.532 3.994 46.55 4.219 ;
      RECT 46.446 3.992 46.532 4.226 ;
      RECT 46.36 3.987 46.446 4.239 ;
      RECT 46.341 3.984 46.36 4.244 ;
      RECT 46.255 3.982 46.341 4.235 ;
      RECT 46.245 3.982 46.255 4.228 ;
      RECT 46.17 3.995 46.245 4.222 ;
      RECT 46.155 4.006 46.165 4.216 ;
      RECT 46.145 4.008 46.155 4.215 ;
      RECT 46.135 4.012 46.145 4.211 ;
      RECT 46.13 4.015 46.135 4.205 ;
      RECT 46.12 4.017 46.13 4.199 ;
      RECT 46.115 4.02 46.12 4.193 ;
      RECT 46.15 10.195 46.325 10.745 ;
      RECT 46.15 7.455 46.32 10.745 ;
      RECT 46.15 7.455 46.325 8.595 ;
      RECT 46.095 4.606 46.1 4.81 ;
      RECT 46.08 4.593 46.095 4.903 ;
      RECT 46.065 4.574 46.08 5.18 ;
      RECT 46.03 4.54 46.065 5.18 ;
      RECT 46.026 4.51 46.03 5.18 ;
      RECT 45.94 4.392 46.026 5.18 ;
      RECT 45.93 4.267 45.94 5.18 ;
      RECT 45.915 4.235 45.93 5.18 ;
      RECT 45.91 4.21 45.915 5.18 ;
      RECT 45.905 4.2 45.91 5.136 ;
      RECT 45.89 4.172 45.905 5.041 ;
      RECT 45.875 4.138 45.89 4.94 ;
      RECT 45.87 4.116 45.875 4.893 ;
      RECT 45.865 4.105 45.87 4.863 ;
      RECT 45.86 4.095 45.865 4.829 ;
      RECT 45.85 4.082 45.86 4.797 ;
      RECT 45.825 4.058 45.85 4.723 ;
      RECT 45.82 4.038 45.825 4.648 ;
      RECT 45.815 4.032 45.82 4.623 ;
      RECT 45.81 4.027 45.815 4.588 ;
      RECT 45.805 4.022 45.81 4.563 ;
      RECT 45.8 4.02 45.805 4.543 ;
      RECT 45.795 4.02 45.8 4.528 ;
      RECT 45.79 4.02 45.795 4.488 ;
      RECT 45.78 4.02 45.79 4.46 ;
      RECT 45.77 4.02 45.78 4.405 ;
      RECT 45.755 4.02 45.77 4.343 ;
      RECT 45.75 4.019 45.755 4.288 ;
      RECT 45.735 4.018 45.75 4.268 ;
      RECT 45.675 4.016 45.735 4.242 ;
      RECT 45.64 4.017 45.675 4.222 ;
      RECT 45.635 4.019 45.64 4.212 ;
      RECT 45.625 4.038 45.635 4.202 ;
      RECT 45.62 4.065 45.625 4.133 ;
      RECT 45.735 3.49 45.905 3.735 ;
      RECT 45.77 3.261 45.905 3.735 ;
      RECT 45.77 3.263 45.915 3.73 ;
      RECT 45.77 3.265 45.94 3.718 ;
      RECT 45.77 3.268 45.965 3.7 ;
      RECT 45.77 3.273 46.015 3.673 ;
      RECT 45.77 3.278 46.035 3.638 ;
      RECT 45.75 3.28 46.045 3.613 ;
      RECT 45.74 3.375 46.045 3.613 ;
      RECT 45.77 3.26 45.88 3.735 ;
      RECT 45.78 3.257 45.875 3.735 ;
      RECT 45.72 7.455 45.89 9.665 ;
      RECT 45.72 7.455 45.895 8.715 ;
      RECT 45.3 4.522 45.49 4.88 ;
      RECT 45.3 4.534 45.525 4.879 ;
      RECT 45.3 4.562 45.545 4.877 ;
      RECT 45.3 4.587 45.55 4.876 ;
      RECT 45.3 4.645 45.565 4.875 ;
      RECT 45.285 4.518 45.445 4.86 ;
      RECT 45.265 4.527 45.49 4.813 ;
      RECT 45.24 4.538 45.525 4.75 ;
      RECT 45.24 4.622 45.56 4.75 ;
      RECT 45.24 4.597 45.555 4.75 ;
      RECT 45.3 4.513 45.445 4.88 ;
      RECT 45.386 4.512 45.445 4.88 ;
      RECT 45.386 4.511 45.43 4.88 ;
      RECT 44.765 10.255 44.94 10.745 ;
      RECT 44.765 7.455 44.935 10.745 ;
      RECT 44.765 9.755 45.175 10.085 ;
      RECT 44.765 8.915 45.175 9.245 ;
      RECT 44.765 7.455 44.94 8.715 ;
      RECT 45.085 4.027 45.09 4.405 ;
      RECT 45.08 3.995 45.085 4.405 ;
      RECT 45.075 3.967 45.08 4.405 ;
      RECT 45.07 3.947 45.075 4.405 ;
      RECT 45.015 3.93 45.07 4.405 ;
      RECT 44.975 3.915 45.015 4.405 ;
      RECT 44.92 3.902 44.975 4.405 ;
      RECT 44.885 3.893 44.92 4.405 ;
      RECT 44.881 3.891 44.885 4.404 ;
      RECT 44.795 3.887 44.881 4.387 ;
      RECT 44.71 3.879 44.795 4.35 ;
      RECT 44.7 3.875 44.71 4.323 ;
      RECT 44.69 3.875 44.7 4.305 ;
      RECT 44.68 3.877 44.69 4.288 ;
      RECT 44.675 3.882 44.68 4.274 ;
      RECT 44.67 3.886 44.675 4.261 ;
      RECT 44.66 3.891 44.67 4.245 ;
      RECT 44.645 3.905 44.66 4.22 ;
      RECT 44.64 3.911 44.645 4.2 ;
      RECT 44.635 3.913 44.64 4.193 ;
      RECT 44.63 3.917 44.635 4.068 ;
      RECT 44.81 4.717 45.055 5.18 ;
      RECT 44.73 4.69 45.05 5.176 ;
      RECT 44.66 4.725 45.055 5.169 ;
      RECT 44.45 4.98 45.055 5.165 ;
      RECT 44.63 4.748 45.055 5.165 ;
      RECT 44.47 4.94 45.055 5.165 ;
      RECT 44.62 4.76 45.055 5.165 ;
      RECT 44.505 4.877 45.055 5.165 ;
      RECT 44.56 4.802 45.055 5.165 ;
      RECT 44.81 4.667 45.05 5.18 ;
      RECT 44.84 4.66 45.05 5.18 ;
      RECT 44.83 4.662 45.05 5.18 ;
      RECT 44.84 4.657 44.97 5.18 ;
      RECT 44.395 3.22 44.481 3.659 ;
      RECT 44.39 3.22 44.481 3.657 ;
      RECT 44.39 3.22 44.55 3.656 ;
      RECT 44.39 3.22 44.58 3.653 ;
      RECT 44.375 3.227 44.58 3.644 ;
      RECT 44.375 3.227 44.585 3.64 ;
      RECT 44.37 3.237 44.585 3.633 ;
      RECT 44.365 3.242 44.585 3.608 ;
      RECT 44.365 3.242 44.6 3.59 ;
      RECT 44.39 3.22 44.62 3.505 ;
      RECT 44.36 3.247 44.62 3.503 ;
      RECT 44.37 3.24 44.625 3.441 ;
      RECT 44.36 3.362 44.63 3.424 ;
      RECT 44.345 3.257 44.625 3.375 ;
      RECT 44.34 3.267 44.625 3.275 ;
      RECT 44.42 4.038 44.425 4.115 ;
      RECT 44.41 4.032 44.42 4.305 ;
      RECT 44.4 4.024 44.41 4.326 ;
      RECT 44.39 4.015 44.4 4.348 ;
      RECT 44.385 4.01 44.39 4.365 ;
      RECT 44.345 4.01 44.385 4.405 ;
      RECT 44.325 4.01 44.345 4.46 ;
      RECT 44.32 4.01 44.325 4.488 ;
      RECT 44.31 4.01 44.32 4.503 ;
      RECT 44.275 4.01 44.31 4.545 ;
      RECT 44.27 4.01 44.275 4.588 ;
      RECT 44.26 4.01 44.27 4.603 ;
      RECT 44.245 4.01 44.26 4.623 ;
      RECT 44.23 4.01 44.245 4.65 ;
      RECT 44.225 4.011 44.23 4.668 ;
      RECT 44.205 4.012 44.225 4.675 ;
      RECT 44.15 4.013 44.205 4.695 ;
      RECT 44.14 4.014 44.15 4.709 ;
      RECT 44.135 4.017 44.14 4.708 ;
      RECT 44.095 4.09 44.135 4.706 ;
      RECT 44.08 4.17 44.095 4.704 ;
      RECT 44.055 4.225 44.08 4.702 ;
      RECT 44.04 4.29 44.055 4.701 ;
      RECT 43.995 4.322 44.04 4.698 ;
      RECT 43.91 4.345 43.995 4.693 ;
      RECT 43.885 4.365 43.91 4.688 ;
      RECT 43.815 4.37 43.885 4.684 ;
      RECT 43.795 4.372 43.815 4.681 ;
      RECT 43.71 4.383 43.795 4.675 ;
      RECT 43.705 4.394 43.71 4.67 ;
      RECT 43.695 4.396 43.705 4.67 ;
      RECT 43.66 4.4 43.695 4.668 ;
      RECT 43.61 4.41 43.66 4.655 ;
      RECT 43.59 4.418 43.61 4.64 ;
      RECT 43.51 4.43 43.59 4.623 ;
      RECT 43.675 3.98 43.845 4.19 ;
      RECT 43.791 3.976 43.845 4.19 ;
      RECT 43.596 3.98 43.845 4.181 ;
      RECT 43.596 3.98 43.85 4.17 ;
      RECT 43.51 3.98 43.85 4.161 ;
      RECT 43.51 3.988 43.86 4.105 ;
      RECT 43.51 4 43.865 4.018 ;
      RECT 43.51 4.007 43.87 4.01 ;
      RECT 43.705 3.978 43.845 4.19 ;
      RECT 43.46 4.923 43.705 5.255 ;
      RECT 43.455 4.915 43.46 5.252 ;
      RECT 43.425 4.935 43.705 5.233 ;
      RECT 43.405 4.967 43.705 5.206 ;
      RECT 43.455 4.92 43.632 5.252 ;
      RECT 43.455 4.917 43.546 5.252 ;
      RECT 43.395 3.265 43.565 3.685 ;
      RECT 43.39 3.265 43.565 3.683 ;
      RECT 43.39 3.265 43.59 3.673 ;
      RECT 43.39 3.265 43.61 3.648 ;
      RECT 43.385 3.265 43.61 3.643 ;
      RECT 43.385 3.265 43.62 3.633 ;
      RECT 43.385 3.265 43.625 3.628 ;
      RECT 43.385 3.27 43.63 3.623 ;
      RECT 43.385 3.302 43.645 3.613 ;
      RECT 43.385 3.372 43.67 3.596 ;
      RECT 43.365 3.372 43.67 3.588 ;
      RECT 43.365 3.432 43.68 3.565 ;
      RECT 43.365 3.472 43.69 3.51 ;
      RECT 43.35 3.265 43.625 3.49 ;
      RECT 43.34 3.28 43.63 3.388 ;
      RECT 42.93 4.67 43.1 5.195 ;
      RECT 42.925 4.67 43.1 5.188 ;
      RECT 42.915 4.67 43.105 5.153 ;
      RECT 42.91 4.68 43.105 5.125 ;
      RECT 42.905 4.7 43.105 5.108 ;
      RECT 42.915 4.675 43.11 5.098 ;
      RECT 42.9 4.72 43.11 5.09 ;
      RECT 42.895 4.74 43.11 5.075 ;
      RECT 42.89 4.77 43.11 5.065 ;
      RECT 42.88 4.815 43.11 5.04 ;
      RECT 42.91 4.685 43.115 5.023 ;
      RECT 42.875 4.867 43.115 5.018 ;
      RECT 42.91 4.695 43.12 4.988 ;
      RECT 42.87 4.9 43.12 4.985 ;
      RECT 42.865 4.925 43.12 4.965 ;
      RECT 42.905 4.712 43.13 4.905 ;
      RECT 42.9 4.734 43.14 4.798 ;
      RECT 42.85 3.981 42.865 4.25 ;
      RECT 42.805 3.965 42.85 4.295 ;
      RECT 42.8 3.953 42.805 4.345 ;
      RECT 42.79 3.949 42.8 4.378 ;
      RECT 42.785 3.946 42.79 4.406 ;
      RECT 42.77 3.948 42.785 4.448 ;
      RECT 42.765 3.952 42.77 4.488 ;
      RECT 42.745 3.957 42.765 4.54 ;
      RECT 42.741 3.962 42.745 4.597 ;
      RECT 42.655 3.981 42.741 4.634 ;
      RECT 42.645 4.002 42.655 4.67 ;
      RECT 42.64 4.01 42.645 4.671 ;
      RECT 42.635 4.052 42.64 4.672 ;
      RECT 42.62 4.14 42.635 4.673 ;
      RECT 42.61 4.29 42.62 4.675 ;
      RECT 42.605 4.335 42.61 4.677 ;
      RECT 42.57 4.377 42.605 4.68 ;
      RECT 42.565 4.395 42.57 4.683 ;
      RECT 42.488 4.401 42.565 4.689 ;
      RECT 42.402 4.415 42.488 4.702 ;
      RECT 42.316 4.429 42.402 4.716 ;
      RECT 42.23 4.443 42.316 4.729 ;
      RECT 42.17 4.455 42.23 4.741 ;
      RECT 42.145 4.462 42.17 4.748 ;
      RECT 42.131 4.465 42.145 4.753 ;
      RECT 42.045 4.473 42.131 4.769 ;
      RECT 42.04 4.48 42.045 4.784 ;
      RECT 42.016 4.48 42.04 4.791 ;
      RECT 41.93 4.483 42.016 4.819 ;
      RECT 41.845 4.487 41.93 4.863 ;
      RECT 41.78 4.491 41.845 4.9 ;
      RECT 41.755 4.494 41.78 4.916 ;
      RECT 41.68 4.507 41.755 4.92 ;
      RECT 41.655 4.525 41.68 4.924 ;
      RECT 41.645 4.532 41.655 4.926 ;
      RECT 41.63 4.535 41.645 4.927 ;
      RECT 41.57 4.547 41.63 4.931 ;
      RECT 41.56 4.561 41.57 4.935 ;
      RECT 41.505 4.571 41.56 4.923 ;
      RECT 41.48 4.592 41.505 4.906 ;
      RECT 41.46 4.612 41.48 4.897 ;
      RECT 41.455 4.625 41.46 4.892 ;
      RECT 41.44 4.637 41.455 4.888 ;
      RECT 42.675 3.292 42.68 3.315 ;
      RECT 42.67 3.283 42.675 3.355 ;
      RECT 42.665 3.281 42.67 3.398 ;
      RECT 42.66 3.272 42.665 3.433 ;
      RECT 42.655 3.262 42.66 3.505 ;
      RECT 42.65 3.252 42.655 3.57 ;
      RECT 42.645 3.249 42.65 3.61 ;
      RECT 42.62 3.243 42.645 3.7 ;
      RECT 42.585 3.231 42.62 3.725 ;
      RECT 42.575 3.222 42.585 3.725 ;
      RECT 42.44 3.22 42.45 3.708 ;
      RECT 42.43 3.22 42.44 3.675 ;
      RECT 42.425 3.22 42.43 3.65 ;
      RECT 42.42 3.22 42.425 3.638 ;
      RECT 42.415 3.22 42.42 3.62 ;
      RECT 42.405 3.22 42.415 3.585 ;
      RECT 42.4 3.222 42.405 3.563 ;
      RECT 42.395 3.228 42.4 3.548 ;
      RECT 42.39 3.234 42.395 3.533 ;
      RECT 42.375 3.246 42.39 3.506 ;
      RECT 42.37 3.257 42.375 3.474 ;
      RECT 42.365 3.267 42.37 3.458 ;
      RECT 42.355 3.275 42.365 3.427 ;
      RECT 42.35 3.285 42.355 3.401 ;
      RECT 42.345 3.342 42.35 3.384 ;
      RECT 42.45 3.22 42.575 3.725 ;
      RECT 42.165 3.907 42.425 4.205 ;
      RECT 42.16 3.914 42.425 4.203 ;
      RECT 42.165 3.909 42.44 4.198 ;
      RECT 42.155 3.922 42.44 4.195 ;
      RECT 42.155 3.927 42.445 4.188 ;
      RECT 42.15 3.935 42.445 4.185 ;
      RECT 42.15 3.952 42.45 3.983 ;
      RECT 42.165 3.904 42.396 4.205 ;
      RECT 42.22 3.903 42.396 4.205 ;
      RECT 42.22 3.9 42.31 4.205 ;
      RECT 42.22 3.897 42.306 4.205 ;
      RECT 41.91 4.17 41.915 4.183 ;
      RECT 41.905 4.137 41.91 4.188 ;
      RECT 41.9 4.092 41.905 4.195 ;
      RECT 41.895 4.047 41.9 4.203 ;
      RECT 41.89 4.015 41.895 4.211 ;
      RECT 41.885 3.975 41.89 4.212 ;
      RECT 41.87 3.955 41.885 4.214 ;
      RECT 41.795 3.937 41.87 4.226 ;
      RECT 41.785 3.93 41.795 4.237 ;
      RECT 41.78 3.93 41.785 4.239 ;
      RECT 41.75 3.936 41.78 4.243 ;
      RECT 41.71 3.949 41.75 4.243 ;
      RECT 41.685 3.96 41.71 4.229 ;
      RECT 41.67 3.966 41.685 4.212 ;
      RECT 41.66 3.968 41.67 4.203 ;
      RECT 41.655 3.969 41.66 4.198 ;
      RECT 41.65 3.97 41.655 4.193 ;
      RECT 41.645 3.971 41.65 4.19 ;
      RECT 41.62 3.976 41.645 4.18 ;
      RECT 41.61 3.992 41.62 4.167 ;
      RECT 41.605 4.012 41.61 4.162 ;
      RECT 41.615 3.405 41.62 3.601 ;
      RECT 41.6 3.369 41.615 3.603 ;
      RECT 41.59 3.351 41.6 3.608 ;
      RECT 41.58 3.337 41.59 3.612 ;
      RECT 41.535 3.321 41.58 3.622 ;
      RECT 41.53 3.311 41.535 3.631 ;
      RECT 41.485 3.3 41.53 3.637 ;
      RECT 41.48 3.288 41.485 3.644 ;
      RECT 41.465 3.283 41.48 3.648 ;
      RECT 41.45 3.275 41.465 3.653 ;
      RECT 41.44 3.268 41.45 3.658 ;
      RECT 41.43 3.265 41.44 3.663 ;
      RECT 41.42 3.265 41.43 3.664 ;
      RECT 41.415 3.262 41.42 3.663 ;
      RECT 41.38 3.257 41.405 3.662 ;
      RECT 41.356 3.253 41.38 3.661 ;
      RECT 41.27 3.244 41.356 3.658 ;
      RECT 41.255 3.236 41.27 3.655 ;
      RECT 41.233 3.235 41.255 3.654 ;
      RECT 41.147 3.235 41.233 3.652 ;
      RECT 41.061 3.235 41.147 3.65 ;
      RECT 40.975 3.235 41.061 3.647 ;
      RECT 40.965 3.235 40.975 3.638 ;
      RECT 40.935 3.235 40.965 3.598 ;
      RECT 40.925 3.245 40.935 3.553 ;
      RECT 40.92 3.285 40.925 3.538 ;
      RECT 40.915 3.3 40.92 3.525 ;
      RECT 40.885 3.38 40.915 3.487 ;
      RECT 41.405 3.26 41.415 3.663 ;
      RECT 41.23 4.025 41.245 4.63 ;
      RECT 41.235 4.02 41.245 4.63 ;
      RECT 41.4 4.02 41.405 4.203 ;
      RECT 41.39 4.02 41.4 4.233 ;
      RECT 41.375 4.02 41.39 4.293 ;
      RECT 41.37 4.02 41.375 4.338 ;
      RECT 41.365 4.02 41.37 4.368 ;
      RECT 41.36 4.02 41.365 4.388 ;
      RECT 41.35 4.02 41.36 4.423 ;
      RECT 41.335 4.02 41.35 4.455 ;
      RECT 41.29 4.02 41.335 4.483 ;
      RECT 41.285 4.02 41.29 4.513 ;
      RECT 41.28 4.02 41.285 4.525 ;
      RECT 41.275 4.02 41.28 4.533 ;
      RECT 41.265 4.02 41.275 4.548 ;
      RECT 41.26 4.02 41.265 4.57 ;
      RECT 41.25 4.02 41.26 4.593 ;
      RECT 41.245 4.02 41.25 4.613 ;
      RECT 41.21 4.035 41.23 4.63 ;
      RECT 41.185 4.052 41.21 4.63 ;
      RECT 41.18 4.062 41.185 4.63 ;
      RECT 41.15 4.077 41.18 4.63 ;
      RECT 41.075 4.119 41.15 4.63 ;
      RECT 41.07 4.15 41.075 4.613 ;
      RECT 41.065 4.154 41.07 4.595 ;
      RECT 41.06 4.158 41.065 4.558 ;
      RECT 41.055 4.342 41.06 4.525 ;
      RECT 40.54 4.531 40.626 5.096 ;
      RECT 40.495 4.533 40.66 5.09 ;
      RECT 40.626 4.53 40.66 5.09 ;
      RECT 40.54 4.532 40.745 5.084 ;
      RECT 40.495 4.542 40.755 5.08 ;
      RECT 40.47 4.534 40.745 5.076 ;
      RECT 40.465 4.537 40.745 5.071 ;
      RECT 40.44 4.552 40.755 5.065 ;
      RECT 40.44 4.577 40.795 5.06 ;
      RECT 40.4 4.585 40.795 5.035 ;
      RECT 40.4 4.612 40.81 5.033 ;
      RECT 40.4 4.642 40.82 5.02 ;
      RECT 40.395 4.787 40.82 5.008 ;
      RECT 40.4 4.716 40.84 5.005 ;
      RECT 40.4 4.773 40.845 4.813 ;
      RECT 40.59 4.052 40.76 4.23 ;
      RECT 40.54 3.991 40.59 4.215 ;
      RECT 40.275 3.971 40.54 4.2 ;
      RECT 40.235 4.035 40.71 4.2 ;
      RECT 40.235 4.025 40.665 4.2 ;
      RECT 40.235 4.022 40.655 4.2 ;
      RECT 40.235 4.01 40.645 4.2 ;
      RECT 40.235 3.995 40.59 4.2 ;
      RECT 40.275 3.967 40.476 4.2 ;
      RECT 40.285 3.945 40.476 4.2 ;
      RECT 40.31 3.93 40.39 4.2 ;
      RECT 40.065 4.46 40.185 4.905 ;
      RECT 40.05 4.46 40.185 4.904 ;
      RECT 40.005 4.482 40.185 4.899 ;
      RECT 39.965 4.531 40.185 4.893 ;
      RECT 39.965 4.531 40.19 4.868 ;
      RECT 39.965 4.531 40.21 4.758 ;
      RECT 39.96 4.561 40.21 4.755 ;
      RECT 40.05 4.46 40.22 4.65 ;
      RECT 39.71 3.245 39.715 3.69 ;
      RECT 39.52 3.245 39.54 3.655 ;
      RECT 39.49 3.245 39.495 3.63 ;
      RECT 40.17 3.552 40.185 3.74 ;
      RECT 40.165 3.537 40.17 3.746 ;
      RECT 40.145 3.51 40.165 3.749 ;
      RECT 40.095 3.477 40.145 3.758 ;
      RECT 40.065 3.457 40.095 3.762 ;
      RECT 40.046 3.445 40.065 3.758 ;
      RECT 39.96 3.417 40.046 3.748 ;
      RECT 39.95 3.392 39.96 3.738 ;
      RECT 39.88 3.36 39.95 3.73 ;
      RECT 39.855 3.32 39.88 3.722 ;
      RECT 39.835 3.302 39.855 3.716 ;
      RECT 39.825 3.292 39.835 3.713 ;
      RECT 39.815 3.285 39.825 3.711 ;
      RECT 39.795 3.272 39.815 3.708 ;
      RECT 39.785 3.262 39.795 3.705 ;
      RECT 39.775 3.255 39.785 3.703 ;
      RECT 39.725 3.247 39.775 3.697 ;
      RECT 39.715 3.245 39.725 3.691 ;
      RECT 39.685 3.245 39.71 3.688 ;
      RECT 39.656 3.245 39.685 3.683 ;
      RECT 39.57 3.245 39.656 3.673 ;
      RECT 39.54 3.245 39.57 3.66 ;
      RECT 39.495 3.245 39.52 3.643 ;
      RECT 39.48 3.245 39.49 3.625 ;
      RECT 39.46 3.252 39.48 3.61 ;
      RECT 39.455 3.267 39.46 3.598 ;
      RECT 39.45 3.272 39.455 3.538 ;
      RECT 39.445 3.277 39.45 3.38 ;
      RECT 39.44 3.28 39.445 3.298 ;
      RECT 39.18 4.57 39.215 4.89 ;
      RECT 39.765 4.755 39.77 4.937 ;
      RECT 39.72 4.637 39.765 4.956 ;
      RECT 39.705 4.614 39.72 4.979 ;
      RECT 39.695 4.604 39.705 4.989 ;
      RECT 39.675 4.599 39.695 5.002 ;
      RECT 39.65 4.597 39.675 5.023 ;
      RECT 39.631 4.596 39.65 5.035 ;
      RECT 39.545 4.593 39.631 5.035 ;
      RECT 39.475 4.588 39.545 5.023 ;
      RECT 39.4 4.584 39.475 4.998 ;
      RECT 39.335 4.58 39.4 4.965 ;
      RECT 39.265 4.577 39.335 4.925 ;
      RECT 39.235 4.573 39.265 4.9 ;
      RECT 39.215 4.571 39.235 4.893 ;
      RECT 39.131 4.569 39.18 4.891 ;
      RECT 39.045 4.566 39.131 4.892 ;
      RECT 38.97 4.565 39.045 4.894 ;
      RECT 38.885 4.565 38.97 4.92 ;
      RECT 38.808 4.566 38.885 4.945 ;
      RECT 38.722 4.567 38.808 4.945 ;
      RECT 38.636 4.567 38.722 4.945 ;
      RECT 38.55 4.568 38.636 4.945 ;
      RECT 38.53 4.569 38.55 4.937 ;
      RECT 38.515 4.575 38.53 4.922 ;
      RECT 38.48 4.595 38.515 4.902 ;
      RECT 38.47 4.615 38.48 4.884 ;
      RECT 39.44 3.92 39.445 4.19 ;
      RECT 39.435 3.911 39.44 4.195 ;
      RECT 39.425 3.901 39.435 4.207 ;
      RECT 39.42 3.89 39.425 4.218 ;
      RECT 39.4 3.884 39.42 4.236 ;
      RECT 39.355 3.881 39.4 4.285 ;
      RECT 39.34 3.88 39.355 4.33 ;
      RECT 39.335 3.88 39.34 4.343 ;
      RECT 39.325 3.88 39.335 4.355 ;
      RECT 39.32 3.881 39.325 4.37 ;
      RECT 39.3 3.889 39.32 4.375 ;
      RECT 39.27 3.905 39.3 4.375 ;
      RECT 39.26 3.917 39.265 4.375 ;
      RECT 39.225 3.932 39.26 4.375 ;
      RECT 39.195 3.952 39.225 4.375 ;
      RECT 39.185 3.977 39.195 4.375 ;
      RECT 39.18 4.005 39.185 4.375 ;
      RECT 39.175 4.035 39.18 4.375 ;
      RECT 39.17 4.052 39.175 4.375 ;
      RECT 39.16 4.08 39.17 4.375 ;
      RECT 39.15 4.115 39.16 4.375 ;
      RECT 39.145 4.15 39.15 4.375 ;
      RECT 39.265 3.915 39.27 4.375 ;
      RECT 38.445 3.975 38.965 4.19 ;
      RECT 38.525 3.915 38.965 4.19 ;
      RECT 38.255 3.245 38.26 3.644 ;
      RECT 38 3.245 38.035 3.642 ;
      RECT 37.595 3.28 37.6 3.636 ;
      RECT 38.34 3.283 38.345 3.538 ;
      RECT 38.335 3.281 38.34 3.544 ;
      RECT 38.33 3.28 38.335 3.551 ;
      RECT 38.305 3.273 38.33 3.575 ;
      RECT 38.3 3.266 38.305 3.599 ;
      RECT 38.295 3.262 38.3 3.608 ;
      RECT 38.285 3.257 38.295 3.621 ;
      RECT 38.28 3.254 38.285 3.63 ;
      RECT 38.275 3.252 38.28 3.635 ;
      RECT 38.26 3.248 38.275 3.645 ;
      RECT 38.245 3.242 38.255 3.644 ;
      RECT 38.207 3.24 38.245 3.644 ;
      RECT 38.121 3.242 38.207 3.644 ;
      RECT 38.035 3.244 38.121 3.643 ;
      RECT 37.964 3.245 38 3.642 ;
      RECT 37.878 3.247 37.964 3.642 ;
      RECT 37.792 3.249 37.878 3.641 ;
      RECT 37.706 3.251 37.792 3.641 ;
      RECT 37.62 3.254 37.706 3.64 ;
      RECT 37.61 3.26 37.62 3.639 ;
      RECT 37.6 3.272 37.61 3.637 ;
      RECT 37.54 3.307 37.595 3.633 ;
      RECT 37.535 3.337 37.54 3.395 ;
      RECT 37.88 4.552 37.885 4.809 ;
      RECT 37.86 4.471 37.88 4.826 ;
      RECT 37.84 4.465 37.86 4.855 ;
      RECT 37.78 4.452 37.84 4.875 ;
      RECT 37.735 4.436 37.78 4.876 ;
      RECT 37.651 4.424 37.735 4.864 ;
      RECT 37.565 4.411 37.651 4.848 ;
      RECT 37.555 4.404 37.565 4.84 ;
      RECT 37.51 4.401 37.555 4.78 ;
      RECT 37.49 4.397 37.51 4.695 ;
      RECT 37.475 4.395 37.49 4.648 ;
      RECT 37.445 4.392 37.475 4.618 ;
      RECT 37.41 4.388 37.445 4.595 ;
      RECT 37.367 4.383 37.41 4.583 ;
      RECT 37.281 4.374 37.367 4.592 ;
      RECT 37.195 4.363 37.281 4.604 ;
      RECT 37.13 4.354 37.195 4.613 ;
      RECT 37.11 4.345 37.13 4.618 ;
      RECT 37.105 4.338 37.11 4.62 ;
      RECT 37.065 4.323 37.105 4.617 ;
      RECT 37.045 4.302 37.065 4.612 ;
      RECT 37.03 4.29 37.045 4.605 ;
      RECT 37.025 4.282 37.03 4.598 ;
      RECT 37.01 4.262 37.025 4.591 ;
      RECT 37.005 4.125 37.01 4.585 ;
      RECT 36.925 4.014 37.005 4.557 ;
      RECT 36.916 4.007 36.925 4.523 ;
      RECT 36.83 4.001 36.916 4.448 ;
      RECT 36.805 3.992 36.83 4.36 ;
      RECT 36.775 3.987 36.805 4.335 ;
      RECT 36.71 3.996 36.775 4.32 ;
      RECT 36.69 4.012 36.71 4.295 ;
      RECT 36.68 4.018 36.69 4.243 ;
      RECT 36.66 4.04 36.68 4.125 ;
      RECT 37.315 4.005 37.485 4.19 ;
      RECT 37.315 4.005 37.52 4.188 ;
      RECT 37.365 3.915 37.535 4.179 ;
      RECT 37.315 4.072 37.54 4.172 ;
      RECT 37.33 3.95 37.535 4.179 ;
      RECT 36.53 4.683 36.595 5.126 ;
      RECT 36.47 4.708 36.595 5.124 ;
      RECT 36.47 4.708 36.65 5.118 ;
      RECT 36.455 4.733 36.65 5.117 ;
      RECT 36.595 4.67 36.67 5.114 ;
      RECT 36.53 4.695 36.75 5.108 ;
      RECT 36.455 4.734 36.795 5.102 ;
      RECT 36.44 4.761 36.795 5.093 ;
      RECT 36.455 4.754 36.815 5.085 ;
      RECT 36.44 4.763 36.82 5.068 ;
      RECT 36.435 4.78 36.82 4.895 ;
      RECT 36.44 3.502 36.475 3.74 ;
      RECT 36.44 3.502 36.505 3.739 ;
      RECT 36.44 3.502 36.62 3.735 ;
      RECT 36.44 3.502 36.675 3.713 ;
      RECT 36.45 3.445 36.73 3.613 ;
      RECT 36.555 3.285 36.585 3.736 ;
      RECT 36.585 3.28 36.765 3.493 ;
      RECT 36.455 3.421 36.765 3.493 ;
      RECT 36.505 3.317 36.555 3.737 ;
      RECT 36.475 3.373 36.765 3.493 ;
      RECT 35.335 7.455 35.505 8.925 ;
      RECT 35.335 7.455 35.51 8.715 ;
      RECT 34.965 9.405 35.435 9.575 ;
      RECT 34.965 8.385 35.135 9.575 ;
      RECT 34.96 3.035 35.13 4.225 ;
      RECT 34.96 3.035 35.43 3.205 ;
      RECT 34.345 3.895 34.52 5.155 ;
      RECT 34.345 3.685 34.515 5.155 ;
      RECT 34.345 7.455 34.515 8.925 ;
      RECT 34.345 7.455 34.52 8.715 ;
      RECT 33.975 3.035 34.145 4.225 ;
      RECT 33.975 3.035 34.445 3.205 ;
      RECT 33.975 9.405 34.445 9.575 ;
      RECT 33.975 8.385 34.145 9.575 ;
      RECT 32.985 4.015 33.16 5.155 ;
      RECT 32.985 1.865 33.155 5.155 ;
      RECT 32.985 1.865 33.16 2.415 ;
      RECT 32.985 10.195 33.16 10.745 ;
      RECT 32.985 7.455 33.155 10.745 ;
      RECT 32.985 7.455 33.16 8.595 ;
      RECT 32.555 3.895 32.73 5.155 ;
      RECT 32.555 2.945 32.725 5.155 ;
      RECT 32.555 7.455 32.725 9.665 ;
      RECT 32.555 7.455 32.73 8.715 ;
      RECT 32.125 3.925 32.295 5.155 ;
      RECT 32.185 2.145 32.355 4.095 ;
      RECT 32.125 1.865 32.295 2.315 ;
      RECT 32.125 10.295 32.295 10.745 ;
      RECT 32.185 8.515 32.355 10.465 ;
      RECT 32.125 7.455 32.295 8.685 ;
      RECT 31.6 3.895 31.775 5.155 ;
      RECT 31.6 1.865 31.77 5.155 ;
      RECT 31.6 3.365 32.01 3.695 ;
      RECT 31.6 2.525 32.01 2.855 ;
      RECT 31.6 1.865 31.775 2.355 ;
      RECT 31.6 10.255 31.775 10.745 ;
      RECT 31.6 7.455 31.77 10.745 ;
      RECT 31.6 9.755 32.01 10.085 ;
      RECT 31.6 8.915 32.01 9.245 ;
      RECT 31.6 7.455 31.775 8.715 ;
      RECT 29.715 4.687 29.73 4.738 ;
      RECT 29.71 4.667 29.715 4.785 ;
      RECT 29.695 4.657 29.71 4.853 ;
      RECT 29.67 4.637 29.695 4.908 ;
      RECT 29.63 4.622 29.67 4.928 ;
      RECT 29.585 4.616 29.63 4.956 ;
      RECT 29.515 4.606 29.585 4.973 ;
      RECT 29.495 4.598 29.515 4.973 ;
      RECT 29.435 4.592 29.495 4.965 ;
      RECT 29.376 4.583 29.435 4.953 ;
      RECT 29.29 4.572 29.376 4.936 ;
      RECT 29.268 4.563 29.29 4.924 ;
      RECT 29.182 4.556 29.268 4.911 ;
      RECT 29.096 4.543 29.182 4.892 ;
      RECT 29.01 4.531 29.096 4.872 ;
      RECT 28.98 4.52 29.01 4.859 ;
      RECT 28.93 4.506 28.98 4.851 ;
      RECT 28.91 4.495 28.93 4.843 ;
      RECT 28.861 4.484 28.91 4.835 ;
      RECT 28.775 4.463 28.861 4.82 ;
      RECT 28.73 4.45 28.775 4.805 ;
      RECT 28.685 4.45 28.73 4.785 ;
      RECT 28.63 4.45 28.685 4.72 ;
      RECT 28.605 4.45 28.63 4.643 ;
      RECT 29.13 4.187 29.3 4.37 ;
      RECT 29.13 4.187 29.315 4.328 ;
      RECT 29.13 4.187 29.32 4.27 ;
      RECT 29.19 3.955 29.325 4.246 ;
      RECT 29.19 3.959 29.33 4.229 ;
      RECT 29.135 4.122 29.33 4.229 ;
      RECT 29.16 3.967 29.3 4.37 ;
      RECT 29.16 3.971 29.34 4.17 ;
      RECT 29.145 4.057 29.34 4.17 ;
      RECT 29.155 3.987 29.3 4.37 ;
      RECT 29.155 3.99 29.35 4.083 ;
      RECT 29.15 4.007 29.35 4.083 ;
      RECT 28.92 3.227 29.09 3.71 ;
      RECT 28.915 3.222 29.065 3.7 ;
      RECT 28.915 3.229 29.095 3.694 ;
      RECT 28.905 3.223 29.065 3.673 ;
      RECT 28.905 3.239 29.11 3.632 ;
      RECT 28.875 3.224 29.065 3.595 ;
      RECT 28.875 3.254 29.12 3.535 ;
      RECT 28.87 3.226 29.065 3.533 ;
      RECT 28.85 3.235 29.095 3.49 ;
      RECT 28.825 3.251 29.11 3.402 ;
      RECT 28.825 3.27 29.135 3.393 ;
      RECT 28.82 3.307 29.135 3.345 ;
      RECT 28.825 3.287 29.14 3.313 ;
      RECT 28.92 3.221 29.03 3.71 ;
      RECT 29.006 3.22 29.03 3.71 ;
      RECT 28.24 4.005 28.245 4.216 ;
      RECT 28.84 4.005 28.845 4.19 ;
      RECT 28.905 4.045 28.91 4.158 ;
      RECT 28.9 4.037 28.905 4.164 ;
      RECT 28.895 4.027 28.9 4.172 ;
      RECT 28.89 4.017 28.895 4.181 ;
      RECT 28.885 4.007 28.89 4.185 ;
      RECT 28.845 4.005 28.885 4.188 ;
      RECT 28.817 4.004 28.84 4.192 ;
      RECT 28.731 4.001 28.817 4.199 ;
      RECT 28.645 3.997 28.731 4.21 ;
      RECT 28.625 3.995 28.645 4.216 ;
      RECT 28.607 3.994 28.625 4.219 ;
      RECT 28.521 3.992 28.607 4.226 ;
      RECT 28.435 3.987 28.521 4.239 ;
      RECT 28.416 3.984 28.435 4.244 ;
      RECT 28.33 3.982 28.416 4.235 ;
      RECT 28.32 3.982 28.33 4.228 ;
      RECT 28.245 3.995 28.32 4.222 ;
      RECT 28.23 4.006 28.24 4.216 ;
      RECT 28.22 4.008 28.23 4.215 ;
      RECT 28.21 4.012 28.22 4.211 ;
      RECT 28.205 4.015 28.21 4.205 ;
      RECT 28.195 4.017 28.205 4.199 ;
      RECT 28.19 4.02 28.195 4.193 ;
      RECT 28.225 10.195 28.4 10.745 ;
      RECT 28.225 7.455 28.395 10.745 ;
      RECT 28.225 7.455 28.4 8.595 ;
      RECT 28.17 4.606 28.175 4.81 ;
      RECT 28.155 4.593 28.17 4.903 ;
      RECT 28.14 4.574 28.155 5.18 ;
      RECT 28.105 4.54 28.14 5.18 ;
      RECT 28.101 4.51 28.105 5.18 ;
      RECT 28.015 4.392 28.101 5.18 ;
      RECT 28.005 4.267 28.015 5.18 ;
      RECT 27.99 4.235 28.005 5.18 ;
      RECT 27.985 4.21 27.99 5.18 ;
      RECT 27.98 4.2 27.985 5.136 ;
      RECT 27.965 4.172 27.98 5.041 ;
      RECT 27.95 4.138 27.965 4.94 ;
      RECT 27.945 4.116 27.95 4.893 ;
      RECT 27.94 4.105 27.945 4.863 ;
      RECT 27.935 4.095 27.94 4.829 ;
      RECT 27.925 4.082 27.935 4.797 ;
      RECT 27.9 4.058 27.925 4.723 ;
      RECT 27.895 4.038 27.9 4.648 ;
      RECT 27.89 4.032 27.895 4.623 ;
      RECT 27.885 4.027 27.89 4.588 ;
      RECT 27.88 4.022 27.885 4.563 ;
      RECT 27.875 4.02 27.88 4.543 ;
      RECT 27.87 4.02 27.875 4.528 ;
      RECT 27.865 4.02 27.87 4.488 ;
      RECT 27.855 4.02 27.865 4.46 ;
      RECT 27.845 4.02 27.855 4.405 ;
      RECT 27.83 4.02 27.845 4.343 ;
      RECT 27.825 4.019 27.83 4.288 ;
      RECT 27.81 4.018 27.825 4.268 ;
      RECT 27.75 4.016 27.81 4.242 ;
      RECT 27.715 4.017 27.75 4.222 ;
      RECT 27.71 4.019 27.715 4.212 ;
      RECT 27.7 4.038 27.71 4.202 ;
      RECT 27.695 4.065 27.7 4.133 ;
      RECT 27.81 3.49 27.98 3.735 ;
      RECT 27.845 3.261 27.98 3.735 ;
      RECT 27.845 3.263 27.99 3.73 ;
      RECT 27.845 3.265 28.015 3.718 ;
      RECT 27.845 3.268 28.04 3.7 ;
      RECT 27.845 3.273 28.09 3.673 ;
      RECT 27.845 3.278 28.11 3.638 ;
      RECT 27.825 3.28 28.12 3.613 ;
      RECT 27.815 3.375 28.12 3.613 ;
      RECT 27.845 3.26 27.955 3.735 ;
      RECT 27.855 3.257 27.95 3.735 ;
      RECT 27.795 7.455 27.965 9.665 ;
      RECT 27.795 7.455 27.97 8.715 ;
      RECT 27.375 4.522 27.565 4.88 ;
      RECT 27.375 4.534 27.6 4.879 ;
      RECT 27.375 4.562 27.62 4.877 ;
      RECT 27.375 4.587 27.625 4.876 ;
      RECT 27.375 4.645 27.64 4.875 ;
      RECT 27.36 4.518 27.52 4.86 ;
      RECT 27.34 4.527 27.565 4.813 ;
      RECT 27.315 4.538 27.6 4.75 ;
      RECT 27.315 4.622 27.635 4.75 ;
      RECT 27.315 4.597 27.63 4.75 ;
      RECT 27.375 4.513 27.52 4.88 ;
      RECT 27.461 4.512 27.52 4.88 ;
      RECT 27.461 4.511 27.505 4.88 ;
      RECT 26.84 10.255 27.015 10.745 ;
      RECT 26.84 7.455 27.01 10.745 ;
      RECT 26.84 9.755 27.25 10.085 ;
      RECT 26.84 8.915 27.25 9.245 ;
      RECT 26.84 7.455 27.015 8.715 ;
      RECT 27.16 4.027 27.165 4.405 ;
      RECT 27.155 3.995 27.16 4.405 ;
      RECT 27.15 3.967 27.155 4.405 ;
      RECT 27.145 3.947 27.15 4.405 ;
      RECT 27.09 3.93 27.145 4.405 ;
      RECT 27.05 3.915 27.09 4.405 ;
      RECT 26.995 3.902 27.05 4.405 ;
      RECT 26.96 3.893 26.995 4.405 ;
      RECT 26.956 3.891 26.96 4.404 ;
      RECT 26.87 3.887 26.956 4.387 ;
      RECT 26.785 3.879 26.87 4.35 ;
      RECT 26.775 3.875 26.785 4.323 ;
      RECT 26.765 3.875 26.775 4.305 ;
      RECT 26.755 3.877 26.765 4.288 ;
      RECT 26.75 3.882 26.755 4.274 ;
      RECT 26.745 3.886 26.75 4.261 ;
      RECT 26.735 3.891 26.745 4.245 ;
      RECT 26.72 3.905 26.735 4.22 ;
      RECT 26.715 3.911 26.72 4.2 ;
      RECT 26.71 3.913 26.715 4.193 ;
      RECT 26.705 3.917 26.71 4.068 ;
      RECT 26.885 4.717 27.13 5.18 ;
      RECT 26.805 4.69 27.125 5.176 ;
      RECT 26.735 4.725 27.13 5.169 ;
      RECT 26.525 4.98 27.13 5.165 ;
      RECT 26.705 4.748 27.13 5.165 ;
      RECT 26.545 4.94 27.13 5.165 ;
      RECT 26.695 4.76 27.13 5.165 ;
      RECT 26.58 4.877 27.13 5.165 ;
      RECT 26.635 4.802 27.13 5.165 ;
      RECT 26.885 4.667 27.125 5.18 ;
      RECT 26.915 4.66 27.125 5.18 ;
      RECT 26.905 4.662 27.125 5.18 ;
      RECT 26.915 4.657 27.045 5.18 ;
      RECT 26.47 3.22 26.556 3.659 ;
      RECT 26.465 3.22 26.556 3.657 ;
      RECT 26.465 3.22 26.625 3.656 ;
      RECT 26.465 3.22 26.655 3.653 ;
      RECT 26.45 3.227 26.655 3.644 ;
      RECT 26.45 3.227 26.66 3.64 ;
      RECT 26.445 3.237 26.66 3.633 ;
      RECT 26.44 3.242 26.66 3.608 ;
      RECT 26.44 3.242 26.675 3.59 ;
      RECT 26.465 3.22 26.695 3.505 ;
      RECT 26.435 3.247 26.695 3.503 ;
      RECT 26.445 3.24 26.7 3.441 ;
      RECT 26.435 3.362 26.705 3.424 ;
      RECT 26.42 3.257 26.7 3.375 ;
      RECT 26.415 3.267 26.7 3.275 ;
      RECT 26.495 4.038 26.5 4.115 ;
      RECT 26.485 4.032 26.495 4.305 ;
      RECT 26.475 4.024 26.485 4.326 ;
      RECT 26.465 4.015 26.475 4.348 ;
      RECT 26.46 4.01 26.465 4.365 ;
      RECT 26.42 4.01 26.46 4.405 ;
      RECT 26.4 4.01 26.42 4.46 ;
      RECT 26.395 4.01 26.4 4.488 ;
      RECT 26.385 4.01 26.395 4.503 ;
      RECT 26.35 4.01 26.385 4.545 ;
      RECT 26.345 4.01 26.35 4.588 ;
      RECT 26.335 4.01 26.345 4.603 ;
      RECT 26.32 4.01 26.335 4.623 ;
      RECT 26.305 4.01 26.32 4.65 ;
      RECT 26.3 4.011 26.305 4.668 ;
      RECT 26.28 4.012 26.3 4.675 ;
      RECT 26.225 4.013 26.28 4.695 ;
      RECT 26.215 4.014 26.225 4.709 ;
      RECT 26.21 4.017 26.215 4.708 ;
      RECT 26.17 4.09 26.21 4.706 ;
      RECT 26.155 4.17 26.17 4.704 ;
      RECT 26.13 4.225 26.155 4.702 ;
      RECT 26.115 4.29 26.13 4.701 ;
      RECT 26.07 4.322 26.115 4.698 ;
      RECT 25.985 4.345 26.07 4.693 ;
      RECT 25.96 4.365 25.985 4.688 ;
      RECT 25.89 4.37 25.96 4.684 ;
      RECT 25.87 4.372 25.89 4.681 ;
      RECT 25.785 4.383 25.87 4.675 ;
      RECT 25.78 4.394 25.785 4.67 ;
      RECT 25.77 4.396 25.78 4.67 ;
      RECT 25.735 4.4 25.77 4.668 ;
      RECT 25.685 4.41 25.735 4.655 ;
      RECT 25.665 4.418 25.685 4.64 ;
      RECT 25.585 4.43 25.665 4.623 ;
      RECT 25.75 3.98 25.92 4.19 ;
      RECT 25.866 3.976 25.92 4.19 ;
      RECT 25.671 3.98 25.92 4.181 ;
      RECT 25.671 3.98 25.925 4.17 ;
      RECT 25.585 3.98 25.925 4.161 ;
      RECT 25.585 3.988 25.935 4.105 ;
      RECT 25.585 4 25.94 4.018 ;
      RECT 25.585 4.007 25.945 4.01 ;
      RECT 25.78 3.978 25.92 4.19 ;
      RECT 25.535 4.923 25.78 5.255 ;
      RECT 25.53 4.915 25.535 5.252 ;
      RECT 25.5 4.935 25.78 5.233 ;
      RECT 25.48 4.967 25.78 5.206 ;
      RECT 25.53 4.92 25.707 5.252 ;
      RECT 25.53 4.917 25.621 5.252 ;
      RECT 25.47 3.265 25.64 3.685 ;
      RECT 25.465 3.265 25.64 3.683 ;
      RECT 25.465 3.265 25.665 3.673 ;
      RECT 25.465 3.265 25.685 3.648 ;
      RECT 25.46 3.265 25.685 3.643 ;
      RECT 25.46 3.265 25.695 3.633 ;
      RECT 25.46 3.265 25.7 3.628 ;
      RECT 25.46 3.27 25.705 3.623 ;
      RECT 25.46 3.302 25.72 3.613 ;
      RECT 25.46 3.372 25.745 3.596 ;
      RECT 25.44 3.372 25.745 3.588 ;
      RECT 25.44 3.432 25.755 3.565 ;
      RECT 25.44 3.472 25.765 3.51 ;
      RECT 25.425 3.265 25.7 3.49 ;
      RECT 25.415 3.28 25.705 3.388 ;
      RECT 25.005 4.67 25.175 5.195 ;
      RECT 25 4.67 25.175 5.188 ;
      RECT 24.99 4.67 25.18 5.153 ;
      RECT 24.985 4.68 25.18 5.125 ;
      RECT 24.98 4.7 25.18 5.108 ;
      RECT 24.99 4.675 25.185 5.098 ;
      RECT 24.975 4.72 25.185 5.09 ;
      RECT 24.97 4.74 25.185 5.075 ;
      RECT 24.965 4.77 25.185 5.065 ;
      RECT 24.955 4.815 25.185 5.04 ;
      RECT 24.985 4.685 25.19 5.023 ;
      RECT 24.95 4.867 25.19 5.018 ;
      RECT 24.985 4.695 25.195 4.988 ;
      RECT 24.945 4.9 25.195 4.985 ;
      RECT 24.94 4.925 25.195 4.965 ;
      RECT 24.98 4.712 25.205 4.905 ;
      RECT 24.975 4.734 25.215 4.798 ;
      RECT 24.925 3.981 24.94 4.25 ;
      RECT 24.88 3.965 24.925 4.295 ;
      RECT 24.875 3.953 24.88 4.345 ;
      RECT 24.865 3.949 24.875 4.378 ;
      RECT 24.86 3.946 24.865 4.406 ;
      RECT 24.845 3.948 24.86 4.448 ;
      RECT 24.84 3.952 24.845 4.488 ;
      RECT 24.82 3.957 24.84 4.54 ;
      RECT 24.816 3.962 24.82 4.597 ;
      RECT 24.73 3.981 24.816 4.634 ;
      RECT 24.72 4.002 24.73 4.67 ;
      RECT 24.715 4.01 24.72 4.671 ;
      RECT 24.71 4.052 24.715 4.672 ;
      RECT 24.695 4.14 24.71 4.673 ;
      RECT 24.685 4.29 24.695 4.675 ;
      RECT 24.68 4.335 24.685 4.677 ;
      RECT 24.645 4.377 24.68 4.68 ;
      RECT 24.64 4.395 24.645 4.683 ;
      RECT 24.563 4.401 24.64 4.689 ;
      RECT 24.477 4.415 24.563 4.702 ;
      RECT 24.391 4.429 24.477 4.716 ;
      RECT 24.305 4.443 24.391 4.729 ;
      RECT 24.245 4.455 24.305 4.741 ;
      RECT 24.22 4.462 24.245 4.748 ;
      RECT 24.206 4.465 24.22 4.753 ;
      RECT 24.12 4.473 24.206 4.769 ;
      RECT 24.115 4.48 24.12 4.784 ;
      RECT 24.091 4.48 24.115 4.791 ;
      RECT 24.005 4.483 24.091 4.819 ;
      RECT 23.92 4.487 24.005 4.863 ;
      RECT 23.855 4.491 23.92 4.9 ;
      RECT 23.83 4.494 23.855 4.916 ;
      RECT 23.755 4.507 23.83 4.92 ;
      RECT 23.73 4.525 23.755 4.924 ;
      RECT 23.72 4.532 23.73 4.926 ;
      RECT 23.705 4.535 23.72 4.927 ;
      RECT 23.645 4.547 23.705 4.931 ;
      RECT 23.635 4.561 23.645 4.935 ;
      RECT 23.58 4.571 23.635 4.923 ;
      RECT 23.555 4.592 23.58 4.906 ;
      RECT 23.535 4.612 23.555 4.897 ;
      RECT 23.53 4.625 23.535 4.892 ;
      RECT 23.515 4.637 23.53 4.888 ;
      RECT 24.75 3.292 24.755 3.315 ;
      RECT 24.745 3.283 24.75 3.355 ;
      RECT 24.74 3.281 24.745 3.398 ;
      RECT 24.735 3.272 24.74 3.433 ;
      RECT 24.73 3.262 24.735 3.505 ;
      RECT 24.725 3.252 24.73 3.57 ;
      RECT 24.72 3.249 24.725 3.61 ;
      RECT 24.695 3.243 24.72 3.7 ;
      RECT 24.66 3.231 24.695 3.725 ;
      RECT 24.65 3.222 24.66 3.725 ;
      RECT 24.515 3.22 24.525 3.708 ;
      RECT 24.505 3.22 24.515 3.675 ;
      RECT 24.5 3.22 24.505 3.65 ;
      RECT 24.495 3.22 24.5 3.638 ;
      RECT 24.49 3.22 24.495 3.62 ;
      RECT 24.48 3.22 24.49 3.585 ;
      RECT 24.475 3.222 24.48 3.563 ;
      RECT 24.47 3.228 24.475 3.548 ;
      RECT 24.465 3.234 24.47 3.533 ;
      RECT 24.45 3.246 24.465 3.506 ;
      RECT 24.445 3.257 24.45 3.474 ;
      RECT 24.44 3.267 24.445 3.458 ;
      RECT 24.43 3.275 24.44 3.427 ;
      RECT 24.425 3.285 24.43 3.401 ;
      RECT 24.42 3.342 24.425 3.384 ;
      RECT 24.525 3.22 24.65 3.725 ;
      RECT 24.24 3.907 24.5 4.205 ;
      RECT 24.235 3.914 24.5 4.203 ;
      RECT 24.24 3.909 24.515 4.198 ;
      RECT 24.23 3.922 24.515 4.195 ;
      RECT 24.23 3.927 24.52 4.188 ;
      RECT 24.225 3.935 24.52 4.185 ;
      RECT 24.225 3.952 24.525 3.983 ;
      RECT 24.24 3.904 24.471 4.205 ;
      RECT 24.295 3.903 24.471 4.205 ;
      RECT 24.295 3.9 24.385 4.205 ;
      RECT 24.295 3.897 24.381 4.205 ;
      RECT 23.985 4.17 23.99 4.183 ;
      RECT 23.98 4.137 23.985 4.188 ;
      RECT 23.975 4.092 23.98 4.195 ;
      RECT 23.97 4.047 23.975 4.203 ;
      RECT 23.965 4.015 23.97 4.211 ;
      RECT 23.96 3.975 23.965 4.212 ;
      RECT 23.945 3.955 23.96 4.214 ;
      RECT 23.87 3.937 23.945 4.226 ;
      RECT 23.86 3.93 23.87 4.237 ;
      RECT 23.855 3.93 23.86 4.239 ;
      RECT 23.825 3.936 23.855 4.243 ;
      RECT 23.785 3.949 23.825 4.243 ;
      RECT 23.76 3.96 23.785 4.229 ;
      RECT 23.745 3.966 23.76 4.212 ;
      RECT 23.735 3.968 23.745 4.203 ;
      RECT 23.73 3.969 23.735 4.198 ;
      RECT 23.725 3.97 23.73 4.193 ;
      RECT 23.72 3.971 23.725 4.19 ;
      RECT 23.695 3.976 23.72 4.18 ;
      RECT 23.685 3.992 23.695 4.167 ;
      RECT 23.68 4.012 23.685 4.162 ;
      RECT 23.69 3.405 23.695 3.601 ;
      RECT 23.675 3.369 23.69 3.603 ;
      RECT 23.665 3.351 23.675 3.608 ;
      RECT 23.655 3.337 23.665 3.612 ;
      RECT 23.61 3.321 23.655 3.622 ;
      RECT 23.605 3.311 23.61 3.631 ;
      RECT 23.56 3.3 23.605 3.637 ;
      RECT 23.555 3.288 23.56 3.644 ;
      RECT 23.54 3.283 23.555 3.648 ;
      RECT 23.525 3.275 23.54 3.653 ;
      RECT 23.515 3.268 23.525 3.658 ;
      RECT 23.505 3.265 23.515 3.663 ;
      RECT 23.495 3.265 23.505 3.664 ;
      RECT 23.49 3.262 23.495 3.663 ;
      RECT 23.455 3.257 23.48 3.662 ;
      RECT 23.431 3.253 23.455 3.661 ;
      RECT 23.345 3.244 23.431 3.658 ;
      RECT 23.33 3.236 23.345 3.655 ;
      RECT 23.308 3.235 23.33 3.654 ;
      RECT 23.222 3.235 23.308 3.652 ;
      RECT 23.136 3.235 23.222 3.65 ;
      RECT 23.05 3.235 23.136 3.647 ;
      RECT 23.04 3.235 23.05 3.638 ;
      RECT 23.01 3.235 23.04 3.598 ;
      RECT 23 3.245 23.01 3.553 ;
      RECT 22.995 3.285 23 3.538 ;
      RECT 22.99 3.3 22.995 3.525 ;
      RECT 22.96 3.38 22.99 3.487 ;
      RECT 23.48 3.26 23.49 3.663 ;
      RECT 23.305 4.025 23.32 4.63 ;
      RECT 23.31 4.02 23.32 4.63 ;
      RECT 23.475 4.02 23.48 4.203 ;
      RECT 23.465 4.02 23.475 4.233 ;
      RECT 23.45 4.02 23.465 4.293 ;
      RECT 23.445 4.02 23.45 4.338 ;
      RECT 23.44 4.02 23.445 4.368 ;
      RECT 23.435 4.02 23.44 4.388 ;
      RECT 23.425 4.02 23.435 4.423 ;
      RECT 23.41 4.02 23.425 4.455 ;
      RECT 23.365 4.02 23.41 4.483 ;
      RECT 23.36 4.02 23.365 4.513 ;
      RECT 23.355 4.02 23.36 4.525 ;
      RECT 23.35 4.02 23.355 4.533 ;
      RECT 23.34 4.02 23.35 4.548 ;
      RECT 23.335 4.02 23.34 4.57 ;
      RECT 23.325 4.02 23.335 4.593 ;
      RECT 23.32 4.02 23.325 4.613 ;
      RECT 23.285 4.035 23.305 4.63 ;
      RECT 23.26 4.052 23.285 4.63 ;
      RECT 23.255 4.062 23.26 4.63 ;
      RECT 23.225 4.077 23.255 4.63 ;
      RECT 23.15 4.119 23.225 4.63 ;
      RECT 23.145 4.15 23.15 4.613 ;
      RECT 23.14 4.154 23.145 4.595 ;
      RECT 23.135 4.158 23.14 4.558 ;
      RECT 23.13 4.342 23.135 4.525 ;
      RECT 22.615 4.531 22.701 5.096 ;
      RECT 22.57 4.533 22.735 5.09 ;
      RECT 22.701 4.53 22.735 5.09 ;
      RECT 22.615 4.532 22.82 5.084 ;
      RECT 22.57 4.542 22.83 5.08 ;
      RECT 22.545 4.534 22.82 5.076 ;
      RECT 22.54 4.537 22.82 5.071 ;
      RECT 22.515 4.552 22.83 5.065 ;
      RECT 22.515 4.577 22.87 5.06 ;
      RECT 22.475 4.585 22.87 5.035 ;
      RECT 22.475 4.612 22.885 5.033 ;
      RECT 22.475 4.642 22.895 5.02 ;
      RECT 22.47 4.787 22.895 5.008 ;
      RECT 22.475 4.716 22.915 5.005 ;
      RECT 22.475 4.773 22.92 4.813 ;
      RECT 22.665 4.052 22.835 4.23 ;
      RECT 22.615 3.991 22.665 4.215 ;
      RECT 22.35 3.971 22.615 4.2 ;
      RECT 22.31 4.035 22.785 4.2 ;
      RECT 22.31 4.025 22.74 4.2 ;
      RECT 22.31 4.022 22.73 4.2 ;
      RECT 22.31 4.01 22.72 4.2 ;
      RECT 22.31 3.995 22.665 4.2 ;
      RECT 22.35 3.967 22.551 4.2 ;
      RECT 22.36 3.945 22.551 4.2 ;
      RECT 22.385 3.93 22.465 4.2 ;
      RECT 22.14 4.46 22.26 4.905 ;
      RECT 22.125 4.46 22.26 4.904 ;
      RECT 22.08 4.482 22.26 4.899 ;
      RECT 22.04 4.531 22.26 4.893 ;
      RECT 22.04 4.531 22.265 4.868 ;
      RECT 22.04 4.531 22.285 4.758 ;
      RECT 22.035 4.561 22.285 4.755 ;
      RECT 22.125 4.46 22.295 4.65 ;
      RECT 21.785 3.245 21.79 3.69 ;
      RECT 21.595 3.245 21.615 3.655 ;
      RECT 21.565 3.245 21.57 3.63 ;
      RECT 22.245 3.552 22.26 3.74 ;
      RECT 22.24 3.537 22.245 3.746 ;
      RECT 22.22 3.51 22.24 3.749 ;
      RECT 22.17 3.477 22.22 3.758 ;
      RECT 22.14 3.457 22.17 3.762 ;
      RECT 22.121 3.445 22.14 3.758 ;
      RECT 22.035 3.417 22.121 3.748 ;
      RECT 22.025 3.392 22.035 3.738 ;
      RECT 21.955 3.36 22.025 3.73 ;
      RECT 21.93 3.32 21.955 3.722 ;
      RECT 21.91 3.302 21.93 3.716 ;
      RECT 21.9 3.292 21.91 3.713 ;
      RECT 21.89 3.285 21.9 3.711 ;
      RECT 21.87 3.272 21.89 3.708 ;
      RECT 21.86 3.262 21.87 3.705 ;
      RECT 21.85 3.255 21.86 3.703 ;
      RECT 21.8 3.247 21.85 3.697 ;
      RECT 21.79 3.245 21.8 3.691 ;
      RECT 21.76 3.245 21.785 3.688 ;
      RECT 21.731 3.245 21.76 3.683 ;
      RECT 21.645 3.245 21.731 3.673 ;
      RECT 21.615 3.245 21.645 3.66 ;
      RECT 21.57 3.245 21.595 3.643 ;
      RECT 21.555 3.245 21.565 3.625 ;
      RECT 21.535 3.252 21.555 3.61 ;
      RECT 21.53 3.267 21.535 3.598 ;
      RECT 21.525 3.272 21.53 3.538 ;
      RECT 21.52 3.277 21.525 3.38 ;
      RECT 21.515 3.28 21.52 3.298 ;
      RECT 21.255 4.57 21.29 4.89 ;
      RECT 21.84 4.755 21.845 4.937 ;
      RECT 21.795 4.637 21.84 4.956 ;
      RECT 21.78 4.614 21.795 4.979 ;
      RECT 21.77 4.604 21.78 4.989 ;
      RECT 21.75 4.599 21.77 5.002 ;
      RECT 21.725 4.597 21.75 5.023 ;
      RECT 21.706 4.596 21.725 5.035 ;
      RECT 21.62 4.593 21.706 5.035 ;
      RECT 21.55 4.588 21.62 5.023 ;
      RECT 21.475 4.584 21.55 4.998 ;
      RECT 21.41 4.58 21.475 4.965 ;
      RECT 21.34 4.577 21.41 4.925 ;
      RECT 21.31 4.573 21.34 4.9 ;
      RECT 21.29 4.571 21.31 4.893 ;
      RECT 21.206 4.569 21.255 4.891 ;
      RECT 21.12 4.566 21.206 4.892 ;
      RECT 21.045 4.565 21.12 4.894 ;
      RECT 20.96 4.565 21.045 4.92 ;
      RECT 20.883 4.566 20.96 4.945 ;
      RECT 20.797 4.567 20.883 4.945 ;
      RECT 20.711 4.567 20.797 4.945 ;
      RECT 20.625 4.568 20.711 4.945 ;
      RECT 20.605 4.569 20.625 4.937 ;
      RECT 20.59 4.575 20.605 4.922 ;
      RECT 20.555 4.595 20.59 4.902 ;
      RECT 20.545 4.615 20.555 4.884 ;
      RECT 21.515 3.92 21.52 4.19 ;
      RECT 21.51 3.911 21.515 4.195 ;
      RECT 21.5 3.901 21.51 4.207 ;
      RECT 21.495 3.89 21.5 4.218 ;
      RECT 21.475 3.884 21.495 4.236 ;
      RECT 21.43 3.881 21.475 4.285 ;
      RECT 21.415 3.88 21.43 4.33 ;
      RECT 21.41 3.88 21.415 4.343 ;
      RECT 21.4 3.88 21.41 4.355 ;
      RECT 21.395 3.881 21.4 4.37 ;
      RECT 21.375 3.889 21.395 4.375 ;
      RECT 21.345 3.905 21.375 4.375 ;
      RECT 21.335 3.917 21.34 4.375 ;
      RECT 21.3 3.932 21.335 4.375 ;
      RECT 21.27 3.952 21.3 4.375 ;
      RECT 21.26 3.977 21.27 4.375 ;
      RECT 21.255 4.005 21.26 4.375 ;
      RECT 21.25 4.035 21.255 4.375 ;
      RECT 21.245 4.052 21.25 4.375 ;
      RECT 21.235 4.08 21.245 4.375 ;
      RECT 21.225 4.115 21.235 4.375 ;
      RECT 21.22 4.15 21.225 4.375 ;
      RECT 21.34 3.915 21.345 4.375 ;
      RECT 20.52 3.975 21.04 4.19 ;
      RECT 20.6 3.915 21.04 4.19 ;
      RECT 20.33 3.245 20.335 3.644 ;
      RECT 20.075 3.245 20.11 3.642 ;
      RECT 19.67 3.28 19.675 3.636 ;
      RECT 20.415 3.283 20.42 3.538 ;
      RECT 20.41 3.281 20.415 3.544 ;
      RECT 20.405 3.28 20.41 3.551 ;
      RECT 20.38 3.273 20.405 3.575 ;
      RECT 20.375 3.266 20.38 3.599 ;
      RECT 20.37 3.262 20.375 3.608 ;
      RECT 20.36 3.257 20.37 3.621 ;
      RECT 20.355 3.254 20.36 3.63 ;
      RECT 20.35 3.252 20.355 3.635 ;
      RECT 20.335 3.248 20.35 3.645 ;
      RECT 20.32 3.242 20.33 3.644 ;
      RECT 20.282 3.24 20.32 3.644 ;
      RECT 20.196 3.242 20.282 3.644 ;
      RECT 20.11 3.244 20.196 3.643 ;
      RECT 20.039 3.245 20.075 3.642 ;
      RECT 19.953 3.247 20.039 3.642 ;
      RECT 19.867 3.249 19.953 3.641 ;
      RECT 19.781 3.251 19.867 3.641 ;
      RECT 19.695 3.254 19.781 3.64 ;
      RECT 19.685 3.26 19.695 3.639 ;
      RECT 19.675 3.272 19.685 3.637 ;
      RECT 19.615 3.307 19.67 3.633 ;
      RECT 19.61 3.337 19.615 3.395 ;
      RECT 19.955 4.552 19.96 4.809 ;
      RECT 19.935 4.471 19.955 4.826 ;
      RECT 19.915 4.465 19.935 4.855 ;
      RECT 19.855 4.452 19.915 4.875 ;
      RECT 19.81 4.436 19.855 4.876 ;
      RECT 19.726 4.424 19.81 4.864 ;
      RECT 19.64 4.411 19.726 4.848 ;
      RECT 19.63 4.404 19.64 4.84 ;
      RECT 19.585 4.401 19.63 4.78 ;
      RECT 19.565 4.397 19.585 4.695 ;
      RECT 19.55 4.395 19.565 4.648 ;
      RECT 19.52 4.392 19.55 4.618 ;
      RECT 19.485 4.388 19.52 4.595 ;
      RECT 19.442 4.383 19.485 4.583 ;
      RECT 19.356 4.374 19.442 4.592 ;
      RECT 19.27 4.363 19.356 4.604 ;
      RECT 19.205 4.354 19.27 4.613 ;
      RECT 19.185 4.345 19.205 4.618 ;
      RECT 19.18 4.338 19.185 4.62 ;
      RECT 19.14 4.323 19.18 4.617 ;
      RECT 19.12 4.302 19.14 4.612 ;
      RECT 19.105 4.29 19.12 4.605 ;
      RECT 19.1 4.282 19.105 4.598 ;
      RECT 19.085 4.262 19.1 4.591 ;
      RECT 19.08 4.125 19.085 4.585 ;
      RECT 19 4.014 19.08 4.557 ;
      RECT 18.991 4.007 19 4.523 ;
      RECT 18.905 4.001 18.991 4.448 ;
      RECT 18.88 3.992 18.905 4.36 ;
      RECT 18.85 3.987 18.88 4.335 ;
      RECT 18.785 3.996 18.85 4.32 ;
      RECT 18.765 4.012 18.785 4.295 ;
      RECT 18.755 4.018 18.765 4.243 ;
      RECT 18.735 4.04 18.755 4.125 ;
      RECT 19.39 4.005 19.56 4.19 ;
      RECT 19.39 4.005 19.595 4.188 ;
      RECT 19.44 3.915 19.61 4.179 ;
      RECT 19.39 4.072 19.615 4.172 ;
      RECT 19.405 3.95 19.61 4.179 ;
      RECT 18.605 4.683 18.67 5.126 ;
      RECT 18.545 4.708 18.67 5.124 ;
      RECT 18.545 4.708 18.725 5.118 ;
      RECT 18.53 4.733 18.725 5.117 ;
      RECT 18.67 4.67 18.745 5.114 ;
      RECT 18.605 4.695 18.825 5.108 ;
      RECT 18.53 4.734 18.87 5.102 ;
      RECT 18.515 4.761 18.87 5.093 ;
      RECT 18.53 4.754 18.89 5.085 ;
      RECT 18.515 4.763 18.895 5.068 ;
      RECT 18.51 4.78 18.895 4.895 ;
      RECT 18.515 3.502 18.55 3.74 ;
      RECT 18.515 3.502 18.58 3.739 ;
      RECT 18.515 3.502 18.695 3.735 ;
      RECT 18.515 3.502 18.75 3.713 ;
      RECT 18.525 3.445 18.805 3.613 ;
      RECT 18.63 3.285 18.66 3.736 ;
      RECT 18.66 3.28 18.84 3.493 ;
      RECT 18.53 3.421 18.84 3.493 ;
      RECT 18.58 3.317 18.63 3.737 ;
      RECT 18.55 3.373 18.84 3.493 ;
      RECT 16.765 7.455 16.935 9.665 ;
      RECT 16.765 7.455 16.94 8.715 ;
      RECT 16.335 10.295 16.505 10.745 ;
      RECT 16.395 8.515 16.565 10.465 ;
      RECT 16.335 7.455 16.505 8.685 ;
      RECT 15.81 10.255 15.985 10.745 ;
      RECT 15.81 7.455 15.98 10.745 ;
      RECT 15.81 9.755 16.22 10.085 ;
      RECT 15.81 8.915 16.22 9.245 ;
      RECT 15.81 7.455 15.985 8.715 ;
      RECT 107.035 10.235 107.21 10.745 ;
      RECT 106.045 1.865 106.22 2.375 ;
      RECT 106.045 10.235 106.22 10.745 ;
      RECT 104.255 1.865 104.43 2.375 ;
      RECT 104.255 10.235 104.43 10.745 ;
      RECT 99.495 10.235 99.67 10.745 ;
      RECT 89.11 10.235 89.285 10.745 ;
      RECT 88.12 1.865 88.295 2.375 ;
      RECT 88.12 10.235 88.295 10.745 ;
      RECT 86.33 1.865 86.505 2.375 ;
      RECT 86.33 10.235 86.505 10.745 ;
      RECT 81.57 10.235 81.745 10.745 ;
      RECT 71.185 10.235 71.36 10.745 ;
      RECT 70.195 1.865 70.37 2.375 ;
      RECT 70.195 10.235 70.37 10.745 ;
      RECT 68.405 1.865 68.58 2.375 ;
      RECT 68.405 10.235 68.58 10.745 ;
      RECT 63.645 10.235 63.82 10.745 ;
      RECT 53.26 10.235 53.435 10.745 ;
      RECT 52.27 1.865 52.445 2.375 ;
      RECT 52.27 10.235 52.445 10.745 ;
      RECT 50.48 1.865 50.655 2.375 ;
      RECT 50.48 10.235 50.655 10.745 ;
      RECT 45.72 10.235 45.895 10.745 ;
      RECT 35.335 10.235 35.51 10.745 ;
      RECT 34.345 1.865 34.52 2.375 ;
      RECT 34.345 10.235 34.52 10.745 ;
      RECT 32.555 1.865 32.73 2.375 ;
      RECT 32.555 10.235 32.73 10.745 ;
      RECT 27.795 10.235 27.97 10.745 ;
      RECT 16.765 10.235 16.94 10.745 ;
  END
END sky130_osu_ring_oscillator_mpr2at_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2ca_8_b0r1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ca_8_b0r1 ;
  SIZE 100.725 BY 12.455 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 33.745 0 34.125 5.26 ;
      LAYER met2 ;
        RECT 33.745 4.88 34.125 5.26 ;
      LAYER li1 ;
        RECT 33.845 1.87 34.02 2.38 ;
        RECT 33.845 3.9 34.02 5.16 ;
        RECT 33.845 3.69 34.015 5.16 ;
      LAYER met1 ;
        RECT 33.76 4.925 34.11 5.215 ;
        RECT 33.785 2.18 34.08 2.41 ;
        RECT 33.785 3.66 34.075 3.89 ;
        RECT 33.845 2.18 34.015 3.89 ;
      LAYER via1 ;
        RECT 33.86 4.995 34.01 5.145 ;
      LAYER via2 ;
        RECT 33.835 4.97 34.035 5.17 ;
      LAYER mcon ;
        RECT 33.845 3.69 34.015 3.86 ;
        RECT 33.845 2.21 34.015 2.38 ;
        RECT 33.85 4.985 34.02 5.155 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 50.33 0 50.71 5.26 ;
      LAYER met2 ;
        RECT 50.33 4.88 50.71 5.26 ;
      LAYER li1 ;
        RECT 50.43 1.87 50.605 2.38 ;
        RECT 50.43 3.9 50.605 5.16 ;
        RECT 50.43 3.69 50.6 5.16 ;
      LAYER met1 ;
        RECT 50.345 4.925 50.695 5.215 ;
        RECT 50.37 2.18 50.665 2.41 ;
        RECT 50.37 3.66 50.66 3.89 ;
        RECT 50.43 2.18 50.6 3.89 ;
      LAYER via1 ;
        RECT 50.445 4.995 50.595 5.145 ;
      LAYER via2 ;
        RECT 50.42 4.97 50.62 5.17 ;
      LAYER mcon ;
        RECT 50.43 3.69 50.6 3.86 ;
        RECT 50.43 2.21 50.6 2.38 ;
        RECT 50.435 4.985 50.605 5.155 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 66.915 0 67.295 5.26 ;
      LAYER met2 ;
        RECT 66.915 4.88 67.295 5.26 ;
      LAYER li1 ;
        RECT 67.015 1.87 67.19 2.38 ;
        RECT 67.015 3.9 67.19 5.16 ;
        RECT 67.015 3.69 67.185 5.16 ;
      LAYER met1 ;
        RECT 66.93 4.925 67.28 5.215 ;
        RECT 66.955 2.18 67.25 2.41 ;
        RECT 66.955 3.66 67.245 3.89 ;
        RECT 67.015 2.18 67.185 3.89 ;
      LAYER via1 ;
        RECT 67.03 4.995 67.18 5.145 ;
      LAYER via2 ;
        RECT 67.005 4.97 67.205 5.17 ;
      LAYER mcon ;
        RECT 67.015 3.69 67.185 3.86 ;
        RECT 67.015 2.21 67.185 2.38 ;
        RECT 67.02 4.985 67.19 5.155 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 83.5 0 83.88 5.26 ;
      LAYER met2 ;
        RECT 83.5 4.88 83.88 5.26 ;
      LAYER li1 ;
        RECT 83.6 1.87 83.775 2.38 ;
        RECT 83.6 3.9 83.775 5.16 ;
        RECT 83.6 3.69 83.77 5.16 ;
      LAYER met1 ;
        RECT 83.515 4.925 83.865 5.215 ;
        RECT 83.54 2.18 83.835 2.41 ;
        RECT 83.54 3.66 83.83 3.89 ;
        RECT 83.6 2.18 83.77 3.89 ;
      LAYER via1 ;
        RECT 83.615 4.995 83.765 5.145 ;
      LAYER via2 ;
        RECT 83.59 4.97 83.79 5.17 ;
      LAYER mcon ;
        RECT 83.6 3.69 83.77 3.86 ;
        RECT 83.6 2.21 83.77 2.38 ;
        RECT 83.605 4.985 83.775 5.155 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 100.08 0 100.46 5.26 ;
      LAYER met2 ;
        RECT 100.08 4.88 100.46 5.26 ;
      LAYER li1 ;
        RECT 100.18 1.87 100.355 2.38 ;
        RECT 100.18 3.9 100.355 5.16 ;
        RECT 100.18 3.69 100.35 5.16 ;
      LAYER met1 ;
        RECT 100.095 4.925 100.445 5.215 ;
        RECT 100.12 2.18 100.415 2.41 ;
        RECT 100.12 3.66 100.41 3.89 ;
        RECT 100.18 2.18 100.35 3.89 ;
      LAYER via1 ;
        RECT 100.195 4.995 100.345 5.145 ;
      LAYER via2 ;
        RECT 100.17 4.97 100.37 5.17 ;
      LAYER mcon ;
        RECT 100.18 3.69 100.35 3.86 ;
        RECT 100.18 2.21 100.35 2.38 ;
        RECT 100.185 4.985 100.355 5.155 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 29.62 8.15 29.945 8.475 ;
        RECT 29.615 4.93 29.94 5.255 ;
        RECT 20.775 9.315 29.86 9.485 ;
        RECT 29.685 4.93 29.86 9.485 ;
        RECT 20.72 8.145 21 8.485 ;
        RECT 20.775 8.145 20.945 9.485 ;
      LAYER li1 ;
        RECT 29.69 2.96 29.86 4.23 ;
        RECT 29.69 8.23 29.86 9.5 ;
        RECT 18.465 8.225 18.635 9.495 ;
      LAYER met1 ;
        RECT 29.63 4.06 30.09 4.23 ;
        RECT 29.615 4.93 29.94 5.255 ;
        RECT 29.63 4.03 29.92 4.26 ;
        RECT 29.69 4.03 29.87 5.255 ;
        RECT 29.62 8.23 30.09 8.4 ;
        RECT 29.62 8.15 29.945 8.475 ;
        RECT 20.69 8.175 21.03 8.455 ;
        RECT 18.405 8.23 21.03 8.4 ;
        RECT 18.405 8.225 18.865 8.4 ;
        RECT 18.405 8.195 18.695 8.425 ;
      LAYER via1 ;
        RECT 20.785 8.24 20.935 8.39 ;
        RECT 29.705 5.015 29.855 5.165 ;
        RECT 29.71 8.235 29.86 8.385 ;
      LAYER mcon ;
        RECT 18.465 8.225 18.635 8.395 ;
        RECT 29.69 8.23 29.86 8.4 ;
        RECT 29.69 4.06 29.86 4.23 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 46.205 8.15 46.53 8.475 ;
        RECT 46.2 4.93 46.525 5.255 ;
        RECT 37.36 9.315 46.445 9.485 ;
        RECT 46.27 4.93 46.445 9.485 ;
        RECT 37.305 8.145 37.585 8.485 ;
        RECT 37.36 8.145 37.53 9.485 ;
      LAYER li1 ;
        RECT 46.275 2.96 46.445 4.23 ;
        RECT 46.275 8.23 46.445 9.5 ;
        RECT 35.05 8.225 35.22 9.495 ;
      LAYER met1 ;
        RECT 46.215 4.06 46.675 4.23 ;
        RECT 46.2 4.93 46.525 5.255 ;
        RECT 46.215 4.03 46.505 4.26 ;
        RECT 46.275 4.03 46.455 5.255 ;
        RECT 46.205 8.23 46.675 8.4 ;
        RECT 46.205 8.15 46.53 8.475 ;
        RECT 37.275 8.175 37.615 8.455 ;
        RECT 34.99 8.23 37.615 8.4 ;
        RECT 34.99 8.225 35.45 8.4 ;
        RECT 34.99 8.195 35.28 8.425 ;
      LAYER via1 ;
        RECT 37.37 8.24 37.52 8.39 ;
        RECT 46.29 5.015 46.44 5.165 ;
        RECT 46.295 8.235 46.445 8.385 ;
      LAYER mcon ;
        RECT 35.05 8.225 35.22 8.395 ;
        RECT 46.275 8.23 46.445 8.4 ;
        RECT 46.275 4.06 46.445 4.23 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 62.79 8.15 63.115 8.475 ;
        RECT 62.785 4.93 63.11 5.255 ;
        RECT 53.945 9.315 63.03 9.485 ;
        RECT 62.855 4.93 63.03 9.485 ;
        RECT 53.89 8.145 54.17 8.485 ;
        RECT 53.945 8.145 54.115 9.485 ;
      LAYER li1 ;
        RECT 62.86 2.96 63.03 4.23 ;
        RECT 62.86 8.23 63.03 9.5 ;
        RECT 51.635 8.225 51.805 9.495 ;
      LAYER met1 ;
        RECT 62.8 4.06 63.26 4.23 ;
        RECT 62.785 4.93 63.11 5.255 ;
        RECT 62.8 4.03 63.09 4.26 ;
        RECT 62.86 4.03 63.04 5.255 ;
        RECT 62.79 8.23 63.26 8.4 ;
        RECT 62.79 8.15 63.115 8.475 ;
        RECT 53.86 8.175 54.2 8.455 ;
        RECT 51.575 8.23 54.2 8.4 ;
        RECT 51.575 8.225 52.035 8.4 ;
        RECT 51.575 8.195 51.865 8.425 ;
      LAYER via1 ;
        RECT 53.955 8.24 54.105 8.39 ;
        RECT 62.875 5.015 63.025 5.165 ;
        RECT 62.88 8.235 63.03 8.385 ;
      LAYER mcon ;
        RECT 51.635 8.225 51.805 8.395 ;
        RECT 62.86 8.23 63.03 8.4 ;
        RECT 62.86 4.06 63.03 4.23 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 79.375 8.15 79.7 8.475 ;
        RECT 79.37 4.93 79.695 5.255 ;
        RECT 70.53 9.315 79.615 9.485 ;
        RECT 79.44 4.93 79.615 9.485 ;
        RECT 70.475 8.145 70.755 8.485 ;
        RECT 70.53 8.145 70.7 9.485 ;
      LAYER li1 ;
        RECT 79.445 2.96 79.615 4.23 ;
        RECT 79.445 8.23 79.615 9.5 ;
        RECT 68.22 8.225 68.39 9.495 ;
      LAYER met1 ;
        RECT 79.385 4.06 79.845 4.23 ;
        RECT 79.37 4.93 79.695 5.255 ;
        RECT 79.385 4.03 79.675 4.26 ;
        RECT 79.445 4.03 79.625 5.255 ;
        RECT 79.375 8.23 79.845 8.4 ;
        RECT 79.375 8.15 79.7 8.475 ;
        RECT 70.445 8.175 70.785 8.455 ;
        RECT 68.16 8.23 70.785 8.4 ;
        RECT 68.16 8.225 68.62 8.4 ;
        RECT 68.16 8.195 68.45 8.425 ;
      LAYER via1 ;
        RECT 70.54 8.24 70.69 8.39 ;
        RECT 79.46 5.015 79.61 5.165 ;
        RECT 79.465 8.235 79.615 8.385 ;
      LAYER mcon ;
        RECT 68.22 8.225 68.39 8.395 ;
        RECT 79.445 8.23 79.615 8.4 ;
        RECT 79.445 4.06 79.615 4.23 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 95.955 8.15 96.28 8.475 ;
        RECT 95.95 4.93 96.275 5.255 ;
        RECT 87.11 9.315 96.195 9.485 ;
        RECT 96.02 4.93 96.195 9.485 ;
        RECT 87.055 8.145 87.335 8.485 ;
        RECT 87.11 8.145 87.28 9.485 ;
      LAYER li1 ;
        RECT 96.025 2.96 96.195 4.23 ;
        RECT 96.025 8.23 96.195 9.5 ;
        RECT 84.8 8.225 84.97 9.495 ;
      LAYER met1 ;
        RECT 95.965 4.06 96.425 4.23 ;
        RECT 95.95 4.93 96.275 5.255 ;
        RECT 95.965 4.03 96.255 4.26 ;
        RECT 96.025 4.03 96.205 5.255 ;
        RECT 95.955 8.23 96.425 8.4 ;
        RECT 95.955 8.15 96.28 8.475 ;
        RECT 87.025 8.175 87.365 8.455 ;
        RECT 84.74 8.23 87.365 8.4 ;
        RECT 84.74 8.225 85.2 8.4 ;
        RECT 84.74 8.195 85.03 8.425 ;
      LAYER via1 ;
        RECT 87.12 8.24 87.27 8.39 ;
        RECT 96.04 5.015 96.19 5.165 ;
        RECT 96.045 8.235 96.195 8.385 ;
      LAYER mcon ;
        RECT 84.8 8.225 84.97 8.395 ;
        RECT 96.025 8.23 96.195 8.4 ;
        RECT 96.025 4.06 96.195 4.23 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 15.235 8.225 15.405 9.495 ;
      LAYER met1 ;
        RECT 15.175 8.225 15.635 8.395 ;
        RECT 15.175 8.195 15.47 8.425 ;
      LAYER mcon ;
        RECT 15.235 8.225 15.405 8.395 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 94.785 5.43 100.725 7.03 ;
        RECT 99.75 4.7 99.92 7.76 ;
        RECT 98.76 4.7 98.93 7.76 ;
        RECT 96.015 4.7 96.185 7.76 ;
        RECT 94.655 5.43 100.725 5.965 ;
        RECT 94.325 4.495 94.655 5.805 ;
        RECT 0 5.635 100.725 5.805 ;
        RECT 92.585 5.095 92.845 5.805 ;
        RECT 92.025 5.635 92.395 6.185 ;
        RECT 91.585 4.715 91.915 4.955 ;
        RECT 91.585 4.715 91.775 4.985 ;
        RECT 91.155 4.985 91.765 5.805 ;
        RECT 91.205 4.985 91.475 6.585 ;
        RECT 90.285 5.095 90.505 5.805 ;
        RECT 90.045 5.635 90.325 6.475 ;
        RECT 89.275 4.765 89.605 4.955 ;
        RECT 88.855 5.135 89.475 5.805 ;
        RECT 89.275 4.765 89.475 5.805 ;
        RECT 89.045 5.135 89.375 6.525 ;
        RECT 87.935 5.125 88.195 5.805 ;
        RECT 78.205 5.43 87.96 7.03 ;
        RECT 83.965 5.425 88.195 5.805 ;
        RECT 84.79 5.425 84.96 7.755 ;
        RECT 83.17 4.7 83.34 7.76 ;
        RECT 82.18 4.7 82.35 7.76 ;
        RECT 79.435 4.7 79.605 7.76 ;
        RECT 78.075 5.43 87.96 5.965 ;
        RECT 77.745 4.495 78.075 5.805 ;
        RECT 76.005 5.095 76.265 5.805 ;
        RECT 75.445 5.635 75.815 6.185 ;
        RECT 75.005 4.715 75.335 4.955 ;
        RECT 75.005 4.715 75.195 4.985 ;
        RECT 74.575 4.985 75.185 5.805 ;
        RECT 74.625 4.985 74.895 6.585 ;
        RECT 73.705 5.095 73.925 5.805 ;
        RECT 73.465 5.635 73.745 6.475 ;
        RECT 72.695 4.765 73.025 4.955 ;
        RECT 72.275 5.135 72.895 5.805 ;
        RECT 72.695 4.765 72.895 5.805 ;
        RECT 72.465 5.135 72.795 6.525 ;
        RECT 71.355 5.125 71.615 5.805 ;
        RECT 61.62 5.43 71.375 7.03 ;
        RECT 67.385 5.425 71.615 5.805 ;
        RECT 68.21 5.425 68.38 7.755 ;
        RECT 66.585 4.7 66.755 7.76 ;
        RECT 65.595 4.7 65.765 7.76 ;
        RECT 62.85 4.7 63.02 7.76 ;
        RECT 61.49 5.43 71.375 5.965 ;
        RECT 61.16 4.495 61.49 5.805 ;
        RECT 59.42 5.095 59.68 5.805 ;
        RECT 58.86 5.635 59.23 6.185 ;
        RECT 58.42 4.715 58.75 4.955 ;
        RECT 58.42 4.715 58.61 4.985 ;
        RECT 57.99 4.985 58.6 5.805 ;
        RECT 58.04 4.985 58.31 6.585 ;
        RECT 57.12 5.095 57.34 5.805 ;
        RECT 56.88 5.635 57.16 6.475 ;
        RECT 56.11 4.765 56.44 4.955 ;
        RECT 55.69 5.135 56.31 5.805 ;
        RECT 56.11 4.765 56.31 5.805 ;
        RECT 55.88 5.135 56.21 6.525 ;
        RECT 54.77 5.125 55.03 5.805 ;
        RECT 45.035 5.43 54.79 7.03 ;
        RECT 50.805 5.425 55.03 5.805 ;
        RECT 51.625 5.425 51.795 7.755 ;
        RECT 50 4.7 50.17 7.76 ;
        RECT 49.01 4.7 49.18 7.76 ;
        RECT 46.265 4.7 46.435 7.76 ;
        RECT 44.905 5.43 54.79 5.965 ;
        RECT 44.575 4.495 44.905 5.805 ;
        RECT 42.835 5.095 43.095 5.805 ;
        RECT 42.275 5.635 42.645 6.185 ;
        RECT 41.835 4.715 42.165 4.955 ;
        RECT 41.835 4.715 42.025 4.985 ;
        RECT 41.405 4.985 42.015 5.805 ;
        RECT 41.455 4.985 41.725 6.585 ;
        RECT 40.535 5.095 40.755 5.805 ;
        RECT 40.295 5.635 40.575 6.475 ;
        RECT 39.525 4.765 39.855 4.955 ;
        RECT 39.105 5.135 39.725 5.805 ;
        RECT 39.525 4.765 39.725 5.805 ;
        RECT 39.295 5.135 39.625 6.525 ;
        RECT 38.185 5.125 38.445 5.805 ;
        RECT 28.45 5.43 38.205 7.03 ;
        RECT 34.225 5.425 38.445 5.805 ;
        RECT 35.04 5.425 35.21 7.755 ;
        RECT 33.415 4.7 33.585 7.76 ;
        RECT 32.425 4.7 32.595 7.76 ;
        RECT 29.68 4.7 29.85 7.76 ;
        RECT 28.32 5.43 38.205 5.965 ;
        RECT 27.99 4.495 28.32 5.805 ;
        RECT 26.25 5.095 26.51 5.805 ;
        RECT 25.69 5.635 26.06 6.185 ;
        RECT 25.25 4.715 25.58 4.955 ;
        RECT 25.25 4.715 25.44 4.985 ;
        RECT 24.82 4.985 25.43 5.805 ;
        RECT 24.87 4.985 25.14 6.585 ;
        RECT 23.95 5.095 24.17 5.805 ;
        RECT 23.71 5.635 23.99 6.475 ;
        RECT 22.94 4.765 23.27 4.955 ;
        RECT 22.52 5.135 23.14 5.805 ;
        RECT 22.94 4.765 23.14 5.805 ;
        RECT 22.71 5.135 23.04 6.525 ;
        RECT 21.6 5.125 21.86 5.805 ;
        RECT 0 5.425 21.62 7.025 ;
        RECT 18.455 5.425 18.625 7.755 ;
        RECT 17.04 10.035 17.215 10.585 ;
        RECT 17.04 7.295 17.215 8.435 ;
        RECT 17.04 5.425 17.21 10.585 ;
        RECT 15.225 5.425 15.395 7.755 ;
      LAYER met1 ;
        RECT 94.785 5.43 100.725 7.03 ;
        RECT 0 5.485 100.725 5.965 ;
        RECT 94.655 5.43 100.725 5.965 ;
        RECT 78.205 5.43 87.96 7.03 ;
        RECT 83.965 5.425 87.955 7.03 ;
        RECT 78.075 5.43 87.96 5.965 ;
        RECT 61.62 5.43 71.375 7.03 ;
        RECT 67.385 5.425 71.375 7.03 ;
        RECT 61.49 5.43 71.375 5.965 ;
        RECT 45.035 5.43 54.79 7.03 ;
        RECT 50.805 5.425 54.79 7.03 ;
        RECT 44.905 5.43 54.79 5.965 ;
        RECT 28.45 5.43 38.205 7.03 ;
        RECT 34.225 5.425 38.205 7.03 ;
        RECT 28.32 5.43 38.205 5.965 ;
        RECT 0 5.425 21.62 7.025 ;
        RECT 16.98 8.935 17.27 9.165 ;
        RECT 16.81 8.965 17.27 9.135 ;
      LAYER mcon ;
        RECT 17.04 8.965 17.21 9.135 ;
        RECT 17.345 6.825 17.515 6.995 ;
        RECT 20.575 6.825 20.745 6.995 ;
        RECT 21.66 5.635 21.83 5.805 ;
        RECT 22.12 5.635 22.29 5.805 ;
        RECT 22.58 5.635 22.75 5.805 ;
        RECT 23.04 5.635 23.21 5.805 ;
        RECT 23.5 5.635 23.67 5.805 ;
        RECT 23.96 5.635 24.13 5.805 ;
        RECT 24.42 5.635 24.59 5.805 ;
        RECT 24.88 5.635 25.05 5.805 ;
        RECT 25.34 5.635 25.51 5.805 ;
        RECT 25.8 5.635 25.97 5.805 ;
        RECT 26.26 5.635 26.43 5.805 ;
        RECT 26.72 5.635 26.89 5.805 ;
        RECT 27.18 5.635 27.35 5.805 ;
        RECT 27.64 5.635 27.81 5.805 ;
        RECT 28.1 5.635 28.27 5.805 ;
        RECT 31.8 6.83 31.97 7 ;
        RECT 31.8 5.46 31.97 5.63 ;
        RECT 32.505 6.83 32.675 7 ;
        RECT 32.505 5.46 32.675 5.63 ;
        RECT 33.495 6.83 33.665 7 ;
        RECT 33.495 5.46 33.665 5.63 ;
        RECT 37.16 6.825 37.33 6.995 ;
        RECT 38.245 5.635 38.415 5.805 ;
        RECT 38.705 5.635 38.875 5.805 ;
        RECT 39.165 5.635 39.335 5.805 ;
        RECT 39.625 5.635 39.795 5.805 ;
        RECT 40.085 5.635 40.255 5.805 ;
        RECT 40.545 5.635 40.715 5.805 ;
        RECT 41.005 5.635 41.175 5.805 ;
        RECT 41.465 5.635 41.635 5.805 ;
        RECT 41.925 5.635 42.095 5.805 ;
        RECT 42.385 5.635 42.555 5.805 ;
        RECT 42.845 5.635 43.015 5.805 ;
        RECT 43.305 5.635 43.475 5.805 ;
        RECT 43.765 5.635 43.935 5.805 ;
        RECT 44.225 5.635 44.395 5.805 ;
        RECT 44.685 5.635 44.855 5.805 ;
        RECT 48.385 6.83 48.555 7 ;
        RECT 48.385 5.46 48.555 5.63 ;
        RECT 49.09 6.83 49.26 7 ;
        RECT 49.09 5.46 49.26 5.63 ;
        RECT 50.08 6.83 50.25 7 ;
        RECT 50.08 5.46 50.25 5.63 ;
        RECT 53.745 6.825 53.915 6.995 ;
        RECT 54.83 5.635 55 5.805 ;
        RECT 55.29 5.635 55.46 5.805 ;
        RECT 55.75 5.635 55.92 5.805 ;
        RECT 56.21 5.635 56.38 5.805 ;
        RECT 56.67 5.635 56.84 5.805 ;
        RECT 57.13 5.635 57.3 5.805 ;
        RECT 57.59 5.635 57.76 5.805 ;
        RECT 58.05 5.635 58.22 5.805 ;
        RECT 58.51 5.635 58.68 5.805 ;
        RECT 58.97 5.635 59.14 5.805 ;
        RECT 59.43 5.635 59.6 5.805 ;
        RECT 59.89 5.635 60.06 5.805 ;
        RECT 60.35 5.635 60.52 5.805 ;
        RECT 60.81 5.635 60.98 5.805 ;
        RECT 61.27 5.635 61.44 5.805 ;
        RECT 64.97 6.83 65.14 7 ;
        RECT 64.97 5.46 65.14 5.63 ;
        RECT 65.675 6.83 65.845 7 ;
        RECT 65.675 5.46 65.845 5.63 ;
        RECT 66.665 6.83 66.835 7 ;
        RECT 66.665 5.46 66.835 5.63 ;
        RECT 70.33 6.825 70.5 6.995 ;
        RECT 71.415 5.635 71.585 5.805 ;
        RECT 71.875 5.635 72.045 5.805 ;
        RECT 72.335 5.635 72.505 5.805 ;
        RECT 72.795 5.635 72.965 5.805 ;
        RECT 73.255 5.635 73.425 5.805 ;
        RECT 73.715 5.635 73.885 5.805 ;
        RECT 74.175 5.635 74.345 5.805 ;
        RECT 74.635 5.635 74.805 5.805 ;
        RECT 75.095 5.635 75.265 5.805 ;
        RECT 75.555 5.635 75.725 5.805 ;
        RECT 76.015 5.635 76.185 5.805 ;
        RECT 76.475 5.635 76.645 5.805 ;
        RECT 76.935 5.635 77.105 5.805 ;
        RECT 77.395 5.635 77.565 5.805 ;
        RECT 77.855 5.635 78.025 5.805 ;
        RECT 81.555 6.83 81.725 7 ;
        RECT 81.555 5.46 81.725 5.63 ;
        RECT 82.26 6.83 82.43 7 ;
        RECT 82.26 5.46 82.43 5.63 ;
        RECT 83.25 6.83 83.42 7 ;
        RECT 83.25 5.46 83.42 5.63 ;
        RECT 86.91 6.825 87.08 6.995 ;
        RECT 87.995 5.635 88.165 5.805 ;
        RECT 88.455 5.635 88.625 5.805 ;
        RECT 88.915 5.635 89.085 5.805 ;
        RECT 89.375 5.635 89.545 5.805 ;
        RECT 89.835 5.635 90.005 5.805 ;
        RECT 90.295 5.635 90.465 5.805 ;
        RECT 90.755 5.635 90.925 5.805 ;
        RECT 91.215 5.635 91.385 5.805 ;
        RECT 91.675 5.635 91.845 5.805 ;
        RECT 92.135 5.635 92.305 5.805 ;
        RECT 92.595 5.635 92.765 5.805 ;
        RECT 93.055 5.635 93.225 5.805 ;
        RECT 93.515 5.635 93.685 5.805 ;
        RECT 93.975 5.635 94.145 5.805 ;
        RECT 94.435 5.635 94.605 5.805 ;
        RECT 98.135 6.83 98.305 7 ;
        RECT 98.135 5.46 98.305 5.63 ;
        RECT 98.84 6.83 99.01 7 ;
        RECT 98.84 5.46 99.01 5.63 ;
        RECT 99.83 6.83 100 7 ;
        RECT 99.83 5.46 100 5.63 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 90.225 7.725 90.56 8.1 ;
        RECT 90.195 7.785 90.535 8.195 ;
        RECT 90.22 7.76 90.56 8.1 ;
        RECT 89.755 7.785 90.56 8.085 ;
        RECT 73.645 7.725 73.98 8.1 ;
        RECT 73.615 7.785 73.955 8.195 ;
        RECT 73.64 7.76 73.98 8.1 ;
        RECT 73.175 7.785 73.98 8.085 ;
        RECT 57.06 7.725 57.395 8.1 ;
        RECT 57.03 7.785 57.37 8.195 ;
        RECT 57.055 7.76 57.395 8.1 ;
        RECT 56.59 7.785 57.395 8.085 ;
        RECT 40.475 7.725 40.81 8.1 ;
        RECT 40.445 7.785 40.785 8.195 ;
        RECT 40.47 7.76 40.81 8.1 ;
        RECT 40.005 7.785 40.81 8.085 ;
        RECT 23.89 7.725 24.225 8.1 ;
        RECT 23.86 7.785 24.2 8.195 ;
        RECT 23.885 7.76 24.225 8.1 ;
        RECT 23.42 7.785 24.225 8.085 ;
      LAYER met2 ;
        RECT 90.255 7.72 90.535 8.095 ;
        RECT 73.675 7.72 73.955 8.095 ;
        RECT 57.09 7.72 57.37 8.095 ;
        RECT 40.505 7.72 40.785 8.095 ;
        RECT 23.92 7.72 24.2 8.095 ;
      LAYER li1 ;
        RECT 0 0 100.725 1.6 ;
        RECT 99.75 0 99.92 2.23 ;
        RECT 98.76 0 98.93 2.23 ;
        RECT 96.015 0 96.185 2.23 ;
        RECT 87.6 0 94.945 3.095 ;
        RECT 94.385 0 94.655 3.895 ;
        RECT 93.475 0 93.715 3.895 ;
        RECT 92.605 0 92.855 3.625 ;
        RECT 90.225 0 90.555 3.545 ;
        RECT 87.935 0 88.195 3.905 ;
        RECT 83.17 0 83.34 2.23 ;
        RECT 82.18 0 82.35 2.23 ;
        RECT 79.435 0 79.605 2.23 ;
        RECT 71.02 0 78.365 3.095 ;
        RECT 77.805 0 78.075 3.895 ;
        RECT 76.895 0 77.135 3.895 ;
        RECT 76.025 0 76.275 3.625 ;
        RECT 73.645 0 73.975 3.545 ;
        RECT 71.355 0 71.615 3.905 ;
        RECT 66.585 0 66.755 2.23 ;
        RECT 65.595 0 65.765 2.23 ;
        RECT 62.85 0 63.02 2.23 ;
        RECT 54.435 0 61.78 3.095 ;
        RECT 61.22 0 61.49 3.895 ;
        RECT 60.31 0 60.55 3.895 ;
        RECT 59.44 0 59.69 3.625 ;
        RECT 57.06 0 57.39 3.545 ;
        RECT 54.77 0 55.03 3.905 ;
        RECT 50 0 50.17 2.23 ;
        RECT 49.01 0 49.18 2.23 ;
        RECT 46.265 0 46.435 2.23 ;
        RECT 37.85 0 45.195 3.095 ;
        RECT 44.635 0 44.905 3.895 ;
        RECT 43.725 0 43.965 3.895 ;
        RECT 42.855 0 43.105 3.625 ;
        RECT 40.475 0 40.805 3.545 ;
        RECT 38.185 0 38.445 3.905 ;
        RECT 33.415 0 33.585 2.23 ;
        RECT 32.425 0 32.595 2.23 ;
        RECT 29.68 0 29.85 2.23 ;
        RECT 21.265 0 28.61 3.095 ;
        RECT 28.05 0 28.32 3.895 ;
        RECT 27.14 0 27.38 3.895 ;
        RECT 26.27 0 26.52 3.625 ;
        RECT 23.89 0 24.22 3.545 ;
        RECT 21.6 0 21.86 3.905 ;
        RECT 0.055 10.855 100.725 12.455 ;
        RECT 99.75 10.23 99.92 12.455 ;
        RECT 98.76 10.23 98.93 12.455 ;
        RECT 96.015 10.23 96.185 12.455 ;
        RECT 87.85 9.465 94.77 12.455 ;
        RECT 87.855 8.355 94.77 12.455 ;
        RECT 93.285 7.845 93.735 12.455 ;
        RECT 91.195 7.955 91.525 12.455 ;
        RECT 89.125 7.895 89.375 12.455 ;
        RECT 84.79 10.225 84.96 12.455 ;
        RECT 83.17 10.23 83.34 12.455 ;
        RECT 82.18 10.23 82.35 12.455 ;
        RECT 79.435 10.23 79.605 12.455 ;
        RECT 71.27 9.465 78.19 12.455 ;
        RECT 71.275 8.355 78.19 12.455 ;
        RECT 76.705 7.845 77.155 12.455 ;
        RECT 74.615 7.955 74.945 12.455 ;
        RECT 72.545 7.895 72.795 12.455 ;
        RECT 68.21 10.225 68.38 12.455 ;
        RECT 66.585 10.23 66.755 12.455 ;
        RECT 65.595 10.23 65.765 12.455 ;
        RECT 62.85 10.23 63.02 12.455 ;
        RECT 54.685 9.465 61.605 12.455 ;
        RECT 54.69 8.355 61.605 12.455 ;
        RECT 60.12 7.845 60.57 12.455 ;
        RECT 58.03 7.955 58.36 12.455 ;
        RECT 55.96 7.895 56.21 12.455 ;
        RECT 51.625 10.225 51.795 12.455 ;
        RECT 50 10.23 50.17 12.455 ;
        RECT 49.01 10.23 49.18 12.455 ;
        RECT 46.265 10.23 46.435 12.455 ;
        RECT 38.1 9.465 45.02 12.455 ;
        RECT 38.105 8.355 45.02 12.455 ;
        RECT 43.535 7.845 43.985 12.455 ;
        RECT 41.445 7.955 41.775 12.455 ;
        RECT 39.375 7.895 39.625 12.455 ;
        RECT 35.04 10.225 35.21 12.455 ;
        RECT 33.415 10.23 33.585 12.455 ;
        RECT 32.425 10.23 32.595 12.455 ;
        RECT 29.68 10.23 29.85 12.455 ;
        RECT 21.515 9.465 28.435 12.455 ;
        RECT 21.52 8.355 28.435 12.455 ;
        RECT 26.95 7.845 27.4 12.455 ;
        RECT 24.86 7.955 25.19 12.455 ;
        RECT 22.79 7.895 23.04 12.455 ;
        RECT 18.455 10.225 18.625 12.455 ;
        RECT 15.225 10.225 15.395 12.455 ;
        RECT 91.495 7.115 91.825 7.445 ;
        RECT 89.275 7.115 89.615 7.365 ;
        RECT 85.805 8.355 85.975 10.305 ;
        RECT 85.745 10.135 85.915 10.585 ;
        RECT 85.745 7.295 85.915 8.525 ;
        RECT 74.915 7.115 75.245 7.445 ;
        RECT 72.695 7.115 73.035 7.365 ;
        RECT 69.225 8.355 69.395 10.305 ;
        RECT 69.165 10.135 69.335 10.585 ;
        RECT 69.165 7.295 69.335 8.525 ;
        RECT 58.33 7.115 58.66 7.445 ;
        RECT 56.11 7.115 56.45 7.365 ;
        RECT 52.64 8.355 52.81 10.305 ;
        RECT 52.58 10.135 52.75 10.585 ;
        RECT 52.58 7.295 52.75 8.525 ;
        RECT 41.745 7.115 42.075 7.445 ;
        RECT 39.525 7.115 39.865 7.365 ;
        RECT 36.055 8.355 36.225 10.305 ;
        RECT 35.995 10.135 36.165 10.585 ;
        RECT 35.995 7.295 36.165 8.525 ;
        RECT 25.16 7.115 25.49 7.445 ;
        RECT 22.94 7.115 23.28 7.365 ;
        RECT 19.47 8.355 19.64 10.305 ;
        RECT 19.41 10.135 19.58 10.585 ;
        RECT 19.41 7.295 19.58 8.525 ;
      LAYER met1 ;
        RECT 0 0 100.725 1.6 ;
        RECT 87.6 0 94.945 3.125 ;
        RECT 71.02 0 78.365 3.125 ;
        RECT 54.435 0 61.78 3.125 ;
        RECT 37.85 0 45.195 3.125 ;
        RECT 21.265 0 28.61 3.125 ;
        RECT 0.055 10.855 100.725 12.455 ;
        RECT 87.85 9.465 94.77 12.455 ;
        RECT 87.855 8.325 94.77 12.455 ;
        RECT 91.445 7.135 91.735 7.365 ;
        RECT 89.315 7.805 91.665 7.945 ;
        RECT 91.525 7.135 91.665 7.945 ;
        RECT 90.245 7.805 90.675 8.045 ;
        RECT 90.255 7.78 90.535 8.045 ;
        RECT 90.275 7.75 90.535 8.045 ;
        RECT 89.235 7.135 89.525 7.365 ;
        RECT 89.315 7.135 89.455 12.455 ;
        RECT 85.745 8.565 86.035 8.795 ;
        RECT 85.58 8.595 85.75 12.455 ;
        RECT 85.57 8.595 86.035 8.765 ;
        RECT 71.27 9.465 78.19 12.455 ;
        RECT 71.275 8.325 78.19 12.455 ;
        RECT 74.865 7.135 75.155 7.365 ;
        RECT 72.735 7.805 75.085 7.945 ;
        RECT 74.945 7.135 75.085 7.945 ;
        RECT 73.665 7.805 74.095 8.045 ;
        RECT 73.675 7.78 73.955 8.045 ;
        RECT 73.695 7.75 73.955 8.045 ;
        RECT 72.655 7.135 72.945 7.365 ;
        RECT 72.735 7.135 72.875 12.455 ;
        RECT 69.165 8.565 69.455 8.795 ;
        RECT 69 8.595 69.17 12.455 ;
        RECT 68.99 8.595 69.455 8.765 ;
        RECT 54.685 9.465 61.605 12.455 ;
        RECT 54.69 8.325 61.605 12.455 ;
        RECT 58.28 7.135 58.57 7.365 ;
        RECT 56.15 7.805 58.5 7.945 ;
        RECT 58.36 7.135 58.5 7.945 ;
        RECT 57.08 7.805 57.51 8.045 ;
        RECT 57.09 7.78 57.37 8.045 ;
        RECT 57.11 7.75 57.37 8.045 ;
        RECT 56.07 7.135 56.36 7.365 ;
        RECT 56.15 7.135 56.29 12.455 ;
        RECT 52.58 8.565 52.87 8.795 ;
        RECT 52.415 8.595 52.585 12.455 ;
        RECT 52.405 8.595 52.87 8.765 ;
        RECT 38.1 9.465 45.02 12.455 ;
        RECT 38.105 8.325 45.02 12.455 ;
        RECT 41.695 7.135 41.985 7.365 ;
        RECT 39.565 7.805 41.915 7.945 ;
        RECT 41.775 7.135 41.915 7.945 ;
        RECT 40.495 7.805 40.925 8.045 ;
        RECT 40.505 7.78 40.785 8.045 ;
        RECT 40.525 7.75 40.785 8.045 ;
        RECT 39.485 7.135 39.775 7.365 ;
        RECT 39.565 7.135 39.705 12.455 ;
        RECT 35.995 8.565 36.285 8.795 ;
        RECT 35.83 8.595 36 12.455 ;
        RECT 35.82 8.595 36.285 8.765 ;
        RECT 21.515 9.465 28.435 12.455 ;
        RECT 21.52 8.325 28.435 12.455 ;
        RECT 25.11 7.135 25.4 7.365 ;
        RECT 22.98 7.805 25.33 7.945 ;
        RECT 25.19 7.135 25.33 7.945 ;
        RECT 23.91 7.805 24.34 8.045 ;
        RECT 23.92 7.78 24.2 8.045 ;
        RECT 23.94 7.75 24.2 8.045 ;
        RECT 22.9 7.135 23.19 7.365 ;
        RECT 22.98 7.135 23.12 12.455 ;
        RECT 19.41 8.565 19.7 8.795 ;
        RECT 19.245 8.595 19.415 12.455 ;
        RECT 19.235 8.595 19.7 8.765 ;
      LAYER via1 ;
        RECT 23.995 7.835 24.145 7.985 ;
        RECT 40.58 7.835 40.73 7.985 ;
        RECT 57.165 7.835 57.315 7.985 ;
        RECT 73.75 7.835 73.9 7.985 ;
        RECT 90.33 7.835 90.48 7.985 ;
      LAYER via2 ;
        RECT 23.96 7.81 24.16 8.01 ;
        RECT 40.545 7.81 40.745 8.01 ;
        RECT 57.13 7.81 57.33 8.01 ;
        RECT 73.715 7.81 73.915 8.01 ;
        RECT 90.295 7.81 90.495 8.01 ;
      LAYER mcon ;
        RECT 15.305 10.885 15.475 11.055 ;
        RECT 15.985 10.885 16.155 11.055 ;
        RECT 16.665 10.885 16.835 11.055 ;
        RECT 17.345 10.885 17.515 11.055 ;
        RECT 18.535 10.885 18.705 11.055 ;
        RECT 19.215 10.885 19.385 11.055 ;
        RECT 19.47 8.595 19.64 8.765 ;
        RECT 19.895 10.885 20.065 11.055 ;
        RECT 20.575 10.885 20.745 11.055 ;
        RECT 21.66 8.355 21.83 8.525 ;
        RECT 21.66 2.925 21.83 3.095 ;
        RECT 22.12 8.355 22.29 8.525 ;
        RECT 22.12 2.925 22.29 3.095 ;
        RECT 22.58 8.355 22.75 8.525 ;
        RECT 22.58 2.925 22.75 3.095 ;
        RECT 22.96 7.165 23.13 7.335 ;
        RECT 23.04 8.355 23.21 8.525 ;
        RECT 23.04 2.925 23.21 3.095 ;
        RECT 23.5 8.355 23.67 8.525 ;
        RECT 23.5 2.925 23.67 3.095 ;
        RECT 23.96 8.355 24.13 8.525 ;
        RECT 23.96 2.925 24.13 3.095 ;
        RECT 24.42 8.355 24.59 8.525 ;
        RECT 24.42 2.925 24.59 3.095 ;
        RECT 24.88 8.355 25.05 8.525 ;
        RECT 24.88 2.925 25.05 3.095 ;
        RECT 25.17 7.165 25.34 7.335 ;
        RECT 25.34 8.355 25.51 8.525 ;
        RECT 25.34 2.925 25.51 3.095 ;
        RECT 25.8 8.355 25.97 8.525 ;
        RECT 25.8 2.925 25.97 3.095 ;
        RECT 26.26 8.355 26.43 8.525 ;
        RECT 26.26 2.925 26.43 3.095 ;
        RECT 26.72 8.355 26.89 8.525 ;
        RECT 26.72 2.925 26.89 3.095 ;
        RECT 27.18 8.355 27.35 8.525 ;
        RECT 27.18 2.925 27.35 3.095 ;
        RECT 27.64 8.355 27.81 8.525 ;
        RECT 27.64 2.925 27.81 3.095 ;
        RECT 28.1 8.355 28.27 8.525 ;
        RECT 28.1 2.925 28.27 3.095 ;
        RECT 29.76 10.89 29.93 11.06 ;
        RECT 29.76 1.4 29.93 1.57 ;
        RECT 30.44 10.89 30.61 11.06 ;
        RECT 30.44 1.4 30.61 1.57 ;
        RECT 31.12 10.89 31.29 11.06 ;
        RECT 31.12 1.4 31.29 1.57 ;
        RECT 31.8 10.89 31.97 11.06 ;
        RECT 31.8 1.4 31.97 1.57 ;
        RECT 32.505 10.89 32.675 11.06 ;
        RECT 32.505 1.4 32.675 1.57 ;
        RECT 33.495 10.89 33.665 11.06 ;
        RECT 33.495 1.4 33.665 1.57 ;
        RECT 35.12 10.885 35.29 11.055 ;
        RECT 35.8 10.885 35.97 11.055 ;
        RECT 36.055 8.595 36.225 8.765 ;
        RECT 36.48 10.885 36.65 11.055 ;
        RECT 37.16 10.885 37.33 11.055 ;
        RECT 38.245 8.355 38.415 8.525 ;
        RECT 38.245 2.925 38.415 3.095 ;
        RECT 38.705 8.355 38.875 8.525 ;
        RECT 38.705 2.925 38.875 3.095 ;
        RECT 39.165 8.355 39.335 8.525 ;
        RECT 39.165 2.925 39.335 3.095 ;
        RECT 39.545 7.165 39.715 7.335 ;
        RECT 39.625 8.355 39.795 8.525 ;
        RECT 39.625 2.925 39.795 3.095 ;
        RECT 40.085 8.355 40.255 8.525 ;
        RECT 40.085 2.925 40.255 3.095 ;
        RECT 40.545 8.355 40.715 8.525 ;
        RECT 40.545 2.925 40.715 3.095 ;
        RECT 41.005 8.355 41.175 8.525 ;
        RECT 41.005 2.925 41.175 3.095 ;
        RECT 41.465 8.355 41.635 8.525 ;
        RECT 41.465 2.925 41.635 3.095 ;
        RECT 41.755 7.165 41.925 7.335 ;
        RECT 41.925 8.355 42.095 8.525 ;
        RECT 41.925 2.925 42.095 3.095 ;
        RECT 42.385 8.355 42.555 8.525 ;
        RECT 42.385 2.925 42.555 3.095 ;
        RECT 42.845 8.355 43.015 8.525 ;
        RECT 42.845 2.925 43.015 3.095 ;
        RECT 43.305 8.355 43.475 8.525 ;
        RECT 43.305 2.925 43.475 3.095 ;
        RECT 43.765 8.355 43.935 8.525 ;
        RECT 43.765 2.925 43.935 3.095 ;
        RECT 44.225 8.355 44.395 8.525 ;
        RECT 44.225 2.925 44.395 3.095 ;
        RECT 44.685 8.355 44.855 8.525 ;
        RECT 44.685 2.925 44.855 3.095 ;
        RECT 46.345 10.89 46.515 11.06 ;
        RECT 46.345 1.4 46.515 1.57 ;
        RECT 47.025 10.89 47.195 11.06 ;
        RECT 47.025 1.4 47.195 1.57 ;
        RECT 47.705 10.89 47.875 11.06 ;
        RECT 47.705 1.4 47.875 1.57 ;
        RECT 48.385 10.89 48.555 11.06 ;
        RECT 48.385 1.4 48.555 1.57 ;
        RECT 49.09 10.89 49.26 11.06 ;
        RECT 49.09 1.4 49.26 1.57 ;
        RECT 50.08 10.89 50.25 11.06 ;
        RECT 50.08 1.4 50.25 1.57 ;
        RECT 51.705 10.885 51.875 11.055 ;
        RECT 52.385 10.885 52.555 11.055 ;
        RECT 52.64 8.595 52.81 8.765 ;
        RECT 53.065 10.885 53.235 11.055 ;
        RECT 53.745 10.885 53.915 11.055 ;
        RECT 54.83 8.355 55 8.525 ;
        RECT 54.83 2.925 55 3.095 ;
        RECT 55.29 8.355 55.46 8.525 ;
        RECT 55.29 2.925 55.46 3.095 ;
        RECT 55.75 8.355 55.92 8.525 ;
        RECT 55.75 2.925 55.92 3.095 ;
        RECT 56.13 7.165 56.3 7.335 ;
        RECT 56.21 8.355 56.38 8.525 ;
        RECT 56.21 2.925 56.38 3.095 ;
        RECT 56.67 8.355 56.84 8.525 ;
        RECT 56.67 2.925 56.84 3.095 ;
        RECT 57.13 8.355 57.3 8.525 ;
        RECT 57.13 2.925 57.3 3.095 ;
        RECT 57.59 8.355 57.76 8.525 ;
        RECT 57.59 2.925 57.76 3.095 ;
        RECT 58.05 8.355 58.22 8.525 ;
        RECT 58.05 2.925 58.22 3.095 ;
        RECT 58.34 7.165 58.51 7.335 ;
        RECT 58.51 8.355 58.68 8.525 ;
        RECT 58.51 2.925 58.68 3.095 ;
        RECT 58.97 8.355 59.14 8.525 ;
        RECT 58.97 2.925 59.14 3.095 ;
        RECT 59.43 8.355 59.6 8.525 ;
        RECT 59.43 2.925 59.6 3.095 ;
        RECT 59.89 8.355 60.06 8.525 ;
        RECT 59.89 2.925 60.06 3.095 ;
        RECT 60.35 8.355 60.52 8.525 ;
        RECT 60.35 2.925 60.52 3.095 ;
        RECT 60.81 8.355 60.98 8.525 ;
        RECT 60.81 2.925 60.98 3.095 ;
        RECT 61.27 8.355 61.44 8.525 ;
        RECT 61.27 2.925 61.44 3.095 ;
        RECT 62.93 10.89 63.1 11.06 ;
        RECT 62.93 1.4 63.1 1.57 ;
        RECT 63.61 10.89 63.78 11.06 ;
        RECT 63.61 1.4 63.78 1.57 ;
        RECT 64.29 10.89 64.46 11.06 ;
        RECT 64.29 1.4 64.46 1.57 ;
        RECT 64.97 10.89 65.14 11.06 ;
        RECT 64.97 1.4 65.14 1.57 ;
        RECT 65.675 10.89 65.845 11.06 ;
        RECT 65.675 1.4 65.845 1.57 ;
        RECT 66.665 10.89 66.835 11.06 ;
        RECT 66.665 1.4 66.835 1.57 ;
        RECT 68.29 10.885 68.46 11.055 ;
        RECT 68.97 10.885 69.14 11.055 ;
        RECT 69.225 8.595 69.395 8.765 ;
        RECT 69.65 10.885 69.82 11.055 ;
        RECT 70.33 10.885 70.5 11.055 ;
        RECT 71.415 8.355 71.585 8.525 ;
        RECT 71.415 2.925 71.585 3.095 ;
        RECT 71.875 8.355 72.045 8.525 ;
        RECT 71.875 2.925 72.045 3.095 ;
        RECT 72.335 8.355 72.505 8.525 ;
        RECT 72.335 2.925 72.505 3.095 ;
        RECT 72.715 7.165 72.885 7.335 ;
        RECT 72.795 8.355 72.965 8.525 ;
        RECT 72.795 2.925 72.965 3.095 ;
        RECT 73.255 8.355 73.425 8.525 ;
        RECT 73.255 2.925 73.425 3.095 ;
        RECT 73.715 8.355 73.885 8.525 ;
        RECT 73.715 2.925 73.885 3.095 ;
        RECT 74.175 8.355 74.345 8.525 ;
        RECT 74.175 2.925 74.345 3.095 ;
        RECT 74.635 8.355 74.805 8.525 ;
        RECT 74.635 2.925 74.805 3.095 ;
        RECT 74.925 7.165 75.095 7.335 ;
        RECT 75.095 8.355 75.265 8.525 ;
        RECT 75.095 2.925 75.265 3.095 ;
        RECT 75.555 8.355 75.725 8.525 ;
        RECT 75.555 2.925 75.725 3.095 ;
        RECT 76.015 8.355 76.185 8.525 ;
        RECT 76.015 2.925 76.185 3.095 ;
        RECT 76.475 8.355 76.645 8.525 ;
        RECT 76.475 2.925 76.645 3.095 ;
        RECT 76.935 8.355 77.105 8.525 ;
        RECT 76.935 2.925 77.105 3.095 ;
        RECT 77.395 8.355 77.565 8.525 ;
        RECT 77.395 2.925 77.565 3.095 ;
        RECT 77.855 8.355 78.025 8.525 ;
        RECT 77.855 2.925 78.025 3.095 ;
        RECT 79.515 10.89 79.685 11.06 ;
        RECT 79.515 1.4 79.685 1.57 ;
        RECT 80.195 10.89 80.365 11.06 ;
        RECT 80.195 1.4 80.365 1.57 ;
        RECT 80.875 10.89 81.045 11.06 ;
        RECT 80.875 1.4 81.045 1.57 ;
        RECT 81.555 10.89 81.725 11.06 ;
        RECT 81.555 1.4 81.725 1.57 ;
        RECT 82.26 10.89 82.43 11.06 ;
        RECT 82.26 1.4 82.43 1.57 ;
        RECT 83.25 10.89 83.42 11.06 ;
        RECT 83.25 1.4 83.42 1.57 ;
        RECT 84.87 10.885 85.04 11.055 ;
        RECT 85.55 10.885 85.72 11.055 ;
        RECT 85.805 8.595 85.975 8.765 ;
        RECT 86.23 10.885 86.4 11.055 ;
        RECT 86.91 10.885 87.08 11.055 ;
        RECT 87.995 8.355 88.165 8.525 ;
        RECT 87.995 2.925 88.165 3.095 ;
        RECT 88.455 8.355 88.625 8.525 ;
        RECT 88.455 2.925 88.625 3.095 ;
        RECT 88.915 8.355 89.085 8.525 ;
        RECT 88.915 2.925 89.085 3.095 ;
        RECT 89.295 7.165 89.465 7.335 ;
        RECT 89.375 8.355 89.545 8.525 ;
        RECT 89.375 2.925 89.545 3.095 ;
        RECT 89.835 8.355 90.005 8.525 ;
        RECT 89.835 2.925 90.005 3.095 ;
        RECT 90.295 8.355 90.465 8.525 ;
        RECT 90.295 2.925 90.465 3.095 ;
        RECT 90.755 8.355 90.925 8.525 ;
        RECT 90.755 2.925 90.925 3.095 ;
        RECT 91.215 8.355 91.385 8.525 ;
        RECT 91.215 2.925 91.385 3.095 ;
        RECT 91.505 7.165 91.675 7.335 ;
        RECT 91.675 8.355 91.845 8.525 ;
        RECT 91.675 2.925 91.845 3.095 ;
        RECT 92.135 8.355 92.305 8.525 ;
        RECT 92.135 2.925 92.305 3.095 ;
        RECT 92.595 8.355 92.765 8.525 ;
        RECT 92.595 2.925 92.765 3.095 ;
        RECT 93.055 8.355 93.225 8.525 ;
        RECT 93.055 2.925 93.225 3.095 ;
        RECT 93.515 8.355 93.685 8.525 ;
        RECT 93.515 2.925 93.685 3.095 ;
        RECT 93.975 8.355 94.145 8.525 ;
        RECT 93.975 2.925 94.145 3.095 ;
        RECT 94.435 8.355 94.605 8.525 ;
        RECT 94.435 2.925 94.605 3.095 ;
        RECT 96.095 10.89 96.265 11.06 ;
        RECT 96.095 1.4 96.265 1.57 ;
        RECT 96.775 10.89 96.945 11.06 ;
        RECT 96.775 1.4 96.945 1.57 ;
        RECT 97.455 10.89 97.625 11.06 ;
        RECT 97.455 1.4 97.625 1.57 ;
        RECT 98.135 10.89 98.305 11.06 ;
        RECT 98.135 1.4 98.305 1.57 ;
        RECT 98.84 10.89 99.01 11.06 ;
        RECT 98.84 1.4 99.01 1.57 ;
        RECT 99.83 10.89 100 11.06 ;
        RECT 99.83 1.4 100 1.57 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 92.62 4.02 92.96 4.36 ;
      RECT 92.62 4.045 93.425 4.345 ;
      RECT 86.075 9.28 86.445 9.65 ;
      RECT 86.075 9.315 91.23 9.615 ;
      RECT 90.925 7.08 91.225 9.615 ;
      RECT 90.3 7.08 91.235 7.425 ;
      RECT 91.94 7.08 92.28 7.42 ;
      RECT 90.3 7.08 91.24 7.42 ;
      RECT 90.3 7.11 92.28 7.41 ;
      RECT 91.73 7.095 92.28 7.41 ;
      RECT 91.73 7.105 92.745 7.405 ;
      RECT 90.3 6.12 90.63 7.425 ;
      RECT 90.3 5.06 90.605 7.425 ;
      RECT 90.3 5.06 90.63 5.805 ;
      RECT 90.3 5.06 92.95 5.39 ;
      RECT 90.3 5.06 92.955 5.385 ;
      RECT 92.615 5.04 92.96 5.38 ;
      RECT 90.3 5.065 93.425 5.365 ;
      RECT 92.635 4.995 92.935 5.39 ;
      RECT 91.925 4.355 92.265 4.705 ;
      RECT 91.455 4.385 92.265 4.685 ;
      RECT 91.26 6.06 91.6 6.4 ;
      RECT 91.26 6.085 92.065 6.385 ;
      RECT 90.58 3.68 90.92 4.02 ;
      RECT 90.115 3.705 90.92 4.005 ;
      RECT 90.475 3.695 90.92 4.005 ;
      RECT 76.04 4.02 76.38 4.36 ;
      RECT 76.04 4.045 76.845 4.345 ;
      RECT 69.495 9.28 69.865 9.65 ;
      RECT 69.495 9.315 74.65 9.615 ;
      RECT 74.345 7.08 74.645 9.615 ;
      RECT 73.72 7.08 74.655 7.425 ;
      RECT 75.36 7.08 75.7 7.42 ;
      RECT 73.72 7.08 74.66 7.42 ;
      RECT 73.72 7.11 75.7 7.41 ;
      RECT 75.15 7.095 75.7 7.41 ;
      RECT 75.15 7.105 76.165 7.405 ;
      RECT 73.72 6.12 74.05 7.425 ;
      RECT 73.72 5.06 74.025 7.425 ;
      RECT 73.72 5.06 74.05 5.805 ;
      RECT 73.72 5.06 76.37 5.39 ;
      RECT 73.72 5.06 76.375 5.385 ;
      RECT 76.035 5.04 76.38 5.38 ;
      RECT 73.72 5.065 76.845 5.365 ;
      RECT 76.055 4.995 76.355 5.39 ;
      RECT 75.345 4.355 75.685 4.705 ;
      RECT 74.875 4.385 75.685 4.685 ;
      RECT 74.68 6.06 75.02 6.4 ;
      RECT 74.68 6.085 75.485 6.385 ;
      RECT 74 3.68 74.34 4.02 ;
      RECT 73.535 3.705 74.34 4.005 ;
      RECT 73.895 3.695 74.34 4.005 ;
      RECT 59.455 4.02 59.795 4.36 ;
      RECT 59.455 4.045 60.26 4.345 ;
      RECT 52.91 9.28 53.28 9.65 ;
      RECT 52.91 9.315 58.065 9.615 ;
      RECT 57.76 7.08 58.06 9.615 ;
      RECT 57.135 7.08 58.07 7.425 ;
      RECT 58.775 7.08 59.115 7.42 ;
      RECT 57.135 7.08 58.075 7.42 ;
      RECT 57.135 7.11 59.115 7.41 ;
      RECT 58.565 7.095 59.115 7.41 ;
      RECT 58.565 7.105 59.58 7.405 ;
      RECT 57.135 6.12 57.465 7.425 ;
      RECT 57.135 5.06 57.44 7.425 ;
      RECT 57.135 5.06 57.465 5.805 ;
      RECT 57.135 5.06 59.785 5.39 ;
      RECT 57.135 5.06 59.79 5.385 ;
      RECT 59.45 5.04 59.795 5.38 ;
      RECT 57.135 5.065 60.26 5.365 ;
      RECT 59.47 4.995 59.77 5.39 ;
      RECT 58.76 4.355 59.1 4.705 ;
      RECT 58.29 4.385 59.1 4.685 ;
      RECT 58.095 6.06 58.435 6.4 ;
      RECT 58.095 6.085 58.9 6.385 ;
      RECT 57.415 3.68 57.755 4.02 ;
      RECT 56.95 3.705 57.755 4.005 ;
      RECT 57.31 3.695 57.755 4.005 ;
      RECT 42.87 4.02 43.21 4.36 ;
      RECT 42.87 4.045 43.675 4.345 ;
      RECT 36.325 9.28 36.695 9.65 ;
      RECT 36.325 9.315 41.48 9.615 ;
      RECT 41.175 7.08 41.475 9.615 ;
      RECT 40.55 7.08 41.485 7.425 ;
      RECT 42.19 7.08 42.53 7.42 ;
      RECT 40.55 7.08 41.49 7.42 ;
      RECT 40.55 7.11 42.53 7.41 ;
      RECT 41.98 7.095 42.53 7.41 ;
      RECT 41.98 7.105 42.995 7.405 ;
      RECT 40.55 6.12 40.88 7.425 ;
      RECT 40.55 5.06 40.855 7.425 ;
      RECT 40.55 5.06 40.88 5.805 ;
      RECT 40.55 5.06 43.2 5.39 ;
      RECT 40.55 5.06 43.205 5.385 ;
      RECT 42.865 5.04 43.21 5.38 ;
      RECT 40.55 5.065 43.675 5.365 ;
      RECT 42.885 4.995 43.185 5.39 ;
      RECT 42.175 4.355 42.515 4.705 ;
      RECT 41.705 4.385 42.515 4.685 ;
      RECT 41.51 6.06 41.85 6.4 ;
      RECT 41.51 6.085 42.315 6.385 ;
      RECT 40.83 3.68 41.17 4.02 ;
      RECT 40.365 3.705 41.17 4.005 ;
      RECT 40.725 3.695 41.17 4.005 ;
      RECT 26.285 4.02 26.625 4.36 ;
      RECT 26.285 4.045 27.09 4.345 ;
      RECT 19.74 9.28 20.11 9.65 ;
      RECT 19.74 9.315 24.895 9.615 ;
      RECT 24.59 7.08 24.89 9.615 ;
      RECT 23.965 7.08 24.9 7.425 ;
      RECT 25.605 7.08 25.945 7.42 ;
      RECT 23.965 7.08 24.905 7.42 ;
      RECT 23.965 7.11 25.945 7.41 ;
      RECT 25.395 7.095 25.945 7.41 ;
      RECT 25.395 7.105 26.41 7.405 ;
      RECT 23.965 6.12 24.295 7.425 ;
      RECT 23.965 5.06 24.27 7.425 ;
      RECT 23.965 5.06 24.295 5.805 ;
      RECT 23.965 5.06 26.615 5.39 ;
      RECT 23.965 5.06 26.62 5.385 ;
      RECT 26.28 5.04 26.625 5.38 ;
      RECT 23.965 5.065 27.09 5.365 ;
      RECT 26.3 4.995 26.6 5.39 ;
      RECT 25.59 4.355 25.93 4.705 ;
      RECT 25.12 4.385 25.93 4.685 ;
      RECT 24.925 6.06 25.265 6.4 ;
      RECT 24.925 6.085 25.73 6.385 ;
      RECT 24.245 3.68 24.585 4.02 ;
      RECT 23.78 3.705 24.585 4.005 ;
      RECT 24.14 3.695 24.585 4.005 ;
      RECT 100.08 7.2 100.46 12.455 ;
      RECT 83.5 7.2 83.88 12.455 ;
      RECT 66.915 7.2 67.295 12.455 ;
      RECT 50.33 7.2 50.71 12.455 ;
      RECT 33.745 7.2 34.125 12.455 ;
    LAYER via2 ;
      RECT 100.17 7.29 100.37 7.49 ;
      RECT 92.695 4.095 92.895 4.295 ;
      RECT 92.695 5.115 92.895 5.315 ;
      RECT 92.015 7.155 92.215 7.355 ;
      RECT 91.995 4.435 92.195 4.635 ;
      RECT 91.335 6.135 91.535 6.335 ;
      RECT 90.965 7.155 91.165 7.355 ;
      RECT 90.655 3.745 90.855 3.945 ;
      RECT 86.16 9.365 86.36 9.565 ;
      RECT 83.59 7.29 83.79 7.49 ;
      RECT 76.115 4.095 76.315 4.295 ;
      RECT 76.115 5.115 76.315 5.315 ;
      RECT 75.435 7.155 75.635 7.355 ;
      RECT 75.415 4.435 75.615 4.635 ;
      RECT 74.755 6.135 74.955 6.335 ;
      RECT 74.385 7.155 74.585 7.355 ;
      RECT 74.075 3.745 74.275 3.945 ;
      RECT 69.58 9.365 69.78 9.565 ;
      RECT 67.005 7.29 67.205 7.49 ;
      RECT 59.53 4.095 59.73 4.295 ;
      RECT 59.53 5.115 59.73 5.315 ;
      RECT 58.85 7.155 59.05 7.355 ;
      RECT 58.83 4.435 59.03 4.635 ;
      RECT 58.17 6.135 58.37 6.335 ;
      RECT 57.8 7.155 58 7.355 ;
      RECT 57.49 3.745 57.69 3.945 ;
      RECT 52.995 9.365 53.195 9.565 ;
      RECT 50.42 7.29 50.62 7.49 ;
      RECT 42.945 4.095 43.145 4.295 ;
      RECT 42.945 5.115 43.145 5.315 ;
      RECT 42.265 7.155 42.465 7.355 ;
      RECT 42.245 4.435 42.445 4.635 ;
      RECT 41.585 6.135 41.785 6.335 ;
      RECT 41.215 7.155 41.415 7.355 ;
      RECT 40.905 3.745 41.105 3.945 ;
      RECT 36.41 9.365 36.61 9.565 ;
      RECT 33.835 7.29 34.035 7.49 ;
      RECT 26.36 4.095 26.56 4.295 ;
      RECT 26.36 5.115 26.56 5.315 ;
      RECT 25.68 7.155 25.88 7.355 ;
      RECT 25.66 4.435 25.86 4.635 ;
      RECT 25 6.135 25.2 6.335 ;
      RECT 24.63 7.155 24.83 7.355 ;
      RECT 24.32 3.745 24.52 3.945 ;
      RECT 19.825 9.365 20.025 9.565 ;
    LAYER met2 ;
      RECT 17.765 10.12 100.355 10.29 ;
      RECT 100.185 9.585 100.355 10.29 ;
      RECT 16.23 10.115 17.765 10.285 ;
      RECT 16.23 8.535 16.4 10.285 ;
      RECT 100.15 9.585 100.475 9.91 ;
      RECT 16.175 8.535 16.455 8.875 ;
      RECT 96.995 8.565 97.315 8.89 ;
      RECT 97.025 7.98 97.195 8.89 ;
      RECT 97.025 7.98 97.2 8.33 ;
      RECT 97.025 7.98 98 8.155 ;
      RECT 97.825 3.26 98 8.155 ;
      RECT 97.77 3.26 98.12 3.61 ;
      RECT 86.66 9.72 96.84 9.89 ;
      RECT 96.68 3.69 96.84 9.89 ;
      RECT 86.66 8.885 86.83 9.89 ;
      RECT 83.605 8.945 83.93 9.27 ;
      RECT 97.795 8.94 98.12 9.265 ;
      RECT 86.605 8.885 86.885 9.225 ;
      RECT 96.68 9.03 98.12 9.2 ;
      RECT 83.605 8.975 84.31 9.145 ;
      RECT 84.31 8.97 86.885 9.14 ;
      RECT 96.995 3.66 97.315 3.98 ;
      RECT 96.68 3.69 97.315 3.86 ;
      RECT 94.74 4.48 95.065 4.805 ;
      RECT 94.74 4.51 95.57 4.695 ;
      RECT 95.4 3.29 95.57 4.695 ;
      RECT 95.325 3.29 95.65 3.615 ;
      RECT 94.355 6.075 94.615 6.395 ;
      RECT 94.415 4.035 94.555 6.395 ;
      RECT 94.355 4.035 94.615 4.355 ;
      RECT 93.335 7.095 93.595 7.415 ;
      RECT 92.715 7.185 93.595 7.325 ;
      RECT 92.715 5.025 92.855 7.325 ;
      RECT 92.655 5.025 92.935 5.4 ;
      RECT 91.975 7.065 92.255 7.44 ;
      RECT 92.035 5.145 92.175 7.44 ;
      RECT 92.035 5.145 92.515 5.285 ;
      RECT 92.375 3.355 92.515 5.285 ;
      RECT 92.315 3.355 92.575 3.695 ;
      RECT 91.295 6.045 91.575 6.42 ;
      RECT 91.355 3.695 91.495 6.42 ;
      RECT 91.295 3.695 91.555 4.015 ;
      RECT 90.925 7.065 91.205 7.44 ;
      RECT 90.925 7.095 91.215 7.415 ;
      RECT 80.415 8.565 80.735 8.89 ;
      RECT 80.445 7.98 80.615 8.89 ;
      RECT 80.445 7.98 80.62 8.33 ;
      RECT 80.445 7.98 81.42 8.155 ;
      RECT 81.245 3.26 81.42 8.155 ;
      RECT 81.19 3.26 81.54 3.61 ;
      RECT 70.08 9.72 80.26 9.89 ;
      RECT 80.1 3.69 80.26 9.89 ;
      RECT 70.08 8.885 70.25 9.89 ;
      RECT 67.02 8.945 67.345 9.27 ;
      RECT 81.215 8.94 81.54 9.265 ;
      RECT 70.025 8.885 70.305 9.225 ;
      RECT 80.1 9.03 81.54 9.2 ;
      RECT 67.02 8.975 67.865 9.145 ;
      RECT 67.865 8.97 70.305 9.14 ;
      RECT 80.415 3.66 80.735 3.98 ;
      RECT 80.1 3.69 80.735 3.86 ;
      RECT 78.16 4.48 78.485 4.805 ;
      RECT 78.16 4.51 78.99 4.695 ;
      RECT 78.82 3.29 78.99 4.695 ;
      RECT 78.745 3.29 79.07 3.615 ;
      RECT 77.775 6.075 78.035 6.395 ;
      RECT 77.835 4.035 77.975 6.395 ;
      RECT 77.775 4.035 78.035 4.355 ;
      RECT 76.755 7.095 77.015 7.415 ;
      RECT 76.135 7.185 77.015 7.325 ;
      RECT 76.135 5.025 76.275 7.325 ;
      RECT 76.075 5.025 76.355 5.4 ;
      RECT 75.395 7.065 75.675 7.44 ;
      RECT 75.455 5.145 75.595 7.44 ;
      RECT 75.455 5.145 75.935 5.285 ;
      RECT 75.795 3.355 75.935 5.285 ;
      RECT 75.735 3.355 75.995 3.695 ;
      RECT 74.715 6.045 74.995 6.42 ;
      RECT 74.775 3.695 74.915 6.42 ;
      RECT 74.715 3.695 74.975 4.015 ;
      RECT 74.345 7.065 74.625 7.44 ;
      RECT 74.345 7.095 74.635 7.415 ;
      RECT 63.83 8.565 64.15 8.89 ;
      RECT 63.86 7.98 64.03 8.89 ;
      RECT 63.86 7.98 64.035 8.33 ;
      RECT 63.86 7.98 64.835 8.155 ;
      RECT 64.66 3.26 64.835 8.155 ;
      RECT 64.605 3.26 64.955 3.61 ;
      RECT 53.495 9.72 63.675 9.89 ;
      RECT 63.515 3.69 63.675 9.89 ;
      RECT 53.495 8.885 53.665 9.89 ;
      RECT 50.435 8.945 50.76 9.27 ;
      RECT 64.63 8.94 64.955 9.265 ;
      RECT 53.44 8.885 53.72 9.225 ;
      RECT 63.515 9.03 64.955 9.2 ;
      RECT 50.435 8.975 51.05 9.145 ;
      RECT 51.05 8.97 53.72 9.14 ;
      RECT 63.83 3.66 64.15 3.98 ;
      RECT 63.515 3.69 64.15 3.86 ;
      RECT 61.575 4.48 61.9 4.805 ;
      RECT 61.575 4.51 62.405 4.695 ;
      RECT 62.235 3.29 62.405 4.695 ;
      RECT 62.16 3.29 62.485 3.615 ;
      RECT 61.19 6.075 61.45 6.395 ;
      RECT 61.25 4.035 61.39 6.395 ;
      RECT 61.19 4.035 61.45 4.355 ;
      RECT 60.17 7.095 60.43 7.415 ;
      RECT 59.55 7.185 60.43 7.325 ;
      RECT 59.55 5.025 59.69 7.325 ;
      RECT 59.49 5.025 59.77 5.4 ;
      RECT 58.81 7.065 59.09 7.44 ;
      RECT 58.87 5.145 59.01 7.44 ;
      RECT 58.87 5.145 59.35 5.285 ;
      RECT 59.21 3.355 59.35 5.285 ;
      RECT 59.15 3.355 59.41 3.695 ;
      RECT 58.13 6.045 58.41 6.42 ;
      RECT 58.19 3.695 58.33 6.42 ;
      RECT 58.13 3.695 58.39 4.015 ;
      RECT 57.76 7.065 58.04 7.44 ;
      RECT 57.76 7.095 58.05 7.415 ;
      RECT 47.245 8.565 47.565 8.89 ;
      RECT 47.275 7.98 47.445 8.89 ;
      RECT 47.275 7.98 47.45 8.33 ;
      RECT 47.275 7.98 48.25 8.155 ;
      RECT 48.075 3.26 48.25 8.155 ;
      RECT 48.02 3.26 48.37 3.61 ;
      RECT 36.91 9.72 47.09 9.89 ;
      RECT 46.93 3.69 47.09 9.89 ;
      RECT 36.91 8.885 37.08 9.89 ;
      RECT 33.85 8.945 34.175 9.27 ;
      RECT 48.045 8.94 48.37 9.265 ;
      RECT 36.855 8.885 37.135 9.225 ;
      RECT 46.93 9.03 48.37 9.2 ;
      RECT 33.85 8.975 34.685 9.145 ;
      RECT 34.685 8.97 37.135 9.14 ;
      RECT 47.245 3.66 47.565 3.98 ;
      RECT 46.93 3.69 47.565 3.86 ;
      RECT 44.99 4.48 45.315 4.805 ;
      RECT 44.99 4.51 45.82 4.695 ;
      RECT 45.65 3.29 45.82 4.695 ;
      RECT 45.575 3.29 45.9 3.615 ;
      RECT 44.605 6.075 44.865 6.395 ;
      RECT 44.665 4.035 44.805 6.395 ;
      RECT 44.605 4.035 44.865 4.355 ;
      RECT 43.585 7.095 43.845 7.415 ;
      RECT 42.965 7.185 43.845 7.325 ;
      RECT 42.965 5.025 43.105 7.325 ;
      RECT 42.905 5.025 43.185 5.4 ;
      RECT 42.225 7.065 42.505 7.44 ;
      RECT 42.285 5.145 42.425 7.44 ;
      RECT 42.285 5.145 42.765 5.285 ;
      RECT 42.625 3.355 42.765 5.285 ;
      RECT 42.565 3.355 42.825 3.695 ;
      RECT 41.545 6.045 41.825 6.42 ;
      RECT 41.605 3.695 41.745 6.42 ;
      RECT 41.545 3.695 41.805 4.015 ;
      RECT 41.175 7.065 41.455 7.44 ;
      RECT 41.175 7.095 41.465 7.415 ;
      RECT 30.66 8.565 30.98 8.89 ;
      RECT 30.69 7.98 30.86 8.89 ;
      RECT 30.69 7.98 30.865 8.33 ;
      RECT 30.69 7.98 31.665 8.155 ;
      RECT 31.49 3.26 31.665 8.155 ;
      RECT 31.435 3.26 31.785 3.61 ;
      RECT 20.325 9.72 30.505 9.89 ;
      RECT 30.345 3.69 30.505 9.89 ;
      RECT 20.325 8.885 20.495 9.89 ;
      RECT 16.55 9.275 16.83 9.615 ;
      RECT 16.55 9.34 17.715 9.51 ;
      RECT 17.545 8.97 17.715 9.51 ;
      RECT 31.46 8.94 31.785 9.265 ;
      RECT 20.27 8.885 20.55 9.225 ;
      RECT 30.345 9.03 31.785 9.2 ;
      RECT 17.545 8.97 17.865 9.145 ;
      RECT 17.545 8.97 20.55 9.14 ;
      RECT 30.66 3.66 30.98 3.98 ;
      RECT 30.345 3.69 30.98 3.86 ;
      RECT 28.405 4.48 28.73 4.805 ;
      RECT 28.405 4.51 29.235 4.695 ;
      RECT 29.065 3.29 29.235 4.695 ;
      RECT 28.99 3.29 29.315 3.615 ;
      RECT 28.02 6.075 28.28 6.395 ;
      RECT 28.08 4.035 28.22 6.395 ;
      RECT 28.02 4.035 28.28 4.355 ;
      RECT 27 7.095 27.26 7.415 ;
      RECT 26.38 7.185 27.26 7.325 ;
      RECT 26.38 5.025 26.52 7.325 ;
      RECT 26.32 5.025 26.6 5.4 ;
      RECT 25.64 7.065 25.92 7.44 ;
      RECT 25.7 5.145 25.84 7.44 ;
      RECT 25.7 5.145 26.18 5.285 ;
      RECT 26.04 3.355 26.18 5.285 ;
      RECT 25.98 3.355 26.24 3.695 ;
      RECT 24.96 6.045 25.24 6.42 ;
      RECT 25.02 3.695 25.16 6.42 ;
      RECT 24.96 3.695 25.22 4.015 ;
      RECT 24.59 7.065 24.87 7.44 ;
      RECT 24.59 7.095 24.88 7.415 ;
      RECT 100.08 7.2 100.46 7.58 ;
      RECT 92.655 4.005 92.935 4.38 ;
      RECT 91.955 4.345 92.235 4.72 ;
      RECT 90.615 3.655 90.895 4.04 ;
      RECT 86.075 9.28 86.45 9.65 ;
      RECT 83.5 7.2 83.88 7.58 ;
      RECT 76.075 4.005 76.355 4.38 ;
      RECT 75.375 4.345 75.655 4.72 ;
      RECT 74.035 3.655 74.315 4.04 ;
      RECT 69.495 9.28 69.865 9.65 ;
      RECT 66.915 7.2 67.295 7.58 ;
      RECT 59.49 4.005 59.77 4.38 ;
      RECT 58.79 4.345 59.07 4.72 ;
      RECT 57.45 3.655 57.73 4.04 ;
      RECT 52.91 9.28 53.28 9.65 ;
      RECT 50.33 7.2 50.71 7.58 ;
      RECT 42.905 4.005 43.185 4.38 ;
      RECT 42.205 4.345 42.485 4.72 ;
      RECT 40.865 3.655 41.145 4.04 ;
      RECT 36.325 9.28 36.695 9.65 ;
      RECT 33.745 7.2 34.125 7.58 ;
      RECT 26.32 4.005 26.6 4.38 ;
      RECT 25.62 4.345 25.9 4.72 ;
      RECT 24.28 3.655 24.56 4.04 ;
      RECT 19.74 9.28 20.11 9.65 ;
    LAYER via1 ;
      RECT 100.24 9.67 100.39 9.82 ;
      RECT 100.195 7.315 100.345 7.465 ;
      RECT 97.885 9.025 98.035 9.175 ;
      RECT 97.87 3.36 98.02 3.51 ;
      RECT 97.08 3.745 97.23 3.895 ;
      RECT 97.08 8.655 97.23 8.805 ;
      RECT 95.415 3.375 95.565 3.525 ;
      RECT 94.83 4.565 94.98 4.715 ;
      RECT 94.41 4.12 94.56 4.27 ;
      RECT 94.41 6.16 94.56 6.31 ;
      RECT 93.39 7.18 93.54 7.33 ;
      RECT 92.71 4.12 92.86 4.27 ;
      RECT 92.71 5.14 92.86 5.29 ;
      RECT 92.37 3.46 92.52 3.61 ;
      RECT 92.03 4.46 92.18 4.61 ;
      RECT 92.03 7.18 92.18 7.33 ;
      RECT 91.35 3.78 91.5 3.93 ;
      RECT 91.35 6.16 91.5 6.31 ;
      RECT 91.01 7.18 91.16 7.33 ;
      RECT 90.67 3.77 90.82 3.92 ;
      RECT 86.67 8.98 86.82 9.13 ;
      RECT 86.185 9.39 86.335 9.54 ;
      RECT 83.695 9.03 83.845 9.18 ;
      RECT 83.615 7.315 83.765 7.465 ;
      RECT 81.305 9.025 81.455 9.175 ;
      RECT 81.29 3.36 81.44 3.51 ;
      RECT 80.5 3.745 80.65 3.895 ;
      RECT 80.5 8.655 80.65 8.805 ;
      RECT 78.835 3.375 78.985 3.525 ;
      RECT 78.25 4.565 78.4 4.715 ;
      RECT 77.83 4.12 77.98 4.27 ;
      RECT 77.83 6.16 77.98 6.31 ;
      RECT 76.81 7.18 76.96 7.33 ;
      RECT 76.13 4.12 76.28 4.27 ;
      RECT 76.13 5.14 76.28 5.29 ;
      RECT 75.79 3.46 75.94 3.61 ;
      RECT 75.45 4.46 75.6 4.61 ;
      RECT 75.45 7.18 75.6 7.33 ;
      RECT 74.77 3.78 74.92 3.93 ;
      RECT 74.77 6.16 74.92 6.31 ;
      RECT 74.43 7.18 74.58 7.33 ;
      RECT 74.09 3.77 74.24 3.92 ;
      RECT 70.09 8.98 70.24 9.13 ;
      RECT 69.605 9.39 69.755 9.54 ;
      RECT 67.11 9.03 67.26 9.18 ;
      RECT 67.03 7.315 67.18 7.465 ;
      RECT 64.72 9.025 64.87 9.175 ;
      RECT 64.705 3.36 64.855 3.51 ;
      RECT 63.915 3.745 64.065 3.895 ;
      RECT 63.915 8.655 64.065 8.805 ;
      RECT 62.25 3.375 62.4 3.525 ;
      RECT 61.665 4.565 61.815 4.715 ;
      RECT 61.245 4.12 61.395 4.27 ;
      RECT 61.245 6.16 61.395 6.31 ;
      RECT 60.225 7.18 60.375 7.33 ;
      RECT 59.545 4.12 59.695 4.27 ;
      RECT 59.545 5.14 59.695 5.29 ;
      RECT 59.205 3.46 59.355 3.61 ;
      RECT 58.865 4.46 59.015 4.61 ;
      RECT 58.865 7.18 59.015 7.33 ;
      RECT 58.185 3.78 58.335 3.93 ;
      RECT 58.185 6.16 58.335 6.31 ;
      RECT 57.845 7.18 57.995 7.33 ;
      RECT 57.505 3.77 57.655 3.92 ;
      RECT 53.505 8.98 53.655 9.13 ;
      RECT 53.02 9.39 53.17 9.54 ;
      RECT 50.525 9.03 50.675 9.18 ;
      RECT 50.445 7.315 50.595 7.465 ;
      RECT 48.135 9.025 48.285 9.175 ;
      RECT 48.12 3.36 48.27 3.51 ;
      RECT 47.33 3.745 47.48 3.895 ;
      RECT 47.33 8.655 47.48 8.805 ;
      RECT 45.665 3.375 45.815 3.525 ;
      RECT 45.08 4.565 45.23 4.715 ;
      RECT 44.66 4.12 44.81 4.27 ;
      RECT 44.66 6.16 44.81 6.31 ;
      RECT 43.64 7.18 43.79 7.33 ;
      RECT 42.96 4.12 43.11 4.27 ;
      RECT 42.96 5.14 43.11 5.29 ;
      RECT 42.62 3.46 42.77 3.61 ;
      RECT 42.28 4.46 42.43 4.61 ;
      RECT 42.28 7.18 42.43 7.33 ;
      RECT 41.6 3.78 41.75 3.93 ;
      RECT 41.6 6.16 41.75 6.31 ;
      RECT 41.26 7.18 41.41 7.33 ;
      RECT 40.92 3.77 41.07 3.92 ;
      RECT 36.92 8.98 37.07 9.13 ;
      RECT 36.435 9.39 36.585 9.54 ;
      RECT 33.94 9.03 34.09 9.18 ;
      RECT 33.86 7.315 34.01 7.465 ;
      RECT 31.55 9.025 31.7 9.175 ;
      RECT 31.535 3.36 31.685 3.51 ;
      RECT 30.745 3.745 30.895 3.895 ;
      RECT 30.745 8.655 30.895 8.805 ;
      RECT 29.08 3.375 29.23 3.525 ;
      RECT 28.495 4.565 28.645 4.715 ;
      RECT 28.075 4.12 28.225 4.27 ;
      RECT 28.075 6.16 28.225 6.31 ;
      RECT 27.055 7.18 27.205 7.33 ;
      RECT 26.375 4.12 26.525 4.27 ;
      RECT 26.375 5.14 26.525 5.29 ;
      RECT 26.035 3.46 26.185 3.61 ;
      RECT 25.695 4.46 25.845 4.61 ;
      RECT 25.695 7.18 25.845 7.33 ;
      RECT 25.015 3.78 25.165 3.93 ;
      RECT 25.015 6.16 25.165 6.31 ;
      RECT 24.675 7.18 24.825 7.33 ;
      RECT 24.335 3.77 24.485 3.92 ;
      RECT 20.335 8.98 20.485 9.13 ;
      RECT 19.85 9.39 20 9.54 ;
      RECT 16.615 9.37 16.765 9.52 ;
      RECT 16.24 8.63 16.39 8.78 ;
    LAYER met1 ;
      RECT 100.12 10.05 100.415 10.28 ;
      RECT 100.18 9.585 100.355 10.28 ;
      RECT 100.15 9.585 100.475 9.91 ;
      RECT 100.18 8.57 100.35 10.28 ;
      RECT 100.12 8.57 100.41 8.8 ;
      RECT 99.715 4.025 100.04 4.26 ;
      RECT 99.715 4.06 100.21 4.23 ;
      RECT 99.715 3.69 99.905 4.26 ;
      RECT 99.13 3.66 99.42 3.89 ;
      RECT 99.13 3.69 99.905 3.86 ;
      RECT 99.19 2.18 99.36 3.89 ;
      RECT 99.13 2.18 99.425 2.41 ;
      RECT 99.13 10.05 99.425 10.28 ;
      RECT 99.19 8.57 99.36 10.28 ;
      RECT 99.13 8.57 99.42 8.8 ;
      RECT 99.13 8.61 99.98 8.77 ;
      RECT 99.815 8.2 99.98 8.77 ;
      RECT 99.13 8.605 99.525 8.77 ;
      RECT 99.815 8.2 99.985 8.435 ;
      RECT 99.75 8.2 100.04 8.43 ;
      RECT 99.75 8.23 100.21 8.4 ;
      RECT 98.76 4.03 99.05 4.26 ;
      RECT 98.76 4.06 99.22 4.23 ;
      RECT 98.825 2.95 98.99 4.26 ;
      RECT 97.34 2.92 97.63 3.15 ;
      RECT 97.34 2.95 98.99 3.12 ;
      RECT 97.4 2.18 97.57 3.15 ;
      RECT 97.34 2.18 97.63 2.41 ;
      RECT 97.34 10.05 97.63 10.28 ;
      RECT 97.4 9.31 97.57 10.28 ;
      RECT 97.4 9.405 98.99 9.575 ;
      RECT 98.82 8.2 98.99 9.575 ;
      RECT 97.34 9.31 97.63 9.54 ;
      RECT 98.76 8.2 99.05 8.43 ;
      RECT 98.76 8.23 99.22 8.4 ;
      RECT 95.325 3.29 95.65 3.615 ;
      RECT 97.77 3.26 98.12 3.61 ;
      RECT 95.325 3.32 98.12 3.49 ;
      RECT 97.795 8.94 98.12 9.265 ;
      RECT 97.77 8.94 98.12 9.17 ;
      RECT 97.6 8.97 98.12 9.14 ;
      RECT 96.995 3.66 97.315 3.98 ;
      RECT 96.97 3.66 97.315 3.89 ;
      RECT 96.68 3.69 97.315 3.86 ;
      RECT 96.995 8.565 97.315 8.89 ;
      RECT 96.97 8.57 97.315 8.8 ;
      RECT 96.795 8.6 97.315 8.77 ;
      RECT 94.74 4.48 95.065 4.805 ;
      RECT 91.945 4.405 92.265 4.665 ;
      RECT 93.915 4.415 94.205 4.645 ;
      RECT 94.64 4.48 95.065 4.62 ;
      RECT 91.945 4.465 94.78 4.605 ;
      RECT 94.325 4.065 94.645 4.325 ;
      RECT 94.045 4.125 94.645 4.265 ;
      RECT 93.305 7.125 93.625 7.385 ;
      RECT 93.305 7.185 93.895 7.325 ;
      RECT 92.625 4.065 92.945 4.325 ;
      RECT 87.885 4.075 88.175 4.305 ;
      RECT 87.885 4.125 92.945 4.265 ;
      RECT 92.715 3.785 92.855 4.325 ;
      RECT 92.715 3.785 93.195 3.925 ;
      RECT 93.055 3.415 93.195 3.925 ;
      RECT 92.975 3.415 93.265 3.645 ;
      RECT 92.625 5.085 92.945 5.345 ;
      RECT 91.955 5.095 92.245 5.325 ;
      RECT 89.745 5.095 90.035 5.325 ;
      RECT 89.745 5.145 92.945 5.285 ;
      RECT 90.925 7.125 91.245 7.385 ;
      RECT 92.635 7.135 92.925 7.365 ;
      RECT 90.255 7.135 90.545 7.365 ;
      RECT 90.255 7.185 91.245 7.325 ;
      RECT 92.715 6.845 92.855 7.365 ;
      RECT 91.015 6.845 91.155 7.385 ;
      RECT 91.015 6.845 92.855 6.985 ;
      RECT 89.915 3.735 90.205 3.965 ;
      RECT 89.995 3.435 90.135 3.965 ;
      RECT 92.315 3.405 92.575 3.695 ;
      RECT 92.285 3.405 92.605 3.665 ;
      RECT 92.185 3.405 92.605 3.645 ;
      RECT 89.995 3.435 92.605 3.575 ;
      RECT 91.265 3.725 91.585 3.985 ;
      RECT 91.265 3.785 91.855 3.925 ;
      RECT 91.265 6.105 91.585 6.365 ;
      RECT 88.555 6.115 88.845 6.345 ;
      RECT 88.555 6.165 91.585 6.305 ;
      RECT 90.585 3.685 90.915 4.015 ;
      RECT 90.585 3.735 91.045 3.965 ;
      RECT 90.585 3.785 91.065 3.925 ;
      RECT 86.575 8.915 86.915 9.195 ;
      RECT 86.545 8.935 86.915 9.165 ;
      RECT 86.375 8.965 86.915 9.135 ;
      RECT 86.115 10.045 86.405 10.275 ;
      RECT 86.175 9.28 86.345 10.275 ;
      RECT 86.075 9.28 86.445 9.65 ;
      RECT 83.54 10.05 83.835 10.28 ;
      RECT 83.6 8.57 83.77 10.28 ;
      RECT 83.6 8.945 83.93 9.27 ;
      RECT 83.54 8.57 83.83 8.8 ;
      RECT 83.135 4.025 83.46 4.26 ;
      RECT 83.135 4.06 83.63 4.23 ;
      RECT 83.135 3.69 83.325 4.26 ;
      RECT 82.55 3.66 82.84 3.89 ;
      RECT 82.55 3.69 83.325 3.86 ;
      RECT 82.61 2.18 82.78 3.89 ;
      RECT 82.55 2.18 82.845 2.41 ;
      RECT 82.55 10.05 82.845 10.28 ;
      RECT 82.61 8.57 82.78 10.28 ;
      RECT 82.55 8.57 82.84 8.8 ;
      RECT 82.55 8.61 83.4 8.77 ;
      RECT 83.235 8.2 83.4 8.77 ;
      RECT 82.55 8.605 82.945 8.77 ;
      RECT 83.235 8.2 83.405 8.435 ;
      RECT 83.17 8.2 83.46 8.43 ;
      RECT 83.17 8.23 83.63 8.4 ;
      RECT 82.18 4.03 82.47 4.26 ;
      RECT 82.18 4.06 82.64 4.23 ;
      RECT 82.245 2.95 82.41 4.26 ;
      RECT 80.76 2.92 81.05 3.15 ;
      RECT 80.76 2.95 82.41 3.12 ;
      RECT 80.82 2.18 80.99 3.15 ;
      RECT 80.76 2.18 81.05 2.41 ;
      RECT 80.76 10.05 81.05 10.28 ;
      RECT 80.82 9.31 80.99 10.28 ;
      RECT 80.82 9.405 82.41 9.575 ;
      RECT 82.24 8.2 82.41 9.575 ;
      RECT 80.76 9.31 81.05 9.54 ;
      RECT 82.18 8.2 82.47 8.43 ;
      RECT 82.18 8.23 82.64 8.4 ;
      RECT 78.745 3.29 79.07 3.615 ;
      RECT 81.19 3.26 81.54 3.61 ;
      RECT 78.745 3.32 81.54 3.49 ;
      RECT 81.215 8.94 81.54 9.265 ;
      RECT 81.19 8.94 81.54 9.17 ;
      RECT 81.02 8.97 81.54 9.14 ;
      RECT 80.415 3.66 80.735 3.98 ;
      RECT 80.39 3.66 80.735 3.89 ;
      RECT 80.1 3.69 80.735 3.86 ;
      RECT 80.415 8.565 80.735 8.89 ;
      RECT 80.39 8.57 80.735 8.8 ;
      RECT 80.215 8.6 80.735 8.77 ;
      RECT 78.16 4.48 78.485 4.805 ;
      RECT 75.365 4.405 75.685 4.665 ;
      RECT 77.335 4.415 77.625 4.645 ;
      RECT 78.06 4.48 78.485 4.62 ;
      RECT 75.365 4.465 78.2 4.605 ;
      RECT 77.745 4.065 78.065 4.325 ;
      RECT 77.465 4.125 78.065 4.265 ;
      RECT 76.725 7.125 77.045 7.385 ;
      RECT 76.725 7.185 77.315 7.325 ;
      RECT 76.045 4.065 76.365 4.325 ;
      RECT 71.305 4.075 71.595 4.305 ;
      RECT 71.305 4.125 76.365 4.265 ;
      RECT 76.135 3.785 76.275 4.325 ;
      RECT 76.135 3.785 76.615 3.925 ;
      RECT 76.475 3.415 76.615 3.925 ;
      RECT 76.395 3.415 76.685 3.645 ;
      RECT 76.045 5.085 76.365 5.345 ;
      RECT 75.375 5.095 75.665 5.325 ;
      RECT 73.165 5.095 73.455 5.325 ;
      RECT 73.165 5.145 76.365 5.285 ;
      RECT 74.345 7.125 74.665 7.385 ;
      RECT 76.055 7.135 76.345 7.365 ;
      RECT 73.675 7.135 73.965 7.365 ;
      RECT 73.675 7.185 74.665 7.325 ;
      RECT 76.135 6.845 76.275 7.365 ;
      RECT 74.435 6.845 74.575 7.385 ;
      RECT 74.435 6.845 76.275 6.985 ;
      RECT 73.335 3.735 73.625 3.965 ;
      RECT 73.415 3.435 73.555 3.965 ;
      RECT 75.735 3.405 75.995 3.695 ;
      RECT 75.705 3.405 76.025 3.665 ;
      RECT 75.605 3.405 76.025 3.645 ;
      RECT 73.415 3.435 76.025 3.575 ;
      RECT 74.685 3.725 75.005 3.985 ;
      RECT 74.685 3.785 75.275 3.925 ;
      RECT 74.685 6.105 75.005 6.365 ;
      RECT 71.975 6.115 72.265 6.345 ;
      RECT 71.975 6.165 75.005 6.305 ;
      RECT 74.005 3.685 74.335 4.015 ;
      RECT 74.005 3.735 74.465 3.965 ;
      RECT 74.005 3.785 74.485 3.925 ;
      RECT 69.995 8.915 70.335 9.195 ;
      RECT 69.965 8.935 70.335 9.165 ;
      RECT 69.795 8.965 70.335 9.135 ;
      RECT 69.535 10.045 69.825 10.275 ;
      RECT 69.595 9.28 69.765 10.275 ;
      RECT 69.495 9.28 69.865 9.65 ;
      RECT 66.955 10.05 67.25 10.28 ;
      RECT 67.015 8.57 67.185 10.28 ;
      RECT 67.015 8.945 67.345 9.27 ;
      RECT 66.955 8.57 67.245 8.8 ;
      RECT 66.55 4.025 66.875 4.26 ;
      RECT 66.55 4.06 67.045 4.23 ;
      RECT 66.55 3.69 66.74 4.26 ;
      RECT 65.965 3.66 66.255 3.89 ;
      RECT 65.965 3.69 66.74 3.86 ;
      RECT 66.025 2.18 66.195 3.89 ;
      RECT 65.965 2.18 66.26 2.41 ;
      RECT 65.965 10.05 66.26 10.28 ;
      RECT 66.025 8.57 66.195 10.28 ;
      RECT 65.965 8.57 66.255 8.8 ;
      RECT 65.965 8.61 66.815 8.77 ;
      RECT 66.65 8.2 66.815 8.77 ;
      RECT 65.965 8.605 66.36 8.77 ;
      RECT 66.65 8.2 66.82 8.435 ;
      RECT 66.585 8.2 66.875 8.43 ;
      RECT 66.585 8.23 67.045 8.4 ;
      RECT 65.595 4.03 65.885 4.26 ;
      RECT 65.595 4.06 66.055 4.23 ;
      RECT 65.66 2.95 65.825 4.26 ;
      RECT 64.175 2.92 64.465 3.15 ;
      RECT 64.175 2.95 65.825 3.12 ;
      RECT 64.235 2.18 64.405 3.15 ;
      RECT 64.175 2.18 64.465 2.41 ;
      RECT 64.175 10.05 64.465 10.28 ;
      RECT 64.235 9.31 64.405 10.28 ;
      RECT 64.235 9.405 65.825 9.575 ;
      RECT 65.655 8.2 65.825 9.575 ;
      RECT 64.175 9.31 64.465 9.54 ;
      RECT 65.595 8.2 65.885 8.43 ;
      RECT 65.595 8.23 66.055 8.4 ;
      RECT 62.16 3.29 62.485 3.615 ;
      RECT 64.605 3.26 64.955 3.61 ;
      RECT 62.16 3.32 64.955 3.49 ;
      RECT 64.63 8.94 64.955 9.265 ;
      RECT 64.605 8.94 64.955 9.17 ;
      RECT 64.435 8.97 64.955 9.14 ;
      RECT 63.83 3.66 64.15 3.98 ;
      RECT 63.805 3.66 64.15 3.89 ;
      RECT 63.515 3.69 64.15 3.86 ;
      RECT 63.83 8.565 64.15 8.89 ;
      RECT 63.805 8.57 64.15 8.8 ;
      RECT 63.63 8.6 64.15 8.77 ;
      RECT 61.575 4.48 61.9 4.805 ;
      RECT 58.78 4.405 59.1 4.665 ;
      RECT 60.75 4.415 61.04 4.645 ;
      RECT 61.475 4.48 61.9 4.62 ;
      RECT 58.78 4.465 61.615 4.605 ;
      RECT 61.16 4.065 61.48 4.325 ;
      RECT 60.88 4.125 61.48 4.265 ;
      RECT 60.14 7.125 60.46 7.385 ;
      RECT 60.14 7.185 60.73 7.325 ;
      RECT 59.46 4.065 59.78 4.325 ;
      RECT 54.72 4.075 55.01 4.305 ;
      RECT 54.72 4.125 59.78 4.265 ;
      RECT 59.55 3.785 59.69 4.325 ;
      RECT 59.55 3.785 60.03 3.925 ;
      RECT 59.89 3.415 60.03 3.925 ;
      RECT 59.81 3.415 60.1 3.645 ;
      RECT 59.46 5.085 59.78 5.345 ;
      RECT 58.79 5.095 59.08 5.325 ;
      RECT 56.58 5.095 56.87 5.325 ;
      RECT 56.58 5.145 59.78 5.285 ;
      RECT 57.76 7.125 58.08 7.385 ;
      RECT 59.47 7.135 59.76 7.365 ;
      RECT 57.09 7.135 57.38 7.365 ;
      RECT 57.09 7.185 58.08 7.325 ;
      RECT 59.55 6.845 59.69 7.365 ;
      RECT 57.85 6.845 57.99 7.385 ;
      RECT 57.85 6.845 59.69 6.985 ;
      RECT 56.75 3.735 57.04 3.965 ;
      RECT 56.83 3.435 56.97 3.965 ;
      RECT 59.15 3.405 59.41 3.695 ;
      RECT 59.12 3.405 59.44 3.665 ;
      RECT 59.02 3.405 59.44 3.645 ;
      RECT 56.83 3.435 59.44 3.575 ;
      RECT 58.1 3.725 58.42 3.985 ;
      RECT 58.1 3.785 58.69 3.925 ;
      RECT 58.1 6.105 58.42 6.365 ;
      RECT 55.39 6.115 55.68 6.345 ;
      RECT 55.39 6.165 58.42 6.305 ;
      RECT 57.42 3.685 57.75 4.015 ;
      RECT 57.42 3.735 57.88 3.965 ;
      RECT 57.42 3.785 57.9 3.925 ;
      RECT 53.41 8.915 53.75 9.195 ;
      RECT 53.38 8.935 53.75 9.165 ;
      RECT 53.21 8.965 53.75 9.135 ;
      RECT 52.95 10.045 53.24 10.275 ;
      RECT 53.01 9.28 53.18 10.275 ;
      RECT 52.91 9.28 53.28 9.65 ;
      RECT 50.37 10.05 50.665 10.28 ;
      RECT 50.43 8.57 50.6 10.28 ;
      RECT 50.43 8.945 50.76 9.27 ;
      RECT 50.37 8.57 50.66 8.8 ;
      RECT 49.965 4.025 50.29 4.26 ;
      RECT 49.965 4.06 50.46 4.23 ;
      RECT 49.965 3.69 50.155 4.26 ;
      RECT 49.38 3.66 49.67 3.89 ;
      RECT 49.38 3.69 50.155 3.86 ;
      RECT 49.44 2.18 49.61 3.89 ;
      RECT 49.38 2.18 49.675 2.41 ;
      RECT 49.38 10.05 49.675 10.28 ;
      RECT 49.44 8.57 49.61 10.28 ;
      RECT 49.38 8.57 49.67 8.8 ;
      RECT 49.38 8.61 50.23 8.77 ;
      RECT 50.065 8.2 50.23 8.77 ;
      RECT 49.38 8.605 49.775 8.77 ;
      RECT 50.065 8.2 50.235 8.435 ;
      RECT 50 8.2 50.29 8.43 ;
      RECT 50 8.23 50.46 8.4 ;
      RECT 49.01 4.03 49.3 4.26 ;
      RECT 49.01 4.06 49.47 4.23 ;
      RECT 49.075 2.95 49.24 4.26 ;
      RECT 47.59 2.92 47.88 3.15 ;
      RECT 47.59 2.95 49.24 3.12 ;
      RECT 47.65 2.18 47.82 3.15 ;
      RECT 47.59 2.18 47.88 2.41 ;
      RECT 47.59 10.05 47.88 10.28 ;
      RECT 47.65 9.31 47.82 10.28 ;
      RECT 47.65 9.405 49.24 9.575 ;
      RECT 49.07 8.2 49.24 9.575 ;
      RECT 47.59 9.31 47.88 9.54 ;
      RECT 49.01 8.2 49.3 8.43 ;
      RECT 49.01 8.23 49.47 8.4 ;
      RECT 45.575 3.29 45.9 3.615 ;
      RECT 48.02 3.26 48.37 3.61 ;
      RECT 45.575 3.32 48.37 3.49 ;
      RECT 48.045 8.94 48.37 9.265 ;
      RECT 48.02 8.94 48.37 9.17 ;
      RECT 47.85 8.97 48.37 9.14 ;
      RECT 47.245 3.66 47.565 3.98 ;
      RECT 47.22 3.66 47.565 3.89 ;
      RECT 46.93 3.69 47.565 3.86 ;
      RECT 47.245 8.565 47.565 8.89 ;
      RECT 47.22 8.57 47.565 8.8 ;
      RECT 47.045 8.6 47.565 8.77 ;
      RECT 44.99 4.48 45.315 4.805 ;
      RECT 42.195 4.405 42.515 4.665 ;
      RECT 44.165 4.415 44.455 4.645 ;
      RECT 44.89 4.48 45.315 4.62 ;
      RECT 42.195 4.465 45.03 4.605 ;
      RECT 44.575 4.065 44.895 4.325 ;
      RECT 44.295 4.125 44.895 4.265 ;
      RECT 43.555 7.125 43.875 7.385 ;
      RECT 43.555 7.185 44.145 7.325 ;
      RECT 42.875 4.065 43.195 4.325 ;
      RECT 38.135 4.075 38.425 4.305 ;
      RECT 38.135 4.125 43.195 4.265 ;
      RECT 42.965 3.785 43.105 4.325 ;
      RECT 42.965 3.785 43.445 3.925 ;
      RECT 43.305 3.415 43.445 3.925 ;
      RECT 43.225 3.415 43.515 3.645 ;
      RECT 42.875 5.085 43.195 5.345 ;
      RECT 42.205 5.095 42.495 5.325 ;
      RECT 39.995 5.095 40.285 5.325 ;
      RECT 39.995 5.145 43.195 5.285 ;
      RECT 41.175 7.125 41.495 7.385 ;
      RECT 42.885 7.135 43.175 7.365 ;
      RECT 40.505 7.135 40.795 7.365 ;
      RECT 40.505 7.185 41.495 7.325 ;
      RECT 42.965 6.845 43.105 7.365 ;
      RECT 41.265 6.845 41.405 7.385 ;
      RECT 41.265 6.845 43.105 6.985 ;
      RECT 40.165 3.735 40.455 3.965 ;
      RECT 40.245 3.435 40.385 3.965 ;
      RECT 42.565 3.405 42.825 3.695 ;
      RECT 42.535 3.405 42.855 3.665 ;
      RECT 42.435 3.405 42.855 3.645 ;
      RECT 40.245 3.435 42.855 3.575 ;
      RECT 41.515 3.725 41.835 3.985 ;
      RECT 41.515 3.785 42.105 3.925 ;
      RECT 41.515 6.105 41.835 6.365 ;
      RECT 38.805 6.115 39.095 6.345 ;
      RECT 38.805 6.165 41.835 6.305 ;
      RECT 40.835 3.685 41.165 4.015 ;
      RECT 40.835 3.735 41.295 3.965 ;
      RECT 40.835 3.785 41.315 3.925 ;
      RECT 36.825 8.915 37.165 9.195 ;
      RECT 36.795 8.935 37.165 9.165 ;
      RECT 36.625 8.965 37.165 9.135 ;
      RECT 36.365 10.045 36.655 10.275 ;
      RECT 36.425 9.28 36.595 10.275 ;
      RECT 36.325 9.28 36.695 9.65 ;
      RECT 33.785 10.05 34.08 10.28 ;
      RECT 33.845 8.57 34.015 10.28 ;
      RECT 33.845 8.945 34.175 9.27 ;
      RECT 33.785 8.57 34.075 8.8 ;
      RECT 33.38 4.025 33.705 4.26 ;
      RECT 33.38 4.06 33.875 4.23 ;
      RECT 33.38 3.69 33.57 4.26 ;
      RECT 32.795 3.66 33.085 3.89 ;
      RECT 32.795 3.69 33.57 3.86 ;
      RECT 32.855 2.18 33.025 3.89 ;
      RECT 32.795 2.18 33.09 2.41 ;
      RECT 32.795 10.05 33.09 10.28 ;
      RECT 32.855 8.57 33.025 10.28 ;
      RECT 32.795 8.57 33.085 8.8 ;
      RECT 32.795 8.61 33.645 8.77 ;
      RECT 33.48 8.2 33.645 8.77 ;
      RECT 32.795 8.605 33.19 8.77 ;
      RECT 33.48 8.2 33.65 8.435 ;
      RECT 33.415 8.2 33.705 8.43 ;
      RECT 33.415 8.23 33.875 8.4 ;
      RECT 32.425 4.03 32.715 4.26 ;
      RECT 32.425 4.06 32.885 4.23 ;
      RECT 32.49 2.95 32.655 4.26 ;
      RECT 31.005 2.92 31.295 3.15 ;
      RECT 31.005 2.95 32.655 3.12 ;
      RECT 31.065 2.18 31.235 3.15 ;
      RECT 31.005 2.18 31.295 2.41 ;
      RECT 31.005 10.05 31.295 10.28 ;
      RECT 31.065 9.31 31.235 10.28 ;
      RECT 31.065 9.405 32.655 9.575 ;
      RECT 32.485 8.2 32.655 9.575 ;
      RECT 31.005 9.31 31.295 9.54 ;
      RECT 32.425 8.2 32.715 8.43 ;
      RECT 32.425 8.23 32.885 8.4 ;
      RECT 28.99 3.29 29.315 3.615 ;
      RECT 31.435 3.26 31.785 3.61 ;
      RECT 28.99 3.32 31.785 3.49 ;
      RECT 31.46 8.94 31.785 9.265 ;
      RECT 31.435 8.94 31.785 9.17 ;
      RECT 31.265 8.97 31.785 9.14 ;
      RECT 30.66 3.66 30.98 3.98 ;
      RECT 30.635 3.66 30.98 3.89 ;
      RECT 30.345 3.69 30.98 3.86 ;
      RECT 30.66 8.565 30.98 8.89 ;
      RECT 30.635 8.57 30.98 8.8 ;
      RECT 30.46 8.6 30.98 8.77 ;
      RECT 28.405 4.48 28.73 4.805 ;
      RECT 25.61 4.405 25.93 4.665 ;
      RECT 27.58 4.415 27.87 4.645 ;
      RECT 28.305 4.48 28.73 4.62 ;
      RECT 25.61 4.465 28.445 4.605 ;
      RECT 27.99 4.065 28.31 4.325 ;
      RECT 27.71 4.125 28.31 4.265 ;
      RECT 26.97 7.125 27.29 7.385 ;
      RECT 26.97 7.185 27.56 7.325 ;
      RECT 26.29 4.065 26.61 4.325 ;
      RECT 21.55 4.075 21.84 4.305 ;
      RECT 21.55 4.125 26.61 4.265 ;
      RECT 26.38 3.785 26.52 4.325 ;
      RECT 26.38 3.785 26.86 3.925 ;
      RECT 26.72 3.415 26.86 3.925 ;
      RECT 26.64 3.415 26.93 3.645 ;
      RECT 26.29 5.085 26.61 5.345 ;
      RECT 25.62 5.095 25.91 5.325 ;
      RECT 23.41 5.095 23.7 5.325 ;
      RECT 23.41 5.145 26.61 5.285 ;
      RECT 24.59 7.125 24.91 7.385 ;
      RECT 26.3 7.135 26.59 7.365 ;
      RECT 23.92 7.135 24.21 7.365 ;
      RECT 23.92 7.185 24.91 7.325 ;
      RECT 26.38 6.845 26.52 7.365 ;
      RECT 24.68 6.845 24.82 7.385 ;
      RECT 24.68 6.845 26.52 6.985 ;
      RECT 23.58 3.735 23.87 3.965 ;
      RECT 23.66 3.435 23.8 3.965 ;
      RECT 25.98 3.405 26.24 3.695 ;
      RECT 25.95 3.405 26.27 3.665 ;
      RECT 25.85 3.405 26.27 3.645 ;
      RECT 23.66 3.435 26.27 3.575 ;
      RECT 24.93 3.725 25.25 3.985 ;
      RECT 24.93 3.785 25.52 3.925 ;
      RECT 24.93 6.105 25.25 6.365 ;
      RECT 22.22 6.115 22.51 6.345 ;
      RECT 22.22 6.165 25.25 6.305 ;
      RECT 24.25 3.685 24.58 4.015 ;
      RECT 24.25 3.735 24.71 3.965 ;
      RECT 24.25 3.785 24.73 3.925 ;
      RECT 20.24 8.915 20.58 9.195 ;
      RECT 20.21 8.935 20.58 9.165 ;
      RECT 20.04 8.965 20.58 9.135 ;
      RECT 19.78 10.045 20.07 10.275 ;
      RECT 19.84 9.28 20.01 10.275 ;
      RECT 19.74 9.28 20.11 9.65 ;
      RECT 16.55 10.045 16.84 10.275 ;
      RECT 16.61 9.305 16.78 10.275 ;
      RECT 16.52 9.305 16.86 9.585 ;
      RECT 16.145 8.565 16.485 8.845 ;
      RECT 16.005 8.595 16.485 8.765 ;
      RECT 100.095 7.245 100.445 7.535 ;
      RECT 93.995 6.105 94.645 6.365 ;
      RECT 91.945 7.125 92.265 7.385 ;
      RECT 83.515 7.245 83.865 7.535 ;
      RECT 77.415 6.105 78.065 6.365 ;
      RECT 75.365 7.125 75.685 7.385 ;
      RECT 66.93 7.245 67.28 7.535 ;
      RECT 60.83 6.105 61.48 6.365 ;
      RECT 58.78 7.125 59.1 7.385 ;
      RECT 50.345 7.245 50.695 7.535 ;
      RECT 44.245 6.105 44.895 6.365 ;
      RECT 42.195 7.125 42.515 7.385 ;
      RECT 33.76 7.245 34.11 7.535 ;
      RECT 27.66 6.105 28.31 6.365 ;
      RECT 25.61 7.125 25.93 7.385 ;
    LAYER mcon ;
      RECT 100.185 7.305 100.355 7.475 ;
      RECT 100.18 8.6 100.35 8.77 ;
      RECT 100.18 10.08 100.35 10.25 ;
      RECT 99.81 4.06 99.98 4.23 ;
      RECT 99.81 8.23 99.98 8.4 ;
      RECT 99.19 2.21 99.36 2.38 ;
      RECT 99.19 3.69 99.36 3.86 ;
      RECT 99.19 8.6 99.36 8.77 ;
      RECT 99.19 10.08 99.36 10.25 ;
      RECT 98.82 4.06 98.99 4.23 ;
      RECT 98.82 8.23 98.99 8.4 ;
      RECT 97.83 3.32 98 3.49 ;
      RECT 97.83 8.97 98 9.14 ;
      RECT 97.4 2.21 97.57 2.38 ;
      RECT 97.4 2.95 97.57 3.12 ;
      RECT 97.4 9.34 97.57 9.51 ;
      RECT 97.4 10.08 97.57 10.25 ;
      RECT 97.03 3.69 97.2 3.86 ;
      RECT 97.03 8.6 97.2 8.77 ;
      RECT 94.395 4.105 94.565 4.275 ;
      RECT 94.055 6.145 94.225 6.315 ;
      RECT 93.975 4.445 94.145 4.615 ;
      RECT 93.375 7.165 93.545 7.335 ;
      RECT 93.035 3.445 93.205 3.615 ;
      RECT 92.695 7.165 92.865 7.335 ;
      RECT 92.245 3.435 92.415 3.605 ;
      RECT 92.015 5.125 92.185 5.295 ;
      RECT 92.015 7.165 92.185 7.335 ;
      RECT 91.335 3.765 91.505 3.935 ;
      RECT 90.815 3.765 90.985 3.935 ;
      RECT 90.315 7.165 90.485 7.335 ;
      RECT 89.975 3.765 90.145 3.935 ;
      RECT 89.805 5.125 89.975 5.295 ;
      RECT 88.615 6.145 88.785 6.315 ;
      RECT 87.945 4.105 88.115 4.275 ;
      RECT 86.605 8.965 86.775 9.135 ;
      RECT 86.175 9.335 86.345 9.505 ;
      RECT 86.175 10.075 86.345 10.245 ;
      RECT 83.605 7.305 83.775 7.475 ;
      RECT 83.6 8.6 83.77 8.77 ;
      RECT 83.6 10.08 83.77 10.25 ;
      RECT 83.23 4.06 83.4 4.23 ;
      RECT 83.23 8.23 83.4 8.4 ;
      RECT 82.61 2.21 82.78 2.38 ;
      RECT 82.61 3.69 82.78 3.86 ;
      RECT 82.61 8.6 82.78 8.77 ;
      RECT 82.61 10.08 82.78 10.25 ;
      RECT 82.24 4.06 82.41 4.23 ;
      RECT 82.24 8.23 82.41 8.4 ;
      RECT 81.25 3.32 81.42 3.49 ;
      RECT 81.25 8.97 81.42 9.14 ;
      RECT 80.82 2.21 80.99 2.38 ;
      RECT 80.82 2.95 80.99 3.12 ;
      RECT 80.82 9.34 80.99 9.51 ;
      RECT 80.82 10.08 80.99 10.25 ;
      RECT 80.45 3.69 80.62 3.86 ;
      RECT 80.45 8.6 80.62 8.77 ;
      RECT 77.815 4.105 77.985 4.275 ;
      RECT 77.475 6.145 77.645 6.315 ;
      RECT 77.395 4.445 77.565 4.615 ;
      RECT 76.795 7.165 76.965 7.335 ;
      RECT 76.455 3.445 76.625 3.615 ;
      RECT 76.115 7.165 76.285 7.335 ;
      RECT 75.665 3.435 75.835 3.605 ;
      RECT 75.435 5.125 75.605 5.295 ;
      RECT 75.435 7.165 75.605 7.335 ;
      RECT 74.755 3.765 74.925 3.935 ;
      RECT 74.235 3.765 74.405 3.935 ;
      RECT 73.735 7.165 73.905 7.335 ;
      RECT 73.395 3.765 73.565 3.935 ;
      RECT 73.225 5.125 73.395 5.295 ;
      RECT 72.035 6.145 72.205 6.315 ;
      RECT 71.365 4.105 71.535 4.275 ;
      RECT 70.025 8.965 70.195 9.135 ;
      RECT 69.595 9.335 69.765 9.505 ;
      RECT 69.595 10.075 69.765 10.245 ;
      RECT 67.02 7.305 67.19 7.475 ;
      RECT 67.015 8.6 67.185 8.77 ;
      RECT 67.015 10.08 67.185 10.25 ;
      RECT 66.645 4.06 66.815 4.23 ;
      RECT 66.645 8.23 66.815 8.4 ;
      RECT 66.025 2.21 66.195 2.38 ;
      RECT 66.025 3.69 66.195 3.86 ;
      RECT 66.025 8.6 66.195 8.77 ;
      RECT 66.025 10.08 66.195 10.25 ;
      RECT 65.655 4.06 65.825 4.23 ;
      RECT 65.655 8.23 65.825 8.4 ;
      RECT 64.665 3.32 64.835 3.49 ;
      RECT 64.665 8.97 64.835 9.14 ;
      RECT 64.235 2.21 64.405 2.38 ;
      RECT 64.235 2.95 64.405 3.12 ;
      RECT 64.235 9.34 64.405 9.51 ;
      RECT 64.235 10.08 64.405 10.25 ;
      RECT 63.865 3.69 64.035 3.86 ;
      RECT 63.865 8.6 64.035 8.77 ;
      RECT 61.23 4.105 61.4 4.275 ;
      RECT 60.89 6.145 61.06 6.315 ;
      RECT 60.81 4.445 60.98 4.615 ;
      RECT 60.21 7.165 60.38 7.335 ;
      RECT 59.87 3.445 60.04 3.615 ;
      RECT 59.53 7.165 59.7 7.335 ;
      RECT 59.08 3.435 59.25 3.605 ;
      RECT 58.85 5.125 59.02 5.295 ;
      RECT 58.85 7.165 59.02 7.335 ;
      RECT 58.17 3.765 58.34 3.935 ;
      RECT 57.65 3.765 57.82 3.935 ;
      RECT 57.15 7.165 57.32 7.335 ;
      RECT 56.81 3.765 56.98 3.935 ;
      RECT 56.64 5.125 56.81 5.295 ;
      RECT 55.45 6.145 55.62 6.315 ;
      RECT 54.78 4.105 54.95 4.275 ;
      RECT 53.44 8.965 53.61 9.135 ;
      RECT 53.01 9.335 53.18 9.505 ;
      RECT 53.01 10.075 53.18 10.245 ;
      RECT 50.435 7.305 50.605 7.475 ;
      RECT 50.43 8.6 50.6 8.77 ;
      RECT 50.43 10.08 50.6 10.25 ;
      RECT 50.06 4.06 50.23 4.23 ;
      RECT 50.06 8.23 50.23 8.4 ;
      RECT 49.44 2.21 49.61 2.38 ;
      RECT 49.44 3.69 49.61 3.86 ;
      RECT 49.44 8.6 49.61 8.77 ;
      RECT 49.44 10.08 49.61 10.25 ;
      RECT 49.07 4.06 49.24 4.23 ;
      RECT 49.07 8.23 49.24 8.4 ;
      RECT 48.08 3.32 48.25 3.49 ;
      RECT 48.08 8.97 48.25 9.14 ;
      RECT 47.65 2.21 47.82 2.38 ;
      RECT 47.65 2.95 47.82 3.12 ;
      RECT 47.65 9.34 47.82 9.51 ;
      RECT 47.65 10.08 47.82 10.25 ;
      RECT 47.28 3.69 47.45 3.86 ;
      RECT 47.28 8.6 47.45 8.77 ;
      RECT 44.645 4.105 44.815 4.275 ;
      RECT 44.305 6.145 44.475 6.315 ;
      RECT 44.225 4.445 44.395 4.615 ;
      RECT 43.625 7.165 43.795 7.335 ;
      RECT 43.285 3.445 43.455 3.615 ;
      RECT 42.945 7.165 43.115 7.335 ;
      RECT 42.495 3.435 42.665 3.605 ;
      RECT 42.265 5.125 42.435 5.295 ;
      RECT 42.265 7.165 42.435 7.335 ;
      RECT 41.585 3.765 41.755 3.935 ;
      RECT 41.065 3.765 41.235 3.935 ;
      RECT 40.565 7.165 40.735 7.335 ;
      RECT 40.225 3.765 40.395 3.935 ;
      RECT 40.055 5.125 40.225 5.295 ;
      RECT 38.865 6.145 39.035 6.315 ;
      RECT 38.195 4.105 38.365 4.275 ;
      RECT 36.855 8.965 37.025 9.135 ;
      RECT 36.425 9.335 36.595 9.505 ;
      RECT 36.425 10.075 36.595 10.245 ;
      RECT 33.85 7.305 34.02 7.475 ;
      RECT 33.845 8.6 34.015 8.77 ;
      RECT 33.845 10.08 34.015 10.25 ;
      RECT 33.475 4.06 33.645 4.23 ;
      RECT 33.475 8.23 33.645 8.4 ;
      RECT 32.855 2.21 33.025 2.38 ;
      RECT 32.855 3.69 33.025 3.86 ;
      RECT 32.855 8.6 33.025 8.77 ;
      RECT 32.855 10.08 33.025 10.25 ;
      RECT 32.485 4.06 32.655 4.23 ;
      RECT 32.485 8.23 32.655 8.4 ;
      RECT 31.495 3.32 31.665 3.49 ;
      RECT 31.495 8.97 31.665 9.14 ;
      RECT 31.065 2.21 31.235 2.38 ;
      RECT 31.065 2.95 31.235 3.12 ;
      RECT 31.065 9.34 31.235 9.51 ;
      RECT 31.065 10.08 31.235 10.25 ;
      RECT 30.695 3.69 30.865 3.86 ;
      RECT 30.695 8.6 30.865 8.77 ;
      RECT 28.06 4.105 28.23 4.275 ;
      RECT 27.72 6.145 27.89 6.315 ;
      RECT 27.64 4.445 27.81 4.615 ;
      RECT 27.04 7.165 27.21 7.335 ;
      RECT 26.7 3.445 26.87 3.615 ;
      RECT 26.36 7.165 26.53 7.335 ;
      RECT 25.91 3.435 26.08 3.605 ;
      RECT 25.68 5.125 25.85 5.295 ;
      RECT 25.68 7.165 25.85 7.335 ;
      RECT 25 3.765 25.17 3.935 ;
      RECT 24.48 3.765 24.65 3.935 ;
      RECT 23.98 7.165 24.15 7.335 ;
      RECT 23.64 3.765 23.81 3.935 ;
      RECT 23.47 5.125 23.64 5.295 ;
      RECT 22.28 6.145 22.45 6.315 ;
      RECT 21.61 4.105 21.78 4.275 ;
      RECT 20.27 8.965 20.44 9.135 ;
      RECT 19.84 9.335 20.01 9.505 ;
      RECT 19.84 10.075 20.01 10.245 ;
      RECT 16.61 9.335 16.78 9.505 ;
      RECT 16.61 10.075 16.78 10.245 ;
      RECT 16.24 8.595 16.41 8.765 ;
    LAYER li1 ;
      RECT 100.18 7.3 100.35 8.77 ;
      RECT 100.18 7.3 100.355 8.56 ;
      RECT 99.81 3.04 99.98 4.23 ;
      RECT 99.81 3.04 100.28 3.21 ;
      RECT 99.81 9.25 100.28 9.42 ;
      RECT 99.81 8.23 99.98 9.42 ;
      RECT 99.19 3.9 99.365 5.16 ;
      RECT 99.19 3.69 99.36 5.16 ;
      RECT 99.19 7.3 99.36 8.77 ;
      RECT 99.19 7.3 99.365 8.56 ;
      RECT 98.82 3.04 98.99 4.23 ;
      RECT 98.82 3.04 99.29 3.21 ;
      RECT 98.82 9.25 99.29 9.42 ;
      RECT 98.82 8.23 98.99 9.42 ;
      RECT 97.83 4.02 98.005 5.16 ;
      RECT 97.83 1.87 98 5.16 ;
      RECT 97.83 1.87 98.005 2.42 ;
      RECT 97.83 10.04 98.005 10.59 ;
      RECT 97.83 7.3 98 10.59 ;
      RECT 97.83 7.3 98.005 8.44 ;
      RECT 97.4 3.9 97.575 5.16 ;
      RECT 97.4 2.95 97.57 5.16 ;
      RECT 97.4 7.3 97.57 9.51 ;
      RECT 97.4 7.3 97.575 8.56 ;
      RECT 96.97 3.93 97.14 5.16 ;
      RECT 97.03 2.15 97.2 4.1 ;
      RECT 96.97 1.87 97.14 2.32 ;
      RECT 96.97 10.14 97.14 10.59 ;
      RECT 97.03 8.36 97.2 10.31 ;
      RECT 96.97 7.3 97.14 8.53 ;
      RECT 96.445 3.9 96.62 5.16 ;
      RECT 96.445 1.87 96.615 5.16 ;
      RECT 96.445 3.37 96.855 3.7 ;
      RECT 96.445 2.53 96.855 2.86 ;
      RECT 96.445 1.87 96.62 2.36 ;
      RECT 96.445 10.1 96.62 10.59 ;
      RECT 96.445 7.3 96.615 10.59 ;
      RECT 96.445 9.6 96.855 9.93 ;
      RECT 96.445 8.76 96.855 9.09 ;
      RECT 96.445 7.3 96.62 8.56 ;
      RECT 91.705 7.935 93.015 8.185 ;
      RECT 91.705 7.615 91.885 8.185 ;
      RECT 91.155 7.615 91.885 7.785 ;
      RECT 91.155 6.775 91.325 7.785 ;
      RECT 91.995 6.815 93.735 6.995 ;
      RECT 93.405 5.975 93.735 6.995 ;
      RECT 91.155 6.775 92.215 6.945 ;
      RECT 93.405 6.145 94.225 6.315 ;
      RECT 92.565 5.975 92.895 6.185 ;
      RECT 92.565 5.975 93.735 6.145 ;
      RECT 93.465 4.495 93.795 5.455 ;
      RECT 93.465 4.495 94.145 4.665 ;
      RECT 93.975 3.265 94.145 4.665 ;
      RECT 93.885 3.265 94.215 3.895 ;
      RECT 93.015 4.765 93.285 5.465 ;
      RECT 93.115 3.265 93.285 5.465 ;
      RECT 93.455 4.075 93.805 4.325 ;
      RECT 93.115 4.105 93.805 4.275 ;
      RECT 93.025 3.265 93.285 3.735 ;
      RECT 92.355 6.405 93.235 6.645 ;
      RECT 93.005 6.315 93.235 6.645 ;
      RECT 91.705 6.405 93.235 6.605 ;
      RECT 92.625 6.355 93.235 6.645 ;
      RECT 91.705 6.275 91.875 6.605 ;
      RECT 92.595 7.165 92.845 7.765 ;
      RECT 92.595 7.165 93.065 7.365 ;
      RECT 92.085 4.385 92.845 4.885 ;
      RECT 91.155 4.195 91.415 4.815 ;
      RECT 92.075 4.325 92.085 4.635 ;
      RECT 92.055 4.385 92.845 4.605 ;
      RECT 92.715 3.995 92.945 4.595 ;
      RECT 92.035 4.315 92.075 4.575 ;
      RECT 92.015 4.385 92.945 4.565 ;
      RECT 91.985 4.385 92.945 4.555 ;
      RECT 91.915 4.385 92.945 4.545 ;
      RECT 91.895 4.385 92.945 4.515 ;
      RECT 91.875 3.295 92.045 4.485 ;
      RECT 91.845 4.385 92.945 4.455 ;
      RECT 91.815 4.385 92.945 4.425 ;
      RECT 91.785 4.375 92.145 4.395 ;
      RECT 91.785 4.365 92.135 4.395 ;
      RECT 91.155 4.195 92.045 4.365 ;
      RECT 91.155 4.355 92.115 4.365 ;
      RECT 91.155 4.345 92.105 4.365 ;
      RECT 91.155 3.295 92.045 3.465 ;
      RECT 92.215 3.795 92.545 4.215 ;
      RECT 92.215 3.305 92.435 4.215 ;
      RECT 92.135 7.165 92.345 7.765 ;
      RECT 91.995 7.165 92.345 7.365 ;
      RECT 90.715 4.765 90.985 5.465 ;
      RECT 90.815 3.265 90.985 5.465 ;
      RECT 90.725 3.265 90.985 3.735 ;
      RECT 88.855 4.425 89.105 4.965 ;
      RECT 89.825 4.425 90.545 4.895 ;
      RECT 88.855 4.425 90.645 4.595 ;
      RECT 90.415 3.995 90.645 4.595 ;
      RECT 89.415 3.305 89.665 4.595 ;
      RECT 88.875 3.305 89.665 3.575 ;
      RECT 89.835 7.115 90.515 7.365 ;
      RECT 90.245 6.755 90.515 7.365 ;
      RECT 89.995 7.535 90.255 8.085 ;
      RECT 89.995 7.535 90.325 8.06 ;
      RECT 88.935 7.535 90.325 7.725 ;
      RECT 88.935 6.695 89.105 7.725 ;
      RECT 88.815 7.115 89.105 7.445 ;
      RECT 88.935 6.695 89.875 6.865 ;
      RECT 89.575 6.145 89.875 6.865 ;
      RECT 89.835 3.725 90.245 4.245 ;
      RECT 89.835 3.305 90.035 4.245 ;
      RECT 88.445 3.485 88.615 5.465 ;
      RECT 88.445 3.995 89.245 4.245 ;
      RECT 88.445 3.485 88.695 4.245 ;
      RECT 88.365 3.485 88.695 3.905 ;
      RECT 88.395 7.895 88.955 8.185 ;
      RECT 88.395 5.975 88.645 8.185 ;
      RECT 88.395 5.975 88.855 6.525 ;
      RECT 86.605 10.035 86.78 10.585 ;
      RECT 86.605 7.295 86.775 10.585 ;
      RECT 86.605 7.295 86.78 8.435 ;
      RECT 86.175 7.295 86.345 9.505 ;
      RECT 86.175 7.295 86.35 8.555 ;
      RECT 85.22 10.095 85.395 10.585 ;
      RECT 85.22 7.295 85.39 10.585 ;
      RECT 85.22 9.595 85.63 9.925 ;
      RECT 85.22 8.755 85.63 9.085 ;
      RECT 85.22 7.295 85.395 8.555 ;
      RECT 83.6 7.3 83.77 8.77 ;
      RECT 83.6 7.3 83.775 8.56 ;
      RECT 83.23 3.04 83.4 4.23 ;
      RECT 83.23 3.04 83.7 3.21 ;
      RECT 83.23 9.25 83.7 9.42 ;
      RECT 83.23 8.23 83.4 9.42 ;
      RECT 82.61 3.9 82.785 5.16 ;
      RECT 82.61 3.69 82.78 5.16 ;
      RECT 82.61 7.3 82.78 8.77 ;
      RECT 82.61 7.3 82.785 8.56 ;
      RECT 82.24 3.04 82.41 4.23 ;
      RECT 82.24 3.04 82.71 3.21 ;
      RECT 82.24 9.25 82.71 9.42 ;
      RECT 82.24 8.23 82.41 9.42 ;
      RECT 81.25 4.02 81.425 5.16 ;
      RECT 81.25 1.87 81.42 5.16 ;
      RECT 81.25 1.87 81.425 2.42 ;
      RECT 81.25 10.04 81.425 10.59 ;
      RECT 81.25 7.3 81.42 10.59 ;
      RECT 81.25 7.3 81.425 8.44 ;
      RECT 80.82 3.9 80.995 5.16 ;
      RECT 80.82 2.95 80.99 5.16 ;
      RECT 80.82 7.3 80.99 9.51 ;
      RECT 80.82 7.3 80.995 8.56 ;
      RECT 80.39 3.93 80.56 5.16 ;
      RECT 80.45 2.15 80.62 4.1 ;
      RECT 80.39 1.87 80.56 2.32 ;
      RECT 80.39 10.14 80.56 10.59 ;
      RECT 80.45 8.36 80.62 10.31 ;
      RECT 80.39 7.3 80.56 8.53 ;
      RECT 79.865 3.9 80.04 5.16 ;
      RECT 79.865 1.87 80.035 5.16 ;
      RECT 79.865 3.37 80.275 3.7 ;
      RECT 79.865 2.53 80.275 2.86 ;
      RECT 79.865 1.87 80.04 2.36 ;
      RECT 79.865 10.1 80.04 10.59 ;
      RECT 79.865 7.3 80.035 10.59 ;
      RECT 79.865 9.6 80.275 9.93 ;
      RECT 79.865 8.76 80.275 9.09 ;
      RECT 79.865 7.3 80.04 8.56 ;
      RECT 75.125 7.935 76.435 8.185 ;
      RECT 75.125 7.615 75.305 8.185 ;
      RECT 74.575 7.615 75.305 7.785 ;
      RECT 74.575 6.775 74.745 7.785 ;
      RECT 75.415 6.815 77.155 6.995 ;
      RECT 76.825 5.975 77.155 6.995 ;
      RECT 74.575 6.775 75.635 6.945 ;
      RECT 76.825 6.145 77.645 6.315 ;
      RECT 75.985 5.975 76.315 6.185 ;
      RECT 75.985 5.975 77.155 6.145 ;
      RECT 76.885 4.495 77.215 5.455 ;
      RECT 76.885 4.495 77.565 4.665 ;
      RECT 77.395 3.265 77.565 4.665 ;
      RECT 77.305 3.265 77.635 3.895 ;
      RECT 76.435 4.765 76.705 5.465 ;
      RECT 76.535 3.265 76.705 5.465 ;
      RECT 76.875 4.075 77.225 4.325 ;
      RECT 76.535 4.105 77.225 4.275 ;
      RECT 76.445 3.265 76.705 3.735 ;
      RECT 75.775 6.405 76.655 6.645 ;
      RECT 76.425 6.315 76.655 6.645 ;
      RECT 75.125 6.405 76.655 6.605 ;
      RECT 76.045 6.355 76.655 6.645 ;
      RECT 75.125 6.275 75.295 6.605 ;
      RECT 76.015 7.165 76.265 7.765 ;
      RECT 76.015 7.165 76.485 7.365 ;
      RECT 75.505 4.385 76.265 4.885 ;
      RECT 74.575 4.195 74.835 4.815 ;
      RECT 75.495 4.325 75.505 4.635 ;
      RECT 75.475 4.385 76.265 4.605 ;
      RECT 76.135 3.995 76.365 4.595 ;
      RECT 75.455 4.315 75.495 4.575 ;
      RECT 75.435 4.385 76.365 4.565 ;
      RECT 75.405 4.385 76.365 4.555 ;
      RECT 75.335 4.385 76.365 4.545 ;
      RECT 75.315 4.385 76.365 4.515 ;
      RECT 75.295 3.295 75.465 4.485 ;
      RECT 75.265 4.385 76.365 4.455 ;
      RECT 75.235 4.385 76.365 4.425 ;
      RECT 75.205 4.375 75.565 4.395 ;
      RECT 75.205 4.365 75.555 4.395 ;
      RECT 74.575 4.195 75.465 4.365 ;
      RECT 74.575 4.355 75.535 4.365 ;
      RECT 74.575 4.345 75.525 4.365 ;
      RECT 74.575 3.295 75.465 3.465 ;
      RECT 75.635 3.795 75.965 4.215 ;
      RECT 75.635 3.305 75.855 4.215 ;
      RECT 75.555 7.165 75.765 7.765 ;
      RECT 75.415 7.165 75.765 7.365 ;
      RECT 74.135 4.765 74.405 5.465 ;
      RECT 74.235 3.265 74.405 5.465 ;
      RECT 74.145 3.265 74.405 3.735 ;
      RECT 72.275 4.425 72.525 4.965 ;
      RECT 73.245 4.425 73.965 4.895 ;
      RECT 72.275 4.425 74.065 4.595 ;
      RECT 73.835 3.995 74.065 4.595 ;
      RECT 72.835 3.305 73.085 4.595 ;
      RECT 72.295 3.305 73.085 3.575 ;
      RECT 73.255 7.115 73.935 7.365 ;
      RECT 73.665 6.755 73.935 7.365 ;
      RECT 73.415 7.535 73.675 8.085 ;
      RECT 73.415 7.535 73.745 8.06 ;
      RECT 72.355 7.535 73.745 7.725 ;
      RECT 72.355 6.695 72.525 7.725 ;
      RECT 72.235 7.115 72.525 7.445 ;
      RECT 72.355 6.695 73.295 6.865 ;
      RECT 72.995 6.145 73.295 6.865 ;
      RECT 73.255 3.725 73.665 4.245 ;
      RECT 73.255 3.305 73.455 4.245 ;
      RECT 71.865 3.485 72.035 5.465 ;
      RECT 71.865 3.995 72.665 4.245 ;
      RECT 71.865 3.485 72.115 4.245 ;
      RECT 71.785 3.485 72.115 3.905 ;
      RECT 71.815 7.895 72.375 8.185 ;
      RECT 71.815 5.975 72.065 8.185 ;
      RECT 71.815 5.975 72.275 6.525 ;
      RECT 70.025 10.035 70.2 10.585 ;
      RECT 70.025 7.295 70.195 10.585 ;
      RECT 70.025 7.295 70.2 8.435 ;
      RECT 69.595 7.295 69.765 9.505 ;
      RECT 69.595 7.295 69.77 8.555 ;
      RECT 68.64 10.095 68.815 10.585 ;
      RECT 68.64 7.295 68.81 10.585 ;
      RECT 68.64 9.595 69.05 9.925 ;
      RECT 68.64 8.755 69.05 9.085 ;
      RECT 68.64 7.295 68.815 8.555 ;
      RECT 67.015 7.3 67.185 8.77 ;
      RECT 67.015 7.3 67.19 8.56 ;
      RECT 66.645 3.04 66.815 4.23 ;
      RECT 66.645 3.04 67.115 3.21 ;
      RECT 66.645 9.25 67.115 9.42 ;
      RECT 66.645 8.23 66.815 9.42 ;
      RECT 66.025 3.9 66.2 5.16 ;
      RECT 66.025 3.69 66.195 5.16 ;
      RECT 66.025 7.3 66.195 8.77 ;
      RECT 66.025 7.3 66.2 8.56 ;
      RECT 65.655 3.04 65.825 4.23 ;
      RECT 65.655 3.04 66.125 3.21 ;
      RECT 65.655 9.25 66.125 9.42 ;
      RECT 65.655 8.23 65.825 9.42 ;
      RECT 64.665 4.02 64.84 5.16 ;
      RECT 64.665 1.87 64.835 5.16 ;
      RECT 64.665 1.87 64.84 2.42 ;
      RECT 64.665 10.04 64.84 10.59 ;
      RECT 64.665 7.3 64.835 10.59 ;
      RECT 64.665 7.3 64.84 8.44 ;
      RECT 64.235 3.9 64.41 5.16 ;
      RECT 64.235 2.95 64.405 5.16 ;
      RECT 64.235 7.3 64.405 9.51 ;
      RECT 64.235 7.3 64.41 8.56 ;
      RECT 63.805 3.93 63.975 5.16 ;
      RECT 63.865 2.15 64.035 4.1 ;
      RECT 63.805 1.87 63.975 2.32 ;
      RECT 63.805 10.14 63.975 10.59 ;
      RECT 63.865 8.36 64.035 10.31 ;
      RECT 63.805 7.3 63.975 8.53 ;
      RECT 63.28 3.9 63.455 5.16 ;
      RECT 63.28 1.87 63.45 5.16 ;
      RECT 63.28 3.37 63.69 3.7 ;
      RECT 63.28 2.53 63.69 2.86 ;
      RECT 63.28 1.87 63.455 2.36 ;
      RECT 63.28 10.1 63.455 10.59 ;
      RECT 63.28 7.3 63.45 10.59 ;
      RECT 63.28 9.6 63.69 9.93 ;
      RECT 63.28 8.76 63.69 9.09 ;
      RECT 63.28 7.3 63.455 8.56 ;
      RECT 58.54 7.935 59.85 8.185 ;
      RECT 58.54 7.615 58.72 8.185 ;
      RECT 57.99 7.615 58.72 7.785 ;
      RECT 57.99 6.775 58.16 7.785 ;
      RECT 58.83 6.815 60.57 6.995 ;
      RECT 60.24 5.975 60.57 6.995 ;
      RECT 57.99 6.775 59.05 6.945 ;
      RECT 60.24 6.145 61.06 6.315 ;
      RECT 59.4 5.975 59.73 6.185 ;
      RECT 59.4 5.975 60.57 6.145 ;
      RECT 60.3 4.495 60.63 5.455 ;
      RECT 60.3 4.495 60.98 4.665 ;
      RECT 60.81 3.265 60.98 4.665 ;
      RECT 60.72 3.265 61.05 3.895 ;
      RECT 59.85 4.765 60.12 5.465 ;
      RECT 59.95 3.265 60.12 5.465 ;
      RECT 60.29 4.075 60.64 4.325 ;
      RECT 59.95 4.105 60.64 4.275 ;
      RECT 59.86 3.265 60.12 3.735 ;
      RECT 59.19 6.405 60.07 6.645 ;
      RECT 59.84 6.315 60.07 6.645 ;
      RECT 58.54 6.405 60.07 6.605 ;
      RECT 59.46 6.355 60.07 6.645 ;
      RECT 58.54 6.275 58.71 6.605 ;
      RECT 59.43 7.165 59.68 7.765 ;
      RECT 59.43 7.165 59.9 7.365 ;
      RECT 58.92 4.385 59.68 4.885 ;
      RECT 57.99 4.195 58.25 4.815 ;
      RECT 58.91 4.325 58.92 4.635 ;
      RECT 58.89 4.385 59.68 4.605 ;
      RECT 59.55 3.995 59.78 4.595 ;
      RECT 58.87 4.315 58.91 4.575 ;
      RECT 58.85 4.385 59.78 4.565 ;
      RECT 58.82 4.385 59.78 4.555 ;
      RECT 58.75 4.385 59.78 4.545 ;
      RECT 58.73 4.385 59.78 4.515 ;
      RECT 58.71 3.295 58.88 4.485 ;
      RECT 58.68 4.385 59.78 4.455 ;
      RECT 58.65 4.385 59.78 4.425 ;
      RECT 58.62 4.375 58.98 4.395 ;
      RECT 58.62 4.365 58.97 4.395 ;
      RECT 57.99 4.195 58.88 4.365 ;
      RECT 57.99 4.355 58.95 4.365 ;
      RECT 57.99 4.345 58.94 4.365 ;
      RECT 57.99 3.295 58.88 3.465 ;
      RECT 59.05 3.795 59.38 4.215 ;
      RECT 59.05 3.305 59.27 4.215 ;
      RECT 58.97 7.165 59.18 7.765 ;
      RECT 58.83 7.165 59.18 7.365 ;
      RECT 57.55 4.765 57.82 5.465 ;
      RECT 57.65 3.265 57.82 5.465 ;
      RECT 57.56 3.265 57.82 3.735 ;
      RECT 55.69 4.425 55.94 4.965 ;
      RECT 56.66 4.425 57.38 4.895 ;
      RECT 55.69 4.425 57.48 4.595 ;
      RECT 57.25 3.995 57.48 4.595 ;
      RECT 56.25 3.305 56.5 4.595 ;
      RECT 55.71 3.305 56.5 3.575 ;
      RECT 56.67 7.115 57.35 7.365 ;
      RECT 57.08 6.755 57.35 7.365 ;
      RECT 56.83 7.535 57.09 8.085 ;
      RECT 56.83 7.535 57.16 8.06 ;
      RECT 55.77 7.535 57.16 7.725 ;
      RECT 55.77 6.695 55.94 7.725 ;
      RECT 55.65 7.115 55.94 7.445 ;
      RECT 55.77 6.695 56.71 6.865 ;
      RECT 56.41 6.145 56.71 6.865 ;
      RECT 56.67 3.725 57.08 4.245 ;
      RECT 56.67 3.305 56.87 4.245 ;
      RECT 55.28 3.485 55.45 5.465 ;
      RECT 55.28 3.995 56.08 4.245 ;
      RECT 55.28 3.485 55.53 4.245 ;
      RECT 55.2 3.485 55.53 3.905 ;
      RECT 55.23 7.895 55.79 8.185 ;
      RECT 55.23 5.975 55.48 8.185 ;
      RECT 55.23 5.975 55.69 6.525 ;
      RECT 53.44 10.035 53.615 10.585 ;
      RECT 53.44 7.295 53.61 10.585 ;
      RECT 53.44 7.295 53.615 8.435 ;
      RECT 53.01 7.295 53.18 9.505 ;
      RECT 53.01 7.295 53.185 8.555 ;
      RECT 52.055 10.095 52.23 10.585 ;
      RECT 52.055 7.295 52.225 10.585 ;
      RECT 52.055 9.595 52.465 9.925 ;
      RECT 52.055 8.755 52.465 9.085 ;
      RECT 52.055 7.295 52.23 8.555 ;
      RECT 50.43 7.3 50.6 8.77 ;
      RECT 50.43 7.3 50.605 8.56 ;
      RECT 50.06 3.04 50.23 4.23 ;
      RECT 50.06 3.04 50.53 3.21 ;
      RECT 50.06 9.25 50.53 9.42 ;
      RECT 50.06 8.23 50.23 9.42 ;
      RECT 49.44 3.9 49.615 5.16 ;
      RECT 49.44 3.69 49.61 5.16 ;
      RECT 49.44 7.3 49.61 8.77 ;
      RECT 49.44 7.3 49.615 8.56 ;
      RECT 49.07 3.04 49.24 4.23 ;
      RECT 49.07 3.04 49.54 3.21 ;
      RECT 49.07 9.25 49.54 9.42 ;
      RECT 49.07 8.23 49.24 9.42 ;
      RECT 48.08 4.02 48.255 5.16 ;
      RECT 48.08 1.87 48.25 5.16 ;
      RECT 48.08 1.87 48.255 2.42 ;
      RECT 48.08 10.04 48.255 10.59 ;
      RECT 48.08 7.3 48.25 10.59 ;
      RECT 48.08 7.3 48.255 8.44 ;
      RECT 47.65 3.9 47.825 5.16 ;
      RECT 47.65 2.95 47.82 5.16 ;
      RECT 47.65 7.3 47.82 9.51 ;
      RECT 47.65 7.3 47.825 8.56 ;
      RECT 47.22 3.93 47.39 5.16 ;
      RECT 47.28 2.15 47.45 4.1 ;
      RECT 47.22 1.87 47.39 2.32 ;
      RECT 47.22 10.14 47.39 10.59 ;
      RECT 47.28 8.36 47.45 10.31 ;
      RECT 47.22 7.3 47.39 8.53 ;
      RECT 46.695 3.9 46.87 5.16 ;
      RECT 46.695 1.87 46.865 5.16 ;
      RECT 46.695 3.37 47.105 3.7 ;
      RECT 46.695 2.53 47.105 2.86 ;
      RECT 46.695 1.87 46.87 2.36 ;
      RECT 46.695 10.1 46.87 10.59 ;
      RECT 46.695 7.3 46.865 10.59 ;
      RECT 46.695 9.6 47.105 9.93 ;
      RECT 46.695 8.76 47.105 9.09 ;
      RECT 46.695 7.3 46.87 8.56 ;
      RECT 41.955 7.935 43.265 8.185 ;
      RECT 41.955 7.615 42.135 8.185 ;
      RECT 41.405 7.615 42.135 7.785 ;
      RECT 41.405 6.775 41.575 7.785 ;
      RECT 42.245 6.815 43.985 6.995 ;
      RECT 43.655 5.975 43.985 6.995 ;
      RECT 41.405 6.775 42.465 6.945 ;
      RECT 43.655 6.145 44.475 6.315 ;
      RECT 42.815 5.975 43.145 6.185 ;
      RECT 42.815 5.975 43.985 6.145 ;
      RECT 43.715 4.495 44.045 5.455 ;
      RECT 43.715 4.495 44.395 4.665 ;
      RECT 44.225 3.265 44.395 4.665 ;
      RECT 44.135 3.265 44.465 3.895 ;
      RECT 43.265 4.765 43.535 5.465 ;
      RECT 43.365 3.265 43.535 5.465 ;
      RECT 43.705 4.075 44.055 4.325 ;
      RECT 43.365 4.105 44.055 4.275 ;
      RECT 43.275 3.265 43.535 3.735 ;
      RECT 42.605 6.405 43.485 6.645 ;
      RECT 43.255 6.315 43.485 6.645 ;
      RECT 41.955 6.405 43.485 6.605 ;
      RECT 42.875 6.355 43.485 6.645 ;
      RECT 41.955 6.275 42.125 6.605 ;
      RECT 42.845 7.165 43.095 7.765 ;
      RECT 42.845 7.165 43.315 7.365 ;
      RECT 42.335 4.385 43.095 4.885 ;
      RECT 41.405 4.195 41.665 4.815 ;
      RECT 42.325 4.325 42.335 4.635 ;
      RECT 42.305 4.385 43.095 4.605 ;
      RECT 42.965 3.995 43.195 4.595 ;
      RECT 42.285 4.315 42.325 4.575 ;
      RECT 42.265 4.385 43.195 4.565 ;
      RECT 42.235 4.385 43.195 4.555 ;
      RECT 42.165 4.385 43.195 4.545 ;
      RECT 42.145 4.385 43.195 4.515 ;
      RECT 42.125 3.295 42.295 4.485 ;
      RECT 42.095 4.385 43.195 4.455 ;
      RECT 42.065 4.385 43.195 4.425 ;
      RECT 42.035 4.375 42.395 4.395 ;
      RECT 42.035 4.365 42.385 4.395 ;
      RECT 41.405 4.195 42.295 4.365 ;
      RECT 41.405 4.355 42.365 4.365 ;
      RECT 41.405 4.345 42.355 4.365 ;
      RECT 41.405 3.295 42.295 3.465 ;
      RECT 42.465 3.795 42.795 4.215 ;
      RECT 42.465 3.305 42.685 4.215 ;
      RECT 42.385 7.165 42.595 7.765 ;
      RECT 42.245 7.165 42.595 7.365 ;
      RECT 40.965 4.765 41.235 5.465 ;
      RECT 41.065 3.265 41.235 5.465 ;
      RECT 40.975 3.265 41.235 3.735 ;
      RECT 39.105 4.425 39.355 4.965 ;
      RECT 40.075 4.425 40.795 4.895 ;
      RECT 39.105 4.425 40.895 4.595 ;
      RECT 40.665 3.995 40.895 4.595 ;
      RECT 39.665 3.305 39.915 4.595 ;
      RECT 39.125 3.305 39.915 3.575 ;
      RECT 40.085 7.115 40.765 7.365 ;
      RECT 40.495 6.755 40.765 7.365 ;
      RECT 40.245 7.535 40.505 8.085 ;
      RECT 40.245 7.535 40.575 8.06 ;
      RECT 39.185 7.535 40.575 7.725 ;
      RECT 39.185 6.695 39.355 7.725 ;
      RECT 39.065 7.115 39.355 7.445 ;
      RECT 39.185 6.695 40.125 6.865 ;
      RECT 39.825 6.145 40.125 6.865 ;
      RECT 40.085 3.725 40.495 4.245 ;
      RECT 40.085 3.305 40.285 4.245 ;
      RECT 38.695 3.485 38.865 5.465 ;
      RECT 38.695 3.995 39.495 4.245 ;
      RECT 38.695 3.485 38.945 4.245 ;
      RECT 38.615 3.485 38.945 3.905 ;
      RECT 38.645 7.895 39.205 8.185 ;
      RECT 38.645 5.975 38.895 8.185 ;
      RECT 38.645 5.975 39.105 6.525 ;
      RECT 36.855 10.035 37.03 10.585 ;
      RECT 36.855 7.295 37.025 10.585 ;
      RECT 36.855 7.295 37.03 8.435 ;
      RECT 36.425 7.295 36.595 9.505 ;
      RECT 36.425 7.295 36.6 8.555 ;
      RECT 35.47 10.095 35.645 10.585 ;
      RECT 35.47 7.295 35.64 10.585 ;
      RECT 35.47 9.595 35.88 9.925 ;
      RECT 35.47 8.755 35.88 9.085 ;
      RECT 35.47 7.295 35.645 8.555 ;
      RECT 33.845 7.3 34.015 8.77 ;
      RECT 33.845 7.3 34.02 8.56 ;
      RECT 33.475 3.04 33.645 4.23 ;
      RECT 33.475 3.04 33.945 3.21 ;
      RECT 33.475 9.25 33.945 9.42 ;
      RECT 33.475 8.23 33.645 9.42 ;
      RECT 32.855 3.9 33.03 5.16 ;
      RECT 32.855 3.69 33.025 5.16 ;
      RECT 32.855 7.3 33.025 8.77 ;
      RECT 32.855 7.3 33.03 8.56 ;
      RECT 32.485 3.04 32.655 4.23 ;
      RECT 32.485 3.04 32.955 3.21 ;
      RECT 32.485 9.25 32.955 9.42 ;
      RECT 32.485 8.23 32.655 9.42 ;
      RECT 31.495 4.02 31.67 5.16 ;
      RECT 31.495 1.87 31.665 5.16 ;
      RECT 31.495 1.87 31.67 2.42 ;
      RECT 31.495 10.04 31.67 10.59 ;
      RECT 31.495 7.3 31.665 10.59 ;
      RECT 31.495 7.3 31.67 8.44 ;
      RECT 31.065 3.9 31.24 5.16 ;
      RECT 31.065 2.95 31.235 5.16 ;
      RECT 31.065 7.3 31.235 9.51 ;
      RECT 31.065 7.3 31.24 8.56 ;
      RECT 30.635 3.93 30.805 5.16 ;
      RECT 30.695 2.15 30.865 4.1 ;
      RECT 30.635 1.87 30.805 2.32 ;
      RECT 30.635 10.14 30.805 10.59 ;
      RECT 30.695 8.36 30.865 10.31 ;
      RECT 30.635 7.3 30.805 8.53 ;
      RECT 30.11 3.9 30.285 5.16 ;
      RECT 30.11 1.87 30.28 5.16 ;
      RECT 30.11 3.37 30.52 3.7 ;
      RECT 30.11 2.53 30.52 2.86 ;
      RECT 30.11 1.87 30.285 2.36 ;
      RECT 30.11 10.1 30.285 10.59 ;
      RECT 30.11 7.3 30.28 10.59 ;
      RECT 30.11 9.6 30.52 9.93 ;
      RECT 30.11 8.76 30.52 9.09 ;
      RECT 30.11 7.3 30.285 8.56 ;
      RECT 25.37 7.935 26.68 8.185 ;
      RECT 25.37 7.615 25.55 8.185 ;
      RECT 24.82 7.615 25.55 7.785 ;
      RECT 24.82 6.775 24.99 7.785 ;
      RECT 25.66 6.815 27.4 6.995 ;
      RECT 27.07 5.975 27.4 6.995 ;
      RECT 24.82 6.775 25.88 6.945 ;
      RECT 27.07 6.145 27.89 6.315 ;
      RECT 26.23 5.975 26.56 6.185 ;
      RECT 26.23 5.975 27.4 6.145 ;
      RECT 27.13 4.495 27.46 5.455 ;
      RECT 27.13 4.495 27.81 4.665 ;
      RECT 27.64 3.265 27.81 4.665 ;
      RECT 27.55 3.265 27.88 3.895 ;
      RECT 26.68 4.765 26.95 5.465 ;
      RECT 26.78 3.265 26.95 5.465 ;
      RECT 27.12 4.075 27.47 4.325 ;
      RECT 26.78 4.105 27.47 4.275 ;
      RECT 26.69 3.265 26.95 3.735 ;
      RECT 26.02 6.405 26.9 6.645 ;
      RECT 26.67 6.315 26.9 6.645 ;
      RECT 25.37 6.405 26.9 6.605 ;
      RECT 26.29 6.355 26.9 6.645 ;
      RECT 25.37 6.275 25.54 6.605 ;
      RECT 26.26 7.165 26.51 7.765 ;
      RECT 26.26 7.165 26.73 7.365 ;
      RECT 25.75 4.385 26.51 4.885 ;
      RECT 24.82 4.195 25.08 4.815 ;
      RECT 25.74 4.325 25.75 4.635 ;
      RECT 25.72 4.385 26.51 4.605 ;
      RECT 26.38 3.995 26.61 4.595 ;
      RECT 25.7 4.315 25.74 4.575 ;
      RECT 25.68 4.385 26.61 4.565 ;
      RECT 25.65 4.385 26.61 4.555 ;
      RECT 25.58 4.385 26.61 4.545 ;
      RECT 25.56 4.385 26.61 4.515 ;
      RECT 25.54 3.295 25.71 4.485 ;
      RECT 25.51 4.385 26.61 4.455 ;
      RECT 25.48 4.385 26.61 4.425 ;
      RECT 25.45 4.375 25.81 4.395 ;
      RECT 25.45 4.365 25.8 4.395 ;
      RECT 24.82 4.195 25.71 4.365 ;
      RECT 24.82 4.355 25.78 4.365 ;
      RECT 24.82 4.345 25.77 4.365 ;
      RECT 24.82 3.295 25.71 3.465 ;
      RECT 25.88 3.795 26.21 4.215 ;
      RECT 25.88 3.305 26.1 4.215 ;
      RECT 25.8 7.165 26.01 7.765 ;
      RECT 25.66 7.165 26.01 7.365 ;
      RECT 24.38 4.765 24.65 5.465 ;
      RECT 24.48 3.265 24.65 5.465 ;
      RECT 24.39 3.265 24.65 3.735 ;
      RECT 22.52 4.425 22.77 4.965 ;
      RECT 23.49 4.425 24.21 4.895 ;
      RECT 22.52 4.425 24.31 4.595 ;
      RECT 24.08 3.995 24.31 4.595 ;
      RECT 23.08 3.305 23.33 4.595 ;
      RECT 22.54 3.305 23.33 3.575 ;
      RECT 23.5 7.115 24.18 7.365 ;
      RECT 23.91 6.755 24.18 7.365 ;
      RECT 23.66 7.535 23.92 8.085 ;
      RECT 23.66 7.535 23.99 8.06 ;
      RECT 22.6 7.535 23.99 7.725 ;
      RECT 22.6 6.695 22.77 7.725 ;
      RECT 22.48 7.115 22.77 7.445 ;
      RECT 22.6 6.695 23.54 6.865 ;
      RECT 23.24 6.145 23.54 6.865 ;
      RECT 23.5 3.725 23.91 4.245 ;
      RECT 23.5 3.305 23.7 4.245 ;
      RECT 22.11 3.485 22.28 5.465 ;
      RECT 22.11 3.995 22.91 4.245 ;
      RECT 22.11 3.485 22.36 4.245 ;
      RECT 22.03 3.485 22.36 3.905 ;
      RECT 22.06 7.895 22.62 8.185 ;
      RECT 22.06 5.975 22.31 8.185 ;
      RECT 22.06 5.975 22.52 6.525 ;
      RECT 20.27 10.035 20.445 10.585 ;
      RECT 20.27 7.295 20.44 10.585 ;
      RECT 20.27 7.295 20.445 8.435 ;
      RECT 19.84 7.295 20.01 9.505 ;
      RECT 19.84 7.295 20.015 8.555 ;
      RECT 18.885 10.095 19.06 10.585 ;
      RECT 18.885 7.295 19.055 10.585 ;
      RECT 18.885 9.595 19.295 9.925 ;
      RECT 18.885 8.755 19.295 9.085 ;
      RECT 18.885 7.295 19.06 8.555 ;
      RECT 16.61 7.295 16.78 9.505 ;
      RECT 16.61 7.295 16.785 8.555 ;
      RECT 16.18 10.135 16.35 10.585 ;
      RECT 16.24 8.355 16.41 10.305 ;
      RECT 16.18 7.295 16.35 8.525 ;
      RECT 15.655 10.095 15.83 10.585 ;
      RECT 15.655 7.295 15.825 10.585 ;
      RECT 15.655 9.595 16.065 9.925 ;
      RECT 15.655 8.755 16.065 9.085 ;
      RECT 15.655 7.295 15.83 8.555 ;
      RECT 100.18 10.08 100.355 10.59 ;
      RECT 99.19 1.87 99.365 2.38 ;
      RECT 99.19 10.08 99.365 10.59 ;
      RECT 97.4 1.87 97.575 2.38 ;
      RECT 97.4 10.08 97.575 10.59 ;
      RECT 94.315 4.075 94.665 4.325 ;
      RECT 93.255 7.165 93.705 7.675 ;
      RECT 91.935 5.125 92.415 5.465 ;
      RECT 91.155 3.635 91.705 4.025 ;
      RECT 89.645 5.125 90.115 5.465 ;
      RECT 87.935 4.075 88.275 4.955 ;
      RECT 86.175 10.075 86.35 10.585 ;
      RECT 83.6 10.08 83.775 10.59 ;
      RECT 82.61 1.87 82.785 2.38 ;
      RECT 82.61 10.08 82.785 10.59 ;
      RECT 80.82 1.87 80.995 2.38 ;
      RECT 80.82 10.08 80.995 10.59 ;
      RECT 77.735 4.075 78.085 4.325 ;
      RECT 76.675 7.165 77.125 7.675 ;
      RECT 75.355 5.125 75.835 5.465 ;
      RECT 74.575 3.635 75.125 4.025 ;
      RECT 73.065 5.125 73.535 5.465 ;
      RECT 71.355 4.075 71.695 4.955 ;
      RECT 69.595 10.075 69.77 10.585 ;
      RECT 67.015 10.08 67.19 10.59 ;
      RECT 66.025 1.87 66.2 2.38 ;
      RECT 66.025 10.08 66.2 10.59 ;
      RECT 64.235 1.87 64.41 2.38 ;
      RECT 64.235 10.08 64.41 10.59 ;
      RECT 61.15 4.075 61.5 4.325 ;
      RECT 60.09 7.165 60.54 7.675 ;
      RECT 58.77 5.125 59.25 5.465 ;
      RECT 57.99 3.635 58.54 4.025 ;
      RECT 56.48 5.125 56.95 5.465 ;
      RECT 54.77 4.075 55.11 4.955 ;
      RECT 53.01 10.075 53.185 10.585 ;
      RECT 50.43 10.08 50.605 10.59 ;
      RECT 49.44 1.87 49.615 2.38 ;
      RECT 49.44 10.08 49.615 10.59 ;
      RECT 47.65 1.87 47.825 2.38 ;
      RECT 47.65 10.08 47.825 10.59 ;
      RECT 44.565 4.075 44.915 4.325 ;
      RECT 43.505 7.165 43.955 7.675 ;
      RECT 42.185 5.125 42.665 5.465 ;
      RECT 41.405 3.635 41.955 4.025 ;
      RECT 39.895 5.125 40.365 5.465 ;
      RECT 38.185 4.075 38.525 4.955 ;
      RECT 36.425 10.075 36.6 10.585 ;
      RECT 33.845 10.08 34.02 10.59 ;
      RECT 32.855 1.87 33.03 2.38 ;
      RECT 32.855 10.08 33.03 10.59 ;
      RECT 31.065 1.87 31.24 2.38 ;
      RECT 31.065 10.08 31.24 10.59 ;
      RECT 27.98 4.075 28.33 4.325 ;
      RECT 26.92 7.165 27.37 7.675 ;
      RECT 25.6 5.125 26.08 5.465 ;
      RECT 24.82 3.635 25.37 4.025 ;
      RECT 23.31 5.125 23.78 5.465 ;
      RECT 21.6 4.075 21.94 4.955 ;
      RECT 19.84 10.075 20.015 10.585 ;
      RECT 16.61 10.075 16.785 10.585 ;
  END
END sky130_osu_ring_oscillator_mpr2ca_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2ca_8_b0r2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ca_8_b0r2 ;
  SIZE 101.085 BY 12.47 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 34.105 0 34.485 5.27 ;
      LAYER met2 ;
        RECT 34.105 4.89 34.485 5.27 ;
      LAYER li1 ;
        RECT 34.205 1.87 34.38 2.38 ;
        RECT 34.205 3.9 34.38 5.16 ;
        RECT 34.205 3.69 34.375 5.16 ;
      LAYER met1 ;
        RECT 34.12 4.935 34.47 5.225 ;
        RECT 34.145 2.18 34.44 2.41 ;
        RECT 34.145 3.66 34.435 3.89 ;
        RECT 34.205 2.18 34.375 3.89 ;
      LAYER via1 ;
        RECT 34.22 5.005 34.37 5.155 ;
      LAYER via2 ;
        RECT 34.195 4.98 34.395 5.18 ;
      LAYER mcon ;
        RECT 34.205 3.69 34.375 3.86 ;
        RECT 34.205 2.21 34.375 2.38 ;
        RECT 34.21 4.99 34.38 5.16 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 50.69 0 51.07 5.27 ;
      LAYER met2 ;
        RECT 50.69 4.89 51.07 5.27 ;
      LAYER li1 ;
        RECT 50.79 1.87 50.965 2.38 ;
        RECT 50.79 3.9 50.965 5.16 ;
        RECT 50.79 3.69 50.96 5.16 ;
      LAYER met1 ;
        RECT 50.705 4.935 51.055 5.225 ;
        RECT 50.73 2.18 51.025 2.41 ;
        RECT 50.73 3.66 51.02 3.89 ;
        RECT 50.79 2.18 50.96 3.89 ;
      LAYER via1 ;
        RECT 50.805 5.005 50.955 5.155 ;
      LAYER via2 ;
        RECT 50.78 4.98 50.98 5.18 ;
      LAYER mcon ;
        RECT 50.79 3.69 50.96 3.86 ;
        RECT 50.79 2.21 50.96 2.38 ;
        RECT 50.795 4.99 50.965 5.16 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 67.275 0.005 67.655 5.275 ;
      LAYER met2 ;
        RECT 67.275 4.895 67.655 5.275 ;
      LAYER li1 ;
        RECT 67.375 1.875 67.55 2.385 ;
        RECT 67.375 3.905 67.55 5.165 ;
        RECT 67.375 3.695 67.545 5.165 ;
      LAYER met1 ;
        RECT 67.29 4.94 67.64 5.23 ;
        RECT 67.315 2.185 67.61 2.415 ;
        RECT 67.315 3.665 67.605 3.895 ;
        RECT 67.375 2.185 67.545 3.895 ;
      LAYER via1 ;
        RECT 67.39 5.01 67.54 5.16 ;
      LAYER via2 ;
        RECT 67.365 4.985 67.565 5.185 ;
      LAYER mcon ;
        RECT 67.375 3.695 67.545 3.865 ;
        RECT 67.375 2.215 67.545 2.385 ;
        RECT 67.38 4.995 67.55 5.165 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 83.86 0.01 84.24 5.28 ;
      LAYER met2 ;
        RECT 83.86 4.9 84.24 5.28 ;
      LAYER li1 ;
        RECT 83.96 1.88 84.135 2.39 ;
        RECT 83.96 3.91 84.135 5.17 ;
        RECT 83.96 3.7 84.13 5.17 ;
      LAYER met1 ;
        RECT 83.875 4.945 84.225 5.235 ;
        RECT 83.9 2.19 84.195 2.42 ;
        RECT 83.9 3.67 84.19 3.9 ;
        RECT 83.96 2.19 84.13 3.9 ;
      LAYER via1 ;
        RECT 83.975 5.015 84.125 5.165 ;
      LAYER via2 ;
        RECT 83.95 4.99 84.15 5.19 ;
      LAYER mcon ;
        RECT 83.96 3.7 84.13 3.87 ;
        RECT 83.96 2.22 84.13 2.39 ;
        RECT 83.965 5 84.135 5.17 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 100.44 0.01 100.82 5.28 ;
      LAYER met2 ;
        RECT 100.44 4.9 100.82 5.28 ;
      LAYER li1 ;
        RECT 100.54 1.88 100.715 2.39 ;
        RECT 100.54 3.91 100.715 5.17 ;
        RECT 100.54 3.7 100.71 5.17 ;
      LAYER met1 ;
        RECT 100.455 4.945 100.805 5.235 ;
        RECT 100.48 2.19 100.775 2.42 ;
        RECT 100.48 3.67 100.77 3.9 ;
        RECT 100.54 2.19 100.71 3.9 ;
      LAYER via1 ;
        RECT 100.555 5.015 100.705 5.165 ;
      LAYER via2 ;
        RECT 100.53 4.99 100.73 5.19 ;
      LAYER mcon ;
        RECT 100.54 3.7 100.71 3.87 ;
        RECT 100.54 2.22 100.71 2.39 ;
        RECT 100.545 5 100.715 5.17 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 29.98 8.15 30.305 8.475 ;
        RECT 29.975 4.93 30.3 5.255 ;
        RECT 21.135 9.3 30.22 9.47 ;
        RECT 30.045 4.93 30.22 9.47 ;
        RECT 21.08 8.145 21.36 8.485 ;
        RECT 21.135 8.145 21.305 9.47 ;
      LAYER li1 ;
        RECT 30.05 2.96 30.22 4.23 ;
        RECT 30.05 8.23 30.22 9.5 ;
        RECT 18.825 8.225 18.995 9.495 ;
      LAYER met1 ;
        RECT 29.99 4.06 30.45 4.23 ;
        RECT 29.975 4.93 30.3 5.255 ;
        RECT 29.99 4.03 30.28 4.26 ;
        RECT 30.05 4.03 30.23 5.255 ;
        RECT 29.98 8.23 30.45 8.4 ;
        RECT 29.98 8.15 30.305 8.475 ;
        RECT 21.05 8.175 21.39 8.455 ;
        RECT 18.765 8.23 21.39 8.4 ;
        RECT 18.765 8.225 19.225 8.4 ;
        RECT 18.765 8.195 19.055 8.425 ;
      LAYER via1 ;
        RECT 21.145 8.24 21.295 8.39 ;
        RECT 30.065 5.015 30.215 5.165 ;
        RECT 30.07 8.235 30.22 8.385 ;
      LAYER mcon ;
        RECT 18.825 8.225 18.995 8.395 ;
        RECT 30.05 8.23 30.22 8.4 ;
        RECT 30.05 4.06 30.22 4.23 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 46.565 8.15 46.89 8.475 ;
        RECT 46.56 4.93 46.885 5.255 ;
        RECT 37.72 9.3 46.805 9.47 ;
        RECT 46.63 4.93 46.805 9.47 ;
        RECT 37.665 8.145 37.945 8.485 ;
        RECT 37.72 8.145 37.89 9.47 ;
      LAYER li1 ;
        RECT 46.635 2.96 46.805 4.23 ;
        RECT 46.635 8.23 46.805 9.5 ;
        RECT 35.41 8.225 35.58 9.495 ;
      LAYER met1 ;
        RECT 46.575 4.06 47.035 4.23 ;
        RECT 46.56 4.93 46.885 5.255 ;
        RECT 46.575 4.03 46.865 4.26 ;
        RECT 46.635 4.03 46.815 5.255 ;
        RECT 46.565 8.23 47.035 8.4 ;
        RECT 46.565 8.15 46.89 8.475 ;
        RECT 37.635 8.175 37.975 8.455 ;
        RECT 35.35 8.23 37.975 8.4 ;
        RECT 35.35 8.225 35.81 8.4 ;
        RECT 35.35 8.195 35.64 8.425 ;
      LAYER via1 ;
        RECT 37.73 8.24 37.88 8.39 ;
        RECT 46.65 5.015 46.8 5.165 ;
        RECT 46.655 8.235 46.805 8.385 ;
      LAYER mcon ;
        RECT 35.41 8.225 35.58 8.395 ;
        RECT 46.635 8.23 46.805 8.4 ;
        RECT 46.635 4.06 46.805 4.23 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 63.15 8.155 63.475 8.48 ;
        RECT 63.145 4.935 63.47 5.26 ;
        RECT 54.305 9.305 63.39 9.475 ;
        RECT 63.215 4.935 63.39 9.475 ;
        RECT 54.25 8.15 54.53 8.49 ;
        RECT 54.305 8.15 54.475 9.475 ;
      LAYER li1 ;
        RECT 63.22 2.965 63.39 4.235 ;
        RECT 63.22 8.235 63.39 9.505 ;
        RECT 51.995 8.23 52.165 9.5 ;
      LAYER met1 ;
        RECT 63.16 4.065 63.62 4.235 ;
        RECT 63.145 4.935 63.47 5.26 ;
        RECT 63.16 4.035 63.45 4.265 ;
        RECT 63.22 4.035 63.4 5.26 ;
        RECT 63.15 8.235 63.62 8.405 ;
        RECT 63.15 8.155 63.475 8.48 ;
        RECT 54.22 8.18 54.56 8.46 ;
        RECT 51.935 8.235 54.56 8.405 ;
        RECT 51.935 8.23 52.395 8.405 ;
        RECT 51.935 8.2 52.225 8.43 ;
      LAYER via1 ;
        RECT 54.315 8.245 54.465 8.395 ;
        RECT 63.235 5.02 63.385 5.17 ;
        RECT 63.24 8.24 63.39 8.39 ;
      LAYER mcon ;
        RECT 51.995 8.23 52.165 8.4 ;
        RECT 63.22 8.235 63.39 8.405 ;
        RECT 63.22 4.065 63.39 4.235 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 79.735 8.16 80.06 8.485 ;
        RECT 79.73 4.94 80.055 5.265 ;
        RECT 70.89 9.31 79.975 9.48 ;
        RECT 79.8 4.94 79.975 9.48 ;
        RECT 70.835 8.155 71.115 8.495 ;
        RECT 70.89 8.155 71.06 9.48 ;
      LAYER li1 ;
        RECT 79.805 2.97 79.975 4.24 ;
        RECT 79.805 8.24 79.975 9.51 ;
        RECT 68.58 8.235 68.75 9.505 ;
      LAYER met1 ;
        RECT 79.745 4.07 80.205 4.24 ;
        RECT 79.73 4.94 80.055 5.265 ;
        RECT 79.745 4.04 80.035 4.27 ;
        RECT 79.805 4.04 79.985 5.265 ;
        RECT 79.735 8.24 80.205 8.41 ;
        RECT 79.735 8.16 80.06 8.485 ;
        RECT 70.805 8.185 71.145 8.465 ;
        RECT 68.52 8.24 71.145 8.41 ;
        RECT 68.52 8.235 68.98 8.41 ;
        RECT 68.52 8.205 68.81 8.435 ;
      LAYER via1 ;
        RECT 70.9 8.25 71.05 8.4 ;
        RECT 79.82 5.025 79.97 5.175 ;
        RECT 79.825 8.245 79.975 8.395 ;
      LAYER mcon ;
        RECT 68.58 8.235 68.75 8.405 ;
        RECT 79.805 8.24 79.975 8.41 ;
        RECT 79.805 4.07 79.975 4.24 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 96.315 8.16 96.64 8.485 ;
        RECT 96.31 4.94 96.635 5.265 ;
        RECT 87.47 9.31 96.555 9.48 ;
        RECT 96.38 4.94 96.555 9.48 ;
        RECT 87.415 8.155 87.695 8.495 ;
        RECT 87.47 8.155 87.64 9.48 ;
      LAYER li1 ;
        RECT 96.385 2.97 96.555 4.24 ;
        RECT 96.385 8.24 96.555 9.51 ;
        RECT 85.16 8.235 85.33 9.505 ;
      LAYER met1 ;
        RECT 96.325 4.07 96.785 4.24 ;
        RECT 96.31 4.94 96.635 5.265 ;
        RECT 96.325 4.04 96.615 4.27 ;
        RECT 96.385 4.04 96.565 5.265 ;
        RECT 96.315 8.24 96.785 8.41 ;
        RECT 96.315 8.16 96.64 8.485 ;
        RECT 87.385 8.185 87.725 8.465 ;
        RECT 85.1 8.24 87.725 8.41 ;
        RECT 85.1 8.235 85.56 8.41 ;
        RECT 85.1 8.205 85.39 8.435 ;
      LAYER via1 ;
        RECT 87.48 8.25 87.63 8.4 ;
        RECT 96.4 5.025 96.55 5.175 ;
        RECT 96.405 8.245 96.555 8.395 ;
      LAYER mcon ;
        RECT 85.16 8.235 85.33 8.405 ;
        RECT 96.385 8.24 96.555 8.41 ;
        RECT 96.385 4.07 96.555 4.24 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 15.595 8.225 15.765 9.495 ;
      LAYER met1 ;
        RECT 15.535 8.225 15.995 8.395 ;
        RECT 15.54 8.2 15.83 8.43 ;
        RECT 15.535 8.195 15.825 8.425 ;
      LAYER mcon ;
        RECT 15.595 8.225 15.765 8.395 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 95.145 5.43 101.085 7.05 ;
        RECT 100.11 4.71 100.28 7.77 ;
        RECT 99.12 4.71 99.29 7.77 ;
        RECT 96.375 4.71 96.545 7.77 ;
        RECT 95.015 5.43 101.085 5.975 ;
        RECT 94.685 4.505 95.015 5.815 ;
        RECT 61.85 5.645 101.085 5.815 ;
        RECT 92.945 5.105 93.205 5.815 ;
        RECT 92.385 5.645 92.755 6.195 ;
        RECT 91.945 4.725 92.275 4.965 ;
        RECT 91.945 4.725 92.135 4.995 ;
        RECT 91.515 4.995 92.125 5.815 ;
        RECT 91.565 4.995 91.835 6.595 ;
        RECT 90.645 5.105 90.865 5.815 ;
        RECT 90.405 5.645 90.685 6.485 ;
        RECT 89.635 4.775 89.965 4.965 ;
        RECT 89.215 5.145 89.835 5.815 ;
        RECT 89.635 4.775 89.835 5.815 ;
        RECT 89.405 5.145 89.735 6.535 ;
        RECT 88.295 5.135 88.555 5.815 ;
        RECT 78.565 5.43 88.33 7.03 ;
        RECT 78.565 5.43 88.075 7.035 ;
        RECT 85.15 5.43 85.32 7.765 ;
        RECT 78.565 5.43 84.505 7.05 ;
        RECT 83.53 4.71 83.7 7.77 ;
        RECT 82.54 4.71 82.71 7.77 ;
        RECT 79.795 4.71 79.965 7.77 ;
        RECT 78.435 5.43 88.33 5.975 ;
        RECT 78.105 4.505 78.435 5.815 ;
        RECT 76.365 5.105 76.625 5.815 ;
        RECT 75.805 5.645 76.175 6.195 ;
        RECT 75.365 4.725 75.695 4.965 ;
        RECT 75.365 4.725 75.555 4.995 ;
        RECT 74.935 4.995 75.545 5.815 ;
        RECT 74.985 4.995 75.255 6.595 ;
        RECT 74.065 5.105 74.285 5.815 ;
        RECT 73.825 5.645 74.105 6.485 ;
        RECT 73.055 4.775 73.385 4.965 ;
        RECT 72.635 5.145 73.255 5.815 ;
        RECT 73.055 4.775 73.255 5.815 ;
        RECT 72.825 5.145 73.155 6.535 ;
        RECT 0 5.64 71.975 5.805 ;
        RECT 71.715 5.135 71.975 5.815 ;
        RECT 61.98 5.43 71.745 7.03 ;
        RECT 61.98 5.43 71.495 7.035 ;
        RECT 68.57 5.43 68.74 7.765 ;
        RECT 61.98 5.43 67.92 7.045 ;
        RECT 66.945 4.705 67.115 7.765 ;
        RECT 65.955 4.705 66.125 7.765 ;
        RECT 63.21 4.705 63.38 7.765 ;
        RECT 61.85 5.43 71.745 5.97 ;
        RECT 61.52 4.5 61.85 5.81 ;
        RECT 45.265 5.645 101.085 5.81 ;
        RECT 59.78 5.1 60.04 5.81 ;
        RECT 59.22 5.64 59.59 6.19 ;
        RECT 58.78 4.72 59.11 4.96 ;
        RECT 58.78 4.72 58.97 4.99 ;
        RECT 58.35 4.99 58.96 5.81 ;
        RECT 58.4 4.99 58.67 6.59 ;
        RECT 57.48 5.1 57.7 5.81 ;
        RECT 57.24 5.64 57.52 6.48 ;
        RECT 56.47 4.77 56.8 4.96 ;
        RECT 56.05 5.14 56.67 5.81 ;
        RECT 56.47 4.77 56.67 5.81 ;
        RECT 56.24 5.14 56.57 6.53 ;
        RECT 0 5.635 55.39 5.805 ;
        RECT 55.13 5.13 55.39 5.81 ;
        RECT 45.395 5.43 55.16 7.03 ;
        RECT 51.985 5.43 52.155 7.76 ;
        RECT 45.395 5.43 51.335 7.04 ;
        RECT 50.36 4.7 50.53 7.76 ;
        RECT 49.37 4.7 49.54 7.76 ;
        RECT 46.625 4.7 46.795 7.76 ;
        RECT 45.265 5.43 55.16 5.965 ;
        RECT 44.935 4.495 45.265 5.805 ;
        RECT 43.195 5.095 43.455 5.805 ;
        RECT 42.635 5.635 43.005 6.185 ;
        RECT 42.195 4.715 42.525 4.955 ;
        RECT 42.195 4.715 42.385 4.985 ;
        RECT 41.765 4.985 42.375 5.805 ;
        RECT 41.815 4.985 42.085 6.585 ;
        RECT 40.895 5.095 41.115 5.805 ;
        RECT 40.655 5.635 40.935 6.475 ;
        RECT 39.885 4.765 40.215 4.955 ;
        RECT 39.465 5.135 40.085 5.805 ;
        RECT 39.885 4.765 40.085 5.805 ;
        RECT 39.655 5.135 39.985 6.525 ;
        RECT 38.545 5.125 38.805 5.805 ;
        RECT 28.81 5.43 38.575 7.03 ;
        RECT 34.75 5.425 38.325 7.03 ;
        RECT 35.4 5.425 35.57 7.755 ;
        RECT 28.81 5.43 34.75 7.04 ;
        RECT 33.775 4.7 33.945 7.76 ;
        RECT 32.785 4.7 32.955 7.76 ;
        RECT 30.04 4.7 30.21 7.76 ;
        RECT 28.68 5.43 38.575 5.965 ;
        RECT 28.35 4.495 28.68 5.805 ;
        RECT 26.61 5.095 26.87 5.805 ;
        RECT 26.05 5.635 26.42 6.185 ;
        RECT 25.61 4.715 25.94 4.955 ;
        RECT 25.61 4.715 25.8 4.985 ;
        RECT 25.18 4.985 25.79 5.805 ;
        RECT 25.23 4.985 25.5 6.585 ;
        RECT 24.31 5.095 24.53 5.805 ;
        RECT 24.07 5.635 24.35 6.475 ;
        RECT 23.3 4.765 23.63 4.955 ;
        RECT 22.88 5.135 23.5 5.805 ;
        RECT 23.3 4.765 23.5 5.805 ;
        RECT 23.07 5.135 23.4 6.525 ;
        RECT 21.96 5.125 22.22 5.805 ;
        RECT 0 5.425 21.965 7.025 ;
        RECT 18.815 5.425 18.985 7.755 ;
        RECT 17.4 10.035 17.575 10.585 ;
        RECT 17.4 7.295 17.575 8.435 ;
        RECT 17.4 5.425 17.57 10.585 ;
        RECT 15.585 5.425 15.755 7.755 ;
      LAYER met1 ;
        RECT 95.145 5.43 101.085 7.05 ;
        RECT 61.98 5.495 101.085 5.975 ;
        RECT 95.02 5.44 101.085 5.975 ;
        RECT 95.015 5.455 101.085 5.975 ;
        RECT 78.565 5.43 88.33 7.03 ;
        RECT 78.565 5.43 88.075 7.035 ;
        RECT 78.565 5.43 84.505 7.05 ;
        RECT 78.435 5.455 88.33 5.975 ;
        RECT 78.44 5.44 88.33 5.975 ;
        RECT 61.98 5.43 71.745 7.03 ;
        RECT 61.98 5.43 71.495 7.035 ;
        RECT 61.98 5.43 67.92 7.045 ;
        RECT 45.395 5.495 101.085 5.97 ;
        RECT 61.855 5.435 71.745 5.97 ;
        RECT 0 5.49 71.745 5.965 ;
        RECT 61.85 5.45 71.745 5.97 ;
        RECT 45.395 5.43 55.16 7.03 ;
        RECT 45.395 5.43 51.335 7.04 ;
        RECT 0 5.485 55.16 5.965 ;
        RECT 45.27 5.43 55.16 5.965 ;
        RECT 45.265 5.445 55.16 5.965 ;
        RECT 28.81 5.43 38.575 7.03 ;
        RECT 34.75 5.425 38.325 7.03 ;
        RECT 28.81 5.43 34.75 7.04 ;
        RECT 28.68 5.445 38.575 5.965 ;
        RECT 28.685 5.43 38.575 5.965 ;
        RECT 0 5.425 21.965 7.025 ;
        RECT 17.34 8.935 17.63 9.165 ;
        RECT 17.17 8.965 17.63 9.135 ;
      LAYER mcon ;
        RECT 17.4 8.965 17.57 9.135 ;
        RECT 17.705 6.825 17.875 6.995 ;
        RECT 20.935 6.825 21.105 6.995 ;
        RECT 22.02 5.635 22.19 5.805 ;
        RECT 22.48 5.635 22.65 5.805 ;
        RECT 22.94 5.635 23.11 5.805 ;
        RECT 23.4 5.635 23.57 5.805 ;
        RECT 23.86 5.635 24.03 5.805 ;
        RECT 24.32 5.635 24.49 5.805 ;
        RECT 24.78 5.635 24.95 5.805 ;
        RECT 25.24 5.635 25.41 5.805 ;
        RECT 25.7 5.635 25.87 5.805 ;
        RECT 26.16 5.635 26.33 5.805 ;
        RECT 26.62 5.635 26.79 5.805 ;
        RECT 27.08 5.635 27.25 5.805 ;
        RECT 27.54 5.635 27.71 5.805 ;
        RECT 28 5.635 28.17 5.805 ;
        RECT 28.46 5.635 28.63 5.805 ;
        RECT 32.16 6.83 32.33 7 ;
        RECT 32.16 5.46 32.33 5.63 ;
        RECT 32.865 6.83 33.035 7 ;
        RECT 32.865 5.46 33.035 5.63 ;
        RECT 33.855 6.83 34.025 7 ;
        RECT 33.855 5.46 34.025 5.63 ;
        RECT 37.52 6.825 37.69 6.995 ;
        RECT 38.605 5.635 38.775 5.805 ;
        RECT 39.065 5.635 39.235 5.805 ;
        RECT 39.525 5.635 39.695 5.805 ;
        RECT 39.985 5.635 40.155 5.805 ;
        RECT 40.445 5.635 40.615 5.805 ;
        RECT 40.905 5.635 41.075 5.805 ;
        RECT 41.365 5.635 41.535 5.805 ;
        RECT 41.825 5.635 41.995 5.805 ;
        RECT 42.285 5.635 42.455 5.805 ;
        RECT 42.745 5.635 42.915 5.805 ;
        RECT 43.205 5.635 43.375 5.805 ;
        RECT 43.665 5.635 43.835 5.805 ;
        RECT 44.125 5.635 44.295 5.805 ;
        RECT 44.585 5.635 44.755 5.805 ;
        RECT 45.045 5.635 45.215 5.805 ;
        RECT 48.745 6.83 48.915 7 ;
        RECT 48.745 5.46 48.915 5.63 ;
        RECT 49.45 6.83 49.62 7 ;
        RECT 49.45 5.46 49.62 5.63 ;
        RECT 50.44 6.83 50.61 7 ;
        RECT 50.44 5.46 50.61 5.63 ;
        RECT 54.105 6.83 54.275 7 ;
        RECT 55.19 5.64 55.36 5.81 ;
        RECT 55.65 5.64 55.82 5.81 ;
        RECT 56.11 5.64 56.28 5.81 ;
        RECT 56.57 5.64 56.74 5.81 ;
        RECT 57.03 5.64 57.2 5.81 ;
        RECT 57.49 5.64 57.66 5.81 ;
        RECT 57.95 5.64 58.12 5.81 ;
        RECT 58.41 5.64 58.58 5.81 ;
        RECT 58.87 5.64 59.04 5.81 ;
        RECT 59.33 5.64 59.5 5.81 ;
        RECT 59.79 5.64 59.96 5.81 ;
        RECT 60.25 5.64 60.42 5.81 ;
        RECT 60.71 5.64 60.88 5.81 ;
        RECT 61.17 5.64 61.34 5.81 ;
        RECT 61.63 5.64 61.8 5.81 ;
        RECT 65.33 6.835 65.5 7.005 ;
        RECT 65.33 5.465 65.5 5.635 ;
        RECT 66.035 6.835 66.205 7.005 ;
        RECT 66.035 5.465 66.205 5.635 ;
        RECT 67.025 6.835 67.195 7.005 ;
        RECT 67.025 5.465 67.195 5.635 ;
        RECT 70.69 6.835 70.86 7.005 ;
        RECT 71.775 5.645 71.945 5.815 ;
        RECT 72.235 5.645 72.405 5.815 ;
        RECT 72.695 5.645 72.865 5.815 ;
        RECT 73.155 5.645 73.325 5.815 ;
        RECT 73.615 5.645 73.785 5.815 ;
        RECT 74.075 5.645 74.245 5.815 ;
        RECT 74.535 5.645 74.705 5.815 ;
        RECT 74.995 5.645 75.165 5.815 ;
        RECT 75.455 5.645 75.625 5.815 ;
        RECT 75.915 5.645 76.085 5.815 ;
        RECT 76.375 5.645 76.545 5.815 ;
        RECT 76.835 5.645 77.005 5.815 ;
        RECT 77.295 5.645 77.465 5.815 ;
        RECT 77.755 5.645 77.925 5.815 ;
        RECT 78.215 5.645 78.385 5.815 ;
        RECT 81.915 6.84 82.085 7.01 ;
        RECT 81.915 5.47 82.085 5.64 ;
        RECT 82.62 6.84 82.79 7.01 ;
        RECT 82.62 5.47 82.79 5.64 ;
        RECT 83.61 6.84 83.78 7.01 ;
        RECT 83.61 5.47 83.78 5.64 ;
        RECT 87.27 6.835 87.44 7.005 ;
        RECT 88.355 5.645 88.525 5.815 ;
        RECT 88.815 5.645 88.985 5.815 ;
        RECT 89.275 5.645 89.445 5.815 ;
        RECT 89.735 5.645 89.905 5.815 ;
        RECT 90.195 5.645 90.365 5.815 ;
        RECT 90.655 5.645 90.825 5.815 ;
        RECT 91.115 5.645 91.285 5.815 ;
        RECT 91.575 5.645 91.745 5.815 ;
        RECT 92.035 5.645 92.205 5.815 ;
        RECT 92.495 5.645 92.665 5.815 ;
        RECT 92.955 5.645 93.125 5.815 ;
        RECT 93.415 5.645 93.585 5.815 ;
        RECT 93.875 5.645 94.045 5.815 ;
        RECT 94.335 5.645 94.505 5.815 ;
        RECT 94.795 5.645 94.965 5.815 ;
        RECT 98.495 6.84 98.665 7.01 ;
        RECT 98.495 5.47 98.665 5.64 ;
        RECT 99.2 6.84 99.37 7.01 ;
        RECT 99.2 5.47 99.37 5.64 ;
        RECT 100.19 6.84 100.36 7.01 ;
        RECT 100.19 5.47 100.36 5.64 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 90.585 7.735 90.92 8.11 ;
        RECT 90.555 7.795 90.895 8.205 ;
        RECT 90.58 7.77 90.92 8.11 ;
        RECT 90.115 7.795 90.92 8.095 ;
        RECT 74.005 7.735 74.34 8.11 ;
        RECT 73.975 7.795 74.315 8.205 ;
        RECT 74 7.77 74.34 8.11 ;
        RECT 73.535 7.795 74.34 8.095 ;
        RECT 57.42 7.73 57.755 8.105 ;
        RECT 57.39 7.79 57.73 8.2 ;
        RECT 57.415 7.765 57.755 8.105 ;
        RECT 56.95 7.79 57.755 8.09 ;
        RECT 40.835 7.725 41.17 8.1 ;
        RECT 40.805 7.785 41.145 8.195 ;
        RECT 40.83 7.76 41.17 8.1 ;
        RECT 40.365 7.785 41.17 8.085 ;
        RECT 24.25 7.725 24.585 8.1 ;
        RECT 24.22 7.785 24.56 8.195 ;
        RECT 24.245 7.76 24.585 8.1 ;
        RECT 23.78 7.785 24.585 8.085 ;
      LAYER met2 ;
        RECT 90.615 7.73 90.895 8.105 ;
        RECT 74.035 7.73 74.315 8.105 ;
        RECT 57.45 7.725 57.73 8.1 ;
        RECT 40.865 7.72 41.145 8.095 ;
        RECT 24.28 7.72 24.56 8.095 ;
      LAYER li1 ;
        RECT 67.92 0 101.085 1.61 ;
        RECT 100.11 0 100.28 2.24 ;
        RECT 99.12 0 99.29 2.24 ;
        RECT 96.375 0 96.545 2.24 ;
        RECT 87.96 0 95.305 3.105 ;
        RECT 94.745 0 95.015 3.905 ;
        RECT 93.835 0 94.075 3.905 ;
        RECT 92.965 0 93.215 3.635 ;
        RECT 90.585 0 90.915 3.555 ;
        RECT 88.295 0 88.555 3.915 ;
        RECT 83.53 0 83.7 2.24 ;
        RECT 82.54 0 82.71 2.24 ;
        RECT 79.795 0 79.965 2.24 ;
        RECT 71.38 0 78.725 3.105 ;
        RECT 78.165 0 78.435 3.905 ;
        RECT 77.255 0 77.495 3.905 ;
        RECT 76.385 0 76.635 3.635 ;
        RECT 74.005 0 74.335 3.555 ;
        RECT 71.715 0 71.975 3.915 ;
        RECT 51.335 0 101.085 1.605 ;
        RECT 66.945 0 67.115 2.235 ;
        RECT 65.955 0 66.125 2.235 ;
        RECT 63.21 0 63.38 2.235 ;
        RECT 54.795 0 62.14 3.1 ;
        RECT 61.58 0 61.85 3.9 ;
        RECT 60.67 0 60.91 3.9 ;
        RECT 59.8 0 60.05 3.63 ;
        RECT 57.42 0 57.75 3.55 ;
        RECT 55.13 0 55.39 3.91 ;
        RECT 0 0 101.085 1.6 ;
        RECT 50.36 0 50.53 2.23 ;
        RECT 49.37 0 49.54 2.23 ;
        RECT 46.625 0 46.795 2.23 ;
        RECT 38.21 0 45.555 3.095 ;
        RECT 44.995 0 45.265 3.895 ;
        RECT 44.085 0 44.325 3.895 ;
        RECT 43.215 0 43.465 3.625 ;
        RECT 40.835 0 41.165 3.545 ;
        RECT 38.545 0 38.805 3.905 ;
        RECT 33.775 0 33.945 2.23 ;
        RECT 32.785 0 32.955 2.23 ;
        RECT 30.04 0 30.21 2.23 ;
        RECT 21.625 0 28.97 3.095 ;
        RECT 28.41 0 28.68 3.895 ;
        RECT 27.5 0 27.74 3.895 ;
        RECT 26.63 0 26.88 3.625 ;
        RECT 24.25 0 24.58 3.545 ;
        RECT 21.96 0 22.22 3.905 ;
        RECT 67.92 10.86 101.085 12.47 ;
        RECT 100.11 10.24 100.28 12.47 ;
        RECT 99.12 10.24 99.29 12.47 ;
        RECT 96.375 10.24 96.545 12.47 ;
        RECT 88.22 9.475 95.12 12.47 ;
        RECT 88.215 8.365 95.115 9.475 ;
        RECT 93.645 7.855 94.095 12.47 ;
        RECT 91.555 7.965 91.885 12.47 ;
        RECT 89.485 7.905 89.735 12.47 ;
        RECT 85.15 10.235 85.32 12.47 ;
        RECT 83.53 10.24 83.7 12.47 ;
        RECT 82.54 10.24 82.71 12.47 ;
        RECT 79.795 10.24 79.965 12.47 ;
        RECT 71.64 9.475 78.54 12.47 ;
        RECT 71.635 8.365 78.535 9.475 ;
        RECT 77.065 7.855 77.515 12.47 ;
        RECT 74.975 7.965 75.305 12.47 ;
        RECT 72.905 7.905 73.155 12.47 ;
        RECT 68.57 10.235 68.74 12.47 ;
        RECT 51.335 10.86 101.085 12.465 ;
        RECT 66.945 10.235 67.115 12.465 ;
        RECT 65.955 10.235 66.125 12.465 ;
        RECT 63.21 10.235 63.38 12.465 ;
        RECT 55.055 9.47 61.955 12.465 ;
        RECT 55.05 8.36 61.95 9.47 ;
        RECT 60.48 7.85 60.93 12.465 ;
        RECT 58.39 7.96 58.72 12.465 ;
        RECT 56.32 7.9 56.57 12.465 ;
        RECT 51.985 10.23 52.155 12.465 ;
        RECT 0 10.86 101.085 12.46 ;
        RECT 50.36 10.23 50.53 12.46 ;
        RECT 49.37 10.23 49.54 12.46 ;
        RECT 46.625 10.23 46.795 12.46 ;
        RECT 38.47 9.465 45.37 12.46 ;
        RECT 38.465 8.355 45.365 9.465 ;
        RECT 43.895 7.845 44.345 12.46 ;
        RECT 41.805 7.955 42.135 12.46 ;
        RECT 39.735 7.895 39.985 12.46 ;
        RECT 35.23 10.855 37.98 12.46 ;
        RECT 35.4 10.225 35.57 12.46 ;
        RECT 33.775 10.23 33.945 12.46 ;
        RECT 32.785 10.23 32.955 12.46 ;
        RECT 30.04 10.23 30.21 12.46 ;
        RECT 21.885 9.465 28.785 12.46 ;
        RECT 21.88 8.355 28.78 9.465 ;
        RECT 27.31 7.845 27.76 12.46 ;
        RECT 25.22 7.955 25.55 12.46 ;
        RECT 23.15 7.895 23.4 12.46 ;
        RECT 18.645 10.855 21.395 12.46 ;
        RECT 18.815 10.225 18.985 12.46 ;
        RECT 15.415 10.855 18.165 12.46 ;
        RECT 15.585 10.225 15.755 12.46 ;
        RECT 91.855 7.125 92.185 7.455 ;
        RECT 89.635 7.125 89.975 7.375 ;
        RECT 86.165 8.365 86.335 10.315 ;
        RECT 86.105 10.145 86.275 10.595 ;
        RECT 86.105 7.305 86.275 8.535 ;
        RECT 75.275 7.125 75.605 7.455 ;
        RECT 73.055 7.125 73.395 7.375 ;
        RECT 69.585 8.365 69.755 10.315 ;
        RECT 69.525 10.145 69.695 10.595 ;
        RECT 69.525 7.305 69.695 8.535 ;
        RECT 58.69 7.12 59.02 7.45 ;
        RECT 56.47 7.12 56.81 7.37 ;
        RECT 53 8.36 53.17 10.31 ;
        RECT 52.94 10.14 53.11 10.59 ;
        RECT 52.94 7.3 53.11 8.53 ;
        RECT 42.105 7.115 42.435 7.445 ;
        RECT 39.885 7.115 40.225 7.365 ;
        RECT 36.415 8.355 36.585 10.305 ;
        RECT 36.355 10.135 36.525 10.585 ;
        RECT 36.355 7.295 36.525 8.525 ;
        RECT 25.52 7.115 25.85 7.445 ;
        RECT 23.3 7.115 23.64 7.365 ;
        RECT 19.83 8.355 20 10.305 ;
        RECT 19.77 10.135 19.94 10.585 ;
        RECT 19.77 7.295 19.94 8.525 ;
      LAYER met1 ;
        RECT 67.92 0 101.085 1.61 ;
        RECT 87.96 0 95.305 3.135 ;
        RECT 71.38 0 78.725 3.135 ;
        RECT 51.335 0 101.085 1.605 ;
        RECT 54.795 0 62.14 3.13 ;
        RECT 0 0 101.085 1.6 ;
        RECT 38.21 0 45.555 3.125 ;
        RECT 21.625 0 28.97 3.125 ;
        RECT 67.92 10.86 101.085 12.47 ;
        RECT 88.22 9.475 95.12 12.47 ;
        RECT 88.215 8.335 95.115 9.475 ;
        RECT 91.805 7.145 92.095 7.375 ;
        RECT 89.675 7.815 92.025 7.955 ;
        RECT 91.885 7.145 92.025 7.955 ;
        RECT 90.605 7.815 91.035 8.055 ;
        RECT 90.64 7.815 90.9 12.47 ;
        RECT 90.615 7.79 90.895 8.055 ;
        RECT 90.635 7.76 90.895 8.055 ;
        RECT 89.595 7.145 89.885 7.375 ;
        RECT 89.675 7.145 89.815 7.955 ;
        RECT 86.105 8.575 86.395 8.805 ;
        RECT 85.94 8.605 86.11 12.47 ;
        RECT 85.93 8.605 86.395 8.775 ;
        RECT 71.64 9.475 78.54 12.47 ;
        RECT 71.635 8.335 78.535 9.475 ;
        RECT 75.225 7.145 75.515 7.375 ;
        RECT 73.095 7.815 75.445 7.955 ;
        RECT 75.305 7.145 75.445 7.955 ;
        RECT 74.025 7.815 74.455 8.055 ;
        RECT 74.06 7.815 74.32 12.47 ;
        RECT 74.035 7.79 74.315 8.055 ;
        RECT 74.055 7.76 74.315 8.055 ;
        RECT 73.015 7.145 73.305 7.375 ;
        RECT 73.095 7.145 73.235 7.955 ;
        RECT 69.525 8.575 69.815 8.805 ;
        RECT 69.36 8.605 69.53 12.47 ;
        RECT 69.35 8.605 69.815 8.775 ;
        RECT 51.335 10.86 101.085 12.465 ;
        RECT 55.055 9.47 61.955 12.465 ;
        RECT 55.05 8.33 61.95 9.47 ;
        RECT 58.64 7.14 58.93 7.37 ;
        RECT 56.51 7.81 58.86 7.95 ;
        RECT 58.72 7.14 58.86 7.95 ;
        RECT 57.44 7.81 57.87 8.05 ;
        RECT 57.475 7.81 57.735 12.465 ;
        RECT 57.45 7.785 57.73 8.05 ;
        RECT 57.47 7.755 57.73 8.05 ;
        RECT 56.43 7.14 56.72 7.37 ;
        RECT 56.51 7.14 56.65 7.95 ;
        RECT 52.94 8.57 53.23 8.8 ;
        RECT 52.775 10.855 52.95 12.465 ;
        RECT 52.775 8.6 52.945 12.465 ;
        RECT 52.765 8.6 53.23 8.77 ;
        RECT 0 10.86 101.085 12.46 ;
        RECT 38.47 9.465 45.37 12.46 ;
        RECT 38.465 8.325 45.365 9.465 ;
        RECT 42.055 7.135 42.345 7.365 ;
        RECT 39.925 7.805 42.275 7.945 ;
        RECT 42.135 7.135 42.275 7.945 ;
        RECT 40.855 7.805 41.285 8.045 ;
        RECT 40.89 7.805 41.15 12.46 ;
        RECT 40.865 7.78 41.145 8.045 ;
        RECT 40.885 7.75 41.145 8.045 ;
        RECT 39.845 7.135 40.135 7.365 ;
        RECT 39.925 7.135 40.065 7.945 ;
        RECT 35.23 10.855 37.98 12.46 ;
        RECT 36.355 8.565 36.645 8.795 ;
        RECT 36.19 10.85 36.365 12.46 ;
        RECT 36.19 8.595 36.36 12.46 ;
        RECT 36.18 8.595 36.645 8.765 ;
        RECT 21.885 9.465 28.785 12.46 ;
        RECT 21.88 8.325 28.78 9.465 ;
        RECT 25.47 7.135 25.76 7.365 ;
        RECT 23.34 7.805 25.69 7.945 ;
        RECT 25.55 7.135 25.69 7.945 ;
        RECT 24.27 7.805 24.7 8.045 ;
        RECT 24.305 7.805 24.565 12.46 ;
        RECT 24.28 7.78 24.56 8.045 ;
        RECT 24.3 7.75 24.56 8.045 ;
        RECT 23.26 7.135 23.55 7.365 ;
        RECT 23.34 7.135 23.48 7.945 ;
        RECT 18.645 10.855 21.395 12.46 ;
        RECT 19.77 8.565 20.06 8.795 ;
        RECT 19.605 10.85 19.78 12.46 ;
        RECT 19.605 8.595 19.775 12.46 ;
        RECT 19.595 8.595 20.06 8.765 ;
        RECT 15.415 10.855 18.165 12.46 ;
      LAYER via1 ;
        RECT 24.355 7.835 24.505 7.985 ;
        RECT 40.94 7.835 41.09 7.985 ;
        RECT 57.525 7.84 57.675 7.99 ;
        RECT 74.11 7.845 74.26 7.995 ;
        RECT 90.69 7.845 90.84 7.995 ;
      LAYER via2 ;
        RECT 24.32 7.81 24.52 8.01 ;
        RECT 40.905 7.81 41.105 8.01 ;
        RECT 57.49 7.815 57.69 8.015 ;
        RECT 74.075 7.82 74.275 8.02 ;
        RECT 90.655 7.82 90.855 8.02 ;
      LAYER mcon ;
        RECT 15.665 10.885 15.835 11.055 ;
        RECT 16.345 10.885 16.515 11.055 ;
        RECT 17.025 10.885 17.195 11.055 ;
        RECT 17.705 10.885 17.875 11.055 ;
        RECT 18.895 10.885 19.065 11.055 ;
        RECT 19.575 10.885 19.745 11.055 ;
        RECT 19.83 8.595 20 8.765 ;
        RECT 20.255 10.885 20.425 11.055 ;
        RECT 20.935 10.885 21.105 11.055 ;
        RECT 22.02 8.355 22.19 8.525 ;
        RECT 22.02 2.925 22.19 3.095 ;
        RECT 22.48 8.355 22.65 8.525 ;
        RECT 22.48 2.925 22.65 3.095 ;
        RECT 22.94 8.355 23.11 8.525 ;
        RECT 22.94 2.925 23.11 3.095 ;
        RECT 23.32 7.165 23.49 7.335 ;
        RECT 23.4 8.355 23.57 8.525 ;
        RECT 23.4 2.925 23.57 3.095 ;
        RECT 23.86 8.355 24.03 8.525 ;
        RECT 23.86 2.925 24.03 3.095 ;
        RECT 24.32 8.355 24.49 8.525 ;
        RECT 24.32 2.925 24.49 3.095 ;
        RECT 24.78 8.355 24.95 8.525 ;
        RECT 24.78 2.925 24.95 3.095 ;
        RECT 25.24 8.355 25.41 8.525 ;
        RECT 25.24 2.925 25.41 3.095 ;
        RECT 25.53 7.165 25.7 7.335 ;
        RECT 25.7 8.355 25.87 8.525 ;
        RECT 25.7 2.925 25.87 3.095 ;
        RECT 26.16 8.355 26.33 8.525 ;
        RECT 26.16 2.925 26.33 3.095 ;
        RECT 26.62 8.355 26.79 8.525 ;
        RECT 26.62 2.925 26.79 3.095 ;
        RECT 27.08 8.355 27.25 8.525 ;
        RECT 27.08 2.925 27.25 3.095 ;
        RECT 27.54 8.355 27.71 8.525 ;
        RECT 27.54 2.925 27.71 3.095 ;
        RECT 28 8.355 28.17 8.525 ;
        RECT 28 2.925 28.17 3.095 ;
        RECT 28.46 8.355 28.63 8.525 ;
        RECT 28.46 2.925 28.63 3.095 ;
        RECT 30.12 10.89 30.29 11.06 ;
        RECT 30.12 1.4 30.29 1.57 ;
        RECT 30.8 10.89 30.97 11.06 ;
        RECT 30.8 1.4 30.97 1.57 ;
        RECT 31.48 10.89 31.65 11.06 ;
        RECT 31.48 1.4 31.65 1.57 ;
        RECT 32.16 10.89 32.33 11.06 ;
        RECT 32.16 1.4 32.33 1.57 ;
        RECT 32.865 10.89 33.035 11.06 ;
        RECT 32.865 1.4 33.035 1.57 ;
        RECT 33.855 10.89 34.025 11.06 ;
        RECT 33.855 1.4 34.025 1.57 ;
        RECT 35.48 10.885 35.65 11.055 ;
        RECT 36.16 10.885 36.33 11.055 ;
        RECT 36.415 8.595 36.585 8.765 ;
        RECT 36.84 10.885 37.01 11.055 ;
        RECT 37.52 10.885 37.69 11.055 ;
        RECT 38.605 8.355 38.775 8.525 ;
        RECT 38.605 2.925 38.775 3.095 ;
        RECT 39.065 8.355 39.235 8.525 ;
        RECT 39.065 2.925 39.235 3.095 ;
        RECT 39.525 8.355 39.695 8.525 ;
        RECT 39.525 2.925 39.695 3.095 ;
        RECT 39.905 7.165 40.075 7.335 ;
        RECT 39.985 8.355 40.155 8.525 ;
        RECT 39.985 2.925 40.155 3.095 ;
        RECT 40.445 8.355 40.615 8.525 ;
        RECT 40.445 2.925 40.615 3.095 ;
        RECT 40.905 8.355 41.075 8.525 ;
        RECT 40.905 2.925 41.075 3.095 ;
        RECT 41.365 8.355 41.535 8.525 ;
        RECT 41.365 2.925 41.535 3.095 ;
        RECT 41.825 8.355 41.995 8.525 ;
        RECT 41.825 2.925 41.995 3.095 ;
        RECT 42.115 7.165 42.285 7.335 ;
        RECT 42.285 8.355 42.455 8.525 ;
        RECT 42.285 2.925 42.455 3.095 ;
        RECT 42.745 8.355 42.915 8.525 ;
        RECT 42.745 2.925 42.915 3.095 ;
        RECT 43.205 8.355 43.375 8.525 ;
        RECT 43.205 2.925 43.375 3.095 ;
        RECT 43.665 8.355 43.835 8.525 ;
        RECT 43.665 2.925 43.835 3.095 ;
        RECT 44.125 8.355 44.295 8.525 ;
        RECT 44.125 2.925 44.295 3.095 ;
        RECT 44.585 8.355 44.755 8.525 ;
        RECT 44.585 2.925 44.755 3.095 ;
        RECT 45.045 8.355 45.215 8.525 ;
        RECT 45.045 2.925 45.215 3.095 ;
        RECT 46.705 10.89 46.875 11.06 ;
        RECT 46.705 1.4 46.875 1.57 ;
        RECT 47.385 10.89 47.555 11.06 ;
        RECT 47.385 1.4 47.555 1.57 ;
        RECT 48.065 10.89 48.235 11.06 ;
        RECT 48.065 1.4 48.235 1.57 ;
        RECT 48.745 10.89 48.915 11.06 ;
        RECT 48.745 1.4 48.915 1.57 ;
        RECT 49.45 10.89 49.62 11.06 ;
        RECT 49.45 1.4 49.62 1.57 ;
        RECT 50.44 10.89 50.61 11.06 ;
        RECT 50.44 1.4 50.61 1.57 ;
        RECT 52.065 10.89 52.235 11.06 ;
        RECT 52.745 10.89 52.915 11.06 ;
        RECT 53 8.6 53.17 8.77 ;
        RECT 53.425 10.89 53.595 11.06 ;
        RECT 54.105 10.89 54.275 11.06 ;
        RECT 55.19 8.36 55.36 8.53 ;
        RECT 55.19 2.93 55.36 3.1 ;
        RECT 55.65 8.36 55.82 8.53 ;
        RECT 55.65 2.93 55.82 3.1 ;
        RECT 56.11 8.36 56.28 8.53 ;
        RECT 56.11 2.93 56.28 3.1 ;
        RECT 56.49 7.17 56.66 7.34 ;
        RECT 56.57 8.36 56.74 8.53 ;
        RECT 56.57 2.93 56.74 3.1 ;
        RECT 57.03 8.36 57.2 8.53 ;
        RECT 57.03 2.93 57.2 3.1 ;
        RECT 57.49 8.36 57.66 8.53 ;
        RECT 57.49 2.93 57.66 3.1 ;
        RECT 57.95 8.36 58.12 8.53 ;
        RECT 57.95 2.93 58.12 3.1 ;
        RECT 58.41 8.36 58.58 8.53 ;
        RECT 58.41 2.93 58.58 3.1 ;
        RECT 58.7 7.17 58.87 7.34 ;
        RECT 58.87 8.36 59.04 8.53 ;
        RECT 58.87 2.93 59.04 3.1 ;
        RECT 59.33 8.36 59.5 8.53 ;
        RECT 59.33 2.93 59.5 3.1 ;
        RECT 59.79 8.36 59.96 8.53 ;
        RECT 59.79 2.93 59.96 3.1 ;
        RECT 60.25 8.36 60.42 8.53 ;
        RECT 60.25 2.93 60.42 3.1 ;
        RECT 60.71 8.36 60.88 8.53 ;
        RECT 60.71 2.93 60.88 3.1 ;
        RECT 61.17 8.36 61.34 8.53 ;
        RECT 61.17 2.93 61.34 3.1 ;
        RECT 61.63 8.36 61.8 8.53 ;
        RECT 61.63 2.93 61.8 3.1 ;
        RECT 63.29 10.895 63.46 11.065 ;
        RECT 63.29 1.405 63.46 1.575 ;
        RECT 63.97 10.895 64.14 11.065 ;
        RECT 63.97 1.405 64.14 1.575 ;
        RECT 64.65 10.895 64.82 11.065 ;
        RECT 64.65 1.405 64.82 1.575 ;
        RECT 65.33 10.895 65.5 11.065 ;
        RECT 65.33 1.405 65.5 1.575 ;
        RECT 66.035 10.895 66.205 11.065 ;
        RECT 66.035 1.405 66.205 1.575 ;
        RECT 67.025 10.895 67.195 11.065 ;
        RECT 67.025 1.405 67.195 1.575 ;
        RECT 68.65 10.895 68.82 11.065 ;
        RECT 69.33 10.895 69.5 11.065 ;
        RECT 69.585 8.605 69.755 8.775 ;
        RECT 70.01 10.895 70.18 11.065 ;
        RECT 70.69 10.895 70.86 11.065 ;
        RECT 71.775 8.365 71.945 8.535 ;
        RECT 71.775 2.935 71.945 3.105 ;
        RECT 72.235 8.365 72.405 8.535 ;
        RECT 72.235 2.935 72.405 3.105 ;
        RECT 72.695 8.365 72.865 8.535 ;
        RECT 72.695 2.935 72.865 3.105 ;
        RECT 73.075 7.175 73.245 7.345 ;
        RECT 73.155 8.365 73.325 8.535 ;
        RECT 73.155 2.935 73.325 3.105 ;
        RECT 73.615 8.365 73.785 8.535 ;
        RECT 73.615 2.935 73.785 3.105 ;
        RECT 74.075 8.365 74.245 8.535 ;
        RECT 74.075 2.935 74.245 3.105 ;
        RECT 74.535 8.365 74.705 8.535 ;
        RECT 74.535 2.935 74.705 3.105 ;
        RECT 74.995 8.365 75.165 8.535 ;
        RECT 74.995 2.935 75.165 3.105 ;
        RECT 75.285 7.175 75.455 7.345 ;
        RECT 75.455 8.365 75.625 8.535 ;
        RECT 75.455 2.935 75.625 3.105 ;
        RECT 75.915 8.365 76.085 8.535 ;
        RECT 75.915 2.935 76.085 3.105 ;
        RECT 76.375 8.365 76.545 8.535 ;
        RECT 76.375 2.935 76.545 3.105 ;
        RECT 76.835 8.365 77.005 8.535 ;
        RECT 76.835 2.935 77.005 3.105 ;
        RECT 77.295 8.365 77.465 8.535 ;
        RECT 77.295 2.935 77.465 3.105 ;
        RECT 77.755 8.365 77.925 8.535 ;
        RECT 77.755 2.935 77.925 3.105 ;
        RECT 78.215 8.365 78.385 8.535 ;
        RECT 78.215 2.935 78.385 3.105 ;
        RECT 79.875 10.9 80.045 11.07 ;
        RECT 79.875 1.41 80.045 1.58 ;
        RECT 80.555 10.9 80.725 11.07 ;
        RECT 80.555 1.41 80.725 1.58 ;
        RECT 81.235 10.9 81.405 11.07 ;
        RECT 81.235 1.41 81.405 1.58 ;
        RECT 81.915 10.9 82.085 11.07 ;
        RECT 81.915 1.41 82.085 1.58 ;
        RECT 82.62 10.9 82.79 11.07 ;
        RECT 82.62 1.41 82.79 1.58 ;
        RECT 83.61 10.9 83.78 11.07 ;
        RECT 83.61 1.41 83.78 1.58 ;
        RECT 85.23 10.895 85.4 11.065 ;
        RECT 85.91 10.895 86.08 11.065 ;
        RECT 86.165 8.605 86.335 8.775 ;
        RECT 86.59 10.895 86.76 11.065 ;
        RECT 87.27 10.895 87.44 11.065 ;
        RECT 88.355 8.365 88.525 8.535 ;
        RECT 88.355 2.935 88.525 3.105 ;
        RECT 88.815 8.365 88.985 8.535 ;
        RECT 88.815 2.935 88.985 3.105 ;
        RECT 89.275 8.365 89.445 8.535 ;
        RECT 89.275 2.935 89.445 3.105 ;
        RECT 89.655 7.175 89.825 7.345 ;
        RECT 89.735 8.365 89.905 8.535 ;
        RECT 89.735 2.935 89.905 3.105 ;
        RECT 90.195 8.365 90.365 8.535 ;
        RECT 90.195 2.935 90.365 3.105 ;
        RECT 90.655 8.365 90.825 8.535 ;
        RECT 90.655 2.935 90.825 3.105 ;
        RECT 91.115 8.365 91.285 8.535 ;
        RECT 91.115 2.935 91.285 3.105 ;
        RECT 91.575 8.365 91.745 8.535 ;
        RECT 91.575 2.935 91.745 3.105 ;
        RECT 91.865 7.175 92.035 7.345 ;
        RECT 92.035 8.365 92.205 8.535 ;
        RECT 92.035 2.935 92.205 3.105 ;
        RECT 92.495 8.365 92.665 8.535 ;
        RECT 92.495 2.935 92.665 3.105 ;
        RECT 92.955 8.365 93.125 8.535 ;
        RECT 92.955 2.935 93.125 3.105 ;
        RECT 93.415 8.365 93.585 8.535 ;
        RECT 93.415 2.935 93.585 3.105 ;
        RECT 93.875 8.365 94.045 8.535 ;
        RECT 93.875 2.935 94.045 3.105 ;
        RECT 94.335 8.365 94.505 8.535 ;
        RECT 94.335 2.935 94.505 3.105 ;
        RECT 94.795 8.365 94.965 8.535 ;
        RECT 94.795 2.935 94.965 3.105 ;
        RECT 96.455 10.9 96.625 11.07 ;
        RECT 96.455 1.41 96.625 1.58 ;
        RECT 97.135 10.9 97.305 11.07 ;
        RECT 97.135 1.41 97.305 1.58 ;
        RECT 97.815 10.9 97.985 11.07 ;
        RECT 97.815 1.41 97.985 1.58 ;
        RECT 98.495 10.9 98.665 11.07 ;
        RECT 98.495 1.41 98.665 1.58 ;
        RECT 99.2 10.9 99.37 11.07 ;
        RECT 99.2 1.41 99.37 1.58 ;
        RECT 100.19 10.9 100.36 11.07 ;
        RECT 100.19 1.41 100.36 1.58 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 92.98 4.03 93.32 4.37 ;
      RECT 92.98 4.055 93.785 4.355 ;
      RECT 86.435 9.29 86.805 9.66 ;
      RECT 86.435 9.325 91.59 9.625 ;
      RECT 91.285 7.09 91.585 9.625 ;
      RECT 92.3 7.09 92.64 7.43 ;
      RECT 90.66 7.09 91.6 7.43 ;
      RECT 90.66 7.115 93.105 7.415 ;
      RECT 90.66 7.1 92.64 7.415 ;
      RECT 90.66 5.07 90.99 7.43 ;
      RECT 90.66 5.07 93.31 5.4 ;
      RECT 90.66 5.07 93.315 5.395 ;
      RECT 92.975 5.05 93.32 5.39 ;
      RECT 90.66 5.075 93.785 5.375 ;
      RECT 92.995 5.005 93.295 5.4 ;
      RECT 92.285 4.365 92.625 4.715 ;
      RECT 91.815 4.395 92.625 4.695 ;
      RECT 91.62 6.07 91.96 6.41 ;
      RECT 91.62 6.095 92.425 6.395 ;
      RECT 90.94 3.69 91.28 4.03 ;
      RECT 90.475 3.715 91.28 4.015 ;
      RECT 90.835 3.705 91.28 4.015 ;
      RECT 76.4 4.03 76.74 4.37 ;
      RECT 76.4 4.055 77.205 4.355 ;
      RECT 69.855 9.29 70.225 9.66 ;
      RECT 69.855 9.325 75.01 9.625 ;
      RECT 74.705 7.09 75.005 9.625 ;
      RECT 75.72 7.09 76.06 7.43 ;
      RECT 74.08 7.09 75.02 7.43 ;
      RECT 74.08 7.115 76.525 7.415 ;
      RECT 74.08 7.1 76.06 7.415 ;
      RECT 74.08 5.07 74.41 7.43 ;
      RECT 74.08 5.07 76.73 5.4 ;
      RECT 74.08 5.07 76.735 5.395 ;
      RECT 76.395 5.05 76.74 5.39 ;
      RECT 74.08 5.075 77.205 5.375 ;
      RECT 76.415 5.005 76.715 5.4 ;
      RECT 75.705 4.365 76.045 4.715 ;
      RECT 75.235 4.395 76.045 4.695 ;
      RECT 75.04 6.07 75.38 6.41 ;
      RECT 75.04 6.095 75.845 6.395 ;
      RECT 74.36 3.69 74.7 4.03 ;
      RECT 73.895 3.715 74.7 4.015 ;
      RECT 74.255 3.705 74.7 4.015 ;
      RECT 59.815 4.025 60.155 4.365 ;
      RECT 59.815 4.05 60.62 4.35 ;
      RECT 53.27 9.285 53.64 9.655 ;
      RECT 53.27 9.32 58.425 9.62 ;
      RECT 58.12 7.085 58.42 9.62 ;
      RECT 59.135 7.085 59.475 7.425 ;
      RECT 57.495 7.085 58.435 7.425 ;
      RECT 57.495 7.11 59.94 7.41 ;
      RECT 57.495 7.095 59.475 7.41 ;
      RECT 57.495 5.065 57.825 7.425 ;
      RECT 57.495 5.065 60.145 5.395 ;
      RECT 57.495 5.065 60.15 5.39 ;
      RECT 59.81 5.045 60.155 5.385 ;
      RECT 57.495 5.07 60.62 5.37 ;
      RECT 59.83 5 60.13 5.395 ;
      RECT 59.12 4.36 59.46 4.71 ;
      RECT 58.65 4.39 59.46 4.69 ;
      RECT 58.455 6.065 58.795 6.405 ;
      RECT 58.455 6.09 59.26 6.39 ;
      RECT 57.775 3.685 58.115 4.025 ;
      RECT 57.31 3.71 58.115 4.01 ;
      RECT 57.67 3.7 58.115 4.01 ;
      RECT 43.23 4.02 43.57 4.36 ;
      RECT 43.23 4.045 44.035 4.345 ;
      RECT 36.685 9.28 37.055 9.65 ;
      RECT 36.685 9.315 41.84 9.615 ;
      RECT 41.535 7.08 41.835 9.615 ;
      RECT 42.55 7.08 42.89 7.42 ;
      RECT 40.91 7.08 41.85 7.42 ;
      RECT 40.91 7.105 43.355 7.405 ;
      RECT 40.91 7.09 42.89 7.405 ;
      RECT 40.91 5.06 41.24 7.42 ;
      RECT 40.91 5.06 43.56 5.39 ;
      RECT 40.91 5.06 43.565 5.385 ;
      RECT 43.225 5.04 43.57 5.38 ;
      RECT 40.91 5.065 44.035 5.365 ;
      RECT 43.245 4.995 43.545 5.39 ;
      RECT 42.535 4.355 42.875 4.705 ;
      RECT 42.065 4.385 42.875 4.685 ;
      RECT 41.87 6.06 42.21 6.4 ;
      RECT 41.87 6.085 42.675 6.385 ;
      RECT 41.19 3.68 41.53 4.02 ;
      RECT 40.725 3.705 41.53 4.005 ;
      RECT 41.085 3.695 41.53 4.005 ;
      RECT 26.645 4.02 26.985 4.36 ;
      RECT 26.645 4.045 27.45 4.345 ;
      RECT 20.1 9.28 20.47 9.65 ;
      RECT 20.1 9.315 25.255 9.615 ;
      RECT 24.95 7.08 25.25 9.615 ;
      RECT 25.965 7.08 26.305 7.42 ;
      RECT 24.325 7.08 25.265 7.42 ;
      RECT 24.325 7.105 26.77 7.405 ;
      RECT 24.325 7.09 26.305 7.405 ;
      RECT 24.325 5.06 24.655 7.42 ;
      RECT 24.325 5.06 26.975 5.39 ;
      RECT 24.325 5.06 26.98 5.385 ;
      RECT 26.64 5.04 26.985 5.38 ;
      RECT 24.325 5.065 27.45 5.365 ;
      RECT 26.66 4.995 26.96 5.39 ;
      RECT 25.95 4.355 26.29 4.705 ;
      RECT 25.48 4.385 26.29 4.685 ;
      RECT 25.285 6.06 25.625 6.4 ;
      RECT 25.285 6.085 26.09 6.385 ;
      RECT 24.605 3.68 24.945 4.02 ;
      RECT 24.14 3.705 24.945 4.005 ;
      RECT 24.5 3.695 24.945 4.005 ;
      RECT 100.44 7.215 100.82 12.47 ;
      RECT 83.86 7.215 84.24 12.47 ;
      RECT 67.275 7.21 67.655 12.465 ;
      RECT 50.69 7.205 51.07 12.46 ;
      RECT 34.105 7.205 34.485 12.46 ;
    LAYER via2 ;
      RECT 100.53 7.305 100.73 7.505 ;
      RECT 93.055 4.105 93.255 4.305 ;
      RECT 93.055 5.125 93.255 5.325 ;
      RECT 92.375 7.165 92.575 7.365 ;
      RECT 92.355 4.445 92.555 4.645 ;
      RECT 91.695 6.145 91.895 6.345 ;
      RECT 91.325 7.165 91.525 7.365 ;
      RECT 91.015 3.755 91.215 3.955 ;
      RECT 86.52 9.375 86.72 9.575 ;
      RECT 83.95 7.305 84.15 7.505 ;
      RECT 76.475 4.105 76.675 4.305 ;
      RECT 76.475 5.125 76.675 5.325 ;
      RECT 75.795 7.165 75.995 7.365 ;
      RECT 75.775 4.445 75.975 4.645 ;
      RECT 75.115 6.145 75.315 6.345 ;
      RECT 74.745 7.165 74.945 7.365 ;
      RECT 74.435 3.755 74.635 3.955 ;
      RECT 69.94 9.375 70.14 9.575 ;
      RECT 67.365 7.3 67.565 7.5 ;
      RECT 59.89 4.1 60.09 4.3 ;
      RECT 59.89 5.12 60.09 5.32 ;
      RECT 59.21 7.16 59.41 7.36 ;
      RECT 59.19 4.44 59.39 4.64 ;
      RECT 58.53 6.14 58.73 6.34 ;
      RECT 58.16 7.16 58.36 7.36 ;
      RECT 57.85 3.75 58.05 3.95 ;
      RECT 53.355 9.37 53.555 9.57 ;
      RECT 50.78 7.295 50.98 7.495 ;
      RECT 43.305 4.095 43.505 4.295 ;
      RECT 43.305 5.115 43.505 5.315 ;
      RECT 42.625 7.155 42.825 7.355 ;
      RECT 42.605 4.435 42.805 4.635 ;
      RECT 41.945 6.135 42.145 6.335 ;
      RECT 41.575 7.155 41.775 7.355 ;
      RECT 41.265 3.745 41.465 3.945 ;
      RECT 36.77 9.365 36.97 9.565 ;
      RECT 34.195 7.295 34.395 7.495 ;
      RECT 26.72 4.095 26.92 4.295 ;
      RECT 26.72 5.115 26.92 5.315 ;
      RECT 26.04 7.155 26.24 7.355 ;
      RECT 26.02 4.435 26.22 4.635 ;
      RECT 25.36 6.135 25.56 6.335 ;
      RECT 24.99 7.155 25.19 7.355 ;
      RECT 24.68 3.745 24.88 3.945 ;
      RECT 20.185 9.365 20.385 9.565 ;
    LAYER met2 ;
      RECT 16.575 10.065 100.715 10.235 ;
      RECT 100.545 9.585 100.715 10.235 ;
      RECT 16.575 8.54 16.745 10.235 ;
      RECT 100.51 9.585 100.835 9.91 ;
      RECT 16.535 8.54 16.815 8.88 ;
      RECT 97.355 8.575 97.675 8.9 ;
      RECT 97.385 7.99 97.555 8.9 ;
      RECT 97.385 7.99 97.56 8.34 ;
      RECT 97.385 7.99 98.36 8.165 ;
      RECT 98.185 3.27 98.36 8.165 ;
      RECT 98.13 3.27 98.48 3.62 ;
      RECT 87.02 9.715 97.2 9.885 ;
      RECT 97.04 3.7 97.2 9.885 ;
      RECT 87.02 8.895 87.19 9.885 ;
      RECT 83.965 8.955 84.29 9.28 ;
      RECT 98.155 8.95 98.48 9.275 ;
      RECT 86.965 8.895 87.245 9.235 ;
      RECT 97.04 9.04 98.48 9.21 ;
      RECT 83.965 8.985 84.84 9.155 ;
      RECT 84.84 8.97 87.245 9.14 ;
      RECT 97.355 3.67 97.675 3.99 ;
      RECT 97.04 3.7 97.675 3.87 ;
      RECT 90.975 3.665 91.255 4.05 ;
      RECT 91.02 2.91 91.19 4.05 ;
      RECT 95.685 3.3 96.01 3.625 ;
      RECT 95.76 2.91 95.93 3.625 ;
      RECT 91.02 2.91 95.93 3.08 ;
      RECT 94.715 6.085 94.975 6.405 ;
      RECT 94.775 4.045 94.915 6.405 ;
      RECT 94.715 4.045 94.975 4.365 ;
      RECT 93.695 7.105 93.955 7.425 ;
      RECT 93.075 7.195 93.955 7.335 ;
      RECT 93.075 5.035 93.215 7.335 ;
      RECT 93.015 5.035 93.295 5.41 ;
      RECT 92.335 7.075 92.615 7.45 ;
      RECT 92.395 5.155 92.535 7.45 ;
      RECT 92.395 5.155 92.875 5.295 ;
      RECT 92.735 3.365 92.875 5.295 ;
      RECT 92.675 3.365 92.935 3.705 ;
      RECT 91.655 6.055 91.935 6.43 ;
      RECT 91.715 3.705 91.855 6.43 ;
      RECT 91.655 3.705 91.915 4.025 ;
      RECT 91.285 7.075 91.565 7.45 ;
      RECT 91.285 7.105 91.575 7.425 ;
      RECT 86.435 9.29 86.81 9.66 ;
      RECT 86.44 9.28 86.81 9.66 ;
      RECT 80.775 8.575 81.095 8.9 ;
      RECT 80.805 7.99 80.975 8.9 ;
      RECT 80.805 7.99 80.98 8.34 ;
      RECT 80.805 7.99 81.78 8.165 ;
      RECT 81.605 3.27 81.78 8.165 ;
      RECT 81.55 3.27 81.9 3.62 ;
      RECT 70.44 9.715 80.62 9.885 ;
      RECT 80.46 3.7 80.62 9.885 ;
      RECT 70.44 8.895 70.61 9.885 ;
      RECT 81.575 8.95 81.9 9.275 ;
      RECT 67.38 8.95 67.705 9.275 ;
      RECT 70.385 8.895 70.665 9.235 ;
      RECT 80.46 9.04 81.9 9.21 ;
      RECT 67.38 8.98 68.305 9.15 ;
      RECT 68.305 8.97 70.665 9.14 ;
      RECT 80.775 3.67 81.095 3.99 ;
      RECT 80.46 3.7 81.095 3.87 ;
      RECT 74.395 3.665 74.675 4.05 ;
      RECT 74.44 2.91 74.61 4.05 ;
      RECT 79.105 3.3 79.43 3.625 ;
      RECT 79.18 2.91 79.35 3.625 ;
      RECT 74.44 2.91 79.35 3.08 ;
      RECT 78.135 6.085 78.395 6.405 ;
      RECT 78.195 4.045 78.335 6.405 ;
      RECT 78.135 4.045 78.395 4.365 ;
      RECT 77.115 7.105 77.375 7.425 ;
      RECT 76.495 7.195 77.375 7.335 ;
      RECT 76.495 5.035 76.635 7.335 ;
      RECT 76.435 5.035 76.715 5.41 ;
      RECT 75.755 7.075 76.035 7.45 ;
      RECT 75.815 5.155 75.955 7.45 ;
      RECT 75.815 5.155 76.295 5.295 ;
      RECT 76.155 3.365 76.295 5.295 ;
      RECT 76.095 3.365 76.355 3.705 ;
      RECT 75.075 6.055 75.355 6.43 ;
      RECT 75.135 3.705 75.275 6.43 ;
      RECT 75.075 3.705 75.335 4.025 ;
      RECT 74.705 7.075 74.985 7.45 ;
      RECT 74.705 7.105 74.995 7.425 ;
      RECT 64.19 8.57 64.51 8.895 ;
      RECT 64.22 7.985 64.39 8.895 ;
      RECT 64.22 7.985 64.395 8.335 ;
      RECT 64.22 7.985 65.195 8.16 ;
      RECT 65.02 3.265 65.195 8.16 ;
      RECT 64.965 3.265 65.315 3.615 ;
      RECT 53.855 9.71 64.035 9.88 ;
      RECT 63.875 3.695 64.035 9.88 ;
      RECT 53.855 8.89 54.025 9.88 ;
      RECT 64.99 8.945 65.315 9.27 ;
      RECT 50.795 8.945 51.12 9.27 ;
      RECT 53.8 8.89 54.08 9.23 ;
      RECT 63.875 9.035 65.315 9.205 ;
      RECT 50.795 8.975 52.075 9.145 ;
      RECT 52.075 8.97 54.08 9.14 ;
      RECT 64.19 3.665 64.51 3.985 ;
      RECT 63.875 3.695 64.51 3.865 ;
      RECT 57.81 3.66 58.09 4.045 ;
      RECT 57.855 2.905 58.025 4.045 ;
      RECT 62.52 3.295 62.845 3.62 ;
      RECT 62.595 2.905 62.765 3.62 ;
      RECT 57.855 2.905 62.765 3.075 ;
      RECT 61.55 6.08 61.81 6.4 ;
      RECT 61.61 4.04 61.75 6.4 ;
      RECT 61.55 4.04 61.81 4.36 ;
      RECT 60.53 7.1 60.79 7.42 ;
      RECT 59.91 7.19 60.79 7.33 ;
      RECT 59.91 5.03 60.05 7.33 ;
      RECT 59.85 5.03 60.13 5.405 ;
      RECT 59.17 7.07 59.45 7.445 ;
      RECT 59.23 5.15 59.37 7.445 ;
      RECT 59.23 5.15 59.71 5.29 ;
      RECT 59.57 3.36 59.71 5.29 ;
      RECT 59.51 3.36 59.77 3.7 ;
      RECT 58.49 6.05 58.77 6.425 ;
      RECT 58.55 3.7 58.69 6.425 ;
      RECT 58.49 3.7 58.75 4.02 ;
      RECT 58.12 7.07 58.4 7.445 ;
      RECT 58.12 7.1 58.41 7.42 ;
      RECT 47.605 8.565 47.925 8.89 ;
      RECT 47.635 7.98 47.805 8.89 ;
      RECT 47.635 7.98 47.81 8.33 ;
      RECT 47.635 7.98 48.61 8.155 ;
      RECT 48.435 3.26 48.61 8.155 ;
      RECT 48.38 3.26 48.73 3.61 ;
      RECT 37.27 9.705 47.45 9.875 ;
      RECT 47.29 3.69 47.45 9.875 ;
      RECT 37.27 8.885 37.44 9.875 ;
      RECT 34.21 8.945 34.535 9.27 ;
      RECT 48.405 8.94 48.73 9.265 ;
      RECT 37.215 8.885 37.495 9.225 ;
      RECT 47.29 9.03 48.73 9.2 ;
      RECT 34.21 8.975 35.26 9.145 ;
      RECT 35.26 8.97 37.495 9.14 ;
      RECT 47.605 3.66 47.925 3.98 ;
      RECT 47.29 3.69 47.925 3.86 ;
      RECT 41.225 3.655 41.505 4.04 ;
      RECT 41.27 2.9 41.44 4.04 ;
      RECT 45.935 3.29 46.26 3.615 ;
      RECT 46.01 2.9 46.18 3.615 ;
      RECT 41.27 2.9 46.18 3.07 ;
      RECT 44.965 6.075 45.225 6.395 ;
      RECT 45.025 4.035 45.165 6.395 ;
      RECT 44.965 4.035 45.225 4.355 ;
      RECT 43.945 7.095 44.205 7.415 ;
      RECT 43.325 7.185 44.205 7.325 ;
      RECT 43.325 5.025 43.465 7.325 ;
      RECT 43.265 5.025 43.545 5.4 ;
      RECT 42.585 7.065 42.865 7.44 ;
      RECT 42.645 5.145 42.785 7.44 ;
      RECT 42.645 5.145 43.125 5.285 ;
      RECT 42.985 3.355 43.125 5.285 ;
      RECT 42.925 3.355 43.185 3.695 ;
      RECT 41.905 6.045 42.185 6.42 ;
      RECT 41.965 3.695 42.105 6.42 ;
      RECT 41.905 3.695 42.165 4.015 ;
      RECT 41.535 7.065 41.815 7.44 ;
      RECT 41.535 7.095 41.825 7.415 ;
      RECT 31.02 8.565 31.34 8.89 ;
      RECT 31.05 7.98 31.22 8.89 ;
      RECT 31.05 7.98 31.225 8.33 ;
      RECT 31.05 7.98 32.025 8.155 ;
      RECT 31.85 3.26 32.025 8.155 ;
      RECT 31.795 3.26 32.145 3.61 ;
      RECT 20.685 9.705 30.865 9.875 ;
      RECT 30.705 3.69 30.865 9.875 ;
      RECT 20.685 8.885 20.855 9.875 ;
      RECT 16.92 9.28 17.2 9.62 ;
      RECT 16.92 9.345 18.11 9.515 ;
      RECT 17.94 8.97 18.11 9.515 ;
      RECT 31.82 8.94 32.145 9.265 ;
      RECT 20.63 8.885 20.91 9.225 ;
      RECT 30.705 9.03 32.145 9.2 ;
      RECT 17.94 8.97 20.91 9.14 ;
      RECT 31.02 3.66 31.34 3.98 ;
      RECT 30.705 3.69 31.34 3.86 ;
      RECT 24.64 3.655 24.92 4.04 ;
      RECT 24.685 2.9 24.855 4.04 ;
      RECT 29.35 3.29 29.675 3.615 ;
      RECT 29.425 2.9 29.595 3.615 ;
      RECT 24.685 2.9 29.595 3.07 ;
      RECT 28.38 6.075 28.64 6.395 ;
      RECT 28.44 4.035 28.58 6.395 ;
      RECT 28.38 4.035 28.64 4.355 ;
      RECT 27.36 7.095 27.62 7.415 ;
      RECT 26.74 7.185 27.62 7.325 ;
      RECT 26.74 5.025 26.88 7.325 ;
      RECT 26.68 5.025 26.96 5.4 ;
      RECT 26 7.065 26.28 7.44 ;
      RECT 26.06 5.145 26.2 7.44 ;
      RECT 26.06 5.145 26.54 5.285 ;
      RECT 26.4 3.355 26.54 5.285 ;
      RECT 26.34 3.355 26.6 3.695 ;
      RECT 25.32 6.045 25.6 6.42 ;
      RECT 25.38 3.695 25.52 6.42 ;
      RECT 25.32 3.695 25.58 4.015 ;
      RECT 24.95 7.065 25.23 7.44 ;
      RECT 24.95 7.095 25.24 7.415 ;
      RECT 100.44 7.215 100.82 7.595 ;
      RECT 93.015 4.015 93.295 4.39 ;
      RECT 92.315 4.355 92.595 4.73 ;
      RECT 83.86 7.215 84.24 7.595 ;
      RECT 76.435 4.015 76.715 4.39 ;
      RECT 75.735 4.355 76.015 4.73 ;
      RECT 69.855 9.28 70.225 9.66 ;
      RECT 67.275 7.21 67.655 7.59 ;
      RECT 59.85 4.01 60.13 4.385 ;
      RECT 59.15 4.35 59.43 4.725 ;
      RECT 53.27 9.28 53.64 9.655 ;
      RECT 50.69 7.205 51.07 7.585 ;
      RECT 43.265 4.005 43.545 4.38 ;
      RECT 42.565 4.345 42.845 4.72 ;
      RECT 36.685 9.28 37.055 9.65 ;
      RECT 34.105 7.205 34.485 7.585 ;
      RECT 26.68 4.005 26.96 4.38 ;
      RECT 25.98 4.345 26.26 4.72 ;
      RECT 20.1 9.28 20.47 9.65 ;
    LAYER via1 ;
      RECT 100.6 9.67 100.75 9.82 ;
      RECT 100.555 7.33 100.705 7.48 ;
      RECT 98.245 9.035 98.395 9.185 ;
      RECT 98.23 3.37 98.38 3.52 ;
      RECT 97.44 3.755 97.59 3.905 ;
      RECT 97.44 8.665 97.59 8.815 ;
      RECT 95.775 3.385 95.925 3.535 ;
      RECT 94.77 4.13 94.92 4.28 ;
      RECT 94.77 6.17 94.92 6.32 ;
      RECT 93.75 7.19 93.9 7.34 ;
      RECT 93.07 4.13 93.22 4.28 ;
      RECT 93.07 5.15 93.22 5.3 ;
      RECT 92.73 3.47 92.88 3.62 ;
      RECT 92.39 4.47 92.54 4.62 ;
      RECT 92.39 7.19 92.54 7.34 ;
      RECT 91.71 3.79 91.86 3.94 ;
      RECT 91.71 6.17 91.86 6.32 ;
      RECT 91.37 7.19 91.52 7.34 ;
      RECT 91.03 3.78 91.18 3.93 ;
      RECT 87.03 8.99 87.18 9.14 ;
      RECT 86.545 9.4 86.695 9.55 ;
      RECT 84.055 9.04 84.205 9.19 ;
      RECT 83.975 7.33 84.125 7.48 ;
      RECT 81.665 9.035 81.815 9.185 ;
      RECT 81.65 3.37 81.8 3.52 ;
      RECT 80.86 3.755 81.01 3.905 ;
      RECT 80.86 8.665 81.01 8.815 ;
      RECT 79.195 3.385 79.345 3.535 ;
      RECT 78.19 4.13 78.34 4.28 ;
      RECT 78.19 6.17 78.34 6.32 ;
      RECT 77.17 7.19 77.32 7.34 ;
      RECT 76.49 4.13 76.64 4.28 ;
      RECT 76.49 5.15 76.64 5.3 ;
      RECT 76.15 3.47 76.3 3.62 ;
      RECT 75.81 4.47 75.96 4.62 ;
      RECT 75.81 7.19 75.96 7.34 ;
      RECT 75.13 3.79 75.28 3.94 ;
      RECT 75.13 6.17 75.28 6.32 ;
      RECT 74.79 7.19 74.94 7.34 ;
      RECT 74.45 3.78 74.6 3.93 ;
      RECT 70.45 8.99 70.6 9.14 ;
      RECT 69.965 9.4 70.115 9.55 ;
      RECT 67.47 9.035 67.62 9.185 ;
      RECT 67.39 7.325 67.54 7.475 ;
      RECT 65.08 9.03 65.23 9.18 ;
      RECT 65.065 3.365 65.215 3.515 ;
      RECT 64.275 3.75 64.425 3.9 ;
      RECT 64.275 8.66 64.425 8.81 ;
      RECT 62.61 3.38 62.76 3.53 ;
      RECT 61.605 4.125 61.755 4.275 ;
      RECT 61.605 6.165 61.755 6.315 ;
      RECT 60.585 7.185 60.735 7.335 ;
      RECT 59.905 4.125 60.055 4.275 ;
      RECT 59.905 5.145 60.055 5.295 ;
      RECT 59.565 3.465 59.715 3.615 ;
      RECT 59.225 4.465 59.375 4.615 ;
      RECT 59.225 7.185 59.375 7.335 ;
      RECT 58.545 3.785 58.695 3.935 ;
      RECT 58.545 6.165 58.695 6.315 ;
      RECT 58.205 7.185 58.355 7.335 ;
      RECT 57.865 3.775 58.015 3.925 ;
      RECT 53.865 8.985 54.015 9.135 ;
      RECT 53.38 9.395 53.53 9.545 ;
      RECT 50.885 9.03 51.035 9.18 ;
      RECT 50.805 7.32 50.955 7.47 ;
      RECT 48.495 9.025 48.645 9.175 ;
      RECT 48.48 3.36 48.63 3.51 ;
      RECT 47.69 3.745 47.84 3.895 ;
      RECT 47.69 8.655 47.84 8.805 ;
      RECT 46.025 3.375 46.175 3.525 ;
      RECT 45.02 4.12 45.17 4.27 ;
      RECT 45.02 6.16 45.17 6.31 ;
      RECT 44 7.18 44.15 7.33 ;
      RECT 43.32 4.12 43.47 4.27 ;
      RECT 43.32 5.14 43.47 5.29 ;
      RECT 42.98 3.46 43.13 3.61 ;
      RECT 42.64 4.46 42.79 4.61 ;
      RECT 42.64 7.18 42.79 7.33 ;
      RECT 41.96 3.78 42.11 3.93 ;
      RECT 41.96 6.16 42.11 6.31 ;
      RECT 41.62 7.18 41.77 7.33 ;
      RECT 41.28 3.77 41.43 3.92 ;
      RECT 37.28 8.98 37.43 9.13 ;
      RECT 36.795 9.39 36.945 9.54 ;
      RECT 34.3 9.03 34.45 9.18 ;
      RECT 34.22 7.32 34.37 7.47 ;
      RECT 31.91 9.025 32.06 9.175 ;
      RECT 31.895 3.36 32.045 3.51 ;
      RECT 31.105 3.745 31.255 3.895 ;
      RECT 31.105 8.655 31.255 8.805 ;
      RECT 29.44 3.375 29.59 3.525 ;
      RECT 28.435 4.12 28.585 4.27 ;
      RECT 28.435 6.16 28.585 6.31 ;
      RECT 27.415 7.18 27.565 7.33 ;
      RECT 26.735 4.12 26.885 4.27 ;
      RECT 26.735 5.14 26.885 5.29 ;
      RECT 26.395 3.46 26.545 3.61 ;
      RECT 26.055 4.46 26.205 4.61 ;
      RECT 26.055 7.18 26.205 7.33 ;
      RECT 25.375 3.78 25.525 3.93 ;
      RECT 25.375 6.16 25.525 6.31 ;
      RECT 25.035 7.18 25.185 7.33 ;
      RECT 24.695 3.77 24.845 3.92 ;
      RECT 20.695 8.98 20.845 9.13 ;
      RECT 20.21 9.39 20.36 9.54 ;
      RECT 16.985 9.375 17.135 9.525 ;
      RECT 16.6 8.635 16.75 8.785 ;
    LAYER met1 ;
      RECT 100.48 10.06 100.775 10.29 ;
      RECT 100.54 9.585 100.715 10.29 ;
      RECT 100.51 9.585 100.835 9.91 ;
      RECT 100.54 8.58 100.71 10.29 ;
      RECT 100.48 8.58 100.77 8.81 ;
      RECT 100.075 4.04 100.4 4.27 ;
      RECT 100.075 4.07 100.57 4.24 ;
      RECT 100.075 3.7 100.265 4.27 ;
      RECT 99.49 3.67 99.78 3.9 ;
      RECT 99.49 3.7 100.265 3.87 ;
      RECT 99.55 2.19 99.72 3.9 ;
      RECT 99.49 2.19 99.785 2.42 ;
      RECT 99.49 10.06 99.785 10.29 ;
      RECT 99.55 8.58 99.72 10.29 ;
      RECT 99.49 8.58 99.78 8.81 ;
      RECT 99.49 8.62 100.34 8.78 ;
      RECT 100.175 8.21 100.34 8.78 ;
      RECT 99.49 8.615 99.885 8.78 ;
      RECT 100.11 8.21 100.4 8.44 ;
      RECT 100.11 8.24 100.57 8.41 ;
      RECT 99.12 4.04 99.41 4.27 ;
      RECT 99.12 4.07 99.58 4.24 ;
      RECT 99.185 2.96 99.35 4.27 ;
      RECT 97.7 2.93 97.99 3.16 ;
      RECT 97.7 2.96 99.35 3.13 ;
      RECT 97.76 2.19 97.93 3.16 ;
      RECT 97.7 2.19 97.99 2.42 ;
      RECT 97.7 10.06 97.99 10.29 ;
      RECT 97.76 9.32 97.93 10.29 ;
      RECT 97.76 9.415 99.35 9.585 ;
      RECT 99.18 8.21 99.35 9.585 ;
      RECT 97.7 9.32 97.99 9.55 ;
      RECT 99.12 8.21 99.41 8.44 ;
      RECT 99.12 8.24 99.58 8.41 ;
      RECT 95.685 3.3 96.01 3.625 ;
      RECT 98.13 3.27 98.48 3.62 ;
      RECT 95.685 3.33 98.48 3.5 ;
      RECT 98.155 8.95 98.48 9.275 ;
      RECT 98.13 8.95 98.48 9.18 ;
      RECT 97.96 8.98 98.48 9.15 ;
      RECT 97.355 3.67 97.675 3.99 ;
      RECT 97.33 3.67 97.675 3.9 ;
      RECT 97.04 3.7 97.675 3.87 ;
      RECT 97.355 8.575 97.675 8.9 ;
      RECT 97.33 8.58 97.675 8.81 ;
      RECT 97.155 8.61 97.675 8.78 ;
      RECT 94.685 4.075 95.005 4.335 ;
      RECT 94.405 4.135 95.005 4.275 ;
      RECT 92.305 4.415 92.625 4.675 ;
      RECT 94.275 4.425 94.565 4.655 ;
      RECT 92.305 4.475 94.57 4.615 ;
      RECT 93.665 7.135 93.985 7.395 ;
      RECT 93.665 7.195 94.255 7.335 ;
      RECT 92.985 4.075 93.305 4.335 ;
      RECT 88.245 4.085 88.535 4.315 ;
      RECT 88.245 4.135 93.305 4.275 ;
      RECT 93.075 3.795 93.215 4.335 ;
      RECT 93.075 3.795 93.555 3.935 ;
      RECT 93.415 3.425 93.555 3.935 ;
      RECT 93.335 3.425 93.625 3.655 ;
      RECT 92.985 5.095 93.305 5.355 ;
      RECT 92.315 5.105 92.605 5.335 ;
      RECT 90.105 5.105 90.395 5.335 ;
      RECT 90.105 5.155 93.305 5.295 ;
      RECT 91.285 7.135 91.605 7.395 ;
      RECT 92.995 7.145 93.285 7.375 ;
      RECT 90.615 7.145 90.905 7.375 ;
      RECT 90.615 7.195 91.605 7.335 ;
      RECT 93.075 6.855 93.215 7.375 ;
      RECT 91.375 6.855 91.515 7.395 ;
      RECT 91.375 6.855 93.215 6.995 ;
      RECT 90.275 3.745 90.565 3.975 ;
      RECT 90.355 3.445 90.495 3.975 ;
      RECT 92.675 3.415 92.935 3.705 ;
      RECT 92.645 3.415 92.965 3.675 ;
      RECT 92.545 3.415 92.965 3.655 ;
      RECT 90.355 3.445 92.965 3.585 ;
      RECT 91.625 3.735 91.945 3.995 ;
      RECT 91.625 3.795 92.215 3.935 ;
      RECT 91.625 6.115 91.945 6.375 ;
      RECT 88.915 6.125 89.205 6.355 ;
      RECT 88.915 6.175 91.945 6.315 ;
      RECT 90.945 3.695 91.275 4.025 ;
      RECT 90.945 3.745 91.405 3.975 ;
      RECT 90.945 3.795 91.425 3.935 ;
      RECT 86.935 8.925 87.275 9.205 ;
      RECT 86.905 8.945 87.275 9.175 ;
      RECT 86.735 8.975 87.275 9.145 ;
      RECT 86.475 10.055 86.765 10.285 ;
      RECT 86.535 9.29 86.705 10.285 ;
      RECT 86.435 9.29 86.805 9.66 ;
      RECT 83.9 10.06 84.195 10.29 ;
      RECT 83.96 8.58 84.13 10.29 ;
      RECT 83.96 8.955 84.29 9.28 ;
      RECT 83.9 8.58 84.19 8.81 ;
      RECT 83.495 4.04 83.82 4.27 ;
      RECT 83.495 4.07 83.99 4.24 ;
      RECT 83.495 3.7 83.685 4.27 ;
      RECT 82.91 3.67 83.2 3.9 ;
      RECT 82.91 3.7 83.685 3.87 ;
      RECT 82.97 2.19 83.14 3.9 ;
      RECT 82.91 2.19 83.205 2.42 ;
      RECT 82.91 10.06 83.205 10.29 ;
      RECT 82.97 8.58 83.14 10.29 ;
      RECT 82.91 8.58 83.2 8.81 ;
      RECT 82.91 8.62 83.76 8.78 ;
      RECT 83.595 8.21 83.76 8.78 ;
      RECT 82.91 8.615 83.305 8.78 ;
      RECT 83.53 8.21 83.82 8.44 ;
      RECT 83.53 8.24 83.99 8.41 ;
      RECT 82.54 4.04 82.83 4.27 ;
      RECT 82.54 4.07 83 4.24 ;
      RECT 82.605 2.96 82.77 4.27 ;
      RECT 81.12 2.93 81.41 3.16 ;
      RECT 81.12 2.96 82.77 3.13 ;
      RECT 81.18 2.19 81.35 3.16 ;
      RECT 81.12 2.19 81.41 2.42 ;
      RECT 81.12 10.06 81.41 10.29 ;
      RECT 81.18 9.32 81.35 10.29 ;
      RECT 81.18 9.415 82.77 9.585 ;
      RECT 82.6 8.21 82.77 9.585 ;
      RECT 81.12 9.32 81.41 9.55 ;
      RECT 82.54 8.21 82.83 8.44 ;
      RECT 82.54 8.24 83 8.41 ;
      RECT 79.105 3.3 79.43 3.625 ;
      RECT 81.55 3.27 81.9 3.62 ;
      RECT 79.105 3.33 81.9 3.5 ;
      RECT 81.575 8.95 81.9 9.275 ;
      RECT 81.55 8.95 81.9 9.18 ;
      RECT 81.38 8.98 81.9 9.15 ;
      RECT 80.775 3.67 81.095 3.99 ;
      RECT 80.75 3.67 81.095 3.9 ;
      RECT 80.46 3.7 81.095 3.87 ;
      RECT 80.775 8.575 81.095 8.9 ;
      RECT 80.75 8.58 81.095 8.81 ;
      RECT 80.575 8.61 81.095 8.78 ;
      RECT 78.105 4.075 78.425 4.335 ;
      RECT 77.825 4.135 78.425 4.275 ;
      RECT 75.725 4.415 76.045 4.675 ;
      RECT 77.695 4.425 77.985 4.655 ;
      RECT 75.725 4.475 77.99 4.615 ;
      RECT 77.085 7.135 77.405 7.395 ;
      RECT 77.085 7.195 77.675 7.335 ;
      RECT 76.405 4.075 76.725 4.335 ;
      RECT 71.665 4.085 71.955 4.315 ;
      RECT 71.665 4.135 76.725 4.275 ;
      RECT 76.495 3.795 76.635 4.335 ;
      RECT 76.495 3.795 76.975 3.935 ;
      RECT 76.835 3.425 76.975 3.935 ;
      RECT 76.755 3.425 77.045 3.655 ;
      RECT 76.405 5.095 76.725 5.355 ;
      RECT 75.735 5.105 76.025 5.335 ;
      RECT 73.525 5.105 73.815 5.335 ;
      RECT 73.525 5.155 76.725 5.295 ;
      RECT 74.705 7.135 75.025 7.395 ;
      RECT 76.415 7.145 76.705 7.375 ;
      RECT 74.035 7.145 74.325 7.375 ;
      RECT 74.035 7.195 75.025 7.335 ;
      RECT 76.495 6.855 76.635 7.375 ;
      RECT 74.795 6.855 74.935 7.395 ;
      RECT 74.795 6.855 76.635 6.995 ;
      RECT 73.695 3.745 73.985 3.975 ;
      RECT 73.775 3.445 73.915 3.975 ;
      RECT 76.095 3.415 76.355 3.705 ;
      RECT 76.065 3.415 76.385 3.675 ;
      RECT 75.965 3.415 76.385 3.655 ;
      RECT 73.775 3.445 76.385 3.585 ;
      RECT 75.045 3.735 75.365 3.995 ;
      RECT 75.045 3.795 75.635 3.935 ;
      RECT 75.045 6.115 75.365 6.375 ;
      RECT 72.335 6.125 72.625 6.355 ;
      RECT 72.335 6.175 75.365 6.315 ;
      RECT 74.365 3.695 74.695 4.025 ;
      RECT 74.365 3.745 74.825 3.975 ;
      RECT 74.365 3.795 74.845 3.935 ;
      RECT 70.355 8.925 70.695 9.205 ;
      RECT 70.325 8.945 70.695 9.175 ;
      RECT 70.155 8.975 70.695 9.145 ;
      RECT 69.895 10.055 70.185 10.285 ;
      RECT 69.955 9.29 70.125 10.285 ;
      RECT 69.855 9.29 70.225 9.66 ;
      RECT 67.315 10.055 67.61 10.285 ;
      RECT 67.375 8.575 67.545 10.285 ;
      RECT 67.375 8.95 67.705 9.275 ;
      RECT 67.315 8.575 67.605 8.805 ;
      RECT 66.91 4.035 67.235 4.265 ;
      RECT 66.91 4.065 67.405 4.235 ;
      RECT 66.91 3.695 67.1 4.265 ;
      RECT 66.325 3.665 66.615 3.895 ;
      RECT 66.325 3.695 67.1 3.865 ;
      RECT 66.385 2.185 66.555 3.895 ;
      RECT 66.325 2.185 66.62 2.415 ;
      RECT 66.325 10.055 66.62 10.285 ;
      RECT 66.385 8.575 66.555 10.285 ;
      RECT 66.325 8.575 66.615 8.805 ;
      RECT 66.325 8.615 67.175 8.775 ;
      RECT 67.01 8.205 67.175 8.775 ;
      RECT 66.325 8.61 66.72 8.775 ;
      RECT 66.945 8.205 67.235 8.435 ;
      RECT 66.945 8.235 67.405 8.405 ;
      RECT 65.955 4.035 66.245 4.265 ;
      RECT 65.955 4.065 66.415 4.235 ;
      RECT 66.02 2.955 66.185 4.265 ;
      RECT 64.535 2.925 64.825 3.155 ;
      RECT 64.535 2.955 66.185 3.125 ;
      RECT 64.595 2.185 64.765 3.155 ;
      RECT 64.535 2.185 64.825 2.415 ;
      RECT 64.535 10.055 64.825 10.285 ;
      RECT 64.595 9.315 64.765 10.285 ;
      RECT 64.595 9.41 66.185 9.58 ;
      RECT 66.015 8.205 66.185 9.58 ;
      RECT 64.535 9.315 64.825 9.545 ;
      RECT 65.955 8.205 66.245 8.435 ;
      RECT 65.955 8.235 66.415 8.405 ;
      RECT 62.52 3.295 62.845 3.62 ;
      RECT 64.965 3.265 65.315 3.615 ;
      RECT 62.52 3.325 65.315 3.495 ;
      RECT 64.99 8.945 65.315 9.27 ;
      RECT 64.965 8.945 65.315 9.175 ;
      RECT 64.795 8.975 65.315 9.145 ;
      RECT 64.19 3.665 64.51 3.985 ;
      RECT 64.165 3.665 64.51 3.895 ;
      RECT 63.875 3.695 64.51 3.865 ;
      RECT 64.19 8.57 64.51 8.895 ;
      RECT 64.165 8.575 64.51 8.805 ;
      RECT 63.99 8.605 64.51 8.775 ;
      RECT 61.52 4.07 61.84 4.33 ;
      RECT 61.24 4.13 61.84 4.27 ;
      RECT 59.14 4.41 59.46 4.67 ;
      RECT 61.11 4.42 61.4 4.65 ;
      RECT 59.14 4.47 61.405 4.61 ;
      RECT 60.5 7.13 60.82 7.39 ;
      RECT 60.5 7.19 61.09 7.33 ;
      RECT 59.82 4.07 60.14 4.33 ;
      RECT 55.08 4.08 55.37 4.31 ;
      RECT 55.08 4.13 60.14 4.27 ;
      RECT 59.91 3.79 60.05 4.33 ;
      RECT 59.91 3.79 60.39 3.93 ;
      RECT 60.25 3.42 60.39 3.93 ;
      RECT 60.17 3.42 60.46 3.65 ;
      RECT 59.82 5.09 60.14 5.35 ;
      RECT 59.15 5.1 59.44 5.33 ;
      RECT 56.94 5.1 57.23 5.33 ;
      RECT 56.94 5.15 60.14 5.29 ;
      RECT 58.12 7.13 58.44 7.39 ;
      RECT 59.83 7.14 60.12 7.37 ;
      RECT 57.45 7.14 57.74 7.37 ;
      RECT 57.45 7.19 58.44 7.33 ;
      RECT 59.91 6.85 60.05 7.37 ;
      RECT 58.21 6.85 58.35 7.39 ;
      RECT 58.21 6.85 60.05 6.99 ;
      RECT 57.11 3.74 57.4 3.97 ;
      RECT 57.19 3.44 57.33 3.97 ;
      RECT 59.51 3.41 59.77 3.7 ;
      RECT 59.48 3.41 59.8 3.67 ;
      RECT 59.38 3.41 59.8 3.65 ;
      RECT 57.19 3.44 59.8 3.58 ;
      RECT 58.46 3.73 58.78 3.99 ;
      RECT 58.46 3.79 59.05 3.93 ;
      RECT 58.46 6.11 58.78 6.37 ;
      RECT 55.75 6.12 56.04 6.35 ;
      RECT 55.75 6.17 58.78 6.31 ;
      RECT 57.78 3.69 58.11 4.02 ;
      RECT 57.78 3.74 58.24 3.97 ;
      RECT 57.78 3.79 58.26 3.93 ;
      RECT 53.8 8.885 54.08 9.23 ;
      RECT 53.77 8.885 54.11 9.2 ;
      RECT 53.74 8.885 54.11 9.17 ;
      RECT 53.57 8.97 54.11 9.14 ;
      RECT 53.31 10.05 53.6 10.28 ;
      RECT 53.37 9.285 53.54 10.28 ;
      RECT 53.27 9.285 53.64 9.655 ;
      RECT 50.73 10.05 51.025 10.28 ;
      RECT 50.79 8.57 50.96 10.28 ;
      RECT 50.79 8.945 51.12 9.27 ;
      RECT 50.73 8.57 51.02 8.8 ;
      RECT 50.325 4.03 50.65 4.26 ;
      RECT 50.325 4.06 50.82 4.23 ;
      RECT 50.325 3.69 50.515 4.26 ;
      RECT 49.74 3.66 50.03 3.89 ;
      RECT 49.74 3.69 50.515 3.86 ;
      RECT 49.8 2.18 49.97 3.89 ;
      RECT 49.74 2.18 50.035 2.41 ;
      RECT 49.74 10.05 50.035 10.28 ;
      RECT 49.8 8.57 49.97 10.28 ;
      RECT 49.74 8.57 50.03 8.8 ;
      RECT 49.74 8.61 50.59 8.77 ;
      RECT 50.425 8.2 50.59 8.77 ;
      RECT 49.74 8.605 50.135 8.77 ;
      RECT 50.36 8.2 50.65 8.43 ;
      RECT 50.36 8.23 50.82 8.4 ;
      RECT 49.37 4.03 49.66 4.26 ;
      RECT 49.37 4.06 49.83 4.23 ;
      RECT 49.435 2.95 49.6 4.26 ;
      RECT 47.95 2.92 48.24 3.15 ;
      RECT 47.95 2.95 49.6 3.12 ;
      RECT 48.01 2.18 48.18 3.15 ;
      RECT 47.95 2.18 48.24 2.41 ;
      RECT 47.95 10.05 48.24 10.28 ;
      RECT 48.01 9.31 48.18 10.28 ;
      RECT 48.01 9.405 49.6 9.575 ;
      RECT 49.43 8.2 49.6 9.575 ;
      RECT 47.95 9.31 48.24 9.54 ;
      RECT 49.37 8.2 49.66 8.43 ;
      RECT 49.37 8.23 49.83 8.4 ;
      RECT 45.935 3.29 46.26 3.615 ;
      RECT 48.38 3.26 48.73 3.61 ;
      RECT 45.935 3.32 48.73 3.49 ;
      RECT 48.405 8.94 48.73 9.265 ;
      RECT 48.38 8.94 48.73 9.17 ;
      RECT 48.21 8.97 48.73 9.14 ;
      RECT 47.605 3.66 47.925 3.98 ;
      RECT 47.58 3.66 47.925 3.89 ;
      RECT 47.29 3.69 47.925 3.86 ;
      RECT 47.605 8.565 47.925 8.89 ;
      RECT 47.58 8.57 47.925 8.8 ;
      RECT 47.405 8.6 47.925 8.77 ;
      RECT 44.935 4.065 45.255 4.325 ;
      RECT 44.655 4.125 45.255 4.265 ;
      RECT 42.555 4.405 42.875 4.665 ;
      RECT 44.525 4.415 44.815 4.645 ;
      RECT 42.555 4.465 44.82 4.605 ;
      RECT 43.915 7.125 44.235 7.385 ;
      RECT 43.915 7.185 44.505 7.325 ;
      RECT 43.235 4.065 43.555 4.325 ;
      RECT 38.495 4.075 38.785 4.305 ;
      RECT 38.495 4.125 43.555 4.265 ;
      RECT 43.325 3.785 43.465 4.325 ;
      RECT 43.325 3.785 43.805 3.925 ;
      RECT 43.665 3.415 43.805 3.925 ;
      RECT 43.585 3.415 43.875 3.645 ;
      RECT 43.235 5.085 43.555 5.345 ;
      RECT 42.565 5.095 42.855 5.325 ;
      RECT 40.355 5.095 40.645 5.325 ;
      RECT 40.355 5.145 43.555 5.285 ;
      RECT 41.535 7.125 41.855 7.385 ;
      RECT 43.245 7.135 43.535 7.365 ;
      RECT 40.865 7.135 41.155 7.365 ;
      RECT 40.865 7.185 41.855 7.325 ;
      RECT 43.325 6.845 43.465 7.365 ;
      RECT 41.625 6.845 41.765 7.385 ;
      RECT 41.625 6.845 43.465 6.985 ;
      RECT 40.525 3.735 40.815 3.965 ;
      RECT 40.605 3.435 40.745 3.965 ;
      RECT 42.925 3.405 43.185 3.695 ;
      RECT 42.895 3.405 43.215 3.665 ;
      RECT 42.795 3.405 43.215 3.645 ;
      RECT 40.605 3.435 43.215 3.575 ;
      RECT 41.875 3.725 42.195 3.985 ;
      RECT 41.875 3.785 42.465 3.925 ;
      RECT 41.875 6.105 42.195 6.365 ;
      RECT 39.165 6.115 39.455 6.345 ;
      RECT 39.165 6.165 42.195 6.305 ;
      RECT 41.195 3.685 41.525 4.015 ;
      RECT 41.195 3.735 41.655 3.965 ;
      RECT 41.195 3.785 41.675 3.925 ;
      RECT 37.185 8.915 37.525 9.195 ;
      RECT 37.155 8.935 37.525 9.165 ;
      RECT 36.985 8.965 37.525 9.135 ;
      RECT 36.725 10.045 37.015 10.275 ;
      RECT 36.785 9.28 36.955 10.275 ;
      RECT 36.685 9.28 37.055 9.65 ;
      RECT 34.145 10.05 34.44 10.28 ;
      RECT 34.205 8.57 34.375 10.28 ;
      RECT 34.205 8.945 34.535 9.27 ;
      RECT 34.145 8.57 34.435 8.8 ;
      RECT 33.74 4.03 34.065 4.26 ;
      RECT 33.74 4.06 34.235 4.23 ;
      RECT 33.74 3.69 33.93 4.26 ;
      RECT 33.155 3.66 33.445 3.89 ;
      RECT 33.155 3.69 33.93 3.86 ;
      RECT 33.215 2.18 33.385 3.89 ;
      RECT 33.155 2.18 33.45 2.41 ;
      RECT 33.155 10.05 33.45 10.28 ;
      RECT 33.215 8.57 33.385 10.28 ;
      RECT 33.155 8.57 33.445 8.8 ;
      RECT 33.155 8.61 34.005 8.77 ;
      RECT 33.84 8.2 34.005 8.77 ;
      RECT 33.155 8.605 33.55 8.77 ;
      RECT 33.775 8.2 34.065 8.43 ;
      RECT 33.775 8.23 34.235 8.4 ;
      RECT 32.785 4.03 33.075 4.26 ;
      RECT 32.785 4.06 33.245 4.23 ;
      RECT 32.85 2.95 33.015 4.26 ;
      RECT 31.365 2.92 31.655 3.15 ;
      RECT 31.365 2.95 33.015 3.12 ;
      RECT 31.425 2.18 31.595 3.15 ;
      RECT 31.365 2.18 31.655 2.41 ;
      RECT 31.365 10.05 31.655 10.28 ;
      RECT 31.425 9.31 31.595 10.28 ;
      RECT 31.425 9.405 33.015 9.575 ;
      RECT 32.845 8.2 33.015 9.575 ;
      RECT 31.365 9.31 31.655 9.54 ;
      RECT 32.785 8.2 33.075 8.43 ;
      RECT 32.785 8.23 33.245 8.4 ;
      RECT 29.35 3.29 29.675 3.615 ;
      RECT 31.795 3.26 32.145 3.61 ;
      RECT 29.35 3.32 32.145 3.49 ;
      RECT 31.82 8.94 32.145 9.265 ;
      RECT 31.795 8.94 32.145 9.17 ;
      RECT 31.625 8.97 32.145 9.14 ;
      RECT 31.02 3.66 31.34 3.98 ;
      RECT 30.995 3.66 31.34 3.89 ;
      RECT 30.705 3.69 31.34 3.86 ;
      RECT 31.02 8.565 31.34 8.89 ;
      RECT 30.995 8.57 31.34 8.8 ;
      RECT 30.82 8.6 31.34 8.77 ;
      RECT 28.35 4.065 28.67 4.325 ;
      RECT 28.07 4.125 28.67 4.265 ;
      RECT 25.97 4.405 26.29 4.665 ;
      RECT 27.94 4.415 28.23 4.645 ;
      RECT 25.97 4.465 28.235 4.605 ;
      RECT 27.33 7.125 27.65 7.385 ;
      RECT 27.33 7.185 27.92 7.325 ;
      RECT 26.65 4.065 26.97 4.325 ;
      RECT 21.91 4.075 22.2 4.305 ;
      RECT 21.91 4.125 26.97 4.265 ;
      RECT 26.74 3.785 26.88 4.325 ;
      RECT 26.74 3.785 27.22 3.925 ;
      RECT 27.08 3.415 27.22 3.925 ;
      RECT 27 3.415 27.29 3.645 ;
      RECT 26.65 5.085 26.97 5.345 ;
      RECT 25.98 5.095 26.27 5.325 ;
      RECT 23.77 5.095 24.06 5.325 ;
      RECT 23.77 5.145 26.97 5.285 ;
      RECT 24.95 7.125 25.27 7.385 ;
      RECT 26.66 7.135 26.95 7.365 ;
      RECT 24.28 7.135 24.57 7.365 ;
      RECT 24.28 7.185 25.27 7.325 ;
      RECT 26.74 6.845 26.88 7.365 ;
      RECT 25.04 6.845 25.18 7.385 ;
      RECT 25.04 6.845 26.88 6.985 ;
      RECT 23.94 3.735 24.23 3.965 ;
      RECT 24.02 3.435 24.16 3.965 ;
      RECT 26.34 3.405 26.6 3.695 ;
      RECT 26.31 3.405 26.63 3.665 ;
      RECT 26.21 3.405 26.63 3.645 ;
      RECT 24.02 3.435 26.63 3.575 ;
      RECT 25.29 3.725 25.61 3.985 ;
      RECT 25.29 3.785 25.88 3.925 ;
      RECT 25.29 6.105 25.61 6.365 ;
      RECT 22.58 6.115 22.87 6.345 ;
      RECT 22.58 6.165 25.61 6.305 ;
      RECT 24.61 3.685 24.94 4.015 ;
      RECT 24.61 3.735 25.07 3.965 ;
      RECT 24.61 3.785 25.09 3.925 ;
      RECT 20.6 8.915 20.94 9.195 ;
      RECT 20.57 8.935 20.94 9.165 ;
      RECT 20.4 8.965 20.94 9.135 ;
      RECT 20.14 10.045 20.43 10.275 ;
      RECT 20.2 9.28 20.37 10.275 ;
      RECT 20.1 9.28 20.47 9.65 ;
      RECT 16.91 10.045 17.2 10.275 ;
      RECT 16.97 9.305 17.14 10.275 ;
      RECT 16.89 9.31 17.23 9.59 ;
      RECT 16.91 9.305 17.2 9.59 ;
      RECT 16.505 8.57 16.845 8.85 ;
      RECT 16.365 8.595 16.845 8.765 ;
      RECT 16.54 8.565 16.83 8.85 ;
      RECT 100.455 7.26 100.805 7.55 ;
      RECT 94.355 6.115 95.005 6.375 ;
      RECT 92.305 7.135 92.625 7.395 ;
      RECT 83.875 7.26 84.225 7.55 ;
      RECT 77.775 6.115 78.425 6.375 ;
      RECT 75.725 7.135 76.045 7.395 ;
      RECT 67.29 7.255 67.64 7.545 ;
      RECT 61.19 6.11 61.84 6.37 ;
      RECT 59.14 7.13 59.46 7.39 ;
      RECT 50.705 7.25 51.055 7.54 ;
      RECT 44.605 6.105 45.255 6.365 ;
      RECT 42.555 7.125 42.875 7.385 ;
      RECT 34.12 7.25 34.47 7.54 ;
      RECT 28.02 6.105 28.67 6.365 ;
      RECT 25.97 7.125 26.29 7.385 ;
    LAYER mcon ;
      RECT 100.545 7.315 100.715 7.485 ;
      RECT 100.54 8.61 100.71 8.78 ;
      RECT 100.54 10.09 100.71 10.26 ;
      RECT 100.17 4.07 100.34 4.24 ;
      RECT 100.17 8.24 100.34 8.41 ;
      RECT 99.55 2.22 99.72 2.39 ;
      RECT 99.55 3.7 99.72 3.87 ;
      RECT 99.55 8.61 99.72 8.78 ;
      RECT 99.55 10.09 99.72 10.26 ;
      RECT 99.18 4.07 99.35 4.24 ;
      RECT 99.18 8.24 99.35 8.41 ;
      RECT 98.19 3.33 98.36 3.5 ;
      RECT 98.19 8.98 98.36 9.15 ;
      RECT 97.76 2.22 97.93 2.39 ;
      RECT 97.76 2.96 97.93 3.13 ;
      RECT 97.76 9.35 97.93 9.52 ;
      RECT 97.76 10.09 97.93 10.26 ;
      RECT 97.39 3.7 97.56 3.87 ;
      RECT 97.39 8.61 97.56 8.78 ;
      RECT 94.755 4.115 94.925 4.285 ;
      RECT 94.415 6.155 94.585 6.325 ;
      RECT 94.335 4.455 94.505 4.625 ;
      RECT 93.735 7.175 93.905 7.345 ;
      RECT 93.395 3.455 93.565 3.625 ;
      RECT 93.055 7.175 93.225 7.345 ;
      RECT 92.605 3.445 92.775 3.615 ;
      RECT 92.375 5.135 92.545 5.305 ;
      RECT 92.375 7.175 92.545 7.345 ;
      RECT 91.695 3.775 91.865 3.945 ;
      RECT 91.175 3.775 91.345 3.945 ;
      RECT 90.675 7.175 90.845 7.345 ;
      RECT 90.335 3.775 90.505 3.945 ;
      RECT 90.165 5.135 90.335 5.305 ;
      RECT 88.975 6.155 89.145 6.325 ;
      RECT 88.305 4.115 88.475 4.285 ;
      RECT 86.965 8.975 87.135 9.145 ;
      RECT 86.535 9.345 86.705 9.515 ;
      RECT 86.535 10.085 86.705 10.255 ;
      RECT 83.965 7.315 84.135 7.485 ;
      RECT 83.96 8.61 84.13 8.78 ;
      RECT 83.96 10.09 84.13 10.26 ;
      RECT 83.59 4.07 83.76 4.24 ;
      RECT 83.59 8.24 83.76 8.41 ;
      RECT 82.97 2.22 83.14 2.39 ;
      RECT 82.97 3.7 83.14 3.87 ;
      RECT 82.97 8.61 83.14 8.78 ;
      RECT 82.97 10.09 83.14 10.26 ;
      RECT 82.6 4.07 82.77 4.24 ;
      RECT 82.6 8.24 82.77 8.41 ;
      RECT 81.61 3.33 81.78 3.5 ;
      RECT 81.61 8.98 81.78 9.15 ;
      RECT 81.18 2.22 81.35 2.39 ;
      RECT 81.18 2.96 81.35 3.13 ;
      RECT 81.18 9.35 81.35 9.52 ;
      RECT 81.18 10.09 81.35 10.26 ;
      RECT 80.81 3.7 80.98 3.87 ;
      RECT 80.81 8.61 80.98 8.78 ;
      RECT 78.175 4.115 78.345 4.285 ;
      RECT 77.835 6.155 78.005 6.325 ;
      RECT 77.755 4.455 77.925 4.625 ;
      RECT 77.155 7.175 77.325 7.345 ;
      RECT 76.815 3.455 76.985 3.625 ;
      RECT 76.475 7.175 76.645 7.345 ;
      RECT 76.025 3.445 76.195 3.615 ;
      RECT 75.795 5.135 75.965 5.305 ;
      RECT 75.795 7.175 75.965 7.345 ;
      RECT 75.115 3.775 75.285 3.945 ;
      RECT 74.595 3.775 74.765 3.945 ;
      RECT 74.095 7.175 74.265 7.345 ;
      RECT 73.755 3.775 73.925 3.945 ;
      RECT 73.585 5.135 73.755 5.305 ;
      RECT 72.395 6.155 72.565 6.325 ;
      RECT 71.725 4.115 71.895 4.285 ;
      RECT 70.385 8.975 70.555 9.145 ;
      RECT 69.955 9.345 70.125 9.515 ;
      RECT 69.955 10.085 70.125 10.255 ;
      RECT 67.38 7.31 67.55 7.48 ;
      RECT 67.375 8.605 67.545 8.775 ;
      RECT 67.375 10.085 67.545 10.255 ;
      RECT 67.005 4.065 67.175 4.235 ;
      RECT 67.005 8.235 67.175 8.405 ;
      RECT 66.385 2.215 66.555 2.385 ;
      RECT 66.385 3.695 66.555 3.865 ;
      RECT 66.385 8.605 66.555 8.775 ;
      RECT 66.385 10.085 66.555 10.255 ;
      RECT 66.015 4.065 66.185 4.235 ;
      RECT 66.015 8.235 66.185 8.405 ;
      RECT 65.025 3.325 65.195 3.495 ;
      RECT 65.025 8.975 65.195 9.145 ;
      RECT 64.595 2.215 64.765 2.385 ;
      RECT 64.595 2.955 64.765 3.125 ;
      RECT 64.595 9.345 64.765 9.515 ;
      RECT 64.595 10.085 64.765 10.255 ;
      RECT 64.225 3.695 64.395 3.865 ;
      RECT 64.225 8.605 64.395 8.775 ;
      RECT 61.59 4.11 61.76 4.28 ;
      RECT 61.25 6.15 61.42 6.32 ;
      RECT 61.17 4.45 61.34 4.62 ;
      RECT 60.57 7.17 60.74 7.34 ;
      RECT 60.23 3.45 60.4 3.62 ;
      RECT 59.89 7.17 60.06 7.34 ;
      RECT 59.44 3.44 59.61 3.61 ;
      RECT 59.21 5.13 59.38 5.3 ;
      RECT 59.21 7.17 59.38 7.34 ;
      RECT 58.53 3.77 58.7 3.94 ;
      RECT 58.01 3.77 58.18 3.94 ;
      RECT 57.51 7.17 57.68 7.34 ;
      RECT 57.17 3.77 57.34 3.94 ;
      RECT 57 5.13 57.17 5.3 ;
      RECT 55.81 6.15 55.98 6.32 ;
      RECT 55.14 4.11 55.31 4.28 ;
      RECT 53.8 8.97 53.97 9.14 ;
      RECT 53.37 9.34 53.54 9.51 ;
      RECT 53.37 10.08 53.54 10.25 ;
      RECT 50.795 7.305 50.965 7.475 ;
      RECT 50.79 8.6 50.96 8.77 ;
      RECT 50.79 10.08 50.96 10.25 ;
      RECT 50.42 4.06 50.59 4.23 ;
      RECT 50.42 8.23 50.59 8.4 ;
      RECT 49.8 2.21 49.97 2.38 ;
      RECT 49.8 3.69 49.97 3.86 ;
      RECT 49.8 8.6 49.97 8.77 ;
      RECT 49.8 10.08 49.97 10.25 ;
      RECT 49.43 4.06 49.6 4.23 ;
      RECT 49.43 8.23 49.6 8.4 ;
      RECT 48.44 3.32 48.61 3.49 ;
      RECT 48.44 8.97 48.61 9.14 ;
      RECT 48.01 2.21 48.18 2.38 ;
      RECT 48.01 2.95 48.18 3.12 ;
      RECT 48.01 9.34 48.18 9.51 ;
      RECT 48.01 10.08 48.18 10.25 ;
      RECT 47.64 3.69 47.81 3.86 ;
      RECT 47.64 8.6 47.81 8.77 ;
      RECT 45.005 4.105 45.175 4.275 ;
      RECT 44.665 6.145 44.835 6.315 ;
      RECT 44.585 4.445 44.755 4.615 ;
      RECT 43.985 7.165 44.155 7.335 ;
      RECT 43.645 3.445 43.815 3.615 ;
      RECT 43.305 7.165 43.475 7.335 ;
      RECT 42.855 3.435 43.025 3.605 ;
      RECT 42.625 5.125 42.795 5.295 ;
      RECT 42.625 7.165 42.795 7.335 ;
      RECT 41.945 3.765 42.115 3.935 ;
      RECT 41.425 3.765 41.595 3.935 ;
      RECT 40.925 7.165 41.095 7.335 ;
      RECT 40.585 3.765 40.755 3.935 ;
      RECT 40.415 5.125 40.585 5.295 ;
      RECT 39.225 6.145 39.395 6.315 ;
      RECT 38.555 4.105 38.725 4.275 ;
      RECT 37.215 8.965 37.385 9.135 ;
      RECT 36.785 9.335 36.955 9.505 ;
      RECT 36.785 10.075 36.955 10.245 ;
      RECT 34.21 7.305 34.38 7.475 ;
      RECT 34.205 8.6 34.375 8.77 ;
      RECT 34.205 10.08 34.375 10.25 ;
      RECT 33.835 4.06 34.005 4.23 ;
      RECT 33.835 8.23 34.005 8.4 ;
      RECT 33.215 2.21 33.385 2.38 ;
      RECT 33.215 3.69 33.385 3.86 ;
      RECT 33.215 8.6 33.385 8.77 ;
      RECT 33.215 10.08 33.385 10.25 ;
      RECT 32.845 4.06 33.015 4.23 ;
      RECT 32.845 8.23 33.015 8.4 ;
      RECT 31.855 3.32 32.025 3.49 ;
      RECT 31.855 8.97 32.025 9.14 ;
      RECT 31.425 2.21 31.595 2.38 ;
      RECT 31.425 2.95 31.595 3.12 ;
      RECT 31.425 9.34 31.595 9.51 ;
      RECT 31.425 10.08 31.595 10.25 ;
      RECT 31.055 3.69 31.225 3.86 ;
      RECT 31.055 8.6 31.225 8.77 ;
      RECT 28.42 4.105 28.59 4.275 ;
      RECT 28.08 6.145 28.25 6.315 ;
      RECT 28 4.445 28.17 4.615 ;
      RECT 27.4 7.165 27.57 7.335 ;
      RECT 27.06 3.445 27.23 3.615 ;
      RECT 26.72 7.165 26.89 7.335 ;
      RECT 26.27 3.435 26.44 3.605 ;
      RECT 26.04 5.125 26.21 5.295 ;
      RECT 26.04 7.165 26.21 7.335 ;
      RECT 25.36 3.765 25.53 3.935 ;
      RECT 24.84 3.765 25.01 3.935 ;
      RECT 24.34 7.165 24.51 7.335 ;
      RECT 24 3.765 24.17 3.935 ;
      RECT 23.83 5.125 24 5.295 ;
      RECT 22.64 6.145 22.81 6.315 ;
      RECT 21.97 4.105 22.14 4.275 ;
      RECT 20.63 8.965 20.8 9.135 ;
      RECT 20.2 9.335 20.37 9.505 ;
      RECT 20.2 10.075 20.37 10.245 ;
      RECT 16.97 9.335 17.14 9.505 ;
      RECT 16.97 10.075 17.14 10.245 ;
      RECT 16.6 8.595 16.77 8.765 ;
    LAYER li1 ;
      RECT 100.54 7.31 100.71 8.78 ;
      RECT 100.54 7.31 100.715 8.57 ;
      RECT 100.17 3.05 100.34 4.24 ;
      RECT 100.17 3.05 100.64 3.22 ;
      RECT 100.17 9.26 100.64 9.43 ;
      RECT 100.17 8.24 100.34 9.43 ;
      RECT 99.55 3.91 99.725 5.17 ;
      RECT 99.55 3.7 99.72 5.17 ;
      RECT 99.55 7.31 99.72 8.78 ;
      RECT 99.55 7.31 99.725 8.57 ;
      RECT 99.18 3.05 99.35 4.24 ;
      RECT 99.18 3.05 99.65 3.22 ;
      RECT 99.18 9.26 99.65 9.43 ;
      RECT 99.18 8.24 99.35 9.43 ;
      RECT 98.19 4.03 98.365 5.17 ;
      RECT 98.19 1.88 98.36 5.17 ;
      RECT 98.19 1.88 98.365 2.43 ;
      RECT 98.19 10.05 98.365 10.6 ;
      RECT 98.19 7.31 98.36 10.6 ;
      RECT 98.19 7.31 98.365 8.45 ;
      RECT 97.76 3.91 97.935 5.17 ;
      RECT 97.76 2.96 97.93 5.17 ;
      RECT 97.76 7.31 97.93 9.52 ;
      RECT 97.76 7.31 97.935 8.57 ;
      RECT 97.33 3.94 97.5 5.17 ;
      RECT 97.39 2.16 97.56 4.11 ;
      RECT 97.33 1.88 97.5 2.33 ;
      RECT 97.33 10.15 97.5 10.6 ;
      RECT 97.39 8.37 97.56 10.32 ;
      RECT 97.33 7.31 97.5 8.54 ;
      RECT 96.805 3.91 96.98 5.17 ;
      RECT 96.805 1.88 96.975 5.17 ;
      RECT 96.805 3.38 97.215 3.71 ;
      RECT 96.805 2.54 97.215 2.87 ;
      RECT 96.805 1.88 96.98 2.37 ;
      RECT 96.805 10.11 96.98 10.6 ;
      RECT 96.805 7.31 96.975 10.6 ;
      RECT 96.805 9.61 97.215 9.94 ;
      RECT 96.805 8.77 97.215 9.1 ;
      RECT 96.805 7.31 96.98 8.57 ;
      RECT 92.065 7.945 93.375 8.195 ;
      RECT 92.065 7.625 92.245 8.195 ;
      RECT 91.515 7.625 92.245 7.795 ;
      RECT 91.515 6.785 91.685 7.795 ;
      RECT 92.355 6.825 94.095 7.005 ;
      RECT 93.765 5.985 94.095 7.005 ;
      RECT 91.515 6.785 92.575 6.955 ;
      RECT 93.765 6.155 94.585 6.325 ;
      RECT 92.925 5.985 93.255 6.195 ;
      RECT 92.925 5.985 94.095 6.155 ;
      RECT 93.825 4.505 94.155 5.465 ;
      RECT 93.825 4.505 94.505 4.675 ;
      RECT 94.335 3.275 94.505 4.675 ;
      RECT 94.245 3.275 94.575 3.905 ;
      RECT 93.375 4.775 93.645 5.475 ;
      RECT 93.475 3.275 93.645 5.475 ;
      RECT 93.815 4.085 94.165 4.335 ;
      RECT 93.475 4.115 94.165 4.285 ;
      RECT 93.385 3.275 93.645 3.745 ;
      RECT 92.715 6.415 93.595 6.655 ;
      RECT 93.365 6.325 93.595 6.655 ;
      RECT 92.065 6.415 93.595 6.615 ;
      RECT 92.985 6.365 93.595 6.655 ;
      RECT 92.065 6.285 92.235 6.615 ;
      RECT 92.955 7.175 93.205 7.775 ;
      RECT 92.955 7.175 93.425 7.375 ;
      RECT 92.445 4.395 93.205 4.895 ;
      RECT 91.515 4.205 91.775 4.825 ;
      RECT 92.435 4.335 92.445 4.645 ;
      RECT 92.415 4.395 93.205 4.615 ;
      RECT 93.075 4.005 93.305 4.605 ;
      RECT 92.395 4.325 92.435 4.585 ;
      RECT 92.375 4.395 93.305 4.575 ;
      RECT 92.345 4.395 93.305 4.565 ;
      RECT 92.275 4.395 93.305 4.555 ;
      RECT 92.255 4.395 93.305 4.525 ;
      RECT 92.235 3.305 92.405 4.495 ;
      RECT 92.205 4.395 93.305 4.465 ;
      RECT 92.175 4.395 93.305 4.435 ;
      RECT 92.145 4.385 92.505 4.405 ;
      RECT 92.145 4.375 92.495 4.405 ;
      RECT 91.515 4.205 92.405 4.375 ;
      RECT 91.515 4.365 92.475 4.375 ;
      RECT 91.515 4.355 92.465 4.375 ;
      RECT 91.515 3.305 92.405 3.475 ;
      RECT 92.575 3.805 92.905 4.225 ;
      RECT 92.575 3.315 92.795 4.225 ;
      RECT 92.495 7.175 92.705 7.775 ;
      RECT 92.355 7.175 92.705 7.375 ;
      RECT 91.075 4.775 91.345 5.475 ;
      RECT 91.175 3.275 91.345 5.475 ;
      RECT 91.085 3.275 91.345 3.745 ;
      RECT 89.215 4.435 89.465 4.975 ;
      RECT 90.185 4.435 90.905 4.905 ;
      RECT 89.215 4.435 91.005 4.605 ;
      RECT 90.775 4.005 91.005 4.605 ;
      RECT 89.775 3.315 90.025 4.605 ;
      RECT 89.235 3.315 90.025 3.585 ;
      RECT 90.195 7.125 90.875 7.375 ;
      RECT 90.605 6.765 90.875 7.375 ;
      RECT 90.355 7.545 90.615 8.095 ;
      RECT 90.355 7.545 90.685 8.07 ;
      RECT 89.295 7.545 90.685 7.735 ;
      RECT 89.295 6.705 89.465 7.735 ;
      RECT 89.175 7.125 89.465 7.455 ;
      RECT 89.295 6.705 90.235 6.875 ;
      RECT 89.935 6.155 90.235 6.875 ;
      RECT 90.195 3.735 90.605 4.255 ;
      RECT 90.195 3.315 90.395 4.255 ;
      RECT 88.805 3.495 88.975 5.475 ;
      RECT 88.805 4.005 89.605 4.255 ;
      RECT 88.805 3.495 89.055 4.255 ;
      RECT 88.725 3.495 89.055 3.915 ;
      RECT 88.755 7.905 89.315 8.195 ;
      RECT 88.755 5.985 89.005 8.195 ;
      RECT 88.755 5.985 89.215 6.535 ;
      RECT 86.965 10.045 87.14 10.595 ;
      RECT 86.965 7.305 87.135 10.595 ;
      RECT 86.965 7.305 87.14 8.445 ;
      RECT 86.535 7.305 86.705 9.515 ;
      RECT 86.535 7.305 86.71 8.565 ;
      RECT 85.58 10.105 85.755 10.595 ;
      RECT 85.58 7.305 85.75 10.595 ;
      RECT 85.58 9.605 85.99 9.935 ;
      RECT 85.58 8.765 85.99 9.095 ;
      RECT 85.58 7.305 85.755 8.565 ;
      RECT 83.96 7.31 84.13 8.78 ;
      RECT 83.96 7.31 84.135 8.57 ;
      RECT 83.59 3.05 83.76 4.24 ;
      RECT 83.59 3.05 84.06 3.22 ;
      RECT 83.59 9.26 84.06 9.43 ;
      RECT 83.59 8.24 83.76 9.43 ;
      RECT 82.97 3.91 83.145 5.17 ;
      RECT 82.97 3.7 83.14 5.17 ;
      RECT 82.97 7.31 83.14 8.78 ;
      RECT 82.97 7.31 83.145 8.57 ;
      RECT 82.6 3.05 82.77 4.24 ;
      RECT 82.6 3.05 83.07 3.22 ;
      RECT 82.6 9.26 83.07 9.43 ;
      RECT 82.6 8.24 82.77 9.43 ;
      RECT 81.61 4.03 81.785 5.17 ;
      RECT 81.61 1.88 81.78 5.17 ;
      RECT 81.61 1.88 81.785 2.43 ;
      RECT 81.61 10.05 81.785 10.6 ;
      RECT 81.61 7.31 81.78 10.6 ;
      RECT 81.61 7.31 81.785 8.45 ;
      RECT 81.18 3.91 81.355 5.17 ;
      RECT 81.18 2.96 81.35 5.17 ;
      RECT 81.18 7.31 81.35 9.52 ;
      RECT 81.18 7.31 81.355 8.57 ;
      RECT 80.75 3.94 80.92 5.17 ;
      RECT 80.81 2.16 80.98 4.11 ;
      RECT 80.75 1.88 80.92 2.33 ;
      RECT 80.75 10.15 80.92 10.6 ;
      RECT 80.81 8.37 80.98 10.32 ;
      RECT 80.75 7.31 80.92 8.54 ;
      RECT 80.225 3.91 80.4 5.17 ;
      RECT 80.225 1.88 80.395 5.17 ;
      RECT 80.225 3.38 80.635 3.71 ;
      RECT 80.225 2.54 80.635 2.87 ;
      RECT 80.225 1.88 80.4 2.37 ;
      RECT 80.225 10.11 80.4 10.6 ;
      RECT 80.225 7.31 80.395 10.6 ;
      RECT 80.225 9.61 80.635 9.94 ;
      RECT 80.225 8.77 80.635 9.1 ;
      RECT 80.225 7.31 80.4 8.57 ;
      RECT 75.485 7.945 76.795 8.195 ;
      RECT 75.485 7.625 75.665 8.195 ;
      RECT 74.935 7.625 75.665 7.795 ;
      RECT 74.935 6.785 75.105 7.795 ;
      RECT 75.775 6.825 77.515 7.005 ;
      RECT 77.185 5.985 77.515 7.005 ;
      RECT 74.935 6.785 75.995 6.955 ;
      RECT 77.185 6.155 78.005 6.325 ;
      RECT 76.345 5.985 76.675 6.195 ;
      RECT 76.345 5.985 77.515 6.155 ;
      RECT 77.245 4.505 77.575 5.465 ;
      RECT 77.245 4.505 77.925 4.675 ;
      RECT 77.755 3.275 77.925 4.675 ;
      RECT 77.665 3.275 77.995 3.905 ;
      RECT 76.795 4.775 77.065 5.475 ;
      RECT 76.895 3.275 77.065 5.475 ;
      RECT 77.235 4.085 77.585 4.335 ;
      RECT 76.895 4.115 77.585 4.285 ;
      RECT 76.805 3.275 77.065 3.745 ;
      RECT 76.135 6.415 77.015 6.655 ;
      RECT 76.785 6.325 77.015 6.655 ;
      RECT 75.485 6.415 77.015 6.615 ;
      RECT 76.405 6.365 77.015 6.655 ;
      RECT 75.485 6.285 75.655 6.615 ;
      RECT 76.375 7.175 76.625 7.775 ;
      RECT 76.375 7.175 76.845 7.375 ;
      RECT 75.865 4.395 76.625 4.895 ;
      RECT 74.935 4.205 75.195 4.825 ;
      RECT 75.855 4.335 75.865 4.645 ;
      RECT 75.835 4.395 76.625 4.615 ;
      RECT 76.495 4.005 76.725 4.605 ;
      RECT 75.815 4.325 75.855 4.585 ;
      RECT 75.795 4.395 76.725 4.575 ;
      RECT 75.765 4.395 76.725 4.565 ;
      RECT 75.695 4.395 76.725 4.555 ;
      RECT 75.675 4.395 76.725 4.525 ;
      RECT 75.655 3.305 75.825 4.495 ;
      RECT 75.625 4.395 76.725 4.465 ;
      RECT 75.595 4.395 76.725 4.435 ;
      RECT 75.565 4.385 75.925 4.405 ;
      RECT 75.565 4.375 75.915 4.405 ;
      RECT 74.935 4.205 75.825 4.375 ;
      RECT 74.935 4.365 75.895 4.375 ;
      RECT 74.935 4.355 75.885 4.375 ;
      RECT 74.935 3.305 75.825 3.475 ;
      RECT 75.995 3.805 76.325 4.225 ;
      RECT 75.995 3.315 76.215 4.225 ;
      RECT 75.915 7.175 76.125 7.775 ;
      RECT 75.775 7.175 76.125 7.375 ;
      RECT 74.495 4.775 74.765 5.475 ;
      RECT 74.595 3.275 74.765 5.475 ;
      RECT 74.505 3.275 74.765 3.745 ;
      RECT 72.635 4.435 72.885 4.975 ;
      RECT 73.605 4.435 74.325 4.905 ;
      RECT 72.635 4.435 74.425 4.605 ;
      RECT 74.195 4.005 74.425 4.605 ;
      RECT 73.195 3.315 73.445 4.605 ;
      RECT 72.655 3.315 73.445 3.585 ;
      RECT 73.615 7.125 74.295 7.375 ;
      RECT 74.025 6.765 74.295 7.375 ;
      RECT 73.775 7.545 74.035 8.095 ;
      RECT 73.775 7.545 74.105 8.07 ;
      RECT 72.715 7.545 74.105 7.735 ;
      RECT 72.715 6.705 72.885 7.735 ;
      RECT 72.595 7.125 72.885 7.455 ;
      RECT 72.715 6.705 73.655 6.875 ;
      RECT 73.355 6.155 73.655 6.875 ;
      RECT 73.615 3.735 74.025 4.255 ;
      RECT 73.615 3.315 73.815 4.255 ;
      RECT 72.225 3.495 72.395 5.475 ;
      RECT 72.225 4.005 73.025 4.255 ;
      RECT 72.225 3.495 72.475 4.255 ;
      RECT 72.145 3.495 72.475 3.915 ;
      RECT 72.175 7.905 72.735 8.195 ;
      RECT 72.175 5.985 72.425 8.195 ;
      RECT 72.175 5.985 72.635 6.535 ;
      RECT 70.385 10.045 70.56 10.595 ;
      RECT 70.385 7.305 70.555 10.595 ;
      RECT 70.385 7.305 70.56 8.445 ;
      RECT 69.955 7.305 70.125 9.515 ;
      RECT 69.955 7.305 70.13 8.565 ;
      RECT 69 10.105 69.175 10.595 ;
      RECT 69 7.305 69.17 10.595 ;
      RECT 69 9.605 69.41 9.935 ;
      RECT 69 8.765 69.41 9.095 ;
      RECT 69 7.305 69.175 8.565 ;
      RECT 67.375 7.305 67.545 8.775 ;
      RECT 67.375 7.305 67.55 8.565 ;
      RECT 67.005 3.045 67.175 4.235 ;
      RECT 67.005 3.045 67.475 3.215 ;
      RECT 67.005 9.255 67.475 9.425 ;
      RECT 67.005 8.235 67.175 9.425 ;
      RECT 66.385 3.905 66.56 5.165 ;
      RECT 66.385 3.695 66.555 5.165 ;
      RECT 66.385 7.305 66.555 8.775 ;
      RECT 66.385 7.305 66.56 8.565 ;
      RECT 66.015 3.045 66.185 4.235 ;
      RECT 66.015 3.045 66.485 3.215 ;
      RECT 66.015 9.255 66.485 9.425 ;
      RECT 66.015 8.235 66.185 9.425 ;
      RECT 65.025 4.025 65.2 5.165 ;
      RECT 65.025 1.875 65.195 5.165 ;
      RECT 65.025 1.875 65.2 2.425 ;
      RECT 65.025 10.045 65.2 10.595 ;
      RECT 65.025 7.305 65.195 10.595 ;
      RECT 65.025 7.305 65.2 8.445 ;
      RECT 64.595 3.905 64.77 5.165 ;
      RECT 64.595 2.955 64.765 5.165 ;
      RECT 64.595 7.305 64.765 9.515 ;
      RECT 64.595 7.305 64.77 8.565 ;
      RECT 64.165 3.935 64.335 5.165 ;
      RECT 64.225 2.155 64.395 4.105 ;
      RECT 64.165 1.875 64.335 2.325 ;
      RECT 64.165 10.145 64.335 10.595 ;
      RECT 64.225 8.365 64.395 10.315 ;
      RECT 64.165 7.305 64.335 8.535 ;
      RECT 63.64 3.905 63.815 5.165 ;
      RECT 63.64 1.875 63.81 5.165 ;
      RECT 63.64 3.375 64.05 3.705 ;
      RECT 63.64 2.535 64.05 2.865 ;
      RECT 63.64 1.875 63.815 2.365 ;
      RECT 63.64 10.105 63.815 10.595 ;
      RECT 63.64 7.305 63.81 10.595 ;
      RECT 63.64 9.605 64.05 9.935 ;
      RECT 63.64 8.765 64.05 9.095 ;
      RECT 63.64 7.305 63.815 8.565 ;
      RECT 58.9 7.94 60.21 8.19 ;
      RECT 58.9 7.62 59.08 8.19 ;
      RECT 58.35 7.62 59.08 7.79 ;
      RECT 58.35 6.78 58.52 7.79 ;
      RECT 59.19 6.82 60.93 7 ;
      RECT 60.6 5.98 60.93 7 ;
      RECT 58.35 6.78 59.41 6.95 ;
      RECT 60.6 6.15 61.42 6.32 ;
      RECT 59.76 5.98 60.09 6.19 ;
      RECT 59.76 5.98 60.93 6.15 ;
      RECT 60.66 4.5 60.99 5.46 ;
      RECT 60.66 4.5 61.34 4.67 ;
      RECT 61.17 3.27 61.34 4.67 ;
      RECT 61.08 3.27 61.41 3.9 ;
      RECT 60.21 4.77 60.48 5.47 ;
      RECT 60.31 3.27 60.48 5.47 ;
      RECT 60.65 4.08 61 4.33 ;
      RECT 60.31 4.11 61 4.28 ;
      RECT 60.22 3.27 60.48 3.74 ;
      RECT 59.55 6.41 60.43 6.65 ;
      RECT 60.2 6.32 60.43 6.65 ;
      RECT 58.9 6.41 60.43 6.61 ;
      RECT 59.82 6.36 60.43 6.65 ;
      RECT 58.9 6.28 59.07 6.61 ;
      RECT 59.79 7.17 60.04 7.77 ;
      RECT 59.79 7.17 60.26 7.37 ;
      RECT 59.28 4.39 60.04 4.89 ;
      RECT 58.35 4.2 58.61 4.82 ;
      RECT 59.27 4.33 59.28 4.64 ;
      RECT 59.25 4.39 60.04 4.61 ;
      RECT 59.91 4 60.14 4.6 ;
      RECT 59.23 4.32 59.27 4.58 ;
      RECT 59.21 4.39 60.14 4.57 ;
      RECT 59.18 4.39 60.14 4.56 ;
      RECT 59.11 4.39 60.14 4.55 ;
      RECT 59.09 4.39 60.14 4.52 ;
      RECT 59.07 3.3 59.24 4.49 ;
      RECT 59.04 4.39 60.14 4.46 ;
      RECT 59.01 4.39 60.14 4.43 ;
      RECT 58.98 4.38 59.34 4.4 ;
      RECT 58.98 4.37 59.33 4.4 ;
      RECT 58.35 4.2 59.24 4.37 ;
      RECT 58.35 4.36 59.31 4.37 ;
      RECT 58.35 4.35 59.3 4.37 ;
      RECT 58.35 3.3 59.24 3.47 ;
      RECT 59.41 3.8 59.74 4.22 ;
      RECT 59.41 3.31 59.63 4.22 ;
      RECT 59.33 7.17 59.54 7.77 ;
      RECT 59.19 7.17 59.54 7.37 ;
      RECT 57.91 4.77 58.18 5.47 ;
      RECT 58.01 3.27 58.18 5.47 ;
      RECT 57.92 3.27 58.18 3.74 ;
      RECT 56.05 4.43 56.3 4.97 ;
      RECT 57.02 4.43 57.74 4.9 ;
      RECT 56.05 4.43 57.84 4.6 ;
      RECT 57.61 4 57.84 4.6 ;
      RECT 56.61 3.31 56.86 4.6 ;
      RECT 56.07 3.31 56.86 3.58 ;
      RECT 57.03 7.12 57.71 7.37 ;
      RECT 57.44 6.76 57.71 7.37 ;
      RECT 57.19 7.54 57.45 8.09 ;
      RECT 57.19 7.54 57.52 8.065 ;
      RECT 56.13 7.54 57.52 7.73 ;
      RECT 56.13 6.7 56.3 7.73 ;
      RECT 56.01 7.12 56.3 7.45 ;
      RECT 56.13 6.7 57.07 6.87 ;
      RECT 56.77 6.15 57.07 6.87 ;
      RECT 57.03 3.73 57.44 4.25 ;
      RECT 57.03 3.31 57.23 4.25 ;
      RECT 55.64 3.49 55.81 5.47 ;
      RECT 55.64 4 56.44 4.25 ;
      RECT 55.64 3.49 55.89 4.25 ;
      RECT 55.56 3.49 55.89 3.91 ;
      RECT 55.59 7.9 56.15 8.19 ;
      RECT 55.59 5.98 55.84 8.19 ;
      RECT 55.59 5.98 56.05 6.53 ;
      RECT 53.8 10.04 53.975 10.59 ;
      RECT 53.8 7.3 53.97 10.59 ;
      RECT 53.8 7.3 53.975 8.44 ;
      RECT 53.37 7.3 53.54 9.51 ;
      RECT 53.37 7.3 53.545 8.56 ;
      RECT 52.415 10.1 52.59 10.59 ;
      RECT 52.415 7.3 52.585 10.59 ;
      RECT 52.415 9.6 52.825 9.93 ;
      RECT 52.415 8.76 52.825 9.09 ;
      RECT 52.415 7.3 52.59 8.56 ;
      RECT 50.79 7.3 50.96 8.77 ;
      RECT 50.79 7.3 50.965 8.56 ;
      RECT 50.42 3.04 50.59 4.23 ;
      RECT 50.42 3.04 50.89 3.21 ;
      RECT 50.42 9.25 50.89 9.42 ;
      RECT 50.42 8.23 50.59 9.42 ;
      RECT 49.8 3.9 49.975 5.16 ;
      RECT 49.8 3.69 49.97 5.16 ;
      RECT 49.8 7.3 49.97 8.77 ;
      RECT 49.8 7.3 49.975 8.56 ;
      RECT 49.43 3.04 49.6 4.23 ;
      RECT 49.43 3.04 49.9 3.21 ;
      RECT 49.43 9.25 49.9 9.42 ;
      RECT 49.43 8.23 49.6 9.42 ;
      RECT 48.44 4.02 48.615 5.16 ;
      RECT 48.44 1.87 48.61 5.16 ;
      RECT 48.44 1.87 48.615 2.42 ;
      RECT 48.44 10.04 48.615 10.59 ;
      RECT 48.44 7.3 48.61 10.59 ;
      RECT 48.44 7.3 48.615 8.44 ;
      RECT 48.01 3.9 48.185 5.16 ;
      RECT 48.01 2.95 48.18 5.16 ;
      RECT 48.01 7.3 48.18 9.51 ;
      RECT 48.01 7.3 48.185 8.56 ;
      RECT 47.58 3.93 47.75 5.16 ;
      RECT 47.64 2.15 47.81 4.1 ;
      RECT 47.58 1.87 47.75 2.32 ;
      RECT 47.58 10.14 47.75 10.59 ;
      RECT 47.64 8.36 47.81 10.31 ;
      RECT 47.58 7.3 47.75 8.53 ;
      RECT 47.055 3.9 47.23 5.16 ;
      RECT 47.055 1.87 47.225 5.16 ;
      RECT 47.055 3.37 47.465 3.7 ;
      RECT 47.055 2.53 47.465 2.86 ;
      RECT 47.055 1.87 47.23 2.36 ;
      RECT 47.055 10.1 47.23 10.59 ;
      RECT 47.055 7.3 47.225 10.59 ;
      RECT 47.055 9.6 47.465 9.93 ;
      RECT 47.055 8.76 47.465 9.09 ;
      RECT 47.055 7.3 47.23 8.56 ;
      RECT 42.315 7.935 43.625 8.185 ;
      RECT 42.315 7.615 42.495 8.185 ;
      RECT 41.765 7.615 42.495 7.785 ;
      RECT 41.765 6.775 41.935 7.785 ;
      RECT 42.605 6.815 44.345 6.995 ;
      RECT 44.015 5.975 44.345 6.995 ;
      RECT 41.765 6.775 42.825 6.945 ;
      RECT 44.015 6.145 44.835 6.315 ;
      RECT 43.175 5.975 43.505 6.185 ;
      RECT 43.175 5.975 44.345 6.145 ;
      RECT 44.075 4.495 44.405 5.455 ;
      RECT 44.075 4.495 44.755 4.665 ;
      RECT 44.585 3.265 44.755 4.665 ;
      RECT 44.495 3.265 44.825 3.895 ;
      RECT 43.625 4.765 43.895 5.465 ;
      RECT 43.725 3.265 43.895 5.465 ;
      RECT 44.065 4.075 44.415 4.325 ;
      RECT 43.725 4.105 44.415 4.275 ;
      RECT 43.635 3.265 43.895 3.735 ;
      RECT 42.965 6.405 43.845 6.645 ;
      RECT 43.615 6.315 43.845 6.645 ;
      RECT 42.315 6.405 43.845 6.605 ;
      RECT 43.235 6.355 43.845 6.645 ;
      RECT 42.315 6.275 42.485 6.605 ;
      RECT 43.205 7.165 43.455 7.765 ;
      RECT 43.205 7.165 43.675 7.365 ;
      RECT 42.695 4.385 43.455 4.885 ;
      RECT 41.765 4.195 42.025 4.815 ;
      RECT 42.685 4.325 42.695 4.635 ;
      RECT 42.665 4.385 43.455 4.605 ;
      RECT 43.325 3.995 43.555 4.595 ;
      RECT 42.645 4.315 42.685 4.575 ;
      RECT 42.625 4.385 43.555 4.565 ;
      RECT 42.595 4.385 43.555 4.555 ;
      RECT 42.525 4.385 43.555 4.545 ;
      RECT 42.505 4.385 43.555 4.515 ;
      RECT 42.485 3.295 42.655 4.485 ;
      RECT 42.455 4.385 43.555 4.455 ;
      RECT 42.425 4.385 43.555 4.425 ;
      RECT 42.395 4.375 42.755 4.395 ;
      RECT 42.395 4.365 42.745 4.395 ;
      RECT 41.765 4.195 42.655 4.365 ;
      RECT 41.765 4.355 42.725 4.365 ;
      RECT 41.765 4.345 42.715 4.365 ;
      RECT 41.765 3.295 42.655 3.465 ;
      RECT 42.825 3.795 43.155 4.215 ;
      RECT 42.825 3.305 43.045 4.215 ;
      RECT 42.745 7.165 42.955 7.765 ;
      RECT 42.605 7.165 42.955 7.365 ;
      RECT 41.325 4.765 41.595 5.465 ;
      RECT 41.425 3.265 41.595 5.465 ;
      RECT 41.335 3.265 41.595 3.735 ;
      RECT 39.465 4.425 39.715 4.965 ;
      RECT 40.435 4.425 41.155 4.895 ;
      RECT 39.465 4.425 41.255 4.595 ;
      RECT 41.025 3.995 41.255 4.595 ;
      RECT 40.025 3.305 40.275 4.595 ;
      RECT 39.485 3.305 40.275 3.575 ;
      RECT 40.445 7.115 41.125 7.365 ;
      RECT 40.855 6.755 41.125 7.365 ;
      RECT 40.605 7.535 40.865 8.085 ;
      RECT 40.605 7.535 40.935 8.06 ;
      RECT 39.545 7.535 40.935 7.725 ;
      RECT 39.545 6.695 39.715 7.725 ;
      RECT 39.425 7.115 39.715 7.445 ;
      RECT 39.545 6.695 40.485 6.865 ;
      RECT 40.185 6.145 40.485 6.865 ;
      RECT 40.445 3.725 40.855 4.245 ;
      RECT 40.445 3.305 40.645 4.245 ;
      RECT 39.055 3.485 39.225 5.465 ;
      RECT 39.055 3.995 39.855 4.245 ;
      RECT 39.055 3.485 39.305 4.245 ;
      RECT 38.975 3.485 39.305 3.905 ;
      RECT 39.005 7.895 39.565 8.185 ;
      RECT 39.005 5.975 39.255 8.185 ;
      RECT 39.005 5.975 39.465 6.525 ;
      RECT 37.215 10.035 37.39 10.585 ;
      RECT 37.215 7.295 37.385 10.585 ;
      RECT 37.215 7.295 37.39 8.435 ;
      RECT 36.785 7.295 36.955 9.505 ;
      RECT 36.785 7.295 36.96 8.555 ;
      RECT 35.83 10.095 36.005 10.585 ;
      RECT 35.83 7.295 36 10.585 ;
      RECT 35.83 9.595 36.24 9.925 ;
      RECT 35.83 8.755 36.24 9.085 ;
      RECT 35.83 7.295 36.005 8.555 ;
      RECT 34.205 7.3 34.375 8.77 ;
      RECT 34.205 7.3 34.38 8.56 ;
      RECT 33.835 3.04 34.005 4.23 ;
      RECT 33.835 3.04 34.305 3.21 ;
      RECT 33.835 9.25 34.305 9.42 ;
      RECT 33.835 8.23 34.005 9.42 ;
      RECT 33.215 3.9 33.39 5.16 ;
      RECT 33.215 3.69 33.385 5.16 ;
      RECT 33.215 7.3 33.385 8.77 ;
      RECT 33.215 7.3 33.39 8.56 ;
      RECT 32.845 3.04 33.015 4.23 ;
      RECT 32.845 3.04 33.315 3.21 ;
      RECT 32.845 9.25 33.315 9.42 ;
      RECT 32.845 8.23 33.015 9.42 ;
      RECT 31.855 4.02 32.03 5.16 ;
      RECT 31.855 1.87 32.025 5.16 ;
      RECT 31.855 1.87 32.03 2.42 ;
      RECT 31.855 10.04 32.03 10.59 ;
      RECT 31.855 7.3 32.025 10.59 ;
      RECT 31.855 7.3 32.03 8.44 ;
      RECT 31.425 3.9 31.6 5.16 ;
      RECT 31.425 2.95 31.595 5.16 ;
      RECT 31.425 7.3 31.595 9.51 ;
      RECT 31.425 7.3 31.6 8.56 ;
      RECT 30.995 3.93 31.165 5.16 ;
      RECT 31.055 2.15 31.225 4.1 ;
      RECT 30.995 1.87 31.165 2.32 ;
      RECT 30.995 10.14 31.165 10.59 ;
      RECT 31.055 8.36 31.225 10.31 ;
      RECT 30.995 7.3 31.165 8.53 ;
      RECT 30.47 3.9 30.645 5.16 ;
      RECT 30.47 1.87 30.64 5.16 ;
      RECT 30.47 3.37 30.88 3.7 ;
      RECT 30.47 2.53 30.88 2.86 ;
      RECT 30.47 1.87 30.645 2.36 ;
      RECT 30.47 10.1 30.645 10.59 ;
      RECT 30.47 7.3 30.64 10.59 ;
      RECT 30.47 9.6 30.88 9.93 ;
      RECT 30.47 8.76 30.88 9.09 ;
      RECT 30.47 7.3 30.645 8.56 ;
      RECT 25.73 7.935 27.04 8.185 ;
      RECT 25.73 7.615 25.91 8.185 ;
      RECT 25.18 7.615 25.91 7.785 ;
      RECT 25.18 6.775 25.35 7.785 ;
      RECT 26.02 6.815 27.76 6.995 ;
      RECT 27.43 5.975 27.76 6.995 ;
      RECT 25.18 6.775 26.24 6.945 ;
      RECT 27.43 6.145 28.25 6.315 ;
      RECT 26.59 5.975 26.92 6.185 ;
      RECT 26.59 5.975 27.76 6.145 ;
      RECT 27.49 4.495 27.82 5.455 ;
      RECT 27.49 4.495 28.17 4.665 ;
      RECT 28 3.265 28.17 4.665 ;
      RECT 27.91 3.265 28.24 3.895 ;
      RECT 27.04 4.765 27.31 5.465 ;
      RECT 27.14 3.265 27.31 5.465 ;
      RECT 27.48 4.075 27.83 4.325 ;
      RECT 27.14 4.105 27.83 4.275 ;
      RECT 27.05 3.265 27.31 3.735 ;
      RECT 26.38 6.405 27.26 6.645 ;
      RECT 27.03 6.315 27.26 6.645 ;
      RECT 25.73 6.405 27.26 6.605 ;
      RECT 26.65 6.355 27.26 6.645 ;
      RECT 25.73 6.275 25.9 6.605 ;
      RECT 26.62 7.165 26.87 7.765 ;
      RECT 26.62 7.165 27.09 7.365 ;
      RECT 26.11 4.385 26.87 4.885 ;
      RECT 25.18 4.195 25.44 4.815 ;
      RECT 26.1 4.325 26.11 4.635 ;
      RECT 26.08 4.385 26.87 4.605 ;
      RECT 26.74 3.995 26.97 4.595 ;
      RECT 26.06 4.315 26.1 4.575 ;
      RECT 26.04 4.385 26.97 4.565 ;
      RECT 26.01 4.385 26.97 4.555 ;
      RECT 25.94 4.385 26.97 4.545 ;
      RECT 25.92 4.385 26.97 4.515 ;
      RECT 25.9 3.295 26.07 4.485 ;
      RECT 25.87 4.385 26.97 4.455 ;
      RECT 25.84 4.385 26.97 4.425 ;
      RECT 25.81 4.375 26.17 4.395 ;
      RECT 25.81 4.365 26.16 4.395 ;
      RECT 25.18 4.195 26.07 4.365 ;
      RECT 25.18 4.355 26.14 4.365 ;
      RECT 25.18 4.345 26.13 4.365 ;
      RECT 25.18 3.295 26.07 3.465 ;
      RECT 26.24 3.795 26.57 4.215 ;
      RECT 26.24 3.305 26.46 4.215 ;
      RECT 26.16 7.165 26.37 7.765 ;
      RECT 26.02 7.165 26.37 7.365 ;
      RECT 24.74 4.765 25.01 5.465 ;
      RECT 24.84 3.265 25.01 5.465 ;
      RECT 24.75 3.265 25.01 3.735 ;
      RECT 22.88 4.425 23.13 4.965 ;
      RECT 23.85 4.425 24.57 4.895 ;
      RECT 22.88 4.425 24.67 4.595 ;
      RECT 24.44 3.995 24.67 4.595 ;
      RECT 23.44 3.305 23.69 4.595 ;
      RECT 22.9 3.305 23.69 3.575 ;
      RECT 23.86 7.115 24.54 7.365 ;
      RECT 24.27 6.755 24.54 7.365 ;
      RECT 24.02 7.535 24.28 8.085 ;
      RECT 24.02 7.535 24.35 8.06 ;
      RECT 22.96 7.535 24.35 7.725 ;
      RECT 22.96 6.695 23.13 7.725 ;
      RECT 22.84 7.115 23.13 7.445 ;
      RECT 22.96 6.695 23.9 6.865 ;
      RECT 23.6 6.145 23.9 6.865 ;
      RECT 23.86 3.725 24.27 4.245 ;
      RECT 23.86 3.305 24.06 4.245 ;
      RECT 22.47 3.485 22.64 5.465 ;
      RECT 22.47 3.995 23.27 4.245 ;
      RECT 22.47 3.485 22.72 4.245 ;
      RECT 22.39 3.485 22.72 3.905 ;
      RECT 22.42 7.895 22.98 8.185 ;
      RECT 22.42 5.975 22.67 8.185 ;
      RECT 22.42 5.975 22.88 6.525 ;
      RECT 20.63 10.035 20.805 10.585 ;
      RECT 20.63 7.295 20.8 10.585 ;
      RECT 20.63 7.295 20.805 8.435 ;
      RECT 20.2 7.295 20.37 9.505 ;
      RECT 20.2 7.295 20.375 8.555 ;
      RECT 19.245 10.095 19.42 10.585 ;
      RECT 19.245 7.295 19.415 10.585 ;
      RECT 19.245 9.595 19.655 9.925 ;
      RECT 19.245 8.755 19.655 9.085 ;
      RECT 19.245 7.295 19.42 8.555 ;
      RECT 16.97 7.295 17.14 9.505 ;
      RECT 16.97 7.295 17.145 8.555 ;
      RECT 16.54 10.135 16.71 10.585 ;
      RECT 16.6 8.355 16.77 10.305 ;
      RECT 16.54 7.295 16.71 8.525 ;
      RECT 16.015 10.095 16.19 10.585 ;
      RECT 16.015 7.295 16.185 10.585 ;
      RECT 16.015 9.595 16.425 9.925 ;
      RECT 16.015 8.755 16.425 9.085 ;
      RECT 16.015 7.295 16.19 8.555 ;
      RECT 100.54 10.09 100.715 10.6 ;
      RECT 99.55 1.88 99.725 2.39 ;
      RECT 99.55 10.09 99.725 10.6 ;
      RECT 97.76 1.88 97.935 2.39 ;
      RECT 97.76 10.09 97.935 10.6 ;
      RECT 94.675 4.085 95.025 4.335 ;
      RECT 93.615 7.175 94.065 7.685 ;
      RECT 92.295 5.135 92.775 5.475 ;
      RECT 91.515 3.645 92.065 4.035 ;
      RECT 90.005 5.135 90.475 5.475 ;
      RECT 88.295 4.085 88.635 4.965 ;
      RECT 86.535 10.085 86.71 10.595 ;
      RECT 83.96 10.09 84.135 10.6 ;
      RECT 82.97 1.88 83.145 2.39 ;
      RECT 82.97 10.09 83.145 10.6 ;
      RECT 81.18 1.88 81.355 2.39 ;
      RECT 81.18 10.09 81.355 10.6 ;
      RECT 78.095 4.085 78.445 4.335 ;
      RECT 77.035 7.175 77.485 7.685 ;
      RECT 75.715 5.135 76.195 5.475 ;
      RECT 74.935 3.645 75.485 4.035 ;
      RECT 73.425 5.135 73.895 5.475 ;
      RECT 71.715 4.085 72.055 4.965 ;
      RECT 69.955 10.085 70.13 10.595 ;
      RECT 67.375 10.085 67.55 10.595 ;
      RECT 66.385 1.875 66.56 2.385 ;
      RECT 66.385 10.085 66.56 10.595 ;
      RECT 64.595 1.875 64.77 2.385 ;
      RECT 64.595 10.085 64.77 10.595 ;
      RECT 61.51 4.08 61.86 4.33 ;
      RECT 60.45 7.17 60.9 7.68 ;
      RECT 59.13 5.13 59.61 5.47 ;
      RECT 58.35 3.64 58.9 4.03 ;
      RECT 56.84 5.13 57.31 5.47 ;
      RECT 55.13 4.08 55.47 4.96 ;
      RECT 53.37 10.08 53.545 10.59 ;
      RECT 50.79 10.08 50.965 10.59 ;
      RECT 49.8 1.87 49.975 2.38 ;
      RECT 49.8 10.08 49.975 10.59 ;
      RECT 48.01 1.87 48.185 2.38 ;
      RECT 48.01 10.08 48.185 10.59 ;
      RECT 44.925 4.075 45.275 4.325 ;
      RECT 43.865 7.165 44.315 7.675 ;
      RECT 42.545 5.125 43.025 5.465 ;
      RECT 41.765 3.635 42.315 4.025 ;
      RECT 40.255 5.125 40.725 5.465 ;
      RECT 38.545 4.075 38.885 4.955 ;
      RECT 36.785 10.075 36.96 10.585 ;
      RECT 34.205 10.08 34.38 10.59 ;
      RECT 33.215 1.87 33.39 2.38 ;
      RECT 33.215 10.08 33.39 10.59 ;
      RECT 31.425 1.87 31.6 2.38 ;
      RECT 31.425 10.08 31.6 10.59 ;
      RECT 28.34 4.075 28.69 4.325 ;
      RECT 27.28 7.165 27.73 7.675 ;
      RECT 25.96 5.125 26.44 5.465 ;
      RECT 25.18 3.635 25.73 4.025 ;
      RECT 23.67 5.125 24.14 5.465 ;
      RECT 21.96 4.075 22.3 4.955 ;
      RECT 20.2 10.075 20.375 10.585 ;
      RECT 16.97 10.075 17.145 10.585 ;
  END
END sky130_osu_ring_oscillator_mpr2ca_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2ct_8_b0r1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ct_8_b0r1 ;
  SIZE 103.925 BY 12.46 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 34.395 0 34.775 5.26 ;
      LAYER met2 ;
        RECT 34.395 4.88 34.775 5.26 ;
      LAYER li1 ;
        RECT 34.495 1.865 34.67 2.375 ;
        RECT 34.495 3.895 34.67 5.155 ;
        RECT 34.495 3.685 34.665 5.155 ;
      LAYER met1 ;
        RECT 34.41 4.925 34.76 5.215 ;
        RECT 34.435 2.175 34.73 2.405 ;
        RECT 34.435 3.655 34.725 3.885 ;
        RECT 34.495 2.175 34.665 3.885 ;
      LAYER via1 ;
        RECT 34.51 4.995 34.66 5.145 ;
      LAYER via2 ;
        RECT 34.485 4.97 34.685 5.17 ;
      LAYER mcon ;
        RECT 34.495 3.685 34.665 3.855 ;
        RECT 34.495 2.205 34.665 2.375 ;
        RECT 34.5 4.985 34.67 5.155 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 51.615 0 51.995 5.26 ;
      LAYER met2 ;
        RECT 51.615 4.88 51.995 5.26 ;
      LAYER li1 ;
        RECT 51.715 1.865 51.89 2.375 ;
        RECT 51.715 3.895 51.89 5.155 ;
        RECT 51.715 3.685 51.885 5.155 ;
      LAYER met1 ;
        RECT 51.63 4.925 51.98 5.215 ;
        RECT 51.655 2.175 51.95 2.405 ;
        RECT 51.655 3.655 51.945 3.885 ;
        RECT 51.715 2.175 51.885 3.885 ;
      LAYER via1 ;
        RECT 51.73 4.995 51.88 5.145 ;
      LAYER via2 ;
        RECT 51.705 4.97 51.905 5.17 ;
      LAYER mcon ;
        RECT 51.715 3.685 51.885 3.855 ;
        RECT 51.715 2.205 51.885 2.375 ;
        RECT 51.72 4.985 51.89 5.155 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 68.835 0 69.215 5.26 ;
      LAYER met2 ;
        RECT 68.835 4.88 69.215 5.26 ;
      LAYER li1 ;
        RECT 68.935 1.865 69.11 2.375 ;
        RECT 68.935 3.895 69.11 5.155 ;
        RECT 68.935 3.685 69.105 5.155 ;
      LAYER met1 ;
        RECT 68.85 4.925 69.2 5.215 ;
        RECT 68.875 2.175 69.17 2.405 ;
        RECT 68.875 3.655 69.165 3.885 ;
        RECT 68.935 2.175 69.105 3.885 ;
      LAYER via1 ;
        RECT 68.95 4.995 69.1 5.145 ;
      LAYER via2 ;
        RECT 68.925 4.97 69.125 5.17 ;
      LAYER mcon ;
        RECT 68.935 3.685 69.105 3.855 ;
        RECT 68.935 2.205 69.105 2.375 ;
        RECT 68.94 4.985 69.11 5.155 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 86.055 0 86.435 5.26 ;
      LAYER met2 ;
        RECT 86.055 4.88 86.435 5.26 ;
      LAYER li1 ;
        RECT 86.155 1.865 86.33 2.375 ;
        RECT 86.155 3.895 86.33 5.155 ;
        RECT 86.155 3.685 86.325 5.155 ;
      LAYER met1 ;
        RECT 86.07 4.925 86.42 5.215 ;
        RECT 86.095 2.175 86.39 2.405 ;
        RECT 86.095 3.655 86.385 3.885 ;
        RECT 86.155 2.175 86.325 3.885 ;
      LAYER via1 ;
        RECT 86.17 4.995 86.32 5.145 ;
      LAYER via2 ;
        RECT 86.145 4.97 86.345 5.17 ;
      LAYER mcon ;
        RECT 86.155 3.685 86.325 3.855 ;
        RECT 86.155 2.205 86.325 2.375 ;
        RECT 86.16 4.985 86.33 5.155 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 103.275 0 103.655 5.26 ;
      LAYER met2 ;
        RECT 103.275 4.88 103.655 5.26 ;
      LAYER li1 ;
        RECT 103.375 1.865 103.55 2.375 ;
        RECT 103.375 3.895 103.55 5.155 ;
        RECT 103.375 3.685 103.545 5.155 ;
      LAYER met1 ;
        RECT 103.29 4.925 103.64 5.215 ;
        RECT 103.315 2.175 103.61 2.405 ;
        RECT 103.315 3.655 103.605 3.885 ;
        RECT 103.375 2.175 103.545 3.885 ;
      LAYER via1 ;
        RECT 103.39 4.995 103.54 5.145 ;
      LAYER via2 ;
        RECT 103.365 4.97 103.565 5.17 ;
      LAYER mcon ;
        RECT 103.375 3.685 103.545 3.855 ;
        RECT 103.375 2.205 103.545 2.375 ;
        RECT 103.38 4.985 103.55 5.155 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 30.27 8.14 30.595 8.465 ;
        RECT 30.27 4.79 30.595 5.115 ;
        RECT 20.97 9.32 30.52 9.49 ;
        RECT 30.35 8.14 30.52 9.49 ;
        RECT 30.34 4.79 30.51 8.465 ;
        RECT 20.915 8.145 21.195 8.485 ;
        RECT 20.97 8.145 21.14 9.49 ;
      LAYER li1 ;
        RECT 30.34 8.225 30.52 8.465 ;
        RECT 30.345 8.225 30.515 9.505 ;
        RECT 30.345 2.955 30.515 4.225 ;
        RECT 18.66 8.235 18.83 9.505 ;
      LAYER met1 ;
        RECT 30.285 4.055 30.745 4.225 ;
        RECT 30.27 4.79 30.595 5.115 ;
        RECT 30.285 4.025 30.575 4.255 ;
        RECT 30.35 4.025 30.52 5.115 ;
        RECT 30.27 8.235 30.745 8.405 ;
        RECT 30.27 8.14 30.595 8.465 ;
        RECT 20.885 8.175 21.225 8.455 ;
        RECT 18.6 8.23 21.225 8.4 ;
        RECT 18.6 8.23 19.06 8.405 ;
        RECT 18.6 8.205 18.89 8.435 ;
      LAYER via1 ;
        RECT 20.98 8.24 21.13 8.39 ;
        RECT 30.36 8.225 30.51 8.375 ;
        RECT 30.36 4.875 30.51 5.025 ;
      LAYER mcon ;
        RECT 18.66 8.235 18.83 8.405 ;
        RECT 30.345 8.235 30.515 8.405 ;
        RECT 30.345 4.055 30.515 4.225 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 47.49 8.14 47.815 8.465 ;
        RECT 47.49 4.79 47.815 5.115 ;
        RECT 38.19 9.32 47.74 9.49 ;
        RECT 47.57 8.14 47.74 9.49 ;
        RECT 47.56 4.79 47.73 8.465 ;
        RECT 38.135 8.145 38.415 8.485 ;
        RECT 38.19 8.145 38.36 9.49 ;
      LAYER li1 ;
        RECT 47.56 8.225 47.74 8.465 ;
        RECT 47.565 8.225 47.735 9.505 ;
        RECT 47.565 2.955 47.735 4.225 ;
        RECT 35.88 8.235 36.05 9.505 ;
      LAYER met1 ;
        RECT 47.505 4.055 47.965 4.225 ;
        RECT 47.49 4.79 47.815 5.115 ;
        RECT 47.505 4.025 47.795 4.255 ;
        RECT 47.57 4.025 47.74 5.115 ;
        RECT 47.49 8.235 47.965 8.405 ;
        RECT 47.49 8.14 47.815 8.465 ;
        RECT 38.105 8.175 38.445 8.455 ;
        RECT 35.82 8.23 38.445 8.4 ;
        RECT 35.82 8.23 36.28 8.405 ;
        RECT 35.82 8.205 36.11 8.435 ;
      LAYER via1 ;
        RECT 38.2 8.24 38.35 8.39 ;
        RECT 47.58 8.225 47.73 8.375 ;
        RECT 47.58 4.875 47.73 5.025 ;
      LAYER mcon ;
        RECT 35.88 8.235 36.05 8.405 ;
        RECT 47.565 8.235 47.735 8.405 ;
        RECT 47.565 4.055 47.735 4.225 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 64.71 8.14 65.035 8.465 ;
        RECT 64.71 4.79 65.035 5.115 ;
        RECT 55.41 9.32 64.96 9.49 ;
        RECT 64.79 8.14 64.96 9.49 ;
        RECT 64.78 4.79 64.95 8.465 ;
        RECT 55.355 8.145 55.635 8.485 ;
        RECT 55.41 8.145 55.58 9.49 ;
      LAYER li1 ;
        RECT 64.78 8.225 64.96 8.465 ;
        RECT 64.785 8.225 64.955 9.505 ;
        RECT 64.785 2.955 64.955 4.225 ;
        RECT 53.1 8.235 53.27 9.505 ;
      LAYER met1 ;
        RECT 64.725 4.055 65.185 4.225 ;
        RECT 64.71 4.79 65.035 5.115 ;
        RECT 64.725 4.025 65.015 4.255 ;
        RECT 64.79 4.025 64.96 5.115 ;
        RECT 64.71 8.235 65.185 8.405 ;
        RECT 64.71 8.14 65.035 8.465 ;
        RECT 55.325 8.175 55.665 8.455 ;
        RECT 53.04 8.23 55.665 8.4 ;
        RECT 53.04 8.23 53.5 8.405 ;
        RECT 53.04 8.205 53.33 8.435 ;
      LAYER via1 ;
        RECT 55.42 8.24 55.57 8.39 ;
        RECT 64.8 8.225 64.95 8.375 ;
        RECT 64.8 4.875 64.95 5.025 ;
      LAYER mcon ;
        RECT 53.1 8.235 53.27 8.405 ;
        RECT 64.785 8.235 64.955 8.405 ;
        RECT 64.785 4.055 64.955 4.225 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 81.93 8.14 82.255 8.465 ;
        RECT 81.93 4.79 82.255 5.115 ;
        RECT 72.63 9.32 82.18 9.49 ;
        RECT 82.01 8.14 82.18 9.49 ;
        RECT 82 4.79 82.17 8.465 ;
        RECT 72.575 8.145 72.855 8.485 ;
        RECT 72.63 8.145 72.8 9.49 ;
      LAYER li1 ;
        RECT 82 8.225 82.18 8.465 ;
        RECT 82.005 8.225 82.175 9.505 ;
        RECT 82.005 2.955 82.175 4.225 ;
        RECT 70.32 8.235 70.49 9.505 ;
      LAYER met1 ;
        RECT 81.945 4.055 82.405 4.225 ;
        RECT 81.93 4.79 82.255 5.115 ;
        RECT 81.945 4.025 82.235 4.255 ;
        RECT 82.01 4.025 82.18 5.115 ;
        RECT 81.93 8.235 82.405 8.405 ;
        RECT 81.93 8.14 82.255 8.465 ;
        RECT 72.545 8.175 72.885 8.455 ;
        RECT 70.26 8.23 72.885 8.4 ;
        RECT 70.26 8.23 70.72 8.405 ;
        RECT 70.26 8.205 70.55 8.435 ;
      LAYER via1 ;
        RECT 72.64 8.24 72.79 8.39 ;
        RECT 82.02 8.225 82.17 8.375 ;
        RECT 82.02 4.875 82.17 5.025 ;
      LAYER mcon ;
        RECT 70.32 8.235 70.49 8.405 ;
        RECT 82.005 8.235 82.175 8.405 ;
        RECT 82.005 4.055 82.175 4.225 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 99.15 8.14 99.475 8.465 ;
        RECT 99.15 4.79 99.475 5.115 ;
        RECT 89.85 9.32 99.4 9.49 ;
        RECT 99.23 8.14 99.4 9.49 ;
        RECT 99.22 4.79 99.39 8.465 ;
        RECT 89.795 8.145 90.075 8.485 ;
        RECT 89.85 8.145 90.02 9.49 ;
      LAYER li1 ;
        RECT 99.22 8.225 99.4 8.465 ;
        RECT 99.225 8.225 99.395 9.505 ;
        RECT 99.225 2.955 99.395 4.225 ;
        RECT 87.54 8.235 87.71 9.505 ;
      LAYER met1 ;
        RECT 99.165 4.055 99.625 4.225 ;
        RECT 99.15 4.79 99.475 5.115 ;
        RECT 99.165 4.025 99.455 4.255 ;
        RECT 99.23 4.025 99.4 5.115 ;
        RECT 99.15 8.235 99.625 8.405 ;
        RECT 99.15 8.14 99.475 8.465 ;
        RECT 89.765 8.175 90.105 8.455 ;
        RECT 87.48 8.23 90.105 8.4 ;
        RECT 87.48 8.23 87.94 8.405 ;
        RECT 87.48 8.205 87.77 8.435 ;
      LAYER via1 ;
        RECT 89.86 8.24 90.01 8.39 ;
        RECT 99.24 8.225 99.39 8.375 ;
        RECT 99.24 4.875 99.39 5.025 ;
      LAYER mcon ;
        RECT 87.54 8.235 87.71 8.405 ;
        RECT 99.225 8.235 99.395 8.405 ;
        RECT 99.225 4.055 99.395 4.225 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 15.25 8.235 15.42 9.505 ;
      LAYER met1 ;
        RECT 15.19 8.235 15.65 8.405 ;
        RECT 15.195 8.2 15.485 8.43 ;
        RECT 15.19 8.205 15.48 8.435 ;
      LAYER mcon ;
        RECT 15.25 8.235 15.42 8.405 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 97.84 5.64 103.925 7.03 ;
        RECT 97.935 5.43 103.925 7.03 ;
        RECT 99.045 5.43 103.77 7.035 ;
        RECT 99.045 5.425 103.765 7.035 ;
        RECT 102.95 5.425 103.12 7.765 ;
        RECT 102.945 4.695 103.115 7.035 ;
        RECT 101.96 4.695 102.13 7.765 ;
        RECT 99.215 4.695 99.385 7.765 ;
        RECT 0.015 5.64 103.925 5.81 ;
        RECT 97.025 5.64 97.305 6.95 ;
        RECT 96.625 4.79 96.795 5.81 ;
        RECT 96.095 5.64 96.355 6.95 ;
        RECT 95.785 5.13 95.955 5.81 ;
        RECT 95.645 5.64 95.925 6.95 ;
        RECT 94.715 5.64 94.975 6.95 ;
        RECT 94.285 5.64 94.545 6.95 ;
        RECT 94.205 4.5 94.535 5.81 ;
        RECT 93.335 5.64 93.615 6.95 ;
        RECT 91.965 4.5 92.295 5.81 ;
        RECT 91.985 4.5 92.245 6.95 ;
        RECT 91.515 4.5 91.745 5.81 ;
        RECT 91.035 5.64 91.315 6.95 ;
        RECT 80.715 5.43 90.845 5.81 ;
        RECT 90.635 4.5 90.845 5.81 ;
        RECT 81.825 5.425 90.845 5.81 ;
        RECT 80.62 5.64 90.505 7 ;
        RECT 87.36 5.425 90.375 7.03 ;
        RECT 87.36 5.425 90.11 7.035 ;
        RECT 87.53 5.425 87.7 7.765 ;
        RECT 80.62 5.64 90.375 7.025 ;
        RECT 80.62 5.64 86.705 7.03 ;
        RECT 81.825 5.425 86.55 7.035 ;
        RECT 85.73 5.425 85.9 7.765 ;
        RECT 85.725 4.695 85.895 7.035 ;
        RECT 84.74 4.695 84.91 7.765 ;
        RECT 81.995 4.695 82.165 7.765 ;
        RECT 79.805 5.64 80.085 6.95 ;
        RECT 79.405 4.79 79.575 5.81 ;
        RECT 78.875 5.64 79.135 6.95 ;
        RECT 78.565 5.13 78.735 5.81 ;
        RECT 78.425 5.64 78.705 6.95 ;
        RECT 77.495 5.64 77.755 6.95 ;
        RECT 77.065 5.64 77.325 6.95 ;
        RECT 76.985 4.5 77.315 5.81 ;
        RECT 76.115 5.64 76.395 6.95 ;
        RECT 74.745 4.5 75.075 5.81 ;
        RECT 74.765 4.5 75.025 6.95 ;
        RECT 74.295 4.5 74.525 5.81 ;
        RECT 73.815 5.64 74.095 6.95 ;
        RECT 63.495 5.43 73.625 5.81 ;
        RECT 73.415 4.5 73.625 5.81 ;
        RECT 64.605 5.425 73.625 5.81 ;
        RECT 63.4 5.64 73.285 7 ;
        RECT 70.14 5.425 73.155 7.03 ;
        RECT 70.14 5.425 72.89 7.035 ;
        RECT 70.31 5.425 70.48 7.765 ;
        RECT 63.4 5.64 73.155 7.025 ;
        RECT 63.4 5.64 69.485 7.03 ;
        RECT 64.605 5.425 69.33 7.035 ;
        RECT 68.51 5.425 68.68 7.765 ;
        RECT 68.505 4.695 68.675 7.035 ;
        RECT 67.52 4.695 67.69 7.765 ;
        RECT 64.775 4.695 64.945 7.765 ;
        RECT 62.585 5.64 62.865 6.95 ;
        RECT 62.185 4.79 62.355 5.81 ;
        RECT 61.655 5.64 61.915 6.95 ;
        RECT 61.345 5.13 61.515 5.81 ;
        RECT 61.205 5.64 61.485 6.95 ;
        RECT 60.275 5.64 60.535 6.95 ;
        RECT 59.845 5.64 60.105 6.95 ;
        RECT 59.765 4.5 60.095 5.81 ;
        RECT 58.895 5.64 59.175 6.95 ;
        RECT 57.525 4.5 57.855 5.81 ;
        RECT 57.545 4.5 57.805 6.95 ;
        RECT 57.075 4.5 57.305 5.81 ;
        RECT 56.595 5.64 56.875 6.95 ;
        RECT 46.275 5.43 56.405 5.81 ;
        RECT 56.195 4.5 56.405 5.81 ;
        RECT 47.385 5.425 56.405 5.81 ;
        RECT 46.18 5.64 56.065 7 ;
        RECT 46.18 5.64 55.935 7.03 ;
        RECT 52.92 5.425 55.67 7.035 ;
        RECT 53.09 5.425 53.26 7.765 ;
        RECT 47.385 5.425 52.11 7.035 ;
        RECT 51.29 5.425 51.46 7.765 ;
        RECT 51.285 4.695 51.455 7.035 ;
        RECT 50.3 4.695 50.47 7.765 ;
        RECT 47.555 4.695 47.725 7.765 ;
        RECT 45.365 5.64 45.645 6.95 ;
        RECT 44.965 4.79 45.135 5.81 ;
        RECT 44.435 5.64 44.695 6.95 ;
        RECT 44.125 5.13 44.295 5.81 ;
        RECT 43.985 5.64 44.265 6.95 ;
        RECT 43.055 5.64 43.315 6.95 ;
        RECT 42.625 5.64 42.885 6.95 ;
        RECT 42.545 4.5 42.875 5.81 ;
        RECT 41.675 5.64 41.955 6.95 ;
        RECT 40.305 4.5 40.635 5.81 ;
        RECT 40.325 4.5 40.585 6.95 ;
        RECT 39.855 4.5 40.085 5.81 ;
        RECT 39.375 5.64 39.655 6.95 ;
        RECT 29.055 5.43 39.185 5.81 ;
        RECT 38.975 4.5 39.185 5.81 ;
        RECT 30.165 5.425 39.185 5.81 ;
        RECT 28.96 5.64 38.845 7 ;
        RECT 35.7 5.425 38.715 7.03 ;
        RECT 35.7 5.425 38.45 7.035 ;
        RECT 35.87 5.425 36.04 7.765 ;
        RECT 28.96 5.64 38.715 7.025 ;
        RECT 28.96 5.64 35.045 7.03 ;
        RECT 30.165 5.425 34.89 7.035 ;
        RECT 34.07 5.425 34.24 7.765 ;
        RECT 34.065 4.695 34.235 7.035 ;
        RECT 33.08 4.695 33.25 7.765 ;
        RECT 30.335 4.695 30.505 7.765 ;
        RECT 28.145 5.64 28.425 6.95 ;
        RECT 27.745 4.79 27.915 5.81 ;
        RECT 27.215 5.64 27.475 6.95 ;
        RECT 26.905 5.13 27.075 5.81 ;
        RECT 26.765 5.64 27.045 6.95 ;
        RECT 25.835 5.64 26.095 6.95 ;
        RECT 25.405 5.64 25.665 6.95 ;
        RECT 25.325 4.5 25.655 5.81 ;
        RECT 24.455 5.64 24.735 6.95 ;
        RECT 23.085 4.5 23.415 5.81 ;
        RECT 23.105 4.5 23.365 6.95 ;
        RECT 22.635 4.5 22.865 5.81 ;
        RECT 22.155 5.64 22.435 6.95 ;
        RECT 0.015 5.425 21.965 5.81 ;
        RECT 21.755 4.5 21.965 5.81 ;
        RECT 0.015 5.425 21.625 7 ;
        RECT 0.015 5.425 21.5 7.025 ;
        RECT 18.48 5.425 21.495 7.03 ;
        RECT 18.48 5.425 21.23 7.035 ;
        RECT 18.65 5.425 18.82 7.765 ;
        RECT 15.07 5.425 17.82 7.035 ;
        RECT 17.055 10.045 17.23 10.595 ;
        RECT 17.055 7.305 17.23 8.445 ;
        RECT 17.055 5.425 17.225 10.595 ;
        RECT 15.24 5.425 15.41 7.765 ;
      LAYER met1 ;
        RECT 97.84 5.485 103.925 7.03 ;
        RECT 97.935 5.43 103.925 7.03 ;
        RECT 99.045 5.43 103.77 7.035 ;
        RECT 99.045 5.425 103.765 7.035 ;
        RECT 0.015 5.485 103.925 5.965 ;
        RECT 80.715 5.43 90.665 5.965 ;
        RECT 81.825 5.425 90.665 5.965 ;
        RECT 80.62 5.485 90.505 7 ;
        RECT 80.62 5.485 90.375 7.03 ;
        RECT 87.36 5.425 90.11 7.035 ;
        RECT 81.825 5.425 86.55 7.035 ;
        RECT 63.495 5.43 73.445 5.965 ;
        RECT 64.605 5.425 73.445 5.965 ;
        RECT 63.4 5.485 73.285 7 ;
        RECT 63.4 5.485 73.155 7.03 ;
        RECT 70.14 5.425 72.89 7.035 ;
        RECT 64.605 5.425 69.33 7.035 ;
        RECT 46.275 5.43 56.225 5.965 ;
        RECT 47.385 5.425 56.225 5.965 ;
        RECT 46.18 5.485 56.065 7 ;
        RECT 46.18 5.485 55.935 7.03 ;
        RECT 52.92 5.425 55.67 7.035 ;
        RECT 47.385 5.425 52.11 7.035 ;
        RECT 29.055 5.43 39.005 5.965 ;
        RECT 30.165 5.425 39.005 5.965 ;
        RECT 28.96 5.485 38.845 7 ;
        RECT 28.96 5.485 38.715 7.03 ;
        RECT 35.7 5.425 38.45 7.035 ;
        RECT 30.165 5.425 34.89 7.035 ;
        RECT 0.015 5.425 21.785 5.965 ;
        RECT 0.015 5.425 21.625 7 ;
        RECT 0.015 5.425 21.5 7.025 ;
        RECT 18.48 5.425 21.495 7.03 ;
        RECT 18.48 5.425 21.23 7.035 ;
        RECT 15.07 5.425 17.82 7.035 ;
        RECT 16.995 8.945 17.285 9.175 ;
        RECT 16.825 8.975 17.285 9.145 ;
      LAYER mcon ;
        RECT 17.055 8.975 17.225 9.145 ;
        RECT 17.36 6.835 17.53 7.005 ;
        RECT 20.77 6.835 20.94 7.005 ;
        RECT 21.755 5.64 21.925 5.81 ;
        RECT 22.215 5.64 22.385 5.81 ;
        RECT 22.675 5.64 22.845 5.81 ;
        RECT 23.135 5.64 23.305 5.81 ;
        RECT 23.595 5.64 23.765 5.81 ;
        RECT 24.055 5.64 24.225 5.81 ;
        RECT 24.515 5.64 24.685 5.81 ;
        RECT 24.975 5.64 25.145 5.81 ;
        RECT 25.435 5.64 25.605 5.81 ;
        RECT 25.895 5.64 26.065 5.81 ;
        RECT 26.355 5.64 26.525 5.81 ;
        RECT 26.815 5.64 26.985 5.81 ;
        RECT 27.275 5.64 27.445 5.81 ;
        RECT 27.735 5.64 27.905 5.81 ;
        RECT 28.195 5.64 28.365 5.81 ;
        RECT 28.655 5.64 28.825 5.81 ;
        RECT 32.455 6.835 32.625 7.005 ;
        RECT 32.455 5.455 32.625 5.625 ;
        RECT 33.16 6.835 33.33 7.005 ;
        RECT 33.16 5.455 33.33 5.625 ;
        RECT 34.145 5.455 34.315 5.625 ;
        RECT 34.15 6.835 34.32 7.005 ;
        RECT 37.99 6.835 38.16 7.005 ;
        RECT 38.975 5.64 39.145 5.81 ;
        RECT 39.435 5.64 39.605 5.81 ;
        RECT 39.895 5.64 40.065 5.81 ;
        RECT 40.355 5.64 40.525 5.81 ;
        RECT 40.815 5.64 40.985 5.81 ;
        RECT 41.275 5.64 41.445 5.81 ;
        RECT 41.735 5.64 41.905 5.81 ;
        RECT 42.195 5.64 42.365 5.81 ;
        RECT 42.655 5.64 42.825 5.81 ;
        RECT 43.115 5.64 43.285 5.81 ;
        RECT 43.575 5.64 43.745 5.81 ;
        RECT 44.035 5.64 44.205 5.81 ;
        RECT 44.495 5.64 44.665 5.81 ;
        RECT 44.955 5.64 45.125 5.81 ;
        RECT 45.415 5.64 45.585 5.81 ;
        RECT 45.875 5.64 46.045 5.81 ;
        RECT 49.675 6.835 49.845 7.005 ;
        RECT 49.675 5.455 49.845 5.625 ;
        RECT 50.38 6.835 50.55 7.005 ;
        RECT 50.38 5.455 50.55 5.625 ;
        RECT 51.365 5.455 51.535 5.625 ;
        RECT 51.37 6.835 51.54 7.005 ;
        RECT 55.21 6.835 55.38 7.005 ;
        RECT 56.195 5.64 56.365 5.81 ;
        RECT 56.655 5.64 56.825 5.81 ;
        RECT 57.115 5.64 57.285 5.81 ;
        RECT 57.575 5.64 57.745 5.81 ;
        RECT 58.035 5.64 58.205 5.81 ;
        RECT 58.495 5.64 58.665 5.81 ;
        RECT 58.955 5.64 59.125 5.81 ;
        RECT 59.415 5.64 59.585 5.81 ;
        RECT 59.875 5.64 60.045 5.81 ;
        RECT 60.335 5.64 60.505 5.81 ;
        RECT 60.795 5.64 60.965 5.81 ;
        RECT 61.255 5.64 61.425 5.81 ;
        RECT 61.715 5.64 61.885 5.81 ;
        RECT 62.175 5.64 62.345 5.81 ;
        RECT 62.635 5.64 62.805 5.81 ;
        RECT 63.095 5.64 63.265 5.81 ;
        RECT 66.895 6.835 67.065 7.005 ;
        RECT 66.895 5.455 67.065 5.625 ;
        RECT 67.6 6.835 67.77 7.005 ;
        RECT 67.6 5.455 67.77 5.625 ;
        RECT 68.585 5.455 68.755 5.625 ;
        RECT 68.59 6.835 68.76 7.005 ;
        RECT 72.43 6.835 72.6 7.005 ;
        RECT 73.415 5.64 73.585 5.81 ;
        RECT 73.875 5.64 74.045 5.81 ;
        RECT 74.335 5.64 74.505 5.81 ;
        RECT 74.795 5.64 74.965 5.81 ;
        RECT 75.255 5.64 75.425 5.81 ;
        RECT 75.715 5.64 75.885 5.81 ;
        RECT 76.175 5.64 76.345 5.81 ;
        RECT 76.635 5.64 76.805 5.81 ;
        RECT 77.095 5.64 77.265 5.81 ;
        RECT 77.555 5.64 77.725 5.81 ;
        RECT 78.015 5.64 78.185 5.81 ;
        RECT 78.475 5.64 78.645 5.81 ;
        RECT 78.935 5.64 79.105 5.81 ;
        RECT 79.395 5.64 79.565 5.81 ;
        RECT 79.855 5.64 80.025 5.81 ;
        RECT 80.315 5.64 80.485 5.81 ;
        RECT 84.115 6.835 84.285 7.005 ;
        RECT 84.115 5.455 84.285 5.625 ;
        RECT 84.82 6.835 84.99 7.005 ;
        RECT 84.82 5.455 84.99 5.625 ;
        RECT 85.805 5.455 85.975 5.625 ;
        RECT 85.81 6.835 85.98 7.005 ;
        RECT 89.65 6.835 89.82 7.005 ;
        RECT 90.635 5.64 90.805 5.81 ;
        RECT 91.095 5.64 91.265 5.81 ;
        RECT 91.555 5.64 91.725 5.81 ;
        RECT 92.015 5.64 92.185 5.81 ;
        RECT 92.475 5.64 92.645 5.81 ;
        RECT 92.935 5.64 93.105 5.81 ;
        RECT 93.395 5.64 93.565 5.81 ;
        RECT 93.855 5.64 94.025 5.81 ;
        RECT 94.315 5.64 94.485 5.81 ;
        RECT 94.775 5.64 94.945 5.81 ;
        RECT 95.235 5.64 95.405 5.81 ;
        RECT 95.695 5.64 95.865 5.81 ;
        RECT 96.155 5.64 96.325 5.81 ;
        RECT 96.615 5.64 96.785 5.81 ;
        RECT 97.075 5.64 97.245 5.81 ;
        RECT 97.535 5.64 97.705 5.81 ;
        RECT 101.335 6.835 101.505 7.005 ;
        RECT 101.335 5.455 101.505 5.625 ;
        RECT 102.04 6.835 102.21 7.005 ;
        RECT 102.04 5.455 102.21 5.625 ;
        RECT 103.025 5.455 103.195 5.625 ;
        RECT 103.03 6.835 103.2 7.005 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 92.875 7.085 93.205 7.415 ;
        RECT 92.405 7.1 93.205 7.4 ;
        RECT 75.655 7.085 75.985 7.415 ;
        RECT 75.185 7.1 75.985 7.4 ;
        RECT 58.435 7.085 58.765 7.415 ;
        RECT 57.965 7.1 58.765 7.4 ;
        RECT 41.215 7.085 41.545 7.415 ;
        RECT 40.745 7.1 41.545 7.4 ;
        RECT 23.995 7.085 24.325 7.415 ;
        RECT 23.525 7.1 24.325 7.4 ;
      LAYER met2 ;
        RECT 92.9 7.065 93.18 7.435 ;
        RECT 75.68 7.065 75.96 7.435 ;
        RECT 58.46 7.065 58.74 7.435 ;
        RECT 41.24 7.065 41.52 7.435 ;
        RECT 24.02 7.065 24.3 7.435 ;
      LAYER li1 ;
        RECT 0.015 0 103.925 1.6 ;
        RECT 102.945 0 103.115 2.225 ;
        RECT 101.96 0 102.13 2.225 ;
        RECT 99.215 0 99.385 2.225 ;
        RECT 90.485 0 98.145 3.09 ;
        RECT 97.385 0 97.715 3.48 ;
        RECT 96.545 0 96.875 3.48 ;
        RECT 94.715 0 95.005 3.925 ;
        RECT 94.265 0 94.535 3.9 ;
        RECT 93.355 0 93.595 3.9 ;
        RECT 92.905 0 93.145 3.9 ;
        RECT 91.965 0 92.235 3.9 ;
        RECT 91.515 0 91.745 3.91 ;
        RECT 90.635 0 90.845 3.91 ;
        RECT 85.725 0 85.895 2.225 ;
        RECT 84.74 0 84.91 2.225 ;
        RECT 81.995 0 82.165 2.225 ;
        RECT 73.265 0 80.925 3.09 ;
        RECT 80.165 0 80.495 3.48 ;
        RECT 79.325 0 79.655 3.48 ;
        RECT 77.495 0 77.785 3.925 ;
        RECT 77.045 0 77.315 3.9 ;
        RECT 76.135 0 76.375 3.9 ;
        RECT 75.685 0 75.925 3.9 ;
        RECT 74.745 0 75.015 3.9 ;
        RECT 74.295 0 74.525 3.91 ;
        RECT 73.415 0 73.625 3.91 ;
        RECT 68.505 0 68.675 2.225 ;
        RECT 67.52 0 67.69 2.225 ;
        RECT 64.775 0 64.945 2.225 ;
        RECT 56.045 0 63.705 3.09 ;
        RECT 62.945 0 63.275 3.48 ;
        RECT 62.105 0 62.435 3.48 ;
        RECT 60.275 0 60.565 3.925 ;
        RECT 59.825 0 60.095 3.9 ;
        RECT 58.915 0 59.155 3.9 ;
        RECT 58.465 0 58.705 3.9 ;
        RECT 57.525 0 57.795 3.9 ;
        RECT 57.075 0 57.305 3.91 ;
        RECT 56.195 0 56.405 3.91 ;
        RECT 51.285 0 51.455 2.225 ;
        RECT 50.3 0 50.47 2.225 ;
        RECT 47.555 0 47.725 2.225 ;
        RECT 38.825 0 46.485 3.09 ;
        RECT 45.725 0 46.055 3.48 ;
        RECT 44.885 0 45.215 3.48 ;
        RECT 43.055 0 43.345 3.925 ;
        RECT 42.605 0 42.875 3.9 ;
        RECT 41.695 0 41.935 3.9 ;
        RECT 41.245 0 41.485 3.9 ;
        RECT 40.305 0 40.575 3.9 ;
        RECT 39.855 0 40.085 3.91 ;
        RECT 38.975 0 39.185 3.91 ;
        RECT 34.065 0 34.235 2.225 ;
        RECT 33.08 0 33.25 2.225 ;
        RECT 30.335 0 30.505 2.225 ;
        RECT 21.605 0 29.265 3.09 ;
        RECT 28.505 0 28.835 3.48 ;
        RECT 27.665 0 27.995 3.48 ;
        RECT 25.835 0 26.125 3.925 ;
        RECT 25.385 0 25.655 3.9 ;
        RECT 24.475 0 24.715 3.9 ;
        RECT 24.025 0 24.265 3.9 ;
        RECT 23.085 0 23.355 3.9 ;
        RECT 22.635 0 22.865 3.91 ;
        RECT 21.755 0 21.965 3.91 ;
        RECT 0 10.86 103.925 12.46 ;
        RECT 102.95 10.235 103.12 12.46 ;
        RECT 101.96 10.235 102.13 12.46 ;
        RECT 99.215 10.235 99.385 12.46 ;
        RECT 90.49 10.855 97.96 12.46 ;
        RECT 90.49 8.36 97.85 12.46 ;
        RECT 96.995 7.56 97.305 12.46 ;
        RECT 95.615 7.56 95.925 12.46 ;
        RECT 93.345 7.12 93.68 7.39 ;
        RECT 93.335 7.56 93.645 12.46 ;
        RECT 92.955 7.17 93.68 7.34 ;
        RECT 92.965 7.17 93.135 12.46 ;
        RECT 91.035 7.56 91.345 12.46 ;
        RECT 87.53 10.235 87.7 12.46 ;
        RECT 85.73 10.235 85.9 12.46 ;
        RECT 84.74 10.235 84.91 12.46 ;
        RECT 81.995 10.235 82.165 12.46 ;
        RECT 73.27 10.855 80.74 12.46 ;
        RECT 73.27 8.36 80.63 12.46 ;
        RECT 79.775 7.56 80.085 12.46 ;
        RECT 78.395 7.56 78.705 12.46 ;
        RECT 76.125 7.12 76.46 7.39 ;
        RECT 76.115 7.56 76.425 12.46 ;
        RECT 75.735 7.17 76.46 7.34 ;
        RECT 75.745 7.17 75.915 12.46 ;
        RECT 73.815 7.56 74.125 12.46 ;
        RECT 70.31 10.235 70.48 12.46 ;
        RECT 68.51 10.235 68.68 12.46 ;
        RECT 67.52 10.235 67.69 12.46 ;
        RECT 64.775 10.235 64.945 12.46 ;
        RECT 56.05 10.855 63.52 12.46 ;
        RECT 56.05 8.36 63.41 12.46 ;
        RECT 62.555 7.56 62.865 12.46 ;
        RECT 61.175 7.56 61.485 12.46 ;
        RECT 58.905 7.12 59.24 7.39 ;
        RECT 58.895 7.56 59.205 12.46 ;
        RECT 58.515 7.17 59.24 7.34 ;
        RECT 58.525 7.17 58.695 12.46 ;
        RECT 56.595 7.56 56.905 12.46 ;
        RECT 53.09 10.235 53.26 12.46 ;
        RECT 51.29 10.235 51.46 12.46 ;
        RECT 50.3 10.235 50.47 12.46 ;
        RECT 47.555 10.235 47.725 12.46 ;
        RECT 38.83 10.855 46.3 12.46 ;
        RECT 38.83 8.36 46.19 12.46 ;
        RECT 45.335 7.56 45.645 12.46 ;
        RECT 43.955 7.56 44.265 12.46 ;
        RECT 41.685 7.12 42.02 7.39 ;
        RECT 41.675 7.56 41.985 12.46 ;
        RECT 41.295 7.17 42.02 7.34 ;
        RECT 41.305 7.17 41.475 12.46 ;
        RECT 39.375 7.56 39.685 12.46 ;
        RECT 35.87 10.235 36.04 12.46 ;
        RECT 34.07 10.235 34.24 12.46 ;
        RECT 33.08 10.235 33.25 12.46 ;
        RECT 30.335 10.235 30.505 12.46 ;
        RECT 21.61 10.855 29.08 12.46 ;
        RECT 21.61 8.36 28.97 12.46 ;
        RECT 28.115 7.56 28.425 12.46 ;
        RECT 26.735 7.56 27.045 12.46 ;
        RECT 24.465 7.12 24.8 7.39 ;
        RECT 24.455 7.56 24.765 12.46 ;
        RECT 24.075 7.17 24.8 7.34 ;
        RECT 24.085 7.17 24.255 12.46 ;
        RECT 22.155 7.56 22.465 12.46 ;
        RECT 18.65 10.235 18.82 12.46 ;
        RECT 15.24 10.235 15.41 12.46 ;
        RECT 91.045 7.12 91.38 7.39 ;
        RECT 90.575 7.17 91.38 7.34 ;
        RECT 88.545 8.365 88.715 10.315 ;
        RECT 88.485 10.145 88.655 10.595 ;
        RECT 88.485 7.305 88.655 8.535 ;
        RECT 73.825 7.12 74.16 7.39 ;
        RECT 73.355 7.17 74.16 7.34 ;
        RECT 71.325 8.365 71.495 10.315 ;
        RECT 71.265 10.145 71.435 10.595 ;
        RECT 71.265 7.305 71.435 8.535 ;
        RECT 56.605 7.12 56.94 7.39 ;
        RECT 56.135 7.17 56.94 7.34 ;
        RECT 54.105 8.365 54.275 10.315 ;
        RECT 54.045 10.145 54.215 10.595 ;
        RECT 54.045 7.305 54.215 8.535 ;
        RECT 39.385 7.12 39.72 7.39 ;
        RECT 38.915 7.17 39.72 7.34 ;
        RECT 36.885 8.365 37.055 10.315 ;
        RECT 36.825 10.145 36.995 10.595 ;
        RECT 36.825 7.305 36.995 8.535 ;
        RECT 22.165 7.12 22.5 7.39 ;
        RECT 21.695 7.17 22.5 7.34 ;
        RECT 19.665 8.365 19.835 10.315 ;
        RECT 19.605 10.145 19.775 10.595 ;
        RECT 19.605 7.305 19.775 8.535 ;
      LAYER met1 ;
        RECT 0.015 0 103.925 1.6 ;
        RECT 90.485 0 98.145 3.12 ;
        RECT 73.265 0 80.925 3.12 ;
        RECT 56.045 0 63.705 3.12 ;
        RECT 38.825 0 46.485 3.12 ;
        RECT 21.605 0 29.265 3.12 ;
        RECT 0 10.86 103.925 12.46 ;
        RECT 90.49 10.855 97.96 12.46 ;
        RECT 90.49 8.33 97.85 12.46 ;
        RECT 88.485 8.575 88.775 8.805 ;
        RECT 88.08 8.6 88.775 8.775 ;
        RECT 88.08 8.6 88.25 12.46 ;
        RECT 73.27 10.855 80.74 12.46 ;
        RECT 73.27 8.33 80.63 12.46 ;
        RECT 71.265 8.575 71.555 8.805 ;
        RECT 70.86 8.6 71.555 8.775 ;
        RECT 70.86 8.6 71.03 12.46 ;
        RECT 56.05 10.855 63.52 12.46 ;
        RECT 56.05 8.33 63.41 12.46 ;
        RECT 54.045 8.575 54.335 8.805 ;
        RECT 53.64 8.6 54.335 8.775 ;
        RECT 53.64 8.6 53.81 12.46 ;
        RECT 38.83 10.855 46.3 12.46 ;
        RECT 38.83 8.33 46.19 12.46 ;
        RECT 36.825 8.575 37.115 8.805 ;
        RECT 36.42 8.6 37.115 8.775 ;
        RECT 36.42 8.6 36.59 12.46 ;
        RECT 21.61 10.855 29.08 12.46 ;
        RECT 21.61 8.33 28.97 12.46 ;
        RECT 19.605 8.575 19.895 8.805 ;
        RECT 19.2 8.6 19.895 8.775 ;
        RECT 19.2 8.6 19.37 12.46 ;
        RECT 92.88 7.125 93.2 7.385 ;
        RECT 90.515 7.185 93.2 7.325 ;
        RECT 90.515 7.14 90.805 7.37 ;
        RECT 75.66 7.125 75.98 7.385 ;
        RECT 73.295 7.185 75.98 7.325 ;
        RECT 73.295 7.14 73.585 7.37 ;
        RECT 58.44 7.125 58.76 7.385 ;
        RECT 56.075 7.185 58.76 7.325 ;
        RECT 56.075 7.14 56.365 7.37 ;
        RECT 41.22 7.125 41.54 7.385 ;
        RECT 38.855 7.185 41.54 7.325 ;
        RECT 38.855 7.14 39.145 7.37 ;
        RECT 24 7.125 24.32 7.385 ;
        RECT 21.635 7.185 24.32 7.325 ;
        RECT 21.635 7.14 21.925 7.37 ;
      LAYER via1 ;
        RECT 24.085 7.18 24.235 7.33 ;
        RECT 41.305 7.18 41.455 7.33 ;
        RECT 58.525 7.18 58.675 7.33 ;
        RECT 75.745 7.18 75.895 7.33 ;
        RECT 92.965 7.18 93.115 7.33 ;
      LAYER via2 ;
        RECT 24.06 7.15 24.26 7.35 ;
        RECT 41.28 7.15 41.48 7.35 ;
        RECT 58.5 7.15 58.7 7.35 ;
        RECT 75.72 7.15 75.92 7.35 ;
        RECT 92.94 7.15 93.14 7.35 ;
      LAYER mcon ;
        RECT 15.32 10.895 15.49 11.065 ;
        RECT 16 10.895 16.17 11.065 ;
        RECT 16.68 10.895 16.85 11.065 ;
        RECT 17.36 10.895 17.53 11.065 ;
        RECT 18.73 10.895 18.9 11.065 ;
        RECT 19.41 10.895 19.58 11.065 ;
        RECT 19.665 8.605 19.835 8.775 ;
        RECT 20.09 10.895 20.26 11.065 ;
        RECT 20.77 10.895 20.94 11.065 ;
        RECT 21.695 7.17 21.865 7.34 ;
        RECT 21.755 8.36 21.925 8.53 ;
        RECT 21.755 2.92 21.925 3.09 ;
        RECT 22.215 8.36 22.385 8.53 ;
        RECT 22.215 2.92 22.385 3.09 ;
        RECT 22.675 8.36 22.845 8.53 ;
        RECT 22.675 2.92 22.845 3.09 ;
        RECT 23.135 8.36 23.305 8.53 ;
        RECT 23.135 2.92 23.305 3.09 ;
        RECT 23.595 8.36 23.765 8.53 ;
        RECT 23.595 2.92 23.765 3.09 ;
        RECT 24.055 8.36 24.225 8.53 ;
        RECT 24.055 2.92 24.225 3.09 ;
        RECT 24.075 7.17 24.245 7.34 ;
        RECT 24.515 8.36 24.685 8.53 ;
        RECT 24.515 2.92 24.685 3.09 ;
        RECT 24.975 8.36 25.145 8.53 ;
        RECT 24.975 2.92 25.145 3.09 ;
        RECT 25.435 8.36 25.605 8.53 ;
        RECT 25.435 2.92 25.605 3.09 ;
        RECT 25.895 8.36 26.065 8.53 ;
        RECT 25.895 2.92 26.065 3.09 ;
        RECT 26.355 8.36 26.525 8.53 ;
        RECT 26.355 2.92 26.525 3.09 ;
        RECT 26.815 8.36 26.985 8.53 ;
        RECT 26.815 2.92 26.985 3.09 ;
        RECT 27.275 8.36 27.445 8.53 ;
        RECT 27.275 2.92 27.445 3.09 ;
        RECT 27.735 8.36 27.905 8.53 ;
        RECT 27.735 2.92 27.905 3.09 ;
        RECT 28.195 8.36 28.365 8.53 ;
        RECT 28.195 2.92 28.365 3.09 ;
        RECT 28.655 8.36 28.825 8.53 ;
        RECT 28.655 2.92 28.825 3.09 ;
        RECT 30.415 10.895 30.585 11.065 ;
        RECT 30.415 1.395 30.585 1.565 ;
        RECT 31.095 10.895 31.265 11.065 ;
        RECT 31.095 1.395 31.265 1.565 ;
        RECT 31.775 10.895 31.945 11.065 ;
        RECT 31.775 1.395 31.945 1.565 ;
        RECT 32.455 10.895 32.625 11.065 ;
        RECT 32.455 1.395 32.625 1.565 ;
        RECT 33.16 10.895 33.33 11.065 ;
        RECT 33.16 1.395 33.33 1.565 ;
        RECT 34.145 1.395 34.315 1.565 ;
        RECT 34.15 10.895 34.32 11.065 ;
        RECT 35.95 10.895 36.12 11.065 ;
        RECT 36.63 10.895 36.8 11.065 ;
        RECT 36.885 8.605 37.055 8.775 ;
        RECT 37.31 10.895 37.48 11.065 ;
        RECT 37.99 10.895 38.16 11.065 ;
        RECT 38.915 7.17 39.085 7.34 ;
        RECT 38.975 8.36 39.145 8.53 ;
        RECT 38.975 2.92 39.145 3.09 ;
        RECT 39.435 8.36 39.605 8.53 ;
        RECT 39.435 2.92 39.605 3.09 ;
        RECT 39.895 8.36 40.065 8.53 ;
        RECT 39.895 2.92 40.065 3.09 ;
        RECT 40.355 8.36 40.525 8.53 ;
        RECT 40.355 2.92 40.525 3.09 ;
        RECT 40.815 8.36 40.985 8.53 ;
        RECT 40.815 2.92 40.985 3.09 ;
        RECT 41.275 8.36 41.445 8.53 ;
        RECT 41.275 2.92 41.445 3.09 ;
        RECT 41.295 7.17 41.465 7.34 ;
        RECT 41.735 8.36 41.905 8.53 ;
        RECT 41.735 2.92 41.905 3.09 ;
        RECT 42.195 8.36 42.365 8.53 ;
        RECT 42.195 2.92 42.365 3.09 ;
        RECT 42.655 8.36 42.825 8.53 ;
        RECT 42.655 2.92 42.825 3.09 ;
        RECT 43.115 8.36 43.285 8.53 ;
        RECT 43.115 2.92 43.285 3.09 ;
        RECT 43.575 8.36 43.745 8.53 ;
        RECT 43.575 2.92 43.745 3.09 ;
        RECT 44.035 8.36 44.205 8.53 ;
        RECT 44.035 2.92 44.205 3.09 ;
        RECT 44.495 8.36 44.665 8.53 ;
        RECT 44.495 2.92 44.665 3.09 ;
        RECT 44.955 8.36 45.125 8.53 ;
        RECT 44.955 2.92 45.125 3.09 ;
        RECT 45.415 8.36 45.585 8.53 ;
        RECT 45.415 2.92 45.585 3.09 ;
        RECT 45.875 8.36 46.045 8.53 ;
        RECT 45.875 2.92 46.045 3.09 ;
        RECT 47.635 10.895 47.805 11.065 ;
        RECT 47.635 1.395 47.805 1.565 ;
        RECT 48.315 10.895 48.485 11.065 ;
        RECT 48.315 1.395 48.485 1.565 ;
        RECT 48.995 10.895 49.165 11.065 ;
        RECT 48.995 1.395 49.165 1.565 ;
        RECT 49.675 10.895 49.845 11.065 ;
        RECT 49.675 1.395 49.845 1.565 ;
        RECT 50.38 10.895 50.55 11.065 ;
        RECT 50.38 1.395 50.55 1.565 ;
        RECT 51.365 1.395 51.535 1.565 ;
        RECT 51.37 10.895 51.54 11.065 ;
        RECT 53.17 10.895 53.34 11.065 ;
        RECT 53.85 10.895 54.02 11.065 ;
        RECT 54.105 8.605 54.275 8.775 ;
        RECT 54.53 10.895 54.7 11.065 ;
        RECT 55.21 10.895 55.38 11.065 ;
        RECT 56.135 7.17 56.305 7.34 ;
        RECT 56.195 8.36 56.365 8.53 ;
        RECT 56.195 2.92 56.365 3.09 ;
        RECT 56.655 8.36 56.825 8.53 ;
        RECT 56.655 2.92 56.825 3.09 ;
        RECT 57.115 8.36 57.285 8.53 ;
        RECT 57.115 2.92 57.285 3.09 ;
        RECT 57.575 8.36 57.745 8.53 ;
        RECT 57.575 2.92 57.745 3.09 ;
        RECT 58.035 8.36 58.205 8.53 ;
        RECT 58.035 2.92 58.205 3.09 ;
        RECT 58.495 8.36 58.665 8.53 ;
        RECT 58.495 2.92 58.665 3.09 ;
        RECT 58.515 7.17 58.685 7.34 ;
        RECT 58.955 8.36 59.125 8.53 ;
        RECT 58.955 2.92 59.125 3.09 ;
        RECT 59.415 8.36 59.585 8.53 ;
        RECT 59.415 2.92 59.585 3.09 ;
        RECT 59.875 8.36 60.045 8.53 ;
        RECT 59.875 2.92 60.045 3.09 ;
        RECT 60.335 8.36 60.505 8.53 ;
        RECT 60.335 2.92 60.505 3.09 ;
        RECT 60.795 8.36 60.965 8.53 ;
        RECT 60.795 2.92 60.965 3.09 ;
        RECT 61.255 8.36 61.425 8.53 ;
        RECT 61.255 2.92 61.425 3.09 ;
        RECT 61.715 8.36 61.885 8.53 ;
        RECT 61.715 2.92 61.885 3.09 ;
        RECT 62.175 8.36 62.345 8.53 ;
        RECT 62.175 2.92 62.345 3.09 ;
        RECT 62.635 8.36 62.805 8.53 ;
        RECT 62.635 2.92 62.805 3.09 ;
        RECT 63.095 8.36 63.265 8.53 ;
        RECT 63.095 2.92 63.265 3.09 ;
        RECT 64.855 10.895 65.025 11.065 ;
        RECT 64.855 1.395 65.025 1.565 ;
        RECT 65.535 10.895 65.705 11.065 ;
        RECT 65.535 1.395 65.705 1.565 ;
        RECT 66.215 10.895 66.385 11.065 ;
        RECT 66.215 1.395 66.385 1.565 ;
        RECT 66.895 10.895 67.065 11.065 ;
        RECT 66.895 1.395 67.065 1.565 ;
        RECT 67.6 10.895 67.77 11.065 ;
        RECT 67.6 1.395 67.77 1.565 ;
        RECT 68.585 1.395 68.755 1.565 ;
        RECT 68.59 10.895 68.76 11.065 ;
        RECT 70.39 10.895 70.56 11.065 ;
        RECT 71.07 10.895 71.24 11.065 ;
        RECT 71.325 8.605 71.495 8.775 ;
        RECT 71.75 10.895 71.92 11.065 ;
        RECT 72.43 10.895 72.6 11.065 ;
        RECT 73.355 7.17 73.525 7.34 ;
        RECT 73.415 8.36 73.585 8.53 ;
        RECT 73.415 2.92 73.585 3.09 ;
        RECT 73.875 8.36 74.045 8.53 ;
        RECT 73.875 2.92 74.045 3.09 ;
        RECT 74.335 8.36 74.505 8.53 ;
        RECT 74.335 2.92 74.505 3.09 ;
        RECT 74.795 8.36 74.965 8.53 ;
        RECT 74.795 2.92 74.965 3.09 ;
        RECT 75.255 8.36 75.425 8.53 ;
        RECT 75.255 2.92 75.425 3.09 ;
        RECT 75.715 8.36 75.885 8.53 ;
        RECT 75.715 2.92 75.885 3.09 ;
        RECT 75.735 7.17 75.905 7.34 ;
        RECT 76.175 8.36 76.345 8.53 ;
        RECT 76.175 2.92 76.345 3.09 ;
        RECT 76.635 8.36 76.805 8.53 ;
        RECT 76.635 2.92 76.805 3.09 ;
        RECT 77.095 8.36 77.265 8.53 ;
        RECT 77.095 2.92 77.265 3.09 ;
        RECT 77.555 8.36 77.725 8.53 ;
        RECT 77.555 2.92 77.725 3.09 ;
        RECT 78.015 8.36 78.185 8.53 ;
        RECT 78.015 2.92 78.185 3.09 ;
        RECT 78.475 8.36 78.645 8.53 ;
        RECT 78.475 2.92 78.645 3.09 ;
        RECT 78.935 8.36 79.105 8.53 ;
        RECT 78.935 2.92 79.105 3.09 ;
        RECT 79.395 8.36 79.565 8.53 ;
        RECT 79.395 2.92 79.565 3.09 ;
        RECT 79.855 8.36 80.025 8.53 ;
        RECT 79.855 2.92 80.025 3.09 ;
        RECT 80.315 8.36 80.485 8.53 ;
        RECT 80.315 2.92 80.485 3.09 ;
        RECT 82.075 10.895 82.245 11.065 ;
        RECT 82.075 1.395 82.245 1.565 ;
        RECT 82.755 10.895 82.925 11.065 ;
        RECT 82.755 1.395 82.925 1.565 ;
        RECT 83.435 10.895 83.605 11.065 ;
        RECT 83.435 1.395 83.605 1.565 ;
        RECT 84.115 10.895 84.285 11.065 ;
        RECT 84.115 1.395 84.285 1.565 ;
        RECT 84.82 10.895 84.99 11.065 ;
        RECT 84.82 1.395 84.99 1.565 ;
        RECT 85.805 1.395 85.975 1.565 ;
        RECT 85.81 10.895 85.98 11.065 ;
        RECT 87.61 10.895 87.78 11.065 ;
        RECT 88.29 10.895 88.46 11.065 ;
        RECT 88.545 8.605 88.715 8.775 ;
        RECT 88.97 10.895 89.14 11.065 ;
        RECT 89.65 10.895 89.82 11.065 ;
        RECT 90.575 7.17 90.745 7.34 ;
        RECT 90.635 8.36 90.805 8.53 ;
        RECT 90.635 2.92 90.805 3.09 ;
        RECT 91.095 8.36 91.265 8.53 ;
        RECT 91.095 2.92 91.265 3.09 ;
        RECT 91.555 8.36 91.725 8.53 ;
        RECT 91.555 2.92 91.725 3.09 ;
        RECT 92.015 8.36 92.185 8.53 ;
        RECT 92.015 2.92 92.185 3.09 ;
        RECT 92.475 8.36 92.645 8.53 ;
        RECT 92.475 2.92 92.645 3.09 ;
        RECT 92.935 8.36 93.105 8.53 ;
        RECT 92.935 2.92 93.105 3.09 ;
        RECT 92.955 7.17 93.125 7.34 ;
        RECT 93.395 8.36 93.565 8.53 ;
        RECT 93.395 2.92 93.565 3.09 ;
        RECT 93.855 8.36 94.025 8.53 ;
        RECT 93.855 2.92 94.025 3.09 ;
        RECT 94.315 8.36 94.485 8.53 ;
        RECT 94.315 2.92 94.485 3.09 ;
        RECT 94.775 8.36 94.945 8.53 ;
        RECT 94.775 2.92 94.945 3.09 ;
        RECT 95.235 8.36 95.405 8.53 ;
        RECT 95.235 2.92 95.405 3.09 ;
        RECT 95.695 8.36 95.865 8.53 ;
        RECT 95.695 2.92 95.865 3.09 ;
        RECT 96.155 8.36 96.325 8.53 ;
        RECT 96.155 2.92 96.325 3.09 ;
        RECT 96.615 8.36 96.785 8.53 ;
        RECT 96.615 2.92 96.785 3.09 ;
        RECT 97.075 8.36 97.245 8.53 ;
        RECT 97.075 2.92 97.245 3.09 ;
        RECT 97.535 8.36 97.705 8.53 ;
        RECT 97.535 2.92 97.705 3.09 ;
        RECT 99.295 10.895 99.465 11.065 ;
        RECT 99.295 1.395 99.465 1.565 ;
        RECT 99.975 10.895 100.145 11.065 ;
        RECT 99.975 1.395 100.145 1.565 ;
        RECT 100.655 10.895 100.825 11.065 ;
        RECT 100.655 1.395 100.825 1.565 ;
        RECT 101.335 10.895 101.505 11.065 ;
        RECT 101.335 1.395 101.505 1.565 ;
        RECT 102.04 10.895 102.21 11.065 ;
        RECT 102.04 1.395 102.21 1.565 ;
        RECT 103.025 1.395 103.195 1.565 ;
        RECT 103.03 10.895 103.2 11.065 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 88.82 9.285 89.19 9.655 ;
      RECT 88.82 9.32 95.97 9.62 ;
      RECT 95.67 7.1 95.97 9.62 ;
      RECT 94.615 7.08 94.915 9.62 ;
      RECT 93.585 7.745 93.885 9.62 ;
      RECT 93.085 7.79 93.885 8.09 ;
      RECT 93.465 7.72 93.765 8.09 ;
      RECT 95.595 7.1 95.97 7.465 ;
      RECT 95.66 7.06 95.96 7.465 ;
      RECT 94.575 7.08 94.915 7.43 ;
      RECT 94.59 7.04 94.89 7.43 ;
      RECT 94.565 7.085 94.915 7.415 ;
      RECT 95.595 7.1 96.405 7.4 ;
      RECT 94.095 7.1 94.915 7.4 ;
      RECT 95.605 7.085 95.96 7.465 ;
      RECT 95.255 5.05 95.585 5.38 ;
      RECT 95.255 5.065 96.055 5.365 ;
      RECT 95.27 5.02 95.57 5.38 ;
      RECT 94.915 4.37 95.245 4.7 ;
      RECT 94.915 4.385 95.715 4.685 ;
      RECT 95 4.36 95.3 4.685 ;
      RECT 94.235 5.45 94.565 5.78 ;
      RECT 92.195 5.45 92.525 5.78 ;
      RECT 92.195 5.465 94.565 5.765 ;
      RECT 93.885 4.71 94.215 5.04 ;
      RECT 93.425 4.725 94.225 5.025 ;
      RECT 93.555 3.52 93.885 3.85 ;
      RECT 93.085 3.535 93.885 3.835 ;
      RECT 93.545 3.53 93.885 3.835 ;
      RECT 71.6 9.285 71.97 9.655 ;
      RECT 71.6 9.32 78.75 9.62 ;
      RECT 78.45 7.1 78.75 9.62 ;
      RECT 77.395 7.08 77.695 9.62 ;
      RECT 76.365 7.745 76.665 9.62 ;
      RECT 75.865 7.79 76.665 8.09 ;
      RECT 76.245 7.72 76.545 8.09 ;
      RECT 78.375 7.1 78.75 7.465 ;
      RECT 78.44 7.06 78.74 7.465 ;
      RECT 77.355 7.08 77.695 7.43 ;
      RECT 77.37 7.04 77.67 7.43 ;
      RECT 77.345 7.085 77.695 7.415 ;
      RECT 78.375 7.1 79.185 7.4 ;
      RECT 76.875 7.1 77.695 7.4 ;
      RECT 78.385 7.085 78.74 7.465 ;
      RECT 78.035 5.05 78.365 5.38 ;
      RECT 78.035 5.065 78.835 5.365 ;
      RECT 78.05 5.02 78.35 5.38 ;
      RECT 77.695 4.37 78.025 4.7 ;
      RECT 77.695 4.385 78.495 4.685 ;
      RECT 77.78 4.36 78.08 4.685 ;
      RECT 77.015 5.45 77.345 5.78 ;
      RECT 74.975 5.45 75.305 5.78 ;
      RECT 74.975 5.465 77.345 5.765 ;
      RECT 76.665 4.71 76.995 5.04 ;
      RECT 76.205 4.725 77.005 5.025 ;
      RECT 76.335 3.52 76.665 3.85 ;
      RECT 75.865 3.535 76.665 3.835 ;
      RECT 76.325 3.53 76.665 3.835 ;
      RECT 54.38 9.285 54.75 9.655 ;
      RECT 54.38 9.32 61.53 9.62 ;
      RECT 61.23 7.1 61.53 9.62 ;
      RECT 60.175 7.08 60.475 9.62 ;
      RECT 59.145 7.745 59.445 9.62 ;
      RECT 58.645 7.79 59.445 8.09 ;
      RECT 59.025 7.72 59.325 8.09 ;
      RECT 61.155 7.1 61.53 7.465 ;
      RECT 61.22 7.06 61.52 7.465 ;
      RECT 60.135 7.08 60.475 7.43 ;
      RECT 60.15 7.04 60.45 7.43 ;
      RECT 60.125 7.085 60.475 7.415 ;
      RECT 61.155 7.1 61.965 7.4 ;
      RECT 59.655 7.1 60.475 7.4 ;
      RECT 61.165 7.085 61.52 7.465 ;
      RECT 60.815 5.05 61.145 5.38 ;
      RECT 60.815 5.065 61.615 5.365 ;
      RECT 60.83 5.02 61.13 5.38 ;
      RECT 60.475 4.37 60.805 4.7 ;
      RECT 60.475 4.385 61.275 4.685 ;
      RECT 60.56 4.36 60.86 4.685 ;
      RECT 59.795 5.45 60.125 5.78 ;
      RECT 57.755 5.45 58.085 5.78 ;
      RECT 57.755 5.465 60.125 5.765 ;
      RECT 59.445 4.71 59.775 5.04 ;
      RECT 58.985 4.725 59.785 5.025 ;
      RECT 59.115 3.52 59.445 3.85 ;
      RECT 58.645 3.535 59.445 3.835 ;
      RECT 59.105 3.53 59.445 3.835 ;
      RECT 37.16 9.285 37.53 9.655 ;
      RECT 37.16 9.32 44.31 9.62 ;
      RECT 44.01 7.1 44.31 9.62 ;
      RECT 42.955 7.08 43.255 9.62 ;
      RECT 41.925 7.745 42.225 9.62 ;
      RECT 41.425 7.79 42.225 8.09 ;
      RECT 41.805 7.72 42.105 8.09 ;
      RECT 43.935 7.1 44.31 7.465 ;
      RECT 44 7.06 44.3 7.465 ;
      RECT 42.915 7.08 43.255 7.43 ;
      RECT 42.93 7.04 43.23 7.43 ;
      RECT 42.905 7.085 43.255 7.415 ;
      RECT 43.935 7.1 44.745 7.4 ;
      RECT 42.435 7.1 43.255 7.4 ;
      RECT 43.945 7.085 44.3 7.465 ;
      RECT 43.595 5.05 43.925 5.38 ;
      RECT 43.595 5.065 44.395 5.365 ;
      RECT 43.61 5.02 43.91 5.38 ;
      RECT 43.255 4.37 43.585 4.7 ;
      RECT 43.255 4.385 44.055 4.685 ;
      RECT 43.34 4.36 43.64 4.685 ;
      RECT 42.575 5.45 42.905 5.78 ;
      RECT 40.535 5.45 40.865 5.78 ;
      RECT 40.535 5.465 42.905 5.765 ;
      RECT 42.225 4.71 42.555 5.04 ;
      RECT 41.765 4.725 42.565 5.025 ;
      RECT 41.895 3.52 42.225 3.85 ;
      RECT 41.425 3.535 42.225 3.835 ;
      RECT 41.885 3.53 42.225 3.835 ;
      RECT 19.94 9.285 20.31 9.655 ;
      RECT 19.94 9.32 27.09 9.62 ;
      RECT 26.79 7.1 27.09 9.62 ;
      RECT 25.735 7.08 26.035 9.62 ;
      RECT 24.705 7.745 25.005 9.62 ;
      RECT 24.205 7.79 25.005 8.09 ;
      RECT 24.585 7.72 24.885 8.09 ;
      RECT 26.715 7.1 27.09 7.465 ;
      RECT 26.78 7.06 27.08 7.465 ;
      RECT 25.695 7.08 26.035 7.43 ;
      RECT 25.71 7.04 26.01 7.43 ;
      RECT 25.685 7.085 26.035 7.415 ;
      RECT 26.715 7.1 27.525 7.4 ;
      RECT 25.215 7.1 26.035 7.4 ;
      RECT 26.725 7.085 27.08 7.465 ;
      RECT 26.375 5.05 26.705 5.38 ;
      RECT 26.375 5.065 27.175 5.365 ;
      RECT 26.39 5.02 26.69 5.38 ;
      RECT 26.035 4.37 26.365 4.7 ;
      RECT 26.035 4.385 26.835 4.685 ;
      RECT 26.12 4.36 26.42 4.685 ;
      RECT 25.355 5.45 25.685 5.78 ;
      RECT 23.315 5.45 23.645 5.78 ;
      RECT 23.315 5.465 25.685 5.765 ;
      RECT 25.005 4.71 25.335 5.04 ;
      RECT 24.545 4.725 25.345 5.025 ;
      RECT 24.675 3.52 25.005 3.85 ;
      RECT 24.205 3.535 25.005 3.835 ;
      RECT 24.665 3.53 25.005 3.835 ;
      RECT 103.28 7.2 103.66 12.46 ;
      RECT 86.06 7.2 86.44 12.46 ;
      RECT 68.84 7.2 69.22 12.46 ;
      RECT 51.62 7.2 52 12.46 ;
      RECT 34.4 7.2 34.78 12.46 ;
    LAYER via2 ;
      RECT 103.37 7.29 103.57 7.49 ;
      RECT 95.67 7.15 95.87 7.35 ;
      RECT 95.32 5.115 95.52 5.315 ;
      RECT 94.98 4.435 95.18 4.635 ;
      RECT 94.63 7.15 94.83 7.35 ;
      RECT 94.3 5.515 94.5 5.715 ;
      RECT 93.95 4.775 94.15 4.975 ;
      RECT 93.62 3.585 93.82 3.785 ;
      RECT 93.62 7.81 93.82 8.01 ;
      RECT 92.26 5.515 92.46 5.715 ;
      RECT 88.905 9.37 89.105 9.57 ;
      RECT 86.15 7.29 86.35 7.49 ;
      RECT 78.45 7.15 78.65 7.35 ;
      RECT 78.1 5.115 78.3 5.315 ;
      RECT 77.76 4.435 77.96 4.635 ;
      RECT 77.41 7.15 77.61 7.35 ;
      RECT 77.08 5.515 77.28 5.715 ;
      RECT 76.73 4.775 76.93 4.975 ;
      RECT 76.4 3.585 76.6 3.785 ;
      RECT 76.4 7.81 76.6 8.01 ;
      RECT 75.04 5.515 75.24 5.715 ;
      RECT 71.685 9.37 71.885 9.57 ;
      RECT 68.93 7.29 69.13 7.49 ;
      RECT 61.23 7.15 61.43 7.35 ;
      RECT 60.88 5.115 61.08 5.315 ;
      RECT 60.54 4.435 60.74 4.635 ;
      RECT 60.19 7.15 60.39 7.35 ;
      RECT 59.86 5.515 60.06 5.715 ;
      RECT 59.51 4.775 59.71 4.975 ;
      RECT 59.18 3.585 59.38 3.785 ;
      RECT 59.18 7.81 59.38 8.01 ;
      RECT 57.82 5.515 58.02 5.715 ;
      RECT 54.465 9.37 54.665 9.57 ;
      RECT 51.71 7.29 51.91 7.49 ;
      RECT 44.01 7.15 44.21 7.35 ;
      RECT 43.66 5.115 43.86 5.315 ;
      RECT 43.32 4.435 43.52 4.635 ;
      RECT 42.97 7.15 43.17 7.35 ;
      RECT 42.64 5.515 42.84 5.715 ;
      RECT 42.29 4.775 42.49 4.975 ;
      RECT 41.96 3.585 42.16 3.785 ;
      RECT 41.96 7.81 42.16 8.01 ;
      RECT 40.6 5.515 40.8 5.715 ;
      RECT 37.245 9.37 37.445 9.57 ;
      RECT 34.49 7.29 34.69 7.49 ;
      RECT 26.79 7.15 26.99 7.35 ;
      RECT 26.44 5.115 26.64 5.315 ;
      RECT 26.1 4.435 26.3 4.635 ;
      RECT 25.75 7.15 25.95 7.35 ;
      RECT 25.42 5.515 25.62 5.715 ;
      RECT 25.07 4.775 25.27 4.975 ;
      RECT 24.74 3.585 24.94 3.785 ;
      RECT 24.74 7.81 24.94 8.01 ;
      RECT 23.38 5.515 23.58 5.715 ;
      RECT 20.025 9.37 20.225 9.57 ;
    LAYER met2 ;
      RECT 16.245 10.065 103.555 10.235 ;
      RECT 103.385 9.585 103.555 10.235 ;
      RECT 16.245 8.54 16.415 10.235 ;
      RECT 103.35 9.585 103.675 9.91 ;
      RECT 16.19 8.54 16.47 8.88 ;
      RECT 100.195 8.565 100.515 8.89 ;
      RECT 100.225 7.98 100.395 8.89 ;
      RECT 100.225 7.98 100.4 8.33 ;
      RECT 100.225 7.98 101.2 8.155 ;
      RECT 101.025 3.26 101.2 8.155 ;
      RECT 94.94 4.35 95.22 4.72 ;
      RECT 95.01 3.64 95.185 4.72 ;
      RECT 95.01 3.64 98.23 3.815 ;
      RECT 98.055 3.32 98.23 3.815 ;
      RECT 98.525 3.29 98.85 3.615 ;
      RECT 100.97 3.26 101.32 3.61 ;
      RECT 98.055 3.32 101.32 3.49 ;
      RECT 89.345 9.65 100.04 9.82 ;
      RECT 99.88 3.69 100.04 9.82 ;
      RECT 89.345 8.83 89.515 9.82 ;
      RECT 86.165 8.945 86.49 9.27 ;
      RECT 100.995 8.94 101.32 9.265 ;
      RECT 99.88 9.03 101.32 9.2 ;
      RECT 89.295 8.83 89.575 9.17 ;
      RECT 86.165 8.975 87.155 9.145 ;
      RECT 87.155 8.97 89.575 9.14 ;
      RECT 100.195 3.66 100.515 3.98 ;
      RECT 99.88 3.69 100.515 3.86 ;
      RECT 96.65 7.76 96.91 8.095 ;
      RECT 96.71 4.035 96.85 8.095 ;
      RECT 96.65 4.035 96.91 4.355 ;
      RECT 95.97 6.075 96.23 6.395 ;
      RECT 96.03 5.055 96.17 6.395 ;
      RECT 95.97 5.055 96.23 5.375 ;
      RECT 94.95 7.76 95.21 8.095 ;
      RECT 94.92 7.805 95.24 8.05 ;
      RECT 95.01 6.505 95.15 8.095 ;
      RECT 94.33 6.505 95.15 6.645 ;
      RECT 94.33 4.035 94.47 6.645 ;
      RECT 94.26 5.43 94.54 5.8 ;
      RECT 94.27 4.035 94.53 4.355 ;
      RECT 92.22 5.43 92.5 5.8 ;
      RECT 92.29 3.695 92.43 5.8 ;
      RECT 92.23 3.695 92.49 4.015 ;
      RECT 91.55 6.075 91.81 6.395 ;
      RECT 91.61 4.035 91.75 6.395 ;
      RECT 91.55 4.035 91.81 4.355 ;
      RECT 82.975 8.565 83.295 8.89 ;
      RECT 83.005 7.98 83.175 8.89 ;
      RECT 83.005 7.98 83.18 8.33 ;
      RECT 83.005 7.98 83.98 8.155 ;
      RECT 83.805 3.26 83.98 8.155 ;
      RECT 77.72 4.35 78 4.72 ;
      RECT 77.79 3.64 77.965 4.72 ;
      RECT 77.79 3.64 81.01 3.815 ;
      RECT 80.835 3.32 81.01 3.815 ;
      RECT 81.305 3.29 81.63 3.615 ;
      RECT 83.75 3.26 84.1 3.61 ;
      RECT 80.835 3.32 84.1 3.49 ;
      RECT 72.125 9.65 82.82 9.82 ;
      RECT 82.66 3.69 82.82 9.82 ;
      RECT 72.125 8.83 72.295 9.82 ;
      RECT 68.945 8.945 69.27 9.27 ;
      RECT 83.775 8.94 84.1 9.265 ;
      RECT 82.66 9.03 84.1 9.2 ;
      RECT 72.075 8.83 72.355 9.17 ;
      RECT 68.945 8.975 69.89 9.145 ;
      RECT 69.89 8.97 72.355 9.14 ;
      RECT 82.975 3.66 83.295 3.98 ;
      RECT 82.66 3.69 83.295 3.86 ;
      RECT 79.43 7.76 79.69 8.095 ;
      RECT 79.49 4.035 79.63 8.095 ;
      RECT 79.43 4.035 79.69 4.355 ;
      RECT 78.75 6.075 79.01 6.395 ;
      RECT 78.81 5.055 78.95 6.395 ;
      RECT 78.75 5.055 79.01 5.375 ;
      RECT 77.73 7.76 77.99 8.095 ;
      RECT 77.7 7.805 78.02 8.05 ;
      RECT 77.79 6.505 77.93 8.095 ;
      RECT 77.11 6.505 77.93 6.645 ;
      RECT 77.11 4.035 77.25 6.645 ;
      RECT 77.04 5.43 77.32 5.8 ;
      RECT 77.05 4.035 77.31 4.355 ;
      RECT 75 5.43 75.28 5.8 ;
      RECT 75.07 3.695 75.21 5.8 ;
      RECT 75.01 3.695 75.27 4.015 ;
      RECT 74.33 6.075 74.59 6.395 ;
      RECT 74.39 4.035 74.53 6.395 ;
      RECT 74.33 4.035 74.59 4.355 ;
      RECT 65.755 8.565 66.075 8.89 ;
      RECT 65.785 7.98 65.955 8.89 ;
      RECT 65.785 7.98 65.96 8.33 ;
      RECT 65.785 7.98 66.76 8.155 ;
      RECT 66.585 3.26 66.76 8.155 ;
      RECT 60.5 4.35 60.78 4.72 ;
      RECT 60.57 3.64 60.745 4.72 ;
      RECT 60.57 3.64 63.79 3.815 ;
      RECT 63.615 3.32 63.79 3.815 ;
      RECT 64.085 3.29 64.41 3.615 ;
      RECT 66.53 3.26 66.88 3.61 ;
      RECT 63.615 3.32 66.88 3.49 ;
      RECT 54.905 9.65 65.6 9.82 ;
      RECT 65.44 3.69 65.6 9.82 ;
      RECT 54.905 8.83 55.075 9.82 ;
      RECT 51.725 8.945 52.05 9.27 ;
      RECT 66.555 8.94 66.88 9.265 ;
      RECT 65.44 9.03 66.88 9.2 ;
      RECT 54.855 8.83 55.135 9.17 ;
      RECT 51.725 8.975 52.65 9.145 ;
      RECT 51.725 8.975 55.145 9.14 ;
      RECT 53.675 8.97 55.145 9.14 ;
      RECT 65.755 3.66 66.075 3.98 ;
      RECT 65.44 3.69 66.075 3.86 ;
      RECT 62.21 7.76 62.47 8.095 ;
      RECT 62.27 4.035 62.41 8.095 ;
      RECT 62.21 4.035 62.47 4.355 ;
      RECT 61.53 6.075 61.79 6.395 ;
      RECT 61.59 5.055 61.73 6.395 ;
      RECT 61.53 5.055 61.79 5.375 ;
      RECT 60.51 7.76 60.77 8.095 ;
      RECT 60.48 7.805 60.8 8.05 ;
      RECT 60.57 6.505 60.71 8.095 ;
      RECT 59.89 6.505 60.71 6.645 ;
      RECT 59.89 4.035 60.03 6.645 ;
      RECT 59.82 5.43 60.1 5.8 ;
      RECT 59.83 4.035 60.09 4.355 ;
      RECT 57.78 5.43 58.06 5.8 ;
      RECT 57.85 3.695 57.99 5.8 ;
      RECT 57.79 3.695 58.05 4.015 ;
      RECT 57.11 6.075 57.37 6.395 ;
      RECT 57.17 4.035 57.31 6.395 ;
      RECT 57.11 4.035 57.37 4.355 ;
      RECT 48.535 8.565 48.855 8.89 ;
      RECT 48.565 7.98 48.735 8.89 ;
      RECT 48.565 7.98 48.74 8.33 ;
      RECT 48.565 7.98 49.54 8.155 ;
      RECT 49.365 3.26 49.54 8.155 ;
      RECT 43.28 4.35 43.56 4.72 ;
      RECT 43.35 3.64 43.525 4.72 ;
      RECT 43.35 3.64 46.57 3.815 ;
      RECT 46.395 3.32 46.57 3.815 ;
      RECT 46.865 3.29 47.19 3.615 ;
      RECT 49.31 3.26 49.66 3.61 ;
      RECT 46.395 3.32 49.66 3.49 ;
      RECT 37.685 9.65 48.38 9.82 ;
      RECT 48.22 3.69 48.38 9.82 ;
      RECT 37.685 8.83 37.855 9.82 ;
      RECT 34.505 8.945 34.83 9.27 ;
      RECT 49.335 8.94 49.66 9.265 ;
      RECT 48.22 9.03 49.66 9.2 ;
      RECT 37.635 8.83 37.915 9.17 ;
      RECT 34.505 8.975 35.415 9.145 ;
      RECT 35.415 8.97 37.915 9.14 ;
      RECT 48.535 3.66 48.855 3.98 ;
      RECT 48.22 3.69 48.855 3.86 ;
      RECT 44.99 7.76 45.25 8.095 ;
      RECT 45.05 4.035 45.19 8.095 ;
      RECT 44.99 4.035 45.25 4.355 ;
      RECT 44.31 6.075 44.57 6.395 ;
      RECT 44.37 5.055 44.51 6.395 ;
      RECT 44.31 5.055 44.57 5.375 ;
      RECT 43.29 7.76 43.55 8.095 ;
      RECT 43.26 7.805 43.58 8.05 ;
      RECT 43.35 6.505 43.49 8.095 ;
      RECT 42.67 6.505 43.49 6.645 ;
      RECT 42.67 4.035 42.81 6.645 ;
      RECT 42.6 5.43 42.88 5.8 ;
      RECT 42.61 4.035 42.87 4.355 ;
      RECT 40.56 5.43 40.84 5.8 ;
      RECT 40.63 3.695 40.77 5.8 ;
      RECT 40.57 3.695 40.83 4.015 ;
      RECT 39.89 6.075 40.15 6.395 ;
      RECT 39.95 4.035 40.09 6.395 ;
      RECT 39.89 4.035 40.15 4.355 ;
      RECT 31.315 8.565 31.635 8.89 ;
      RECT 31.345 7.98 31.515 8.89 ;
      RECT 31.345 7.98 31.52 8.33 ;
      RECT 31.345 7.98 32.32 8.155 ;
      RECT 32.145 3.26 32.32 8.155 ;
      RECT 26.06 4.35 26.34 4.72 ;
      RECT 26.13 3.64 26.305 4.72 ;
      RECT 26.13 3.64 29.35 3.815 ;
      RECT 29.175 3.32 29.35 3.815 ;
      RECT 29.645 3.29 29.97 3.615 ;
      RECT 32.09 3.26 32.44 3.61 ;
      RECT 29.175 3.32 32.44 3.49 ;
      RECT 20.465 9.65 31.16 9.82 ;
      RECT 31 3.69 31.16 9.82 ;
      RECT 20.465 8.83 20.635 9.82 ;
      RECT 16.565 9.28 16.845 9.62 ;
      RECT 16.565 9.345 17.775 9.515 ;
      RECT 17.605 8.97 17.775 9.515 ;
      RECT 32.115 8.94 32.44 9.265 ;
      RECT 31 9.03 32.44 9.2 ;
      RECT 20.415 8.83 20.695 9.17 ;
      RECT 17.605 8.97 20.695 9.14 ;
      RECT 31.315 3.66 31.635 3.98 ;
      RECT 31 3.69 31.635 3.86 ;
      RECT 27.77 7.76 28.03 8.095 ;
      RECT 27.83 4.035 27.97 8.095 ;
      RECT 27.77 4.035 28.03 4.355 ;
      RECT 27.09 6.075 27.35 6.395 ;
      RECT 27.15 5.055 27.29 6.395 ;
      RECT 27.09 5.055 27.35 5.375 ;
      RECT 26.07 7.76 26.33 8.095 ;
      RECT 26.04 7.805 26.36 8.05 ;
      RECT 26.13 6.505 26.27 8.095 ;
      RECT 25.45 6.505 26.27 6.645 ;
      RECT 25.45 4.035 25.59 6.645 ;
      RECT 25.38 5.43 25.66 5.8 ;
      RECT 25.39 4.035 25.65 4.355 ;
      RECT 23.34 5.43 23.62 5.8 ;
      RECT 23.41 3.695 23.55 5.8 ;
      RECT 23.35 3.695 23.61 4.015 ;
      RECT 22.67 6.075 22.93 6.395 ;
      RECT 22.73 4.035 22.87 6.395 ;
      RECT 22.67 4.035 22.93 4.355 ;
      RECT 103.28 7.2 103.66 7.58 ;
      RECT 95.63 7.065 95.91 7.435 ;
      RECT 95.28 5.03 95.56 5.4 ;
      RECT 94.59 7.065 94.87 7.435 ;
      RECT 93.91 4.69 94.19 5.06 ;
      RECT 93.58 3.5 93.86 3.87 ;
      RECT 93.58 7.725 93.86 8.095 ;
      RECT 88.82 9.285 89.19 9.655 ;
      RECT 86.06 7.2 86.44 7.58 ;
      RECT 78.41 7.065 78.69 7.435 ;
      RECT 78.06 5.03 78.34 5.4 ;
      RECT 77.37 7.065 77.65 7.435 ;
      RECT 76.69 4.69 76.97 5.06 ;
      RECT 76.36 3.5 76.64 3.87 ;
      RECT 76.36 7.725 76.64 8.095 ;
      RECT 71.6 9.285 71.97 9.655 ;
      RECT 68.84 7.2 69.22 7.58 ;
      RECT 61.19 7.065 61.47 7.435 ;
      RECT 60.84 5.03 61.12 5.4 ;
      RECT 60.15 7.065 60.43 7.435 ;
      RECT 59.47 4.69 59.75 5.06 ;
      RECT 59.14 3.5 59.42 3.87 ;
      RECT 59.14 7.725 59.42 8.095 ;
      RECT 54.38 9.285 54.75 9.655 ;
      RECT 51.62 7.2 52 7.58 ;
      RECT 43.97 7.065 44.25 7.435 ;
      RECT 43.62 5.03 43.9 5.4 ;
      RECT 42.93 7.065 43.21 7.435 ;
      RECT 42.25 4.69 42.53 5.06 ;
      RECT 41.92 3.5 42.2 3.87 ;
      RECT 41.92 7.725 42.2 8.095 ;
      RECT 37.16 9.285 37.53 9.655 ;
      RECT 34.4 7.2 34.78 7.58 ;
      RECT 26.75 7.065 27.03 7.435 ;
      RECT 26.4 5.03 26.68 5.4 ;
      RECT 25.71 7.065 25.99 7.435 ;
      RECT 25.03 4.69 25.31 5.06 ;
      RECT 24.7 3.5 24.98 3.87 ;
      RECT 24.7 7.725 24.98 8.095 ;
      RECT 19.94 9.285 20.31 9.655 ;
    LAYER via1 ;
      RECT 103.44 9.67 103.59 9.82 ;
      RECT 103.395 7.315 103.545 7.465 ;
      RECT 101.085 9.025 101.235 9.175 ;
      RECT 101.07 3.36 101.22 3.51 ;
      RECT 100.28 3.745 100.43 3.895 ;
      RECT 100.28 8.655 100.43 8.805 ;
      RECT 98.615 3.375 98.765 3.525 ;
      RECT 96.705 4.12 96.855 4.27 ;
      RECT 96.705 7.845 96.855 7.995 ;
      RECT 96.025 5.14 96.175 5.29 ;
      RECT 96.025 6.16 96.175 6.31 ;
      RECT 95.685 7.165 95.835 7.315 ;
      RECT 95.345 5.14 95.495 5.29 ;
      RECT 95.005 4.46 95.155 4.61 ;
      RECT 95.005 7.845 95.155 7.995 ;
      RECT 94.655 7.165 94.805 7.315 ;
      RECT 94.325 4.12 94.475 4.27 ;
      RECT 93.985 4.8 94.135 4.95 ;
      RECT 93.645 3.61 93.795 3.76 ;
      RECT 93.645 7.83 93.795 7.98 ;
      RECT 92.285 3.78 92.435 3.93 ;
      RECT 91.605 4.12 91.755 4.27 ;
      RECT 91.605 6.16 91.755 6.31 ;
      RECT 89.36 8.925 89.51 9.075 ;
      RECT 88.93 9.395 89.08 9.545 ;
      RECT 86.255 9.03 86.405 9.18 ;
      RECT 86.175 7.315 86.325 7.465 ;
      RECT 83.865 9.025 84.015 9.175 ;
      RECT 83.85 3.36 84 3.51 ;
      RECT 83.06 3.745 83.21 3.895 ;
      RECT 83.06 8.655 83.21 8.805 ;
      RECT 81.395 3.375 81.545 3.525 ;
      RECT 79.485 4.12 79.635 4.27 ;
      RECT 79.485 7.845 79.635 7.995 ;
      RECT 78.805 5.14 78.955 5.29 ;
      RECT 78.805 6.16 78.955 6.31 ;
      RECT 78.465 7.165 78.615 7.315 ;
      RECT 78.125 5.14 78.275 5.29 ;
      RECT 77.785 4.46 77.935 4.61 ;
      RECT 77.785 7.845 77.935 7.995 ;
      RECT 77.435 7.165 77.585 7.315 ;
      RECT 77.105 4.12 77.255 4.27 ;
      RECT 76.765 4.8 76.915 4.95 ;
      RECT 76.425 3.61 76.575 3.76 ;
      RECT 76.425 7.83 76.575 7.98 ;
      RECT 75.065 3.78 75.215 3.93 ;
      RECT 74.385 4.12 74.535 4.27 ;
      RECT 74.385 6.16 74.535 6.31 ;
      RECT 72.14 8.925 72.29 9.075 ;
      RECT 71.71 9.395 71.86 9.545 ;
      RECT 69.035 9.03 69.185 9.18 ;
      RECT 68.955 7.315 69.105 7.465 ;
      RECT 66.645 9.025 66.795 9.175 ;
      RECT 66.63 3.36 66.78 3.51 ;
      RECT 65.84 3.745 65.99 3.895 ;
      RECT 65.84 8.655 65.99 8.805 ;
      RECT 64.175 3.375 64.325 3.525 ;
      RECT 62.265 4.12 62.415 4.27 ;
      RECT 62.265 7.845 62.415 7.995 ;
      RECT 61.585 5.14 61.735 5.29 ;
      RECT 61.585 6.16 61.735 6.31 ;
      RECT 61.245 7.165 61.395 7.315 ;
      RECT 60.905 5.14 61.055 5.29 ;
      RECT 60.565 4.46 60.715 4.61 ;
      RECT 60.565 7.845 60.715 7.995 ;
      RECT 60.215 7.165 60.365 7.315 ;
      RECT 59.885 4.12 60.035 4.27 ;
      RECT 59.545 4.8 59.695 4.95 ;
      RECT 59.205 3.61 59.355 3.76 ;
      RECT 59.205 7.83 59.355 7.98 ;
      RECT 57.845 3.78 57.995 3.93 ;
      RECT 57.165 4.12 57.315 4.27 ;
      RECT 57.165 6.16 57.315 6.31 ;
      RECT 54.92 8.925 55.07 9.075 ;
      RECT 54.49 9.395 54.64 9.545 ;
      RECT 51.815 9.03 51.965 9.18 ;
      RECT 51.735 7.315 51.885 7.465 ;
      RECT 49.425 9.025 49.575 9.175 ;
      RECT 49.41 3.36 49.56 3.51 ;
      RECT 48.62 3.745 48.77 3.895 ;
      RECT 48.62 8.655 48.77 8.805 ;
      RECT 46.955 3.375 47.105 3.525 ;
      RECT 45.045 4.12 45.195 4.27 ;
      RECT 45.045 7.845 45.195 7.995 ;
      RECT 44.365 5.14 44.515 5.29 ;
      RECT 44.365 6.16 44.515 6.31 ;
      RECT 44.025 7.165 44.175 7.315 ;
      RECT 43.685 5.14 43.835 5.29 ;
      RECT 43.345 4.46 43.495 4.61 ;
      RECT 43.345 7.845 43.495 7.995 ;
      RECT 42.995 7.165 43.145 7.315 ;
      RECT 42.665 4.12 42.815 4.27 ;
      RECT 42.325 4.8 42.475 4.95 ;
      RECT 41.985 3.61 42.135 3.76 ;
      RECT 41.985 7.83 42.135 7.98 ;
      RECT 40.625 3.78 40.775 3.93 ;
      RECT 39.945 4.12 40.095 4.27 ;
      RECT 39.945 6.16 40.095 6.31 ;
      RECT 37.7 8.925 37.85 9.075 ;
      RECT 37.27 9.395 37.42 9.545 ;
      RECT 34.595 9.03 34.745 9.18 ;
      RECT 34.515 7.315 34.665 7.465 ;
      RECT 32.205 9.025 32.355 9.175 ;
      RECT 32.19 3.36 32.34 3.51 ;
      RECT 31.4 3.745 31.55 3.895 ;
      RECT 31.4 8.655 31.55 8.805 ;
      RECT 29.735 3.375 29.885 3.525 ;
      RECT 27.825 4.12 27.975 4.27 ;
      RECT 27.825 7.845 27.975 7.995 ;
      RECT 27.145 5.14 27.295 5.29 ;
      RECT 27.145 6.16 27.295 6.31 ;
      RECT 26.805 7.165 26.955 7.315 ;
      RECT 26.465 5.14 26.615 5.29 ;
      RECT 26.125 4.46 26.275 4.61 ;
      RECT 26.125 7.845 26.275 7.995 ;
      RECT 25.775 7.165 25.925 7.315 ;
      RECT 25.445 4.12 25.595 4.27 ;
      RECT 25.105 4.8 25.255 4.95 ;
      RECT 24.765 3.61 24.915 3.76 ;
      RECT 24.765 7.83 24.915 7.98 ;
      RECT 23.405 3.78 23.555 3.93 ;
      RECT 22.725 4.12 22.875 4.27 ;
      RECT 22.725 6.16 22.875 6.31 ;
      RECT 20.48 8.925 20.63 9.075 ;
      RECT 20.05 9.395 20.2 9.545 ;
      RECT 16.63 9.375 16.78 9.525 ;
      RECT 16.255 8.635 16.405 8.785 ;
    LAYER met1 ;
      RECT 103.32 10.055 103.615 10.285 ;
      RECT 103.38 9.585 103.555 10.285 ;
      RECT 103.35 9.585 103.675 9.91 ;
      RECT 103.38 8.575 103.55 10.285 ;
      RECT 103.32 8.575 103.61 8.805 ;
      RECT 102.33 10.055 102.625 10.285 ;
      RECT 102.39 8.575 102.56 10.285 ;
      RECT 102.33 8.575 102.62 8.805 ;
      RECT 102.33 8.61 103.18 8.77 ;
      RECT 103.015 8.205 103.18 8.77 ;
      RECT 102.33 8.605 102.725 8.77 ;
      RECT 102.95 8.205 103.24 8.435 ;
      RECT 102.95 8.235 103.41 8.405 ;
      RECT 102.915 4.025 103.235 4.26 ;
      RECT 102.915 4.055 103.405 4.225 ;
      RECT 102.915 3.69 103.105 4.26 ;
      RECT 102.33 3.655 102.62 3.885 ;
      RECT 102.33 3.69 103.105 3.86 ;
      RECT 102.39 2.175 102.56 3.885 ;
      RECT 102.33 2.175 102.625 2.405 ;
      RECT 101.96 4.025 102.25 4.255 ;
      RECT 101.96 4.055 102.42 4.225 ;
      RECT 102.025 2.95 102.19 4.255 ;
      RECT 100.54 2.915 100.83 3.145 ;
      RECT 100.54 2.95 102.19 3.12 ;
      RECT 100.6 2.175 100.77 3.145 ;
      RECT 100.54 2.175 100.83 2.405 ;
      RECT 100.54 10.055 100.83 10.285 ;
      RECT 100.6 9.315 100.77 10.285 ;
      RECT 100.6 9.405 102.19 9.575 ;
      RECT 102.02 8.205 102.19 9.575 ;
      RECT 100.54 9.315 100.83 9.545 ;
      RECT 101.96 8.205 102.25 8.435 ;
      RECT 101.96 8.235 102.42 8.405 ;
      RECT 100.97 3.26 101.32 3.61 ;
      RECT 100.8 3.315 101.32 3.485 ;
      RECT 100.995 8.94 101.32 9.265 ;
      RECT 100.97 8.945 101.32 9.175 ;
      RECT 100.8 8.975 101.32 9.145 ;
      RECT 100.195 3.66 100.515 3.98 ;
      RECT 100.17 3.655 100.46 3.885 ;
      RECT 99.88 3.69 100.515 3.86 ;
      RECT 99.995 3.685 100.515 3.86 ;
      RECT 100.195 8.565 100.515 8.89 ;
      RECT 100.17 8.575 100.515 8.805 ;
      RECT 99.995 8.605 100.515 8.775 ;
      RECT 95.94 5.085 96.26 5.345 ;
      RECT 96.975 5.1 97.265 5.33 ;
      RECT 95.94 5.145 97.265 5.285 ;
      RECT 96.975 7.14 97.265 7.37 ;
      RECT 95.6 7.11 95.92 7.37 ;
      RECT 97.05 6.83 97.19 7.37 ;
      RECT 95.69 6.83 95.83 7.37 ;
      RECT 95.69 6.83 97.19 6.97 ;
      RECT 96.62 4.065 96.94 4.325 ;
      RECT 96.345 4.125 96.94 4.265 ;
      RECT 96.295 7.805 96.94 8.05 ;
      RECT 96.62 7.775 96.94 8.05 ;
      RECT 92.555 7.82 92.845 8.05 ;
      RECT 93.56 7.775 93.88 8.035 ;
      RECT 92.555 7.865 94.47 8.005 ;
      RECT 94.33 7.51 94.47 8.005 ;
      RECT 93.555 7.835 93.885 8.005 ;
      RECT 94.33 7.51 96.34 7.65 ;
      RECT 96.2 7.14 96.34 7.65 ;
      RECT 96.125 7.14 96.415 7.37 ;
      RECT 95.94 6.105 96.26 6.365 ;
      RECT 93.795 6.12 94.085 6.35 ;
      RECT 93.795 6.165 96.26 6.305 ;
      RECT 95.26 5.085 95.58 5.345 ;
      RECT 92.895 5.1 93.185 5.33 ;
      RECT 92.895 5.145 95.58 5.285 ;
      RECT 94.92 7.79 95.24 8.05 ;
      RECT 94.92 7.865 95.515 8.005 ;
      RECT 94.92 4.405 95.24 4.665 ;
      RECT 94.645 4.465 95.24 4.605 ;
      RECT 94.245 7.125 94.89 7.37 ;
      RECT 94.57 7.11 94.89 7.37 ;
      RECT 94.24 4.065 94.56 4.325 ;
      RECT 93.965 4.125 94.56 4.265 ;
      RECT 93.9 4.745 94.22 5.005 ;
      RECT 91.025 4.76 91.315 4.99 ;
      RECT 91.025 4.805 94.22 4.945 ;
      RECT 93.48 4.085 93.62 4.945 ;
      RECT 93.405 4.085 93.695 4.315 ;
      RECT 93.56 3.555 93.88 3.815 ;
      RECT 93.56 3.57 94.065 3.8 ;
      RECT 93.47 3.615 94.065 3.755 ;
      RECT 92.895 4.085 93.185 4.315 ;
      RECT 92.29 4.13 93.185 4.27 ;
      RECT 92.29 3.725 92.43 4.27 ;
      RECT 92.2 3.725 92.52 3.985 ;
      RECT 91.52 4.065 91.84 4.325 ;
      RECT 91.245 4.125 91.84 4.265 ;
      RECT 91.52 6.105 91.84 6.365 ;
      RECT 91.245 6.165 91.84 6.305 ;
      RECT 89.285 8.86 89.575 9.175 ;
      RECT 89.115 8.975 89.575 9.145 ;
      RECT 89.265 8.86 89.605 9.14 ;
      RECT 88.855 10.055 89.145 10.285 ;
      RECT 88.915 9.285 89.085 10.285 ;
      RECT 88.82 9.285 89.19 9.655 ;
      RECT 86.1 10.055 86.395 10.285 ;
      RECT 86.16 8.575 86.33 10.285 ;
      RECT 86.16 8.945 86.49 9.27 ;
      RECT 86.1 8.575 86.39 8.805 ;
      RECT 85.11 10.055 85.405 10.285 ;
      RECT 85.17 8.575 85.34 10.285 ;
      RECT 85.11 8.575 85.4 8.805 ;
      RECT 85.11 8.61 85.96 8.77 ;
      RECT 85.795 8.205 85.96 8.77 ;
      RECT 85.11 8.605 85.505 8.77 ;
      RECT 85.73 8.205 86.02 8.435 ;
      RECT 85.73 8.235 86.19 8.405 ;
      RECT 85.695 4.025 86.015 4.26 ;
      RECT 85.695 4.055 86.185 4.225 ;
      RECT 85.695 3.69 85.885 4.26 ;
      RECT 85.11 3.655 85.4 3.885 ;
      RECT 85.11 3.69 85.885 3.86 ;
      RECT 85.17 2.175 85.34 3.885 ;
      RECT 85.11 2.175 85.405 2.405 ;
      RECT 84.74 4.025 85.03 4.255 ;
      RECT 84.74 4.055 85.2 4.225 ;
      RECT 84.805 2.95 84.97 4.255 ;
      RECT 83.32 2.915 83.61 3.145 ;
      RECT 83.32 2.95 84.97 3.12 ;
      RECT 83.38 2.175 83.55 3.145 ;
      RECT 83.32 2.175 83.61 2.405 ;
      RECT 83.32 10.055 83.61 10.285 ;
      RECT 83.38 9.315 83.55 10.285 ;
      RECT 83.38 9.405 84.97 9.575 ;
      RECT 84.8 8.205 84.97 9.575 ;
      RECT 83.32 9.315 83.61 9.545 ;
      RECT 84.74 8.205 85.03 8.435 ;
      RECT 84.74 8.235 85.2 8.405 ;
      RECT 83.75 3.26 84.1 3.61 ;
      RECT 83.58 3.315 84.1 3.485 ;
      RECT 83.775 8.94 84.1 9.265 ;
      RECT 83.75 8.945 84.1 9.175 ;
      RECT 83.58 8.975 84.1 9.145 ;
      RECT 82.975 3.66 83.295 3.98 ;
      RECT 82.95 3.655 83.24 3.885 ;
      RECT 82.66 3.69 83.295 3.86 ;
      RECT 82.775 3.685 83.295 3.86 ;
      RECT 82.975 8.565 83.295 8.89 ;
      RECT 82.95 8.575 83.295 8.805 ;
      RECT 82.775 8.605 83.295 8.775 ;
      RECT 78.72 5.085 79.04 5.345 ;
      RECT 79.755 5.1 80.045 5.33 ;
      RECT 78.72 5.145 80.045 5.285 ;
      RECT 79.755 7.14 80.045 7.37 ;
      RECT 78.38 7.11 78.7 7.37 ;
      RECT 79.83 6.83 79.97 7.37 ;
      RECT 78.47 6.83 78.61 7.37 ;
      RECT 78.47 6.83 79.97 6.97 ;
      RECT 79.4 4.065 79.72 4.325 ;
      RECT 79.125 4.125 79.72 4.265 ;
      RECT 79.075 7.805 79.72 8.05 ;
      RECT 79.4 7.775 79.72 8.05 ;
      RECT 75.335 7.82 75.625 8.05 ;
      RECT 76.34 7.775 76.66 8.035 ;
      RECT 75.335 7.865 77.25 8.005 ;
      RECT 77.11 7.51 77.25 8.005 ;
      RECT 76.335 7.835 76.665 8.005 ;
      RECT 77.11 7.51 79.12 7.65 ;
      RECT 78.98 7.14 79.12 7.65 ;
      RECT 78.905 7.14 79.195 7.37 ;
      RECT 78.72 6.105 79.04 6.365 ;
      RECT 76.575 6.12 76.865 6.35 ;
      RECT 76.575 6.165 79.04 6.305 ;
      RECT 78.04 5.085 78.36 5.345 ;
      RECT 75.675 5.1 75.965 5.33 ;
      RECT 75.675 5.145 78.36 5.285 ;
      RECT 77.7 7.79 78.02 8.05 ;
      RECT 77.7 7.865 78.295 8.005 ;
      RECT 77.7 4.405 78.02 4.665 ;
      RECT 77.425 4.465 78.02 4.605 ;
      RECT 77.025 7.125 77.67 7.37 ;
      RECT 77.35 7.11 77.67 7.37 ;
      RECT 77.02 4.065 77.34 4.325 ;
      RECT 76.745 4.125 77.34 4.265 ;
      RECT 76.68 4.745 77 5.005 ;
      RECT 73.805 4.76 74.095 4.99 ;
      RECT 73.805 4.805 77 4.945 ;
      RECT 76.26 4.085 76.4 4.945 ;
      RECT 76.185 4.085 76.475 4.315 ;
      RECT 76.34 3.555 76.66 3.815 ;
      RECT 76.34 3.57 76.845 3.8 ;
      RECT 76.25 3.615 76.845 3.755 ;
      RECT 75.675 4.085 75.965 4.315 ;
      RECT 75.07 4.13 75.965 4.27 ;
      RECT 75.07 3.725 75.21 4.27 ;
      RECT 74.98 3.725 75.3 3.985 ;
      RECT 74.3 4.065 74.62 4.325 ;
      RECT 74.025 4.125 74.62 4.265 ;
      RECT 74.3 6.105 74.62 6.365 ;
      RECT 74.025 6.165 74.62 6.305 ;
      RECT 72.065 8.86 72.355 9.175 ;
      RECT 71.895 8.975 72.355 9.145 ;
      RECT 72.045 8.86 72.385 9.14 ;
      RECT 71.635 10.055 71.925 10.285 ;
      RECT 71.695 9.285 71.865 10.285 ;
      RECT 71.6 9.285 71.97 9.655 ;
      RECT 68.88 10.055 69.175 10.285 ;
      RECT 68.94 8.575 69.11 10.285 ;
      RECT 68.94 8.945 69.27 9.27 ;
      RECT 68.88 8.575 69.17 8.805 ;
      RECT 67.89 10.055 68.185 10.285 ;
      RECT 67.95 8.575 68.12 10.285 ;
      RECT 67.89 8.575 68.18 8.805 ;
      RECT 67.89 8.61 68.74 8.77 ;
      RECT 68.575 8.205 68.74 8.77 ;
      RECT 67.89 8.605 68.285 8.77 ;
      RECT 68.51 8.205 68.8 8.435 ;
      RECT 68.51 8.235 68.97 8.405 ;
      RECT 68.475 4.025 68.795 4.26 ;
      RECT 68.475 4.055 68.965 4.225 ;
      RECT 68.475 3.69 68.665 4.26 ;
      RECT 67.89 3.655 68.18 3.885 ;
      RECT 67.89 3.69 68.665 3.86 ;
      RECT 67.95 2.175 68.12 3.885 ;
      RECT 67.89 2.175 68.185 2.405 ;
      RECT 67.52 4.025 67.81 4.255 ;
      RECT 67.52 4.055 67.98 4.225 ;
      RECT 67.585 2.95 67.75 4.255 ;
      RECT 66.1 2.915 66.39 3.145 ;
      RECT 66.1 2.95 67.75 3.12 ;
      RECT 66.16 2.175 66.33 3.145 ;
      RECT 66.1 2.175 66.39 2.405 ;
      RECT 66.1 10.055 66.39 10.285 ;
      RECT 66.16 9.315 66.33 10.285 ;
      RECT 66.16 9.405 67.75 9.575 ;
      RECT 67.58 8.205 67.75 9.575 ;
      RECT 66.1 9.315 66.39 9.545 ;
      RECT 67.52 8.205 67.81 8.435 ;
      RECT 67.52 8.235 67.98 8.405 ;
      RECT 66.53 3.26 66.88 3.61 ;
      RECT 66.36 3.315 66.88 3.485 ;
      RECT 66.555 8.94 66.88 9.265 ;
      RECT 66.53 8.945 66.88 9.175 ;
      RECT 66.36 8.975 66.88 9.145 ;
      RECT 65.755 3.66 66.075 3.98 ;
      RECT 65.73 3.655 66.02 3.885 ;
      RECT 65.44 3.69 66.075 3.86 ;
      RECT 65.555 3.685 66.075 3.86 ;
      RECT 65.755 8.565 66.075 8.89 ;
      RECT 65.73 8.575 66.075 8.805 ;
      RECT 65.555 8.605 66.075 8.775 ;
      RECT 61.5 5.085 61.82 5.345 ;
      RECT 62.535 5.1 62.825 5.33 ;
      RECT 61.5 5.145 62.825 5.285 ;
      RECT 62.535 7.14 62.825 7.37 ;
      RECT 61.16 7.11 61.48 7.37 ;
      RECT 62.61 6.83 62.75 7.37 ;
      RECT 61.25 6.83 61.39 7.37 ;
      RECT 61.25 6.83 62.75 6.97 ;
      RECT 62.18 4.065 62.5 4.325 ;
      RECT 61.905 4.125 62.5 4.265 ;
      RECT 61.855 7.805 62.5 8.05 ;
      RECT 62.18 7.775 62.5 8.05 ;
      RECT 58.115 7.82 58.405 8.05 ;
      RECT 59.12 7.775 59.44 8.035 ;
      RECT 58.115 7.865 60.03 8.005 ;
      RECT 59.89 7.51 60.03 8.005 ;
      RECT 59.115 7.835 59.445 8.005 ;
      RECT 59.89 7.51 61.9 7.65 ;
      RECT 61.76 7.14 61.9 7.65 ;
      RECT 61.685 7.14 61.975 7.37 ;
      RECT 61.5 6.105 61.82 6.365 ;
      RECT 59.355 6.12 59.645 6.35 ;
      RECT 59.355 6.165 61.82 6.305 ;
      RECT 60.82 5.085 61.14 5.345 ;
      RECT 58.455 5.1 58.745 5.33 ;
      RECT 58.455 5.145 61.14 5.285 ;
      RECT 60.48 7.79 60.8 8.05 ;
      RECT 60.48 7.865 61.075 8.005 ;
      RECT 60.48 4.405 60.8 4.665 ;
      RECT 60.205 4.465 60.8 4.605 ;
      RECT 59.805 7.125 60.45 7.37 ;
      RECT 60.13 7.11 60.45 7.37 ;
      RECT 59.8 4.065 60.12 4.325 ;
      RECT 59.525 4.125 60.12 4.265 ;
      RECT 59.46 4.745 59.78 5.005 ;
      RECT 56.585 4.76 56.875 4.99 ;
      RECT 56.585 4.805 59.78 4.945 ;
      RECT 59.04 4.085 59.18 4.945 ;
      RECT 58.965 4.085 59.255 4.315 ;
      RECT 59.12 3.555 59.44 3.815 ;
      RECT 59.12 3.57 59.625 3.8 ;
      RECT 59.03 3.615 59.625 3.755 ;
      RECT 58.455 4.085 58.745 4.315 ;
      RECT 57.85 4.13 58.745 4.27 ;
      RECT 57.85 3.725 57.99 4.27 ;
      RECT 57.76 3.725 58.08 3.985 ;
      RECT 57.08 4.065 57.4 4.325 ;
      RECT 56.805 4.125 57.4 4.265 ;
      RECT 57.08 6.105 57.4 6.365 ;
      RECT 56.805 6.165 57.4 6.305 ;
      RECT 54.845 8.86 55.135 9.175 ;
      RECT 54.675 8.975 55.135 9.145 ;
      RECT 54.825 8.86 55.165 9.14 ;
      RECT 54.415 10.055 54.705 10.285 ;
      RECT 54.475 9.285 54.645 10.285 ;
      RECT 54.38 9.285 54.75 9.655 ;
      RECT 51.66 10.055 51.955 10.285 ;
      RECT 51.72 8.575 51.89 10.285 ;
      RECT 51.72 8.945 52.05 9.27 ;
      RECT 51.66 8.575 51.95 8.805 ;
      RECT 50.67 10.055 50.965 10.285 ;
      RECT 50.73 8.575 50.9 10.285 ;
      RECT 50.67 8.575 50.96 8.805 ;
      RECT 50.67 8.61 51.52 8.77 ;
      RECT 51.355 8.205 51.52 8.77 ;
      RECT 50.67 8.605 51.065 8.77 ;
      RECT 51.29 8.205 51.58 8.435 ;
      RECT 51.29 8.235 51.75 8.405 ;
      RECT 51.255 4.025 51.575 4.26 ;
      RECT 51.255 4.055 51.745 4.225 ;
      RECT 51.255 3.69 51.445 4.26 ;
      RECT 50.67 3.655 50.96 3.885 ;
      RECT 50.67 3.69 51.445 3.86 ;
      RECT 50.73 2.175 50.9 3.885 ;
      RECT 50.67 2.175 50.965 2.405 ;
      RECT 50.3 4.025 50.59 4.255 ;
      RECT 50.3 4.055 50.76 4.225 ;
      RECT 50.365 2.95 50.53 4.255 ;
      RECT 48.88 2.915 49.17 3.145 ;
      RECT 48.88 2.95 50.53 3.12 ;
      RECT 48.94 2.175 49.11 3.145 ;
      RECT 48.88 2.175 49.17 2.405 ;
      RECT 48.88 10.055 49.17 10.285 ;
      RECT 48.94 9.315 49.11 10.285 ;
      RECT 48.94 9.405 50.53 9.575 ;
      RECT 50.36 8.205 50.53 9.575 ;
      RECT 48.88 9.315 49.17 9.545 ;
      RECT 50.3 8.205 50.59 8.435 ;
      RECT 50.3 8.235 50.76 8.405 ;
      RECT 49.31 3.26 49.66 3.61 ;
      RECT 49.14 3.315 49.66 3.485 ;
      RECT 49.335 8.94 49.66 9.265 ;
      RECT 49.31 8.945 49.66 9.175 ;
      RECT 49.14 8.975 49.66 9.145 ;
      RECT 48.535 3.66 48.855 3.98 ;
      RECT 48.51 3.655 48.8 3.885 ;
      RECT 48.22 3.69 48.855 3.86 ;
      RECT 48.335 3.685 48.855 3.86 ;
      RECT 48.535 8.565 48.855 8.89 ;
      RECT 48.51 8.575 48.855 8.805 ;
      RECT 48.335 8.605 48.855 8.775 ;
      RECT 44.28 5.085 44.6 5.345 ;
      RECT 45.315 5.1 45.605 5.33 ;
      RECT 44.28 5.145 45.605 5.285 ;
      RECT 45.315 7.14 45.605 7.37 ;
      RECT 43.94 7.11 44.26 7.37 ;
      RECT 45.39 6.83 45.53 7.37 ;
      RECT 44.03 6.83 44.17 7.37 ;
      RECT 44.03 6.83 45.53 6.97 ;
      RECT 44.96 4.065 45.28 4.325 ;
      RECT 44.685 4.125 45.28 4.265 ;
      RECT 44.635 7.805 45.28 8.05 ;
      RECT 44.96 7.775 45.28 8.05 ;
      RECT 40.895 7.82 41.185 8.05 ;
      RECT 41.9 7.775 42.22 8.035 ;
      RECT 40.895 7.865 42.81 8.005 ;
      RECT 42.67 7.51 42.81 8.005 ;
      RECT 41.895 7.835 42.225 8.005 ;
      RECT 42.67 7.51 44.68 7.65 ;
      RECT 44.54 7.14 44.68 7.65 ;
      RECT 44.465 7.14 44.755 7.37 ;
      RECT 44.28 6.105 44.6 6.365 ;
      RECT 42.135 6.12 42.425 6.35 ;
      RECT 42.135 6.165 44.6 6.305 ;
      RECT 43.6 5.085 43.92 5.345 ;
      RECT 41.235 5.1 41.525 5.33 ;
      RECT 41.235 5.145 43.92 5.285 ;
      RECT 43.26 7.79 43.58 8.05 ;
      RECT 43.26 7.865 43.855 8.005 ;
      RECT 43.26 4.405 43.58 4.665 ;
      RECT 42.985 4.465 43.58 4.605 ;
      RECT 42.585 7.125 43.23 7.37 ;
      RECT 42.91 7.11 43.23 7.37 ;
      RECT 42.58 4.065 42.9 4.325 ;
      RECT 42.305 4.125 42.9 4.265 ;
      RECT 42.24 4.745 42.56 5.005 ;
      RECT 39.365 4.76 39.655 4.99 ;
      RECT 39.365 4.805 42.56 4.945 ;
      RECT 41.82 4.085 41.96 4.945 ;
      RECT 41.745 4.085 42.035 4.315 ;
      RECT 41.9 3.555 42.22 3.815 ;
      RECT 41.9 3.57 42.405 3.8 ;
      RECT 41.81 3.615 42.405 3.755 ;
      RECT 41.235 4.085 41.525 4.315 ;
      RECT 40.63 4.13 41.525 4.27 ;
      RECT 40.63 3.725 40.77 4.27 ;
      RECT 40.54 3.725 40.86 3.985 ;
      RECT 39.86 4.065 40.18 4.325 ;
      RECT 39.585 4.125 40.18 4.265 ;
      RECT 39.86 6.105 40.18 6.365 ;
      RECT 39.585 6.165 40.18 6.305 ;
      RECT 37.625 8.86 37.915 9.175 ;
      RECT 37.455 8.975 37.915 9.145 ;
      RECT 37.605 8.86 37.945 9.14 ;
      RECT 37.195 10.055 37.485 10.285 ;
      RECT 37.255 9.285 37.425 10.285 ;
      RECT 37.16 9.285 37.53 9.655 ;
      RECT 34.44 10.055 34.735 10.285 ;
      RECT 34.5 8.575 34.67 10.285 ;
      RECT 34.5 8.945 34.83 9.27 ;
      RECT 34.44 8.575 34.73 8.805 ;
      RECT 33.45 10.055 33.745 10.285 ;
      RECT 33.51 8.575 33.68 10.285 ;
      RECT 33.45 8.575 33.74 8.805 ;
      RECT 33.45 8.61 34.3 8.77 ;
      RECT 34.135 8.205 34.3 8.77 ;
      RECT 33.45 8.605 33.845 8.77 ;
      RECT 34.07 8.205 34.36 8.435 ;
      RECT 34.07 8.235 34.53 8.405 ;
      RECT 34.035 4.025 34.355 4.26 ;
      RECT 34.035 4.055 34.525 4.225 ;
      RECT 34.035 3.69 34.225 4.26 ;
      RECT 33.45 3.655 33.74 3.885 ;
      RECT 33.45 3.69 34.225 3.86 ;
      RECT 33.51 2.175 33.68 3.885 ;
      RECT 33.45 2.175 33.745 2.405 ;
      RECT 33.08 4.025 33.37 4.255 ;
      RECT 33.08 4.055 33.54 4.225 ;
      RECT 33.145 2.95 33.31 4.255 ;
      RECT 31.66 2.915 31.95 3.145 ;
      RECT 31.66 2.95 33.31 3.12 ;
      RECT 31.72 2.175 31.89 3.145 ;
      RECT 31.66 2.175 31.95 2.405 ;
      RECT 31.66 10.055 31.95 10.285 ;
      RECT 31.72 9.315 31.89 10.285 ;
      RECT 31.72 9.405 33.31 9.575 ;
      RECT 33.14 8.205 33.31 9.575 ;
      RECT 31.66 9.315 31.95 9.545 ;
      RECT 33.08 8.205 33.37 8.435 ;
      RECT 33.08 8.235 33.54 8.405 ;
      RECT 32.09 3.26 32.44 3.61 ;
      RECT 31.92 3.315 32.44 3.485 ;
      RECT 32.115 8.94 32.44 9.265 ;
      RECT 32.09 8.945 32.44 9.175 ;
      RECT 31.92 8.975 32.44 9.145 ;
      RECT 31.315 3.66 31.635 3.98 ;
      RECT 31.29 3.655 31.58 3.885 ;
      RECT 31 3.69 31.635 3.86 ;
      RECT 31.115 3.685 31.635 3.86 ;
      RECT 31.315 8.565 31.635 8.89 ;
      RECT 31.29 8.575 31.635 8.805 ;
      RECT 31.115 8.605 31.635 8.775 ;
      RECT 27.06 5.085 27.38 5.345 ;
      RECT 28.095 5.1 28.385 5.33 ;
      RECT 27.06 5.145 28.385 5.285 ;
      RECT 28.095 7.14 28.385 7.37 ;
      RECT 26.72 7.11 27.04 7.37 ;
      RECT 28.17 6.83 28.31 7.37 ;
      RECT 26.81 6.83 26.95 7.37 ;
      RECT 26.81 6.83 28.31 6.97 ;
      RECT 27.74 4.065 28.06 4.325 ;
      RECT 27.465 4.125 28.06 4.265 ;
      RECT 27.415 7.805 28.06 8.05 ;
      RECT 27.74 7.775 28.06 8.05 ;
      RECT 23.675 7.82 23.965 8.05 ;
      RECT 24.68 7.775 25 8.035 ;
      RECT 23.675 7.865 25.59 8.005 ;
      RECT 25.45 7.51 25.59 8.005 ;
      RECT 24.675 7.835 25.005 8.005 ;
      RECT 25.45 7.51 27.46 7.65 ;
      RECT 27.32 7.14 27.46 7.65 ;
      RECT 27.245 7.14 27.535 7.37 ;
      RECT 27.06 6.105 27.38 6.365 ;
      RECT 24.915 6.12 25.205 6.35 ;
      RECT 24.915 6.165 27.38 6.305 ;
      RECT 26.38 5.085 26.7 5.345 ;
      RECT 24.015 5.1 24.305 5.33 ;
      RECT 24.015 5.145 26.7 5.285 ;
      RECT 26.04 7.79 26.36 8.05 ;
      RECT 26.04 7.865 26.635 8.005 ;
      RECT 26.04 4.405 26.36 4.665 ;
      RECT 25.765 4.465 26.36 4.605 ;
      RECT 25.365 7.125 26.01 7.37 ;
      RECT 25.69 7.11 26.01 7.37 ;
      RECT 25.36 4.065 25.68 4.325 ;
      RECT 25.085 4.125 25.68 4.265 ;
      RECT 25.02 4.745 25.34 5.005 ;
      RECT 22.145 4.76 22.435 4.99 ;
      RECT 22.145 4.805 25.34 4.945 ;
      RECT 24.6 4.085 24.74 4.945 ;
      RECT 24.525 4.085 24.815 4.315 ;
      RECT 24.68 3.555 25 3.815 ;
      RECT 24.68 3.57 25.185 3.8 ;
      RECT 24.59 3.615 25.185 3.755 ;
      RECT 24.015 4.085 24.305 4.315 ;
      RECT 23.41 4.13 24.305 4.27 ;
      RECT 23.41 3.725 23.55 4.27 ;
      RECT 23.32 3.725 23.64 3.985 ;
      RECT 22.64 4.065 22.96 4.325 ;
      RECT 22.365 4.125 22.96 4.265 ;
      RECT 22.64 6.105 22.96 6.365 ;
      RECT 22.365 6.165 22.96 6.305 ;
      RECT 20.405 8.86 20.695 9.175 ;
      RECT 20.235 8.975 20.695 9.145 ;
      RECT 20.385 8.86 20.725 9.14 ;
      RECT 19.975 10.055 20.265 10.285 ;
      RECT 20.035 9.285 20.205 10.285 ;
      RECT 19.94 9.285 20.31 9.655 ;
      RECT 16.565 10.055 16.855 10.285 ;
      RECT 16.625 9.31 16.795 10.285 ;
      RECT 16.535 9.31 16.875 9.59 ;
      RECT 16.16 8.57 16.5 8.85 ;
      RECT 16.02 8.605 16.5 8.775 ;
      RECT 103.295 7.245 103.645 7.535 ;
      RECT 98.525 3.29 98.85 3.615 ;
      RECT 86.075 7.245 86.425 7.535 ;
      RECT 81.305 3.29 81.63 3.615 ;
      RECT 68.855 7.245 69.205 7.535 ;
      RECT 64.085 3.29 64.41 3.615 ;
      RECT 51.635 7.245 51.985 7.535 ;
      RECT 46.865 3.29 47.19 3.615 ;
      RECT 34.415 7.245 34.765 7.535 ;
      RECT 29.645 3.29 29.97 3.615 ;
    LAYER mcon ;
      RECT 103.385 7.305 103.555 7.475 ;
      RECT 103.38 8.605 103.55 8.775 ;
      RECT 103.38 10.085 103.55 10.255 ;
      RECT 103.01 8.235 103.18 8.405 ;
      RECT 103.005 4.055 103.175 4.225 ;
      RECT 102.39 2.205 102.56 2.375 ;
      RECT 102.39 3.685 102.56 3.855 ;
      RECT 102.39 8.605 102.56 8.775 ;
      RECT 102.39 10.085 102.56 10.255 ;
      RECT 102.02 4.055 102.19 4.225 ;
      RECT 102.02 8.235 102.19 8.405 ;
      RECT 101.03 3.315 101.2 3.485 ;
      RECT 101.03 8.975 101.2 9.145 ;
      RECT 100.6 2.205 100.77 2.375 ;
      RECT 100.6 2.945 100.77 3.115 ;
      RECT 100.6 9.345 100.77 9.515 ;
      RECT 100.6 10.085 100.77 10.255 ;
      RECT 100.23 3.685 100.4 3.855 ;
      RECT 100.23 8.605 100.4 8.775 ;
      RECT 97.035 5.13 97.205 5.3 ;
      RECT 97.035 7.17 97.205 7.34 ;
      RECT 96.695 4.11 96.865 4.28 ;
      RECT 96.355 7.85 96.525 8.02 ;
      RECT 96.185 7.17 96.355 7.34 ;
      RECT 95.675 7.17 95.845 7.34 ;
      RECT 94.995 4.45 95.165 4.62 ;
      RECT 94.995 7.85 95.165 8.02 ;
      RECT 94.315 4.11 94.485 4.28 ;
      RECT 94.305 7.17 94.475 7.34 ;
      RECT 93.855 6.15 94.025 6.32 ;
      RECT 93.835 3.6 94.005 3.77 ;
      RECT 93.465 4.115 93.635 4.285 ;
      RECT 92.955 4.115 93.125 4.285 ;
      RECT 92.955 5.13 93.125 5.3 ;
      RECT 92.615 7.85 92.785 8.02 ;
      RECT 91.595 4.11 91.765 4.28 ;
      RECT 91.595 6.15 91.765 6.32 ;
      RECT 91.085 4.79 91.255 4.96 ;
      RECT 89.345 8.975 89.515 9.145 ;
      RECT 88.915 9.345 89.085 9.515 ;
      RECT 88.915 10.085 89.085 10.255 ;
      RECT 86.165 7.305 86.335 7.475 ;
      RECT 86.16 8.605 86.33 8.775 ;
      RECT 86.16 10.085 86.33 10.255 ;
      RECT 85.79 8.235 85.96 8.405 ;
      RECT 85.785 4.055 85.955 4.225 ;
      RECT 85.17 2.205 85.34 2.375 ;
      RECT 85.17 3.685 85.34 3.855 ;
      RECT 85.17 8.605 85.34 8.775 ;
      RECT 85.17 10.085 85.34 10.255 ;
      RECT 84.8 4.055 84.97 4.225 ;
      RECT 84.8 8.235 84.97 8.405 ;
      RECT 83.81 3.315 83.98 3.485 ;
      RECT 83.81 8.975 83.98 9.145 ;
      RECT 83.38 2.205 83.55 2.375 ;
      RECT 83.38 2.945 83.55 3.115 ;
      RECT 83.38 9.345 83.55 9.515 ;
      RECT 83.38 10.085 83.55 10.255 ;
      RECT 83.01 3.685 83.18 3.855 ;
      RECT 83.01 8.605 83.18 8.775 ;
      RECT 79.815 5.13 79.985 5.3 ;
      RECT 79.815 7.17 79.985 7.34 ;
      RECT 79.475 4.11 79.645 4.28 ;
      RECT 79.135 7.85 79.305 8.02 ;
      RECT 78.965 7.17 79.135 7.34 ;
      RECT 78.455 7.17 78.625 7.34 ;
      RECT 77.775 4.45 77.945 4.62 ;
      RECT 77.775 7.85 77.945 8.02 ;
      RECT 77.095 4.11 77.265 4.28 ;
      RECT 77.085 7.17 77.255 7.34 ;
      RECT 76.635 6.15 76.805 6.32 ;
      RECT 76.615 3.6 76.785 3.77 ;
      RECT 76.245 4.115 76.415 4.285 ;
      RECT 75.735 4.115 75.905 4.285 ;
      RECT 75.735 5.13 75.905 5.3 ;
      RECT 75.395 7.85 75.565 8.02 ;
      RECT 74.375 4.11 74.545 4.28 ;
      RECT 74.375 6.15 74.545 6.32 ;
      RECT 73.865 4.79 74.035 4.96 ;
      RECT 72.125 8.975 72.295 9.145 ;
      RECT 71.695 9.345 71.865 9.515 ;
      RECT 71.695 10.085 71.865 10.255 ;
      RECT 68.945 7.305 69.115 7.475 ;
      RECT 68.94 8.605 69.11 8.775 ;
      RECT 68.94 10.085 69.11 10.255 ;
      RECT 68.57 8.235 68.74 8.405 ;
      RECT 68.565 4.055 68.735 4.225 ;
      RECT 67.95 2.205 68.12 2.375 ;
      RECT 67.95 3.685 68.12 3.855 ;
      RECT 67.95 8.605 68.12 8.775 ;
      RECT 67.95 10.085 68.12 10.255 ;
      RECT 67.58 4.055 67.75 4.225 ;
      RECT 67.58 8.235 67.75 8.405 ;
      RECT 66.59 3.315 66.76 3.485 ;
      RECT 66.59 8.975 66.76 9.145 ;
      RECT 66.16 2.205 66.33 2.375 ;
      RECT 66.16 2.945 66.33 3.115 ;
      RECT 66.16 9.345 66.33 9.515 ;
      RECT 66.16 10.085 66.33 10.255 ;
      RECT 65.79 3.685 65.96 3.855 ;
      RECT 65.79 8.605 65.96 8.775 ;
      RECT 62.595 5.13 62.765 5.3 ;
      RECT 62.595 7.17 62.765 7.34 ;
      RECT 62.255 4.11 62.425 4.28 ;
      RECT 61.915 7.85 62.085 8.02 ;
      RECT 61.745 7.17 61.915 7.34 ;
      RECT 61.235 7.17 61.405 7.34 ;
      RECT 60.555 4.45 60.725 4.62 ;
      RECT 60.555 7.85 60.725 8.02 ;
      RECT 59.875 4.11 60.045 4.28 ;
      RECT 59.865 7.17 60.035 7.34 ;
      RECT 59.415 6.15 59.585 6.32 ;
      RECT 59.395 3.6 59.565 3.77 ;
      RECT 59.025 4.115 59.195 4.285 ;
      RECT 58.515 4.115 58.685 4.285 ;
      RECT 58.515 5.13 58.685 5.3 ;
      RECT 58.175 7.85 58.345 8.02 ;
      RECT 57.155 4.11 57.325 4.28 ;
      RECT 57.155 6.15 57.325 6.32 ;
      RECT 56.645 4.79 56.815 4.96 ;
      RECT 54.905 8.975 55.075 9.145 ;
      RECT 54.475 9.345 54.645 9.515 ;
      RECT 54.475 10.085 54.645 10.255 ;
      RECT 51.725 7.305 51.895 7.475 ;
      RECT 51.72 8.605 51.89 8.775 ;
      RECT 51.72 10.085 51.89 10.255 ;
      RECT 51.35 8.235 51.52 8.405 ;
      RECT 51.345 4.055 51.515 4.225 ;
      RECT 50.73 2.205 50.9 2.375 ;
      RECT 50.73 3.685 50.9 3.855 ;
      RECT 50.73 8.605 50.9 8.775 ;
      RECT 50.73 10.085 50.9 10.255 ;
      RECT 50.36 4.055 50.53 4.225 ;
      RECT 50.36 8.235 50.53 8.405 ;
      RECT 49.37 3.315 49.54 3.485 ;
      RECT 49.37 8.975 49.54 9.145 ;
      RECT 48.94 2.205 49.11 2.375 ;
      RECT 48.94 2.945 49.11 3.115 ;
      RECT 48.94 9.345 49.11 9.515 ;
      RECT 48.94 10.085 49.11 10.255 ;
      RECT 48.57 3.685 48.74 3.855 ;
      RECT 48.57 8.605 48.74 8.775 ;
      RECT 45.375 5.13 45.545 5.3 ;
      RECT 45.375 7.17 45.545 7.34 ;
      RECT 45.035 4.11 45.205 4.28 ;
      RECT 44.695 7.85 44.865 8.02 ;
      RECT 44.525 7.17 44.695 7.34 ;
      RECT 44.015 7.17 44.185 7.34 ;
      RECT 43.335 4.45 43.505 4.62 ;
      RECT 43.335 7.85 43.505 8.02 ;
      RECT 42.655 4.11 42.825 4.28 ;
      RECT 42.645 7.17 42.815 7.34 ;
      RECT 42.195 6.15 42.365 6.32 ;
      RECT 42.175 3.6 42.345 3.77 ;
      RECT 41.805 4.115 41.975 4.285 ;
      RECT 41.295 4.115 41.465 4.285 ;
      RECT 41.295 5.13 41.465 5.3 ;
      RECT 40.955 7.85 41.125 8.02 ;
      RECT 39.935 4.11 40.105 4.28 ;
      RECT 39.935 6.15 40.105 6.32 ;
      RECT 39.425 4.79 39.595 4.96 ;
      RECT 37.685 8.975 37.855 9.145 ;
      RECT 37.255 9.345 37.425 9.515 ;
      RECT 37.255 10.085 37.425 10.255 ;
      RECT 34.505 7.305 34.675 7.475 ;
      RECT 34.5 8.605 34.67 8.775 ;
      RECT 34.5 10.085 34.67 10.255 ;
      RECT 34.13 8.235 34.3 8.405 ;
      RECT 34.125 4.055 34.295 4.225 ;
      RECT 33.51 2.205 33.68 2.375 ;
      RECT 33.51 3.685 33.68 3.855 ;
      RECT 33.51 8.605 33.68 8.775 ;
      RECT 33.51 10.085 33.68 10.255 ;
      RECT 33.14 4.055 33.31 4.225 ;
      RECT 33.14 8.235 33.31 8.405 ;
      RECT 32.15 3.315 32.32 3.485 ;
      RECT 32.15 8.975 32.32 9.145 ;
      RECT 31.72 2.205 31.89 2.375 ;
      RECT 31.72 2.945 31.89 3.115 ;
      RECT 31.72 9.345 31.89 9.515 ;
      RECT 31.72 10.085 31.89 10.255 ;
      RECT 31.35 3.685 31.52 3.855 ;
      RECT 31.35 8.605 31.52 8.775 ;
      RECT 28.155 5.13 28.325 5.3 ;
      RECT 28.155 7.17 28.325 7.34 ;
      RECT 27.815 4.11 27.985 4.28 ;
      RECT 27.475 7.85 27.645 8.02 ;
      RECT 27.305 7.17 27.475 7.34 ;
      RECT 26.795 7.17 26.965 7.34 ;
      RECT 26.115 4.45 26.285 4.62 ;
      RECT 26.115 7.85 26.285 8.02 ;
      RECT 25.435 4.11 25.605 4.28 ;
      RECT 25.425 7.17 25.595 7.34 ;
      RECT 24.975 6.15 25.145 6.32 ;
      RECT 24.955 3.6 25.125 3.77 ;
      RECT 24.585 4.115 24.755 4.285 ;
      RECT 24.075 4.115 24.245 4.285 ;
      RECT 24.075 5.13 24.245 5.3 ;
      RECT 23.735 7.85 23.905 8.02 ;
      RECT 22.715 4.11 22.885 4.28 ;
      RECT 22.715 6.15 22.885 6.32 ;
      RECT 22.205 4.79 22.375 4.96 ;
      RECT 20.465 8.975 20.635 9.145 ;
      RECT 20.035 9.345 20.205 9.515 ;
      RECT 20.035 10.085 20.205 10.255 ;
      RECT 16.625 9.345 16.795 9.515 ;
      RECT 16.625 10.085 16.795 10.255 ;
      RECT 16.255 8.605 16.425 8.775 ;
    LAYER li1 ;
      RECT 103.38 7.305 103.55 8.775 ;
      RECT 103.38 7.305 103.555 8.565 ;
      RECT 103.01 9.255 103.48 9.425 ;
      RECT 103.01 8.235 103.18 9.425 ;
      RECT 103.005 3.035 103.175 4.225 ;
      RECT 103.005 3.035 103.475 3.205 ;
      RECT 102.39 3.895 102.565 5.155 ;
      RECT 102.39 3.685 102.56 5.155 ;
      RECT 102.39 7.305 102.56 8.775 ;
      RECT 102.39 7.305 102.565 8.565 ;
      RECT 102.02 3.035 102.19 4.225 ;
      RECT 102.02 3.035 102.49 3.205 ;
      RECT 102.02 9.255 102.49 9.425 ;
      RECT 102.02 8.235 102.19 9.425 ;
      RECT 101.03 4.015 101.205 5.155 ;
      RECT 101.03 1.865 101.2 5.155 ;
      RECT 101.03 1.865 101.205 2.415 ;
      RECT 101.03 10.045 101.205 10.595 ;
      RECT 101.03 7.305 101.2 10.595 ;
      RECT 101.03 7.305 101.205 8.445 ;
      RECT 100.6 3.895 100.775 5.155 ;
      RECT 100.6 2.945 100.77 5.155 ;
      RECT 100.6 7.305 100.77 9.515 ;
      RECT 100.6 7.305 100.775 8.565 ;
      RECT 100.17 3.925 100.34 5.155 ;
      RECT 100.23 2.145 100.4 4.095 ;
      RECT 100.17 1.865 100.34 2.315 ;
      RECT 100.17 10.145 100.34 10.595 ;
      RECT 100.23 8.365 100.4 10.315 ;
      RECT 100.17 7.305 100.34 8.535 ;
      RECT 99.645 3.895 99.82 5.155 ;
      RECT 99.645 1.865 99.815 5.155 ;
      RECT 99.645 3.365 100.055 3.695 ;
      RECT 99.645 2.525 100.055 2.855 ;
      RECT 99.645 1.865 99.82 2.355 ;
      RECT 99.645 10.105 99.82 10.595 ;
      RECT 99.645 7.305 99.815 10.595 ;
      RECT 99.645 9.605 100.055 9.935 ;
      RECT 99.645 8.765 100.055 9.095 ;
      RECT 99.645 7.305 99.82 8.565 ;
      RECT 97.385 4.79 97.765 5.47 ;
      RECT 97.595 3.66 97.765 5.47 ;
      RECT 95.515 3.66 95.745 4.33 ;
      RECT 95.515 3.66 97.765 3.83 ;
      RECT 97.045 3.34 97.215 3.83 ;
      RECT 97.035 4.45 97.205 5.3 ;
      RECT 96.12 4.45 97.425 4.62 ;
      RECT 97.18 4 97.425 4.62 ;
      RECT 96.12 4.08 96.29 4.62 ;
      RECT 95.915 4.08 96.29 4.25 ;
      RECT 96.095 7.56 96.79 8.19 ;
      RECT 96.62 5.98 96.79 8.19 ;
      RECT 96.525 5.98 96.855 6.96 ;
      RECT 96.125 4.79 96.455 5.47 ;
      RECT 95.215 4.79 95.615 5.47 ;
      RECT 95.215 4.79 96.455 4.96 ;
      RECT 94.715 4.37 95.035 5.47 ;
      RECT 94.715 4.37 95.165 4.62 ;
      RECT 94.715 4.37 95.345 4.54 ;
      RECT 95.175 3.32 95.345 4.54 ;
      RECT 95.175 3.32 96.13 3.49 ;
      RECT 94.715 7.56 95.41 8.19 ;
      RECT 95.24 5.98 95.41 8.19 ;
      RECT 95.145 5.98 95.475 6.96 ;
      RECT 94.735 7.12 95.07 7.37 ;
      RECT 94.19 7.12 94.525 7.37 ;
      RECT 94.19 7.17 95.07 7.34 ;
      RECT 93.85 7.56 94.545 8.19 ;
      RECT 93.85 5.98 94.02 8.19 ;
      RECT 93.785 5.98 94.115 6.96 ;
      RECT 93.345 4.5 93.675 5.455 ;
      RECT 93.345 4.5 94.025 4.67 ;
      RECT 93.855 3.26 94.025 4.67 ;
      RECT 93.765 3.26 94.095 3.9 ;
      RECT 92.825 4.5 93.155 5.455 ;
      RECT 92.475 4.5 93.155 4.67 ;
      RECT 92.475 3.26 92.645 4.67 ;
      RECT 92.405 3.26 92.735 3.9 ;
      RECT 92.615 7.17 92.785 8.02 ;
      RECT 91.89 7.12 92.225 7.37 ;
      RECT 91.89 7.17 92.785 7.34 ;
      RECT 91.955 4.08 92.305 4.33 ;
      RECT 91.435 4.08 91.765 4.33 ;
      RECT 91.435 4.11 92.305 4.28 ;
      RECT 91.55 7.56 92.245 8.19 ;
      RECT 91.55 5.98 91.72 8.19 ;
      RECT 91.485 5.98 91.815 6.96 ;
      RECT 91.015 4.49 91.345 5.47 ;
      RECT 91.015 3.26 91.265 5.47 ;
      RECT 91.015 3.26 91.345 3.89 ;
      RECT 89.345 10.045 89.52 10.595 ;
      RECT 89.345 7.305 89.515 10.595 ;
      RECT 89.345 7.305 89.52 8.445 ;
      RECT 88.915 7.305 89.085 9.515 ;
      RECT 88.915 7.305 89.09 8.565 ;
      RECT 87.96 10.105 88.135 10.595 ;
      RECT 87.96 7.305 88.13 10.595 ;
      RECT 87.96 9.605 88.37 9.935 ;
      RECT 87.96 8.765 88.37 9.095 ;
      RECT 87.96 7.305 88.135 8.565 ;
      RECT 86.16 7.305 86.33 8.775 ;
      RECT 86.16 7.305 86.335 8.565 ;
      RECT 85.79 9.255 86.26 9.425 ;
      RECT 85.79 8.235 85.96 9.425 ;
      RECT 85.785 3.035 85.955 4.225 ;
      RECT 85.785 3.035 86.255 3.205 ;
      RECT 85.17 3.895 85.345 5.155 ;
      RECT 85.17 3.685 85.34 5.155 ;
      RECT 85.17 7.305 85.34 8.775 ;
      RECT 85.17 7.305 85.345 8.565 ;
      RECT 84.8 3.035 84.97 4.225 ;
      RECT 84.8 3.035 85.27 3.205 ;
      RECT 84.8 9.255 85.27 9.425 ;
      RECT 84.8 8.235 84.97 9.425 ;
      RECT 83.81 4.015 83.985 5.155 ;
      RECT 83.81 1.865 83.98 5.155 ;
      RECT 83.81 1.865 83.985 2.415 ;
      RECT 83.81 10.045 83.985 10.595 ;
      RECT 83.81 7.305 83.98 10.595 ;
      RECT 83.81 7.305 83.985 8.445 ;
      RECT 83.38 3.895 83.555 5.155 ;
      RECT 83.38 2.945 83.55 5.155 ;
      RECT 83.38 7.305 83.55 9.515 ;
      RECT 83.38 7.305 83.555 8.565 ;
      RECT 82.95 3.925 83.12 5.155 ;
      RECT 83.01 2.145 83.18 4.095 ;
      RECT 82.95 1.865 83.12 2.315 ;
      RECT 82.95 10.145 83.12 10.595 ;
      RECT 83.01 8.365 83.18 10.315 ;
      RECT 82.95 7.305 83.12 8.535 ;
      RECT 82.425 3.895 82.6 5.155 ;
      RECT 82.425 1.865 82.595 5.155 ;
      RECT 82.425 3.365 82.835 3.695 ;
      RECT 82.425 2.525 82.835 2.855 ;
      RECT 82.425 1.865 82.6 2.355 ;
      RECT 82.425 10.105 82.6 10.595 ;
      RECT 82.425 7.305 82.595 10.595 ;
      RECT 82.425 9.605 82.835 9.935 ;
      RECT 82.425 8.765 82.835 9.095 ;
      RECT 82.425 7.305 82.6 8.565 ;
      RECT 80.165 4.79 80.545 5.47 ;
      RECT 80.375 3.66 80.545 5.47 ;
      RECT 78.295 3.66 78.525 4.33 ;
      RECT 78.295 3.66 80.545 3.83 ;
      RECT 79.825 3.34 79.995 3.83 ;
      RECT 79.815 4.45 79.985 5.3 ;
      RECT 78.9 4.45 80.205 4.62 ;
      RECT 79.96 4 80.205 4.62 ;
      RECT 78.9 4.08 79.07 4.62 ;
      RECT 78.695 4.08 79.07 4.25 ;
      RECT 78.875 7.56 79.57 8.19 ;
      RECT 79.4 5.98 79.57 8.19 ;
      RECT 79.305 5.98 79.635 6.96 ;
      RECT 78.905 4.79 79.235 5.47 ;
      RECT 77.995 4.79 78.395 5.47 ;
      RECT 77.995 4.79 79.235 4.96 ;
      RECT 77.495 4.37 77.815 5.47 ;
      RECT 77.495 4.37 77.945 4.62 ;
      RECT 77.495 4.37 78.125 4.54 ;
      RECT 77.955 3.32 78.125 4.54 ;
      RECT 77.955 3.32 78.91 3.49 ;
      RECT 77.495 7.56 78.19 8.19 ;
      RECT 78.02 5.98 78.19 8.19 ;
      RECT 77.925 5.98 78.255 6.96 ;
      RECT 77.515 7.12 77.85 7.37 ;
      RECT 76.97 7.12 77.305 7.37 ;
      RECT 76.97 7.17 77.85 7.34 ;
      RECT 76.63 7.56 77.325 8.19 ;
      RECT 76.63 5.98 76.8 8.19 ;
      RECT 76.565 5.98 76.895 6.96 ;
      RECT 76.125 4.5 76.455 5.455 ;
      RECT 76.125 4.5 76.805 4.67 ;
      RECT 76.635 3.26 76.805 4.67 ;
      RECT 76.545 3.26 76.875 3.9 ;
      RECT 75.605 4.5 75.935 5.455 ;
      RECT 75.255 4.5 75.935 4.67 ;
      RECT 75.255 3.26 75.425 4.67 ;
      RECT 75.185 3.26 75.515 3.9 ;
      RECT 75.395 7.17 75.565 8.02 ;
      RECT 74.67 7.12 75.005 7.37 ;
      RECT 74.67 7.17 75.565 7.34 ;
      RECT 74.735 4.08 75.085 4.33 ;
      RECT 74.215 4.08 74.545 4.33 ;
      RECT 74.215 4.11 75.085 4.28 ;
      RECT 74.33 7.56 75.025 8.19 ;
      RECT 74.33 5.98 74.5 8.19 ;
      RECT 74.265 5.98 74.595 6.96 ;
      RECT 73.795 4.49 74.125 5.47 ;
      RECT 73.795 3.26 74.045 5.47 ;
      RECT 73.795 3.26 74.125 3.89 ;
      RECT 72.125 10.045 72.3 10.595 ;
      RECT 72.125 7.305 72.295 10.595 ;
      RECT 72.125 7.305 72.3 8.445 ;
      RECT 71.695 7.305 71.865 9.515 ;
      RECT 71.695 7.305 71.87 8.565 ;
      RECT 70.74 10.105 70.915 10.595 ;
      RECT 70.74 7.305 70.91 10.595 ;
      RECT 70.74 9.605 71.15 9.935 ;
      RECT 70.74 8.765 71.15 9.095 ;
      RECT 70.74 7.305 70.915 8.565 ;
      RECT 68.94 7.305 69.11 8.775 ;
      RECT 68.94 7.305 69.115 8.565 ;
      RECT 68.57 9.255 69.04 9.425 ;
      RECT 68.57 8.235 68.74 9.425 ;
      RECT 68.565 3.035 68.735 4.225 ;
      RECT 68.565 3.035 69.035 3.205 ;
      RECT 67.95 3.895 68.125 5.155 ;
      RECT 67.95 3.685 68.12 5.155 ;
      RECT 67.95 7.305 68.12 8.775 ;
      RECT 67.95 7.305 68.125 8.565 ;
      RECT 67.58 3.035 67.75 4.225 ;
      RECT 67.58 3.035 68.05 3.205 ;
      RECT 67.58 9.255 68.05 9.425 ;
      RECT 67.58 8.235 67.75 9.425 ;
      RECT 66.59 4.015 66.765 5.155 ;
      RECT 66.59 1.865 66.76 5.155 ;
      RECT 66.59 1.865 66.765 2.415 ;
      RECT 66.59 10.045 66.765 10.595 ;
      RECT 66.59 7.305 66.76 10.595 ;
      RECT 66.59 7.305 66.765 8.445 ;
      RECT 66.16 3.895 66.335 5.155 ;
      RECT 66.16 2.945 66.33 5.155 ;
      RECT 66.16 7.305 66.33 9.515 ;
      RECT 66.16 7.305 66.335 8.565 ;
      RECT 65.73 3.925 65.9 5.155 ;
      RECT 65.79 2.145 65.96 4.095 ;
      RECT 65.73 1.865 65.9 2.315 ;
      RECT 65.73 10.145 65.9 10.595 ;
      RECT 65.79 8.365 65.96 10.315 ;
      RECT 65.73 7.305 65.9 8.535 ;
      RECT 65.205 3.895 65.38 5.155 ;
      RECT 65.205 1.865 65.375 5.155 ;
      RECT 65.205 3.365 65.615 3.695 ;
      RECT 65.205 2.525 65.615 2.855 ;
      RECT 65.205 1.865 65.38 2.355 ;
      RECT 65.205 10.105 65.38 10.595 ;
      RECT 65.205 7.305 65.375 10.595 ;
      RECT 65.205 9.605 65.615 9.935 ;
      RECT 65.205 8.765 65.615 9.095 ;
      RECT 65.205 7.305 65.38 8.565 ;
      RECT 62.945 4.79 63.325 5.47 ;
      RECT 63.155 3.66 63.325 5.47 ;
      RECT 61.075 3.66 61.305 4.33 ;
      RECT 61.075 3.66 63.325 3.83 ;
      RECT 62.605 3.34 62.775 3.83 ;
      RECT 62.595 4.45 62.765 5.3 ;
      RECT 61.68 4.45 62.985 4.62 ;
      RECT 62.74 4 62.985 4.62 ;
      RECT 61.68 4.08 61.85 4.62 ;
      RECT 61.475 4.08 61.85 4.25 ;
      RECT 61.655 7.56 62.35 8.19 ;
      RECT 62.18 5.98 62.35 8.19 ;
      RECT 62.085 5.98 62.415 6.96 ;
      RECT 61.685 4.79 62.015 5.47 ;
      RECT 60.775 4.79 61.175 5.47 ;
      RECT 60.775 4.79 62.015 4.96 ;
      RECT 60.275 4.37 60.595 5.47 ;
      RECT 60.275 4.37 60.725 4.62 ;
      RECT 60.275 4.37 60.905 4.54 ;
      RECT 60.735 3.32 60.905 4.54 ;
      RECT 60.735 3.32 61.69 3.49 ;
      RECT 60.275 7.56 60.97 8.19 ;
      RECT 60.8 5.98 60.97 8.19 ;
      RECT 60.705 5.98 61.035 6.96 ;
      RECT 60.295 7.12 60.63 7.37 ;
      RECT 59.75 7.12 60.085 7.37 ;
      RECT 59.75 7.17 60.63 7.34 ;
      RECT 59.41 7.56 60.105 8.19 ;
      RECT 59.41 5.98 59.58 8.19 ;
      RECT 59.345 5.98 59.675 6.96 ;
      RECT 58.905 4.5 59.235 5.455 ;
      RECT 58.905 4.5 59.585 4.67 ;
      RECT 59.415 3.26 59.585 4.67 ;
      RECT 59.325 3.26 59.655 3.9 ;
      RECT 58.385 4.5 58.715 5.455 ;
      RECT 58.035 4.5 58.715 4.67 ;
      RECT 58.035 3.26 58.205 4.67 ;
      RECT 57.965 3.26 58.295 3.9 ;
      RECT 58.175 7.17 58.345 8.02 ;
      RECT 57.45 7.12 57.785 7.37 ;
      RECT 57.45 7.17 58.345 7.34 ;
      RECT 57.515 4.08 57.865 4.33 ;
      RECT 56.995 4.08 57.325 4.33 ;
      RECT 56.995 4.11 57.865 4.28 ;
      RECT 57.11 7.56 57.805 8.19 ;
      RECT 57.11 5.98 57.28 8.19 ;
      RECT 57.045 5.98 57.375 6.96 ;
      RECT 56.575 4.49 56.905 5.47 ;
      RECT 56.575 3.26 56.825 5.47 ;
      RECT 56.575 3.26 56.905 3.89 ;
      RECT 54.905 10.045 55.08 10.595 ;
      RECT 54.905 7.305 55.075 10.595 ;
      RECT 54.905 7.305 55.08 8.445 ;
      RECT 54.475 7.305 54.645 9.515 ;
      RECT 54.475 7.305 54.65 8.565 ;
      RECT 53.52 10.105 53.695 10.595 ;
      RECT 53.52 7.305 53.69 10.595 ;
      RECT 53.52 9.605 53.93 9.935 ;
      RECT 53.52 8.765 53.93 9.095 ;
      RECT 53.52 7.305 53.695 8.565 ;
      RECT 51.72 7.305 51.89 8.775 ;
      RECT 51.72 7.305 51.895 8.565 ;
      RECT 51.35 9.255 51.82 9.425 ;
      RECT 51.35 8.235 51.52 9.425 ;
      RECT 51.345 3.035 51.515 4.225 ;
      RECT 51.345 3.035 51.815 3.205 ;
      RECT 50.73 3.895 50.905 5.155 ;
      RECT 50.73 3.685 50.9 5.155 ;
      RECT 50.73 7.305 50.9 8.775 ;
      RECT 50.73 7.305 50.905 8.565 ;
      RECT 50.36 3.035 50.53 4.225 ;
      RECT 50.36 3.035 50.83 3.205 ;
      RECT 50.36 9.255 50.83 9.425 ;
      RECT 50.36 8.235 50.53 9.425 ;
      RECT 49.37 4.015 49.545 5.155 ;
      RECT 49.37 1.865 49.54 5.155 ;
      RECT 49.37 1.865 49.545 2.415 ;
      RECT 49.37 10.045 49.545 10.595 ;
      RECT 49.37 7.305 49.54 10.595 ;
      RECT 49.37 7.305 49.545 8.445 ;
      RECT 48.94 3.895 49.115 5.155 ;
      RECT 48.94 2.945 49.11 5.155 ;
      RECT 48.94 7.305 49.11 9.515 ;
      RECT 48.94 7.305 49.115 8.565 ;
      RECT 48.51 3.925 48.68 5.155 ;
      RECT 48.57 2.145 48.74 4.095 ;
      RECT 48.51 1.865 48.68 2.315 ;
      RECT 48.51 10.145 48.68 10.595 ;
      RECT 48.57 8.365 48.74 10.315 ;
      RECT 48.51 7.305 48.68 8.535 ;
      RECT 47.985 3.895 48.16 5.155 ;
      RECT 47.985 1.865 48.155 5.155 ;
      RECT 47.985 3.365 48.395 3.695 ;
      RECT 47.985 2.525 48.395 2.855 ;
      RECT 47.985 1.865 48.16 2.355 ;
      RECT 47.985 10.105 48.16 10.595 ;
      RECT 47.985 7.305 48.155 10.595 ;
      RECT 47.985 9.605 48.395 9.935 ;
      RECT 47.985 8.765 48.395 9.095 ;
      RECT 47.985 7.305 48.16 8.565 ;
      RECT 45.725 4.79 46.105 5.47 ;
      RECT 45.935 3.66 46.105 5.47 ;
      RECT 43.855 3.66 44.085 4.33 ;
      RECT 43.855 3.66 46.105 3.83 ;
      RECT 45.385 3.34 45.555 3.83 ;
      RECT 45.375 4.45 45.545 5.3 ;
      RECT 44.46 4.45 45.765 4.62 ;
      RECT 45.52 4 45.765 4.62 ;
      RECT 44.46 4.08 44.63 4.62 ;
      RECT 44.255 4.08 44.63 4.25 ;
      RECT 44.435 7.56 45.13 8.19 ;
      RECT 44.96 5.98 45.13 8.19 ;
      RECT 44.865 5.98 45.195 6.96 ;
      RECT 44.465 4.79 44.795 5.47 ;
      RECT 43.555 4.79 43.955 5.47 ;
      RECT 43.555 4.79 44.795 4.96 ;
      RECT 43.055 4.37 43.375 5.47 ;
      RECT 43.055 4.37 43.505 4.62 ;
      RECT 43.055 4.37 43.685 4.54 ;
      RECT 43.515 3.32 43.685 4.54 ;
      RECT 43.515 3.32 44.47 3.49 ;
      RECT 43.055 7.56 43.75 8.19 ;
      RECT 43.58 5.98 43.75 8.19 ;
      RECT 43.485 5.98 43.815 6.96 ;
      RECT 43.075 7.12 43.41 7.37 ;
      RECT 42.53 7.12 42.865 7.37 ;
      RECT 42.53 7.17 43.41 7.34 ;
      RECT 42.19 7.56 42.885 8.19 ;
      RECT 42.19 5.98 42.36 8.19 ;
      RECT 42.125 5.98 42.455 6.96 ;
      RECT 41.685 4.5 42.015 5.455 ;
      RECT 41.685 4.5 42.365 4.67 ;
      RECT 42.195 3.26 42.365 4.67 ;
      RECT 42.105 3.26 42.435 3.9 ;
      RECT 41.165 4.5 41.495 5.455 ;
      RECT 40.815 4.5 41.495 4.67 ;
      RECT 40.815 3.26 40.985 4.67 ;
      RECT 40.745 3.26 41.075 3.9 ;
      RECT 40.955 7.17 41.125 8.02 ;
      RECT 40.23 7.12 40.565 7.37 ;
      RECT 40.23 7.17 41.125 7.34 ;
      RECT 40.295 4.08 40.645 4.33 ;
      RECT 39.775 4.08 40.105 4.33 ;
      RECT 39.775 4.11 40.645 4.28 ;
      RECT 39.89 7.56 40.585 8.19 ;
      RECT 39.89 5.98 40.06 8.19 ;
      RECT 39.825 5.98 40.155 6.96 ;
      RECT 39.355 4.49 39.685 5.47 ;
      RECT 39.355 3.26 39.605 5.47 ;
      RECT 39.355 3.26 39.685 3.89 ;
      RECT 37.685 10.045 37.86 10.595 ;
      RECT 37.685 7.305 37.855 10.595 ;
      RECT 37.685 7.305 37.86 8.445 ;
      RECT 37.255 7.305 37.425 9.515 ;
      RECT 37.255 7.305 37.43 8.565 ;
      RECT 36.3 10.105 36.475 10.595 ;
      RECT 36.3 7.305 36.47 10.595 ;
      RECT 36.3 9.605 36.71 9.935 ;
      RECT 36.3 8.765 36.71 9.095 ;
      RECT 36.3 7.305 36.475 8.565 ;
      RECT 34.5 7.305 34.67 8.775 ;
      RECT 34.5 7.305 34.675 8.565 ;
      RECT 34.13 9.255 34.6 9.425 ;
      RECT 34.13 8.235 34.3 9.425 ;
      RECT 34.125 3.035 34.295 4.225 ;
      RECT 34.125 3.035 34.595 3.205 ;
      RECT 33.51 3.895 33.685 5.155 ;
      RECT 33.51 3.685 33.68 5.155 ;
      RECT 33.51 7.305 33.68 8.775 ;
      RECT 33.51 7.305 33.685 8.565 ;
      RECT 33.14 3.035 33.31 4.225 ;
      RECT 33.14 3.035 33.61 3.205 ;
      RECT 33.14 9.255 33.61 9.425 ;
      RECT 33.14 8.235 33.31 9.425 ;
      RECT 32.15 4.015 32.325 5.155 ;
      RECT 32.15 1.865 32.32 5.155 ;
      RECT 32.15 1.865 32.325 2.415 ;
      RECT 32.15 10.045 32.325 10.595 ;
      RECT 32.15 7.305 32.32 10.595 ;
      RECT 32.15 7.305 32.325 8.445 ;
      RECT 31.72 3.895 31.895 5.155 ;
      RECT 31.72 2.945 31.89 5.155 ;
      RECT 31.72 7.305 31.89 9.515 ;
      RECT 31.72 7.305 31.895 8.565 ;
      RECT 31.29 3.925 31.46 5.155 ;
      RECT 31.35 2.145 31.52 4.095 ;
      RECT 31.29 1.865 31.46 2.315 ;
      RECT 31.29 10.145 31.46 10.595 ;
      RECT 31.35 8.365 31.52 10.315 ;
      RECT 31.29 7.305 31.46 8.535 ;
      RECT 30.765 3.895 30.94 5.155 ;
      RECT 30.765 1.865 30.935 5.155 ;
      RECT 30.765 3.365 31.175 3.695 ;
      RECT 30.765 2.525 31.175 2.855 ;
      RECT 30.765 1.865 30.94 2.355 ;
      RECT 30.765 10.105 30.94 10.595 ;
      RECT 30.765 7.305 30.935 10.595 ;
      RECT 30.765 9.605 31.175 9.935 ;
      RECT 30.765 8.765 31.175 9.095 ;
      RECT 30.765 7.305 30.94 8.565 ;
      RECT 28.505 4.79 28.885 5.47 ;
      RECT 28.715 3.66 28.885 5.47 ;
      RECT 26.635 3.66 26.865 4.33 ;
      RECT 26.635 3.66 28.885 3.83 ;
      RECT 28.165 3.34 28.335 3.83 ;
      RECT 28.155 4.45 28.325 5.3 ;
      RECT 27.24 4.45 28.545 4.62 ;
      RECT 28.3 4 28.545 4.62 ;
      RECT 27.24 4.08 27.41 4.62 ;
      RECT 27.035 4.08 27.41 4.25 ;
      RECT 27.215 7.56 27.91 8.19 ;
      RECT 27.74 5.98 27.91 8.19 ;
      RECT 27.645 5.98 27.975 6.96 ;
      RECT 27.245 4.79 27.575 5.47 ;
      RECT 26.335 4.79 26.735 5.47 ;
      RECT 26.335 4.79 27.575 4.96 ;
      RECT 25.835 4.37 26.155 5.47 ;
      RECT 25.835 4.37 26.285 4.62 ;
      RECT 25.835 4.37 26.465 4.54 ;
      RECT 26.295 3.32 26.465 4.54 ;
      RECT 26.295 3.32 27.25 3.49 ;
      RECT 25.835 7.56 26.53 8.19 ;
      RECT 26.36 5.98 26.53 8.19 ;
      RECT 26.265 5.98 26.595 6.96 ;
      RECT 25.855 7.12 26.19 7.37 ;
      RECT 25.31 7.12 25.645 7.37 ;
      RECT 25.31 7.17 26.19 7.34 ;
      RECT 24.97 7.56 25.665 8.19 ;
      RECT 24.97 5.98 25.14 8.19 ;
      RECT 24.905 5.98 25.235 6.96 ;
      RECT 24.465 4.5 24.795 5.455 ;
      RECT 24.465 4.5 25.145 4.67 ;
      RECT 24.975 3.26 25.145 4.67 ;
      RECT 24.885 3.26 25.215 3.9 ;
      RECT 23.945 4.5 24.275 5.455 ;
      RECT 23.595 4.5 24.275 4.67 ;
      RECT 23.595 3.26 23.765 4.67 ;
      RECT 23.525 3.26 23.855 3.9 ;
      RECT 23.735 7.17 23.905 8.02 ;
      RECT 23.01 7.12 23.345 7.37 ;
      RECT 23.01 7.17 23.905 7.34 ;
      RECT 23.075 4.08 23.425 4.33 ;
      RECT 22.555 4.08 22.885 4.33 ;
      RECT 22.555 4.11 23.425 4.28 ;
      RECT 22.67 7.56 23.365 8.19 ;
      RECT 22.67 5.98 22.84 8.19 ;
      RECT 22.605 5.98 22.935 6.96 ;
      RECT 22.135 4.49 22.465 5.47 ;
      RECT 22.135 3.26 22.385 5.47 ;
      RECT 22.135 3.26 22.465 3.89 ;
      RECT 20.465 10.045 20.64 10.595 ;
      RECT 20.465 7.305 20.635 10.595 ;
      RECT 20.465 7.305 20.64 8.445 ;
      RECT 20.035 7.305 20.205 9.515 ;
      RECT 20.035 7.305 20.21 8.565 ;
      RECT 19.08 10.105 19.255 10.595 ;
      RECT 19.08 7.305 19.25 10.595 ;
      RECT 19.08 9.605 19.49 9.935 ;
      RECT 19.08 8.765 19.49 9.095 ;
      RECT 19.08 7.305 19.255 8.565 ;
      RECT 16.625 7.305 16.795 9.515 ;
      RECT 16.625 7.305 16.8 8.565 ;
      RECT 16.195 10.145 16.365 10.595 ;
      RECT 16.255 8.365 16.425 10.315 ;
      RECT 16.195 7.305 16.365 8.535 ;
      RECT 15.67 10.105 15.845 10.595 ;
      RECT 15.67 7.305 15.84 10.595 ;
      RECT 15.67 9.605 16.08 9.935 ;
      RECT 15.67 8.765 16.08 9.095 ;
      RECT 15.67 7.305 15.845 8.565 ;
      RECT 103.38 10.085 103.555 10.595 ;
      RECT 102.39 1.865 102.565 2.375 ;
      RECT 102.39 10.085 102.565 10.595 ;
      RECT 100.6 1.865 100.775 2.375 ;
      RECT 100.6 10.085 100.775 10.595 ;
      RECT 96.96 7.12 97.295 7.39 ;
      RECT 96.46 4.08 97.01 4.28 ;
      RECT 96.115 7.12 96.45 7.37 ;
      RECT 95.58 7.12 95.915 7.39 ;
      RECT 94.195 4.08 94.545 4.33 ;
      RECT 93.335 4.08 93.685 4.33 ;
      RECT 92.815 4.08 93.165 4.33 ;
      RECT 88.915 10.085 89.09 10.595 ;
      RECT 86.16 10.085 86.335 10.595 ;
      RECT 85.17 1.865 85.345 2.375 ;
      RECT 85.17 10.085 85.345 10.595 ;
      RECT 83.38 1.865 83.555 2.375 ;
      RECT 83.38 10.085 83.555 10.595 ;
      RECT 79.74 7.12 80.075 7.39 ;
      RECT 79.24 4.08 79.79 4.28 ;
      RECT 78.895 7.12 79.23 7.37 ;
      RECT 78.36 7.12 78.695 7.39 ;
      RECT 76.975 4.08 77.325 4.33 ;
      RECT 76.115 4.08 76.465 4.33 ;
      RECT 75.595 4.08 75.945 4.33 ;
      RECT 71.695 10.085 71.87 10.595 ;
      RECT 68.94 10.085 69.115 10.595 ;
      RECT 67.95 1.865 68.125 2.375 ;
      RECT 67.95 10.085 68.125 10.595 ;
      RECT 66.16 1.865 66.335 2.375 ;
      RECT 66.16 10.085 66.335 10.595 ;
      RECT 62.52 7.12 62.855 7.39 ;
      RECT 62.02 4.08 62.57 4.28 ;
      RECT 61.675 7.12 62.01 7.37 ;
      RECT 61.14 7.12 61.475 7.39 ;
      RECT 59.755 4.08 60.105 4.33 ;
      RECT 58.895 4.08 59.245 4.33 ;
      RECT 58.375 4.08 58.725 4.33 ;
      RECT 54.475 10.085 54.65 10.595 ;
      RECT 51.72 10.085 51.895 10.595 ;
      RECT 50.73 1.865 50.905 2.375 ;
      RECT 50.73 10.085 50.905 10.595 ;
      RECT 48.94 1.865 49.115 2.375 ;
      RECT 48.94 10.085 49.115 10.595 ;
      RECT 45.3 7.12 45.635 7.39 ;
      RECT 44.8 4.08 45.35 4.28 ;
      RECT 44.455 7.12 44.79 7.37 ;
      RECT 43.92 7.12 44.255 7.39 ;
      RECT 42.535 4.08 42.885 4.33 ;
      RECT 41.675 4.08 42.025 4.33 ;
      RECT 41.155 4.08 41.505 4.33 ;
      RECT 37.255 10.085 37.43 10.595 ;
      RECT 34.5 10.085 34.675 10.595 ;
      RECT 33.51 1.865 33.685 2.375 ;
      RECT 33.51 10.085 33.685 10.595 ;
      RECT 31.72 1.865 31.895 2.375 ;
      RECT 31.72 10.085 31.895 10.595 ;
      RECT 28.08 7.12 28.415 7.39 ;
      RECT 27.58 4.08 28.13 4.28 ;
      RECT 27.235 7.12 27.57 7.37 ;
      RECT 26.7 7.12 27.035 7.39 ;
      RECT 25.315 4.08 25.665 4.33 ;
      RECT 24.455 4.08 24.805 4.33 ;
      RECT 23.935 4.08 24.285 4.33 ;
      RECT 20.035 10.085 20.21 10.595 ;
      RECT 16.625 10.085 16.8 10.595 ;
  END
END sky130_osu_ring_oscillator_mpr2ct_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2ct_8_b0r2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ct_8_b0r2 ;
  SIZE 103.915 BY 12.465 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 34.37 0 34.75 5.265 ;
      LAYER met2 ;
        RECT 34.37 4.885 34.75 5.265 ;
      LAYER li1 ;
        RECT 34.47 1.865 34.645 2.375 ;
        RECT 34.47 3.895 34.645 5.155 ;
        RECT 34.47 3.685 34.64 5.155 ;
      LAYER met1 ;
        RECT 34.385 4.93 34.735 5.22 ;
        RECT 34.41 2.175 34.705 2.405 ;
        RECT 34.41 3.655 34.7 3.885 ;
        RECT 34.47 2.175 34.64 3.885 ;
      LAYER via1 ;
        RECT 34.485 5 34.635 5.15 ;
      LAYER via2 ;
        RECT 34.46 4.975 34.66 5.175 ;
      LAYER mcon ;
        RECT 34.47 3.685 34.64 3.855 ;
        RECT 34.47 2.205 34.64 2.375 ;
        RECT 34.475 4.985 34.645 5.155 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 51.59 0 51.97 5.265 ;
      LAYER met2 ;
        RECT 51.59 4.885 51.97 5.265 ;
      LAYER li1 ;
        RECT 51.69 1.865 51.865 2.375 ;
        RECT 51.69 3.895 51.865 5.155 ;
        RECT 51.69 3.685 51.86 5.155 ;
      LAYER met1 ;
        RECT 51.605 4.93 51.955 5.22 ;
        RECT 51.63 2.175 51.925 2.405 ;
        RECT 51.63 3.655 51.92 3.885 ;
        RECT 51.69 2.175 51.86 3.885 ;
      LAYER via1 ;
        RECT 51.705 5 51.855 5.15 ;
      LAYER via2 ;
        RECT 51.68 4.975 51.88 5.175 ;
      LAYER mcon ;
        RECT 51.69 3.685 51.86 3.855 ;
        RECT 51.69 2.205 51.86 2.375 ;
        RECT 51.695 4.985 51.865 5.155 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 68.81 0.005 69.19 5.27 ;
      LAYER met2 ;
        RECT 68.81 4.89 69.19 5.27 ;
      LAYER li1 ;
        RECT 68.91 1.87 69.085 2.38 ;
        RECT 68.91 3.9 69.085 5.16 ;
        RECT 68.91 3.69 69.08 5.16 ;
      LAYER met1 ;
        RECT 68.825 4.935 69.175 5.225 ;
        RECT 68.85 2.18 69.145 2.41 ;
        RECT 68.85 3.66 69.14 3.89 ;
        RECT 68.91 2.18 69.08 3.89 ;
      LAYER via1 ;
        RECT 68.925 5.005 69.075 5.155 ;
      LAYER via2 ;
        RECT 68.9 4.98 69.1 5.18 ;
      LAYER mcon ;
        RECT 68.91 3.69 69.08 3.86 ;
        RECT 68.91 2.21 69.08 2.38 ;
        RECT 68.915 4.99 69.085 5.16 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 86.03 0 86.41 5.265 ;
      LAYER met2 ;
        RECT 86.03 4.885 86.41 5.265 ;
      LAYER li1 ;
        RECT 86.13 1.865 86.305 2.375 ;
        RECT 86.13 3.895 86.305 5.155 ;
        RECT 86.13 3.685 86.3 5.155 ;
      LAYER met1 ;
        RECT 86.045 4.93 86.395 5.22 ;
        RECT 86.07 2.175 86.365 2.405 ;
        RECT 86.07 3.655 86.36 3.885 ;
        RECT 86.13 3.2 86.31 3.37 ;
        RECT 86.13 2.175 86.3 3.885 ;
      LAYER via1 ;
        RECT 86.145 5 86.295 5.15 ;
      LAYER via2 ;
        RECT 86.12 4.975 86.32 5.175 ;
      LAYER mcon ;
        RECT 86.13 3.685 86.3 3.855 ;
        RECT 86.13 2.205 86.3 2.375 ;
        RECT 86.135 4.985 86.305 5.155 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 103.25 0 103.63 5.265 ;
      LAYER met2 ;
        RECT 103.25 4.885 103.63 5.265 ;
      LAYER li1 ;
        RECT 103.35 1.865 103.525 2.375 ;
        RECT 103.35 3.895 103.525 5.155 ;
        RECT 103.35 3.685 103.52 5.155 ;
      LAYER met1 ;
        RECT 103.265 4.93 103.615 5.22 ;
        RECT 103.29 2.175 103.585 2.405 ;
        RECT 103.29 3.655 103.58 3.885 ;
        RECT 103.35 2.175 103.52 3.885 ;
      LAYER via1 ;
        RECT 103.365 5 103.515 5.15 ;
      LAYER via2 ;
        RECT 103.34 4.975 103.54 5.175 ;
      LAYER mcon ;
        RECT 103.35 3.685 103.52 3.855 ;
        RECT 103.35 2.205 103.52 2.375 ;
        RECT 103.355 4.985 103.525 5.155 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 30.245 8.14 30.57 8.465 ;
        RECT 30.245 4.79 30.57 5.115 ;
        RECT 20.945 9.24 30.495 9.41 ;
        RECT 30.325 8.14 30.495 9.41 ;
        RECT 30.315 4.79 30.485 8.465 ;
        RECT 20.89 8.145 21.17 8.485 ;
        RECT 20.945 8.145 21.115 9.41 ;
      LAYER li1 ;
        RECT 30.315 8.225 30.495 8.465 ;
        RECT 30.32 8.225 30.49 9.505 ;
        RECT 30.32 2.955 30.49 4.225 ;
        RECT 18.635 8.235 18.805 9.505 ;
      LAYER met1 ;
        RECT 30.26 4.055 30.72 4.225 ;
        RECT 30.245 4.79 30.57 5.115 ;
        RECT 30.26 4.025 30.55 4.255 ;
        RECT 30.325 4.025 30.495 5.115 ;
        RECT 30.245 8.235 30.72 8.405 ;
        RECT 30.245 8.14 30.57 8.465 ;
        RECT 20.86 8.175 21.2 8.455 ;
        RECT 18.575 8.23 21.2 8.4 ;
        RECT 18.575 8.23 19.035 8.405 ;
        RECT 18.575 8.205 18.865 8.435 ;
      LAYER via1 ;
        RECT 20.955 8.24 21.105 8.39 ;
        RECT 30.335 8.225 30.485 8.375 ;
        RECT 30.335 4.875 30.485 5.025 ;
      LAYER mcon ;
        RECT 18.635 8.235 18.805 8.405 ;
        RECT 30.32 8.235 30.49 8.405 ;
        RECT 30.32 4.055 30.49 4.225 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 47.465 8.14 47.79 8.465 ;
        RECT 47.465 4.79 47.79 5.115 ;
        RECT 38.165 9.24 47.715 9.41 ;
        RECT 47.545 8.14 47.715 9.41 ;
        RECT 47.535 4.79 47.705 8.465 ;
        RECT 38.11 8.145 38.39 8.485 ;
        RECT 38.165 8.145 38.335 9.41 ;
      LAYER li1 ;
        RECT 47.535 8.225 47.715 8.465 ;
        RECT 47.54 8.225 47.71 9.505 ;
        RECT 47.54 2.955 47.71 4.225 ;
        RECT 35.855 8.235 36.025 9.505 ;
      LAYER met1 ;
        RECT 47.48 4.055 47.94 4.225 ;
        RECT 47.465 4.79 47.79 5.115 ;
        RECT 47.48 4.025 47.77 4.255 ;
        RECT 47.545 4.025 47.715 5.115 ;
        RECT 47.465 8.235 47.94 8.405 ;
        RECT 47.465 8.14 47.79 8.465 ;
        RECT 38.08 8.175 38.42 8.455 ;
        RECT 35.795 8.23 38.42 8.4 ;
        RECT 35.795 8.23 36.255 8.405 ;
        RECT 35.795 8.205 36.085 8.435 ;
      LAYER via1 ;
        RECT 38.175 8.24 38.325 8.39 ;
        RECT 47.555 8.225 47.705 8.375 ;
        RECT 47.555 4.875 47.705 5.025 ;
      LAYER mcon ;
        RECT 35.855 8.235 36.025 8.405 ;
        RECT 47.54 8.235 47.71 8.405 ;
        RECT 47.54 4.055 47.71 4.225 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 64.685 8.145 65.01 8.47 ;
        RECT 64.685 4.795 65.01 5.12 ;
        RECT 55.385 9.245 64.935 9.415 ;
        RECT 64.765 8.145 64.935 9.415 ;
        RECT 64.755 4.795 64.925 8.47 ;
        RECT 55.33 8.15 55.61 8.49 ;
        RECT 55.385 8.15 55.555 9.415 ;
      LAYER li1 ;
        RECT 64.755 8.23 64.935 8.47 ;
        RECT 64.76 8.23 64.93 9.51 ;
        RECT 64.76 2.96 64.93 4.23 ;
        RECT 53.075 8.24 53.245 9.51 ;
      LAYER met1 ;
        RECT 64.7 4.06 65.16 4.23 ;
        RECT 64.685 4.795 65.01 5.12 ;
        RECT 64.7 4.03 64.99 4.26 ;
        RECT 64.765 4.03 64.935 5.12 ;
        RECT 64.685 8.24 65.16 8.41 ;
        RECT 64.685 8.145 65.01 8.47 ;
        RECT 55.3 8.18 55.64 8.46 ;
        RECT 53.015 8.235 55.64 8.405 ;
        RECT 53.015 8.235 53.475 8.41 ;
        RECT 53.015 8.21 53.305 8.44 ;
      LAYER via1 ;
        RECT 55.395 8.245 55.545 8.395 ;
        RECT 64.775 8.23 64.925 8.38 ;
        RECT 64.775 4.88 64.925 5.03 ;
      LAYER mcon ;
        RECT 53.075 8.24 53.245 8.41 ;
        RECT 64.76 8.24 64.93 8.41 ;
        RECT 64.76 4.06 64.93 4.23 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 81.905 8.14 82.23 8.465 ;
        RECT 81.905 4.79 82.23 5.115 ;
        RECT 72.605 9.24 82.155 9.41 ;
        RECT 81.985 8.14 82.155 9.41 ;
        RECT 81.975 4.79 82.145 8.465 ;
        RECT 72.55 8.145 72.83 8.485 ;
        RECT 72.605 8.145 72.775 9.41 ;
      LAYER li1 ;
        RECT 81.975 8.225 82.155 8.465 ;
        RECT 81.98 8.225 82.15 9.505 ;
        RECT 81.98 2.955 82.15 4.225 ;
        RECT 70.295 8.235 70.465 9.505 ;
      LAYER met1 ;
        RECT 81.92 4.055 82.38 4.225 ;
        RECT 81.905 4.79 82.23 5.115 ;
        RECT 81.92 4.025 82.21 4.255 ;
        RECT 81.985 4.025 82.155 5.115 ;
        RECT 81.905 8.235 82.38 8.405 ;
        RECT 81.905 8.14 82.23 8.465 ;
        RECT 72.52 8.175 72.86 8.455 ;
        RECT 70.235 8.23 72.86 8.4 ;
        RECT 70.235 8.23 70.695 8.405 ;
        RECT 70.235 8.205 70.525 8.435 ;
      LAYER via1 ;
        RECT 72.615 8.24 72.765 8.39 ;
        RECT 81.995 8.225 82.145 8.375 ;
        RECT 81.995 4.875 82.145 5.025 ;
      LAYER mcon ;
        RECT 70.295 8.235 70.465 8.405 ;
        RECT 81.98 8.235 82.15 8.405 ;
        RECT 81.98 4.055 82.15 4.225 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 99.125 8.14 99.45 8.465 ;
        RECT 99.125 4.79 99.45 5.115 ;
        RECT 89.825 9.24 99.375 9.41 ;
        RECT 99.205 8.14 99.375 9.41 ;
        RECT 99.195 4.79 99.365 8.465 ;
        RECT 89.77 8.145 90.05 8.485 ;
        RECT 89.825 8.145 89.995 9.41 ;
      LAYER li1 ;
        RECT 99.195 8.225 99.375 8.465 ;
        RECT 99.2 8.225 99.37 9.505 ;
        RECT 99.2 2.955 99.37 4.225 ;
        RECT 87.515 8.235 87.685 9.505 ;
      LAYER met1 ;
        RECT 99.14 4.055 99.6 4.225 ;
        RECT 99.125 4.79 99.45 5.115 ;
        RECT 99.14 4.025 99.43 4.255 ;
        RECT 99.205 4.025 99.375 5.115 ;
        RECT 99.125 8.235 99.6 8.405 ;
        RECT 99.125 8.14 99.45 8.465 ;
        RECT 89.74 8.175 90.08 8.455 ;
        RECT 87.455 8.23 90.08 8.4 ;
        RECT 87.455 8.23 87.915 8.405 ;
        RECT 87.455 8.205 87.745 8.435 ;
      LAYER via1 ;
        RECT 89.835 8.24 89.985 8.39 ;
        RECT 99.215 8.225 99.365 8.375 ;
        RECT 99.215 4.875 99.365 5.025 ;
      LAYER mcon ;
        RECT 87.515 8.235 87.685 8.405 ;
        RECT 99.2 8.235 99.37 8.405 ;
        RECT 99.2 4.055 99.37 4.225 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 15.225 8.235 15.395 9.505 ;
      LAYER met1 ;
        RECT 15.165 8.235 15.625 8.405 ;
        RECT 15.17 8.2 15.46 8.43 ;
        RECT 15.165 8.205 15.455 8.435 ;
      LAYER mcon ;
        RECT 15.225 8.235 15.395 8.405 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 97.915 5.43 103.9 7.03 ;
        RECT 99.02 5.43 103.745 7.035 ;
        RECT 99.02 5.425 103.74 7.035 ;
        RECT 102.925 5.425 103.095 7.765 ;
        RECT 102.92 4.695 103.09 7.035 ;
        RECT 101.935 4.695 102.105 7.765 ;
        RECT 99.19 4.695 99.36 7.765 ;
        RECT 97.815 5.64 103.9 6.8 ;
        RECT 97.91 5.43 103.9 6.8 ;
        RECT 63.47 5.64 103.9 5.81 ;
        RECT 97 5.64 97.28 6.95 ;
        RECT 96.6 4.79 96.77 5.81 ;
        RECT 96.07 5.64 96.33 6.95 ;
        RECT 95.76 5.13 95.93 5.81 ;
        RECT 95.62 5.64 95.9 6.95 ;
        RECT 94.69 5.64 94.95 6.95 ;
        RECT 94.26 5.64 94.52 6.95 ;
        RECT 94.18 4.5 94.51 5.81 ;
        RECT 93.31 5.64 93.59 6.95 ;
        RECT 91.94 4.5 92.27 5.81 ;
        RECT 91.96 4.5 92.22 6.95 ;
        RECT 91.49 4.5 91.72 5.81 ;
        RECT 91.01 5.64 91.29 6.95 ;
        RECT 80.595 5.64 90.825 6.8 ;
        RECT 80.69 5.43 90.82 6.8 ;
        RECT 90.61 4.5 90.82 6.8 ;
        RECT 81.8 5.425 90.82 6.8 ;
        RECT 80.695 5.43 90.245 7.03 ;
        RECT 87.335 5.425 90.085 7.035 ;
        RECT 87.505 5.425 87.675 7.765 ;
        RECT 81.8 5.425 86.525 7.035 ;
        RECT 85.705 5.425 85.875 7.765 ;
        RECT 85.7 4.695 85.87 7.035 ;
        RECT 84.715 4.695 84.885 7.765 ;
        RECT 81.97 4.695 82.14 7.765 ;
        RECT 79.78 5.64 80.06 6.95 ;
        RECT 79.38 4.79 79.55 5.81 ;
        RECT 78.85 5.64 79.11 6.95 ;
        RECT 78.54 5.13 78.71 5.81 ;
        RECT 78.4 5.64 78.68 6.95 ;
        RECT 77.47 5.64 77.73 6.95 ;
        RECT 77.04 5.64 77.3 6.95 ;
        RECT 76.96 4.5 77.29 5.81 ;
        RECT 76.09 5.64 76.37 6.95 ;
        RECT 74.72 4.5 75.05 5.81 ;
        RECT 74.74 4.5 75 6.95 ;
        RECT 74.27 4.5 74.5 5.81 ;
        RECT 73.79 5.64 74.07 6.95 ;
        RECT 63.375 5.645 73.605 6.8 ;
        RECT 63.47 5.435 73.6 6.8 ;
        RECT 73.39 4.5 73.6 6.8 ;
        RECT 69.455 5.425 73.6 6.8 ;
        RECT 63.475 5.43 73.025 7.03 ;
        RECT 70.115 5.425 72.865 7.035 ;
        RECT 70.285 5.425 70.455 7.765 ;
        RECT 63.475 5.43 69.46 7.035 ;
        RECT 64.58 5.43 69.305 7.04 ;
        RECT 68.485 5.43 68.655 7.77 ;
        RECT 68.48 4.7 68.65 7.04 ;
        RECT 67.495 4.7 67.665 7.77 ;
        RECT 64.75 4.7 64.92 7.77 ;
        RECT 63.375 5.645 73.025 6.805 ;
        RECT 46.155 5.645 73.605 5.815 ;
        RECT 62.56 5.645 62.84 6.955 ;
        RECT 62.16 4.795 62.33 5.815 ;
        RECT 61.63 5.645 61.89 6.955 ;
        RECT 61.32 5.135 61.49 5.815 ;
        RECT 61.18 5.645 61.46 6.955 ;
        RECT 60.25 5.645 60.51 6.955 ;
        RECT 59.82 5.645 60.08 6.955 ;
        RECT 59.74 4.505 60.07 5.815 ;
        RECT 58.87 5.645 59.15 6.955 ;
        RECT 57.5 4.505 57.83 5.815 ;
        RECT 57.52 4.505 57.78 6.955 ;
        RECT 57.05 4.505 57.28 5.815 ;
        RECT 56.57 5.645 56.85 6.955 ;
        RECT 46.255 5.645 56.385 6.805 ;
        RECT 0 5.64 56.38 5.81 ;
        RECT 56.17 4.505 56.38 6.805 ;
        RECT 46.25 5.43 56.38 6.8 ;
        RECT 46.255 5.43 55.805 7.03 ;
        RECT 52.895 5.43 55.645 7.04 ;
        RECT 53.065 5.43 53.235 7.77 ;
        RECT 47.36 5.43 52.085 7.035 ;
        RECT 47.36 5.425 52.08 7.035 ;
        RECT 51.265 5.425 51.435 7.765 ;
        RECT 51.26 4.695 51.43 7.035 ;
        RECT 50.275 4.695 50.445 7.765 ;
        RECT 47.53 4.695 47.7 7.765 ;
        RECT 46.155 5.645 56.385 6.8 ;
        RECT 45.34 5.64 45.62 6.95 ;
        RECT 44.94 4.79 45.11 5.81 ;
        RECT 44.41 5.64 44.67 6.95 ;
        RECT 44.1 5.13 44.27 5.81 ;
        RECT 43.96 5.64 44.24 6.95 ;
        RECT 43.03 5.64 43.29 6.95 ;
        RECT 42.6 5.64 42.86 6.95 ;
        RECT 42.52 4.5 42.85 5.81 ;
        RECT 41.65 5.64 41.93 6.95 ;
        RECT 40.28 4.5 40.61 5.81 ;
        RECT 40.3 4.5 40.56 6.95 ;
        RECT 39.83 4.5 40.06 5.81 ;
        RECT 39.35 5.64 39.63 6.95 ;
        RECT 28.935 5.64 39.165 6.8 ;
        RECT 29.03 5.43 39.16 6.8 ;
        RECT 38.95 4.5 39.16 6.8 ;
        RECT 30.14 5.425 39.16 6.8 ;
        RECT 29.035 5.43 38.585 7.005 ;
        RECT 29.035 5.43 38.58 7.03 ;
        RECT 35.675 5.425 38.425 7.035 ;
        RECT 35.845 5.425 36.015 7.765 ;
        RECT 30.14 5.425 34.865 7.035 ;
        RECT 34.045 5.425 34.215 7.765 ;
        RECT 34.04 4.695 34.21 7.035 ;
        RECT 33.055 4.695 33.225 7.765 ;
        RECT 30.31 4.695 30.48 7.765 ;
        RECT 28.12 5.64 28.4 6.95 ;
        RECT 27.72 4.79 27.89 5.81 ;
        RECT 27.19 5.64 27.45 6.95 ;
        RECT 26.88 5.13 27.05 5.81 ;
        RECT 26.74 5.64 27.02 6.95 ;
        RECT 25.81 5.64 26.07 6.95 ;
        RECT 25.38 5.64 25.64 6.95 ;
        RECT 25.3 4.5 25.63 5.81 ;
        RECT 24.43 5.64 24.71 6.95 ;
        RECT 23.06 4.5 23.39 5.81 ;
        RECT 23.08 4.5 23.34 6.95 ;
        RECT 22.61 4.5 22.84 5.81 ;
        RECT 22.13 5.64 22.41 6.95 ;
        RECT 0 5.64 21.945 6.8 ;
        RECT 0 5.425 21.94 7 ;
        RECT 21.73 4.5 21.94 7 ;
        RECT 0 5.425 21.47 7.025 ;
        RECT 18.455 5.425 21.205 7.035 ;
        RECT 18.625 5.425 18.795 7.765 ;
        RECT 15.045 5.425 17.795 7.035 ;
        RECT 17.03 10.045 17.205 10.595 ;
        RECT 17.03 7.305 17.205 8.445 ;
        RECT 17.03 5.425 17.2 10.595 ;
        RECT 15.215 5.425 15.385 7.765 ;
      LAYER met1 ;
        RECT 97.915 5.43 103.9 7.03 ;
        RECT 99.02 5.43 103.745 7.035 ;
        RECT 99.02 5.425 103.74 7.035 ;
        RECT 97.825 5.485 103.9 6.955 ;
        RECT 97.91 5.43 103.9 6.955 ;
        RECT 97.815 5.485 103.9 6.8 ;
        RECT 63.47 5.485 103.9 5.965 ;
        RECT 80.595 5.485 90.825 6.8 ;
        RECT 80.69 5.43 90.82 6.8 ;
        RECT 81.8 5.425 90.82 6.8 ;
        RECT 80.695 5.43 90.245 7.03 ;
        RECT 87.335 5.425 90.085 7.035 ;
        RECT 81.8 5.425 86.525 7.035 ;
        RECT 80.605 5.485 90.245 6.955 ;
        RECT 63.375 5.49 73.605 6.8 ;
        RECT 63.47 5.435 73.6 6.8 ;
        RECT 69.455 5.425 73.6 6.8 ;
        RECT 63.475 5.43 73.025 7.03 ;
        RECT 70.115 5.425 72.865 7.035 ;
        RECT 63.475 5.43 69.46 7.035 ;
        RECT 64.58 5.43 69.305 7.04 ;
        RECT 63.385 5.49 73.025 6.96 ;
        RECT 63.375 5.49 73.025 6.805 ;
        RECT 46.155 5.49 73.605 5.97 ;
        RECT 46.165 5.49 56.385 6.805 ;
        RECT 0 5.485 56.38 5.965 ;
        RECT 46.25 5.43 56.38 6.805 ;
        RECT 46.255 5.43 55.805 7.03 ;
        RECT 52.895 5.43 55.645 7.04 ;
        RECT 47.36 5.43 52.085 7.035 ;
        RECT 47.36 5.425 52.08 7.035 ;
        RECT 46.165 5.485 55.805 6.955 ;
        RECT 46.155 5.49 56.385 6.8 ;
        RECT 28.935 5.485 39.165 6.8 ;
        RECT 29.03 5.43 39.16 6.8 ;
        RECT 30.14 5.425 39.16 6.8 ;
        RECT 29.035 5.43 38.585 7.005 ;
        RECT 29.035 5.43 38.58 7.03 ;
        RECT 35.675 5.425 38.425 7.035 ;
        RECT 30.14 5.425 34.865 7.035 ;
        RECT 28.945 5.485 38.585 6.955 ;
        RECT 0 5.485 21.945 6.8 ;
        RECT 0 5.425 21.94 7 ;
        RECT 0 5.425 21.47 7.025 ;
        RECT 18.455 5.425 21.205 7.035 ;
        RECT 15.045 5.425 17.795 7.035 ;
        RECT 16.97 8.945 17.26 9.175 ;
        RECT 16.8 8.975 17.26 9.145 ;
      LAYER mcon ;
        RECT 17.03 8.975 17.2 9.145 ;
        RECT 17.335 6.835 17.505 7.005 ;
        RECT 20.745 6.835 20.915 7.005 ;
        RECT 21.73 5.64 21.9 5.81 ;
        RECT 22.19 5.64 22.36 5.81 ;
        RECT 22.65 5.64 22.82 5.81 ;
        RECT 23.11 5.64 23.28 5.81 ;
        RECT 23.57 5.64 23.74 5.81 ;
        RECT 24.03 5.64 24.2 5.81 ;
        RECT 24.49 5.64 24.66 5.81 ;
        RECT 24.95 5.64 25.12 5.81 ;
        RECT 25.41 5.64 25.58 5.81 ;
        RECT 25.87 5.64 26.04 5.81 ;
        RECT 26.33 5.64 26.5 5.81 ;
        RECT 26.79 5.64 26.96 5.81 ;
        RECT 27.25 5.64 27.42 5.81 ;
        RECT 27.71 5.64 27.88 5.81 ;
        RECT 28.17 5.64 28.34 5.81 ;
        RECT 28.63 5.64 28.8 5.81 ;
        RECT 32.43 6.835 32.6 7.005 ;
        RECT 32.43 5.455 32.6 5.625 ;
        RECT 33.135 6.835 33.305 7.005 ;
        RECT 33.135 5.455 33.305 5.625 ;
        RECT 34.12 5.455 34.29 5.625 ;
        RECT 34.125 6.835 34.295 7.005 ;
        RECT 37.965 6.835 38.135 7.005 ;
        RECT 38.95 5.64 39.12 5.81 ;
        RECT 39.41 5.64 39.58 5.81 ;
        RECT 39.87 5.64 40.04 5.81 ;
        RECT 40.33 5.64 40.5 5.81 ;
        RECT 40.79 5.64 40.96 5.81 ;
        RECT 41.25 5.64 41.42 5.81 ;
        RECT 41.71 5.64 41.88 5.81 ;
        RECT 42.17 5.64 42.34 5.81 ;
        RECT 42.63 5.64 42.8 5.81 ;
        RECT 43.09 5.64 43.26 5.81 ;
        RECT 43.55 5.64 43.72 5.81 ;
        RECT 44.01 5.64 44.18 5.81 ;
        RECT 44.47 5.64 44.64 5.81 ;
        RECT 44.93 5.64 45.1 5.81 ;
        RECT 45.39 5.64 45.56 5.81 ;
        RECT 45.85 5.64 46.02 5.81 ;
        RECT 49.65 6.835 49.82 7.005 ;
        RECT 49.65 5.455 49.82 5.625 ;
        RECT 50.355 6.835 50.525 7.005 ;
        RECT 50.355 5.455 50.525 5.625 ;
        RECT 51.34 5.455 51.51 5.625 ;
        RECT 51.345 6.835 51.515 7.005 ;
        RECT 55.185 6.84 55.355 7.01 ;
        RECT 56.17 5.645 56.34 5.815 ;
        RECT 56.63 5.645 56.8 5.815 ;
        RECT 57.09 5.645 57.26 5.815 ;
        RECT 57.55 5.645 57.72 5.815 ;
        RECT 58.01 5.645 58.18 5.815 ;
        RECT 58.47 5.645 58.64 5.815 ;
        RECT 58.93 5.645 59.1 5.815 ;
        RECT 59.39 5.645 59.56 5.815 ;
        RECT 59.85 5.645 60.02 5.815 ;
        RECT 60.31 5.645 60.48 5.815 ;
        RECT 60.77 5.645 60.94 5.815 ;
        RECT 61.23 5.645 61.4 5.815 ;
        RECT 61.69 5.645 61.86 5.815 ;
        RECT 62.15 5.645 62.32 5.815 ;
        RECT 62.61 5.645 62.78 5.815 ;
        RECT 63.07 5.645 63.24 5.815 ;
        RECT 66.87 6.84 67.04 7.01 ;
        RECT 66.87 5.46 67.04 5.63 ;
        RECT 67.575 6.84 67.745 7.01 ;
        RECT 67.575 5.46 67.745 5.63 ;
        RECT 68.56 5.46 68.73 5.63 ;
        RECT 68.565 6.84 68.735 7.01 ;
        RECT 72.405 6.835 72.575 7.005 ;
        RECT 73.39 5.64 73.56 5.81 ;
        RECT 73.85 5.64 74.02 5.81 ;
        RECT 74.31 5.64 74.48 5.81 ;
        RECT 74.77 5.64 74.94 5.81 ;
        RECT 75.23 5.64 75.4 5.81 ;
        RECT 75.69 5.64 75.86 5.81 ;
        RECT 76.15 5.64 76.32 5.81 ;
        RECT 76.61 5.64 76.78 5.81 ;
        RECT 77.07 5.64 77.24 5.81 ;
        RECT 77.53 5.64 77.7 5.81 ;
        RECT 77.99 5.64 78.16 5.81 ;
        RECT 78.45 5.64 78.62 5.81 ;
        RECT 78.91 5.64 79.08 5.81 ;
        RECT 79.37 5.64 79.54 5.81 ;
        RECT 79.83 5.64 80 5.81 ;
        RECT 80.29 5.64 80.46 5.81 ;
        RECT 84.09 6.835 84.26 7.005 ;
        RECT 84.09 5.455 84.26 5.625 ;
        RECT 84.795 6.835 84.965 7.005 ;
        RECT 84.795 5.455 84.965 5.625 ;
        RECT 85.78 5.455 85.95 5.625 ;
        RECT 85.785 6.835 85.955 7.005 ;
        RECT 89.625 6.835 89.795 7.005 ;
        RECT 90.61 5.64 90.78 5.81 ;
        RECT 91.07 5.64 91.24 5.81 ;
        RECT 91.53 5.64 91.7 5.81 ;
        RECT 91.99 5.64 92.16 5.81 ;
        RECT 92.45 5.64 92.62 5.81 ;
        RECT 92.91 5.64 93.08 5.81 ;
        RECT 93.37 5.64 93.54 5.81 ;
        RECT 93.83 5.64 94 5.81 ;
        RECT 94.29 5.64 94.46 5.81 ;
        RECT 94.75 5.64 94.92 5.81 ;
        RECT 95.21 5.64 95.38 5.81 ;
        RECT 95.67 5.64 95.84 5.81 ;
        RECT 96.13 5.64 96.3 5.81 ;
        RECT 96.59 5.64 96.76 5.81 ;
        RECT 97.05 5.64 97.22 5.81 ;
        RECT 97.51 5.64 97.68 5.81 ;
        RECT 101.31 6.835 101.48 7.005 ;
        RECT 101.31 5.455 101.48 5.625 ;
        RECT 102.015 6.835 102.185 7.005 ;
        RECT 102.015 5.455 102.185 5.625 ;
        RECT 103 5.455 103.17 5.625 ;
        RECT 103.005 6.835 103.175 7.005 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 92.85 7.085 93.18 7.415 ;
        RECT 92.38 7.1 93.18 7.4 ;
        RECT 75.63 7.085 75.96 7.415 ;
        RECT 75.16 7.1 75.96 7.4 ;
        RECT 58.41 7.09 58.74 7.42 ;
        RECT 57.94 7.105 58.74 7.405 ;
        RECT 41.19 7.085 41.52 7.415 ;
        RECT 40.72 7.1 41.52 7.4 ;
        RECT 23.97 7.085 24.3 7.415 ;
        RECT 23.5 7.1 24.3 7.4 ;
      LAYER met2 ;
        RECT 92.875 7.065 93.155 7.435 ;
        RECT 75.655 7.065 75.935 7.435 ;
        RECT 58.435 7.07 58.715 7.44 ;
        RECT 41.215 7.065 41.495 7.435 ;
        RECT 23.995 7.065 24.275 7.435 ;
      LAYER li1 ;
        RECT 0.045 0 103.915 1.6 ;
        RECT 102.92 0 103.09 2.225 ;
        RECT 101.935 0 102.105 2.225 ;
        RECT 99.19 0 99.36 2.225 ;
        RECT 90.46 0 98.12 3.09 ;
        RECT 97.36 0 97.69 3.48 ;
        RECT 96.52 0 96.85 3.48 ;
        RECT 94.69 0 94.98 3.925 ;
        RECT 94.24 0 94.51 3.9 ;
        RECT 93.33 0 93.57 3.9 ;
        RECT 92.88 0 93.12 3.9 ;
        RECT 91.94 0 92.21 3.9 ;
        RECT 91.49 0 91.72 3.91 ;
        RECT 90.61 0 90.82 3.91 ;
        RECT 85.7 0 85.87 2.225 ;
        RECT 84.715 0 84.885 2.225 ;
        RECT 81.97 0 82.14 2.225 ;
        RECT 73.24 0 80.9 3.09 ;
        RECT 80.14 0 80.47 3.48 ;
        RECT 79.3 0 79.63 3.48 ;
        RECT 77.47 0 77.76 3.925 ;
        RECT 77.02 0 77.29 3.9 ;
        RECT 76.11 0 76.35 3.9 ;
        RECT 75.66 0 75.9 3.9 ;
        RECT 74.72 0 74.99 3.9 ;
        RECT 74.27 0 74.5 3.91 ;
        RECT 73.39 0 73.6 3.91 ;
        RECT 52.235 0 69.475 1.605 ;
        RECT 68.48 0 68.65 2.23 ;
        RECT 67.495 0 67.665 2.23 ;
        RECT 64.75 0 64.92 2.23 ;
        RECT 56.02 0 63.68 3.095 ;
        RECT 62.92 0 63.25 3.485 ;
        RECT 62.08 0 62.41 3.485 ;
        RECT 60.25 0 60.54 3.93 ;
        RECT 59.8 0 60.07 3.905 ;
        RECT 58.89 0 59.13 3.905 ;
        RECT 58.44 0 58.68 3.905 ;
        RECT 57.5 0 57.77 3.905 ;
        RECT 57.05 0 57.28 3.915 ;
        RECT 56.17 0 56.38 3.915 ;
        RECT 51.26 0 51.43 2.225 ;
        RECT 50.275 0 50.445 2.225 ;
        RECT 47.53 0 47.7 2.225 ;
        RECT 38.8 0 46.46 3.09 ;
        RECT 45.7 0 46.03 3.48 ;
        RECT 44.86 0 45.19 3.48 ;
        RECT 43.03 0 43.32 3.925 ;
        RECT 42.58 0 42.85 3.9 ;
        RECT 41.67 0 41.91 3.9 ;
        RECT 41.22 0 41.46 3.9 ;
        RECT 40.28 0 40.55 3.9 ;
        RECT 39.83 0 40.06 3.91 ;
        RECT 38.95 0 39.16 3.91 ;
        RECT 34.04 0 34.21 2.225 ;
        RECT 33.055 0 33.225 2.225 ;
        RECT 30.31 0 30.48 2.225 ;
        RECT 21.58 0 29.24 3.09 ;
        RECT 28.48 0 28.81 3.48 ;
        RECT 27.64 0 27.97 3.48 ;
        RECT 25.81 0 26.1 3.925 ;
        RECT 25.36 0 25.63 3.9 ;
        RECT 24.45 0 24.69 3.9 ;
        RECT 24 0 24.24 3.9 ;
        RECT 23.06 0 23.33 3.9 ;
        RECT 22.61 0 22.84 3.91 ;
        RECT 21.73 0 21.94 3.91 ;
        RECT 0.045 10.86 103.915 12.46 ;
        RECT 102.925 10.235 103.095 12.46 ;
        RECT 101.935 10.235 102.105 12.46 ;
        RECT 99.19 10.235 99.36 12.46 ;
        RECT 90.465 8.36 97.825 12.46 ;
        RECT 96.97 7.56 97.28 12.46 ;
        RECT 95.59 7.56 95.9 12.46 ;
        RECT 93.32 7.12 93.655 7.39 ;
        RECT 93.31 7.56 93.62 12.46 ;
        RECT 92.93 7.17 93.655 7.34 ;
        RECT 92.94 7.17 93.11 12.46 ;
        RECT 91.01 7.56 91.32 12.46 ;
        RECT 87.505 10.235 87.675 12.46 ;
        RECT 85.705 10.235 85.875 12.46 ;
        RECT 84.715 10.235 84.885 12.46 ;
        RECT 81.97 10.235 82.14 12.46 ;
        RECT 73.245 8.36 80.605 12.46 ;
        RECT 79.75 7.56 80.06 12.46 ;
        RECT 78.37 7.56 78.68 12.46 ;
        RECT 76.1 7.12 76.435 7.39 ;
        RECT 76.09 7.56 76.4 12.46 ;
        RECT 75.71 7.17 76.435 7.34 ;
        RECT 75.72 7.17 75.89 12.46 ;
        RECT 73.79 7.56 74.1 12.46 ;
        RECT 70.285 10.235 70.455 12.46 ;
        RECT 52.235 10.86 69.475 12.465 ;
        RECT 68.485 10.24 68.655 12.465 ;
        RECT 67.495 10.24 67.665 12.465 ;
        RECT 64.75 10.24 64.92 12.465 ;
        RECT 56.025 8.365 63.385 12.465 ;
        RECT 62.53 7.565 62.84 12.465 ;
        RECT 61.15 7.565 61.46 12.465 ;
        RECT 58.88 7.125 59.215 7.395 ;
        RECT 58.87 7.565 59.18 12.465 ;
        RECT 58.49 7.175 59.215 7.345 ;
        RECT 58.5 7.175 58.67 12.465 ;
        RECT 56.57 7.565 56.88 12.465 ;
        RECT 53.065 10.24 53.235 12.465 ;
        RECT 51.265 10.235 51.435 12.46 ;
        RECT 50.275 10.235 50.445 12.46 ;
        RECT 47.53 10.235 47.7 12.46 ;
        RECT 38.805 8.36 46.165 12.46 ;
        RECT 45.31 7.56 45.62 12.46 ;
        RECT 43.93 7.56 44.24 12.46 ;
        RECT 41.66 7.12 41.995 7.39 ;
        RECT 41.65 7.56 41.96 12.46 ;
        RECT 41.27 7.17 41.995 7.34 ;
        RECT 41.28 7.17 41.45 12.46 ;
        RECT 39.35 7.56 39.66 12.46 ;
        RECT 35.845 10.235 36.015 12.46 ;
        RECT 34.045 10.235 34.215 12.46 ;
        RECT 33.055 10.235 33.225 12.46 ;
        RECT 30.31 10.235 30.48 12.46 ;
        RECT 21.585 8.36 28.945 12.46 ;
        RECT 28.09 7.56 28.4 12.46 ;
        RECT 26.71 7.56 27.02 12.46 ;
        RECT 24.44 7.12 24.775 7.39 ;
        RECT 24.43 7.56 24.74 12.46 ;
        RECT 24.05 7.17 24.775 7.34 ;
        RECT 24.06 7.17 24.23 12.46 ;
        RECT 22.13 7.56 22.44 12.46 ;
        RECT 18.625 10.235 18.795 12.46 ;
        RECT 15.215 10.235 15.385 12.46 ;
        RECT 91.02 7.12 91.355 7.39 ;
        RECT 90.55 7.17 91.355 7.34 ;
        RECT 88.52 8.365 88.69 10.315 ;
        RECT 88.46 10.145 88.63 10.595 ;
        RECT 88.46 7.305 88.63 8.535 ;
        RECT 73.8 7.12 74.135 7.39 ;
        RECT 73.33 7.17 74.135 7.34 ;
        RECT 71.3 8.365 71.47 10.315 ;
        RECT 71.24 10.145 71.41 10.595 ;
        RECT 71.24 7.305 71.41 8.535 ;
        RECT 56.58 7.125 56.915 7.395 ;
        RECT 56.11 7.175 56.915 7.345 ;
        RECT 54.08 8.37 54.25 10.32 ;
        RECT 54.02 10.15 54.19 10.6 ;
        RECT 54.02 7.31 54.19 8.54 ;
        RECT 39.36 7.12 39.695 7.39 ;
        RECT 38.89 7.17 39.695 7.34 ;
        RECT 36.86 8.365 37.03 10.315 ;
        RECT 36.8 10.145 36.97 10.595 ;
        RECT 36.8 7.305 36.97 8.535 ;
        RECT 22.14 7.12 22.475 7.39 ;
        RECT 21.67 7.17 22.475 7.34 ;
        RECT 19.64 8.365 19.81 10.315 ;
        RECT 19.58 10.145 19.75 10.595 ;
        RECT 19.58 7.305 19.75 8.535 ;
      LAYER met1 ;
        RECT 0.045 0 103.915 1.6 ;
        RECT 90.46 0 98.12 3.12 ;
        RECT 73.24 0 80.9 3.12 ;
        RECT 52.235 0 69.475 1.605 ;
        RECT 56.02 0 63.68 3.125 ;
        RECT 38.8 0 46.46 3.12 ;
        RECT 21.58 0 29.24 3.12 ;
        RECT 0.045 10.86 103.915 12.46 ;
        RECT 90.465 8.33 97.825 12.46 ;
        RECT 88.46 8.575 88.75 8.805 ;
        RECT 88.055 8.6 88.75 8.775 ;
        RECT 88.055 8.6 88.225 12.46 ;
        RECT 73.245 8.33 80.605 12.46 ;
        RECT 71.24 8.575 71.53 8.805 ;
        RECT 70.835 8.6 71.53 8.775 ;
        RECT 70.835 8.6 71.005 12.46 ;
        RECT 52.235 10.86 69.475 12.465 ;
        RECT 56.025 8.335 63.385 12.465 ;
        RECT 54.02 8.58 54.31 8.81 ;
        RECT 53.615 8.605 54.31 8.78 ;
        RECT 53.615 8.605 53.785 12.465 ;
        RECT 38.805 8.33 46.165 12.46 ;
        RECT 36.8 8.575 37.09 8.805 ;
        RECT 36.395 8.6 37.09 8.775 ;
        RECT 36.395 8.6 36.565 12.46 ;
        RECT 21.585 8.33 28.945 12.46 ;
        RECT 19.58 8.575 19.87 8.805 ;
        RECT 19.175 8.6 19.87 8.775 ;
        RECT 19.175 8.6 19.345 12.46 ;
        RECT 92.855 7.125 93.175 7.385 ;
        RECT 90.49 7.185 93.175 7.325 ;
        RECT 90.49 7.14 90.78 7.37 ;
        RECT 75.635 7.125 75.955 7.385 ;
        RECT 73.27 7.185 75.955 7.325 ;
        RECT 73.27 7.14 73.56 7.37 ;
        RECT 58.415 7.13 58.735 7.39 ;
        RECT 56.05 7.19 58.735 7.33 ;
        RECT 56.05 7.145 56.34 7.375 ;
        RECT 41.195 7.125 41.515 7.385 ;
        RECT 38.83 7.185 41.515 7.325 ;
        RECT 38.83 7.14 39.12 7.37 ;
        RECT 23.975 7.125 24.295 7.385 ;
        RECT 21.61 7.185 24.295 7.325 ;
        RECT 21.61 7.14 21.9 7.37 ;
      LAYER via1 ;
        RECT 24.06 7.18 24.21 7.33 ;
        RECT 41.28 7.18 41.43 7.33 ;
        RECT 58.5 7.185 58.65 7.335 ;
        RECT 75.72 7.18 75.87 7.33 ;
        RECT 92.94 7.18 93.09 7.33 ;
      LAYER via2 ;
        RECT 24.035 7.15 24.235 7.35 ;
        RECT 41.255 7.15 41.455 7.35 ;
        RECT 58.475 7.155 58.675 7.355 ;
        RECT 75.695 7.15 75.895 7.35 ;
        RECT 92.915 7.15 93.115 7.35 ;
      LAYER mcon ;
        RECT 15.295 10.895 15.465 11.065 ;
        RECT 15.975 10.895 16.145 11.065 ;
        RECT 16.655 10.895 16.825 11.065 ;
        RECT 17.335 10.895 17.505 11.065 ;
        RECT 18.705 10.895 18.875 11.065 ;
        RECT 19.385 10.895 19.555 11.065 ;
        RECT 19.64 8.605 19.81 8.775 ;
        RECT 20.065 10.895 20.235 11.065 ;
        RECT 20.745 10.895 20.915 11.065 ;
        RECT 21.67 7.17 21.84 7.34 ;
        RECT 21.73 8.36 21.9 8.53 ;
        RECT 21.73 2.92 21.9 3.09 ;
        RECT 22.19 8.36 22.36 8.53 ;
        RECT 22.19 2.92 22.36 3.09 ;
        RECT 22.65 8.36 22.82 8.53 ;
        RECT 22.65 2.92 22.82 3.09 ;
        RECT 23.11 8.36 23.28 8.53 ;
        RECT 23.11 2.92 23.28 3.09 ;
        RECT 23.57 8.36 23.74 8.53 ;
        RECT 23.57 2.92 23.74 3.09 ;
        RECT 24.03 8.36 24.2 8.53 ;
        RECT 24.03 2.92 24.2 3.09 ;
        RECT 24.05 7.17 24.22 7.34 ;
        RECT 24.49 8.36 24.66 8.53 ;
        RECT 24.49 2.92 24.66 3.09 ;
        RECT 24.95 8.36 25.12 8.53 ;
        RECT 24.95 2.92 25.12 3.09 ;
        RECT 25.41 8.36 25.58 8.53 ;
        RECT 25.41 2.92 25.58 3.09 ;
        RECT 25.87 8.36 26.04 8.53 ;
        RECT 25.87 2.92 26.04 3.09 ;
        RECT 26.33 8.36 26.5 8.53 ;
        RECT 26.33 2.92 26.5 3.09 ;
        RECT 26.79 8.36 26.96 8.53 ;
        RECT 26.79 2.92 26.96 3.09 ;
        RECT 27.25 8.36 27.42 8.53 ;
        RECT 27.25 2.92 27.42 3.09 ;
        RECT 27.71 8.36 27.88 8.53 ;
        RECT 27.71 2.92 27.88 3.09 ;
        RECT 28.17 8.36 28.34 8.53 ;
        RECT 28.17 2.92 28.34 3.09 ;
        RECT 28.63 8.36 28.8 8.53 ;
        RECT 28.63 2.92 28.8 3.09 ;
        RECT 30.39 10.895 30.56 11.065 ;
        RECT 30.39 1.395 30.56 1.565 ;
        RECT 31.07 10.895 31.24 11.065 ;
        RECT 31.07 1.395 31.24 1.565 ;
        RECT 31.75 10.895 31.92 11.065 ;
        RECT 31.75 1.395 31.92 1.565 ;
        RECT 32.43 10.895 32.6 11.065 ;
        RECT 32.43 1.395 32.6 1.565 ;
        RECT 33.135 10.895 33.305 11.065 ;
        RECT 33.135 1.395 33.305 1.565 ;
        RECT 34.12 1.395 34.29 1.565 ;
        RECT 34.125 10.895 34.295 11.065 ;
        RECT 35.925 10.895 36.095 11.065 ;
        RECT 36.605 10.895 36.775 11.065 ;
        RECT 36.86 8.605 37.03 8.775 ;
        RECT 37.285 10.895 37.455 11.065 ;
        RECT 37.965 10.895 38.135 11.065 ;
        RECT 38.89 7.17 39.06 7.34 ;
        RECT 38.95 8.36 39.12 8.53 ;
        RECT 38.95 2.92 39.12 3.09 ;
        RECT 39.41 8.36 39.58 8.53 ;
        RECT 39.41 2.92 39.58 3.09 ;
        RECT 39.87 8.36 40.04 8.53 ;
        RECT 39.87 2.92 40.04 3.09 ;
        RECT 40.33 8.36 40.5 8.53 ;
        RECT 40.33 2.92 40.5 3.09 ;
        RECT 40.79 8.36 40.96 8.53 ;
        RECT 40.79 2.92 40.96 3.09 ;
        RECT 41.25 8.36 41.42 8.53 ;
        RECT 41.25 2.92 41.42 3.09 ;
        RECT 41.27 7.17 41.44 7.34 ;
        RECT 41.71 8.36 41.88 8.53 ;
        RECT 41.71 2.92 41.88 3.09 ;
        RECT 42.17 8.36 42.34 8.53 ;
        RECT 42.17 2.92 42.34 3.09 ;
        RECT 42.63 8.36 42.8 8.53 ;
        RECT 42.63 2.92 42.8 3.09 ;
        RECT 43.09 8.36 43.26 8.53 ;
        RECT 43.09 2.92 43.26 3.09 ;
        RECT 43.55 8.36 43.72 8.53 ;
        RECT 43.55 2.92 43.72 3.09 ;
        RECT 44.01 8.36 44.18 8.53 ;
        RECT 44.01 2.92 44.18 3.09 ;
        RECT 44.47 8.36 44.64 8.53 ;
        RECT 44.47 2.92 44.64 3.09 ;
        RECT 44.93 8.36 45.1 8.53 ;
        RECT 44.93 2.92 45.1 3.09 ;
        RECT 45.39 8.36 45.56 8.53 ;
        RECT 45.39 2.92 45.56 3.09 ;
        RECT 45.85 8.36 46.02 8.53 ;
        RECT 45.85 2.92 46.02 3.09 ;
        RECT 47.61 10.895 47.78 11.065 ;
        RECT 47.61 1.395 47.78 1.565 ;
        RECT 48.29 10.895 48.46 11.065 ;
        RECT 48.29 1.395 48.46 1.565 ;
        RECT 48.97 10.895 49.14 11.065 ;
        RECT 48.97 1.395 49.14 1.565 ;
        RECT 49.65 10.895 49.82 11.065 ;
        RECT 49.65 1.395 49.82 1.565 ;
        RECT 50.355 10.895 50.525 11.065 ;
        RECT 50.355 1.395 50.525 1.565 ;
        RECT 51.34 1.395 51.51 1.565 ;
        RECT 51.345 10.895 51.515 11.065 ;
        RECT 53.145 10.9 53.315 11.07 ;
        RECT 53.825 10.9 53.995 11.07 ;
        RECT 54.08 8.61 54.25 8.78 ;
        RECT 54.505 10.9 54.675 11.07 ;
        RECT 55.185 10.9 55.355 11.07 ;
        RECT 56.11 7.175 56.28 7.345 ;
        RECT 56.17 8.365 56.34 8.535 ;
        RECT 56.17 2.925 56.34 3.095 ;
        RECT 56.63 8.365 56.8 8.535 ;
        RECT 56.63 2.925 56.8 3.095 ;
        RECT 57.09 8.365 57.26 8.535 ;
        RECT 57.09 2.925 57.26 3.095 ;
        RECT 57.55 8.365 57.72 8.535 ;
        RECT 57.55 2.925 57.72 3.095 ;
        RECT 58.01 8.365 58.18 8.535 ;
        RECT 58.01 2.925 58.18 3.095 ;
        RECT 58.47 8.365 58.64 8.535 ;
        RECT 58.47 2.925 58.64 3.095 ;
        RECT 58.49 7.175 58.66 7.345 ;
        RECT 58.93 8.365 59.1 8.535 ;
        RECT 58.93 2.925 59.1 3.095 ;
        RECT 59.39 8.365 59.56 8.535 ;
        RECT 59.39 2.925 59.56 3.095 ;
        RECT 59.85 8.365 60.02 8.535 ;
        RECT 59.85 2.925 60.02 3.095 ;
        RECT 60.31 8.365 60.48 8.535 ;
        RECT 60.31 2.925 60.48 3.095 ;
        RECT 60.77 8.365 60.94 8.535 ;
        RECT 60.77 2.925 60.94 3.095 ;
        RECT 61.23 8.365 61.4 8.535 ;
        RECT 61.23 2.925 61.4 3.095 ;
        RECT 61.69 8.365 61.86 8.535 ;
        RECT 61.69 2.925 61.86 3.095 ;
        RECT 62.15 8.365 62.32 8.535 ;
        RECT 62.15 2.925 62.32 3.095 ;
        RECT 62.61 8.365 62.78 8.535 ;
        RECT 62.61 2.925 62.78 3.095 ;
        RECT 63.07 8.365 63.24 8.535 ;
        RECT 63.07 2.925 63.24 3.095 ;
        RECT 64.83 10.9 65 11.07 ;
        RECT 64.83 1.4 65 1.57 ;
        RECT 65.51 10.9 65.68 11.07 ;
        RECT 65.51 1.4 65.68 1.57 ;
        RECT 66.19 10.9 66.36 11.07 ;
        RECT 66.19 1.4 66.36 1.57 ;
        RECT 66.87 10.9 67.04 11.07 ;
        RECT 66.87 1.4 67.04 1.57 ;
        RECT 67.575 10.9 67.745 11.07 ;
        RECT 67.575 1.4 67.745 1.57 ;
        RECT 68.56 1.4 68.73 1.57 ;
        RECT 68.565 10.9 68.735 11.07 ;
        RECT 70.365 10.895 70.535 11.065 ;
        RECT 71.045 10.895 71.215 11.065 ;
        RECT 71.3 8.605 71.47 8.775 ;
        RECT 71.725 10.895 71.895 11.065 ;
        RECT 72.405 10.895 72.575 11.065 ;
        RECT 73.33 7.17 73.5 7.34 ;
        RECT 73.39 8.36 73.56 8.53 ;
        RECT 73.39 2.92 73.56 3.09 ;
        RECT 73.85 8.36 74.02 8.53 ;
        RECT 73.85 2.92 74.02 3.09 ;
        RECT 74.31 8.36 74.48 8.53 ;
        RECT 74.31 2.92 74.48 3.09 ;
        RECT 74.77 8.36 74.94 8.53 ;
        RECT 74.77 2.92 74.94 3.09 ;
        RECT 75.23 8.36 75.4 8.53 ;
        RECT 75.23 2.92 75.4 3.09 ;
        RECT 75.69 8.36 75.86 8.53 ;
        RECT 75.69 2.92 75.86 3.09 ;
        RECT 75.71 7.17 75.88 7.34 ;
        RECT 76.15 8.36 76.32 8.53 ;
        RECT 76.15 2.92 76.32 3.09 ;
        RECT 76.61 8.36 76.78 8.53 ;
        RECT 76.61 2.92 76.78 3.09 ;
        RECT 77.07 8.36 77.24 8.53 ;
        RECT 77.07 2.92 77.24 3.09 ;
        RECT 77.53 8.36 77.7 8.53 ;
        RECT 77.53 2.92 77.7 3.09 ;
        RECT 77.99 8.36 78.16 8.53 ;
        RECT 77.99 2.92 78.16 3.09 ;
        RECT 78.45 8.36 78.62 8.53 ;
        RECT 78.45 2.92 78.62 3.09 ;
        RECT 78.91 8.36 79.08 8.53 ;
        RECT 78.91 2.92 79.08 3.09 ;
        RECT 79.37 8.36 79.54 8.53 ;
        RECT 79.37 2.92 79.54 3.09 ;
        RECT 79.83 8.36 80 8.53 ;
        RECT 79.83 2.92 80 3.09 ;
        RECT 80.29 8.36 80.46 8.53 ;
        RECT 80.29 2.92 80.46 3.09 ;
        RECT 82.05 10.895 82.22 11.065 ;
        RECT 82.05 1.395 82.22 1.565 ;
        RECT 82.73 10.895 82.9 11.065 ;
        RECT 82.73 1.395 82.9 1.565 ;
        RECT 83.41 10.895 83.58 11.065 ;
        RECT 83.41 1.395 83.58 1.565 ;
        RECT 84.09 10.895 84.26 11.065 ;
        RECT 84.09 1.395 84.26 1.565 ;
        RECT 84.795 10.895 84.965 11.065 ;
        RECT 84.795 1.395 84.965 1.565 ;
        RECT 85.78 1.395 85.95 1.565 ;
        RECT 85.785 10.895 85.955 11.065 ;
        RECT 87.585 10.895 87.755 11.065 ;
        RECT 88.265 10.895 88.435 11.065 ;
        RECT 88.52 8.605 88.69 8.775 ;
        RECT 88.945 10.895 89.115 11.065 ;
        RECT 89.625 10.895 89.795 11.065 ;
        RECT 90.55 7.17 90.72 7.34 ;
        RECT 90.61 8.36 90.78 8.53 ;
        RECT 90.61 2.92 90.78 3.09 ;
        RECT 91.07 8.36 91.24 8.53 ;
        RECT 91.07 2.92 91.24 3.09 ;
        RECT 91.53 8.36 91.7 8.53 ;
        RECT 91.53 2.92 91.7 3.09 ;
        RECT 91.99 8.36 92.16 8.53 ;
        RECT 91.99 2.92 92.16 3.09 ;
        RECT 92.45 8.36 92.62 8.53 ;
        RECT 92.45 2.92 92.62 3.09 ;
        RECT 92.91 8.36 93.08 8.53 ;
        RECT 92.91 2.92 93.08 3.09 ;
        RECT 92.93 7.17 93.1 7.34 ;
        RECT 93.37 8.36 93.54 8.53 ;
        RECT 93.37 2.92 93.54 3.09 ;
        RECT 93.83 8.36 94 8.53 ;
        RECT 93.83 2.92 94 3.09 ;
        RECT 94.29 8.36 94.46 8.53 ;
        RECT 94.29 2.92 94.46 3.09 ;
        RECT 94.75 8.36 94.92 8.53 ;
        RECT 94.75 2.92 94.92 3.09 ;
        RECT 95.21 8.36 95.38 8.53 ;
        RECT 95.21 2.92 95.38 3.09 ;
        RECT 95.67 8.36 95.84 8.53 ;
        RECT 95.67 2.92 95.84 3.09 ;
        RECT 96.13 8.36 96.3 8.53 ;
        RECT 96.13 2.92 96.3 3.09 ;
        RECT 96.59 8.36 96.76 8.53 ;
        RECT 96.59 2.92 96.76 3.09 ;
        RECT 97.05 8.36 97.22 8.53 ;
        RECT 97.05 2.92 97.22 3.09 ;
        RECT 97.51 8.36 97.68 8.53 ;
        RECT 97.51 2.92 97.68 3.09 ;
        RECT 99.27 10.895 99.44 11.065 ;
        RECT 99.27 1.395 99.44 1.565 ;
        RECT 99.95 10.895 100.12 11.065 ;
        RECT 99.95 1.395 100.12 1.565 ;
        RECT 100.63 10.895 100.8 11.065 ;
        RECT 100.63 1.395 100.8 1.565 ;
        RECT 101.31 10.895 101.48 11.065 ;
        RECT 101.31 1.395 101.48 1.565 ;
        RECT 102.015 10.895 102.185 11.065 ;
        RECT 102.015 1.395 102.185 1.565 ;
        RECT 103 1.395 103.17 1.565 ;
        RECT 103.005 10.895 103.175 11.065 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 88.795 9.285 89.165 9.655 ;
      RECT 88.795 9.32 95.945 9.62 ;
      RECT 95.645 7.1 95.945 9.62 ;
      RECT 94.59 7.08 94.89 9.62 ;
      RECT 93.56 7.745 93.86 9.62 ;
      RECT 93.06 7.79 93.86 8.09 ;
      RECT 93.44 7.72 93.74 8.09 ;
      RECT 95.57 7.1 95.945 7.465 ;
      RECT 95.635 7.06 95.935 7.465 ;
      RECT 94.55 7.08 94.89 7.43 ;
      RECT 94.565 7.04 94.865 7.43 ;
      RECT 94.54 7.085 94.89 7.415 ;
      RECT 95.57 7.1 96.38 7.4 ;
      RECT 94.07 7.1 94.89 7.4 ;
      RECT 95.58 7.085 95.935 7.465 ;
      RECT 95.23 5.05 95.56 5.38 ;
      RECT 95.23 5.065 96.03 5.365 ;
      RECT 95.245 5.02 95.545 5.38 ;
      RECT 94.89 4.37 95.22 4.7 ;
      RECT 94.89 4.385 95.69 4.685 ;
      RECT 94.975 4.36 95.275 4.685 ;
      RECT 94.21 5.45 94.54 5.78 ;
      RECT 92.17 5.45 92.5 5.78 ;
      RECT 92.17 5.465 94.54 5.765 ;
      RECT 93.86 4.71 94.19 5.04 ;
      RECT 93.4 4.725 94.2 5.025 ;
      RECT 93.53 3.52 93.86 3.85 ;
      RECT 93.06 3.535 93.86 3.835 ;
      RECT 93.52 3.53 93.86 3.835 ;
      RECT 71.575 9.285 71.945 9.655 ;
      RECT 71.575 9.32 78.725 9.62 ;
      RECT 78.425 7.1 78.725 9.62 ;
      RECT 77.37 7.08 77.67 9.62 ;
      RECT 76.34 7.745 76.64 9.62 ;
      RECT 75.84 7.79 76.64 8.09 ;
      RECT 76.22 7.72 76.52 8.09 ;
      RECT 78.35 7.1 78.725 7.465 ;
      RECT 78.415 7.06 78.715 7.465 ;
      RECT 77.33 7.08 77.67 7.43 ;
      RECT 77.345 7.04 77.645 7.43 ;
      RECT 77.32 7.085 77.67 7.415 ;
      RECT 78.35 7.1 79.16 7.4 ;
      RECT 76.85 7.1 77.67 7.4 ;
      RECT 78.36 7.085 78.715 7.465 ;
      RECT 78.01 5.05 78.34 5.38 ;
      RECT 78.01 5.065 78.81 5.365 ;
      RECT 78.025 5.02 78.325 5.38 ;
      RECT 77.67 4.37 78 4.7 ;
      RECT 77.67 4.385 78.47 4.685 ;
      RECT 77.755 4.36 78.055 4.685 ;
      RECT 76.99 5.45 77.32 5.78 ;
      RECT 74.95 5.45 75.28 5.78 ;
      RECT 74.95 5.465 77.32 5.765 ;
      RECT 76.64 4.71 76.97 5.04 ;
      RECT 76.18 4.725 76.98 5.025 ;
      RECT 76.31 3.52 76.64 3.85 ;
      RECT 75.84 3.535 76.64 3.835 ;
      RECT 76.3 3.53 76.64 3.835 ;
      RECT 54.355 9.29 54.725 9.66 ;
      RECT 54.355 9.325 61.505 9.625 ;
      RECT 61.205 7.105 61.505 9.625 ;
      RECT 60.15 7.085 60.45 9.625 ;
      RECT 59.12 7.75 59.42 9.625 ;
      RECT 58.62 7.795 59.42 8.095 ;
      RECT 59 7.725 59.3 8.095 ;
      RECT 61.13 7.105 61.505 7.47 ;
      RECT 61.195 7.065 61.495 7.47 ;
      RECT 60.11 7.085 60.45 7.435 ;
      RECT 60.125 7.045 60.425 7.435 ;
      RECT 60.1 7.09 60.45 7.42 ;
      RECT 61.13 7.105 61.94 7.405 ;
      RECT 59.63 7.105 60.45 7.405 ;
      RECT 61.14 7.09 61.495 7.47 ;
      RECT 60.79 5.055 61.12 5.385 ;
      RECT 60.79 5.07 61.59 5.37 ;
      RECT 60.805 5.025 61.105 5.385 ;
      RECT 60.45 4.375 60.78 4.705 ;
      RECT 60.45 4.39 61.25 4.69 ;
      RECT 60.535 4.365 60.835 4.69 ;
      RECT 59.77 5.455 60.1 5.785 ;
      RECT 57.73 5.455 58.06 5.785 ;
      RECT 57.73 5.47 60.1 5.77 ;
      RECT 59.42 4.715 59.75 5.045 ;
      RECT 58.96 4.73 59.76 5.03 ;
      RECT 59.09 3.525 59.42 3.855 ;
      RECT 58.62 3.54 59.42 3.84 ;
      RECT 59.08 3.535 59.42 3.84 ;
      RECT 37.135 9.285 37.505 9.655 ;
      RECT 37.135 9.32 44.285 9.62 ;
      RECT 43.985 7.1 44.285 9.62 ;
      RECT 42.93 7.08 43.23 9.62 ;
      RECT 41.9 7.745 42.2 9.62 ;
      RECT 41.4 7.79 42.2 8.09 ;
      RECT 41.78 7.72 42.08 8.09 ;
      RECT 43.91 7.1 44.285 7.465 ;
      RECT 43.975 7.06 44.275 7.465 ;
      RECT 42.89 7.08 43.23 7.43 ;
      RECT 42.905 7.04 43.205 7.43 ;
      RECT 42.88 7.085 43.23 7.415 ;
      RECT 43.91 7.1 44.72 7.4 ;
      RECT 42.41 7.1 43.23 7.4 ;
      RECT 43.92 7.085 44.275 7.465 ;
      RECT 43.57 5.05 43.9 5.38 ;
      RECT 43.57 5.065 44.37 5.365 ;
      RECT 43.585 5.02 43.885 5.38 ;
      RECT 43.23 4.37 43.56 4.7 ;
      RECT 43.23 4.385 44.03 4.685 ;
      RECT 43.315 4.36 43.615 4.685 ;
      RECT 42.55 5.45 42.88 5.78 ;
      RECT 40.51 5.45 40.84 5.78 ;
      RECT 40.51 5.465 42.88 5.765 ;
      RECT 42.2 4.71 42.53 5.04 ;
      RECT 41.74 4.725 42.54 5.025 ;
      RECT 41.87 3.52 42.2 3.85 ;
      RECT 41.4 3.535 42.2 3.835 ;
      RECT 41.86 3.53 42.2 3.835 ;
      RECT 19.915 9.285 20.285 9.655 ;
      RECT 19.915 9.32 27.065 9.62 ;
      RECT 26.765 7.1 27.065 9.62 ;
      RECT 25.71 7.08 26.01 9.62 ;
      RECT 24.68 7.745 24.98 9.62 ;
      RECT 24.18 7.79 24.98 8.09 ;
      RECT 24.56 7.72 24.86 8.09 ;
      RECT 26.69 7.1 27.065 7.465 ;
      RECT 26.755 7.06 27.055 7.465 ;
      RECT 25.67 7.08 26.01 7.43 ;
      RECT 25.685 7.04 25.985 7.43 ;
      RECT 25.66 7.085 26.01 7.415 ;
      RECT 26.69 7.1 27.5 7.4 ;
      RECT 25.19 7.1 26.01 7.4 ;
      RECT 26.7 7.085 27.055 7.465 ;
      RECT 26.35 5.05 26.68 5.38 ;
      RECT 26.35 5.065 27.15 5.365 ;
      RECT 26.365 5.02 26.665 5.38 ;
      RECT 26.01 4.37 26.34 4.7 ;
      RECT 26.01 4.385 26.81 4.685 ;
      RECT 26.095 4.36 26.395 4.685 ;
      RECT 25.33 5.45 25.66 5.78 ;
      RECT 23.29 5.45 23.62 5.78 ;
      RECT 23.29 5.465 25.66 5.765 ;
      RECT 24.98 4.71 25.31 5.04 ;
      RECT 24.52 4.725 25.32 5.025 ;
      RECT 24.65 3.52 24.98 3.85 ;
      RECT 24.18 3.535 24.98 3.835 ;
      RECT 24.64 3.53 24.98 3.835 ;
      RECT 103.255 7.2 103.635 12.46 ;
      RECT 86.035 7.2 86.415 12.46 ;
      RECT 68.815 7.205 69.195 12.465 ;
      RECT 51.595 7.2 51.975 12.46 ;
      RECT 34.375 7.2 34.755 12.46 ;
    LAYER via2 ;
      RECT 103.345 7.29 103.545 7.49 ;
      RECT 95.645 7.15 95.845 7.35 ;
      RECT 95.295 5.115 95.495 5.315 ;
      RECT 94.955 4.435 95.155 4.635 ;
      RECT 94.605 7.15 94.805 7.35 ;
      RECT 94.275 5.515 94.475 5.715 ;
      RECT 93.925 4.775 94.125 4.975 ;
      RECT 93.595 3.585 93.795 3.785 ;
      RECT 93.595 7.81 93.795 8.01 ;
      RECT 92.235 5.515 92.435 5.715 ;
      RECT 88.88 9.37 89.08 9.57 ;
      RECT 86.125 7.29 86.325 7.49 ;
      RECT 78.425 7.15 78.625 7.35 ;
      RECT 78.075 5.115 78.275 5.315 ;
      RECT 77.735 4.435 77.935 4.635 ;
      RECT 77.385 7.15 77.585 7.35 ;
      RECT 77.055 5.515 77.255 5.715 ;
      RECT 76.705 4.775 76.905 4.975 ;
      RECT 76.375 3.585 76.575 3.785 ;
      RECT 76.375 7.81 76.575 8.01 ;
      RECT 75.015 5.515 75.215 5.715 ;
      RECT 71.66 9.37 71.86 9.57 ;
      RECT 68.905 7.295 69.105 7.495 ;
      RECT 61.205 7.155 61.405 7.355 ;
      RECT 60.855 5.12 61.055 5.32 ;
      RECT 60.515 4.44 60.715 4.64 ;
      RECT 60.165 7.155 60.365 7.355 ;
      RECT 59.835 5.52 60.035 5.72 ;
      RECT 59.485 4.78 59.685 4.98 ;
      RECT 59.155 3.59 59.355 3.79 ;
      RECT 59.155 7.815 59.355 8.015 ;
      RECT 57.795 5.52 57.995 5.72 ;
      RECT 54.44 9.375 54.64 9.575 ;
      RECT 51.685 7.29 51.885 7.49 ;
      RECT 43.985 7.15 44.185 7.35 ;
      RECT 43.635 5.115 43.835 5.315 ;
      RECT 43.295 4.435 43.495 4.635 ;
      RECT 42.945 7.15 43.145 7.35 ;
      RECT 42.615 5.515 42.815 5.715 ;
      RECT 42.265 4.775 42.465 4.975 ;
      RECT 41.935 3.585 42.135 3.785 ;
      RECT 41.935 7.81 42.135 8.01 ;
      RECT 40.575 5.515 40.775 5.715 ;
      RECT 37.22 9.37 37.42 9.57 ;
      RECT 34.465 7.29 34.665 7.49 ;
      RECT 26.765 7.15 26.965 7.35 ;
      RECT 26.415 5.115 26.615 5.315 ;
      RECT 26.075 4.435 26.275 4.635 ;
      RECT 25.725 7.15 25.925 7.35 ;
      RECT 25.395 5.515 25.595 5.715 ;
      RECT 25.045 4.775 25.245 4.975 ;
      RECT 24.715 3.585 24.915 3.785 ;
      RECT 24.715 7.81 24.915 8.01 ;
      RECT 23.355 5.515 23.555 5.715 ;
      RECT 20 9.37 20.2 9.57 ;
    LAYER met2 ;
      RECT 16.21 10.055 103.53 10.225 ;
      RECT 103.36 9.585 103.53 10.225 ;
      RECT 16.21 8.54 16.38 10.225 ;
      RECT 103.325 9.585 103.65 9.91 ;
      RECT 16.165 8.54 16.445 8.88 ;
      RECT 100.17 8.565 100.49 8.89 ;
      RECT 100.2 7.98 100.37 8.89 ;
      RECT 100.2 7.98 100.375 8.33 ;
      RECT 100.2 7.98 101.175 8.155 ;
      RECT 101 3.26 101.175 8.155 ;
      RECT 93.555 3.5 93.835 3.87 ;
      RECT 93.555 3.64 98.205 3.815 ;
      RECT 98.03 3.32 98.205 3.815 ;
      RECT 98.5 3.29 98.825 3.615 ;
      RECT 100.945 3.26 101.295 3.61 ;
      RECT 98.03 3.32 101.295 3.49 ;
      RECT 89.32 9.55 100.015 9.72 ;
      RECT 99.855 3.69 100.015 9.72 ;
      RECT 89.32 8.83 89.49 9.72 ;
      RECT 86.14 8.945 86.465 9.27 ;
      RECT 100.97 8.94 101.295 9.265 ;
      RECT 99.855 9.03 101.295 9.2 ;
      RECT 89.27 8.83 89.55 9.17 ;
      RECT 86.14 8.975 86.925 9.145 ;
      RECT 86.925 8.97 89.55 9.14 ;
      RECT 100.17 3.66 100.49 3.98 ;
      RECT 99.855 3.69 100.49 3.86 ;
      RECT 96.625 7.76 96.885 8.095 ;
      RECT 96.685 4.035 96.825 8.095 ;
      RECT 96.625 4.035 96.885 4.355 ;
      RECT 95.945 6.075 96.205 6.395 ;
      RECT 96.005 5.055 96.145 6.395 ;
      RECT 95.945 5.055 96.205 5.375 ;
      RECT 94.925 7.76 95.185 8.095 ;
      RECT 94.895 7.805 95.215 8.05 ;
      RECT 94.985 6.505 95.125 8.095 ;
      RECT 94.305 6.505 95.125 6.645 ;
      RECT 94.305 4.035 94.445 6.645 ;
      RECT 94.235 5.43 94.515 5.8 ;
      RECT 94.245 4.035 94.505 4.355 ;
      RECT 92.195 5.43 92.475 5.8 ;
      RECT 92.265 3.695 92.405 5.8 ;
      RECT 92.205 3.695 92.465 4.015 ;
      RECT 91.525 6.075 91.785 6.395 ;
      RECT 91.585 4.035 91.725 6.395 ;
      RECT 91.525 4.035 91.785 4.355 ;
      RECT 82.95 8.565 83.27 8.89 ;
      RECT 82.98 7.98 83.15 8.89 ;
      RECT 82.98 7.98 83.155 8.33 ;
      RECT 82.98 7.98 83.955 8.155 ;
      RECT 83.78 3.26 83.955 8.155 ;
      RECT 76.335 3.5 76.615 3.87 ;
      RECT 76.335 3.64 80.985 3.815 ;
      RECT 80.81 3.32 80.985 3.815 ;
      RECT 81.28 3.29 81.605 3.615 ;
      RECT 83.725 3.26 84.075 3.61 ;
      RECT 80.81 3.32 84.075 3.49 ;
      RECT 72.1 9.55 82.795 9.72 ;
      RECT 82.635 3.69 82.795 9.72 ;
      RECT 72.1 8.83 72.27 9.72 ;
      RECT 68.92 8.95 69.245 9.275 ;
      RECT 83.75 8.94 84.075 9.265 ;
      RECT 82.635 9.03 84.075 9.2 ;
      RECT 72.05 8.83 72.33 9.17 ;
      RECT 68.92 8.98 69.97 9.15 ;
      RECT 68.92 8.98 70.045 9.145 ;
      RECT 70.045 8.97 72.33 9.14 ;
      RECT 69.97 8.975 72.33 9.14 ;
      RECT 82.95 3.66 83.27 3.98 ;
      RECT 82.635 3.69 83.27 3.86 ;
      RECT 79.405 7.76 79.665 8.095 ;
      RECT 79.465 4.035 79.605 8.095 ;
      RECT 79.405 4.035 79.665 4.355 ;
      RECT 78.725 6.075 78.985 6.395 ;
      RECT 78.785 5.055 78.925 6.395 ;
      RECT 78.725 5.055 78.985 5.375 ;
      RECT 77.705 7.76 77.965 8.095 ;
      RECT 77.675 7.805 77.995 8.05 ;
      RECT 77.765 6.505 77.905 8.095 ;
      RECT 77.085 6.505 77.905 6.645 ;
      RECT 77.085 4.035 77.225 6.645 ;
      RECT 77.015 5.43 77.295 5.8 ;
      RECT 77.025 4.035 77.285 4.355 ;
      RECT 74.975 5.43 75.255 5.8 ;
      RECT 75.045 3.695 75.185 5.8 ;
      RECT 74.985 3.695 75.245 4.015 ;
      RECT 74.305 6.075 74.565 6.395 ;
      RECT 74.365 4.035 74.505 6.395 ;
      RECT 74.305 4.035 74.565 4.355 ;
      RECT 65.73 8.57 66.05 8.895 ;
      RECT 65.76 7.985 65.93 8.895 ;
      RECT 65.76 7.985 65.935 8.335 ;
      RECT 65.76 7.985 66.735 8.16 ;
      RECT 66.56 3.265 66.735 8.16 ;
      RECT 59.115 3.505 59.395 3.875 ;
      RECT 59.115 3.645 63.765 3.82 ;
      RECT 63.59 3.325 63.765 3.82 ;
      RECT 64.06 3.295 64.385 3.62 ;
      RECT 66.505 3.265 66.855 3.615 ;
      RECT 63.59 3.325 66.855 3.495 ;
      RECT 54.88 9.555 65.575 9.725 ;
      RECT 65.415 3.695 65.575 9.725 ;
      RECT 54.88 8.835 55.05 9.725 ;
      RECT 66.53 8.945 66.855 9.27 ;
      RECT 51.7 8.945 52.025 9.27 ;
      RECT 65.415 9.035 66.855 9.205 ;
      RECT 54.83 8.835 55.11 9.175 ;
      RECT 51.7 8.975 52.885 9.145 ;
      RECT 52.885 8.97 55.12 9.14 ;
      RECT 65.73 3.665 66.05 3.985 ;
      RECT 65.415 3.695 66.05 3.865 ;
      RECT 62.185 7.765 62.445 8.1 ;
      RECT 62.245 4.04 62.385 8.1 ;
      RECT 62.185 4.04 62.445 4.36 ;
      RECT 61.505 6.08 61.765 6.4 ;
      RECT 61.565 5.06 61.705 6.4 ;
      RECT 61.505 5.06 61.765 5.38 ;
      RECT 60.485 7.765 60.745 8.1 ;
      RECT 60.455 7.81 60.775 8.055 ;
      RECT 60.545 6.51 60.685 8.1 ;
      RECT 59.865 6.51 60.685 6.65 ;
      RECT 59.865 4.04 60.005 6.65 ;
      RECT 59.795 5.435 60.075 5.805 ;
      RECT 59.805 4.04 60.065 4.36 ;
      RECT 57.755 5.435 58.035 5.805 ;
      RECT 57.825 3.7 57.965 5.805 ;
      RECT 57.765 3.7 58.025 4.02 ;
      RECT 57.085 6.08 57.345 6.4 ;
      RECT 57.145 4.04 57.285 6.4 ;
      RECT 57.085 4.04 57.345 4.36 ;
      RECT 48.51 8.565 48.83 8.89 ;
      RECT 48.54 7.98 48.71 8.89 ;
      RECT 48.54 7.98 48.715 8.33 ;
      RECT 48.54 7.98 49.515 8.155 ;
      RECT 49.34 3.26 49.515 8.155 ;
      RECT 41.895 3.5 42.175 3.87 ;
      RECT 41.895 3.64 46.545 3.815 ;
      RECT 46.37 3.32 46.545 3.815 ;
      RECT 46.84 3.29 47.165 3.615 ;
      RECT 49.285 3.26 49.635 3.61 ;
      RECT 46.37 3.32 49.635 3.49 ;
      RECT 37.66 9.55 48.355 9.72 ;
      RECT 48.195 3.69 48.355 9.72 ;
      RECT 37.66 8.83 37.83 9.72 ;
      RECT 34.48 8.945 34.805 9.27 ;
      RECT 49.31 8.94 49.635 9.265 ;
      RECT 48.195 9.03 49.635 9.2 ;
      RECT 37.61 8.83 37.89 9.17 ;
      RECT 34.48 8.975 35.715 9.145 ;
      RECT 35.715 8.97 37.89 9.14 ;
      RECT 48.51 3.66 48.83 3.98 ;
      RECT 48.195 3.69 48.83 3.86 ;
      RECT 44.965 7.76 45.225 8.095 ;
      RECT 45.025 4.035 45.165 8.095 ;
      RECT 44.965 4.035 45.225 4.355 ;
      RECT 44.285 6.075 44.545 6.395 ;
      RECT 44.345 5.055 44.485 6.395 ;
      RECT 44.285 5.055 44.545 5.375 ;
      RECT 43.265 7.76 43.525 8.095 ;
      RECT 43.235 7.805 43.555 8.05 ;
      RECT 43.325 6.505 43.465 8.095 ;
      RECT 42.645 6.505 43.465 6.645 ;
      RECT 42.645 4.035 42.785 6.645 ;
      RECT 42.575 5.43 42.855 5.8 ;
      RECT 42.585 4.035 42.845 4.355 ;
      RECT 40.535 5.43 40.815 5.8 ;
      RECT 40.605 3.695 40.745 5.8 ;
      RECT 40.545 3.695 40.805 4.015 ;
      RECT 39.865 6.075 40.125 6.395 ;
      RECT 39.925 4.035 40.065 6.395 ;
      RECT 39.865 4.035 40.125 4.355 ;
      RECT 31.29 8.565 31.61 8.89 ;
      RECT 31.32 7.98 31.49 8.89 ;
      RECT 31.32 7.98 31.495 8.33 ;
      RECT 31.32 7.98 32.295 8.155 ;
      RECT 32.12 3.26 32.295 8.155 ;
      RECT 24.675 3.5 24.955 3.87 ;
      RECT 24.675 3.64 29.325 3.815 ;
      RECT 29.15 3.32 29.325 3.815 ;
      RECT 29.62 3.29 29.945 3.615 ;
      RECT 32.065 3.26 32.415 3.61 ;
      RECT 29.15 3.32 32.415 3.49 ;
      RECT 20.44 9.55 31.135 9.72 ;
      RECT 30.975 3.69 31.135 9.72 ;
      RECT 16.54 9.28 16.82 9.62 ;
      RECT 20.44 8.83 20.61 9.72 ;
      RECT 16.54 9.345 17.745 9.515 ;
      RECT 17.575 8.97 17.745 9.515 ;
      RECT 32.09 8.94 32.415 9.265 ;
      RECT 30.975 9.03 32.415 9.2 ;
      RECT 20.39 8.83 20.67 9.17 ;
      RECT 17.575 8.97 20.67 9.14 ;
      RECT 31.29 3.66 31.61 3.98 ;
      RECT 30.975 3.69 31.61 3.86 ;
      RECT 27.745 7.76 28.005 8.095 ;
      RECT 27.805 4.035 27.945 8.095 ;
      RECT 27.745 4.035 28.005 4.355 ;
      RECT 27.065 6.075 27.325 6.395 ;
      RECT 27.125 5.055 27.265 6.395 ;
      RECT 27.065 5.055 27.325 5.375 ;
      RECT 26.045 7.76 26.305 8.095 ;
      RECT 26.015 7.805 26.335 8.05 ;
      RECT 26.105 6.505 26.245 8.095 ;
      RECT 25.425 6.505 26.245 6.645 ;
      RECT 25.425 4.035 25.565 6.645 ;
      RECT 25.355 5.43 25.635 5.8 ;
      RECT 25.365 4.035 25.625 4.355 ;
      RECT 23.315 5.43 23.595 5.8 ;
      RECT 23.385 3.695 23.525 5.8 ;
      RECT 23.325 3.695 23.585 4.015 ;
      RECT 22.645 6.075 22.905 6.395 ;
      RECT 22.705 4.035 22.845 6.395 ;
      RECT 22.645 4.035 22.905 4.355 ;
      RECT 103.255 7.2 103.635 7.58 ;
      RECT 95.605 7.065 95.885 7.435 ;
      RECT 95.255 5.03 95.535 5.4 ;
      RECT 94.915 4.35 95.195 4.72 ;
      RECT 94.565 7.065 94.845 7.435 ;
      RECT 93.885 4.69 94.165 5.06 ;
      RECT 93.555 7.725 93.835 8.095 ;
      RECT 88.795 9.285 89.165 9.655 ;
      RECT 86.035 7.2 86.415 7.58 ;
      RECT 78.385 7.065 78.665 7.435 ;
      RECT 78.035 5.03 78.315 5.4 ;
      RECT 77.695 4.35 77.975 4.72 ;
      RECT 77.345 7.065 77.625 7.435 ;
      RECT 76.665 4.69 76.945 5.06 ;
      RECT 76.335 7.725 76.615 8.095 ;
      RECT 71.575 9.285 71.945 9.655 ;
      RECT 68.815 7.205 69.195 7.585 ;
      RECT 61.165 7.07 61.445 7.44 ;
      RECT 60.815 5.035 61.095 5.405 ;
      RECT 60.475 4.355 60.755 4.725 ;
      RECT 60.125 7.07 60.405 7.44 ;
      RECT 59.445 4.695 59.725 5.065 ;
      RECT 59.115 7.73 59.395 8.1 ;
      RECT 54.355 9.29 54.725 9.66 ;
      RECT 51.595 7.2 51.975 7.58 ;
      RECT 43.945 7.065 44.225 7.435 ;
      RECT 43.595 5.03 43.875 5.4 ;
      RECT 43.255 4.35 43.535 4.72 ;
      RECT 42.905 7.065 43.185 7.435 ;
      RECT 42.225 4.69 42.505 5.06 ;
      RECT 41.895 7.725 42.175 8.095 ;
      RECT 37.135 9.285 37.505 9.655 ;
      RECT 34.375 7.2 34.755 7.58 ;
      RECT 26.725 7.065 27.005 7.435 ;
      RECT 26.375 5.03 26.655 5.4 ;
      RECT 26.035 4.35 26.315 4.72 ;
      RECT 25.685 7.065 25.965 7.435 ;
      RECT 25.005 4.69 25.285 5.06 ;
      RECT 24.675 7.725 24.955 8.095 ;
      RECT 19.915 9.285 20.285 9.655 ;
    LAYER via1 ;
      RECT 103.415 9.67 103.565 9.82 ;
      RECT 103.37 7.315 103.52 7.465 ;
      RECT 101.06 9.025 101.21 9.175 ;
      RECT 101.045 3.36 101.195 3.51 ;
      RECT 100.255 3.745 100.405 3.895 ;
      RECT 100.255 8.655 100.405 8.805 ;
      RECT 98.59 3.375 98.74 3.525 ;
      RECT 96.68 4.12 96.83 4.27 ;
      RECT 96.68 7.845 96.83 7.995 ;
      RECT 96 5.14 96.15 5.29 ;
      RECT 96 6.16 96.15 6.31 ;
      RECT 95.66 7.165 95.81 7.315 ;
      RECT 95.32 5.14 95.47 5.29 ;
      RECT 94.98 4.46 95.13 4.61 ;
      RECT 94.98 7.845 95.13 7.995 ;
      RECT 94.63 7.165 94.78 7.315 ;
      RECT 94.3 4.12 94.45 4.27 ;
      RECT 93.96 4.8 94.11 4.95 ;
      RECT 93.62 3.61 93.77 3.76 ;
      RECT 93.62 7.83 93.77 7.98 ;
      RECT 92.26 3.78 92.41 3.93 ;
      RECT 91.58 4.12 91.73 4.27 ;
      RECT 91.58 6.16 91.73 6.31 ;
      RECT 89.335 8.925 89.485 9.075 ;
      RECT 88.905 9.395 89.055 9.545 ;
      RECT 86.23 9.03 86.38 9.18 ;
      RECT 86.15 7.315 86.3 7.465 ;
      RECT 83.84 9.025 83.99 9.175 ;
      RECT 83.825 3.36 83.975 3.51 ;
      RECT 83.035 3.745 83.185 3.895 ;
      RECT 83.035 8.655 83.185 8.805 ;
      RECT 81.37 3.375 81.52 3.525 ;
      RECT 79.46 4.12 79.61 4.27 ;
      RECT 79.46 7.845 79.61 7.995 ;
      RECT 78.78 5.14 78.93 5.29 ;
      RECT 78.78 6.16 78.93 6.31 ;
      RECT 78.44 7.165 78.59 7.315 ;
      RECT 78.1 5.14 78.25 5.29 ;
      RECT 77.76 4.46 77.91 4.61 ;
      RECT 77.76 7.845 77.91 7.995 ;
      RECT 77.41 7.165 77.56 7.315 ;
      RECT 77.08 4.12 77.23 4.27 ;
      RECT 76.74 4.8 76.89 4.95 ;
      RECT 76.4 3.61 76.55 3.76 ;
      RECT 76.4 7.83 76.55 7.98 ;
      RECT 75.04 3.78 75.19 3.93 ;
      RECT 74.36 4.12 74.51 4.27 ;
      RECT 74.36 6.16 74.51 6.31 ;
      RECT 72.115 8.925 72.265 9.075 ;
      RECT 71.685 9.395 71.835 9.545 ;
      RECT 69.01 9.035 69.16 9.185 ;
      RECT 68.93 7.32 69.08 7.47 ;
      RECT 66.62 9.03 66.77 9.18 ;
      RECT 66.605 3.365 66.755 3.515 ;
      RECT 65.815 3.75 65.965 3.9 ;
      RECT 65.815 8.66 65.965 8.81 ;
      RECT 64.15 3.38 64.3 3.53 ;
      RECT 62.24 4.125 62.39 4.275 ;
      RECT 62.24 7.85 62.39 8 ;
      RECT 61.56 5.145 61.71 5.295 ;
      RECT 61.56 6.165 61.71 6.315 ;
      RECT 61.22 7.17 61.37 7.32 ;
      RECT 60.88 5.145 61.03 5.295 ;
      RECT 60.54 4.465 60.69 4.615 ;
      RECT 60.54 7.85 60.69 8 ;
      RECT 60.19 7.17 60.34 7.32 ;
      RECT 59.86 4.125 60.01 4.275 ;
      RECT 59.52 4.805 59.67 4.955 ;
      RECT 59.18 3.615 59.33 3.765 ;
      RECT 59.18 7.835 59.33 7.985 ;
      RECT 57.82 3.785 57.97 3.935 ;
      RECT 57.14 4.125 57.29 4.275 ;
      RECT 57.14 6.165 57.29 6.315 ;
      RECT 54.895 8.93 55.045 9.08 ;
      RECT 54.465 9.4 54.615 9.55 ;
      RECT 51.79 9.03 51.94 9.18 ;
      RECT 51.71 7.315 51.86 7.465 ;
      RECT 49.4 9.025 49.55 9.175 ;
      RECT 49.385 3.36 49.535 3.51 ;
      RECT 48.595 3.745 48.745 3.895 ;
      RECT 48.595 8.655 48.745 8.805 ;
      RECT 46.93 3.375 47.08 3.525 ;
      RECT 45.02 4.12 45.17 4.27 ;
      RECT 45.02 7.845 45.17 7.995 ;
      RECT 44.34 5.14 44.49 5.29 ;
      RECT 44.34 6.16 44.49 6.31 ;
      RECT 44 7.165 44.15 7.315 ;
      RECT 43.66 5.14 43.81 5.29 ;
      RECT 43.32 4.46 43.47 4.61 ;
      RECT 43.32 7.845 43.47 7.995 ;
      RECT 42.97 7.165 43.12 7.315 ;
      RECT 42.64 4.12 42.79 4.27 ;
      RECT 42.3 4.8 42.45 4.95 ;
      RECT 41.96 3.61 42.11 3.76 ;
      RECT 41.96 7.83 42.11 7.98 ;
      RECT 40.6 3.78 40.75 3.93 ;
      RECT 39.92 4.12 40.07 4.27 ;
      RECT 39.92 6.16 40.07 6.31 ;
      RECT 37.675 8.925 37.825 9.075 ;
      RECT 37.245 9.395 37.395 9.545 ;
      RECT 34.57 9.03 34.72 9.18 ;
      RECT 34.49 7.315 34.64 7.465 ;
      RECT 32.18 9.025 32.33 9.175 ;
      RECT 32.165 3.36 32.315 3.51 ;
      RECT 31.375 3.745 31.525 3.895 ;
      RECT 31.375 8.655 31.525 8.805 ;
      RECT 29.71 3.375 29.86 3.525 ;
      RECT 27.8 4.12 27.95 4.27 ;
      RECT 27.8 7.845 27.95 7.995 ;
      RECT 27.12 5.14 27.27 5.29 ;
      RECT 27.12 6.16 27.27 6.31 ;
      RECT 26.78 7.165 26.93 7.315 ;
      RECT 26.44 5.14 26.59 5.29 ;
      RECT 26.1 4.46 26.25 4.61 ;
      RECT 26.1 7.845 26.25 7.995 ;
      RECT 25.75 7.165 25.9 7.315 ;
      RECT 25.42 4.12 25.57 4.27 ;
      RECT 25.08 4.8 25.23 4.95 ;
      RECT 24.74 3.61 24.89 3.76 ;
      RECT 24.74 7.83 24.89 7.98 ;
      RECT 23.38 3.78 23.53 3.93 ;
      RECT 22.7 4.12 22.85 4.27 ;
      RECT 22.7 6.16 22.85 6.31 ;
      RECT 20.455 8.925 20.605 9.075 ;
      RECT 20.025 9.395 20.175 9.545 ;
      RECT 16.605 9.375 16.755 9.525 ;
      RECT 16.23 8.635 16.38 8.785 ;
    LAYER met1 ;
      RECT 103.295 10.055 103.59 10.285 ;
      RECT 103.355 9.585 103.53 10.285 ;
      RECT 103.325 9.585 103.65 9.91 ;
      RECT 103.355 8.575 103.525 10.285 ;
      RECT 103.295 8.575 103.585 8.805 ;
      RECT 102.305 10.055 102.6 10.285 ;
      RECT 102.365 8.575 102.535 10.285 ;
      RECT 102.305 8.575 102.595 8.805 ;
      RECT 102.305 8.61 103.155 8.77 ;
      RECT 102.99 8.205 103.155 8.77 ;
      RECT 102.305 8.605 102.7 8.77 ;
      RECT 102.925 8.205 103.215 8.435 ;
      RECT 102.925 8.235 103.385 8.405 ;
      RECT 102.885 4.025 103.21 4.26 ;
      RECT 102.885 4.055 103.38 4.225 ;
      RECT 102.89 3.69 103.08 4.26 ;
      RECT 102.305 3.655 102.595 3.885 ;
      RECT 102.305 3.69 103.08 3.86 ;
      RECT 102.365 2.175 102.535 3.885 ;
      RECT 102.305 2.175 102.6 2.405 ;
      RECT 101.935 4.025 102.225 4.255 ;
      RECT 101.935 4.055 102.395 4.225 ;
      RECT 102 2.95 102.165 4.255 ;
      RECT 100.515 2.915 100.805 3.145 ;
      RECT 100.515 2.95 102.165 3.12 ;
      RECT 100.575 2.175 100.745 3.145 ;
      RECT 100.515 2.175 100.805 2.405 ;
      RECT 100.515 10.055 100.805 10.285 ;
      RECT 100.575 9.315 100.745 10.285 ;
      RECT 100.575 9.405 102.165 9.575 ;
      RECT 101.995 8.205 102.165 9.575 ;
      RECT 100.515 9.315 100.805 9.545 ;
      RECT 101.935 8.205 102.225 8.435 ;
      RECT 101.935 8.235 102.395 8.405 ;
      RECT 100.945 3.26 101.295 3.61 ;
      RECT 100.775 3.315 101.295 3.485 ;
      RECT 100.97 8.94 101.295 9.265 ;
      RECT 100.945 8.945 101.295 9.175 ;
      RECT 100.775 8.975 101.295 9.145 ;
      RECT 100.17 3.66 100.49 3.98 ;
      RECT 100.145 3.655 100.435 3.885 ;
      RECT 99.855 3.69 100.49 3.86 ;
      RECT 99.97 3.685 100.49 3.86 ;
      RECT 100.17 8.565 100.49 8.89 ;
      RECT 100.145 8.575 100.49 8.805 ;
      RECT 99.97 8.605 100.49 8.775 ;
      RECT 95.915 5.085 96.235 5.345 ;
      RECT 96.95 5.1 97.24 5.33 ;
      RECT 95.915 5.145 97.24 5.285 ;
      RECT 96.95 7.14 97.24 7.37 ;
      RECT 95.575 7.11 95.895 7.37 ;
      RECT 97.025 6.83 97.165 7.37 ;
      RECT 95.665 6.83 95.805 7.37 ;
      RECT 95.665 6.83 97.165 6.97 ;
      RECT 96.595 4.065 96.915 4.325 ;
      RECT 96.32 4.125 96.915 4.265 ;
      RECT 96.27 7.805 96.915 8.05 ;
      RECT 96.595 7.775 96.915 8.05 ;
      RECT 92.53 7.82 92.82 8.05 ;
      RECT 93.535 7.775 93.855 8.035 ;
      RECT 92.53 7.865 94.445 8.005 ;
      RECT 94.305 7.51 94.445 8.005 ;
      RECT 93.53 7.835 93.86 8.005 ;
      RECT 94.305 7.51 96.315 7.65 ;
      RECT 96.175 7.14 96.315 7.65 ;
      RECT 96.1 7.14 96.39 7.37 ;
      RECT 95.915 6.105 96.235 6.365 ;
      RECT 93.77 6.12 94.06 6.35 ;
      RECT 93.77 6.165 96.235 6.305 ;
      RECT 95.235 5.085 95.555 5.345 ;
      RECT 92.87 5.1 93.16 5.33 ;
      RECT 92.87 5.145 95.555 5.285 ;
      RECT 94.895 7.79 95.215 8.05 ;
      RECT 94.895 7.865 95.49 8.005 ;
      RECT 94.895 4.405 95.215 4.665 ;
      RECT 94.62 4.465 95.215 4.605 ;
      RECT 94.22 7.125 94.865 7.37 ;
      RECT 94.545 7.11 94.865 7.37 ;
      RECT 94.215 4.065 94.535 4.325 ;
      RECT 93.94 4.125 94.535 4.265 ;
      RECT 93.875 4.745 94.195 5.005 ;
      RECT 91 4.76 91.29 4.99 ;
      RECT 91 4.805 94.195 4.945 ;
      RECT 93.455 4.085 93.595 4.945 ;
      RECT 93.38 4.085 93.67 4.315 ;
      RECT 93.535 3.555 93.855 3.815 ;
      RECT 93.535 3.57 94.04 3.8 ;
      RECT 93.445 3.615 94.04 3.755 ;
      RECT 92.87 4.085 93.16 4.315 ;
      RECT 92.265 4.13 93.16 4.27 ;
      RECT 92.265 3.725 92.405 4.27 ;
      RECT 92.175 3.725 92.495 3.985 ;
      RECT 91.495 4.065 91.815 4.325 ;
      RECT 91.22 4.125 91.815 4.265 ;
      RECT 91.495 6.105 91.815 6.365 ;
      RECT 91.22 6.165 91.815 6.305 ;
      RECT 89.26 8.86 89.55 9.175 ;
      RECT 89.09 8.975 89.55 9.145 ;
      RECT 89.24 8.86 89.58 9.14 ;
      RECT 88.83 10.055 89.12 10.285 ;
      RECT 88.89 9.285 89.06 10.285 ;
      RECT 88.795 9.285 89.165 9.655 ;
      RECT 86.075 10.055 86.37 10.285 ;
      RECT 86.135 8.575 86.305 10.285 ;
      RECT 86.135 8.945 86.465 9.27 ;
      RECT 86.075 8.575 86.365 8.805 ;
      RECT 85.085 10.055 85.38 10.285 ;
      RECT 85.145 8.575 85.315 10.285 ;
      RECT 85.085 8.575 85.375 8.805 ;
      RECT 85.085 8.61 85.935 8.77 ;
      RECT 85.77 8.205 85.935 8.77 ;
      RECT 85.085 8.605 85.48 8.77 ;
      RECT 85.705 8.205 85.995 8.435 ;
      RECT 85.705 8.235 86.165 8.405 ;
      RECT 85.665 4.025 85.99 4.26 ;
      RECT 85.665 4.055 86.16 4.225 ;
      RECT 85.67 3.69 85.86 4.26 ;
      RECT 85.085 3.655 85.375 3.885 ;
      RECT 85.085 3.69 85.86 3.86 ;
      RECT 85.145 2.175 85.315 3.885 ;
      RECT 85.085 2.175 85.38 2.405 ;
      RECT 84.715 4.025 85.005 4.255 ;
      RECT 84.715 4.055 85.175 4.225 ;
      RECT 84.78 2.95 84.945 4.255 ;
      RECT 83.295 2.915 83.585 3.145 ;
      RECT 83.295 2.95 84.945 3.12 ;
      RECT 83.355 2.175 83.525 3.145 ;
      RECT 83.295 2.175 83.585 2.405 ;
      RECT 83.295 10.055 83.585 10.285 ;
      RECT 83.355 9.315 83.525 10.285 ;
      RECT 83.355 9.405 84.945 9.575 ;
      RECT 84.775 8.205 84.945 9.575 ;
      RECT 83.295 9.315 83.585 9.545 ;
      RECT 84.715 8.205 85.005 8.435 ;
      RECT 84.715 8.235 85.175 8.405 ;
      RECT 83.725 3.26 84.075 3.61 ;
      RECT 83.555 3.315 84.075 3.485 ;
      RECT 83.75 8.94 84.075 9.265 ;
      RECT 83.725 8.945 84.075 9.175 ;
      RECT 83.555 8.975 84.075 9.145 ;
      RECT 82.95 3.66 83.27 3.98 ;
      RECT 82.925 3.655 83.215 3.885 ;
      RECT 82.635 3.69 83.27 3.86 ;
      RECT 82.75 3.685 83.27 3.86 ;
      RECT 82.95 8.565 83.27 8.89 ;
      RECT 82.925 8.575 83.27 8.805 ;
      RECT 82.75 8.605 83.27 8.775 ;
      RECT 78.695 5.085 79.015 5.345 ;
      RECT 79.73 5.1 80.02 5.33 ;
      RECT 78.695 5.145 80.02 5.285 ;
      RECT 79.73 7.14 80.02 7.37 ;
      RECT 78.355 7.11 78.675 7.37 ;
      RECT 79.805 6.83 79.945 7.37 ;
      RECT 78.445 6.83 78.585 7.37 ;
      RECT 78.445 6.83 79.945 6.97 ;
      RECT 79.375 4.065 79.695 4.325 ;
      RECT 79.1 4.125 79.695 4.265 ;
      RECT 79.05 7.805 79.695 8.05 ;
      RECT 79.375 7.775 79.695 8.05 ;
      RECT 75.31 7.82 75.6 8.05 ;
      RECT 76.315 7.775 76.635 8.035 ;
      RECT 75.31 7.865 77.225 8.005 ;
      RECT 77.085 7.51 77.225 8.005 ;
      RECT 76.31 7.835 76.64 8.005 ;
      RECT 77.085 7.51 79.095 7.65 ;
      RECT 78.955 7.14 79.095 7.65 ;
      RECT 78.88 7.14 79.17 7.37 ;
      RECT 78.695 6.105 79.015 6.365 ;
      RECT 76.55 6.12 76.84 6.35 ;
      RECT 76.55 6.165 79.015 6.305 ;
      RECT 78.015 5.085 78.335 5.345 ;
      RECT 75.65 5.1 75.94 5.33 ;
      RECT 75.65 5.145 78.335 5.285 ;
      RECT 77.675 7.79 77.995 8.05 ;
      RECT 77.675 7.865 78.27 8.005 ;
      RECT 77.675 4.405 77.995 4.665 ;
      RECT 77.4 4.465 77.995 4.605 ;
      RECT 77 7.125 77.645 7.37 ;
      RECT 77.325 7.11 77.645 7.37 ;
      RECT 76.995 4.065 77.315 4.325 ;
      RECT 76.72 4.125 77.315 4.265 ;
      RECT 76.655 4.745 76.975 5.005 ;
      RECT 73.78 4.76 74.07 4.99 ;
      RECT 73.78 4.805 76.975 4.945 ;
      RECT 76.235 4.085 76.375 4.945 ;
      RECT 76.16 4.085 76.45 4.315 ;
      RECT 76.315 3.555 76.635 3.815 ;
      RECT 76.315 3.57 76.82 3.8 ;
      RECT 76.225 3.615 76.82 3.755 ;
      RECT 75.65 4.085 75.94 4.315 ;
      RECT 75.045 4.13 75.94 4.27 ;
      RECT 75.045 3.725 75.185 4.27 ;
      RECT 74.955 3.725 75.275 3.985 ;
      RECT 74.275 4.065 74.595 4.325 ;
      RECT 74 4.125 74.595 4.265 ;
      RECT 74.275 6.105 74.595 6.365 ;
      RECT 74 6.165 74.595 6.305 ;
      RECT 72.04 8.86 72.33 9.175 ;
      RECT 71.87 8.975 72.33 9.145 ;
      RECT 72.02 8.86 72.36 9.14 ;
      RECT 71.61 10.055 71.9 10.285 ;
      RECT 71.67 9.285 71.84 10.285 ;
      RECT 71.575 9.285 71.945 9.655 ;
      RECT 68.855 10.06 69.15 10.29 ;
      RECT 68.915 8.58 69.085 10.29 ;
      RECT 68.915 8.95 69.245 9.275 ;
      RECT 68.855 8.58 69.145 8.81 ;
      RECT 67.865 10.06 68.16 10.29 ;
      RECT 67.925 8.58 68.095 10.29 ;
      RECT 67.865 8.58 68.155 8.81 ;
      RECT 67.865 8.615 68.715 8.775 ;
      RECT 68.55 8.21 68.715 8.775 ;
      RECT 67.865 8.61 68.26 8.775 ;
      RECT 68.485 8.21 68.775 8.44 ;
      RECT 68.485 8.24 68.945 8.41 ;
      RECT 68.445 4.03 68.77 4.265 ;
      RECT 68.445 4.06 68.94 4.23 ;
      RECT 68.45 3.695 68.64 4.265 ;
      RECT 67.865 3.66 68.155 3.89 ;
      RECT 67.865 3.695 68.64 3.865 ;
      RECT 67.925 2.18 68.095 3.89 ;
      RECT 67.865 2.18 68.16 2.41 ;
      RECT 67.495 4.03 67.785 4.26 ;
      RECT 67.495 4.06 67.955 4.23 ;
      RECT 67.56 2.955 67.725 4.26 ;
      RECT 66.075 2.92 66.365 3.15 ;
      RECT 66.075 2.955 67.725 3.125 ;
      RECT 66.135 2.18 66.305 3.15 ;
      RECT 66.075 2.18 66.365 2.41 ;
      RECT 66.075 10.06 66.365 10.29 ;
      RECT 66.135 9.32 66.305 10.29 ;
      RECT 66.135 9.41 67.725 9.58 ;
      RECT 67.555 8.21 67.725 9.58 ;
      RECT 66.075 9.32 66.365 9.55 ;
      RECT 67.495 8.21 67.785 8.44 ;
      RECT 67.495 8.24 67.955 8.41 ;
      RECT 66.505 3.265 66.855 3.615 ;
      RECT 66.335 3.32 66.855 3.49 ;
      RECT 66.53 8.945 66.855 9.27 ;
      RECT 66.505 8.95 66.855 9.18 ;
      RECT 66.335 8.98 66.855 9.15 ;
      RECT 65.73 3.665 66.05 3.985 ;
      RECT 65.705 3.66 65.995 3.89 ;
      RECT 65.415 3.695 66.05 3.865 ;
      RECT 65.53 3.69 66.05 3.865 ;
      RECT 65.73 8.57 66.05 8.895 ;
      RECT 65.705 8.58 66.05 8.81 ;
      RECT 65.53 8.61 66.05 8.78 ;
      RECT 61.475 5.09 61.795 5.35 ;
      RECT 62.51 5.105 62.8 5.335 ;
      RECT 61.475 5.15 62.8 5.29 ;
      RECT 62.51 7.145 62.8 7.375 ;
      RECT 61.135 7.115 61.455 7.375 ;
      RECT 62.585 6.835 62.725 7.375 ;
      RECT 61.225 6.835 61.365 7.375 ;
      RECT 61.225 6.835 62.725 6.975 ;
      RECT 62.155 4.07 62.475 4.33 ;
      RECT 61.88 4.13 62.475 4.27 ;
      RECT 61.83 7.81 62.475 8.055 ;
      RECT 62.155 7.78 62.475 8.055 ;
      RECT 58.09 7.825 58.38 8.055 ;
      RECT 59.095 7.78 59.415 8.04 ;
      RECT 58.09 7.87 60.005 8.01 ;
      RECT 59.865 7.515 60.005 8.01 ;
      RECT 59.09 7.84 59.42 8.01 ;
      RECT 59.865 7.515 61.875 7.655 ;
      RECT 61.735 7.145 61.875 7.655 ;
      RECT 61.66 7.145 61.95 7.375 ;
      RECT 61.475 6.11 61.795 6.37 ;
      RECT 59.33 6.125 59.62 6.355 ;
      RECT 59.33 6.17 61.795 6.31 ;
      RECT 60.795 5.09 61.115 5.35 ;
      RECT 58.43 5.105 58.72 5.335 ;
      RECT 58.43 5.15 61.115 5.29 ;
      RECT 60.455 7.795 60.775 8.055 ;
      RECT 60.455 7.87 61.05 8.01 ;
      RECT 60.455 4.41 60.775 4.67 ;
      RECT 60.18 4.47 60.775 4.61 ;
      RECT 59.78 7.13 60.425 7.375 ;
      RECT 60.105 7.115 60.425 7.375 ;
      RECT 59.775 4.07 60.095 4.33 ;
      RECT 59.5 4.13 60.095 4.27 ;
      RECT 59.435 4.75 59.755 5.01 ;
      RECT 56.56 4.765 56.85 4.995 ;
      RECT 56.56 4.81 59.755 4.95 ;
      RECT 59.015 4.09 59.155 4.95 ;
      RECT 58.94 4.09 59.23 4.32 ;
      RECT 59.095 3.56 59.415 3.82 ;
      RECT 59.095 3.575 59.6 3.805 ;
      RECT 59.005 3.62 59.6 3.76 ;
      RECT 58.43 4.09 58.72 4.32 ;
      RECT 57.825 4.135 58.72 4.275 ;
      RECT 57.825 3.73 57.965 4.275 ;
      RECT 57.735 3.73 58.055 3.99 ;
      RECT 57.055 4.07 57.375 4.33 ;
      RECT 56.78 4.13 57.375 4.27 ;
      RECT 57.055 6.11 57.375 6.37 ;
      RECT 56.78 6.17 57.375 6.31 ;
      RECT 54.82 8.865 55.11 9.18 ;
      RECT 54.65 8.98 55.11 9.15 ;
      RECT 54.8 8.865 55.14 9.145 ;
      RECT 54.39 10.06 54.68 10.29 ;
      RECT 54.45 9.29 54.62 10.29 ;
      RECT 54.355 9.29 54.725 9.66 ;
      RECT 51.635 10.055 51.93 10.285 ;
      RECT 51.695 8.575 51.865 10.285 ;
      RECT 51.695 8.945 52.025 9.27 ;
      RECT 51.635 8.575 51.925 8.805 ;
      RECT 50.645 10.055 50.94 10.285 ;
      RECT 50.705 8.575 50.875 10.285 ;
      RECT 50.645 8.575 50.935 8.805 ;
      RECT 50.645 8.61 51.495 8.77 ;
      RECT 51.33 8.205 51.495 8.77 ;
      RECT 50.645 8.605 51.04 8.77 ;
      RECT 51.265 8.205 51.555 8.435 ;
      RECT 51.265 8.235 51.725 8.405 ;
      RECT 51.225 4.025 51.55 4.26 ;
      RECT 51.225 4.055 51.72 4.225 ;
      RECT 51.23 3.69 51.42 4.26 ;
      RECT 50.645 3.655 50.935 3.885 ;
      RECT 50.645 3.69 51.42 3.86 ;
      RECT 50.705 2.175 50.875 3.885 ;
      RECT 50.645 2.175 50.94 2.405 ;
      RECT 50.275 4.025 50.565 4.255 ;
      RECT 50.275 4.055 50.735 4.225 ;
      RECT 50.34 2.95 50.505 4.255 ;
      RECT 48.855 2.915 49.145 3.145 ;
      RECT 48.855 2.95 50.505 3.12 ;
      RECT 48.915 2.175 49.085 3.145 ;
      RECT 48.855 2.175 49.145 2.405 ;
      RECT 48.855 10.055 49.145 10.285 ;
      RECT 48.915 9.315 49.085 10.285 ;
      RECT 48.915 9.405 50.505 9.575 ;
      RECT 50.335 8.205 50.505 9.575 ;
      RECT 48.855 9.315 49.145 9.545 ;
      RECT 50.275 8.205 50.565 8.435 ;
      RECT 50.275 8.235 50.735 8.405 ;
      RECT 49.285 3.26 49.635 3.61 ;
      RECT 49.115 3.315 49.635 3.485 ;
      RECT 49.31 8.94 49.635 9.265 ;
      RECT 49.285 8.945 49.635 9.175 ;
      RECT 49.115 8.975 49.635 9.145 ;
      RECT 48.51 3.66 48.83 3.98 ;
      RECT 48.485 3.655 48.775 3.885 ;
      RECT 48.195 3.69 48.83 3.86 ;
      RECT 48.31 3.685 48.83 3.86 ;
      RECT 48.51 8.565 48.83 8.89 ;
      RECT 48.485 8.575 48.83 8.805 ;
      RECT 48.31 8.605 48.83 8.775 ;
      RECT 44.255 5.085 44.575 5.345 ;
      RECT 45.29 5.1 45.58 5.33 ;
      RECT 44.255 5.145 45.58 5.285 ;
      RECT 45.29 7.14 45.58 7.37 ;
      RECT 43.915 7.11 44.235 7.37 ;
      RECT 45.365 6.83 45.505 7.37 ;
      RECT 44.005 6.83 44.145 7.37 ;
      RECT 44.005 6.83 45.505 6.97 ;
      RECT 44.935 4.065 45.255 4.325 ;
      RECT 44.66 4.125 45.255 4.265 ;
      RECT 44.61 7.805 45.255 8.05 ;
      RECT 44.935 7.775 45.255 8.05 ;
      RECT 40.87 7.82 41.16 8.05 ;
      RECT 41.875 7.775 42.195 8.035 ;
      RECT 40.87 7.865 42.785 8.005 ;
      RECT 42.645 7.51 42.785 8.005 ;
      RECT 41.87 7.835 42.2 8.005 ;
      RECT 42.645 7.51 44.655 7.65 ;
      RECT 44.515 7.14 44.655 7.65 ;
      RECT 44.44 7.14 44.73 7.37 ;
      RECT 44.255 6.105 44.575 6.365 ;
      RECT 42.11 6.12 42.4 6.35 ;
      RECT 42.11 6.165 44.575 6.305 ;
      RECT 43.575 5.085 43.895 5.345 ;
      RECT 41.21 5.1 41.5 5.33 ;
      RECT 41.21 5.145 43.895 5.285 ;
      RECT 43.235 7.79 43.555 8.05 ;
      RECT 43.235 7.865 43.83 8.005 ;
      RECT 43.235 4.405 43.555 4.665 ;
      RECT 42.96 4.465 43.555 4.605 ;
      RECT 42.56 7.125 43.205 7.37 ;
      RECT 42.885 7.11 43.205 7.37 ;
      RECT 42.555 4.065 42.875 4.325 ;
      RECT 42.28 4.125 42.875 4.265 ;
      RECT 42.215 4.745 42.535 5.005 ;
      RECT 39.34 4.76 39.63 4.99 ;
      RECT 39.34 4.805 42.535 4.945 ;
      RECT 41.795 4.085 41.935 4.945 ;
      RECT 41.72 4.085 42.01 4.315 ;
      RECT 41.875 3.555 42.195 3.815 ;
      RECT 41.875 3.57 42.38 3.8 ;
      RECT 41.785 3.615 42.38 3.755 ;
      RECT 41.21 4.085 41.5 4.315 ;
      RECT 40.605 4.13 41.5 4.27 ;
      RECT 40.605 3.725 40.745 4.27 ;
      RECT 40.515 3.725 40.835 3.985 ;
      RECT 39.835 4.065 40.155 4.325 ;
      RECT 39.56 4.125 40.155 4.265 ;
      RECT 39.835 6.105 40.155 6.365 ;
      RECT 39.56 6.165 40.155 6.305 ;
      RECT 37.6 8.86 37.89 9.175 ;
      RECT 37.43 8.975 37.89 9.145 ;
      RECT 37.58 8.86 37.92 9.14 ;
      RECT 37.17 10.055 37.46 10.285 ;
      RECT 37.23 9.285 37.4 10.285 ;
      RECT 37.135 9.285 37.505 9.655 ;
      RECT 34.415 10.055 34.71 10.285 ;
      RECT 34.475 8.575 34.645 10.285 ;
      RECT 34.475 8.945 34.805 9.27 ;
      RECT 34.415 8.575 34.705 8.805 ;
      RECT 33.425 10.055 33.72 10.285 ;
      RECT 33.485 8.575 33.655 10.285 ;
      RECT 33.425 8.575 33.715 8.805 ;
      RECT 33.425 8.61 34.275 8.77 ;
      RECT 34.11 8.205 34.275 8.77 ;
      RECT 33.425 8.605 33.82 8.77 ;
      RECT 34.045 8.205 34.335 8.435 ;
      RECT 34.045 8.235 34.505 8.405 ;
      RECT 34.005 4.025 34.33 4.26 ;
      RECT 34.005 4.055 34.5 4.225 ;
      RECT 34.01 3.69 34.2 4.26 ;
      RECT 33.425 3.655 33.715 3.885 ;
      RECT 33.425 3.69 34.2 3.86 ;
      RECT 33.485 2.175 33.655 3.885 ;
      RECT 33.425 2.175 33.72 2.405 ;
      RECT 33.055 4.025 33.345 4.255 ;
      RECT 33.055 4.055 33.515 4.225 ;
      RECT 33.12 2.95 33.285 4.255 ;
      RECT 31.635 2.915 31.925 3.145 ;
      RECT 31.635 2.95 33.285 3.12 ;
      RECT 31.695 2.175 31.865 3.145 ;
      RECT 31.635 2.175 31.925 2.405 ;
      RECT 31.635 10.055 31.925 10.285 ;
      RECT 31.695 9.315 31.865 10.285 ;
      RECT 31.695 9.405 33.285 9.575 ;
      RECT 33.115 8.205 33.285 9.575 ;
      RECT 31.635 9.315 31.925 9.545 ;
      RECT 33.055 8.205 33.345 8.435 ;
      RECT 33.055 8.235 33.515 8.405 ;
      RECT 32.065 3.26 32.415 3.61 ;
      RECT 31.895 3.315 32.415 3.485 ;
      RECT 32.09 8.94 32.415 9.265 ;
      RECT 32.065 8.945 32.415 9.175 ;
      RECT 31.895 8.975 32.415 9.145 ;
      RECT 31.29 3.66 31.61 3.98 ;
      RECT 31.265 3.655 31.555 3.885 ;
      RECT 30.975 3.69 31.61 3.86 ;
      RECT 31.09 3.685 31.61 3.86 ;
      RECT 31.29 8.565 31.61 8.89 ;
      RECT 31.265 8.575 31.61 8.805 ;
      RECT 31.09 8.605 31.61 8.775 ;
      RECT 27.035 5.085 27.355 5.345 ;
      RECT 28.07 5.1 28.36 5.33 ;
      RECT 27.035 5.145 28.36 5.285 ;
      RECT 28.07 7.14 28.36 7.37 ;
      RECT 26.695 7.11 27.015 7.37 ;
      RECT 28.145 6.83 28.285 7.37 ;
      RECT 26.785 6.83 26.925 7.37 ;
      RECT 26.785 6.83 28.285 6.97 ;
      RECT 27.715 4.065 28.035 4.325 ;
      RECT 27.44 4.125 28.035 4.265 ;
      RECT 27.39 7.805 28.035 8.05 ;
      RECT 27.715 7.775 28.035 8.05 ;
      RECT 23.65 7.82 23.94 8.05 ;
      RECT 24.655 7.775 24.975 8.035 ;
      RECT 23.65 7.865 25.565 8.005 ;
      RECT 25.425 7.51 25.565 8.005 ;
      RECT 24.65 7.835 24.98 8.005 ;
      RECT 25.425 7.51 27.435 7.65 ;
      RECT 27.295 7.14 27.435 7.65 ;
      RECT 27.22 7.14 27.51 7.37 ;
      RECT 27.035 6.105 27.355 6.365 ;
      RECT 24.89 6.12 25.18 6.35 ;
      RECT 24.89 6.165 27.355 6.305 ;
      RECT 26.355 5.085 26.675 5.345 ;
      RECT 23.99 5.1 24.28 5.33 ;
      RECT 23.99 5.145 26.675 5.285 ;
      RECT 26.015 7.79 26.335 8.05 ;
      RECT 26.015 7.865 26.61 8.005 ;
      RECT 26.015 4.405 26.335 4.665 ;
      RECT 25.74 4.465 26.335 4.605 ;
      RECT 25.34 7.125 25.985 7.37 ;
      RECT 25.665 7.11 25.985 7.37 ;
      RECT 25.335 4.065 25.655 4.325 ;
      RECT 25.06 4.125 25.655 4.265 ;
      RECT 24.995 4.745 25.315 5.005 ;
      RECT 22.12 4.76 22.41 4.99 ;
      RECT 22.12 4.805 25.315 4.945 ;
      RECT 24.575 4.085 24.715 4.945 ;
      RECT 24.5 4.085 24.79 4.315 ;
      RECT 24.655 3.555 24.975 3.815 ;
      RECT 24.655 3.57 25.16 3.8 ;
      RECT 24.565 3.615 25.16 3.755 ;
      RECT 23.99 4.085 24.28 4.315 ;
      RECT 23.385 4.13 24.28 4.27 ;
      RECT 23.385 3.725 23.525 4.27 ;
      RECT 23.295 3.725 23.615 3.985 ;
      RECT 22.615 4.065 22.935 4.325 ;
      RECT 22.34 4.125 22.935 4.265 ;
      RECT 22.615 6.105 22.935 6.365 ;
      RECT 22.34 6.165 22.935 6.305 ;
      RECT 20.38 8.86 20.67 9.175 ;
      RECT 20.21 8.975 20.67 9.145 ;
      RECT 20.36 8.86 20.7 9.14 ;
      RECT 19.95 10.055 20.24 10.285 ;
      RECT 20.01 9.285 20.18 10.285 ;
      RECT 19.915 9.285 20.285 9.655 ;
      RECT 16.54 10.055 16.83 10.285 ;
      RECT 16.6 9.31 16.77 10.285 ;
      RECT 16.51 9.31 16.85 9.59 ;
      RECT 16.135 8.57 16.475 8.85 ;
      RECT 15.995 8.605 16.475 8.775 ;
      RECT 103.27 7.245 103.62 7.535 ;
      RECT 98.5 3.29 98.825 3.615 ;
      RECT 86.05 7.245 86.4 7.535 ;
      RECT 81.28 3.29 81.605 3.615 ;
      RECT 68.83 7.25 69.18 7.54 ;
      RECT 64.06 3.295 64.385 3.62 ;
      RECT 51.61 7.245 51.96 7.535 ;
      RECT 46.84 3.29 47.165 3.615 ;
      RECT 34.39 7.245 34.74 7.535 ;
      RECT 29.62 3.29 29.945 3.615 ;
    LAYER mcon ;
      RECT 103.36 7.305 103.53 7.475 ;
      RECT 103.355 8.605 103.525 8.775 ;
      RECT 103.355 10.085 103.525 10.255 ;
      RECT 102.985 8.235 103.155 8.405 ;
      RECT 102.98 4.055 103.15 4.225 ;
      RECT 102.365 2.205 102.535 2.375 ;
      RECT 102.365 3.685 102.535 3.855 ;
      RECT 102.365 8.605 102.535 8.775 ;
      RECT 102.365 10.085 102.535 10.255 ;
      RECT 101.995 4.055 102.165 4.225 ;
      RECT 101.995 8.235 102.165 8.405 ;
      RECT 101.005 3.315 101.175 3.485 ;
      RECT 101.005 8.975 101.175 9.145 ;
      RECT 100.575 2.205 100.745 2.375 ;
      RECT 100.575 2.945 100.745 3.115 ;
      RECT 100.575 9.345 100.745 9.515 ;
      RECT 100.575 10.085 100.745 10.255 ;
      RECT 100.205 3.685 100.375 3.855 ;
      RECT 100.205 8.605 100.375 8.775 ;
      RECT 97.01 5.13 97.18 5.3 ;
      RECT 97.01 7.17 97.18 7.34 ;
      RECT 96.67 4.11 96.84 4.28 ;
      RECT 96.33 7.85 96.5 8.02 ;
      RECT 96.16 7.17 96.33 7.34 ;
      RECT 95.65 7.17 95.82 7.34 ;
      RECT 94.97 4.45 95.14 4.62 ;
      RECT 94.97 7.85 95.14 8.02 ;
      RECT 94.29 4.11 94.46 4.28 ;
      RECT 94.28 7.17 94.45 7.34 ;
      RECT 93.83 6.15 94 6.32 ;
      RECT 93.81 3.6 93.98 3.77 ;
      RECT 93.44 4.115 93.61 4.285 ;
      RECT 92.93 4.115 93.1 4.285 ;
      RECT 92.93 5.13 93.1 5.3 ;
      RECT 92.59 7.85 92.76 8.02 ;
      RECT 91.57 4.11 91.74 4.28 ;
      RECT 91.57 6.15 91.74 6.32 ;
      RECT 91.06 4.79 91.23 4.96 ;
      RECT 89.32 8.975 89.49 9.145 ;
      RECT 88.89 9.345 89.06 9.515 ;
      RECT 88.89 10.085 89.06 10.255 ;
      RECT 86.14 7.305 86.31 7.475 ;
      RECT 86.135 8.605 86.305 8.775 ;
      RECT 86.135 10.085 86.305 10.255 ;
      RECT 85.765 8.235 85.935 8.405 ;
      RECT 85.76 4.055 85.93 4.225 ;
      RECT 85.145 2.205 85.315 2.375 ;
      RECT 85.145 3.685 85.315 3.855 ;
      RECT 85.145 8.605 85.315 8.775 ;
      RECT 85.145 10.085 85.315 10.255 ;
      RECT 84.775 4.055 84.945 4.225 ;
      RECT 84.775 8.235 84.945 8.405 ;
      RECT 83.785 3.315 83.955 3.485 ;
      RECT 83.785 8.975 83.955 9.145 ;
      RECT 83.355 2.205 83.525 2.375 ;
      RECT 83.355 2.945 83.525 3.115 ;
      RECT 83.355 9.345 83.525 9.515 ;
      RECT 83.355 10.085 83.525 10.255 ;
      RECT 82.985 3.685 83.155 3.855 ;
      RECT 82.985 8.605 83.155 8.775 ;
      RECT 79.79 5.13 79.96 5.3 ;
      RECT 79.79 7.17 79.96 7.34 ;
      RECT 79.45 4.11 79.62 4.28 ;
      RECT 79.11 7.85 79.28 8.02 ;
      RECT 78.94 7.17 79.11 7.34 ;
      RECT 78.43 7.17 78.6 7.34 ;
      RECT 77.75 4.45 77.92 4.62 ;
      RECT 77.75 7.85 77.92 8.02 ;
      RECT 77.07 4.11 77.24 4.28 ;
      RECT 77.06 7.17 77.23 7.34 ;
      RECT 76.61 6.15 76.78 6.32 ;
      RECT 76.59 3.6 76.76 3.77 ;
      RECT 76.22 4.115 76.39 4.285 ;
      RECT 75.71 4.115 75.88 4.285 ;
      RECT 75.71 5.13 75.88 5.3 ;
      RECT 75.37 7.85 75.54 8.02 ;
      RECT 74.35 4.11 74.52 4.28 ;
      RECT 74.35 6.15 74.52 6.32 ;
      RECT 73.84 4.79 74.01 4.96 ;
      RECT 72.1 8.975 72.27 9.145 ;
      RECT 71.67 9.345 71.84 9.515 ;
      RECT 71.67 10.085 71.84 10.255 ;
      RECT 68.92 7.31 69.09 7.48 ;
      RECT 68.915 8.61 69.085 8.78 ;
      RECT 68.915 10.09 69.085 10.26 ;
      RECT 68.545 8.24 68.715 8.41 ;
      RECT 68.54 4.06 68.71 4.23 ;
      RECT 67.925 2.21 68.095 2.38 ;
      RECT 67.925 3.69 68.095 3.86 ;
      RECT 67.925 8.61 68.095 8.78 ;
      RECT 67.925 10.09 68.095 10.26 ;
      RECT 67.555 4.06 67.725 4.23 ;
      RECT 67.555 8.24 67.725 8.41 ;
      RECT 66.565 3.32 66.735 3.49 ;
      RECT 66.565 8.98 66.735 9.15 ;
      RECT 66.135 2.21 66.305 2.38 ;
      RECT 66.135 2.95 66.305 3.12 ;
      RECT 66.135 9.35 66.305 9.52 ;
      RECT 66.135 10.09 66.305 10.26 ;
      RECT 65.765 3.69 65.935 3.86 ;
      RECT 65.765 8.61 65.935 8.78 ;
      RECT 62.57 5.135 62.74 5.305 ;
      RECT 62.57 7.175 62.74 7.345 ;
      RECT 62.23 4.115 62.4 4.285 ;
      RECT 61.89 7.855 62.06 8.025 ;
      RECT 61.72 7.175 61.89 7.345 ;
      RECT 61.21 7.175 61.38 7.345 ;
      RECT 60.53 4.455 60.7 4.625 ;
      RECT 60.53 7.855 60.7 8.025 ;
      RECT 59.85 4.115 60.02 4.285 ;
      RECT 59.84 7.175 60.01 7.345 ;
      RECT 59.39 6.155 59.56 6.325 ;
      RECT 59.37 3.605 59.54 3.775 ;
      RECT 59 4.12 59.17 4.29 ;
      RECT 58.49 4.12 58.66 4.29 ;
      RECT 58.49 5.135 58.66 5.305 ;
      RECT 58.15 7.855 58.32 8.025 ;
      RECT 57.13 4.115 57.3 4.285 ;
      RECT 57.13 6.155 57.3 6.325 ;
      RECT 56.62 4.795 56.79 4.965 ;
      RECT 54.88 8.98 55.05 9.15 ;
      RECT 54.45 9.35 54.62 9.52 ;
      RECT 54.45 10.09 54.62 10.26 ;
      RECT 51.7 7.305 51.87 7.475 ;
      RECT 51.695 8.605 51.865 8.775 ;
      RECT 51.695 10.085 51.865 10.255 ;
      RECT 51.325 8.235 51.495 8.405 ;
      RECT 51.32 4.055 51.49 4.225 ;
      RECT 50.705 2.205 50.875 2.375 ;
      RECT 50.705 3.685 50.875 3.855 ;
      RECT 50.705 8.605 50.875 8.775 ;
      RECT 50.705 10.085 50.875 10.255 ;
      RECT 50.335 4.055 50.505 4.225 ;
      RECT 50.335 8.235 50.505 8.405 ;
      RECT 49.345 3.315 49.515 3.485 ;
      RECT 49.345 8.975 49.515 9.145 ;
      RECT 48.915 2.205 49.085 2.375 ;
      RECT 48.915 2.945 49.085 3.115 ;
      RECT 48.915 9.345 49.085 9.515 ;
      RECT 48.915 10.085 49.085 10.255 ;
      RECT 48.545 3.685 48.715 3.855 ;
      RECT 48.545 8.605 48.715 8.775 ;
      RECT 45.35 5.13 45.52 5.3 ;
      RECT 45.35 7.17 45.52 7.34 ;
      RECT 45.01 4.11 45.18 4.28 ;
      RECT 44.67 7.85 44.84 8.02 ;
      RECT 44.5 7.17 44.67 7.34 ;
      RECT 43.99 7.17 44.16 7.34 ;
      RECT 43.31 4.45 43.48 4.62 ;
      RECT 43.31 7.85 43.48 8.02 ;
      RECT 42.63 4.11 42.8 4.28 ;
      RECT 42.62 7.17 42.79 7.34 ;
      RECT 42.17 6.15 42.34 6.32 ;
      RECT 42.15 3.6 42.32 3.77 ;
      RECT 41.78 4.115 41.95 4.285 ;
      RECT 41.27 4.115 41.44 4.285 ;
      RECT 41.27 5.13 41.44 5.3 ;
      RECT 40.93 7.85 41.1 8.02 ;
      RECT 39.91 4.11 40.08 4.28 ;
      RECT 39.91 6.15 40.08 6.32 ;
      RECT 39.4 4.79 39.57 4.96 ;
      RECT 37.66 8.975 37.83 9.145 ;
      RECT 37.23 9.345 37.4 9.515 ;
      RECT 37.23 10.085 37.4 10.255 ;
      RECT 34.48 7.305 34.65 7.475 ;
      RECT 34.475 8.605 34.645 8.775 ;
      RECT 34.475 10.085 34.645 10.255 ;
      RECT 34.105 8.235 34.275 8.405 ;
      RECT 34.1 4.055 34.27 4.225 ;
      RECT 33.485 2.205 33.655 2.375 ;
      RECT 33.485 3.685 33.655 3.855 ;
      RECT 33.485 8.605 33.655 8.775 ;
      RECT 33.485 10.085 33.655 10.255 ;
      RECT 33.115 4.055 33.285 4.225 ;
      RECT 33.115 8.235 33.285 8.405 ;
      RECT 32.125 3.315 32.295 3.485 ;
      RECT 32.125 8.975 32.295 9.145 ;
      RECT 31.695 2.205 31.865 2.375 ;
      RECT 31.695 2.945 31.865 3.115 ;
      RECT 31.695 9.345 31.865 9.515 ;
      RECT 31.695 10.085 31.865 10.255 ;
      RECT 31.325 3.685 31.495 3.855 ;
      RECT 31.325 8.605 31.495 8.775 ;
      RECT 28.13 5.13 28.3 5.3 ;
      RECT 28.13 7.17 28.3 7.34 ;
      RECT 27.79 4.11 27.96 4.28 ;
      RECT 27.45 7.85 27.62 8.02 ;
      RECT 27.28 7.17 27.45 7.34 ;
      RECT 26.77 7.17 26.94 7.34 ;
      RECT 26.09 4.45 26.26 4.62 ;
      RECT 26.09 7.85 26.26 8.02 ;
      RECT 25.41 4.11 25.58 4.28 ;
      RECT 25.4 7.17 25.57 7.34 ;
      RECT 24.95 6.15 25.12 6.32 ;
      RECT 24.93 3.6 25.1 3.77 ;
      RECT 24.56 4.115 24.73 4.285 ;
      RECT 24.05 4.115 24.22 4.285 ;
      RECT 24.05 5.13 24.22 5.3 ;
      RECT 23.71 7.85 23.88 8.02 ;
      RECT 22.69 4.11 22.86 4.28 ;
      RECT 22.69 6.15 22.86 6.32 ;
      RECT 22.18 4.79 22.35 4.96 ;
      RECT 20.44 8.975 20.61 9.145 ;
      RECT 20.01 9.345 20.18 9.515 ;
      RECT 20.01 10.085 20.18 10.255 ;
      RECT 16.6 9.345 16.77 9.515 ;
      RECT 16.6 10.085 16.77 10.255 ;
      RECT 16.23 8.605 16.4 8.775 ;
    LAYER li1 ;
      RECT 103.355 7.305 103.525 8.775 ;
      RECT 103.355 7.305 103.53 8.565 ;
      RECT 102.985 9.255 103.455 9.425 ;
      RECT 102.985 8.235 103.155 9.425 ;
      RECT 102.98 3.035 103.15 4.225 ;
      RECT 102.98 3.035 103.45 3.205 ;
      RECT 102.365 3.895 102.54 5.155 ;
      RECT 102.365 3.685 102.535 5.155 ;
      RECT 102.365 7.305 102.535 8.775 ;
      RECT 102.365 7.305 102.54 8.565 ;
      RECT 101.995 3.035 102.165 4.225 ;
      RECT 101.995 3.035 102.465 3.205 ;
      RECT 101.995 9.255 102.465 9.425 ;
      RECT 101.995 8.235 102.165 9.425 ;
      RECT 101.005 4.015 101.18 5.155 ;
      RECT 101.005 1.865 101.175 5.155 ;
      RECT 101.005 1.865 101.18 2.415 ;
      RECT 101.005 10.045 101.18 10.595 ;
      RECT 101.005 7.305 101.175 10.595 ;
      RECT 101.005 7.305 101.18 8.445 ;
      RECT 100.575 3.895 100.75 5.155 ;
      RECT 100.575 2.945 100.745 5.155 ;
      RECT 100.575 7.305 100.745 9.515 ;
      RECT 100.575 7.305 100.75 8.565 ;
      RECT 100.145 3.925 100.315 5.155 ;
      RECT 100.205 2.145 100.375 4.095 ;
      RECT 100.145 1.865 100.315 2.315 ;
      RECT 100.145 10.145 100.315 10.595 ;
      RECT 100.205 8.365 100.375 10.315 ;
      RECT 100.145 7.305 100.315 8.535 ;
      RECT 99.62 3.895 99.795 5.155 ;
      RECT 99.62 1.865 99.79 5.155 ;
      RECT 99.62 3.365 100.03 3.695 ;
      RECT 99.62 2.525 100.03 2.855 ;
      RECT 99.62 1.865 99.795 2.355 ;
      RECT 99.62 10.105 99.795 10.595 ;
      RECT 99.62 7.305 99.79 10.595 ;
      RECT 99.62 9.605 100.03 9.935 ;
      RECT 99.62 8.765 100.03 9.095 ;
      RECT 99.62 7.305 99.795 8.565 ;
      RECT 97.36 4.79 97.74 5.47 ;
      RECT 97.57 3.66 97.74 5.47 ;
      RECT 95.49 3.66 95.72 4.33 ;
      RECT 95.49 3.66 97.74 3.83 ;
      RECT 97.02 3.34 97.19 3.83 ;
      RECT 97.01 4.45 97.18 5.3 ;
      RECT 96.095 4.45 97.4 4.62 ;
      RECT 97.155 4 97.4 4.62 ;
      RECT 96.095 4.08 96.265 4.62 ;
      RECT 95.89 4.08 96.265 4.25 ;
      RECT 96.07 7.56 96.765 8.19 ;
      RECT 96.595 5.98 96.765 8.19 ;
      RECT 96.5 5.98 96.83 6.96 ;
      RECT 96.1 4.79 96.43 5.47 ;
      RECT 95.19 4.79 95.59 5.47 ;
      RECT 95.19 4.79 96.43 4.96 ;
      RECT 94.69 4.37 95.01 5.47 ;
      RECT 94.69 4.37 95.14 4.62 ;
      RECT 94.69 4.37 95.32 4.54 ;
      RECT 95.15 3.32 95.32 4.54 ;
      RECT 95.15 3.32 96.105 3.49 ;
      RECT 94.69 7.56 95.385 8.19 ;
      RECT 95.215 5.98 95.385 8.19 ;
      RECT 95.12 5.98 95.45 6.96 ;
      RECT 94.71 7.12 95.045 7.37 ;
      RECT 94.165 7.12 94.5 7.37 ;
      RECT 94.165 7.17 95.045 7.34 ;
      RECT 93.825 7.56 94.52 8.19 ;
      RECT 93.825 5.98 93.995 8.19 ;
      RECT 93.76 5.98 94.09 6.96 ;
      RECT 93.32 4.5 93.65 5.455 ;
      RECT 93.32 4.5 94 4.67 ;
      RECT 93.83 3.26 94 4.67 ;
      RECT 93.74 3.26 94.07 3.9 ;
      RECT 92.8 4.5 93.13 5.455 ;
      RECT 92.45 4.5 93.13 4.67 ;
      RECT 92.45 3.26 92.62 4.67 ;
      RECT 92.38 3.26 92.71 3.9 ;
      RECT 92.59 7.17 92.76 8.02 ;
      RECT 91.865 7.12 92.2 7.37 ;
      RECT 91.865 7.17 92.76 7.34 ;
      RECT 91.93 4.08 92.28 4.33 ;
      RECT 91.41 4.08 91.74 4.33 ;
      RECT 91.41 4.11 92.28 4.28 ;
      RECT 91.525 7.56 92.22 8.19 ;
      RECT 91.525 5.98 91.695 8.19 ;
      RECT 91.46 5.98 91.79 6.96 ;
      RECT 90.99 4.49 91.32 5.47 ;
      RECT 90.99 3.26 91.24 5.47 ;
      RECT 90.99 3.26 91.32 3.89 ;
      RECT 89.32 10.045 89.495 10.595 ;
      RECT 89.32 7.305 89.49 10.595 ;
      RECT 89.32 7.305 89.495 8.445 ;
      RECT 88.89 7.305 89.06 9.515 ;
      RECT 88.89 7.305 89.065 8.565 ;
      RECT 87.935 10.105 88.11 10.595 ;
      RECT 87.935 7.305 88.105 10.595 ;
      RECT 87.935 9.605 88.345 9.935 ;
      RECT 87.935 8.765 88.345 9.095 ;
      RECT 87.935 7.305 88.11 8.565 ;
      RECT 86.135 7.305 86.305 8.775 ;
      RECT 86.135 7.305 86.31 8.565 ;
      RECT 85.765 9.255 86.235 9.425 ;
      RECT 85.765 8.235 85.935 9.425 ;
      RECT 85.76 3.035 85.93 4.225 ;
      RECT 85.76 3.035 86.23 3.205 ;
      RECT 85.145 3.895 85.32 5.155 ;
      RECT 85.145 3.685 85.315 5.155 ;
      RECT 85.145 7.305 85.315 8.775 ;
      RECT 85.145 7.305 85.32 8.565 ;
      RECT 84.775 3.035 84.945 4.225 ;
      RECT 84.775 3.035 85.245 3.205 ;
      RECT 84.775 9.255 85.245 9.425 ;
      RECT 84.775 8.235 84.945 9.425 ;
      RECT 83.785 4.015 83.96 5.155 ;
      RECT 83.785 1.865 83.955 5.155 ;
      RECT 83.785 1.865 83.96 2.415 ;
      RECT 83.785 10.045 83.96 10.595 ;
      RECT 83.785 7.305 83.955 10.595 ;
      RECT 83.785 7.305 83.96 8.445 ;
      RECT 83.355 3.895 83.53 5.155 ;
      RECT 83.355 2.945 83.525 5.155 ;
      RECT 83.355 7.305 83.525 9.515 ;
      RECT 83.355 7.305 83.53 8.565 ;
      RECT 82.925 3.925 83.095 5.155 ;
      RECT 82.985 2.145 83.155 4.095 ;
      RECT 82.925 1.865 83.095 2.315 ;
      RECT 82.925 10.145 83.095 10.595 ;
      RECT 82.985 8.365 83.155 10.315 ;
      RECT 82.925 7.305 83.095 8.535 ;
      RECT 82.4 3.895 82.575 5.155 ;
      RECT 82.4 1.865 82.57 5.155 ;
      RECT 82.4 3.365 82.81 3.695 ;
      RECT 82.4 2.525 82.81 2.855 ;
      RECT 82.4 1.865 82.575 2.355 ;
      RECT 82.4 10.105 82.575 10.595 ;
      RECT 82.4 7.305 82.57 10.595 ;
      RECT 82.4 9.605 82.81 9.935 ;
      RECT 82.4 8.765 82.81 9.095 ;
      RECT 82.4 7.305 82.575 8.565 ;
      RECT 80.14 4.79 80.52 5.47 ;
      RECT 80.35 3.66 80.52 5.47 ;
      RECT 78.27 3.66 78.5 4.33 ;
      RECT 78.27 3.66 80.52 3.83 ;
      RECT 79.8 3.34 79.97 3.83 ;
      RECT 79.79 4.45 79.96 5.3 ;
      RECT 78.875 4.45 80.18 4.62 ;
      RECT 79.935 4 80.18 4.62 ;
      RECT 78.875 4.08 79.045 4.62 ;
      RECT 78.67 4.08 79.045 4.25 ;
      RECT 78.85 7.56 79.545 8.19 ;
      RECT 79.375 5.98 79.545 8.19 ;
      RECT 79.28 5.98 79.61 6.96 ;
      RECT 78.88 4.79 79.21 5.47 ;
      RECT 77.97 4.79 78.37 5.47 ;
      RECT 77.97 4.79 79.21 4.96 ;
      RECT 77.47 4.37 77.79 5.47 ;
      RECT 77.47 4.37 77.92 4.62 ;
      RECT 77.47 4.37 78.1 4.54 ;
      RECT 77.93 3.32 78.1 4.54 ;
      RECT 77.93 3.32 78.885 3.49 ;
      RECT 77.47 7.56 78.165 8.19 ;
      RECT 77.995 5.98 78.165 8.19 ;
      RECT 77.9 5.98 78.23 6.96 ;
      RECT 77.49 7.12 77.825 7.37 ;
      RECT 76.945 7.12 77.28 7.37 ;
      RECT 76.945 7.17 77.825 7.34 ;
      RECT 76.605 7.56 77.3 8.19 ;
      RECT 76.605 5.98 76.775 8.19 ;
      RECT 76.54 5.98 76.87 6.96 ;
      RECT 76.1 4.5 76.43 5.455 ;
      RECT 76.1 4.5 76.78 4.67 ;
      RECT 76.61 3.26 76.78 4.67 ;
      RECT 76.52 3.26 76.85 3.9 ;
      RECT 75.58 4.5 75.91 5.455 ;
      RECT 75.23 4.5 75.91 4.67 ;
      RECT 75.23 3.26 75.4 4.67 ;
      RECT 75.16 3.26 75.49 3.9 ;
      RECT 75.37 7.17 75.54 8.02 ;
      RECT 74.645 7.12 74.98 7.37 ;
      RECT 74.645 7.17 75.54 7.34 ;
      RECT 74.71 4.08 75.06 4.33 ;
      RECT 74.19 4.08 74.52 4.33 ;
      RECT 74.19 4.11 75.06 4.28 ;
      RECT 74.305 7.56 75 8.19 ;
      RECT 74.305 5.98 74.475 8.19 ;
      RECT 74.24 5.98 74.57 6.96 ;
      RECT 73.77 4.49 74.1 5.47 ;
      RECT 73.77 3.26 74.02 5.47 ;
      RECT 73.77 3.26 74.1 3.89 ;
      RECT 72.1 10.045 72.275 10.595 ;
      RECT 72.1 7.305 72.27 10.595 ;
      RECT 72.1 7.305 72.275 8.445 ;
      RECT 71.67 7.305 71.84 9.515 ;
      RECT 71.67 7.305 71.845 8.565 ;
      RECT 70.715 10.105 70.89 10.595 ;
      RECT 70.715 7.305 70.885 10.595 ;
      RECT 70.715 9.605 71.125 9.935 ;
      RECT 70.715 8.765 71.125 9.095 ;
      RECT 70.715 7.305 70.89 8.565 ;
      RECT 68.915 7.31 69.085 8.78 ;
      RECT 68.915 7.31 69.09 8.57 ;
      RECT 68.545 9.26 69.015 9.43 ;
      RECT 68.545 8.24 68.715 9.43 ;
      RECT 68.54 3.04 68.71 4.23 ;
      RECT 68.54 3.04 69.01 3.21 ;
      RECT 67.925 3.9 68.1 5.16 ;
      RECT 67.925 3.69 68.095 5.16 ;
      RECT 67.925 7.31 68.095 8.78 ;
      RECT 67.925 7.31 68.1 8.57 ;
      RECT 67.555 3.04 67.725 4.23 ;
      RECT 67.555 3.04 68.025 3.21 ;
      RECT 67.555 9.26 68.025 9.43 ;
      RECT 67.555 8.24 67.725 9.43 ;
      RECT 66.565 4.02 66.74 5.16 ;
      RECT 66.565 1.87 66.735 5.16 ;
      RECT 66.565 1.87 66.74 2.42 ;
      RECT 66.565 10.05 66.74 10.6 ;
      RECT 66.565 7.31 66.735 10.6 ;
      RECT 66.565 7.31 66.74 8.45 ;
      RECT 66.135 3.9 66.31 5.16 ;
      RECT 66.135 2.95 66.305 5.16 ;
      RECT 66.135 7.31 66.305 9.52 ;
      RECT 66.135 7.31 66.31 8.57 ;
      RECT 65.705 3.93 65.875 5.16 ;
      RECT 65.765 2.15 65.935 4.1 ;
      RECT 65.705 1.87 65.875 2.32 ;
      RECT 65.705 10.15 65.875 10.6 ;
      RECT 65.765 8.37 65.935 10.32 ;
      RECT 65.705 7.31 65.875 8.54 ;
      RECT 65.18 3.9 65.355 5.16 ;
      RECT 65.18 1.87 65.35 5.16 ;
      RECT 65.18 3.37 65.59 3.7 ;
      RECT 65.18 2.53 65.59 2.86 ;
      RECT 65.18 1.87 65.355 2.36 ;
      RECT 65.18 10.11 65.355 10.6 ;
      RECT 65.18 7.31 65.35 10.6 ;
      RECT 65.18 9.61 65.59 9.94 ;
      RECT 65.18 8.77 65.59 9.1 ;
      RECT 65.18 7.31 65.355 8.57 ;
      RECT 62.92 4.795 63.3 5.475 ;
      RECT 63.13 3.665 63.3 5.475 ;
      RECT 61.05 3.665 61.28 4.335 ;
      RECT 61.05 3.665 63.3 3.835 ;
      RECT 62.58 3.345 62.75 3.835 ;
      RECT 62.57 4.455 62.74 5.305 ;
      RECT 61.655 4.455 62.96 4.625 ;
      RECT 62.715 4.005 62.96 4.625 ;
      RECT 61.655 4.085 61.825 4.625 ;
      RECT 61.45 4.085 61.825 4.255 ;
      RECT 61.63 7.565 62.325 8.195 ;
      RECT 62.155 5.985 62.325 8.195 ;
      RECT 62.06 5.985 62.39 6.965 ;
      RECT 61.66 4.795 61.99 5.475 ;
      RECT 60.75 4.795 61.15 5.475 ;
      RECT 60.75 4.795 61.99 4.965 ;
      RECT 60.25 4.375 60.57 5.475 ;
      RECT 60.25 4.375 60.7 4.625 ;
      RECT 60.25 4.375 60.88 4.545 ;
      RECT 60.71 3.325 60.88 4.545 ;
      RECT 60.71 3.325 61.665 3.495 ;
      RECT 60.25 7.565 60.945 8.195 ;
      RECT 60.775 5.985 60.945 8.195 ;
      RECT 60.68 5.985 61.01 6.965 ;
      RECT 60.27 7.125 60.605 7.375 ;
      RECT 59.725 7.125 60.06 7.375 ;
      RECT 59.725 7.175 60.605 7.345 ;
      RECT 59.385 7.565 60.08 8.195 ;
      RECT 59.385 5.985 59.555 8.195 ;
      RECT 59.32 5.985 59.65 6.965 ;
      RECT 58.88 4.505 59.21 5.46 ;
      RECT 58.88 4.505 59.56 4.675 ;
      RECT 59.39 3.265 59.56 4.675 ;
      RECT 59.3 3.265 59.63 3.905 ;
      RECT 58.36 4.505 58.69 5.46 ;
      RECT 58.01 4.505 58.69 4.675 ;
      RECT 58.01 3.265 58.18 4.675 ;
      RECT 57.94 3.265 58.27 3.905 ;
      RECT 58.15 7.175 58.32 8.025 ;
      RECT 57.425 7.125 57.76 7.375 ;
      RECT 57.425 7.175 58.32 7.345 ;
      RECT 57.49 4.085 57.84 4.335 ;
      RECT 56.97 4.085 57.3 4.335 ;
      RECT 56.97 4.115 57.84 4.285 ;
      RECT 57.085 7.565 57.78 8.195 ;
      RECT 57.085 5.985 57.255 8.195 ;
      RECT 57.02 5.985 57.35 6.965 ;
      RECT 56.55 4.495 56.88 5.475 ;
      RECT 56.55 3.265 56.8 5.475 ;
      RECT 56.55 3.265 56.88 3.895 ;
      RECT 54.88 10.05 55.055 10.6 ;
      RECT 54.88 7.31 55.05 10.6 ;
      RECT 54.88 7.31 55.055 8.45 ;
      RECT 54.45 7.31 54.62 9.52 ;
      RECT 54.45 7.31 54.625 8.57 ;
      RECT 53.495 10.11 53.67 10.6 ;
      RECT 53.495 7.31 53.665 10.6 ;
      RECT 53.495 9.61 53.905 9.94 ;
      RECT 53.495 8.77 53.905 9.1 ;
      RECT 53.495 7.31 53.67 8.57 ;
      RECT 51.695 7.305 51.865 8.775 ;
      RECT 51.695 7.305 51.87 8.565 ;
      RECT 51.325 9.255 51.795 9.425 ;
      RECT 51.325 8.235 51.495 9.425 ;
      RECT 51.32 3.035 51.49 4.225 ;
      RECT 51.32 3.035 51.79 3.205 ;
      RECT 50.705 3.895 50.88 5.155 ;
      RECT 50.705 3.685 50.875 5.155 ;
      RECT 50.705 7.305 50.875 8.775 ;
      RECT 50.705 7.305 50.88 8.565 ;
      RECT 50.335 3.035 50.505 4.225 ;
      RECT 50.335 3.035 50.805 3.205 ;
      RECT 50.335 9.255 50.805 9.425 ;
      RECT 50.335 8.235 50.505 9.425 ;
      RECT 49.345 4.015 49.52 5.155 ;
      RECT 49.345 1.865 49.515 5.155 ;
      RECT 49.345 1.865 49.52 2.415 ;
      RECT 49.345 10.045 49.52 10.595 ;
      RECT 49.345 7.305 49.515 10.595 ;
      RECT 49.345 7.305 49.52 8.445 ;
      RECT 48.915 3.895 49.09 5.155 ;
      RECT 48.915 2.945 49.085 5.155 ;
      RECT 48.915 7.305 49.085 9.515 ;
      RECT 48.915 7.305 49.09 8.565 ;
      RECT 48.485 3.925 48.655 5.155 ;
      RECT 48.545 2.145 48.715 4.095 ;
      RECT 48.485 1.865 48.655 2.315 ;
      RECT 48.485 10.145 48.655 10.595 ;
      RECT 48.545 8.365 48.715 10.315 ;
      RECT 48.485 7.305 48.655 8.535 ;
      RECT 47.96 3.895 48.135 5.155 ;
      RECT 47.96 1.865 48.13 5.155 ;
      RECT 47.96 3.365 48.37 3.695 ;
      RECT 47.96 2.525 48.37 2.855 ;
      RECT 47.96 1.865 48.135 2.355 ;
      RECT 47.96 10.105 48.135 10.595 ;
      RECT 47.96 7.305 48.13 10.595 ;
      RECT 47.96 9.605 48.37 9.935 ;
      RECT 47.96 8.765 48.37 9.095 ;
      RECT 47.96 7.305 48.135 8.565 ;
      RECT 45.7 4.79 46.08 5.47 ;
      RECT 45.91 3.66 46.08 5.47 ;
      RECT 43.83 3.66 44.06 4.33 ;
      RECT 43.83 3.66 46.08 3.83 ;
      RECT 45.36 3.34 45.53 3.83 ;
      RECT 45.35 4.45 45.52 5.3 ;
      RECT 44.435 4.45 45.74 4.62 ;
      RECT 45.495 4 45.74 4.62 ;
      RECT 44.435 4.08 44.605 4.62 ;
      RECT 44.23 4.08 44.605 4.25 ;
      RECT 44.41 7.56 45.105 8.19 ;
      RECT 44.935 5.98 45.105 8.19 ;
      RECT 44.84 5.98 45.17 6.96 ;
      RECT 44.44 4.79 44.77 5.47 ;
      RECT 43.53 4.79 43.93 5.47 ;
      RECT 43.53 4.79 44.77 4.96 ;
      RECT 43.03 4.37 43.35 5.47 ;
      RECT 43.03 4.37 43.48 4.62 ;
      RECT 43.03 4.37 43.66 4.54 ;
      RECT 43.49 3.32 43.66 4.54 ;
      RECT 43.49 3.32 44.445 3.49 ;
      RECT 43.03 7.56 43.725 8.19 ;
      RECT 43.555 5.98 43.725 8.19 ;
      RECT 43.46 5.98 43.79 6.96 ;
      RECT 43.05 7.12 43.385 7.37 ;
      RECT 42.505 7.12 42.84 7.37 ;
      RECT 42.505 7.17 43.385 7.34 ;
      RECT 42.165 7.56 42.86 8.19 ;
      RECT 42.165 5.98 42.335 8.19 ;
      RECT 42.1 5.98 42.43 6.96 ;
      RECT 41.66 4.5 41.99 5.455 ;
      RECT 41.66 4.5 42.34 4.67 ;
      RECT 42.17 3.26 42.34 4.67 ;
      RECT 42.08 3.26 42.41 3.9 ;
      RECT 41.14 4.5 41.47 5.455 ;
      RECT 40.79 4.5 41.47 4.67 ;
      RECT 40.79 3.26 40.96 4.67 ;
      RECT 40.72 3.26 41.05 3.9 ;
      RECT 40.93 7.17 41.1 8.02 ;
      RECT 40.205 7.12 40.54 7.37 ;
      RECT 40.205 7.17 41.1 7.34 ;
      RECT 40.27 4.08 40.62 4.33 ;
      RECT 39.75 4.08 40.08 4.33 ;
      RECT 39.75 4.11 40.62 4.28 ;
      RECT 39.865 7.56 40.56 8.19 ;
      RECT 39.865 5.98 40.035 8.19 ;
      RECT 39.8 5.98 40.13 6.96 ;
      RECT 39.33 4.49 39.66 5.47 ;
      RECT 39.33 3.26 39.58 5.47 ;
      RECT 39.33 3.26 39.66 3.89 ;
      RECT 37.66 10.045 37.835 10.595 ;
      RECT 37.66 7.305 37.83 10.595 ;
      RECT 37.66 7.305 37.835 8.445 ;
      RECT 37.23 7.305 37.4 9.515 ;
      RECT 37.23 7.305 37.405 8.565 ;
      RECT 36.275 10.105 36.45 10.595 ;
      RECT 36.275 7.305 36.445 10.595 ;
      RECT 36.275 9.605 36.685 9.935 ;
      RECT 36.275 8.765 36.685 9.095 ;
      RECT 36.275 7.305 36.45 8.565 ;
      RECT 34.475 7.305 34.645 8.775 ;
      RECT 34.475 7.305 34.65 8.565 ;
      RECT 34.105 9.255 34.575 9.425 ;
      RECT 34.105 8.235 34.275 9.425 ;
      RECT 34.1 3.035 34.27 4.225 ;
      RECT 34.1 3.035 34.57 3.205 ;
      RECT 33.485 3.895 33.66 5.155 ;
      RECT 33.485 3.685 33.655 5.155 ;
      RECT 33.485 7.305 33.655 8.775 ;
      RECT 33.485 7.305 33.66 8.565 ;
      RECT 33.115 3.035 33.285 4.225 ;
      RECT 33.115 3.035 33.585 3.205 ;
      RECT 33.115 9.255 33.585 9.425 ;
      RECT 33.115 8.235 33.285 9.425 ;
      RECT 32.125 4.015 32.3 5.155 ;
      RECT 32.125 1.865 32.295 5.155 ;
      RECT 32.125 1.865 32.3 2.415 ;
      RECT 32.125 10.045 32.3 10.595 ;
      RECT 32.125 7.305 32.295 10.595 ;
      RECT 32.125 7.305 32.3 8.445 ;
      RECT 31.695 3.895 31.87 5.155 ;
      RECT 31.695 2.945 31.865 5.155 ;
      RECT 31.695 7.305 31.865 9.515 ;
      RECT 31.695 7.305 31.87 8.565 ;
      RECT 31.265 3.925 31.435 5.155 ;
      RECT 31.325 2.145 31.495 4.095 ;
      RECT 31.265 1.865 31.435 2.315 ;
      RECT 31.265 10.145 31.435 10.595 ;
      RECT 31.325 8.365 31.495 10.315 ;
      RECT 31.265 7.305 31.435 8.535 ;
      RECT 30.74 3.895 30.915 5.155 ;
      RECT 30.74 1.865 30.91 5.155 ;
      RECT 30.74 3.365 31.15 3.695 ;
      RECT 30.74 2.525 31.15 2.855 ;
      RECT 30.74 1.865 30.915 2.355 ;
      RECT 30.74 10.105 30.915 10.595 ;
      RECT 30.74 7.305 30.91 10.595 ;
      RECT 30.74 9.605 31.15 9.935 ;
      RECT 30.74 8.765 31.15 9.095 ;
      RECT 30.74 7.305 30.915 8.565 ;
      RECT 28.48 4.79 28.86 5.47 ;
      RECT 28.69 3.66 28.86 5.47 ;
      RECT 26.61 3.66 26.84 4.33 ;
      RECT 26.61 3.66 28.86 3.83 ;
      RECT 28.14 3.34 28.31 3.83 ;
      RECT 28.13 4.45 28.3 5.3 ;
      RECT 27.215 4.45 28.52 4.62 ;
      RECT 28.275 4 28.52 4.62 ;
      RECT 27.215 4.08 27.385 4.62 ;
      RECT 27.01 4.08 27.385 4.25 ;
      RECT 27.19 7.56 27.885 8.19 ;
      RECT 27.715 5.98 27.885 8.19 ;
      RECT 27.62 5.98 27.95 6.96 ;
      RECT 27.22 4.79 27.55 5.47 ;
      RECT 26.31 4.79 26.71 5.47 ;
      RECT 26.31 4.79 27.55 4.96 ;
      RECT 25.81 4.37 26.13 5.47 ;
      RECT 25.81 4.37 26.26 4.62 ;
      RECT 25.81 4.37 26.44 4.54 ;
      RECT 26.27 3.32 26.44 4.54 ;
      RECT 26.27 3.32 27.225 3.49 ;
      RECT 25.81 7.56 26.505 8.19 ;
      RECT 26.335 5.98 26.505 8.19 ;
      RECT 26.24 5.98 26.57 6.96 ;
      RECT 25.83 7.12 26.165 7.37 ;
      RECT 25.285 7.12 25.62 7.37 ;
      RECT 25.285 7.17 26.165 7.34 ;
      RECT 24.945 7.56 25.64 8.19 ;
      RECT 24.945 5.98 25.115 8.19 ;
      RECT 24.88 5.98 25.21 6.96 ;
      RECT 24.44 4.5 24.77 5.455 ;
      RECT 24.44 4.5 25.12 4.67 ;
      RECT 24.95 3.26 25.12 4.67 ;
      RECT 24.86 3.26 25.19 3.9 ;
      RECT 23.92 4.5 24.25 5.455 ;
      RECT 23.57 4.5 24.25 4.67 ;
      RECT 23.57 3.26 23.74 4.67 ;
      RECT 23.5 3.26 23.83 3.9 ;
      RECT 23.71 7.17 23.88 8.02 ;
      RECT 22.985 7.12 23.32 7.37 ;
      RECT 22.985 7.17 23.88 7.34 ;
      RECT 23.05 4.08 23.4 4.33 ;
      RECT 22.53 4.08 22.86 4.33 ;
      RECT 22.53 4.11 23.4 4.28 ;
      RECT 22.645 7.56 23.34 8.19 ;
      RECT 22.645 5.98 22.815 8.19 ;
      RECT 22.58 5.98 22.91 6.96 ;
      RECT 22.11 4.49 22.44 5.47 ;
      RECT 22.11 3.26 22.36 5.47 ;
      RECT 22.11 3.26 22.44 3.89 ;
      RECT 20.44 10.045 20.615 10.595 ;
      RECT 20.44 7.305 20.61 10.595 ;
      RECT 20.44 7.305 20.615 8.445 ;
      RECT 20.01 7.305 20.18 9.515 ;
      RECT 20.01 7.305 20.185 8.565 ;
      RECT 19.055 10.105 19.23 10.595 ;
      RECT 19.055 7.305 19.225 10.595 ;
      RECT 19.055 9.605 19.465 9.935 ;
      RECT 19.055 8.765 19.465 9.095 ;
      RECT 19.055 7.305 19.23 8.565 ;
      RECT 16.6 7.305 16.77 9.515 ;
      RECT 16.6 7.305 16.775 8.565 ;
      RECT 16.17 10.145 16.34 10.595 ;
      RECT 16.23 8.365 16.4 10.315 ;
      RECT 16.17 7.305 16.34 8.535 ;
      RECT 15.645 10.105 15.82 10.595 ;
      RECT 15.645 7.305 15.815 10.595 ;
      RECT 15.645 9.605 16.055 9.935 ;
      RECT 15.645 8.765 16.055 9.095 ;
      RECT 15.645 7.305 15.82 8.565 ;
      RECT 103.355 10.085 103.53 10.595 ;
      RECT 102.365 1.865 102.54 2.375 ;
      RECT 102.365 10.085 102.54 10.595 ;
      RECT 100.575 1.865 100.75 2.375 ;
      RECT 100.575 10.085 100.75 10.595 ;
      RECT 96.935 7.12 97.27 7.39 ;
      RECT 96.435 4.08 96.985 4.28 ;
      RECT 96.09 7.12 96.425 7.37 ;
      RECT 95.555 7.12 95.89 7.39 ;
      RECT 94.17 4.08 94.52 4.33 ;
      RECT 93.31 4.08 93.66 4.33 ;
      RECT 92.79 4.08 93.14 4.33 ;
      RECT 88.89 10.085 89.065 10.595 ;
      RECT 86.135 10.085 86.31 10.595 ;
      RECT 85.145 1.865 85.32 2.375 ;
      RECT 85.145 10.085 85.32 10.595 ;
      RECT 83.355 1.865 83.53 2.375 ;
      RECT 83.355 10.085 83.53 10.595 ;
      RECT 79.715 7.12 80.05 7.39 ;
      RECT 79.215 4.08 79.765 4.28 ;
      RECT 78.87 7.12 79.205 7.37 ;
      RECT 78.335 7.12 78.67 7.39 ;
      RECT 76.95 4.08 77.3 4.33 ;
      RECT 76.09 4.08 76.44 4.33 ;
      RECT 75.57 4.08 75.92 4.33 ;
      RECT 71.67 10.085 71.845 10.595 ;
      RECT 68.915 10.09 69.09 10.6 ;
      RECT 67.925 1.87 68.1 2.38 ;
      RECT 67.925 10.09 68.1 10.6 ;
      RECT 66.135 1.87 66.31 2.38 ;
      RECT 66.135 10.09 66.31 10.6 ;
      RECT 62.495 7.125 62.83 7.395 ;
      RECT 61.995 4.085 62.545 4.285 ;
      RECT 61.65 7.125 61.985 7.375 ;
      RECT 61.115 7.125 61.45 7.395 ;
      RECT 59.73 4.085 60.08 4.335 ;
      RECT 58.87 4.085 59.22 4.335 ;
      RECT 58.35 4.085 58.7 4.335 ;
      RECT 54.45 10.09 54.625 10.6 ;
      RECT 51.695 10.085 51.87 10.595 ;
      RECT 50.705 1.865 50.88 2.375 ;
      RECT 50.705 10.085 50.88 10.595 ;
      RECT 48.915 1.865 49.09 2.375 ;
      RECT 48.915 10.085 49.09 10.595 ;
      RECT 45.275 7.12 45.61 7.39 ;
      RECT 44.775 4.08 45.325 4.28 ;
      RECT 44.43 7.12 44.765 7.37 ;
      RECT 43.895 7.12 44.23 7.39 ;
      RECT 42.51 4.08 42.86 4.33 ;
      RECT 41.65 4.08 42 4.33 ;
      RECT 41.13 4.08 41.48 4.33 ;
      RECT 37.23 10.085 37.405 10.595 ;
      RECT 34.475 10.085 34.65 10.595 ;
      RECT 33.485 1.865 33.66 2.375 ;
      RECT 33.485 10.085 33.66 10.595 ;
      RECT 31.695 1.865 31.87 2.375 ;
      RECT 31.695 10.085 31.87 10.595 ;
      RECT 28.055 7.12 28.39 7.39 ;
      RECT 27.555 4.08 28.105 4.28 ;
      RECT 27.21 7.12 27.545 7.37 ;
      RECT 26.675 7.12 27.01 7.39 ;
      RECT 25.29 4.08 25.64 4.33 ;
      RECT 24.43 4.08 24.78 4.33 ;
      RECT 23.91 4.08 24.26 4.33 ;
      RECT 20.01 10.085 20.185 10.595 ;
      RECT 16.6 10.085 16.775 10.595 ;
  END
END sky130_osu_ring_oscillator_mpr2ct_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2ea_8_b0r1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ea_8_b0r1 ;
  SIZE 99.43 BY 12.46 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 33.48 0 33.86 5.265 ;
      LAYER met2 ;
        RECT 33.48 4.885 33.86 5.265 ;
      LAYER li1 ;
        RECT 33.58 1.87 33.755 2.38 ;
        RECT 33.58 3.9 33.755 5.16 ;
        RECT 33.58 3.69 33.75 5.16 ;
      LAYER met1 ;
        RECT 33.495 4.93 33.845 5.22 ;
        RECT 33.52 2.18 33.815 2.41 ;
        RECT 33.52 3.66 33.81 3.89 ;
        RECT 33.58 2.18 33.75 3.89 ;
      LAYER via1 ;
        RECT 33.595 5 33.745 5.15 ;
      LAYER via2 ;
        RECT 33.57 4.975 33.77 5.175 ;
      LAYER mcon ;
        RECT 33.58 3.69 33.75 3.86 ;
        RECT 33.58 2.21 33.75 2.38 ;
        RECT 33.585 4.99 33.755 5.16 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 49.805 0 50.185 5.265 ;
      LAYER met2 ;
        RECT 49.805 4.885 50.185 5.265 ;
      LAYER li1 ;
        RECT 49.905 1.87 50.08 2.38 ;
        RECT 49.905 3.9 50.08 5.16 ;
        RECT 49.905 3.69 50.075 5.16 ;
      LAYER met1 ;
        RECT 49.82 4.93 50.17 5.22 ;
        RECT 49.845 2.18 50.14 2.41 ;
        RECT 49.845 3.66 50.135 3.89 ;
        RECT 49.905 2.18 50.075 3.89 ;
      LAYER via1 ;
        RECT 49.92 5 50.07 5.15 ;
      LAYER via2 ;
        RECT 49.895 4.975 50.095 5.175 ;
      LAYER mcon ;
        RECT 49.905 3.69 50.075 3.86 ;
        RECT 49.905 2.21 50.075 2.38 ;
        RECT 49.91 4.99 50.08 5.16 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 66.13 0 66.51 5.265 ;
      LAYER met2 ;
        RECT 66.13 4.885 66.51 5.265 ;
      LAYER li1 ;
        RECT 66.23 1.87 66.405 2.38 ;
        RECT 66.23 3.9 66.405 5.16 ;
        RECT 66.23 3.69 66.4 5.16 ;
      LAYER met1 ;
        RECT 66.145 4.93 66.495 5.22 ;
        RECT 66.17 2.18 66.465 2.41 ;
        RECT 66.17 3.66 66.46 3.89 ;
        RECT 66.23 2.18 66.4 3.89 ;
      LAYER via1 ;
        RECT 66.245 5 66.395 5.15 ;
      LAYER via2 ;
        RECT 66.22 4.975 66.42 5.175 ;
      LAYER mcon ;
        RECT 66.23 3.69 66.4 3.86 ;
        RECT 66.23 2.21 66.4 2.38 ;
        RECT 66.235 4.99 66.405 5.16 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 82.455 0 82.835 5.265 ;
      LAYER met2 ;
        RECT 82.455 4.885 82.835 5.265 ;
      LAYER li1 ;
        RECT 82.555 1.87 82.73 2.38 ;
        RECT 82.555 3.9 82.73 5.16 ;
        RECT 82.555 3.69 82.725 5.16 ;
      LAYER met1 ;
        RECT 82.47 4.93 82.82 5.22 ;
        RECT 82.495 2.18 82.79 2.41 ;
        RECT 82.495 3.66 82.785 3.89 ;
        RECT 82.555 2.18 82.725 3.89 ;
      LAYER via1 ;
        RECT 82.57 5 82.72 5.15 ;
      LAYER via2 ;
        RECT 82.545 4.975 82.745 5.175 ;
      LAYER mcon ;
        RECT 82.555 3.69 82.725 3.86 ;
        RECT 82.555 2.21 82.725 2.38 ;
        RECT 82.56 4.99 82.73 5.16 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 98.78 0 99.16 5.265 ;
      LAYER met2 ;
        RECT 98.78 4.885 99.16 5.265 ;
      LAYER li1 ;
        RECT 98.88 1.87 99.055 2.38 ;
        RECT 98.88 3.9 99.055 5.16 ;
        RECT 98.88 3.69 99.05 5.16 ;
      LAYER met1 ;
        RECT 98.795 4.93 99.145 5.22 ;
        RECT 98.82 2.18 99.115 2.41 ;
        RECT 98.82 3.66 99.11 3.89 ;
        RECT 98.88 2.18 99.05 3.89 ;
      LAYER via1 ;
        RECT 98.895 5 99.045 5.15 ;
      LAYER via2 ;
        RECT 98.87 4.975 99.07 5.175 ;
      LAYER mcon ;
        RECT 98.88 3.69 99.05 3.86 ;
        RECT 98.88 2.21 99.05 2.38 ;
        RECT 98.885 4.99 99.055 5.16 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 29.355 4 29.695 4.35 ;
        RECT 29.345 8.125 29.685 8.475 ;
        RECT 29.43 4 29.6 8.475 ;
      LAYER li1 ;
        RECT 29.425 2.955 29.595 4.225 ;
        RECT 29.425 8.235 29.595 9.505 ;
        RECT 23.81 8.235 23.98 9.505 ;
      LAYER met1 ;
        RECT 29.355 4.055 29.825 4.225 ;
        RECT 29.355 4 29.695 4.35 ;
        RECT 29.345 8.235 29.825 8.405 ;
        RECT 29.345 8.125 29.685 8.475 ;
        RECT 23.75 8.23 29.685 8.4 ;
        RECT 23.75 8.23 24.21 8.405 ;
        RECT 23.75 8.205 24.04 8.435 ;
      LAYER via1 ;
        RECT 29.445 8.225 29.595 8.375 ;
        RECT 29.455 4.1 29.605 4.25 ;
      LAYER mcon ;
        RECT 23.81 8.235 23.98 8.405 ;
        RECT 29.425 8.235 29.595 8.405 ;
        RECT 29.425 4.055 29.595 4.225 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 45.68 4 46.02 4.35 ;
        RECT 45.67 8.125 46.01 8.475 ;
        RECT 45.755 4 45.925 8.475 ;
      LAYER li1 ;
        RECT 45.75 2.955 45.92 4.225 ;
        RECT 45.75 8.235 45.92 9.505 ;
        RECT 40.135 8.235 40.305 9.505 ;
      LAYER met1 ;
        RECT 45.68 4.055 46.15 4.225 ;
        RECT 45.68 4 46.02 4.35 ;
        RECT 45.67 8.235 46.15 8.405 ;
        RECT 45.67 8.125 46.01 8.475 ;
        RECT 40.075 8.23 46.01 8.4 ;
        RECT 40.075 8.23 40.535 8.405 ;
        RECT 40.075 8.205 40.365 8.435 ;
      LAYER via1 ;
        RECT 45.77 8.225 45.92 8.375 ;
        RECT 45.78 4.1 45.93 4.25 ;
      LAYER mcon ;
        RECT 40.135 8.235 40.305 8.405 ;
        RECT 45.75 8.235 45.92 8.405 ;
        RECT 45.75 4.055 45.92 4.225 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 62.005 4 62.345 4.35 ;
        RECT 61.995 8.125 62.335 8.475 ;
        RECT 62.08 4 62.25 8.475 ;
      LAYER li1 ;
        RECT 62.075 2.955 62.245 4.225 ;
        RECT 62.075 8.235 62.245 9.505 ;
        RECT 56.46 8.235 56.63 9.505 ;
      LAYER met1 ;
        RECT 62.005 4.055 62.475 4.225 ;
        RECT 62.005 4 62.345 4.35 ;
        RECT 61.995 8.235 62.475 8.405 ;
        RECT 61.995 8.125 62.335 8.475 ;
        RECT 56.4 8.23 62.335 8.4 ;
        RECT 56.4 8.23 56.86 8.405 ;
        RECT 56.4 8.205 56.69 8.435 ;
      LAYER via1 ;
        RECT 62.095 8.225 62.245 8.375 ;
        RECT 62.105 4.1 62.255 4.25 ;
      LAYER mcon ;
        RECT 56.46 8.235 56.63 8.405 ;
        RECT 62.075 8.235 62.245 8.405 ;
        RECT 62.075 4.055 62.245 4.225 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 78.33 4 78.67 4.35 ;
        RECT 78.32 8.125 78.66 8.475 ;
        RECT 78.405 4 78.575 8.475 ;
      LAYER li1 ;
        RECT 78.4 2.955 78.57 4.225 ;
        RECT 78.4 8.235 78.57 9.505 ;
        RECT 72.785 8.235 72.955 9.505 ;
      LAYER met1 ;
        RECT 78.33 4.055 78.8 4.225 ;
        RECT 78.33 4 78.67 4.35 ;
        RECT 78.32 8.235 78.8 8.405 ;
        RECT 78.32 8.125 78.66 8.475 ;
        RECT 72.725 8.23 78.66 8.4 ;
        RECT 72.725 8.23 73.185 8.405 ;
        RECT 72.725 8.205 73.015 8.435 ;
      LAYER via1 ;
        RECT 78.42 8.225 78.57 8.375 ;
        RECT 78.43 4.1 78.58 4.25 ;
      LAYER mcon ;
        RECT 72.785 8.235 72.955 8.405 ;
        RECT 78.4 8.235 78.57 8.405 ;
        RECT 78.4 4.055 78.57 4.225 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 94.655 4 94.995 4.35 ;
        RECT 94.645 8.125 94.985 8.475 ;
        RECT 94.73 4 94.9 8.475 ;
      LAYER li1 ;
        RECT 94.725 2.955 94.895 4.225 ;
        RECT 94.725 8.235 94.895 9.505 ;
        RECT 89.11 8.235 89.28 9.505 ;
      LAYER met1 ;
        RECT 94.655 4.055 95.125 4.225 ;
        RECT 94.655 4 94.995 4.35 ;
        RECT 94.645 8.235 95.125 8.405 ;
        RECT 94.645 8.125 94.985 8.475 ;
        RECT 89.05 8.23 94.985 8.4 ;
        RECT 89.05 8.23 89.51 8.405 ;
        RECT 89.05 8.205 89.34 8.435 ;
      LAYER via1 ;
        RECT 94.745 8.225 94.895 8.375 ;
        RECT 94.755 4.1 94.905 4.25 ;
      LAYER mcon ;
        RECT 89.11 8.235 89.28 8.405 ;
        RECT 94.725 8.235 94.895 8.405 ;
        RECT 94.725 4.055 94.895 4.225 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 15.23 8.235 15.4 9.505 ;
      LAYER met1 ;
        RECT 15.17 8.235 15.63 8.405 ;
        RECT 15.175 8.2 15.465 8.43 ;
        RECT 15.17 8.205 15.46 8.435 ;
      LAYER mcon ;
        RECT 15.23 8.235 15.4 8.405 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.005 5.43 99.425 7.03 ;
        RECT 98.455 5.43 98.625 7.76 ;
        RECT 98.45 4.7 98.62 7.03 ;
        RECT 94.545 5.425 98.28 7.035 ;
        RECT 97.46 4.695 97.63 7.765 ;
        RECT 94.715 4.695 94.885 7.765 ;
        RECT 92.93 4.93 93.1 7.03 ;
        RECT 91.97 4.93 92.14 7.03 ;
        RECT 88.93 5.43 91.68 7.035 ;
        RECT 89.53 4.93 89.7 7.035 ;
        RECT 89.1 5.43 89.27 7.765 ;
        RECT 88.53 4.93 88.7 7.03 ;
        RECT 87.57 4.93 87.74 7.03 ;
        RECT 85.13 4.93 85.3 7.03 ;
        RECT 82.13 5.43 82.3 7.76 ;
        RECT 82.125 4.7 82.295 7.03 ;
        RECT 78.22 5.425 81.955 7.035 ;
        RECT 81.135 4.695 81.305 7.765 ;
        RECT 78.39 4.695 78.56 7.765 ;
        RECT 76.605 4.93 76.775 7.03 ;
        RECT 75.645 4.93 75.815 7.03 ;
        RECT 72.605 5.43 75.355 7.035 ;
        RECT 73.205 4.93 73.375 7.035 ;
        RECT 72.775 5.43 72.945 7.765 ;
        RECT 72.205 4.93 72.375 7.03 ;
        RECT 71.245 4.93 71.415 7.03 ;
        RECT 68.805 4.93 68.975 7.03 ;
        RECT 65.805 5.43 65.975 7.76 ;
        RECT 65.8 4.7 65.97 7.03 ;
        RECT 61.895 5.425 65.63 7.035 ;
        RECT 64.81 4.695 64.98 7.765 ;
        RECT 62.065 4.695 62.235 7.765 ;
        RECT 60.28 4.93 60.45 7.03 ;
        RECT 59.32 4.93 59.49 7.03 ;
        RECT 56.28 5.43 59.03 7.035 ;
        RECT 56.88 4.93 57.05 7.035 ;
        RECT 56.45 5.43 56.62 7.765 ;
        RECT 55.88 4.93 56.05 7.03 ;
        RECT 54.92 4.93 55.09 7.03 ;
        RECT 52.48 4.93 52.65 7.03 ;
        RECT 49.48 5.43 49.65 7.76 ;
        RECT 49.475 4.7 49.645 7.03 ;
        RECT 45.57 5.425 49.305 7.035 ;
        RECT 48.485 4.695 48.655 7.765 ;
        RECT 45.74 4.695 45.91 7.765 ;
        RECT 43.955 4.93 44.125 7.03 ;
        RECT 42.995 4.93 43.165 7.03 ;
        RECT 39.955 5.43 42.705 7.035 ;
        RECT 40.555 4.93 40.725 7.035 ;
        RECT 40.125 5.43 40.295 7.765 ;
        RECT 39.555 4.93 39.725 7.03 ;
        RECT 38.595 4.93 38.765 7.03 ;
        RECT 36.155 4.93 36.325 7.03 ;
        RECT 33.155 5.43 33.325 7.76 ;
        RECT 33.15 4.7 33.32 7.03 ;
        RECT 29.245 5.425 32.98 7.035 ;
        RECT 32.16 4.695 32.33 7.765 ;
        RECT 29.415 4.695 29.585 7.765 ;
        RECT 27.63 4.93 27.8 7.03 ;
        RECT 26.67 4.93 26.84 7.03 ;
        RECT 23.63 5.43 26.38 7.035 ;
        RECT 24.23 4.93 24.4 7.035 ;
        RECT 23.8 5.43 23.97 7.765 ;
        RECT 23.23 4.93 23.4 7.03 ;
        RECT 22.27 4.93 22.44 7.03 ;
        RECT 19.83 4.93 20 7.03 ;
        RECT 15.05 5.43 17.8 7.035 ;
        RECT 17.035 10.045 17.21 10.595 ;
        RECT 17.035 7.305 17.21 8.445 ;
        RECT 17.035 5.43 17.205 10.595 ;
        RECT 15.22 5.43 15.39 7.765 ;
      LAYER met1 ;
        RECT 0.005 5.43 99.425 7.03 ;
        RECT 94.545 5.425 98.28 7.035 ;
        RECT 83.84 5.4 93.5 7.03 ;
        RECT 88.93 5.4 91.68 7.035 ;
        RECT 78.22 5.425 81.955 7.035 ;
        RECT 67.515 5.4 77.175 7.03 ;
        RECT 72.605 5.4 75.355 7.035 ;
        RECT 61.895 5.425 65.63 7.035 ;
        RECT 51.19 5.4 60.85 7.03 ;
        RECT 56.28 5.4 59.03 7.035 ;
        RECT 45.57 5.425 49.305 7.035 ;
        RECT 34.865 5.4 44.525 7.03 ;
        RECT 39.955 5.4 42.705 7.035 ;
        RECT 29.245 5.425 32.98 7.035 ;
        RECT 18.54 5.4 28.2 7.03 ;
        RECT 23.63 5.4 26.38 7.035 ;
        RECT 15.05 5.43 17.8 7.035 ;
        RECT 16.975 8.945 17.265 9.175 ;
        RECT 16.805 8.975 17.265 9.145 ;
      LAYER mcon ;
        RECT 17.035 8.975 17.205 9.145 ;
        RECT 17.34 6.835 17.51 7.005 ;
        RECT 18.685 5.43 18.855 5.6 ;
        RECT 19.145 5.43 19.315 5.6 ;
        RECT 19.605 5.43 19.775 5.6 ;
        RECT 20.065 5.43 20.235 5.6 ;
        RECT 20.525 5.43 20.695 5.6 ;
        RECT 20.985 5.43 21.155 5.6 ;
        RECT 21.445 5.43 21.615 5.6 ;
        RECT 21.905 5.43 22.075 5.6 ;
        RECT 22.365 5.43 22.535 5.6 ;
        RECT 22.825 5.43 22.995 5.6 ;
        RECT 23.285 5.43 23.455 5.6 ;
        RECT 23.745 5.43 23.915 5.6 ;
        RECT 24.205 5.43 24.375 5.6 ;
        RECT 24.665 5.43 24.835 5.6 ;
        RECT 25.125 5.43 25.295 5.6 ;
        RECT 25.585 5.43 25.755 5.6 ;
        RECT 25.92 6.835 26.09 7.005 ;
        RECT 26.045 5.43 26.215 5.6 ;
        RECT 26.505 5.43 26.675 5.6 ;
        RECT 26.965 5.43 27.135 5.6 ;
        RECT 27.425 5.43 27.595 5.6 ;
        RECT 27.885 5.43 28.055 5.6 ;
        RECT 31.535 6.835 31.705 7.005 ;
        RECT 31.535 5.455 31.705 5.625 ;
        RECT 32.24 6.835 32.41 7.005 ;
        RECT 32.24 5.455 32.41 5.625 ;
        RECT 33.23 5.46 33.4 5.63 ;
        RECT 33.235 6.83 33.405 7 ;
        RECT 35.01 5.43 35.18 5.6 ;
        RECT 35.47 5.43 35.64 5.6 ;
        RECT 35.93 5.43 36.1 5.6 ;
        RECT 36.39 5.43 36.56 5.6 ;
        RECT 36.85 5.43 37.02 5.6 ;
        RECT 37.31 5.43 37.48 5.6 ;
        RECT 37.77 5.43 37.94 5.6 ;
        RECT 38.23 5.43 38.4 5.6 ;
        RECT 38.69 5.43 38.86 5.6 ;
        RECT 39.15 5.43 39.32 5.6 ;
        RECT 39.61 5.43 39.78 5.6 ;
        RECT 40.07 5.43 40.24 5.6 ;
        RECT 40.53 5.43 40.7 5.6 ;
        RECT 40.99 5.43 41.16 5.6 ;
        RECT 41.45 5.43 41.62 5.6 ;
        RECT 41.91 5.43 42.08 5.6 ;
        RECT 42.245 6.835 42.415 7.005 ;
        RECT 42.37 5.43 42.54 5.6 ;
        RECT 42.83 5.43 43 5.6 ;
        RECT 43.29 5.43 43.46 5.6 ;
        RECT 43.75 5.43 43.92 5.6 ;
        RECT 44.21 5.43 44.38 5.6 ;
        RECT 47.86 6.835 48.03 7.005 ;
        RECT 47.86 5.455 48.03 5.625 ;
        RECT 48.565 6.835 48.735 7.005 ;
        RECT 48.565 5.455 48.735 5.625 ;
        RECT 49.555 5.46 49.725 5.63 ;
        RECT 49.56 6.83 49.73 7 ;
        RECT 51.335 5.43 51.505 5.6 ;
        RECT 51.795 5.43 51.965 5.6 ;
        RECT 52.255 5.43 52.425 5.6 ;
        RECT 52.715 5.43 52.885 5.6 ;
        RECT 53.175 5.43 53.345 5.6 ;
        RECT 53.635 5.43 53.805 5.6 ;
        RECT 54.095 5.43 54.265 5.6 ;
        RECT 54.555 5.43 54.725 5.6 ;
        RECT 55.015 5.43 55.185 5.6 ;
        RECT 55.475 5.43 55.645 5.6 ;
        RECT 55.935 5.43 56.105 5.6 ;
        RECT 56.395 5.43 56.565 5.6 ;
        RECT 56.855 5.43 57.025 5.6 ;
        RECT 57.315 5.43 57.485 5.6 ;
        RECT 57.775 5.43 57.945 5.6 ;
        RECT 58.235 5.43 58.405 5.6 ;
        RECT 58.57 6.835 58.74 7.005 ;
        RECT 58.695 5.43 58.865 5.6 ;
        RECT 59.155 5.43 59.325 5.6 ;
        RECT 59.615 5.43 59.785 5.6 ;
        RECT 60.075 5.43 60.245 5.6 ;
        RECT 60.535 5.43 60.705 5.6 ;
        RECT 64.185 6.835 64.355 7.005 ;
        RECT 64.185 5.455 64.355 5.625 ;
        RECT 64.89 6.835 65.06 7.005 ;
        RECT 64.89 5.455 65.06 5.625 ;
        RECT 65.88 5.46 66.05 5.63 ;
        RECT 65.885 6.83 66.055 7 ;
        RECT 67.66 5.43 67.83 5.6 ;
        RECT 68.12 5.43 68.29 5.6 ;
        RECT 68.58 5.43 68.75 5.6 ;
        RECT 69.04 5.43 69.21 5.6 ;
        RECT 69.5 5.43 69.67 5.6 ;
        RECT 69.96 5.43 70.13 5.6 ;
        RECT 70.42 5.43 70.59 5.6 ;
        RECT 70.88 5.43 71.05 5.6 ;
        RECT 71.34 5.43 71.51 5.6 ;
        RECT 71.8 5.43 71.97 5.6 ;
        RECT 72.26 5.43 72.43 5.6 ;
        RECT 72.72 5.43 72.89 5.6 ;
        RECT 73.18 5.43 73.35 5.6 ;
        RECT 73.64 5.43 73.81 5.6 ;
        RECT 74.1 5.43 74.27 5.6 ;
        RECT 74.56 5.43 74.73 5.6 ;
        RECT 74.895 6.835 75.065 7.005 ;
        RECT 75.02 5.43 75.19 5.6 ;
        RECT 75.48 5.43 75.65 5.6 ;
        RECT 75.94 5.43 76.11 5.6 ;
        RECT 76.4 5.43 76.57 5.6 ;
        RECT 76.86 5.43 77.03 5.6 ;
        RECT 80.51 6.835 80.68 7.005 ;
        RECT 80.51 5.455 80.68 5.625 ;
        RECT 81.215 6.835 81.385 7.005 ;
        RECT 81.215 5.455 81.385 5.625 ;
        RECT 82.205 5.46 82.375 5.63 ;
        RECT 82.21 6.83 82.38 7 ;
        RECT 83.985 5.43 84.155 5.6 ;
        RECT 84.445 5.43 84.615 5.6 ;
        RECT 84.905 5.43 85.075 5.6 ;
        RECT 85.365 5.43 85.535 5.6 ;
        RECT 85.825 5.43 85.995 5.6 ;
        RECT 86.285 5.43 86.455 5.6 ;
        RECT 86.745 5.43 86.915 5.6 ;
        RECT 87.205 5.43 87.375 5.6 ;
        RECT 87.665 5.43 87.835 5.6 ;
        RECT 88.125 5.43 88.295 5.6 ;
        RECT 88.585 5.43 88.755 5.6 ;
        RECT 89.045 5.43 89.215 5.6 ;
        RECT 89.505 5.43 89.675 5.6 ;
        RECT 89.965 5.43 90.135 5.6 ;
        RECT 90.425 5.43 90.595 5.6 ;
        RECT 90.885 5.43 91.055 5.6 ;
        RECT 91.22 6.835 91.39 7.005 ;
        RECT 91.345 5.43 91.515 5.6 ;
        RECT 91.805 5.43 91.975 5.6 ;
        RECT 92.265 5.43 92.435 5.6 ;
        RECT 92.725 5.43 92.895 5.6 ;
        RECT 93.185 5.43 93.355 5.6 ;
        RECT 96.835 6.835 97.005 7.005 ;
        RECT 96.835 5.455 97.005 5.625 ;
        RECT 97.54 6.835 97.71 7.005 ;
        RECT 97.54 5.455 97.71 5.625 ;
        RECT 98.53 5.46 98.7 5.63 ;
        RECT 98.535 6.83 98.705 7 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 92.73 4.27 93.06 5 ;
        RECT 76.405 4.27 76.735 5 ;
        RECT 60.08 4.27 60.41 5 ;
        RECT 43.755 4.27 44.085 5 ;
        RECT 27.43 4.27 27.76 5 ;
      LAYER met2 ;
        RECT 92.755 4.25 93.035 4.62 ;
        RECT 92.765 3.995 93.025 4.62 ;
        RECT 76.43 4.25 76.71 4.62 ;
        RECT 76.44 3.995 76.7 4.62 ;
        RECT 60.105 4.25 60.385 4.62 ;
        RECT 60.115 3.995 60.375 4.62 ;
        RECT 43.78 4.25 44.06 4.62 ;
        RECT 43.79 3.995 44.05 4.62 ;
        RECT 27.455 4.25 27.735 4.62 ;
        RECT 27.465 3.995 27.725 4.62 ;
      LAYER li1 ;
        RECT 0.05 10.86 99.43 12.46 ;
        RECT 98.455 10.23 98.625 12.46 ;
        RECT 97.46 10.235 97.63 12.46 ;
        RECT 94.715 10.235 94.885 12.46 ;
        RECT 89.1 10.235 89.27 12.46 ;
        RECT 82.13 10.23 82.3 12.46 ;
        RECT 81.135 10.235 81.305 12.46 ;
        RECT 78.39 10.235 78.56 12.46 ;
        RECT 72.775 10.235 72.945 12.46 ;
        RECT 65.805 10.23 65.975 12.46 ;
        RECT 64.81 10.235 64.98 12.46 ;
        RECT 62.065 10.235 62.235 12.46 ;
        RECT 56.45 10.235 56.62 12.46 ;
        RECT 49.48 10.23 49.65 12.46 ;
        RECT 48.485 10.235 48.655 12.46 ;
        RECT 45.74 10.235 45.91 12.46 ;
        RECT 40.125 10.235 40.295 12.46 ;
        RECT 33.155 10.23 33.325 12.46 ;
        RECT 32.16 10.235 32.33 12.46 ;
        RECT 29.415 10.235 29.585 12.46 ;
        RECT 23.8 10.235 23.97 12.46 ;
        RECT 15.22 10.235 15.39 12.46 ;
        RECT 0 0 99.425 1.6 ;
        RECT 98.45 0 98.62 2.23 ;
        RECT 97.46 0 97.63 2.225 ;
        RECT 94.715 0 94.885 2.225 ;
        RECT 83.84 0 93.655 2.88 ;
        RECT 91.97 0 92.14 3.38 ;
        RECT 90.01 0 90.18 3.38 ;
        RECT 89.94 0 90.18 2.89 ;
        RECT 88.39 0 88.585 2.89 ;
        RECT 87.57 0 87.74 3.38 ;
        RECT 86.61 0 86.78 3.38 ;
        RECT 86.09 0 86.78 2.89 ;
        RECT 86.09 0 86.26 3.38 ;
        RECT 85.13 0 85.3 3.38 ;
        RECT 84.17 0 84.34 3.38 ;
        RECT 83.965 0 84.34 2.89 ;
        RECT 82.125 0 82.295 2.23 ;
        RECT 81.135 0 81.305 2.225 ;
        RECT 78.39 0 78.56 2.225 ;
        RECT 67.515 0 77.33 2.88 ;
        RECT 75.645 0 75.815 3.38 ;
        RECT 73.685 0 73.855 3.38 ;
        RECT 73.615 0 73.855 2.89 ;
        RECT 72.065 0 72.26 2.89 ;
        RECT 71.245 0 71.415 3.38 ;
        RECT 70.285 0 70.455 3.38 ;
        RECT 69.765 0 70.455 2.89 ;
        RECT 69.765 0 69.935 3.38 ;
        RECT 68.805 0 68.975 3.38 ;
        RECT 67.845 0 68.015 3.38 ;
        RECT 67.64 0 68.015 2.89 ;
        RECT 65.8 0 65.97 2.23 ;
        RECT 64.81 0 64.98 2.225 ;
        RECT 62.065 0 62.235 2.225 ;
        RECT 51.19 0 61.005 2.88 ;
        RECT 59.32 0 59.49 3.38 ;
        RECT 57.36 0 57.53 3.38 ;
        RECT 57.29 0 57.53 2.89 ;
        RECT 55.74 0 55.935 2.89 ;
        RECT 54.92 0 55.09 3.38 ;
        RECT 53.96 0 54.13 3.38 ;
        RECT 53.44 0 54.13 2.89 ;
        RECT 53.44 0 53.61 3.38 ;
        RECT 52.48 0 52.65 3.38 ;
        RECT 51.52 0 51.69 3.38 ;
        RECT 51.315 0 51.69 2.89 ;
        RECT 49.475 0 49.645 2.23 ;
        RECT 48.485 0 48.655 2.225 ;
        RECT 45.74 0 45.91 2.225 ;
        RECT 34.865 0 44.68 2.88 ;
        RECT 42.995 0 43.165 3.38 ;
        RECT 41.035 0 41.205 3.38 ;
        RECT 40.965 0 41.205 2.89 ;
        RECT 39.415 0 39.61 2.89 ;
        RECT 38.595 0 38.765 3.38 ;
        RECT 37.635 0 37.805 3.38 ;
        RECT 37.115 0 37.805 2.89 ;
        RECT 37.115 0 37.285 3.38 ;
        RECT 36.155 0 36.325 3.38 ;
        RECT 35.195 0 35.365 3.38 ;
        RECT 34.99 0 35.365 2.89 ;
        RECT 33.15 0 33.32 2.23 ;
        RECT 32.16 0 32.33 2.225 ;
        RECT 29.415 0 29.585 2.225 ;
        RECT 18.54 0 28.355 2.88 ;
        RECT 26.67 0 26.84 3.38 ;
        RECT 24.71 0 24.88 3.38 ;
        RECT 24.64 0 24.88 2.89 ;
        RECT 23.09 0 23.285 2.89 ;
        RECT 22.27 0 22.44 3.38 ;
        RECT 21.31 0 21.48 3.38 ;
        RECT 20.79 0 21.48 2.89 ;
        RECT 20.79 0 20.96 3.38 ;
        RECT 19.83 0 20 3.38 ;
        RECT 18.87 0 19.04 3.38 ;
        RECT 18.665 0 19.04 2.89 ;
        RECT 92.93 3.87 93.1 4.24 ;
        RECT 92.61 3.87 93.1 4.04 ;
        RECT 90.97 3.87 91.14 4.24 ;
        RECT 90.65 3.87 91.14 4.04 ;
        RECT 90.115 8.365 90.285 10.315 ;
        RECT 90.055 10.145 90.225 10.595 ;
        RECT 90.055 7.305 90.225 8.535 ;
        RECT 76.605 3.87 76.775 4.24 ;
        RECT 76.285 3.87 76.775 4.04 ;
        RECT 74.645 3.87 74.815 4.24 ;
        RECT 74.325 3.87 74.815 4.04 ;
        RECT 73.79 8.365 73.96 10.315 ;
        RECT 73.73 10.145 73.9 10.595 ;
        RECT 73.73 7.305 73.9 8.535 ;
        RECT 60.28 3.87 60.45 4.24 ;
        RECT 59.96 3.87 60.45 4.04 ;
        RECT 58.32 3.87 58.49 4.24 ;
        RECT 58 3.87 58.49 4.04 ;
        RECT 57.465 8.365 57.635 10.315 ;
        RECT 57.405 10.145 57.575 10.595 ;
        RECT 57.405 7.305 57.575 8.535 ;
        RECT 43.955 3.87 44.125 4.24 ;
        RECT 43.635 3.87 44.125 4.04 ;
        RECT 41.995 3.87 42.165 4.24 ;
        RECT 41.675 3.87 42.165 4.04 ;
        RECT 41.14 8.365 41.31 10.315 ;
        RECT 41.08 10.145 41.25 10.595 ;
        RECT 41.08 7.305 41.25 8.535 ;
        RECT 27.63 3.87 27.8 4.24 ;
        RECT 27.31 3.87 27.8 4.04 ;
        RECT 25.67 3.87 25.84 4.24 ;
        RECT 25.35 3.87 25.84 4.04 ;
        RECT 24.815 8.365 24.985 10.315 ;
        RECT 24.755 10.145 24.925 10.595 ;
        RECT 24.755 7.305 24.925 8.535 ;
      LAYER met1 ;
        RECT 0.05 10.86 99.43 12.46 ;
        RECT 90.055 8.575 90.345 8.805 ;
        RECT 89.675 8.6 90.345 8.775 ;
        RECT 89.675 8.6 89.85 12.46 ;
        RECT 73.73 8.575 74.02 8.805 ;
        RECT 73.35 8.6 74.02 8.775 ;
        RECT 73.35 8.6 73.525 12.46 ;
        RECT 57.405 8.575 57.695 8.805 ;
        RECT 57.025 8.6 57.695 8.775 ;
        RECT 57.025 8.6 57.2 12.46 ;
        RECT 41.08 8.575 41.37 8.805 ;
        RECT 40.7 8.6 41.37 8.775 ;
        RECT 40.7 8.6 40.875 12.46 ;
        RECT 24.755 8.575 25.045 8.805 ;
        RECT 24.375 8.6 25.045 8.775 ;
        RECT 24.375 8.6 24.55 12.46 ;
        RECT 0 0 99.425 1.6 ;
        RECT 93.47 0 93.655 4.24 ;
        RECT 92.705 4.085 93.655 4.24 ;
        RECT 92.735 4.055 93.655 4.24 ;
        RECT 83.84 0 93.655 2.91 ;
        RECT 92.735 4.04 93.16 4.27 ;
        RECT 92.735 4.025 93.055 4.285 ;
        RECT 91.245 4.225 93.01 4.35 ;
        RECT 91.245 4.225 92.845 4.365 ;
        RECT 90.91 4.085 91.385 4.27 ;
        RECT 90.91 4.04 91.2 4.27 ;
        RECT 77.145 0 77.33 4.24 ;
        RECT 76.38 4.085 77.33 4.24 ;
        RECT 76.41 4.055 77.33 4.24 ;
        RECT 67.515 0 77.33 2.91 ;
        RECT 76.41 4.04 76.835 4.27 ;
        RECT 76.41 4.025 76.73 4.285 ;
        RECT 74.92 4.225 76.685 4.35 ;
        RECT 74.92 4.225 76.52 4.365 ;
        RECT 74.585 4.085 75.06 4.27 ;
        RECT 74.585 4.04 74.875 4.27 ;
        RECT 60.82 0 61.005 4.24 ;
        RECT 60.055 4.085 61.005 4.24 ;
        RECT 60.085 4.055 61.005 4.24 ;
        RECT 51.19 0 61.005 2.91 ;
        RECT 60.085 4.04 60.51 4.27 ;
        RECT 60.085 4.025 60.405 4.285 ;
        RECT 58.595 4.225 60.36 4.35 ;
        RECT 58.595 4.225 60.195 4.365 ;
        RECT 58.26 4.085 58.735 4.27 ;
        RECT 58.26 4.04 58.55 4.27 ;
        RECT 44.495 0 44.68 4.24 ;
        RECT 43.73 4.085 44.68 4.24 ;
        RECT 43.76 4.055 44.68 4.24 ;
        RECT 34.865 0 44.68 2.91 ;
        RECT 43.76 4.04 44.185 4.27 ;
        RECT 43.76 4.025 44.08 4.285 ;
        RECT 42.27 4.225 44.035 4.35 ;
        RECT 42.27 4.225 43.87 4.365 ;
        RECT 41.935 4.085 42.41 4.27 ;
        RECT 41.935 4.04 42.225 4.27 ;
        RECT 28.17 0 28.355 4.24 ;
        RECT 27.405 4.085 28.355 4.24 ;
        RECT 27.435 4.055 28.355 4.24 ;
        RECT 18.54 0 28.355 2.91 ;
        RECT 27.435 4.04 27.86 4.27 ;
        RECT 27.435 4.025 27.755 4.285 ;
        RECT 25.945 4.225 27.71 4.35 ;
        RECT 25.945 4.225 27.545 4.365 ;
        RECT 25.61 4.085 26.085 4.27 ;
        RECT 25.61 4.04 25.9 4.27 ;
      LAYER via1 ;
        RECT 27.52 4.08 27.67 4.23 ;
        RECT 43.845 4.08 43.995 4.23 ;
        RECT 60.17 4.08 60.32 4.23 ;
        RECT 76.495 4.08 76.645 4.23 ;
        RECT 92.82 4.08 92.97 4.23 ;
      LAYER via2 ;
        RECT 27.495 4.335 27.695 4.535 ;
        RECT 43.82 4.335 44.02 4.535 ;
        RECT 60.145 4.335 60.345 4.535 ;
        RECT 76.47 4.335 76.67 4.535 ;
        RECT 92.795 4.335 92.995 4.535 ;
      LAYER mcon ;
        RECT 15.3 10.895 15.47 11.065 ;
        RECT 15.98 10.895 16.15 11.065 ;
        RECT 16.66 10.895 16.83 11.065 ;
        RECT 17.34 10.895 17.51 11.065 ;
        RECT 18.685 2.71 18.855 2.88 ;
        RECT 19.145 2.71 19.315 2.88 ;
        RECT 19.605 2.71 19.775 2.88 ;
        RECT 20.065 2.71 20.235 2.88 ;
        RECT 20.525 2.71 20.695 2.88 ;
        RECT 20.985 2.71 21.155 2.88 ;
        RECT 21.445 2.71 21.615 2.88 ;
        RECT 21.905 2.71 22.075 2.88 ;
        RECT 22.365 2.71 22.535 2.88 ;
        RECT 22.825 2.71 22.995 2.88 ;
        RECT 23.285 2.71 23.455 2.88 ;
        RECT 23.745 2.71 23.915 2.88 ;
        RECT 23.88 10.895 24.05 11.065 ;
        RECT 24.205 2.71 24.375 2.88 ;
        RECT 24.56 10.895 24.73 11.065 ;
        RECT 24.665 2.71 24.835 2.88 ;
        RECT 24.815 8.605 24.985 8.775 ;
        RECT 25.125 2.71 25.295 2.88 ;
        RECT 25.24 10.895 25.41 11.065 ;
        RECT 25.585 2.71 25.755 2.88 ;
        RECT 25.67 4.07 25.84 4.24 ;
        RECT 25.92 10.895 26.09 11.065 ;
        RECT 26.045 2.71 26.215 2.88 ;
        RECT 26.505 2.71 26.675 2.88 ;
        RECT 26.965 2.71 27.135 2.88 ;
        RECT 27.425 2.71 27.595 2.88 ;
        RECT 27.63 4.07 27.8 4.24 ;
        RECT 27.885 2.71 28.055 2.88 ;
        RECT 29.495 10.895 29.665 11.065 ;
        RECT 29.495 1.395 29.665 1.565 ;
        RECT 30.175 10.895 30.345 11.065 ;
        RECT 30.175 1.395 30.345 1.565 ;
        RECT 30.855 10.895 31.025 11.065 ;
        RECT 30.855 1.395 31.025 1.565 ;
        RECT 31.535 10.895 31.705 11.065 ;
        RECT 31.535 1.395 31.705 1.565 ;
        RECT 32.24 10.895 32.41 11.065 ;
        RECT 32.24 1.395 32.41 1.565 ;
        RECT 33.23 1.4 33.4 1.57 ;
        RECT 33.235 10.89 33.405 11.06 ;
        RECT 35.01 2.71 35.18 2.88 ;
        RECT 35.47 2.71 35.64 2.88 ;
        RECT 35.93 2.71 36.1 2.88 ;
        RECT 36.39 2.71 36.56 2.88 ;
        RECT 36.85 2.71 37.02 2.88 ;
        RECT 37.31 2.71 37.48 2.88 ;
        RECT 37.77 2.71 37.94 2.88 ;
        RECT 38.23 2.71 38.4 2.88 ;
        RECT 38.69 2.71 38.86 2.88 ;
        RECT 39.15 2.71 39.32 2.88 ;
        RECT 39.61 2.71 39.78 2.88 ;
        RECT 40.07 2.71 40.24 2.88 ;
        RECT 40.205 10.895 40.375 11.065 ;
        RECT 40.53 2.71 40.7 2.88 ;
        RECT 40.885 10.895 41.055 11.065 ;
        RECT 40.99 2.71 41.16 2.88 ;
        RECT 41.14 8.605 41.31 8.775 ;
        RECT 41.45 2.71 41.62 2.88 ;
        RECT 41.565 10.895 41.735 11.065 ;
        RECT 41.91 2.71 42.08 2.88 ;
        RECT 41.995 4.07 42.165 4.24 ;
        RECT 42.245 10.895 42.415 11.065 ;
        RECT 42.37 2.71 42.54 2.88 ;
        RECT 42.83 2.71 43 2.88 ;
        RECT 43.29 2.71 43.46 2.88 ;
        RECT 43.75 2.71 43.92 2.88 ;
        RECT 43.955 4.07 44.125 4.24 ;
        RECT 44.21 2.71 44.38 2.88 ;
        RECT 45.82 10.895 45.99 11.065 ;
        RECT 45.82 1.395 45.99 1.565 ;
        RECT 46.5 10.895 46.67 11.065 ;
        RECT 46.5 1.395 46.67 1.565 ;
        RECT 47.18 10.895 47.35 11.065 ;
        RECT 47.18 1.395 47.35 1.565 ;
        RECT 47.86 10.895 48.03 11.065 ;
        RECT 47.86 1.395 48.03 1.565 ;
        RECT 48.565 10.895 48.735 11.065 ;
        RECT 48.565 1.395 48.735 1.565 ;
        RECT 49.555 1.4 49.725 1.57 ;
        RECT 49.56 10.89 49.73 11.06 ;
        RECT 51.335 2.71 51.505 2.88 ;
        RECT 51.795 2.71 51.965 2.88 ;
        RECT 52.255 2.71 52.425 2.88 ;
        RECT 52.715 2.71 52.885 2.88 ;
        RECT 53.175 2.71 53.345 2.88 ;
        RECT 53.635 2.71 53.805 2.88 ;
        RECT 54.095 2.71 54.265 2.88 ;
        RECT 54.555 2.71 54.725 2.88 ;
        RECT 55.015 2.71 55.185 2.88 ;
        RECT 55.475 2.71 55.645 2.88 ;
        RECT 55.935 2.71 56.105 2.88 ;
        RECT 56.395 2.71 56.565 2.88 ;
        RECT 56.53 10.895 56.7 11.065 ;
        RECT 56.855 2.71 57.025 2.88 ;
        RECT 57.21 10.895 57.38 11.065 ;
        RECT 57.315 2.71 57.485 2.88 ;
        RECT 57.465 8.605 57.635 8.775 ;
        RECT 57.775 2.71 57.945 2.88 ;
        RECT 57.89 10.895 58.06 11.065 ;
        RECT 58.235 2.71 58.405 2.88 ;
        RECT 58.32 4.07 58.49 4.24 ;
        RECT 58.57 10.895 58.74 11.065 ;
        RECT 58.695 2.71 58.865 2.88 ;
        RECT 59.155 2.71 59.325 2.88 ;
        RECT 59.615 2.71 59.785 2.88 ;
        RECT 60.075 2.71 60.245 2.88 ;
        RECT 60.28 4.07 60.45 4.24 ;
        RECT 60.535 2.71 60.705 2.88 ;
        RECT 62.145 10.895 62.315 11.065 ;
        RECT 62.145 1.395 62.315 1.565 ;
        RECT 62.825 10.895 62.995 11.065 ;
        RECT 62.825 1.395 62.995 1.565 ;
        RECT 63.505 10.895 63.675 11.065 ;
        RECT 63.505 1.395 63.675 1.565 ;
        RECT 64.185 10.895 64.355 11.065 ;
        RECT 64.185 1.395 64.355 1.565 ;
        RECT 64.89 10.895 65.06 11.065 ;
        RECT 64.89 1.395 65.06 1.565 ;
        RECT 65.88 1.4 66.05 1.57 ;
        RECT 65.885 10.89 66.055 11.06 ;
        RECT 67.66 2.71 67.83 2.88 ;
        RECT 68.12 2.71 68.29 2.88 ;
        RECT 68.58 2.71 68.75 2.88 ;
        RECT 69.04 2.71 69.21 2.88 ;
        RECT 69.5 2.71 69.67 2.88 ;
        RECT 69.96 2.71 70.13 2.88 ;
        RECT 70.42 2.71 70.59 2.88 ;
        RECT 70.88 2.71 71.05 2.88 ;
        RECT 71.34 2.71 71.51 2.88 ;
        RECT 71.8 2.71 71.97 2.88 ;
        RECT 72.26 2.71 72.43 2.88 ;
        RECT 72.72 2.71 72.89 2.88 ;
        RECT 72.855 10.895 73.025 11.065 ;
        RECT 73.18 2.71 73.35 2.88 ;
        RECT 73.535 10.895 73.705 11.065 ;
        RECT 73.64 2.71 73.81 2.88 ;
        RECT 73.79 8.605 73.96 8.775 ;
        RECT 74.1 2.71 74.27 2.88 ;
        RECT 74.215 10.895 74.385 11.065 ;
        RECT 74.56 2.71 74.73 2.88 ;
        RECT 74.645 4.07 74.815 4.24 ;
        RECT 74.895 10.895 75.065 11.065 ;
        RECT 75.02 2.71 75.19 2.88 ;
        RECT 75.48 2.71 75.65 2.88 ;
        RECT 75.94 2.71 76.11 2.88 ;
        RECT 76.4 2.71 76.57 2.88 ;
        RECT 76.605 4.07 76.775 4.24 ;
        RECT 76.86 2.71 77.03 2.88 ;
        RECT 78.47 10.895 78.64 11.065 ;
        RECT 78.47 1.395 78.64 1.565 ;
        RECT 79.15 10.895 79.32 11.065 ;
        RECT 79.15 1.395 79.32 1.565 ;
        RECT 79.83 10.895 80 11.065 ;
        RECT 79.83 1.395 80 1.565 ;
        RECT 80.51 10.895 80.68 11.065 ;
        RECT 80.51 1.395 80.68 1.565 ;
        RECT 81.215 10.895 81.385 11.065 ;
        RECT 81.215 1.395 81.385 1.565 ;
        RECT 82.205 1.4 82.375 1.57 ;
        RECT 82.21 10.89 82.38 11.06 ;
        RECT 83.985 2.71 84.155 2.88 ;
        RECT 84.445 2.71 84.615 2.88 ;
        RECT 84.905 2.71 85.075 2.88 ;
        RECT 85.365 2.71 85.535 2.88 ;
        RECT 85.825 2.71 85.995 2.88 ;
        RECT 86.285 2.71 86.455 2.88 ;
        RECT 86.745 2.71 86.915 2.88 ;
        RECT 87.205 2.71 87.375 2.88 ;
        RECT 87.665 2.71 87.835 2.88 ;
        RECT 88.125 2.71 88.295 2.88 ;
        RECT 88.585 2.71 88.755 2.88 ;
        RECT 89.045 2.71 89.215 2.88 ;
        RECT 89.18 10.895 89.35 11.065 ;
        RECT 89.505 2.71 89.675 2.88 ;
        RECT 89.86 10.895 90.03 11.065 ;
        RECT 89.965 2.71 90.135 2.88 ;
        RECT 90.115 8.605 90.285 8.775 ;
        RECT 90.425 2.71 90.595 2.88 ;
        RECT 90.54 10.895 90.71 11.065 ;
        RECT 90.885 2.71 91.055 2.88 ;
        RECT 90.97 4.07 91.14 4.24 ;
        RECT 91.22 10.895 91.39 11.065 ;
        RECT 91.345 2.71 91.515 2.88 ;
        RECT 91.805 2.71 91.975 2.88 ;
        RECT 92.265 2.71 92.435 2.88 ;
        RECT 92.725 2.71 92.895 2.88 ;
        RECT 92.93 4.07 93.1 4.24 ;
        RECT 93.185 2.71 93.355 2.88 ;
        RECT 94.795 10.895 94.965 11.065 ;
        RECT 94.795 1.395 94.965 1.565 ;
        RECT 95.475 10.895 95.645 11.065 ;
        RECT 95.475 1.395 95.645 1.565 ;
        RECT 96.155 10.895 96.325 11.065 ;
        RECT 96.155 1.395 96.325 1.565 ;
        RECT 96.835 10.895 97.005 11.065 ;
        RECT 96.835 1.395 97.005 1.565 ;
        RECT 97.54 10.895 97.71 11.065 ;
        RECT 97.54 1.395 97.71 1.565 ;
        RECT 98.53 1.4 98.7 1.57 ;
        RECT 98.535 10.89 98.705 11.06 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 90.405 9.34 90.775 9.71 ;
      RECT 90.405 9.375 92.39 9.675 ;
      RECT 92.09 3.575 92.39 9.675 ;
      RECT 89.09 3.31 89.42 4.04 ;
      RECT 88.21 3.31 88.54 4.04 ;
      RECT 91.29 3.575 92.58 3.875 ;
      RECT 92.25 3.145 92.58 3.875 ;
      RECT 88.21 3.575 90.35 3.875 ;
      RECT 90.05 3.26 90.35 3.875 ;
      RECT 91.29 3.275 91.595 3.875 ;
      RECT 90.05 3.26 91.41 3.57 ;
      RECT 88.71 4.83 89.04 5.16 ;
      RECT 87.505 4.845 89.04 5.145 ;
      RECT 87.505 3.725 87.805 5.145 ;
      RECT 87.25 3.71 87.58 4.04 ;
      RECT 74.08 9.34 74.45 9.71 ;
      RECT 74.08 9.375 76.065 9.675 ;
      RECT 75.765 3.575 76.065 9.675 ;
      RECT 72.765 3.31 73.095 4.04 ;
      RECT 71.885 3.31 72.215 4.04 ;
      RECT 74.965 3.575 76.255 3.875 ;
      RECT 75.925 3.145 76.255 3.875 ;
      RECT 71.885 3.575 74.025 3.875 ;
      RECT 73.725 3.26 74.025 3.875 ;
      RECT 74.965 3.275 75.27 3.875 ;
      RECT 73.725 3.26 75.085 3.57 ;
      RECT 72.385 4.83 72.715 5.16 ;
      RECT 71.18 4.845 72.715 5.145 ;
      RECT 71.18 3.725 71.48 5.145 ;
      RECT 70.925 3.71 71.255 4.04 ;
      RECT 57.755 9.34 58.125 9.71 ;
      RECT 57.755 9.375 59.74 9.675 ;
      RECT 59.44 3.575 59.74 9.675 ;
      RECT 56.44 3.31 56.77 4.04 ;
      RECT 55.56 3.31 55.89 4.04 ;
      RECT 58.64 3.575 59.93 3.875 ;
      RECT 59.6 3.145 59.93 3.875 ;
      RECT 55.56 3.575 57.7 3.875 ;
      RECT 57.4 3.26 57.7 3.875 ;
      RECT 58.64 3.275 58.945 3.875 ;
      RECT 57.4 3.26 58.76 3.57 ;
      RECT 56.06 4.83 56.39 5.16 ;
      RECT 54.855 4.845 56.39 5.145 ;
      RECT 54.855 3.725 55.155 5.145 ;
      RECT 54.6 3.71 54.93 4.04 ;
      RECT 41.43 9.34 41.8 9.71 ;
      RECT 41.43 9.375 43.415 9.675 ;
      RECT 43.115 3.575 43.415 9.675 ;
      RECT 40.115 3.31 40.445 4.04 ;
      RECT 39.235 3.31 39.565 4.04 ;
      RECT 42.315 3.575 43.605 3.875 ;
      RECT 43.275 3.145 43.605 3.875 ;
      RECT 39.235 3.575 41.375 3.875 ;
      RECT 41.075 3.26 41.375 3.875 ;
      RECT 42.315 3.275 42.62 3.875 ;
      RECT 41.075 3.26 42.435 3.57 ;
      RECT 39.735 4.83 40.065 5.16 ;
      RECT 38.53 4.845 40.065 5.145 ;
      RECT 38.53 3.725 38.83 5.145 ;
      RECT 38.275 3.71 38.605 4.04 ;
      RECT 25.105 9.34 25.475 9.71 ;
      RECT 25.105 9.375 27.09 9.675 ;
      RECT 26.79 3.575 27.09 9.675 ;
      RECT 23.79 3.31 24.12 4.04 ;
      RECT 22.91 3.31 23.24 4.04 ;
      RECT 25.99 3.575 27.28 3.875 ;
      RECT 26.95 3.145 27.28 3.875 ;
      RECT 22.91 3.575 25.05 3.875 ;
      RECT 24.75 3.26 25.05 3.875 ;
      RECT 25.99 3.275 26.295 3.875 ;
      RECT 24.75 3.26 26.11 3.57 ;
      RECT 23.41 4.83 23.74 5.16 ;
      RECT 22.205 4.845 23.74 5.145 ;
      RECT 22.205 3.725 22.505 5.145 ;
      RECT 21.95 3.71 22.28 4.04 ;
      RECT 98.785 7.195 99.165 12.46 ;
      RECT 90.65 3.87 90.98 4.6 ;
      RECT 86.53 3.71 86.86 4.44 ;
      RECT 85.53 3.15 85.86 3.88 ;
      RECT 84.09 3.87 84.42 4.6 ;
      RECT 82.46 7.195 82.84 12.46 ;
      RECT 74.325 3.87 74.655 4.6 ;
      RECT 70.205 3.71 70.535 4.44 ;
      RECT 69.205 3.15 69.535 3.88 ;
      RECT 67.765 3.87 68.095 4.6 ;
      RECT 66.135 7.195 66.515 12.46 ;
      RECT 58 3.87 58.33 4.6 ;
      RECT 53.88 3.71 54.21 4.44 ;
      RECT 52.88 3.15 53.21 3.88 ;
      RECT 51.44 3.87 51.77 4.6 ;
      RECT 49.81 7.195 50.19 12.46 ;
      RECT 41.675 3.87 42.005 4.6 ;
      RECT 37.555 3.71 37.885 4.44 ;
      RECT 36.555 3.15 36.885 3.88 ;
      RECT 35.115 3.87 35.445 4.6 ;
      RECT 33.485 7.195 33.865 12.46 ;
      RECT 25.35 3.87 25.68 4.6 ;
      RECT 21.23 3.71 21.56 4.44 ;
      RECT 20.23 3.15 20.56 3.88 ;
      RECT 18.79 3.87 19.12 4.6 ;
    LAYER via2 ;
      RECT 98.875 7.285 99.075 7.485 ;
      RECT 92.315 3.61 92.515 3.81 ;
      RECT 90.715 4.335 90.915 4.535 ;
      RECT 90.49 9.425 90.69 9.625 ;
      RECT 89.155 3.775 89.355 3.975 ;
      RECT 88.775 4.895 88.975 5.095 ;
      RECT 88.275 3.775 88.475 3.975 ;
      RECT 87.315 3.775 87.515 3.975 ;
      RECT 86.595 3.775 86.795 3.975 ;
      RECT 85.595 3.215 85.795 3.415 ;
      RECT 84.155 4.335 84.355 4.535 ;
      RECT 82.55 7.285 82.75 7.485 ;
      RECT 75.99 3.61 76.19 3.81 ;
      RECT 74.39 4.335 74.59 4.535 ;
      RECT 74.165 9.425 74.365 9.625 ;
      RECT 72.83 3.775 73.03 3.975 ;
      RECT 72.45 4.895 72.65 5.095 ;
      RECT 71.95 3.775 72.15 3.975 ;
      RECT 70.99 3.775 71.19 3.975 ;
      RECT 70.27 3.775 70.47 3.975 ;
      RECT 69.27 3.215 69.47 3.415 ;
      RECT 67.83 4.335 68.03 4.535 ;
      RECT 66.225 7.285 66.425 7.485 ;
      RECT 59.665 3.61 59.865 3.81 ;
      RECT 58.065 4.335 58.265 4.535 ;
      RECT 57.84 9.425 58.04 9.625 ;
      RECT 56.505 3.775 56.705 3.975 ;
      RECT 56.125 4.895 56.325 5.095 ;
      RECT 55.625 3.775 55.825 3.975 ;
      RECT 54.665 3.775 54.865 3.975 ;
      RECT 53.945 3.775 54.145 3.975 ;
      RECT 52.945 3.215 53.145 3.415 ;
      RECT 51.505 4.335 51.705 4.535 ;
      RECT 49.9 7.285 50.1 7.485 ;
      RECT 43.34 3.61 43.54 3.81 ;
      RECT 41.74 4.335 41.94 4.535 ;
      RECT 41.515 9.425 41.715 9.625 ;
      RECT 40.18 3.775 40.38 3.975 ;
      RECT 39.8 4.895 40 5.095 ;
      RECT 39.3 3.775 39.5 3.975 ;
      RECT 38.34 3.775 38.54 3.975 ;
      RECT 37.62 3.775 37.82 3.975 ;
      RECT 36.62 3.215 36.82 3.415 ;
      RECT 35.18 4.335 35.38 4.535 ;
      RECT 33.575 7.285 33.775 7.485 ;
      RECT 27.015 3.61 27.215 3.81 ;
      RECT 25.415 4.335 25.615 4.535 ;
      RECT 25.19 9.425 25.39 9.625 ;
      RECT 23.855 3.775 24.055 3.975 ;
      RECT 23.475 4.895 23.675 5.095 ;
      RECT 22.975 3.775 23.175 3.975 ;
      RECT 22.015 3.775 22.215 3.975 ;
      RECT 21.295 3.775 21.495 3.975 ;
      RECT 20.295 3.215 20.495 3.415 ;
      RECT 18.855 4.335 19.055 4.535 ;
    LAYER met2 ;
      RECT 16.23 10.685 99.055 10.855 ;
      RECT 98.885 9.56 99.055 10.855 ;
      RECT 16.23 8.54 16.4 10.855 ;
      RECT 98.855 9.56 99.205 9.91 ;
      RECT 16.17 8.54 16.46 8.89 ;
      RECT 95.695 8.505 96.015 8.83 ;
      RECT 95.725 7.98 95.895 8.83 ;
      RECT 95.725 7.98 95.9 8.33 ;
      RECT 95.725 7.98 96.7 8.155 ;
      RECT 96.525 3.26 96.7 8.155 ;
      RECT 96.47 3.26 96.82 3.61 ;
      RECT 96.495 8.94 96.82 9.265 ;
      RECT 95.38 9.03 96.82 9.2 ;
      RECT 95.38 3.69 95.54 9.2 ;
      RECT 95.695 3.66 96.015 3.98 ;
      RECT 95.38 3.69 96.015 3.86 ;
      RECT 85.555 3.13 85.835 3.5 ;
      RECT 85.59 2.565 85.76 3.5 ;
      RECT 94.165 2.565 94.335 3.11 ;
      RECT 94.075 2.755 94.415 3.105 ;
      RECT 94.075 2.565 94.335 3.105 ;
      RECT 85.59 2.565 94.335 2.735 ;
      RECT 90.795 3.69 91.075 4.06 ;
      RECT 89.725 3.715 89.985 4.035 ;
      RECT 92.275 3.525 92.555 3.895 ;
      RECT 92.885 3.435 93.145 3.755 ;
      RECT 89.785 2.875 89.925 4.035 ;
      RECT 90.865 2.875 91.005 4.06 ;
      RECT 91.985 3.525 93.145 3.665 ;
      RECT 91.985 2.875 92.125 3.665 ;
      RECT 89.785 2.875 92.125 3.015 ;
      RECT 89.815 5.015 91.99 5.18 ;
      RECT 91.845 3.895 91.99 5.18 ;
      RECT 88.735 4.81 89.015 5.18 ;
      RECT 88.735 4.925 89.955 5.065 ;
      RECT 91.565 3.895 91.99 4.035 ;
      RECT 91.565 3.715 91.825 4.035 ;
      RECT 84.905 5.295 88.565 5.435 ;
      RECT 88.425 4.48 88.565 5.435 ;
      RECT 84.905 4.365 85.045 5.435 ;
      RECT 91.445 4.555 91.705 4.875 ;
      RECT 88.425 4.48 90.955 4.62 ;
      RECT 90.675 4.25 90.955 4.62 ;
      RECT 84.905 4.365 85.355 4.62 ;
      RECT 85.075 4.25 85.355 4.62 ;
      RECT 91.445 4.365 91.645 4.875 ;
      RECT 90.675 4.365 91.645 4.505 ;
      RECT 91.245 3.155 91.385 4.505 ;
      RECT 91.185 3.155 91.445 3.475 ;
      RECT 82.505 8.94 82.855 9.29 ;
      RECT 91.06 8.895 91.41 9.245 ;
      RECT 82.505 8.97 91.41 9.17 ;
      RECT 85.085 3.715 85.345 4.035 ;
      RECT 85.085 3.805 86.125 3.945 ;
      RECT 85.985 3.015 86.125 3.945 ;
      RECT 88.745 3.155 89.005 3.475 ;
      RECT 85.985 3.015 88.945 3.155 ;
      RECT 88.125 3.995 88.385 4.315 ;
      RECT 88.125 3.995 88.445 4.225 ;
      RECT 88.235 3.69 88.515 4.06 ;
      RECT 87.825 4.555 88.145 4.875 ;
      RECT 87.825 3.435 87.965 4.875 ;
      RECT 87.765 3.435 88.025 3.755 ;
      RECT 85.325 4.835 85.585 5.155 ;
      RECT 85.325 4.925 87.005 5.065 ;
      RECT 86.865 4.645 87.005 5.065 ;
      RECT 86.865 4.645 87.305 4.875 ;
      RECT 87.045 4.555 87.305 4.875 ;
      RECT 86.365 3.715 86.765 4.225 ;
      RECT 86.555 3.69 86.835 4.06 ;
      RECT 86.305 3.715 86.835 4.035 ;
      RECT 79.37 8.505 79.69 8.83 ;
      RECT 79.4 7.98 79.57 8.83 ;
      RECT 79.4 7.98 79.575 8.33 ;
      RECT 79.4 7.98 80.375 8.155 ;
      RECT 80.2 3.26 80.375 8.155 ;
      RECT 80.145 3.26 80.495 3.61 ;
      RECT 80.17 8.94 80.495 9.265 ;
      RECT 79.055 9.03 80.495 9.2 ;
      RECT 79.055 3.69 79.215 9.2 ;
      RECT 79.37 3.66 79.69 3.98 ;
      RECT 79.055 3.69 79.69 3.86 ;
      RECT 69.23 3.13 69.51 3.5 ;
      RECT 69.265 2.565 69.435 3.5 ;
      RECT 77.84 2.565 78.01 3.11 ;
      RECT 77.75 2.755 78.09 3.105 ;
      RECT 77.75 2.565 78.01 3.105 ;
      RECT 69.265 2.565 78.01 2.735 ;
      RECT 74.47 3.69 74.75 4.06 ;
      RECT 73.4 3.715 73.66 4.035 ;
      RECT 75.95 3.525 76.23 3.895 ;
      RECT 76.56 3.435 76.82 3.755 ;
      RECT 73.46 2.875 73.6 4.035 ;
      RECT 74.54 2.875 74.68 4.06 ;
      RECT 75.66 3.525 76.82 3.665 ;
      RECT 75.66 2.875 75.8 3.665 ;
      RECT 73.46 2.875 75.8 3.015 ;
      RECT 73.49 5.015 75.665 5.18 ;
      RECT 75.52 3.895 75.665 5.18 ;
      RECT 72.41 4.81 72.69 5.18 ;
      RECT 72.41 4.925 73.63 5.065 ;
      RECT 75.24 3.895 75.665 4.035 ;
      RECT 75.24 3.715 75.5 4.035 ;
      RECT 68.58 5.295 72.24 5.435 ;
      RECT 72.1 4.48 72.24 5.435 ;
      RECT 68.58 4.365 68.72 5.435 ;
      RECT 75.12 4.555 75.38 4.875 ;
      RECT 72.1 4.48 74.63 4.62 ;
      RECT 74.35 4.25 74.63 4.62 ;
      RECT 68.58 4.365 69.03 4.62 ;
      RECT 68.75 4.25 69.03 4.62 ;
      RECT 75.12 4.365 75.32 4.875 ;
      RECT 74.35 4.365 75.32 4.505 ;
      RECT 74.92 3.155 75.06 4.505 ;
      RECT 74.86 3.155 75.12 3.475 ;
      RECT 66.18 8.94 66.53 9.29 ;
      RECT 74.73 8.895 75.08 9.245 ;
      RECT 66.18 8.97 75.08 9.17 ;
      RECT 68.76 3.715 69.02 4.035 ;
      RECT 68.76 3.805 69.8 3.945 ;
      RECT 69.66 3.015 69.8 3.945 ;
      RECT 72.42 3.155 72.68 3.475 ;
      RECT 69.66 3.015 72.62 3.155 ;
      RECT 71.8 3.995 72.06 4.315 ;
      RECT 71.8 3.995 72.12 4.225 ;
      RECT 71.91 3.69 72.19 4.06 ;
      RECT 71.5 4.555 71.82 4.875 ;
      RECT 71.5 3.435 71.64 4.875 ;
      RECT 71.44 3.435 71.7 3.755 ;
      RECT 69 4.835 69.26 5.155 ;
      RECT 69 4.925 70.68 5.065 ;
      RECT 70.54 4.645 70.68 5.065 ;
      RECT 70.54 4.645 70.98 4.875 ;
      RECT 70.72 4.555 70.98 4.875 ;
      RECT 70.04 3.715 70.44 4.225 ;
      RECT 70.23 3.69 70.51 4.06 ;
      RECT 69.98 3.715 70.51 4.035 ;
      RECT 63.045 8.505 63.365 8.83 ;
      RECT 63.075 7.98 63.245 8.83 ;
      RECT 63.075 7.98 63.25 8.33 ;
      RECT 63.075 7.98 64.05 8.155 ;
      RECT 63.875 3.26 64.05 8.155 ;
      RECT 63.82 3.26 64.17 3.61 ;
      RECT 63.845 8.94 64.17 9.265 ;
      RECT 62.73 9.03 64.17 9.2 ;
      RECT 62.73 3.69 62.89 9.2 ;
      RECT 63.045 3.66 63.365 3.98 ;
      RECT 62.73 3.69 63.365 3.86 ;
      RECT 52.905 3.13 53.185 3.5 ;
      RECT 52.94 2.565 53.11 3.5 ;
      RECT 61.515 2.565 61.685 3.11 ;
      RECT 61.425 2.755 61.765 3.105 ;
      RECT 61.425 2.565 61.685 3.105 ;
      RECT 52.94 2.565 61.685 2.735 ;
      RECT 58.145 3.69 58.425 4.06 ;
      RECT 57.075 3.715 57.335 4.035 ;
      RECT 59.625 3.525 59.905 3.895 ;
      RECT 60.235 3.435 60.495 3.755 ;
      RECT 57.135 2.875 57.275 4.035 ;
      RECT 58.215 2.875 58.355 4.06 ;
      RECT 59.335 3.525 60.495 3.665 ;
      RECT 59.335 2.875 59.475 3.665 ;
      RECT 57.135 2.875 59.475 3.015 ;
      RECT 57.165 5.015 59.34 5.18 ;
      RECT 59.195 3.895 59.34 5.18 ;
      RECT 56.085 4.81 56.365 5.18 ;
      RECT 56.085 4.925 57.305 5.065 ;
      RECT 58.915 3.895 59.34 4.035 ;
      RECT 58.915 3.715 59.175 4.035 ;
      RECT 52.255 5.295 55.915 5.435 ;
      RECT 55.775 4.48 55.915 5.435 ;
      RECT 52.255 4.365 52.395 5.435 ;
      RECT 58.795 4.555 59.055 4.875 ;
      RECT 55.775 4.48 58.305 4.62 ;
      RECT 58.025 4.25 58.305 4.62 ;
      RECT 52.255 4.365 52.705 4.62 ;
      RECT 52.425 4.25 52.705 4.62 ;
      RECT 58.795 4.365 58.995 4.875 ;
      RECT 58.025 4.365 58.995 4.505 ;
      RECT 58.595 3.155 58.735 4.505 ;
      RECT 58.535 3.155 58.795 3.475 ;
      RECT 49.9 8.945 50.25 9.295 ;
      RECT 58.405 8.9 58.755 9.25 ;
      RECT 49.9 8.975 58.755 9.175 ;
      RECT 52.435 3.715 52.695 4.035 ;
      RECT 52.435 3.805 53.475 3.945 ;
      RECT 53.335 3.015 53.475 3.945 ;
      RECT 56.095 3.155 56.355 3.475 ;
      RECT 53.335 3.015 56.295 3.155 ;
      RECT 55.475 3.995 55.735 4.315 ;
      RECT 55.475 3.995 55.795 4.225 ;
      RECT 55.585 3.69 55.865 4.06 ;
      RECT 55.175 4.555 55.495 4.875 ;
      RECT 55.175 3.435 55.315 4.875 ;
      RECT 55.115 3.435 55.375 3.755 ;
      RECT 52.675 4.835 52.935 5.155 ;
      RECT 52.675 4.925 54.355 5.065 ;
      RECT 54.215 4.645 54.355 5.065 ;
      RECT 54.215 4.645 54.655 4.875 ;
      RECT 54.395 4.555 54.655 4.875 ;
      RECT 53.715 3.715 54.115 4.225 ;
      RECT 53.905 3.69 54.185 4.06 ;
      RECT 53.655 3.715 54.185 4.035 ;
      RECT 46.72 8.505 47.04 8.83 ;
      RECT 46.75 7.98 46.92 8.83 ;
      RECT 46.75 7.98 46.925 8.33 ;
      RECT 46.75 7.98 47.725 8.155 ;
      RECT 47.55 3.26 47.725 8.155 ;
      RECT 47.495 3.26 47.845 3.61 ;
      RECT 47.52 8.94 47.845 9.265 ;
      RECT 46.405 9.03 47.845 9.2 ;
      RECT 46.405 3.69 46.565 9.2 ;
      RECT 46.72 3.66 47.04 3.98 ;
      RECT 46.405 3.69 47.04 3.86 ;
      RECT 36.58 3.13 36.86 3.5 ;
      RECT 36.615 2.565 36.785 3.5 ;
      RECT 45.19 2.565 45.36 3.11 ;
      RECT 45.1 2.755 45.44 3.105 ;
      RECT 45.1 2.565 45.36 3.105 ;
      RECT 36.615 2.565 45.36 2.735 ;
      RECT 41.82 3.69 42.1 4.06 ;
      RECT 40.75 3.715 41.01 4.035 ;
      RECT 43.3 3.525 43.58 3.895 ;
      RECT 43.91 3.435 44.17 3.755 ;
      RECT 40.81 2.875 40.95 4.035 ;
      RECT 41.89 2.875 42.03 4.06 ;
      RECT 43.01 3.525 44.17 3.665 ;
      RECT 43.01 2.875 43.15 3.665 ;
      RECT 40.81 2.875 43.15 3.015 ;
      RECT 40.84 5.015 43.015 5.18 ;
      RECT 42.87 3.895 43.015 5.18 ;
      RECT 39.76 4.81 40.04 5.18 ;
      RECT 39.76 4.925 40.98 5.065 ;
      RECT 42.59 3.895 43.015 4.035 ;
      RECT 42.59 3.715 42.85 4.035 ;
      RECT 35.93 5.295 39.59 5.435 ;
      RECT 39.45 4.48 39.59 5.435 ;
      RECT 35.93 4.365 36.07 5.435 ;
      RECT 42.47 4.555 42.73 4.875 ;
      RECT 39.45 4.48 41.98 4.62 ;
      RECT 41.7 4.25 41.98 4.62 ;
      RECT 35.93 4.365 36.38 4.62 ;
      RECT 36.1 4.25 36.38 4.62 ;
      RECT 42.47 4.365 42.67 4.875 ;
      RECT 41.7 4.365 42.67 4.505 ;
      RECT 42.27 3.155 42.41 4.505 ;
      RECT 42.21 3.155 42.47 3.475 ;
      RECT 33.575 8.94 33.925 9.29 ;
      RECT 42.08 8.895 42.43 9.245 ;
      RECT 33.575 8.97 42.43 9.17 ;
      RECT 36.11 3.715 36.37 4.035 ;
      RECT 36.11 3.805 37.15 3.945 ;
      RECT 37.01 3.015 37.15 3.945 ;
      RECT 39.77 3.155 40.03 3.475 ;
      RECT 37.01 3.015 39.97 3.155 ;
      RECT 39.15 3.995 39.41 4.315 ;
      RECT 39.15 3.995 39.47 4.225 ;
      RECT 39.26 3.69 39.54 4.06 ;
      RECT 38.85 4.555 39.17 4.875 ;
      RECT 38.85 3.435 38.99 4.875 ;
      RECT 38.79 3.435 39.05 3.755 ;
      RECT 36.35 4.835 36.61 5.155 ;
      RECT 36.35 4.925 38.03 5.065 ;
      RECT 37.89 4.645 38.03 5.065 ;
      RECT 37.89 4.645 38.33 4.875 ;
      RECT 38.07 4.555 38.33 4.875 ;
      RECT 37.39 3.715 37.79 4.225 ;
      RECT 37.58 3.69 37.86 4.06 ;
      RECT 37.33 3.715 37.86 4.035 ;
      RECT 30.395 8.505 30.715 8.83 ;
      RECT 30.425 7.98 30.595 8.83 ;
      RECT 30.425 7.98 30.6 8.33 ;
      RECT 30.425 7.98 31.4 8.155 ;
      RECT 31.225 3.26 31.4 8.155 ;
      RECT 31.17 3.26 31.52 3.61 ;
      RECT 31.195 8.94 31.52 9.265 ;
      RECT 30.08 9.03 31.52 9.2 ;
      RECT 30.08 3.69 30.24 9.2 ;
      RECT 30.395 3.66 30.715 3.98 ;
      RECT 30.08 3.69 30.715 3.86 ;
      RECT 20.255 3.13 20.535 3.5 ;
      RECT 20.29 2.565 20.46 3.5 ;
      RECT 28.865 2.565 29.035 3.11 ;
      RECT 28.775 2.755 29.115 3.105 ;
      RECT 28.775 2.565 29.035 3.105 ;
      RECT 20.29 2.565 29.035 2.735 ;
      RECT 25.495 3.69 25.775 4.06 ;
      RECT 24.425 3.715 24.685 4.035 ;
      RECT 26.975 3.525 27.255 3.895 ;
      RECT 27.585 3.435 27.845 3.755 ;
      RECT 24.485 2.875 24.625 4.035 ;
      RECT 25.565 2.875 25.705 4.06 ;
      RECT 26.685 3.525 27.845 3.665 ;
      RECT 26.685 2.875 26.825 3.665 ;
      RECT 24.485 2.875 26.825 3.015 ;
      RECT 16.545 9.28 16.835 9.63 ;
      RECT 16.545 9.335 17.83 9.51 ;
      RECT 17.655 8.97 17.83 9.51 ;
      RECT 26.59 8.89 26.94 9.24 ;
      RECT 17.655 8.97 26.94 9.145 ;
      RECT 24.515 5.015 26.69 5.18 ;
      RECT 26.545 3.895 26.69 5.18 ;
      RECT 23.435 4.81 23.715 5.18 ;
      RECT 23.435 4.925 24.655 5.065 ;
      RECT 26.265 3.895 26.69 4.035 ;
      RECT 26.265 3.715 26.525 4.035 ;
      RECT 19.605 5.295 23.265 5.435 ;
      RECT 23.125 4.48 23.265 5.435 ;
      RECT 19.605 4.365 19.745 5.435 ;
      RECT 26.145 4.555 26.405 4.875 ;
      RECT 23.125 4.48 25.655 4.62 ;
      RECT 25.375 4.25 25.655 4.62 ;
      RECT 19.605 4.365 20.055 4.62 ;
      RECT 19.775 4.25 20.055 4.62 ;
      RECT 26.145 4.365 26.345 4.875 ;
      RECT 25.375 4.365 26.345 4.505 ;
      RECT 25.945 3.155 26.085 4.505 ;
      RECT 25.885 3.155 26.145 3.475 ;
      RECT 19.785 3.715 20.045 4.035 ;
      RECT 19.785 3.805 20.825 3.945 ;
      RECT 20.685 3.015 20.825 3.945 ;
      RECT 23.445 3.155 23.705 3.475 ;
      RECT 20.685 3.015 23.645 3.155 ;
      RECT 22.825 3.995 23.085 4.315 ;
      RECT 22.825 3.995 23.145 4.225 ;
      RECT 22.935 3.69 23.215 4.06 ;
      RECT 22.525 4.555 22.845 4.875 ;
      RECT 22.525 3.435 22.665 4.875 ;
      RECT 22.465 3.435 22.725 3.755 ;
      RECT 20.025 4.835 20.285 5.155 ;
      RECT 20.025 4.925 21.705 5.065 ;
      RECT 21.565 4.645 21.705 5.065 ;
      RECT 21.565 4.645 22.005 4.875 ;
      RECT 21.745 4.555 22.005 4.875 ;
      RECT 21.065 3.715 21.465 4.225 ;
      RECT 21.255 3.69 21.535 4.06 ;
      RECT 21.005 3.715 21.535 4.035 ;
      RECT 98.785 7.195 99.165 7.575 ;
      RECT 90.405 9.34 90.775 9.71 ;
      RECT 89.115 3.69 89.395 4.06 ;
      RECT 87.275 3.69 87.555 4.06 ;
      RECT 84.115 4.25 84.395 4.62 ;
      RECT 82.46 7.195 82.84 7.575 ;
      RECT 74.08 9.34 74.45 9.71 ;
      RECT 72.79 3.69 73.07 4.06 ;
      RECT 70.95 3.69 71.23 4.06 ;
      RECT 67.79 4.25 68.07 4.62 ;
      RECT 66.135 7.195 66.515 7.575 ;
      RECT 57.755 9.34 58.125 9.71 ;
      RECT 56.465 3.69 56.745 4.06 ;
      RECT 54.625 3.69 54.905 4.06 ;
      RECT 51.465 4.25 51.745 4.62 ;
      RECT 49.81 7.195 50.19 7.575 ;
      RECT 41.43 9.34 41.8 9.71 ;
      RECT 40.14 3.69 40.42 4.06 ;
      RECT 38.3 3.69 38.58 4.06 ;
      RECT 35.14 4.25 35.42 4.62 ;
      RECT 33.485 7.195 33.865 7.575 ;
      RECT 25.105 9.34 25.475 9.71 ;
      RECT 23.815 3.69 24.095 4.06 ;
      RECT 21.975 3.69 22.255 4.06 ;
      RECT 18.815 4.25 19.095 4.62 ;
    LAYER via1 ;
      RECT 98.955 9.66 99.105 9.81 ;
      RECT 98.9 7.31 99.05 7.46 ;
      RECT 96.585 9.025 96.735 9.175 ;
      RECT 96.57 3.36 96.72 3.51 ;
      RECT 95.78 3.745 95.93 3.895 ;
      RECT 95.78 8.61 95.93 8.76 ;
      RECT 94.175 2.855 94.325 3.005 ;
      RECT 92.94 3.52 93.09 3.67 ;
      RECT 91.62 3.8 91.77 3.95 ;
      RECT 91.5 4.64 91.65 4.79 ;
      RECT 91.24 3.24 91.39 3.39 ;
      RECT 91.16 8.995 91.31 9.145 ;
      RECT 90.515 9.45 90.665 9.6 ;
      RECT 89.78 3.8 89.93 3.95 ;
      RECT 89.18 3.8 89.33 3.95 ;
      RECT 88.8 3.24 88.95 3.39 ;
      RECT 88.18 4.08 88.33 4.23 ;
      RECT 87.94 4.64 88.09 4.79 ;
      RECT 87.82 3.52 87.97 3.67 ;
      RECT 87.34 3.8 87.49 3.95 ;
      RECT 87.1 4.64 87.25 4.79 ;
      RECT 86.36 3.8 86.51 3.95 ;
      RECT 85.62 3.24 85.77 3.39 ;
      RECT 85.38 4.92 85.53 5.07 ;
      RECT 85.14 3.8 85.29 3.95 ;
      RECT 85.14 4.36 85.29 4.51 ;
      RECT 84.18 4.36 84.33 4.51 ;
      RECT 82.605 9.04 82.755 9.19 ;
      RECT 82.575 7.31 82.725 7.46 ;
      RECT 80.26 9.025 80.41 9.175 ;
      RECT 80.245 3.36 80.395 3.51 ;
      RECT 79.455 3.745 79.605 3.895 ;
      RECT 79.455 8.61 79.605 8.76 ;
      RECT 77.85 2.855 78 3.005 ;
      RECT 76.615 3.52 76.765 3.67 ;
      RECT 75.295 3.8 75.445 3.95 ;
      RECT 75.175 4.64 75.325 4.79 ;
      RECT 74.915 3.24 75.065 3.39 ;
      RECT 74.83 8.995 74.98 9.145 ;
      RECT 74.19 9.45 74.34 9.6 ;
      RECT 73.455 3.8 73.605 3.95 ;
      RECT 72.855 3.8 73.005 3.95 ;
      RECT 72.475 3.24 72.625 3.39 ;
      RECT 71.855 4.08 72.005 4.23 ;
      RECT 71.615 4.64 71.765 4.79 ;
      RECT 71.495 3.52 71.645 3.67 ;
      RECT 71.015 3.8 71.165 3.95 ;
      RECT 70.775 4.64 70.925 4.79 ;
      RECT 70.035 3.8 70.185 3.95 ;
      RECT 69.295 3.24 69.445 3.39 ;
      RECT 69.055 4.92 69.205 5.07 ;
      RECT 68.815 3.8 68.965 3.95 ;
      RECT 68.815 4.36 68.965 4.51 ;
      RECT 67.855 4.36 68.005 4.51 ;
      RECT 66.28 9.04 66.43 9.19 ;
      RECT 66.25 7.31 66.4 7.46 ;
      RECT 63.935 9.025 64.085 9.175 ;
      RECT 63.92 3.36 64.07 3.51 ;
      RECT 63.13 3.745 63.28 3.895 ;
      RECT 63.13 8.61 63.28 8.76 ;
      RECT 61.525 2.855 61.675 3.005 ;
      RECT 60.29 3.52 60.44 3.67 ;
      RECT 58.97 3.8 59.12 3.95 ;
      RECT 58.85 4.64 59 4.79 ;
      RECT 58.59 3.24 58.74 3.39 ;
      RECT 58.505 9 58.655 9.15 ;
      RECT 57.865 9.45 58.015 9.6 ;
      RECT 57.13 3.8 57.28 3.95 ;
      RECT 56.53 3.8 56.68 3.95 ;
      RECT 56.15 3.24 56.3 3.39 ;
      RECT 55.53 4.08 55.68 4.23 ;
      RECT 55.29 4.64 55.44 4.79 ;
      RECT 55.17 3.52 55.32 3.67 ;
      RECT 54.69 3.8 54.84 3.95 ;
      RECT 54.45 4.64 54.6 4.79 ;
      RECT 53.71 3.8 53.86 3.95 ;
      RECT 52.97 3.24 53.12 3.39 ;
      RECT 52.73 4.92 52.88 5.07 ;
      RECT 52.49 3.8 52.64 3.95 ;
      RECT 52.49 4.36 52.64 4.51 ;
      RECT 51.53 4.36 51.68 4.51 ;
      RECT 50 9.045 50.15 9.195 ;
      RECT 49.925 7.31 50.075 7.46 ;
      RECT 47.61 9.025 47.76 9.175 ;
      RECT 47.595 3.36 47.745 3.51 ;
      RECT 46.805 3.745 46.955 3.895 ;
      RECT 46.805 8.61 46.955 8.76 ;
      RECT 45.2 2.855 45.35 3.005 ;
      RECT 43.965 3.52 44.115 3.67 ;
      RECT 42.645 3.8 42.795 3.95 ;
      RECT 42.525 4.64 42.675 4.79 ;
      RECT 42.265 3.24 42.415 3.39 ;
      RECT 42.18 8.995 42.33 9.145 ;
      RECT 41.54 9.45 41.69 9.6 ;
      RECT 40.805 3.8 40.955 3.95 ;
      RECT 40.205 3.8 40.355 3.95 ;
      RECT 39.825 3.24 39.975 3.39 ;
      RECT 39.205 4.08 39.355 4.23 ;
      RECT 38.965 4.64 39.115 4.79 ;
      RECT 38.845 3.52 38.995 3.67 ;
      RECT 38.365 3.8 38.515 3.95 ;
      RECT 38.125 4.64 38.275 4.79 ;
      RECT 37.385 3.8 37.535 3.95 ;
      RECT 36.645 3.24 36.795 3.39 ;
      RECT 36.405 4.92 36.555 5.07 ;
      RECT 36.165 3.8 36.315 3.95 ;
      RECT 36.165 4.36 36.315 4.51 ;
      RECT 35.205 4.36 35.355 4.51 ;
      RECT 33.675 9.04 33.825 9.19 ;
      RECT 33.6 7.31 33.75 7.46 ;
      RECT 31.285 9.025 31.435 9.175 ;
      RECT 31.27 3.36 31.42 3.51 ;
      RECT 30.48 3.745 30.63 3.895 ;
      RECT 30.48 8.61 30.63 8.76 ;
      RECT 28.875 2.855 29.025 3.005 ;
      RECT 27.64 3.52 27.79 3.67 ;
      RECT 26.69 8.99 26.84 9.14 ;
      RECT 26.32 3.8 26.47 3.95 ;
      RECT 26.2 4.64 26.35 4.79 ;
      RECT 25.94 3.24 26.09 3.39 ;
      RECT 25.215 9.45 25.365 9.6 ;
      RECT 24.48 3.8 24.63 3.95 ;
      RECT 23.88 3.8 24.03 3.95 ;
      RECT 23.5 3.24 23.65 3.39 ;
      RECT 22.88 4.08 23.03 4.23 ;
      RECT 22.64 4.64 22.79 4.79 ;
      RECT 22.52 3.52 22.67 3.67 ;
      RECT 22.04 3.8 22.19 3.95 ;
      RECT 21.8 4.64 21.95 4.79 ;
      RECT 21.06 3.8 21.21 3.95 ;
      RECT 20.32 3.24 20.47 3.39 ;
      RECT 20.08 4.92 20.23 5.07 ;
      RECT 19.84 3.8 19.99 3.95 ;
      RECT 19.84 4.36 19.99 4.51 ;
      RECT 18.88 4.36 19.03 4.51 ;
      RECT 16.615 9.38 16.765 9.53 ;
      RECT 16.24 8.64 16.39 8.79 ;
    LAYER met1 ;
      RECT 98.825 10.05 99.12 10.28 ;
      RECT 98.885 9.56 99.06 10.28 ;
      RECT 98.855 9.56 99.205 9.91 ;
      RECT 98.885 8.57 99.055 10.28 ;
      RECT 98.825 8.57 99.115 8.8 ;
      RECT 97.83 10.055 98.125 10.285 ;
      RECT 97.89 8.575 98.06 10.285 ;
      RECT 97.83 8.575 98.12 8.805 ;
      RECT 97.83 8.61 98.685 8.77 ;
      RECT 98.515 8.2 98.685 8.77 ;
      RECT 97.83 8.605 98.225 8.77 ;
      RECT 98.455 8.2 98.745 8.43 ;
      RECT 98.455 8.23 98.915 8.4 ;
      RECT 98.415 4.03 98.74 4.26 ;
      RECT 98.415 4.06 98.91 4.23 ;
      RECT 98.415 3.69 98.605 4.26 ;
      RECT 97.83 3.655 98.12 3.885 ;
      RECT 97.83 3.69 98.605 3.86 ;
      RECT 97.89 2.175 98.06 3.885 ;
      RECT 97.83 2.175 98.125 2.405 ;
      RECT 97.46 4.025 97.75 4.255 ;
      RECT 97.46 4.055 97.92 4.225 ;
      RECT 97.525 2.95 97.69 4.255 ;
      RECT 96.04 2.915 96.33 3.145 ;
      RECT 96.04 2.95 97.69 3.12 ;
      RECT 96.1 2.175 96.27 3.145 ;
      RECT 96.04 2.175 96.33 2.405 ;
      RECT 96.04 10.055 96.33 10.285 ;
      RECT 96.1 9.315 96.27 10.285 ;
      RECT 96.1 9.405 97.69 9.575 ;
      RECT 97.52 8.205 97.69 9.575 ;
      RECT 96.04 9.315 96.33 9.545 ;
      RECT 97.46 8.205 97.75 8.435 ;
      RECT 97.46 8.235 97.92 8.405 ;
      RECT 96.47 3.26 96.82 3.61 ;
      RECT 94.165 3.32 96.82 3.49 ;
      RECT 96.3 3.315 96.82 3.49 ;
      RECT 94.165 2.755 94.335 3.49 ;
      RECT 94.075 2.755 94.415 3.105 ;
      RECT 96.495 8.94 96.82 9.265 ;
      RECT 91.06 8.895 91.41 9.245 ;
      RECT 96.47 8.945 96.82 9.175 ;
      RECT 90.855 8.945 91.41 9.175 ;
      RECT 96.3 8.97 96.82 9.145 ;
      RECT 90.685 8.975 91.41 9.145 ;
      RECT 90.855 8.97 96.82 9.14 ;
      RECT 95.695 3.66 96.015 3.98 ;
      RECT 95.67 3.655 95.96 3.885 ;
      RECT 95.665 3.685 96.015 3.86 ;
      RECT 95.495 3.685 96.015 3.855 ;
      RECT 95.695 8.54 96.015 8.83 ;
      RECT 95.67 8.575 96.015 8.805 ;
      RECT 95.495 8.605 96.015 8.775 ;
      RECT 92.15 3.76 92.44 3.99 ;
      RECT 92.15 3.76 92.605 3.945 ;
      RECT 92.465 3.665 93.085 3.805 ;
      RECT 92.855 3.465 93.175 3.725 ;
      RECT 91.535 3.745 91.855 4.005 ;
      RECT 91.535 3.745 92 3.99 ;
      RECT 91.86 3.365 92 3.99 ;
      RECT 91.86 3.365 92.125 3.505 ;
      RECT 92.39 3.2 92.68 3.43 ;
      RECT 91.985 3.245 92.68 3.385 ;
      RECT 91.43 4.585 91.72 5.11 ;
      RECT 91.415 4.585 91.735 4.845 ;
      RECT 91.155 3.185 91.475 3.445 ;
      RECT 91.155 3.2 91.72 3.43 ;
      RECT 90.43 4.88 90.72 5.11 ;
      RECT 90.625 3.525 90.765 5.065 ;
      RECT 90.67 3.48 90.96 3.71 ;
      RECT 90.265 3.525 90.96 3.665 ;
      RECT 90.265 3.365 90.405 3.665 ;
      RECT 88.805 3.365 90.405 3.505 ;
      RECT 88.715 3.185 89.035 3.445 ;
      RECT 88.715 3.2 89.28 3.445 ;
      RECT 90.425 10.055 90.715 10.285 ;
      RECT 90.485 9.315 90.655 10.285 ;
      RECT 90.405 9.36 90.775 9.71 ;
      RECT 90.405 9.34 90.715 9.71 ;
      RECT 90.425 9.315 90.715 9.71 ;
      RECT 87.825 4.225 90.405 4.365 ;
      RECT 90.19 4.04 90.48 4.27 ;
      RECT 87.75 4.04 88.415 4.27 ;
      RECT 88.095 4.025 88.415 4.365 ;
      RECT 89.095 3.745 89.415 4.005 ;
      RECT 89.095 3.76 89.52 3.99 ;
      RECT 87.735 3.465 88.055 3.725 ;
      RECT 88.23 3.48 88.52 3.71 ;
      RECT 87.735 3.525 88.52 3.665 ;
      RECT 87.855 4.585 88.175 4.845 ;
      RECT 87.015 4.585 87.335 4.845 ;
      RECT 87.855 4.6 88.28 4.83 ;
      RECT 87.015 4.645 88.28 4.785 ;
      RECT 86.55 4.32 86.84 4.55 ;
      RECT 86.625 3.245 86.765 4.55 ;
      RECT 86.275 3.745 86.765 4.005 ;
      RECT 86.03 3.76 86.765 3.99 ;
      RECT 87.03 3.2 87.32 3.43 ;
      RECT 86.625 3.245 87.32 3.385 ;
      RECT 85.79 4.6 86.08 4.83 ;
      RECT 85.79 4.6 86.245 4.785 ;
      RECT 86.105 4.225 86.245 4.785 ;
      RECT 85.745 4.225 86.245 4.365 ;
      RECT 85.745 3.245 85.885 4.365 ;
      RECT 85.535 3.185 85.855 3.445 ;
      RECT 85.295 4.865 85.615 5.125 ;
      RECT 84.59 4.88 84.88 5.11 ;
      RECT 84.59 4.925 85.615 5.065 ;
      RECT 84.665 4.875 84.925 5.065 ;
      RECT 85.055 3.745 85.375 4.005 ;
      RECT 85.055 3.76 85.6 3.99 ;
      RECT 85.055 4.305 85.375 4.565 ;
      RECT 85.055 4.32 85.6 4.55 ;
      RECT 84.095 4.305 84.415 4.565 ;
      RECT 84.185 3.245 84.325 4.565 ;
      RECT 84.59 3.2 84.88 3.43 ;
      RECT 84.185 3.245 84.88 3.385 ;
      RECT 82.5 10.05 82.795 10.28 ;
      RECT 82.56 8.57 82.73 10.28 ;
      RECT 82.505 8.94 82.855 9.29 ;
      RECT 82.5 8.57 82.79 8.8 ;
      RECT 81.505 10.055 81.8 10.285 ;
      RECT 81.565 8.575 81.735 10.285 ;
      RECT 81.505 8.575 81.795 8.805 ;
      RECT 81.505 8.61 82.36 8.77 ;
      RECT 82.19 8.2 82.36 8.77 ;
      RECT 81.505 8.605 81.9 8.77 ;
      RECT 82.13 8.2 82.42 8.43 ;
      RECT 82.13 8.23 82.59 8.4 ;
      RECT 82.09 4.03 82.415 4.26 ;
      RECT 82.09 4.06 82.585 4.23 ;
      RECT 82.09 3.69 82.28 4.26 ;
      RECT 81.505 3.655 81.795 3.885 ;
      RECT 81.505 3.69 82.28 3.86 ;
      RECT 81.565 2.175 81.735 3.885 ;
      RECT 81.505 2.175 81.8 2.405 ;
      RECT 81.135 4.025 81.425 4.255 ;
      RECT 81.135 4.055 81.595 4.225 ;
      RECT 81.2 2.95 81.365 4.255 ;
      RECT 79.715 2.915 80.005 3.145 ;
      RECT 79.715 2.95 81.365 3.12 ;
      RECT 79.775 2.175 79.945 3.145 ;
      RECT 79.715 2.175 80.005 2.405 ;
      RECT 79.715 10.055 80.005 10.285 ;
      RECT 79.775 9.315 79.945 10.285 ;
      RECT 79.775 9.405 81.365 9.575 ;
      RECT 81.195 8.205 81.365 9.575 ;
      RECT 79.715 9.315 80.005 9.545 ;
      RECT 81.135 8.205 81.425 8.435 ;
      RECT 81.135 8.235 81.595 8.405 ;
      RECT 80.145 3.26 80.495 3.61 ;
      RECT 77.84 3.32 80.495 3.49 ;
      RECT 79.975 3.315 80.495 3.49 ;
      RECT 77.84 2.755 78.01 3.49 ;
      RECT 77.75 2.755 78.09 3.105 ;
      RECT 80.17 8.94 80.495 9.265 ;
      RECT 74.73 8.895 75.08 9.245 ;
      RECT 80.145 8.945 80.495 9.175 ;
      RECT 74.53 8.945 75.08 9.175 ;
      RECT 79.975 8.97 80.495 9.145 ;
      RECT 74.36 8.975 75.08 9.145 ;
      RECT 74.53 8.97 80.495 9.14 ;
      RECT 79.37 3.66 79.69 3.98 ;
      RECT 79.345 3.655 79.635 3.885 ;
      RECT 79.34 3.685 79.69 3.86 ;
      RECT 79.17 3.685 79.69 3.855 ;
      RECT 79.37 8.54 79.69 8.83 ;
      RECT 79.345 8.575 79.69 8.805 ;
      RECT 79.17 8.605 79.69 8.775 ;
      RECT 75.825 3.76 76.115 3.99 ;
      RECT 75.825 3.76 76.28 3.945 ;
      RECT 76.14 3.665 76.76 3.805 ;
      RECT 76.53 3.465 76.85 3.725 ;
      RECT 75.21 3.745 75.53 4.005 ;
      RECT 75.21 3.745 75.675 3.99 ;
      RECT 75.535 3.365 75.675 3.99 ;
      RECT 75.535 3.365 75.8 3.505 ;
      RECT 76.065 3.2 76.355 3.43 ;
      RECT 75.66 3.245 76.355 3.385 ;
      RECT 75.105 4.585 75.395 5.11 ;
      RECT 75.09 4.585 75.41 4.845 ;
      RECT 74.83 3.185 75.15 3.445 ;
      RECT 74.83 3.2 75.395 3.43 ;
      RECT 74.105 4.88 74.395 5.11 ;
      RECT 74.3 3.525 74.44 5.065 ;
      RECT 74.345 3.48 74.635 3.71 ;
      RECT 73.94 3.525 74.635 3.665 ;
      RECT 73.94 3.365 74.08 3.665 ;
      RECT 72.48 3.365 74.08 3.505 ;
      RECT 72.39 3.185 72.71 3.445 ;
      RECT 72.39 3.2 72.955 3.445 ;
      RECT 74.1 10.055 74.39 10.285 ;
      RECT 74.16 9.315 74.33 10.285 ;
      RECT 74.08 9.36 74.45 9.71 ;
      RECT 74.08 9.34 74.39 9.71 ;
      RECT 74.1 9.315 74.39 9.71 ;
      RECT 71.5 4.225 74.08 4.365 ;
      RECT 73.865 4.04 74.155 4.27 ;
      RECT 71.425 4.04 72.09 4.27 ;
      RECT 71.77 4.025 72.09 4.365 ;
      RECT 72.77 3.745 73.09 4.005 ;
      RECT 72.77 3.76 73.195 3.99 ;
      RECT 71.41 3.465 71.73 3.725 ;
      RECT 71.905 3.48 72.195 3.71 ;
      RECT 71.41 3.525 72.195 3.665 ;
      RECT 71.53 4.585 71.85 4.845 ;
      RECT 70.69 4.585 71.01 4.845 ;
      RECT 71.53 4.6 71.955 4.83 ;
      RECT 70.69 4.645 71.955 4.785 ;
      RECT 70.225 4.32 70.515 4.55 ;
      RECT 70.3 3.245 70.44 4.55 ;
      RECT 69.95 3.745 70.44 4.005 ;
      RECT 69.705 3.76 70.44 3.99 ;
      RECT 70.705 3.2 70.995 3.43 ;
      RECT 70.3 3.245 70.995 3.385 ;
      RECT 69.465 4.6 69.755 4.83 ;
      RECT 69.465 4.6 69.92 4.785 ;
      RECT 69.78 4.225 69.92 4.785 ;
      RECT 69.42 4.225 69.92 4.365 ;
      RECT 69.42 3.245 69.56 4.365 ;
      RECT 69.21 3.185 69.53 3.445 ;
      RECT 68.97 4.865 69.29 5.125 ;
      RECT 68.265 4.88 68.555 5.11 ;
      RECT 68.265 4.925 69.29 5.065 ;
      RECT 68.34 4.875 68.6 5.065 ;
      RECT 68.73 3.745 69.05 4.005 ;
      RECT 68.73 3.76 69.275 3.99 ;
      RECT 68.73 4.305 69.05 4.565 ;
      RECT 68.73 4.32 69.275 4.55 ;
      RECT 67.77 4.305 68.09 4.565 ;
      RECT 67.86 3.245 68 4.565 ;
      RECT 68.265 3.2 68.555 3.43 ;
      RECT 67.86 3.245 68.555 3.385 ;
      RECT 66.175 10.05 66.47 10.28 ;
      RECT 66.235 8.57 66.405 10.28 ;
      RECT 66.18 8.94 66.53 9.29 ;
      RECT 66.175 8.57 66.465 8.8 ;
      RECT 65.18 10.055 65.475 10.285 ;
      RECT 65.24 8.575 65.41 10.285 ;
      RECT 65.18 8.575 65.47 8.805 ;
      RECT 65.18 8.61 66.035 8.77 ;
      RECT 65.865 8.2 66.035 8.77 ;
      RECT 65.18 8.605 65.575 8.77 ;
      RECT 65.805 8.2 66.095 8.43 ;
      RECT 65.805 8.23 66.265 8.4 ;
      RECT 65.765 4.03 66.09 4.26 ;
      RECT 65.765 4.06 66.26 4.23 ;
      RECT 65.765 3.69 65.955 4.26 ;
      RECT 65.18 3.655 65.47 3.885 ;
      RECT 65.18 3.69 65.955 3.86 ;
      RECT 65.24 2.175 65.41 3.885 ;
      RECT 65.18 2.175 65.475 2.405 ;
      RECT 64.81 4.025 65.1 4.255 ;
      RECT 64.81 4.055 65.27 4.225 ;
      RECT 64.875 2.95 65.04 4.255 ;
      RECT 63.39 2.915 63.68 3.145 ;
      RECT 63.39 2.95 65.04 3.12 ;
      RECT 63.45 2.175 63.62 3.145 ;
      RECT 63.39 2.175 63.68 2.405 ;
      RECT 63.39 10.055 63.68 10.285 ;
      RECT 63.45 9.315 63.62 10.285 ;
      RECT 63.45 9.405 65.04 9.575 ;
      RECT 64.87 8.205 65.04 9.575 ;
      RECT 63.39 9.315 63.68 9.545 ;
      RECT 64.81 8.205 65.1 8.435 ;
      RECT 64.81 8.235 65.27 8.405 ;
      RECT 63.82 3.26 64.17 3.61 ;
      RECT 61.515 3.32 64.17 3.49 ;
      RECT 63.65 3.315 64.17 3.49 ;
      RECT 61.515 2.755 61.685 3.49 ;
      RECT 61.425 2.755 61.765 3.105 ;
      RECT 63.845 8.94 64.17 9.265 ;
      RECT 58.405 8.9 58.755 9.25 ;
      RECT 63.82 8.945 64.17 9.175 ;
      RECT 58.205 8.945 58.755 9.175 ;
      RECT 63.65 8.97 64.17 9.145 ;
      RECT 58.035 8.975 58.755 9.145 ;
      RECT 58.205 8.97 64.17 9.14 ;
      RECT 63.045 3.66 63.365 3.98 ;
      RECT 63.02 3.655 63.31 3.885 ;
      RECT 63.015 3.685 63.365 3.86 ;
      RECT 62.845 3.685 63.365 3.855 ;
      RECT 63.045 8.54 63.365 8.83 ;
      RECT 63.02 8.575 63.365 8.805 ;
      RECT 62.845 8.605 63.365 8.775 ;
      RECT 59.5 3.76 59.79 3.99 ;
      RECT 59.5 3.76 59.955 3.945 ;
      RECT 59.815 3.665 60.435 3.805 ;
      RECT 60.205 3.465 60.525 3.725 ;
      RECT 58.885 3.745 59.205 4.005 ;
      RECT 58.885 3.745 59.35 3.99 ;
      RECT 59.21 3.365 59.35 3.99 ;
      RECT 59.21 3.365 59.475 3.505 ;
      RECT 59.74 3.2 60.03 3.43 ;
      RECT 59.335 3.245 60.03 3.385 ;
      RECT 58.78 4.585 59.07 5.11 ;
      RECT 58.765 4.585 59.085 4.845 ;
      RECT 58.505 3.185 58.825 3.445 ;
      RECT 58.505 3.2 59.07 3.43 ;
      RECT 57.78 4.88 58.07 5.11 ;
      RECT 57.975 3.525 58.115 5.065 ;
      RECT 58.02 3.48 58.31 3.71 ;
      RECT 57.615 3.525 58.31 3.665 ;
      RECT 57.615 3.365 57.755 3.665 ;
      RECT 56.155 3.365 57.755 3.505 ;
      RECT 56.065 3.185 56.385 3.445 ;
      RECT 56.065 3.2 56.63 3.445 ;
      RECT 57.775 10.055 58.065 10.285 ;
      RECT 57.835 9.315 58.005 10.285 ;
      RECT 57.755 9.36 58.125 9.71 ;
      RECT 57.755 9.34 58.065 9.71 ;
      RECT 57.775 9.315 58.065 9.71 ;
      RECT 55.175 4.225 57.755 4.365 ;
      RECT 57.54 4.04 57.83 4.27 ;
      RECT 55.1 4.04 55.765 4.27 ;
      RECT 55.445 4.025 55.765 4.365 ;
      RECT 56.445 3.745 56.765 4.005 ;
      RECT 56.445 3.76 56.87 3.99 ;
      RECT 55.085 3.465 55.405 3.725 ;
      RECT 55.58 3.48 55.87 3.71 ;
      RECT 55.085 3.525 55.87 3.665 ;
      RECT 55.205 4.585 55.525 4.845 ;
      RECT 54.365 4.585 54.685 4.845 ;
      RECT 55.205 4.6 55.63 4.83 ;
      RECT 54.365 4.645 55.63 4.785 ;
      RECT 53.9 4.32 54.19 4.55 ;
      RECT 53.975 3.245 54.115 4.55 ;
      RECT 53.625 3.745 54.115 4.005 ;
      RECT 53.38 3.76 54.115 3.99 ;
      RECT 54.38 3.2 54.67 3.43 ;
      RECT 53.975 3.245 54.67 3.385 ;
      RECT 53.14 4.6 53.43 4.83 ;
      RECT 53.14 4.6 53.595 4.785 ;
      RECT 53.455 4.225 53.595 4.785 ;
      RECT 53.095 4.225 53.595 4.365 ;
      RECT 53.095 3.245 53.235 4.365 ;
      RECT 52.885 3.185 53.205 3.445 ;
      RECT 52.645 4.865 52.965 5.125 ;
      RECT 51.94 4.88 52.23 5.11 ;
      RECT 51.94 4.925 52.965 5.065 ;
      RECT 52.015 4.875 52.275 5.065 ;
      RECT 52.405 3.745 52.725 4.005 ;
      RECT 52.405 3.76 52.95 3.99 ;
      RECT 52.405 4.305 52.725 4.565 ;
      RECT 52.405 4.32 52.95 4.55 ;
      RECT 51.445 4.305 51.765 4.565 ;
      RECT 51.535 3.245 51.675 4.565 ;
      RECT 51.94 3.2 52.23 3.43 ;
      RECT 51.535 3.245 52.23 3.385 ;
      RECT 49.85 10.05 50.145 10.28 ;
      RECT 49.91 8.57 50.08 10.28 ;
      RECT 49.895 8.945 50.25 9.3 ;
      RECT 49.85 8.57 50.14 8.8 ;
      RECT 48.855 10.055 49.15 10.285 ;
      RECT 48.915 8.575 49.085 10.285 ;
      RECT 48.855 8.575 49.145 8.805 ;
      RECT 48.855 8.61 49.71 8.77 ;
      RECT 49.54 8.2 49.71 8.77 ;
      RECT 48.855 8.605 49.25 8.77 ;
      RECT 49.48 8.2 49.77 8.43 ;
      RECT 49.48 8.23 49.94 8.4 ;
      RECT 49.44 4.03 49.765 4.26 ;
      RECT 49.44 4.06 49.935 4.23 ;
      RECT 49.44 3.69 49.63 4.26 ;
      RECT 48.855 3.655 49.145 3.885 ;
      RECT 48.855 3.69 49.63 3.86 ;
      RECT 48.915 2.175 49.085 3.885 ;
      RECT 48.855 2.175 49.15 2.405 ;
      RECT 48.485 4.025 48.775 4.255 ;
      RECT 48.485 4.055 48.945 4.225 ;
      RECT 48.55 2.95 48.715 4.255 ;
      RECT 47.065 2.915 47.355 3.145 ;
      RECT 47.065 2.95 48.715 3.12 ;
      RECT 47.125 2.175 47.295 3.145 ;
      RECT 47.065 2.175 47.355 2.405 ;
      RECT 47.065 10.055 47.355 10.285 ;
      RECT 47.125 9.315 47.295 10.285 ;
      RECT 47.125 9.405 48.715 9.575 ;
      RECT 48.545 8.205 48.715 9.575 ;
      RECT 47.065 9.315 47.355 9.545 ;
      RECT 48.485 8.205 48.775 8.435 ;
      RECT 48.485 8.235 48.945 8.405 ;
      RECT 47.495 3.26 47.845 3.61 ;
      RECT 45.19 3.32 47.845 3.49 ;
      RECT 47.325 3.315 47.845 3.49 ;
      RECT 45.19 2.755 45.36 3.49 ;
      RECT 45.1 2.755 45.44 3.105 ;
      RECT 47.52 8.94 47.845 9.265 ;
      RECT 42.08 8.895 42.43 9.245 ;
      RECT 47.495 8.945 47.845 9.175 ;
      RECT 41.88 8.945 42.43 9.175 ;
      RECT 47.325 8.97 47.845 9.145 ;
      RECT 41.71 8.975 42.43 9.145 ;
      RECT 41.88 8.97 47.845 9.14 ;
      RECT 46.72 3.66 47.04 3.98 ;
      RECT 46.695 3.655 46.985 3.885 ;
      RECT 46.69 3.685 47.04 3.86 ;
      RECT 46.52 3.685 47.04 3.855 ;
      RECT 46.72 8.54 47.04 8.83 ;
      RECT 46.695 8.575 47.04 8.805 ;
      RECT 46.52 8.605 47.04 8.775 ;
      RECT 43.175 3.76 43.465 3.99 ;
      RECT 43.175 3.76 43.63 3.945 ;
      RECT 43.49 3.665 44.11 3.805 ;
      RECT 43.88 3.465 44.2 3.725 ;
      RECT 42.56 3.745 42.88 4.005 ;
      RECT 42.56 3.745 43.025 3.99 ;
      RECT 42.885 3.365 43.025 3.99 ;
      RECT 42.885 3.365 43.15 3.505 ;
      RECT 43.415 3.2 43.705 3.43 ;
      RECT 43.01 3.245 43.705 3.385 ;
      RECT 42.455 4.585 42.745 5.11 ;
      RECT 42.44 4.585 42.76 4.845 ;
      RECT 42.18 3.185 42.5 3.445 ;
      RECT 42.18 3.2 42.745 3.43 ;
      RECT 41.455 4.88 41.745 5.11 ;
      RECT 41.65 3.525 41.79 5.065 ;
      RECT 41.695 3.48 41.985 3.71 ;
      RECT 41.29 3.525 41.985 3.665 ;
      RECT 41.29 3.365 41.43 3.665 ;
      RECT 39.83 3.365 41.43 3.505 ;
      RECT 39.74 3.185 40.06 3.445 ;
      RECT 39.74 3.2 40.305 3.445 ;
      RECT 41.45 10.055 41.74 10.285 ;
      RECT 41.51 9.315 41.68 10.285 ;
      RECT 41.43 9.36 41.8 9.71 ;
      RECT 41.43 9.34 41.74 9.71 ;
      RECT 41.45 9.315 41.74 9.71 ;
      RECT 38.85 4.225 41.43 4.365 ;
      RECT 41.215 4.04 41.505 4.27 ;
      RECT 38.775 4.04 39.44 4.27 ;
      RECT 39.12 4.025 39.44 4.365 ;
      RECT 40.12 3.745 40.44 4.005 ;
      RECT 40.12 3.76 40.545 3.99 ;
      RECT 38.76 3.465 39.08 3.725 ;
      RECT 39.255 3.48 39.545 3.71 ;
      RECT 38.76 3.525 39.545 3.665 ;
      RECT 38.88 4.585 39.2 4.845 ;
      RECT 38.04 4.585 38.36 4.845 ;
      RECT 38.88 4.6 39.305 4.83 ;
      RECT 38.04 4.645 39.305 4.785 ;
      RECT 37.575 4.32 37.865 4.55 ;
      RECT 37.65 3.245 37.79 4.55 ;
      RECT 37.3 3.745 37.79 4.005 ;
      RECT 37.055 3.76 37.79 3.99 ;
      RECT 38.055 3.2 38.345 3.43 ;
      RECT 37.65 3.245 38.345 3.385 ;
      RECT 36.815 4.6 37.105 4.83 ;
      RECT 36.815 4.6 37.27 4.785 ;
      RECT 37.13 4.225 37.27 4.785 ;
      RECT 36.77 4.225 37.27 4.365 ;
      RECT 36.77 3.245 36.91 4.365 ;
      RECT 36.56 3.185 36.88 3.445 ;
      RECT 36.32 4.865 36.64 5.125 ;
      RECT 35.615 4.88 35.905 5.11 ;
      RECT 35.615 4.925 36.64 5.065 ;
      RECT 35.69 4.875 35.95 5.065 ;
      RECT 36.08 3.745 36.4 4.005 ;
      RECT 36.08 3.76 36.625 3.99 ;
      RECT 36.08 4.305 36.4 4.565 ;
      RECT 36.08 4.32 36.625 4.55 ;
      RECT 35.12 4.305 35.44 4.565 ;
      RECT 35.21 3.245 35.35 4.565 ;
      RECT 35.615 3.2 35.905 3.43 ;
      RECT 35.21 3.245 35.905 3.385 ;
      RECT 33.525 10.05 33.82 10.28 ;
      RECT 33.585 8.57 33.755 10.28 ;
      RECT 33.575 8.94 33.925 9.29 ;
      RECT 33.525 8.57 33.815 8.8 ;
      RECT 32.53 10.055 32.825 10.285 ;
      RECT 32.59 8.575 32.76 10.285 ;
      RECT 32.53 8.575 32.82 8.805 ;
      RECT 32.53 8.61 33.385 8.77 ;
      RECT 33.215 8.2 33.385 8.77 ;
      RECT 32.53 8.605 32.925 8.77 ;
      RECT 33.155 8.2 33.445 8.43 ;
      RECT 33.155 8.23 33.615 8.4 ;
      RECT 33.115 4.03 33.44 4.26 ;
      RECT 33.115 4.06 33.61 4.23 ;
      RECT 33.115 3.69 33.305 4.26 ;
      RECT 32.53 3.655 32.82 3.885 ;
      RECT 32.53 3.69 33.305 3.86 ;
      RECT 32.59 2.175 32.76 3.885 ;
      RECT 32.53 2.175 32.825 2.405 ;
      RECT 32.16 4.025 32.45 4.255 ;
      RECT 32.16 4.055 32.62 4.225 ;
      RECT 32.225 2.95 32.39 4.255 ;
      RECT 30.74 2.915 31.03 3.145 ;
      RECT 30.74 2.95 32.39 3.12 ;
      RECT 30.8 2.175 30.97 3.145 ;
      RECT 30.74 2.175 31.03 2.405 ;
      RECT 30.74 10.055 31.03 10.285 ;
      RECT 30.8 9.315 30.97 10.285 ;
      RECT 30.8 9.405 32.39 9.575 ;
      RECT 32.22 8.205 32.39 9.575 ;
      RECT 30.74 9.315 31.03 9.545 ;
      RECT 32.16 8.205 32.45 8.435 ;
      RECT 32.16 8.235 32.62 8.405 ;
      RECT 31.17 3.26 31.52 3.61 ;
      RECT 28.865 3.32 31.52 3.49 ;
      RECT 31 3.315 31.52 3.49 ;
      RECT 28.865 2.755 29.035 3.49 ;
      RECT 28.775 2.755 29.115 3.105 ;
      RECT 31.195 8.94 31.52 9.265 ;
      RECT 26.59 8.89 26.94 9.24 ;
      RECT 31.17 8.945 31.52 9.175 ;
      RECT 25.555 8.945 25.845 9.175 ;
      RECT 31 8.97 31.52 9.145 ;
      RECT 25.385 8.975 25.845 9.145 ;
      RECT 25.555 8.97 31.52 9.14 ;
      RECT 30.395 3.66 30.715 3.98 ;
      RECT 30.37 3.655 30.66 3.885 ;
      RECT 30.365 3.685 30.715 3.86 ;
      RECT 30.195 3.685 30.715 3.855 ;
      RECT 30.395 8.54 30.715 8.83 ;
      RECT 30.37 8.575 30.715 8.805 ;
      RECT 30.195 8.605 30.715 8.775 ;
      RECT 26.85 3.76 27.14 3.99 ;
      RECT 26.85 3.76 27.305 3.945 ;
      RECT 27.165 3.665 27.785 3.805 ;
      RECT 27.555 3.465 27.875 3.725 ;
      RECT 26.235 3.745 26.555 4.005 ;
      RECT 26.235 3.745 26.7 3.99 ;
      RECT 26.56 3.365 26.7 3.99 ;
      RECT 26.56 3.365 26.825 3.505 ;
      RECT 27.09 3.2 27.38 3.43 ;
      RECT 26.685 3.245 27.38 3.385 ;
      RECT 26.13 4.585 26.42 5.11 ;
      RECT 26.115 4.585 26.435 4.845 ;
      RECT 25.855 3.185 26.175 3.445 ;
      RECT 25.855 3.2 26.42 3.43 ;
      RECT 25.13 4.88 25.42 5.11 ;
      RECT 25.325 3.525 25.465 5.065 ;
      RECT 25.37 3.48 25.66 3.71 ;
      RECT 24.965 3.525 25.66 3.665 ;
      RECT 24.965 3.365 25.105 3.665 ;
      RECT 23.505 3.365 25.105 3.505 ;
      RECT 23.415 3.185 23.735 3.445 ;
      RECT 23.415 3.2 23.98 3.445 ;
      RECT 25.125 10.055 25.415 10.285 ;
      RECT 25.185 9.315 25.355 10.285 ;
      RECT 25.105 9.36 25.475 9.71 ;
      RECT 25.105 9.34 25.415 9.71 ;
      RECT 25.125 9.315 25.415 9.71 ;
      RECT 22.525 4.225 25.105 4.365 ;
      RECT 24.89 4.04 25.18 4.27 ;
      RECT 22.45 4.04 23.115 4.27 ;
      RECT 22.795 4.025 23.115 4.365 ;
      RECT 23.795 3.745 24.115 4.005 ;
      RECT 23.795 3.76 24.22 3.99 ;
      RECT 22.435 3.465 22.755 3.725 ;
      RECT 22.93 3.48 23.22 3.71 ;
      RECT 22.435 3.525 23.22 3.665 ;
      RECT 22.555 4.585 22.875 4.845 ;
      RECT 21.715 4.585 22.035 4.845 ;
      RECT 22.555 4.6 22.98 4.83 ;
      RECT 21.715 4.645 22.98 4.785 ;
      RECT 21.25 4.32 21.54 4.55 ;
      RECT 21.325 3.245 21.465 4.55 ;
      RECT 20.975 3.745 21.465 4.005 ;
      RECT 20.73 3.76 21.465 3.99 ;
      RECT 21.73 3.2 22.02 3.43 ;
      RECT 21.325 3.245 22.02 3.385 ;
      RECT 20.49 4.6 20.78 4.83 ;
      RECT 20.49 4.6 20.945 4.785 ;
      RECT 20.805 4.225 20.945 4.785 ;
      RECT 20.445 4.225 20.945 4.365 ;
      RECT 20.445 3.245 20.585 4.365 ;
      RECT 20.235 3.185 20.555 3.445 ;
      RECT 19.995 4.865 20.315 5.125 ;
      RECT 19.29 4.88 19.58 5.11 ;
      RECT 19.29 4.925 20.315 5.065 ;
      RECT 19.365 4.875 19.625 5.065 ;
      RECT 19.755 3.745 20.075 4.005 ;
      RECT 19.755 3.76 20.3 3.99 ;
      RECT 19.755 4.305 20.075 4.565 ;
      RECT 19.755 4.32 20.3 4.55 ;
      RECT 18.795 4.305 19.115 4.565 ;
      RECT 18.885 3.245 19.025 4.565 ;
      RECT 19.29 3.2 19.58 3.43 ;
      RECT 18.885 3.245 19.58 3.385 ;
      RECT 16.545 10.055 16.835 10.285 ;
      RECT 16.605 9.31 16.775 10.285 ;
      RECT 16.515 9.31 16.865 9.6 ;
      RECT 16.14 8.57 16.49 8.86 ;
      RECT 16 8.605 16.49 8.775 ;
      RECT 98.8 7.24 99.15 7.53 ;
      RECT 89.695 3.745 90.015 4.005 ;
      RECT 87.255 3.745 87.575 4.005 ;
      RECT 82.475 7.24 82.825 7.53 ;
      RECT 73.37 3.745 73.69 4.005 ;
      RECT 70.93 3.745 71.25 4.005 ;
      RECT 66.15 7.24 66.5 7.53 ;
      RECT 57.045 3.745 57.365 4.005 ;
      RECT 54.605 3.745 54.925 4.005 ;
      RECT 49.825 7.24 50.175 7.53 ;
      RECT 40.72 3.745 41.04 4.005 ;
      RECT 38.28 3.745 38.6 4.005 ;
      RECT 33.5 7.24 33.85 7.53 ;
      RECT 24.395 3.745 24.715 4.005 ;
      RECT 21.955 3.745 22.275 4.005 ;
    LAYER mcon ;
      RECT 98.89 7.3 99.06 7.47 ;
      RECT 98.885 8.6 99.055 8.77 ;
      RECT 98.885 10.08 99.055 10.25 ;
      RECT 98.515 8.23 98.685 8.4 ;
      RECT 98.51 4.06 98.68 4.23 ;
      RECT 97.89 2.205 98.06 2.375 ;
      RECT 97.89 3.685 98.06 3.855 ;
      RECT 97.89 8.605 98.06 8.775 ;
      RECT 97.89 10.085 98.06 10.255 ;
      RECT 97.52 4.055 97.69 4.225 ;
      RECT 97.52 8.235 97.69 8.405 ;
      RECT 96.53 3.315 96.7 3.485 ;
      RECT 96.53 8.975 96.7 9.145 ;
      RECT 96.1 2.205 96.27 2.375 ;
      RECT 96.1 2.945 96.27 3.115 ;
      RECT 96.1 9.345 96.27 9.515 ;
      RECT 96.1 10.085 96.27 10.255 ;
      RECT 95.73 3.685 95.9 3.855 ;
      RECT 95.73 8.605 95.9 8.775 ;
      RECT 92.45 3.23 92.62 3.4 ;
      RECT 92.21 3.79 92.38 3.96 ;
      RECT 91.73 3.79 91.9 3.96 ;
      RECT 91.49 3.23 91.66 3.4 ;
      RECT 91.49 4.91 91.66 5.08 ;
      RECT 90.915 8.975 91.085 9.145 ;
      RECT 90.73 3.51 90.9 3.68 ;
      RECT 90.49 4.91 90.66 5.08 ;
      RECT 90.485 9.345 90.655 9.515 ;
      RECT 90.485 10.085 90.655 10.255 ;
      RECT 90.25 4.07 90.42 4.24 ;
      RECT 89.77 3.79 89.94 3.96 ;
      RECT 89.29 3.79 89.46 3.96 ;
      RECT 89.05 3.23 89.22 3.4 ;
      RECT 88.29 3.51 88.46 3.68 ;
      RECT 88.05 4.63 88.22 4.8 ;
      RECT 87.81 4.07 87.98 4.24 ;
      RECT 87.33 3.79 87.5 3.96 ;
      RECT 87.09 3.23 87.26 3.4 ;
      RECT 87.09 4.63 87.26 4.8 ;
      RECT 86.61 4.35 86.78 4.52 ;
      RECT 86.09 3.79 86.26 3.96 ;
      RECT 85.85 4.63 86.02 4.8 ;
      RECT 85.61 3.23 85.78 3.4 ;
      RECT 85.37 3.79 85.54 3.96 ;
      RECT 85.37 4.35 85.54 4.52 ;
      RECT 84.65 3.23 84.82 3.4 ;
      RECT 84.65 4.91 84.82 5.08 ;
      RECT 84.17 4.35 84.34 4.52 ;
      RECT 82.565 7.3 82.735 7.47 ;
      RECT 82.56 8.6 82.73 8.77 ;
      RECT 82.56 10.08 82.73 10.25 ;
      RECT 82.19 8.23 82.36 8.4 ;
      RECT 82.185 4.06 82.355 4.23 ;
      RECT 81.565 2.205 81.735 2.375 ;
      RECT 81.565 3.685 81.735 3.855 ;
      RECT 81.565 8.605 81.735 8.775 ;
      RECT 81.565 10.085 81.735 10.255 ;
      RECT 81.195 4.055 81.365 4.225 ;
      RECT 81.195 8.235 81.365 8.405 ;
      RECT 80.205 3.315 80.375 3.485 ;
      RECT 80.205 8.975 80.375 9.145 ;
      RECT 79.775 2.205 79.945 2.375 ;
      RECT 79.775 2.945 79.945 3.115 ;
      RECT 79.775 9.345 79.945 9.515 ;
      RECT 79.775 10.085 79.945 10.255 ;
      RECT 79.405 3.685 79.575 3.855 ;
      RECT 79.405 8.605 79.575 8.775 ;
      RECT 76.125 3.23 76.295 3.4 ;
      RECT 75.885 3.79 76.055 3.96 ;
      RECT 75.405 3.79 75.575 3.96 ;
      RECT 75.165 3.23 75.335 3.4 ;
      RECT 75.165 4.91 75.335 5.08 ;
      RECT 74.59 8.975 74.76 9.145 ;
      RECT 74.405 3.51 74.575 3.68 ;
      RECT 74.165 4.91 74.335 5.08 ;
      RECT 74.16 9.345 74.33 9.515 ;
      RECT 74.16 10.085 74.33 10.255 ;
      RECT 73.925 4.07 74.095 4.24 ;
      RECT 73.445 3.79 73.615 3.96 ;
      RECT 72.965 3.79 73.135 3.96 ;
      RECT 72.725 3.23 72.895 3.4 ;
      RECT 71.965 3.51 72.135 3.68 ;
      RECT 71.725 4.63 71.895 4.8 ;
      RECT 71.485 4.07 71.655 4.24 ;
      RECT 71.005 3.79 71.175 3.96 ;
      RECT 70.765 3.23 70.935 3.4 ;
      RECT 70.765 4.63 70.935 4.8 ;
      RECT 70.285 4.35 70.455 4.52 ;
      RECT 69.765 3.79 69.935 3.96 ;
      RECT 69.525 4.63 69.695 4.8 ;
      RECT 69.285 3.23 69.455 3.4 ;
      RECT 69.045 3.79 69.215 3.96 ;
      RECT 69.045 4.35 69.215 4.52 ;
      RECT 68.325 3.23 68.495 3.4 ;
      RECT 68.325 4.91 68.495 5.08 ;
      RECT 67.845 4.35 68.015 4.52 ;
      RECT 66.24 7.3 66.41 7.47 ;
      RECT 66.235 8.6 66.405 8.77 ;
      RECT 66.235 10.08 66.405 10.25 ;
      RECT 65.865 8.23 66.035 8.4 ;
      RECT 65.86 4.06 66.03 4.23 ;
      RECT 65.24 2.205 65.41 2.375 ;
      RECT 65.24 3.685 65.41 3.855 ;
      RECT 65.24 8.605 65.41 8.775 ;
      RECT 65.24 10.085 65.41 10.255 ;
      RECT 64.87 4.055 65.04 4.225 ;
      RECT 64.87 8.235 65.04 8.405 ;
      RECT 63.88 3.315 64.05 3.485 ;
      RECT 63.88 8.975 64.05 9.145 ;
      RECT 63.45 2.205 63.62 2.375 ;
      RECT 63.45 2.945 63.62 3.115 ;
      RECT 63.45 9.345 63.62 9.515 ;
      RECT 63.45 10.085 63.62 10.255 ;
      RECT 63.08 3.685 63.25 3.855 ;
      RECT 63.08 8.605 63.25 8.775 ;
      RECT 59.8 3.23 59.97 3.4 ;
      RECT 59.56 3.79 59.73 3.96 ;
      RECT 59.08 3.79 59.25 3.96 ;
      RECT 58.84 3.23 59.01 3.4 ;
      RECT 58.84 4.91 59.01 5.08 ;
      RECT 58.265 8.975 58.435 9.145 ;
      RECT 58.08 3.51 58.25 3.68 ;
      RECT 57.84 4.91 58.01 5.08 ;
      RECT 57.835 9.345 58.005 9.515 ;
      RECT 57.835 10.085 58.005 10.255 ;
      RECT 57.6 4.07 57.77 4.24 ;
      RECT 57.12 3.79 57.29 3.96 ;
      RECT 56.64 3.79 56.81 3.96 ;
      RECT 56.4 3.23 56.57 3.4 ;
      RECT 55.64 3.51 55.81 3.68 ;
      RECT 55.4 4.63 55.57 4.8 ;
      RECT 55.16 4.07 55.33 4.24 ;
      RECT 54.68 3.79 54.85 3.96 ;
      RECT 54.44 3.23 54.61 3.4 ;
      RECT 54.44 4.63 54.61 4.8 ;
      RECT 53.96 4.35 54.13 4.52 ;
      RECT 53.44 3.79 53.61 3.96 ;
      RECT 53.2 4.63 53.37 4.8 ;
      RECT 52.96 3.23 53.13 3.4 ;
      RECT 52.72 3.79 52.89 3.96 ;
      RECT 52.72 4.35 52.89 4.52 ;
      RECT 52 3.23 52.17 3.4 ;
      RECT 52 4.91 52.17 5.08 ;
      RECT 51.52 4.35 51.69 4.52 ;
      RECT 49.915 7.3 50.085 7.47 ;
      RECT 49.91 8.6 50.08 8.77 ;
      RECT 49.91 10.08 50.08 10.25 ;
      RECT 49.54 8.23 49.71 8.4 ;
      RECT 49.535 4.06 49.705 4.23 ;
      RECT 48.915 2.205 49.085 2.375 ;
      RECT 48.915 3.685 49.085 3.855 ;
      RECT 48.915 8.605 49.085 8.775 ;
      RECT 48.915 10.085 49.085 10.255 ;
      RECT 48.545 4.055 48.715 4.225 ;
      RECT 48.545 8.235 48.715 8.405 ;
      RECT 47.555 3.315 47.725 3.485 ;
      RECT 47.555 8.975 47.725 9.145 ;
      RECT 47.125 2.205 47.295 2.375 ;
      RECT 47.125 2.945 47.295 3.115 ;
      RECT 47.125 9.345 47.295 9.515 ;
      RECT 47.125 10.085 47.295 10.255 ;
      RECT 46.755 3.685 46.925 3.855 ;
      RECT 46.755 8.605 46.925 8.775 ;
      RECT 43.475 3.23 43.645 3.4 ;
      RECT 43.235 3.79 43.405 3.96 ;
      RECT 42.755 3.79 42.925 3.96 ;
      RECT 42.515 3.23 42.685 3.4 ;
      RECT 42.515 4.91 42.685 5.08 ;
      RECT 41.94 8.975 42.11 9.145 ;
      RECT 41.755 3.51 41.925 3.68 ;
      RECT 41.515 4.91 41.685 5.08 ;
      RECT 41.51 9.345 41.68 9.515 ;
      RECT 41.51 10.085 41.68 10.255 ;
      RECT 41.275 4.07 41.445 4.24 ;
      RECT 40.795 3.79 40.965 3.96 ;
      RECT 40.315 3.79 40.485 3.96 ;
      RECT 40.075 3.23 40.245 3.4 ;
      RECT 39.315 3.51 39.485 3.68 ;
      RECT 39.075 4.63 39.245 4.8 ;
      RECT 38.835 4.07 39.005 4.24 ;
      RECT 38.355 3.79 38.525 3.96 ;
      RECT 38.115 3.23 38.285 3.4 ;
      RECT 38.115 4.63 38.285 4.8 ;
      RECT 37.635 4.35 37.805 4.52 ;
      RECT 37.115 3.79 37.285 3.96 ;
      RECT 36.875 4.63 37.045 4.8 ;
      RECT 36.635 3.23 36.805 3.4 ;
      RECT 36.395 3.79 36.565 3.96 ;
      RECT 36.395 4.35 36.565 4.52 ;
      RECT 35.675 3.23 35.845 3.4 ;
      RECT 35.675 4.91 35.845 5.08 ;
      RECT 35.195 4.35 35.365 4.52 ;
      RECT 33.59 7.3 33.76 7.47 ;
      RECT 33.585 8.6 33.755 8.77 ;
      RECT 33.585 10.08 33.755 10.25 ;
      RECT 33.215 8.23 33.385 8.4 ;
      RECT 33.21 4.06 33.38 4.23 ;
      RECT 32.59 2.205 32.76 2.375 ;
      RECT 32.59 3.685 32.76 3.855 ;
      RECT 32.59 8.605 32.76 8.775 ;
      RECT 32.59 10.085 32.76 10.255 ;
      RECT 32.22 4.055 32.39 4.225 ;
      RECT 32.22 8.235 32.39 8.405 ;
      RECT 31.23 3.315 31.4 3.485 ;
      RECT 31.23 8.975 31.4 9.145 ;
      RECT 30.8 2.205 30.97 2.375 ;
      RECT 30.8 2.945 30.97 3.115 ;
      RECT 30.8 9.345 30.97 9.515 ;
      RECT 30.8 10.085 30.97 10.255 ;
      RECT 30.43 3.685 30.6 3.855 ;
      RECT 30.43 8.605 30.6 8.775 ;
      RECT 27.15 3.23 27.32 3.4 ;
      RECT 26.91 3.79 27.08 3.96 ;
      RECT 26.43 3.79 26.6 3.96 ;
      RECT 26.19 3.23 26.36 3.4 ;
      RECT 26.19 4.91 26.36 5.08 ;
      RECT 25.615 8.975 25.785 9.145 ;
      RECT 25.43 3.51 25.6 3.68 ;
      RECT 25.19 4.91 25.36 5.08 ;
      RECT 25.185 9.345 25.355 9.515 ;
      RECT 25.185 10.085 25.355 10.255 ;
      RECT 24.95 4.07 25.12 4.24 ;
      RECT 24.47 3.79 24.64 3.96 ;
      RECT 23.99 3.79 24.16 3.96 ;
      RECT 23.75 3.23 23.92 3.4 ;
      RECT 22.99 3.51 23.16 3.68 ;
      RECT 22.75 4.63 22.92 4.8 ;
      RECT 22.51 4.07 22.68 4.24 ;
      RECT 22.03 3.79 22.2 3.96 ;
      RECT 21.79 3.23 21.96 3.4 ;
      RECT 21.79 4.63 21.96 4.8 ;
      RECT 21.31 4.35 21.48 4.52 ;
      RECT 20.79 3.79 20.96 3.96 ;
      RECT 20.55 4.63 20.72 4.8 ;
      RECT 20.31 3.23 20.48 3.4 ;
      RECT 20.07 3.79 20.24 3.96 ;
      RECT 20.07 4.35 20.24 4.52 ;
      RECT 19.35 3.23 19.52 3.4 ;
      RECT 19.35 4.91 19.52 5.08 ;
      RECT 18.87 4.35 19.04 4.52 ;
      RECT 16.605 9.345 16.775 9.515 ;
      RECT 16.605 10.085 16.775 10.255 ;
      RECT 16.235 8.605 16.405 8.775 ;
    LAYER li1 ;
      RECT 98.885 7.3 99.055 8.77 ;
      RECT 98.885 7.3 99.06 8.56 ;
      RECT 98.515 9.25 98.985 9.42 ;
      RECT 98.515 8.23 98.685 9.42 ;
      RECT 98.51 3.04 98.68 4.23 ;
      RECT 98.51 3.04 98.98 3.21 ;
      RECT 97.89 3.895 98.065 5.155 ;
      RECT 97.89 3.685 98.06 5.155 ;
      RECT 97.89 7.305 98.06 8.775 ;
      RECT 97.89 7.305 98.065 8.565 ;
      RECT 97.52 3.035 97.69 4.225 ;
      RECT 97.52 3.035 97.99 3.205 ;
      RECT 97.52 9.255 97.99 9.425 ;
      RECT 97.52 8.235 97.69 9.425 ;
      RECT 96.53 4.015 96.705 5.155 ;
      RECT 96.53 1.865 96.7 5.155 ;
      RECT 96.53 1.865 96.705 2.415 ;
      RECT 96.53 10.045 96.705 10.595 ;
      RECT 96.53 7.305 96.7 10.595 ;
      RECT 96.53 7.305 96.705 8.445 ;
      RECT 96.1 3.895 96.275 5.155 ;
      RECT 96.1 2.945 96.27 5.155 ;
      RECT 96.1 7.305 96.27 9.515 ;
      RECT 96.1 7.305 96.275 8.565 ;
      RECT 95.67 3.925 95.84 5.155 ;
      RECT 95.73 2.145 95.9 4.095 ;
      RECT 95.67 1.865 95.84 2.315 ;
      RECT 95.67 10.145 95.84 10.595 ;
      RECT 95.73 8.365 95.9 10.315 ;
      RECT 95.67 7.305 95.84 8.535 ;
      RECT 95.145 3.895 95.32 5.155 ;
      RECT 95.145 1.865 95.315 5.155 ;
      RECT 95.145 3.365 95.555 3.695 ;
      RECT 95.145 2.525 95.555 2.855 ;
      RECT 95.145 1.865 95.32 2.355 ;
      RECT 95.145 10.105 95.32 10.595 ;
      RECT 95.145 7.305 95.315 10.595 ;
      RECT 95.145 9.605 95.555 9.935 ;
      RECT 95.145 8.765 95.555 9.095 ;
      RECT 95.145 7.305 95.32 8.565 ;
      RECT 92.45 3.13 92.62 3.4 ;
      RECT 92.45 3.13 93.18 3.3 ;
      RECT 92.37 4.52 92.7 4.69 ;
      RECT 91.61 4.35 92.62 4.52 ;
      RECT 91.61 3.87 91.78 4.52 ;
      RECT 91.73 3.79 91.9 4.12 ;
      RECT 90.89 4.52 91.22 4.69 ;
      RECT 88.97 4.52 90.26 4.69 ;
      RECT 90.01 4.435 91.14 4.605 ;
      RECT 90.73 3.51 91.14 3.68 ;
      RECT 90.97 3.05 91.14 3.68 ;
      RECT 90.915 10.045 91.09 10.595 ;
      RECT 90.915 7.305 91.085 10.595 ;
      RECT 90.915 7.305 91.09 8.445 ;
      RECT 90.485 7.305 90.655 9.515 ;
      RECT 90.485 7.305 90.66 8.565 ;
      RECT 89.53 10.105 89.705 10.595 ;
      RECT 89.53 7.305 89.7 10.595 ;
      RECT 89.53 9.605 89.94 9.935 ;
      RECT 89.53 8.765 89.94 9.095 ;
      RECT 89.53 7.305 89.705 8.565 ;
      RECT 88.21 3.87 89.54 4.04 ;
      RECT 89.29 3.79 89.46 4.04 ;
      RECT 88.29 3.47 88.46 3.68 ;
      RECT 88.29 3.47 88.78 3.64 ;
      RECT 86.97 4.63 87.26 4.8 ;
      RECT 86.97 3.87 87.14 4.8 ;
      RECT 86.77 3.87 87.14 4.04 ;
      RECT 85.77 3.87 86.26 4.04 ;
      RECT 86.09 3.79 86.26 4.04 ;
      RECT 85.85 4.63 86.26 4.8 ;
      RECT 86.09 4.44 86.26 4.8 ;
      RECT 84.89 4.35 85.54 4.52 ;
      RECT 84.89 3.79 85.06 4.52 ;
      RECT 84.53 4.91 84.82 5.08 ;
      RECT 84.53 3.87 84.7 5.08 ;
      RECT 84.33 3.87 84.7 4.04 ;
      RECT 82.56 7.3 82.73 8.77 ;
      RECT 82.56 7.3 82.735 8.56 ;
      RECT 82.19 9.25 82.66 9.42 ;
      RECT 82.19 8.23 82.36 9.42 ;
      RECT 82.185 3.04 82.355 4.23 ;
      RECT 82.185 3.04 82.655 3.21 ;
      RECT 81.565 3.895 81.74 5.155 ;
      RECT 81.565 3.685 81.735 5.155 ;
      RECT 81.565 7.305 81.735 8.775 ;
      RECT 81.565 7.305 81.74 8.565 ;
      RECT 81.195 3.035 81.365 4.225 ;
      RECT 81.195 3.035 81.665 3.205 ;
      RECT 81.195 9.255 81.665 9.425 ;
      RECT 81.195 8.235 81.365 9.425 ;
      RECT 80.205 4.015 80.38 5.155 ;
      RECT 80.205 1.865 80.375 5.155 ;
      RECT 80.205 1.865 80.38 2.415 ;
      RECT 80.205 10.045 80.38 10.595 ;
      RECT 80.205 7.305 80.375 10.595 ;
      RECT 80.205 7.305 80.38 8.445 ;
      RECT 79.775 3.895 79.95 5.155 ;
      RECT 79.775 2.945 79.945 5.155 ;
      RECT 79.775 7.305 79.945 9.515 ;
      RECT 79.775 7.305 79.95 8.565 ;
      RECT 79.345 3.925 79.515 5.155 ;
      RECT 79.405 2.145 79.575 4.095 ;
      RECT 79.345 1.865 79.515 2.315 ;
      RECT 79.345 10.145 79.515 10.595 ;
      RECT 79.405 8.365 79.575 10.315 ;
      RECT 79.345 7.305 79.515 8.535 ;
      RECT 78.82 3.895 78.995 5.155 ;
      RECT 78.82 1.865 78.99 5.155 ;
      RECT 78.82 3.365 79.23 3.695 ;
      RECT 78.82 2.525 79.23 2.855 ;
      RECT 78.82 1.865 78.995 2.355 ;
      RECT 78.82 10.105 78.995 10.595 ;
      RECT 78.82 7.305 78.99 10.595 ;
      RECT 78.82 9.605 79.23 9.935 ;
      RECT 78.82 8.765 79.23 9.095 ;
      RECT 78.82 7.305 78.995 8.565 ;
      RECT 76.125 3.13 76.295 3.4 ;
      RECT 76.125 3.13 76.855 3.3 ;
      RECT 76.045 4.52 76.375 4.69 ;
      RECT 75.285 4.35 76.295 4.52 ;
      RECT 75.285 3.87 75.455 4.52 ;
      RECT 75.405 3.79 75.575 4.12 ;
      RECT 74.565 4.52 74.895 4.69 ;
      RECT 72.645 4.52 73.935 4.69 ;
      RECT 73.685 4.435 74.815 4.605 ;
      RECT 74.405 3.51 74.815 3.68 ;
      RECT 74.645 3.05 74.815 3.68 ;
      RECT 74.59 10.045 74.765 10.595 ;
      RECT 74.59 7.305 74.76 10.595 ;
      RECT 74.59 7.305 74.765 8.445 ;
      RECT 74.16 7.305 74.33 9.515 ;
      RECT 74.16 7.305 74.335 8.565 ;
      RECT 73.205 10.105 73.38 10.595 ;
      RECT 73.205 7.305 73.375 10.595 ;
      RECT 73.205 9.605 73.615 9.935 ;
      RECT 73.205 8.765 73.615 9.095 ;
      RECT 73.205 7.305 73.38 8.565 ;
      RECT 71.885 3.87 73.215 4.04 ;
      RECT 72.965 3.79 73.135 4.04 ;
      RECT 71.965 3.47 72.135 3.68 ;
      RECT 71.965 3.47 72.455 3.64 ;
      RECT 70.645 4.63 70.935 4.8 ;
      RECT 70.645 3.87 70.815 4.8 ;
      RECT 70.445 3.87 70.815 4.04 ;
      RECT 69.445 3.87 69.935 4.04 ;
      RECT 69.765 3.79 69.935 4.04 ;
      RECT 69.525 4.63 69.935 4.8 ;
      RECT 69.765 4.44 69.935 4.8 ;
      RECT 68.565 4.35 69.215 4.52 ;
      RECT 68.565 3.79 68.735 4.52 ;
      RECT 68.205 4.91 68.495 5.08 ;
      RECT 68.205 3.87 68.375 5.08 ;
      RECT 68.005 3.87 68.375 4.04 ;
      RECT 66.235 7.3 66.405 8.77 ;
      RECT 66.235 7.3 66.41 8.56 ;
      RECT 65.865 9.25 66.335 9.42 ;
      RECT 65.865 8.23 66.035 9.42 ;
      RECT 65.86 3.04 66.03 4.23 ;
      RECT 65.86 3.04 66.33 3.21 ;
      RECT 65.24 3.895 65.415 5.155 ;
      RECT 65.24 3.685 65.41 5.155 ;
      RECT 65.24 7.305 65.41 8.775 ;
      RECT 65.24 7.305 65.415 8.565 ;
      RECT 64.87 3.035 65.04 4.225 ;
      RECT 64.87 3.035 65.34 3.205 ;
      RECT 64.87 9.255 65.34 9.425 ;
      RECT 64.87 8.235 65.04 9.425 ;
      RECT 63.88 4.015 64.055 5.155 ;
      RECT 63.88 1.865 64.05 5.155 ;
      RECT 63.88 1.865 64.055 2.415 ;
      RECT 63.88 10.045 64.055 10.595 ;
      RECT 63.88 7.305 64.05 10.595 ;
      RECT 63.88 7.305 64.055 8.445 ;
      RECT 63.45 3.895 63.625 5.155 ;
      RECT 63.45 2.945 63.62 5.155 ;
      RECT 63.45 7.305 63.62 9.515 ;
      RECT 63.45 7.305 63.625 8.565 ;
      RECT 63.02 3.925 63.19 5.155 ;
      RECT 63.08 2.145 63.25 4.095 ;
      RECT 63.02 1.865 63.19 2.315 ;
      RECT 63.02 10.145 63.19 10.595 ;
      RECT 63.08 8.365 63.25 10.315 ;
      RECT 63.02 7.305 63.19 8.535 ;
      RECT 62.495 3.895 62.67 5.155 ;
      RECT 62.495 1.865 62.665 5.155 ;
      RECT 62.495 3.365 62.905 3.695 ;
      RECT 62.495 2.525 62.905 2.855 ;
      RECT 62.495 1.865 62.67 2.355 ;
      RECT 62.495 10.105 62.67 10.595 ;
      RECT 62.495 7.305 62.665 10.595 ;
      RECT 62.495 9.605 62.905 9.935 ;
      RECT 62.495 8.765 62.905 9.095 ;
      RECT 62.495 7.305 62.67 8.565 ;
      RECT 59.8 3.13 59.97 3.4 ;
      RECT 59.8 3.13 60.53 3.3 ;
      RECT 59.72 4.52 60.05 4.69 ;
      RECT 58.96 4.35 59.97 4.52 ;
      RECT 58.96 3.87 59.13 4.52 ;
      RECT 59.08 3.79 59.25 4.12 ;
      RECT 58.24 4.52 58.57 4.69 ;
      RECT 56.32 4.52 57.61 4.69 ;
      RECT 57.36 4.435 58.49 4.605 ;
      RECT 58.08 3.51 58.49 3.68 ;
      RECT 58.32 3.05 58.49 3.68 ;
      RECT 58.265 10.045 58.44 10.595 ;
      RECT 58.265 7.305 58.435 10.595 ;
      RECT 58.265 7.305 58.44 8.445 ;
      RECT 57.835 7.305 58.005 9.515 ;
      RECT 57.835 7.305 58.01 8.565 ;
      RECT 56.88 10.105 57.055 10.595 ;
      RECT 56.88 7.305 57.05 10.595 ;
      RECT 56.88 9.605 57.29 9.935 ;
      RECT 56.88 8.765 57.29 9.095 ;
      RECT 56.88 7.305 57.055 8.565 ;
      RECT 55.56 3.87 56.89 4.04 ;
      RECT 56.64 3.79 56.81 4.04 ;
      RECT 55.64 3.47 55.81 3.68 ;
      RECT 55.64 3.47 56.13 3.64 ;
      RECT 54.32 4.63 54.61 4.8 ;
      RECT 54.32 3.87 54.49 4.8 ;
      RECT 54.12 3.87 54.49 4.04 ;
      RECT 53.12 3.87 53.61 4.04 ;
      RECT 53.44 3.79 53.61 4.04 ;
      RECT 53.2 4.63 53.61 4.8 ;
      RECT 53.44 4.44 53.61 4.8 ;
      RECT 52.24 4.35 52.89 4.52 ;
      RECT 52.24 3.79 52.41 4.52 ;
      RECT 51.88 4.91 52.17 5.08 ;
      RECT 51.88 3.87 52.05 5.08 ;
      RECT 51.68 3.87 52.05 4.04 ;
      RECT 49.91 7.3 50.08 8.77 ;
      RECT 49.91 7.3 50.085 8.56 ;
      RECT 49.54 9.25 50.01 9.42 ;
      RECT 49.54 8.23 49.71 9.42 ;
      RECT 49.535 3.04 49.705 4.23 ;
      RECT 49.535 3.04 50.005 3.21 ;
      RECT 48.915 3.895 49.09 5.155 ;
      RECT 48.915 3.685 49.085 5.155 ;
      RECT 48.915 7.305 49.085 8.775 ;
      RECT 48.915 7.305 49.09 8.565 ;
      RECT 48.545 3.035 48.715 4.225 ;
      RECT 48.545 3.035 49.015 3.205 ;
      RECT 48.545 9.255 49.015 9.425 ;
      RECT 48.545 8.235 48.715 9.425 ;
      RECT 47.555 4.015 47.73 5.155 ;
      RECT 47.555 1.865 47.725 5.155 ;
      RECT 47.555 1.865 47.73 2.415 ;
      RECT 47.555 10.045 47.73 10.595 ;
      RECT 47.555 7.305 47.725 10.595 ;
      RECT 47.555 7.305 47.73 8.445 ;
      RECT 47.125 3.895 47.3 5.155 ;
      RECT 47.125 2.945 47.295 5.155 ;
      RECT 47.125 7.305 47.295 9.515 ;
      RECT 47.125 7.305 47.3 8.565 ;
      RECT 46.695 3.925 46.865 5.155 ;
      RECT 46.755 2.145 46.925 4.095 ;
      RECT 46.695 1.865 46.865 2.315 ;
      RECT 46.695 10.145 46.865 10.595 ;
      RECT 46.755 8.365 46.925 10.315 ;
      RECT 46.695 7.305 46.865 8.535 ;
      RECT 46.17 3.895 46.345 5.155 ;
      RECT 46.17 1.865 46.34 5.155 ;
      RECT 46.17 3.365 46.58 3.695 ;
      RECT 46.17 2.525 46.58 2.855 ;
      RECT 46.17 1.865 46.345 2.355 ;
      RECT 46.17 10.105 46.345 10.595 ;
      RECT 46.17 7.305 46.34 10.595 ;
      RECT 46.17 9.605 46.58 9.935 ;
      RECT 46.17 8.765 46.58 9.095 ;
      RECT 46.17 7.305 46.345 8.565 ;
      RECT 43.475 3.13 43.645 3.4 ;
      RECT 43.475 3.13 44.205 3.3 ;
      RECT 43.395 4.52 43.725 4.69 ;
      RECT 42.635 4.35 43.645 4.52 ;
      RECT 42.635 3.87 42.805 4.52 ;
      RECT 42.755 3.79 42.925 4.12 ;
      RECT 41.915 4.52 42.245 4.69 ;
      RECT 39.995 4.52 41.285 4.69 ;
      RECT 41.035 4.435 42.165 4.605 ;
      RECT 41.755 3.51 42.165 3.68 ;
      RECT 41.995 3.05 42.165 3.68 ;
      RECT 41.94 10.045 42.115 10.595 ;
      RECT 41.94 7.305 42.11 10.595 ;
      RECT 41.94 7.305 42.115 8.445 ;
      RECT 41.51 7.305 41.68 9.515 ;
      RECT 41.51 7.305 41.685 8.565 ;
      RECT 40.555 10.105 40.73 10.595 ;
      RECT 40.555 7.305 40.725 10.595 ;
      RECT 40.555 9.605 40.965 9.935 ;
      RECT 40.555 8.765 40.965 9.095 ;
      RECT 40.555 7.305 40.73 8.565 ;
      RECT 39.235 3.87 40.565 4.04 ;
      RECT 40.315 3.79 40.485 4.04 ;
      RECT 39.315 3.47 39.485 3.68 ;
      RECT 39.315 3.47 39.805 3.64 ;
      RECT 37.995 4.63 38.285 4.8 ;
      RECT 37.995 3.87 38.165 4.8 ;
      RECT 37.795 3.87 38.165 4.04 ;
      RECT 36.795 3.87 37.285 4.04 ;
      RECT 37.115 3.79 37.285 4.04 ;
      RECT 36.875 4.63 37.285 4.8 ;
      RECT 37.115 4.44 37.285 4.8 ;
      RECT 35.915 4.35 36.565 4.52 ;
      RECT 35.915 3.79 36.085 4.52 ;
      RECT 35.555 4.91 35.845 5.08 ;
      RECT 35.555 3.87 35.725 5.08 ;
      RECT 35.355 3.87 35.725 4.04 ;
      RECT 33.585 7.3 33.755 8.77 ;
      RECT 33.585 7.3 33.76 8.56 ;
      RECT 33.215 9.25 33.685 9.42 ;
      RECT 33.215 8.23 33.385 9.42 ;
      RECT 33.21 3.04 33.38 4.23 ;
      RECT 33.21 3.04 33.68 3.21 ;
      RECT 32.59 3.895 32.765 5.155 ;
      RECT 32.59 3.685 32.76 5.155 ;
      RECT 32.59 7.305 32.76 8.775 ;
      RECT 32.59 7.305 32.765 8.565 ;
      RECT 32.22 3.035 32.39 4.225 ;
      RECT 32.22 3.035 32.69 3.205 ;
      RECT 32.22 9.255 32.69 9.425 ;
      RECT 32.22 8.235 32.39 9.425 ;
      RECT 31.23 4.015 31.405 5.155 ;
      RECT 31.23 1.865 31.4 5.155 ;
      RECT 31.23 1.865 31.405 2.415 ;
      RECT 31.23 10.045 31.405 10.595 ;
      RECT 31.23 7.305 31.4 10.595 ;
      RECT 31.23 7.305 31.405 8.445 ;
      RECT 30.8 3.895 30.975 5.155 ;
      RECT 30.8 2.945 30.97 5.155 ;
      RECT 30.8 7.305 30.97 9.515 ;
      RECT 30.8 7.305 30.975 8.565 ;
      RECT 30.37 3.925 30.54 5.155 ;
      RECT 30.43 2.145 30.6 4.095 ;
      RECT 30.37 1.865 30.54 2.315 ;
      RECT 30.37 10.145 30.54 10.595 ;
      RECT 30.43 8.365 30.6 10.315 ;
      RECT 30.37 7.305 30.54 8.535 ;
      RECT 29.845 3.895 30.02 5.155 ;
      RECT 29.845 1.865 30.015 5.155 ;
      RECT 29.845 3.365 30.255 3.695 ;
      RECT 29.845 2.525 30.255 2.855 ;
      RECT 29.845 1.865 30.02 2.355 ;
      RECT 29.845 10.105 30.02 10.595 ;
      RECT 29.845 7.305 30.015 10.595 ;
      RECT 29.845 9.605 30.255 9.935 ;
      RECT 29.845 8.765 30.255 9.095 ;
      RECT 29.845 7.305 30.02 8.565 ;
      RECT 27.15 3.13 27.32 3.4 ;
      RECT 27.15 3.13 27.88 3.3 ;
      RECT 27.07 4.52 27.4 4.69 ;
      RECT 26.31 4.35 27.32 4.52 ;
      RECT 26.31 3.87 26.48 4.52 ;
      RECT 26.43 3.79 26.6 4.12 ;
      RECT 25.59 4.52 25.92 4.69 ;
      RECT 23.67 4.52 24.96 4.69 ;
      RECT 24.71 4.435 25.84 4.605 ;
      RECT 25.43 3.51 25.84 3.68 ;
      RECT 25.67 3.05 25.84 3.68 ;
      RECT 25.615 10.045 25.79 10.595 ;
      RECT 25.615 7.305 25.785 10.595 ;
      RECT 25.615 7.305 25.79 8.445 ;
      RECT 25.185 7.305 25.355 9.515 ;
      RECT 25.185 7.305 25.36 8.565 ;
      RECT 24.23 10.105 24.405 10.595 ;
      RECT 24.23 7.305 24.4 10.595 ;
      RECT 24.23 9.605 24.64 9.935 ;
      RECT 24.23 8.765 24.64 9.095 ;
      RECT 24.23 7.305 24.405 8.565 ;
      RECT 22.91 3.87 24.24 4.04 ;
      RECT 23.99 3.79 24.16 4.04 ;
      RECT 22.99 3.47 23.16 3.68 ;
      RECT 22.99 3.47 23.48 3.64 ;
      RECT 21.67 4.63 21.96 4.8 ;
      RECT 21.67 3.87 21.84 4.8 ;
      RECT 21.47 3.87 21.84 4.04 ;
      RECT 20.47 3.87 20.96 4.04 ;
      RECT 20.79 3.79 20.96 4.04 ;
      RECT 20.55 4.63 20.96 4.8 ;
      RECT 20.79 4.44 20.96 4.8 ;
      RECT 19.59 4.35 20.24 4.52 ;
      RECT 19.59 3.79 19.76 4.52 ;
      RECT 19.23 4.91 19.52 5.08 ;
      RECT 19.23 3.87 19.4 5.08 ;
      RECT 19.03 3.87 19.4 4.04 ;
      RECT 16.605 7.305 16.775 9.515 ;
      RECT 16.605 7.305 16.78 8.565 ;
      RECT 16.175 10.145 16.345 10.595 ;
      RECT 16.235 8.365 16.405 10.315 ;
      RECT 16.175 7.305 16.345 8.535 ;
      RECT 15.65 10.105 15.825 10.595 ;
      RECT 15.65 7.305 15.82 10.595 ;
      RECT 15.65 9.605 16.06 9.935 ;
      RECT 15.65 8.765 16.06 9.095 ;
      RECT 15.65 7.305 15.825 8.565 ;
      RECT 98.885 10.08 99.06 10.59 ;
      RECT 97.89 1.865 98.065 2.375 ;
      RECT 97.89 10.085 98.065 10.595 ;
      RECT 96.1 1.865 96.275 2.375 ;
      RECT 96.1 10.085 96.275 10.595 ;
      RECT 92.21 3.79 92.38 4.12 ;
      RECT 91.49 3.05 91.66 3.4 ;
      RECT 91.49 4.78 91.66 5.11 ;
      RECT 90.49 4.78 90.66 5.11 ;
      RECT 90.485 10.085 90.66 10.595 ;
      RECT 90.25 3.79 90.42 4.24 ;
      RECT 89.77 3.79 89.94 4.12 ;
      RECT 89.05 3.05 89.22 3.4 ;
      RECT 88.05 4.44 88.22 4.8 ;
      RECT 87.81 3.79 87.98 4.24 ;
      RECT 87.33 3.79 87.5 4.12 ;
      RECT 87.09 3.05 87.26 3.4 ;
      RECT 86.61 4.35 86.78 4.77 ;
      RECT 85.61 3.05 85.78 3.4 ;
      RECT 85.37 3.79 85.54 4.12 ;
      RECT 84.65 3.05 84.82 3.4 ;
      RECT 84.17 4.35 84.34 4.77 ;
      RECT 82.56 10.08 82.735 10.59 ;
      RECT 81.565 1.865 81.74 2.375 ;
      RECT 81.565 10.085 81.74 10.595 ;
      RECT 79.775 1.865 79.95 2.375 ;
      RECT 79.775 10.085 79.95 10.595 ;
      RECT 75.885 3.79 76.055 4.12 ;
      RECT 75.165 3.05 75.335 3.4 ;
      RECT 75.165 4.78 75.335 5.11 ;
      RECT 74.165 4.78 74.335 5.11 ;
      RECT 74.16 10.085 74.335 10.595 ;
      RECT 73.925 3.79 74.095 4.24 ;
      RECT 73.445 3.79 73.615 4.12 ;
      RECT 72.725 3.05 72.895 3.4 ;
      RECT 71.725 4.44 71.895 4.8 ;
      RECT 71.485 3.79 71.655 4.24 ;
      RECT 71.005 3.79 71.175 4.12 ;
      RECT 70.765 3.05 70.935 3.4 ;
      RECT 70.285 4.35 70.455 4.77 ;
      RECT 69.285 3.05 69.455 3.4 ;
      RECT 69.045 3.79 69.215 4.12 ;
      RECT 68.325 3.05 68.495 3.4 ;
      RECT 67.845 4.35 68.015 4.77 ;
      RECT 66.235 10.08 66.41 10.59 ;
      RECT 65.24 1.865 65.415 2.375 ;
      RECT 65.24 10.085 65.415 10.595 ;
      RECT 63.45 1.865 63.625 2.375 ;
      RECT 63.45 10.085 63.625 10.595 ;
      RECT 59.56 3.79 59.73 4.12 ;
      RECT 58.84 3.05 59.01 3.4 ;
      RECT 58.84 4.78 59.01 5.11 ;
      RECT 57.84 4.78 58.01 5.11 ;
      RECT 57.835 10.085 58.01 10.595 ;
      RECT 57.6 3.79 57.77 4.24 ;
      RECT 57.12 3.79 57.29 4.12 ;
      RECT 56.4 3.05 56.57 3.4 ;
      RECT 55.4 4.44 55.57 4.8 ;
      RECT 55.16 3.79 55.33 4.24 ;
      RECT 54.68 3.79 54.85 4.12 ;
      RECT 54.44 3.05 54.61 3.4 ;
      RECT 53.96 4.35 54.13 4.77 ;
      RECT 52.96 3.05 53.13 3.4 ;
      RECT 52.72 3.79 52.89 4.12 ;
      RECT 52 3.05 52.17 3.4 ;
      RECT 51.52 4.35 51.69 4.77 ;
      RECT 49.91 10.08 50.085 10.59 ;
      RECT 48.915 1.865 49.09 2.375 ;
      RECT 48.915 10.085 49.09 10.595 ;
      RECT 47.125 1.865 47.3 2.375 ;
      RECT 47.125 10.085 47.3 10.595 ;
      RECT 43.235 3.79 43.405 4.12 ;
      RECT 42.515 3.05 42.685 3.4 ;
      RECT 42.515 4.78 42.685 5.11 ;
      RECT 41.515 4.78 41.685 5.11 ;
      RECT 41.51 10.085 41.685 10.595 ;
      RECT 41.275 3.79 41.445 4.24 ;
      RECT 40.795 3.79 40.965 4.12 ;
      RECT 40.075 3.05 40.245 3.4 ;
      RECT 39.075 4.44 39.245 4.8 ;
      RECT 38.835 3.79 39.005 4.24 ;
      RECT 38.355 3.79 38.525 4.12 ;
      RECT 38.115 3.05 38.285 3.4 ;
      RECT 37.635 4.35 37.805 4.77 ;
      RECT 36.635 3.05 36.805 3.4 ;
      RECT 36.395 3.79 36.565 4.12 ;
      RECT 35.675 3.05 35.845 3.4 ;
      RECT 35.195 4.35 35.365 4.77 ;
      RECT 33.585 10.08 33.76 10.59 ;
      RECT 32.59 1.865 32.765 2.375 ;
      RECT 32.59 10.085 32.765 10.595 ;
      RECT 30.8 1.865 30.975 2.375 ;
      RECT 30.8 10.085 30.975 10.595 ;
      RECT 26.91 3.79 27.08 4.12 ;
      RECT 26.19 3.05 26.36 3.4 ;
      RECT 26.19 4.78 26.36 5.11 ;
      RECT 25.19 4.78 25.36 5.11 ;
      RECT 25.185 10.085 25.36 10.595 ;
      RECT 24.95 3.79 25.12 4.24 ;
      RECT 24.47 3.79 24.64 4.12 ;
      RECT 23.75 3.05 23.92 3.4 ;
      RECT 22.75 4.44 22.92 4.8 ;
      RECT 22.51 3.79 22.68 4.24 ;
      RECT 22.03 3.79 22.2 4.12 ;
      RECT 21.79 3.05 21.96 3.4 ;
      RECT 21.31 4.35 21.48 4.77 ;
      RECT 20.31 3.05 20.48 3.4 ;
      RECT 20.07 3.79 20.24 4.12 ;
      RECT 19.35 3.05 19.52 3.4 ;
      RECT 18.87 4.35 19.04 4.77 ;
      RECT 16.605 10.085 16.78 10.595 ;
  END
END sky130_osu_ring_oscillator_mpr2ea_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2ea_8_b0r2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ea_8_b0r2 ;
  SIZE 99.425 BY 12.46 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.47965 ;
    PORT
      LAYER li1 ;
        RECT 33.575 1.87 33.75 2.38 ;
        RECT 33.575 3.9 33.75 5.16 ;
        RECT 33.575 3.69 33.745 5.16 ;
      LAYER met1 ;
        RECT 33.515 2.18 33.81 2.41 ;
        RECT 33.515 3.66 33.805 3.89 ;
        RECT 33.575 2.18 33.745 3.89 ;
      LAYER mcon ;
        RECT 33.575 3.69 33.745 3.86 ;
        RECT 33.575 2.21 33.745 2.38 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.47965 ;
    PORT
      LAYER li1 ;
        RECT 49.9 1.87 50.075 2.38 ;
        RECT 49.9 3.9 50.075 5.16 ;
        RECT 49.9 3.69 50.07 5.16 ;
      LAYER met1 ;
        RECT 49.84 2.18 50.135 2.41 ;
        RECT 49.84 3.66 50.13 3.89 ;
        RECT 49.9 2.18 50.07 3.89 ;
      LAYER mcon ;
        RECT 49.9 3.69 50.07 3.86 ;
        RECT 49.9 2.21 50.07 2.38 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.47965 ;
    PORT
      LAYER li1 ;
        RECT 66.225 1.87 66.4 2.38 ;
        RECT 66.225 3.9 66.4 5.16 ;
        RECT 66.225 3.69 66.395 5.16 ;
      LAYER met1 ;
        RECT 66.165 2.18 66.46 2.41 ;
        RECT 66.165 3.66 66.455 3.89 ;
        RECT 66.225 2.18 66.395 3.89 ;
      LAYER mcon ;
        RECT 66.225 3.69 66.395 3.86 ;
        RECT 66.225 2.21 66.395 2.38 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.47965 ;
    PORT
      LAYER li1 ;
        RECT 82.55 1.87 82.725 2.38 ;
        RECT 82.55 3.9 82.725 5.16 ;
        RECT 82.55 3.69 82.72 5.16 ;
      LAYER met1 ;
        RECT 82.49 2.18 82.785 2.41 ;
        RECT 82.49 3.66 82.78 3.89 ;
        RECT 82.55 2.18 82.72 3.89 ;
      LAYER mcon ;
        RECT 82.55 3.69 82.72 3.86 ;
        RECT 82.55 2.21 82.72 2.38 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.47965 ;
    PORT
      LAYER li1 ;
        RECT 98.875 1.87 99.05 2.38 ;
        RECT 98.875 3.9 99.05 5.16 ;
        RECT 98.875 3.69 99.045 5.16 ;
      LAYER met1 ;
        RECT 98.815 2.18 99.11 2.41 ;
        RECT 98.815 3.66 99.105 3.89 ;
        RECT 98.875 2.18 99.045 3.89 ;
      LAYER mcon ;
        RECT 98.875 3.69 99.045 3.86 ;
        RECT 98.875 2.21 99.045 2.38 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 29.35 4 29.69 4.35 ;
        RECT 29.34 8.125 29.68 8.475 ;
        RECT 29.425 4 29.595 8.475 ;
      LAYER li1 ;
        RECT 29.42 2.955 29.59 4.225 ;
        RECT 29.42 8.235 29.59 9.505 ;
        RECT 23.805 8.235 23.975 9.505 ;
      LAYER met1 ;
        RECT 29.35 4.055 29.82 4.225 ;
        RECT 29.35 4 29.69 4.35 ;
        RECT 29.34 8.235 29.82 8.405 ;
        RECT 29.34 8.125 29.68 8.475 ;
        RECT 23.745 8.23 29.68 8.4 ;
        RECT 23.745 8.23 24.205 8.405 ;
        RECT 23.745 8.205 24.035 8.435 ;
      LAYER via1 ;
        RECT 29.44 8.225 29.59 8.375 ;
        RECT 29.45 4.1 29.6 4.25 ;
      LAYER mcon ;
        RECT 23.805 8.235 23.975 8.405 ;
        RECT 29.42 8.235 29.59 8.405 ;
        RECT 29.42 4.055 29.59 4.225 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 45.675 4 46.015 4.35 ;
        RECT 45.665 8.125 46.005 8.475 ;
        RECT 45.75 4 45.92 8.475 ;
      LAYER li1 ;
        RECT 45.745 2.955 45.915 4.225 ;
        RECT 45.745 8.235 45.915 9.505 ;
        RECT 40.13 8.235 40.3 9.505 ;
      LAYER met1 ;
        RECT 45.675 4.055 46.145 4.225 ;
        RECT 45.675 4 46.015 4.35 ;
        RECT 45.665 8.235 46.145 8.405 ;
        RECT 45.665 8.125 46.005 8.475 ;
        RECT 40.07 8.23 46.005 8.4 ;
        RECT 40.07 8.23 40.53 8.405 ;
        RECT 40.07 8.205 40.36 8.435 ;
      LAYER via1 ;
        RECT 45.765 8.225 45.915 8.375 ;
        RECT 45.775 4.1 45.925 4.25 ;
      LAYER mcon ;
        RECT 40.13 8.235 40.3 8.405 ;
        RECT 45.745 8.235 45.915 8.405 ;
        RECT 45.745 4.055 45.915 4.225 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 62 4 62.34 4.35 ;
        RECT 61.99 8.125 62.33 8.475 ;
        RECT 62.075 4 62.245 8.475 ;
      LAYER li1 ;
        RECT 62.07 2.955 62.24 4.225 ;
        RECT 62.07 8.235 62.24 9.505 ;
        RECT 56.455 8.235 56.625 9.505 ;
      LAYER met1 ;
        RECT 62 4.055 62.47 4.225 ;
        RECT 62 4 62.34 4.35 ;
        RECT 61.99 8.235 62.47 8.405 ;
        RECT 61.99 8.125 62.33 8.475 ;
        RECT 56.395 8.23 62.33 8.4 ;
        RECT 56.395 8.23 56.855 8.405 ;
        RECT 56.395 8.205 56.685 8.435 ;
      LAYER via1 ;
        RECT 62.09 8.225 62.24 8.375 ;
        RECT 62.1 4.1 62.25 4.25 ;
      LAYER mcon ;
        RECT 56.455 8.235 56.625 8.405 ;
        RECT 62.07 8.235 62.24 8.405 ;
        RECT 62.07 4.055 62.24 4.225 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 78.325 4 78.665 4.35 ;
        RECT 78.315 8.125 78.655 8.475 ;
        RECT 78.4 4 78.57 8.475 ;
      LAYER li1 ;
        RECT 78.395 2.955 78.565 4.225 ;
        RECT 78.395 8.235 78.565 9.505 ;
        RECT 72.78 8.235 72.95 9.505 ;
      LAYER met1 ;
        RECT 78.325 4.055 78.795 4.225 ;
        RECT 78.325 4 78.665 4.35 ;
        RECT 78.315 8.235 78.795 8.405 ;
        RECT 78.315 8.125 78.655 8.475 ;
        RECT 72.72 8.23 78.655 8.4 ;
        RECT 72.72 8.23 73.18 8.405 ;
        RECT 72.72 8.205 73.01 8.435 ;
      LAYER via1 ;
        RECT 78.415 8.225 78.565 8.375 ;
        RECT 78.425 4.1 78.575 4.25 ;
      LAYER mcon ;
        RECT 72.78 8.235 72.95 8.405 ;
        RECT 78.395 8.235 78.565 8.405 ;
        RECT 78.395 4.055 78.565 4.225 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 94.65 4 94.99 4.35 ;
        RECT 94.64 8.125 94.98 8.475 ;
        RECT 94.725 4 94.895 8.475 ;
      LAYER li1 ;
        RECT 94.72 2.955 94.89 4.225 ;
        RECT 94.72 8.235 94.89 9.505 ;
        RECT 89.105 8.235 89.275 9.505 ;
      LAYER met1 ;
        RECT 94.65 4.055 95.12 4.225 ;
        RECT 94.65 4 94.99 4.35 ;
        RECT 94.64 8.235 95.12 8.405 ;
        RECT 94.64 8.125 94.98 8.475 ;
        RECT 89.045 8.23 94.98 8.4 ;
        RECT 89.045 8.23 89.505 8.405 ;
        RECT 89.045 8.205 89.335 8.435 ;
      LAYER via1 ;
        RECT 94.74 8.225 94.89 8.375 ;
        RECT 94.75 4.1 94.9 4.25 ;
      LAYER mcon ;
        RECT 89.105 8.235 89.275 8.405 ;
        RECT 94.72 8.235 94.89 8.405 ;
        RECT 94.72 4.055 94.89 4.225 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 15.225 8.235 15.395 9.505 ;
      LAYER met1 ;
        RECT 15.165 8.235 15.625 8.405 ;
        RECT 15.17 8.2 15.46 8.43 ;
        RECT 15.165 8.205 15.455 8.435 ;
      LAYER mcon ;
        RECT 15.225 8.235 15.395 8.405 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 5.435 99.42 7.035 ;
        RECT 17.79 5.43 99.42 7.035 ;
        RECT 98.45 5.43 98.62 7.76 ;
        RECT 98.445 4.7 98.615 7.035 ;
        RECT 94.54 5.425 98.275 7.035 ;
        RECT 97.455 4.695 97.625 7.765 ;
        RECT 94.71 4.695 94.88 7.765 ;
        RECT 83.835 5.33 93.495 7.035 ;
        RECT 92.925 4.83 93.095 7.035 ;
        RECT 91.965 4.83 92.135 7.035 ;
        RECT 89.525 4.83 89.695 7.035 ;
        RECT 89.095 5.33 89.265 7.765 ;
        RECT 88.525 4.83 88.695 7.035 ;
        RECT 87.565 4.83 87.735 7.035 ;
        RECT 85.125 4.83 85.295 7.035 ;
        RECT 82.125 5.43 82.295 7.76 ;
        RECT 82.12 4.7 82.29 7.035 ;
        RECT 78.215 5.425 81.95 7.035 ;
        RECT 81.13 4.695 81.3 7.765 ;
        RECT 78.385 4.695 78.555 7.765 ;
        RECT 67.51 5.33 77.17 7.035 ;
        RECT 76.6 4.83 76.77 7.035 ;
        RECT 75.64 4.83 75.81 7.035 ;
        RECT 73.2 4.83 73.37 7.035 ;
        RECT 72.77 5.33 72.94 7.765 ;
        RECT 72.2 4.83 72.37 7.035 ;
        RECT 71.24 4.83 71.41 7.035 ;
        RECT 68.8 4.83 68.97 7.035 ;
        RECT 65.8 5.43 65.97 7.76 ;
        RECT 65.795 4.7 65.965 7.035 ;
        RECT 61.89 5.425 65.625 7.035 ;
        RECT 64.805 4.695 64.975 7.765 ;
        RECT 62.06 4.695 62.23 7.765 ;
        RECT 51.185 5.33 60.845 7.035 ;
        RECT 60.275 4.83 60.445 7.035 ;
        RECT 59.315 4.83 59.485 7.035 ;
        RECT 56.875 4.83 57.045 7.035 ;
        RECT 56.445 5.33 56.615 7.765 ;
        RECT 55.875 4.83 56.045 7.035 ;
        RECT 54.915 4.83 55.085 7.035 ;
        RECT 52.475 4.83 52.645 7.035 ;
        RECT 49.475 5.43 49.645 7.76 ;
        RECT 49.47 4.7 49.64 7.035 ;
        RECT 45.565 5.425 49.3 7.035 ;
        RECT 48.48 4.695 48.65 7.765 ;
        RECT 45.735 4.695 45.905 7.765 ;
        RECT 34.86 5.33 44.52 7.035 ;
        RECT 43.95 4.83 44.12 7.035 ;
        RECT 42.99 4.83 43.16 7.035 ;
        RECT 40.55 4.83 40.72 7.035 ;
        RECT 40.12 5.33 40.29 7.765 ;
        RECT 39.55 4.83 39.72 7.035 ;
        RECT 38.59 4.83 38.76 7.035 ;
        RECT 36.15 4.83 36.32 7.035 ;
        RECT 33.15 5.43 33.32 7.76 ;
        RECT 33.145 4.7 33.315 7.035 ;
        RECT 29.24 5.425 32.975 7.035 ;
        RECT 32.155 4.695 32.325 7.765 ;
        RECT 29.41 4.695 29.58 7.765 ;
        RECT 18.535 5.33 28.195 7.035 ;
        RECT 27.625 4.83 27.795 7.035 ;
        RECT 26.665 4.83 26.835 7.035 ;
        RECT 24.225 4.83 24.395 7.035 ;
        RECT 23.795 5.33 23.965 7.765 ;
        RECT 23.225 4.83 23.395 7.035 ;
        RECT 22.265 4.83 22.435 7.035 ;
        RECT 19.825 4.83 19.995 7.035 ;
        RECT 17.03 10.045 17.205 10.595 ;
        RECT 17.03 7.305 17.205 8.445 ;
        RECT 17.03 5.435 17.2 10.595 ;
        RECT 15.215 5.435 15.385 7.765 ;
      LAYER met1 ;
        RECT 0 5.435 99.42 7.035 ;
        RECT 17.79 5.43 99.42 7.035 ;
        RECT 94.54 5.425 98.275 7.035 ;
        RECT 83.835 5.3 93.495 7.035 ;
        RECT 78.215 5.425 81.95 7.035 ;
        RECT 67.51 5.3 77.17 7.035 ;
        RECT 61.89 5.425 65.625 7.035 ;
        RECT 51.185 5.3 60.845 7.035 ;
        RECT 45.565 5.425 49.3 7.035 ;
        RECT 34.86 5.3 44.52 7.035 ;
        RECT 29.24 5.425 32.975 7.035 ;
        RECT 18.535 5.3 28.195 7.035 ;
        RECT 16.97 8.945 17.26 9.175 ;
        RECT 16.8 8.975 17.26 9.145 ;
      LAYER mcon ;
        RECT 17.03 8.975 17.2 9.145 ;
        RECT 17.335 6.835 17.505 7.005 ;
        RECT 18.68 5.33 18.85 5.5 ;
        RECT 19.14 5.33 19.31 5.5 ;
        RECT 19.6 5.33 19.77 5.5 ;
        RECT 20.06 5.33 20.23 5.5 ;
        RECT 20.52 5.33 20.69 5.5 ;
        RECT 20.98 5.33 21.15 5.5 ;
        RECT 21.44 5.33 21.61 5.5 ;
        RECT 21.9 5.33 22.07 5.5 ;
        RECT 22.36 5.33 22.53 5.5 ;
        RECT 22.82 5.33 22.99 5.5 ;
        RECT 23.28 5.33 23.45 5.5 ;
        RECT 23.74 5.33 23.91 5.5 ;
        RECT 24.2 5.33 24.37 5.5 ;
        RECT 24.66 5.33 24.83 5.5 ;
        RECT 25.12 5.33 25.29 5.5 ;
        RECT 25.58 5.33 25.75 5.5 ;
        RECT 25.915 6.835 26.085 7.005 ;
        RECT 26.04 5.33 26.21 5.5 ;
        RECT 26.5 5.33 26.67 5.5 ;
        RECT 26.96 5.33 27.13 5.5 ;
        RECT 27.42 5.33 27.59 5.5 ;
        RECT 27.88 5.33 28.05 5.5 ;
        RECT 31.53 6.835 31.7 7.005 ;
        RECT 31.53 5.455 31.7 5.625 ;
        RECT 32.235 6.835 32.405 7.005 ;
        RECT 32.235 5.455 32.405 5.625 ;
        RECT 33.225 5.46 33.395 5.63 ;
        RECT 33.23 6.83 33.4 7 ;
        RECT 35.005 5.33 35.175 5.5 ;
        RECT 35.465 5.33 35.635 5.5 ;
        RECT 35.925 5.33 36.095 5.5 ;
        RECT 36.385 5.33 36.555 5.5 ;
        RECT 36.845 5.33 37.015 5.5 ;
        RECT 37.305 5.33 37.475 5.5 ;
        RECT 37.765 5.33 37.935 5.5 ;
        RECT 38.225 5.33 38.395 5.5 ;
        RECT 38.685 5.33 38.855 5.5 ;
        RECT 39.145 5.33 39.315 5.5 ;
        RECT 39.605 5.33 39.775 5.5 ;
        RECT 40.065 5.33 40.235 5.5 ;
        RECT 40.525 5.33 40.695 5.5 ;
        RECT 40.985 5.33 41.155 5.5 ;
        RECT 41.445 5.33 41.615 5.5 ;
        RECT 41.905 5.33 42.075 5.5 ;
        RECT 42.24 6.835 42.41 7.005 ;
        RECT 42.365 5.33 42.535 5.5 ;
        RECT 42.825 5.33 42.995 5.5 ;
        RECT 43.285 5.33 43.455 5.5 ;
        RECT 43.745 5.33 43.915 5.5 ;
        RECT 44.205 5.33 44.375 5.5 ;
        RECT 47.855 6.835 48.025 7.005 ;
        RECT 47.855 5.455 48.025 5.625 ;
        RECT 48.56 6.835 48.73 7.005 ;
        RECT 48.56 5.455 48.73 5.625 ;
        RECT 49.55 5.46 49.72 5.63 ;
        RECT 49.555 6.83 49.725 7 ;
        RECT 51.33 5.33 51.5 5.5 ;
        RECT 51.79 5.33 51.96 5.5 ;
        RECT 52.25 5.33 52.42 5.5 ;
        RECT 52.71 5.33 52.88 5.5 ;
        RECT 53.17 5.33 53.34 5.5 ;
        RECT 53.63 5.33 53.8 5.5 ;
        RECT 54.09 5.33 54.26 5.5 ;
        RECT 54.55 5.33 54.72 5.5 ;
        RECT 55.01 5.33 55.18 5.5 ;
        RECT 55.47 5.33 55.64 5.5 ;
        RECT 55.93 5.33 56.1 5.5 ;
        RECT 56.39 5.33 56.56 5.5 ;
        RECT 56.85 5.33 57.02 5.5 ;
        RECT 57.31 5.33 57.48 5.5 ;
        RECT 57.77 5.33 57.94 5.5 ;
        RECT 58.23 5.33 58.4 5.5 ;
        RECT 58.565 6.835 58.735 7.005 ;
        RECT 58.69 5.33 58.86 5.5 ;
        RECT 59.15 5.33 59.32 5.5 ;
        RECT 59.61 5.33 59.78 5.5 ;
        RECT 60.07 5.33 60.24 5.5 ;
        RECT 60.53 5.33 60.7 5.5 ;
        RECT 64.18 6.835 64.35 7.005 ;
        RECT 64.18 5.455 64.35 5.625 ;
        RECT 64.885 6.835 65.055 7.005 ;
        RECT 64.885 5.455 65.055 5.625 ;
        RECT 65.875 5.46 66.045 5.63 ;
        RECT 65.88 6.83 66.05 7 ;
        RECT 67.655 5.33 67.825 5.5 ;
        RECT 68.115 5.33 68.285 5.5 ;
        RECT 68.575 5.33 68.745 5.5 ;
        RECT 69.035 5.33 69.205 5.5 ;
        RECT 69.495 5.33 69.665 5.5 ;
        RECT 69.955 5.33 70.125 5.5 ;
        RECT 70.415 5.33 70.585 5.5 ;
        RECT 70.875 5.33 71.045 5.5 ;
        RECT 71.335 5.33 71.505 5.5 ;
        RECT 71.795 5.33 71.965 5.5 ;
        RECT 72.255 5.33 72.425 5.5 ;
        RECT 72.715 5.33 72.885 5.5 ;
        RECT 73.175 5.33 73.345 5.5 ;
        RECT 73.635 5.33 73.805 5.5 ;
        RECT 74.095 5.33 74.265 5.5 ;
        RECT 74.555 5.33 74.725 5.5 ;
        RECT 74.89 6.835 75.06 7.005 ;
        RECT 75.015 5.33 75.185 5.5 ;
        RECT 75.475 5.33 75.645 5.5 ;
        RECT 75.935 5.33 76.105 5.5 ;
        RECT 76.395 5.33 76.565 5.5 ;
        RECT 76.855 5.33 77.025 5.5 ;
        RECT 80.505 6.835 80.675 7.005 ;
        RECT 80.505 5.455 80.675 5.625 ;
        RECT 81.21 6.835 81.38 7.005 ;
        RECT 81.21 5.455 81.38 5.625 ;
        RECT 82.2 5.46 82.37 5.63 ;
        RECT 82.205 6.83 82.375 7 ;
        RECT 83.98 5.33 84.15 5.5 ;
        RECT 84.44 5.33 84.61 5.5 ;
        RECT 84.9 5.33 85.07 5.5 ;
        RECT 85.36 5.33 85.53 5.5 ;
        RECT 85.82 5.33 85.99 5.5 ;
        RECT 86.28 5.33 86.45 5.5 ;
        RECT 86.74 5.33 86.91 5.5 ;
        RECT 87.2 5.33 87.37 5.5 ;
        RECT 87.66 5.33 87.83 5.5 ;
        RECT 88.12 5.33 88.29 5.5 ;
        RECT 88.58 5.33 88.75 5.5 ;
        RECT 89.04 5.33 89.21 5.5 ;
        RECT 89.5 5.33 89.67 5.5 ;
        RECT 89.96 5.33 90.13 5.5 ;
        RECT 90.42 5.33 90.59 5.5 ;
        RECT 90.88 5.33 91.05 5.5 ;
        RECT 91.215 6.835 91.385 7.005 ;
        RECT 91.34 5.33 91.51 5.5 ;
        RECT 91.8 5.33 91.97 5.5 ;
        RECT 92.26 5.33 92.43 5.5 ;
        RECT 92.72 5.33 92.89 5.5 ;
        RECT 93.18 5.33 93.35 5.5 ;
        RECT 96.83 6.835 97 7.005 ;
        RECT 96.83 5.455 97 5.625 ;
        RECT 97.535 6.835 97.705 7.005 ;
        RECT 97.535 5.455 97.705 5.625 ;
        RECT 98.525 5.46 98.695 5.63 ;
        RECT 98.53 6.83 98.7 7 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 92.725 4.17 93.055 4.9 ;
        RECT 76.4 4.17 76.73 4.9 ;
        RECT 60.075 4.17 60.405 4.9 ;
        RECT 43.75 4.17 44.08 4.9 ;
        RECT 27.425 4.17 27.755 4.9 ;
      LAYER met2 ;
        RECT 92.75 4.15 93.03 4.52 ;
        RECT 92.76 3.895 93.02 4.52 ;
        RECT 76.425 4.15 76.705 4.52 ;
        RECT 76.435 3.895 76.695 4.52 ;
        RECT 60.1 4.15 60.38 4.52 ;
        RECT 60.11 3.895 60.37 4.52 ;
        RECT 43.775 4.15 44.055 4.52 ;
        RECT 43.785 3.895 44.045 4.52 ;
        RECT 27.45 4.15 27.73 4.52 ;
        RECT 27.46 3.895 27.72 4.52 ;
      LAYER li1 ;
        RECT 0 10.86 99.425 12.46 ;
        RECT 98.45 10.23 98.62 12.46 ;
        RECT 97.455 10.235 97.625 12.46 ;
        RECT 94.71 10.235 94.88 12.46 ;
        RECT 89.095 10.235 89.265 12.46 ;
        RECT 82.125 10.23 82.295 12.46 ;
        RECT 81.13 10.235 81.3 12.46 ;
        RECT 78.385 10.235 78.555 12.46 ;
        RECT 72.77 10.235 72.94 12.46 ;
        RECT 65.8 10.23 65.97 12.46 ;
        RECT 64.805 10.235 64.975 12.46 ;
        RECT 62.06 10.235 62.23 12.46 ;
        RECT 56.445 10.235 56.615 12.46 ;
        RECT 49.475 10.23 49.645 12.46 ;
        RECT 48.48 10.235 48.65 12.46 ;
        RECT 45.735 10.235 45.905 12.46 ;
        RECT 40.12 10.235 40.29 12.46 ;
        RECT 33.15 10.23 33.32 12.46 ;
        RECT 32.155 10.235 32.325 12.46 ;
        RECT 29.41 10.235 29.58 12.46 ;
        RECT 23.795 10.235 23.965 12.46 ;
        RECT 15.215 10.235 15.385 12.46 ;
        RECT 0 0 99.42 1.6 ;
        RECT 98.445 0 98.615 2.23 ;
        RECT 97.455 0 97.625 2.225 ;
        RECT 94.71 0 94.88 2.225 ;
        RECT 93.46 0 93.65 2.88 ;
        RECT 93.455 0 93.65 2.86 ;
        RECT 83.835 0 93.65 2.78 ;
        RECT 91.965 0 92.135 3.28 ;
        RECT 90.005 0 90.175 3.28 ;
        RECT 89.935 0 90.175 2.89 ;
        RECT 88.095 0 88.29 2.86 ;
        RECT 87.565 0 87.735 3.28 ;
        RECT 86.605 0 86.775 3.28 ;
        RECT 86.085 0 86.255 3.28 ;
        RECT 85.125 0 85.295 3.28 ;
        RECT 84.165 0 84.335 3.28 ;
        RECT 82.12 0 82.29 2.23 ;
        RECT 81.13 0 81.3 2.225 ;
        RECT 78.385 0 78.555 2.225 ;
        RECT 77.135 0 77.325 2.88 ;
        RECT 77.13 0 77.325 2.86 ;
        RECT 67.51 0 77.325 2.78 ;
        RECT 75.64 0 75.81 3.28 ;
        RECT 73.68 0 73.85 3.28 ;
        RECT 73.61 0 73.85 2.89 ;
        RECT 71.77 0 71.965 2.86 ;
        RECT 71.24 0 71.41 3.28 ;
        RECT 70.28 0 70.45 3.28 ;
        RECT 69.76 0 69.93 3.28 ;
        RECT 68.8 0 68.97 3.28 ;
        RECT 67.84 0 68.01 3.28 ;
        RECT 65.795 0 65.965 2.23 ;
        RECT 64.805 0 64.975 2.225 ;
        RECT 62.06 0 62.23 2.225 ;
        RECT 60.81 0 61 2.88 ;
        RECT 60.805 0 61 2.86 ;
        RECT 51.185 0 61 2.78 ;
        RECT 59.315 0 59.485 3.28 ;
        RECT 57.355 0 57.525 3.28 ;
        RECT 57.285 0 57.525 2.89 ;
        RECT 55.445 0 55.64 2.86 ;
        RECT 54.915 0 55.085 3.28 ;
        RECT 53.955 0 54.125 3.28 ;
        RECT 53.435 0 53.605 3.28 ;
        RECT 52.475 0 52.645 3.28 ;
        RECT 51.515 0 51.685 3.28 ;
        RECT 49.47 0 49.64 2.23 ;
        RECT 48.48 0 48.65 2.225 ;
        RECT 45.735 0 45.905 2.225 ;
        RECT 44.485 0 44.675 2.88 ;
        RECT 44.48 0 44.675 2.86 ;
        RECT 34.86 0 44.675 2.78 ;
        RECT 42.99 0 43.16 3.28 ;
        RECT 41.03 0 41.2 3.28 ;
        RECT 40.96 0 41.2 2.89 ;
        RECT 39.12 0 39.315 2.86 ;
        RECT 38.59 0 38.76 3.28 ;
        RECT 37.63 0 37.8 3.28 ;
        RECT 37.11 0 37.28 3.28 ;
        RECT 36.15 0 36.32 3.28 ;
        RECT 35.19 0 35.36 3.28 ;
        RECT 33.145 0 33.315 2.23 ;
        RECT 32.155 0 32.325 2.225 ;
        RECT 29.41 0 29.58 2.225 ;
        RECT 28.16 0 28.35 2.88 ;
        RECT 28.155 0 28.35 2.86 ;
        RECT 18.535 0 28.35 2.78 ;
        RECT 26.665 0 26.835 3.28 ;
        RECT 24.705 0 24.875 3.28 ;
        RECT 24.635 0 24.875 2.89 ;
        RECT 22.795 0 22.99 2.86 ;
        RECT 22.265 0 22.435 3.28 ;
        RECT 21.305 0 21.475 3.28 ;
        RECT 20.785 0 20.955 3.28 ;
        RECT 19.825 0 19.995 3.28 ;
        RECT 18.865 0 19.035 3.28 ;
        RECT 92.925 3.77 93.095 4.14 ;
        RECT 92.605 3.77 93.095 3.94 ;
        RECT 90.965 3.77 91.135 4.14 ;
        RECT 90.645 3.77 91.135 3.94 ;
        RECT 90.11 8.365 90.28 10.315 ;
        RECT 90.05 10.145 90.22 10.595 ;
        RECT 90.05 7.305 90.22 8.535 ;
        RECT 76.6 3.77 76.77 4.14 ;
        RECT 76.28 3.77 76.77 3.94 ;
        RECT 74.64 3.77 74.81 4.14 ;
        RECT 74.32 3.77 74.81 3.94 ;
        RECT 73.785 8.365 73.955 10.315 ;
        RECT 73.725 10.145 73.895 10.595 ;
        RECT 73.725 7.305 73.895 8.535 ;
        RECT 60.275 3.77 60.445 4.14 ;
        RECT 59.955 3.77 60.445 3.94 ;
        RECT 58.315 3.77 58.485 4.14 ;
        RECT 57.995 3.77 58.485 3.94 ;
        RECT 57.46 8.365 57.63 10.315 ;
        RECT 57.4 10.145 57.57 10.595 ;
        RECT 57.4 7.305 57.57 8.535 ;
        RECT 43.95 3.77 44.12 4.14 ;
        RECT 43.63 3.77 44.12 3.94 ;
        RECT 41.99 3.77 42.16 4.14 ;
        RECT 41.67 3.77 42.16 3.94 ;
        RECT 41.135 8.365 41.305 10.315 ;
        RECT 41.075 10.145 41.245 10.595 ;
        RECT 41.075 7.305 41.245 8.535 ;
        RECT 27.625 3.77 27.795 4.14 ;
        RECT 27.305 3.77 27.795 3.94 ;
        RECT 25.665 3.77 25.835 4.14 ;
        RECT 25.345 3.77 25.835 3.94 ;
        RECT 24.81 8.365 24.98 10.315 ;
        RECT 24.75 10.145 24.92 10.595 ;
        RECT 24.75 7.305 24.92 8.535 ;
      LAYER met1 ;
        RECT 0 10.86 99.425 12.46 ;
        RECT 90.05 8.575 90.34 8.805 ;
        RECT 89.67 8.6 90.34 8.775 ;
        RECT 89.67 8.6 89.845 12.46 ;
        RECT 73.725 8.575 74.015 8.805 ;
        RECT 73.345 8.6 74.015 8.775 ;
        RECT 73.345 8.6 73.52 12.46 ;
        RECT 57.4 8.575 57.69 8.805 ;
        RECT 57.02 8.6 57.69 8.775 ;
        RECT 57.02 8.6 57.195 12.46 ;
        RECT 41.075 8.575 41.365 8.805 ;
        RECT 40.695 8.6 41.365 8.775 ;
        RECT 40.695 8.6 40.87 12.46 ;
        RECT 24.75 8.575 25.04 8.805 ;
        RECT 24.37 8.6 25.04 8.775 ;
        RECT 24.37 8.6 24.545 12.46 ;
        RECT 0 0 99.42 1.6 ;
        RECT 93.465 0 93.65 4.24 ;
        RECT 92.7 4.055 93.65 4.24 ;
        RECT 93.46 0 93.65 2.88 ;
        RECT 93.455 0 93.65 2.86 ;
        RECT 83.835 0 93.65 2.81 ;
        RECT 92.7 3.985 93.155 4.24 ;
        RECT 92.73 3.94 93.155 4.24 ;
        RECT 92.73 3.925 93.05 4.24 ;
        RECT 92.765 3.925 93.005 4.35 ;
        RECT 91.24 4.125 93.005 4.265 ;
        RECT 90.905 3.985 91.38 4.17 ;
        RECT 90.905 3.94 91.195 4.17 ;
        RECT 89.935 0 90.13 2.89 ;
        RECT 88.095 0 88.29 2.86 ;
        RECT 86.26 0 86.455 2.89 ;
        RECT 83.96 0 84.155 2.89 ;
        RECT 77.14 0 77.325 4.24 ;
        RECT 76.375 4.055 77.325 4.24 ;
        RECT 77.135 0 77.325 2.88 ;
        RECT 77.13 0 77.325 2.86 ;
        RECT 67.51 0 77.325 2.81 ;
        RECT 76.375 3.985 76.83 4.24 ;
        RECT 76.405 3.94 76.83 4.24 ;
        RECT 76.405 3.925 76.725 4.24 ;
        RECT 76.44 3.925 76.68 4.35 ;
        RECT 74.915 4.125 76.68 4.265 ;
        RECT 74.58 3.985 75.055 4.17 ;
        RECT 74.58 3.94 74.87 4.17 ;
        RECT 73.61 0 73.805 2.89 ;
        RECT 71.77 0 71.965 2.86 ;
        RECT 69.935 0 70.13 2.89 ;
        RECT 67.635 0 67.83 2.89 ;
        RECT 60.815 0 61 4.24 ;
        RECT 60.05 4.055 61 4.24 ;
        RECT 60.81 0 61 2.88 ;
        RECT 60.805 0 61 2.86 ;
        RECT 51.185 0 61 2.81 ;
        RECT 60.05 3.985 60.505 4.24 ;
        RECT 60.08 3.94 60.505 4.24 ;
        RECT 60.08 3.925 60.4 4.24 ;
        RECT 60.115 3.925 60.355 4.35 ;
        RECT 58.59 4.125 60.355 4.265 ;
        RECT 58.255 3.985 58.73 4.17 ;
        RECT 58.255 3.94 58.545 4.17 ;
        RECT 57.285 0 57.48 2.89 ;
        RECT 55.445 0 55.64 2.86 ;
        RECT 53.61 0 53.805 2.89 ;
        RECT 51.31 0 51.505 2.89 ;
        RECT 44.49 0 44.675 4.24 ;
        RECT 43.725 4.055 44.675 4.24 ;
        RECT 44.485 0 44.675 2.88 ;
        RECT 44.48 0 44.675 2.86 ;
        RECT 34.86 0 44.675 2.81 ;
        RECT 43.725 3.985 44.18 4.24 ;
        RECT 43.755 3.94 44.18 4.24 ;
        RECT 43.755 3.925 44.075 4.24 ;
        RECT 43.79 3.925 44.03 4.35 ;
        RECT 42.265 4.125 44.03 4.265 ;
        RECT 41.93 3.985 42.405 4.17 ;
        RECT 41.93 3.94 42.22 4.17 ;
        RECT 40.96 0 41.155 2.89 ;
        RECT 39.12 0 39.315 2.86 ;
        RECT 37.285 0 37.48 2.89 ;
        RECT 34.985 0 35.18 2.89 ;
        RECT 28.165 0 28.35 4.24 ;
        RECT 27.4 4.055 28.35 4.24 ;
        RECT 28.16 0 28.35 2.88 ;
        RECT 28.155 0 28.35 2.86 ;
        RECT 18.535 0 28.35 2.81 ;
        RECT 27.4 3.985 27.855 4.24 ;
        RECT 27.43 3.94 27.855 4.24 ;
        RECT 27.43 3.925 27.75 4.24 ;
        RECT 27.465 3.925 27.705 4.35 ;
        RECT 25.94 4.125 27.705 4.265 ;
        RECT 25.605 3.985 26.08 4.17 ;
        RECT 25.605 3.94 25.895 4.17 ;
        RECT 24.635 0 24.83 2.89 ;
        RECT 22.795 0 22.99 2.86 ;
        RECT 20.96 0 21.155 2.89 ;
        RECT 18.66 0 18.855 2.89 ;
      LAYER via1 ;
        RECT 27.515 3.98 27.665 4.13 ;
        RECT 43.84 3.98 43.99 4.13 ;
        RECT 60.165 3.98 60.315 4.13 ;
        RECT 76.49 3.98 76.64 4.13 ;
        RECT 92.815 3.98 92.965 4.13 ;
      LAYER via2 ;
        RECT 27.49 4.235 27.69 4.435 ;
        RECT 43.815 4.235 44.015 4.435 ;
        RECT 60.14 4.235 60.34 4.435 ;
        RECT 76.465 4.235 76.665 4.435 ;
        RECT 92.79 4.235 92.99 4.435 ;
      LAYER mcon ;
        RECT 15.295 10.895 15.465 11.065 ;
        RECT 15.975 10.895 16.145 11.065 ;
        RECT 16.655 10.895 16.825 11.065 ;
        RECT 17.335 10.895 17.505 11.065 ;
        RECT 18.68 2.61 18.85 2.78 ;
        RECT 19.14 2.61 19.31 2.78 ;
        RECT 19.6 2.61 19.77 2.78 ;
        RECT 20.06 2.61 20.23 2.78 ;
        RECT 20.52 2.61 20.69 2.78 ;
        RECT 20.98 2.61 21.15 2.78 ;
        RECT 21.44 2.61 21.61 2.78 ;
        RECT 21.9 2.61 22.07 2.78 ;
        RECT 22.36 2.61 22.53 2.78 ;
        RECT 22.82 2.61 22.99 2.78 ;
        RECT 23.28 2.61 23.45 2.78 ;
        RECT 23.74 2.61 23.91 2.78 ;
        RECT 23.875 10.895 24.045 11.065 ;
        RECT 24.2 2.61 24.37 2.78 ;
        RECT 24.555 10.895 24.725 11.065 ;
        RECT 24.66 2.61 24.83 2.78 ;
        RECT 24.81 8.605 24.98 8.775 ;
        RECT 25.12 2.61 25.29 2.78 ;
        RECT 25.235 10.895 25.405 11.065 ;
        RECT 25.58 2.61 25.75 2.78 ;
        RECT 25.665 3.97 25.835 4.14 ;
        RECT 25.915 10.895 26.085 11.065 ;
        RECT 26.04 2.61 26.21 2.78 ;
        RECT 26.5 2.61 26.67 2.78 ;
        RECT 26.96 2.61 27.13 2.78 ;
        RECT 27.42 2.61 27.59 2.78 ;
        RECT 27.625 3.97 27.795 4.14 ;
        RECT 27.88 2.61 28.05 2.78 ;
        RECT 29.49 10.895 29.66 11.065 ;
        RECT 29.49 1.395 29.66 1.565 ;
        RECT 30.17 10.895 30.34 11.065 ;
        RECT 30.17 1.395 30.34 1.565 ;
        RECT 30.85 10.895 31.02 11.065 ;
        RECT 30.85 1.395 31.02 1.565 ;
        RECT 31.53 10.895 31.7 11.065 ;
        RECT 31.53 1.395 31.7 1.565 ;
        RECT 32.235 10.895 32.405 11.065 ;
        RECT 32.235 1.395 32.405 1.565 ;
        RECT 33.225 1.4 33.395 1.57 ;
        RECT 33.23 10.89 33.4 11.06 ;
        RECT 35.005 2.61 35.175 2.78 ;
        RECT 35.465 2.61 35.635 2.78 ;
        RECT 35.925 2.61 36.095 2.78 ;
        RECT 36.385 2.61 36.555 2.78 ;
        RECT 36.845 2.61 37.015 2.78 ;
        RECT 37.305 2.61 37.475 2.78 ;
        RECT 37.765 2.61 37.935 2.78 ;
        RECT 38.225 2.61 38.395 2.78 ;
        RECT 38.685 2.61 38.855 2.78 ;
        RECT 39.145 2.61 39.315 2.78 ;
        RECT 39.605 2.61 39.775 2.78 ;
        RECT 40.065 2.61 40.235 2.78 ;
        RECT 40.2 10.895 40.37 11.065 ;
        RECT 40.525 2.61 40.695 2.78 ;
        RECT 40.88 10.895 41.05 11.065 ;
        RECT 40.985 2.61 41.155 2.78 ;
        RECT 41.135 8.605 41.305 8.775 ;
        RECT 41.445 2.61 41.615 2.78 ;
        RECT 41.56 10.895 41.73 11.065 ;
        RECT 41.905 2.61 42.075 2.78 ;
        RECT 41.99 3.97 42.16 4.14 ;
        RECT 42.24 10.895 42.41 11.065 ;
        RECT 42.365 2.61 42.535 2.78 ;
        RECT 42.825 2.61 42.995 2.78 ;
        RECT 43.285 2.61 43.455 2.78 ;
        RECT 43.745 2.61 43.915 2.78 ;
        RECT 43.95 3.97 44.12 4.14 ;
        RECT 44.205 2.61 44.375 2.78 ;
        RECT 45.815 10.895 45.985 11.065 ;
        RECT 45.815 1.395 45.985 1.565 ;
        RECT 46.495 10.895 46.665 11.065 ;
        RECT 46.495 1.395 46.665 1.565 ;
        RECT 47.175 10.895 47.345 11.065 ;
        RECT 47.175 1.395 47.345 1.565 ;
        RECT 47.855 10.895 48.025 11.065 ;
        RECT 47.855 1.395 48.025 1.565 ;
        RECT 48.56 10.895 48.73 11.065 ;
        RECT 48.56 1.395 48.73 1.565 ;
        RECT 49.55 1.4 49.72 1.57 ;
        RECT 49.555 10.89 49.725 11.06 ;
        RECT 51.33 2.61 51.5 2.78 ;
        RECT 51.79 2.61 51.96 2.78 ;
        RECT 52.25 2.61 52.42 2.78 ;
        RECT 52.71 2.61 52.88 2.78 ;
        RECT 53.17 2.61 53.34 2.78 ;
        RECT 53.63 2.61 53.8 2.78 ;
        RECT 54.09 2.61 54.26 2.78 ;
        RECT 54.55 2.61 54.72 2.78 ;
        RECT 55.01 2.61 55.18 2.78 ;
        RECT 55.47 2.61 55.64 2.78 ;
        RECT 55.93 2.61 56.1 2.78 ;
        RECT 56.39 2.61 56.56 2.78 ;
        RECT 56.525 10.895 56.695 11.065 ;
        RECT 56.85 2.61 57.02 2.78 ;
        RECT 57.205 10.895 57.375 11.065 ;
        RECT 57.31 2.61 57.48 2.78 ;
        RECT 57.46 8.605 57.63 8.775 ;
        RECT 57.77 2.61 57.94 2.78 ;
        RECT 57.885 10.895 58.055 11.065 ;
        RECT 58.23 2.61 58.4 2.78 ;
        RECT 58.315 3.97 58.485 4.14 ;
        RECT 58.565 10.895 58.735 11.065 ;
        RECT 58.69 2.61 58.86 2.78 ;
        RECT 59.15 2.61 59.32 2.78 ;
        RECT 59.61 2.61 59.78 2.78 ;
        RECT 60.07 2.61 60.24 2.78 ;
        RECT 60.275 3.97 60.445 4.14 ;
        RECT 60.53 2.61 60.7 2.78 ;
        RECT 62.14 10.895 62.31 11.065 ;
        RECT 62.14 1.395 62.31 1.565 ;
        RECT 62.82 10.895 62.99 11.065 ;
        RECT 62.82 1.395 62.99 1.565 ;
        RECT 63.5 10.895 63.67 11.065 ;
        RECT 63.5 1.395 63.67 1.565 ;
        RECT 64.18 10.895 64.35 11.065 ;
        RECT 64.18 1.395 64.35 1.565 ;
        RECT 64.885 10.895 65.055 11.065 ;
        RECT 64.885 1.395 65.055 1.565 ;
        RECT 65.875 1.4 66.045 1.57 ;
        RECT 65.88 10.89 66.05 11.06 ;
        RECT 67.655 2.61 67.825 2.78 ;
        RECT 68.115 2.61 68.285 2.78 ;
        RECT 68.575 2.61 68.745 2.78 ;
        RECT 69.035 2.61 69.205 2.78 ;
        RECT 69.495 2.61 69.665 2.78 ;
        RECT 69.955 2.61 70.125 2.78 ;
        RECT 70.415 2.61 70.585 2.78 ;
        RECT 70.875 2.61 71.045 2.78 ;
        RECT 71.335 2.61 71.505 2.78 ;
        RECT 71.795 2.61 71.965 2.78 ;
        RECT 72.255 2.61 72.425 2.78 ;
        RECT 72.715 2.61 72.885 2.78 ;
        RECT 72.85 10.895 73.02 11.065 ;
        RECT 73.175 2.61 73.345 2.78 ;
        RECT 73.53 10.895 73.7 11.065 ;
        RECT 73.635 2.61 73.805 2.78 ;
        RECT 73.785 8.605 73.955 8.775 ;
        RECT 74.095 2.61 74.265 2.78 ;
        RECT 74.21 10.895 74.38 11.065 ;
        RECT 74.555 2.61 74.725 2.78 ;
        RECT 74.64 3.97 74.81 4.14 ;
        RECT 74.89 10.895 75.06 11.065 ;
        RECT 75.015 2.61 75.185 2.78 ;
        RECT 75.475 2.61 75.645 2.78 ;
        RECT 75.935 2.61 76.105 2.78 ;
        RECT 76.395 2.61 76.565 2.78 ;
        RECT 76.6 3.97 76.77 4.14 ;
        RECT 76.855 2.61 77.025 2.78 ;
        RECT 78.465 10.895 78.635 11.065 ;
        RECT 78.465 1.395 78.635 1.565 ;
        RECT 79.145 10.895 79.315 11.065 ;
        RECT 79.145 1.395 79.315 1.565 ;
        RECT 79.825 10.895 79.995 11.065 ;
        RECT 79.825 1.395 79.995 1.565 ;
        RECT 80.505 10.895 80.675 11.065 ;
        RECT 80.505 1.395 80.675 1.565 ;
        RECT 81.21 10.895 81.38 11.065 ;
        RECT 81.21 1.395 81.38 1.565 ;
        RECT 82.2 1.4 82.37 1.57 ;
        RECT 82.205 10.89 82.375 11.06 ;
        RECT 83.98 2.61 84.15 2.78 ;
        RECT 84.44 2.61 84.61 2.78 ;
        RECT 84.9 2.61 85.07 2.78 ;
        RECT 85.36 2.61 85.53 2.78 ;
        RECT 85.82 2.61 85.99 2.78 ;
        RECT 86.28 2.61 86.45 2.78 ;
        RECT 86.74 2.61 86.91 2.78 ;
        RECT 87.2 2.61 87.37 2.78 ;
        RECT 87.66 2.61 87.83 2.78 ;
        RECT 88.12 2.61 88.29 2.78 ;
        RECT 88.58 2.61 88.75 2.78 ;
        RECT 89.04 2.61 89.21 2.78 ;
        RECT 89.175 10.895 89.345 11.065 ;
        RECT 89.5 2.61 89.67 2.78 ;
        RECT 89.855 10.895 90.025 11.065 ;
        RECT 89.96 2.61 90.13 2.78 ;
        RECT 90.11 8.605 90.28 8.775 ;
        RECT 90.42 2.61 90.59 2.78 ;
        RECT 90.535 10.895 90.705 11.065 ;
        RECT 90.88 2.61 91.05 2.78 ;
        RECT 90.965 3.97 91.135 4.14 ;
        RECT 91.215 10.895 91.385 11.065 ;
        RECT 91.34 2.61 91.51 2.78 ;
        RECT 91.8 2.61 91.97 2.78 ;
        RECT 92.26 2.61 92.43 2.78 ;
        RECT 92.72 2.61 92.89 2.78 ;
        RECT 92.925 3.97 93.095 4.14 ;
        RECT 93.18 2.61 93.35 2.78 ;
        RECT 94.79 10.895 94.96 11.065 ;
        RECT 94.79 1.395 94.96 1.565 ;
        RECT 95.47 10.895 95.64 11.065 ;
        RECT 95.47 1.395 95.64 1.565 ;
        RECT 96.15 10.895 96.32 11.065 ;
        RECT 96.15 1.395 96.32 1.565 ;
        RECT 96.83 10.895 97 11.065 ;
        RECT 96.83 1.395 97 1.565 ;
        RECT 97.535 10.895 97.705 11.065 ;
        RECT 97.535 1.395 97.705 1.565 ;
        RECT 98.525 1.4 98.695 1.57 ;
        RECT 98.53 10.89 98.7 11.06 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 90.4 9.34 90.77 9.71 ;
      RECT 90.4 9.375 92.385 9.675 ;
      RECT 92.085 3.575 92.385 9.675 ;
      RECT 89.085 3.21 89.415 3.94 ;
      RECT 88.205 3.21 88.535 3.94 ;
      RECT 91.285 3.575 92.575 3.875 ;
      RECT 92.245 3.045 92.575 3.875 ;
      RECT 88.205 3.575 90.345 3.875 ;
      RECT 90.045 3.16 90.345 3.875 ;
      RECT 91.285 3.16 91.59 3.875 ;
      RECT 90.045 3.16 91.59 3.47 ;
      RECT 88.705 4.73 89.035 5.06 ;
      RECT 87.5 4.745 89.035 5.045 ;
      RECT 87.5 3.625 87.8 5.045 ;
      RECT 87.245 3.61 87.575 3.94 ;
      RECT 74.075 9.34 74.445 9.71 ;
      RECT 74.075 9.375 76.06 9.675 ;
      RECT 75.76 3.575 76.06 9.675 ;
      RECT 72.76 3.21 73.09 3.94 ;
      RECT 71.88 3.21 72.21 3.94 ;
      RECT 74.96 3.575 76.25 3.875 ;
      RECT 75.92 3.045 76.25 3.875 ;
      RECT 71.88 3.575 74.02 3.875 ;
      RECT 73.72 3.16 74.02 3.875 ;
      RECT 74.96 3.16 75.265 3.875 ;
      RECT 73.72 3.16 75.265 3.47 ;
      RECT 72.38 4.73 72.71 5.06 ;
      RECT 71.175 4.745 72.71 5.045 ;
      RECT 71.175 3.625 71.475 5.045 ;
      RECT 70.92 3.61 71.25 3.94 ;
      RECT 57.75 9.34 58.12 9.71 ;
      RECT 57.75 9.375 59.735 9.675 ;
      RECT 59.435 3.575 59.735 9.675 ;
      RECT 56.435 3.21 56.765 3.94 ;
      RECT 55.555 3.21 55.885 3.94 ;
      RECT 58.635 3.575 59.925 3.875 ;
      RECT 59.595 3.045 59.925 3.875 ;
      RECT 55.555 3.575 57.695 3.875 ;
      RECT 57.395 3.16 57.695 3.875 ;
      RECT 58.635 3.16 58.94 3.875 ;
      RECT 57.395 3.16 58.94 3.47 ;
      RECT 56.055 4.73 56.385 5.06 ;
      RECT 54.85 4.745 56.385 5.045 ;
      RECT 54.85 3.625 55.15 5.045 ;
      RECT 54.595 3.61 54.925 3.94 ;
      RECT 41.425 9.34 41.795 9.71 ;
      RECT 41.425 9.375 43.41 9.675 ;
      RECT 43.11 3.575 43.41 9.675 ;
      RECT 40.11 3.21 40.44 3.94 ;
      RECT 39.23 3.21 39.56 3.94 ;
      RECT 42.31 3.575 43.6 3.875 ;
      RECT 43.27 3.045 43.6 3.875 ;
      RECT 39.23 3.575 41.37 3.875 ;
      RECT 41.07 3.16 41.37 3.875 ;
      RECT 42.31 3.16 42.615 3.875 ;
      RECT 41.07 3.16 42.615 3.47 ;
      RECT 39.73 4.73 40.06 5.06 ;
      RECT 38.525 4.745 40.06 5.045 ;
      RECT 38.525 3.625 38.825 5.045 ;
      RECT 38.27 3.61 38.6 3.94 ;
      RECT 25.1 9.34 25.47 9.71 ;
      RECT 25.1 9.375 27.085 9.675 ;
      RECT 26.785 3.575 27.085 9.675 ;
      RECT 23.785 3.21 24.115 3.94 ;
      RECT 22.905 3.21 23.235 3.94 ;
      RECT 25.985 3.575 27.275 3.875 ;
      RECT 26.945 3.045 27.275 3.875 ;
      RECT 22.905 3.575 25.045 3.875 ;
      RECT 24.745 3.16 25.045 3.875 ;
      RECT 25.985 3.16 26.29 3.875 ;
      RECT 24.745 3.16 26.29 3.47 ;
      RECT 23.405 4.73 23.735 5.06 ;
      RECT 22.2 4.745 23.735 5.045 ;
      RECT 22.2 3.625 22.5 5.045 ;
      RECT 21.945 3.61 22.275 3.94 ;
      RECT 90.645 3.77 90.975 4.5 ;
      RECT 86.525 3.61 86.855 4.34 ;
      RECT 85.525 3.05 85.855 3.78 ;
      RECT 84.085 3.77 84.415 4.5 ;
      RECT 74.32 3.77 74.65 4.5 ;
      RECT 70.2 3.61 70.53 4.34 ;
      RECT 69.2 3.05 69.53 3.78 ;
      RECT 67.76 3.77 68.09 4.5 ;
      RECT 57.995 3.77 58.325 4.5 ;
      RECT 53.875 3.61 54.205 4.34 ;
      RECT 52.875 3.05 53.205 3.78 ;
      RECT 51.435 3.77 51.765 4.5 ;
      RECT 41.67 3.77 42 4.5 ;
      RECT 37.55 3.61 37.88 4.34 ;
      RECT 36.55 3.05 36.88 3.78 ;
      RECT 35.11 3.77 35.44 4.5 ;
      RECT 25.345 3.77 25.675 4.5 ;
      RECT 21.225 3.61 21.555 4.34 ;
      RECT 20.225 3.05 20.555 3.78 ;
      RECT 18.785 3.77 19.115 4.5 ;
    LAYER via2 ;
      RECT 92.31 3.51 92.51 3.71 ;
      RECT 90.71 4.235 90.91 4.435 ;
      RECT 90.485 9.425 90.685 9.625 ;
      RECT 89.15 3.675 89.35 3.875 ;
      RECT 88.77 4.795 88.97 4.995 ;
      RECT 88.27 3.675 88.47 3.875 ;
      RECT 87.31 3.675 87.51 3.875 ;
      RECT 86.59 3.675 86.79 3.875 ;
      RECT 85.59 3.115 85.79 3.315 ;
      RECT 84.15 4.235 84.35 4.435 ;
      RECT 75.985 3.51 76.185 3.71 ;
      RECT 74.385 4.235 74.585 4.435 ;
      RECT 74.16 9.425 74.36 9.625 ;
      RECT 72.825 3.675 73.025 3.875 ;
      RECT 72.445 4.795 72.645 4.995 ;
      RECT 71.945 3.675 72.145 3.875 ;
      RECT 70.985 3.675 71.185 3.875 ;
      RECT 70.265 3.675 70.465 3.875 ;
      RECT 69.265 3.115 69.465 3.315 ;
      RECT 67.825 4.235 68.025 4.435 ;
      RECT 59.66 3.51 59.86 3.71 ;
      RECT 58.06 4.235 58.26 4.435 ;
      RECT 57.835 9.425 58.035 9.625 ;
      RECT 56.5 3.675 56.7 3.875 ;
      RECT 56.12 4.795 56.32 4.995 ;
      RECT 55.62 3.675 55.82 3.875 ;
      RECT 54.66 3.675 54.86 3.875 ;
      RECT 53.94 3.675 54.14 3.875 ;
      RECT 52.94 3.115 53.14 3.315 ;
      RECT 51.5 4.235 51.7 4.435 ;
      RECT 43.335 3.51 43.535 3.71 ;
      RECT 41.735 4.235 41.935 4.435 ;
      RECT 41.51 9.425 41.71 9.625 ;
      RECT 40.175 3.675 40.375 3.875 ;
      RECT 39.795 4.795 39.995 4.995 ;
      RECT 39.295 3.675 39.495 3.875 ;
      RECT 38.335 3.675 38.535 3.875 ;
      RECT 37.615 3.675 37.815 3.875 ;
      RECT 36.615 3.115 36.815 3.315 ;
      RECT 35.175 4.235 35.375 4.435 ;
      RECT 27.01 3.51 27.21 3.71 ;
      RECT 25.41 4.235 25.61 4.435 ;
      RECT 25.185 9.425 25.385 9.625 ;
      RECT 23.85 3.675 24.05 3.875 ;
      RECT 23.47 4.795 23.67 4.995 ;
      RECT 22.97 3.675 23.17 3.875 ;
      RECT 22.01 3.675 22.21 3.875 ;
      RECT 21.29 3.675 21.49 3.875 ;
      RECT 20.29 3.115 20.49 3.315 ;
      RECT 18.85 4.235 19.05 4.435 ;
    LAYER met2 ;
      RECT 16.225 10.685 99.05 10.855 ;
      RECT 98.88 9.56 99.05 10.855 ;
      RECT 16.225 8.54 16.395 10.855 ;
      RECT 98.85 9.56 99.2 9.91 ;
      RECT 16.165 8.54 16.455 8.89 ;
      RECT 95.69 8.505 96.01 8.83 ;
      RECT 95.72 7.98 95.89 8.83 ;
      RECT 95.72 7.98 95.895 8.33 ;
      RECT 95.72 7.98 96.695 8.155 ;
      RECT 96.52 3.26 96.695 8.155 ;
      RECT 96.465 3.26 96.815 3.61 ;
      RECT 96.49 8.94 96.815 9.265 ;
      RECT 95.375 9.03 96.815 9.2 ;
      RECT 95.375 3.69 95.535 9.2 ;
      RECT 95.69 3.66 96.01 3.98 ;
      RECT 95.375 3.69 96.01 3.86 ;
      RECT 84.11 4.15 84.39 4.52 ;
      RECT 84.165 2.355 84.335 4.52 ;
      RECT 94.16 2.35 94.33 3.11 ;
      RECT 94.07 2.755 94.41 3.105 ;
      RECT 94.07 2.355 94.33 3.105 ;
      RECT 94.105 2.35 94.33 3.105 ;
      RECT 84.165 2.355 94.33 2.515 ;
      RECT 90.79 3.59 91.07 3.96 ;
      RECT 89.72 3.615 89.98 3.935 ;
      RECT 92.27 3.425 92.55 3.795 ;
      RECT 92.88 3.335 93.14 3.655 ;
      RECT 89.78 2.775 89.92 3.935 ;
      RECT 90.86 2.775 91 3.96 ;
      RECT 91.98 3.425 93.14 3.565 ;
      RECT 91.98 2.775 92.12 3.565 ;
      RECT 89.78 2.775 92.12 2.915 ;
      RECT 89.81 4.915 91.985 5.08 ;
      RECT 91.84 3.795 91.985 5.08 ;
      RECT 88.73 4.71 89.01 5.08 ;
      RECT 88.73 4.825 89.95 4.965 ;
      RECT 91.56 3.795 91.985 3.935 ;
      RECT 91.56 3.615 91.82 3.935 ;
      RECT 84.9 5.195 88.56 5.335 ;
      RECT 88.42 4.38 88.56 5.335 ;
      RECT 84.9 4.265 85.04 5.335 ;
      RECT 91.44 4.455 91.7 4.775 ;
      RECT 88.42 4.38 90.95 4.52 ;
      RECT 90.67 4.15 90.95 4.52 ;
      RECT 84.9 4.265 85.35 4.52 ;
      RECT 85.07 4.15 85.35 4.52 ;
      RECT 91.44 4.265 91.64 4.775 ;
      RECT 90.67 4.265 91.64 4.405 ;
      RECT 91.24 3.055 91.38 4.405 ;
      RECT 91.18 3.055 91.44 3.375 ;
      RECT 82.5 8.94 82.85 9.29 ;
      RECT 91.055 8.895 91.405 9.245 ;
      RECT 82.5 8.97 91.405 9.17 ;
      RECT 85.08 3.615 85.34 3.935 ;
      RECT 85.08 3.705 86.12 3.845 ;
      RECT 85.98 2.915 86.12 3.845 ;
      RECT 88.74 3.055 89 3.375 ;
      RECT 85.98 2.915 88.94 3.055 ;
      RECT 88.12 3.895 88.38 4.215 ;
      RECT 88.12 3.895 88.44 4.125 ;
      RECT 88.23 3.59 88.51 3.96 ;
      RECT 87.82 4.455 88.14 4.775 ;
      RECT 87.82 3.335 87.96 4.775 ;
      RECT 87.76 3.335 88.02 3.655 ;
      RECT 85.32 4.735 85.58 5.055 ;
      RECT 85.32 4.825 87 4.965 ;
      RECT 86.86 4.545 87 4.965 ;
      RECT 86.86 4.545 87.3 4.775 ;
      RECT 87.04 4.455 87.3 4.775 ;
      RECT 86.36 3.615 86.76 4.125 ;
      RECT 86.55 3.59 86.83 3.96 ;
      RECT 86.3 3.615 86.83 3.935 ;
      RECT 79.365 8.505 79.685 8.83 ;
      RECT 79.395 7.98 79.565 8.83 ;
      RECT 79.395 7.98 79.57 8.33 ;
      RECT 79.395 7.98 80.37 8.155 ;
      RECT 80.195 3.26 80.37 8.155 ;
      RECT 80.14 3.26 80.49 3.61 ;
      RECT 80.165 8.94 80.49 9.265 ;
      RECT 79.05 9.03 80.49 9.2 ;
      RECT 79.05 3.69 79.21 9.2 ;
      RECT 79.365 3.66 79.685 3.98 ;
      RECT 79.05 3.69 79.685 3.86 ;
      RECT 67.785 4.15 68.065 4.52 ;
      RECT 67.84 2.355 68.01 4.52 ;
      RECT 77.835 2.35 78.005 3.11 ;
      RECT 77.745 2.755 78.085 3.105 ;
      RECT 77.745 2.355 78.005 3.105 ;
      RECT 77.78 2.35 78.005 3.105 ;
      RECT 67.84 2.355 78.005 2.515 ;
      RECT 74.465 3.59 74.745 3.96 ;
      RECT 73.395 3.615 73.655 3.935 ;
      RECT 75.945 3.425 76.225 3.795 ;
      RECT 76.555 3.335 76.815 3.655 ;
      RECT 73.455 2.775 73.595 3.935 ;
      RECT 74.535 2.775 74.675 3.96 ;
      RECT 75.655 3.425 76.815 3.565 ;
      RECT 75.655 2.775 75.795 3.565 ;
      RECT 73.455 2.775 75.795 2.915 ;
      RECT 73.485 4.915 75.66 5.08 ;
      RECT 75.515 3.795 75.66 5.08 ;
      RECT 72.405 4.71 72.685 5.08 ;
      RECT 72.405 4.825 73.625 4.965 ;
      RECT 75.235 3.795 75.66 3.935 ;
      RECT 75.235 3.615 75.495 3.935 ;
      RECT 68.575 5.195 72.235 5.335 ;
      RECT 72.095 4.38 72.235 5.335 ;
      RECT 68.575 4.265 68.715 5.335 ;
      RECT 75.115 4.455 75.375 4.775 ;
      RECT 72.095 4.38 74.625 4.52 ;
      RECT 74.345 4.15 74.625 4.52 ;
      RECT 68.575 4.265 69.025 4.52 ;
      RECT 68.745 4.15 69.025 4.52 ;
      RECT 75.115 4.265 75.315 4.775 ;
      RECT 74.345 4.265 75.315 4.405 ;
      RECT 74.915 3.055 75.055 4.405 ;
      RECT 74.855 3.055 75.115 3.375 ;
      RECT 66.175 8.94 66.525 9.29 ;
      RECT 74.725 8.895 75.075 9.245 ;
      RECT 66.175 8.97 75.075 9.17 ;
      RECT 68.755 3.615 69.015 3.935 ;
      RECT 68.755 3.705 69.795 3.845 ;
      RECT 69.655 2.915 69.795 3.845 ;
      RECT 72.415 3.055 72.675 3.375 ;
      RECT 69.655 2.915 72.615 3.055 ;
      RECT 71.795 3.895 72.055 4.215 ;
      RECT 71.795 3.895 72.115 4.125 ;
      RECT 71.905 3.59 72.185 3.96 ;
      RECT 71.495 4.455 71.815 4.775 ;
      RECT 71.495 3.335 71.635 4.775 ;
      RECT 71.435 3.335 71.695 3.655 ;
      RECT 68.995 4.735 69.255 5.055 ;
      RECT 68.995 4.825 70.675 4.965 ;
      RECT 70.535 4.545 70.675 4.965 ;
      RECT 70.535 4.545 70.975 4.775 ;
      RECT 70.715 4.455 70.975 4.775 ;
      RECT 70.035 3.615 70.435 4.125 ;
      RECT 70.225 3.59 70.505 3.96 ;
      RECT 69.975 3.615 70.505 3.935 ;
      RECT 63.04 8.505 63.36 8.83 ;
      RECT 63.07 7.98 63.24 8.83 ;
      RECT 63.07 7.98 63.245 8.33 ;
      RECT 63.07 7.98 64.045 8.155 ;
      RECT 63.87 3.26 64.045 8.155 ;
      RECT 63.815 3.26 64.165 3.61 ;
      RECT 63.84 8.94 64.165 9.265 ;
      RECT 62.725 9.03 64.165 9.2 ;
      RECT 62.725 3.69 62.885 9.2 ;
      RECT 63.04 3.66 63.36 3.98 ;
      RECT 62.725 3.69 63.36 3.86 ;
      RECT 51.46 4.15 51.74 4.52 ;
      RECT 51.515 2.355 51.685 4.52 ;
      RECT 61.51 2.35 61.68 3.11 ;
      RECT 61.42 2.755 61.76 3.105 ;
      RECT 61.42 2.355 61.68 3.105 ;
      RECT 61.455 2.35 61.68 3.105 ;
      RECT 51.515 2.355 61.68 2.515 ;
      RECT 58.14 3.59 58.42 3.96 ;
      RECT 57.07 3.615 57.33 3.935 ;
      RECT 59.62 3.425 59.9 3.795 ;
      RECT 60.23 3.335 60.49 3.655 ;
      RECT 57.13 2.775 57.27 3.935 ;
      RECT 58.21 2.775 58.35 3.96 ;
      RECT 59.33 3.425 60.49 3.565 ;
      RECT 59.33 2.775 59.47 3.565 ;
      RECT 57.13 2.775 59.47 2.915 ;
      RECT 57.16 4.915 59.335 5.08 ;
      RECT 59.19 3.795 59.335 5.08 ;
      RECT 56.08 4.71 56.36 5.08 ;
      RECT 56.08 4.825 57.3 4.965 ;
      RECT 58.91 3.795 59.335 3.935 ;
      RECT 58.91 3.615 59.17 3.935 ;
      RECT 52.25 5.195 55.91 5.335 ;
      RECT 55.77 4.38 55.91 5.335 ;
      RECT 52.25 4.265 52.39 5.335 ;
      RECT 58.79 4.455 59.05 4.775 ;
      RECT 55.77 4.38 58.3 4.52 ;
      RECT 58.02 4.15 58.3 4.52 ;
      RECT 52.25 4.265 52.7 4.52 ;
      RECT 52.42 4.15 52.7 4.52 ;
      RECT 58.79 4.265 58.99 4.775 ;
      RECT 58.02 4.265 58.99 4.405 ;
      RECT 58.59 3.055 58.73 4.405 ;
      RECT 58.53 3.055 58.79 3.375 ;
      RECT 49.895 8.945 50.245 9.295 ;
      RECT 58.4 8.9 58.75 9.25 ;
      RECT 49.895 8.975 58.75 9.175 ;
      RECT 52.43 3.615 52.69 3.935 ;
      RECT 52.43 3.705 53.47 3.845 ;
      RECT 53.33 2.915 53.47 3.845 ;
      RECT 56.09 3.055 56.35 3.375 ;
      RECT 53.33 2.915 56.29 3.055 ;
      RECT 55.47 3.895 55.73 4.215 ;
      RECT 55.47 3.895 55.79 4.125 ;
      RECT 55.58 3.59 55.86 3.96 ;
      RECT 55.17 4.455 55.49 4.775 ;
      RECT 55.17 3.335 55.31 4.775 ;
      RECT 55.11 3.335 55.37 3.655 ;
      RECT 52.67 4.735 52.93 5.055 ;
      RECT 52.67 4.825 54.35 4.965 ;
      RECT 54.21 4.545 54.35 4.965 ;
      RECT 54.21 4.545 54.65 4.775 ;
      RECT 54.39 4.455 54.65 4.775 ;
      RECT 53.71 3.615 54.11 4.125 ;
      RECT 53.9 3.59 54.18 3.96 ;
      RECT 53.65 3.615 54.18 3.935 ;
      RECT 46.715 8.505 47.035 8.83 ;
      RECT 46.745 7.98 46.915 8.83 ;
      RECT 46.745 7.98 46.92 8.33 ;
      RECT 46.745 7.98 47.72 8.155 ;
      RECT 47.545 3.26 47.72 8.155 ;
      RECT 47.49 3.26 47.84 3.61 ;
      RECT 47.515 8.94 47.84 9.265 ;
      RECT 46.4 9.03 47.84 9.2 ;
      RECT 46.4 3.69 46.56 9.2 ;
      RECT 46.715 3.66 47.035 3.98 ;
      RECT 46.4 3.69 47.035 3.86 ;
      RECT 35.135 4.15 35.415 4.52 ;
      RECT 35.19 2.355 35.36 4.52 ;
      RECT 45.185 2.35 45.355 3.11 ;
      RECT 45.095 2.755 45.435 3.105 ;
      RECT 45.095 2.355 45.355 3.105 ;
      RECT 45.13 2.35 45.355 3.105 ;
      RECT 35.19 2.355 45.355 2.515 ;
      RECT 41.815 3.59 42.095 3.96 ;
      RECT 40.745 3.615 41.005 3.935 ;
      RECT 43.295 3.425 43.575 3.795 ;
      RECT 43.905 3.335 44.165 3.655 ;
      RECT 40.805 2.775 40.945 3.935 ;
      RECT 41.885 2.775 42.025 3.96 ;
      RECT 43.005 3.425 44.165 3.565 ;
      RECT 43.005 2.775 43.145 3.565 ;
      RECT 40.805 2.775 43.145 2.915 ;
      RECT 40.835 4.915 43.01 5.08 ;
      RECT 42.865 3.795 43.01 5.08 ;
      RECT 39.755 4.71 40.035 5.08 ;
      RECT 39.755 4.825 40.975 4.965 ;
      RECT 42.585 3.795 43.01 3.935 ;
      RECT 42.585 3.615 42.845 3.935 ;
      RECT 35.925 5.195 39.585 5.335 ;
      RECT 39.445 4.38 39.585 5.335 ;
      RECT 35.925 4.265 36.065 5.335 ;
      RECT 42.465 4.455 42.725 4.775 ;
      RECT 39.445 4.38 41.975 4.52 ;
      RECT 41.695 4.15 41.975 4.52 ;
      RECT 35.925 4.265 36.375 4.52 ;
      RECT 36.095 4.15 36.375 4.52 ;
      RECT 42.465 4.265 42.665 4.775 ;
      RECT 41.695 4.265 42.665 4.405 ;
      RECT 42.265 3.055 42.405 4.405 ;
      RECT 42.205 3.055 42.465 3.375 ;
      RECT 33.57 8.94 33.92 9.29 ;
      RECT 42.075 8.895 42.425 9.245 ;
      RECT 33.57 8.97 42.425 9.17 ;
      RECT 36.105 3.615 36.365 3.935 ;
      RECT 36.105 3.705 37.145 3.845 ;
      RECT 37.005 2.915 37.145 3.845 ;
      RECT 39.765 3.055 40.025 3.375 ;
      RECT 37.005 2.915 39.965 3.055 ;
      RECT 39.145 3.895 39.405 4.215 ;
      RECT 39.145 3.895 39.465 4.125 ;
      RECT 39.255 3.59 39.535 3.96 ;
      RECT 38.845 4.455 39.165 4.775 ;
      RECT 38.845 3.335 38.985 4.775 ;
      RECT 38.785 3.335 39.045 3.655 ;
      RECT 36.345 4.735 36.605 5.055 ;
      RECT 36.345 4.825 38.025 4.965 ;
      RECT 37.885 4.545 38.025 4.965 ;
      RECT 37.885 4.545 38.325 4.775 ;
      RECT 38.065 4.455 38.325 4.775 ;
      RECT 37.385 3.615 37.785 4.125 ;
      RECT 37.575 3.59 37.855 3.96 ;
      RECT 37.325 3.615 37.855 3.935 ;
      RECT 30.39 8.505 30.71 8.83 ;
      RECT 30.42 7.98 30.59 8.83 ;
      RECT 30.42 7.98 30.595 8.33 ;
      RECT 30.42 7.98 31.395 8.155 ;
      RECT 31.22 3.26 31.395 8.155 ;
      RECT 31.165 3.26 31.515 3.61 ;
      RECT 31.19 8.94 31.515 9.265 ;
      RECT 30.075 9.03 31.515 9.2 ;
      RECT 30.075 3.69 30.235 9.2 ;
      RECT 30.39 3.66 30.71 3.98 ;
      RECT 30.075 3.69 30.71 3.86 ;
      RECT 18.81 4.15 19.09 4.52 ;
      RECT 18.865 2.355 19.035 4.52 ;
      RECT 28.86 2.35 29.03 3.11 ;
      RECT 28.77 2.755 29.11 3.105 ;
      RECT 28.77 2.355 29.03 3.105 ;
      RECT 28.805 2.35 29.03 3.105 ;
      RECT 18.865 2.355 29.03 2.515 ;
      RECT 25.49 3.59 25.77 3.96 ;
      RECT 24.42 3.615 24.68 3.935 ;
      RECT 26.97 3.425 27.25 3.795 ;
      RECT 27.58 3.335 27.84 3.655 ;
      RECT 24.48 2.775 24.62 3.935 ;
      RECT 25.56 2.775 25.7 3.96 ;
      RECT 26.68 3.425 27.84 3.565 ;
      RECT 26.68 2.775 26.82 3.565 ;
      RECT 24.48 2.775 26.82 2.915 ;
      RECT 16.54 9.28 16.83 9.63 ;
      RECT 16.54 9.335 17.88 9.505 ;
      RECT 17.71 8.97 17.88 9.505 ;
      RECT 26.585 8.89 26.935 9.24 ;
      RECT 17.71 8.97 26.935 9.14 ;
      RECT 24.51 4.915 26.685 5.08 ;
      RECT 26.54 3.795 26.685 5.08 ;
      RECT 23.43 4.71 23.71 5.08 ;
      RECT 23.43 4.825 24.65 4.965 ;
      RECT 26.26 3.795 26.685 3.935 ;
      RECT 26.26 3.615 26.52 3.935 ;
      RECT 19.6 5.195 23.26 5.335 ;
      RECT 23.12 4.38 23.26 5.335 ;
      RECT 19.6 4.265 19.74 5.335 ;
      RECT 26.14 4.455 26.4 4.775 ;
      RECT 23.12 4.38 25.65 4.52 ;
      RECT 25.37 4.15 25.65 4.52 ;
      RECT 19.6 4.265 20.05 4.52 ;
      RECT 19.77 4.15 20.05 4.52 ;
      RECT 26.14 4.265 26.34 4.775 ;
      RECT 25.37 4.265 26.34 4.405 ;
      RECT 25.94 3.055 26.08 4.405 ;
      RECT 25.88 3.055 26.14 3.375 ;
      RECT 19.78 3.615 20.04 3.935 ;
      RECT 19.78 3.705 20.82 3.845 ;
      RECT 20.68 2.915 20.82 3.845 ;
      RECT 23.44 3.055 23.7 3.375 ;
      RECT 20.68 2.915 23.64 3.055 ;
      RECT 22.82 3.895 23.08 4.215 ;
      RECT 22.82 3.895 23.14 4.125 ;
      RECT 22.93 3.59 23.21 3.96 ;
      RECT 22.52 4.455 22.84 4.775 ;
      RECT 22.52 3.335 22.66 4.775 ;
      RECT 22.46 3.335 22.72 3.655 ;
      RECT 20.02 4.735 20.28 5.055 ;
      RECT 20.02 4.825 21.7 4.965 ;
      RECT 21.56 4.545 21.7 4.965 ;
      RECT 21.56 4.545 22 4.775 ;
      RECT 21.74 4.455 22 4.775 ;
      RECT 21.06 3.615 21.46 4.125 ;
      RECT 21.25 3.59 21.53 3.96 ;
      RECT 21 3.615 21.53 3.935 ;
      RECT 90.4 9.34 90.77 9.71 ;
      RECT 89.11 3.59 89.39 3.96 ;
      RECT 87.27 3.59 87.55 3.96 ;
      RECT 85.55 3.03 85.83 3.4 ;
      RECT 74.075 9.34 74.445 9.71 ;
      RECT 72.785 3.59 73.065 3.96 ;
      RECT 70.945 3.59 71.225 3.96 ;
      RECT 69.225 3.03 69.505 3.4 ;
      RECT 57.75 9.34 58.12 9.71 ;
      RECT 56.46 3.59 56.74 3.96 ;
      RECT 54.62 3.59 54.9 3.96 ;
      RECT 52.9 3.03 53.18 3.4 ;
      RECT 41.425 9.34 41.795 9.71 ;
      RECT 40.135 3.59 40.415 3.96 ;
      RECT 38.295 3.59 38.575 3.96 ;
      RECT 36.575 3.03 36.855 3.4 ;
      RECT 25.1 9.34 25.47 9.71 ;
      RECT 23.81 3.59 24.09 3.96 ;
      RECT 21.97 3.59 22.25 3.96 ;
      RECT 20.25 3.03 20.53 3.4 ;
    LAYER via1 ;
      RECT 98.95 9.66 99.1 9.81 ;
      RECT 96.58 9.025 96.73 9.175 ;
      RECT 96.565 3.36 96.715 3.51 ;
      RECT 95.775 3.745 95.925 3.895 ;
      RECT 95.775 8.61 95.925 8.76 ;
      RECT 94.17 2.855 94.32 3.005 ;
      RECT 92.935 3.42 93.085 3.57 ;
      RECT 91.615 3.7 91.765 3.85 ;
      RECT 91.495 4.54 91.645 4.69 ;
      RECT 91.235 3.14 91.385 3.29 ;
      RECT 91.155 8.995 91.305 9.145 ;
      RECT 90.51 9.45 90.66 9.6 ;
      RECT 89.775 3.7 89.925 3.85 ;
      RECT 89.175 3.7 89.325 3.85 ;
      RECT 88.795 3.14 88.945 3.29 ;
      RECT 88.175 3.98 88.325 4.13 ;
      RECT 87.935 4.54 88.085 4.69 ;
      RECT 87.815 3.42 87.965 3.57 ;
      RECT 87.335 3.7 87.485 3.85 ;
      RECT 87.095 4.54 87.245 4.69 ;
      RECT 86.355 3.7 86.505 3.85 ;
      RECT 85.615 3.14 85.765 3.29 ;
      RECT 85.375 4.82 85.525 4.97 ;
      RECT 85.135 3.7 85.285 3.85 ;
      RECT 85.135 4.26 85.285 4.41 ;
      RECT 84.175 4.26 84.325 4.41 ;
      RECT 82.6 9.04 82.75 9.19 ;
      RECT 80.255 9.025 80.405 9.175 ;
      RECT 80.24 3.36 80.39 3.51 ;
      RECT 79.45 3.745 79.6 3.895 ;
      RECT 79.45 8.61 79.6 8.76 ;
      RECT 77.845 2.855 77.995 3.005 ;
      RECT 76.61 3.42 76.76 3.57 ;
      RECT 75.29 3.7 75.44 3.85 ;
      RECT 75.17 4.54 75.32 4.69 ;
      RECT 74.91 3.14 75.06 3.29 ;
      RECT 74.825 8.995 74.975 9.145 ;
      RECT 74.185 9.45 74.335 9.6 ;
      RECT 73.45 3.7 73.6 3.85 ;
      RECT 72.85 3.7 73 3.85 ;
      RECT 72.47 3.14 72.62 3.29 ;
      RECT 71.85 3.98 72 4.13 ;
      RECT 71.61 4.54 71.76 4.69 ;
      RECT 71.49 3.42 71.64 3.57 ;
      RECT 71.01 3.7 71.16 3.85 ;
      RECT 70.77 4.54 70.92 4.69 ;
      RECT 70.03 3.7 70.18 3.85 ;
      RECT 69.29 3.14 69.44 3.29 ;
      RECT 69.05 4.82 69.2 4.97 ;
      RECT 68.81 3.7 68.96 3.85 ;
      RECT 68.81 4.26 68.96 4.41 ;
      RECT 67.85 4.26 68 4.41 ;
      RECT 66.275 9.04 66.425 9.19 ;
      RECT 63.93 9.025 64.08 9.175 ;
      RECT 63.915 3.36 64.065 3.51 ;
      RECT 63.125 3.745 63.275 3.895 ;
      RECT 63.125 8.61 63.275 8.76 ;
      RECT 61.52 2.855 61.67 3.005 ;
      RECT 60.285 3.42 60.435 3.57 ;
      RECT 58.965 3.7 59.115 3.85 ;
      RECT 58.845 4.54 58.995 4.69 ;
      RECT 58.585 3.14 58.735 3.29 ;
      RECT 58.5 9 58.65 9.15 ;
      RECT 57.86 9.45 58.01 9.6 ;
      RECT 57.125 3.7 57.275 3.85 ;
      RECT 56.525 3.7 56.675 3.85 ;
      RECT 56.145 3.14 56.295 3.29 ;
      RECT 55.525 3.98 55.675 4.13 ;
      RECT 55.285 4.54 55.435 4.69 ;
      RECT 55.165 3.42 55.315 3.57 ;
      RECT 54.685 3.7 54.835 3.85 ;
      RECT 54.445 4.54 54.595 4.69 ;
      RECT 53.705 3.7 53.855 3.85 ;
      RECT 52.965 3.14 53.115 3.29 ;
      RECT 52.725 4.82 52.875 4.97 ;
      RECT 52.485 3.7 52.635 3.85 ;
      RECT 52.485 4.26 52.635 4.41 ;
      RECT 51.525 4.26 51.675 4.41 ;
      RECT 49.995 9.045 50.145 9.195 ;
      RECT 47.605 9.025 47.755 9.175 ;
      RECT 47.59 3.36 47.74 3.51 ;
      RECT 46.8 3.745 46.95 3.895 ;
      RECT 46.8 8.61 46.95 8.76 ;
      RECT 45.195 2.855 45.345 3.005 ;
      RECT 43.96 3.42 44.11 3.57 ;
      RECT 42.64 3.7 42.79 3.85 ;
      RECT 42.52 4.54 42.67 4.69 ;
      RECT 42.26 3.14 42.41 3.29 ;
      RECT 42.175 8.995 42.325 9.145 ;
      RECT 41.535 9.45 41.685 9.6 ;
      RECT 40.8 3.7 40.95 3.85 ;
      RECT 40.2 3.7 40.35 3.85 ;
      RECT 39.82 3.14 39.97 3.29 ;
      RECT 39.2 3.98 39.35 4.13 ;
      RECT 38.96 4.54 39.11 4.69 ;
      RECT 38.84 3.42 38.99 3.57 ;
      RECT 38.36 3.7 38.51 3.85 ;
      RECT 38.12 4.54 38.27 4.69 ;
      RECT 37.38 3.7 37.53 3.85 ;
      RECT 36.64 3.14 36.79 3.29 ;
      RECT 36.4 4.82 36.55 4.97 ;
      RECT 36.16 3.7 36.31 3.85 ;
      RECT 36.16 4.26 36.31 4.41 ;
      RECT 35.2 4.26 35.35 4.41 ;
      RECT 33.67 9.04 33.82 9.19 ;
      RECT 31.28 9.025 31.43 9.175 ;
      RECT 31.265 3.36 31.415 3.51 ;
      RECT 30.475 3.745 30.625 3.895 ;
      RECT 30.475 8.61 30.625 8.76 ;
      RECT 28.87 2.855 29.02 3.005 ;
      RECT 27.635 3.42 27.785 3.57 ;
      RECT 26.685 8.99 26.835 9.14 ;
      RECT 26.315 3.7 26.465 3.85 ;
      RECT 26.195 4.54 26.345 4.69 ;
      RECT 25.935 3.14 26.085 3.29 ;
      RECT 25.21 9.45 25.36 9.6 ;
      RECT 24.475 3.7 24.625 3.85 ;
      RECT 23.875 3.7 24.025 3.85 ;
      RECT 23.495 3.14 23.645 3.29 ;
      RECT 22.875 3.98 23.025 4.13 ;
      RECT 22.635 4.54 22.785 4.69 ;
      RECT 22.515 3.42 22.665 3.57 ;
      RECT 22.035 3.7 22.185 3.85 ;
      RECT 21.795 4.54 21.945 4.69 ;
      RECT 21.055 3.7 21.205 3.85 ;
      RECT 20.315 3.14 20.465 3.29 ;
      RECT 20.075 4.82 20.225 4.97 ;
      RECT 19.835 3.7 19.985 3.85 ;
      RECT 19.835 4.26 19.985 4.41 ;
      RECT 18.875 4.26 19.025 4.41 ;
      RECT 16.61 9.38 16.76 9.53 ;
      RECT 16.235 8.64 16.385 8.79 ;
    LAYER met1 ;
      RECT 98.82 10.05 99.115 10.28 ;
      RECT 98.88 9.56 99.055 10.28 ;
      RECT 98.85 9.56 99.2 9.91 ;
      RECT 98.88 8.57 99.05 10.28 ;
      RECT 98.82 8.57 99.11 8.8 ;
      RECT 97.825 10.055 98.12 10.285 ;
      RECT 97.885 8.575 98.055 10.285 ;
      RECT 97.825 8.575 98.115 8.805 ;
      RECT 97.825 8.61 98.68 8.77 ;
      RECT 98.51 8.2 98.68 8.77 ;
      RECT 97.825 8.605 98.22 8.77 ;
      RECT 98.45 8.2 98.74 8.43 ;
      RECT 98.45 8.23 98.91 8.4 ;
      RECT 98.41 4.03 98.735 4.26 ;
      RECT 98.41 4.06 98.905 4.23 ;
      RECT 98.41 3.69 98.6 4.26 ;
      RECT 97.825 3.655 98.115 3.885 ;
      RECT 97.825 3.69 98.6 3.86 ;
      RECT 97.885 2.175 98.055 3.885 ;
      RECT 97.825 2.175 98.12 2.405 ;
      RECT 97.455 4.025 97.745 4.255 ;
      RECT 97.455 4.055 97.915 4.225 ;
      RECT 97.52 2.95 97.685 4.255 ;
      RECT 96.035 2.915 96.325 3.145 ;
      RECT 96.035 2.95 97.685 3.12 ;
      RECT 96.095 2.175 96.265 3.145 ;
      RECT 96.035 2.175 96.325 2.405 ;
      RECT 96.035 10.055 96.325 10.285 ;
      RECT 96.095 9.315 96.265 10.285 ;
      RECT 96.095 9.405 97.685 9.575 ;
      RECT 97.515 8.205 97.685 9.575 ;
      RECT 96.035 9.315 96.325 9.545 ;
      RECT 97.455 8.205 97.745 8.435 ;
      RECT 97.455 8.235 97.915 8.405 ;
      RECT 96.465 3.26 96.815 3.61 ;
      RECT 94.16 3.32 96.815 3.49 ;
      RECT 96.295 3.315 96.815 3.49 ;
      RECT 94.16 2.755 94.33 3.49 ;
      RECT 94.07 2.755 94.41 3.105 ;
      RECT 96.49 8.94 96.815 9.265 ;
      RECT 91.055 8.895 91.405 9.245 ;
      RECT 96.465 8.945 96.815 9.175 ;
      RECT 90.85 8.945 91.405 9.175 ;
      RECT 96.295 8.97 96.815 9.145 ;
      RECT 90.68 8.975 91.405 9.145 ;
      RECT 90.85 8.97 96.815 9.14 ;
      RECT 95.69 3.66 96.01 3.98 ;
      RECT 95.665 3.655 95.955 3.885 ;
      RECT 95.66 3.685 96.01 3.86 ;
      RECT 95.49 3.685 96.01 3.855 ;
      RECT 95.69 8.54 96.01 8.83 ;
      RECT 95.665 8.575 96.01 8.805 ;
      RECT 95.49 8.605 96.01 8.775 ;
      RECT 92.145 3.66 92.435 3.89 ;
      RECT 92.145 3.66 92.6 3.845 ;
      RECT 92.46 3.565 93.08 3.705 ;
      RECT 92.85 3.365 93.17 3.625 ;
      RECT 91.53 3.645 91.85 3.905 ;
      RECT 91.53 3.645 91.995 3.89 ;
      RECT 91.855 3.265 91.995 3.89 ;
      RECT 91.855 3.265 92.12 3.405 ;
      RECT 92.385 3.1 92.675 3.33 ;
      RECT 91.98 3.145 92.675 3.285 ;
      RECT 91.425 4.485 91.715 5.01 ;
      RECT 91.41 4.485 91.73 4.745 ;
      RECT 91.15 3.085 91.47 3.345 ;
      RECT 91.15 3.1 91.715 3.33 ;
      RECT 90.425 4.78 90.715 5.01 ;
      RECT 90.62 3.425 90.76 4.965 ;
      RECT 90.665 3.38 90.955 3.61 ;
      RECT 90.26 3.425 90.955 3.565 ;
      RECT 90.26 3.265 90.4 3.565 ;
      RECT 88.8 3.265 90.4 3.405 ;
      RECT 88.71 3.085 89.03 3.345 ;
      RECT 88.71 3.1 89.275 3.345 ;
      RECT 90.42 10.055 90.71 10.285 ;
      RECT 90.48 9.315 90.65 10.285 ;
      RECT 90.4 9.36 90.77 9.71 ;
      RECT 90.4 9.34 90.71 9.71 ;
      RECT 90.42 9.315 90.71 9.71 ;
      RECT 87.82 4.125 90.4 4.265 ;
      RECT 90.185 3.94 90.475 4.17 ;
      RECT 87.745 3.94 88.41 4.17 ;
      RECT 88.09 3.925 88.41 4.265 ;
      RECT 89.09 3.645 89.41 3.905 ;
      RECT 89.09 3.66 89.515 3.89 ;
      RECT 87.73 3.365 88.05 3.625 ;
      RECT 88.225 3.38 88.515 3.61 ;
      RECT 87.73 3.425 88.515 3.565 ;
      RECT 87.85 4.485 88.17 4.745 ;
      RECT 87.01 4.485 87.33 4.745 ;
      RECT 87.85 4.5 88.275 4.73 ;
      RECT 87.01 4.545 88.275 4.685 ;
      RECT 86.545 4.22 86.835 4.45 ;
      RECT 86.62 3.145 86.76 4.45 ;
      RECT 86.27 3.645 86.76 3.905 ;
      RECT 86.025 3.66 86.76 3.89 ;
      RECT 87.025 3.1 87.315 3.33 ;
      RECT 86.62 3.145 87.315 3.285 ;
      RECT 85.785 4.5 86.075 4.73 ;
      RECT 85.785 4.5 86.24 4.685 ;
      RECT 86.1 4.125 86.24 4.685 ;
      RECT 85.74 4.125 86.24 4.265 ;
      RECT 85.74 3.145 85.88 4.265 ;
      RECT 85.53 3.085 85.85 3.345 ;
      RECT 85.29 4.765 85.61 5.025 ;
      RECT 84.585 4.78 84.875 5.01 ;
      RECT 84.585 4.825 85.61 4.965 ;
      RECT 84.66 4.775 84.92 4.965 ;
      RECT 85.05 3.645 85.37 3.905 ;
      RECT 85.05 3.66 85.595 3.89 ;
      RECT 85.05 4.205 85.37 4.465 ;
      RECT 85.05 4.22 85.595 4.45 ;
      RECT 84.09 4.205 84.41 4.465 ;
      RECT 84.18 3.145 84.32 4.465 ;
      RECT 84.585 3.1 84.875 3.33 ;
      RECT 84.18 3.145 84.875 3.285 ;
      RECT 82.495 10.05 82.79 10.28 ;
      RECT 82.555 8.57 82.725 10.28 ;
      RECT 82.5 8.94 82.85 9.29 ;
      RECT 82.495 8.57 82.785 8.8 ;
      RECT 81.5 10.055 81.795 10.285 ;
      RECT 81.56 8.575 81.73 10.285 ;
      RECT 81.5 8.575 81.79 8.805 ;
      RECT 81.5 8.61 82.355 8.77 ;
      RECT 82.185 8.2 82.355 8.77 ;
      RECT 81.5 8.605 81.895 8.77 ;
      RECT 82.125 8.2 82.415 8.43 ;
      RECT 82.125 8.23 82.585 8.4 ;
      RECT 82.085 4.03 82.41 4.26 ;
      RECT 82.085 4.06 82.58 4.23 ;
      RECT 82.085 3.69 82.275 4.26 ;
      RECT 81.5 3.655 81.79 3.885 ;
      RECT 81.5 3.69 82.275 3.86 ;
      RECT 81.56 2.175 81.73 3.885 ;
      RECT 81.5 2.175 81.795 2.405 ;
      RECT 81.13 4.025 81.42 4.255 ;
      RECT 81.13 4.055 81.59 4.225 ;
      RECT 81.195 2.95 81.36 4.255 ;
      RECT 79.71 2.915 80 3.145 ;
      RECT 79.71 2.95 81.36 3.12 ;
      RECT 79.77 2.175 79.94 3.145 ;
      RECT 79.71 2.175 80 2.405 ;
      RECT 79.71 10.055 80 10.285 ;
      RECT 79.77 9.315 79.94 10.285 ;
      RECT 79.77 9.405 81.36 9.575 ;
      RECT 81.19 8.205 81.36 9.575 ;
      RECT 79.71 9.315 80 9.545 ;
      RECT 81.13 8.205 81.42 8.435 ;
      RECT 81.13 8.235 81.59 8.405 ;
      RECT 80.14 3.26 80.49 3.61 ;
      RECT 77.835 3.32 80.49 3.49 ;
      RECT 79.97 3.315 80.49 3.49 ;
      RECT 77.835 2.755 78.005 3.49 ;
      RECT 77.745 2.755 78.085 3.105 ;
      RECT 80.165 8.94 80.49 9.265 ;
      RECT 74.725 8.895 75.075 9.245 ;
      RECT 80.14 8.945 80.49 9.175 ;
      RECT 74.525 8.945 75.075 9.175 ;
      RECT 79.97 8.97 80.49 9.145 ;
      RECT 74.355 8.975 75.075 9.145 ;
      RECT 74.525 8.97 80.49 9.14 ;
      RECT 79.365 3.66 79.685 3.98 ;
      RECT 79.34 3.655 79.63 3.885 ;
      RECT 79.335 3.685 79.685 3.86 ;
      RECT 79.165 3.685 79.685 3.855 ;
      RECT 79.365 8.54 79.685 8.83 ;
      RECT 79.34 8.575 79.685 8.805 ;
      RECT 79.165 8.605 79.685 8.775 ;
      RECT 75.82 3.66 76.11 3.89 ;
      RECT 75.82 3.66 76.275 3.845 ;
      RECT 76.135 3.565 76.755 3.705 ;
      RECT 76.525 3.365 76.845 3.625 ;
      RECT 75.205 3.645 75.525 3.905 ;
      RECT 75.205 3.645 75.67 3.89 ;
      RECT 75.53 3.265 75.67 3.89 ;
      RECT 75.53 3.265 75.795 3.405 ;
      RECT 76.06 3.1 76.35 3.33 ;
      RECT 75.655 3.145 76.35 3.285 ;
      RECT 75.1 4.485 75.39 5.01 ;
      RECT 75.085 4.485 75.405 4.745 ;
      RECT 74.825 3.085 75.145 3.345 ;
      RECT 74.825 3.1 75.39 3.33 ;
      RECT 74.1 4.78 74.39 5.01 ;
      RECT 74.295 3.425 74.435 4.965 ;
      RECT 74.34 3.38 74.63 3.61 ;
      RECT 73.935 3.425 74.63 3.565 ;
      RECT 73.935 3.265 74.075 3.565 ;
      RECT 72.475 3.265 74.075 3.405 ;
      RECT 72.385 3.085 72.705 3.345 ;
      RECT 72.385 3.1 72.95 3.345 ;
      RECT 74.095 10.055 74.385 10.285 ;
      RECT 74.155 9.315 74.325 10.285 ;
      RECT 74.075 9.36 74.445 9.71 ;
      RECT 74.075 9.34 74.385 9.71 ;
      RECT 74.095 9.315 74.385 9.71 ;
      RECT 71.495 4.125 74.075 4.265 ;
      RECT 73.86 3.94 74.15 4.17 ;
      RECT 71.42 3.94 72.085 4.17 ;
      RECT 71.765 3.925 72.085 4.265 ;
      RECT 72.765 3.645 73.085 3.905 ;
      RECT 72.765 3.66 73.19 3.89 ;
      RECT 71.405 3.365 71.725 3.625 ;
      RECT 71.9 3.38 72.19 3.61 ;
      RECT 71.405 3.425 72.19 3.565 ;
      RECT 71.525 4.485 71.845 4.745 ;
      RECT 70.685 4.485 71.005 4.745 ;
      RECT 71.525 4.5 71.95 4.73 ;
      RECT 70.685 4.545 71.95 4.685 ;
      RECT 70.22 4.22 70.51 4.45 ;
      RECT 70.295 3.145 70.435 4.45 ;
      RECT 69.945 3.645 70.435 3.905 ;
      RECT 69.7 3.66 70.435 3.89 ;
      RECT 70.7 3.1 70.99 3.33 ;
      RECT 70.295 3.145 70.99 3.285 ;
      RECT 69.46 4.5 69.75 4.73 ;
      RECT 69.46 4.5 69.915 4.685 ;
      RECT 69.775 4.125 69.915 4.685 ;
      RECT 69.415 4.125 69.915 4.265 ;
      RECT 69.415 3.145 69.555 4.265 ;
      RECT 69.205 3.085 69.525 3.345 ;
      RECT 68.965 4.765 69.285 5.025 ;
      RECT 68.26 4.78 68.55 5.01 ;
      RECT 68.26 4.825 69.285 4.965 ;
      RECT 68.335 4.775 68.595 4.965 ;
      RECT 68.725 3.645 69.045 3.905 ;
      RECT 68.725 3.66 69.27 3.89 ;
      RECT 68.725 4.205 69.045 4.465 ;
      RECT 68.725 4.22 69.27 4.45 ;
      RECT 67.765 4.205 68.085 4.465 ;
      RECT 67.855 3.145 67.995 4.465 ;
      RECT 68.26 3.1 68.55 3.33 ;
      RECT 67.855 3.145 68.55 3.285 ;
      RECT 66.17 10.05 66.465 10.28 ;
      RECT 66.23 8.57 66.4 10.28 ;
      RECT 66.175 8.94 66.525 9.29 ;
      RECT 66.17 8.57 66.46 8.8 ;
      RECT 65.175 10.055 65.47 10.285 ;
      RECT 65.235 8.575 65.405 10.285 ;
      RECT 65.175 8.575 65.465 8.805 ;
      RECT 65.175 8.61 66.03 8.77 ;
      RECT 65.86 8.2 66.03 8.77 ;
      RECT 65.175 8.605 65.57 8.77 ;
      RECT 65.8 8.2 66.09 8.43 ;
      RECT 65.8 8.23 66.26 8.4 ;
      RECT 65.76 4.03 66.085 4.26 ;
      RECT 65.76 4.06 66.255 4.23 ;
      RECT 65.76 3.69 65.95 4.26 ;
      RECT 65.175 3.655 65.465 3.885 ;
      RECT 65.175 3.69 65.95 3.86 ;
      RECT 65.235 2.175 65.405 3.885 ;
      RECT 65.175 2.175 65.47 2.405 ;
      RECT 64.805 4.025 65.095 4.255 ;
      RECT 64.805 4.055 65.265 4.225 ;
      RECT 64.87 2.95 65.035 4.255 ;
      RECT 63.385 2.915 63.675 3.145 ;
      RECT 63.385 2.95 65.035 3.12 ;
      RECT 63.445 2.175 63.615 3.145 ;
      RECT 63.385 2.175 63.675 2.405 ;
      RECT 63.385 10.055 63.675 10.285 ;
      RECT 63.445 9.315 63.615 10.285 ;
      RECT 63.445 9.405 65.035 9.575 ;
      RECT 64.865 8.205 65.035 9.575 ;
      RECT 63.385 9.315 63.675 9.545 ;
      RECT 64.805 8.205 65.095 8.435 ;
      RECT 64.805 8.235 65.265 8.405 ;
      RECT 63.815 3.26 64.165 3.61 ;
      RECT 61.51 3.32 64.165 3.49 ;
      RECT 63.645 3.315 64.165 3.49 ;
      RECT 61.51 2.755 61.68 3.49 ;
      RECT 61.42 2.755 61.76 3.105 ;
      RECT 63.84 8.94 64.165 9.265 ;
      RECT 58.4 8.9 58.75 9.25 ;
      RECT 63.815 8.945 64.165 9.175 ;
      RECT 58.2 8.945 58.75 9.175 ;
      RECT 63.645 8.97 64.165 9.145 ;
      RECT 58.03 8.975 58.75 9.145 ;
      RECT 58.2 8.97 64.165 9.14 ;
      RECT 63.04 3.66 63.36 3.98 ;
      RECT 63.015 3.655 63.305 3.885 ;
      RECT 63.01 3.685 63.36 3.86 ;
      RECT 62.84 3.685 63.36 3.855 ;
      RECT 63.04 8.54 63.36 8.83 ;
      RECT 63.015 8.575 63.36 8.805 ;
      RECT 62.84 8.605 63.36 8.775 ;
      RECT 59.495 3.66 59.785 3.89 ;
      RECT 59.495 3.66 59.95 3.845 ;
      RECT 59.81 3.565 60.43 3.705 ;
      RECT 60.2 3.365 60.52 3.625 ;
      RECT 58.88 3.645 59.2 3.905 ;
      RECT 58.88 3.645 59.345 3.89 ;
      RECT 59.205 3.265 59.345 3.89 ;
      RECT 59.205 3.265 59.47 3.405 ;
      RECT 59.735 3.1 60.025 3.33 ;
      RECT 59.33 3.145 60.025 3.285 ;
      RECT 58.775 4.485 59.065 5.01 ;
      RECT 58.76 4.485 59.08 4.745 ;
      RECT 58.5 3.085 58.82 3.345 ;
      RECT 58.5 3.1 59.065 3.33 ;
      RECT 57.775 4.78 58.065 5.01 ;
      RECT 57.97 3.425 58.11 4.965 ;
      RECT 58.015 3.38 58.305 3.61 ;
      RECT 57.61 3.425 58.305 3.565 ;
      RECT 57.61 3.265 57.75 3.565 ;
      RECT 56.15 3.265 57.75 3.405 ;
      RECT 56.06 3.085 56.38 3.345 ;
      RECT 56.06 3.1 56.625 3.345 ;
      RECT 57.77 10.055 58.06 10.285 ;
      RECT 57.83 9.315 58 10.285 ;
      RECT 57.75 9.36 58.12 9.71 ;
      RECT 57.75 9.34 58.06 9.71 ;
      RECT 57.77 9.315 58.06 9.71 ;
      RECT 55.17 4.125 57.75 4.265 ;
      RECT 57.535 3.94 57.825 4.17 ;
      RECT 55.095 3.94 55.76 4.17 ;
      RECT 55.44 3.925 55.76 4.265 ;
      RECT 56.44 3.645 56.76 3.905 ;
      RECT 56.44 3.66 56.865 3.89 ;
      RECT 55.08 3.365 55.4 3.625 ;
      RECT 55.575 3.38 55.865 3.61 ;
      RECT 55.08 3.425 55.865 3.565 ;
      RECT 55.2 4.485 55.52 4.745 ;
      RECT 54.36 4.485 54.68 4.745 ;
      RECT 55.2 4.5 55.625 4.73 ;
      RECT 54.36 4.545 55.625 4.685 ;
      RECT 53.895 4.22 54.185 4.45 ;
      RECT 53.97 3.145 54.11 4.45 ;
      RECT 53.62 3.645 54.11 3.905 ;
      RECT 53.375 3.66 54.11 3.89 ;
      RECT 54.375 3.1 54.665 3.33 ;
      RECT 53.97 3.145 54.665 3.285 ;
      RECT 53.135 4.5 53.425 4.73 ;
      RECT 53.135 4.5 53.59 4.685 ;
      RECT 53.45 4.125 53.59 4.685 ;
      RECT 53.09 4.125 53.59 4.265 ;
      RECT 53.09 3.145 53.23 4.265 ;
      RECT 52.88 3.085 53.2 3.345 ;
      RECT 52.64 4.765 52.96 5.025 ;
      RECT 51.935 4.78 52.225 5.01 ;
      RECT 51.935 4.825 52.96 4.965 ;
      RECT 52.01 4.775 52.27 4.965 ;
      RECT 52.4 3.645 52.72 3.905 ;
      RECT 52.4 3.66 52.945 3.89 ;
      RECT 52.4 4.205 52.72 4.465 ;
      RECT 52.4 4.22 52.945 4.45 ;
      RECT 51.44 4.205 51.76 4.465 ;
      RECT 51.53 3.145 51.67 4.465 ;
      RECT 51.935 3.1 52.225 3.33 ;
      RECT 51.53 3.145 52.225 3.285 ;
      RECT 49.845 10.05 50.14 10.28 ;
      RECT 49.905 8.57 50.075 10.28 ;
      RECT 49.89 8.945 50.245 9.3 ;
      RECT 49.845 8.57 50.135 8.8 ;
      RECT 48.85 10.055 49.145 10.285 ;
      RECT 48.91 8.575 49.08 10.285 ;
      RECT 48.85 8.575 49.14 8.805 ;
      RECT 48.85 8.61 49.705 8.77 ;
      RECT 49.535 8.2 49.705 8.77 ;
      RECT 48.85 8.605 49.245 8.77 ;
      RECT 49.475 8.2 49.765 8.43 ;
      RECT 49.475 8.23 49.935 8.4 ;
      RECT 49.435 4.03 49.76 4.26 ;
      RECT 49.435 4.06 49.93 4.23 ;
      RECT 49.435 3.69 49.625 4.26 ;
      RECT 48.85 3.655 49.14 3.885 ;
      RECT 48.85 3.69 49.625 3.86 ;
      RECT 48.91 2.175 49.08 3.885 ;
      RECT 48.85 2.175 49.145 2.405 ;
      RECT 48.48 4.025 48.77 4.255 ;
      RECT 48.48 4.055 48.94 4.225 ;
      RECT 48.545 2.95 48.71 4.255 ;
      RECT 47.06 2.915 47.35 3.145 ;
      RECT 47.06 2.95 48.71 3.12 ;
      RECT 47.12 2.175 47.29 3.145 ;
      RECT 47.06 2.175 47.35 2.405 ;
      RECT 47.06 10.055 47.35 10.285 ;
      RECT 47.12 9.315 47.29 10.285 ;
      RECT 47.12 9.405 48.71 9.575 ;
      RECT 48.54 8.205 48.71 9.575 ;
      RECT 47.06 9.315 47.35 9.545 ;
      RECT 48.48 8.205 48.77 8.435 ;
      RECT 48.48 8.235 48.94 8.405 ;
      RECT 47.49 3.26 47.84 3.61 ;
      RECT 45.185 3.32 47.84 3.49 ;
      RECT 47.32 3.315 47.84 3.49 ;
      RECT 45.185 2.755 45.355 3.49 ;
      RECT 45.095 2.755 45.435 3.105 ;
      RECT 47.515 8.94 47.84 9.265 ;
      RECT 42.075 8.895 42.425 9.245 ;
      RECT 47.49 8.945 47.84 9.175 ;
      RECT 41.875 8.945 42.425 9.175 ;
      RECT 47.32 8.97 47.84 9.145 ;
      RECT 41.705 8.975 42.425 9.145 ;
      RECT 41.875 8.97 47.84 9.14 ;
      RECT 46.715 3.66 47.035 3.98 ;
      RECT 46.69 3.655 46.98 3.885 ;
      RECT 46.685 3.685 47.035 3.86 ;
      RECT 46.515 3.685 47.035 3.855 ;
      RECT 46.715 8.54 47.035 8.83 ;
      RECT 46.69 8.575 47.035 8.805 ;
      RECT 46.515 8.605 47.035 8.775 ;
      RECT 43.17 3.66 43.46 3.89 ;
      RECT 43.17 3.66 43.625 3.845 ;
      RECT 43.485 3.565 44.105 3.705 ;
      RECT 43.875 3.365 44.195 3.625 ;
      RECT 42.555 3.645 42.875 3.905 ;
      RECT 42.555 3.645 43.02 3.89 ;
      RECT 42.88 3.265 43.02 3.89 ;
      RECT 42.88 3.265 43.145 3.405 ;
      RECT 43.41 3.1 43.7 3.33 ;
      RECT 43.005 3.145 43.7 3.285 ;
      RECT 42.45 4.485 42.74 5.01 ;
      RECT 42.435 4.485 42.755 4.745 ;
      RECT 42.175 3.085 42.495 3.345 ;
      RECT 42.175 3.1 42.74 3.33 ;
      RECT 41.45 4.78 41.74 5.01 ;
      RECT 41.645 3.425 41.785 4.965 ;
      RECT 41.69 3.38 41.98 3.61 ;
      RECT 41.285 3.425 41.98 3.565 ;
      RECT 41.285 3.265 41.425 3.565 ;
      RECT 39.825 3.265 41.425 3.405 ;
      RECT 39.735 3.085 40.055 3.345 ;
      RECT 39.735 3.1 40.3 3.345 ;
      RECT 41.445 10.055 41.735 10.285 ;
      RECT 41.505 9.315 41.675 10.285 ;
      RECT 41.425 9.36 41.795 9.71 ;
      RECT 41.425 9.34 41.735 9.71 ;
      RECT 41.445 9.315 41.735 9.71 ;
      RECT 38.845 4.125 41.425 4.265 ;
      RECT 41.21 3.94 41.5 4.17 ;
      RECT 38.77 3.94 39.435 4.17 ;
      RECT 39.115 3.925 39.435 4.265 ;
      RECT 40.115 3.645 40.435 3.905 ;
      RECT 40.115 3.66 40.54 3.89 ;
      RECT 38.755 3.365 39.075 3.625 ;
      RECT 39.25 3.38 39.54 3.61 ;
      RECT 38.755 3.425 39.54 3.565 ;
      RECT 38.875 4.485 39.195 4.745 ;
      RECT 38.035 4.485 38.355 4.745 ;
      RECT 38.875 4.5 39.3 4.73 ;
      RECT 38.035 4.545 39.3 4.685 ;
      RECT 37.57 4.22 37.86 4.45 ;
      RECT 37.645 3.145 37.785 4.45 ;
      RECT 37.295 3.645 37.785 3.905 ;
      RECT 37.05 3.66 37.785 3.89 ;
      RECT 38.05 3.1 38.34 3.33 ;
      RECT 37.645 3.145 38.34 3.285 ;
      RECT 36.81 4.5 37.1 4.73 ;
      RECT 36.81 4.5 37.265 4.685 ;
      RECT 37.125 4.125 37.265 4.685 ;
      RECT 36.765 4.125 37.265 4.265 ;
      RECT 36.765 3.145 36.905 4.265 ;
      RECT 36.555 3.085 36.875 3.345 ;
      RECT 36.315 4.765 36.635 5.025 ;
      RECT 35.61 4.78 35.9 5.01 ;
      RECT 35.61 4.825 36.635 4.965 ;
      RECT 35.685 4.775 35.945 4.965 ;
      RECT 36.075 3.645 36.395 3.905 ;
      RECT 36.075 3.66 36.62 3.89 ;
      RECT 36.075 4.205 36.395 4.465 ;
      RECT 36.075 4.22 36.62 4.45 ;
      RECT 35.115 4.205 35.435 4.465 ;
      RECT 35.205 3.145 35.345 4.465 ;
      RECT 35.61 3.1 35.9 3.33 ;
      RECT 35.205 3.145 35.9 3.285 ;
      RECT 33.52 10.05 33.815 10.28 ;
      RECT 33.58 8.57 33.75 10.28 ;
      RECT 33.57 8.94 33.92 9.29 ;
      RECT 33.52 8.57 33.81 8.8 ;
      RECT 32.525 10.055 32.82 10.285 ;
      RECT 32.585 8.575 32.755 10.285 ;
      RECT 32.525 8.575 32.815 8.805 ;
      RECT 32.525 8.61 33.38 8.77 ;
      RECT 33.21 8.2 33.38 8.77 ;
      RECT 32.525 8.605 32.92 8.77 ;
      RECT 33.15 8.2 33.44 8.43 ;
      RECT 33.15 8.23 33.61 8.4 ;
      RECT 33.11 4.03 33.435 4.26 ;
      RECT 33.11 4.06 33.605 4.23 ;
      RECT 33.11 3.69 33.3 4.26 ;
      RECT 32.525 3.655 32.815 3.885 ;
      RECT 32.525 3.69 33.3 3.86 ;
      RECT 32.585 2.175 32.755 3.885 ;
      RECT 32.525 2.175 32.82 2.405 ;
      RECT 32.155 4.025 32.445 4.255 ;
      RECT 32.155 4.055 32.615 4.225 ;
      RECT 32.22 2.95 32.385 4.255 ;
      RECT 30.735 2.915 31.025 3.145 ;
      RECT 30.735 2.95 32.385 3.12 ;
      RECT 30.795 2.175 30.965 3.145 ;
      RECT 30.735 2.175 31.025 2.405 ;
      RECT 30.735 10.055 31.025 10.285 ;
      RECT 30.795 9.315 30.965 10.285 ;
      RECT 30.795 9.405 32.385 9.575 ;
      RECT 32.215 8.205 32.385 9.575 ;
      RECT 30.735 9.315 31.025 9.545 ;
      RECT 32.155 8.205 32.445 8.435 ;
      RECT 32.155 8.235 32.615 8.405 ;
      RECT 31.165 3.26 31.515 3.61 ;
      RECT 28.86 3.32 31.515 3.49 ;
      RECT 30.995 3.315 31.515 3.49 ;
      RECT 28.86 2.755 29.03 3.49 ;
      RECT 28.77 2.755 29.11 3.105 ;
      RECT 31.19 8.94 31.515 9.265 ;
      RECT 26.585 8.89 26.935 9.24 ;
      RECT 31.165 8.945 31.515 9.175 ;
      RECT 25.55 8.945 25.84 9.175 ;
      RECT 30.995 8.97 31.515 9.145 ;
      RECT 25.38 8.975 25.84 9.145 ;
      RECT 25.55 8.97 31.515 9.14 ;
      RECT 30.39 3.66 30.71 3.98 ;
      RECT 30.365 3.655 30.655 3.885 ;
      RECT 30.36 3.685 30.71 3.86 ;
      RECT 30.19 3.685 30.71 3.855 ;
      RECT 30.39 8.54 30.71 8.83 ;
      RECT 30.365 8.575 30.71 8.805 ;
      RECT 30.19 8.605 30.71 8.775 ;
      RECT 26.845 3.66 27.135 3.89 ;
      RECT 26.845 3.66 27.3 3.845 ;
      RECT 27.16 3.565 27.78 3.705 ;
      RECT 27.55 3.365 27.87 3.625 ;
      RECT 26.23 3.645 26.55 3.905 ;
      RECT 26.23 3.645 26.695 3.89 ;
      RECT 26.555 3.265 26.695 3.89 ;
      RECT 26.555 3.265 26.82 3.405 ;
      RECT 27.085 3.1 27.375 3.33 ;
      RECT 26.68 3.145 27.375 3.285 ;
      RECT 26.125 4.485 26.415 5.01 ;
      RECT 26.11 4.485 26.43 4.745 ;
      RECT 25.85 3.085 26.17 3.345 ;
      RECT 25.85 3.1 26.415 3.33 ;
      RECT 25.125 4.78 25.415 5.01 ;
      RECT 25.32 3.425 25.46 4.965 ;
      RECT 25.365 3.38 25.655 3.61 ;
      RECT 24.96 3.425 25.655 3.565 ;
      RECT 24.96 3.265 25.1 3.565 ;
      RECT 23.5 3.265 25.1 3.405 ;
      RECT 23.41 3.085 23.73 3.345 ;
      RECT 23.41 3.1 23.975 3.345 ;
      RECT 25.12 10.055 25.41 10.285 ;
      RECT 25.18 9.315 25.35 10.285 ;
      RECT 25.1 9.36 25.47 9.71 ;
      RECT 25.1 9.34 25.41 9.71 ;
      RECT 25.12 9.315 25.41 9.71 ;
      RECT 22.52 4.125 25.1 4.265 ;
      RECT 24.885 3.94 25.175 4.17 ;
      RECT 22.445 3.94 23.11 4.17 ;
      RECT 22.79 3.925 23.11 4.265 ;
      RECT 23.79 3.645 24.11 3.905 ;
      RECT 23.79 3.66 24.215 3.89 ;
      RECT 22.43 3.365 22.75 3.625 ;
      RECT 22.925 3.38 23.215 3.61 ;
      RECT 22.43 3.425 23.215 3.565 ;
      RECT 22.55 4.485 22.87 4.745 ;
      RECT 21.71 4.485 22.03 4.745 ;
      RECT 22.55 4.5 22.975 4.73 ;
      RECT 21.71 4.545 22.975 4.685 ;
      RECT 21.245 4.22 21.535 4.45 ;
      RECT 21.32 3.145 21.46 4.45 ;
      RECT 20.97 3.645 21.46 3.905 ;
      RECT 20.725 3.66 21.46 3.89 ;
      RECT 21.725 3.1 22.015 3.33 ;
      RECT 21.32 3.145 22.015 3.285 ;
      RECT 20.485 4.5 20.775 4.73 ;
      RECT 20.485 4.5 20.94 4.685 ;
      RECT 20.8 4.125 20.94 4.685 ;
      RECT 20.44 4.125 20.94 4.265 ;
      RECT 20.44 3.145 20.58 4.265 ;
      RECT 20.23 3.085 20.55 3.345 ;
      RECT 19.99 4.765 20.31 5.025 ;
      RECT 19.285 4.78 19.575 5.01 ;
      RECT 19.285 4.825 20.31 4.965 ;
      RECT 19.36 4.775 19.62 4.965 ;
      RECT 19.75 3.645 20.07 3.905 ;
      RECT 19.75 3.66 20.295 3.89 ;
      RECT 19.75 4.205 20.07 4.465 ;
      RECT 19.75 4.22 20.295 4.45 ;
      RECT 18.79 4.205 19.11 4.465 ;
      RECT 18.88 3.145 19.02 4.465 ;
      RECT 19.285 3.1 19.575 3.33 ;
      RECT 18.88 3.145 19.575 3.285 ;
      RECT 16.54 10.055 16.83 10.285 ;
      RECT 16.6 9.31 16.77 10.285 ;
      RECT 16.51 9.31 16.86 9.6 ;
      RECT 16.135 8.57 16.485 8.86 ;
      RECT 15.995 8.605 16.485 8.775 ;
      RECT 89.69 3.645 90.01 3.905 ;
      RECT 87.25 3.645 87.57 3.905 ;
      RECT 73.365 3.645 73.685 3.905 ;
      RECT 70.925 3.645 71.245 3.905 ;
      RECT 57.04 3.645 57.36 3.905 ;
      RECT 54.6 3.645 54.92 3.905 ;
      RECT 40.715 3.645 41.035 3.905 ;
      RECT 38.275 3.645 38.595 3.905 ;
      RECT 24.39 3.645 24.71 3.905 ;
      RECT 21.95 3.645 22.27 3.905 ;
    LAYER mcon ;
      RECT 98.88 8.6 99.05 8.77 ;
      RECT 98.88 10.08 99.05 10.25 ;
      RECT 98.51 8.23 98.68 8.4 ;
      RECT 98.505 4.06 98.675 4.23 ;
      RECT 97.885 2.205 98.055 2.375 ;
      RECT 97.885 3.685 98.055 3.855 ;
      RECT 97.885 8.605 98.055 8.775 ;
      RECT 97.885 10.085 98.055 10.255 ;
      RECT 97.515 4.055 97.685 4.225 ;
      RECT 97.515 8.235 97.685 8.405 ;
      RECT 96.525 3.315 96.695 3.485 ;
      RECT 96.525 8.975 96.695 9.145 ;
      RECT 96.095 2.205 96.265 2.375 ;
      RECT 96.095 2.945 96.265 3.115 ;
      RECT 96.095 9.345 96.265 9.515 ;
      RECT 96.095 10.085 96.265 10.255 ;
      RECT 95.725 3.685 95.895 3.855 ;
      RECT 95.725 8.605 95.895 8.775 ;
      RECT 92.445 3.13 92.615 3.3 ;
      RECT 92.205 3.69 92.375 3.86 ;
      RECT 91.725 3.69 91.895 3.86 ;
      RECT 91.485 3.13 91.655 3.3 ;
      RECT 91.485 4.81 91.655 4.98 ;
      RECT 90.91 8.975 91.08 9.145 ;
      RECT 90.725 3.41 90.895 3.58 ;
      RECT 90.485 4.81 90.655 4.98 ;
      RECT 90.48 9.345 90.65 9.515 ;
      RECT 90.48 10.085 90.65 10.255 ;
      RECT 90.245 3.97 90.415 4.14 ;
      RECT 89.765 3.69 89.935 3.86 ;
      RECT 89.285 3.69 89.455 3.86 ;
      RECT 89.045 3.13 89.215 3.3 ;
      RECT 88.285 3.41 88.455 3.58 ;
      RECT 88.045 4.53 88.215 4.7 ;
      RECT 87.805 3.97 87.975 4.14 ;
      RECT 87.325 3.69 87.495 3.86 ;
      RECT 87.085 3.13 87.255 3.3 ;
      RECT 87.085 4.53 87.255 4.7 ;
      RECT 86.605 4.25 86.775 4.42 ;
      RECT 86.085 3.69 86.255 3.86 ;
      RECT 85.845 4.53 86.015 4.7 ;
      RECT 85.605 3.13 85.775 3.3 ;
      RECT 85.365 3.69 85.535 3.86 ;
      RECT 85.365 4.25 85.535 4.42 ;
      RECT 84.645 3.13 84.815 3.3 ;
      RECT 84.645 4.81 84.815 4.98 ;
      RECT 84.165 4.25 84.335 4.42 ;
      RECT 82.555 8.6 82.725 8.77 ;
      RECT 82.555 10.08 82.725 10.25 ;
      RECT 82.185 8.23 82.355 8.4 ;
      RECT 82.18 4.06 82.35 4.23 ;
      RECT 81.56 2.205 81.73 2.375 ;
      RECT 81.56 3.685 81.73 3.855 ;
      RECT 81.56 8.605 81.73 8.775 ;
      RECT 81.56 10.085 81.73 10.255 ;
      RECT 81.19 4.055 81.36 4.225 ;
      RECT 81.19 8.235 81.36 8.405 ;
      RECT 80.2 3.315 80.37 3.485 ;
      RECT 80.2 8.975 80.37 9.145 ;
      RECT 79.77 2.205 79.94 2.375 ;
      RECT 79.77 2.945 79.94 3.115 ;
      RECT 79.77 9.345 79.94 9.515 ;
      RECT 79.77 10.085 79.94 10.255 ;
      RECT 79.4 3.685 79.57 3.855 ;
      RECT 79.4 8.605 79.57 8.775 ;
      RECT 76.12 3.13 76.29 3.3 ;
      RECT 75.88 3.69 76.05 3.86 ;
      RECT 75.4 3.69 75.57 3.86 ;
      RECT 75.16 3.13 75.33 3.3 ;
      RECT 75.16 4.81 75.33 4.98 ;
      RECT 74.585 8.975 74.755 9.145 ;
      RECT 74.4 3.41 74.57 3.58 ;
      RECT 74.16 4.81 74.33 4.98 ;
      RECT 74.155 9.345 74.325 9.515 ;
      RECT 74.155 10.085 74.325 10.255 ;
      RECT 73.92 3.97 74.09 4.14 ;
      RECT 73.44 3.69 73.61 3.86 ;
      RECT 72.96 3.69 73.13 3.86 ;
      RECT 72.72 3.13 72.89 3.3 ;
      RECT 71.96 3.41 72.13 3.58 ;
      RECT 71.72 4.53 71.89 4.7 ;
      RECT 71.48 3.97 71.65 4.14 ;
      RECT 71 3.69 71.17 3.86 ;
      RECT 70.76 3.13 70.93 3.3 ;
      RECT 70.76 4.53 70.93 4.7 ;
      RECT 70.28 4.25 70.45 4.42 ;
      RECT 69.76 3.69 69.93 3.86 ;
      RECT 69.52 4.53 69.69 4.7 ;
      RECT 69.28 3.13 69.45 3.3 ;
      RECT 69.04 3.69 69.21 3.86 ;
      RECT 69.04 4.25 69.21 4.42 ;
      RECT 68.32 3.13 68.49 3.3 ;
      RECT 68.32 4.81 68.49 4.98 ;
      RECT 67.84 4.25 68.01 4.42 ;
      RECT 66.23 8.6 66.4 8.77 ;
      RECT 66.23 10.08 66.4 10.25 ;
      RECT 65.86 8.23 66.03 8.4 ;
      RECT 65.855 4.06 66.025 4.23 ;
      RECT 65.235 2.205 65.405 2.375 ;
      RECT 65.235 3.685 65.405 3.855 ;
      RECT 65.235 8.605 65.405 8.775 ;
      RECT 65.235 10.085 65.405 10.255 ;
      RECT 64.865 4.055 65.035 4.225 ;
      RECT 64.865 8.235 65.035 8.405 ;
      RECT 63.875 3.315 64.045 3.485 ;
      RECT 63.875 8.975 64.045 9.145 ;
      RECT 63.445 2.205 63.615 2.375 ;
      RECT 63.445 2.945 63.615 3.115 ;
      RECT 63.445 9.345 63.615 9.515 ;
      RECT 63.445 10.085 63.615 10.255 ;
      RECT 63.075 3.685 63.245 3.855 ;
      RECT 63.075 8.605 63.245 8.775 ;
      RECT 59.795 3.13 59.965 3.3 ;
      RECT 59.555 3.69 59.725 3.86 ;
      RECT 59.075 3.69 59.245 3.86 ;
      RECT 58.835 3.13 59.005 3.3 ;
      RECT 58.835 4.81 59.005 4.98 ;
      RECT 58.26 8.975 58.43 9.145 ;
      RECT 58.075 3.41 58.245 3.58 ;
      RECT 57.835 4.81 58.005 4.98 ;
      RECT 57.83 9.345 58 9.515 ;
      RECT 57.83 10.085 58 10.255 ;
      RECT 57.595 3.97 57.765 4.14 ;
      RECT 57.115 3.69 57.285 3.86 ;
      RECT 56.635 3.69 56.805 3.86 ;
      RECT 56.395 3.13 56.565 3.3 ;
      RECT 55.635 3.41 55.805 3.58 ;
      RECT 55.395 4.53 55.565 4.7 ;
      RECT 55.155 3.97 55.325 4.14 ;
      RECT 54.675 3.69 54.845 3.86 ;
      RECT 54.435 3.13 54.605 3.3 ;
      RECT 54.435 4.53 54.605 4.7 ;
      RECT 53.955 4.25 54.125 4.42 ;
      RECT 53.435 3.69 53.605 3.86 ;
      RECT 53.195 4.53 53.365 4.7 ;
      RECT 52.955 3.13 53.125 3.3 ;
      RECT 52.715 3.69 52.885 3.86 ;
      RECT 52.715 4.25 52.885 4.42 ;
      RECT 51.995 3.13 52.165 3.3 ;
      RECT 51.995 4.81 52.165 4.98 ;
      RECT 51.515 4.25 51.685 4.42 ;
      RECT 49.905 8.6 50.075 8.77 ;
      RECT 49.905 10.08 50.075 10.25 ;
      RECT 49.535 8.23 49.705 8.4 ;
      RECT 49.53 4.06 49.7 4.23 ;
      RECT 48.91 2.205 49.08 2.375 ;
      RECT 48.91 3.685 49.08 3.855 ;
      RECT 48.91 8.605 49.08 8.775 ;
      RECT 48.91 10.085 49.08 10.255 ;
      RECT 48.54 4.055 48.71 4.225 ;
      RECT 48.54 8.235 48.71 8.405 ;
      RECT 47.55 3.315 47.72 3.485 ;
      RECT 47.55 8.975 47.72 9.145 ;
      RECT 47.12 2.205 47.29 2.375 ;
      RECT 47.12 2.945 47.29 3.115 ;
      RECT 47.12 9.345 47.29 9.515 ;
      RECT 47.12 10.085 47.29 10.255 ;
      RECT 46.75 3.685 46.92 3.855 ;
      RECT 46.75 8.605 46.92 8.775 ;
      RECT 43.47 3.13 43.64 3.3 ;
      RECT 43.23 3.69 43.4 3.86 ;
      RECT 42.75 3.69 42.92 3.86 ;
      RECT 42.51 3.13 42.68 3.3 ;
      RECT 42.51 4.81 42.68 4.98 ;
      RECT 41.935 8.975 42.105 9.145 ;
      RECT 41.75 3.41 41.92 3.58 ;
      RECT 41.51 4.81 41.68 4.98 ;
      RECT 41.505 9.345 41.675 9.515 ;
      RECT 41.505 10.085 41.675 10.255 ;
      RECT 41.27 3.97 41.44 4.14 ;
      RECT 40.79 3.69 40.96 3.86 ;
      RECT 40.31 3.69 40.48 3.86 ;
      RECT 40.07 3.13 40.24 3.3 ;
      RECT 39.31 3.41 39.48 3.58 ;
      RECT 39.07 4.53 39.24 4.7 ;
      RECT 38.83 3.97 39 4.14 ;
      RECT 38.35 3.69 38.52 3.86 ;
      RECT 38.11 3.13 38.28 3.3 ;
      RECT 38.11 4.53 38.28 4.7 ;
      RECT 37.63 4.25 37.8 4.42 ;
      RECT 37.11 3.69 37.28 3.86 ;
      RECT 36.87 4.53 37.04 4.7 ;
      RECT 36.63 3.13 36.8 3.3 ;
      RECT 36.39 3.69 36.56 3.86 ;
      RECT 36.39 4.25 36.56 4.42 ;
      RECT 35.67 3.13 35.84 3.3 ;
      RECT 35.67 4.81 35.84 4.98 ;
      RECT 35.19 4.25 35.36 4.42 ;
      RECT 33.58 8.6 33.75 8.77 ;
      RECT 33.58 10.08 33.75 10.25 ;
      RECT 33.21 8.23 33.38 8.4 ;
      RECT 33.205 4.06 33.375 4.23 ;
      RECT 32.585 2.205 32.755 2.375 ;
      RECT 32.585 3.685 32.755 3.855 ;
      RECT 32.585 8.605 32.755 8.775 ;
      RECT 32.585 10.085 32.755 10.255 ;
      RECT 32.215 4.055 32.385 4.225 ;
      RECT 32.215 8.235 32.385 8.405 ;
      RECT 31.225 3.315 31.395 3.485 ;
      RECT 31.225 8.975 31.395 9.145 ;
      RECT 30.795 2.205 30.965 2.375 ;
      RECT 30.795 2.945 30.965 3.115 ;
      RECT 30.795 9.345 30.965 9.515 ;
      RECT 30.795 10.085 30.965 10.255 ;
      RECT 30.425 3.685 30.595 3.855 ;
      RECT 30.425 8.605 30.595 8.775 ;
      RECT 27.145 3.13 27.315 3.3 ;
      RECT 26.905 3.69 27.075 3.86 ;
      RECT 26.425 3.69 26.595 3.86 ;
      RECT 26.185 3.13 26.355 3.3 ;
      RECT 26.185 4.81 26.355 4.98 ;
      RECT 25.61 8.975 25.78 9.145 ;
      RECT 25.425 3.41 25.595 3.58 ;
      RECT 25.185 4.81 25.355 4.98 ;
      RECT 25.18 9.345 25.35 9.515 ;
      RECT 25.18 10.085 25.35 10.255 ;
      RECT 24.945 3.97 25.115 4.14 ;
      RECT 24.465 3.69 24.635 3.86 ;
      RECT 23.985 3.69 24.155 3.86 ;
      RECT 23.745 3.13 23.915 3.3 ;
      RECT 22.985 3.41 23.155 3.58 ;
      RECT 22.745 4.53 22.915 4.7 ;
      RECT 22.505 3.97 22.675 4.14 ;
      RECT 22.025 3.69 22.195 3.86 ;
      RECT 21.785 3.13 21.955 3.3 ;
      RECT 21.785 4.53 21.955 4.7 ;
      RECT 21.305 4.25 21.475 4.42 ;
      RECT 20.785 3.69 20.955 3.86 ;
      RECT 20.545 4.53 20.715 4.7 ;
      RECT 20.305 3.13 20.475 3.3 ;
      RECT 20.065 3.69 20.235 3.86 ;
      RECT 20.065 4.25 20.235 4.42 ;
      RECT 19.345 3.13 19.515 3.3 ;
      RECT 19.345 4.81 19.515 4.98 ;
      RECT 18.865 4.25 19.035 4.42 ;
      RECT 16.6 9.345 16.77 9.515 ;
      RECT 16.6 10.085 16.77 10.255 ;
      RECT 16.23 8.605 16.4 8.775 ;
    LAYER li1 ;
      RECT 98.88 7.3 99.05 8.77 ;
      RECT 98.88 7.3 99.055 8.56 ;
      RECT 98.51 9.25 98.98 9.42 ;
      RECT 98.51 8.23 98.68 9.42 ;
      RECT 98.505 3.04 98.675 4.23 ;
      RECT 98.505 3.04 98.975 3.21 ;
      RECT 97.885 3.895 98.06 5.155 ;
      RECT 97.885 3.685 98.055 5.155 ;
      RECT 97.885 7.305 98.055 8.775 ;
      RECT 97.885 7.305 98.06 8.565 ;
      RECT 97.515 3.035 97.685 4.225 ;
      RECT 97.515 3.035 97.985 3.205 ;
      RECT 97.515 9.255 97.985 9.425 ;
      RECT 97.515 8.235 97.685 9.425 ;
      RECT 96.525 4.015 96.7 5.155 ;
      RECT 96.525 1.865 96.695 5.155 ;
      RECT 96.525 1.865 96.7 2.415 ;
      RECT 96.525 10.045 96.7 10.595 ;
      RECT 96.525 7.305 96.695 10.595 ;
      RECT 96.525 7.305 96.7 8.445 ;
      RECT 96.095 3.895 96.27 5.155 ;
      RECT 96.095 2.945 96.265 5.155 ;
      RECT 96.095 7.305 96.265 9.515 ;
      RECT 96.095 7.305 96.27 8.565 ;
      RECT 95.665 3.925 95.835 5.155 ;
      RECT 95.725 2.145 95.895 4.095 ;
      RECT 95.665 1.865 95.835 2.315 ;
      RECT 95.665 10.145 95.835 10.595 ;
      RECT 95.725 8.365 95.895 10.315 ;
      RECT 95.665 7.305 95.835 8.535 ;
      RECT 95.14 3.895 95.315 5.155 ;
      RECT 95.14 1.865 95.31 5.155 ;
      RECT 95.14 3.365 95.55 3.695 ;
      RECT 95.14 2.525 95.55 2.855 ;
      RECT 95.14 1.865 95.315 2.355 ;
      RECT 95.14 10.105 95.315 10.595 ;
      RECT 95.14 7.305 95.31 10.595 ;
      RECT 95.14 9.605 95.55 9.935 ;
      RECT 95.14 8.765 95.55 9.095 ;
      RECT 95.14 7.305 95.315 8.565 ;
      RECT 92.445 3.03 92.615 3.3 ;
      RECT 92.445 3.03 93.175 3.2 ;
      RECT 92.365 4.42 92.695 4.59 ;
      RECT 91.605 4.25 92.615 4.42 ;
      RECT 91.605 3.77 91.775 4.42 ;
      RECT 91.725 3.69 91.895 4.02 ;
      RECT 90.885 4.42 91.215 4.59 ;
      RECT 88.965 4.42 90.255 4.59 ;
      RECT 90.005 4.335 91.135 4.505 ;
      RECT 90.725 3.41 91.135 3.58 ;
      RECT 90.965 2.95 91.135 3.58 ;
      RECT 90.91 10.045 91.085 10.595 ;
      RECT 90.91 7.305 91.08 10.595 ;
      RECT 90.91 7.305 91.085 8.445 ;
      RECT 90.48 7.305 90.65 9.515 ;
      RECT 90.48 7.305 90.655 8.565 ;
      RECT 89.525 10.105 89.7 10.595 ;
      RECT 89.525 7.305 89.695 10.595 ;
      RECT 89.525 9.605 89.935 9.935 ;
      RECT 89.525 8.765 89.935 9.095 ;
      RECT 89.525 7.305 89.7 8.565 ;
      RECT 88.205 3.77 89.535 3.94 ;
      RECT 89.285 3.69 89.455 3.94 ;
      RECT 88.285 3.37 88.455 3.58 ;
      RECT 88.285 3.37 88.775 3.54 ;
      RECT 86.965 4.53 87.255 4.7 ;
      RECT 86.965 3.77 87.135 4.7 ;
      RECT 86.765 3.77 87.135 3.94 ;
      RECT 85.765 3.77 86.255 3.94 ;
      RECT 86.085 3.69 86.255 3.94 ;
      RECT 85.845 4.53 86.255 4.7 ;
      RECT 86.085 4.34 86.255 4.7 ;
      RECT 84.885 4.25 85.535 4.42 ;
      RECT 84.885 3.69 85.055 4.42 ;
      RECT 84.525 4.81 84.815 4.98 ;
      RECT 84.525 3.77 84.695 4.98 ;
      RECT 84.325 3.77 84.695 3.94 ;
      RECT 82.555 7.3 82.725 8.77 ;
      RECT 82.555 7.3 82.73 8.56 ;
      RECT 82.185 9.25 82.655 9.42 ;
      RECT 82.185 8.23 82.355 9.42 ;
      RECT 82.18 3.04 82.35 4.23 ;
      RECT 82.18 3.04 82.65 3.21 ;
      RECT 81.56 3.895 81.735 5.155 ;
      RECT 81.56 3.685 81.73 5.155 ;
      RECT 81.56 7.305 81.73 8.775 ;
      RECT 81.56 7.305 81.735 8.565 ;
      RECT 81.19 3.035 81.36 4.225 ;
      RECT 81.19 3.035 81.66 3.205 ;
      RECT 81.19 9.255 81.66 9.425 ;
      RECT 81.19 8.235 81.36 9.425 ;
      RECT 80.2 4.015 80.375 5.155 ;
      RECT 80.2 1.865 80.37 5.155 ;
      RECT 80.2 1.865 80.375 2.415 ;
      RECT 80.2 10.045 80.375 10.595 ;
      RECT 80.2 7.305 80.37 10.595 ;
      RECT 80.2 7.305 80.375 8.445 ;
      RECT 79.77 3.895 79.945 5.155 ;
      RECT 79.77 2.945 79.94 5.155 ;
      RECT 79.77 7.305 79.94 9.515 ;
      RECT 79.77 7.305 79.945 8.565 ;
      RECT 79.34 3.925 79.51 5.155 ;
      RECT 79.4 2.145 79.57 4.095 ;
      RECT 79.34 1.865 79.51 2.315 ;
      RECT 79.34 10.145 79.51 10.595 ;
      RECT 79.4 8.365 79.57 10.315 ;
      RECT 79.34 7.305 79.51 8.535 ;
      RECT 78.815 3.895 78.99 5.155 ;
      RECT 78.815 1.865 78.985 5.155 ;
      RECT 78.815 3.365 79.225 3.695 ;
      RECT 78.815 2.525 79.225 2.855 ;
      RECT 78.815 1.865 78.99 2.355 ;
      RECT 78.815 10.105 78.99 10.595 ;
      RECT 78.815 7.305 78.985 10.595 ;
      RECT 78.815 9.605 79.225 9.935 ;
      RECT 78.815 8.765 79.225 9.095 ;
      RECT 78.815 7.305 78.99 8.565 ;
      RECT 76.12 3.03 76.29 3.3 ;
      RECT 76.12 3.03 76.85 3.2 ;
      RECT 76.04 4.42 76.37 4.59 ;
      RECT 75.28 4.25 76.29 4.42 ;
      RECT 75.28 3.77 75.45 4.42 ;
      RECT 75.4 3.69 75.57 4.02 ;
      RECT 74.56 4.42 74.89 4.59 ;
      RECT 72.64 4.42 73.93 4.59 ;
      RECT 73.68 4.335 74.81 4.505 ;
      RECT 74.4 3.41 74.81 3.58 ;
      RECT 74.64 2.95 74.81 3.58 ;
      RECT 74.585 10.045 74.76 10.595 ;
      RECT 74.585 7.305 74.755 10.595 ;
      RECT 74.585 7.305 74.76 8.445 ;
      RECT 74.155 7.305 74.325 9.515 ;
      RECT 74.155 7.305 74.33 8.565 ;
      RECT 73.2 10.105 73.375 10.595 ;
      RECT 73.2 7.305 73.37 10.595 ;
      RECT 73.2 9.605 73.61 9.935 ;
      RECT 73.2 8.765 73.61 9.095 ;
      RECT 73.2 7.305 73.375 8.565 ;
      RECT 71.88 3.77 73.21 3.94 ;
      RECT 72.96 3.69 73.13 3.94 ;
      RECT 71.96 3.37 72.13 3.58 ;
      RECT 71.96 3.37 72.45 3.54 ;
      RECT 70.64 4.53 70.93 4.7 ;
      RECT 70.64 3.77 70.81 4.7 ;
      RECT 70.44 3.77 70.81 3.94 ;
      RECT 69.44 3.77 69.93 3.94 ;
      RECT 69.76 3.69 69.93 3.94 ;
      RECT 69.52 4.53 69.93 4.7 ;
      RECT 69.76 4.34 69.93 4.7 ;
      RECT 68.56 4.25 69.21 4.42 ;
      RECT 68.56 3.69 68.73 4.42 ;
      RECT 68.2 4.81 68.49 4.98 ;
      RECT 68.2 3.77 68.37 4.98 ;
      RECT 68 3.77 68.37 3.94 ;
      RECT 66.23 7.3 66.4 8.77 ;
      RECT 66.23 7.3 66.405 8.56 ;
      RECT 65.86 9.25 66.33 9.42 ;
      RECT 65.86 8.23 66.03 9.42 ;
      RECT 65.855 3.04 66.025 4.23 ;
      RECT 65.855 3.04 66.325 3.21 ;
      RECT 65.235 3.895 65.41 5.155 ;
      RECT 65.235 3.685 65.405 5.155 ;
      RECT 65.235 7.305 65.405 8.775 ;
      RECT 65.235 7.305 65.41 8.565 ;
      RECT 64.865 3.035 65.035 4.225 ;
      RECT 64.865 3.035 65.335 3.205 ;
      RECT 64.865 9.255 65.335 9.425 ;
      RECT 64.865 8.235 65.035 9.425 ;
      RECT 63.875 4.015 64.05 5.155 ;
      RECT 63.875 1.865 64.045 5.155 ;
      RECT 63.875 1.865 64.05 2.415 ;
      RECT 63.875 10.045 64.05 10.595 ;
      RECT 63.875 7.305 64.045 10.595 ;
      RECT 63.875 7.305 64.05 8.445 ;
      RECT 63.445 3.895 63.62 5.155 ;
      RECT 63.445 2.945 63.615 5.155 ;
      RECT 63.445 7.305 63.615 9.515 ;
      RECT 63.445 7.305 63.62 8.565 ;
      RECT 63.015 3.925 63.185 5.155 ;
      RECT 63.075 2.145 63.245 4.095 ;
      RECT 63.015 1.865 63.185 2.315 ;
      RECT 63.015 10.145 63.185 10.595 ;
      RECT 63.075 8.365 63.245 10.315 ;
      RECT 63.015 7.305 63.185 8.535 ;
      RECT 62.49 3.895 62.665 5.155 ;
      RECT 62.49 1.865 62.66 5.155 ;
      RECT 62.49 3.365 62.9 3.695 ;
      RECT 62.49 2.525 62.9 2.855 ;
      RECT 62.49 1.865 62.665 2.355 ;
      RECT 62.49 10.105 62.665 10.595 ;
      RECT 62.49 7.305 62.66 10.595 ;
      RECT 62.49 9.605 62.9 9.935 ;
      RECT 62.49 8.765 62.9 9.095 ;
      RECT 62.49 7.305 62.665 8.565 ;
      RECT 59.795 3.03 59.965 3.3 ;
      RECT 59.795 3.03 60.525 3.2 ;
      RECT 59.715 4.42 60.045 4.59 ;
      RECT 58.955 4.25 59.965 4.42 ;
      RECT 58.955 3.77 59.125 4.42 ;
      RECT 59.075 3.69 59.245 4.02 ;
      RECT 58.235 4.42 58.565 4.59 ;
      RECT 56.315 4.42 57.605 4.59 ;
      RECT 57.355 4.335 58.485 4.505 ;
      RECT 58.075 3.41 58.485 3.58 ;
      RECT 58.315 2.95 58.485 3.58 ;
      RECT 58.26 10.045 58.435 10.595 ;
      RECT 58.26 7.305 58.43 10.595 ;
      RECT 58.26 7.305 58.435 8.445 ;
      RECT 57.83 7.305 58 9.515 ;
      RECT 57.83 7.305 58.005 8.565 ;
      RECT 56.875 10.105 57.05 10.595 ;
      RECT 56.875 7.305 57.045 10.595 ;
      RECT 56.875 9.605 57.285 9.935 ;
      RECT 56.875 8.765 57.285 9.095 ;
      RECT 56.875 7.305 57.05 8.565 ;
      RECT 55.555 3.77 56.885 3.94 ;
      RECT 56.635 3.69 56.805 3.94 ;
      RECT 55.635 3.37 55.805 3.58 ;
      RECT 55.635 3.37 56.125 3.54 ;
      RECT 54.315 4.53 54.605 4.7 ;
      RECT 54.315 3.77 54.485 4.7 ;
      RECT 54.115 3.77 54.485 3.94 ;
      RECT 53.115 3.77 53.605 3.94 ;
      RECT 53.435 3.69 53.605 3.94 ;
      RECT 53.195 4.53 53.605 4.7 ;
      RECT 53.435 4.34 53.605 4.7 ;
      RECT 52.235 4.25 52.885 4.42 ;
      RECT 52.235 3.69 52.405 4.42 ;
      RECT 51.875 4.81 52.165 4.98 ;
      RECT 51.875 3.77 52.045 4.98 ;
      RECT 51.675 3.77 52.045 3.94 ;
      RECT 49.905 7.3 50.075 8.77 ;
      RECT 49.905 7.3 50.08 8.56 ;
      RECT 49.535 9.25 50.005 9.42 ;
      RECT 49.535 8.23 49.705 9.42 ;
      RECT 49.53 3.04 49.7 4.23 ;
      RECT 49.53 3.04 50 3.21 ;
      RECT 48.91 3.895 49.085 5.155 ;
      RECT 48.91 3.685 49.08 5.155 ;
      RECT 48.91 7.305 49.08 8.775 ;
      RECT 48.91 7.305 49.085 8.565 ;
      RECT 48.54 3.035 48.71 4.225 ;
      RECT 48.54 3.035 49.01 3.205 ;
      RECT 48.54 9.255 49.01 9.425 ;
      RECT 48.54 8.235 48.71 9.425 ;
      RECT 47.55 4.015 47.725 5.155 ;
      RECT 47.55 1.865 47.72 5.155 ;
      RECT 47.55 1.865 47.725 2.415 ;
      RECT 47.55 10.045 47.725 10.595 ;
      RECT 47.55 7.305 47.72 10.595 ;
      RECT 47.55 7.305 47.725 8.445 ;
      RECT 47.12 3.895 47.295 5.155 ;
      RECT 47.12 2.945 47.29 5.155 ;
      RECT 47.12 7.305 47.29 9.515 ;
      RECT 47.12 7.305 47.295 8.565 ;
      RECT 46.69 3.925 46.86 5.155 ;
      RECT 46.75 2.145 46.92 4.095 ;
      RECT 46.69 1.865 46.86 2.315 ;
      RECT 46.69 10.145 46.86 10.595 ;
      RECT 46.75 8.365 46.92 10.315 ;
      RECT 46.69 7.305 46.86 8.535 ;
      RECT 46.165 3.895 46.34 5.155 ;
      RECT 46.165 1.865 46.335 5.155 ;
      RECT 46.165 3.365 46.575 3.695 ;
      RECT 46.165 2.525 46.575 2.855 ;
      RECT 46.165 1.865 46.34 2.355 ;
      RECT 46.165 10.105 46.34 10.595 ;
      RECT 46.165 7.305 46.335 10.595 ;
      RECT 46.165 9.605 46.575 9.935 ;
      RECT 46.165 8.765 46.575 9.095 ;
      RECT 46.165 7.305 46.34 8.565 ;
      RECT 43.47 3.03 43.64 3.3 ;
      RECT 43.47 3.03 44.2 3.2 ;
      RECT 43.39 4.42 43.72 4.59 ;
      RECT 42.63 4.25 43.64 4.42 ;
      RECT 42.63 3.77 42.8 4.42 ;
      RECT 42.75 3.69 42.92 4.02 ;
      RECT 41.91 4.42 42.24 4.59 ;
      RECT 39.99 4.42 41.28 4.59 ;
      RECT 41.03 4.335 42.16 4.505 ;
      RECT 41.75 3.41 42.16 3.58 ;
      RECT 41.99 2.95 42.16 3.58 ;
      RECT 41.935 10.045 42.11 10.595 ;
      RECT 41.935 7.305 42.105 10.595 ;
      RECT 41.935 7.305 42.11 8.445 ;
      RECT 41.505 7.305 41.675 9.515 ;
      RECT 41.505 7.305 41.68 8.565 ;
      RECT 40.55 10.105 40.725 10.595 ;
      RECT 40.55 7.305 40.72 10.595 ;
      RECT 40.55 9.605 40.96 9.935 ;
      RECT 40.55 8.765 40.96 9.095 ;
      RECT 40.55 7.305 40.725 8.565 ;
      RECT 39.23 3.77 40.56 3.94 ;
      RECT 40.31 3.69 40.48 3.94 ;
      RECT 39.31 3.37 39.48 3.58 ;
      RECT 39.31 3.37 39.8 3.54 ;
      RECT 37.99 4.53 38.28 4.7 ;
      RECT 37.99 3.77 38.16 4.7 ;
      RECT 37.79 3.77 38.16 3.94 ;
      RECT 36.79 3.77 37.28 3.94 ;
      RECT 37.11 3.69 37.28 3.94 ;
      RECT 36.87 4.53 37.28 4.7 ;
      RECT 37.11 4.34 37.28 4.7 ;
      RECT 35.91 4.25 36.56 4.42 ;
      RECT 35.91 3.69 36.08 4.42 ;
      RECT 35.55 4.81 35.84 4.98 ;
      RECT 35.55 3.77 35.72 4.98 ;
      RECT 35.35 3.77 35.72 3.94 ;
      RECT 33.58 7.3 33.75 8.77 ;
      RECT 33.58 7.3 33.755 8.56 ;
      RECT 33.21 9.25 33.68 9.42 ;
      RECT 33.21 8.23 33.38 9.42 ;
      RECT 33.205 3.04 33.375 4.23 ;
      RECT 33.205 3.04 33.675 3.21 ;
      RECT 32.585 3.895 32.76 5.155 ;
      RECT 32.585 3.685 32.755 5.155 ;
      RECT 32.585 7.305 32.755 8.775 ;
      RECT 32.585 7.305 32.76 8.565 ;
      RECT 32.215 3.035 32.385 4.225 ;
      RECT 32.215 3.035 32.685 3.205 ;
      RECT 32.215 9.255 32.685 9.425 ;
      RECT 32.215 8.235 32.385 9.425 ;
      RECT 31.225 4.015 31.4 5.155 ;
      RECT 31.225 1.865 31.395 5.155 ;
      RECT 31.225 1.865 31.4 2.415 ;
      RECT 31.225 10.045 31.4 10.595 ;
      RECT 31.225 7.305 31.395 10.595 ;
      RECT 31.225 7.305 31.4 8.445 ;
      RECT 30.795 3.895 30.97 5.155 ;
      RECT 30.795 2.945 30.965 5.155 ;
      RECT 30.795 7.305 30.965 9.515 ;
      RECT 30.795 7.305 30.97 8.565 ;
      RECT 30.365 3.925 30.535 5.155 ;
      RECT 30.425 2.145 30.595 4.095 ;
      RECT 30.365 1.865 30.535 2.315 ;
      RECT 30.365 10.145 30.535 10.595 ;
      RECT 30.425 8.365 30.595 10.315 ;
      RECT 30.365 7.305 30.535 8.535 ;
      RECT 29.84 3.895 30.015 5.155 ;
      RECT 29.84 1.865 30.01 5.155 ;
      RECT 29.84 3.365 30.25 3.695 ;
      RECT 29.84 2.525 30.25 2.855 ;
      RECT 29.84 1.865 30.015 2.355 ;
      RECT 29.84 10.105 30.015 10.595 ;
      RECT 29.84 7.305 30.01 10.595 ;
      RECT 29.84 9.605 30.25 9.935 ;
      RECT 29.84 8.765 30.25 9.095 ;
      RECT 29.84 7.305 30.015 8.565 ;
      RECT 27.145 3.03 27.315 3.3 ;
      RECT 27.145 3.03 27.875 3.2 ;
      RECT 27.065 4.42 27.395 4.59 ;
      RECT 26.305 4.25 27.315 4.42 ;
      RECT 26.305 3.77 26.475 4.42 ;
      RECT 26.425 3.69 26.595 4.02 ;
      RECT 25.585 4.42 25.915 4.59 ;
      RECT 23.665 4.42 24.955 4.59 ;
      RECT 24.705 4.335 25.835 4.505 ;
      RECT 25.425 3.41 25.835 3.58 ;
      RECT 25.665 2.95 25.835 3.58 ;
      RECT 25.61 10.045 25.785 10.595 ;
      RECT 25.61 7.305 25.78 10.595 ;
      RECT 25.61 7.305 25.785 8.445 ;
      RECT 25.18 7.305 25.35 9.515 ;
      RECT 25.18 7.305 25.355 8.565 ;
      RECT 24.225 10.105 24.4 10.595 ;
      RECT 24.225 7.305 24.395 10.595 ;
      RECT 24.225 9.605 24.635 9.935 ;
      RECT 24.225 8.765 24.635 9.095 ;
      RECT 24.225 7.305 24.4 8.565 ;
      RECT 22.905 3.77 24.235 3.94 ;
      RECT 23.985 3.69 24.155 3.94 ;
      RECT 22.985 3.37 23.155 3.58 ;
      RECT 22.985 3.37 23.475 3.54 ;
      RECT 21.665 4.53 21.955 4.7 ;
      RECT 21.665 3.77 21.835 4.7 ;
      RECT 21.465 3.77 21.835 3.94 ;
      RECT 20.465 3.77 20.955 3.94 ;
      RECT 20.785 3.69 20.955 3.94 ;
      RECT 20.545 4.53 20.955 4.7 ;
      RECT 20.785 4.34 20.955 4.7 ;
      RECT 19.585 4.25 20.235 4.42 ;
      RECT 19.585 3.69 19.755 4.42 ;
      RECT 19.225 4.81 19.515 4.98 ;
      RECT 19.225 3.77 19.395 4.98 ;
      RECT 19.025 3.77 19.395 3.94 ;
      RECT 16.6 7.305 16.77 9.515 ;
      RECT 16.6 7.305 16.775 8.565 ;
      RECT 16.17 10.145 16.34 10.595 ;
      RECT 16.23 8.365 16.4 10.315 ;
      RECT 16.17 7.305 16.34 8.535 ;
      RECT 15.645 10.105 15.82 10.595 ;
      RECT 15.645 7.305 15.815 10.595 ;
      RECT 15.645 9.605 16.055 9.935 ;
      RECT 15.645 8.765 16.055 9.095 ;
      RECT 15.645 7.305 15.82 8.565 ;
      RECT 98.88 10.08 99.055 10.59 ;
      RECT 97.885 1.865 98.06 2.375 ;
      RECT 97.885 10.085 98.06 10.595 ;
      RECT 96.095 1.865 96.27 2.375 ;
      RECT 96.095 10.085 96.27 10.595 ;
      RECT 92.205 3.69 92.375 4.02 ;
      RECT 91.485 2.95 91.655 3.3 ;
      RECT 91.485 4.68 91.655 5.01 ;
      RECT 90.485 4.68 90.655 5.01 ;
      RECT 90.48 10.085 90.655 10.595 ;
      RECT 90.245 3.69 90.415 4.14 ;
      RECT 89.765 3.69 89.935 4.02 ;
      RECT 89.045 2.95 89.215 3.3 ;
      RECT 88.045 4.34 88.215 4.7 ;
      RECT 87.805 3.69 87.975 4.14 ;
      RECT 87.325 3.69 87.495 4.02 ;
      RECT 87.085 2.95 87.255 3.3 ;
      RECT 86.605 4.25 86.775 4.67 ;
      RECT 85.605 2.95 85.775 3.3 ;
      RECT 85.365 3.69 85.535 4.02 ;
      RECT 84.645 2.95 84.815 3.3 ;
      RECT 84.165 4.25 84.335 4.67 ;
      RECT 82.555 10.08 82.73 10.59 ;
      RECT 81.56 1.865 81.735 2.375 ;
      RECT 81.56 10.085 81.735 10.595 ;
      RECT 79.77 1.865 79.945 2.375 ;
      RECT 79.77 10.085 79.945 10.595 ;
      RECT 75.88 3.69 76.05 4.02 ;
      RECT 75.16 2.95 75.33 3.3 ;
      RECT 75.16 4.68 75.33 5.01 ;
      RECT 74.16 4.68 74.33 5.01 ;
      RECT 74.155 10.085 74.33 10.595 ;
      RECT 73.92 3.69 74.09 4.14 ;
      RECT 73.44 3.69 73.61 4.02 ;
      RECT 72.72 2.95 72.89 3.3 ;
      RECT 71.72 4.34 71.89 4.7 ;
      RECT 71.48 3.69 71.65 4.14 ;
      RECT 71 3.69 71.17 4.02 ;
      RECT 70.76 2.95 70.93 3.3 ;
      RECT 70.28 4.25 70.45 4.67 ;
      RECT 69.28 2.95 69.45 3.3 ;
      RECT 69.04 3.69 69.21 4.02 ;
      RECT 68.32 2.95 68.49 3.3 ;
      RECT 67.84 4.25 68.01 4.67 ;
      RECT 66.23 10.08 66.405 10.59 ;
      RECT 65.235 1.865 65.41 2.375 ;
      RECT 65.235 10.085 65.41 10.595 ;
      RECT 63.445 1.865 63.62 2.375 ;
      RECT 63.445 10.085 63.62 10.595 ;
      RECT 59.555 3.69 59.725 4.02 ;
      RECT 58.835 2.95 59.005 3.3 ;
      RECT 58.835 4.68 59.005 5.01 ;
      RECT 57.835 4.68 58.005 5.01 ;
      RECT 57.83 10.085 58.005 10.595 ;
      RECT 57.595 3.69 57.765 4.14 ;
      RECT 57.115 3.69 57.285 4.02 ;
      RECT 56.395 2.95 56.565 3.3 ;
      RECT 55.395 4.34 55.565 4.7 ;
      RECT 55.155 3.69 55.325 4.14 ;
      RECT 54.675 3.69 54.845 4.02 ;
      RECT 54.435 2.95 54.605 3.3 ;
      RECT 53.955 4.25 54.125 4.67 ;
      RECT 52.955 2.95 53.125 3.3 ;
      RECT 52.715 3.69 52.885 4.02 ;
      RECT 51.995 2.95 52.165 3.3 ;
      RECT 51.515 4.25 51.685 4.67 ;
      RECT 49.905 10.08 50.08 10.59 ;
      RECT 48.91 1.865 49.085 2.375 ;
      RECT 48.91 10.085 49.085 10.595 ;
      RECT 47.12 1.865 47.295 2.375 ;
      RECT 47.12 10.085 47.295 10.595 ;
      RECT 43.23 3.69 43.4 4.02 ;
      RECT 42.51 2.95 42.68 3.3 ;
      RECT 42.51 4.68 42.68 5.01 ;
      RECT 41.51 4.68 41.68 5.01 ;
      RECT 41.505 10.085 41.68 10.595 ;
      RECT 41.27 3.69 41.44 4.14 ;
      RECT 40.79 3.69 40.96 4.02 ;
      RECT 40.07 2.95 40.24 3.3 ;
      RECT 39.07 4.34 39.24 4.7 ;
      RECT 38.83 3.69 39 4.14 ;
      RECT 38.35 3.69 38.52 4.02 ;
      RECT 38.11 2.95 38.28 3.3 ;
      RECT 37.63 4.25 37.8 4.67 ;
      RECT 36.63 2.95 36.8 3.3 ;
      RECT 36.39 3.69 36.56 4.02 ;
      RECT 35.67 2.95 35.84 3.3 ;
      RECT 35.19 4.25 35.36 4.67 ;
      RECT 33.58 10.08 33.755 10.59 ;
      RECT 32.585 1.865 32.76 2.375 ;
      RECT 32.585 10.085 32.76 10.595 ;
      RECT 30.795 1.865 30.97 2.375 ;
      RECT 30.795 10.085 30.97 10.595 ;
      RECT 26.905 3.69 27.075 4.02 ;
      RECT 26.185 2.95 26.355 3.3 ;
      RECT 26.185 4.68 26.355 5.01 ;
      RECT 25.185 4.68 25.355 5.01 ;
      RECT 25.18 10.085 25.355 10.595 ;
      RECT 24.945 3.69 25.115 4.14 ;
      RECT 24.465 3.69 24.635 4.02 ;
      RECT 23.745 2.95 23.915 3.3 ;
      RECT 22.745 4.34 22.915 4.7 ;
      RECT 22.505 3.69 22.675 4.14 ;
      RECT 22.025 3.69 22.195 4.02 ;
      RECT 21.785 2.95 21.955 3.3 ;
      RECT 21.305 4.25 21.475 4.67 ;
      RECT 20.305 2.95 20.475 3.3 ;
      RECT 20.065 3.69 20.235 4.02 ;
      RECT 19.345 2.95 19.515 3.3 ;
      RECT 18.865 4.25 19.035 4.67 ;
      RECT 16.6 10.085 16.775 10.595 ;
  END
END sky130_osu_ring_oscillator_mpr2ea_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2et_8_b0r1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2et_8_b0r1 ;
  SIZE 110.615 BY 12.465 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 35.71 0 36.09 5.27 ;
      LAYER met2 ;
        RECT 35.71 4.89 36.09 5.27 ;
      LAYER li1 ;
        RECT 35.81 1.87 35.985 2.38 ;
        RECT 35.81 3.9 35.985 5.16 ;
        RECT 35.81 3.69 35.98 5.16 ;
      LAYER met1 ;
        RECT 35.725 4.935 36.075 5.225 ;
        RECT 35.75 2.18 36.045 2.41 ;
        RECT 35.75 3.66 36.04 3.89 ;
        RECT 35.81 2.18 35.98 3.89 ;
      LAYER via1 ;
        RECT 35.825 5.005 35.975 5.155 ;
      LAYER via2 ;
        RECT 35.8 4.98 36 5.18 ;
      LAYER mcon ;
        RECT 35.81 3.69 35.98 3.86 ;
        RECT 35.81 2.21 35.98 2.38 ;
        RECT 35.815 4.99 35.985 5.16 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 54.27 0 54.65 5.27 ;
      LAYER met2 ;
        RECT 54.27 4.89 54.65 5.27 ;
      LAYER li1 ;
        RECT 54.37 1.87 54.545 2.38 ;
        RECT 54.37 3.9 54.545 5.16 ;
        RECT 54.37 3.69 54.54 5.16 ;
      LAYER met1 ;
        RECT 54.285 4.935 54.635 5.225 ;
        RECT 54.31 2.18 54.605 2.41 ;
        RECT 54.31 3.66 54.6 3.89 ;
        RECT 54.37 2.18 54.54 3.89 ;
      LAYER via1 ;
        RECT 54.385 5.005 54.535 5.155 ;
      LAYER via2 ;
        RECT 54.36 4.98 54.56 5.18 ;
      LAYER mcon ;
        RECT 54.37 3.69 54.54 3.86 ;
        RECT 54.37 2.21 54.54 2.38 ;
        RECT 54.375 4.99 54.545 5.16 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 72.83 0 73.21 5.27 ;
      LAYER met2 ;
        RECT 72.83 4.89 73.21 5.27 ;
      LAYER li1 ;
        RECT 72.93 1.87 73.105 2.38 ;
        RECT 72.93 3.9 73.105 5.16 ;
        RECT 72.93 3.69 73.1 5.16 ;
      LAYER met1 ;
        RECT 72.845 4.935 73.195 5.225 ;
        RECT 72.87 2.18 73.165 2.41 ;
        RECT 72.87 3.66 73.16 3.89 ;
        RECT 72.93 2.18 73.1 3.89 ;
      LAYER via1 ;
        RECT 72.945 5.005 73.095 5.155 ;
      LAYER via2 ;
        RECT 72.92 4.98 73.12 5.18 ;
      LAYER mcon ;
        RECT 72.93 3.69 73.1 3.86 ;
        RECT 72.93 2.21 73.1 2.38 ;
        RECT 72.935 4.99 73.105 5.16 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 91.39 0 91.77 5.27 ;
      LAYER met2 ;
        RECT 91.39 4.89 91.77 5.27 ;
      LAYER li1 ;
        RECT 91.49 1.87 91.665 2.38 ;
        RECT 91.49 3.9 91.665 5.16 ;
        RECT 91.49 3.69 91.66 5.16 ;
      LAYER met1 ;
        RECT 91.405 4.935 91.755 5.225 ;
        RECT 91.43 2.18 91.725 2.41 ;
        RECT 91.43 3.66 91.72 3.89 ;
        RECT 91.49 2.18 91.66 3.89 ;
      LAYER via1 ;
        RECT 91.505 5.005 91.655 5.155 ;
      LAYER via2 ;
        RECT 91.48 4.98 91.68 5.18 ;
      LAYER mcon ;
        RECT 91.49 3.69 91.66 3.86 ;
        RECT 91.49 2.21 91.66 2.38 ;
        RECT 91.495 4.99 91.665 5.16 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 109.95 0 110.33 5.27 ;
      LAYER met2 ;
        RECT 109.95 4.89 110.33 5.27 ;
      LAYER li1 ;
        RECT 110.05 1.87 110.225 2.38 ;
        RECT 110.05 3.9 110.225 5.16 ;
        RECT 110.05 3.69 110.22 5.16 ;
      LAYER met1 ;
        RECT 109.965 4.935 110.315 5.225 ;
        RECT 109.99 2.18 110.285 2.41 ;
        RECT 109.99 3.66 110.28 3.89 ;
        RECT 110.05 2.18 110.22 3.89 ;
      LAYER via1 ;
        RECT 110.065 5.005 110.215 5.155 ;
      LAYER via2 ;
        RECT 110.04 4.98 110.24 5.18 ;
      LAYER mcon ;
        RECT 110.05 3.69 110.22 3.86 ;
        RECT 110.05 2.21 110.22 2.38 ;
        RECT 110.055 4.99 110.225 5.16 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 31.59 4 31.93 4.35 ;
        RECT 31.58 8.135 31.92 8.485 ;
        RECT 31.665 4 31.835 8.485 ;
      LAYER li1 ;
        RECT 31.66 2.955 31.83 4.225 ;
        RECT 31.66 8.24 31.83 9.51 ;
        RECT 26.045 8.24 26.215 9.51 ;
      LAYER met1 ;
        RECT 25.985 8.235 32.065 8.405 ;
        RECT 31.58 8.235 32.06 8.41 ;
        RECT 31.58 8.135 31.92 8.485 ;
        RECT 25.985 8.235 26.445 8.41 ;
        RECT 25.985 8.21 26.275 8.44 ;
        RECT 31.59 4.055 32.06 4.225 ;
        RECT 31.59 4 31.93 4.35 ;
      LAYER via1 ;
        RECT 31.68 8.235 31.83 8.385 ;
        RECT 31.69 4.1 31.84 4.25 ;
      LAYER mcon ;
        RECT 26.045 8.24 26.215 8.41 ;
        RECT 31.66 8.24 31.83 8.41 ;
        RECT 31.66 4.055 31.83 4.225 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 50.15 4 50.49 4.35 ;
        RECT 50.14 8.135 50.48 8.485 ;
        RECT 50.225 4 50.395 8.485 ;
      LAYER li1 ;
        RECT 50.22 2.955 50.39 4.225 ;
        RECT 50.22 8.24 50.39 9.51 ;
        RECT 44.605 8.24 44.775 9.51 ;
      LAYER met1 ;
        RECT 44.545 8.235 50.625 8.405 ;
        RECT 50.14 8.235 50.62 8.41 ;
        RECT 50.14 8.135 50.48 8.485 ;
        RECT 44.545 8.235 45.005 8.41 ;
        RECT 44.545 8.21 44.835 8.44 ;
        RECT 50.15 4.055 50.62 4.225 ;
        RECT 50.15 4 50.49 4.35 ;
      LAYER via1 ;
        RECT 50.24 8.235 50.39 8.385 ;
        RECT 50.25 4.1 50.4 4.25 ;
      LAYER mcon ;
        RECT 44.605 8.24 44.775 8.41 ;
        RECT 50.22 8.24 50.39 8.41 ;
        RECT 50.22 4.055 50.39 4.225 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 68.71 4 69.05 4.35 ;
        RECT 68.7 8.135 69.04 8.485 ;
        RECT 68.785 4 68.955 8.485 ;
      LAYER li1 ;
        RECT 68.78 2.955 68.95 4.225 ;
        RECT 68.78 8.24 68.95 9.51 ;
        RECT 63.165 8.24 63.335 9.51 ;
      LAYER met1 ;
        RECT 63.105 8.235 69.185 8.405 ;
        RECT 68.7 8.235 69.18 8.41 ;
        RECT 68.7 8.135 69.04 8.485 ;
        RECT 63.105 8.235 63.565 8.41 ;
        RECT 63.105 8.21 63.395 8.44 ;
        RECT 68.71 4.055 69.18 4.225 ;
        RECT 68.71 4 69.05 4.35 ;
      LAYER via1 ;
        RECT 68.8 8.235 68.95 8.385 ;
        RECT 68.81 4.1 68.96 4.25 ;
      LAYER mcon ;
        RECT 63.165 8.24 63.335 8.41 ;
        RECT 68.78 8.24 68.95 8.41 ;
        RECT 68.78 4.055 68.95 4.225 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 87.27 4 87.61 4.35 ;
        RECT 87.26 8.135 87.6 8.485 ;
        RECT 87.345 4 87.515 8.485 ;
      LAYER li1 ;
        RECT 87.34 2.955 87.51 4.225 ;
        RECT 87.34 8.24 87.51 9.51 ;
        RECT 81.725 8.24 81.895 9.51 ;
      LAYER met1 ;
        RECT 81.665 8.235 87.745 8.405 ;
        RECT 87.26 8.235 87.74 8.41 ;
        RECT 87.26 8.135 87.6 8.485 ;
        RECT 81.665 8.235 82.125 8.41 ;
        RECT 81.665 8.21 81.955 8.44 ;
        RECT 87.27 4.055 87.74 4.225 ;
        RECT 87.27 4 87.61 4.35 ;
      LAYER via1 ;
        RECT 87.36 8.235 87.51 8.385 ;
        RECT 87.37 4.1 87.52 4.25 ;
      LAYER mcon ;
        RECT 81.725 8.24 81.895 8.41 ;
        RECT 87.34 8.24 87.51 8.41 ;
        RECT 87.34 4.055 87.51 4.225 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 105.83 4 106.17 4.35 ;
        RECT 105.82 8.135 106.16 8.485 ;
        RECT 105.905 4 106.075 8.485 ;
      LAYER li1 ;
        RECT 105.9 2.955 106.07 4.225 ;
        RECT 105.9 8.24 106.07 9.51 ;
        RECT 100.285 8.24 100.455 9.51 ;
      LAYER met1 ;
        RECT 100.225 8.235 106.305 8.405 ;
        RECT 105.82 8.235 106.3 8.41 ;
        RECT 105.82 8.135 106.16 8.485 ;
        RECT 100.225 8.235 100.685 8.41 ;
        RECT 100.225 8.21 100.515 8.44 ;
        RECT 105.83 4.055 106.3 4.225 ;
        RECT 105.83 4 106.17 4.35 ;
      LAYER via1 ;
        RECT 105.92 8.235 106.07 8.385 ;
        RECT 105.93 4.1 106.08 4.25 ;
      LAYER mcon ;
        RECT 100.285 8.24 100.455 8.41 ;
        RECT 105.9 8.24 106.07 8.41 ;
        RECT 105.9 4.055 106.07 4.225 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 15.23 8.24 15.4 9.51 ;
      LAYER met1 ;
        RECT 15.17 8.24 15.63 8.41 ;
        RECT 15.175 8.205 15.465 8.435 ;
        RECT 15.17 8.21 15.46 8.44 ;
      LAYER mcon ;
        RECT 15.23 8.24 15.4 8.41 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 5.45 110.6 7.05 ;
        RECT 92.785 5.43 110.6 7.05 ;
        RECT 109.625 5.43 109.795 7.765 ;
        RECT 109.62 4.7 109.79 7.05 ;
        RECT 108.635 4.7 108.805 7.765 ;
        RECT 105.72 5.425 108.805 7.05 ;
        RECT 105.89 4.695 106.06 7.77 ;
        RECT 102.875 4.93 103.045 7.05 ;
        RECT 100.435 4.93 100.605 7.05 ;
        RECT 100.275 5.43 100.445 7.77 ;
        RECT 98.475 4.93 98.645 7.05 ;
        RECT 97.515 4.93 97.685 7.05 ;
        RECT 95.555 4.93 95.725 7.05 ;
        RECT 94.555 4.93 94.725 7.05 ;
        RECT 93.595 4.93 93.765 7.05 ;
        RECT 17.8 5.435 110.6 7.05 ;
        RECT 74.225 5.43 92.04 7.05 ;
        RECT 91.065 5.43 91.235 7.765 ;
        RECT 91.06 4.7 91.23 7.05 ;
        RECT 90.075 4.7 90.245 7.765 ;
        RECT 87.16 5.425 90.245 7.05 ;
        RECT 87.33 4.695 87.5 7.77 ;
        RECT 84.315 4.93 84.485 7.05 ;
        RECT 81.875 4.93 82.045 7.05 ;
        RECT 81.715 5.43 81.885 7.77 ;
        RECT 79.915 4.93 80.085 7.05 ;
        RECT 78.955 4.93 79.125 7.05 ;
        RECT 76.995 4.93 77.165 7.05 ;
        RECT 75.995 4.93 76.165 7.05 ;
        RECT 75.035 4.93 75.205 7.05 ;
        RECT 55.665 5.43 73.48 7.05 ;
        RECT 72.505 5.43 72.675 7.765 ;
        RECT 72.5 4.7 72.67 7.05 ;
        RECT 71.515 4.7 71.685 7.765 ;
        RECT 68.6 5.425 71.685 7.05 ;
        RECT 68.77 4.695 68.94 7.77 ;
        RECT 65.755 4.93 65.925 7.05 ;
        RECT 63.315 4.93 63.485 7.05 ;
        RECT 63.155 5.43 63.325 7.77 ;
        RECT 61.355 4.93 61.525 7.05 ;
        RECT 60.395 4.93 60.565 7.05 ;
        RECT 58.435 4.93 58.605 7.05 ;
        RECT 57.435 4.93 57.605 7.05 ;
        RECT 56.475 4.93 56.645 7.05 ;
        RECT 37.105 5.43 54.92 7.05 ;
        RECT 53.945 5.43 54.115 7.765 ;
        RECT 53.94 4.7 54.11 7.05 ;
        RECT 52.955 4.7 53.125 7.765 ;
        RECT 50.04 5.425 53.125 7.05 ;
        RECT 50.21 4.695 50.38 7.77 ;
        RECT 47.195 4.93 47.365 7.05 ;
        RECT 44.755 4.93 44.925 7.05 ;
        RECT 44.595 5.43 44.765 7.77 ;
        RECT 42.795 4.93 42.965 7.05 ;
        RECT 41.835 4.93 42.005 7.05 ;
        RECT 39.875 4.93 40.045 7.05 ;
        RECT 38.875 4.93 39.045 7.05 ;
        RECT 37.915 4.93 38.085 7.05 ;
        RECT 18.545 5.43 36.36 7.05 ;
        RECT 35.385 5.43 35.555 7.765 ;
        RECT 35.38 4.7 35.55 7.05 ;
        RECT 34.395 4.7 34.565 7.765 ;
        RECT 31.48 5.425 34.565 7.05 ;
        RECT 31.65 4.695 31.82 7.77 ;
        RECT 28.635 4.93 28.805 7.05 ;
        RECT 26.195 4.93 26.365 7.05 ;
        RECT 26.035 5.43 26.205 7.77 ;
        RECT 24.235 4.93 24.405 7.05 ;
        RECT 23.275 4.93 23.445 7.05 ;
        RECT 21.315 4.93 21.485 7.05 ;
        RECT 20.315 4.93 20.485 7.05 ;
        RECT 19.355 4.93 19.525 7.05 ;
        RECT 17.035 10.05 17.21 10.6 ;
        RECT 17.035 7.31 17.21 8.45 ;
        RECT 17.035 5.45 17.205 10.6 ;
        RECT 15.22 5.45 15.39 7.77 ;
      LAYER met1 ;
        RECT 17.815 5.425 110.615 7.025 ;
        RECT 0 5.45 110.6 7.05 ;
        RECT 92.785 5.4 104.745 7.05 ;
        RECT 74.225 5.4 86.185 7.05 ;
        RECT 55.665 5.4 67.625 7.05 ;
        RECT 37.105 5.4 49.065 7.05 ;
        RECT 18.545 5.4 30.505 7.05 ;
        RECT 16.975 8.95 17.265 9.18 ;
        RECT 16.805 8.98 17.265 9.15 ;
      LAYER mcon ;
        RECT 17.035 8.98 17.205 9.15 ;
        RECT 17.34 6.84 17.51 7.01 ;
        RECT 18.69 5.43 18.86 5.6 ;
        RECT 19.15 5.43 19.32 5.6 ;
        RECT 19.61 5.43 19.78 5.6 ;
        RECT 20.07 5.43 20.24 5.6 ;
        RECT 20.53 5.43 20.7 5.6 ;
        RECT 20.99 5.43 21.16 5.6 ;
        RECT 21.45 5.43 21.62 5.6 ;
        RECT 21.91 5.43 22.08 5.6 ;
        RECT 22.37 5.43 22.54 5.6 ;
        RECT 22.83 5.43 23 5.6 ;
        RECT 23.29 5.43 23.46 5.6 ;
        RECT 23.75 5.43 23.92 5.6 ;
        RECT 24.21 5.43 24.38 5.6 ;
        RECT 24.67 5.43 24.84 5.6 ;
        RECT 25.13 5.43 25.3 5.6 ;
        RECT 25.59 5.43 25.76 5.6 ;
        RECT 26.05 5.43 26.22 5.6 ;
        RECT 26.51 5.43 26.68 5.6 ;
        RECT 26.97 5.43 27.14 5.6 ;
        RECT 27.43 5.43 27.6 5.6 ;
        RECT 27.89 5.43 28.06 5.6 ;
        RECT 28.155 6.84 28.325 7.01 ;
        RECT 28.35 5.43 28.52 5.6 ;
        RECT 28.81 5.43 28.98 5.6 ;
        RECT 29.27 5.43 29.44 5.6 ;
        RECT 29.73 5.43 29.9 5.6 ;
        RECT 30.19 5.43 30.36 5.6 ;
        RECT 33.77 6.84 33.94 7.01 ;
        RECT 33.77 5.455 33.94 5.625 ;
        RECT 34.475 6.835 34.645 7.005 ;
        RECT 34.475 5.46 34.645 5.63 ;
        RECT 35.46 5.46 35.63 5.63 ;
        RECT 35.465 6.835 35.635 7.005 ;
        RECT 37.25 5.43 37.42 5.6 ;
        RECT 37.71 5.43 37.88 5.6 ;
        RECT 38.17 5.43 38.34 5.6 ;
        RECT 38.63 5.43 38.8 5.6 ;
        RECT 39.09 5.43 39.26 5.6 ;
        RECT 39.55 5.43 39.72 5.6 ;
        RECT 40.01 5.43 40.18 5.6 ;
        RECT 40.47 5.43 40.64 5.6 ;
        RECT 40.93 5.43 41.1 5.6 ;
        RECT 41.39 5.43 41.56 5.6 ;
        RECT 41.85 5.43 42.02 5.6 ;
        RECT 42.31 5.43 42.48 5.6 ;
        RECT 42.77 5.43 42.94 5.6 ;
        RECT 43.23 5.43 43.4 5.6 ;
        RECT 43.69 5.43 43.86 5.6 ;
        RECT 44.15 5.43 44.32 5.6 ;
        RECT 44.61 5.43 44.78 5.6 ;
        RECT 45.07 5.43 45.24 5.6 ;
        RECT 45.53 5.43 45.7 5.6 ;
        RECT 45.99 5.43 46.16 5.6 ;
        RECT 46.45 5.43 46.62 5.6 ;
        RECT 46.715 6.84 46.885 7.01 ;
        RECT 46.91 5.43 47.08 5.6 ;
        RECT 47.37 5.43 47.54 5.6 ;
        RECT 47.83 5.43 48 5.6 ;
        RECT 48.29 5.43 48.46 5.6 ;
        RECT 48.75 5.43 48.92 5.6 ;
        RECT 52.33 6.84 52.5 7.01 ;
        RECT 52.33 5.455 52.5 5.625 ;
        RECT 53.035 6.835 53.205 7.005 ;
        RECT 53.035 5.46 53.205 5.63 ;
        RECT 54.02 5.46 54.19 5.63 ;
        RECT 54.025 6.835 54.195 7.005 ;
        RECT 55.81 5.43 55.98 5.6 ;
        RECT 56.27 5.43 56.44 5.6 ;
        RECT 56.73 5.43 56.9 5.6 ;
        RECT 57.19 5.43 57.36 5.6 ;
        RECT 57.65 5.43 57.82 5.6 ;
        RECT 58.11 5.43 58.28 5.6 ;
        RECT 58.57 5.43 58.74 5.6 ;
        RECT 59.03 5.43 59.2 5.6 ;
        RECT 59.49 5.43 59.66 5.6 ;
        RECT 59.95 5.43 60.12 5.6 ;
        RECT 60.41 5.43 60.58 5.6 ;
        RECT 60.87 5.43 61.04 5.6 ;
        RECT 61.33 5.43 61.5 5.6 ;
        RECT 61.79 5.43 61.96 5.6 ;
        RECT 62.25 5.43 62.42 5.6 ;
        RECT 62.71 5.43 62.88 5.6 ;
        RECT 63.17 5.43 63.34 5.6 ;
        RECT 63.63 5.43 63.8 5.6 ;
        RECT 64.09 5.43 64.26 5.6 ;
        RECT 64.55 5.43 64.72 5.6 ;
        RECT 65.01 5.43 65.18 5.6 ;
        RECT 65.275 6.84 65.445 7.01 ;
        RECT 65.47 5.43 65.64 5.6 ;
        RECT 65.93 5.43 66.1 5.6 ;
        RECT 66.39 5.43 66.56 5.6 ;
        RECT 66.85 5.43 67.02 5.6 ;
        RECT 67.31 5.43 67.48 5.6 ;
        RECT 70.89 6.84 71.06 7.01 ;
        RECT 70.89 5.455 71.06 5.625 ;
        RECT 71.595 6.835 71.765 7.005 ;
        RECT 71.595 5.46 71.765 5.63 ;
        RECT 72.58 5.46 72.75 5.63 ;
        RECT 72.585 6.835 72.755 7.005 ;
        RECT 74.37 5.43 74.54 5.6 ;
        RECT 74.83 5.43 75 5.6 ;
        RECT 75.29 5.43 75.46 5.6 ;
        RECT 75.75 5.43 75.92 5.6 ;
        RECT 76.21 5.43 76.38 5.6 ;
        RECT 76.67 5.43 76.84 5.6 ;
        RECT 77.13 5.43 77.3 5.6 ;
        RECT 77.59 5.43 77.76 5.6 ;
        RECT 78.05 5.43 78.22 5.6 ;
        RECT 78.51 5.43 78.68 5.6 ;
        RECT 78.97 5.43 79.14 5.6 ;
        RECT 79.43 5.43 79.6 5.6 ;
        RECT 79.89 5.43 80.06 5.6 ;
        RECT 80.35 5.43 80.52 5.6 ;
        RECT 80.81 5.43 80.98 5.6 ;
        RECT 81.27 5.43 81.44 5.6 ;
        RECT 81.73 5.43 81.9 5.6 ;
        RECT 82.19 5.43 82.36 5.6 ;
        RECT 82.65 5.43 82.82 5.6 ;
        RECT 83.11 5.43 83.28 5.6 ;
        RECT 83.57 5.43 83.74 5.6 ;
        RECT 83.835 6.84 84.005 7.01 ;
        RECT 84.03 5.43 84.2 5.6 ;
        RECT 84.49 5.43 84.66 5.6 ;
        RECT 84.95 5.43 85.12 5.6 ;
        RECT 85.41 5.43 85.58 5.6 ;
        RECT 85.87 5.43 86.04 5.6 ;
        RECT 89.45 6.84 89.62 7.01 ;
        RECT 89.45 5.455 89.62 5.625 ;
        RECT 90.155 6.835 90.325 7.005 ;
        RECT 90.155 5.46 90.325 5.63 ;
        RECT 91.14 5.46 91.31 5.63 ;
        RECT 91.145 6.835 91.315 7.005 ;
        RECT 92.93 5.43 93.1 5.6 ;
        RECT 93.39 5.43 93.56 5.6 ;
        RECT 93.85 5.43 94.02 5.6 ;
        RECT 94.31 5.43 94.48 5.6 ;
        RECT 94.77 5.43 94.94 5.6 ;
        RECT 95.23 5.43 95.4 5.6 ;
        RECT 95.69 5.43 95.86 5.6 ;
        RECT 96.15 5.43 96.32 5.6 ;
        RECT 96.61 5.43 96.78 5.6 ;
        RECT 97.07 5.43 97.24 5.6 ;
        RECT 97.53 5.43 97.7 5.6 ;
        RECT 97.99 5.43 98.16 5.6 ;
        RECT 98.45 5.43 98.62 5.6 ;
        RECT 98.91 5.43 99.08 5.6 ;
        RECT 99.37 5.43 99.54 5.6 ;
        RECT 99.83 5.43 100 5.6 ;
        RECT 100.29 5.43 100.46 5.6 ;
        RECT 100.75 5.43 100.92 5.6 ;
        RECT 101.21 5.43 101.38 5.6 ;
        RECT 101.67 5.43 101.84 5.6 ;
        RECT 102.13 5.43 102.3 5.6 ;
        RECT 102.395 6.84 102.565 7.01 ;
        RECT 102.59 5.43 102.76 5.6 ;
        RECT 103.05 5.43 103.22 5.6 ;
        RECT 103.51 5.43 103.68 5.6 ;
        RECT 103.97 5.43 104.14 5.6 ;
        RECT 104.43 5.43 104.6 5.6 ;
        RECT 108.01 6.84 108.18 7.01 ;
        RECT 108.01 5.455 108.18 5.625 ;
        RECT 108.715 6.835 108.885 7.005 ;
        RECT 108.715 5.46 108.885 5.63 ;
        RECT 109.7 5.46 109.87 5.63 ;
        RECT 109.705 6.835 109.875 7.005 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 94.4 3.71 95.13 4.04 ;
        RECT 75.84 3.71 76.57 4.04 ;
        RECT 57.28 3.71 58.01 4.04 ;
        RECT 38.72 3.71 39.45 4.04 ;
        RECT 20.16 3.71 20.89 4.04 ;
      LAYER met2 ;
        RECT 96.23 3.715 96.49 4.035 ;
        RECT 94.45 3.805 96.49 3.945 ;
        RECT 94.83 2.295 95.17 2.635 ;
        RECT 94.76 3.69 95.04 4.06 ;
        RECT 94.855 2.295 95.025 4.06 ;
        RECT 94.51 4.275 94.77 4.595 ;
        RECT 94.45 3.805 94.59 4.505 ;
        RECT 77.67 3.715 77.93 4.035 ;
        RECT 75.89 3.805 77.93 3.945 ;
        RECT 76.27 2.295 76.61 2.635 ;
        RECT 76.2 3.69 76.48 4.06 ;
        RECT 76.295 2.295 76.465 4.06 ;
        RECT 75.95 4.275 76.21 4.595 ;
        RECT 75.89 3.805 76.03 4.505 ;
        RECT 59.11 3.715 59.37 4.035 ;
        RECT 57.33 3.805 59.37 3.945 ;
        RECT 57.71 2.295 58.05 2.635 ;
        RECT 57.64 3.69 57.92 4.06 ;
        RECT 57.735 2.295 57.905 4.06 ;
        RECT 57.39 4.275 57.65 4.595 ;
        RECT 57.33 3.805 57.47 4.505 ;
        RECT 40.55 3.715 40.81 4.035 ;
        RECT 38.77 3.805 40.81 3.945 ;
        RECT 39.15 2.295 39.49 2.635 ;
        RECT 39.08 3.69 39.36 4.06 ;
        RECT 39.175 2.295 39.345 4.06 ;
        RECT 38.83 4.275 39.09 4.595 ;
        RECT 38.77 3.805 38.91 4.505 ;
        RECT 21.99 3.715 22.25 4.035 ;
        RECT 20.21 3.805 22.25 3.945 ;
        RECT 20.59 2.295 20.93 2.635 ;
        RECT 20.52 3.69 20.8 4.06 ;
        RECT 20.615 2.295 20.785 4.06 ;
        RECT 20.27 4.275 20.53 4.595 ;
        RECT 20.21 3.805 20.35 4.505 ;
      LAYER li1 ;
        RECT 0.005 10.865 110.605 12.465 ;
        RECT 109.625 10.235 109.795 12.465 ;
        RECT 108.635 10.235 108.805 12.465 ;
        RECT 105.89 10.24 106.06 12.465 ;
        RECT 100.275 10.24 100.445 12.465 ;
        RECT 91.065 10.235 91.235 12.465 ;
        RECT 90.075 10.235 90.245 12.465 ;
        RECT 87.33 10.24 87.5 12.465 ;
        RECT 81.715 10.24 81.885 12.465 ;
        RECT 72.505 10.235 72.675 12.465 ;
        RECT 71.515 10.235 71.685 12.465 ;
        RECT 68.77 10.24 68.94 12.465 ;
        RECT 63.155 10.24 63.325 12.465 ;
        RECT 53.945 10.235 54.115 12.465 ;
        RECT 52.955 10.235 53.125 12.465 ;
        RECT 50.21 10.24 50.38 12.465 ;
        RECT 44.595 10.24 44.765 12.465 ;
        RECT 35.385 10.235 35.555 12.465 ;
        RECT 34.395 10.235 34.565 12.465 ;
        RECT 31.65 10.24 31.82 12.465 ;
        RECT 26.035 10.24 26.205 12.465 ;
        RECT 15.22 10.24 15.39 12.465 ;
        RECT 0.005 0 110.6 1.6 ;
        RECT 109.62 0 109.79 2.23 ;
        RECT 108.635 0 108.805 2.23 ;
        RECT 105.89 0 106.06 2.225 ;
        RECT 92.785 0 104.83 2.88 ;
        RECT 103.835 0 104.005 3.38 ;
        RECT 102.875 0 103.045 3.38 ;
        RECT 101.915 0 102.085 3.38 ;
        RECT 101.395 0 101.565 3.38 ;
        RECT 100.435 0 100.605 3.38 ;
        RECT 99.435 0 99.605 3.38 ;
        RECT 98.475 0 98.645 3.38 ;
        RECT 97.44 0 97.635 2.89 ;
        RECT 96.995 0 97.165 3.38 ;
        RECT 95.075 0 95.335 2.89 ;
        RECT 95.075 0 95.245 3.38 ;
        RECT 93.595 0 93.765 3.38 ;
        RECT 91.06 0 91.23 2.23 ;
        RECT 90.075 0 90.245 2.23 ;
        RECT 87.33 0 87.5 2.225 ;
        RECT 74.225 0 86.27 2.88 ;
        RECT 85.275 0 85.445 3.38 ;
        RECT 84.315 0 84.485 3.38 ;
        RECT 83.355 0 83.525 3.38 ;
        RECT 82.835 0 83.005 3.38 ;
        RECT 81.875 0 82.045 3.38 ;
        RECT 80.875 0 81.045 3.38 ;
        RECT 79.915 0 80.085 3.38 ;
        RECT 78.88 0 79.075 2.89 ;
        RECT 78.435 0 78.605 3.38 ;
        RECT 76.515 0 76.775 2.89 ;
        RECT 76.515 0 76.685 3.38 ;
        RECT 75.035 0 75.205 3.38 ;
        RECT 72.5 0 72.67 2.23 ;
        RECT 71.515 0 71.685 2.23 ;
        RECT 68.77 0 68.94 2.225 ;
        RECT 55.665 0 67.71 2.88 ;
        RECT 66.715 0 66.885 3.38 ;
        RECT 65.755 0 65.925 3.38 ;
        RECT 64.795 0 64.965 3.38 ;
        RECT 64.275 0 64.445 3.38 ;
        RECT 63.315 0 63.485 3.38 ;
        RECT 62.315 0 62.485 3.38 ;
        RECT 61.355 0 61.525 3.38 ;
        RECT 60.32 0 60.515 2.89 ;
        RECT 59.875 0 60.045 3.38 ;
        RECT 57.955 0 58.215 2.89 ;
        RECT 57.955 0 58.125 3.38 ;
        RECT 56.475 0 56.645 3.38 ;
        RECT 53.94 0 54.11 2.23 ;
        RECT 52.955 0 53.125 2.23 ;
        RECT 50.21 0 50.38 2.225 ;
        RECT 37.105 0 49.15 2.88 ;
        RECT 48.155 0 48.325 3.38 ;
        RECT 47.195 0 47.365 3.38 ;
        RECT 46.235 0 46.405 3.38 ;
        RECT 45.715 0 45.885 3.38 ;
        RECT 44.755 0 44.925 3.38 ;
        RECT 43.755 0 43.925 3.38 ;
        RECT 42.795 0 42.965 3.38 ;
        RECT 41.76 0 41.955 2.89 ;
        RECT 41.315 0 41.485 3.38 ;
        RECT 39.395 0 39.655 2.89 ;
        RECT 39.395 0 39.565 3.38 ;
        RECT 37.915 0 38.085 3.38 ;
        RECT 35.38 0 35.55 2.23 ;
        RECT 34.395 0 34.565 2.23 ;
        RECT 31.65 0 31.82 2.225 ;
        RECT 18.545 0 30.59 2.88 ;
        RECT 29.595 0 29.765 3.38 ;
        RECT 28.635 0 28.805 3.38 ;
        RECT 27.675 0 27.845 3.38 ;
        RECT 27.155 0 27.325 3.38 ;
        RECT 26.195 0 26.365 3.38 ;
        RECT 25.195 0 25.365 3.38 ;
        RECT 24.235 0 24.405 3.38 ;
        RECT 23.2 0 23.395 2.89 ;
        RECT 22.755 0 22.925 3.38 ;
        RECT 20.835 0 21.095 2.89 ;
        RECT 20.835 0 21.005 3.38 ;
        RECT 19.355 0 19.525 3.38 ;
        RECT 101.29 8.37 101.46 10.32 ;
        RECT 101.23 10.15 101.4 10.6 ;
        RECT 101.23 7.31 101.4 8.54 ;
        RECT 96.275 3.79 96.445 4.12 ;
        RECT 94.435 4.35 94.725 4.52 ;
        RECT 94.435 3.87 94.605 4.52 ;
        RECT 94.235 3.87 94.605 4.04 ;
        RECT 82.73 8.37 82.9 10.32 ;
        RECT 82.67 10.15 82.84 10.6 ;
        RECT 82.67 7.31 82.84 8.54 ;
        RECT 77.715 3.79 77.885 4.12 ;
        RECT 75.875 4.35 76.165 4.52 ;
        RECT 75.875 3.87 76.045 4.52 ;
        RECT 75.675 3.87 76.045 4.04 ;
        RECT 64.17 8.37 64.34 10.32 ;
        RECT 64.11 10.15 64.28 10.6 ;
        RECT 64.11 7.31 64.28 8.54 ;
        RECT 59.155 3.79 59.325 4.12 ;
        RECT 57.315 4.35 57.605 4.52 ;
        RECT 57.315 3.87 57.485 4.52 ;
        RECT 57.115 3.87 57.485 4.04 ;
        RECT 45.61 8.37 45.78 10.32 ;
        RECT 45.55 10.15 45.72 10.6 ;
        RECT 45.55 7.31 45.72 8.54 ;
        RECT 40.595 3.79 40.765 4.12 ;
        RECT 38.755 4.35 39.045 4.52 ;
        RECT 38.755 3.87 38.925 4.52 ;
        RECT 38.555 3.87 38.925 4.04 ;
        RECT 27.05 8.37 27.22 10.32 ;
        RECT 26.99 10.15 27.16 10.6 ;
        RECT 26.99 7.31 27.16 8.54 ;
        RECT 22.035 3.79 22.205 4.12 ;
        RECT 20.195 4.35 20.485 4.52 ;
        RECT 20.195 3.87 20.365 4.52 ;
        RECT 19.995 3.87 20.365 4.04 ;
      LAYER met1 ;
        RECT 0.005 0 110.605 1.6 ;
        RECT 92.785 0 104.83 2.88 ;
        RECT 92.785 0 104.745 2.91 ;
        RECT 74.225 0 86.27 2.88 ;
        RECT 74.225 0 86.185 2.91 ;
        RECT 55.665 0 67.71 2.88 ;
        RECT 55.665 0 67.625 2.91 ;
        RECT 37.105 0 49.15 2.88 ;
        RECT 37.105 0 49.065 2.91 ;
        RECT 18.545 0 30.59 2.88 ;
        RECT 18.545 0 30.505 2.91 ;
        RECT 0.005 10.865 110.605 12.465 ;
        RECT 101.23 8.58 101.52 8.81 ;
        RECT 100.79 8.605 101.52 8.78 ;
        RECT 100.79 8.605 100.96 12.465 ;
        RECT 82.67 8.58 82.96 8.81 ;
        RECT 82.23 8.605 82.96 8.78 ;
        RECT 82.23 8.605 82.4 12.465 ;
        RECT 64.11 8.58 64.4 8.81 ;
        RECT 63.67 8.605 64.4 8.78 ;
        RECT 63.67 8.605 63.84 12.465 ;
        RECT 45.55 8.58 45.84 8.81 ;
        RECT 45.11 8.605 45.84 8.78 ;
        RECT 45.11 8.605 45.28 12.465 ;
        RECT 26.99 8.58 27.28 8.81 ;
        RECT 26.55 8.605 27.28 8.78 ;
        RECT 26.55 8.605 26.72 12.465 ;
        RECT 96.215 3.665 96.505 4.035 ;
        RECT 95.45 3.665 96.505 3.805 ;
        RECT 94.48 4.305 94.8 4.565 ;
        RECT 77.655 3.665 77.945 4.035 ;
        RECT 76.89 3.665 77.945 3.805 ;
        RECT 75.92 4.305 76.24 4.565 ;
        RECT 59.095 3.665 59.385 4.035 ;
        RECT 58.33 3.665 59.385 3.805 ;
        RECT 57.36 4.305 57.68 4.565 ;
        RECT 40.535 3.665 40.825 4.035 ;
        RECT 39.77 3.665 40.825 3.805 ;
        RECT 38.8 4.305 39.12 4.565 ;
        RECT 21.975 3.665 22.265 4.035 ;
        RECT 21.21 3.665 22.265 3.805 ;
        RECT 20.24 4.305 20.56 4.565 ;
      LAYER via1 ;
        RECT 20.325 4.36 20.475 4.51 ;
        RECT 20.685 2.39 20.835 2.54 ;
        RECT 22.045 3.8 22.195 3.95 ;
        RECT 38.885 4.36 39.035 4.51 ;
        RECT 39.245 2.39 39.395 2.54 ;
        RECT 40.605 3.8 40.755 3.95 ;
        RECT 57.445 4.36 57.595 4.51 ;
        RECT 57.805 2.39 57.955 2.54 ;
        RECT 59.165 3.8 59.315 3.95 ;
        RECT 76.005 4.36 76.155 4.51 ;
        RECT 76.365 2.39 76.515 2.54 ;
        RECT 77.725 3.8 77.875 3.95 ;
        RECT 94.565 4.36 94.715 4.51 ;
        RECT 94.925 2.39 95.075 2.54 ;
        RECT 96.285 3.8 96.435 3.95 ;
      LAYER via2 ;
        RECT 20.56 3.775 20.76 3.975 ;
        RECT 39.12 3.775 39.32 3.975 ;
        RECT 57.68 3.775 57.88 3.975 ;
        RECT 76.24 3.775 76.44 3.975 ;
        RECT 94.8 3.775 95 3.975 ;
      LAYER mcon ;
        RECT 15.3 10.9 15.47 11.07 ;
        RECT 15.98 10.9 16.15 11.07 ;
        RECT 16.66 10.9 16.83 11.07 ;
        RECT 17.34 10.9 17.51 11.07 ;
        RECT 18.69 2.71 18.86 2.88 ;
        RECT 19.15 2.71 19.32 2.88 ;
        RECT 19.61 2.71 19.78 2.88 ;
        RECT 20.07 2.71 20.24 2.88 ;
        RECT 20.315 4.35 20.485 4.52 ;
        RECT 20.53 2.71 20.7 2.88 ;
        RECT 20.99 2.71 21.16 2.88 ;
        RECT 21.45 2.71 21.62 2.88 ;
        RECT 21.91 2.71 22.08 2.88 ;
        RECT 22.035 3.79 22.205 3.96 ;
        RECT 22.37 2.71 22.54 2.88 ;
        RECT 22.83 2.71 23 2.88 ;
        RECT 23.29 2.71 23.46 2.88 ;
        RECT 23.75 2.71 23.92 2.88 ;
        RECT 24.21 2.71 24.38 2.88 ;
        RECT 24.67 2.71 24.84 2.88 ;
        RECT 25.13 2.71 25.3 2.88 ;
        RECT 25.59 2.71 25.76 2.88 ;
        RECT 26.05 2.71 26.22 2.88 ;
        RECT 26.115 10.9 26.285 11.07 ;
        RECT 26.51 2.71 26.68 2.88 ;
        RECT 26.795 10.9 26.965 11.07 ;
        RECT 26.97 2.71 27.14 2.88 ;
        RECT 27.05 8.61 27.22 8.78 ;
        RECT 27.43 2.71 27.6 2.88 ;
        RECT 27.475 10.9 27.645 11.07 ;
        RECT 27.89 2.71 28.06 2.88 ;
        RECT 28.155 10.9 28.325 11.07 ;
        RECT 28.35 2.71 28.52 2.88 ;
        RECT 28.81 2.71 28.98 2.88 ;
        RECT 29.27 2.71 29.44 2.88 ;
        RECT 29.73 2.71 29.9 2.88 ;
        RECT 30.19 2.71 30.36 2.88 ;
        RECT 31.73 10.9 31.9 11.07 ;
        RECT 31.73 1.395 31.9 1.565 ;
        RECT 32.41 10.9 32.58 11.07 ;
        RECT 32.41 1.395 32.58 1.565 ;
        RECT 33.09 10.9 33.26 11.07 ;
        RECT 33.09 1.395 33.26 1.565 ;
        RECT 33.77 10.9 33.94 11.07 ;
        RECT 33.77 1.395 33.94 1.565 ;
        RECT 34.475 10.895 34.645 11.065 ;
        RECT 34.475 1.4 34.645 1.57 ;
        RECT 35.46 1.4 35.63 1.57 ;
        RECT 35.465 10.895 35.635 11.065 ;
        RECT 37.25 2.71 37.42 2.88 ;
        RECT 37.71 2.71 37.88 2.88 ;
        RECT 38.17 2.71 38.34 2.88 ;
        RECT 38.63 2.71 38.8 2.88 ;
        RECT 38.875 4.35 39.045 4.52 ;
        RECT 39.09 2.71 39.26 2.88 ;
        RECT 39.55 2.71 39.72 2.88 ;
        RECT 40.01 2.71 40.18 2.88 ;
        RECT 40.47 2.71 40.64 2.88 ;
        RECT 40.595 3.79 40.765 3.96 ;
        RECT 40.93 2.71 41.1 2.88 ;
        RECT 41.39 2.71 41.56 2.88 ;
        RECT 41.85 2.71 42.02 2.88 ;
        RECT 42.31 2.71 42.48 2.88 ;
        RECT 42.77 2.71 42.94 2.88 ;
        RECT 43.23 2.71 43.4 2.88 ;
        RECT 43.69 2.71 43.86 2.88 ;
        RECT 44.15 2.71 44.32 2.88 ;
        RECT 44.61 2.71 44.78 2.88 ;
        RECT 44.675 10.9 44.845 11.07 ;
        RECT 45.07 2.71 45.24 2.88 ;
        RECT 45.355 10.9 45.525 11.07 ;
        RECT 45.53 2.71 45.7 2.88 ;
        RECT 45.61 8.61 45.78 8.78 ;
        RECT 45.99 2.71 46.16 2.88 ;
        RECT 46.035 10.9 46.205 11.07 ;
        RECT 46.45 2.71 46.62 2.88 ;
        RECT 46.715 10.9 46.885 11.07 ;
        RECT 46.91 2.71 47.08 2.88 ;
        RECT 47.37 2.71 47.54 2.88 ;
        RECT 47.83 2.71 48 2.88 ;
        RECT 48.29 2.71 48.46 2.88 ;
        RECT 48.75 2.71 48.92 2.88 ;
        RECT 50.29 10.9 50.46 11.07 ;
        RECT 50.29 1.395 50.46 1.565 ;
        RECT 50.97 10.9 51.14 11.07 ;
        RECT 50.97 1.395 51.14 1.565 ;
        RECT 51.65 10.9 51.82 11.07 ;
        RECT 51.65 1.395 51.82 1.565 ;
        RECT 52.33 10.9 52.5 11.07 ;
        RECT 52.33 1.395 52.5 1.565 ;
        RECT 53.035 10.895 53.205 11.065 ;
        RECT 53.035 1.4 53.205 1.57 ;
        RECT 54.02 1.4 54.19 1.57 ;
        RECT 54.025 10.895 54.195 11.065 ;
        RECT 55.81 2.71 55.98 2.88 ;
        RECT 56.27 2.71 56.44 2.88 ;
        RECT 56.73 2.71 56.9 2.88 ;
        RECT 57.19 2.71 57.36 2.88 ;
        RECT 57.435 4.35 57.605 4.52 ;
        RECT 57.65 2.71 57.82 2.88 ;
        RECT 58.11 2.71 58.28 2.88 ;
        RECT 58.57 2.71 58.74 2.88 ;
        RECT 59.03 2.71 59.2 2.88 ;
        RECT 59.155 3.79 59.325 3.96 ;
        RECT 59.49 2.71 59.66 2.88 ;
        RECT 59.95 2.71 60.12 2.88 ;
        RECT 60.41 2.71 60.58 2.88 ;
        RECT 60.87 2.71 61.04 2.88 ;
        RECT 61.33 2.71 61.5 2.88 ;
        RECT 61.79 2.71 61.96 2.88 ;
        RECT 62.25 2.71 62.42 2.88 ;
        RECT 62.71 2.71 62.88 2.88 ;
        RECT 63.17 2.71 63.34 2.88 ;
        RECT 63.235 10.9 63.405 11.07 ;
        RECT 63.63 2.71 63.8 2.88 ;
        RECT 63.915 10.9 64.085 11.07 ;
        RECT 64.09 2.71 64.26 2.88 ;
        RECT 64.17 8.61 64.34 8.78 ;
        RECT 64.55 2.71 64.72 2.88 ;
        RECT 64.595 10.9 64.765 11.07 ;
        RECT 65.01 2.71 65.18 2.88 ;
        RECT 65.275 10.9 65.445 11.07 ;
        RECT 65.47 2.71 65.64 2.88 ;
        RECT 65.93 2.71 66.1 2.88 ;
        RECT 66.39 2.71 66.56 2.88 ;
        RECT 66.85 2.71 67.02 2.88 ;
        RECT 67.31 2.71 67.48 2.88 ;
        RECT 68.85 10.9 69.02 11.07 ;
        RECT 68.85 1.395 69.02 1.565 ;
        RECT 69.53 10.9 69.7 11.07 ;
        RECT 69.53 1.395 69.7 1.565 ;
        RECT 70.21 10.9 70.38 11.07 ;
        RECT 70.21 1.395 70.38 1.565 ;
        RECT 70.89 10.9 71.06 11.07 ;
        RECT 70.89 1.395 71.06 1.565 ;
        RECT 71.595 10.895 71.765 11.065 ;
        RECT 71.595 1.4 71.765 1.57 ;
        RECT 72.58 1.4 72.75 1.57 ;
        RECT 72.585 10.895 72.755 11.065 ;
        RECT 74.37 2.71 74.54 2.88 ;
        RECT 74.83 2.71 75 2.88 ;
        RECT 75.29 2.71 75.46 2.88 ;
        RECT 75.75 2.71 75.92 2.88 ;
        RECT 75.995 4.35 76.165 4.52 ;
        RECT 76.21 2.71 76.38 2.88 ;
        RECT 76.67 2.71 76.84 2.88 ;
        RECT 77.13 2.71 77.3 2.88 ;
        RECT 77.59 2.71 77.76 2.88 ;
        RECT 77.715 3.79 77.885 3.96 ;
        RECT 78.05 2.71 78.22 2.88 ;
        RECT 78.51 2.71 78.68 2.88 ;
        RECT 78.97 2.71 79.14 2.88 ;
        RECT 79.43 2.71 79.6 2.88 ;
        RECT 79.89 2.71 80.06 2.88 ;
        RECT 80.35 2.71 80.52 2.88 ;
        RECT 80.81 2.71 80.98 2.88 ;
        RECT 81.27 2.71 81.44 2.88 ;
        RECT 81.73 2.71 81.9 2.88 ;
        RECT 81.795 10.9 81.965 11.07 ;
        RECT 82.19 2.71 82.36 2.88 ;
        RECT 82.475 10.9 82.645 11.07 ;
        RECT 82.65 2.71 82.82 2.88 ;
        RECT 82.73 8.61 82.9 8.78 ;
        RECT 83.11 2.71 83.28 2.88 ;
        RECT 83.155 10.9 83.325 11.07 ;
        RECT 83.57 2.71 83.74 2.88 ;
        RECT 83.835 10.9 84.005 11.07 ;
        RECT 84.03 2.71 84.2 2.88 ;
        RECT 84.49 2.71 84.66 2.88 ;
        RECT 84.95 2.71 85.12 2.88 ;
        RECT 85.41 2.71 85.58 2.88 ;
        RECT 85.87 2.71 86.04 2.88 ;
        RECT 87.41 10.9 87.58 11.07 ;
        RECT 87.41 1.395 87.58 1.565 ;
        RECT 88.09 10.9 88.26 11.07 ;
        RECT 88.09 1.395 88.26 1.565 ;
        RECT 88.77 10.9 88.94 11.07 ;
        RECT 88.77 1.395 88.94 1.565 ;
        RECT 89.45 10.9 89.62 11.07 ;
        RECT 89.45 1.395 89.62 1.565 ;
        RECT 90.155 10.895 90.325 11.065 ;
        RECT 90.155 1.4 90.325 1.57 ;
        RECT 91.14 1.4 91.31 1.57 ;
        RECT 91.145 10.895 91.315 11.065 ;
        RECT 92.93 2.71 93.1 2.88 ;
        RECT 93.39 2.71 93.56 2.88 ;
        RECT 93.85 2.71 94.02 2.88 ;
        RECT 94.31 2.71 94.48 2.88 ;
        RECT 94.555 4.35 94.725 4.52 ;
        RECT 94.77 2.71 94.94 2.88 ;
        RECT 95.23 2.71 95.4 2.88 ;
        RECT 95.69 2.71 95.86 2.88 ;
        RECT 96.15 2.71 96.32 2.88 ;
        RECT 96.275 3.79 96.445 3.96 ;
        RECT 96.61 2.71 96.78 2.88 ;
        RECT 97.07 2.71 97.24 2.88 ;
        RECT 97.53 2.71 97.7 2.88 ;
        RECT 97.99 2.71 98.16 2.88 ;
        RECT 98.45 2.71 98.62 2.88 ;
        RECT 98.91 2.71 99.08 2.88 ;
        RECT 99.37 2.71 99.54 2.88 ;
        RECT 99.83 2.71 100 2.88 ;
        RECT 100.29 2.71 100.46 2.88 ;
        RECT 100.355 10.9 100.525 11.07 ;
        RECT 100.75 2.71 100.92 2.88 ;
        RECT 101.035 10.9 101.205 11.07 ;
        RECT 101.21 2.71 101.38 2.88 ;
        RECT 101.29 8.61 101.46 8.78 ;
        RECT 101.67 2.71 101.84 2.88 ;
        RECT 101.715 10.9 101.885 11.07 ;
        RECT 102.13 2.71 102.3 2.88 ;
        RECT 102.395 10.9 102.565 11.07 ;
        RECT 102.59 2.71 102.76 2.88 ;
        RECT 103.05 2.71 103.22 2.88 ;
        RECT 103.51 2.71 103.68 2.88 ;
        RECT 103.97 2.71 104.14 2.88 ;
        RECT 104.43 2.71 104.6 2.88 ;
        RECT 105.97 10.9 106.14 11.07 ;
        RECT 105.97 1.395 106.14 1.565 ;
        RECT 106.65 10.9 106.82 11.07 ;
        RECT 106.65 1.395 106.82 1.565 ;
        RECT 107.33 10.9 107.5 11.07 ;
        RECT 107.33 1.395 107.5 1.565 ;
        RECT 108.01 10.9 108.18 11.07 ;
        RECT 108.01 1.395 108.18 1.565 ;
        RECT 108.715 10.895 108.885 11.065 ;
        RECT 108.715 1.4 108.885 1.57 ;
        RECT 109.7 1.4 109.87 1.57 ;
        RECT 109.705 10.895 109.875 11.065 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 102.09 4.83 102.645 5.16 ;
      RECT 102.09 3.165 102.39 5.16 ;
      RECT 98.155 4.27 98.71 4.6 ;
      RECT 98.41 3.165 98.71 4.6 ;
      RECT 98.41 3.165 102.39 3.465 ;
      RECT 101.56 9.345 101.935 9.715 ;
      RECT 101.56 9.385 102.565 9.685 ;
      RECT 102.265 5.7 102.565 9.685 ;
      RECT 92.435 5.7 102.565 6.995 ;
      RECT 92.04 5.435 92.88 5.925 ;
      RECT 96.94 3.71 97.24 6.995 ;
      RECT 95.505 4.27 95.805 6.995 ;
      RECT 92.435 3.715 92.735 6.995 ;
      RECT 95.475 4.27 96.205 4.6 ;
      RECT 96.915 3.71 97.645 4.04 ;
      RECT 93.365 3.71 94.095 4.04 ;
      RECT 92.435 3.715 94.095 4.015 ;
      RECT 83.53 4.83 84.085 5.16 ;
      RECT 83.53 3.165 83.83 5.16 ;
      RECT 79.595 4.27 80.15 4.6 ;
      RECT 79.85 3.165 80.15 4.6 ;
      RECT 79.85 3.165 83.83 3.465 ;
      RECT 83 9.345 83.375 9.715 ;
      RECT 83 9.385 84.005 9.685 ;
      RECT 83.705 5.7 84.005 9.685 ;
      RECT 73.875 5.7 84.005 6.995 ;
      RECT 73.48 5.435 74.32 5.925 ;
      RECT 78.38 3.71 78.68 6.995 ;
      RECT 76.945 4.27 77.245 6.995 ;
      RECT 73.875 3.715 74.175 6.995 ;
      RECT 76.915 4.27 77.645 4.6 ;
      RECT 78.355 3.71 79.085 4.04 ;
      RECT 74.805 3.71 75.535 4.04 ;
      RECT 73.875 3.715 75.535 4.015 ;
      RECT 64.97 4.83 65.525 5.16 ;
      RECT 64.97 3.165 65.27 5.16 ;
      RECT 61.035 4.27 61.59 4.6 ;
      RECT 61.29 3.165 61.59 4.6 ;
      RECT 61.29 3.165 65.27 3.465 ;
      RECT 64.44 9.345 64.815 9.715 ;
      RECT 64.44 9.385 65.445 9.685 ;
      RECT 65.145 5.7 65.445 9.685 ;
      RECT 55.315 5.7 65.445 6.995 ;
      RECT 54.92 5.435 55.76 5.925 ;
      RECT 59.82 3.71 60.12 6.995 ;
      RECT 58.385 4.27 58.685 6.995 ;
      RECT 55.315 3.715 55.615 6.995 ;
      RECT 58.355 4.27 59.085 4.6 ;
      RECT 59.795 3.71 60.525 4.04 ;
      RECT 56.245 3.71 56.975 4.04 ;
      RECT 55.315 3.715 56.975 4.015 ;
      RECT 46.41 4.83 46.965 5.16 ;
      RECT 46.41 3.165 46.71 5.16 ;
      RECT 42.475 4.27 43.03 4.6 ;
      RECT 42.73 3.165 43.03 4.6 ;
      RECT 42.73 3.165 46.71 3.465 ;
      RECT 45.88 9.345 46.255 9.715 ;
      RECT 45.88 9.385 46.885 9.685 ;
      RECT 46.585 5.7 46.885 9.685 ;
      RECT 36.755 5.7 46.885 6.995 ;
      RECT 36.36 5.435 37.2 5.925 ;
      RECT 41.26 3.71 41.56 6.995 ;
      RECT 39.825 4.27 40.125 6.995 ;
      RECT 36.755 3.715 37.055 6.995 ;
      RECT 39.795 4.27 40.525 4.6 ;
      RECT 41.235 3.71 41.965 4.04 ;
      RECT 37.685 3.71 38.415 4.04 ;
      RECT 36.755 3.715 38.415 4.015 ;
      RECT 27.85 4.83 28.405 5.16 ;
      RECT 27.85 3.165 28.15 5.16 ;
      RECT 23.915 4.27 24.47 4.6 ;
      RECT 24.17 3.165 24.47 4.6 ;
      RECT 24.17 3.165 28.15 3.465 ;
      RECT 27.32 9.345 27.695 9.715 ;
      RECT 27.32 9.385 28.325 9.685 ;
      RECT 28.025 5.7 28.325 9.685 ;
      RECT 18.195 5.7 28.325 6.995 ;
      RECT 17.8 5.435 18.64 5.925 ;
      RECT 22.7 3.71 23 6.995 ;
      RECT 21.265 4.27 21.565 6.995 ;
      RECT 18.195 3.715 18.495 6.995 ;
      RECT 21.235 4.27 21.965 4.6 ;
      RECT 22.675 3.71 23.405 4.04 ;
      RECT 19.125 3.71 19.855 4.04 ;
      RECT 18.195 3.715 19.855 4.015 ;
      RECT 109.955 7.2 110.335 12.465 ;
      RECT 103.275 3.15 104.005 3.48 ;
      RECT 101.055 4.83 101.785 5.16 ;
      RECT 99.355 4.83 100.085 5.16 ;
      RECT 93.035 4.83 93.765 5.16 ;
      RECT 91.395 7.2 91.775 12.465 ;
      RECT 84.715 3.15 85.445 3.48 ;
      RECT 82.495 4.83 83.225 5.16 ;
      RECT 80.795 4.83 81.525 5.16 ;
      RECT 74.475 4.83 75.205 5.16 ;
      RECT 72.835 7.2 73.215 12.465 ;
      RECT 66.155 3.15 66.885 3.48 ;
      RECT 63.935 4.83 64.665 5.16 ;
      RECT 62.235 4.83 62.965 5.16 ;
      RECT 55.915 4.83 56.645 5.16 ;
      RECT 54.275 7.2 54.655 12.465 ;
      RECT 47.595 3.15 48.325 3.48 ;
      RECT 45.375 4.83 46.105 5.16 ;
      RECT 43.675 4.83 44.405 5.16 ;
      RECT 37.355 4.83 38.085 5.16 ;
      RECT 35.715 7.2 36.095 12.465 ;
      RECT 29.035 3.15 29.765 3.48 ;
      RECT 26.815 4.83 27.545 5.16 ;
      RECT 25.115 4.83 25.845 5.16 ;
      RECT 18.795 4.83 19.525 5.16 ;
    LAYER via2 ;
      RECT 110.045 7.29 110.245 7.49 ;
      RECT 103.34 3.215 103.54 3.415 ;
      RECT 102.38 4.895 102.58 5.095 ;
      RECT 101.645 9.43 101.845 9.63 ;
      RECT 101.38 4.895 101.58 5.095 ;
      RECT 99.42 4.895 99.62 5.095 ;
      RECT 98.22 4.335 98.42 4.535 ;
      RECT 96.98 3.775 97.18 3.975 ;
      RECT 95.54 4.335 95.74 4.535 ;
      RECT 93.58 3.775 93.78 3.975 ;
      RECT 93.1 4.895 93.3 5.095 ;
      RECT 91.485 7.29 91.685 7.49 ;
      RECT 84.78 3.215 84.98 3.415 ;
      RECT 83.82 4.895 84.02 5.095 ;
      RECT 83.085 9.43 83.285 9.63 ;
      RECT 82.82 4.895 83.02 5.095 ;
      RECT 80.86 4.895 81.06 5.095 ;
      RECT 79.66 4.335 79.86 4.535 ;
      RECT 78.42 3.775 78.62 3.975 ;
      RECT 76.98 4.335 77.18 4.535 ;
      RECT 75.02 3.775 75.22 3.975 ;
      RECT 74.54 4.895 74.74 5.095 ;
      RECT 72.925 7.29 73.125 7.49 ;
      RECT 66.22 3.215 66.42 3.415 ;
      RECT 65.26 4.895 65.46 5.095 ;
      RECT 64.525 9.43 64.725 9.63 ;
      RECT 64.26 4.895 64.46 5.095 ;
      RECT 62.3 4.895 62.5 5.095 ;
      RECT 61.1 4.335 61.3 4.535 ;
      RECT 59.86 3.775 60.06 3.975 ;
      RECT 58.42 4.335 58.62 4.535 ;
      RECT 56.46 3.775 56.66 3.975 ;
      RECT 55.98 4.895 56.18 5.095 ;
      RECT 54.365 7.29 54.565 7.49 ;
      RECT 47.66 3.215 47.86 3.415 ;
      RECT 46.7 4.895 46.9 5.095 ;
      RECT 45.965 9.43 46.165 9.63 ;
      RECT 45.7 4.895 45.9 5.095 ;
      RECT 43.74 4.895 43.94 5.095 ;
      RECT 42.54 4.335 42.74 4.535 ;
      RECT 41.3 3.775 41.5 3.975 ;
      RECT 39.86 4.335 40.06 4.535 ;
      RECT 37.9 3.775 38.1 3.975 ;
      RECT 37.42 4.895 37.62 5.095 ;
      RECT 35.805 7.29 36.005 7.49 ;
      RECT 29.1 3.215 29.3 3.415 ;
      RECT 28.14 4.895 28.34 5.095 ;
      RECT 27.405 9.43 27.605 9.63 ;
      RECT 27.14 4.895 27.34 5.095 ;
      RECT 25.18 4.895 25.38 5.095 ;
      RECT 23.98 4.335 24.18 4.535 ;
      RECT 22.74 3.775 22.94 3.975 ;
      RECT 21.3 4.335 21.5 4.535 ;
      RECT 19.34 3.775 19.54 3.975 ;
      RECT 18.86 4.895 19.06 5.095 ;
    LAYER met2 ;
      RECT 16.235 10.69 110.23 10.86 ;
      RECT 110.06 9.565 110.23 10.86 ;
      RECT 16.235 8.545 16.405 10.86 ;
      RECT 110.03 9.565 110.38 9.915 ;
      RECT 16.17 8.545 16.46 8.895 ;
      RECT 106.87 8.51 107.19 8.835 ;
      RECT 106.9 7.985 107.07 8.835 ;
      RECT 106.9 7.985 107.075 8.335 ;
      RECT 106.9 7.985 107.875 8.16 ;
      RECT 107.7 3.26 107.875 8.16 ;
      RECT 107.645 3.26 107.995 3.61 ;
      RECT 107.67 8.945 107.995 9.27 ;
      RECT 106.555 9.035 107.995 9.205 ;
      RECT 106.555 3.69 106.715 9.205 ;
      RECT 106.87 3.66 107.19 3.98 ;
      RECT 106.555 3.69 107.19 3.86 ;
      RECT 101.39 5.43 105.525 5.62 ;
      RECT 105.355 4.44 105.525 5.62 ;
      RECT 105.335 4.445 105.525 5.62 ;
      RECT 101.39 4.81 101.58 5.62 ;
      RECT 101.34 4.81 101.62 5.18 ;
      RECT 105.265 4.445 105.605 4.795 ;
      RECT 91.445 8.945 91.795 9.295 ;
      RECT 102.23 8.9 102.58 9.25 ;
      RECT 91.445 8.975 102.58 9.175 ;
      RECT 101.87 4.275 102.13 4.595 ;
      RECT 101.93 3.155 102.07 4.595 ;
      RECT 101.87 3.155 102.13 3.475 ;
      RECT 100.87 4.835 101.13 5.155 ;
      RECT 100.87 4.25 101.07 5.155 ;
      RECT 100.81 3.155 100.95 4.785 ;
      RECT 100.81 4.25 101.31 4.62 ;
      RECT 100.75 3.155 101.01 3.475 ;
      RECT 100.39 4.835 100.65 5.155 ;
      RECT 100.45 3.245 100.59 5.155 ;
      RECT 100.15 3.245 100.59 3.475 ;
      RECT 100.15 3.155 100.41 3.475 ;
      RECT 99.91 3.715 100.17 4.035 ;
      RECT 99.33 3.805 100.17 3.945 ;
      RECT 99.33 2.865 99.47 3.945 ;
      RECT 95.99 3.155 96.25 3.475 ;
      RECT 95.99 3.245 97.03 3.385 ;
      RECT 96.89 2.865 97.03 3.385 ;
      RECT 96.89 2.865 99.47 3.005 ;
      RECT 99.38 4.81 99.66 5.18 ;
      RECT 99.45 4.365 99.59 5.18 ;
      RECT 99.26 4.25 99.54 4.62 ;
      RECT 98.97 4.365 99.59 4.505 ;
      RECT 98.97 3.155 99.11 4.505 ;
      RECT 98.91 3.155 99.17 3.475 ;
      RECT 98.18 4.25 98.46 4.62 ;
      RECT 98.25 3.155 98.39 4.62 ;
      RECT 98.19 3.155 98.45 3.475 ;
      RECT 97.83 4.835 98.09 5.155 ;
      RECT 97.89 3.245 98.03 5.155 ;
      RECT 97.47 3.155 97.73 3.475 ;
      RECT 97.47 3.245 98.03 3.385 ;
      RECT 95.5 4.25 95.78 4.62 ;
      RECT 97.47 4.275 97.73 4.595 ;
      RECT 95.15 4.275 95.78 4.595 ;
      RECT 95.15 4.365 97.73 4.505 ;
      RECT 96.94 3.69 97.22 4.06 ;
      RECT 96.94 3.715 97.47 4.035 ;
      RECT 94.03 4.275 94.29 4.595 ;
      RECT 94.09 3.155 94.23 4.595 ;
      RECT 94.03 3.155 94.29 3.475 ;
      RECT 93.06 4.81 93.34 5.18 ;
      RECT 93.07 4.555 93.33 5.18 ;
      RECT 88.31 8.51 88.63 8.835 ;
      RECT 88.34 7.985 88.51 8.835 ;
      RECT 88.34 7.985 88.515 8.335 ;
      RECT 88.34 7.985 89.315 8.16 ;
      RECT 89.14 3.26 89.315 8.16 ;
      RECT 89.085 3.26 89.435 3.61 ;
      RECT 89.11 8.945 89.435 9.27 ;
      RECT 87.995 9.035 89.435 9.205 ;
      RECT 87.995 3.69 88.155 9.205 ;
      RECT 88.31 3.66 88.63 3.98 ;
      RECT 87.995 3.69 88.63 3.86 ;
      RECT 82.83 5.43 86.965 5.62 ;
      RECT 86.795 4.44 86.965 5.62 ;
      RECT 86.775 4.445 86.965 5.62 ;
      RECT 82.83 4.81 83.02 5.62 ;
      RECT 82.78 4.81 83.06 5.18 ;
      RECT 86.705 4.445 87.045 4.795 ;
      RECT 72.885 8.945 73.235 9.295 ;
      RECT 83.67 8.9 84.02 9.25 ;
      RECT 72.885 8.975 84.02 9.175 ;
      RECT 83.31 4.275 83.57 4.595 ;
      RECT 83.37 3.155 83.51 4.595 ;
      RECT 83.31 3.155 83.57 3.475 ;
      RECT 82.31 4.835 82.57 5.155 ;
      RECT 82.31 4.25 82.51 5.155 ;
      RECT 82.25 3.155 82.39 4.785 ;
      RECT 82.25 4.25 82.75 4.62 ;
      RECT 82.19 3.155 82.45 3.475 ;
      RECT 81.83 4.835 82.09 5.155 ;
      RECT 81.89 3.245 82.03 5.155 ;
      RECT 81.59 3.245 82.03 3.475 ;
      RECT 81.59 3.155 81.85 3.475 ;
      RECT 81.35 3.715 81.61 4.035 ;
      RECT 80.77 3.805 81.61 3.945 ;
      RECT 80.77 2.865 80.91 3.945 ;
      RECT 77.43 3.155 77.69 3.475 ;
      RECT 77.43 3.245 78.47 3.385 ;
      RECT 78.33 2.865 78.47 3.385 ;
      RECT 78.33 2.865 80.91 3.005 ;
      RECT 80.82 4.81 81.1 5.18 ;
      RECT 80.89 4.365 81.03 5.18 ;
      RECT 80.7 4.25 80.98 4.62 ;
      RECT 80.41 4.365 81.03 4.505 ;
      RECT 80.41 3.155 80.55 4.505 ;
      RECT 80.35 3.155 80.61 3.475 ;
      RECT 79.62 4.25 79.9 4.62 ;
      RECT 79.69 3.155 79.83 4.62 ;
      RECT 79.63 3.155 79.89 3.475 ;
      RECT 79.27 4.835 79.53 5.155 ;
      RECT 79.33 3.245 79.47 5.155 ;
      RECT 78.91 3.155 79.17 3.475 ;
      RECT 78.91 3.245 79.47 3.385 ;
      RECT 76.94 4.25 77.22 4.62 ;
      RECT 78.91 4.275 79.17 4.595 ;
      RECT 76.59 4.275 77.22 4.595 ;
      RECT 76.59 4.365 79.17 4.505 ;
      RECT 78.38 3.69 78.66 4.06 ;
      RECT 78.38 3.715 78.91 4.035 ;
      RECT 75.47 4.275 75.73 4.595 ;
      RECT 75.53 3.155 75.67 4.595 ;
      RECT 75.47 3.155 75.73 3.475 ;
      RECT 74.5 4.81 74.78 5.18 ;
      RECT 74.51 4.555 74.77 5.18 ;
      RECT 69.75 8.51 70.07 8.835 ;
      RECT 69.78 7.985 69.95 8.835 ;
      RECT 69.78 7.985 69.955 8.335 ;
      RECT 69.78 7.985 70.755 8.16 ;
      RECT 70.58 3.26 70.755 8.16 ;
      RECT 70.525 3.26 70.875 3.61 ;
      RECT 70.55 8.945 70.875 9.27 ;
      RECT 69.435 9.035 70.875 9.205 ;
      RECT 69.435 3.69 69.595 9.205 ;
      RECT 69.75 3.66 70.07 3.98 ;
      RECT 69.435 3.69 70.07 3.86 ;
      RECT 64.27 5.43 68.405 5.62 ;
      RECT 68.235 4.44 68.405 5.62 ;
      RECT 68.215 4.445 68.405 5.62 ;
      RECT 64.27 4.81 64.46 5.62 ;
      RECT 64.22 4.81 64.5 5.18 ;
      RECT 68.145 4.445 68.485 4.795 ;
      RECT 54.37 8.95 54.72 9.3 ;
      RECT 65.11 8.905 65.46 9.255 ;
      RECT 54.37 8.98 65.46 9.18 ;
      RECT 64.75 4.275 65.01 4.595 ;
      RECT 64.81 3.155 64.95 4.595 ;
      RECT 64.75 3.155 65.01 3.475 ;
      RECT 63.75 4.835 64.01 5.155 ;
      RECT 63.75 4.25 63.95 5.155 ;
      RECT 63.69 3.155 63.83 4.785 ;
      RECT 63.69 4.25 64.19 4.62 ;
      RECT 63.63 3.155 63.89 3.475 ;
      RECT 63.27 4.835 63.53 5.155 ;
      RECT 63.33 3.245 63.47 5.155 ;
      RECT 63.03 3.245 63.47 3.475 ;
      RECT 63.03 3.155 63.29 3.475 ;
      RECT 62.79 3.715 63.05 4.035 ;
      RECT 62.21 3.805 63.05 3.945 ;
      RECT 62.21 2.865 62.35 3.945 ;
      RECT 58.87 3.155 59.13 3.475 ;
      RECT 58.87 3.245 59.91 3.385 ;
      RECT 59.77 2.865 59.91 3.385 ;
      RECT 59.77 2.865 62.35 3.005 ;
      RECT 62.26 4.81 62.54 5.18 ;
      RECT 62.33 4.365 62.47 5.18 ;
      RECT 62.14 4.25 62.42 4.62 ;
      RECT 61.85 4.365 62.47 4.505 ;
      RECT 61.85 3.155 61.99 4.505 ;
      RECT 61.79 3.155 62.05 3.475 ;
      RECT 61.06 4.25 61.34 4.62 ;
      RECT 61.13 3.155 61.27 4.62 ;
      RECT 61.07 3.155 61.33 3.475 ;
      RECT 60.71 4.835 60.97 5.155 ;
      RECT 60.77 3.245 60.91 5.155 ;
      RECT 60.35 3.155 60.61 3.475 ;
      RECT 60.35 3.245 60.91 3.385 ;
      RECT 58.38 4.25 58.66 4.62 ;
      RECT 60.35 4.275 60.61 4.595 ;
      RECT 58.03 4.275 58.66 4.595 ;
      RECT 58.03 4.365 60.61 4.505 ;
      RECT 59.82 3.69 60.1 4.06 ;
      RECT 59.82 3.715 60.35 4.035 ;
      RECT 56.91 4.275 57.17 4.595 ;
      RECT 56.97 3.155 57.11 4.595 ;
      RECT 56.91 3.155 57.17 3.475 ;
      RECT 55.94 4.81 56.22 5.18 ;
      RECT 55.95 4.555 56.21 5.18 ;
      RECT 51.19 8.51 51.51 8.835 ;
      RECT 51.22 7.985 51.39 8.835 ;
      RECT 51.22 7.985 51.395 8.335 ;
      RECT 51.22 7.985 52.195 8.16 ;
      RECT 52.02 3.26 52.195 8.16 ;
      RECT 51.965 3.26 52.315 3.61 ;
      RECT 51.99 8.945 52.315 9.27 ;
      RECT 50.875 9.035 52.315 9.205 ;
      RECT 50.875 3.69 51.035 9.205 ;
      RECT 51.19 3.66 51.51 3.98 ;
      RECT 50.875 3.69 51.51 3.86 ;
      RECT 45.71 5.43 49.845 5.62 ;
      RECT 49.675 4.44 49.845 5.62 ;
      RECT 49.655 4.445 49.845 5.62 ;
      RECT 45.71 4.81 45.9 5.62 ;
      RECT 45.66 4.81 45.94 5.18 ;
      RECT 49.585 4.445 49.925 4.795 ;
      RECT 35.81 8.945 36.16 9.295 ;
      RECT 46.555 8.9 46.905 9.25 ;
      RECT 35.81 8.975 46.905 9.175 ;
      RECT 46.19 4.275 46.45 4.595 ;
      RECT 46.25 3.155 46.39 4.595 ;
      RECT 46.19 3.155 46.45 3.475 ;
      RECT 45.19 4.835 45.45 5.155 ;
      RECT 45.19 4.25 45.39 5.155 ;
      RECT 45.13 3.155 45.27 4.785 ;
      RECT 45.13 4.25 45.63 4.62 ;
      RECT 45.07 3.155 45.33 3.475 ;
      RECT 44.71 4.835 44.97 5.155 ;
      RECT 44.77 3.245 44.91 5.155 ;
      RECT 44.47 3.245 44.91 3.475 ;
      RECT 44.47 3.155 44.73 3.475 ;
      RECT 44.23 3.715 44.49 4.035 ;
      RECT 43.65 3.805 44.49 3.945 ;
      RECT 43.65 2.865 43.79 3.945 ;
      RECT 40.31 3.155 40.57 3.475 ;
      RECT 40.31 3.245 41.35 3.385 ;
      RECT 41.21 2.865 41.35 3.385 ;
      RECT 41.21 2.865 43.79 3.005 ;
      RECT 43.7 4.81 43.98 5.18 ;
      RECT 43.77 4.365 43.91 5.18 ;
      RECT 43.58 4.25 43.86 4.62 ;
      RECT 43.29 4.365 43.91 4.505 ;
      RECT 43.29 3.155 43.43 4.505 ;
      RECT 43.23 3.155 43.49 3.475 ;
      RECT 42.5 4.25 42.78 4.62 ;
      RECT 42.57 3.155 42.71 4.62 ;
      RECT 42.51 3.155 42.77 3.475 ;
      RECT 42.15 4.835 42.41 5.155 ;
      RECT 42.21 3.245 42.35 5.155 ;
      RECT 41.79 3.155 42.05 3.475 ;
      RECT 41.79 3.245 42.35 3.385 ;
      RECT 39.82 4.25 40.1 4.62 ;
      RECT 41.79 4.275 42.05 4.595 ;
      RECT 39.47 4.275 40.1 4.595 ;
      RECT 39.47 4.365 42.05 4.505 ;
      RECT 41.26 3.69 41.54 4.06 ;
      RECT 41.26 3.715 41.79 4.035 ;
      RECT 38.35 4.275 38.61 4.595 ;
      RECT 38.41 3.155 38.55 4.595 ;
      RECT 38.35 3.155 38.61 3.475 ;
      RECT 37.38 4.81 37.66 5.18 ;
      RECT 37.39 4.555 37.65 5.18 ;
      RECT 32.63 8.51 32.95 8.835 ;
      RECT 32.66 7.985 32.83 8.835 ;
      RECT 32.66 7.985 32.835 8.335 ;
      RECT 32.66 7.985 33.635 8.16 ;
      RECT 33.46 3.26 33.635 8.16 ;
      RECT 33.405 3.26 33.755 3.61 ;
      RECT 33.43 8.945 33.755 9.27 ;
      RECT 32.315 9.035 33.755 9.205 ;
      RECT 32.315 3.69 32.475 9.205 ;
      RECT 32.63 3.66 32.95 3.98 ;
      RECT 32.315 3.69 32.95 3.86 ;
      RECT 27.15 5.43 31.285 5.62 ;
      RECT 31.115 4.44 31.285 5.62 ;
      RECT 31.095 4.445 31.285 5.62 ;
      RECT 27.15 4.81 27.34 5.62 ;
      RECT 27.1 4.81 27.38 5.18 ;
      RECT 31.025 4.445 31.365 4.795 ;
      RECT 16.545 9.285 16.835 9.635 ;
      RECT 16.545 9.34 17.86 9.51 ;
      RECT 17.69 8.975 17.86 9.51 ;
      RECT 27.995 8.895 28.345 9.245 ;
      RECT 17.69 8.975 28.345 9.145 ;
      RECT 27.63 4.275 27.89 4.595 ;
      RECT 27.69 3.155 27.83 4.595 ;
      RECT 27.63 3.155 27.89 3.475 ;
      RECT 26.63 4.835 26.89 5.155 ;
      RECT 26.63 4.25 26.83 5.155 ;
      RECT 26.57 3.155 26.71 4.785 ;
      RECT 26.57 4.25 27.07 4.62 ;
      RECT 26.51 3.155 26.77 3.475 ;
      RECT 26.15 4.835 26.41 5.155 ;
      RECT 26.21 3.245 26.35 5.155 ;
      RECT 25.91 3.245 26.35 3.475 ;
      RECT 25.91 3.155 26.17 3.475 ;
      RECT 25.67 3.715 25.93 4.035 ;
      RECT 25.09 3.805 25.93 3.945 ;
      RECT 25.09 2.865 25.23 3.945 ;
      RECT 21.75 3.155 22.01 3.475 ;
      RECT 21.75 3.245 22.79 3.385 ;
      RECT 22.65 2.865 22.79 3.385 ;
      RECT 22.65 2.865 25.23 3.005 ;
      RECT 25.14 4.81 25.42 5.18 ;
      RECT 25.21 4.365 25.35 5.18 ;
      RECT 25.02 4.25 25.3 4.62 ;
      RECT 24.73 4.365 25.35 4.505 ;
      RECT 24.73 3.155 24.87 4.505 ;
      RECT 24.67 3.155 24.93 3.475 ;
      RECT 23.94 4.25 24.22 4.62 ;
      RECT 24.01 3.155 24.15 4.62 ;
      RECT 23.95 3.155 24.21 3.475 ;
      RECT 23.59 4.835 23.85 5.155 ;
      RECT 23.65 3.245 23.79 5.155 ;
      RECT 23.23 3.155 23.49 3.475 ;
      RECT 23.23 3.245 23.79 3.385 ;
      RECT 21.26 4.25 21.54 4.62 ;
      RECT 23.23 4.275 23.49 4.595 ;
      RECT 20.91 4.275 21.54 4.595 ;
      RECT 20.91 4.365 23.49 4.505 ;
      RECT 22.7 3.69 22.98 4.06 ;
      RECT 22.7 3.715 23.23 4.035 ;
      RECT 19.79 4.275 20.05 4.595 ;
      RECT 19.85 3.155 19.99 4.595 ;
      RECT 19.79 3.155 20.05 3.475 ;
      RECT 18.82 4.81 19.1 5.18 ;
      RECT 18.83 4.555 19.09 5.18 ;
      RECT 109.955 7.2 110.335 7.58 ;
      RECT 103.3 3.13 103.58 3.5 ;
      RECT 102.34 4.81 102.62 5.18 ;
      RECT 101.56 9.345 101.935 9.715 ;
      RECT 93.54 3.69 93.82 4.06 ;
      RECT 91.395 7.2 91.775 7.58 ;
      RECT 84.74 3.13 85.02 3.5 ;
      RECT 83.78 4.81 84.06 5.18 ;
      RECT 83 9.345 83.375 9.715 ;
      RECT 74.98 3.69 75.26 4.06 ;
      RECT 72.835 7.2 73.215 7.58 ;
      RECT 66.18 3.13 66.46 3.5 ;
      RECT 65.22 4.81 65.5 5.18 ;
      RECT 64.44 9.345 64.815 9.715 ;
      RECT 56.42 3.69 56.7 4.06 ;
      RECT 54.275 7.2 54.655 7.58 ;
      RECT 47.62 3.13 47.9 3.5 ;
      RECT 46.66 4.81 46.94 5.18 ;
      RECT 45.88 9.345 46.255 9.715 ;
      RECT 37.86 3.69 38.14 4.06 ;
      RECT 35.715 7.2 36.095 7.58 ;
      RECT 29.06 3.13 29.34 3.5 ;
      RECT 28.1 4.81 28.38 5.18 ;
      RECT 27.32 9.345 27.695 9.715 ;
      RECT 19.3 3.69 19.58 4.06 ;
    LAYER via1 ;
      RECT 110.13 9.665 110.28 9.815 ;
      RECT 110.07 7.315 110.22 7.465 ;
      RECT 107.76 9.03 107.91 9.18 ;
      RECT 107.745 3.36 107.895 3.51 ;
      RECT 106.955 3.745 107.105 3.895 ;
      RECT 106.955 8.615 107.105 8.765 ;
      RECT 105.365 4.545 105.515 4.695 ;
      RECT 103.365 3.24 103.515 3.39 ;
      RECT 102.405 4.92 102.555 5.07 ;
      RECT 102.33 9 102.48 9.15 ;
      RECT 101.925 3.24 102.075 3.39 ;
      RECT 101.925 4.36 102.075 4.51 ;
      RECT 101.67 9.455 101.82 9.605 ;
      RECT 101.405 4.92 101.555 5.07 ;
      RECT 100.925 4.92 101.075 5.07 ;
      RECT 100.805 3.24 100.955 3.39 ;
      RECT 100.445 4.92 100.595 5.07 ;
      RECT 100.205 3.24 100.355 3.39 ;
      RECT 99.965 3.8 100.115 3.95 ;
      RECT 99.445 4.92 99.595 5.07 ;
      RECT 98.965 3.24 99.115 3.39 ;
      RECT 98.245 3.24 98.395 3.39 ;
      RECT 98.245 4.36 98.395 4.51 ;
      RECT 97.885 4.92 98.035 5.07 ;
      RECT 97.525 3.24 97.675 3.39 ;
      RECT 97.525 4.36 97.675 4.51 ;
      RECT 97.265 3.8 97.415 3.95 ;
      RECT 96.045 3.24 96.195 3.39 ;
      RECT 95.205 4.36 95.355 4.51 ;
      RECT 94.085 3.24 94.235 3.39 ;
      RECT 94.085 4.36 94.235 4.51 ;
      RECT 93.605 3.8 93.755 3.95 ;
      RECT 93.125 4.64 93.275 4.79 ;
      RECT 91.545 9.045 91.695 9.195 ;
      RECT 91.51 7.315 91.66 7.465 ;
      RECT 89.2 9.03 89.35 9.18 ;
      RECT 89.185 3.36 89.335 3.51 ;
      RECT 88.395 3.745 88.545 3.895 ;
      RECT 88.395 8.615 88.545 8.765 ;
      RECT 86.805 4.545 86.955 4.695 ;
      RECT 84.805 3.24 84.955 3.39 ;
      RECT 83.845 4.92 83.995 5.07 ;
      RECT 83.77 9 83.92 9.15 ;
      RECT 83.365 3.24 83.515 3.39 ;
      RECT 83.365 4.36 83.515 4.51 ;
      RECT 83.11 9.455 83.26 9.605 ;
      RECT 82.845 4.92 82.995 5.07 ;
      RECT 82.365 4.92 82.515 5.07 ;
      RECT 82.245 3.24 82.395 3.39 ;
      RECT 81.885 4.92 82.035 5.07 ;
      RECT 81.645 3.24 81.795 3.39 ;
      RECT 81.405 3.8 81.555 3.95 ;
      RECT 80.885 4.92 81.035 5.07 ;
      RECT 80.405 3.24 80.555 3.39 ;
      RECT 79.685 3.24 79.835 3.39 ;
      RECT 79.685 4.36 79.835 4.51 ;
      RECT 79.325 4.92 79.475 5.07 ;
      RECT 78.965 3.24 79.115 3.39 ;
      RECT 78.965 4.36 79.115 4.51 ;
      RECT 78.705 3.8 78.855 3.95 ;
      RECT 77.485 3.24 77.635 3.39 ;
      RECT 76.645 4.36 76.795 4.51 ;
      RECT 75.525 3.24 75.675 3.39 ;
      RECT 75.525 4.36 75.675 4.51 ;
      RECT 75.045 3.8 75.195 3.95 ;
      RECT 74.565 4.64 74.715 4.79 ;
      RECT 72.985 9.045 73.135 9.195 ;
      RECT 72.95 7.315 73.1 7.465 ;
      RECT 70.64 9.03 70.79 9.18 ;
      RECT 70.625 3.36 70.775 3.51 ;
      RECT 69.835 3.745 69.985 3.895 ;
      RECT 69.835 8.615 69.985 8.765 ;
      RECT 68.245 4.545 68.395 4.695 ;
      RECT 66.245 3.24 66.395 3.39 ;
      RECT 65.285 4.92 65.435 5.07 ;
      RECT 65.21 9.005 65.36 9.155 ;
      RECT 64.805 3.24 64.955 3.39 ;
      RECT 64.805 4.36 64.955 4.51 ;
      RECT 64.55 9.455 64.7 9.605 ;
      RECT 64.285 4.92 64.435 5.07 ;
      RECT 63.805 4.92 63.955 5.07 ;
      RECT 63.685 3.24 63.835 3.39 ;
      RECT 63.325 4.92 63.475 5.07 ;
      RECT 63.085 3.24 63.235 3.39 ;
      RECT 62.845 3.8 62.995 3.95 ;
      RECT 62.325 4.92 62.475 5.07 ;
      RECT 61.845 3.24 61.995 3.39 ;
      RECT 61.125 3.24 61.275 3.39 ;
      RECT 61.125 4.36 61.275 4.51 ;
      RECT 60.765 4.92 60.915 5.07 ;
      RECT 60.405 3.24 60.555 3.39 ;
      RECT 60.405 4.36 60.555 4.51 ;
      RECT 60.145 3.8 60.295 3.95 ;
      RECT 58.925 3.24 59.075 3.39 ;
      RECT 58.085 4.36 58.235 4.51 ;
      RECT 56.965 3.24 57.115 3.39 ;
      RECT 56.965 4.36 57.115 4.51 ;
      RECT 56.485 3.8 56.635 3.95 ;
      RECT 56.005 4.64 56.155 4.79 ;
      RECT 54.47 9.05 54.62 9.2 ;
      RECT 54.39 7.315 54.54 7.465 ;
      RECT 52.08 9.03 52.23 9.18 ;
      RECT 52.065 3.36 52.215 3.51 ;
      RECT 51.275 3.745 51.425 3.895 ;
      RECT 51.275 8.615 51.425 8.765 ;
      RECT 49.685 4.545 49.835 4.695 ;
      RECT 47.685 3.24 47.835 3.39 ;
      RECT 46.725 4.92 46.875 5.07 ;
      RECT 46.655 9 46.805 9.15 ;
      RECT 46.245 3.24 46.395 3.39 ;
      RECT 46.245 4.36 46.395 4.51 ;
      RECT 45.99 9.455 46.14 9.605 ;
      RECT 45.725 4.92 45.875 5.07 ;
      RECT 45.245 4.92 45.395 5.07 ;
      RECT 45.125 3.24 45.275 3.39 ;
      RECT 44.765 4.92 44.915 5.07 ;
      RECT 44.525 3.24 44.675 3.39 ;
      RECT 44.285 3.8 44.435 3.95 ;
      RECT 43.765 4.92 43.915 5.07 ;
      RECT 43.285 3.24 43.435 3.39 ;
      RECT 42.565 3.24 42.715 3.39 ;
      RECT 42.565 4.36 42.715 4.51 ;
      RECT 42.205 4.92 42.355 5.07 ;
      RECT 41.845 3.24 41.995 3.39 ;
      RECT 41.845 4.36 41.995 4.51 ;
      RECT 41.585 3.8 41.735 3.95 ;
      RECT 40.365 3.24 40.515 3.39 ;
      RECT 39.525 4.36 39.675 4.51 ;
      RECT 38.405 3.24 38.555 3.39 ;
      RECT 38.405 4.36 38.555 4.51 ;
      RECT 37.925 3.8 38.075 3.95 ;
      RECT 37.445 4.64 37.595 4.79 ;
      RECT 35.91 9.045 36.06 9.195 ;
      RECT 35.83 7.315 35.98 7.465 ;
      RECT 33.52 9.03 33.67 9.18 ;
      RECT 33.505 3.36 33.655 3.51 ;
      RECT 32.715 3.745 32.865 3.895 ;
      RECT 32.715 8.615 32.865 8.765 ;
      RECT 31.125 4.545 31.275 4.695 ;
      RECT 29.125 3.24 29.275 3.39 ;
      RECT 28.165 4.92 28.315 5.07 ;
      RECT 28.095 8.995 28.245 9.145 ;
      RECT 27.685 3.24 27.835 3.39 ;
      RECT 27.685 4.36 27.835 4.51 ;
      RECT 27.43 9.455 27.58 9.605 ;
      RECT 27.165 4.92 27.315 5.07 ;
      RECT 26.685 4.92 26.835 5.07 ;
      RECT 26.565 3.24 26.715 3.39 ;
      RECT 26.205 4.92 26.355 5.07 ;
      RECT 25.965 3.24 26.115 3.39 ;
      RECT 25.725 3.8 25.875 3.95 ;
      RECT 25.205 4.92 25.355 5.07 ;
      RECT 24.725 3.24 24.875 3.39 ;
      RECT 24.005 3.24 24.155 3.39 ;
      RECT 24.005 4.36 24.155 4.51 ;
      RECT 23.645 4.92 23.795 5.07 ;
      RECT 23.285 3.24 23.435 3.39 ;
      RECT 23.285 4.36 23.435 4.51 ;
      RECT 23.025 3.8 23.175 3.95 ;
      RECT 21.805 3.24 21.955 3.39 ;
      RECT 20.965 4.36 21.115 4.51 ;
      RECT 19.845 3.24 19.995 3.39 ;
      RECT 19.845 4.36 19.995 4.51 ;
      RECT 19.365 3.8 19.515 3.95 ;
      RECT 18.885 4.64 19.035 4.79 ;
      RECT 16.615 9.385 16.765 9.535 ;
      RECT 16.24 8.645 16.39 8.795 ;
    LAYER met1 ;
      RECT 109.995 10.055 110.29 10.285 ;
      RECT 110.055 9.565 110.23 10.285 ;
      RECT 110.03 9.565 110.38 9.915 ;
      RECT 110.055 8.575 110.225 10.285 ;
      RECT 109.995 8.575 110.285 8.805 ;
      RECT 109.005 10.055 109.3 10.285 ;
      RECT 109.065 8.575 109.235 10.285 ;
      RECT 109.065 8.81 109.855 8.97 ;
      RECT 109.7 8.205 109.855 8.97 ;
      RECT 109.69 8.63 109.855 8.97 ;
      RECT 109.065 8.575 109.295 8.97 ;
      RECT 109.005 8.575 109.295 8.805 ;
      RECT 109.625 8.205 109.915 8.435 ;
      RECT 109.625 8.235 110.085 8.405 ;
      RECT 109.62 4.03 109.91 4.26 ;
      RECT 109.59 3.725 109.78 4.255 ;
      RECT 109.59 4.06 110.08 4.23 ;
      RECT 109.235 3.725 109.78 3.895 ;
      RECT 109.065 2.18 109.235 3.89 ;
      RECT 109.005 3.66 109.295 3.89 ;
      RECT 109.005 2.18 109.3 2.41 ;
      RECT 108.7 4.03 108.87 4.335 ;
      RECT 108.635 4.03 108.925 4.26 ;
      RECT 108.635 4.06 109.095 4.23 ;
      RECT 108.7 2.95 108.865 4.335 ;
      RECT 107.215 2.915 107.505 3.145 ;
      RECT 107.215 2.95 108.865 3.12 ;
      RECT 107.275 2.175 107.445 3.145 ;
      RECT 107.215 2.175 107.505 2.405 ;
      RECT 107.215 10.06 107.505 10.29 ;
      RECT 107.275 9.32 107.445 10.29 ;
      RECT 107.275 9.41 108.865 9.58 ;
      RECT 108.695 8.205 108.865 9.58 ;
      RECT 107.215 9.32 107.505 9.55 ;
      RECT 108.635 8.205 108.925 8.435 ;
      RECT 108.635 8.235 109.095 8.405 ;
      RECT 105.265 4.445 105.605 4.795 ;
      RECT 105.355 3.32 105.525 4.795 ;
      RECT 107.645 3.26 107.995 3.61 ;
      RECT 105.355 3.32 107.995 3.49 ;
      RECT 107.475 3.315 107.995 3.49 ;
      RECT 107.67 8.945 107.995 9.27 ;
      RECT 102.23 8.9 102.58 9.25 ;
      RECT 107.645 8.95 107.995 9.18 ;
      RECT 102.03 8.95 102.58 9.18 ;
      RECT 107.475 8.975 107.995 9.15 ;
      RECT 101.86 8.975 102.58 9.15 ;
      RECT 101.86 8.975 107.995 9.145 ;
      RECT 106.87 3.66 107.19 3.98 ;
      RECT 106.845 3.655 107.135 3.885 ;
      RECT 106.84 3.685 107.19 3.86 ;
      RECT 106.67 3.685 107.19 3.855 ;
      RECT 106.87 8.545 107.19 8.835 ;
      RECT 106.845 8.58 107.19 8.81 ;
      RECT 106.67 8.61 107.19 8.78 ;
      RECT 102.32 4.865 102.64 5.125 ;
      RECT 103.61 4.04 103.75 4.9 ;
      RECT 102.41 4.76 103.75 4.9 ;
      RECT 102.41 4.32 102.55 5.125 ;
      RECT 102.335 4.32 102.625 4.55 ;
      RECT 103.535 4.04 103.825 4.27 ;
      RECT 103.055 4.32 103.345 4.55 ;
      RECT 103.25 3.245 103.39 4.505 ;
      RECT 103.28 3.185 103.6 3.445 ;
      RECT 99.88 3.745 100.2 4.005 ;
      RECT 102.575 3.76 102.865 3.99 ;
      RECT 99.97 3.665 102.79 3.805 ;
      RECT 101.84 3.185 102.16 3.445 ;
      RECT 102.335 3.2 102.625 3.43 ;
      RECT 101.84 3.245 102.625 3.385 ;
      RECT 101.84 4.305 102.16 4.565 ;
      RECT 101.84 4.085 102.07 4.565 ;
      RECT 101.335 4.04 101.625 4.27 ;
      RECT 101.335 4.085 102.07 4.225 ;
      RECT 101.6 10.06 101.89 10.29 ;
      RECT 101.66 9.32 101.83 10.29 ;
      RECT 101.56 9.345 101.94 9.715 ;
      RECT 101.6 9.32 101.89 9.715 ;
      RECT 100.36 4.865 100.68 5.125 ;
      RECT 99.895 4.88 100.185 5.11 ;
      RECT 99.895 4.925 100.68 5.065 ;
      RECT 98.655 3.76 98.945 3.99 ;
      RECT 98.655 3.805 99.59 3.945 ;
      RECT 99.45 3.245 99.59 3.945 ;
      RECT 100.12 3.185 100.44 3.445 ;
      RECT 99.895 3.2 100.44 3.43 ;
      RECT 99.45 3.245 100.44 3.385 ;
      RECT 97.8 4.865 98.12 5.125 ;
      RECT 97.8 4.925 98.87 5.065 ;
      RECT 98.73 4.365 98.87 5.065 ;
      RECT 99.895 4.32 100.185 4.55 ;
      RECT 98.73 4.365 100.185 4.505 ;
      RECT 98.16 3.185 98.48 3.445 ;
      RECT 97.935 3.2 98.48 3.43 ;
      RECT 97.18 3.745 97.5 4.005 ;
      RECT 98.175 3.76 98.465 3.99 ;
      RECT 96.935 3.76 97.5 3.99 ;
      RECT 96.935 3.805 98.465 3.945 ;
      RECT 96.455 4.32 96.745 4.55 ;
      RECT 96.65 3.245 96.79 4.505 ;
      RECT 97.44 3.185 97.76 3.445 ;
      RECT 96.455 3.2 96.745 3.43 ;
      RECT 96.455 3.245 97.76 3.385 ;
      RECT 96.05 4.76 97.15 4.9 ;
      RECT 96.935 4.6 97.225 4.83 ;
      RECT 95.975 4.6 96.265 4.83 ;
      RECT 95.96 3.185 96.28 3.445 ;
      RECT 94 3.185 94.32 3.445 ;
      RECT 94 3.245 96.28 3.385 ;
      RECT 95.12 4.305 95.44 4.565 ;
      RECT 95.12 4.305 95.95 4.445 ;
      RECT 95.735 4.04 95.95 4.445 ;
      RECT 95.735 4.04 96.025 4.27 ;
      RECT 93.52 3.745 93.84 4.005 ;
      RECT 94.93 3.76 95.22 3.99 ;
      RECT 93.52 3.76 94.065 3.99 ;
      RECT 93.52 3.845 94.47 3.985 ;
      RECT 94.33 3.665 94.47 3.985 ;
      RECT 94.83 3.76 95.22 3.945 ;
      RECT 94.33 3.665 94.97 3.805 ;
      RECT 93.04 4.555 93.36 4.97 ;
      RECT 93.12 3.2 93.275 4.97 ;
      RECT 93.055 3.2 93.345 3.43 ;
      RECT 91.435 10.055 91.73 10.285 ;
      RECT 91.495 8.575 91.665 10.285 ;
      RECT 91.445 8.945 91.795 9.295 ;
      RECT 91.435 8.575 91.725 8.805 ;
      RECT 90.445 10.055 90.74 10.285 ;
      RECT 90.505 8.575 90.675 10.285 ;
      RECT 90.505 8.81 91.295 8.97 ;
      RECT 91.14 8.205 91.295 8.97 ;
      RECT 91.13 8.63 91.295 8.97 ;
      RECT 90.505 8.575 90.735 8.97 ;
      RECT 90.445 8.575 90.735 8.805 ;
      RECT 91.065 8.205 91.355 8.435 ;
      RECT 91.065 8.235 91.525 8.405 ;
      RECT 91.06 4.03 91.35 4.26 ;
      RECT 91.03 3.725 91.22 4.255 ;
      RECT 91.03 4.06 91.52 4.23 ;
      RECT 90.675 3.725 91.22 3.895 ;
      RECT 90.505 2.18 90.675 3.89 ;
      RECT 90.445 3.66 90.735 3.89 ;
      RECT 90.445 2.18 90.74 2.41 ;
      RECT 90.14 4.03 90.31 4.335 ;
      RECT 90.075 4.03 90.365 4.26 ;
      RECT 90.075 4.06 90.535 4.23 ;
      RECT 90.14 2.95 90.305 4.335 ;
      RECT 88.655 2.915 88.945 3.145 ;
      RECT 88.655 2.95 90.305 3.12 ;
      RECT 88.715 2.175 88.885 3.145 ;
      RECT 88.655 2.175 88.945 2.405 ;
      RECT 88.655 10.06 88.945 10.29 ;
      RECT 88.715 9.32 88.885 10.29 ;
      RECT 88.715 9.41 90.305 9.58 ;
      RECT 90.135 8.205 90.305 9.58 ;
      RECT 88.655 9.32 88.945 9.55 ;
      RECT 90.075 8.205 90.365 8.435 ;
      RECT 90.075 8.235 90.535 8.405 ;
      RECT 86.705 4.445 87.045 4.795 ;
      RECT 86.795 3.32 86.965 4.795 ;
      RECT 89.085 3.26 89.435 3.61 ;
      RECT 86.795 3.32 89.435 3.49 ;
      RECT 88.915 3.315 89.435 3.49 ;
      RECT 89.11 8.945 89.435 9.27 ;
      RECT 83.67 8.9 84.02 9.25 ;
      RECT 89.085 8.95 89.435 9.18 ;
      RECT 83.47 8.95 84.02 9.18 ;
      RECT 88.915 8.975 89.435 9.15 ;
      RECT 83.3 8.975 84.02 9.15 ;
      RECT 83.3 8.975 89.435 9.145 ;
      RECT 88.31 3.66 88.63 3.98 ;
      RECT 88.285 3.655 88.575 3.885 ;
      RECT 88.28 3.685 88.63 3.86 ;
      RECT 88.11 3.685 88.63 3.855 ;
      RECT 88.31 8.545 88.63 8.835 ;
      RECT 88.285 8.58 88.63 8.81 ;
      RECT 88.11 8.61 88.63 8.78 ;
      RECT 83.76 4.865 84.08 5.125 ;
      RECT 85.05 4.04 85.19 4.9 ;
      RECT 83.85 4.76 85.19 4.9 ;
      RECT 83.85 4.32 83.99 5.125 ;
      RECT 83.775 4.32 84.065 4.55 ;
      RECT 84.975 4.04 85.265 4.27 ;
      RECT 84.495 4.32 84.785 4.55 ;
      RECT 84.69 3.245 84.83 4.505 ;
      RECT 84.72 3.185 85.04 3.445 ;
      RECT 81.32 3.745 81.64 4.005 ;
      RECT 84.015 3.76 84.305 3.99 ;
      RECT 81.41 3.665 84.23 3.805 ;
      RECT 83.28 3.185 83.6 3.445 ;
      RECT 83.775 3.2 84.065 3.43 ;
      RECT 83.28 3.245 84.065 3.385 ;
      RECT 83.28 4.305 83.6 4.565 ;
      RECT 83.28 4.085 83.51 4.565 ;
      RECT 82.775 4.04 83.065 4.27 ;
      RECT 82.775 4.085 83.51 4.225 ;
      RECT 83.04 10.06 83.33 10.29 ;
      RECT 83.1 9.32 83.27 10.29 ;
      RECT 83 9.345 83.38 9.715 ;
      RECT 83.04 9.32 83.33 9.715 ;
      RECT 81.8 4.865 82.12 5.125 ;
      RECT 81.335 4.88 81.625 5.11 ;
      RECT 81.335 4.925 82.12 5.065 ;
      RECT 80.095 3.76 80.385 3.99 ;
      RECT 80.095 3.805 81.03 3.945 ;
      RECT 80.89 3.245 81.03 3.945 ;
      RECT 81.56 3.185 81.88 3.445 ;
      RECT 81.335 3.2 81.88 3.43 ;
      RECT 80.89 3.245 81.88 3.385 ;
      RECT 79.24 4.865 79.56 5.125 ;
      RECT 79.24 4.925 80.31 5.065 ;
      RECT 80.17 4.365 80.31 5.065 ;
      RECT 81.335 4.32 81.625 4.55 ;
      RECT 80.17 4.365 81.625 4.505 ;
      RECT 79.6 3.185 79.92 3.445 ;
      RECT 79.375 3.2 79.92 3.43 ;
      RECT 78.62 3.745 78.94 4.005 ;
      RECT 79.615 3.76 79.905 3.99 ;
      RECT 78.375 3.76 78.94 3.99 ;
      RECT 78.375 3.805 79.905 3.945 ;
      RECT 77.895 4.32 78.185 4.55 ;
      RECT 78.09 3.245 78.23 4.505 ;
      RECT 78.88 3.185 79.2 3.445 ;
      RECT 77.895 3.2 78.185 3.43 ;
      RECT 77.895 3.245 79.2 3.385 ;
      RECT 77.49 4.76 78.59 4.9 ;
      RECT 78.375 4.6 78.665 4.83 ;
      RECT 77.415 4.6 77.705 4.83 ;
      RECT 77.4 3.185 77.72 3.445 ;
      RECT 75.44 3.185 75.76 3.445 ;
      RECT 75.44 3.245 77.72 3.385 ;
      RECT 76.56 4.305 76.88 4.565 ;
      RECT 76.56 4.305 77.39 4.445 ;
      RECT 77.175 4.04 77.39 4.445 ;
      RECT 77.175 4.04 77.465 4.27 ;
      RECT 74.96 3.745 75.28 4.005 ;
      RECT 76.37 3.76 76.66 3.99 ;
      RECT 74.96 3.76 75.505 3.99 ;
      RECT 74.96 3.845 75.91 3.985 ;
      RECT 75.77 3.665 75.91 3.985 ;
      RECT 76.27 3.76 76.66 3.945 ;
      RECT 75.77 3.665 76.41 3.805 ;
      RECT 74.48 4.555 74.8 4.97 ;
      RECT 74.56 3.2 74.715 4.97 ;
      RECT 74.495 3.2 74.785 3.43 ;
      RECT 72.875 10.055 73.17 10.285 ;
      RECT 72.935 8.575 73.105 10.285 ;
      RECT 72.885 8.945 73.235 9.295 ;
      RECT 72.875 8.575 73.165 8.805 ;
      RECT 71.885 10.055 72.18 10.285 ;
      RECT 71.945 8.575 72.115 10.285 ;
      RECT 71.945 8.81 72.735 8.97 ;
      RECT 72.58 8.205 72.735 8.97 ;
      RECT 72.57 8.63 72.735 8.97 ;
      RECT 71.945 8.575 72.175 8.97 ;
      RECT 71.885 8.575 72.175 8.805 ;
      RECT 72.505 8.205 72.795 8.435 ;
      RECT 72.505 8.235 72.965 8.405 ;
      RECT 72.5 4.03 72.79 4.26 ;
      RECT 72.47 3.725 72.66 4.255 ;
      RECT 72.47 4.06 72.96 4.23 ;
      RECT 72.115 3.725 72.66 3.895 ;
      RECT 71.945 2.18 72.115 3.89 ;
      RECT 71.885 3.66 72.175 3.89 ;
      RECT 71.885 2.18 72.18 2.41 ;
      RECT 71.58 4.03 71.75 4.335 ;
      RECT 71.515 4.03 71.805 4.26 ;
      RECT 71.515 4.06 71.975 4.23 ;
      RECT 71.58 2.95 71.745 4.335 ;
      RECT 70.095 2.915 70.385 3.145 ;
      RECT 70.095 2.95 71.745 3.12 ;
      RECT 70.155 2.175 70.325 3.145 ;
      RECT 70.095 2.175 70.385 2.405 ;
      RECT 70.095 10.06 70.385 10.29 ;
      RECT 70.155 9.32 70.325 10.29 ;
      RECT 70.155 9.41 71.745 9.58 ;
      RECT 71.575 8.205 71.745 9.58 ;
      RECT 70.095 9.32 70.385 9.55 ;
      RECT 71.515 8.205 71.805 8.435 ;
      RECT 71.515 8.235 71.975 8.405 ;
      RECT 68.145 4.445 68.485 4.795 ;
      RECT 68.235 3.32 68.405 4.795 ;
      RECT 70.525 3.26 70.875 3.61 ;
      RECT 68.235 3.32 70.875 3.49 ;
      RECT 70.355 3.315 70.875 3.49 ;
      RECT 70.55 8.945 70.875 9.27 ;
      RECT 65.11 8.905 65.46 9.255 ;
      RECT 70.525 8.95 70.875 9.18 ;
      RECT 64.91 8.95 65.46 9.18 ;
      RECT 70.355 8.975 70.875 9.15 ;
      RECT 64.74 8.975 65.46 9.15 ;
      RECT 64.74 8.975 70.875 9.145 ;
      RECT 69.75 3.66 70.07 3.98 ;
      RECT 69.725 3.655 70.015 3.885 ;
      RECT 69.72 3.685 70.07 3.86 ;
      RECT 69.55 3.685 70.07 3.855 ;
      RECT 69.75 8.545 70.07 8.835 ;
      RECT 69.725 8.58 70.07 8.81 ;
      RECT 69.55 8.61 70.07 8.78 ;
      RECT 65.2 4.865 65.52 5.125 ;
      RECT 66.49 4.04 66.63 4.9 ;
      RECT 65.29 4.76 66.63 4.9 ;
      RECT 65.29 4.32 65.43 5.125 ;
      RECT 65.215 4.32 65.505 4.55 ;
      RECT 66.415 4.04 66.705 4.27 ;
      RECT 65.935 4.32 66.225 4.55 ;
      RECT 66.13 3.245 66.27 4.505 ;
      RECT 66.16 3.185 66.48 3.445 ;
      RECT 62.76 3.745 63.08 4.005 ;
      RECT 65.455 3.76 65.745 3.99 ;
      RECT 62.85 3.665 65.67 3.805 ;
      RECT 64.72 3.185 65.04 3.445 ;
      RECT 65.215 3.2 65.505 3.43 ;
      RECT 64.72 3.245 65.505 3.385 ;
      RECT 64.72 4.305 65.04 4.565 ;
      RECT 64.72 4.085 64.95 4.565 ;
      RECT 64.215 4.04 64.505 4.27 ;
      RECT 64.215 4.085 64.95 4.225 ;
      RECT 64.48 10.06 64.77 10.29 ;
      RECT 64.54 9.32 64.71 10.29 ;
      RECT 64.44 9.345 64.82 9.715 ;
      RECT 64.48 9.32 64.77 9.715 ;
      RECT 63.24 4.865 63.56 5.125 ;
      RECT 62.775 4.88 63.065 5.11 ;
      RECT 62.775 4.925 63.56 5.065 ;
      RECT 61.535 3.76 61.825 3.99 ;
      RECT 61.535 3.805 62.47 3.945 ;
      RECT 62.33 3.245 62.47 3.945 ;
      RECT 63 3.185 63.32 3.445 ;
      RECT 62.775 3.2 63.32 3.43 ;
      RECT 62.33 3.245 63.32 3.385 ;
      RECT 60.68 4.865 61 5.125 ;
      RECT 60.68 4.925 61.75 5.065 ;
      RECT 61.61 4.365 61.75 5.065 ;
      RECT 62.775 4.32 63.065 4.55 ;
      RECT 61.61 4.365 63.065 4.505 ;
      RECT 61.04 3.185 61.36 3.445 ;
      RECT 60.815 3.2 61.36 3.43 ;
      RECT 60.06 3.745 60.38 4.005 ;
      RECT 61.055 3.76 61.345 3.99 ;
      RECT 59.815 3.76 60.38 3.99 ;
      RECT 59.815 3.805 61.345 3.945 ;
      RECT 59.335 4.32 59.625 4.55 ;
      RECT 59.53 3.245 59.67 4.505 ;
      RECT 60.32 3.185 60.64 3.445 ;
      RECT 59.335 3.2 59.625 3.43 ;
      RECT 59.335 3.245 60.64 3.385 ;
      RECT 58.93 4.76 60.03 4.9 ;
      RECT 59.815 4.6 60.105 4.83 ;
      RECT 58.855 4.6 59.145 4.83 ;
      RECT 58.84 3.185 59.16 3.445 ;
      RECT 56.88 3.185 57.2 3.445 ;
      RECT 56.88 3.245 59.16 3.385 ;
      RECT 58 4.305 58.32 4.565 ;
      RECT 58 4.305 58.83 4.445 ;
      RECT 58.615 4.04 58.83 4.445 ;
      RECT 58.615 4.04 58.905 4.27 ;
      RECT 56.4 3.745 56.72 4.005 ;
      RECT 57.81 3.76 58.1 3.99 ;
      RECT 56.4 3.76 56.945 3.99 ;
      RECT 56.4 3.845 57.35 3.985 ;
      RECT 57.21 3.665 57.35 3.985 ;
      RECT 57.71 3.76 58.1 3.945 ;
      RECT 57.21 3.665 57.85 3.805 ;
      RECT 55.92 4.555 56.24 4.97 ;
      RECT 56 3.2 56.155 4.97 ;
      RECT 55.935 3.2 56.225 3.43 ;
      RECT 54.315 10.055 54.61 10.285 ;
      RECT 54.375 8.575 54.545 10.285 ;
      RECT 54.365 8.95 54.72 9.305 ;
      RECT 54.315 8.575 54.605 8.805 ;
      RECT 53.325 10.055 53.62 10.285 ;
      RECT 53.385 8.575 53.555 10.285 ;
      RECT 53.385 8.81 54.175 8.97 ;
      RECT 54.02 8.205 54.175 8.97 ;
      RECT 54.01 8.63 54.175 8.97 ;
      RECT 53.385 8.575 53.615 8.97 ;
      RECT 53.325 8.575 53.615 8.805 ;
      RECT 53.945 8.205 54.235 8.435 ;
      RECT 53.945 8.235 54.405 8.405 ;
      RECT 53.94 4.03 54.23 4.26 ;
      RECT 53.91 3.725 54.1 4.255 ;
      RECT 53.91 4.06 54.4 4.23 ;
      RECT 53.555 3.725 54.1 3.895 ;
      RECT 53.385 2.18 53.555 3.89 ;
      RECT 53.325 3.66 53.615 3.89 ;
      RECT 53.325 2.18 53.62 2.41 ;
      RECT 53.02 4.03 53.19 4.335 ;
      RECT 52.955 4.03 53.245 4.26 ;
      RECT 52.955 4.06 53.415 4.23 ;
      RECT 53.02 2.95 53.185 4.335 ;
      RECT 51.535 2.915 51.825 3.145 ;
      RECT 51.535 2.95 53.185 3.12 ;
      RECT 51.595 2.175 51.765 3.145 ;
      RECT 51.535 2.175 51.825 2.405 ;
      RECT 51.535 10.06 51.825 10.29 ;
      RECT 51.595 9.32 51.765 10.29 ;
      RECT 51.595 9.41 53.185 9.58 ;
      RECT 53.015 8.205 53.185 9.58 ;
      RECT 51.535 9.32 51.825 9.55 ;
      RECT 52.955 8.205 53.245 8.435 ;
      RECT 52.955 8.235 53.415 8.405 ;
      RECT 49.585 4.445 49.925 4.795 ;
      RECT 49.675 3.32 49.845 4.795 ;
      RECT 51.965 3.26 52.315 3.61 ;
      RECT 49.675 3.32 52.315 3.49 ;
      RECT 51.795 3.315 52.315 3.49 ;
      RECT 51.99 8.945 52.315 9.27 ;
      RECT 46.555 8.9 46.905 9.25 ;
      RECT 51.965 8.95 52.315 9.18 ;
      RECT 46.35 8.95 46.905 9.18 ;
      RECT 51.795 8.975 52.315 9.15 ;
      RECT 46.18 8.975 46.905 9.15 ;
      RECT 46.18 8.975 52.315 9.145 ;
      RECT 51.19 3.66 51.51 3.98 ;
      RECT 51.165 3.655 51.455 3.885 ;
      RECT 51.16 3.685 51.51 3.86 ;
      RECT 50.99 3.685 51.51 3.855 ;
      RECT 51.19 8.545 51.51 8.835 ;
      RECT 51.165 8.58 51.51 8.81 ;
      RECT 50.99 8.61 51.51 8.78 ;
      RECT 46.64 4.865 46.96 5.125 ;
      RECT 47.93 4.04 48.07 4.9 ;
      RECT 46.73 4.76 48.07 4.9 ;
      RECT 46.73 4.32 46.87 5.125 ;
      RECT 46.655 4.32 46.945 4.55 ;
      RECT 47.855 4.04 48.145 4.27 ;
      RECT 47.375 4.32 47.665 4.55 ;
      RECT 47.57 3.245 47.71 4.505 ;
      RECT 47.6 3.185 47.92 3.445 ;
      RECT 44.2 3.745 44.52 4.005 ;
      RECT 46.895 3.76 47.185 3.99 ;
      RECT 44.29 3.665 47.11 3.805 ;
      RECT 46.16 3.185 46.48 3.445 ;
      RECT 46.655 3.2 46.945 3.43 ;
      RECT 46.16 3.245 46.945 3.385 ;
      RECT 46.16 4.305 46.48 4.565 ;
      RECT 46.16 4.085 46.39 4.565 ;
      RECT 45.655 4.04 45.945 4.27 ;
      RECT 45.655 4.085 46.39 4.225 ;
      RECT 45.92 10.06 46.21 10.29 ;
      RECT 45.98 9.32 46.15 10.29 ;
      RECT 45.88 9.345 46.26 9.715 ;
      RECT 45.92 9.32 46.21 9.715 ;
      RECT 44.68 4.865 45 5.125 ;
      RECT 44.215 4.88 44.505 5.11 ;
      RECT 44.215 4.925 45 5.065 ;
      RECT 42.975 3.76 43.265 3.99 ;
      RECT 42.975 3.805 43.91 3.945 ;
      RECT 43.77 3.245 43.91 3.945 ;
      RECT 44.44 3.185 44.76 3.445 ;
      RECT 44.215 3.2 44.76 3.43 ;
      RECT 43.77 3.245 44.76 3.385 ;
      RECT 42.12 4.865 42.44 5.125 ;
      RECT 42.12 4.925 43.19 5.065 ;
      RECT 43.05 4.365 43.19 5.065 ;
      RECT 44.215 4.32 44.505 4.55 ;
      RECT 43.05 4.365 44.505 4.505 ;
      RECT 42.48 3.185 42.8 3.445 ;
      RECT 42.255 3.2 42.8 3.43 ;
      RECT 41.5 3.745 41.82 4.005 ;
      RECT 42.495 3.76 42.785 3.99 ;
      RECT 41.255 3.76 41.82 3.99 ;
      RECT 41.255 3.805 42.785 3.945 ;
      RECT 40.775 4.32 41.065 4.55 ;
      RECT 40.97 3.245 41.11 4.505 ;
      RECT 41.76 3.185 42.08 3.445 ;
      RECT 40.775 3.2 41.065 3.43 ;
      RECT 40.775 3.245 42.08 3.385 ;
      RECT 40.37 4.76 41.47 4.9 ;
      RECT 41.255 4.6 41.545 4.83 ;
      RECT 40.295 4.6 40.585 4.83 ;
      RECT 40.28 3.185 40.6 3.445 ;
      RECT 38.32 3.185 38.64 3.445 ;
      RECT 38.32 3.245 40.6 3.385 ;
      RECT 39.44 4.305 39.76 4.565 ;
      RECT 39.44 4.305 40.27 4.445 ;
      RECT 40.055 4.04 40.27 4.445 ;
      RECT 40.055 4.04 40.345 4.27 ;
      RECT 37.84 3.745 38.16 4.005 ;
      RECT 39.25 3.76 39.54 3.99 ;
      RECT 37.84 3.76 38.385 3.99 ;
      RECT 37.84 3.845 38.79 3.985 ;
      RECT 38.65 3.665 38.79 3.985 ;
      RECT 39.15 3.76 39.54 3.945 ;
      RECT 38.65 3.665 39.29 3.805 ;
      RECT 37.36 4.555 37.68 4.97 ;
      RECT 37.44 3.2 37.595 4.97 ;
      RECT 37.375 3.2 37.665 3.43 ;
      RECT 35.755 10.055 36.05 10.285 ;
      RECT 35.815 8.575 35.985 10.285 ;
      RECT 35.81 8.945 36.16 9.295 ;
      RECT 35.755 8.575 36.045 8.805 ;
      RECT 34.765 10.055 35.06 10.285 ;
      RECT 34.825 8.575 34.995 10.285 ;
      RECT 34.825 8.81 35.615 8.97 ;
      RECT 35.46 8.205 35.615 8.97 ;
      RECT 35.45 8.63 35.615 8.97 ;
      RECT 34.825 8.575 35.055 8.97 ;
      RECT 34.765 8.575 35.055 8.805 ;
      RECT 35.385 8.205 35.675 8.435 ;
      RECT 35.385 8.235 35.845 8.405 ;
      RECT 35.38 4.03 35.67 4.26 ;
      RECT 35.35 3.725 35.54 4.255 ;
      RECT 35.35 4.06 35.84 4.23 ;
      RECT 34.995 3.725 35.54 3.895 ;
      RECT 34.825 2.18 34.995 3.89 ;
      RECT 34.765 3.66 35.055 3.89 ;
      RECT 34.765 2.18 35.06 2.41 ;
      RECT 34.46 4.03 34.63 4.335 ;
      RECT 34.395 4.03 34.685 4.26 ;
      RECT 34.395 4.06 34.855 4.23 ;
      RECT 34.46 2.95 34.625 4.335 ;
      RECT 32.975 2.915 33.265 3.145 ;
      RECT 32.975 2.95 34.625 3.12 ;
      RECT 33.035 2.175 33.205 3.145 ;
      RECT 32.975 2.175 33.265 2.405 ;
      RECT 32.975 10.06 33.265 10.29 ;
      RECT 33.035 9.32 33.205 10.29 ;
      RECT 33.035 9.41 34.625 9.58 ;
      RECT 34.455 8.205 34.625 9.58 ;
      RECT 32.975 9.32 33.265 9.55 ;
      RECT 34.395 8.205 34.685 8.435 ;
      RECT 34.395 8.235 34.855 8.405 ;
      RECT 31.025 4.445 31.365 4.795 ;
      RECT 31.115 3.32 31.285 4.795 ;
      RECT 33.405 3.26 33.755 3.61 ;
      RECT 31.115 3.32 33.755 3.49 ;
      RECT 33.235 3.315 33.755 3.49 ;
      RECT 33.43 8.945 33.755 9.27 ;
      RECT 27.995 8.895 28.345 9.245 ;
      RECT 33.405 8.95 33.755 9.18 ;
      RECT 27.79 8.95 28.345 9.18 ;
      RECT 33.235 8.975 33.755 9.15 ;
      RECT 27.62 8.975 28.345 9.15 ;
      RECT 27.62 8.975 33.755 9.145 ;
      RECT 32.63 3.66 32.95 3.98 ;
      RECT 32.605 3.655 32.895 3.885 ;
      RECT 32.6 3.685 32.95 3.86 ;
      RECT 32.43 3.685 32.95 3.855 ;
      RECT 32.63 8.545 32.95 8.835 ;
      RECT 32.605 8.58 32.95 8.81 ;
      RECT 32.43 8.61 32.95 8.78 ;
      RECT 28.08 4.865 28.4 5.125 ;
      RECT 29.37 4.04 29.51 4.9 ;
      RECT 28.17 4.76 29.51 4.9 ;
      RECT 28.17 4.32 28.31 5.125 ;
      RECT 28.095 4.32 28.385 4.55 ;
      RECT 29.295 4.04 29.585 4.27 ;
      RECT 28.815 4.32 29.105 4.55 ;
      RECT 29.01 3.245 29.15 4.505 ;
      RECT 29.04 3.185 29.36 3.445 ;
      RECT 25.64 3.745 25.96 4.005 ;
      RECT 28.335 3.76 28.625 3.99 ;
      RECT 25.73 3.665 28.55 3.805 ;
      RECT 27.6 3.185 27.92 3.445 ;
      RECT 28.095 3.2 28.385 3.43 ;
      RECT 27.6 3.245 28.385 3.385 ;
      RECT 27.6 4.305 27.92 4.565 ;
      RECT 27.6 4.085 27.83 4.565 ;
      RECT 27.095 4.04 27.385 4.27 ;
      RECT 27.095 4.085 27.83 4.225 ;
      RECT 27.36 10.06 27.65 10.29 ;
      RECT 27.42 9.32 27.59 10.29 ;
      RECT 27.32 9.345 27.7 9.715 ;
      RECT 27.36 9.32 27.65 9.715 ;
      RECT 26.12 4.865 26.44 5.125 ;
      RECT 25.655 4.88 25.945 5.11 ;
      RECT 25.655 4.925 26.44 5.065 ;
      RECT 24.415 3.76 24.705 3.99 ;
      RECT 24.415 3.805 25.35 3.945 ;
      RECT 25.21 3.245 25.35 3.945 ;
      RECT 25.88 3.185 26.2 3.445 ;
      RECT 25.655 3.2 26.2 3.43 ;
      RECT 25.21 3.245 26.2 3.385 ;
      RECT 23.56 4.865 23.88 5.125 ;
      RECT 23.56 4.925 24.63 5.065 ;
      RECT 24.49 4.365 24.63 5.065 ;
      RECT 25.655 4.32 25.945 4.55 ;
      RECT 24.49 4.365 25.945 4.505 ;
      RECT 23.92 3.185 24.24 3.445 ;
      RECT 23.695 3.2 24.24 3.43 ;
      RECT 22.94 3.745 23.26 4.005 ;
      RECT 23.935 3.76 24.225 3.99 ;
      RECT 22.695 3.76 23.26 3.99 ;
      RECT 22.695 3.805 24.225 3.945 ;
      RECT 22.215 4.32 22.505 4.55 ;
      RECT 22.41 3.245 22.55 4.505 ;
      RECT 23.2 3.185 23.52 3.445 ;
      RECT 22.215 3.2 22.505 3.43 ;
      RECT 22.215 3.245 23.52 3.385 ;
      RECT 21.81 4.76 22.91 4.9 ;
      RECT 22.695 4.6 22.985 4.83 ;
      RECT 21.735 4.6 22.025 4.83 ;
      RECT 21.72 3.185 22.04 3.445 ;
      RECT 19.76 3.185 20.08 3.445 ;
      RECT 19.76 3.245 22.04 3.385 ;
      RECT 20.88 4.305 21.2 4.565 ;
      RECT 20.88 4.305 21.71 4.445 ;
      RECT 21.495 4.04 21.71 4.445 ;
      RECT 21.495 4.04 21.785 4.27 ;
      RECT 19.28 3.745 19.6 4.005 ;
      RECT 20.69 3.76 20.98 3.99 ;
      RECT 19.28 3.76 19.825 3.99 ;
      RECT 19.28 3.845 20.23 3.985 ;
      RECT 20.09 3.665 20.23 3.985 ;
      RECT 20.59 3.76 20.98 3.945 ;
      RECT 20.09 3.665 20.73 3.805 ;
      RECT 18.8 4.555 19.12 4.97 ;
      RECT 18.88 3.2 19.035 4.97 ;
      RECT 18.815 3.2 19.105 3.43 ;
      RECT 16.545 10.06 16.835 10.29 ;
      RECT 16.605 9.315 16.775 10.29 ;
      RECT 16.515 9.315 16.865 9.605 ;
      RECT 16.14 8.575 16.49 8.865 ;
      RECT 16 8.61 16.49 8.78 ;
      RECT 109.97 7.245 110.32 7.535 ;
      RECT 101.32 4.865 101.64 5.125 ;
      RECT 100.72 3.185 101.4 3.445 ;
      RECT 100.84 4.865 101.16 5.125 ;
      RECT 99.36 4.865 99.68 5.125 ;
      RECT 98.88 3.185 99.2 3.445 ;
      RECT 98.16 4.305 98.48 4.565 ;
      RECT 97.44 4.305 97.76 4.565 ;
      RECT 94 4.305 94.32 4.565 ;
      RECT 91.41 7.245 91.76 7.535 ;
      RECT 82.76 4.865 83.08 5.125 ;
      RECT 82.16 3.185 82.84 3.445 ;
      RECT 82.28 4.865 82.6 5.125 ;
      RECT 80.8 4.865 81.12 5.125 ;
      RECT 80.32 3.185 80.64 3.445 ;
      RECT 79.6 4.305 79.92 4.565 ;
      RECT 78.88 4.305 79.2 4.565 ;
      RECT 75.44 4.305 75.76 4.565 ;
      RECT 72.85 7.245 73.2 7.535 ;
      RECT 64.2 4.865 64.52 5.125 ;
      RECT 63.6 3.185 64.28 3.445 ;
      RECT 63.72 4.865 64.04 5.125 ;
      RECT 62.24 4.865 62.56 5.125 ;
      RECT 61.76 3.185 62.08 3.445 ;
      RECT 61.04 4.305 61.36 4.565 ;
      RECT 60.32 4.305 60.64 4.565 ;
      RECT 56.88 4.305 57.2 4.565 ;
      RECT 54.29 7.245 54.64 7.535 ;
      RECT 45.64 4.865 45.96 5.125 ;
      RECT 45.04 3.185 45.72 3.445 ;
      RECT 45.16 4.865 45.48 5.125 ;
      RECT 43.68 4.865 44 5.125 ;
      RECT 43.2 3.185 43.52 3.445 ;
      RECT 42.48 4.305 42.8 4.565 ;
      RECT 41.76 4.305 42.08 4.565 ;
      RECT 38.32 4.305 38.64 4.565 ;
      RECT 35.73 7.245 36.08 7.535 ;
      RECT 27.08 4.865 27.4 5.125 ;
      RECT 26.48 3.185 27.16 3.445 ;
      RECT 26.6 4.865 26.92 5.125 ;
      RECT 25.12 4.865 25.44 5.125 ;
      RECT 24.64 3.185 24.96 3.445 ;
      RECT 23.92 4.305 24.24 4.565 ;
      RECT 23.2 4.305 23.52 4.565 ;
      RECT 19.76 4.305 20.08 4.565 ;
    LAYER mcon ;
      RECT 110.06 7.305 110.23 7.475 ;
      RECT 110.055 8.605 110.225 8.775 ;
      RECT 110.055 10.085 110.225 10.255 ;
      RECT 109.685 8.235 109.855 8.405 ;
      RECT 109.68 4.06 109.85 4.23 ;
      RECT 109.065 2.21 109.235 2.38 ;
      RECT 109.065 3.69 109.235 3.86 ;
      RECT 109.065 8.605 109.235 8.775 ;
      RECT 109.065 10.085 109.235 10.255 ;
      RECT 108.695 4.06 108.865 4.23 ;
      RECT 108.695 8.235 108.865 8.405 ;
      RECT 107.705 3.315 107.875 3.485 ;
      RECT 107.705 8.98 107.875 9.15 ;
      RECT 107.275 2.205 107.445 2.375 ;
      RECT 107.275 2.945 107.445 3.115 ;
      RECT 107.275 9.35 107.445 9.52 ;
      RECT 107.275 10.09 107.445 10.26 ;
      RECT 106.905 3.685 107.075 3.855 ;
      RECT 106.905 8.61 107.075 8.78 ;
      RECT 103.595 4.07 103.765 4.24 ;
      RECT 103.355 3.23 103.525 3.4 ;
      RECT 103.115 4.35 103.285 4.52 ;
      RECT 102.635 3.79 102.805 3.96 ;
      RECT 102.395 3.23 102.565 3.4 ;
      RECT 102.395 4.35 102.565 4.52 ;
      RECT 102.395 4.91 102.565 5.08 ;
      RECT 102.09 8.98 102.26 9.15 ;
      RECT 101.915 4.35 102.085 4.52 ;
      RECT 101.66 9.35 101.83 9.52 ;
      RECT 101.66 10.09 101.83 10.26 ;
      RECT 101.395 4.07 101.565 4.24 ;
      RECT 101.395 4.91 101.565 5.08 ;
      RECT 100.915 3.23 101.085 3.4 ;
      RECT 100.915 4.91 101.085 5.08 ;
      RECT 99.955 3.23 100.125 3.4 ;
      RECT 99.955 3.79 100.125 3.96 ;
      RECT 99.955 4.35 100.125 4.52 ;
      RECT 99.955 4.91 100.125 5.08 ;
      RECT 99.435 4.91 99.605 5.08 ;
      RECT 98.955 3.23 99.125 3.4 ;
      RECT 98.715 3.79 98.885 3.96 ;
      RECT 98.235 3.79 98.405 3.96 ;
      RECT 98.235 4.35 98.405 4.52 ;
      RECT 97.995 3.23 98.165 3.4 ;
      RECT 97.515 4.35 97.685 4.52 ;
      RECT 96.995 3.79 97.165 3.96 ;
      RECT 96.995 4.63 97.165 4.8 ;
      RECT 96.515 3.23 96.685 3.4 ;
      RECT 96.515 4.35 96.685 4.52 ;
      RECT 96.035 4.63 96.205 4.8 ;
      RECT 95.795 4.07 95.965 4.24 ;
      RECT 94.99 3.79 95.16 3.96 ;
      RECT 94.075 3.23 94.245 3.4 ;
      RECT 94.075 4.35 94.245 4.52 ;
      RECT 93.835 3.79 94.005 3.96 ;
      RECT 93.115 3.23 93.285 3.4 ;
      RECT 93.115 4.77 93.285 4.94 ;
      RECT 91.5 7.305 91.67 7.475 ;
      RECT 91.495 8.605 91.665 8.775 ;
      RECT 91.495 10.085 91.665 10.255 ;
      RECT 91.125 8.235 91.295 8.405 ;
      RECT 91.12 4.06 91.29 4.23 ;
      RECT 90.505 2.21 90.675 2.38 ;
      RECT 90.505 3.69 90.675 3.86 ;
      RECT 90.505 8.605 90.675 8.775 ;
      RECT 90.505 10.085 90.675 10.255 ;
      RECT 90.135 4.06 90.305 4.23 ;
      RECT 90.135 8.235 90.305 8.405 ;
      RECT 89.145 3.315 89.315 3.485 ;
      RECT 89.145 8.98 89.315 9.15 ;
      RECT 88.715 2.205 88.885 2.375 ;
      RECT 88.715 2.945 88.885 3.115 ;
      RECT 88.715 9.35 88.885 9.52 ;
      RECT 88.715 10.09 88.885 10.26 ;
      RECT 88.345 3.685 88.515 3.855 ;
      RECT 88.345 8.61 88.515 8.78 ;
      RECT 85.035 4.07 85.205 4.24 ;
      RECT 84.795 3.23 84.965 3.4 ;
      RECT 84.555 4.35 84.725 4.52 ;
      RECT 84.075 3.79 84.245 3.96 ;
      RECT 83.835 3.23 84.005 3.4 ;
      RECT 83.835 4.35 84.005 4.52 ;
      RECT 83.835 4.91 84.005 5.08 ;
      RECT 83.53 8.98 83.7 9.15 ;
      RECT 83.355 4.35 83.525 4.52 ;
      RECT 83.1 9.35 83.27 9.52 ;
      RECT 83.1 10.09 83.27 10.26 ;
      RECT 82.835 4.07 83.005 4.24 ;
      RECT 82.835 4.91 83.005 5.08 ;
      RECT 82.355 3.23 82.525 3.4 ;
      RECT 82.355 4.91 82.525 5.08 ;
      RECT 81.395 3.23 81.565 3.4 ;
      RECT 81.395 3.79 81.565 3.96 ;
      RECT 81.395 4.35 81.565 4.52 ;
      RECT 81.395 4.91 81.565 5.08 ;
      RECT 80.875 4.91 81.045 5.08 ;
      RECT 80.395 3.23 80.565 3.4 ;
      RECT 80.155 3.79 80.325 3.96 ;
      RECT 79.675 3.79 79.845 3.96 ;
      RECT 79.675 4.35 79.845 4.52 ;
      RECT 79.435 3.23 79.605 3.4 ;
      RECT 78.955 4.35 79.125 4.52 ;
      RECT 78.435 3.79 78.605 3.96 ;
      RECT 78.435 4.63 78.605 4.8 ;
      RECT 77.955 3.23 78.125 3.4 ;
      RECT 77.955 4.35 78.125 4.52 ;
      RECT 77.475 4.63 77.645 4.8 ;
      RECT 77.235 4.07 77.405 4.24 ;
      RECT 76.43 3.79 76.6 3.96 ;
      RECT 75.515 3.23 75.685 3.4 ;
      RECT 75.515 4.35 75.685 4.52 ;
      RECT 75.275 3.79 75.445 3.96 ;
      RECT 74.555 3.23 74.725 3.4 ;
      RECT 74.555 4.77 74.725 4.94 ;
      RECT 72.94 7.305 73.11 7.475 ;
      RECT 72.935 8.605 73.105 8.775 ;
      RECT 72.935 10.085 73.105 10.255 ;
      RECT 72.565 8.235 72.735 8.405 ;
      RECT 72.56 4.06 72.73 4.23 ;
      RECT 71.945 2.21 72.115 2.38 ;
      RECT 71.945 3.69 72.115 3.86 ;
      RECT 71.945 8.605 72.115 8.775 ;
      RECT 71.945 10.085 72.115 10.255 ;
      RECT 71.575 4.06 71.745 4.23 ;
      RECT 71.575 8.235 71.745 8.405 ;
      RECT 70.585 3.315 70.755 3.485 ;
      RECT 70.585 8.98 70.755 9.15 ;
      RECT 70.155 2.205 70.325 2.375 ;
      RECT 70.155 2.945 70.325 3.115 ;
      RECT 70.155 9.35 70.325 9.52 ;
      RECT 70.155 10.09 70.325 10.26 ;
      RECT 69.785 3.685 69.955 3.855 ;
      RECT 69.785 8.61 69.955 8.78 ;
      RECT 66.475 4.07 66.645 4.24 ;
      RECT 66.235 3.23 66.405 3.4 ;
      RECT 65.995 4.35 66.165 4.52 ;
      RECT 65.515 3.79 65.685 3.96 ;
      RECT 65.275 3.23 65.445 3.4 ;
      RECT 65.275 4.35 65.445 4.52 ;
      RECT 65.275 4.91 65.445 5.08 ;
      RECT 64.97 8.98 65.14 9.15 ;
      RECT 64.795 4.35 64.965 4.52 ;
      RECT 64.54 9.35 64.71 9.52 ;
      RECT 64.54 10.09 64.71 10.26 ;
      RECT 64.275 4.07 64.445 4.24 ;
      RECT 64.275 4.91 64.445 5.08 ;
      RECT 63.795 3.23 63.965 3.4 ;
      RECT 63.795 4.91 63.965 5.08 ;
      RECT 62.835 3.23 63.005 3.4 ;
      RECT 62.835 3.79 63.005 3.96 ;
      RECT 62.835 4.35 63.005 4.52 ;
      RECT 62.835 4.91 63.005 5.08 ;
      RECT 62.315 4.91 62.485 5.08 ;
      RECT 61.835 3.23 62.005 3.4 ;
      RECT 61.595 3.79 61.765 3.96 ;
      RECT 61.115 3.79 61.285 3.96 ;
      RECT 61.115 4.35 61.285 4.52 ;
      RECT 60.875 3.23 61.045 3.4 ;
      RECT 60.395 4.35 60.565 4.52 ;
      RECT 59.875 3.79 60.045 3.96 ;
      RECT 59.875 4.63 60.045 4.8 ;
      RECT 59.395 3.23 59.565 3.4 ;
      RECT 59.395 4.35 59.565 4.52 ;
      RECT 58.915 4.63 59.085 4.8 ;
      RECT 58.675 4.07 58.845 4.24 ;
      RECT 57.87 3.79 58.04 3.96 ;
      RECT 56.955 3.23 57.125 3.4 ;
      RECT 56.955 4.35 57.125 4.52 ;
      RECT 56.715 3.79 56.885 3.96 ;
      RECT 55.995 3.23 56.165 3.4 ;
      RECT 55.995 4.77 56.165 4.94 ;
      RECT 54.38 7.305 54.55 7.475 ;
      RECT 54.375 8.605 54.545 8.775 ;
      RECT 54.375 10.085 54.545 10.255 ;
      RECT 54.005 8.235 54.175 8.405 ;
      RECT 54 4.06 54.17 4.23 ;
      RECT 53.385 2.21 53.555 2.38 ;
      RECT 53.385 3.69 53.555 3.86 ;
      RECT 53.385 8.605 53.555 8.775 ;
      RECT 53.385 10.085 53.555 10.255 ;
      RECT 53.015 4.06 53.185 4.23 ;
      RECT 53.015 8.235 53.185 8.405 ;
      RECT 52.025 3.315 52.195 3.485 ;
      RECT 52.025 8.98 52.195 9.15 ;
      RECT 51.595 2.205 51.765 2.375 ;
      RECT 51.595 2.945 51.765 3.115 ;
      RECT 51.595 9.35 51.765 9.52 ;
      RECT 51.595 10.09 51.765 10.26 ;
      RECT 51.225 3.685 51.395 3.855 ;
      RECT 51.225 8.61 51.395 8.78 ;
      RECT 47.915 4.07 48.085 4.24 ;
      RECT 47.675 3.23 47.845 3.4 ;
      RECT 47.435 4.35 47.605 4.52 ;
      RECT 46.955 3.79 47.125 3.96 ;
      RECT 46.715 3.23 46.885 3.4 ;
      RECT 46.715 4.35 46.885 4.52 ;
      RECT 46.715 4.91 46.885 5.08 ;
      RECT 46.41 8.98 46.58 9.15 ;
      RECT 46.235 4.35 46.405 4.52 ;
      RECT 45.98 9.35 46.15 9.52 ;
      RECT 45.98 10.09 46.15 10.26 ;
      RECT 45.715 4.07 45.885 4.24 ;
      RECT 45.715 4.91 45.885 5.08 ;
      RECT 45.235 3.23 45.405 3.4 ;
      RECT 45.235 4.91 45.405 5.08 ;
      RECT 44.275 3.23 44.445 3.4 ;
      RECT 44.275 3.79 44.445 3.96 ;
      RECT 44.275 4.35 44.445 4.52 ;
      RECT 44.275 4.91 44.445 5.08 ;
      RECT 43.755 4.91 43.925 5.08 ;
      RECT 43.275 3.23 43.445 3.4 ;
      RECT 43.035 3.79 43.205 3.96 ;
      RECT 42.555 3.79 42.725 3.96 ;
      RECT 42.555 4.35 42.725 4.52 ;
      RECT 42.315 3.23 42.485 3.4 ;
      RECT 41.835 4.35 42.005 4.52 ;
      RECT 41.315 3.79 41.485 3.96 ;
      RECT 41.315 4.63 41.485 4.8 ;
      RECT 40.835 3.23 41.005 3.4 ;
      RECT 40.835 4.35 41.005 4.52 ;
      RECT 40.355 4.63 40.525 4.8 ;
      RECT 40.115 4.07 40.285 4.24 ;
      RECT 39.31 3.79 39.48 3.96 ;
      RECT 38.395 3.23 38.565 3.4 ;
      RECT 38.395 4.35 38.565 4.52 ;
      RECT 38.155 3.79 38.325 3.96 ;
      RECT 37.435 3.23 37.605 3.4 ;
      RECT 37.435 4.77 37.605 4.94 ;
      RECT 35.82 7.305 35.99 7.475 ;
      RECT 35.815 8.605 35.985 8.775 ;
      RECT 35.815 10.085 35.985 10.255 ;
      RECT 35.445 8.235 35.615 8.405 ;
      RECT 35.44 4.06 35.61 4.23 ;
      RECT 34.825 2.21 34.995 2.38 ;
      RECT 34.825 3.69 34.995 3.86 ;
      RECT 34.825 8.605 34.995 8.775 ;
      RECT 34.825 10.085 34.995 10.255 ;
      RECT 34.455 4.06 34.625 4.23 ;
      RECT 34.455 8.235 34.625 8.405 ;
      RECT 33.465 3.315 33.635 3.485 ;
      RECT 33.465 8.98 33.635 9.15 ;
      RECT 33.035 2.205 33.205 2.375 ;
      RECT 33.035 2.945 33.205 3.115 ;
      RECT 33.035 9.35 33.205 9.52 ;
      RECT 33.035 10.09 33.205 10.26 ;
      RECT 32.665 3.685 32.835 3.855 ;
      RECT 32.665 8.61 32.835 8.78 ;
      RECT 29.355 4.07 29.525 4.24 ;
      RECT 29.115 3.23 29.285 3.4 ;
      RECT 28.875 4.35 29.045 4.52 ;
      RECT 28.395 3.79 28.565 3.96 ;
      RECT 28.155 3.23 28.325 3.4 ;
      RECT 28.155 4.35 28.325 4.52 ;
      RECT 28.155 4.91 28.325 5.08 ;
      RECT 27.85 8.98 28.02 9.15 ;
      RECT 27.675 4.35 27.845 4.52 ;
      RECT 27.42 9.35 27.59 9.52 ;
      RECT 27.42 10.09 27.59 10.26 ;
      RECT 27.155 4.07 27.325 4.24 ;
      RECT 27.155 4.91 27.325 5.08 ;
      RECT 26.675 3.23 26.845 3.4 ;
      RECT 26.675 4.91 26.845 5.08 ;
      RECT 25.715 3.23 25.885 3.4 ;
      RECT 25.715 3.79 25.885 3.96 ;
      RECT 25.715 4.35 25.885 4.52 ;
      RECT 25.715 4.91 25.885 5.08 ;
      RECT 25.195 4.91 25.365 5.08 ;
      RECT 24.715 3.23 24.885 3.4 ;
      RECT 24.475 3.79 24.645 3.96 ;
      RECT 23.995 3.79 24.165 3.96 ;
      RECT 23.995 4.35 24.165 4.52 ;
      RECT 23.755 3.23 23.925 3.4 ;
      RECT 23.275 4.35 23.445 4.52 ;
      RECT 22.755 3.79 22.925 3.96 ;
      RECT 22.755 4.63 22.925 4.8 ;
      RECT 22.275 3.23 22.445 3.4 ;
      RECT 22.275 4.35 22.445 4.52 ;
      RECT 21.795 4.63 21.965 4.8 ;
      RECT 21.555 4.07 21.725 4.24 ;
      RECT 20.75 3.79 20.92 3.96 ;
      RECT 19.835 3.23 20.005 3.4 ;
      RECT 19.835 4.35 20.005 4.52 ;
      RECT 19.595 3.79 19.765 3.96 ;
      RECT 18.875 3.23 19.045 3.4 ;
      RECT 18.875 4.77 19.045 4.94 ;
      RECT 16.605 9.35 16.775 9.52 ;
      RECT 16.605 10.09 16.775 10.26 ;
      RECT 16.235 8.61 16.405 8.78 ;
    LAYER li1 ;
      RECT 110.055 7.305 110.225 8.775 ;
      RECT 110.055 7.305 110.23 8.565 ;
      RECT 109.685 9.255 110.155 9.425 ;
      RECT 109.685 8.235 109.855 9.425 ;
      RECT 109.68 3.04 109.85 4.23 ;
      RECT 109.68 3.04 110.15 3.21 ;
      RECT 109.065 3.9 109.24 5.16 ;
      RECT 109.065 3.69 109.235 5.16 ;
      RECT 109.065 7.305 109.235 8.775 ;
      RECT 109.065 7.305 109.24 8.565 ;
      RECT 108.695 3.04 108.865 4.23 ;
      RECT 108.695 3.04 109.165 3.21 ;
      RECT 108.695 9.255 109.165 9.425 ;
      RECT 108.695 8.235 108.865 9.425 ;
      RECT 107.705 4.015 107.88 5.155 ;
      RECT 107.705 1.865 107.875 5.155 ;
      RECT 107.705 1.865 107.88 2.415 ;
      RECT 107.705 10.05 107.88 10.6 ;
      RECT 107.705 7.31 107.875 10.6 ;
      RECT 107.705 7.31 107.88 8.45 ;
      RECT 107.275 3.895 107.45 5.155 ;
      RECT 107.275 2.945 107.445 5.155 ;
      RECT 107.275 7.31 107.445 9.52 ;
      RECT 107.275 7.31 107.45 8.57 ;
      RECT 106.845 3.925 107.015 5.155 ;
      RECT 106.905 2.145 107.075 4.095 ;
      RECT 106.845 1.865 107.015 2.315 ;
      RECT 106.845 10.15 107.015 10.6 ;
      RECT 106.905 8.37 107.075 10.32 ;
      RECT 106.845 7.31 107.015 8.54 ;
      RECT 106.32 3.895 106.495 5.155 ;
      RECT 106.32 1.865 106.49 5.155 ;
      RECT 106.32 3.365 106.73 3.695 ;
      RECT 106.32 2.525 106.73 2.855 ;
      RECT 106.32 1.865 106.495 2.355 ;
      RECT 106.32 10.11 106.495 10.6 ;
      RECT 106.32 7.31 106.49 10.6 ;
      RECT 106.32 9.61 106.73 9.94 ;
      RECT 106.32 8.77 106.73 9.1 ;
      RECT 106.32 7.31 106.495 8.57 ;
      RECT 103.115 4.52 104.085 4.69 ;
      RECT 103.115 4.35 103.285 4.69 ;
      RECT 102.635 3.79 102.805 4.12 ;
      RECT 102.635 3.87 103.365 4.04 ;
      RECT 102.275 4.91 102.565 5.08 ;
      RECT 102.275 3.87 102.445 5.08 ;
      RECT 102.275 4.35 102.565 4.52 ;
      RECT 102.075 3.87 102.445 4.04 ;
      RECT 102.09 10.05 102.265 10.6 ;
      RECT 102.09 7.31 102.26 10.6 ;
      RECT 102.09 7.31 102.265 8.45 ;
      RECT 101.66 7.31 101.83 9.52 ;
      RECT 101.66 7.31 101.835 8.57 ;
      RECT 101.395 3.97 101.565 4.24 ;
      RECT 101.155 3.97 101.565 4.14 ;
      RECT 101.075 3.87 101.405 4.04 ;
      RECT 100.915 4.91 101.565 5.08 ;
      RECT 101.395 4.44 101.565 5.08 ;
      RECT 101.275 4.52 101.565 5.08 ;
      RECT 100.705 10.11 100.88 10.6 ;
      RECT 100.705 7.31 100.875 10.6 ;
      RECT 100.705 9.61 101.115 9.94 ;
      RECT 100.705 8.77 101.115 9.1 ;
      RECT 100.705 7.31 100.88 8.57 ;
      RECT 99.955 4.21 100.125 4.52 ;
      RECT 99.955 4.21 100.845 4.38 ;
      RECT 100.675 3.79 100.845 4.38 ;
      RECT 99.955 3.87 100.445 4.04 ;
      RECT 99.955 3.79 100.125 4.04 ;
      RECT 97.915 4.52 98.405 4.69 ;
      RECT 99.075 3.87 99.245 4.52 ;
      RECT 98.235 4.35 99.245 4.52 ;
      RECT 99.195 3.79 99.365 4.12 ;
      RECT 97.995 3.13 98.165 3.4 ;
      RECT 97.435 3.13 98.165 3.3 ;
      RECT 97.515 3.87 97.685 4.52 ;
      RECT 97.515 3.87 98.005 4.04 ;
      RECT 96.675 3.87 97.165 4.04 ;
      RECT 96.995 3.79 97.165 4.04 ;
      RECT 96.515 3.13 96.685 3.4 ;
      RECT 95.955 3.13 96.685 3.3 ;
      RECT 96.035 4.52 96.205 4.8 ;
      RECT 94.995 4.52 96.285 4.69 ;
      RECT 94.99 3.87 95.565 4.04 ;
      RECT 94.99 3.79 95.16 4.04 ;
      RECT 94.075 3.13 94.245 3.4 ;
      RECT 94.075 3.13 94.805 3.3 ;
      RECT 94.075 4.35 94.245 4.77 ;
      RECT 93.455 4.435 94.245 4.605 ;
      RECT 93.455 4.21 93.625 4.605 ;
      RECT 93.355 3.79 93.525 4.38 ;
      RECT 93.115 3.87 93.525 4.14 ;
      RECT 91.495 7.305 91.665 8.775 ;
      RECT 91.495 7.305 91.67 8.565 ;
      RECT 91.125 9.255 91.595 9.425 ;
      RECT 91.125 8.235 91.295 9.425 ;
      RECT 91.12 3.04 91.29 4.23 ;
      RECT 91.12 3.04 91.59 3.21 ;
      RECT 90.505 3.9 90.68 5.16 ;
      RECT 90.505 3.69 90.675 5.16 ;
      RECT 90.505 7.305 90.675 8.775 ;
      RECT 90.505 7.305 90.68 8.565 ;
      RECT 90.135 3.04 90.305 4.23 ;
      RECT 90.135 3.04 90.605 3.21 ;
      RECT 90.135 9.255 90.605 9.425 ;
      RECT 90.135 8.235 90.305 9.425 ;
      RECT 89.145 4.015 89.32 5.155 ;
      RECT 89.145 1.865 89.315 5.155 ;
      RECT 89.145 1.865 89.32 2.415 ;
      RECT 89.145 10.05 89.32 10.6 ;
      RECT 89.145 7.31 89.315 10.6 ;
      RECT 89.145 7.31 89.32 8.45 ;
      RECT 88.715 3.895 88.89 5.155 ;
      RECT 88.715 2.945 88.885 5.155 ;
      RECT 88.715 7.31 88.885 9.52 ;
      RECT 88.715 7.31 88.89 8.57 ;
      RECT 88.285 3.925 88.455 5.155 ;
      RECT 88.345 2.145 88.515 4.095 ;
      RECT 88.285 1.865 88.455 2.315 ;
      RECT 88.285 10.15 88.455 10.6 ;
      RECT 88.345 8.37 88.515 10.32 ;
      RECT 88.285 7.31 88.455 8.54 ;
      RECT 87.76 3.895 87.935 5.155 ;
      RECT 87.76 1.865 87.93 5.155 ;
      RECT 87.76 3.365 88.17 3.695 ;
      RECT 87.76 2.525 88.17 2.855 ;
      RECT 87.76 1.865 87.935 2.355 ;
      RECT 87.76 10.11 87.935 10.6 ;
      RECT 87.76 7.31 87.93 10.6 ;
      RECT 87.76 9.61 88.17 9.94 ;
      RECT 87.76 8.77 88.17 9.1 ;
      RECT 87.76 7.31 87.935 8.57 ;
      RECT 84.555 4.52 85.525 4.69 ;
      RECT 84.555 4.35 84.725 4.69 ;
      RECT 84.075 3.79 84.245 4.12 ;
      RECT 84.075 3.87 84.805 4.04 ;
      RECT 83.715 4.91 84.005 5.08 ;
      RECT 83.715 3.87 83.885 5.08 ;
      RECT 83.715 4.35 84.005 4.52 ;
      RECT 83.515 3.87 83.885 4.04 ;
      RECT 83.53 10.05 83.705 10.6 ;
      RECT 83.53 7.31 83.7 10.6 ;
      RECT 83.53 7.31 83.705 8.45 ;
      RECT 83.1 7.31 83.27 9.52 ;
      RECT 83.1 7.31 83.275 8.57 ;
      RECT 82.835 3.97 83.005 4.24 ;
      RECT 82.595 3.97 83.005 4.14 ;
      RECT 82.515 3.87 82.845 4.04 ;
      RECT 82.355 4.91 83.005 5.08 ;
      RECT 82.835 4.44 83.005 5.08 ;
      RECT 82.715 4.52 83.005 5.08 ;
      RECT 82.145 10.11 82.32 10.6 ;
      RECT 82.145 7.31 82.315 10.6 ;
      RECT 82.145 9.61 82.555 9.94 ;
      RECT 82.145 8.77 82.555 9.1 ;
      RECT 82.145 7.31 82.32 8.57 ;
      RECT 81.395 4.21 81.565 4.52 ;
      RECT 81.395 4.21 82.285 4.38 ;
      RECT 82.115 3.79 82.285 4.38 ;
      RECT 81.395 3.87 81.885 4.04 ;
      RECT 81.395 3.79 81.565 4.04 ;
      RECT 79.355 4.52 79.845 4.69 ;
      RECT 80.515 3.87 80.685 4.52 ;
      RECT 79.675 4.35 80.685 4.52 ;
      RECT 80.635 3.79 80.805 4.12 ;
      RECT 79.435 3.13 79.605 3.4 ;
      RECT 78.875 3.13 79.605 3.3 ;
      RECT 78.955 3.87 79.125 4.52 ;
      RECT 78.955 3.87 79.445 4.04 ;
      RECT 78.115 3.87 78.605 4.04 ;
      RECT 78.435 3.79 78.605 4.04 ;
      RECT 77.955 3.13 78.125 3.4 ;
      RECT 77.395 3.13 78.125 3.3 ;
      RECT 77.475 4.52 77.645 4.8 ;
      RECT 76.435 4.52 77.725 4.69 ;
      RECT 76.43 3.87 77.005 4.04 ;
      RECT 76.43 3.79 76.6 4.04 ;
      RECT 75.515 3.13 75.685 3.4 ;
      RECT 75.515 3.13 76.245 3.3 ;
      RECT 75.515 4.35 75.685 4.77 ;
      RECT 74.895 4.435 75.685 4.605 ;
      RECT 74.895 4.21 75.065 4.605 ;
      RECT 74.795 3.79 74.965 4.38 ;
      RECT 74.555 3.87 74.965 4.14 ;
      RECT 72.935 7.305 73.105 8.775 ;
      RECT 72.935 7.305 73.11 8.565 ;
      RECT 72.565 9.255 73.035 9.425 ;
      RECT 72.565 8.235 72.735 9.425 ;
      RECT 72.56 3.04 72.73 4.23 ;
      RECT 72.56 3.04 73.03 3.21 ;
      RECT 71.945 3.9 72.12 5.16 ;
      RECT 71.945 3.69 72.115 5.16 ;
      RECT 71.945 7.305 72.115 8.775 ;
      RECT 71.945 7.305 72.12 8.565 ;
      RECT 71.575 3.04 71.745 4.23 ;
      RECT 71.575 3.04 72.045 3.21 ;
      RECT 71.575 9.255 72.045 9.425 ;
      RECT 71.575 8.235 71.745 9.425 ;
      RECT 70.585 4.015 70.76 5.155 ;
      RECT 70.585 1.865 70.755 5.155 ;
      RECT 70.585 1.865 70.76 2.415 ;
      RECT 70.585 10.05 70.76 10.6 ;
      RECT 70.585 7.31 70.755 10.6 ;
      RECT 70.585 7.31 70.76 8.45 ;
      RECT 70.155 3.895 70.33 5.155 ;
      RECT 70.155 2.945 70.325 5.155 ;
      RECT 70.155 7.31 70.325 9.52 ;
      RECT 70.155 7.31 70.33 8.57 ;
      RECT 69.725 3.925 69.895 5.155 ;
      RECT 69.785 2.145 69.955 4.095 ;
      RECT 69.725 1.865 69.895 2.315 ;
      RECT 69.725 10.15 69.895 10.6 ;
      RECT 69.785 8.37 69.955 10.32 ;
      RECT 69.725 7.31 69.895 8.54 ;
      RECT 69.2 3.895 69.375 5.155 ;
      RECT 69.2 1.865 69.37 5.155 ;
      RECT 69.2 3.365 69.61 3.695 ;
      RECT 69.2 2.525 69.61 2.855 ;
      RECT 69.2 1.865 69.375 2.355 ;
      RECT 69.2 10.11 69.375 10.6 ;
      RECT 69.2 7.31 69.37 10.6 ;
      RECT 69.2 9.61 69.61 9.94 ;
      RECT 69.2 8.77 69.61 9.1 ;
      RECT 69.2 7.31 69.375 8.57 ;
      RECT 65.995 4.52 66.965 4.69 ;
      RECT 65.995 4.35 66.165 4.69 ;
      RECT 65.515 3.79 65.685 4.12 ;
      RECT 65.515 3.87 66.245 4.04 ;
      RECT 65.155 4.91 65.445 5.08 ;
      RECT 65.155 3.87 65.325 5.08 ;
      RECT 65.155 4.35 65.445 4.52 ;
      RECT 64.955 3.87 65.325 4.04 ;
      RECT 64.97 10.05 65.145 10.6 ;
      RECT 64.97 7.31 65.14 10.6 ;
      RECT 64.97 7.31 65.145 8.45 ;
      RECT 64.54 7.31 64.71 9.52 ;
      RECT 64.54 7.31 64.715 8.57 ;
      RECT 64.275 3.97 64.445 4.24 ;
      RECT 64.035 3.97 64.445 4.14 ;
      RECT 63.955 3.87 64.285 4.04 ;
      RECT 63.795 4.91 64.445 5.08 ;
      RECT 64.275 4.44 64.445 5.08 ;
      RECT 64.155 4.52 64.445 5.08 ;
      RECT 63.585 10.11 63.76 10.6 ;
      RECT 63.585 7.31 63.755 10.6 ;
      RECT 63.585 9.61 63.995 9.94 ;
      RECT 63.585 8.77 63.995 9.1 ;
      RECT 63.585 7.31 63.76 8.57 ;
      RECT 62.835 4.21 63.005 4.52 ;
      RECT 62.835 4.21 63.725 4.38 ;
      RECT 63.555 3.79 63.725 4.38 ;
      RECT 62.835 3.87 63.325 4.04 ;
      RECT 62.835 3.79 63.005 4.04 ;
      RECT 60.795 4.52 61.285 4.69 ;
      RECT 61.955 3.87 62.125 4.52 ;
      RECT 61.115 4.35 62.125 4.52 ;
      RECT 62.075 3.79 62.245 4.12 ;
      RECT 60.875 3.13 61.045 3.4 ;
      RECT 60.315 3.13 61.045 3.3 ;
      RECT 60.395 3.87 60.565 4.52 ;
      RECT 60.395 3.87 60.885 4.04 ;
      RECT 59.555 3.87 60.045 4.04 ;
      RECT 59.875 3.79 60.045 4.04 ;
      RECT 59.395 3.13 59.565 3.4 ;
      RECT 58.835 3.13 59.565 3.3 ;
      RECT 58.915 4.52 59.085 4.8 ;
      RECT 57.875 4.52 59.165 4.69 ;
      RECT 57.87 3.87 58.445 4.04 ;
      RECT 57.87 3.79 58.04 4.04 ;
      RECT 56.955 3.13 57.125 3.4 ;
      RECT 56.955 3.13 57.685 3.3 ;
      RECT 56.955 4.35 57.125 4.77 ;
      RECT 56.335 4.435 57.125 4.605 ;
      RECT 56.335 4.21 56.505 4.605 ;
      RECT 56.235 3.79 56.405 4.38 ;
      RECT 55.995 3.87 56.405 4.14 ;
      RECT 54.375 7.305 54.545 8.775 ;
      RECT 54.375 7.305 54.55 8.565 ;
      RECT 54.005 9.255 54.475 9.425 ;
      RECT 54.005 8.235 54.175 9.425 ;
      RECT 54 3.04 54.17 4.23 ;
      RECT 54 3.04 54.47 3.21 ;
      RECT 53.385 3.9 53.56 5.16 ;
      RECT 53.385 3.69 53.555 5.16 ;
      RECT 53.385 7.305 53.555 8.775 ;
      RECT 53.385 7.305 53.56 8.565 ;
      RECT 53.015 3.04 53.185 4.23 ;
      RECT 53.015 3.04 53.485 3.21 ;
      RECT 53.015 9.255 53.485 9.425 ;
      RECT 53.015 8.235 53.185 9.425 ;
      RECT 52.025 4.015 52.2 5.155 ;
      RECT 52.025 1.865 52.195 5.155 ;
      RECT 52.025 1.865 52.2 2.415 ;
      RECT 52.025 10.05 52.2 10.6 ;
      RECT 52.025 7.31 52.195 10.6 ;
      RECT 52.025 7.31 52.2 8.45 ;
      RECT 51.595 3.895 51.77 5.155 ;
      RECT 51.595 2.945 51.765 5.155 ;
      RECT 51.595 7.31 51.765 9.52 ;
      RECT 51.595 7.31 51.77 8.57 ;
      RECT 51.165 3.925 51.335 5.155 ;
      RECT 51.225 2.145 51.395 4.095 ;
      RECT 51.165 1.865 51.335 2.315 ;
      RECT 51.165 10.15 51.335 10.6 ;
      RECT 51.225 8.37 51.395 10.32 ;
      RECT 51.165 7.31 51.335 8.54 ;
      RECT 50.64 3.895 50.815 5.155 ;
      RECT 50.64 1.865 50.81 5.155 ;
      RECT 50.64 3.365 51.05 3.695 ;
      RECT 50.64 2.525 51.05 2.855 ;
      RECT 50.64 1.865 50.815 2.355 ;
      RECT 50.64 10.11 50.815 10.6 ;
      RECT 50.64 7.31 50.81 10.6 ;
      RECT 50.64 9.61 51.05 9.94 ;
      RECT 50.64 8.77 51.05 9.1 ;
      RECT 50.64 7.31 50.815 8.57 ;
      RECT 47.435 4.52 48.405 4.69 ;
      RECT 47.435 4.35 47.605 4.69 ;
      RECT 46.955 3.79 47.125 4.12 ;
      RECT 46.955 3.87 47.685 4.04 ;
      RECT 46.595 4.91 46.885 5.08 ;
      RECT 46.595 3.87 46.765 5.08 ;
      RECT 46.595 4.35 46.885 4.52 ;
      RECT 46.395 3.87 46.765 4.04 ;
      RECT 46.41 10.05 46.585 10.6 ;
      RECT 46.41 7.31 46.58 10.6 ;
      RECT 46.41 7.31 46.585 8.45 ;
      RECT 45.98 7.31 46.15 9.52 ;
      RECT 45.98 7.31 46.155 8.57 ;
      RECT 45.715 3.97 45.885 4.24 ;
      RECT 45.475 3.97 45.885 4.14 ;
      RECT 45.395 3.87 45.725 4.04 ;
      RECT 45.235 4.91 45.885 5.08 ;
      RECT 45.715 4.44 45.885 5.08 ;
      RECT 45.595 4.52 45.885 5.08 ;
      RECT 45.025 10.11 45.2 10.6 ;
      RECT 45.025 7.31 45.195 10.6 ;
      RECT 45.025 9.61 45.435 9.94 ;
      RECT 45.025 8.77 45.435 9.1 ;
      RECT 45.025 7.31 45.2 8.57 ;
      RECT 44.275 4.21 44.445 4.52 ;
      RECT 44.275 4.21 45.165 4.38 ;
      RECT 44.995 3.79 45.165 4.38 ;
      RECT 44.275 3.87 44.765 4.04 ;
      RECT 44.275 3.79 44.445 4.04 ;
      RECT 42.235 4.52 42.725 4.69 ;
      RECT 43.395 3.87 43.565 4.52 ;
      RECT 42.555 4.35 43.565 4.52 ;
      RECT 43.515 3.79 43.685 4.12 ;
      RECT 42.315 3.13 42.485 3.4 ;
      RECT 41.755 3.13 42.485 3.3 ;
      RECT 41.835 3.87 42.005 4.52 ;
      RECT 41.835 3.87 42.325 4.04 ;
      RECT 40.995 3.87 41.485 4.04 ;
      RECT 41.315 3.79 41.485 4.04 ;
      RECT 40.835 3.13 41.005 3.4 ;
      RECT 40.275 3.13 41.005 3.3 ;
      RECT 40.355 4.52 40.525 4.8 ;
      RECT 39.315 4.52 40.605 4.69 ;
      RECT 39.31 3.87 39.885 4.04 ;
      RECT 39.31 3.79 39.48 4.04 ;
      RECT 38.395 3.13 38.565 3.4 ;
      RECT 38.395 3.13 39.125 3.3 ;
      RECT 38.395 4.35 38.565 4.77 ;
      RECT 37.775 4.435 38.565 4.605 ;
      RECT 37.775 4.21 37.945 4.605 ;
      RECT 37.675 3.79 37.845 4.38 ;
      RECT 37.435 3.87 37.845 4.14 ;
      RECT 35.815 7.305 35.985 8.775 ;
      RECT 35.815 7.305 35.99 8.565 ;
      RECT 35.445 9.255 35.915 9.425 ;
      RECT 35.445 8.235 35.615 9.425 ;
      RECT 35.44 3.04 35.61 4.23 ;
      RECT 35.44 3.04 35.91 3.21 ;
      RECT 34.825 3.9 35 5.16 ;
      RECT 34.825 3.69 34.995 5.16 ;
      RECT 34.825 7.305 34.995 8.775 ;
      RECT 34.825 7.305 35 8.565 ;
      RECT 34.455 3.04 34.625 4.23 ;
      RECT 34.455 3.04 34.925 3.21 ;
      RECT 34.455 9.255 34.925 9.425 ;
      RECT 34.455 8.235 34.625 9.425 ;
      RECT 33.465 4.015 33.64 5.155 ;
      RECT 33.465 1.865 33.635 5.155 ;
      RECT 33.465 1.865 33.64 2.415 ;
      RECT 33.465 10.05 33.64 10.6 ;
      RECT 33.465 7.31 33.635 10.6 ;
      RECT 33.465 7.31 33.64 8.45 ;
      RECT 33.035 3.895 33.21 5.155 ;
      RECT 33.035 2.945 33.205 5.155 ;
      RECT 33.035 7.31 33.205 9.52 ;
      RECT 33.035 7.31 33.21 8.57 ;
      RECT 32.605 3.925 32.775 5.155 ;
      RECT 32.665 2.145 32.835 4.095 ;
      RECT 32.605 1.865 32.775 2.315 ;
      RECT 32.605 10.15 32.775 10.6 ;
      RECT 32.665 8.37 32.835 10.32 ;
      RECT 32.605 7.31 32.775 8.54 ;
      RECT 32.08 3.895 32.255 5.155 ;
      RECT 32.08 1.865 32.25 5.155 ;
      RECT 32.08 3.365 32.49 3.695 ;
      RECT 32.08 2.525 32.49 2.855 ;
      RECT 32.08 1.865 32.255 2.355 ;
      RECT 32.08 10.11 32.255 10.6 ;
      RECT 32.08 7.31 32.25 10.6 ;
      RECT 32.08 9.61 32.49 9.94 ;
      RECT 32.08 8.77 32.49 9.1 ;
      RECT 32.08 7.31 32.255 8.57 ;
      RECT 28.875 4.52 29.845 4.69 ;
      RECT 28.875 4.35 29.045 4.69 ;
      RECT 28.395 3.79 28.565 4.12 ;
      RECT 28.395 3.87 29.125 4.04 ;
      RECT 28.035 4.91 28.325 5.08 ;
      RECT 28.035 3.87 28.205 5.08 ;
      RECT 28.035 4.35 28.325 4.52 ;
      RECT 27.835 3.87 28.205 4.04 ;
      RECT 27.85 10.05 28.025 10.6 ;
      RECT 27.85 7.31 28.02 10.6 ;
      RECT 27.85 7.31 28.025 8.45 ;
      RECT 27.42 7.31 27.59 9.52 ;
      RECT 27.42 7.31 27.595 8.57 ;
      RECT 27.155 3.97 27.325 4.24 ;
      RECT 26.915 3.97 27.325 4.14 ;
      RECT 26.835 3.87 27.165 4.04 ;
      RECT 26.675 4.91 27.325 5.08 ;
      RECT 27.155 4.44 27.325 5.08 ;
      RECT 27.035 4.52 27.325 5.08 ;
      RECT 26.465 10.11 26.64 10.6 ;
      RECT 26.465 7.31 26.635 10.6 ;
      RECT 26.465 9.61 26.875 9.94 ;
      RECT 26.465 8.77 26.875 9.1 ;
      RECT 26.465 7.31 26.64 8.57 ;
      RECT 25.715 4.21 25.885 4.52 ;
      RECT 25.715 4.21 26.605 4.38 ;
      RECT 26.435 3.79 26.605 4.38 ;
      RECT 25.715 3.87 26.205 4.04 ;
      RECT 25.715 3.79 25.885 4.04 ;
      RECT 23.675 4.52 24.165 4.69 ;
      RECT 24.835 3.87 25.005 4.52 ;
      RECT 23.995 4.35 25.005 4.52 ;
      RECT 24.955 3.79 25.125 4.12 ;
      RECT 23.755 3.13 23.925 3.4 ;
      RECT 23.195 3.13 23.925 3.3 ;
      RECT 23.275 3.87 23.445 4.52 ;
      RECT 23.275 3.87 23.765 4.04 ;
      RECT 22.435 3.87 22.925 4.04 ;
      RECT 22.755 3.79 22.925 4.04 ;
      RECT 22.275 3.13 22.445 3.4 ;
      RECT 21.715 3.13 22.445 3.3 ;
      RECT 21.795 4.52 21.965 4.8 ;
      RECT 20.755 4.52 22.045 4.69 ;
      RECT 20.75 3.87 21.325 4.04 ;
      RECT 20.75 3.79 20.92 4.04 ;
      RECT 19.835 3.13 20.005 3.4 ;
      RECT 19.835 3.13 20.565 3.3 ;
      RECT 19.835 4.35 20.005 4.77 ;
      RECT 19.215 4.435 20.005 4.605 ;
      RECT 19.215 4.21 19.385 4.605 ;
      RECT 19.115 3.79 19.285 4.38 ;
      RECT 18.875 3.87 19.285 4.14 ;
      RECT 16.605 7.31 16.775 9.52 ;
      RECT 16.605 7.31 16.78 8.57 ;
      RECT 16.175 10.15 16.345 10.6 ;
      RECT 16.235 8.37 16.405 10.32 ;
      RECT 16.175 7.31 16.345 8.54 ;
      RECT 15.65 10.11 15.825 10.6 ;
      RECT 15.65 7.31 15.82 10.6 ;
      RECT 15.65 9.61 16.06 9.94 ;
      RECT 15.65 8.77 16.06 9.1 ;
      RECT 15.65 7.31 15.825 8.57 ;
      RECT 110.055 10.085 110.23 10.595 ;
      RECT 109.065 1.87 109.24 2.38 ;
      RECT 109.065 10.085 109.24 10.595 ;
      RECT 107.275 1.865 107.45 2.375 ;
      RECT 107.275 10.09 107.45 10.6 ;
      RECT 103.595 3.79 103.765 4.24 ;
      RECT 103.355 3.05 103.525 3.4 ;
      RECT 102.395 3.05 102.565 3.4 ;
      RECT 101.915 4.35 102.085 4.77 ;
      RECT 101.66 10.09 101.835 10.6 ;
      RECT 100.915 3.05 101.085 3.4 ;
      RECT 99.955 3.05 100.125 3.4 ;
      RECT 99.955 4.78 100.125 5.11 ;
      RECT 99.435 4.44 99.605 5.08 ;
      RECT 98.955 3.05 99.125 3.4 ;
      RECT 98.715 3.79 98.885 4.12 ;
      RECT 98.235 3.79 98.405 4.12 ;
      RECT 96.995 4.44 97.165 4.8 ;
      RECT 96.515 4.35 96.685 4.77 ;
      RECT 95.795 3.79 95.965 4.24 ;
      RECT 93.835 3.79 94.005 4.12 ;
      RECT 93.115 3.05 93.285 3.4 ;
      RECT 93.115 4.58 93.285 4.94 ;
      RECT 91.495 10.085 91.67 10.595 ;
      RECT 90.505 1.87 90.68 2.38 ;
      RECT 90.505 10.085 90.68 10.595 ;
      RECT 88.715 1.865 88.89 2.375 ;
      RECT 88.715 10.09 88.89 10.6 ;
      RECT 85.035 3.79 85.205 4.24 ;
      RECT 84.795 3.05 84.965 3.4 ;
      RECT 83.835 3.05 84.005 3.4 ;
      RECT 83.355 4.35 83.525 4.77 ;
      RECT 83.1 10.09 83.275 10.6 ;
      RECT 82.355 3.05 82.525 3.4 ;
      RECT 81.395 3.05 81.565 3.4 ;
      RECT 81.395 4.78 81.565 5.11 ;
      RECT 80.875 4.44 81.045 5.08 ;
      RECT 80.395 3.05 80.565 3.4 ;
      RECT 80.155 3.79 80.325 4.12 ;
      RECT 79.675 3.79 79.845 4.12 ;
      RECT 78.435 4.44 78.605 4.8 ;
      RECT 77.955 4.35 78.125 4.77 ;
      RECT 77.235 3.79 77.405 4.24 ;
      RECT 75.275 3.79 75.445 4.12 ;
      RECT 74.555 3.05 74.725 3.4 ;
      RECT 74.555 4.58 74.725 4.94 ;
      RECT 72.935 10.085 73.11 10.595 ;
      RECT 71.945 1.87 72.12 2.38 ;
      RECT 71.945 10.085 72.12 10.595 ;
      RECT 70.155 1.865 70.33 2.375 ;
      RECT 70.155 10.09 70.33 10.6 ;
      RECT 66.475 3.79 66.645 4.24 ;
      RECT 66.235 3.05 66.405 3.4 ;
      RECT 65.275 3.05 65.445 3.4 ;
      RECT 64.795 4.35 64.965 4.77 ;
      RECT 64.54 10.09 64.715 10.6 ;
      RECT 63.795 3.05 63.965 3.4 ;
      RECT 62.835 3.05 63.005 3.4 ;
      RECT 62.835 4.78 63.005 5.11 ;
      RECT 62.315 4.44 62.485 5.08 ;
      RECT 61.835 3.05 62.005 3.4 ;
      RECT 61.595 3.79 61.765 4.12 ;
      RECT 61.115 3.79 61.285 4.12 ;
      RECT 59.875 4.44 60.045 4.8 ;
      RECT 59.395 4.35 59.565 4.77 ;
      RECT 58.675 3.79 58.845 4.24 ;
      RECT 56.715 3.79 56.885 4.12 ;
      RECT 55.995 3.05 56.165 3.4 ;
      RECT 55.995 4.58 56.165 4.94 ;
      RECT 54.375 10.085 54.55 10.595 ;
      RECT 53.385 1.87 53.56 2.38 ;
      RECT 53.385 10.085 53.56 10.595 ;
      RECT 51.595 1.865 51.77 2.375 ;
      RECT 51.595 10.09 51.77 10.6 ;
      RECT 47.915 3.79 48.085 4.24 ;
      RECT 47.675 3.05 47.845 3.4 ;
      RECT 46.715 3.05 46.885 3.4 ;
      RECT 46.235 4.35 46.405 4.77 ;
      RECT 45.98 10.09 46.155 10.6 ;
      RECT 45.235 3.05 45.405 3.4 ;
      RECT 44.275 3.05 44.445 3.4 ;
      RECT 44.275 4.78 44.445 5.11 ;
      RECT 43.755 4.44 43.925 5.08 ;
      RECT 43.275 3.05 43.445 3.4 ;
      RECT 43.035 3.79 43.205 4.12 ;
      RECT 42.555 3.79 42.725 4.12 ;
      RECT 41.315 4.44 41.485 4.8 ;
      RECT 40.835 4.35 41.005 4.77 ;
      RECT 40.115 3.79 40.285 4.24 ;
      RECT 38.155 3.79 38.325 4.12 ;
      RECT 37.435 3.05 37.605 3.4 ;
      RECT 37.435 4.58 37.605 4.94 ;
      RECT 35.815 10.085 35.99 10.595 ;
      RECT 34.825 1.87 35 2.38 ;
      RECT 34.825 10.085 35 10.595 ;
      RECT 33.035 1.865 33.21 2.375 ;
      RECT 33.035 10.09 33.21 10.6 ;
      RECT 29.355 3.79 29.525 4.24 ;
      RECT 29.115 3.05 29.285 3.4 ;
      RECT 28.155 3.05 28.325 3.4 ;
      RECT 27.675 4.35 27.845 4.77 ;
      RECT 27.42 10.09 27.595 10.6 ;
      RECT 26.675 3.05 26.845 3.4 ;
      RECT 25.715 3.05 25.885 3.4 ;
      RECT 25.715 4.78 25.885 5.11 ;
      RECT 25.195 4.44 25.365 5.08 ;
      RECT 24.715 3.05 24.885 3.4 ;
      RECT 24.475 3.79 24.645 4.12 ;
      RECT 23.995 3.79 24.165 4.12 ;
      RECT 22.755 4.44 22.925 4.8 ;
      RECT 22.275 4.35 22.445 4.77 ;
      RECT 21.555 3.79 21.725 4.24 ;
      RECT 19.595 3.79 19.765 4.12 ;
      RECT 18.875 3.05 19.045 3.4 ;
      RECT 18.875 4.58 19.045 4.94 ;
      RECT 16.605 10.09 16.78 10.6 ;
  END
END sky130_osu_ring_oscillator_mpr2et_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2et_8_b0r2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2et_8_b0r2 ;
  SIZE 110.6 BY 12.465 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 35.71 0 36.09 5.265 ;
      LAYER met2 ;
        RECT 35.71 4.885 36.09 5.265 ;
      LAYER li1 ;
        RECT 35.81 1.87 35.985 2.38 ;
        RECT 35.81 3.9 35.985 5.16 ;
        RECT 35.81 3.69 35.98 5.16 ;
      LAYER met1 ;
        RECT 35.725 4.93 36.075 5.22 ;
        RECT 35.75 2.18 36.045 2.41 ;
        RECT 35.75 3.66 36.04 3.89 ;
        RECT 35.81 2.18 35.98 3.89 ;
      LAYER via1 ;
        RECT 35.825 5 35.975 5.15 ;
      LAYER via2 ;
        RECT 35.8 4.975 36 5.175 ;
      LAYER mcon ;
        RECT 35.81 3.69 35.98 3.86 ;
        RECT 35.81 2.21 35.98 2.38 ;
        RECT 35.815 4.99 35.985 5.16 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 54.27 0 54.65 5.265 ;
      LAYER met2 ;
        RECT 54.27 4.885 54.65 5.265 ;
      LAYER li1 ;
        RECT 54.37 1.87 54.545 2.38 ;
        RECT 54.37 3.9 54.545 5.16 ;
        RECT 54.37 3.69 54.54 5.16 ;
      LAYER met1 ;
        RECT 54.285 4.93 54.635 5.22 ;
        RECT 54.31 2.18 54.605 2.41 ;
        RECT 54.31 3.66 54.6 3.89 ;
        RECT 54.37 2.18 54.54 3.89 ;
      LAYER via1 ;
        RECT 54.385 5 54.535 5.15 ;
      LAYER via2 ;
        RECT 54.36 4.975 54.56 5.175 ;
      LAYER mcon ;
        RECT 54.37 3.69 54.54 3.86 ;
        RECT 54.37 2.21 54.54 2.38 ;
        RECT 54.375 4.99 54.545 5.16 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 72.83 0 73.21 5.265 ;
      LAYER met2 ;
        RECT 72.83 4.885 73.21 5.265 ;
      LAYER li1 ;
        RECT 72.93 1.87 73.105 2.38 ;
        RECT 72.93 3.9 73.105 5.16 ;
        RECT 72.93 3.69 73.1 5.16 ;
      LAYER met1 ;
        RECT 72.845 4.93 73.195 5.22 ;
        RECT 72.87 2.18 73.165 2.41 ;
        RECT 72.87 3.66 73.16 3.89 ;
        RECT 72.93 2.18 73.1 3.89 ;
      LAYER via1 ;
        RECT 72.945 5 73.095 5.15 ;
      LAYER via2 ;
        RECT 72.92 4.975 73.12 5.175 ;
      LAYER mcon ;
        RECT 72.93 3.69 73.1 3.86 ;
        RECT 72.93 2.21 73.1 2.38 ;
        RECT 72.935 4.99 73.105 5.16 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 91.39 0 91.77 5.265 ;
      LAYER met2 ;
        RECT 91.39 4.885 91.77 5.265 ;
      LAYER li1 ;
        RECT 91.49 1.87 91.665 2.38 ;
        RECT 91.49 3.9 91.665 5.16 ;
        RECT 91.49 3.69 91.66 5.16 ;
      LAYER met1 ;
        RECT 91.405 4.93 91.755 5.22 ;
        RECT 91.43 2.18 91.725 2.41 ;
        RECT 91.43 3.66 91.72 3.89 ;
        RECT 91.49 2.18 91.66 3.89 ;
      LAYER via1 ;
        RECT 91.505 5 91.655 5.15 ;
      LAYER via2 ;
        RECT 91.48 4.975 91.68 5.175 ;
      LAYER mcon ;
        RECT 91.49 3.69 91.66 3.86 ;
        RECT 91.49 2.21 91.66 2.38 ;
        RECT 91.495 4.99 91.665 5.16 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 109.95 0 110.33 5.265 ;
      LAYER met2 ;
        RECT 109.95 4.885 110.33 5.265 ;
      LAYER li1 ;
        RECT 110.05 1.87 110.225 2.38 ;
        RECT 110.05 3.9 110.225 5.16 ;
        RECT 110.05 3.69 110.22 5.16 ;
      LAYER met1 ;
        RECT 109.965 4.93 110.315 5.22 ;
        RECT 109.99 2.18 110.285 2.41 ;
        RECT 109.99 3.66 110.28 3.89 ;
        RECT 110.05 2.18 110.22 3.89 ;
      LAYER via1 ;
        RECT 110.065 5 110.215 5.15 ;
      LAYER via2 ;
        RECT 110.04 4.975 110.24 5.175 ;
      LAYER mcon ;
        RECT 110.05 3.69 110.22 3.86 ;
        RECT 110.05 2.21 110.22 2.38 ;
        RECT 110.055 4.99 110.225 5.16 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 31.585 4 31.925 4.35 ;
        RECT 31.575 8.135 31.915 8.485 ;
        RECT 31.66 4 31.83 8.485 ;
      LAYER li1 ;
        RECT 31.655 2.955 31.825 4.225 ;
        RECT 31.655 8.24 31.825 9.51 ;
        RECT 26.04 8.24 26.21 9.51 ;
      LAYER met1 ;
        RECT 25.98 8.235 32.06 8.405 ;
        RECT 31.575 8.235 32.055 8.41 ;
        RECT 31.575 8.135 31.915 8.485 ;
        RECT 25.98 8.235 26.44 8.41 ;
        RECT 25.98 8.21 26.27 8.44 ;
        RECT 31.585 4.055 32.055 4.225 ;
        RECT 31.585 4 31.925 4.35 ;
      LAYER via1 ;
        RECT 31.675 8.235 31.825 8.385 ;
        RECT 31.685 4.1 31.835 4.25 ;
      LAYER mcon ;
        RECT 26.04 8.24 26.21 8.41 ;
        RECT 31.655 8.24 31.825 8.41 ;
        RECT 31.655 4.055 31.825 4.225 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 50.145 4 50.485 4.35 ;
        RECT 50.135 8.135 50.475 8.485 ;
        RECT 50.22 4 50.39 8.485 ;
      LAYER li1 ;
        RECT 50.215 2.955 50.385 4.225 ;
        RECT 50.215 8.24 50.385 9.51 ;
        RECT 44.6 8.24 44.77 9.51 ;
      LAYER met1 ;
        RECT 44.54 8.235 50.62 8.405 ;
        RECT 50.135 8.235 50.615 8.41 ;
        RECT 50.135 8.135 50.475 8.485 ;
        RECT 44.54 8.235 45 8.41 ;
        RECT 44.54 8.21 44.83 8.44 ;
        RECT 50.145 4.055 50.615 4.225 ;
        RECT 50.145 4 50.485 4.35 ;
      LAYER via1 ;
        RECT 50.235 8.235 50.385 8.385 ;
        RECT 50.245 4.1 50.395 4.25 ;
      LAYER mcon ;
        RECT 44.6 8.24 44.77 8.41 ;
        RECT 50.215 8.24 50.385 8.41 ;
        RECT 50.215 4.055 50.385 4.225 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 68.705 4 69.045 4.35 ;
        RECT 68.695 8.135 69.035 8.485 ;
        RECT 68.78 4 68.95 8.485 ;
      LAYER li1 ;
        RECT 68.775 2.955 68.945 4.225 ;
        RECT 68.775 8.24 68.945 9.51 ;
        RECT 63.16 8.24 63.33 9.51 ;
      LAYER met1 ;
        RECT 63.1 8.235 69.18 8.405 ;
        RECT 68.695 8.235 69.175 8.41 ;
        RECT 68.695 8.135 69.035 8.485 ;
        RECT 63.1 8.235 63.56 8.41 ;
        RECT 63.1 8.21 63.39 8.44 ;
        RECT 68.705 4.055 69.175 4.225 ;
        RECT 68.705 4 69.045 4.35 ;
      LAYER via1 ;
        RECT 68.795 8.235 68.945 8.385 ;
        RECT 68.805 4.1 68.955 4.25 ;
      LAYER mcon ;
        RECT 63.16 8.24 63.33 8.41 ;
        RECT 68.775 8.24 68.945 8.41 ;
        RECT 68.775 4.055 68.945 4.225 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 87.265 4 87.605 4.35 ;
        RECT 87.255 8.135 87.595 8.485 ;
        RECT 87.34 4 87.51 8.485 ;
      LAYER li1 ;
        RECT 87.335 2.955 87.505 4.225 ;
        RECT 87.335 8.24 87.505 9.51 ;
        RECT 81.72 8.24 81.89 9.51 ;
      LAYER met1 ;
        RECT 81.66 8.235 87.74 8.405 ;
        RECT 87.255 8.235 87.735 8.41 ;
        RECT 87.255 8.135 87.595 8.485 ;
        RECT 81.66 8.235 82.12 8.41 ;
        RECT 81.66 8.21 81.95 8.44 ;
        RECT 87.265 4.055 87.735 4.225 ;
        RECT 87.265 4 87.605 4.35 ;
      LAYER via1 ;
        RECT 87.355 8.235 87.505 8.385 ;
        RECT 87.365 4.1 87.515 4.25 ;
      LAYER mcon ;
        RECT 81.72 8.24 81.89 8.41 ;
        RECT 87.335 8.24 87.505 8.41 ;
        RECT 87.335 4.055 87.505 4.225 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 105.825 4 106.165 4.35 ;
        RECT 105.815 8.135 106.155 8.485 ;
        RECT 105.9 4 106.07 8.485 ;
      LAYER li1 ;
        RECT 105.895 2.955 106.065 4.225 ;
        RECT 105.895 8.24 106.065 9.51 ;
        RECT 100.28 8.24 100.45 9.51 ;
      LAYER met1 ;
        RECT 100.22 8.235 106.3 8.405 ;
        RECT 105.815 8.235 106.295 8.41 ;
        RECT 105.815 8.135 106.155 8.485 ;
        RECT 100.22 8.235 100.68 8.41 ;
        RECT 100.22 8.21 100.51 8.44 ;
        RECT 105.825 4.055 106.295 4.225 ;
        RECT 105.825 4 106.165 4.35 ;
      LAYER via1 ;
        RECT 105.915 8.235 106.065 8.385 ;
        RECT 105.925 4.1 106.075 4.25 ;
      LAYER mcon ;
        RECT 100.28 8.24 100.45 8.41 ;
        RECT 105.895 8.24 106.065 8.41 ;
        RECT 105.895 4.055 106.065 4.225 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 15.225 8.24 15.395 9.51 ;
      LAYER met1 ;
        RECT 15.14 8.24 15.625 8.41 ;
        RECT 15.14 8.195 15.48 8.455 ;
      LAYER mcon ;
        RECT 15.225 8.24 15.395 8.41 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 92.78 5.43 110.595 7.035 ;
        RECT 0 5.44 110.495 7.04 ;
        RECT 109.625 5.43 109.795 7.765 ;
        RECT 109.62 4.7 109.79 7.04 ;
        RECT 105.715 5.425 109.45 7.04 ;
        RECT 108.63 4.695 108.8 7.77 ;
        RECT 105.885 4.695 106.055 7.77 ;
        RECT 102.87 4.93 103.04 7.04 ;
        RECT 100.43 4.93 100.6 7.04 ;
        RECT 100.27 5.43 100.44 7.77 ;
        RECT 98.47 4.93 98.64 7.04 ;
        RECT 97.51 4.93 97.68 7.04 ;
        RECT 95.55 4.93 95.72 7.04 ;
        RECT 94.55 4.93 94.72 7.04 ;
        RECT 93.59 4.93 93.76 7.04 ;
        RECT 74.22 5.43 92.035 7.04 ;
        RECT 91.065 5.43 91.235 7.765 ;
        RECT 91.06 4.7 91.23 7.04 ;
        RECT 87.155 5.425 90.89 7.04 ;
        RECT 90.07 4.695 90.24 7.77 ;
        RECT 87.325 4.695 87.495 7.77 ;
        RECT 84.31 4.93 84.48 7.04 ;
        RECT 81.87 4.93 82.04 7.04 ;
        RECT 81.71 5.43 81.88 7.77 ;
        RECT 79.91 4.93 80.08 7.04 ;
        RECT 78.95 4.93 79.12 7.04 ;
        RECT 76.99 4.93 77.16 7.04 ;
        RECT 75.99 4.93 76.16 7.04 ;
        RECT 75.03 4.93 75.2 7.04 ;
        RECT 55.66 5.43 73.475 7.04 ;
        RECT 72.505 5.43 72.675 7.765 ;
        RECT 72.5 4.7 72.67 7.04 ;
        RECT 68.595 5.425 72.33 7.04 ;
        RECT 71.51 4.695 71.68 7.77 ;
        RECT 68.765 4.695 68.935 7.77 ;
        RECT 65.75 4.93 65.92 7.04 ;
        RECT 63.31 4.93 63.48 7.04 ;
        RECT 63.15 5.43 63.32 7.77 ;
        RECT 61.35 4.93 61.52 7.04 ;
        RECT 60.39 4.93 60.56 7.04 ;
        RECT 58.43 4.93 58.6 7.04 ;
        RECT 57.43 4.93 57.6 7.04 ;
        RECT 56.47 4.93 56.64 7.04 ;
        RECT 37.1 5.43 54.915 7.04 ;
        RECT 53.945 5.43 54.115 7.765 ;
        RECT 53.94 4.7 54.11 7.04 ;
        RECT 50.035 5.425 53.77 7.04 ;
        RECT 52.95 4.695 53.12 7.77 ;
        RECT 50.205 4.695 50.375 7.77 ;
        RECT 47.19 4.93 47.36 7.04 ;
        RECT 44.75 4.93 44.92 7.04 ;
        RECT 44.59 5.43 44.76 7.77 ;
        RECT 42.79 4.93 42.96 7.04 ;
        RECT 41.83 4.93 42 7.04 ;
        RECT 39.87 4.93 40.04 7.04 ;
        RECT 38.87 4.93 39.04 7.04 ;
        RECT 37.91 4.93 38.08 7.04 ;
        RECT 18.54 5.43 36.355 7.04 ;
        RECT 35.385 5.43 35.555 7.765 ;
        RECT 35.38 4.7 35.55 7.04 ;
        RECT 31.475 5.425 35.21 7.04 ;
        RECT 34.39 4.695 34.56 7.77 ;
        RECT 31.645 4.695 31.815 7.77 ;
        RECT 28.63 4.93 28.8 7.04 ;
        RECT 26.19 4.93 26.36 7.04 ;
        RECT 26.03 5.43 26.2 7.77 ;
        RECT 24.23 4.93 24.4 7.04 ;
        RECT 23.27 4.93 23.44 7.04 ;
        RECT 21.31 4.93 21.48 7.04 ;
        RECT 20.31 4.93 20.48 7.04 ;
        RECT 19.35 4.93 19.52 7.04 ;
        RECT 17.03 10.05 17.205 10.6 ;
        RECT 17.03 7.31 17.205 8.45 ;
        RECT 17.03 5.44 17.2 10.6 ;
        RECT 15.215 5.44 15.385 7.77 ;
      LAYER met1 ;
        RECT 92.78 5.43 110.595 7.035 ;
        RECT 0 5.44 110.495 7.04 ;
        RECT 105.715 5.425 109.45 7.04 ;
        RECT 92.78 5.4 104.74 7.04 ;
        RECT 74.22 5.43 92.035 7.04 ;
        RECT 87.155 5.425 90.89 7.04 ;
        RECT 74.22 5.4 86.18 7.04 ;
        RECT 55.66 5.43 73.475 7.04 ;
        RECT 68.595 5.425 72.33 7.04 ;
        RECT 55.66 5.4 67.62 7.04 ;
        RECT 37.1 5.43 54.915 7.04 ;
        RECT 50.035 5.425 53.77 7.04 ;
        RECT 37.1 5.4 49.06 7.04 ;
        RECT 18.54 5.43 36.355 7.04 ;
        RECT 31.475 5.425 35.21 7.04 ;
        RECT 18.54 5.4 30.5 7.04 ;
        RECT 16.97 8.95 17.26 9.18 ;
        RECT 16.8 8.98 17.26 9.15 ;
      LAYER mcon ;
        RECT 17.03 8.98 17.2 9.15 ;
        RECT 17.335 6.84 17.505 7.01 ;
        RECT 18.685 5.43 18.855 5.6 ;
        RECT 19.145 5.43 19.315 5.6 ;
        RECT 19.605 5.43 19.775 5.6 ;
        RECT 20.065 5.43 20.235 5.6 ;
        RECT 20.525 5.43 20.695 5.6 ;
        RECT 20.985 5.43 21.155 5.6 ;
        RECT 21.445 5.43 21.615 5.6 ;
        RECT 21.905 5.43 22.075 5.6 ;
        RECT 22.365 5.43 22.535 5.6 ;
        RECT 22.825 5.43 22.995 5.6 ;
        RECT 23.285 5.43 23.455 5.6 ;
        RECT 23.745 5.43 23.915 5.6 ;
        RECT 24.205 5.43 24.375 5.6 ;
        RECT 24.665 5.43 24.835 5.6 ;
        RECT 25.125 5.43 25.295 5.6 ;
        RECT 25.585 5.43 25.755 5.6 ;
        RECT 26.045 5.43 26.215 5.6 ;
        RECT 26.505 5.43 26.675 5.6 ;
        RECT 26.965 5.43 27.135 5.6 ;
        RECT 27.425 5.43 27.595 5.6 ;
        RECT 27.885 5.43 28.055 5.6 ;
        RECT 28.15 6.84 28.32 7.01 ;
        RECT 28.345 5.43 28.515 5.6 ;
        RECT 28.805 5.43 28.975 5.6 ;
        RECT 29.265 5.43 29.435 5.6 ;
        RECT 29.725 5.43 29.895 5.6 ;
        RECT 30.185 5.43 30.355 5.6 ;
        RECT 33.765 6.84 33.935 7.01 ;
        RECT 33.765 5.455 33.935 5.625 ;
        RECT 34.47 6.84 34.64 7.01 ;
        RECT 34.47 5.455 34.64 5.625 ;
        RECT 35.46 5.46 35.63 5.63 ;
        RECT 35.465 6.835 35.635 7.005 ;
        RECT 37.245 5.43 37.415 5.6 ;
        RECT 37.705 5.43 37.875 5.6 ;
        RECT 38.165 5.43 38.335 5.6 ;
        RECT 38.625 5.43 38.795 5.6 ;
        RECT 39.085 5.43 39.255 5.6 ;
        RECT 39.545 5.43 39.715 5.6 ;
        RECT 40.005 5.43 40.175 5.6 ;
        RECT 40.465 5.43 40.635 5.6 ;
        RECT 40.925 5.43 41.095 5.6 ;
        RECT 41.385 5.43 41.555 5.6 ;
        RECT 41.845 5.43 42.015 5.6 ;
        RECT 42.305 5.43 42.475 5.6 ;
        RECT 42.765 5.43 42.935 5.6 ;
        RECT 43.225 5.43 43.395 5.6 ;
        RECT 43.685 5.43 43.855 5.6 ;
        RECT 44.145 5.43 44.315 5.6 ;
        RECT 44.605 5.43 44.775 5.6 ;
        RECT 45.065 5.43 45.235 5.6 ;
        RECT 45.525 5.43 45.695 5.6 ;
        RECT 45.985 5.43 46.155 5.6 ;
        RECT 46.445 5.43 46.615 5.6 ;
        RECT 46.71 6.84 46.88 7.01 ;
        RECT 46.905 5.43 47.075 5.6 ;
        RECT 47.365 5.43 47.535 5.6 ;
        RECT 47.825 5.43 47.995 5.6 ;
        RECT 48.285 5.43 48.455 5.6 ;
        RECT 48.745 5.43 48.915 5.6 ;
        RECT 52.325 6.84 52.495 7.01 ;
        RECT 52.325 5.455 52.495 5.625 ;
        RECT 53.03 6.84 53.2 7.01 ;
        RECT 53.03 5.455 53.2 5.625 ;
        RECT 54.02 5.46 54.19 5.63 ;
        RECT 54.025 6.835 54.195 7.005 ;
        RECT 55.805 5.43 55.975 5.6 ;
        RECT 56.265 5.43 56.435 5.6 ;
        RECT 56.725 5.43 56.895 5.6 ;
        RECT 57.185 5.43 57.355 5.6 ;
        RECT 57.645 5.43 57.815 5.6 ;
        RECT 58.105 5.43 58.275 5.6 ;
        RECT 58.565 5.43 58.735 5.6 ;
        RECT 59.025 5.43 59.195 5.6 ;
        RECT 59.485 5.43 59.655 5.6 ;
        RECT 59.945 5.43 60.115 5.6 ;
        RECT 60.405 5.43 60.575 5.6 ;
        RECT 60.865 5.43 61.035 5.6 ;
        RECT 61.325 5.43 61.495 5.6 ;
        RECT 61.785 5.43 61.955 5.6 ;
        RECT 62.245 5.43 62.415 5.6 ;
        RECT 62.705 5.43 62.875 5.6 ;
        RECT 63.165 5.43 63.335 5.6 ;
        RECT 63.625 5.43 63.795 5.6 ;
        RECT 64.085 5.43 64.255 5.6 ;
        RECT 64.545 5.43 64.715 5.6 ;
        RECT 65.005 5.43 65.175 5.6 ;
        RECT 65.27 6.84 65.44 7.01 ;
        RECT 65.465 5.43 65.635 5.6 ;
        RECT 65.925 5.43 66.095 5.6 ;
        RECT 66.385 5.43 66.555 5.6 ;
        RECT 66.845 5.43 67.015 5.6 ;
        RECT 67.305 5.43 67.475 5.6 ;
        RECT 70.885 6.84 71.055 7.01 ;
        RECT 70.885 5.455 71.055 5.625 ;
        RECT 71.59 6.84 71.76 7.01 ;
        RECT 71.59 5.455 71.76 5.625 ;
        RECT 72.58 5.46 72.75 5.63 ;
        RECT 72.585 6.835 72.755 7.005 ;
        RECT 74.365 5.43 74.535 5.6 ;
        RECT 74.825 5.43 74.995 5.6 ;
        RECT 75.285 5.43 75.455 5.6 ;
        RECT 75.745 5.43 75.915 5.6 ;
        RECT 76.205 5.43 76.375 5.6 ;
        RECT 76.665 5.43 76.835 5.6 ;
        RECT 77.125 5.43 77.295 5.6 ;
        RECT 77.585 5.43 77.755 5.6 ;
        RECT 78.045 5.43 78.215 5.6 ;
        RECT 78.505 5.43 78.675 5.6 ;
        RECT 78.965 5.43 79.135 5.6 ;
        RECT 79.425 5.43 79.595 5.6 ;
        RECT 79.885 5.43 80.055 5.6 ;
        RECT 80.345 5.43 80.515 5.6 ;
        RECT 80.805 5.43 80.975 5.6 ;
        RECT 81.265 5.43 81.435 5.6 ;
        RECT 81.725 5.43 81.895 5.6 ;
        RECT 82.185 5.43 82.355 5.6 ;
        RECT 82.645 5.43 82.815 5.6 ;
        RECT 83.105 5.43 83.275 5.6 ;
        RECT 83.565 5.43 83.735 5.6 ;
        RECT 83.83 6.84 84 7.01 ;
        RECT 84.025 5.43 84.195 5.6 ;
        RECT 84.485 5.43 84.655 5.6 ;
        RECT 84.945 5.43 85.115 5.6 ;
        RECT 85.405 5.43 85.575 5.6 ;
        RECT 85.865 5.43 86.035 5.6 ;
        RECT 89.445 6.84 89.615 7.01 ;
        RECT 89.445 5.455 89.615 5.625 ;
        RECT 90.15 6.84 90.32 7.01 ;
        RECT 90.15 5.455 90.32 5.625 ;
        RECT 91.14 5.46 91.31 5.63 ;
        RECT 91.145 6.835 91.315 7.005 ;
        RECT 92.925 5.43 93.095 5.6 ;
        RECT 93.385 5.43 93.555 5.6 ;
        RECT 93.845 5.43 94.015 5.6 ;
        RECT 94.305 5.43 94.475 5.6 ;
        RECT 94.765 5.43 94.935 5.6 ;
        RECT 95.225 5.43 95.395 5.6 ;
        RECT 95.685 5.43 95.855 5.6 ;
        RECT 96.145 5.43 96.315 5.6 ;
        RECT 96.605 5.43 96.775 5.6 ;
        RECT 97.065 5.43 97.235 5.6 ;
        RECT 97.525 5.43 97.695 5.6 ;
        RECT 97.985 5.43 98.155 5.6 ;
        RECT 98.445 5.43 98.615 5.6 ;
        RECT 98.905 5.43 99.075 5.6 ;
        RECT 99.365 5.43 99.535 5.6 ;
        RECT 99.825 5.43 99.995 5.6 ;
        RECT 100.285 5.43 100.455 5.6 ;
        RECT 100.745 5.43 100.915 5.6 ;
        RECT 101.205 5.43 101.375 5.6 ;
        RECT 101.665 5.43 101.835 5.6 ;
        RECT 102.125 5.43 102.295 5.6 ;
        RECT 102.39 6.84 102.56 7.01 ;
        RECT 102.585 5.43 102.755 5.6 ;
        RECT 103.045 5.43 103.215 5.6 ;
        RECT 103.505 5.43 103.675 5.6 ;
        RECT 103.965 5.43 104.135 5.6 ;
        RECT 104.425 5.43 104.595 5.6 ;
        RECT 108.005 6.84 108.175 7.01 ;
        RECT 108.005 5.455 108.175 5.625 ;
        RECT 108.71 6.84 108.88 7.01 ;
        RECT 108.71 5.455 108.88 5.625 ;
        RECT 109.7 5.46 109.87 5.63 ;
        RECT 109.705 6.835 109.875 7.005 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 94.395 3.71 95.125 4.04 ;
        RECT 75.835 3.71 76.565 4.04 ;
        RECT 57.275 3.71 58.005 4.04 ;
        RECT 38.715 3.71 39.445 4.04 ;
        RECT 20.155 3.71 20.885 4.04 ;
      LAYER met2 ;
        RECT 96.225 3.715 96.485 4.035 ;
        RECT 94.445 3.805 96.485 3.945 ;
        RECT 94.825 2.295 95.165 2.635 ;
        RECT 94.755 3.69 95.035 4.06 ;
        RECT 94.85 2.295 95.02 4.06 ;
        RECT 94.505 4.275 94.765 4.595 ;
        RECT 94.445 3.805 94.585 4.505 ;
        RECT 77.665 3.715 77.925 4.035 ;
        RECT 75.885 3.805 77.925 3.945 ;
        RECT 76.265 2.295 76.605 2.635 ;
        RECT 76.195 3.69 76.475 4.06 ;
        RECT 76.29 2.295 76.46 4.06 ;
        RECT 75.945 4.275 76.205 4.595 ;
        RECT 75.885 3.805 76.025 4.505 ;
        RECT 59.105 3.715 59.365 4.035 ;
        RECT 57.325 3.805 59.365 3.945 ;
        RECT 57.705 2.295 58.045 2.635 ;
        RECT 57.635 3.69 57.915 4.06 ;
        RECT 57.73 2.295 57.9 4.06 ;
        RECT 57.385 4.275 57.645 4.595 ;
        RECT 57.325 3.805 57.465 4.505 ;
        RECT 40.545 3.715 40.805 4.035 ;
        RECT 38.765 3.805 40.805 3.945 ;
        RECT 39.145 2.295 39.485 2.635 ;
        RECT 39.075 3.69 39.355 4.06 ;
        RECT 39.17 2.295 39.34 4.06 ;
        RECT 38.825 4.275 39.085 4.595 ;
        RECT 38.765 3.805 38.905 4.505 ;
        RECT 21.985 3.715 22.245 4.035 ;
        RECT 20.205 3.805 22.245 3.945 ;
        RECT 20.585 2.295 20.925 2.635 ;
        RECT 20.515 3.69 20.795 4.06 ;
        RECT 20.61 2.295 20.78 4.06 ;
        RECT 20.265 4.275 20.525 4.595 ;
        RECT 20.205 3.805 20.345 4.505 ;
      LAYER li1 ;
        RECT 0 10.865 110.6 12.465 ;
        RECT 109.625 10.235 109.795 12.465 ;
        RECT 108.63 10.24 108.8 12.465 ;
        RECT 105.885 10.24 106.055 12.465 ;
        RECT 100.27 10.24 100.44 12.465 ;
        RECT 91.065 10.235 91.235 12.465 ;
        RECT 90.07 10.24 90.24 12.465 ;
        RECT 87.325 10.24 87.495 12.465 ;
        RECT 81.71 10.24 81.88 12.465 ;
        RECT 72.505 10.235 72.675 12.465 ;
        RECT 71.51 10.24 71.68 12.465 ;
        RECT 68.765 10.24 68.935 12.465 ;
        RECT 63.15 10.24 63.32 12.465 ;
        RECT 53.945 10.235 54.115 12.465 ;
        RECT 52.95 10.24 53.12 12.465 ;
        RECT 50.205 10.24 50.375 12.465 ;
        RECT 44.59 10.24 44.76 12.465 ;
        RECT 35.385 10.235 35.555 12.465 ;
        RECT 34.39 10.24 34.56 12.465 ;
        RECT 31.645 10.24 31.815 12.465 ;
        RECT 26.03 10.24 26.2 12.465 ;
        RECT 15.215 10.24 15.385 12.465 ;
        RECT 0 0 110.595 1.6 ;
        RECT 109.62 0 109.79 2.23 ;
        RECT 108.63 0 108.8 2.225 ;
        RECT 105.885 0 106.055 2.225 ;
        RECT 92.78 0 104.825 2.88 ;
        RECT 103.83 0 104 3.38 ;
        RECT 102.87 0 103.04 3.38 ;
        RECT 101.91 0 102.08 3.38 ;
        RECT 101.39 0 101.56 3.38 ;
        RECT 100.43 0 100.6 3.38 ;
        RECT 99.43 0 99.6 3.38 ;
        RECT 98.47 0 98.64 3.38 ;
        RECT 97.435 0 97.63 2.89 ;
        RECT 96.99 0 97.16 3.38 ;
        RECT 95.07 0 95.33 2.89 ;
        RECT 95.07 0 95.24 3.38 ;
        RECT 93.59 0 93.76 3.38 ;
        RECT 91.06 0 91.23 2.23 ;
        RECT 90.07 0 90.24 2.225 ;
        RECT 87.325 0 87.495 2.225 ;
        RECT 74.22 0 86.265 2.88 ;
        RECT 85.27 0 85.44 3.38 ;
        RECT 84.31 0 84.48 3.38 ;
        RECT 83.35 0 83.52 3.38 ;
        RECT 82.83 0 83 3.38 ;
        RECT 81.87 0 82.04 3.38 ;
        RECT 80.87 0 81.04 3.38 ;
        RECT 79.91 0 80.08 3.38 ;
        RECT 78.875 0 79.07 2.89 ;
        RECT 78.43 0 78.6 3.38 ;
        RECT 76.51 0 76.77 2.89 ;
        RECT 76.51 0 76.68 3.38 ;
        RECT 75.03 0 75.2 3.38 ;
        RECT 72.5 0 72.67 2.23 ;
        RECT 71.51 0 71.68 2.225 ;
        RECT 68.765 0 68.935 2.225 ;
        RECT 55.66 0 67.705 2.88 ;
        RECT 66.71 0 66.88 3.38 ;
        RECT 65.75 0 65.92 3.38 ;
        RECT 64.79 0 64.96 3.38 ;
        RECT 64.27 0 64.44 3.38 ;
        RECT 63.31 0 63.48 3.38 ;
        RECT 62.31 0 62.48 3.38 ;
        RECT 61.35 0 61.52 3.38 ;
        RECT 60.315 0 60.51 2.89 ;
        RECT 59.87 0 60.04 3.38 ;
        RECT 57.95 0 58.21 2.89 ;
        RECT 57.95 0 58.12 3.38 ;
        RECT 56.47 0 56.64 3.38 ;
        RECT 53.94 0 54.11 2.23 ;
        RECT 52.95 0 53.12 2.225 ;
        RECT 50.205 0 50.375 2.225 ;
        RECT 37.1 0 49.145 2.88 ;
        RECT 48.15 0 48.32 3.38 ;
        RECT 47.19 0 47.36 3.38 ;
        RECT 46.23 0 46.4 3.38 ;
        RECT 45.71 0 45.88 3.38 ;
        RECT 44.75 0 44.92 3.38 ;
        RECT 43.75 0 43.92 3.38 ;
        RECT 42.79 0 42.96 3.38 ;
        RECT 41.755 0 41.95 2.89 ;
        RECT 41.31 0 41.48 3.38 ;
        RECT 39.39 0 39.65 2.89 ;
        RECT 39.39 0 39.56 3.38 ;
        RECT 37.91 0 38.08 3.38 ;
        RECT 35.38 0 35.55 2.23 ;
        RECT 34.39 0 34.56 2.225 ;
        RECT 31.645 0 31.815 2.225 ;
        RECT 18.54 0 30.585 2.88 ;
        RECT 29.59 0 29.76 3.38 ;
        RECT 28.63 0 28.8 3.38 ;
        RECT 27.67 0 27.84 3.38 ;
        RECT 27.15 0 27.32 3.38 ;
        RECT 26.19 0 26.36 3.38 ;
        RECT 25.19 0 25.36 3.38 ;
        RECT 24.23 0 24.4 3.38 ;
        RECT 23.195 0 23.39 2.89 ;
        RECT 22.75 0 22.92 3.38 ;
        RECT 20.83 0 21.09 2.89 ;
        RECT 20.83 0 21 3.38 ;
        RECT 19.35 0 19.52 3.38 ;
        RECT 101.285 8.37 101.455 10.32 ;
        RECT 101.225 10.15 101.395 10.6 ;
        RECT 101.225 7.31 101.395 8.54 ;
        RECT 96.27 3.79 96.44 4.12 ;
        RECT 94.43 4.35 94.72 4.52 ;
        RECT 94.43 3.87 94.6 4.52 ;
        RECT 94.23 3.87 94.6 4.04 ;
        RECT 82.725 8.37 82.895 10.32 ;
        RECT 82.665 10.15 82.835 10.6 ;
        RECT 82.665 7.31 82.835 8.54 ;
        RECT 77.71 3.79 77.88 4.12 ;
        RECT 75.87 4.35 76.16 4.52 ;
        RECT 75.87 3.87 76.04 4.52 ;
        RECT 75.67 3.87 76.04 4.04 ;
        RECT 64.165 8.37 64.335 10.32 ;
        RECT 64.105 10.15 64.275 10.6 ;
        RECT 64.105 7.31 64.275 8.54 ;
        RECT 59.15 3.79 59.32 4.12 ;
        RECT 57.31 4.35 57.6 4.52 ;
        RECT 57.31 3.87 57.48 4.52 ;
        RECT 57.11 3.87 57.48 4.04 ;
        RECT 45.605 8.37 45.775 10.32 ;
        RECT 45.545 10.15 45.715 10.6 ;
        RECT 45.545 7.31 45.715 8.54 ;
        RECT 40.59 3.79 40.76 4.12 ;
        RECT 38.75 4.35 39.04 4.52 ;
        RECT 38.75 3.87 38.92 4.52 ;
        RECT 38.55 3.87 38.92 4.04 ;
        RECT 27.045 8.37 27.215 10.32 ;
        RECT 26.985 10.15 27.155 10.6 ;
        RECT 26.985 7.31 27.155 8.54 ;
        RECT 22.03 3.79 22.2 4.12 ;
        RECT 20.19 4.35 20.48 4.52 ;
        RECT 20.19 3.87 20.36 4.52 ;
        RECT 19.99 3.87 20.36 4.04 ;
      LAYER met1 ;
        RECT 0 10.865 110.6 12.465 ;
        RECT 101.225 8.58 101.515 8.81 ;
        RECT 100.785 8.605 101.515 8.78 ;
        RECT 100.785 8.605 100.955 12.465 ;
        RECT 82.665 8.58 82.955 8.81 ;
        RECT 82.225 8.605 82.955 8.78 ;
        RECT 82.225 8.605 82.395 12.465 ;
        RECT 64.105 8.58 64.395 8.81 ;
        RECT 63.665 8.605 64.395 8.78 ;
        RECT 63.665 8.605 63.835 12.465 ;
        RECT 45.545 8.58 45.835 8.81 ;
        RECT 45.105 8.605 45.835 8.78 ;
        RECT 45.105 8.605 45.275 12.465 ;
        RECT 26.985 8.58 27.275 8.81 ;
        RECT 26.545 8.605 27.275 8.78 ;
        RECT 26.545 8.605 26.715 12.465 ;
        RECT 0 0 110.595 1.6 ;
        RECT 92.78 0 104.825 2.88 ;
        RECT 92.78 0 104.74 2.91 ;
        RECT 74.22 0 86.265 2.88 ;
        RECT 74.22 0 86.18 2.91 ;
        RECT 55.66 0 67.705 2.88 ;
        RECT 55.66 0 67.62 2.91 ;
        RECT 37.1 0 49.145 2.88 ;
        RECT 37.1 0 49.06 2.91 ;
        RECT 18.54 0 30.585 2.88 ;
        RECT 18.54 0 30.5 2.91 ;
        RECT 96.21 3.665 96.5 4.035 ;
        RECT 95.445 3.665 96.5 3.805 ;
        RECT 94.475 4.305 94.795 4.565 ;
        RECT 77.65 3.665 77.94 4.035 ;
        RECT 76.885 3.665 77.94 3.805 ;
        RECT 75.915 4.305 76.235 4.565 ;
        RECT 59.09 3.665 59.38 4.035 ;
        RECT 58.325 3.665 59.38 3.805 ;
        RECT 57.355 4.305 57.675 4.565 ;
        RECT 40.53 3.665 40.82 4.035 ;
        RECT 39.765 3.665 40.82 3.805 ;
        RECT 38.795 4.305 39.115 4.565 ;
        RECT 21.97 3.665 22.26 4.035 ;
        RECT 21.205 3.665 22.26 3.805 ;
        RECT 20.235 4.305 20.555 4.565 ;
      LAYER via1 ;
        RECT 20.32 4.36 20.47 4.51 ;
        RECT 20.68 2.39 20.83 2.54 ;
        RECT 22.04 3.8 22.19 3.95 ;
        RECT 38.88 4.36 39.03 4.51 ;
        RECT 39.24 2.39 39.39 2.54 ;
        RECT 40.6 3.8 40.75 3.95 ;
        RECT 57.44 4.36 57.59 4.51 ;
        RECT 57.8 2.39 57.95 2.54 ;
        RECT 59.16 3.8 59.31 3.95 ;
        RECT 76 4.36 76.15 4.51 ;
        RECT 76.36 2.39 76.51 2.54 ;
        RECT 77.72 3.8 77.87 3.95 ;
        RECT 94.56 4.36 94.71 4.51 ;
        RECT 94.92 2.39 95.07 2.54 ;
        RECT 96.28 3.8 96.43 3.95 ;
      LAYER via2 ;
        RECT 20.555 3.775 20.755 3.975 ;
        RECT 39.115 3.775 39.315 3.975 ;
        RECT 57.675 3.775 57.875 3.975 ;
        RECT 76.235 3.775 76.435 3.975 ;
        RECT 94.795 3.775 94.995 3.975 ;
      LAYER mcon ;
        RECT 15.295 10.9 15.465 11.07 ;
        RECT 15.975 10.9 16.145 11.07 ;
        RECT 16.655 10.9 16.825 11.07 ;
        RECT 17.335 10.9 17.505 11.07 ;
        RECT 18.685 2.71 18.855 2.88 ;
        RECT 19.145 2.71 19.315 2.88 ;
        RECT 19.605 2.71 19.775 2.88 ;
        RECT 20.065 2.71 20.235 2.88 ;
        RECT 20.31 4.35 20.48 4.52 ;
        RECT 20.525 2.71 20.695 2.88 ;
        RECT 20.985 2.71 21.155 2.88 ;
        RECT 21.445 2.71 21.615 2.88 ;
        RECT 21.905 2.71 22.075 2.88 ;
        RECT 22.03 3.79 22.2 3.96 ;
        RECT 22.365 2.71 22.535 2.88 ;
        RECT 22.825 2.71 22.995 2.88 ;
        RECT 23.285 2.71 23.455 2.88 ;
        RECT 23.745 2.71 23.915 2.88 ;
        RECT 24.205 2.71 24.375 2.88 ;
        RECT 24.665 2.71 24.835 2.88 ;
        RECT 25.125 2.71 25.295 2.88 ;
        RECT 25.585 2.71 25.755 2.88 ;
        RECT 26.045 2.71 26.215 2.88 ;
        RECT 26.11 10.9 26.28 11.07 ;
        RECT 26.505 2.71 26.675 2.88 ;
        RECT 26.79 10.9 26.96 11.07 ;
        RECT 26.965 2.71 27.135 2.88 ;
        RECT 27.045 8.61 27.215 8.78 ;
        RECT 27.425 2.71 27.595 2.88 ;
        RECT 27.47 10.9 27.64 11.07 ;
        RECT 27.885 2.71 28.055 2.88 ;
        RECT 28.15 10.9 28.32 11.07 ;
        RECT 28.345 2.71 28.515 2.88 ;
        RECT 28.805 2.71 28.975 2.88 ;
        RECT 29.265 2.71 29.435 2.88 ;
        RECT 29.725 2.71 29.895 2.88 ;
        RECT 30.185 2.71 30.355 2.88 ;
        RECT 31.725 10.9 31.895 11.07 ;
        RECT 31.725 1.395 31.895 1.565 ;
        RECT 32.405 10.9 32.575 11.07 ;
        RECT 32.405 1.395 32.575 1.565 ;
        RECT 33.085 10.9 33.255 11.07 ;
        RECT 33.085 1.395 33.255 1.565 ;
        RECT 33.765 10.9 33.935 11.07 ;
        RECT 33.765 1.395 33.935 1.565 ;
        RECT 34.47 10.9 34.64 11.07 ;
        RECT 34.47 1.395 34.64 1.565 ;
        RECT 35.46 1.4 35.63 1.57 ;
        RECT 35.465 10.895 35.635 11.065 ;
        RECT 37.245 2.71 37.415 2.88 ;
        RECT 37.705 2.71 37.875 2.88 ;
        RECT 38.165 2.71 38.335 2.88 ;
        RECT 38.625 2.71 38.795 2.88 ;
        RECT 38.87 4.35 39.04 4.52 ;
        RECT 39.085 2.71 39.255 2.88 ;
        RECT 39.545 2.71 39.715 2.88 ;
        RECT 40.005 2.71 40.175 2.88 ;
        RECT 40.465 2.71 40.635 2.88 ;
        RECT 40.59 3.79 40.76 3.96 ;
        RECT 40.925 2.71 41.095 2.88 ;
        RECT 41.385 2.71 41.555 2.88 ;
        RECT 41.845 2.71 42.015 2.88 ;
        RECT 42.305 2.71 42.475 2.88 ;
        RECT 42.765 2.71 42.935 2.88 ;
        RECT 43.225 2.71 43.395 2.88 ;
        RECT 43.685 2.71 43.855 2.88 ;
        RECT 44.145 2.71 44.315 2.88 ;
        RECT 44.605 2.71 44.775 2.88 ;
        RECT 44.67 10.9 44.84 11.07 ;
        RECT 45.065 2.71 45.235 2.88 ;
        RECT 45.35 10.9 45.52 11.07 ;
        RECT 45.525 2.71 45.695 2.88 ;
        RECT 45.605 8.61 45.775 8.78 ;
        RECT 45.985 2.71 46.155 2.88 ;
        RECT 46.03 10.9 46.2 11.07 ;
        RECT 46.445 2.71 46.615 2.88 ;
        RECT 46.71 10.9 46.88 11.07 ;
        RECT 46.905 2.71 47.075 2.88 ;
        RECT 47.365 2.71 47.535 2.88 ;
        RECT 47.825 2.71 47.995 2.88 ;
        RECT 48.285 2.71 48.455 2.88 ;
        RECT 48.745 2.71 48.915 2.88 ;
        RECT 50.285 10.9 50.455 11.07 ;
        RECT 50.285 1.395 50.455 1.565 ;
        RECT 50.965 10.9 51.135 11.07 ;
        RECT 50.965 1.395 51.135 1.565 ;
        RECT 51.645 10.9 51.815 11.07 ;
        RECT 51.645 1.395 51.815 1.565 ;
        RECT 52.325 10.9 52.495 11.07 ;
        RECT 52.325 1.395 52.495 1.565 ;
        RECT 53.03 10.9 53.2 11.07 ;
        RECT 53.03 1.395 53.2 1.565 ;
        RECT 54.02 1.4 54.19 1.57 ;
        RECT 54.025 10.895 54.195 11.065 ;
        RECT 55.805 2.71 55.975 2.88 ;
        RECT 56.265 2.71 56.435 2.88 ;
        RECT 56.725 2.71 56.895 2.88 ;
        RECT 57.185 2.71 57.355 2.88 ;
        RECT 57.43 4.35 57.6 4.52 ;
        RECT 57.645 2.71 57.815 2.88 ;
        RECT 58.105 2.71 58.275 2.88 ;
        RECT 58.565 2.71 58.735 2.88 ;
        RECT 59.025 2.71 59.195 2.88 ;
        RECT 59.15 3.79 59.32 3.96 ;
        RECT 59.485 2.71 59.655 2.88 ;
        RECT 59.945 2.71 60.115 2.88 ;
        RECT 60.405 2.71 60.575 2.88 ;
        RECT 60.865 2.71 61.035 2.88 ;
        RECT 61.325 2.71 61.495 2.88 ;
        RECT 61.785 2.71 61.955 2.88 ;
        RECT 62.245 2.71 62.415 2.88 ;
        RECT 62.705 2.71 62.875 2.88 ;
        RECT 63.165 2.71 63.335 2.88 ;
        RECT 63.23 10.9 63.4 11.07 ;
        RECT 63.625 2.71 63.795 2.88 ;
        RECT 63.91 10.9 64.08 11.07 ;
        RECT 64.085 2.71 64.255 2.88 ;
        RECT 64.165 8.61 64.335 8.78 ;
        RECT 64.545 2.71 64.715 2.88 ;
        RECT 64.59 10.9 64.76 11.07 ;
        RECT 65.005 2.71 65.175 2.88 ;
        RECT 65.27 10.9 65.44 11.07 ;
        RECT 65.465 2.71 65.635 2.88 ;
        RECT 65.925 2.71 66.095 2.88 ;
        RECT 66.385 2.71 66.555 2.88 ;
        RECT 66.845 2.71 67.015 2.88 ;
        RECT 67.305 2.71 67.475 2.88 ;
        RECT 68.845 10.9 69.015 11.07 ;
        RECT 68.845 1.395 69.015 1.565 ;
        RECT 69.525 10.9 69.695 11.07 ;
        RECT 69.525 1.395 69.695 1.565 ;
        RECT 70.205 10.9 70.375 11.07 ;
        RECT 70.205 1.395 70.375 1.565 ;
        RECT 70.885 10.9 71.055 11.07 ;
        RECT 70.885 1.395 71.055 1.565 ;
        RECT 71.59 10.9 71.76 11.07 ;
        RECT 71.59 1.395 71.76 1.565 ;
        RECT 72.58 1.4 72.75 1.57 ;
        RECT 72.585 10.895 72.755 11.065 ;
        RECT 74.365 2.71 74.535 2.88 ;
        RECT 74.825 2.71 74.995 2.88 ;
        RECT 75.285 2.71 75.455 2.88 ;
        RECT 75.745 2.71 75.915 2.88 ;
        RECT 75.99 4.35 76.16 4.52 ;
        RECT 76.205 2.71 76.375 2.88 ;
        RECT 76.665 2.71 76.835 2.88 ;
        RECT 77.125 2.71 77.295 2.88 ;
        RECT 77.585 2.71 77.755 2.88 ;
        RECT 77.71 3.79 77.88 3.96 ;
        RECT 78.045 2.71 78.215 2.88 ;
        RECT 78.505 2.71 78.675 2.88 ;
        RECT 78.965 2.71 79.135 2.88 ;
        RECT 79.425 2.71 79.595 2.88 ;
        RECT 79.885 2.71 80.055 2.88 ;
        RECT 80.345 2.71 80.515 2.88 ;
        RECT 80.805 2.71 80.975 2.88 ;
        RECT 81.265 2.71 81.435 2.88 ;
        RECT 81.725 2.71 81.895 2.88 ;
        RECT 81.79 10.9 81.96 11.07 ;
        RECT 82.185 2.71 82.355 2.88 ;
        RECT 82.47 10.9 82.64 11.07 ;
        RECT 82.645 2.71 82.815 2.88 ;
        RECT 82.725 8.61 82.895 8.78 ;
        RECT 83.105 2.71 83.275 2.88 ;
        RECT 83.15 10.9 83.32 11.07 ;
        RECT 83.565 2.71 83.735 2.88 ;
        RECT 83.83 10.9 84 11.07 ;
        RECT 84.025 2.71 84.195 2.88 ;
        RECT 84.485 2.71 84.655 2.88 ;
        RECT 84.945 2.71 85.115 2.88 ;
        RECT 85.405 2.71 85.575 2.88 ;
        RECT 85.865 2.71 86.035 2.88 ;
        RECT 87.405 10.9 87.575 11.07 ;
        RECT 87.405 1.395 87.575 1.565 ;
        RECT 88.085 10.9 88.255 11.07 ;
        RECT 88.085 1.395 88.255 1.565 ;
        RECT 88.765 10.9 88.935 11.07 ;
        RECT 88.765 1.395 88.935 1.565 ;
        RECT 89.445 10.9 89.615 11.07 ;
        RECT 89.445 1.395 89.615 1.565 ;
        RECT 90.15 10.9 90.32 11.07 ;
        RECT 90.15 1.395 90.32 1.565 ;
        RECT 91.14 1.4 91.31 1.57 ;
        RECT 91.145 10.895 91.315 11.065 ;
        RECT 92.925 2.71 93.095 2.88 ;
        RECT 93.385 2.71 93.555 2.88 ;
        RECT 93.845 2.71 94.015 2.88 ;
        RECT 94.305 2.71 94.475 2.88 ;
        RECT 94.55 4.35 94.72 4.52 ;
        RECT 94.765 2.71 94.935 2.88 ;
        RECT 95.225 2.71 95.395 2.88 ;
        RECT 95.685 2.71 95.855 2.88 ;
        RECT 96.145 2.71 96.315 2.88 ;
        RECT 96.27 3.79 96.44 3.96 ;
        RECT 96.605 2.71 96.775 2.88 ;
        RECT 97.065 2.71 97.235 2.88 ;
        RECT 97.525 2.71 97.695 2.88 ;
        RECT 97.985 2.71 98.155 2.88 ;
        RECT 98.445 2.71 98.615 2.88 ;
        RECT 98.905 2.71 99.075 2.88 ;
        RECT 99.365 2.71 99.535 2.88 ;
        RECT 99.825 2.71 99.995 2.88 ;
        RECT 100.285 2.71 100.455 2.88 ;
        RECT 100.35 10.9 100.52 11.07 ;
        RECT 100.745 2.71 100.915 2.88 ;
        RECT 101.03 10.9 101.2 11.07 ;
        RECT 101.205 2.71 101.375 2.88 ;
        RECT 101.285 8.61 101.455 8.78 ;
        RECT 101.665 2.71 101.835 2.88 ;
        RECT 101.71 10.9 101.88 11.07 ;
        RECT 102.125 2.71 102.295 2.88 ;
        RECT 102.39 10.9 102.56 11.07 ;
        RECT 102.585 2.71 102.755 2.88 ;
        RECT 103.045 2.71 103.215 2.88 ;
        RECT 103.505 2.71 103.675 2.88 ;
        RECT 103.965 2.71 104.135 2.88 ;
        RECT 104.425 2.71 104.595 2.88 ;
        RECT 105.965 10.9 106.135 11.07 ;
        RECT 105.965 1.395 106.135 1.565 ;
        RECT 106.645 10.9 106.815 11.07 ;
        RECT 106.645 1.395 106.815 1.565 ;
        RECT 107.325 10.9 107.495 11.07 ;
        RECT 107.325 1.395 107.495 1.565 ;
        RECT 108.005 10.9 108.175 11.07 ;
        RECT 108.005 1.395 108.175 1.565 ;
        RECT 108.71 10.9 108.88 11.07 ;
        RECT 108.71 1.395 108.88 1.565 ;
        RECT 109.7 1.4 109.87 1.57 ;
        RECT 109.705 10.895 109.875 11.065 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 102.085 4.83 102.64 5.16 ;
      RECT 102.085 3.165 102.385 5.16 ;
      RECT 98.15 4.27 98.705 4.6 ;
      RECT 98.405 3.165 98.705 4.6 ;
      RECT 98.405 3.165 102.385 3.465 ;
      RECT 101.555 9.345 101.93 9.715 ;
      RECT 101.555 9.385 102.56 9.685 ;
      RECT 102.26 6.695 102.56 9.685 ;
      RECT 92.43 6.695 102.56 6.995 ;
      RECT 96.935 3.71 97.235 6.995 ;
      RECT 95.5 4.27 95.8 6.995 ;
      RECT 92.43 3.715 92.73 6.995 ;
      RECT 95.47 4.27 96.2 4.6 ;
      RECT 96.91 3.71 97.64 4.04 ;
      RECT 93.36 3.71 94.09 4.04 ;
      RECT 92.43 3.715 94.09 4.015 ;
      RECT 83.525 4.83 84.08 5.16 ;
      RECT 83.525 3.165 83.825 5.16 ;
      RECT 79.59 4.27 80.145 4.6 ;
      RECT 79.845 3.165 80.145 4.6 ;
      RECT 79.845 3.165 83.825 3.465 ;
      RECT 82.995 9.345 83.37 9.715 ;
      RECT 82.995 9.385 84 9.685 ;
      RECT 83.7 6.695 84 9.685 ;
      RECT 73.87 6.695 84 6.995 ;
      RECT 78.375 3.71 78.675 6.995 ;
      RECT 76.94 4.27 77.24 6.995 ;
      RECT 73.87 3.715 74.17 6.995 ;
      RECT 76.91 4.27 77.64 4.6 ;
      RECT 78.35 3.71 79.08 4.04 ;
      RECT 74.8 3.71 75.53 4.04 ;
      RECT 73.87 3.715 75.53 4.015 ;
      RECT 64.965 4.83 65.52 5.16 ;
      RECT 64.965 3.165 65.265 5.16 ;
      RECT 61.03 4.27 61.585 4.6 ;
      RECT 61.285 3.165 61.585 4.6 ;
      RECT 61.285 3.165 65.265 3.465 ;
      RECT 64.435 9.345 64.81 9.715 ;
      RECT 64.435 9.385 65.44 9.685 ;
      RECT 65.14 6.695 65.44 9.685 ;
      RECT 55.31 6.695 65.44 6.995 ;
      RECT 59.815 3.71 60.115 6.995 ;
      RECT 58.38 4.27 58.68 6.995 ;
      RECT 55.31 3.715 55.61 6.995 ;
      RECT 58.35 4.27 59.08 4.6 ;
      RECT 59.79 3.71 60.52 4.04 ;
      RECT 56.24 3.71 56.97 4.04 ;
      RECT 55.31 3.715 56.97 4.015 ;
      RECT 46.405 4.83 46.96 5.16 ;
      RECT 46.405 3.165 46.705 5.16 ;
      RECT 42.47 4.27 43.025 4.6 ;
      RECT 42.725 3.165 43.025 4.6 ;
      RECT 42.725 3.165 46.705 3.465 ;
      RECT 45.875 9.345 46.25 9.715 ;
      RECT 45.875 9.385 46.88 9.685 ;
      RECT 46.58 6.695 46.88 9.685 ;
      RECT 36.75 6.695 46.88 6.995 ;
      RECT 41.255 3.71 41.555 6.995 ;
      RECT 39.82 4.27 40.12 6.995 ;
      RECT 36.75 3.715 37.05 6.995 ;
      RECT 39.79 4.27 40.52 4.6 ;
      RECT 41.23 3.71 41.96 4.04 ;
      RECT 37.68 3.71 38.41 4.04 ;
      RECT 36.75 3.715 38.41 4.015 ;
      RECT 27.845 4.83 28.4 5.16 ;
      RECT 27.845 3.165 28.145 5.16 ;
      RECT 23.91 4.27 24.465 4.6 ;
      RECT 24.165 3.165 24.465 4.6 ;
      RECT 24.165 3.165 28.145 3.465 ;
      RECT 27.315 9.345 27.69 9.715 ;
      RECT 27.315 9.385 28.32 9.685 ;
      RECT 28.02 6.695 28.32 9.685 ;
      RECT 18.19 6.695 28.32 6.995 ;
      RECT 22.695 3.71 22.995 6.995 ;
      RECT 21.26 4.27 21.56 6.995 ;
      RECT 18.19 3.715 18.49 6.995 ;
      RECT 21.23 4.27 21.96 4.6 ;
      RECT 22.67 3.71 23.4 4.04 ;
      RECT 19.12 3.71 19.85 4.04 ;
      RECT 18.19 3.715 19.85 4.015 ;
      RECT 109.955 7.2 110.335 12.465 ;
      RECT 103.27 3.15 104 3.48 ;
      RECT 101.05 4.83 101.78 5.16 ;
      RECT 99.35 4.83 100.08 5.16 ;
      RECT 93.03 4.83 93.76 5.16 ;
      RECT 91.395 7.2 91.775 12.465 ;
      RECT 84.71 3.15 85.44 3.48 ;
      RECT 82.49 4.83 83.22 5.16 ;
      RECT 80.79 4.83 81.52 5.16 ;
      RECT 74.47 4.83 75.2 5.16 ;
      RECT 72.835 7.2 73.215 12.465 ;
      RECT 66.15 3.15 66.88 3.48 ;
      RECT 63.93 4.83 64.66 5.16 ;
      RECT 62.23 4.83 62.96 5.16 ;
      RECT 55.91 4.83 56.64 5.16 ;
      RECT 54.275 7.2 54.655 12.465 ;
      RECT 47.59 3.15 48.32 3.48 ;
      RECT 45.37 4.83 46.1 5.16 ;
      RECT 43.67 4.83 44.4 5.16 ;
      RECT 37.35 4.83 38.08 5.16 ;
      RECT 35.715 7.2 36.095 12.465 ;
      RECT 29.03 3.15 29.76 3.48 ;
      RECT 26.81 4.83 27.54 5.16 ;
      RECT 25.11 4.83 25.84 5.16 ;
      RECT 18.79 4.83 19.52 5.16 ;
    LAYER via2 ;
      RECT 110.045 7.29 110.245 7.49 ;
      RECT 103.335 3.215 103.535 3.415 ;
      RECT 102.375 4.895 102.575 5.095 ;
      RECT 101.64 9.43 101.84 9.63 ;
      RECT 101.375 4.895 101.575 5.095 ;
      RECT 99.415 4.895 99.615 5.095 ;
      RECT 98.215 4.335 98.415 4.535 ;
      RECT 96.975 3.775 97.175 3.975 ;
      RECT 95.535 4.335 95.735 4.535 ;
      RECT 93.575 3.775 93.775 3.975 ;
      RECT 93.095 4.895 93.295 5.095 ;
      RECT 91.485 7.29 91.685 7.49 ;
      RECT 84.775 3.215 84.975 3.415 ;
      RECT 83.815 4.895 84.015 5.095 ;
      RECT 83.08 9.43 83.28 9.63 ;
      RECT 82.815 4.895 83.015 5.095 ;
      RECT 80.855 4.895 81.055 5.095 ;
      RECT 79.655 4.335 79.855 4.535 ;
      RECT 78.415 3.775 78.615 3.975 ;
      RECT 76.975 4.335 77.175 4.535 ;
      RECT 75.015 3.775 75.215 3.975 ;
      RECT 74.535 4.895 74.735 5.095 ;
      RECT 72.925 7.29 73.125 7.49 ;
      RECT 66.215 3.215 66.415 3.415 ;
      RECT 65.255 4.895 65.455 5.095 ;
      RECT 64.52 9.43 64.72 9.63 ;
      RECT 64.255 4.895 64.455 5.095 ;
      RECT 62.295 4.895 62.495 5.095 ;
      RECT 61.095 4.335 61.295 4.535 ;
      RECT 59.855 3.775 60.055 3.975 ;
      RECT 58.415 4.335 58.615 4.535 ;
      RECT 56.455 3.775 56.655 3.975 ;
      RECT 55.975 4.895 56.175 5.095 ;
      RECT 54.365 7.29 54.565 7.49 ;
      RECT 47.655 3.215 47.855 3.415 ;
      RECT 46.695 4.895 46.895 5.095 ;
      RECT 45.96 9.43 46.16 9.63 ;
      RECT 45.695 4.895 45.895 5.095 ;
      RECT 43.735 4.895 43.935 5.095 ;
      RECT 42.535 4.335 42.735 4.535 ;
      RECT 41.295 3.775 41.495 3.975 ;
      RECT 39.855 4.335 40.055 4.535 ;
      RECT 37.895 3.775 38.095 3.975 ;
      RECT 37.415 4.895 37.615 5.095 ;
      RECT 35.805 7.29 36.005 7.49 ;
      RECT 29.095 3.215 29.295 3.415 ;
      RECT 28.135 4.895 28.335 5.095 ;
      RECT 27.4 9.43 27.6 9.63 ;
      RECT 27.135 4.895 27.335 5.095 ;
      RECT 25.175 4.895 25.375 5.095 ;
      RECT 23.975 4.335 24.175 4.535 ;
      RECT 22.735 3.775 22.935 3.975 ;
      RECT 21.295 4.335 21.495 4.535 ;
      RECT 19.335 3.775 19.535 3.975 ;
      RECT 18.855 4.895 19.055 5.095 ;
    LAYER met2 ;
      RECT 16.225 10.69 110.225 10.86 ;
      RECT 110.055 9.565 110.225 10.86 ;
      RECT 16.225 8.545 16.395 10.86 ;
      RECT 110.025 9.565 110.375 9.915 ;
      RECT 16.165 8.545 16.455 8.895 ;
      RECT 106.865 8.51 107.185 8.835 ;
      RECT 106.895 7.985 107.065 8.835 ;
      RECT 106.895 7.985 107.07 8.335 ;
      RECT 106.895 7.985 107.87 8.16 ;
      RECT 107.695 3.26 107.87 8.16 ;
      RECT 107.64 3.26 107.99 3.61 ;
      RECT 107.665 8.945 107.99 9.27 ;
      RECT 106.55 9.035 107.99 9.205 ;
      RECT 106.55 3.69 106.71 9.205 ;
      RECT 106.865 3.66 107.185 3.98 ;
      RECT 106.55 3.69 107.185 3.86 ;
      RECT 99.43 5.43 105.52 5.62 ;
      RECT 105.35 4.44 105.52 5.62 ;
      RECT 105.33 4.445 105.52 5.62 ;
      RECT 99.43 4.81 99.6 5.62 ;
      RECT 99.375 4.81 99.655 5.18 ;
      RECT 99.445 4.365 99.585 5.62 ;
      RECT 105.26 4.445 105.6 4.795 ;
      RECT 99.255 4.25 99.535 4.62 ;
      RECT 98.965 4.365 99.585 4.505 ;
      RECT 98.965 3.155 99.105 4.505 ;
      RECT 98.905 3.155 99.165 3.475 ;
      RECT 91.44 8.945 91.79 9.295 ;
      RECT 102.225 8.9 102.575 9.25 ;
      RECT 91.44 8.975 102.575 9.175 ;
      RECT 101.865 4.275 102.125 4.595 ;
      RECT 101.925 3.155 102.065 4.595 ;
      RECT 101.865 3.155 102.125 3.475 ;
      RECT 100.865 4.835 101.125 5.155 ;
      RECT 100.865 4.25 101.065 5.155 ;
      RECT 100.805 3.155 100.945 4.785 ;
      RECT 100.805 4.25 101.305 4.62 ;
      RECT 100.745 3.155 101.005 3.475 ;
      RECT 100.385 4.835 100.645 5.155 ;
      RECT 100.445 3.245 100.585 5.155 ;
      RECT 100.145 3.245 100.585 3.475 ;
      RECT 100.145 3.155 100.405 3.475 ;
      RECT 99.905 3.715 100.165 4.035 ;
      RECT 99.325 3.805 100.165 3.945 ;
      RECT 99.325 2.865 99.465 3.945 ;
      RECT 95.985 3.155 96.245 3.475 ;
      RECT 95.985 3.245 97.025 3.385 ;
      RECT 96.885 2.865 97.025 3.385 ;
      RECT 96.885 2.865 99.465 3.005 ;
      RECT 98.175 4.25 98.455 4.62 ;
      RECT 98.245 3.155 98.385 4.62 ;
      RECT 98.185 3.155 98.445 3.475 ;
      RECT 97.825 4.835 98.085 5.155 ;
      RECT 97.885 3.245 98.025 5.155 ;
      RECT 97.465 3.155 97.725 3.475 ;
      RECT 97.465 3.245 98.025 3.385 ;
      RECT 95.495 4.25 95.775 4.62 ;
      RECT 97.465 4.275 97.725 4.595 ;
      RECT 95.145 4.275 95.775 4.595 ;
      RECT 95.145 4.365 97.725 4.505 ;
      RECT 96.935 3.69 97.215 4.06 ;
      RECT 96.935 3.715 97.465 4.035 ;
      RECT 94.025 4.275 94.285 4.595 ;
      RECT 94.085 3.155 94.225 4.595 ;
      RECT 94.025 3.155 94.285 3.475 ;
      RECT 93.055 4.81 93.335 5.18 ;
      RECT 93.065 4.555 93.325 5.18 ;
      RECT 88.305 8.51 88.625 8.835 ;
      RECT 88.335 7.985 88.505 8.835 ;
      RECT 88.335 7.985 88.51 8.335 ;
      RECT 88.335 7.985 89.31 8.16 ;
      RECT 89.135 3.26 89.31 8.16 ;
      RECT 89.08 3.26 89.43 3.61 ;
      RECT 89.105 8.945 89.43 9.27 ;
      RECT 87.99 9.035 89.43 9.205 ;
      RECT 87.99 3.69 88.15 9.205 ;
      RECT 88.305 3.66 88.625 3.98 ;
      RECT 87.99 3.69 88.625 3.86 ;
      RECT 80.87 5.43 86.96 5.62 ;
      RECT 86.79 4.44 86.96 5.62 ;
      RECT 86.77 4.445 86.96 5.62 ;
      RECT 80.87 4.81 81.04 5.62 ;
      RECT 80.815 4.81 81.095 5.18 ;
      RECT 80.885 4.365 81.025 5.62 ;
      RECT 86.7 4.445 87.04 4.795 ;
      RECT 80.695 4.25 80.975 4.62 ;
      RECT 80.405 4.365 81.025 4.505 ;
      RECT 80.405 3.155 80.545 4.505 ;
      RECT 80.345 3.155 80.605 3.475 ;
      RECT 72.88 8.945 73.23 9.295 ;
      RECT 83.665 8.9 84.015 9.25 ;
      RECT 72.88 8.975 84.015 9.175 ;
      RECT 83.305 4.275 83.565 4.595 ;
      RECT 83.365 3.155 83.505 4.595 ;
      RECT 83.305 3.155 83.565 3.475 ;
      RECT 82.305 4.835 82.565 5.155 ;
      RECT 82.305 4.25 82.505 5.155 ;
      RECT 82.245 3.155 82.385 4.785 ;
      RECT 82.245 4.25 82.745 4.62 ;
      RECT 82.185 3.155 82.445 3.475 ;
      RECT 81.825 4.835 82.085 5.155 ;
      RECT 81.885 3.245 82.025 5.155 ;
      RECT 81.585 3.245 82.025 3.475 ;
      RECT 81.585 3.155 81.845 3.475 ;
      RECT 81.345 3.715 81.605 4.035 ;
      RECT 80.765 3.805 81.605 3.945 ;
      RECT 80.765 2.865 80.905 3.945 ;
      RECT 77.425 3.155 77.685 3.475 ;
      RECT 77.425 3.245 78.465 3.385 ;
      RECT 78.325 2.865 78.465 3.385 ;
      RECT 78.325 2.865 80.905 3.005 ;
      RECT 79.615 4.25 79.895 4.62 ;
      RECT 79.685 3.155 79.825 4.62 ;
      RECT 79.625 3.155 79.885 3.475 ;
      RECT 79.265 4.835 79.525 5.155 ;
      RECT 79.325 3.245 79.465 5.155 ;
      RECT 78.905 3.155 79.165 3.475 ;
      RECT 78.905 3.245 79.465 3.385 ;
      RECT 76.935 4.25 77.215 4.62 ;
      RECT 78.905 4.275 79.165 4.595 ;
      RECT 76.585 4.275 77.215 4.595 ;
      RECT 76.585 4.365 79.165 4.505 ;
      RECT 78.375 3.69 78.655 4.06 ;
      RECT 78.375 3.715 78.905 4.035 ;
      RECT 75.465 4.275 75.725 4.595 ;
      RECT 75.525 3.155 75.665 4.595 ;
      RECT 75.465 3.155 75.725 3.475 ;
      RECT 74.495 4.81 74.775 5.18 ;
      RECT 74.505 4.555 74.765 5.18 ;
      RECT 69.745 8.51 70.065 8.835 ;
      RECT 69.775 7.985 69.945 8.835 ;
      RECT 69.775 7.985 69.95 8.335 ;
      RECT 69.775 7.985 70.75 8.16 ;
      RECT 70.575 3.26 70.75 8.16 ;
      RECT 70.52 3.26 70.87 3.61 ;
      RECT 70.545 8.945 70.87 9.27 ;
      RECT 69.43 9.035 70.87 9.205 ;
      RECT 69.43 3.69 69.59 9.205 ;
      RECT 69.745 3.66 70.065 3.98 ;
      RECT 69.43 3.69 70.065 3.86 ;
      RECT 62.31 5.43 68.4 5.62 ;
      RECT 68.23 4.44 68.4 5.62 ;
      RECT 68.21 4.445 68.4 5.62 ;
      RECT 62.31 4.81 62.48 5.62 ;
      RECT 62.255 4.81 62.535 5.18 ;
      RECT 62.325 4.365 62.465 5.62 ;
      RECT 68.14 4.445 68.48 4.795 ;
      RECT 62.135 4.25 62.415 4.62 ;
      RECT 61.845 4.365 62.465 4.505 ;
      RECT 61.845 3.155 61.985 4.505 ;
      RECT 61.785 3.155 62.045 3.475 ;
      RECT 54.365 8.95 54.715 9.3 ;
      RECT 65.105 8.905 65.455 9.255 ;
      RECT 54.365 8.98 65.455 9.18 ;
      RECT 64.745 4.275 65.005 4.595 ;
      RECT 64.805 3.155 64.945 4.595 ;
      RECT 64.745 3.155 65.005 3.475 ;
      RECT 63.745 4.835 64.005 5.155 ;
      RECT 63.745 4.25 63.945 5.155 ;
      RECT 63.685 3.155 63.825 4.785 ;
      RECT 63.685 4.25 64.185 4.62 ;
      RECT 63.625 3.155 63.885 3.475 ;
      RECT 63.265 4.835 63.525 5.155 ;
      RECT 63.325 3.245 63.465 5.155 ;
      RECT 63.025 3.245 63.465 3.475 ;
      RECT 63.025 3.155 63.285 3.475 ;
      RECT 62.785 3.715 63.045 4.035 ;
      RECT 62.205 3.805 63.045 3.945 ;
      RECT 62.205 2.865 62.345 3.945 ;
      RECT 58.865 3.155 59.125 3.475 ;
      RECT 58.865 3.245 59.905 3.385 ;
      RECT 59.765 2.865 59.905 3.385 ;
      RECT 59.765 2.865 62.345 3.005 ;
      RECT 61.055 4.25 61.335 4.62 ;
      RECT 61.125 3.155 61.265 4.62 ;
      RECT 61.065 3.155 61.325 3.475 ;
      RECT 60.705 4.835 60.965 5.155 ;
      RECT 60.765 3.245 60.905 5.155 ;
      RECT 60.345 3.155 60.605 3.475 ;
      RECT 60.345 3.245 60.905 3.385 ;
      RECT 58.375 4.25 58.655 4.62 ;
      RECT 60.345 4.275 60.605 4.595 ;
      RECT 58.025 4.275 58.655 4.595 ;
      RECT 58.025 4.365 60.605 4.505 ;
      RECT 59.815 3.69 60.095 4.06 ;
      RECT 59.815 3.715 60.345 4.035 ;
      RECT 56.905 4.275 57.165 4.595 ;
      RECT 56.965 3.155 57.105 4.595 ;
      RECT 56.905 3.155 57.165 3.475 ;
      RECT 55.935 4.81 56.215 5.18 ;
      RECT 55.945 4.555 56.205 5.18 ;
      RECT 51.185 8.51 51.505 8.835 ;
      RECT 51.215 7.985 51.385 8.835 ;
      RECT 51.215 7.985 51.39 8.335 ;
      RECT 51.215 7.985 52.19 8.16 ;
      RECT 52.015 3.26 52.19 8.16 ;
      RECT 51.96 3.26 52.31 3.61 ;
      RECT 51.985 8.945 52.31 9.27 ;
      RECT 50.87 9.035 52.31 9.205 ;
      RECT 50.87 3.69 51.03 9.205 ;
      RECT 51.185 3.66 51.505 3.98 ;
      RECT 50.87 3.69 51.505 3.86 ;
      RECT 43.75 5.43 49.84 5.62 ;
      RECT 49.67 4.44 49.84 5.62 ;
      RECT 49.65 4.445 49.84 5.62 ;
      RECT 43.75 4.81 43.92 5.62 ;
      RECT 43.695 4.81 43.975 5.18 ;
      RECT 43.765 4.365 43.905 5.62 ;
      RECT 49.58 4.445 49.92 4.795 ;
      RECT 43.575 4.25 43.855 4.62 ;
      RECT 43.285 4.365 43.905 4.505 ;
      RECT 43.285 3.155 43.425 4.505 ;
      RECT 43.225 3.155 43.485 3.475 ;
      RECT 35.805 8.945 36.155 9.295 ;
      RECT 46.55 8.9 46.9 9.25 ;
      RECT 35.805 8.975 46.9 9.175 ;
      RECT 46.185 4.275 46.445 4.595 ;
      RECT 46.245 3.155 46.385 4.595 ;
      RECT 46.185 3.155 46.445 3.475 ;
      RECT 45.185 4.835 45.445 5.155 ;
      RECT 45.185 4.25 45.385 5.155 ;
      RECT 45.125 3.155 45.265 4.785 ;
      RECT 45.125 4.25 45.625 4.62 ;
      RECT 45.065 3.155 45.325 3.475 ;
      RECT 44.705 4.835 44.965 5.155 ;
      RECT 44.765 3.245 44.905 5.155 ;
      RECT 44.465 3.245 44.905 3.475 ;
      RECT 44.465 3.155 44.725 3.475 ;
      RECT 44.225 3.715 44.485 4.035 ;
      RECT 43.645 3.805 44.485 3.945 ;
      RECT 43.645 2.865 43.785 3.945 ;
      RECT 40.305 3.155 40.565 3.475 ;
      RECT 40.305 3.245 41.345 3.385 ;
      RECT 41.205 2.865 41.345 3.385 ;
      RECT 41.205 2.865 43.785 3.005 ;
      RECT 42.495 4.25 42.775 4.62 ;
      RECT 42.565 3.155 42.705 4.62 ;
      RECT 42.505 3.155 42.765 3.475 ;
      RECT 42.145 4.835 42.405 5.155 ;
      RECT 42.205 3.245 42.345 5.155 ;
      RECT 41.785 3.155 42.045 3.475 ;
      RECT 41.785 3.245 42.345 3.385 ;
      RECT 39.815 4.25 40.095 4.62 ;
      RECT 41.785 4.275 42.045 4.595 ;
      RECT 39.465 4.275 40.095 4.595 ;
      RECT 39.465 4.365 42.045 4.505 ;
      RECT 41.255 3.69 41.535 4.06 ;
      RECT 41.255 3.715 41.785 4.035 ;
      RECT 38.345 4.275 38.605 4.595 ;
      RECT 38.405 3.155 38.545 4.595 ;
      RECT 38.345 3.155 38.605 3.475 ;
      RECT 37.375 4.81 37.655 5.18 ;
      RECT 37.385 4.555 37.645 5.18 ;
      RECT 32.625 8.51 32.945 8.835 ;
      RECT 32.655 7.985 32.825 8.835 ;
      RECT 32.655 7.985 32.83 8.335 ;
      RECT 32.655 7.985 33.63 8.16 ;
      RECT 33.455 3.26 33.63 8.16 ;
      RECT 33.4 3.26 33.75 3.61 ;
      RECT 33.425 8.945 33.75 9.27 ;
      RECT 32.31 9.035 33.75 9.205 ;
      RECT 32.31 3.69 32.47 9.205 ;
      RECT 32.625 3.66 32.945 3.98 ;
      RECT 32.31 3.69 32.945 3.86 ;
      RECT 25.19 5.43 31.28 5.62 ;
      RECT 31.11 4.44 31.28 5.62 ;
      RECT 31.09 4.445 31.28 5.62 ;
      RECT 25.19 4.81 25.36 5.62 ;
      RECT 25.135 4.81 25.415 5.18 ;
      RECT 25.205 4.365 25.345 5.62 ;
      RECT 31.02 4.445 31.36 4.795 ;
      RECT 25.015 4.25 25.295 4.62 ;
      RECT 24.725 4.365 25.345 4.505 ;
      RECT 24.725 3.155 24.865 4.505 ;
      RECT 24.665 3.155 24.925 3.475 ;
      RECT 16.54 9.285 16.83 9.635 ;
      RECT 16.54 9.345 17.73 9.515 ;
      RECT 17.56 8.975 17.73 9.515 ;
      RECT 27.99 8.895 28.34 9.245 ;
      RECT 17.56 8.975 28.34 9.145 ;
      RECT 27.625 4.275 27.885 4.595 ;
      RECT 27.685 3.155 27.825 4.595 ;
      RECT 27.625 3.155 27.885 3.475 ;
      RECT 26.625 4.835 26.885 5.155 ;
      RECT 26.625 4.25 26.825 5.155 ;
      RECT 26.565 3.155 26.705 4.785 ;
      RECT 26.565 4.25 27.065 4.62 ;
      RECT 26.505 3.155 26.765 3.475 ;
      RECT 26.145 4.835 26.405 5.155 ;
      RECT 26.205 3.245 26.345 5.155 ;
      RECT 25.905 3.245 26.345 3.475 ;
      RECT 25.905 3.155 26.165 3.475 ;
      RECT 25.665 3.715 25.925 4.035 ;
      RECT 25.085 3.805 25.925 3.945 ;
      RECT 25.085 2.865 25.225 3.945 ;
      RECT 21.745 3.155 22.005 3.475 ;
      RECT 21.745 3.245 22.785 3.385 ;
      RECT 22.645 2.865 22.785 3.385 ;
      RECT 22.645 2.865 25.225 3.005 ;
      RECT 23.935 4.25 24.215 4.62 ;
      RECT 24.005 3.155 24.145 4.62 ;
      RECT 23.945 3.155 24.205 3.475 ;
      RECT 23.585 4.835 23.845 5.155 ;
      RECT 23.645 3.245 23.785 5.155 ;
      RECT 23.225 3.155 23.485 3.475 ;
      RECT 23.225 3.245 23.785 3.385 ;
      RECT 21.255 4.25 21.535 4.62 ;
      RECT 23.225 4.275 23.485 4.595 ;
      RECT 20.905 4.275 21.535 4.595 ;
      RECT 20.905 4.365 23.485 4.505 ;
      RECT 22.695 3.69 22.975 4.06 ;
      RECT 22.695 3.715 23.225 4.035 ;
      RECT 19.785 4.275 20.045 4.595 ;
      RECT 19.845 3.155 19.985 4.595 ;
      RECT 19.785 3.155 20.045 3.475 ;
      RECT 18.815 4.81 19.095 5.18 ;
      RECT 18.825 4.555 19.085 5.18 ;
      RECT 109.955 7.2 110.335 7.58 ;
      RECT 103.295 3.13 103.575 3.5 ;
      RECT 102.335 4.81 102.615 5.18 ;
      RECT 101.555 9.345 101.93 9.715 ;
      RECT 101.335 4.81 101.615 5.18 ;
      RECT 93.535 3.69 93.815 4.06 ;
      RECT 91.395 7.2 91.775 7.58 ;
      RECT 84.735 3.13 85.015 3.5 ;
      RECT 83.775 4.81 84.055 5.18 ;
      RECT 82.995 9.345 83.37 9.715 ;
      RECT 82.775 4.81 83.055 5.18 ;
      RECT 74.975 3.69 75.255 4.06 ;
      RECT 72.835 7.2 73.215 7.58 ;
      RECT 66.175 3.13 66.455 3.5 ;
      RECT 65.215 4.81 65.495 5.18 ;
      RECT 64.435 9.345 64.81 9.715 ;
      RECT 64.215 4.81 64.495 5.18 ;
      RECT 56.415 3.69 56.695 4.06 ;
      RECT 54.275 7.2 54.655 7.58 ;
      RECT 47.615 3.13 47.895 3.5 ;
      RECT 46.655 4.81 46.935 5.18 ;
      RECT 45.875 9.345 46.25 9.715 ;
      RECT 45.655 4.81 45.935 5.18 ;
      RECT 37.855 3.69 38.135 4.06 ;
      RECT 35.715 7.2 36.095 7.58 ;
      RECT 29.055 3.13 29.335 3.5 ;
      RECT 28.095 4.81 28.375 5.18 ;
      RECT 27.315 9.345 27.69 9.715 ;
      RECT 27.095 4.81 27.375 5.18 ;
      RECT 19.295 3.69 19.575 4.06 ;
    LAYER via1 ;
      RECT 110.125 9.665 110.275 9.815 ;
      RECT 110.07 7.315 110.22 7.465 ;
      RECT 107.755 9.03 107.905 9.18 ;
      RECT 107.74 3.36 107.89 3.51 ;
      RECT 106.95 3.745 107.1 3.895 ;
      RECT 106.95 8.615 107.1 8.765 ;
      RECT 105.36 4.545 105.51 4.695 ;
      RECT 103.36 3.24 103.51 3.39 ;
      RECT 102.4 4.92 102.55 5.07 ;
      RECT 102.325 9 102.475 9.15 ;
      RECT 101.92 3.24 102.07 3.39 ;
      RECT 101.92 4.36 102.07 4.51 ;
      RECT 101.665 9.455 101.815 9.605 ;
      RECT 101.4 4.92 101.55 5.07 ;
      RECT 100.92 4.92 101.07 5.07 ;
      RECT 100.8 3.24 100.95 3.39 ;
      RECT 100.44 4.92 100.59 5.07 ;
      RECT 100.2 3.24 100.35 3.39 ;
      RECT 99.96 3.8 100.11 3.95 ;
      RECT 99.44 4.92 99.59 5.07 ;
      RECT 98.96 3.24 99.11 3.39 ;
      RECT 98.24 3.24 98.39 3.39 ;
      RECT 98.24 4.36 98.39 4.51 ;
      RECT 97.88 4.92 98.03 5.07 ;
      RECT 97.52 3.24 97.67 3.39 ;
      RECT 97.52 4.36 97.67 4.51 ;
      RECT 97.26 3.8 97.41 3.95 ;
      RECT 96.04 3.24 96.19 3.39 ;
      RECT 95.2 4.36 95.35 4.51 ;
      RECT 94.08 3.24 94.23 3.39 ;
      RECT 94.08 4.36 94.23 4.51 ;
      RECT 93.6 3.8 93.75 3.95 ;
      RECT 93.12 4.64 93.27 4.79 ;
      RECT 91.54 9.045 91.69 9.195 ;
      RECT 91.51 7.315 91.66 7.465 ;
      RECT 89.195 9.03 89.345 9.18 ;
      RECT 89.18 3.36 89.33 3.51 ;
      RECT 88.39 3.745 88.54 3.895 ;
      RECT 88.39 8.615 88.54 8.765 ;
      RECT 86.8 4.545 86.95 4.695 ;
      RECT 84.8 3.24 84.95 3.39 ;
      RECT 83.84 4.92 83.99 5.07 ;
      RECT 83.765 9 83.915 9.15 ;
      RECT 83.36 3.24 83.51 3.39 ;
      RECT 83.36 4.36 83.51 4.51 ;
      RECT 83.105 9.455 83.255 9.605 ;
      RECT 82.84 4.92 82.99 5.07 ;
      RECT 82.36 4.92 82.51 5.07 ;
      RECT 82.24 3.24 82.39 3.39 ;
      RECT 81.88 4.92 82.03 5.07 ;
      RECT 81.64 3.24 81.79 3.39 ;
      RECT 81.4 3.8 81.55 3.95 ;
      RECT 80.88 4.92 81.03 5.07 ;
      RECT 80.4 3.24 80.55 3.39 ;
      RECT 79.68 3.24 79.83 3.39 ;
      RECT 79.68 4.36 79.83 4.51 ;
      RECT 79.32 4.92 79.47 5.07 ;
      RECT 78.96 3.24 79.11 3.39 ;
      RECT 78.96 4.36 79.11 4.51 ;
      RECT 78.7 3.8 78.85 3.95 ;
      RECT 77.48 3.24 77.63 3.39 ;
      RECT 76.64 4.36 76.79 4.51 ;
      RECT 75.52 3.24 75.67 3.39 ;
      RECT 75.52 4.36 75.67 4.51 ;
      RECT 75.04 3.8 75.19 3.95 ;
      RECT 74.56 4.64 74.71 4.79 ;
      RECT 72.98 9.045 73.13 9.195 ;
      RECT 72.95 7.315 73.1 7.465 ;
      RECT 70.635 9.03 70.785 9.18 ;
      RECT 70.62 3.36 70.77 3.51 ;
      RECT 69.83 3.745 69.98 3.895 ;
      RECT 69.83 8.615 69.98 8.765 ;
      RECT 68.24 4.545 68.39 4.695 ;
      RECT 66.24 3.24 66.39 3.39 ;
      RECT 65.28 4.92 65.43 5.07 ;
      RECT 65.205 9.005 65.355 9.155 ;
      RECT 64.8 3.24 64.95 3.39 ;
      RECT 64.8 4.36 64.95 4.51 ;
      RECT 64.545 9.455 64.695 9.605 ;
      RECT 64.28 4.92 64.43 5.07 ;
      RECT 63.8 4.92 63.95 5.07 ;
      RECT 63.68 3.24 63.83 3.39 ;
      RECT 63.32 4.92 63.47 5.07 ;
      RECT 63.08 3.24 63.23 3.39 ;
      RECT 62.84 3.8 62.99 3.95 ;
      RECT 62.32 4.92 62.47 5.07 ;
      RECT 61.84 3.24 61.99 3.39 ;
      RECT 61.12 3.24 61.27 3.39 ;
      RECT 61.12 4.36 61.27 4.51 ;
      RECT 60.76 4.92 60.91 5.07 ;
      RECT 60.4 3.24 60.55 3.39 ;
      RECT 60.4 4.36 60.55 4.51 ;
      RECT 60.14 3.8 60.29 3.95 ;
      RECT 58.92 3.24 59.07 3.39 ;
      RECT 58.08 4.36 58.23 4.51 ;
      RECT 56.96 3.24 57.11 3.39 ;
      RECT 56.96 4.36 57.11 4.51 ;
      RECT 56.48 3.8 56.63 3.95 ;
      RECT 56 4.64 56.15 4.79 ;
      RECT 54.465 9.05 54.615 9.2 ;
      RECT 54.39 7.315 54.54 7.465 ;
      RECT 52.075 9.03 52.225 9.18 ;
      RECT 52.06 3.36 52.21 3.51 ;
      RECT 51.27 3.745 51.42 3.895 ;
      RECT 51.27 8.615 51.42 8.765 ;
      RECT 49.68 4.545 49.83 4.695 ;
      RECT 47.68 3.24 47.83 3.39 ;
      RECT 46.72 4.92 46.87 5.07 ;
      RECT 46.65 9 46.8 9.15 ;
      RECT 46.24 3.24 46.39 3.39 ;
      RECT 46.24 4.36 46.39 4.51 ;
      RECT 45.985 9.455 46.135 9.605 ;
      RECT 45.72 4.92 45.87 5.07 ;
      RECT 45.24 4.92 45.39 5.07 ;
      RECT 45.12 3.24 45.27 3.39 ;
      RECT 44.76 4.92 44.91 5.07 ;
      RECT 44.52 3.24 44.67 3.39 ;
      RECT 44.28 3.8 44.43 3.95 ;
      RECT 43.76 4.92 43.91 5.07 ;
      RECT 43.28 3.24 43.43 3.39 ;
      RECT 42.56 3.24 42.71 3.39 ;
      RECT 42.56 4.36 42.71 4.51 ;
      RECT 42.2 4.92 42.35 5.07 ;
      RECT 41.84 3.24 41.99 3.39 ;
      RECT 41.84 4.36 41.99 4.51 ;
      RECT 41.58 3.8 41.73 3.95 ;
      RECT 40.36 3.24 40.51 3.39 ;
      RECT 39.52 4.36 39.67 4.51 ;
      RECT 38.4 3.24 38.55 3.39 ;
      RECT 38.4 4.36 38.55 4.51 ;
      RECT 37.92 3.8 38.07 3.95 ;
      RECT 37.44 4.64 37.59 4.79 ;
      RECT 35.905 9.045 36.055 9.195 ;
      RECT 35.83 7.315 35.98 7.465 ;
      RECT 33.515 9.03 33.665 9.18 ;
      RECT 33.5 3.36 33.65 3.51 ;
      RECT 32.71 3.745 32.86 3.895 ;
      RECT 32.71 8.615 32.86 8.765 ;
      RECT 31.12 4.545 31.27 4.695 ;
      RECT 29.12 3.24 29.27 3.39 ;
      RECT 28.16 4.92 28.31 5.07 ;
      RECT 28.09 8.995 28.24 9.145 ;
      RECT 27.68 3.24 27.83 3.39 ;
      RECT 27.68 4.36 27.83 4.51 ;
      RECT 27.425 9.455 27.575 9.605 ;
      RECT 27.16 4.92 27.31 5.07 ;
      RECT 26.68 4.92 26.83 5.07 ;
      RECT 26.56 3.24 26.71 3.39 ;
      RECT 26.2 4.92 26.35 5.07 ;
      RECT 25.96 3.24 26.11 3.39 ;
      RECT 25.72 3.8 25.87 3.95 ;
      RECT 25.2 4.92 25.35 5.07 ;
      RECT 24.72 3.24 24.87 3.39 ;
      RECT 24 3.24 24.15 3.39 ;
      RECT 24 4.36 24.15 4.51 ;
      RECT 23.64 4.92 23.79 5.07 ;
      RECT 23.28 3.24 23.43 3.39 ;
      RECT 23.28 4.36 23.43 4.51 ;
      RECT 23.02 3.8 23.17 3.95 ;
      RECT 21.8 3.24 21.95 3.39 ;
      RECT 20.96 4.36 21.11 4.51 ;
      RECT 19.84 3.24 19.99 3.39 ;
      RECT 19.84 4.36 19.99 4.51 ;
      RECT 19.36 3.8 19.51 3.95 ;
      RECT 18.88 4.64 19.03 4.79 ;
      RECT 16.61 9.385 16.76 9.535 ;
      RECT 16.235 8.645 16.385 8.795 ;
    LAYER met1 ;
      RECT 109.995 10.055 110.29 10.285 ;
      RECT 110.055 9.565 110.23 10.285 ;
      RECT 110.025 9.565 110.375 9.915 ;
      RECT 110.055 8.575 110.225 10.285 ;
      RECT 109.995 8.575 110.285 8.805 ;
      RECT 109 10.06 109.295 10.29 ;
      RECT 109.06 8.58 109.23 10.29 ;
      RECT 109 8.58 109.29 8.81 ;
      RECT 109 8.615 109.855 8.775 ;
      RECT 109.685 8.205 109.855 8.775 ;
      RECT 109 8.61 109.395 8.775 ;
      RECT 109.625 8.205 109.915 8.435 ;
      RECT 109.625 8.235 110.085 8.405 ;
      RECT 109.585 4.03 109.91 4.26 ;
      RECT 109.585 4.06 110.08 4.23 ;
      RECT 109.585 3.69 109.775 4.26 ;
      RECT 109 3.655 109.29 3.885 ;
      RECT 109 3.69 109.775 3.86 ;
      RECT 109.06 2.175 109.23 3.885 ;
      RECT 109 2.175 109.295 2.405 ;
      RECT 108.63 4.025 108.92 4.255 ;
      RECT 108.63 4.055 109.09 4.225 ;
      RECT 108.695 2.95 108.86 4.255 ;
      RECT 107.21 2.915 107.5 3.145 ;
      RECT 107.21 2.95 108.86 3.12 ;
      RECT 107.27 2.175 107.44 3.145 ;
      RECT 107.21 2.175 107.5 2.405 ;
      RECT 107.21 10.06 107.5 10.29 ;
      RECT 107.27 9.32 107.44 10.29 ;
      RECT 107.27 9.41 108.86 9.58 ;
      RECT 108.69 8.21 108.86 9.58 ;
      RECT 107.21 9.32 107.5 9.55 ;
      RECT 108.63 8.21 108.92 8.44 ;
      RECT 108.63 8.24 109.09 8.41 ;
      RECT 105.26 4.445 105.6 4.795 ;
      RECT 105.35 3.32 105.52 4.795 ;
      RECT 107.64 3.26 107.99 3.61 ;
      RECT 105.35 3.32 107.99 3.49 ;
      RECT 107.47 3.315 107.99 3.49 ;
      RECT 107.665 8.945 107.99 9.27 ;
      RECT 102.225 8.9 102.575 9.25 ;
      RECT 107.64 8.95 107.99 9.18 ;
      RECT 102.025 8.95 102.575 9.18 ;
      RECT 107.47 8.975 107.99 9.15 ;
      RECT 101.855 8.975 102.575 9.15 ;
      RECT 101.855 8.975 107.99 9.145 ;
      RECT 106.865 3.66 107.185 3.98 ;
      RECT 106.84 3.655 107.13 3.885 ;
      RECT 106.835 3.685 107.185 3.86 ;
      RECT 106.665 3.685 107.185 3.855 ;
      RECT 106.865 8.545 107.185 8.835 ;
      RECT 106.84 8.58 107.185 8.81 ;
      RECT 106.665 8.61 107.185 8.78 ;
      RECT 102.315 4.865 102.635 5.125 ;
      RECT 103.605 4.04 103.745 4.9 ;
      RECT 102.405 4.76 103.745 4.9 ;
      RECT 102.405 4.32 102.545 5.125 ;
      RECT 102.33 4.32 102.62 4.55 ;
      RECT 103.53 4.04 103.82 4.27 ;
      RECT 103.05 4.32 103.34 4.55 ;
      RECT 103.245 3.245 103.385 4.505 ;
      RECT 103.275 3.185 103.595 3.445 ;
      RECT 99.875 3.745 100.195 4.005 ;
      RECT 102.57 3.76 102.86 3.99 ;
      RECT 99.965 3.665 102.785 3.805 ;
      RECT 101.835 3.185 102.155 3.445 ;
      RECT 102.33 3.2 102.62 3.43 ;
      RECT 101.835 3.245 102.62 3.385 ;
      RECT 101.835 4.305 102.155 4.565 ;
      RECT 101.835 4.085 102.065 4.565 ;
      RECT 101.33 4.04 101.62 4.27 ;
      RECT 101.33 4.085 102.065 4.225 ;
      RECT 101.595 10.06 101.885 10.29 ;
      RECT 101.655 9.32 101.825 10.29 ;
      RECT 101.555 9.345 101.935 9.715 ;
      RECT 101.595 9.32 101.885 9.715 ;
      RECT 100.355 4.865 100.675 5.125 ;
      RECT 99.89 4.88 100.18 5.11 ;
      RECT 99.89 4.925 100.675 5.065 ;
      RECT 98.65 3.76 98.94 3.99 ;
      RECT 98.65 3.805 99.585 3.945 ;
      RECT 99.445 3.245 99.585 3.945 ;
      RECT 100.115 3.185 100.435 3.445 ;
      RECT 99.89 3.2 100.435 3.43 ;
      RECT 99.445 3.245 100.435 3.385 ;
      RECT 97.795 4.865 98.115 5.125 ;
      RECT 97.795 4.925 98.865 5.065 ;
      RECT 98.725 4.365 98.865 5.065 ;
      RECT 99.89 4.32 100.18 4.55 ;
      RECT 98.725 4.365 100.18 4.505 ;
      RECT 98.155 3.185 98.475 3.445 ;
      RECT 97.93 3.2 98.475 3.43 ;
      RECT 97.175 3.745 97.495 4.005 ;
      RECT 98.17 3.76 98.46 3.99 ;
      RECT 96.93 3.76 97.495 3.99 ;
      RECT 96.93 3.805 98.46 3.945 ;
      RECT 96.45 4.32 96.74 4.55 ;
      RECT 96.645 3.245 96.785 4.505 ;
      RECT 97.435 3.185 97.755 3.445 ;
      RECT 96.45 3.2 96.74 3.43 ;
      RECT 96.45 3.245 97.755 3.385 ;
      RECT 96.045 4.76 97.145 4.9 ;
      RECT 96.93 4.6 97.22 4.83 ;
      RECT 95.97 4.6 96.26 4.83 ;
      RECT 95.955 3.185 96.275 3.445 ;
      RECT 93.995 3.185 94.315 3.445 ;
      RECT 93.995 3.245 96.275 3.385 ;
      RECT 95.115 4.305 95.435 4.565 ;
      RECT 95.115 4.305 95.945 4.445 ;
      RECT 95.73 4.04 95.945 4.445 ;
      RECT 95.73 4.04 96.02 4.27 ;
      RECT 93.515 3.745 93.835 4.005 ;
      RECT 94.925 3.76 95.215 3.99 ;
      RECT 93.515 3.76 94.06 3.99 ;
      RECT 93.515 3.845 94.465 3.985 ;
      RECT 94.325 3.665 94.465 3.985 ;
      RECT 94.825 3.76 95.215 3.945 ;
      RECT 94.325 3.665 94.965 3.805 ;
      RECT 93.035 4.555 93.355 4.97 ;
      RECT 93.115 3.2 93.27 4.97 ;
      RECT 93.05 3.2 93.34 3.43 ;
      RECT 91.435 10.055 91.73 10.285 ;
      RECT 91.495 8.575 91.665 10.285 ;
      RECT 91.44 8.945 91.79 9.295 ;
      RECT 91.435 8.575 91.725 8.805 ;
      RECT 90.44 10.06 90.735 10.29 ;
      RECT 90.5 8.58 90.67 10.29 ;
      RECT 90.44 8.58 90.73 8.81 ;
      RECT 90.44 8.615 91.295 8.775 ;
      RECT 91.125 8.205 91.295 8.775 ;
      RECT 90.44 8.61 90.835 8.775 ;
      RECT 91.065 8.205 91.355 8.435 ;
      RECT 91.065 8.235 91.525 8.405 ;
      RECT 91.025 4.03 91.35 4.26 ;
      RECT 91.025 4.06 91.52 4.23 ;
      RECT 91.025 3.69 91.215 4.26 ;
      RECT 90.44 3.655 90.73 3.885 ;
      RECT 90.44 3.69 91.215 3.86 ;
      RECT 90.5 2.175 90.67 3.885 ;
      RECT 90.44 2.175 90.735 2.405 ;
      RECT 90.07 4.025 90.36 4.255 ;
      RECT 90.07 4.055 90.53 4.225 ;
      RECT 90.135 2.95 90.3 4.255 ;
      RECT 88.65 2.915 88.94 3.145 ;
      RECT 88.65 2.95 90.3 3.12 ;
      RECT 88.71 2.175 88.88 3.145 ;
      RECT 88.65 2.175 88.94 2.405 ;
      RECT 88.65 10.06 88.94 10.29 ;
      RECT 88.71 9.32 88.88 10.29 ;
      RECT 88.71 9.41 90.3 9.58 ;
      RECT 90.13 8.21 90.3 9.58 ;
      RECT 88.65 9.32 88.94 9.55 ;
      RECT 90.07 8.21 90.36 8.44 ;
      RECT 90.07 8.24 90.53 8.41 ;
      RECT 86.7 4.445 87.04 4.795 ;
      RECT 86.79 3.32 86.96 4.795 ;
      RECT 89.08 3.26 89.43 3.61 ;
      RECT 86.79 3.32 89.43 3.49 ;
      RECT 88.91 3.315 89.43 3.49 ;
      RECT 89.105 8.945 89.43 9.27 ;
      RECT 83.665 8.9 84.015 9.25 ;
      RECT 89.08 8.95 89.43 9.18 ;
      RECT 83.465 8.95 84.015 9.18 ;
      RECT 88.91 8.975 89.43 9.15 ;
      RECT 83.295 8.975 84.015 9.15 ;
      RECT 83.295 8.975 89.43 9.145 ;
      RECT 88.305 3.66 88.625 3.98 ;
      RECT 88.28 3.655 88.57 3.885 ;
      RECT 88.275 3.685 88.625 3.86 ;
      RECT 88.105 3.685 88.625 3.855 ;
      RECT 88.305 8.545 88.625 8.835 ;
      RECT 88.28 8.58 88.625 8.81 ;
      RECT 88.105 8.61 88.625 8.78 ;
      RECT 83.755 4.865 84.075 5.125 ;
      RECT 85.045 4.04 85.185 4.9 ;
      RECT 83.845 4.76 85.185 4.9 ;
      RECT 83.845 4.32 83.985 5.125 ;
      RECT 83.77 4.32 84.06 4.55 ;
      RECT 84.97 4.04 85.26 4.27 ;
      RECT 84.49 4.32 84.78 4.55 ;
      RECT 84.685 3.245 84.825 4.505 ;
      RECT 84.715 3.185 85.035 3.445 ;
      RECT 81.315 3.745 81.635 4.005 ;
      RECT 84.01 3.76 84.3 3.99 ;
      RECT 81.405 3.665 84.225 3.805 ;
      RECT 83.275 3.185 83.595 3.445 ;
      RECT 83.77 3.2 84.06 3.43 ;
      RECT 83.275 3.245 84.06 3.385 ;
      RECT 83.275 4.305 83.595 4.565 ;
      RECT 83.275 4.085 83.505 4.565 ;
      RECT 82.77 4.04 83.06 4.27 ;
      RECT 82.77 4.085 83.505 4.225 ;
      RECT 83.035 10.06 83.325 10.29 ;
      RECT 83.095 9.32 83.265 10.29 ;
      RECT 82.995 9.345 83.375 9.715 ;
      RECT 83.035 9.32 83.325 9.715 ;
      RECT 81.795 4.865 82.115 5.125 ;
      RECT 81.33 4.88 81.62 5.11 ;
      RECT 81.33 4.925 82.115 5.065 ;
      RECT 80.09 3.76 80.38 3.99 ;
      RECT 80.09 3.805 81.025 3.945 ;
      RECT 80.885 3.245 81.025 3.945 ;
      RECT 81.555 3.185 81.875 3.445 ;
      RECT 81.33 3.2 81.875 3.43 ;
      RECT 80.885 3.245 81.875 3.385 ;
      RECT 79.235 4.865 79.555 5.125 ;
      RECT 79.235 4.925 80.305 5.065 ;
      RECT 80.165 4.365 80.305 5.065 ;
      RECT 81.33 4.32 81.62 4.55 ;
      RECT 80.165 4.365 81.62 4.505 ;
      RECT 79.595 3.185 79.915 3.445 ;
      RECT 79.37 3.2 79.915 3.43 ;
      RECT 78.615 3.745 78.935 4.005 ;
      RECT 79.61 3.76 79.9 3.99 ;
      RECT 78.37 3.76 78.935 3.99 ;
      RECT 78.37 3.805 79.9 3.945 ;
      RECT 77.89 4.32 78.18 4.55 ;
      RECT 78.085 3.245 78.225 4.505 ;
      RECT 78.875 3.185 79.195 3.445 ;
      RECT 77.89 3.2 78.18 3.43 ;
      RECT 77.89 3.245 79.195 3.385 ;
      RECT 77.485 4.76 78.585 4.9 ;
      RECT 78.37 4.6 78.66 4.83 ;
      RECT 77.41 4.6 77.7 4.83 ;
      RECT 77.395 3.185 77.715 3.445 ;
      RECT 75.435 3.185 75.755 3.445 ;
      RECT 75.435 3.245 77.715 3.385 ;
      RECT 76.555 4.305 76.875 4.565 ;
      RECT 76.555 4.305 77.385 4.445 ;
      RECT 77.17 4.04 77.385 4.445 ;
      RECT 77.17 4.04 77.46 4.27 ;
      RECT 74.955 3.745 75.275 4.005 ;
      RECT 76.365 3.76 76.655 3.99 ;
      RECT 74.955 3.76 75.5 3.99 ;
      RECT 74.955 3.845 75.905 3.985 ;
      RECT 75.765 3.665 75.905 3.985 ;
      RECT 76.265 3.76 76.655 3.945 ;
      RECT 75.765 3.665 76.405 3.805 ;
      RECT 74.475 4.555 74.795 4.97 ;
      RECT 74.555 3.2 74.71 4.97 ;
      RECT 74.49 3.2 74.78 3.43 ;
      RECT 72.875 10.055 73.17 10.285 ;
      RECT 72.935 8.575 73.105 10.285 ;
      RECT 72.88 8.945 73.23 9.295 ;
      RECT 72.875 8.575 73.165 8.805 ;
      RECT 71.88 10.06 72.175 10.29 ;
      RECT 71.94 8.58 72.11 10.29 ;
      RECT 71.88 8.58 72.17 8.81 ;
      RECT 71.88 8.615 72.735 8.775 ;
      RECT 72.565 8.205 72.735 8.775 ;
      RECT 71.88 8.61 72.275 8.775 ;
      RECT 72.505 8.205 72.795 8.435 ;
      RECT 72.505 8.235 72.965 8.405 ;
      RECT 72.465 4.03 72.79 4.26 ;
      RECT 72.465 4.06 72.96 4.23 ;
      RECT 72.465 3.69 72.655 4.26 ;
      RECT 71.88 3.655 72.17 3.885 ;
      RECT 71.88 3.69 72.655 3.86 ;
      RECT 71.94 2.175 72.11 3.885 ;
      RECT 71.88 2.175 72.175 2.405 ;
      RECT 71.51 4.025 71.8 4.255 ;
      RECT 71.51 4.055 71.97 4.225 ;
      RECT 71.575 2.95 71.74 4.255 ;
      RECT 70.09 2.915 70.38 3.145 ;
      RECT 70.09 2.95 71.74 3.12 ;
      RECT 70.15 2.175 70.32 3.145 ;
      RECT 70.09 2.175 70.38 2.405 ;
      RECT 70.09 10.06 70.38 10.29 ;
      RECT 70.15 9.32 70.32 10.29 ;
      RECT 70.15 9.41 71.74 9.58 ;
      RECT 71.57 8.21 71.74 9.58 ;
      RECT 70.09 9.32 70.38 9.55 ;
      RECT 71.51 8.21 71.8 8.44 ;
      RECT 71.51 8.24 71.97 8.41 ;
      RECT 68.14 4.445 68.48 4.795 ;
      RECT 68.23 3.32 68.4 4.795 ;
      RECT 70.52 3.26 70.87 3.61 ;
      RECT 68.23 3.32 70.87 3.49 ;
      RECT 70.35 3.315 70.87 3.49 ;
      RECT 70.545 8.945 70.87 9.27 ;
      RECT 65.105 8.905 65.455 9.255 ;
      RECT 70.52 8.95 70.87 9.18 ;
      RECT 64.905 8.95 65.455 9.18 ;
      RECT 70.35 8.975 70.87 9.15 ;
      RECT 64.735 8.975 65.455 9.15 ;
      RECT 64.735 8.975 70.87 9.145 ;
      RECT 69.745 3.66 70.065 3.98 ;
      RECT 69.72 3.655 70.01 3.885 ;
      RECT 69.715 3.685 70.065 3.86 ;
      RECT 69.545 3.685 70.065 3.855 ;
      RECT 69.745 8.545 70.065 8.835 ;
      RECT 69.72 8.58 70.065 8.81 ;
      RECT 69.545 8.61 70.065 8.78 ;
      RECT 65.195 4.865 65.515 5.125 ;
      RECT 66.485 4.04 66.625 4.9 ;
      RECT 65.285 4.76 66.625 4.9 ;
      RECT 65.285 4.32 65.425 5.125 ;
      RECT 65.21 4.32 65.5 4.55 ;
      RECT 66.41 4.04 66.7 4.27 ;
      RECT 65.93 4.32 66.22 4.55 ;
      RECT 66.125 3.245 66.265 4.505 ;
      RECT 66.155 3.185 66.475 3.445 ;
      RECT 62.755 3.745 63.075 4.005 ;
      RECT 65.45 3.76 65.74 3.99 ;
      RECT 62.845 3.665 65.665 3.805 ;
      RECT 64.715 3.185 65.035 3.445 ;
      RECT 65.21 3.2 65.5 3.43 ;
      RECT 64.715 3.245 65.5 3.385 ;
      RECT 64.715 4.305 65.035 4.565 ;
      RECT 64.715 4.085 64.945 4.565 ;
      RECT 64.21 4.04 64.5 4.27 ;
      RECT 64.21 4.085 64.945 4.225 ;
      RECT 64.475 10.06 64.765 10.29 ;
      RECT 64.535 9.32 64.705 10.29 ;
      RECT 64.435 9.345 64.815 9.715 ;
      RECT 64.475 9.32 64.765 9.715 ;
      RECT 63.235 4.865 63.555 5.125 ;
      RECT 62.77 4.88 63.06 5.11 ;
      RECT 62.77 4.925 63.555 5.065 ;
      RECT 61.53 3.76 61.82 3.99 ;
      RECT 61.53 3.805 62.465 3.945 ;
      RECT 62.325 3.245 62.465 3.945 ;
      RECT 62.995 3.185 63.315 3.445 ;
      RECT 62.77 3.2 63.315 3.43 ;
      RECT 62.325 3.245 63.315 3.385 ;
      RECT 60.675 4.865 60.995 5.125 ;
      RECT 60.675 4.925 61.745 5.065 ;
      RECT 61.605 4.365 61.745 5.065 ;
      RECT 62.77 4.32 63.06 4.55 ;
      RECT 61.605 4.365 63.06 4.505 ;
      RECT 61.035 3.185 61.355 3.445 ;
      RECT 60.81 3.2 61.355 3.43 ;
      RECT 60.055 3.745 60.375 4.005 ;
      RECT 61.05 3.76 61.34 3.99 ;
      RECT 59.81 3.76 60.375 3.99 ;
      RECT 59.81 3.805 61.34 3.945 ;
      RECT 59.33 4.32 59.62 4.55 ;
      RECT 59.525 3.245 59.665 4.505 ;
      RECT 60.315 3.185 60.635 3.445 ;
      RECT 59.33 3.2 59.62 3.43 ;
      RECT 59.33 3.245 60.635 3.385 ;
      RECT 58.925 4.76 60.025 4.9 ;
      RECT 59.81 4.6 60.1 4.83 ;
      RECT 58.85 4.6 59.14 4.83 ;
      RECT 58.835 3.185 59.155 3.445 ;
      RECT 56.875 3.185 57.195 3.445 ;
      RECT 56.875 3.245 59.155 3.385 ;
      RECT 57.995 4.305 58.315 4.565 ;
      RECT 57.995 4.305 58.825 4.445 ;
      RECT 58.61 4.04 58.825 4.445 ;
      RECT 58.61 4.04 58.9 4.27 ;
      RECT 56.395 3.745 56.715 4.005 ;
      RECT 57.805 3.76 58.095 3.99 ;
      RECT 56.395 3.76 56.94 3.99 ;
      RECT 56.395 3.845 57.345 3.985 ;
      RECT 57.205 3.665 57.345 3.985 ;
      RECT 57.705 3.76 58.095 3.945 ;
      RECT 57.205 3.665 57.845 3.805 ;
      RECT 55.915 4.555 56.235 4.97 ;
      RECT 55.995 3.2 56.15 4.97 ;
      RECT 55.93 3.2 56.22 3.43 ;
      RECT 54.315 10.055 54.61 10.285 ;
      RECT 54.375 8.575 54.545 10.285 ;
      RECT 54.36 8.95 54.715 9.305 ;
      RECT 54.315 8.575 54.605 8.805 ;
      RECT 53.32 10.06 53.615 10.29 ;
      RECT 53.38 8.58 53.55 10.29 ;
      RECT 53.32 8.58 53.61 8.81 ;
      RECT 53.32 8.615 54.175 8.775 ;
      RECT 54.005 8.205 54.175 8.775 ;
      RECT 53.32 8.61 53.715 8.775 ;
      RECT 53.945 8.205 54.235 8.435 ;
      RECT 53.945 8.235 54.405 8.405 ;
      RECT 53.905 4.03 54.23 4.26 ;
      RECT 53.905 4.06 54.4 4.23 ;
      RECT 53.905 3.69 54.095 4.26 ;
      RECT 53.32 3.655 53.61 3.885 ;
      RECT 53.32 3.69 54.095 3.86 ;
      RECT 53.38 2.175 53.55 3.885 ;
      RECT 53.32 2.175 53.615 2.405 ;
      RECT 52.95 4.025 53.24 4.255 ;
      RECT 52.95 4.055 53.41 4.225 ;
      RECT 53.015 2.95 53.18 4.255 ;
      RECT 51.53 2.915 51.82 3.145 ;
      RECT 51.53 2.95 53.18 3.12 ;
      RECT 51.59 2.175 51.76 3.145 ;
      RECT 51.53 2.175 51.82 2.405 ;
      RECT 51.53 10.06 51.82 10.29 ;
      RECT 51.59 9.32 51.76 10.29 ;
      RECT 51.59 9.41 53.18 9.58 ;
      RECT 53.01 8.21 53.18 9.58 ;
      RECT 51.53 9.32 51.82 9.55 ;
      RECT 52.95 8.21 53.24 8.44 ;
      RECT 52.95 8.24 53.41 8.41 ;
      RECT 49.58 4.445 49.92 4.795 ;
      RECT 49.67 3.32 49.84 4.795 ;
      RECT 51.96 3.26 52.31 3.61 ;
      RECT 49.67 3.32 52.31 3.49 ;
      RECT 51.79 3.315 52.31 3.49 ;
      RECT 51.985 8.945 52.31 9.27 ;
      RECT 46.55 8.9 46.9 9.25 ;
      RECT 51.96 8.95 52.31 9.18 ;
      RECT 46.345 8.95 46.9 9.18 ;
      RECT 51.79 8.975 52.31 9.15 ;
      RECT 46.175 8.975 46.9 9.15 ;
      RECT 46.175 8.975 52.31 9.145 ;
      RECT 51.185 3.66 51.505 3.98 ;
      RECT 51.16 3.655 51.45 3.885 ;
      RECT 51.155 3.685 51.505 3.86 ;
      RECT 50.985 3.685 51.505 3.855 ;
      RECT 51.185 8.545 51.505 8.835 ;
      RECT 51.16 8.58 51.505 8.81 ;
      RECT 50.985 8.61 51.505 8.78 ;
      RECT 46.635 4.865 46.955 5.125 ;
      RECT 47.925 4.04 48.065 4.9 ;
      RECT 46.725 4.76 48.065 4.9 ;
      RECT 46.725 4.32 46.865 5.125 ;
      RECT 46.65 4.32 46.94 4.55 ;
      RECT 47.85 4.04 48.14 4.27 ;
      RECT 47.37 4.32 47.66 4.55 ;
      RECT 47.565 3.245 47.705 4.505 ;
      RECT 47.595 3.185 47.915 3.445 ;
      RECT 44.195 3.745 44.515 4.005 ;
      RECT 46.89 3.76 47.18 3.99 ;
      RECT 44.285 3.665 47.105 3.805 ;
      RECT 46.155 3.185 46.475 3.445 ;
      RECT 46.65 3.2 46.94 3.43 ;
      RECT 46.155 3.245 46.94 3.385 ;
      RECT 46.155 4.305 46.475 4.565 ;
      RECT 46.155 4.085 46.385 4.565 ;
      RECT 45.65 4.04 45.94 4.27 ;
      RECT 45.65 4.085 46.385 4.225 ;
      RECT 45.915 10.06 46.205 10.29 ;
      RECT 45.975 9.32 46.145 10.29 ;
      RECT 45.875 9.345 46.255 9.715 ;
      RECT 45.915 9.32 46.205 9.715 ;
      RECT 44.675 4.865 44.995 5.125 ;
      RECT 44.21 4.88 44.5 5.11 ;
      RECT 44.21 4.925 44.995 5.065 ;
      RECT 42.97 3.76 43.26 3.99 ;
      RECT 42.97 3.805 43.905 3.945 ;
      RECT 43.765 3.245 43.905 3.945 ;
      RECT 44.435 3.185 44.755 3.445 ;
      RECT 44.21 3.2 44.755 3.43 ;
      RECT 43.765 3.245 44.755 3.385 ;
      RECT 42.115 4.865 42.435 5.125 ;
      RECT 42.115 4.925 43.185 5.065 ;
      RECT 43.045 4.365 43.185 5.065 ;
      RECT 44.21 4.32 44.5 4.55 ;
      RECT 43.045 4.365 44.5 4.505 ;
      RECT 42.475 3.185 42.795 3.445 ;
      RECT 42.25 3.2 42.795 3.43 ;
      RECT 41.495 3.745 41.815 4.005 ;
      RECT 42.49 3.76 42.78 3.99 ;
      RECT 41.25 3.76 41.815 3.99 ;
      RECT 41.25 3.805 42.78 3.945 ;
      RECT 40.77 4.32 41.06 4.55 ;
      RECT 40.965 3.245 41.105 4.505 ;
      RECT 41.755 3.185 42.075 3.445 ;
      RECT 40.77 3.2 41.06 3.43 ;
      RECT 40.77 3.245 42.075 3.385 ;
      RECT 40.365 4.76 41.465 4.9 ;
      RECT 41.25 4.6 41.54 4.83 ;
      RECT 40.29 4.6 40.58 4.83 ;
      RECT 40.275 3.185 40.595 3.445 ;
      RECT 38.315 3.185 38.635 3.445 ;
      RECT 38.315 3.245 40.595 3.385 ;
      RECT 39.435 4.305 39.755 4.565 ;
      RECT 39.435 4.305 40.265 4.445 ;
      RECT 40.05 4.04 40.265 4.445 ;
      RECT 40.05 4.04 40.34 4.27 ;
      RECT 37.835 3.745 38.155 4.005 ;
      RECT 39.245 3.76 39.535 3.99 ;
      RECT 37.835 3.76 38.38 3.99 ;
      RECT 37.835 3.845 38.785 3.985 ;
      RECT 38.645 3.665 38.785 3.985 ;
      RECT 39.145 3.76 39.535 3.945 ;
      RECT 38.645 3.665 39.285 3.805 ;
      RECT 37.355 4.555 37.675 4.97 ;
      RECT 37.435 3.2 37.59 4.97 ;
      RECT 37.37 3.2 37.66 3.43 ;
      RECT 35.755 10.055 36.05 10.285 ;
      RECT 35.815 8.575 35.985 10.285 ;
      RECT 35.805 8.945 36.155 9.295 ;
      RECT 35.755 8.575 36.045 8.805 ;
      RECT 34.76 10.06 35.055 10.29 ;
      RECT 34.82 8.58 34.99 10.29 ;
      RECT 34.76 8.58 35.05 8.81 ;
      RECT 34.76 8.615 35.615 8.775 ;
      RECT 35.445 8.205 35.615 8.775 ;
      RECT 34.76 8.61 35.155 8.775 ;
      RECT 35.385 8.205 35.675 8.435 ;
      RECT 35.385 8.235 35.845 8.405 ;
      RECT 35.345 4.03 35.67 4.26 ;
      RECT 35.345 4.06 35.84 4.23 ;
      RECT 35.345 3.69 35.535 4.26 ;
      RECT 34.76 3.655 35.05 3.885 ;
      RECT 34.76 3.69 35.535 3.86 ;
      RECT 34.82 2.175 34.99 3.885 ;
      RECT 34.76 2.175 35.055 2.405 ;
      RECT 34.39 4.025 34.68 4.255 ;
      RECT 34.39 4.055 34.85 4.225 ;
      RECT 34.455 2.95 34.62 4.255 ;
      RECT 32.97 2.915 33.26 3.145 ;
      RECT 32.97 2.95 34.62 3.12 ;
      RECT 33.03 2.175 33.2 3.145 ;
      RECT 32.97 2.175 33.26 2.405 ;
      RECT 32.97 10.06 33.26 10.29 ;
      RECT 33.03 9.32 33.2 10.29 ;
      RECT 33.03 9.41 34.62 9.58 ;
      RECT 34.45 8.21 34.62 9.58 ;
      RECT 32.97 9.32 33.26 9.55 ;
      RECT 34.39 8.21 34.68 8.44 ;
      RECT 34.39 8.24 34.85 8.41 ;
      RECT 31.02 4.445 31.36 4.795 ;
      RECT 31.11 3.32 31.28 4.795 ;
      RECT 33.4 3.26 33.75 3.61 ;
      RECT 31.11 3.32 33.75 3.49 ;
      RECT 33.23 3.315 33.75 3.49 ;
      RECT 33.425 8.945 33.75 9.27 ;
      RECT 27.99 8.895 28.34 9.245 ;
      RECT 33.4 8.95 33.75 9.18 ;
      RECT 27.785 8.95 28.34 9.18 ;
      RECT 33.23 8.975 33.75 9.15 ;
      RECT 27.615 8.975 28.34 9.15 ;
      RECT 27.615 8.975 33.75 9.145 ;
      RECT 32.625 3.66 32.945 3.98 ;
      RECT 32.6 3.655 32.89 3.885 ;
      RECT 32.595 3.685 32.945 3.86 ;
      RECT 32.425 3.685 32.945 3.855 ;
      RECT 32.625 8.545 32.945 8.835 ;
      RECT 32.6 8.58 32.945 8.81 ;
      RECT 32.425 8.61 32.945 8.78 ;
      RECT 28.075 4.865 28.395 5.125 ;
      RECT 29.365 4.04 29.505 4.9 ;
      RECT 28.165 4.76 29.505 4.9 ;
      RECT 28.165 4.32 28.305 5.125 ;
      RECT 28.09 4.32 28.38 4.55 ;
      RECT 29.29 4.04 29.58 4.27 ;
      RECT 28.81 4.32 29.1 4.55 ;
      RECT 29.005 3.245 29.145 4.505 ;
      RECT 29.035 3.185 29.355 3.445 ;
      RECT 25.635 3.745 25.955 4.005 ;
      RECT 28.33 3.76 28.62 3.99 ;
      RECT 25.725 3.665 28.545 3.805 ;
      RECT 27.595 3.185 27.915 3.445 ;
      RECT 28.09 3.2 28.38 3.43 ;
      RECT 27.595 3.245 28.38 3.385 ;
      RECT 27.595 4.305 27.915 4.565 ;
      RECT 27.595 4.085 27.825 4.565 ;
      RECT 27.09 4.04 27.38 4.27 ;
      RECT 27.09 4.085 27.825 4.225 ;
      RECT 27.355 10.06 27.645 10.29 ;
      RECT 27.415 9.32 27.585 10.29 ;
      RECT 27.315 9.345 27.695 9.715 ;
      RECT 27.355 9.32 27.645 9.715 ;
      RECT 26.115 4.865 26.435 5.125 ;
      RECT 25.65 4.88 25.94 5.11 ;
      RECT 25.65 4.925 26.435 5.065 ;
      RECT 24.41 3.76 24.7 3.99 ;
      RECT 24.41 3.805 25.345 3.945 ;
      RECT 25.205 3.245 25.345 3.945 ;
      RECT 25.875 3.185 26.195 3.445 ;
      RECT 25.65 3.2 26.195 3.43 ;
      RECT 25.205 3.245 26.195 3.385 ;
      RECT 23.555 4.865 23.875 5.125 ;
      RECT 23.555 4.925 24.625 5.065 ;
      RECT 24.485 4.365 24.625 5.065 ;
      RECT 25.65 4.32 25.94 4.55 ;
      RECT 24.485 4.365 25.94 4.505 ;
      RECT 23.915 3.185 24.235 3.445 ;
      RECT 23.69 3.2 24.235 3.43 ;
      RECT 22.935 3.745 23.255 4.005 ;
      RECT 23.93 3.76 24.22 3.99 ;
      RECT 22.69 3.76 23.255 3.99 ;
      RECT 22.69 3.805 24.22 3.945 ;
      RECT 22.21 4.32 22.5 4.55 ;
      RECT 22.405 3.245 22.545 4.505 ;
      RECT 23.195 3.185 23.515 3.445 ;
      RECT 22.21 3.2 22.5 3.43 ;
      RECT 22.21 3.245 23.515 3.385 ;
      RECT 21.805 4.76 22.905 4.9 ;
      RECT 22.69 4.6 22.98 4.83 ;
      RECT 21.73 4.6 22.02 4.83 ;
      RECT 21.715 3.185 22.035 3.445 ;
      RECT 19.755 3.185 20.075 3.445 ;
      RECT 19.755 3.245 22.035 3.385 ;
      RECT 20.875 4.305 21.195 4.565 ;
      RECT 20.875 4.305 21.705 4.445 ;
      RECT 21.49 4.04 21.705 4.445 ;
      RECT 21.49 4.04 21.78 4.27 ;
      RECT 19.275 3.745 19.595 4.005 ;
      RECT 20.685 3.76 20.975 3.99 ;
      RECT 19.275 3.76 19.82 3.99 ;
      RECT 19.275 3.845 20.225 3.985 ;
      RECT 20.085 3.665 20.225 3.985 ;
      RECT 20.585 3.76 20.975 3.945 ;
      RECT 20.085 3.665 20.725 3.805 ;
      RECT 18.795 4.555 19.115 4.97 ;
      RECT 18.875 3.2 19.03 4.97 ;
      RECT 18.81 3.2 19.1 3.43 ;
      RECT 16.54 10.06 16.83 10.29 ;
      RECT 16.6 9.315 16.77 10.29 ;
      RECT 16.51 9.315 16.86 9.605 ;
      RECT 16.135 8.575 16.485 8.865 ;
      RECT 15.995 8.61 16.485 8.78 ;
      RECT 109.97 7.245 110.32 7.535 ;
      RECT 101.315 4.865 101.635 5.125 ;
      RECT 100.715 3.185 101.395 3.445 ;
      RECT 100.835 4.865 101.155 5.125 ;
      RECT 99.355 4.865 99.675 5.125 ;
      RECT 98.875 3.185 99.195 3.445 ;
      RECT 98.155 4.305 98.475 4.565 ;
      RECT 97.435 4.305 97.755 4.565 ;
      RECT 93.995 4.305 94.315 4.565 ;
      RECT 91.41 7.245 91.76 7.535 ;
      RECT 82.755 4.865 83.075 5.125 ;
      RECT 82.155 3.185 82.835 3.445 ;
      RECT 82.275 4.865 82.595 5.125 ;
      RECT 80.795 4.865 81.115 5.125 ;
      RECT 80.315 3.185 80.635 3.445 ;
      RECT 79.595 4.305 79.915 4.565 ;
      RECT 78.875 4.305 79.195 4.565 ;
      RECT 75.435 4.305 75.755 4.565 ;
      RECT 72.85 7.245 73.2 7.535 ;
      RECT 64.195 4.865 64.515 5.125 ;
      RECT 63.595 3.185 64.275 3.445 ;
      RECT 63.715 4.865 64.035 5.125 ;
      RECT 62.235 4.865 62.555 5.125 ;
      RECT 61.755 3.185 62.075 3.445 ;
      RECT 61.035 4.305 61.355 4.565 ;
      RECT 60.315 4.305 60.635 4.565 ;
      RECT 56.875 4.305 57.195 4.565 ;
      RECT 54.29 7.245 54.64 7.535 ;
      RECT 45.635 4.865 45.955 5.125 ;
      RECT 45.035 3.185 45.715 3.445 ;
      RECT 45.155 4.865 45.475 5.125 ;
      RECT 43.675 4.865 43.995 5.125 ;
      RECT 43.195 3.185 43.515 3.445 ;
      RECT 42.475 4.305 42.795 4.565 ;
      RECT 41.755 4.305 42.075 4.565 ;
      RECT 38.315 4.305 38.635 4.565 ;
      RECT 35.73 7.245 36.08 7.535 ;
      RECT 27.075 4.865 27.395 5.125 ;
      RECT 26.475 3.185 27.155 3.445 ;
      RECT 26.595 4.865 26.915 5.125 ;
      RECT 25.115 4.865 25.435 5.125 ;
      RECT 24.635 3.185 24.955 3.445 ;
      RECT 23.915 4.305 24.235 4.565 ;
      RECT 23.195 4.305 23.515 4.565 ;
      RECT 19.755 4.305 20.075 4.565 ;
    LAYER mcon ;
      RECT 110.06 7.305 110.23 7.475 ;
      RECT 110.055 8.605 110.225 8.775 ;
      RECT 110.055 10.085 110.225 10.255 ;
      RECT 109.685 8.235 109.855 8.405 ;
      RECT 109.68 4.06 109.85 4.23 ;
      RECT 109.06 2.205 109.23 2.375 ;
      RECT 109.06 3.685 109.23 3.855 ;
      RECT 109.06 8.61 109.23 8.78 ;
      RECT 109.06 10.09 109.23 10.26 ;
      RECT 108.69 4.055 108.86 4.225 ;
      RECT 108.69 8.24 108.86 8.41 ;
      RECT 107.7 3.315 107.87 3.485 ;
      RECT 107.7 8.98 107.87 9.15 ;
      RECT 107.27 2.205 107.44 2.375 ;
      RECT 107.27 2.945 107.44 3.115 ;
      RECT 107.27 9.35 107.44 9.52 ;
      RECT 107.27 10.09 107.44 10.26 ;
      RECT 106.9 3.685 107.07 3.855 ;
      RECT 106.9 8.61 107.07 8.78 ;
      RECT 103.59 4.07 103.76 4.24 ;
      RECT 103.35 3.23 103.52 3.4 ;
      RECT 103.11 4.35 103.28 4.52 ;
      RECT 102.63 3.79 102.8 3.96 ;
      RECT 102.39 3.23 102.56 3.4 ;
      RECT 102.39 4.35 102.56 4.52 ;
      RECT 102.39 4.91 102.56 5.08 ;
      RECT 102.085 8.98 102.255 9.15 ;
      RECT 101.91 4.35 102.08 4.52 ;
      RECT 101.655 9.35 101.825 9.52 ;
      RECT 101.655 10.09 101.825 10.26 ;
      RECT 101.39 4.07 101.56 4.24 ;
      RECT 101.39 4.91 101.56 5.08 ;
      RECT 100.91 3.23 101.08 3.4 ;
      RECT 100.91 4.91 101.08 5.08 ;
      RECT 99.95 3.23 100.12 3.4 ;
      RECT 99.95 3.79 100.12 3.96 ;
      RECT 99.95 4.35 100.12 4.52 ;
      RECT 99.95 4.91 100.12 5.08 ;
      RECT 99.43 4.91 99.6 5.08 ;
      RECT 98.95 3.23 99.12 3.4 ;
      RECT 98.71 3.79 98.88 3.96 ;
      RECT 98.23 3.79 98.4 3.96 ;
      RECT 98.23 4.35 98.4 4.52 ;
      RECT 97.99 3.23 98.16 3.4 ;
      RECT 97.51 4.35 97.68 4.52 ;
      RECT 96.99 3.79 97.16 3.96 ;
      RECT 96.99 4.63 97.16 4.8 ;
      RECT 96.51 3.23 96.68 3.4 ;
      RECT 96.51 4.35 96.68 4.52 ;
      RECT 96.03 4.63 96.2 4.8 ;
      RECT 95.79 4.07 95.96 4.24 ;
      RECT 94.985 3.79 95.155 3.96 ;
      RECT 94.07 3.23 94.24 3.4 ;
      RECT 94.07 4.35 94.24 4.52 ;
      RECT 93.83 3.79 94 3.96 ;
      RECT 93.11 3.23 93.28 3.4 ;
      RECT 93.11 4.77 93.28 4.94 ;
      RECT 91.5 7.305 91.67 7.475 ;
      RECT 91.495 8.605 91.665 8.775 ;
      RECT 91.495 10.085 91.665 10.255 ;
      RECT 91.125 8.235 91.295 8.405 ;
      RECT 91.12 4.06 91.29 4.23 ;
      RECT 90.5 2.205 90.67 2.375 ;
      RECT 90.5 3.685 90.67 3.855 ;
      RECT 90.5 8.61 90.67 8.78 ;
      RECT 90.5 10.09 90.67 10.26 ;
      RECT 90.13 4.055 90.3 4.225 ;
      RECT 90.13 8.24 90.3 8.41 ;
      RECT 89.14 3.315 89.31 3.485 ;
      RECT 89.14 8.98 89.31 9.15 ;
      RECT 88.71 2.205 88.88 2.375 ;
      RECT 88.71 2.945 88.88 3.115 ;
      RECT 88.71 9.35 88.88 9.52 ;
      RECT 88.71 10.09 88.88 10.26 ;
      RECT 88.34 3.685 88.51 3.855 ;
      RECT 88.34 8.61 88.51 8.78 ;
      RECT 85.03 4.07 85.2 4.24 ;
      RECT 84.79 3.23 84.96 3.4 ;
      RECT 84.55 4.35 84.72 4.52 ;
      RECT 84.07 3.79 84.24 3.96 ;
      RECT 83.83 3.23 84 3.4 ;
      RECT 83.83 4.35 84 4.52 ;
      RECT 83.83 4.91 84 5.08 ;
      RECT 83.525 8.98 83.695 9.15 ;
      RECT 83.35 4.35 83.52 4.52 ;
      RECT 83.095 9.35 83.265 9.52 ;
      RECT 83.095 10.09 83.265 10.26 ;
      RECT 82.83 4.07 83 4.24 ;
      RECT 82.83 4.91 83 5.08 ;
      RECT 82.35 3.23 82.52 3.4 ;
      RECT 82.35 4.91 82.52 5.08 ;
      RECT 81.39 3.23 81.56 3.4 ;
      RECT 81.39 3.79 81.56 3.96 ;
      RECT 81.39 4.35 81.56 4.52 ;
      RECT 81.39 4.91 81.56 5.08 ;
      RECT 80.87 4.91 81.04 5.08 ;
      RECT 80.39 3.23 80.56 3.4 ;
      RECT 80.15 3.79 80.32 3.96 ;
      RECT 79.67 3.79 79.84 3.96 ;
      RECT 79.67 4.35 79.84 4.52 ;
      RECT 79.43 3.23 79.6 3.4 ;
      RECT 78.95 4.35 79.12 4.52 ;
      RECT 78.43 3.79 78.6 3.96 ;
      RECT 78.43 4.63 78.6 4.8 ;
      RECT 77.95 3.23 78.12 3.4 ;
      RECT 77.95 4.35 78.12 4.52 ;
      RECT 77.47 4.63 77.64 4.8 ;
      RECT 77.23 4.07 77.4 4.24 ;
      RECT 76.425 3.79 76.595 3.96 ;
      RECT 75.51 3.23 75.68 3.4 ;
      RECT 75.51 4.35 75.68 4.52 ;
      RECT 75.27 3.79 75.44 3.96 ;
      RECT 74.55 3.23 74.72 3.4 ;
      RECT 74.55 4.77 74.72 4.94 ;
      RECT 72.94 7.305 73.11 7.475 ;
      RECT 72.935 8.605 73.105 8.775 ;
      RECT 72.935 10.085 73.105 10.255 ;
      RECT 72.565 8.235 72.735 8.405 ;
      RECT 72.56 4.06 72.73 4.23 ;
      RECT 71.94 2.205 72.11 2.375 ;
      RECT 71.94 3.685 72.11 3.855 ;
      RECT 71.94 8.61 72.11 8.78 ;
      RECT 71.94 10.09 72.11 10.26 ;
      RECT 71.57 4.055 71.74 4.225 ;
      RECT 71.57 8.24 71.74 8.41 ;
      RECT 70.58 3.315 70.75 3.485 ;
      RECT 70.58 8.98 70.75 9.15 ;
      RECT 70.15 2.205 70.32 2.375 ;
      RECT 70.15 2.945 70.32 3.115 ;
      RECT 70.15 9.35 70.32 9.52 ;
      RECT 70.15 10.09 70.32 10.26 ;
      RECT 69.78 3.685 69.95 3.855 ;
      RECT 69.78 8.61 69.95 8.78 ;
      RECT 66.47 4.07 66.64 4.24 ;
      RECT 66.23 3.23 66.4 3.4 ;
      RECT 65.99 4.35 66.16 4.52 ;
      RECT 65.51 3.79 65.68 3.96 ;
      RECT 65.27 3.23 65.44 3.4 ;
      RECT 65.27 4.35 65.44 4.52 ;
      RECT 65.27 4.91 65.44 5.08 ;
      RECT 64.965 8.98 65.135 9.15 ;
      RECT 64.79 4.35 64.96 4.52 ;
      RECT 64.535 9.35 64.705 9.52 ;
      RECT 64.535 10.09 64.705 10.26 ;
      RECT 64.27 4.07 64.44 4.24 ;
      RECT 64.27 4.91 64.44 5.08 ;
      RECT 63.79 3.23 63.96 3.4 ;
      RECT 63.79 4.91 63.96 5.08 ;
      RECT 62.83 3.23 63 3.4 ;
      RECT 62.83 3.79 63 3.96 ;
      RECT 62.83 4.35 63 4.52 ;
      RECT 62.83 4.91 63 5.08 ;
      RECT 62.31 4.91 62.48 5.08 ;
      RECT 61.83 3.23 62 3.4 ;
      RECT 61.59 3.79 61.76 3.96 ;
      RECT 61.11 3.79 61.28 3.96 ;
      RECT 61.11 4.35 61.28 4.52 ;
      RECT 60.87 3.23 61.04 3.4 ;
      RECT 60.39 4.35 60.56 4.52 ;
      RECT 59.87 3.79 60.04 3.96 ;
      RECT 59.87 4.63 60.04 4.8 ;
      RECT 59.39 3.23 59.56 3.4 ;
      RECT 59.39 4.35 59.56 4.52 ;
      RECT 58.91 4.63 59.08 4.8 ;
      RECT 58.67 4.07 58.84 4.24 ;
      RECT 57.865 3.79 58.035 3.96 ;
      RECT 56.95 3.23 57.12 3.4 ;
      RECT 56.95 4.35 57.12 4.52 ;
      RECT 56.71 3.79 56.88 3.96 ;
      RECT 55.99 3.23 56.16 3.4 ;
      RECT 55.99 4.77 56.16 4.94 ;
      RECT 54.38 7.305 54.55 7.475 ;
      RECT 54.375 8.605 54.545 8.775 ;
      RECT 54.375 10.085 54.545 10.255 ;
      RECT 54.005 8.235 54.175 8.405 ;
      RECT 54 4.06 54.17 4.23 ;
      RECT 53.38 2.205 53.55 2.375 ;
      RECT 53.38 3.685 53.55 3.855 ;
      RECT 53.38 8.61 53.55 8.78 ;
      RECT 53.38 10.09 53.55 10.26 ;
      RECT 53.01 4.055 53.18 4.225 ;
      RECT 53.01 8.24 53.18 8.41 ;
      RECT 52.02 3.315 52.19 3.485 ;
      RECT 52.02 8.98 52.19 9.15 ;
      RECT 51.59 2.205 51.76 2.375 ;
      RECT 51.59 2.945 51.76 3.115 ;
      RECT 51.59 9.35 51.76 9.52 ;
      RECT 51.59 10.09 51.76 10.26 ;
      RECT 51.22 3.685 51.39 3.855 ;
      RECT 51.22 8.61 51.39 8.78 ;
      RECT 47.91 4.07 48.08 4.24 ;
      RECT 47.67 3.23 47.84 3.4 ;
      RECT 47.43 4.35 47.6 4.52 ;
      RECT 46.95 3.79 47.12 3.96 ;
      RECT 46.71 3.23 46.88 3.4 ;
      RECT 46.71 4.35 46.88 4.52 ;
      RECT 46.71 4.91 46.88 5.08 ;
      RECT 46.405 8.98 46.575 9.15 ;
      RECT 46.23 4.35 46.4 4.52 ;
      RECT 45.975 9.35 46.145 9.52 ;
      RECT 45.975 10.09 46.145 10.26 ;
      RECT 45.71 4.07 45.88 4.24 ;
      RECT 45.71 4.91 45.88 5.08 ;
      RECT 45.23 3.23 45.4 3.4 ;
      RECT 45.23 4.91 45.4 5.08 ;
      RECT 44.27 3.23 44.44 3.4 ;
      RECT 44.27 3.79 44.44 3.96 ;
      RECT 44.27 4.35 44.44 4.52 ;
      RECT 44.27 4.91 44.44 5.08 ;
      RECT 43.75 4.91 43.92 5.08 ;
      RECT 43.27 3.23 43.44 3.4 ;
      RECT 43.03 3.79 43.2 3.96 ;
      RECT 42.55 3.79 42.72 3.96 ;
      RECT 42.55 4.35 42.72 4.52 ;
      RECT 42.31 3.23 42.48 3.4 ;
      RECT 41.83 4.35 42 4.52 ;
      RECT 41.31 3.79 41.48 3.96 ;
      RECT 41.31 4.63 41.48 4.8 ;
      RECT 40.83 3.23 41 3.4 ;
      RECT 40.83 4.35 41 4.52 ;
      RECT 40.35 4.63 40.52 4.8 ;
      RECT 40.11 4.07 40.28 4.24 ;
      RECT 39.305 3.79 39.475 3.96 ;
      RECT 38.39 3.23 38.56 3.4 ;
      RECT 38.39 4.35 38.56 4.52 ;
      RECT 38.15 3.79 38.32 3.96 ;
      RECT 37.43 3.23 37.6 3.4 ;
      RECT 37.43 4.77 37.6 4.94 ;
      RECT 35.82 7.305 35.99 7.475 ;
      RECT 35.815 8.605 35.985 8.775 ;
      RECT 35.815 10.085 35.985 10.255 ;
      RECT 35.445 8.235 35.615 8.405 ;
      RECT 35.44 4.06 35.61 4.23 ;
      RECT 34.82 2.205 34.99 2.375 ;
      RECT 34.82 3.685 34.99 3.855 ;
      RECT 34.82 8.61 34.99 8.78 ;
      RECT 34.82 10.09 34.99 10.26 ;
      RECT 34.45 4.055 34.62 4.225 ;
      RECT 34.45 8.24 34.62 8.41 ;
      RECT 33.46 3.315 33.63 3.485 ;
      RECT 33.46 8.98 33.63 9.15 ;
      RECT 33.03 2.205 33.2 2.375 ;
      RECT 33.03 2.945 33.2 3.115 ;
      RECT 33.03 9.35 33.2 9.52 ;
      RECT 33.03 10.09 33.2 10.26 ;
      RECT 32.66 3.685 32.83 3.855 ;
      RECT 32.66 8.61 32.83 8.78 ;
      RECT 29.35 4.07 29.52 4.24 ;
      RECT 29.11 3.23 29.28 3.4 ;
      RECT 28.87 4.35 29.04 4.52 ;
      RECT 28.39 3.79 28.56 3.96 ;
      RECT 28.15 3.23 28.32 3.4 ;
      RECT 28.15 4.35 28.32 4.52 ;
      RECT 28.15 4.91 28.32 5.08 ;
      RECT 27.845 8.98 28.015 9.15 ;
      RECT 27.67 4.35 27.84 4.52 ;
      RECT 27.415 9.35 27.585 9.52 ;
      RECT 27.415 10.09 27.585 10.26 ;
      RECT 27.15 4.07 27.32 4.24 ;
      RECT 27.15 4.91 27.32 5.08 ;
      RECT 26.67 3.23 26.84 3.4 ;
      RECT 26.67 4.91 26.84 5.08 ;
      RECT 25.71 3.23 25.88 3.4 ;
      RECT 25.71 3.79 25.88 3.96 ;
      RECT 25.71 4.35 25.88 4.52 ;
      RECT 25.71 4.91 25.88 5.08 ;
      RECT 25.19 4.91 25.36 5.08 ;
      RECT 24.71 3.23 24.88 3.4 ;
      RECT 24.47 3.79 24.64 3.96 ;
      RECT 23.99 3.79 24.16 3.96 ;
      RECT 23.99 4.35 24.16 4.52 ;
      RECT 23.75 3.23 23.92 3.4 ;
      RECT 23.27 4.35 23.44 4.52 ;
      RECT 22.75 3.79 22.92 3.96 ;
      RECT 22.75 4.63 22.92 4.8 ;
      RECT 22.27 3.23 22.44 3.4 ;
      RECT 22.27 4.35 22.44 4.52 ;
      RECT 21.79 4.63 21.96 4.8 ;
      RECT 21.55 4.07 21.72 4.24 ;
      RECT 20.745 3.79 20.915 3.96 ;
      RECT 19.83 3.23 20 3.4 ;
      RECT 19.83 4.35 20 4.52 ;
      RECT 19.59 3.79 19.76 3.96 ;
      RECT 18.87 3.23 19.04 3.4 ;
      RECT 18.87 4.77 19.04 4.94 ;
      RECT 16.6 9.35 16.77 9.52 ;
      RECT 16.6 10.09 16.77 10.26 ;
      RECT 16.23 8.61 16.4 8.78 ;
    LAYER li1 ;
      RECT 110.055 7.305 110.225 8.775 ;
      RECT 110.055 7.305 110.23 8.565 ;
      RECT 109.685 9.255 110.155 9.425 ;
      RECT 109.685 8.235 109.855 9.425 ;
      RECT 109.68 3.04 109.85 4.23 ;
      RECT 109.68 3.04 110.15 3.21 ;
      RECT 109.06 3.895 109.235 5.155 ;
      RECT 109.06 3.685 109.23 5.155 ;
      RECT 109.06 7.31 109.23 8.78 ;
      RECT 109.06 7.31 109.235 8.57 ;
      RECT 108.69 3.035 108.86 4.225 ;
      RECT 108.69 3.035 109.16 3.205 ;
      RECT 108.69 9.26 109.16 9.43 ;
      RECT 108.69 8.24 108.86 9.43 ;
      RECT 107.7 4.015 107.875 5.155 ;
      RECT 107.7 1.865 107.87 5.155 ;
      RECT 107.7 1.865 107.875 2.415 ;
      RECT 107.7 10.05 107.875 10.6 ;
      RECT 107.7 7.31 107.87 10.6 ;
      RECT 107.7 7.31 107.875 8.45 ;
      RECT 107.27 3.895 107.445 5.155 ;
      RECT 107.27 2.945 107.44 5.155 ;
      RECT 107.27 7.31 107.44 9.52 ;
      RECT 107.27 7.31 107.445 8.57 ;
      RECT 106.84 3.925 107.01 5.155 ;
      RECT 106.9 2.145 107.07 4.095 ;
      RECT 106.84 1.865 107.01 2.315 ;
      RECT 106.84 10.15 107.01 10.6 ;
      RECT 106.9 8.37 107.07 10.32 ;
      RECT 106.84 7.31 107.01 8.54 ;
      RECT 106.315 3.895 106.49 5.155 ;
      RECT 106.315 1.865 106.485 5.155 ;
      RECT 106.315 3.365 106.725 3.695 ;
      RECT 106.315 2.525 106.725 2.855 ;
      RECT 106.315 1.865 106.49 2.355 ;
      RECT 106.315 10.11 106.49 10.6 ;
      RECT 106.315 7.31 106.485 10.6 ;
      RECT 106.315 9.61 106.725 9.94 ;
      RECT 106.315 8.77 106.725 9.1 ;
      RECT 106.315 7.31 106.49 8.57 ;
      RECT 103.11 4.52 104.08 4.69 ;
      RECT 103.11 4.35 103.28 4.69 ;
      RECT 102.63 3.79 102.8 4.12 ;
      RECT 102.63 3.87 103.36 4.04 ;
      RECT 102.27 4.91 102.56 5.08 ;
      RECT 102.27 3.87 102.44 5.08 ;
      RECT 102.27 4.35 102.56 4.52 ;
      RECT 102.07 3.87 102.44 4.04 ;
      RECT 102.085 10.05 102.26 10.6 ;
      RECT 102.085 7.31 102.255 10.6 ;
      RECT 102.085 7.31 102.26 8.45 ;
      RECT 101.655 7.31 101.825 9.52 ;
      RECT 101.655 7.31 101.83 8.57 ;
      RECT 101.39 3.97 101.56 4.24 ;
      RECT 101.15 3.97 101.56 4.14 ;
      RECT 101.07 3.87 101.4 4.04 ;
      RECT 100.91 4.91 101.56 5.08 ;
      RECT 101.39 4.44 101.56 5.08 ;
      RECT 101.27 4.52 101.56 5.08 ;
      RECT 100.7 10.11 100.875 10.6 ;
      RECT 100.7 7.31 100.87 10.6 ;
      RECT 100.7 9.61 101.11 9.94 ;
      RECT 100.7 8.77 101.11 9.1 ;
      RECT 100.7 7.31 100.875 8.57 ;
      RECT 99.95 4.21 100.12 4.52 ;
      RECT 99.95 4.21 100.84 4.38 ;
      RECT 100.67 3.79 100.84 4.38 ;
      RECT 99.95 3.87 100.44 4.04 ;
      RECT 99.95 3.79 100.12 4.04 ;
      RECT 97.91 4.52 98.4 4.69 ;
      RECT 99.07 3.87 99.24 4.52 ;
      RECT 98.23 4.35 99.24 4.52 ;
      RECT 99.19 3.79 99.36 4.12 ;
      RECT 97.99 3.13 98.16 3.4 ;
      RECT 97.43 3.13 98.16 3.3 ;
      RECT 97.51 3.87 97.68 4.52 ;
      RECT 97.51 3.87 98 4.04 ;
      RECT 96.67 3.87 97.16 4.04 ;
      RECT 96.99 3.79 97.16 4.04 ;
      RECT 96.51 3.13 96.68 3.4 ;
      RECT 95.95 3.13 96.68 3.3 ;
      RECT 96.03 4.52 96.2 4.8 ;
      RECT 94.99 4.52 96.28 4.69 ;
      RECT 94.985 3.87 95.56 4.04 ;
      RECT 94.985 3.79 95.155 4.04 ;
      RECT 94.07 3.13 94.24 3.4 ;
      RECT 94.07 3.13 94.8 3.3 ;
      RECT 94.07 4.35 94.24 4.77 ;
      RECT 93.45 4.435 94.24 4.605 ;
      RECT 93.45 4.21 93.62 4.605 ;
      RECT 93.35 3.79 93.52 4.38 ;
      RECT 93.11 3.87 93.52 4.14 ;
      RECT 91.495 7.305 91.665 8.775 ;
      RECT 91.495 7.305 91.67 8.565 ;
      RECT 91.125 9.255 91.595 9.425 ;
      RECT 91.125 8.235 91.295 9.425 ;
      RECT 91.12 3.04 91.29 4.23 ;
      RECT 91.12 3.04 91.59 3.21 ;
      RECT 90.5 3.895 90.675 5.155 ;
      RECT 90.5 3.685 90.67 5.155 ;
      RECT 90.5 7.31 90.67 8.78 ;
      RECT 90.5 7.31 90.675 8.57 ;
      RECT 90.13 3.035 90.3 4.225 ;
      RECT 90.13 3.035 90.6 3.205 ;
      RECT 90.13 9.26 90.6 9.43 ;
      RECT 90.13 8.24 90.3 9.43 ;
      RECT 89.14 4.015 89.315 5.155 ;
      RECT 89.14 1.865 89.31 5.155 ;
      RECT 89.14 1.865 89.315 2.415 ;
      RECT 89.14 10.05 89.315 10.6 ;
      RECT 89.14 7.31 89.31 10.6 ;
      RECT 89.14 7.31 89.315 8.45 ;
      RECT 88.71 3.895 88.885 5.155 ;
      RECT 88.71 2.945 88.88 5.155 ;
      RECT 88.71 7.31 88.88 9.52 ;
      RECT 88.71 7.31 88.885 8.57 ;
      RECT 88.28 3.925 88.45 5.155 ;
      RECT 88.34 2.145 88.51 4.095 ;
      RECT 88.28 1.865 88.45 2.315 ;
      RECT 88.28 10.15 88.45 10.6 ;
      RECT 88.34 8.37 88.51 10.32 ;
      RECT 88.28 7.31 88.45 8.54 ;
      RECT 87.755 3.895 87.93 5.155 ;
      RECT 87.755 1.865 87.925 5.155 ;
      RECT 87.755 3.365 88.165 3.695 ;
      RECT 87.755 2.525 88.165 2.855 ;
      RECT 87.755 1.865 87.93 2.355 ;
      RECT 87.755 10.11 87.93 10.6 ;
      RECT 87.755 7.31 87.925 10.6 ;
      RECT 87.755 9.61 88.165 9.94 ;
      RECT 87.755 8.77 88.165 9.1 ;
      RECT 87.755 7.31 87.93 8.57 ;
      RECT 84.55 4.52 85.52 4.69 ;
      RECT 84.55 4.35 84.72 4.69 ;
      RECT 84.07 3.79 84.24 4.12 ;
      RECT 84.07 3.87 84.8 4.04 ;
      RECT 83.71 4.91 84 5.08 ;
      RECT 83.71 3.87 83.88 5.08 ;
      RECT 83.71 4.35 84 4.52 ;
      RECT 83.51 3.87 83.88 4.04 ;
      RECT 83.525 10.05 83.7 10.6 ;
      RECT 83.525 7.31 83.695 10.6 ;
      RECT 83.525 7.31 83.7 8.45 ;
      RECT 83.095 7.31 83.265 9.52 ;
      RECT 83.095 7.31 83.27 8.57 ;
      RECT 82.83 3.97 83 4.24 ;
      RECT 82.59 3.97 83 4.14 ;
      RECT 82.51 3.87 82.84 4.04 ;
      RECT 82.35 4.91 83 5.08 ;
      RECT 82.83 4.44 83 5.08 ;
      RECT 82.71 4.52 83 5.08 ;
      RECT 82.14 10.11 82.315 10.6 ;
      RECT 82.14 7.31 82.31 10.6 ;
      RECT 82.14 9.61 82.55 9.94 ;
      RECT 82.14 8.77 82.55 9.1 ;
      RECT 82.14 7.31 82.315 8.57 ;
      RECT 81.39 4.21 81.56 4.52 ;
      RECT 81.39 4.21 82.28 4.38 ;
      RECT 82.11 3.79 82.28 4.38 ;
      RECT 81.39 3.87 81.88 4.04 ;
      RECT 81.39 3.79 81.56 4.04 ;
      RECT 79.35 4.52 79.84 4.69 ;
      RECT 80.51 3.87 80.68 4.52 ;
      RECT 79.67 4.35 80.68 4.52 ;
      RECT 80.63 3.79 80.8 4.12 ;
      RECT 79.43 3.13 79.6 3.4 ;
      RECT 78.87 3.13 79.6 3.3 ;
      RECT 78.95 3.87 79.12 4.52 ;
      RECT 78.95 3.87 79.44 4.04 ;
      RECT 78.11 3.87 78.6 4.04 ;
      RECT 78.43 3.79 78.6 4.04 ;
      RECT 77.95 3.13 78.12 3.4 ;
      RECT 77.39 3.13 78.12 3.3 ;
      RECT 77.47 4.52 77.64 4.8 ;
      RECT 76.43 4.52 77.72 4.69 ;
      RECT 76.425 3.87 77 4.04 ;
      RECT 76.425 3.79 76.595 4.04 ;
      RECT 75.51 3.13 75.68 3.4 ;
      RECT 75.51 3.13 76.24 3.3 ;
      RECT 75.51 4.35 75.68 4.77 ;
      RECT 74.89 4.435 75.68 4.605 ;
      RECT 74.89 4.21 75.06 4.605 ;
      RECT 74.79 3.79 74.96 4.38 ;
      RECT 74.55 3.87 74.96 4.14 ;
      RECT 72.935 7.305 73.105 8.775 ;
      RECT 72.935 7.305 73.11 8.565 ;
      RECT 72.565 9.255 73.035 9.425 ;
      RECT 72.565 8.235 72.735 9.425 ;
      RECT 72.56 3.04 72.73 4.23 ;
      RECT 72.56 3.04 73.03 3.21 ;
      RECT 71.94 3.895 72.115 5.155 ;
      RECT 71.94 3.685 72.11 5.155 ;
      RECT 71.94 7.31 72.11 8.78 ;
      RECT 71.94 7.31 72.115 8.57 ;
      RECT 71.57 3.035 71.74 4.225 ;
      RECT 71.57 3.035 72.04 3.205 ;
      RECT 71.57 9.26 72.04 9.43 ;
      RECT 71.57 8.24 71.74 9.43 ;
      RECT 70.58 4.015 70.755 5.155 ;
      RECT 70.58 1.865 70.75 5.155 ;
      RECT 70.58 1.865 70.755 2.415 ;
      RECT 70.58 10.05 70.755 10.6 ;
      RECT 70.58 7.31 70.75 10.6 ;
      RECT 70.58 7.31 70.755 8.45 ;
      RECT 70.15 3.895 70.325 5.155 ;
      RECT 70.15 2.945 70.32 5.155 ;
      RECT 70.15 7.31 70.32 9.52 ;
      RECT 70.15 7.31 70.325 8.57 ;
      RECT 69.72 3.925 69.89 5.155 ;
      RECT 69.78 2.145 69.95 4.095 ;
      RECT 69.72 1.865 69.89 2.315 ;
      RECT 69.72 10.15 69.89 10.6 ;
      RECT 69.78 8.37 69.95 10.32 ;
      RECT 69.72 7.31 69.89 8.54 ;
      RECT 69.195 3.895 69.37 5.155 ;
      RECT 69.195 1.865 69.365 5.155 ;
      RECT 69.195 3.365 69.605 3.695 ;
      RECT 69.195 2.525 69.605 2.855 ;
      RECT 69.195 1.865 69.37 2.355 ;
      RECT 69.195 10.11 69.37 10.6 ;
      RECT 69.195 7.31 69.365 10.6 ;
      RECT 69.195 9.61 69.605 9.94 ;
      RECT 69.195 8.77 69.605 9.1 ;
      RECT 69.195 7.31 69.37 8.57 ;
      RECT 65.99 4.52 66.96 4.69 ;
      RECT 65.99 4.35 66.16 4.69 ;
      RECT 65.51 3.79 65.68 4.12 ;
      RECT 65.51 3.87 66.24 4.04 ;
      RECT 65.15 4.91 65.44 5.08 ;
      RECT 65.15 3.87 65.32 5.08 ;
      RECT 65.15 4.35 65.44 4.52 ;
      RECT 64.95 3.87 65.32 4.04 ;
      RECT 64.965 10.05 65.14 10.6 ;
      RECT 64.965 7.31 65.135 10.6 ;
      RECT 64.965 7.31 65.14 8.45 ;
      RECT 64.535 7.31 64.705 9.52 ;
      RECT 64.535 7.31 64.71 8.57 ;
      RECT 64.27 3.97 64.44 4.24 ;
      RECT 64.03 3.97 64.44 4.14 ;
      RECT 63.95 3.87 64.28 4.04 ;
      RECT 63.79 4.91 64.44 5.08 ;
      RECT 64.27 4.44 64.44 5.08 ;
      RECT 64.15 4.52 64.44 5.08 ;
      RECT 63.58 10.11 63.755 10.6 ;
      RECT 63.58 7.31 63.75 10.6 ;
      RECT 63.58 9.61 63.99 9.94 ;
      RECT 63.58 8.77 63.99 9.1 ;
      RECT 63.58 7.31 63.755 8.57 ;
      RECT 62.83 4.21 63 4.52 ;
      RECT 62.83 4.21 63.72 4.38 ;
      RECT 63.55 3.79 63.72 4.38 ;
      RECT 62.83 3.87 63.32 4.04 ;
      RECT 62.83 3.79 63 4.04 ;
      RECT 60.79 4.52 61.28 4.69 ;
      RECT 61.95 3.87 62.12 4.52 ;
      RECT 61.11 4.35 62.12 4.52 ;
      RECT 62.07 3.79 62.24 4.12 ;
      RECT 60.87 3.13 61.04 3.4 ;
      RECT 60.31 3.13 61.04 3.3 ;
      RECT 60.39 3.87 60.56 4.52 ;
      RECT 60.39 3.87 60.88 4.04 ;
      RECT 59.55 3.87 60.04 4.04 ;
      RECT 59.87 3.79 60.04 4.04 ;
      RECT 59.39 3.13 59.56 3.4 ;
      RECT 58.83 3.13 59.56 3.3 ;
      RECT 58.91 4.52 59.08 4.8 ;
      RECT 57.87 4.52 59.16 4.69 ;
      RECT 57.865 3.87 58.44 4.04 ;
      RECT 57.865 3.79 58.035 4.04 ;
      RECT 56.95 3.13 57.12 3.4 ;
      RECT 56.95 3.13 57.68 3.3 ;
      RECT 56.95 4.35 57.12 4.77 ;
      RECT 56.33 4.435 57.12 4.605 ;
      RECT 56.33 4.21 56.5 4.605 ;
      RECT 56.23 3.79 56.4 4.38 ;
      RECT 55.99 3.87 56.4 4.14 ;
      RECT 54.375 7.305 54.545 8.775 ;
      RECT 54.375 7.305 54.55 8.565 ;
      RECT 54.005 9.255 54.475 9.425 ;
      RECT 54.005 8.235 54.175 9.425 ;
      RECT 54 3.04 54.17 4.23 ;
      RECT 54 3.04 54.47 3.21 ;
      RECT 53.38 3.895 53.555 5.155 ;
      RECT 53.38 3.685 53.55 5.155 ;
      RECT 53.38 7.31 53.55 8.78 ;
      RECT 53.38 7.31 53.555 8.57 ;
      RECT 53.01 3.035 53.18 4.225 ;
      RECT 53.01 3.035 53.48 3.205 ;
      RECT 53.01 9.26 53.48 9.43 ;
      RECT 53.01 8.24 53.18 9.43 ;
      RECT 52.02 4.015 52.195 5.155 ;
      RECT 52.02 1.865 52.19 5.155 ;
      RECT 52.02 1.865 52.195 2.415 ;
      RECT 52.02 10.05 52.195 10.6 ;
      RECT 52.02 7.31 52.19 10.6 ;
      RECT 52.02 7.31 52.195 8.45 ;
      RECT 51.59 3.895 51.765 5.155 ;
      RECT 51.59 2.945 51.76 5.155 ;
      RECT 51.59 7.31 51.76 9.52 ;
      RECT 51.59 7.31 51.765 8.57 ;
      RECT 51.16 3.925 51.33 5.155 ;
      RECT 51.22 2.145 51.39 4.095 ;
      RECT 51.16 1.865 51.33 2.315 ;
      RECT 51.16 10.15 51.33 10.6 ;
      RECT 51.22 8.37 51.39 10.32 ;
      RECT 51.16 7.31 51.33 8.54 ;
      RECT 50.635 3.895 50.81 5.155 ;
      RECT 50.635 1.865 50.805 5.155 ;
      RECT 50.635 3.365 51.045 3.695 ;
      RECT 50.635 2.525 51.045 2.855 ;
      RECT 50.635 1.865 50.81 2.355 ;
      RECT 50.635 10.11 50.81 10.6 ;
      RECT 50.635 7.31 50.805 10.6 ;
      RECT 50.635 9.61 51.045 9.94 ;
      RECT 50.635 8.77 51.045 9.1 ;
      RECT 50.635 7.31 50.81 8.57 ;
      RECT 47.43 4.52 48.4 4.69 ;
      RECT 47.43 4.35 47.6 4.69 ;
      RECT 46.95 3.79 47.12 4.12 ;
      RECT 46.95 3.87 47.68 4.04 ;
      RECT 46.59 4.91 46.88 5.08 ;
      RECT 46.59 3.87 46.76 5.08 ;
      RECT 46.59 4.35 46.88 4.52 ;
      RECT 46.39 3.87 46.76 4.04 ;
      RECT 46.405 10.05 46.58 10.6 ;
      RECT 46.405 7.31 46.575 10.6 ;
      RECT 46.405 7.31 46.58 8.45 ;
      RECT 45.975 7.31 46.145 9.52 ;
      RECT 45.975 7.31 46.15 8.57 ;
      RECT 45.71 3.97 45.88 4.24 ;
      RECT 45.47 3.97 45.88 4.14 ;
      RECT 45.39 3.87 45.72 4.04 ;
      RECT 45.23 4.91 45.88 5.08 ;
      RECT 45.71 4.44 45.88 5.08 ;
      RECT 45.59 4.52 45.88 5.08 ;
      RECT 45.02 10.11 45.195 10.6 ;
      RECT 45.02 7.31 45.19 10.6 ;
      RECT 45.02 9.61 45.43 9.94 ;
      RECT 45.02 8.77 45.43 9.1 ;
      RECT 45.02 7.31 45.195 8.57 ;
      RECT 44.27 4.21 44.44 4.52 ;
      RECT 44.27 4.21 45.16 4.38 ;
      RECT 44.99 3.79 45.16 4.38 ;
      RECT 44.27 3.87 44.76 4.04 ;
      RECT 44.27 3.79 44.44 4.04 ;
      RECT 42.23 4.52 42.72 4.69 ;
      RECT 43.39 3.87 43.56 4.52 ;
      RECT 42.55 4.35 43.56 4.52 ;
      RECT 43.51 3.79 43.68 4.12 ;
      RECT 42.31 3.13 42.48 3.4 ;
      RECT 41.75 3.13 42.48 3.3 ;
      RECT 41.83 3.87 42 4.52 ;
      RECT 41.83 3.87 42.32 4.04 ;
      RECT 40.99 3.87 41.48 4.04 ;
      RECT 41.31 3.79 41.48 4.04 ;
      RECT 40.83 3.13 41 3.4 ;
      RECT 40.27 3.13 41 3.3 ;
      RECT 40.35 4.52 40.52 4.8 ;
      RECT 39.31 4.52 40.6 4.69 ;
      RECT 39.305 3.87 39.88 4.04 ;
      RECT 39.305 3.79 39.475 4.04 ;
      RECT 38.39 3.13 38.56 3.4 ;
      RECT 38.39 3.13 39.12 3.3 ;
      RECT 38.39 4.35 38.56 4.77 ;
      RECT 37.77 4.435 38.56 4.605 ;
      RECT 37.77 4.21 37.94 4.605 ;
      RECT 37.67 3.79 37.84 4.38 ;
      RECT 37.43 3.87 37.84 4.14 ;
      RECT 35.815 7.305 35.985 8.775 ;
      RECT 35.815 7.305 35.99 8.565 ;
      RECT 35.445 9.255 35.915 9.425 ;
      RECT 35.445 8.235 35.615 9.425 ;
      RECT 35.44 3.04 35.61 4.23 ;
      RECT 35.44 3.04 35.91 3.21 ;
      RECT 34.82 3.895 34.995 5.155 ;
      RECT 34.82 3.685 34.99 5.155 ;
      RECT 34.82 7.31 34.99 8.78 ;
      RECT 34.82 7.31 34.995 8.57 ;
      RECT 34.45 3.035 34.62 4.225 ;
      RECT 34.45 3.035 34.92 3.205 ;
      RECT 34.45 9.26 34.92 9.43 ;
      RECT 34.45 8.24 34.62 9.43 ;
      RECT 33.46 4.015 33.635 5.155 ;
      RECT 33.46 1.865 33.63 5.155 ;
      RECT 33.46 1.865 33.635 2.415 ;
      RECT 33.46 10.05 33.635 10.6 ;
      RECT 33.46 7.31 33.63 10.6 ;
      RECT 33.46 7.31 33.635 8.45 ;
      RECT 33.03 3.895 33.205 5.155 ;
      RECT 33.03 2.945 33.2 5.155 ;
      RECT 33.03 7.31 33.2 9.52 ;
      RECT 33.03 7.31 33.205 8.57 ;
      RECT 32.6 3.925 32.77 5.155 ;
      RECT 32.66 2.145 32.83 4.095 ;
      RECT 32.6 1.865 32.77 2.315 ;
      RECT 32.6 10.15 32.77 10.6 ;
      RECT 32.66 8.37 32.83 10.32 ;
      RECT 32.6 7.31 32.77 8.54 ;
      RECT 32.075 3.895 32.25 5.155 ;
      RECT 32.075 1.865 32.245 5.155 ;
      RECT 32.075 3.365 32.485 3.695 ;
      RECT 32.075 2.525 32.485 2.855 ;
      RECT 32.075 1.865 32.25 2.355 ;
      RECT 32.075 10.11 32.25 10.6 ;
      RECT 32.075 7.31 32.245 10.6 ;
      RECT 32.075 9.61 32.485 9.94 ;
      RECT 32.075 8.77 32.485 9.1 ;
      RECT 32.075 7.31 32.25 8.57 ;
      RECT 28.87 4.52 29.84 4.69 ;
      RECT 28.87 4.35 29.04 4.69 ;
      RECT 28.39 3.79 28.56 4.12 ;
      RECT 28.39 3.87 29.12 4.04 ;
      RECT 28.03 4.91 28.32 5.08 ;
      RECT 28.03 3.87 28.2 5.08 ;
      RECT 28.03 4.35 28.32 4.52 ;
      RECT 27.83 3.87 28.2 4.04 ;
      RECT 27.845 10.05 28.02 10.6 ;
      RECT 27.845 7.31 28.015 10.6 ;
      RECT 27.845 7.31 28.02 8.45 ;
      RECT 27.415 7.31 27.585 9.52 ;
      RECT 27.415 7.31 27.59 8.57 ;
      RECT 27.15 3.97 27.32 4.24 ;
      RECT 26.91 3.97 27.32 4.14 ;
      RECT 26.83 3.87 27.16 4.04 ;
      RECT 26.67 4.91 27.32 5.08 ;
      RECT 27.15 4.44 27.32 5.08 ;
      RECT 27.03 4.52 27.32 5.08 ;
      RECT 26.46 10.11 26.635 10.6 ;
      RECT 26.46 7.31 26.63 10.6 ;
      RECT 26.46 9.61 26.87 9.94 ;
      RECT 26.46 8.77 26.87 9.1 ;
      RECT 26.46 7.31 26.635 8.57 ;
      RECT 25.71 4.21 25.88 4.52 ;
      RECT 25.71 4.21 26.6 4.38 ;
      RECT 26.43 3.79 26.6 4.38 ;
      RECT 25.71 3.87 26.2 4.04 ;
      RECT 25.71 3.79 25.88 4.04 ;
      RECT 23.67 4.52 24.16 4.69 ;
      RECT 24.83 3.87 25 4.52 ;
      RECT 23.99 4.35 25 4.52 ;
      RECT 24.95 3.79 25.12 4.12 ;
      RECT 23.75 3.13 23.92 3.4 ;
      RECT 23.19 3.13 23.92 3.3 ;
      RECT 23.27 3.87 23.44 4.52 ;
      RECT 23.27 3.87 23.76 4.04 ;
      RECT 22.43 3.87 22.92 4.04 ;
      RECT 22.75 3.79 22.92 4.04 ;
      RECT 22.27 3.13 22.44 3.4 ;
      RECT 21.71 3.13 22.44 3.3 ;
      RECT 21.79 4.52 21.96 4.8 ;
      RECT 20.75 4.52 22.04 4.69 ;
      RECT 20.745 3.87 21.32 4.04 ;
      RECT 20.745 3.79 20.915 4.04 ;
      RECT 19.83 3.13 20 3.4 ;
      RECT 19.83 3.13 20.56 3.3 ;
      RECT 19.83 4.35 20 4.77 ;
      RECT 19.21 4.435 20 4.605 ;
      RECT 19.21 4.21 19.38 4.605 ;
      RECT 19.11 3.79 19.28 4.38 ;
      RECT 18.87 3.87 19.28 4.14 ;
      RECT 16.6 7.31 16.77 9.52 ;
      RECT 16.6 7.31 16.775 8.57 ;
      RECT 16.17 10.15 16.34 10.6 ;
      RECT 16.23 8.37 16.4 10.32 ;
      RECT 16.17 7.31 16.34 8.54 ;
      RECT 15.645 10.11 15.82 10.6 ;
      RECT 15.645 7.31 15.815 10.6 ;
      RECT 15.645 9.61 16.055 9.94 ;
      RECT 15.645 8.77 16.055 9.1 ;
      RECT 15.645 7.31 15.82 8.57 ;
      RECT 110.055 10.085 110.23 10.595 ;
      RECT 109.06 1.865 109.235 2.375 ;
      RECT 109.06 10.09 109.235 10.6 ;
      RECT 107.27 1.865 107.445 2.375 ;
      RECT 107.27 10.09 107.445 10.6 ;
      RECT 103.59 3.79 103.76 4.24 ;
      RECT 103.35 3.05 103.52 3.4 ;
      RECT 102.39 3.05 102.56 3.4 ;
      RECT 101.91 4.35 102.08 4.77 ;
      RECT 101.655 10.09 101.83 10.6 ;
      RECT 100.91 3.05 101.08 3.4 ;
      RECT 99.95 3.05 100.12 3.4 ;
      RECT 99.95 4.78 100.12 5.11 ;
      RECT 99.43 4.44 99.6 5.08 ;
      RECT 98.95 3.05 99.12 3.4 ;
      RECT 98.71 3.79 98.88 4.12 ;
      RECT 98.23 3.79 98.4 4.12 ;
      RECT 96.99 4.44 97.16 4.8 ;
      RECT 96.51 4.35 96.68 4.77 ;
      RECT 95.79 3.79 95.96 4.24 ;
      RECT 93.83 3.79 94 4.12 ;
      RECT 93.11 3.05 93.28 3.4 ;
      RECT 93.11 4.58 93.28 4.94 ;
      RECT 91.495 10.085 91.67 10.595 ;
      RECT 90.5 1.865 90.675 2.375 ;
      RECT 90.5 10.09 90.675 10.6 ;
      RECT 88.71 1.865 88.885 2.375 ;
      RECT 88.71 10.09 88.885 10.6 ;
      RECT 85.03 3.79 85.2 4.24 ;
      RECT 84.79 3.05 84.96 3.4 ;
      RECT 83.83 3.05 84 3.4 ;
      RECT 83.35 4.35 83.52 4.77 ;
      RECT 83.095 10.09 83.27 10.6 ;
      RECT 82.35 3.05 82.52 3.4 ;
      RECT 81.39 3.05 81.56 3.4 ;
      RECT 81.39 4.78 81.56 5.11 ;
      RECT 80.87 4.44 81.04 5.08 ;
      RECT 80.39 3.05 80.56 3.4 ;
      RECT 80.15 3.79 80.32 4.12 ;
      RECT 79.67 3.79 79.84 4.12 ;
      RECT 78.43 4.44 78.6 4.8 ;
      RECT 77.95 4.35 78.12 4.77 ;
      RECT 77.23 3.79 77.4 4.24 ;
      RECT 75.27 3.79 75.44 4.12 ;
      RECT 74.55 3.05 74.72 3.4 ;
      RECT 74.55 4.58 74.72 4.94 ;
      RECT 72.935 10.085 73.11 10.595 ;
      RECT 71.94 1.865 72.115 2.375 ;
      RECT 71.94 10.09 72.115 10.6 ;
      RECT 70.15 1.865 70.325 2.375 ;
      RECT 70.15 10.09 70.325 10.6 ;
      RECT 66.47 3.79 66.64 4.24 ;
      RECT 66.23 3.05 66.4 3.4 ;
      RECT 65.27 3.05 65.44 3.4 ;
      RECT 64.79 4.35 64.96 4.77 ;
      RECT 64.535 10.09 64.71 10.6 ;
      RECT 63.79 3.05 63.96 3.4 ;
      RECT 62.83 3.05 63 3.4 ;
      RECT 62.83 4.78 63 5.11 ;
      RECT 62.31 4.44 62.48 5.08 ;
      RECT 61.83 3.05 62 3.4 ;
      RECT 61.59 3.79 61.76 4.12 ;
      RECT 61.11 3.79 61.28 4.12 ;
      RECT 59.87 4.44 60.04 4.8 ;
      RECT 59.39 4.35 59.56 4.77 ;
      RECT 58.67 3.79 58.84 4.24 ;
      RECT 56.71 3.79 56.88 4.12 ;
      RECT 55.99 3.05 56.16 3.4 ;
      RECT 55.99 4.58 56.16 4.94 ;
      RECT 54.375 10.085 54.55 10.595 ;
      RECT 53.38 1.865 53.555 2.375 ;
      RECT 53.38 10.09 53.555 10.6 ;
      RECT 51.59 1.865 51.765 2.375 ;
      RECT 51.59 10.09 51.765 10.6 ;
      RECT 47.91 3.79 48.08 4.24 ;
      RECT 47.67 3.05 47.84 3.4 ;
      RECT 46.71 3.05 46.88 3.4 ;
      RECT 46.23 4.35 46.4 4.77 ;
      RECT 45.975 10.09 46.15 10.6 ;
      RECT 45.23 3.05 45.4 3.4 ;
      RECT 44.27 3.05 44.44 3.4 ;
      RECT 44.27 4.78 44.44 5.11 ;
      RECT 43.75 4.44 43.92 5.08 ;
      RECT 43.27 3.05 43.44 3.4 ;
      RECT 43.03 3.79 43.2 4.12 ;
      RECT 42.55 3.79 42.72 4.12 ;
      RECT 41.31 4.44 41.48 4.8 ;
      RECT 40.83 4.35 41 4.77 ;
      RECT 40.11 3.79 40.28 4.24 ;
      RECT 38.15 3.79 38.32 4.12 ;
      RECT 37.43 3.05 37.6 3.4 ;
      RECT 37.43 4.58 37.6 4.94 ;
      RECT 35.815 10.085 35.99 10.595 ;
      RECT 34.82 1.865 34.995 2.375 ;
      RECT 34.82 10.09 34.995 10.6 ;
      RECT 33.03 1.865 33.205 2.375 ;
      RECT 33.03 10.09 33.205 10.6 ;
      RECT 29.35 3.79 29.52 4.24 ;
      RECT 29.11 3.05 29.28 3.4 ;
      RECT 28.15 3.05 28.32 3.4 ;
      RECT 27.67 4.35 27.84 4.77 ;
      RECT 27.415 10.09 27.59 10.6 ;
      RECT 26.67 3.05 26.84 3.4 ;
      RECT 25.71 3.05 25.88 3.4 ;
      RECT 25.71 4.78 25.88 5.11 ;
      RECT 25.19 4.44 25.36 5.08 ;
      RECT 24.71 3.05 24.88 3.4 ;
      RECT 24.47 3.79 24.64 4.12 ;
      RECT 23.99 3.79 24.16 4.12 ;
      RECT 22.75 4.44 22.92 4.8 ;
      RECT 22.27 4.35 22.44 4.77 ;
      RECT 21.55 3.79 21.72 4.24 ;
      RECT 19.59 3.79 19.76 4.12 ;
      RECT 18.87 3.05 19.04 3.4 ;
      RECT 18.87 4.58 19.04 4.94 ;
      RECT 16.6 10.09 16.775 10.6 ;
  END
END sky130_osu_ring_oscillator_mpr2et_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2xa_8_b0r1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2xa_8_b0r1 ;
  SIZE 104.045 BY 12.465 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 42.355 0 42.735 5.26 ;
      LAYER met2 ;
        RECT 42.355 4.88 42.735 5.26 ;
      LAYER li1 ;
        RECT 42.455 1.865 42.63 2.375 ;
        RECT 42.455 3.895 42.63 5.155 ;
        RECT 42.455 3.685 42.625 5.155 ;
      LAYER met1 ;
        RECT 42.37 4.925 42.72 5.215 ;
        RECT 42.395 2.175 42.69 2.405 ;
        RECT 42.395 3.655 42.685 3.885 ;
        RECT 42.455 2.175 42.625 3.885 ;
      LAYER via1 ;
        RECT 42.47 4.995 42.62 5.145 ;
      LAYER via2 ;
        RECT 42.445 4.97 42.645 5.17 ;
      LAYER mcon ;
        RECT 42.455 3.685 42.625 3.855 ;
        RECT 42.455 2.205 42.625 2.375 ;
        RECT 42.46 4.985 42.63 5.155 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 57.615 0 57.995 5.26 ;
      LAYER met2 ;
        RECT 57.615 4.88 57.995 5.26 ;
      LAYER li1 ;
        RECT 57.715 1.865 57.89 2.375 ;
        RECT 57.715 3.895 57.89 5.155 ;
        RECT 57.715 3.685 57.885 5.155 ;
      LAYER met1 ;
        RECT 57.63 4.925 57.98 5.215 ;
        RECT 57.655 2.175 57.95 2.405 ;
        RECT 57.655 3.655 57.945 3.885 ;
        RECT 57.715 2.175 57.885 3.885 ;
      LAYER via1 ;
        RECT 57.73 4.995 57.88 5.145 ;
      LAYER via2 ;
        RECT 57.705 4.97 57.905 5.17 ;
      LAYER mcon ;
        RECT 57.715 3.685 57.885 3.855 ;
        RECT 57.715 2.205 57.885 2.375 ;
        RECT 57.72 4.985 57.89 5.155 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 72.875 0 73.255 5.26 ;
      LAYER met2 ;
        RECT 72.875 4.88 73.255 5.26 ;
      LAYER li1 ;
        RECT 72.975 1.865 73.15 2.375 ;
        RECT 72.975 3.895 73.15 5.155 ;
        RECT 72.975 3.685 73.145 5.155 ;
      LAYER met1 ;
        RECT 72.89 4.925 73.24 5.215 ;
        RECT 72.915 2.175 73.21 2.405 ;
        RECT 72.915 3.655 73.205 3.885 ;
        RECT 72.975 2.175 73.145 3.885 ;
      LAYER via1 ;
        RECT 72.99 4.995 73.14 5.145 ;
      LAYER via2 ;
        RECT 72.965 4.97 73.165 5.17 ;
      LAYER mcon ;
        RECT 72.975 3.685 73.145 3.855 ;
        RECT 72.975 2.205 73.145 2.375 ;
        RECT 72.98 4.985 73.15 5.155 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 88.135 0 88.515 5.26 ;
      LAYER met2 ;
        RECT 88.135 4.88 88.515 5.26 ;
      LAYER li1 ;
        RECT 88.235 1.865 88.41 2.375 ;
        RECT 88.235 3.895 88.41 5.155 ;
        RECT 88.235 3.685 88.405 5.155 ;
      LAYER met1 ;
        RECT 88.15 4.925 88.5 5.215 ;
        RECT 88.175 2.175 88.47 2.405 ;
        RECT 88.175 3.655 88.465 3.885 ;
        RECT 88.235 2.175 88.405 3.885 ;
      LAYER via1 ;
        RECT 88.25 4.995 88.4 5.145 ;
      LAYER via2 ;
        RECT 88.225 4.97 88.425 5.17 ;
      LAYER mcon ;
        RECT 88.235 3.685 88.405 3.855 ;
        RECT 88.235 2.205 88.405 2.375 ;
        RECT 88.24 4.985 88.41 5.155 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 103.395 0 103.775 5.26 ;
      LAYER met2 ;
        RECT 103.395 4.88 103.775 5.26 ;
      LAYER li1 ;
        RECT 103.495 1.865 103.67 2.375 ;
        RECT 103.495 3.895 103.67 5.155 ;
        RECT 103.495 3.685 103.665 5.155 ;
      LAYER met1 ;
        RECT 103.41 4.925 103.76 5.215 ;
        RECT 103.435 2.175 103.73 2.405 ;
        RECT 103.435 3.655 103.725 3.885 ;
        RECT 103.495 2.175 103.665 3.885 ;
      LAYER via1 ;
        RECT 103.51 4.995 103.66 5.145 ;
      LAYER via2 ;
        RECT 103.485 4.97 103.685 5.17 ;
      LAYER mcon ;
        RECT 103.495 3.685 103.665 3.855 ;
        RECT 103.495 2.205 103.665 2.375 ;
        RECT 103.5 4.985 103.67 5.155 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 38.23 8.15 38.57 8.5 ;
        RECT 38.23 4 38.57 4.35 ;
        RECT 38.31 4 38.48 8.5 ;
      LAYER li1 ;
        RECT 38.305 2.955 38.475 4.225 ;
        RECT 38.305 8.24 38.475 9.51 ;
        RECT 32.69 8.24 32.86 9.51 ;
      LAYER met1 ;
        RECT 38.23 4.055 38.705 4.225 ;
        RECT 38.23 4 38.57 4.35 ;
        RECT 38.23 8.24 38.705 8.41 ;
        RECT 38.23 8.15 38.57 8.5 ;
        RECT 32.63 8.235 38.57 8.405 ;
        RECT 32.63 8.235 33.09 8.41 ;
        RECT 32.63 8.21 32.92 8.44 ;
      LAYER via1 ;
        RECT 38.33 8.25 38.48 8.4 ;
        RECT 38.33 4.1 38.48 4.25 ;
      LAYER mcon ;
        RECT 32.69 8.24 32.86 8.41 ;
        RECT 38.305 8.24 38.475 8.41 ;
        RECT 38.305 4.055 38.475 4.225 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 53.49 8.15 53.83 8.5 ;
        RECT 53.49 4 53.83 4.35 ;
        RECT 53.57 4 53.74 8.5 ;
      LAYER li1 ;
        RECT 53.565 2.955 53.735 4.225 ;
        RECT 53.565 8.24 53.735 9.51 ;
        RECT 47.95 8.24 48.12 9.51 ;
      LAYER met1 ;
        RECT 53.49 4.055 53.965 4.225 ;
        RECT 53.49 4 53.83 4.35 ;
        RECT 53.49 8.24 53.965 8.41 ;
        RECT 53.49 8.15 53.83 8.5 ;
        RECT 47.89 8.235 53.83 8.405 ;
        RECT 47.89 8.235 48.35 8.41 ;
        RECT 47.89 8.21 48.18 8.44 ;
      LAYER via1 ;
        RECT 53.59 8.25 53.74 8.4 ;
        RECT 53.59 4.1 53.74 4.25 ;
      LAYER mcon ;
        RECT 47.95 8.24 48.12 8.41 ;
        RECT 53.565 8.24 53.735 8.41 ;
        RECT 53.565 4.055 53.735 4.225 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 68.75 8.15 69.09 8.5 ;
        RECT 68.75 4 69.09 4.35 ;
        RECT 68.83 4 69 8.5 ;
      LAYER li1 ;
        RECT 68.825 2.955 68.995 4.225 ;
        RECT 68.825 8.24 68.995 9.51 ;
        RECT 63.21 8.24 63.38 9.51 ;
      LAYER met1 ;
        RECT 68.75 4.055 69.225 4.225 ;
        RECT 68.75 4 69.09 4.35 ;
        RECT 68.75 8.24 69.225 8.41 ;
        RECT 68.75 8.15 69.09 8.5 ;
        RECT 63.15 8.235 69.09 8.405 ;
        RECT 63.15 8.235 63.61 8.41 ;
        RECT 63.15 8.21 63.44 8.44 ;
      LAYER via1 ;
        RECT 68.85 8.25 69 8.4 ;
        RECT 68.85 4.1 69 4.25 ;
      LAYER mcon ;
        RECT 63.21 8.24 63.38 8.41 ;
        RECT 68.825 8.24 68.995 8.41 ;
        RECT 68.825 4.055 68.995 4.225 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 84.01 8.15 84.35 8.5 ;
        RECT 84.01 4 84.35 4.35 ;
        RECT 84.09 4 84.26 8.5 ;
      LAYER li1 ;
        RECT 84.085 2.955 84.255 4.225 ;
        RECT 84.085 8.24 84.255 9.51 ;
        RECT 78.47 8.24 78.64 9.51 ;
      LAYER met1 ;
        RECT 84.01 4.055 84.485 4.225 ;
        RECT 84.01 4 84.35 4.35 ;
        RECT 84.01 8.24 84.485 8.41 ;
        RECT 84.01 8.15 84.35 8.5 ;
        RECT 78.41 8.235 84.35 8.405 ;
        RECT 78.41 8.235 78.87 8.41 ;
        RECT 78.41 8.21 78.7 8.44 ;
      LAYER via1 ;
        RECT 84.11 8.25 84.26 8.4 ;
        RECT 84.11 4.1 84.26 4.25 ;
      LAYER mcon ;
        RECT 78.47 8.24 78.64 8.41 ;
        RECT 84.085 8.24 84.255 8.41 ;
        RECT 84.085 4.055 84.255 4.225 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 99.27 8.15 99.61 8.5 ;
        RECT 99.27 4 99.61 4.35 ;
        RECT 99.35 4 99.52 8.5 ;
      LAYER li1 ;
        RECT 99.345 2.955 99.515 4.225 ;
        RECT 99.345 8.24 99.515 9.51 ;
        RECT 93.73 8.24 93.9 9.51 ;
      LAYER met1 ;
        RECT 99.27 4.055 99.745 4.225 ;
        RECT 99.27 4 99.61 4.35 ;
        RECT 99.27 8.24 99.745 8.41 ;
        RECT 99.27 8.15 99.61 8.5 ;
        RECT 93.67 8.235 99.61 8.405 ;
        RECT 93.67 8.235 94.13 8.41 ;
        RECT 93.67 8.21 93.96 8.44 ;
      LAYER via1 ;
        RECT 99.37 8.25 99.52 8.4 ;
        RECT 99.37 4.1 99.52 4.25 ;
      LAYER mcon ;
        RECT 93.73 8.24 93.9 8.41 ;
        RECT 99.345 8.24 99.515 8.41 ;
        RECT 99.345 4.055 99.515 4.225 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 25.175 8.24 25.345 9.51 ;
      LAYER met1 ;
        RECT 25.115 8.24 25.575 8.41 ;
        RECT 25.12 8.205 25.41 8.435 ;
        RECT 25.115 8.21 25.405 8.44 ;
      LAYER mcon ;
        RECT 25.175 8.24 25.345 8.41 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 5.435 104.045 7.035 ;
        RECT 89.535 5.43 104.045 7.035 ;
        RECT 99.165 5.43 103.89 7.04 ;
        RECT 99.165 5.425 103.885 7.04 ;
        RECT 103.07 5.425 103.24 7.77 ;
        RECT 103.065 4.695 103.235 7.04 ;
        RECT 102.08 4.695 102.25 7.77 ;
        RECT 99.335 4.695 99.505 7.77 ;
        RECT 96.565 4.93 96.735 7.035 ;
        RECT 93.55 5.43 96.3 7.04 ;
        RECT 94.645 4.93 94.815 7.04 ;
        RECT 93.72 5.43 93.89 7.77 ;
        RECT 93.705 4.93 93.875 7.04 ;
        RECT 92.245 4.93 92.415 7.035 ;
        RECT 90.325 4.93 90.495 7.035 ;
        RECT 74.275 5.43 88.785 7.035 ;
        RECT 83.905 5.43 88.63 7.04 ;
        RECT 83.905 5.425 88.625 7.04 ;
        RECT 87.81 5.425 87.98 7.77 ;
        RECT 87.805 4.695 87.975 7.04 ;
        RECT 86.82 4.695 86.99 7.77 ;
        RECT 84.075 4.695 84.245 7.77 ;
        RECT 81.305 4.93 81.475 7.035 ;
        RECT 78.29 5.43 81.04 7.04 ;
        RECT 79.385 4.93 79.555 7.04 ;
        RECT 78.46 5.43 78.63 7.77 ;
        RECT 78.445 4.93 78.615 7.04 ;
        RECT 76.985 4.93 77.155 7.035 ;
        RECT 75.065 4.93 75.235 7.035 ;
        RECT 59.015 5.43 73.525 7.035 ;
        RECT 68.645 5.43 73.37 7.04 ;
        RECT 68.645 5.425 73.365 7.04 ;
        RECT 72.55 5.425 72.72 7.77 ;
        RECT 72.545 4.695 72.715 7.04 ;
        RECT 71.56 4.695 71.73 7.77 ;
        RECT 68.815 4.695 68.985 7.77 ;
        RECT 66.045 4.93 66.215 7.035 ;
        RECT 63.03 5.43 65.78 7.04 ;
        RECT 64.125 4.93 64.295 7.04 ;
        RECT 63.2 5.43 63.37 7.77 ;
        RECT 63.185 4.93 63.355 7.04 ;
        RECT 61.725 4.93 61.895 7.035 ;
        RECT 59.805 4.93 59.975 7.035 ;
        RECT 43.755 5.43 58.265 7.035 ;
        RECT 53.385 5.43 58.11 7.04 ;
        RECT 53.385 5.425 58.105 7.04 ;
        RECT 57.29 5.425 57.46 7.77 ;
        RECT 57.285 4.695 57.455 7.04 ;
        RECT 56.3 4.695 56.47 7.77 ;
        RECT 53.555 4.695 53.725 7.77 ;
        RECT 50.785 4.93 50.955 7.035 ;
        RECT 47.77 5.43 50.52 7.04 ;
        RECT 48.865 4.93 49.035 7.04 ;
        RECT 47.94 5.43 48.11 7.77 ;
        RECT 47.925 4.93 48.095 7.04 ;
        RECT 46.465 4.93 46.635 7.035 ;
        RECT 44.545 4.93 44.715 7.035 ;
        RECT 28.495 5.43 43.005 7.035 ;
        RECT 38.125 5.43 42.85 7.04 ;
        RECT 38.125 5.425 42.845 7.04 ;
        RECT 42.03 5.425 42.2 7.77 ;
        RECT 42.025 4.695 42.195 7.04 ;
        RECT 41.04 4.695 41.21 7.77 ;
        RECT 38.295 4.695 38.465 7.77 ;
        RECT 35.525 4.93 35.695 7.035 ;
        RECT 32.51 5.43 35.26 7.04 ;
        RECT 33.605 4.93 33.775 7.04 ;
        RECT 32.68 5.43 32.85 7.77 ;
        RECT 32.665 4.93 32.835 7.04 ;
        RECT 31.205 4.93 31.375 7.035 ;
        RECT 29.285 4.93 29.455 7.035 ;
        RECT 24.995 5.435 27.745 7.04 ;
        RECT 26.98 10.05 27.155 10.6 ;
        RECT 26.98 7.31 27.155 8.45 ;
        RECT 26.98 5.435 27.15 10.6 ;
        RECT 25.165 5.435 25.335 7.77 ;
      LAYER met1 ;
        RECT 0 5.435 104.045 7.035 ;
        RECT 89.535 5.43 104.045 7.035 ;
        RECT 99.165 5.43 103.89 7.04 ;
        RECT 99.165 5.425 103.885 7.04 ;
        RECT 89.535 5.4 98.275 7.035 ;
        RECT 93.55 5.4 96.3 7.04 ;
        RECT 74.275 5.43 88.785 7.035 ;
        RECT 83.905 5.43 88.63 7.04 ;
        RECT 83.905 5.425 88.625 7.04 ;
        RECT 74.275 5.4 83.015 7.035 ;
        RECT 78.29 5.4 81.04 7.04 ;
        RECT 59.015 5.43 73.525 7.035 ;
        RECT 68.645 5.43 73.37 7.04 ;
        RECT 68.645 5.425 73.365 7.04 ;
        RECT 59.015 5.4 67.755 7.035 ;
        RECT 63.03 5.4 65.78 7.04 ;
        RECT 43.755 5.43 58.265 7.035 ;
        RECT 53.385 5.43 58.11 7.04 ;
        RECT 53.385 5.425 58.105 7.04 ;
        RECT 43.755 5.4 52.495 7.035 ;
        RECT 47.77 5.4 50.52 7.04 ;
        RECT 28.495 5.43 43.005 7.035 ;
        RECT 38.125 5.43 42.85 7.04 ;
        RECT 38.125 5.425 42.845 7.04 ;
        RECT 28.495 5.4 37.235 7.035 ;
        RECT 32.51 5.4 35.26 7.04 ;
        RECT 24.995 5.435 27.745 7.04 ;
        RECT 26.92 8.95 27.21 9.18 ;
        RECT 26.75 8.98 27.21 9.15 ;
      LAYER mcon ;
        RECT 26.98 8.98 27.15 9.15 ;
        RECT 27.285 6.84 27.455 7.01 ;
        RECT 28.64 5.43 28.81 5.6 ;
        RECT 29.1 5.43 29.27 5.6 ;
        RECT 29.56 5.43 29.73 5.6 ;
        RECT 30.02 5.43 30.19 5.6 ;
        RECT 30.48 5.43 30.65 5.6 ;
        RECT 30.94 5.43 31.11 5.6 ;
        RECT 31.4 5.43 31.57 5.6 ;
        RECT 31.86 5.43 32.03 5.6 ;
        RECT 32.32 5.43 32.49 5.6 ;
        RECT 32.78 5.43 32.95 5.6 ;
        RECT 33.24 5.43 33.41 5.6 ;
        RECT 33.7 5.43 33.87 5.6 ;
        RECT 34.16 5.43 34.33 5.6 ;
        RECT 34.62 5.43 34.79 5.6 ;
        RECT 34.8 6.84 34.97 7.01 ;
        RECT 35.08 5.43 35.25 5.6 ;
        RECT 35.54 5.43 35.71 5.6 ;
        RECT 36 5.43 36.17 5.6 ;
        RECT 36.46 5.43 36.63 5.6 ;
        RECT 36.92 5.43 37.09 5.6 ;
        RECT 40.415 6.84 40.585 7.01 ;
        RECT 40.415 5.455 40.585 5.625 ;
        RECT 41.12 6.84 41.29 7.01 ;
        RECT 41.12 5.455 41.29 5.625 ;
        RECT 42.105 5.455 42.275 5.625 ;
        RECT 42.11 6.84 42.28 7.01 ;
        RECT 43.9 5.43 44.07 5.6 ;
        RECT 44.36 5.43 44.53 5.6 ;
        RECT 44.82 5.43 44.99 5.6 ;
        RECT 45.28 5.43 45.45 5.6 ;
        RECT 45.74 5.43 45.91 5.6 ;
        RECT 46.2 5.43 46.37 5.6 ;
        RECT 46.66 5.43 46.83 5.6 ;
        RECT 47.12 5.43 47.29 5.6 ;
        RECT 47.58 5.43 47.75 5.6 ;
        RECT 48.04 5.43 48.21 5.6 ;
        RECT 48.5 5.43 48.67 5.6 ;
        RECT 48.96 5.43 49.13 5.6 ;
        RECT 49.42 5.43 49.59 5.6 ;
        RECT 49.88 5.43 50.05 5.6 ;
        RECT 50.06 6.84 50.23 7.01 ;
        RECT 50.34 5.43 50.51 5.6 ;
        RECT 50.8 5.43 50.97 5.6 ;
        RECT 51.26 5.43 51.43 5.6 ;
        RECT 51.72 5.43 51.89 5.6 ;
        RECT 52.18 5.43 52.35 5.6 ;
        RECT 55.675 6.84 55.845 7.01 ;
        RECT 55.675 5.455 55.845 5.625 ;
        RECT 56.38 6.84 56.55 7.01 ;
        RECT 56.38 5.455 56.55 5.625 ;
        RECT 57.365 5.455 57.535 5.625 ;
        RECT 57.37 6.84 57.54 7.01 ;
        RECT 59.16 5.43 59.33 5.6 ;
        RECT 59.62 5.43 59.79 5.6 ;
        RECT 60.08 5.43 60.25 5.6 ;
        RECT 60.54 5.43 60.71 5.6 ;
        RECT 61 5.43 61.17 5.6 ;
        RECT 61.46 5.43 61.63 5.6 ;
        RECT 61.92 5.43 62.09 5.6 ;
        RECT 62.38 5.43 62.55 5.6 ;
        RECT 62.84 5.43 63.01 5.6 ;
        RECT 63.3 5.43 63.47 5.6 ;
        RECT 63.76 5.43 63.93 5.6 ;
        RECT 64.22 5.43 64.39 5.6 ;
        RECT 64.68 5.43 64.85 5.6 ;
        RECT 65.14 5.43 65.31 5.6 ;
        RECT 65.32 6.84 65.49 7.01 ;
        RECT 65.6 5.43 65.77 5.6 ;
        RECT 66.06 5.43 66.23 5.6 ;
        RECT 66.52 5.43 66.69 5.6 ;
        RECT 66.98 5.43 67.15 5.6 ;
        RECT 67.44 5.43 67.61 5.6 ;
        RECT 70.935 6.84 71.105 7.01 ;
        RECT 70.935 5.455 71.105 5.625 ;
        RECT 71.64 6.84 71.81 7.01 ;
        RECT 71.64 5.455 71.81 5.625 ;
        RECT 72.625 5.455 72.795 5.625 ;
        RECT 72.63 6.84 72.8 7.01 ;
        RECT 74.42 5.43 74.59 5.6 ;
        RECT 74.88 5.43 75.05 5.6 ;
        RECT 75.34 5.43 75.51 5.6 ;
        RECT 75.8 5.43 75.97 5.6 ;
        RECT 76.26 5.43 76.43 5.6 ;
        RECT 76.72 5.43 76.89 5.6 ;
        RECT 77.18 5.43 77.35 5.6 ;
        RECT 77.64 5.43 77.81 5.6 ;
        RECT 78.1 5.43 78.27 5.6 ;
        RECT 78.56 5.43 78.73 5.6 ;
        RECT 79.02 5.43 79.19 5.6 ;
        RECT 79.48 5.43 79.65 5.6 ;
        RECT 79.94 5.43 80.11 5.6 ;
        RECT 80.4 5.43 80.57 5.6 ;
        RECT 80.58 6.84 80.75 7.01 ;
        RECT 80.86 5.43 81.03 5.6 ;
        RECT 81.32 5.43 81.49 5.6 ;
        RECT 81.78 5.43 81.95 5.6 ;
        RECT 82.24 5.43 82.41 5.6 ;
        RECT 82.7 5.43 82.87 5.6 ;
        RECT 86.195 6.84 86.365 7.01 ;
        RECT 86.195 5.455 86.365 5.625 ;
        RECT 86.9 6.84 87.07 7.01 ;
        RECT 86.9 5.455 87.07 5.625 ;
        RECT 87.885 5.455 88.055 5.625 ;
        RECT 87.89 6.84 88.06 7.01 ;
        RECT 89.68 5.43 89.85 5.6 ;
        RECT 90.14 5.43 90.31 5.6 ;
        RECT 90.6 5.43 90.77 5.6 ;
        RECT 91.06 5.43 91.23 5.6 ;
        RECT 91.52 5.43 91.69 5.6 ;
        RECT 91.98 5.43 92.15 5.6 ;
        RECT 92.44 5.43 92.61 5.6 ;
        RECT 92.9 5.43 93.07 5.6 ;
        RECT 93.36 5.43 93.53 5.6 ;
        RECT 93.82 5.43 93.99 5.6 ;
        RECT 94.28 5.43 94.45 5.6 ;
        RECT 94.74 5.43 94.91 5.6 ;
        RECT 95.2 5.43 95.37 5.6 ;
        RECT 95.66 5.43 95.83 5.6 ;
        RECT 95.84 6.84 96.01 7.01 ;
        RECT 96.12 5.43 96.29 5.6 ;
        RECT 96.58 5.43 96.75 5.6 ;
        RECT 97.04 5.43 97.21 5.6 ;
        RECT 97.5 5.43 97.67 5.6 ;
        RECT 97.96 5.43 98.13 5.6 ;
        RECT 101.455 6.84 101.625 7.01 ;
        RECT 101.455 5.455 101.625 5.625 ;
        RECT 102.16 6.84 102.33 7.01 ;
        RECT 102.16 5.455 102.33 5.625 ;
        RECT 103.145 5.455 103.315 5.625 ;
        RECT 103.15 6.84 103.32 7.01 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 90.365 3.15 91.095 3.48 ;
        RECT 75.105 3.15 75.835 3.48 ;
        RECT 59.845 3.15 60.575 3.48 ;
        RECT 44.585 3.15 45.315 3.48 ;
        RECT 29.325 3.15 30.055 3.48 ;
      LAYER met2 ;
        RECT 90.51 3.155 90.9 3.475 ;
        RECT 90.51 3.13 90.79 3.5 ;
        RECT 75.25 3.155 75.64 3.475 ;
        RECT 75.25 3.13 75.53 3.5 ;
        RECT 59.99 3.155 60.38 3.475 ;
        RECT 59.99 3.13 60.27 3.5 ;
        RECT 44.73 3.155 45.12 3.475 ;
        RECT 44.73 3.13 45.01 3.5 ;
        RECT 29.47 3.155 29.86 3.475 ;
        RECT 29.47 3.13 29.75 3.5 ;
      LAYER li1 ;
        RECT 0 0 104.045 1.6 ;
        RECT 103.065 0 103.235 2.225 ;
        RECT 102.08 0 102.25 2.225 ;
        RECT 99.335 0 99.505 2.225 ;
        RECT 89.535 0 98.275 2.88 ;
        RECT 97.505 0 97.675 3.38 ;
        RECT 96.565 0 96.735 3.38 ;
        RECT 95.605 0 95.775 3.38 ;
        RECT 94.56 0 94.755 2.89 ;
        RECT 93.685 0 93.855 3.38 ;
        RECT 92.725 0 92.895 3.38 ;
        RECT 90.805 0 91.08 2.89 ;
        RECT 90.805 0 90.975 3.38 ;
        RECT 87.805 0 87.975 2.225 ;
        RECT 86.82 0 86.99 2.225 ;
        RECT 84.075 0 84.245 2.225 ;
        RECT 74.275 0 83.015 2.88 ;
        RECT 82.245 0 82.415 3.38 ;
        RECT 81.305 0 81.475 3.38 ;
        RECT 80.345 0 80.515 3.38 ;
        RECT 79.3 0 79.495 2.89 ;
        RECT 78.425 0 78.595 3.38 ;
        RECT 77.465 0 77.635 3.38 ;
        RECT 75.545 0 75.82 2.89 ;
        RECT 75.545 0 75.715 3.38 ;
        RECT 72.545 0 72.715 2.225 ;
        RECT 71.56 0 71.73 2.225 ;
        RECT 68.815 0 68.985 2.225 ;
        RECT 59.015 0 67.755 2.88 ;
        RECT 66.985 0 67.155 3.38 ;
        RECT 66.045 0 66.215 3.38 ;
        RECT 65.085 0 65.255 3.38 ;
        RECT 64.04 0 64.235 2.89 ;
        RECT 63.165 0 63.335 3.38 ;
        RECT 62.205 0 62.375 3.38 ;
        RECT 60.285 0 60.56 2.89 ;
        RECT 60.285 0 60.455 3.38 ;
        RECT 57.285 0 57.455 2.225 ;
        RECT 56.3 0 56.47 2.225 ;
        RECT 53.555 0 53.725 2.225 ;
        RECT 43.755 0 52.495 2.88 ;
        RECT 51.725 0 51.895 3.38 ;
        RECT 50.785 0 50.955 3.38 ;
        RECT 49.825 0 49.995 3.38 ;
        RECT 48.78 0 48.975 2.89 ;
        RECT 47.905 0 48.075 3.38 ;
        RECT 46.945 0 47.115 3.38 ;
        RECT 45.025 0 45.3 2.89 ;
        RECT 45.025 0 45.195 3.38 ;
        RECT 42.025 0 42.195 2.225 ;
        RECT 41.04 0 41.21 2.225 ;
        RECT 38.295 0 38.465 2.225 ;
        RECT 28.495 0 37.235 2.88 ;
        RECT 36.465 0 36.635 3.38 ;
        RECT 35.525 0 35.695 3.38 ;
        RECT 34.565 0 34.735 3.38 ;
        RECT 33.52 0 33.715 2.89 ;
        RECT 32.645 0 32.815 3.38 ;
        RECT 31.685 0 31.855 3.38 ;
        RECT 29.765 0 30.04 2.89 ;
        RECT 29.765 0 29.935 3.38 ;
        RECT 0 10.865 104.045 12.465 ;
        RECT 103.07 10.24 103.24 12.465 ;
        RECT 102.08 10.24 102.25 12.465 ;
        RECT 99.335 10.24 99.505 12.465 ;
        RECT 93.72 10.24 93.89 12.465 ;
        RECT 87.81 10.24 87.98 12.465 ;
        RECT 86.82 10.24 86.99 12.465 ;
        RECT 84.075 10.24 84.245 12.465 ;
        RECT 78.46 10.24 78.63 12.465 ;
        RECT 72.55 10.24 72.72 12.465 ;
        RECT 71.56 10.24 71.73 12.465 ;
        RECT 68.815 10.24 68.985 12.465 ;
        RECT 63.2 10.24 63.37 12.465 ;
        RECT 57.29 10.24 57.46 12.465 ;
        RECT 56.3 10.24 56.47 12.465 ;
        RECT 53.555 10.24 53.725 12.465 ;
        RECT 47.94 10.24 48.11 12.465 ;
        RECT 42.03 10.24 42.2 12.465 ;
        RECT 41.04 10.24 41.21 12.465 ;
        RECT 38.295 10.24 38.465 12.465 ;
        RECT 32.68 10.24 32.85 12.465 ;
        RECT 25.165 10.24 25.335 12.465 ;
        RECT 94.735 8.37 94.905 10.32 ;
        RECT 94.675 10.15 94.845 10.6 ;
        RECT 94.675 7.31 94.845 8.54 ;
        RECT 91.405 3.87 91.775 4.04 ;
        RECT 91.405 3.23 91.575 4.04 ;
        RECT 91.285 3.23 91.575 3.4 ;
        RECT 90.085 3.79 90.255 4.24 ;
        RECT 79.475 8.37 79.645 10.32 ;
        RECT 79.415 10.15 79.585 10.6 ;
        RECT 79.415 7.31 79.585 8.54 ;
        RECT 76.145 3.87 76.515 4.04 ;
        RECT 76.145 3.23 76.315 4.04 ;
        RECT 76.025 3.23 76.315 3.4 ;
        RECT 74.825 3.79 74.995 4.24 ;
        RECT 64.215 8.37 64.385 10.32 ;
        RECT 64.155 10.15 64.325 10.6 ;
        RECT 64.155 7.31 64.325 8.54 ;
        RECT 60.885 3.87 61.255 4.04 ;
        RECT 60.885 3.23 61.055 4.04 ;
        RECT 60.765 3.23 61.055 3.4 ;
        RECT 59.565 3.79 59.735 4.24 ;
        RECT 48.955 8.37 49.125 10.32 ;
        RECT 48.895 10.15 49.065 10.6 ;
        RECT 48.895 7.31 49.065 8.54 ;
        RECT 45.625 3.87 45.995 4.04 ;
        RECT 45.625 3.23 45.795 4.04 ;
        RECT 45.505 3.23 45.795 3.4 ;
        RECT 44.305 3.79 44.475 4.24 ;
        RECT 33.695 8.37 33.865 10.32 ;
        RECT 33.635 10.15 33.805 10.6 ;
        RECT 33.635 7.31 33.805 8.54 ;
        RECT 30.365 3.87 30.735 4.04 ;
        RECT 30.365 3.23 30.535 4.04 ;
        RECT 30.245 3.23 30.535 3.4 ;
        RECT 29.045 3.79 29.215 4.24 ;
      LAYER met1 ;
        RECT 0 0 104.045 1.6 ;
        RECT 98.08 0 98.275 2.92 ;
        RECT 89.535 0 98.275 2.915 ;
        RECT 91.225 3.2 91.515 3.43 ;
        RECT 90.34 3.245 91.515 3.385 ;
        RECT 90.52 3.185 90.93 3.445 ;
        RECT 90.52 0 90.81 3.445 ;
        RECT 90.1 3.665 90.72 3.805 ;
        RECT 90.58 0 90.72 3.805 ;
        RECT 90.34 3.245 90.72 3.505 ;
        RECT 90.025 4.04 90.315 4.27 ;
        RECT 90.1 3.665 90.24 4.27 ;
        RECT 82.82 0 83.015 2.92 ;
        RECT 74.275 0 83.015 2.915 ;
        RECT 75.965 3.2 76.255 3.43 ;
        RECT 75.08 3.245 76.255 3.385 ;
        RECT 75.26 3.185 75.67 3.445 ;
        RECT 75.26 0 75.55 3.445 ;
        RECT 74.84 3.665 75.46 3.805 ;
        RECT 75.32 0 75.46 3.805 ;
        RECT 75.08 3.245 75.46 3.505 ;
        RECT 74.765 4.04 75.055 4.27 ;
        RECT 74.84 3.665 74.98 4.27 ;
        RECT 67.56 0 67.755 2.92 ;
        RECT 59.015 0 67.755 2.915 ;
        RECT 60.705 3.2 60.995 3.43 ;
        RECT 59.82 3.245 60.995 3.385 ;
        RECT 60 3.185 60.41 3.445 ;
        RECT 60 0 60.29 3.445 ;
        RECT 59.58 3.665 60.2 3.805 ;
        RECT 60.06 0 60.2 3.805 ;
        RECT 59.82 3.245 60.2 3.505 ;
        RECT 59.505 4.04 59.795 4.27 ;
        RECT 59.58 3.665 59.72 4.27 ;
        RECT 52.3 0 52.495 2.92 ;
        RECT 43.755 0 52.495 2.915 ;
        RECT 45.445 3.2 45.735 3.43 ;
        RECT 44.56 3.245 45.735 3.385 ;
        RECT 44.74 3.185 45.15 3.445 ;
        RECT 44.74 0 45.03 3.445 ;
        RECT 44.32 3.665 44.94 3.805 ;
        RECT 44.8 0 44.94 3.805 ;
        RECT 44.56 3.245 44.94 3.505 ;
        RECT 44.245 4.04 44.535 4.27 ;
        RECT 44.32 3.665 44.46 4.27 ;
        RECT 37.04 0 37.235 2.92 ;
        RECT 28.495 0 37.235 2.915 ;
        RECT 30.185 3.2 30.475 3.43 ;
        RECT 29.3 3.245 30.475 3.385 ;
        RECT 29.48 3.185 29.89 3.445 ;
        RECT 29.48 0 29.77 3.445 ;
        RECT 29.06 3.665 29.68 3.805 ;
        RECT 29.54 0 29.68 3.805 ;
        RECT 29.3 3.245 29.68 3.505 ;
        RECT 28.985 4.04 29.275 4.27 ;
        RECT 29.06 3.665 29.2 4.27 ;
        RECT 0 10.865 104.045 12.465 ;
        RECT 94.675 8.58 94.965 8.81 ;
        RECT 94.505 8.605 94.675 12.465 ;
        RECT 94.5 8.61 94.965 8.78 ;
        RECT 79.415 8.58 79.705 8.81 ;
        RECT 79.245 8.605 79.415 12.465 ;
        RECT 79.24 8.61 79.705 8.78 ;
        RECT 64.155 8.58 64.445 8.81 ;
        RECT 63.985 8.605 64.155 12.465 ;
        RECT 63.98 8.61 64.445 8.78 ;
        RECT 48.895 8.58 49.185 8.81 ;
        RECT 48.725 8.605 48.895 12.465 ;
        RECT 48.72 8.61 49.185 8.78 ;
        RECT 33.635 8.58 33.925 8.81 ;
        RECT 33.465 8.605 33.635 12.465 ;
        RECT 33.46 8.61 33.925 8.78 ;
      LAYER via1 ;
        RECT 29.655 3.24 29.805 3.39 ;
        RECT 44.915 3.24 45.065 3.39 ;
        RECT 60.175 3.24 60.325 3.39 ;
        RECT 75.435 3.24 75.585 3.39 ;
        RECT 90.695 3.24 90.845 3.39 ;
      LAYER via2 ;
        RECT 29.51 3.215 29.71 3.415 ;
        RECT 44.77 3.215 44.97 3.415 ;
        RECT 60.03 3.215 60.23 3.415 ;
        RECT 75.29 3.215 75.49 3.415 ;
        RECT 90.55 3.215 90.75 3.415 ;
      LAYER mcon ;
        RECT 25.245 10.9 25.415 11.07 ;
        RECT 25.925 10.9 26.095 11.07 ;
        RECT 26.605 10.9 26.775 11.07 ;
        RECT 27.285 10.9 27.455 11.07 ;
        RECT 28.64 2.71 28.81 2.88 ;
        RECT 29.045 4.07 29.215 4.24 ;
        RECT 29.1 2.71 29.27 2.88 ;
        RECT 29.56 2.71 29.73 2.88 ;
        RECT 30.02 2.71 30.19 2.88 ;
        RECT 30.245 3.23 30.415 3.4 ;
        RECT 30.48 2.71 30.65 2.88 ;
        RECT 30.94 2.71 31.11 2.88 ;
        RECT 31.4 2.71 31.57 2.88 ;
        RECT 31.86 2.71 32.03 2.88 ;
        RECT 32.32 2.71 32.49 2.88 ;
        RECT 32.76 10.9 32.93 11.07 ;
        RECT 32.78 2.71 32.95 2.88 ;
        RECT 33.24 2.71 33.41 2.88 ;
        RECT 33.44 10.9 33.61 11.07 ;
        RECT 33.695 8.61 33.865 8.78 ;
        RECT 33.7 2.71 33.87 2.88 ;
        RECT 34.12 10.9 34.29 11.07 ;
        RECT 34.16 2.71 34.33 2.88 ;
        RECT 34.62 2.71 34.79 2.88 ;
        RECT 34.8 10.9 34.97 11.07 ;
        RECT 35.08 2.71 35.25 2.88 ;
        RECT 35.54 2.71 35.71 2.88 ;
        RECT 36 2.71 36.17 2.88 ;
        RECT 36.46 2.71 36.63 2.88 ;
        RECT 36.92 2.71 37.09 2.88 ;
        RECT 38.375 10.9 38.545 11.07 ;
        RECT 38.375 1.395 38.545 1.565 ;
        RECT 39.055 10.9 39.225 11.07 ;
        RECT 39.055 1.395 39.225 1.565 ;
        RECT 39.735 10.9 39.905 11.07 ;
        RECT 39.735 1.395 39.905 1.565 ;
        RECT 40.415 10.9 40.585 11.07 ;
        RECT 40.415 1.395 40.585 1.565 ;
        RECT 41.12 10.9 41.29 11.07 ;
        RECT 41.12 1.395 41.29 1.565 ;
        RECT 42.105 1.395 42.275 1.565 ;
        RECT 42.11 10.9 42.28 11.07 ;
        RECT 43.9 2.71 44.07 2.88 ;
        RECT 44.305 4.07 44.475 4.24 ;
        RECT 44.36 2.71 44.53 2.88 ;
        RECT 44.82 2.71 44.99 2.88 ;
        RECT 45.28 2.71 45.45 2.88 ;
        RECT 45.505 3.23 45.675 3.4 ;
        RECT 45.74 2.71 45.91 2.88 ;
        RECT 46.2 2.71 46.37 2.88 ;
        RECT 46.66 2.71 46.83 2.88 ;
        RECT 47.12 2.71 47.29 2.88 ;
        RECT 47.58 2.71 47.75 2.88 ;
        RECT 48.02 10.9 48.19 11.07 ;
        RECT 48.04 2.71 48.21 2.88 ;
        RECT 48.5 2.71 48.67 2.88 ;
        RECT 48.7 10.9 48.87 11.07 ;
        RECT 48.955 8.61 49.125 8.78 ;
        RECT 48.96 2.71 49.13 2.88 ;
        RECT 49.38 10.9 49.55 11.07 ;
        RECT 49.42 2.71 49.59 2.88 ;
        RECT 49.88 2.71 50.05 2.88 ;
        RECT 50.06 10.9 50.23 11.07 ;
        RECT 50.34 2.71 50.51 2.88 ;
        RECT 50.8 2.71 50.97 2.88 ;
        RECT 51.26 2.71 51.43 2.88 ;
        RECT 51.72 2.71 51.89 2.88 ;
        RECT 52.18 2.71 52.35 2.88 ;
        RECT 53.635 10.9 53.805 11.07 ;
        RECT 53.635 1.395 53.805 1.565 ;
        RECT 54.315 10.9 54.485 11.07 ;
        RECT 54.315 1.395 54.485 1.565 ;
        RECT 54.995 10.9 55.165 11.07 ;
        RECT 54.995 1.395 55.165 1.565 ;
        RECT 55.675 10.9 55.845 11.07 ;
        RECT 55.675 1.395 55.845 1.565 ;
        RECT 56.38 10.9 56.55 11.07 ;
        RECT 56.38 1.395 56.55 1.565 ;
        RECT 57.365 1.395 57.535 1.565 ;
        RECT 57.37 10.9 57.54 11.07 ;
        RECT 59.16 2.71 59.33 2.88 ;
        RECT 59.565 4.07 59.735 4.24 ;
        RECT 59.62 2.71 59.79 2.88 ;
        RECT 60.08 2.71 60.25 2.88 ;
        RECT 60.54 2.71 60.71 2.88 ;
        RECT 60.765 3.23 60.935 3.4 ;
        RECT 61 2.71 61.17 2.88 ;
        RECT 61.46 2.71 61.63 2.88 ;
        RECT 61.92 2.71 62.09 2.88 ;
        RECT 62.38 2.71 62.55 2.88 ;
        RECT 62.84 2.71 63.01 2.88 ;
        RECT 63.28 10.9 63.45 11.07 ;
        RECT 63.3 2.71 63.47 2.88 ;
        RECT 63.76 2.71 63.93 2.88 ;
        RECT 63.96 10.9 64.13 11.07 ;
        RECT 64.215 8.61 64.385 8.78 ;
        RECT 64.22 2.71 64.39 2.88 ;
        RECT 64.64 10.9 64.81 11.07 ;
        RECT 64.68 2.71 64.85 2.88 ;
        RECT 65.14 2.71 65.31 2.88 ;
        RECT 65.32 10.9 65.49 11.07 ;
        RECT 65.6 2.71 65.77 2.88 ;
        RECT 66.06 2.71 66.23 2.88 ;
        RECT 66.52 2.71 66.69 2.88 ;
        RECT 66.98 2.71 67.15 2.88 ;
        RECT 67.44 2.71 67.61 2.88 ;
        RECT 68.895 10.9 69.065 11.07 ;
        RECT 68.895 1.395 69.065 1.565 ;
        RECT 69.575 10.9 69.745 11.07 ;
        RECT 69.575 1.395 69.745 1.565 ;
        RECT 70.255 10.9 70.425 11.07 ;
        RECT 70.255 1.395 70.425 1.565 ;
        RECT 70.935 10.9 71.105 11.07 ;
        RECT 70.935 1.395 71.105 1.565 ;
        RECT 71.64 10.9 71.81 11.07 ;
        RECT 71.64 1.395 71.81 1.565 ;
        RECT 72.625 1.395 72.795 1.565 ;
        RECT 72.63 10.9 72.8 11.07 ;
        RECT 74.42 2.71 74.59 2.88 ;
        RECT 74.825 4.07 74.995 4.24 ;
        RECT 74.88 2.71 75.05 2.88 ;
        RECT 75.34 2.71 75.51 2.88 ;
        RECT 75.8 2.71 75.97 2.88 ;
        RECT 76.025 3.23 76.195 3.4 ;
        RECT 76.26 2.71 76.43 2.88 ;
        RECT 76.72 2.71 76.89 2.88 ;
        RECT 77.18 2.71 77.35 2.88 ;
        RECT 77.64 2.71 77.81 2.88 ;
        RECT 78.1 2.71 78.27 2.88 ;
        RECT 78.54 10.9 78.71 11.07 ;
        RECT 78.56 2.71 78.73 2.88 ;
        RECT 79.02 2.71 79.19 2.88 ;
        RECT 79.22 10.9 79.39 11.07 ;
        RECT 79.475 8.61 79.645 8.78 ;
        RECT 79.48 2.71 79.65 2.88 ;
        RECT 79.9 10.9 80.07 11.07 ;
        RECT 79.94 2.71 80.11 2.88 ;
        RECT 80.4 2.71 80.57 2.88 ;
        RECT 80.58 10.9 80.75 11.07 ;
        RECT 80.86 2.71 81.03 2.88 ;
        RECT 81.32 2.71 81.49 2.88 ;
        RECT 81.78 2.71 81.95 2.88 ;
        RECT 82.24 2.71 82.41 2.88 ;
        RECT 82.7 2.71 82.87 2.88 ;
        RECT 84.155 10.9 84.325 11.07 ;
        RECT 84.155 1.395 84.325 1.565 ;
        RECT 84.835 10.9 85.005 11.07 ;
        RECT 84.835 1.395 85.005 1.565 ;
        RECT 85.515 10.9 85.685 11.07 ;
        RECT 85.515 1.395 85.685 1.565 ;
        RECT 86.195 10.9 86.365 11.07 ;
        RECT 86.195 1.395 86.365 1.565 ;
        RECT 86.9 10.9 87.07 11.07 ;
        RECT 86.9 1.395 87.07 1.565 ;
        RECT 87.885 1.395 88.055 1.565 ;
        RECT 87.89 10.9 88.06 11.07 ;
        RECT 89.68 2.71 89.85 2.88 ;
        RECT 90.085 4.07 90.255 4.24 ;
        RECT 90.14 2.71 90.31 2.88 ;
        RECT 90.6 2.71 90.77 2.88 ;
        RECT 91.06 2.71 91.23 2.88 ;
        RECT 91.285 3.23 91.455 3.4 ;
        RECT 91.52 2.71 91.69 2.88 ;
        RECT 91.98 2.71 92.15 2.88 ;
        RECT 92.44 2.71 92.61 2.88 ;
        RECT 92.9 2.71 93.07 2.88 ;
        RECT 93.36 2.71 93.53 2.88 ;
        RECT 93.8 10.9 93.97 11.07 ;
        RECT 93.82 2.71 93.99 2.88 ;
        RECT 94.28 2.71 94.45 2.88 ;
        RECT 94.48 10.9 94.65 11.07 ;
        RECT 94.735 8.61 94.905 8.78 ;
        RECT 94.74 2.71 94.91 2.88 ;
        RECT 95.16 10.9 95.33 11.07 ;
        RECT 95.2 2.71 95.37 2.88 ;
        RECT 95.66 2.71 95.83 2.88 ;
        RECT 95.84 10.9 96.01 11.07 ;
        RECT 96.12 2.71 96.29 2.88 ;
        RECT 96.58 2.71 96.75 2.88 ;
        RECT 97.04 2.71 97.21 2.88 ;
        RECT 97.5 2.71 97.67 2.88 ;
        RECT 97.96 2.71 98.13 2.88 ;
        RECT 99.415 10.9 99.585 11.07 ;
        RECT 99.415 1.395 99.585 1.565 ;
        RECT 100.095 10.9 100.265 11.07 ;
        RECT 100.095 1.395 100.265 1.565 ;
        RECT 100.775 10.9 100.945 11.07 ;
        RECT 100.775 1.395 100.945 1.565 ;
        RECT 101.455 10.9 101.625 11.07 ;
        RECT 101.455 1.395 101.625 1.565 ;
        RECT 102.16 10.9 102.33 11.07 ;
        RECT 102.16 1.395 102.33 1.565 ;
        RECT 103.145 1.395 103.315 1.565 ;
        RECT 103.15 10.9 103.32 11.07 ;
    END
  END vssd1
  OBS
    LAYER met4 ;
      RECT 91.685 4.27 92.015 4.6 ;
      RECT 91.7 3.795 92.015 4.6 ;
      RECT 93.845 3.78 94.175 4.135 ;
      RECT 91.7 3.795 94.175 4.095 ;
      RECT 76.425 4.27 76.755 4.6 ;
      RECT 76.44 3.795 76.755 4.6 ;
      RECT 78.585 3.78 78.915 4.135 ;
      RECT 76.44 3.795 78.915 4.095 ;
      RECT 61.165 4.27 61.495 4.6 ;
      RECT 61.18 3.795 61.495 4.6 ;
      RECT 63.325 3.78 63.655 4.135 ;
      RECT 61.18 3.795 63.655 4.095 ;
      RECT 45.905 4.27 46.235 4.6 ;
      RECT 45.92 3.795 46.235 4.6 ;
      RECT 48.065 3.78 48.395 4.135 ;
      RECT 45.92 3.795 48.395 4.095 ;
      RECT 30.645 4.27 30.975 4.6 ;
      RECT 30.66 3.795 30.975 4.6 ;
      RECT 32.805 3.78 33.135 4.135 ;
      RECT 30.66 3.795 33.135 4.095 ;
    LAYER via3 ;
      RECT 93.91 3.87 94.11 4.07 ;
      RECT 91.75 4.335 91.95 4.535 ;
      RECT 78.65 3.87 78.85 4.07 ;
      RECT 76.49 4.335 76.69 4.535 ;
      RECT 63.39 3.87 63.59 4.07 ;
      RECT 61.23 4.335 61.43 4.535 ;
      RECT 48.13 3.87 48.33 4.07 ;
      RECT 45.97 4.335 46.17 4.535 ;
      RECT 32.87 3.87 33.07 4.07 ;
      RECT 30.71 4.335 30.91 4.535 ;
    LAYER met3 ;
      RECT 95.005 9.345 95.375 9.715 ;
      RECT 95.04 6.175 95.34 9.715 ;
      RECT 95.035 5.47 95.335 6.53 ;
      RECT 90.805 5.47 95.335 5.77 ;
      RECT 93.6 3.81 93.9 5.77 ;
      RECT 90.805 4.27 91.105 5.77 ;
      RECT 94.325 4.805 94.655 5.16 ;
      RECT 92.42 4.845 94.655 5.145 ;
      RECT 92.42 3.71 92.72 5.145 ;
      RECT 90.5 4.27 91.23 4.6 ;
      RECT 93.395 3.815 94.175 4.16 ;
      RECT 93.85 3.78 94.175 4.16 ;
      RECT 92.405 3.71 92.735 4.04 ;
      RECT 91.69 3.71 92.01 4.625 ;
      RECT 91.69 3.71 92.02 4.245 ;
      RECT 79.745 9.345 80.115 9.715 ;
      RECT 79.78 6.175 80.08 9.715 ;
      RECT 79.775 5.47 80.075 6.53 ;
      RECT 75.545 5.47 80.075 5.77 ;
      RECT 78.34 3.81 78.64 5.77 ;
      RECT 75.545 4.27 75.845 5.77 ;
      RECT 79.065 4.805 79.395 5.16 ;
      RECT 77.16 4.845 79.395 5.145 ;
      RECT 77.16 3.71 77.46 5.145 ;
      RECT 75.24 4.27 75.97 4.6 ;
      RECT 78.135 3.815 78.915 4.16 ;
      RECT 78.59 3.78 78.915 4.16 ;
      RECT 77.145 3.71 77.475 4.04 ;
      RECT 76.43 3.71 76.75 4.625 ;
      RECT 76.43 3.71 76.76 4.245 ;
      RECT 64.485 9.345 64.855 9.715 ;
      RECT 64.52 6.175 64.82 9.715 ;
      RECT 64.515 5.47 64.815 6.53 ;
      RECT 60.285 5.47 64.815 5.77 ;
      RECT 63.08 3.81 63.38 5.77 ;
      RECT 60.285 4.27 60.585 5.77 ;
      RECT 63.805 4.805 64.135 5.16 ;
      RECT 61.9 4.845 64.135 5.145 ;
      RECT 61.9 3.71 62.2 5.145 ;
      RECT 59.98 4.27 60.71 4.6 ;
      RECT 62.875 3.815 63.655 4.16 ;
      RECT 63.33 3.78 63.655 4.16 ;
      RECT 61.885 3.71 62.215 4.04 ;
      RECT 61.17 3.71 61.49 4.625 ;
      RECT 61.17 3.71 61.5 4.245 ;
      RECT 49.225 9.345 49.595 9.715 ;
      RECT 49.26 6.175 49.56 9.715 ;
      RECT 49.255 5.47 49.555 6.53 ;
      RECT 45.025 5.47 49.555 5.77 ;
      RECT 47.82 3.81 48.12 5.77 ;
      RECT 45.025 4.27 45.325 5.77 ;
      RECT 48.545 4.805 48.875 5.16 ;
      RECT 46.64 4.845 48.875 5.145 ;
      RECT 46.64 3.71 46.94 5.145 ;
      RECT 44.72 4.27 45.45 4.6 ;
      RECT 47.615 3.815 48.395 4.16 ;
      RECT 48.07 3.78 48.395 4.16 ;
      RECT 46.625 3.71 46.955 4.04 ;
      RECT 45.91 3.71 46.23 4.625 ;
      RECT 45.91 3.71 46.24 4.245 ;
      RECT 33.965 9.345 34.335 9.715 ;
      RECT 34 6.175 34.3 9.715 ;
      RECT 33.995 5.47 34.295 6.53 ;
      RECT 29.765 5.47 34.295 5.77 ;
      RECT 32.56 3.81 32.86 5.77 ;
      RECT 29.765 4.27 30.065 5.77 ;
      RECT 33.285 4.805 33.615 5.16 ;
      RECT 31.38 4.845 33.615 5.145 ;
      RECT 31.38 3.71 31.68 5.145 ;
      RECT 29.46 4.27 30.19 4.6 ;
      RECT 32.355 3.815 33.135 4.16 ;
      RECT 32.81 3.78 33.135 4.16 ;
      RECT 31.365 3.71 31.695 4.04 ;
      RECT 30.65 3.71 30.97 4.625 ;
      RECT 30.65 3.71 30.98 4.245 ;
      RECT 103.4 7.205 103.78 12.465 ;
      RECT 97.245 3.15 97.975 3.48 ;
      RECT 95.555 3.165 96.285 3.495 ;
      RECT 94.52 3.15 95.25 3.5 ;
      RECT 92.97 3.175 93.7 3.505 ;
      RECT 88.14 7.205 88.52 12.465 ;
      RECT 81.985 3.15 82.715 3.48 ;
      RECT 80.295 3.165 81.025 3.495 ;
      RECT 79.26 3.15 79.99 3.5 ;
      RECT 77.71 3.175 78.44 3.505 ;
      RECT 72.88 7.205 73.26 12.465 ;
      RECT 66.725 3.15 67.455 3.48 ;
      RECT 65.035 3.165 65.765 3.495 ;
      RECT 64 3.15 64.73 3.5 ;
      RECT 62.45 3.175 63.18 3.505 ;
      RECT 57.62 7.205 58 12.465 ;
      RECT 51.465 3.15 52.195 3.48 ;
      RECT 49.775 3.165 50.505 3.495 ;
      RECT 48.74 3.15 49.47 3.5 ;
      RECT 47.19 3.175 47.92 3.505 ;
      RECT 42.36 7.205 42.74 12.465 ;
      RECT 36.205 3.15 36.935 3.48 ;
      RECT 34.515 3.165 35.245 3.495 ;
      RECT 33.48 3.15 34.21 3.5 ;
      RECT 31.93 3.175 32.66 3.505 ;
    LAYER via2 ;
      RECT 103.49 7.295 103.69 7.495 ;
      RECT 97.48 3.215 97.68 3.415 ;
      RECT 95.62 3.23 95.82 3.43 ;
      RECT 95.09 9.43 95.29 9.63 ;
      RECT 94.6 3.235 94.8 3.435 ;
      RECT 94.39 4.87 94.59 5.07 ;
      RECT 93.91 3.87 94.11 4.07 ;
      RECT 93.16 3.24 93.36 3.44 ;
      RECT 92.47 3.775 92.67 3.975 ;
      RECT 91.755 3.775 91.955 3.975 ;
      RECT 90.79 4.335 90.99 4.535 ;
      RECT 88.23 7.295 88.43 7.495 ;
      RECT 82.22 3.215 82.42 3.415 ;
      RECT 80.36 3.23 80.56 3.43 ;
      RECT 79.83 9.43 80.03 9.63 ;
      RECT 79.34 3.235 79.54 3.435 ;
      RECT 79.13 4.87 79.33 5.07 ;
      RECT 78.65 3.87 78.85 4.07 ;
      RECT 77.9 3.24 78.1 3.44 ;
      RECT 77.21 3.775 77.41 3.975 ;
      RECT 76.495 3.775 76.695 3.975 ;
      RECT 75.53 4.335 75.73 4.535 ;
      RECT 72.97 7.295 73.17 7.495 ;
      RECT 66.96 3.215 67.16 3.415 ;
      RECT 65.1 3.23 65.3 3.43 ;
      RECT 64.57 9.43 64.77 9.63 ;
      RECT 64.08 3.235 64.28 3.435 ;
      RECT 63.87 4.87 64.07 5.07 ;
      RECT 63.39 3.87 63.59 4.07 ;
      RECT 62.64 3.24 62.84 3.44 ;
      RECT 61.95 3.775 62.15 3.975 ;
      RECT 61.235 3.775 61.435 3.975 ;
      RECT 60.27 4.335 60.47 4.535 ;
      RECT 57.71 7.295 57.91 7.495 ;
      RECT 51.7 3.215 51.9 3.415 ;
      RECT 49.84 3.23 50.04 3.43 ;
      RECT 49.31 9.43 49.51 9.63 ;
      RECT 48.82 3.235 49.02 3.435 ;
      RECT 48.61 4.87 48.81 5.07 ;
      RECT 48.13 3.87 48.33 4.07 ;
      RECT 47.38 3.24 47.58 3.44 ;
      RECT 46.69 3.775 46.89 3.975 ;
      RECT 45.975 3.775 46.175 3.975 ;
      RECT 45.01 4.335 45.21 4.535 ;
      RECT 42.45 7.295 42.65 7.495 ;
      RECT 36.44 3.215 36.64 3.415 ;
      RECT 34.58 3.23 34.78 3.43 ;
      RECT 34.05 9.43 34.25 9.63 ;
      RECT 33.56 3.235 33.76 3.435 ;
      RECT 33.35 4.87 33.55 5.07 ;
      RECT 32.87 3.87 33.07 4.07 ;
      RECT 32.12 3.24 32.32 3.44 ;
      RECT 31.43 3.775 31.63 3.975 ;
      RECT 30.715 3.775 30.915 3.975 ;
      RECT 29.75 4.335 29.95 4.535 ;
    LAYER met2 ;
      RECT 26.175 10.69 103.675 10.86 ;
      RECT 103.505 9.565 103.675 10.86 ;
      RECT 26.175 8.545 26.345 10.86 ;
      RECT 103.475 9.565 103.825 9.915 ;
      RECT 26.115 8.545 26.405 8.895 ;
      RECT 100.315 8.51 100.635 8.835 ;
      RECT 100.345 7.985 100.515 8.835 ;
      RECT 100.345 7.985 100.52 8.335 ;
      RECT 100.345 7.985 101.32 8.16 ;
      RECT 101.145 3.26 101.32 8.16 ;
      RECT 101.09 3.26 101.44 3.61 ;
      RECT 101.115 8.945 101.44 9.27 ;
      RECT 100 9.035 101.44 9.205 ;
      RECT 100 3.69 100.16 9.205 ;
      RECT 100.315 3.66 100.635 3.98 ;
      RECT 100 3.69 100.635 3.86 ;
      RECT 97.45 4.835 97.71 5.155 ;
      RECT 97.51 3.13 97.65 5.155 ;
      RECT 98.71 3.995 99.05 4.345 ;
      RECT 98.085 4.065 99.05 4.265 ;
      RECT 98.085 3.235 98.285 4.265 ;
      RECT 97.335 3.69 97.65 4.06 ;
      RECT 98.8 3.99 98.97 4.345 ;
      RECT 97.405 3.245 97.65 4.06 ;
      RECT 97.44 3.13 97.72 3.5 ;
      RECT 97.44 3.235 98.285 3.435 ;
      RECT 96.76 3.715 97.02 4.035 ;
      RECT 96.1 3.805 97.02 3.945 ;
      RECT 96.1 2.865 96.24 3.945 ;
      RECT 92.56 3.155 92.82 3.475 ;
      RECT 92.74 2.865 92.88 3.385 ;
      RECT 92.74 2.865 96.24 3.005 ;
      RECT 88.19 8.95 88.54 9.3 ;
      RECT 95.675 8.905 96.025 9.255 ;
      RECT 88.19 8.98 96.025 9.18 ;
      RECT 95.59 4.555 95.85 4.875 ;
      RECT 95.65 3.145 95.79 4.875 ;
      RECT 95.58 3.145 95.86 3.515 ;
      RECT 92.98 5.305 95.415 5.445 ;
      RECT 95.275 3.995 95.415 5.445 ;
      RECT 92.98 4.925 93.12 5.445 ;
      RECT 92.68 4.925 93.12 5.155 ;
      RECT 90.34 4.925 93.12 5.065 ;
      RECT 92.68 4.835 92.94 5.155 ;
      RECT 90.34 4.645 90.48 5.065 ;
      RECT 89.83 4.555 90.09 4.875 ;
      RECT 89.83 4.645 90.48 4.785 ;
      RECT 89.885 4.435 90.03 4.875 ;
      RECT 89.89 3.155 90.03 4.875 ;
      RECT 95.215 3.995 95.475 4.315 ;
      RECT 89.885 3.155 90.03 3.615 ;
      RECT 89.825 3.155 90.09 3.475 ;
      RECT 94.84 4.835 95.105 5.155 ;
      RECT 94.9 3.245 95.04 5.155 ;
      RECT 94.56 3.245 95.04 3.52 ;
      RECT 94.36 3.15 94.84 3.495 ;
      RECT 94.35 4.785 94.63 5.155 ;
      RECT 94.42 3.69 94.56 5.155 ;
      RECT 94.36 3.69 94.62 4.315 ;
      RECT 94.35 3.69 94.63 4.06 ;
      RECT 93.28 4.835 93.54 5.155 ;
      RECT 93.28 4.645 93.48 5.155 ;
      RECT 93.085 4.645 93.48 4.785 ;
      RECT 93.085 3.155 93.225 4.785 ;
      RECT 93.085 3.155 93.4 3.525 ;
      RECT 93.025 3.155 93.4 3.475 ;
      RECT 90.75 4.25 91.03 4.62 ;
      RECT 92.2 4.275 92.46 4.595 ;
      RECT 90.58 4.365 92.46 4.505 ;
      RECT 90.58 4.25 91.03 4.505 ;
      RECT 90.52 3.69 90.78 4.315 ;
      RECT 90.51 3.69 90.79 4.06 ;
      RECT 91.59 3.69 92 4.06 ;
      RECT 91 3.715 91.26 4.035 ;
      RECT 91 3.805 92 3.945 ;
      RECT 85.055 8.51 85.375 8.835 ;
      RECT 85.085 7.985 85.255 8.835 ;
      RECT 85.085 7.985 85.26 8.335 ;
      RECT 85.085 7.985 86.06 8.16 ;
      RECT 85.885 3.26 86.06 8.16 ;
      RECT 85.83 3.26 86.18 3.61 ;
      RECT 85.855 8.945 86.18 9.27 ;
      RECT 84.74 9.035 86.18 9.205 ;
      RECT 84.74 3.69 84.9 9.205 ;
      RECT 85.055 3.66 85.375 3.98 ;
      RECT 84.74 3.69 85.375 3.86 ;
      RECT 82.19 4.835 82.45 5.155 ;
      RECT 82.25 3.13 82.39 5.155 ;
      RECT 83.45 3.995 83.79 4.345 ;
      RECT 82.825 4.065 83.79 4.265 ;
      RECT 82.825 3.235 83.025 4.265 ;
      RECT 82.075 3.69 82.39 4.06 ;
      RECT 83.54 3.99 83.71 4.345 ;
      RECT 82.145 3.245 82.39 4.06 ;
      RECT 82.18 3.13 82.46 3.5 ;
      RECT 82.18 3.235 83.025 3.435 ;
      RECT 81.5 3.715 81.76 4.035 ;
      RECT 80.84 3.805 81.76 3.945 ;
      RECT 80.84 2.865 80.98 3.945 ;
      RECT 77.3 3.155 77.56 3.475 ;
      RECT 77.48 2.865 77.62 3.385 ;
      RECT 77.48 2.865 80.98 3.005 ;
      RECT 72.93 8.95 73.28 9.3 ;
      RECT 80.42 8.905 80.77 9.255 ;
      RECT 72.93 8.98 80.77 9.18 ;
      RECT 80.33 4.555 80.59 4.875 ;
      RECT 80.39 3.145 80.53 4.875 ;
      RECT 80.32 3.145 80.6 3.515 ;
      RECT 77.72 5.305 80.155 5.445 ;
      RECT 80.015 3.995 80.155 5.445 ;
      RECT 77.72 4.925 77.86 5.445 ;
      RECT 77.42 4.925 77.86 5.155 ;
      RECT 75.08 4.925 77.86 5.065 ;
      RECT 77.42 4.835 77.68 5.155 ;
      RECT 75.08 4.645 75.22 5.065 ;
      RECT 74.57 4.555 74.83 4.875 ;
      RECT 74.57 4.645 75.22 4.785 ;
      RECT 74.625 4.435 74.77 4.875 ;
      RECT 74.63 3.155 74.77 4.875 ;
      RECT 79.955 3.995 80.215 4.315 ;
      RECT 74.625 3.155 74.77 3.615 ;
      RECT 74.565 3.155 74.83 3.475 ;
      RECT 79.58 4.835 79.845 5.155 ;
      RECT 79.64 3.245 79.78 5.155 ;
      RECT 79.3 3.245 79.78 3.52 ;
      RECT 79.1 3.15 79.58 3.495 ;
      RECT 79.09 4.785 79.37 5.155 ;
      RECT 79.16 3.69 79.3 5.155 ;
      RECT 79.1 3.69 79.36 4.315 ;
      RECT 79.09 3.69 79.37 4.06 ;
      RECT 78.02 4.835 78.28 5.155 ;
      RECT 78.02 4.645 78.22 5.155 ;
      RECT 77.825 4.645 78.22 4.785 ;
      RECT 77.825 3.155 77.965 4.785 ;
      RECT 77.825 3.155 78.14 3.525 ;
      RECT 77.765 3.155 78.14 3.475 ;
      RECT 75.49 4.25 75.77 4.62 ;
      RECT 76.94 4.275 77.2 4.595 ;
      RECT 75.32 4.365 77.2 4.505 ;
      RECT 75.32 4.25 75.77 4.505 ;
      RECT 75.26 3.69 75.52 4.315 ;
      RECT 75.25 3.69 75.53 4.06 ;
      RECT 76.33 3.69 76.74 4.06 ;
      RECT 75.74 3.715 76 4.035 ;
      RECT 75.74 3.805 76.74 3.945 ;
      RECT 69.795 8.51 70.115 8.835 ;
      RECT 69.825 7.985 69.995 8.835 ;
      RECT 69.825 7.985 70 8.335 ;
      RECT 69.825 7.985 70.8 8.16 ;
      RECT 70.625 3.26 70.8 8.16 ;
      RECT 70.57 3.26 70.92 3.61 ;
      RECT 70.595 8.945 70.92 9.27 ;
      RECT 69.48 9.035 70.92 9.205 ;
      RECT 69.48 3.69 69.64 9.205 ;
      RECT 69.795 3.66 70.115 3.98 ;
      RECT 69.48 3.69 70.115 3.86 ;
      RECT 66.93 4.835 67.19 5.155 ;
      RECT 66.99 3.13 67.13 5.155 ;
      RECT 68.19 3.995 68.53 4.345 ;
      RECT 67.565 4.065 68.53 4.265 ;
      RECT 67.565 3.235 67.765 4.265 ;
      RECT 66.815 3.69 67.13 4.06 ;
      RECT 68.28 3.99 68.45 4.345 ;
      RECT 66.885 3.245 67.13 4.06 ;
      RECT 66.92 3.13 67.2 3.5 ;
      RECT 66.92 3.235 67.765 3.435 ;
      RECT 66.24 3.715 66.5 4.035 ;
      RECT 65.58 3.805 66.5 3.945 ;
      RECT 65.58 2.865 65.72 3.945 ;
      RECT 62.04 3.155 62.3 3.475 ;
      RECT 62.22 2.865 62.36 3.385 ;
      RECT 62.22 2.865 65.72 3.005 ;
      RECT 57.715 8.95 58.065 9.3 ;
      RECT 65.155 8.905 65.505 9.255 ;
      RECT 57.715 8.98 65.505 9.18 ;
      RECT 65.07 4.555 65.33 4.875 ;
      RECT 65.13 3.145 65.27 4.875 ;
      RECT 65.06 3.145 65.34 3.515 ;
      RECT 62.46 5.305 64.895 5.445 ;
      RECT 64.755 3.995 64.895 5.445 ;
      RECT 62.46 4.925 62.6 5.445 ;
      RECT 62.16 4.925 62.6 5.155 ;
      RECT 59.82 4.925 62.6 5.065 ;
      RECT 62.16 4.835 62.42 5.155 ;
      RECT 59.82 4.645 59.96 5.065 ;
      RECT 59.31 4.555 59.57 4.875 ;
      RECT 59.31 4.645 59.96 4.785 ;
      RECT 59.365 4.435 59.51 4.875 ;
      RECT 59.37 3.155 59.51 4.875 ;
      RECT 64.695 3.995 64.955 4.315 ;
      RECT 59.365 3.155 59.51 3.615 ;
      RECT 59.305 3.155 59.57 3.475 ;
      RECT 64.32 4.835 64.585 5.155 ;
      RECT 64.38 3.245 64.52 5.155 ;
      RECT 64.04 3.245 64.52 3.52 ;
      RECT 63.84 3.15 64.32 3.495 ;
      RECT 63.83 4.785 64.11 5.155 ;
      RECT 63.9 3.69 64.04 5.155 ;
      RECT 63.84 3.69 64.1 4.315 ;
      RECT 63.83 3.69 64.11 4.06 ;
      RECT 62.76 4.835 63.02 5.155 ;
      RECT 62.76 4.645 62.96 5.155 ;
      RECT 62.565 4.645 62.96 4.785 ;
      RECT 62.565 3.155 62.705 4.785 ;
      RECT 62.565 3.155 62.88 3.525 ;
      RECT 62.505 3.155 62.88 3.475 ;
      RECT 60.23 4.25 60.51 4.62 ;
      RECT 61.68 4.275 61.94 4.595 ;
      RECT 60.06 4.365 61.94 4.505 ;
      RECT 60.06 4.25 60.51 4.505 ;
      RECT 60 3.69 60.26 4.315 ;
      RECT 59.99 3.69 60.27 4.06 ;
      RECT 61.07 3.69 61.48 4.06 ;
      RECT 60.48 3.715 60.74 4.035 ;
      RECT 60.48 3.805 61.48 3.945 ;
      RECT 54.535 8.51 54.855 8.835 ;
      RECT 54.565 7.985 54.735 8.835 ;
      RECT 54.565 7.985 54.74 8.335 ;
      RECT 54.565 7.985 55.54 8.16 ;
      RECT 55.365 3.26 55.54 8.16 ;
      RECT 55.31 3.26 55.66 3.61 ;
      RECT 55.335 8.945 55.66 9.27 ;
      RECT 54.22 9.035 55.66 9.205 ;
      RECT 54.22 3.69 54.38 9.205 ;
      RECT 54.535 3.66 54.855 3.98 ;
      RECT 54.22 3.69 54.855 3.86 ;
      RECT 51.67 4.835 51.93 5.155 ;
      RECT 51.73 3.13 51.87 5.155 ;
      RECT 52.93 3.995 53.27 4.345 ;
      RECT 52.305 4.065 53.27 4.265 ;
      RECT 52.305 3.235 52.505 4.265 ;
      RECT 51.555 3.69 51.87 4.06 ;
      RECT 53.02 3.99 53.19 4.345 ;
      RECT 51.625 3.245 51.87 4.06 ;
      RECT 51.66 3.13 51.94 3.5 ;
      RECT 51.66 3.235 52.505 3.435 ;
      RECT 50.98 3.715 51.24 4.035 ;
      RECT 50.32 3.805 51.24 3.945 ;
      RECT 50.32 2.865 50.46 3.945 ;
      RECT 46.78 3.155 47.04 3.475 ;
      RECT 46.96 2.865 47.1 3.385 ;
      RECT 46.96 2.865 50.46 3.005 ;
      RECT 42.455 8.95 42.805 9.3 ;
      RECT 49.895 8.905 50.245 9.255 ;
      RECT 42.455 8.98 50.245 9.18 ;
      RECT 49.81 4.555 50.07 4.875 ;
      RECT 49.87 3.145 50.01 4.875 ;
      RECT 49.8 3.145 50.08 3.515 ;
      RECT 47.2 5.305 49.635 5.445 ;
      RECT 49.495 3.995 49.635 5.445 ;
      RECT 47.2 4.925 47.34 5.445 ;
      RECT 46.9 4.925 47.34 5.155 ;
      RECT 44.56 4.925 47.34 5.065 ;
      RECT 46.9 4.835 47.16 5.155 ;
      RECT 44.56 4.645 44.7 5.065 ;
      RECT 44.05 4.555 44.31 4.875 ;
      RECT 44.05 4.645 44.7 4.785 ;
      RECT 44.105 4.435 44.25 4.875 ;
      RECT 44.11 3.155 44.25 4.875 ;
      RECT 49.435 3.995 49.695 4.315 ;
      RECT 44.105 3.155 44.25 3.615 ;
      RECT 44.045 3.155 44.31 3.475 ;
      RECT 49.06 4.835 49.325 5.155 ;
      RECT 49.12 3.245 49.26 5.155 ;
      RECT 48.78 3.245 49.26 3.52 ;
      RECT 48.58 3.15 49.06 3.495 ;
      RECT 48.57 4.785 48.85 5.155 ;
      RECT 48.64 3.69 48.78 5.155 ;
      RECT 48.58 3.69 48.84 4.315 ;
      RECT 48.57 3.69 48.85 4.06 ;
      RECT 47.5 4.835 47.76 5.155 ;
      RECT 47.5 4.645 47.7 5.155 ;
      RECT 47.305 4.645 47.7 4.785 ;
      RECT 47.305 3.155 47.445 4.785 ;
      RECT 47.305 3.155 47.62 3.525 ;
      RECT 47.245 3.155 47.62 3.475 ;
      RECT 44.97 4.25 45.25 4.62 ;
      RECT 46.42 4.275 46.68 4.595 ;
      RECT 44.8 4.365 46.68 4.505 ;
      RECT 44.8 4.25 45.25 4.505 ;
      RECT 44.74 3.69 45 4.315 ;
      RECT 44.73 3.69 45.01 4.06 ;
      RECT 45.81 3.69 46.22 4.06 ;
      RECT 45.22 3.715 45.48 4.035 ;
      RECT 45.22 3.805 46.22 3.945 ;
      RECT 39.275 8.51 39.595 8.835 ;
      RECT 39.305 7.985 39.475 8.835 ;
      RECT 39.305 7.985 39.48 8.335 ;
      RECT 39.305 7.985 40.28 8.16 ;
      RECT 40.105 3.26 40.28 8.16 ;
      RECT 40.05 3.26 40.4 3.61 ;
      RECT 40.075 8.945 40.4 9.27 ;
      RECT 38.96 9.035 40.4 9.205 ;
      RECT 38.96 3.69 39.12 9.205 ;
      RECT 39.275 3.66 39.595 3.98 ;
      RECT 38.96 3.69 39.595 3.86 ;
      RECT 36.41 4.835 36.67 5.155 ;
      RECT 36.47 3.13 36.61 5.155 ;
      RECT 37.67 3.995 38.01 4.345 ;
      RECT 37.045 4.065 38.01 4.265 ;
      RECT 37.045 3.235 37.245 4.265 ;
      RECT 36.295 3.69 36.61 4.06 ;
      RECT 37.76 3.99 37.93 4.345 ;
      RECT 36.365 3.245 36.61 4.06 ;
      RECT 36.4 3.13 36.68 3.5 ;
      RECT 36.4 3.235 37.245 3.435 ;
      RECT 35.72 3.715 35.98 4.035 ;
      RECT 35.06 3.805 35.98 3.945 ;
      RECT 35.06 2.865 35.2 3.945 ;
      RECT 31.52 3.155 31.78 3.475 ;
      RECT 31.7 2.865 31.84 3.385 ;
      RECT 31.7 2.865 35.2 3.005 ;
      RECT 26.49 9.285 26.78 9.635 ;
      RECT 26.49 9.355 27.71 9.525 ;
      RECT 27.54 8.975 27.71 9.525 ;
      RECT 34.635 8.895 34.985 9.245 ;
      RECT 27.54 8.975 34.985 9.145 ;
      RECT 34.55 4.555 34.81 4.875 ;
      RECT 34.61 3.145 34.75 4.875 ;
      RECT 34.54 3.145 34.82 3.515 ;
      RECT 31.94 5.305 34.375 5.445 ;
      RECT 34.235 3.995 34.375 5.445 ;
      RECT 31.94 4.925 32.08 5.445 ;
      RECT 31.64 4.925 32.08 5.155 ;
      RECT 29.3 4.925 32.08 5.065 ;
      RECT 31.64 4.835 31.9 5.155 ;
      RECT 29.3 4.645 29.44 5.065 ;
      RECT 28.79 4.555 29.05 4.875 ;
      RECT 28.79 4.645 29.44 4.785 ;
      RECT 28.845 4.435 28.99 4.875 ;
      RECT 28.85 3.155 28.99 4.875 ;
      RECT 34.175 3.995 34.435 4.315 ;
      RECT 28.845 3.155 28.99 3.615 ;
      RECT 28.785 3.155 29.05 3.475 ;
      RECT 33.8 4.835 34.065 5.155 ;
      RECT 33.86 3.245 34 5.155 ;
      RECT 33.52 3.245 34 3.52 ;
      RECT 33.32 3.15 33.8 3.495 ;
      RECT 33.31 4.785 33.59 5.155 ;
      RECT 33.38 3.69 33.52 5.155 ;
      RECT 33.32 3.69 33.58 4.315 ;
      RECT 33.31 3.69 33.59 4.06 ;
      RECT 32.24 4.835 32.5 5.155 ;
      RECT 32.24 4.645 32.44 5.155 ;
      RECT 32.045 4.645 32.44 4.785 ;
      RECT 32.045 3.155 32.185 4.785 ;
      RECT 32.045 3.155 32.36 3.525 ;
      RECT 31.985 3.155 32.36 3.475 ;
      RECT 29.71 4.25 29.99 4.62 ;
      RECT 31.16 4.275 31.42 4.595 ;
      RECT 29.54 4.365 31.42 4.505 ;
      RECT 29.54 4.25 29.99 4.505 ;
      RECT 29.48 3.69 29.74 4.315 ;
      RECT 29.47 3.69 29.75 4.06 ;
      RECT 30.55 3.69 30.96 4.06 ;
      RECT 29.96 3.715 30.22 4.035 ;
      RECT 29.96 3.805 30.96 3.945 ;
      RECT 103.4 7.205 103.78 7.585 ;
      RECT 95.005 9.345 95.375 9.715 ;
      RECT 93.87 3.69 94.15 4.155 ;
      RECT 93.63 3.155 93.91 3.5 ;
      RECT 92.43 3.69 92.71 4.06 ;
      RECT 88.14 7.205 88.52 7.585 ;
      RECT 79.745 9.345 80.115 9.715 ;
      RECT 78.61 3.69 78.89 4.155 ;
      RECT 78.37 3.155 78.65 3.5 ;
      RECT 77.17 3.69 77.45 4.06 ;
      RECT 72.88 7.205 73.26 7.585 ;
      RECT 64.485 9.345 64.855 9.715 ;
      RECT 63.35 3.69 63.63 4.155 ;
      RECT 63.11 3.155 63.39 3.5 ;
      RECT 61.91 3.69 62.19 4.06 ;
      RECT 57.62 7.205 58 7.585 ;
      RECT 49.225 9.345 49.595 9.715 ;
      RECT 48.09 3.69 48.37 4.155 ;
      RECT 47.85 3.155 48.13 3.5 ;
      RECT 46.65 3.69 46.93 4.06 ;
      RECT 42.36 7.205 42.74 7.585 ;
      RECT 33.965 9.345 34.335 9.715 ;
      RECT 32.83 3.69 33.11 4.155 ;
      RECT 32.59 3.155 32.87 3.5 ;
      RECT 31.39 3.69 31.67 4.06 ;
    LAYER via1 ;
      RECT 103.575 9.665 103.725 9.815 ;
      RECT 103.515 7.32 103.665 7.47 ;
      RECT 101.205 9.03 101.355 9.18 ;
      RECT 101.19 3.36 101.34 3.51 ;
      RECT 100.4 3.745 100.55 3.895 ;
      RECT 100.4 8.615 100.55 8.765 ;
      RECT 98.81 4.095 98.96 4.245 ;
      RECT 97.505 3.24 97.655 3.39 ;
      RECT 97.505 4.92 97.655 5.07 ;
      RECT 96.815 3.8 96.965 3.95 ;
      RECT 95.775 9.005 95.925 9.155 ;
      RECT 95.645 3.24 95.795 3.39 ;
      RECT 95.645 4.64 95.795 4.79 ;
      RECT 95.27 4.08 95.42 4.23 ;
      RECT 95.115 9.455 95.265 9.605 ;
      RECT 94.895 4.92 95.045 5.07 ;
      RECT 94.415 3.24 94.565 3.39 ;
      RECT 94.415 4.08 94.565 4.23 ;
      RECT 93.935 3.8 94.085 3.95 ;
      RECT 93.695 3.24 93.845 3.39 ;
      RECT 93.335 4.92 93.485 5.07 ;
      RECT 93.08 3.24 93.23 3.39 ;
      RECT 92.735 4.92 92.885 5.07 ;
      RECT 92.615 3.24 92.765 3.39 ;
      RECT 92.495 3.8 92.645 3.95 ;
      RECT 92.255 4.36 92.405 4.51 ;
      RECT 91.055 3.8 91.205 3.95 ;
      RECT 90.575 4.08 90.725 4.23 ;
      RECT 89.885 4.64 90.035 4.79 ;
      RECT 89.88 3.24 90.03 3.39 ;
      RECT 88.29 9.05 88.44 9.2 ;
      RECT 88.255 7.32 88.405 7.47 ;
      RECT 85.945 9.03 86.095 9.18 ;
      RECT 85.93 3.36 86.08 3.51 ;
      RECT 85.14 3.745 85.29 3.895 ;
      RECT 85.14 8.615 85.29 8.765 ;
      RECT 83.55 4.095 83.7 4.245 ;
      RECT 82.245 3.24 82.395 3.39 ;
      RECT 82.245 4.92 82.395 5.07 ;
      RECT 81.555 3.8 81.705 3.95 ;
      RECT 80.52 9.005 80.67 9.155 ;
      RECT 80.385 3.24 80.535 3.39 ;
      RECT 80.385 4.64 80.535 4.79 ;
      RECT 80.01 4.08 80.16 4.23 ;
      RECT 79.855 9.455 80.005 9.605 ;
      RECT 79.635 4.92 79.785 5.07 ;
      RECT 79.155 3.24 79.305 3.39 ;
      RECT 79.155 4.08 79.305 4.23 ;
      RECT 78.675 3.8 78.825 3.95 ;
      RECT 78.435 3.24 78.585 3.39 ;
      RECT 78.075 4.92 78.225 5.07 ;
      RECT 77.82 3.24 77.97 3.39 ;
      RECT 77.475 4.92 77.625 5.07 ;
      RECT 77.355 3.24 77.505 3.39 ;
      RECT 77.235 3.8 77.385 3.95 ;
      RECT 76.995 4.36 77.145 4.51 ;
      RECT 75.795 3.8 75.945 3.95 ;
      RECT 75.315 4.08 75.465 4.23 ;
      RECT 74.625 4.64 74.775 4.79 ;
      RECT 74.62 3.24 74.77 3.39 ;
      RECT 73.03 9.05 73.18 9.2 ;
      RECT 72.995 7.32 73.145 7.47 ;
      RECT 70.685 9.03 70.835 9.18 ;
      RECT 70.67 3.36 70.82 3.51 ;
      RECT 69.88 3.745 70.03 3.895 ;
      RECT 69.88 8.615 70.03 8.765 ;
      RECT 68.29 4.095 68.44 4.245 ;
      RECT 66.985 3.24 67.135 3.39 ;
      RECT 66.985 4.92 67.135 5.07 ;
      RECT 66.295 3.8 66.445 3.95 ;
      RECT 65.255 9.005 65.405 9.155 ;
      RECT 65.125 3.24 65.275 3.39 ;
      RECT 65.125 4.64 65.275 4.79 ;
      RECT 64.75 4.08 64.9 4.23 ;
      RECT 64.595 9.455 64.745 9.605 ;
      RECT 64.375 4.92 64.525 5.07 ;
      RECT 63.895 3.24 64.045 3.39 ;
      RECT 63.895 4.08 64.045 4.23 ;
      RECT 63.415 3.8 63.565 3.95 ;
      RECT 63.175 3.24 63.325 3.39 ;
      RECT 62.815 4.92 62.965 5.07 ;
      RECT 62.56 3.24 62.71 3.39 ;
      RECT 62.215 4.92 62.365 5.07 ;
      RECT 62.095 3.24 62.245 3.39 ;
      RECT 61.975 3.8 62.125 3.95 ;
      RECT 61.735 4.36 61.885 4.51 ;
      RECT 60.535 3.8 60.685 3.95 ;
      RECT 60.055 4.08 60.205 4.23 ;
      RECT 59.365 4.64 59.515 4.79 ;
      RECT 59.36 3.24 59.51 3.39 ;
      RECT 57.815 9.05 57.965 9.2 ;
      RECT 57.735 7.32 57.885 7.47 ;
      RECT 55.425 9.03 55.575 9.18 ;
      RECT 55.41 3.36 55.56 3.51 ;
      RECT 54.62 3.745 54.77 3.895 ;
      RECT 54.62 8.615 54.77 8.765 ;
      RECT 53.03 4.095 53.18 4.245 ;
      RECT 51.725 3.24 51.875 3.39 ;
      RECT 51.725 4.92 51.875 5.07 ;
      RECT 51.035 3.8 51.185 3.95 ;
      RECT 49.995 9.005 50.145 9.155 ;
      RECT 49.865 3.24 50.015 3.39 ;
      RECT 49.865 4.64 50.015 4.79 ;
      RECT 49.49 4.08 49.64 4.23 ;
      RECT 49.335 9.455 49.485 9.605 ;
      RECT 49.115 4.92 49.265 5.07 ;
      RECT 48.635 3.24 48.785 3.39 ;
      RECT 48.635 4.08 48.785 4.23 ;
      RECT 48.155 3.8 48.305 3.95 ;
      RECT 47.915 3.24 48.065 3.39 ;
      RECT 47.555 4.92 47.705 5.07 ;
      RECT 47.3 3.24 47.45 3.39 ;
      RECT 46.955 4.92 47.105 5.07 ;
      RECT 46.835 3.24 46.985 3.39 ;
      RECT 46.715 3.8 46.865 3.95 ;
      RECT 46.475 4.36 46.625 4.51 ;
      RECT 45.275 3.8 45.425 3.95 ;
      RECT 44.795 4.08 44.945 4.23 ;
      RECT 44.105 4.64 44.255 4.79 ;
      RECT 44.1 3.24 44.25 3.39 ;
      RECT 42.555 9.05 42.705 9.2 ;
      RECT 42.475 7.32 42.625 7.47 ;
      RECT 40.165 9.03 40.315 9.18 ;
      RECT 40.15 3.36 40.3 3.51 ;
      RECT 39.36 3.745 39.51 3.895 ;
      RECT 39.36 8.615 39.51 8.765 ;
      RECT 37.77 4.095 37.92 4.245 ;
      RECT 36.465 3.24 36.615 3.39 ;
      RECT 36.465 4.92 36.615 5.07 ;
      RECT 35.775 3.8 35.925 3.95 ;
      RECT 34.735 8.995 34.885 9.145 ;
      RECT 34.605 3.24 34.755 3.39 ;
      RECT 34.605 4.64 34.755 4.79 ;
      RECT 34.23 4.08 34.38 4.23 ;
      RECT 34.075 9.455 34.225 9.605 ;
      RECT 33.855 4.92 34.005 5.07 ;
      RECT 33.375 3.24 33.525 3.39 ;
      RECT 33.375 4.08 33.525 4.23 ;
      RECT 32.895 3.8 33.045 3.95 ;
      RECT 32.655 3.24 32.805 3.39 ;
      RECT 32.295 4.92 32.445 5.07 ;
      RECT 32.04 3.24 32.19 3.39 ;
      RECT 31.695 4.92 31.845 5.07 ;
      RECT 31.575 3.24 31.725 3.39 ;
      RECT 31.455 3.8 31.605 3.95 ;
      RECT 31.215 4.36 31.365 4.51 ;
      RECT 30.015 3.8 30.165 3.95 ;
      RECT 29.535 4.08 29.685 4.23 ;
      RECT 28.845 4.64 28.995 4.79 ;
      RECT 28.84 3.24 28.99 3.39 ;
      RECT 26.56 9.385 26.71 9.535 ;
      RECT 26.185 8.645 26.335 8.795 ;
    LAYER met1 ;
      RECT 103.44 10.06 103.735 10.29 ;
      RECT 103.5 9.565 103.675 10.29 ;
      RECT 103.475 9.565 103.825 9.915 ;
      RECT 103.5 8.58 103.67 10.29 ;
      RECT 103.44 8.58 103.73 8.81 ;
      RECT 102.45 10.06 102.745 10.29 ;
      RECT 102.51 8.58 102.68 10.29 ;
      RECT 102.45 8.58 102.74 8.81 ;
      RECT 102.45 8.615 103.3 8.775 ;
      RECT 103.135 8.21 103.3 8.775 ;
      RECT 102.45 8.61 102.845 8.775 ;
      RECT 103.07 8.21 103.36 8.44 ;
      RECT 103.07 8.24 103.53 8.41 ;
      RECT 103.035 4.025 103.355 4.26 ;
      RECT 103.035 4.055 103.525 4.225 ;
      RECT 103.035 3.69 103.225 4.26 ;
      RECT 102.45 3.655 102.74 3.885 ;
      RECT 102.45 3.69 103.225 3.86 ;
      RECT 102.51 2.175 102.68 3.885 ;
      RECT 102.45 2.175 102.745 2.405 ;
      RECT 102.08 4.025 102.37 4.255 ;
      RECT 102.08 4.055 102.54 4.225 ;
      RECT 102.145 2.95 102.31 4.255 ;
      RECT 100.66 2.915 100.95 3.145 ;
      RECT 100.66 2.95 102.31 3.12 ;
      RECT 100.72 2.175 100.89 3.145 ;
      RECT 100.66 2.175 100.95 2.405 ;
      RECT 100.66 10.06 100.95 10.29 ;
      RECT 100.72 9.32 100.89 10.29 ;
      RECT 100.72 9.41 102.31 9.58 ;
      RECT 102.14 8.21 102.31 9.58 ;
      RECT 100.66 9.32 100.95 9.55 ;
      RECT 102.08 8.21 102.37 8.44 ;
      RECT 102.08 8.24 102.54 8.41 ;
      RECT 98.71 3.995 99.05 4.345 ;
      RECT 98.8 3.32 98.97 4.345 ;
      RECT 101.09 3.26 101.44 3.61 ;
      RECT 98.8 3.32 101.44 3.49 ;
      RECT 100.92 3.315 101.44 3.49 ;
      RECT 101.115 8.945 101.44 9.27 ;
      RECT 95.675 8.905 96.025 9.255 ;
      RECT 101.09 8.95 101.44 9.18 ;
      RECT 95.475 8.95 96.025 9.18 ;
      RECT 100.92 8.975 101.44 9.15 ;
      RECT 95.305 8.98 96.025 9.15 ;
      RECT 95.365 8.975 101.44 9.145 ;
      RECT 100.315 3.66 100.635 3.98 ;
      RECT 100.29 3.655 100.58 3.885 ;
      RECT 100.28 3.685 100.635 3.86 ;
      RECT 100.115 3.685 100.635 3.855 ;
      RECT 100.315 8.545 100.635 8.835 ;
      RECT 100.29 8.58 100.635 8.81 ;
      RECT 100.115 8.61 100.635 8.78 ;
      RECT 97.42 3.185 97.74 3.445 ;
      RECT 96.985 3.2 97.275 3.43 ;
      RECT 96.985 3.245 97.74 3.385 ;
      RECT 97.42 4.865 97.74 5.125 ;
      RECT 96.985 4.88 97.275 5.11 ;
      RECT 96.985 4.925 97.74 5.065 ;
      RECT 96.745 4.32 97.035 4.55 ;
      RECT 96.745 4.365 97.32 4.505 ;
      RECT 97.18 4.225 97.44 4.365 ;
      RECT 97.225 4.04 97.515 4.27 ;
      RECT 95.38 4.225 96.48 4.365 ;
      RECT 95.185 4.025 95.505 4.285 ;
      RECT 96.265 4.04 96.555 4.27 ;
      RECT 95.185 4.04 95.595 4.285 ;
      RECT 95.56 3.185 95.88 3.445 ;
      RECT 96.025 3.2 96.315 3.43 ;
      RECT 95.56 3.245 96.315 3.385 ;
      RECT 93.175 4.365 93.35 4.69 ;
      RECT 92.86 4.45 95.04 4.59 ;
      RECT 94.9 3.46 95.04 4.59 ;
      RECT 92.86 4.365 94.155 4.59 ;
      RECT 93.865 4.32 94.155 4.59 ;
      RECT 92.86 4.085 93.195 4.59 ;
      RECT 92.905 4.04 93.195 4.59 ;
      RECT 95.785 3.76 96.075 3.99 ;
      RECT 94.9 3.665 96 3.805 ;
      RECT 94.825 3.46 95.115 3.71 ;
      RECT 95.045 10.06 95.335 10.29 ;
      RECT 95.105 9.32 95.275 10.29 ;
      RECT 95.005 9.345 95.375 9.715 ;
      RECT 95.045 9.32 95.335 9.715 ;
      RECT 94.81 4.865 95.135 5.125 ;
      RECT 94.81 4.88 95.33 5.11 ;
      RECT 93.385 3.76 93.675 3.99 ;
      RECT 93.535 3.365 93.675 3.99 ;
      RECT 93.535 3.365 93.84 3.505 ;
      RECT 94.33 3.185 94.65 3.445 ;
      RECT 93.61 3.185 93.93 3.445 ;
      RECT 94.105 3.2 94.65 3.43 ;
      RECT 93.61 3.245 94.65 3.385 ;
      RECT 93.25 4.865 93.57 5.125 ;
      RECT 93.145 4.88 93.57 5.11 ;
      RECT 91.225 4.32 91.515 4.55 ;
      RECT 91.225 4.32 91.68 4.505 ;
      RECT 91.54 3.845 91.68 4.505 ;
      RECT 91.66 3.245 91.8 3.985 ;
      RECT 92.53 3.185 92.85 3.445 ;
      RECT 91.705 3.2 91.995 3.43 ;
      RECT 91.66 3.245 92.85 3.385 ;
      RECT 92.41 3.745 92.73 4.005 ;
      RECT 91.945 3.76 92.235 3.99 ;
      RECT 91.945 3.805 92.73 3.945 ;
      RECT 92.17 4.305 92.49 4.565 ;
      RECT 92.17 4.32 92.715 4.55 ;
      RECT 91.705 4.88 91.995 5.11 ;
      RECT 90.82 4.76 91.92 4.9 ;
      RECT 90.745 4.6 91.035 4.83 ;
      RECT 88.18 10.06 88.475 10.29 ;
      RECT 88.24 8.58 88.41 10.29 ;
      RECT 88.19 8.95 88.54 9.3 ;
      RECT 88.18 8.58 88.47 8.81 ;
      RECT 87.19 10.06 87.485 10.29 ;
      RECT 87.25 8.58 87.42 10.29 ;
      RECT 87.19 8.58 87.48 8.81 ;
      RECT 87.19 8.615 88.04 8.775 ;
      RECT 87.875 8.21 88.04 8.775 ;
      RECT 87.19 8.61 87.585 8.775 ;
      RECT 87.81 8.21 88.1 8.44 ;
      RECT 87.81 8.24 88.27 8.41 ;
      RECT 87.775 4.025 88.095 4.26 ;
      RECT 87.775 4.055 88.265 4.225 ;
      RECT 87.775 3.69 87.965 4.26 ;
      RECT 87.19 3.655 87.48 3.885 ;
      RECT 87.19 3.69 87.965 3.86 ;
      RECT 87.25 2.175 87.42 3.885 ;
      RECT 87.19 2.175 87.485 2.405 ;
      RECT 86.82 4.025 87.11 4.255 ;
      RECT 86.82 4.055 87.28 4.225 ;
      RECT 86.885 2.95 87.05 4.255 ;
      RECT 85.4 2.915 85.69 3.145 ;
      RECT 85.4 2.95 87.05 3.12 ;
      RECT 85.46 2.175 85.63 3.145 ;
      RECT 85.4 2.175 85.69 2.405 ;
      RECT 85.4 10.06 85.69 10.29 ;
      RECT 85.46 9.32 85.63 10.29 ;
      RECT 85.46 9.41 87.05 9.58 ;
      RECT 86.88 8.21 87.05 9.58 ;
      RECT 85.4 9.32 85.69 9.55 ;
      RECT 86.82 8.21 87.11 8.44 ;
      RECT 86.82 8.24 87.28 8.41 ;
      RECT 83.45 3.995 83.79 4.345 ;
      RECT 83.54 3.32 83.71 4.345 ;
      RECT 85.83 3.26 86.18 3.61 ;
      RECT 83.54 3.32 86.18 3.49 ;
      RECT 85.66 3.315 86.18 3.49 ;
      RECT 85.855 8.945 86.18 9.27 ;
      RECT 80.42 8.905 80.77 9.255 ;
      RECT 85.83 8.95 86.18 9.18 ;
      RECT 80.215 8.95 80.77 9.18 ;
      RECT 85.66 8.975 86.18 9.15 ;
      RECT 80.045 8.98 80.77 9.15 ;
      RECT 80.105 8.975 86.18 9.145 ;
      RECT 85.055 3.66 85.375 3.98 ;
      RECT 85.03 3.655 85.32 3.885 ;
      RECT 85.02 3.685 85.375 3.86 ;
      RECT 84.855 3.685 85.375 3.855 ;
      RECT 85.055 8.545 85.375 8.835 ;
      RECT 85.03 8.58 85.375 8.81 ;
      RECT 84.855 8.61 85.375 8.78 ;
      RECT 82.16 3.185 82.48 3.445 ;
      RECT 81.725 3.2 82.015 3.43 ;
      RECT 81.725 3.245 82.48 3.385 ;
      RECT 82.16 4.865 82.48 5.125 ;
      RECT 81.725 4.88 82.015 5.11 ;
      RECT 81.725 4.925 82.48 5.065 ;
      RECT 81.485 4.32 81.775 4.55 ;
      RECT 81.485 4.365 82.06 4.505 ;
      RECT 81.92 4.225 82.18 4.365 ;
      RECT 81.965 4.04 82.255 4.27 ;
      RECT 80.12 4.225 81.22 4.365 ;
      RECT 79.925 4.025 80.245 4.285 ;
      RECT 81.005 4.04 81.295 4.27 ;
      RECT 79.925 4.04 80.335 4.285 ;
      RECT 80.3 3.185 80.62 3.445 ;
      RECT 80.765 3.2 81.055 3.43 ;
      RECT 80.3 3.245 81.055 3.385 ;
      RECT 77.915 4.365 78.09 4.69 ;
      RECT 77.6 4.45 79.78 4.59 ;
      RECT 79.64 3.46 79.78 4.59 ;
      RECT 77.6 4.365 78.895 4.59 ;
      RECT 78.605 4.32 78.895 4.59 ;
      RECT 77.6 4.085 77.935 4.59 ;
      RECT 77.645 4.04 77.935 4.59 ;
      RECT 80.525 3.76 80.815 3.99 ;
      RECT 79.64 3.665 80.74 3.805 ;
      RECT 79.565 3.46 79.855 3.71 ;
      RECT 79.785 10.06 80.075 10.29 ;
      RECT 79.845 9.32 80.015 10.29 ;
      RECT 79.745 9.345 80.115 9.715 ;
      RECT 79.785 9.32 80.075 9.715 ;
      RECT 79.55 4.865 79.875 5.125 ;
      RECT 79.55 4.88 80.07 5.11 ;
      RECT 78.125 3.76 78.415 3.99 ;
      RECT 78.275 3.365 78.415 3.99 ;
      RECT 78.275 3.365 78.58 3.505 ;
      RECT 79.07 3.185 79.39 3.445 ;
      RECT 78.35 3.185 78.67 3.445 ;
      RECT 78.845 3.2 79.39 3.43 ;
      RECT 78.35 3.245 79.39 3.385 ;
      RECT 77.99 4.865 78.31 5.125 ;
      RECT 77.885 4.88 78.31 5.11 ;
      RECT 75.965 4.32 76.255 4.55 ;
      RECT 75.965 4.32 76.42 4.505 ;
      RECT 76.28 3.845 76.42 4.505 ;
      RECT 76.4 3.245 76.54 3.985 ;
      RECT 77.27 3.185 77.59 3.445 ;
      RECT 76.445 3.2 76.735 3.43 ;
      RECT 76.4 3.245 77.59 3.385 ;
      RECT 77.15 3.745 77.47 4.005 ;
      RECT 76.685 3.76 76.975 3.99 ;
      RECT 76.685 3.805 77.47 3.945 ;
      RECT 76.91 4.305 77.23 4.565 ;
      RECT 76.91 4.32 77.455 4.55 ;
      RECT 76.445 4.88 76.735 5.11 ;
      RECT 75.56 4.76 76.66 4.9 ;
      RECT 75.485 4.6 75.775 4.83 ;
      RECT 72.92 10.06 73.215 10.29 ;
      RECT 72.98 8.58 73.15 10.29 ;
      RECT 72.93 8.95 73.28 9.3 ;
      RECT 72.92 8.58 73.21 8.81 ;
      RECT 71.93 10.06 72.225 10.29 ;
      RECT 71.99 8.58 72.16 10.29 ;
      RECT 71.93 8.58 72.22 8.81 ;
      RECT 71.93 8.615 72.78 8.775 ;
      RECT 72.615 8.21 72.78 8.775 ;
      RECT 71.93 8.61 72.325 8.775 ;
      RECT 72.55 8.21 72.84 8.44 ;
      RECT 72.55 8.24 73.01 8.41 ;
      RECT 72.515 4.025 72.835 4.26 ;
      RECT 72.515 4.055 73.005 4.225 ;
      RECT 72.515 3.69 72.705 4.26 ;
      RECT 71.93 3.655 72.22 3.885 ;
      RECT 71.93 3.69 72.705 3.86 ;
      RECT 71.99 2.175 72.16 3.885 ;
      RECT 71.93 2.175 72.225 2.405 ;
      RECT 71.56 4.025 71.85 4.255 ;
      RECT 71.56 4.055 72.02 4.225 ;
      RECT 71.625 2.95 71.79 4.255 ;
      RECT 70.14 2.915 70.43 3.145 ;
      RECT 70.14 2.95 71.79 3.12 ;
      RECT 70.2 2.175 70.37 3.145 ;
      RECT 70.14 2.175 70.43 2.405 ;
      RECT 70.14 10.06 70.43 10.29 ;
      RECT 70.2 9.32 70.37 10.29 ;
      RECT 70.2 9.41 71.79 9.58 ;
      RECT 71.62 8.21 71.79 9.58 ;
      RECT 70.14 9.32 70.43 9.55 ;
      RECT 71.56 8.21 71.85 8.44 ;
      RECT 71.56 8.24 72.02 8.41 ;
      RECT 68.19 3.995 68.53 4.345 ;
      RECT 68.28 3.32 68.45 4.345 ;
      RECT 70.57 3.26 70.92 3.61 ;
      RECT 68.28 3.32 70.92 3.49 ;
      RECT 70.4 3.315 70.92 3.49 ;
      RECT 70.595 8.945 70.92 9.27 ;
      RECT 65.155 8.905 65.505 9.255 ;
      RECT 70.57 8.95 70.92 9.18 ;
      RECT 64.955 8.95 65.505 9.18 ;
      RECT 70.4 8.975 70.92 9.15 ;
      RECT 64.785 8.98 65.505 9.15 ;
      RECT 64.845 8.975 70.92 9.145 ;
      RECT 69.795 3.66 70.115 3.98 ;
      RECT 69.77 3.655 70.06 3.885 ;
      RECT 69.76 3.685 70.115 3.86 ;
      RECT 69.595 3.685 70.115 3.855 ;
      RECT 69.795 8.545 70.115 8.835 ;
      RECT 69.77 8.58 70.115 8.81 ;
      RECT 69.595 8.61 70.115 8.78 ;
      RECT 66.9 3.185 67.22 3.445 ;
      RECT 66.465 3.2 66.755 3.43 ;
      RECT 66.465 3.245 67.22 3.385 ;
      RECT 66.9 4.865 67.22 5.125 ;
      RECT 66.465 4.88 66.755 5.11 ;
      RECT 66.465 4.925 67.22 5.065 ;
      RECT 66.225 4.32 66.515 4.55 ;
      RECT 66.225 4.365 66.8 4.505 ;
      RECT 66.66 4.225 66.92 4.365 ;
      RECT 66.705 4.04 66.995 4.27 ;
      RECT 64.86 4.225 65.96 4.365 ;
      RECT 64.665 4.025 64.985 4.285 ;
      RECT 65.745 4.04 66.035 4.27 ;
      RECT 64.665 4.04 65.075 4.285 ;
      RECT 65.04 3.185 65.36 3.445 ;
      RECT 65.505 3.2 65.795 3.43 ;
      RECT 65.04 3.245 65.795 3.385 ;
      RECT 62.655 4.365 62.83 4.69 ;
      RECT 62.34 4.45 64.52 4.59 ;
      RECT 64.38 3.46 64.52 4.59 ;
      RECT 62.34 4.365 63.635 4.59 ;
      RECT 63.345 4.32 63.635 4.59 ;
      RECT 62.34 4.085 62.675 4.59 ;
      RECT 62.385 4.04 62.675 4.59 ;
      RECT 65.265 3.76 65.555 3.99 ;
      RECT 64.38 3.665 65.48 3.805 ;
      RECT 64.305 3.46 64.595 3.71 ;
      RECT 64.525 10.06 64.815 10.29 ;
      RECT 64.585 9.32 64.755 10.29 ;
      RECT 64.485 9.345 64.855 9.715 ;
      RECT 64.525 9.32 64.815 9.715 ;
      RECT 64.29 4.865 64.615 5.125 ;
      RECT 64.29 4.88 64.81 5.11 ;
      RECT 62.865 3.76 63.155 3.99 ;
      RECT 63.015 3.365 63.155 3.99 ;
      RECT 63.015 3.365 63.32 3.505 ;
      RECT 63.81 3.185 64.13 3.445 ;
      RECT 63.09 3.185 63.41 3.445 ;
      RECT 63.585 3.2 64.13 3.43 ;
      RECT 63.09 3.245 64.13 3.385 ;
      RECT 62.73 4.865 63.05 5.125 ;
      RECT 62.625 4.88 63.05 5.11 ;
      RECT 60.705 4.32 60.995 4.55 ;
      RECT 60.705 4.32 61.16 4.505 ;
      RECT 61.02 3.845 61.16 4.505 ;
      RECT 61.14 3.245 61.28 3.985 ;
      RECT 62.01 3.185 62.33 3.445 ;
      RECT 61.185 3.2 61.475 3.43 ;
      RECT 61.14 3.245 62.33 3.385 ;
      RECT 61.89 3.745 62.21 4.005 ;
      RECT 61.425 3.76 61.715 3.99 ;
      RECT 61.425 3.805 62.21 3.945 ;
      RECT 61.65 4.305 61.97 4.565 ;
      RECT 61.65 4.32 62.195 4.55 ;
      RECT 61.185 4.88 61.475 5.11 ;
      RECT 60.3 4.76 61.4 4.9 ;
      RECT 60.225 4.6 60.515 4.83 ;
      RECT 57.66 10.06 57.955 10.29 ;
      RECT 57.72 8.58 57.89 10.29 ;
      RECT 57.71 8.95 58.065 9.305 ;
      RECT 57.66 8.58 57.95 8.81 ;
      RECT 56.67 10.06 56.965 10.29 ;
      RECT 56.73 8.58 56.9 10.29 ;
      RECT 56.67 8.58 56.96 8.81 ;
      RECT 56.67 8.615 57.52 8.775 ;
      RECT 57.355 8.21 57.52 8.775 ;
      RECT 56.67 8.61 57.065 8.775 ;
      RECT 57.29 8.21 57.58 8.44 ;
      RECT 57.29 8.24 57.75 8.41 ;
      RECT 57.255 4.025 57.575 4.26 ;
      RECT 57.255 4.055 57.745 4.225 ;
      RECT 57.255 3.69 57.445 4.26 ;
      RECT 56.67 3.655 56.96 3.885 ;
      RECT 56.67 3.69 57.445 3.86 ;
      RECT 56.73 2.175 56.9 3.885 ;
      RECT 56.67 2.175 56.965 2.405 ;
      RECT 56.3 4.025 56.59 4.255 ;
      RECT 56.3 4.055 56.76 4.225 ;
      RECT 56.365 2.95 56.53 4.255 ;
      RECT 54.88 2.915 55.17 3.145 ;
      RECT 54.88 2.95 56.53 3.12 ;
      RECT 54.94 2.175 55.11 3.145 ;
      RECT 54.88 2.175 55.17 2.405 ;
      RECT 54.88 10.06 55.17 10.29 ;
      RECT 54.94 9.32 55.11 10.29 ;
      RECT 54.94 9.41 56.53 9.58 ;
      RECT 56.36 8.21 56.53 9.58 ;
      RECT 54.88 9.32 55.17 9.55 ;
      RECT 56.3 8.21 56.59 8.44 ;
      RECT 56.3 8.24 56.76 8.41 ;
      RECT 52.93 3.995 53.27 4.345 ;
      RECT 53.02 3.32 53.19 4.345 ;
      RECT 55.31 3.26 55.66 3.61 ;
      RECT 53.02 3.32 55.66 3.49 ;
      RECT 55.14 3.315 55.66 3.49 ;
      RECT 55.335 8.945 55.66 9.27 ;
      RECT 49.895 8.905 50.245 9.255 ;
      RECT 55.31 8.95 55.66 9.18 ;
      RECT 49.695 8.95 50.245 9.18 ;
      RECT 55.14 8.975 55.66 9.15 ;
      RECT 49.525 8.98 50.245 9.15 ;
      RECT 49.585 8.975 55.66 9.145 ;
      RECT 54.535 3.66 54.855 3.98 ;
      RECT 54.51 3.655 54.8 3.885 ;
      RECT 54.5 3.685 54.855 3.86 ;
      RECT 54.335 3.685 54.855 3.855 ;
      RECT 54.535 8.545 54.855 8.835 ;
      RECT 54.51 8.58 54.855 8.81 ;
      RECT 54.335 8.61 54.855 8.78 ;
      RECT 51.64 3.185 51.96 3.445 ;
      RECT 51.205 3.2 51.495 3.43 ;
      RECT 51.205 3.245 51.96 3.385 ;
      RECT 51.64 4.865 51.96 5.125 ;
      RECT 51.205 4.88 51.495 5.11 ;
      RECT 51.205 4.925 51.96 5.065 ;
      RECT 50.965 4.32 51.255 4.55 ;
      RECT 50.965 4.365 51.54 4.505 ;
      RECT 51.4 4.225 51.66 4.365 ;
      RECT 51.445 4.04 51.735 4.27 ;
      RECT 49.6 4.225 50.7 4.365 ;
      RECT 49.405 4.025 49.725 4.285 ;
      RECT 50.485 4.04 50.775 4.27 ;
      RECT 49.405 4.04 49.815 4.285 ;
      RECT 49.78 3.185 50.1 3.445 ;
      RECT 50.245 3.2 50.535 3.43 ;
      RECT 49.78 3.245 50.535 3.385 ;
      RECT 47.395 4.365 47.57 4.69 ;
      RECT 47.08 4.45 49.26 4.59 ;
      RECT 49.12 3.46 49.26 4.59 ;
      RECT 47.08 4.365 48.375 4.59 ;
      RECT 48.085 4.32 48.375 4.59 ;
      RECT 47.08 4.085 47.415 4.59 ;
      RECT 47.125 4.04 47.415 4.59 ;
      RECT 50.005 3.76 50.295 3.99 ;
      RECT 49.12 3.665 50.22 3.805 ;
      RECT 49.045 3.46 49.335 3.71 ;
      RECT 49.265 10.06 49.555 10.29 ;
      RECT 49.325 9.32 49.495 10.29 ;
      RECT 49.225 9.345 49.595 9.715 ;
      RECT 49.265 9.32 49.555 9.715 ;
      RECT 49.03 4.865 49.355 5.125 ;
      RECT 49.03 4.88 49.55 5.11 ;
      RECT 47.605 3.76 47.895 3.99 ;
      RECT 47.755 3.365 47.895 3.99 ;
      RECT 47.755 3.365 48.06 3.505 ;
      RECT 48.55 3.185 48.87 3.445 ;
      RECT 47.83 3.185 48.15 3.445 ;
      RECT 48.325 3.2 48.87 3.43 ;
      RECT 47.83 3.245 48.87 3.385 ;
      RECT 47.47 4.865 47.79 5.125 ;
      RECT 47.365 4.88 47.79 5.11 ;
      RECT 45.445 4.32 45.735 4.55 ;
      RECT 45.445 4.32 45.9 4.505 ;
      RECT 45.76 3.845 45.9 4.505 ;
      RECT 45.88 3.245 46.02 3.985 ;
      RECT 46.75 3.185 47.07 3.445 ;
      RECT 45.925 3.2 46.215 3.43 ;
      RECT 45.88 3.245 47.07 3.385 ;
      RECT 46.63 3.745 46.95 4.005 ;
      RECT 46.165 3.76 46.455 3.99 ;
      RECT 46.165 3.805 46.95 3.945 ;
      RECT 46.39 4.305 46.71 4.565 ;
      RECT 46.39 4.32 46.935 4.55 ;
      RECT 45.925 4.88 46.215 5.11 ;
      RECT 45.04 4.76 46.14 4.9 ;
      RECT 44.965 4.6 45.255 4.83 ;
      RECT 42.4 10.06 42.695 10.29 ;
      RECT 42.46 8.58 42.63 10.29 ;
      RECT 42.455 8.95 42.805 9.3 ;
      RECT 42.4 8.58 42.69 8.81 ;
      RECT 41.41 10.06 41.705 10.29 ;
      RECT 41.47 8.58 41.64 10.29 ;
      RECT 41.41 8.58 41.7 8.81 ;
      RECT 41.41 8.615 42.26 8.775 ;
      RECT 42.095 8.21 42.26 8.775 ;
      RECT 41.41 8.61 41.805 8.775 ;
      RECT 42.03 8.21 42.32 8.44 ;
      RECT 42.03 8.24 42.49 8.41 ;
      RECT 41.995 4.025 42.315 4.26 ;
      RECT 41.995 4.055 42.485 4.225 ;
      RECT 41.995 3.69 42.185 4.26 ;
      RECT 41.41 3.655 41.7 3.885 ;
      RECT 41.41 3.69 42.185 3.86 ;
      RECT 41.47 2.175 41.64 3.885 ;
      RECT 41.41 2.175 41.705 2.405 ;
      RECT 41.04 4.025 41.33 4.255 ;
      RECT 41.04 4.055 41.5 4.225 ;
      RECT 41.105 2.95 41.27 4.255 ;
      RECT 39.62 2.915 39.91 3.145 ;
      RECT 39.62 2.95 41.27 3.12 ;
      RECT 39.68 2.175 39.85 3.145 ;
      RECT 39.62 2.175 39.91 2.405 ;
      RECT 39.62 10.06 39.91 10.29 ;
      RECT 39.68 9.32 39.85 10.29 ;
      RECT 39.68 9.41 41.27 9.58 ;
      RECT 41.1 8.21 41.27 9.58 ;
      RECT 39.62 9.32 39.91 9.55 ;
      RECT 41.04 8.21 41.33 8.44 ;
      RECT 41.04 8.24 41.5 8.41 ;
      RECT 37.67 3.995 38.01 4.345 ;
      RECT 37.76 3.32 37.93 4.345 ;
      RECT 40.05 3.26 40.4 3.61 ;
      RECT 37.76 3.32 40.4 3.49 ;
      RECT 39.88 3.315 40.4 3.49 ;
      RECT 40.075 8.945 40.4 9.27 ;
      RECT 34.635 8.895 34.985 9.245 ;
      RECT 40.05 8.95 40.4 9.18 ;
      RECT 34.435 8.95 34.985 9.18 ;
      RECT 39.88 8.975 40.4 9.15 ;
      RECT 34.265 8.98 34.985 9.15 ;
      RECT 34.325 8.975 40.4 9.145 ;
      RECT 39.275 3.66 39.595 3.98 ;
      RECT 39.25 3.655 39.54 3.885 ;
      RECT 39.24 3.685 39.595 3.86 ;
      RECT 39.075 3.685 39.595 3.855 ;
      RECT 39.275 8.545 39.595 8.835 ;
      RECT 39.25 8.58 39.595 8.81 ;
      RECT 39.075 8.61 39.595 8.78 ;
      RECT 36.38 3.185 36.7 3.445 ;
      RECT 35.945 3.2 36.235 3.43 ;
      RECT 35.945 3.245 36.7 3.385 ;
      RECT 36.38 4.865 36.7 5.125 ;
      RECT 35.945 4.88 36.235 5.11 ;
      RECT 35.945 4.925 36.7 5.065 ;
      RECT 35.705 4.32 35.995 4.55 ;
      RECT 35.705 4.365 36.28 4.505 ;
      RECT 36.14 4.225 36.4 4.365 ;
      RECT 36.185 4.04 36.475 4.27 ;
      RECT 34.34 4.225 35.44 4.365 ;
      RECT 34.145 4.025 34.465 4.285 ;
      RECT 35.225 4.04 35.515 4.27 ;
      RECT 34.145 4.04 34.555 4.285 ;
      RECT 34.52 3.185 34.84 3.445 ;
      RECT 34.985 3.2 35.275 3.43 ;
      RECT 34.52 3.245 35.275 3.385 ;
      RECT 32.135 4.365 32.31 4.69 ;
      RECT 31.82 4.45 34 4.59 ;
      RECT 33.86 3.46 34 4.59 ;
      RECT 31.82 4.365 33.115 4.59 ;
      RECT 32.825 4.32 33.115 4.59 ;
      RECT 31.82 4.085 32.155 4.59 ;
      RECT 31.865 4.04 32.155 4.59 ;
      RECT 34.745 3.76 35.035 3.99 ;
      RECT 33.86 3.665 34.96 3.805 ;
      RECT 33.785 3.46 34.075 3.71 ;
      RECT 34.005 10.06 34.295 10.29 ;
      RECT 34.065 9.32 34.235 10.29 ;
      RECT 33.965 9.345 34.335 9.715 ;
      RECT 34.005 9.32 34.295 9.715 ;
      RECT 33.77 4.865 34.095 5.125 ;
      RECT 33.77 4.88 34.29 5.11 ;
      RECT 32.345 3.76 32.635 3.99 ;
      RECT 32.495 3.365 32.635 3.99 ;
      RECT 32.495 3.365 32.8 3.505 ;
      RECT 33.29 3.185 33.61 3.445 ;
      RECT 32.57 3.185 32.89 3.445 ;
      RECT 33.065 3.2 33.61 3.43 ;
      RECT 32.57 3.245 33.61 3.385 ;
      RECT 32.21 4.865 32.53 5.125 ;
      RECT 32.105 4.88 32.53 5.11 ;
      RECT 30.185 4.32 30.475 4.55 ;
      RECT 30.185 4.32 30.64 4.505 ;
      RECT 30.5 3.845 30.64 4.505 ;
      RECT 30.62 3.245 30.76 3.985 ;
      RECT 31.49 3.185 31.81 3.445 ;
      RECT 30.665 3.2 30.955 3.43 ;
      RECT 30.62 3.245 31.81 3.385 ;
      RECT 31.37 3.745 31.69 4.005 ;
      RECT 30.905 3.76 31.195 3.99 ;
      RECT 30.905 3.805 31.69 3.945 ;
      RECT 31.13 4.305 31.45 4.565 ;
      RECT 31.13 4.32 31.675 4.55 ;
      RECT 30.665 4.88 30.955 5.11 ;
      RECT 29.78 4.76 30.88 4.9 ;
      RECT 29.705 4.6 29.995 4.83 ;
      RECT 26.49 10.06 26.78 10.29 ;
      RECT 26.55 9.315 26.72 10.29 ;
      RECT 26.46 9.315 26.81 9.605 ;
      RECT 26.085 8.575 26.435 8.865 ;
      RECT 25.945 8.61 26.435 8.78 ;
      RECT 103.415 7.25 103.765 7.54 ;
      RECT 96.73 3.745 97.05 4.005 ;
      RECT 95.56 4.585 95.88 4.845 ;
      RECT 94.33 4.025 94.65 4.285 ;
      RECT 93.85 3.745 94.17 4.005 ;
      RECT 92.995 3.185 93.395 3.445 ;
      RECT 92.65 4.865 92.97 5.125 ;
      RECT 90.97 3.745 91.29 4.005 ;
      RECT 90.49 4.025 90.81 4.285 ;
      RECT 89.795 3.185 90.12 3.445 ;
      RECT 89.8 4.585 90.12 4.845 ;
      RECT 88.155 7.25 88.505 7.54 ;
      RECT 81.47 3.745 81.79 4.005 ;
      RECT 80.3 4.585 80.62 4.845 ;
      RECT 79.07 4.025 79.39 4.285 ;
      RECT 78.59 3.745 78.91 4.005 ;
      RECT 77.735 3.185 78.135 3.445 ;
      RECT 77.39 4.865 77.71 5.125 ;
      RECT 75.71 3.745 76.03 4.005 ;
      RECT 75.23 4.025 75.55 4.285 ;
      RECT 74.535 3.185 74.86 3.445 ;
      RECT 74.54 4.585 74.86 4.845 ;
      RECT 72.895 7.25 73.245 7.54 ;
      RECT 66.21 3.745 66.53 4.005 ;
      RECT 65.04 4.585 65.36 4.845 ;
      RECT 63.81 4.025 64.13 4.285 ;
      RECT 63.33 3.745 63.65 4.005 ;
      RECT 62.475 3.185 62.875 3.445 ;
      RECT 62.13 4.865 62.45 5.125 ;
      RECT 60.45 3.745 60.77 4.005 ;
      RECT 59.97 4.025 60.29 4.285 ;
      RECT 59.275 3.185 59.6 3.445 ;
      RECT 59.28 4.585 59.6 4.845 ;
      RECT 57.635 7.25 57.985 7.54 ;
      RECT 50.95 3.745 51.27 4.005 ;
      RECT 49.78 4.585 50.1 4.845 ;
      RECT 48.55 4.025 48.87 4.285 ;
      RECT 48.07 3.745 48.39 4.005 ;
      RECT 47.215 3.185 47.615 3.445 ;
      RECT 46.87 4.865 47.19 5.125 ;
      RECT 45.19 3.745 45.51 4.005 ;
      RECT 44.71 4.025 45.03 4.285 ;
      RECT 44.015 3.185 44.34 3.445 ;
      RECT 44.02 4.585 44.34 4.845 ;
      RECT 42.375 7.25 42.725 7.54 ;
      RECT 35.69 3.745 36.01 4.005 ;
      RECT 34.52 4.585 34.84 4.845 ;
      RECT 33.29 4.025 33.61 4.285 ;
      RECT 32.81 3.745 33.13 4.005 ;
      RECT 31.955 3.185 32.355 3.445 ;
      RECT 31.61 4.865 31.93 5.125 ;
      RECT 29.93 3.745 30.25 4.005 ;
      RECT 29.45 4.025 29.77 4.285 ;
      RECT 28.755 3.185 29.08 3.445 ;
      RECT 28.76 4.585 29.08 4.845 ;
    LAYER mcon ;
      RECT 103.505 7.31 103.675 7.48 ;
      RECT 103.5 8.61 103.67 8.78 ;
      RECT 103.5 10.09 103.67 10.26 ;
      RECT 103.13 8.24 103.3 8.41 ;
      RECT 103.125 4.055 103.295 4.225 ;
      RECT 102.51 2.205 102.68 2.375 ;
      RECT 102.51 3.685 102.68 3.855 ;
      RECT 102.51 8.61 102.68 8.78 ;
      RECT 102.51 10.09 102.68 10.26 ;
      RECT 102.14 4.055 102.31 4.225 ;
      RECT 102.14 8.24 102.31 8.41 ;
      RECT 101.15 3.315 101.32 3.485 ;
      RECT 101.15 8.98 101.32 9.15 ;
      RECT 100.72 2.205 100.89 2.375 ;
      RECT 100.72 2.945 100.89 3.115 ;
      RECT 100.72 9.35 100.89 9.52 ;
      RECT 100.72 10.09 100.89 10.26 ;
      RECT 100.35 3.685 100.52 3.855 ;
      RECT 100.35 8.61 100.52 8.78 ;
      RECT 97.285 4.07 97.455 4.24 ;
      RECT 97.045 3.23 97.215 3.4 ;
      RECT 97.045 4.91 97.215 5.08 ;
      RECT 96.805 3.79 96.975 3.96 ;
      RECT 96.805 4.35 96.975 4.52 ;
      RECT 96.325 4.07 96.495 4.24 ;
      RECT 96.085 3.23 96.255 3.4 ;
      RECT 95.845 3.79 96.015 3.96 ;
      RECT 95.635 4.63 95.805 4.8 ;
      RECT 95.535 8.98 95.705 9.15 ;
      RECT 95.365 4.07 95.535 4.24 ;
      RECT 95.105 9.35 95.275 9.52 ;
      RECT 95.105 10.09 95.275 10.26 ;
      RECT 95.1 4.91 95.27 5.08 ;
      RECT 94.885 3.49 95.055 3.66 ;
      RECT 94.405 4.07 94.575 4.24 ;
      RECT 94.165 3.23 94.335 3.4 ;
      RECT 93.925 3.79 94.095 3.96 ;
      RECT 93.925 4.35 94.095 4.52 ;
      RECT 93.445 3.79 93.615 3.96 ;
      RECT 93.205 4.91 93.375 5.08 ;
      RECT 93.165 3.23 93.335 3.4 ;
      RECT 92.965 4.07 93.135 4.24 ;
      RECT 92.725 4.91 92.895 5.08 ;
      RECT 92.485 4.35 92.655 4.52 ;
      RECT 92.005 3.79 92.175 3.96 ;
      RECT 91.765 3.23 91.935 3.4 ;
      RECT 91.765 4.91 91.935 5.08 ;
      RECT 91.285 4.35 91.455 4.52 ;
      RECT 91.045 3.79 91.215 3.96 ;
      RECT 90.805 4.63 90.975 4.8 ;
      RECT 90.565 4.07 90.735 4.24 ;
      RECT 89.87 3.23 90.04 3.4 ;
      RECT 89.87 4.63 90.04 4.8 ;
      RECT 88.245 7.31 88.415 7.48 ;
      RECT 88.24 8.61 88.41 8.78 ;
      RECT 88.24 10.09 88.41 10.26 ;
      RECT 87.87 8.24 88.04 8.41 ;
      RECT 87.865 4.055 88.035 4.225 ;
      RECT 87.25 2.205 87.42 2.375 ;
      RECT 87.25 3.685 87.42 3.855 ;
      RECT 87.25 8.61 87.42 8.78 ;
      RECT 87.25 10.09 87.42 10.26 ;
      RECT 86.88 4.055 87.05 4.225 ;
      RECT 86.88 8.24 87.05 8.41 ;
      RECT 85.89 3.315 86.06 3.485 ;
      RECT 85.89 8.98 86.06 9.15 ;
      RECT 85.46 2.205 85.63 2.375 ;
      RECT 85.46 2.945 85.63 3.115 ;
      RECT 85.46 9.35 85.63 9.52 ;
      RECT 85.46 10.09 85.63 10.26 ;
      RECT 85.09 3.685 85.26 3.855 ;
      RECT 85.09 8.61 85.26 8.78 ;
      RECT 82.025 4.07 82.195 4.24 ;
      RECT 81.785 3.23 81.955 3.4 ;
      RECT 81.785 4.91 81.955 5.08 ;
      RECT 81.545 3.79 81.715 3.96 ;
      RECT 81.545 4.35 81.715 4.52 ;
      RECT 81.065 4.07 81.235 4.24 ;
      RECT 80.825 3.23 80.995 3.4 ;
      RECT 80.585 3.79 80.755 3.96 ;
      RECT 80.375 4.63 80.545 4.8 ;
      RECT 80.275 8.98 80.445 9.15 ;
      RECT 80.105 4.07 80.275 4.24 ;
      RECT 79.845 9.35 80.015 9.52 ;
      RECT 79.845 10.09 80.015 10.26 ;
      RECT 79.84 4.91 80.01 5.08 ;
      RECT 79.625 3.49 79.795 3.66 ;
      RECT 79.145 4.07 79.315 4.24 ;
      RECT 78.905 3.23 79.075 3.4 ;
      RECT 78.665 3.79 78.835 3.96 ;
      RECT 78.665 4.35 78.835 4.52 ;
      RECT 78.185 3.79 78.355 3.96 ;
      RECT 77.945 4.91 78.115 5.08 ;
      RECT 77.905 3.23 78.075 3.4 ;
      RECT 77.705 4.07 77.875 4.24 ;
      RECT 77.465 4.91 77.635 5.08 ;
      RECT 77.225 4.35 77.395 4.52 ;
      RECT 76.745 3.79 76.915 3.96 ;
      RECT 76.505 3.23 76.675 3.4 ;
      RECT 76.505 4.91 76.675 5.08 ;
      RECT 76.025 4.35 76.195 4.52 ;
      RECT 75.785 3.79 75.955 3.96 ;
      RECT 75.545 4.63 75.715 4.8 ;
      RECT 75.305 4.07 75.475 4.24 ;
      RECT 74.61 3.23 74.78 3.4 ;
      RECT 74.61 4.63 74.78 4.8 ;
      RECT 72.985 7.31 73.155 7.48 ;
      RECT 72.98 8.61 73.15 8.78 ;
      RECT 72.98 10.09 73.15 10.26 ;
      RECT 72.61 8.24 72.78 8.41 ;
      RECT 72.605 4.055 72.775 4.225 ;
      RECT 71.99 2.205 72.16 2.375 ;
      RECT 71.99 3.685 72.16 3.855 ;
      RECT 71.99 8.61 72.16 8.78 ;
      RECT 71.99 10.09 72.16 10.26 ;
      RECT 71.62 4.055 71.79 4.225 ;
      RECT 71.62 8.24 71.79 8.41 ;
      RECT 70.63 3.315 70.8 3.485 ;
      RECT 70.63 8.98 70.8 9.15 ;
      RECT 70.2 2.205 70.37 2.375 ;
      RECT 70.2 2.945 70.37 3.115 ;
      RECT 70.2 9.35 70.37 9.52 ;
      RECT 70.2 10.09 70.37 10.26 ;
      RECT 69.83 3.685 70 3.855 ;
      RECT 69.83 8.61 70 8.78 ;
      RECT 66.765 4.07 66.935 4.24 ;
      RECT 66.525 3.23 66.695 3.4 ;
      RECT 66.525 4.91 66.695 5.08 ;
      RECT 66.285 3.79 66.455 3.96 ;
      RECT 66.285 4.35 66.455 4.52 ;
      RECT 65.805 4.07 65.975 4.24 ;
      RECT 65.565 3.23 65.735 3.4 ;
      RECT 65.325 3.79 65.495 3.96 ;
      RECT 65.115 4.63 65.285 4.8 ;
      RECT 65.015 8.98 65.185 9.15 ;
      RECT 64.845 4.07 65.015 4.24 ;
      RECT 64.585 9.35 64.755 9.52 ;
      RECT 64.585 10.09 64.755 10.26 ;
      RECT 64.58 4.91 64.75 5.08 ;
      RECT 64.365 3.49 64.535 3.66 ;
      RECT 63.885 4.07 64.055 4.24 ;
      RECT 63.645 3.23 63.815 3.4 ;
      RECT 63.405 3.79 63.575 3.96 ;
      RECT 63.405 4.35 63.575 4.52 ;
      RECT 62.925 3.79 63.095 3.96 ;
      RECT 62.685 4.91 62.855 5.08 ;
      RECT 62.645 3.23 62.815 3.4 ;
      RECT 62.445 4.07 62.615 4.24 ;
      RECT 62.205 4.91 62.375 5.08 ;
      RECT 61.965 4.35 62.135 4.52 ;
      RECT 61.485 3.79 61.655 3.96 ;
      RECT 61.245 3.23 61.415 3.4 ;
      RECT 61.245 4.91 61.415 5.08 ;
      RECT 60.765 4.35 60.935 4.52 ;
      RECT 60.525 3.79 60.695 3.96 ;
      RECT 60.285 4.63 60.455 4.8 ;
      RECT 60.045 4.07 60.215 4.24 ;
      RECT 59.35 3.23 59.52 3.4 ;
      RECT 59.35 4.63 59.52 4.8 ;
      RECT 57.725 7.31 57.895 7.48 ;
      RECT 57.72 8.61 57.89 8.78 ;
      RECT 57.72 10.09 57.89 10.26 ;
      RECT 57.35 8.24 57.52 8.41 ;
      RECT 57.345 4.055 57.515 4.225 ;
      RECT 56.73 2.205 56.9 2.375 ;
      RECT 56.73 3.685 56.9 3.855 ;
      RECT 56.73 8.61 56.9 8.78 ;
      RECT 56.73 10.09 56.9 10.26 ;
      RECT 56.36 4.055 56.53 4.225 ;
      RECT 56.36 8.24 56.53 8.41 ;
      RECT 55.37 3.315 55.54 3.485 ;
      RECT 55.37 8.98 55.54 9.15 ;
      RECT 54.94 2.205 55.11 2.375 ;
      RECT 54.94 2.945 55.11 3.115 ;
      RECT 54.94 9.35 55.11 9.52 ;
      RECT 54.94 10.09 55.11 10.26 ;
      RECT 54.57 3.685 54.74 3.855 ;
      RECT 54.57 8.61 54.74 8.78 ;
      RECT 51.505 4.07 51.675 4.24 ;
      RECT 51.265 3.23 51.435 3.4 ;
      RECT 51.265 4.91 51.435 5.08 ;
      RECT 51.025 3.79 51.195 3.96 ;
      RECT 51.025 4.35 51.195 4.52 ;
      RECT 50.545 4.07 50.715 4.24 ;
      RECT 50.305 3.23 50.475 3.4 ;
      RECT 50.065 3.79 50.235 3.96 ;
      RECT 49.855 4.63 50.025 4.8 ;
      RECT 49.755 8.98 49.925 9.15 ;
      RECT 49.585 4.07 49.755 4.24 ;
      RECT 49.325 9.35 49.495 9.52 ;
      RECT 49.325 10.09 49.495 10.26 ;
      RECT 49.32 4.91 49.49 5.08 ;
      RECT 49.105 3.49 49.275 3.66 ;
      RECT 48.625 4.07 48.795 4.24 ;
      RECT 48.385 3.23 48.555 3.4 ;
      RECT 48.145 3.79 48.315 3.96 ;
      RECT 48.145 4.35 48.315 4.52 ;
      RECT 47.665 3.79 47.835 3.96 ;
      RECT 47.425 4.91 47.595 5.08 ;
      RECT 47.385 3.23 47.555 3.4 ;
      RECT 47.185 4.07 47.355 4.24 ;
      RECT 46.945 4.91 47.115 5.08 ;
      RECT 46.705 4.35 46.875 4.52 ;
      RECT 46.225 3.79 46.395 3.96 ;
      RECT 45.985 3.23 46.155 3.4 ;
      RECT 45.985 4.91 46.155 5.08 ;
      RECT 45.505 4.35 45.675 4.52 ;
      RECT 45.265 3.79 45.435 3.96 ;
      RECT 45.025 4.63 45.195 4.8 ;
      RECT 44.785 4.07 44.955 4.24 ;
      RECT 44.09 3.23 44.26 3.4 ;
      RECT 44.09 4.63 44.26 4.8 ;
      RECT 42.465 7.31 42.635 7.48 ;
      RECT 42.46 8.61 42.63 8.78 ;
      RECT 42.46 10.09 42.63 10.26 ;
      RECT 42.09 8.24 42.26 8.41 ;
      RECT 42.085 4.055 42.255 4.225 ;
      RECT 41.47 2.205 41.64 2.375 ;
      RECT 41.47 3.685 41.64 3.855 ;
      RECT 41.47 8.61 41.64 8.78 ;
      RECT 41.47 10.09 41.64 10.26 ;
      RECT 41.1 4.055 41.27 4.225 ;
      RECT 41.1 8.24 41.27 8.41 ;
      RECT 40.11 3.315 40.28 3.485 ;
      RECT 40.11 8.98 40.28 9.15 ;
      RECT 39.68 2.205 39.85 2.375 ;
      RECT 39.68 2.945 39.85 3.115 ;
      RECT 39.68 9.35 39.85 9.52 ;
      RECT 39.68 10.09 39.85 10.26 ;
      RECT 39.31 3.685 39.48 3.855 ;
      RECT 39.31 8.61 39.48 8.78 ;
      RECT 36.245 4.07 36.415 4.24 ;
      RECT 36.005 3.23 36.175 3.4 ;
      RECT 36.005 4.91 36.175 5.08 ;
      RECT 35.765 3.79 35.935 3.96 ;
      RECT 35.765 4.35 35.935 4.52 ;
      RECT 35.285 4.07 35.455 4.24 ;
      RECT 35.045 3.23 35.215 3.4 ;
      RECT 34.805 3.79 34.975 3.96 ;
      RECT 34.595 4.63 34.765 4.8 ;
      RECT 34.495 8.98 34.665 9.15 ;
      RECT 34.325 4.07 34.495 4.24 ;
      RECT 34.065 9.35 34.235 9.52 ;
      RECT 34.065 10.09 34.235 10.26 ;
      RECT 34.06 4.91 34.23 5.08 ;
      RECT 33.845 3.49 34.015 3.66 ;
      RECT 33.365 4.07 33.535 4.24 ;
      RECT 33.125 3.23 33.295 3.4 ;
      RECT 32.885 3.79 33.055 3.96 ;
      RECT 32.885 4.35 33.055 4.52 ;
      RECT 32.405 3.79 32.575 3.96 ;
      RECT 32.165 4.91 32.335 5.08 ;
      RECT 32.125 3.23 32.295 3.4 ;
      RECT 31.925 4.07 32.095 4.24 ;
      RECT 31.685 4.91 31.855 5.08 ;
      RECT 31.445 4.35 31.615 4.52 ;
      RECT 30.965 3.79 31.135 3.96 ;
      RECT 30.725 3.23 30.895 3.4 ;
      RECT 30.725 4.91 30.895 5.08 ;
      RECT 30.245 4.35 30.415 4.52 ;
      RECT 30.005 3.79 30.175 3.96 ;
      RECT 29.765 4.63 29.935 4.8 ;
      RECT 29.525 4.07 29.695 4.24 ;
      RECT 28.83 3.23 29 3.4 ;
      RECT 28.83 4.63 29 4.8 ;
      RECT 26.55 9.35 26.72 9.52 ;
      RECT 26.55 10.09 26.72 10.26 ;
      RECT 26.18 8.61 26.35 8.78 ;
    LAYER li1 ;
      RECT 103.5 7.31 103.67 8.78 ;
      RECT 103.5 7.31 103.675 8.57 ;
      RECT 103.13 9.26 103.6 9.43 ;
      RECT 103.13 8.24 103.3 9.43 ;
      RECT 103.125 3.035 103.295 4.225 ;
      RECT 103.125 3.035 103.595 3.205 ;
      RECT 102.51 3.895 102.685 5.155 ;
      RECT 102.51 3.685 102.68 5.155 ;
      RECT 102.51 7.31 102.68 8.78 ;
      RECT 102.51 7.31 102.685 8.57 ;
      RECT 102.14 3.035 102.31 4.225 ;
      RECT 102.14 3.035 102.61 3.205 ;
      RECT 102.14 9.26 102.61 9.43 ;
      RECT 102.14 8.24 102.31 9.43 ;
      RECT 101.15 4.015 101.325 5.155 ;
      RECT 101.15 1.865 101.32 5.155 ;
      RECT 101.15 1.865 101.325 2.415 ;
      RECT 101.15 10.05 101.325 10.6 ;
      RECT 101.15 7.31 101.32 10.6 ;
      RECT 101.15 7.31 101.325 8.45 ;
      RECT 100.72 3.895 100.895 5.155 ;
      RECT 100.72 2.945 100.89 5.155 ;
      RECT 100.72 7.31 100.89 9.52 ;
      RECT 100.72 7.31 100.895 8.57 ;
      RECT 100.29 3.925 100.46 5.155 ;
      RECT 100.35 2.145 100.52 4.095 ;
      RECT 100.29 1.865 100.46 2.315 ;
      RECT 100.29 10.15 100.46 10.6 ;
      RECT 100.35 8.37 100.52 10.32 ;
      RECT 100.29 7.31 100.46 8.54 ;
      RECT 99.765 3.895 99.94 5.155 ;
      RECT 99.765 1.865 99.935 5.155 ;
      RECT 99.765 3.365 100.175 3.695 ;
      RECT 99.765 2.525 100.175 2.855 ;
      RECT 99.765 1.865 99.94 2.355 ;
      RECT 99.765 10.11 99.94 10.6 ;
      RECT 99.765 7.31 99.935 10.6 ;
      RECT 99.765 9.61 100.175 9.94 ;
      RECT 99.765 8.77 100.175 9.1 ;
      RECT 99.765 7.31 99.94 8.57 ;
      RECT 97.045 4.91 97.56 5.08 ;
      RECT 97.39 4.52 97.56 5.08 ;
      RECT 97.495 4.44 97.67 4.77 ;
      RECT 97.285 3.83 97.56 4.24 ;
      RECT 97.165 3.83 97.56 4.04 ;
      RECT 95.63 4.44 95.805 4.8 ;
      RECT 95.63 4.52 96.975 4.69 ;
      RECT 96.805 4.35 96.975 4.69 ;
      RECT 95.535 10.05 95.71 10.6 ;
      RECT 95.535 7.31 95.705 10.6 ;
      RECT 95.535 7.31 95.71 8.45 ;
      RECT 95.365 3.87 95.535 4.24 ;
      RECT 94.885 3.87 95.535 4.14 ;
      RECT 94.805 3.87 95.615 4.04 ;
      RECT 94.165 3.11 94.335 3.4 ;
      RECT 94.165 3.11 95.405 3.28 ;
      RECT 95.105 7.31 95.275 9.52 ;
      RECT 95.105 7.31 95.28 8.57 ;
      RECT 94.885 3.45 95.055 3.66 ;
      RECT 94.525 3.45 95.055 3.62 ;
      RECT 94.15 10.11 94.325 10.6 ;
      RECT 94.15 7.31 94.32 10.6 ;
      RECT 94.15 9.61 94.56 9.94 ;
      RECT 94.15 8.77 94.56 9.1 ;
      RECT 94.15 7.31 94.325 8.57 ;
      RECT 93.925 4.52 94.415 4.69 ;
      RECT 93.925 4.35 94.095 4.69 ;
      RECT 93.205 4.52 93.375 5.08 ;
      RECT 93.1 4.52 93.43 4.69 ;
      RECT 93.165 3.13 93.335 3.4 ;
      RECT 93.205 3.05 93.375 3.38 ;
      RECT 93.07 3.13 93.375 3.35 ;
      RECT 91.645 4.52 91.935 5.08 ;
      RECT 91.765 4.44 91.935 5.08 ;
      RECT 88.24 7.31 88.41 8.78 ;
      RECT 88.24 7.31 88.415 8.57 ;
      RECT 87.87 9.26 88.34 9.43 ;
      RECT 87.87 8.24 88.04 9.43 ;
      RECT 87.865 3.035 88.035 4.225 ;
      RECT 87.865 3.035 88.335 3.205 ;
      RECT 87.25 3.895 87.425 5.155 ;
      RECT 87.25 3.685 87.42 5.155 ;
      RECT 87.25 7.31 87.42 8.78 ;
      RECT 87.25 7.31 87.425 8.57 ;
      RECT 86.88 3.035 87.05 4.225 ;
      RECT 86.88 3.035 87.35 3.205 ;
      RECT 86.88 9.26 87.35 9.43 ;
      RECT 86.88 8.24 87.05 9.43 ;
      RECT 85.89 4.015 86.065 5.155 ;
      RECT 85.89 1.865 86.06 5.155 ;
      RECT 85.89 1.865 86.065 2.415 ;
      RECT 85.89 10.05 86.065 10.6 ;
      RECT 85.89 7.31 86.06 10.6 ;
      RECT 85.89 7.31 86.065 8.45 ;
      RECT 85.46 3.895 85.635 5.155 ;
      RECT 85.46 2.945 85.63 5.155 ;
      RECT 85.46 7.31 85.63 9.52 ;
      RECT 85.46 7.31 85.635 8.57 ;
      RECT 85.03 3.925 85.2 5.155 ;
      RECT 85.09 2.145 85.26 4.095 ;
      RECT 85.03 1.865 85.2 2.315 ;
      RECT 85.03 10.15 85.2 10.6 ;
      RECT 85.09 8.37 85.26 10.32 ;
      RECT 85.03 7.31 85.2 8.54 ;
      RECT 84.505 3.895 84.68 5.155 ;
      RECT 84.505 1.865 84.675 5.155 ;
      RECT 84.505 3.365 84.915 3.695 ;
      RECT 84.505 2.525 84.915 2.855 ;
      RECT 84.505 1.865 84.68 2.355 ;
      RECT 84.505 10.11 84.68 10.6 ;
      RECT 84.505 7.31 84.675 10.6 ;
      RECT 84.505 9.61 84.915 9.94 ;
      RECT 84.505 8.77 84.915 9.1 ;
      RECT 84.505 7.31 84.68 8.57 ;
      RECT 81.785 4.91 82.3 5.08 ;
      RECT 82.13 4.52 82.3 5.08 ;
      RECT 82.235 4.44 82.41 4.77 ;
      RECT 82.025 3.83 82.3 4.24 ;
      RECT 81.905 3.83 82.3 4.04 ;
      RECT 80.37 4.44 80.545 4.8 ;
      RECT 80.37 4.52 81.715 4.69 ;
      RECT 81.545 4.35 81.715 4.69 ;
      RECT 80.275 10.05 80.45 10.6 ;
      RECT 80.275 7.31 80.445 10.6 ;
      RECT 80.275 7.31 80.45 8.45 ;
      RECT 80.105 3.87 80.275 4.24 ;
      RECT 79.625 3.87 80.275 4.14 ;
      RECT 79.545 3.87 80.355 4.04 ;
      RECT 78.905 3.11 79.075 3.4 ;
      RECT 78.905 3.11 80.145 3.28 ;
      RECT 79.845 7.31 80.015 9.52 ;
      RECT 79.845 7.31 80.02 8.57 ;
      RECT 79.625 3.45 79.795 3.66 ;
      RECT 79.265 3.45 79.795 3.62 ;
      RECT 78.89 10.11 79.065 10.6 ;
      RECT 78.89 7.31 79.06 10.6 ;
      RECT 78.89 9.61 79.3 9.94 ;
      RECT 78.89 8.77 79.3 9.1 ;
      RECT 78.89 7.31 79.065 8.57 ;
      RECT 78.665 4.52 79.155 4.69 ;
      RECT 78.665 4.35 78.835 4.69 ;
      RECT 77.945 4.52 78.115 5.08 ;
      RECT 77.84 4.52 78.17 4.69 ;
      RECT 77.905 3.13 78.075 3.4 ;
      RECT 77.945 3.05 78.115 3.38 ;
      RECT 77.81 3.13 78.115 3.35 ;
      RECT 76.385 4.52 76.675 5.08 ;
      RECT 76.505 4.44 76.675 5.08 ;
      RECT 72.98 7.31 73.15 8.78 ;
      RECT 72.98 7.31 73.155 8.57 ;
      RECT 72.61 9.26 73.08 9.43 ;
      RECT 72.61 8.24 72.78 9.43 ;
      RECT 72.605 3.035 72.775 4.225 ;
      RECT 72.605 3.035 73.075 3.205 ;
      RECT 71.99 3.895 72.165 5.155 ;
      RECT 71.99 3.685 72.16 5.155 ;
      RECT 71.99 7.31 72.16 8.78 ;
      RECT 71.99 7.31 72.165 8.57 ;
      RECT 71.62 3.035 71.79 4.225 ;
      RECT 71.62 3.035 72.09 3.205 ;
      RECT 71.62 9.26 72.09 9.43 ;
      RECT 71.62 8.24 71.79 9.43 ;
      RECT 70.63 4.015 70.805 5.155 ;
      RECT 70.63 1.865 70.8 5.155 ;
      RECT 70.63 1.865 70.805 2.415 ;
      RECT 70.63 10.05 70.805 10.6 ;
      RECT 70.63 7.31 70.8 10.6 ;
      RECT 70.63 7.31 70.805 8.45 ;
      RECT 70.2 3.895 70.375 5.155 ;
      RECT 70.2 2.945 70.37 5.155 ;
      RECT 70.2 7.31 70.37 9.52 ;
      RECT 70.2 7.31 70.375 8.57 ;
      RECT 69.77 3.925 69.94 5.155 ;
      RECT 69.83 2.145 70 4.095 ;
      RECT 69.77 1.865 69.94 2.315 ;
      RECT 69.77 10.15 69.94 10.6 ;
      RECT 69.83 8.37 70 10.32 ;
      RECT 69.77 7.31 69.94 8.54 ;
      RECT 69.245 3.895 69.42 5.155 ;
      RECT 69.245 1.865 69.415 5.155 ;
      RECT 69.245 3.365 69.655 3.695 ;
      RECT 69.245 2.525 69.655 2.855 ;
      RECT 69.245 1.865 69.42 2.355 ;
      RECT 69.245 10.11 69.42 10.6 ;
      RECT 69.245 7.31 69.415 10.6 ;
      RECT 69.245 9.61 69.655 9.94 ;
      RECT 69.245 8.77 69.655 9.1 ;
      RECT 69.245 7.31 69.42 8.57 ;
      RECT 66.525 4.91 67.04 5.08 ;
      RECT 66.87 4.52 67.04 5.08 ;
      RECT 66.975 4.44 67.15 4.77 ;
      RECT 66.765 3.83 67.04 4.24 ;
      RECT 66.645 3.83 67.04 4.04 ;
      RECT 65.11 4.44 65.285 4.8 ;
      RECT 65.11 4.52 66.455 4.69 ;
      RECT 66.285 4.35 66.455 4.69 ;
      RECT 65.015 10.05 65.19 10.6 ;
      RECT 65.015 7.31 65.185 10.6 ;
      RECT 65.015 7.31 65.19 8.45 ;
      RECT 64.845 3.87 65.015 4.24 ;
      RECT 64.365 3.87 65.015 4.14 ;
      RECT 64.285 3.87 65.095 4.04 ;
      RECT 63.645 3.11 63.815 3.4 ;
      RECT 63.645 3.11 64.885 3.28 ;
      RECT 64.585 7.31 64.755 9.52 ;
      RECT 64.585 7.31 64.76 8.57 ;
      RECT 64.365 3.45 64.535 3.66 ;
      RECT 64.005 3.45 64.535 3.62 ;
      RECT 63.63 10.11 63.805 10.6 ;
      RECT 63.63 7.31 63.8 10.6 ;
      RECT 63.63 9.61 64.04 9.94 ;
      RECT 63.63 8.77 64.04 9.1 ;
      RECT 63.63 7.31 63.805 8.57 ;
      RECT 63.405 4.52 63.895 4.69 ;
      RECT 63.405 4.35 63.575 4.69 ;
      RECT 62.685 4.52 62.855 5.08 ;
      RECT 62.58 4.52 62.91 4.69 ;
      RECT 62.645 3.13 62.815 3.4 ;
      RECT 62.685 3.05 62.855 3.38 ;
      RECT 62.55 3.13 62.855 3.35 ;
      RECT 61.125 4.52 61.415 5.08 ;
      RECT 61.245 4.44 61.415 5.08 ;
      RECT 57.72 7.31 57.89 8.78 ;
      RECT 57.72 7.31 57.895 8.57 ;
      RECT 57.35 9.26 57.82 9.43 ;
      RECT 57.35 8.24 57.52 9.43 ;
      RECT 57.345 3.035 57.515 4.225 ;
      RECT 57.345 3.035 57.815 3.205 ;
      RECT 56.73 3.895 56.905 5.155 ;
      RECT 56.73 3.685 56.9 5.155 ;
      RECT 56.73 7.31 56.9 8.78 ;
      RECT 56.73 7.31 56.905 8.57 ;
      RECT 56.36 3.035 56.53 4.225 ;
      RECT 56.36 3.035 56.83 3.205 ;
      RECT 56.36 9.26 56.83 9.43 ;
      RECT 56.36 8.24 56.53 9.43 ;
      RECT 55.37 4.015 55.545 5.155 ;
      RECT 55.37 1.865 55.54 5.155 ;
      RECT 55.37 1.865 55.545 2.415 ;
      RECT 55.37 10.05 55.545 10.6 ;
      RECT 55.37 7.31 55.54 10.6 ;
      RECT 55.37 7.31 55.545 8.45 ;
      RECT 54.94 3.895 55.115 5.155 ;
      RECT 54.94 2.945 55.11 5.155 ;
      RECT 54.94 7.31 55.11 9.52 ;
      RECT 54.94 7.31 55.115 8.57 ;
      RECT 54.51 3.925 54.68 5.155 ;
      RECT 54.57 2.145 54.74 4.095 ;
      RECT 54.51 1.865 54.68 2.315 ;
      RECT 54.51 10.15 54.68 10.6 ;
      RECT 54.57 8.37 54.74 10.32 ;
      RECT 54.51 7.31 54.68 8.54 ;
      RECT 53.985 3.895 54.16 5.155 ;
      RECT 53.985 1.865 54.155 5.155 ;
      RECT 53.985 3.365 54.395 3.695 ;
      RECT 53.985 2.525 54.395 2.855 ;
      RECT 53.985 1.865 54.16 2.355 ;
      RECT 53.985 10.11 54.16 10.6 ;
      RECT 53.985 7.31 54.155 10.6 ;
      RECT 53.985 9.61 54.395 9.94 ;
      RECT 53.985 8.77 54.395 9.1 ;
      RECT 53.985 7.31 54.16 8.57 ;
      RECT 51.265 4.91 51.78 5.08 ;
      RECT 51.61 4.52 51.78 5.08 ;
      RECT 51.715 4.44 51.89 4.77 ;
      RECT 51.505 3.83 51.78 4.24 ;
      RECT 51.385 3.83 51.78 4.04 ;
      RECT 49.85 4.44 50.025 4.8 ;
      RECT 49.85 4.52 51.195 4.69 ;
      RECT 51.025 4.35 51.195 4.69 ;
      RECT 49.755 10.05 49.93 10.6 ;
      RECT 49.755 7.31 49.925 10.6 ;
      RECT 49.755 7.31 49.93 8.45 ;
      RECT 49.585 3.87 49.755 4.24 ;
      RECT 49.105 3.87 49.755 4.14 ;
      RECT 49.025 3.87 49.835 4.04 ;
      RECT 48.385 3.11 48.555 3.4 ;
      RECT 48.385 3.11 49.625 3.28 ;
      RECT 49.325 7.31 49.495 9.52 ;
      RECT 49.325 7.31 49.5 8.57 ;
      RECT 49.105 3.45 49.275 3.66 ;
      RECT 48.745 3.45 49.275 3.62 ;
      RECT 48.37 10.11 48.545 10.6 ;
      RECT 48.37 7.31 48.54 10.6 ;
      RECT 48.37 9.61 48.78 9.94 ;
      RECT 48.37 8.77 48.78 9.1 ;
      RECT 48.37 7.31 48.545 8.57 ;
      RECT 48.145 4.52 48.635 4.69 ;
      RECT 48.145 4.35 48.315 4.69 ;
      RECT 47.425 4.52 47.595 5.08 ;
      RECT 47.32 4.52 47.65 4.69 ;
      RECT 47.385 3.13 47.555 3.4 ;
      RECT 47.425 3.05 47.595 3.38 ;
      RECT 47.29 3.13 47.595 3.35 ;
      RECT 45.865 4.52 46.155 5.08 ;
      RECT 45.985 4.44 46.155 5.08 ;
      RECT 42.46 7.31 42.63 8.78 ;
      RECT 42.46 7.31 42.635 8.57 ;
      RECT 42.09 9.26 42.56 9.43 ;
      RECT 42.09 8.24 42.26 9.43 ;
      RECT 42.085 3.035 42.255 4.225 ;
      RECT 42.085 3.035 42.555 3.205 ;
      RECT 41.47 3.895 41.645 5.155 ;
      RECT 41.47 3.685 41.64 5.155 ;
      RECT 41.47 7.31 41.64 8.78 ;
      RECT 41.47 7.31 41.645 8.57 ;
      RECT 41.1 3.035 41.27 4.225 ;
      RECT 41.1 3.035 41.57 3.205 ;
      RECT 41.1 9.26 41.57 9.43 ;
      RECT 41.1 8.24 41.27 9.43 ;
      RECT 40.11 4.015 40.285 5.155 ;
      RECT 40.11 1.865 40.28 5.155 ;
      RECT 40.11 1.865 40.285 2.415 ;
      RECT 40.11 10.05 40.285 10.6 ;
      RECT 40.11 7.31 40.28 10.6 ;
      RECT 40.11 7.31 40.285 8.45 ;
      RECT 39.68 3.895 39.855 5.155 ;
      RECT 39.68 2.945 39.85 5.155 ;
      RECT 39.68 7.31 39.85 9.52 ;
      RECT 39.68 7.31 39.855 8.57 ;
      RECT 39.25 3.925 39.42 5.155 ;
      RECT 39.31 2.145 39.48 4.095 ;
      RECT 39.25 1.865 39.42 2.315 ;
      RECT 39.25 10.15 39.42 10.6 ;
      RECT 39.31 8.37 39.48 10.32 ;
      RECT 39.25 7.31 39.42 8.54 ;
      RECT 38.725 3.895 38.9 5.155 ;
      RECT 38.725 1.865 38.895 5.155 ;
      RECT 38.725 3.365 39.135 3.695 ;
      RECT 38.725 2.525 39.135 2.855 ;
      RECT 38.725 1.865 38.9 2.355 ;
      RECT 38.725 10.11 38.9 10.6 ;
      RECT 38.725 7.31 38.895 10.6 ;
      RECT 38.725 9.61 39.135 9.94 ;
      RECT 38.725 8.77 39.135 9.1 ;
      RECT 38.725 7.31 38.9 8.57 ;
      RECT 36.005 4.91 36.52 5.08 ;
      RECT 36.35 4.52 36.52 5.08 ;
      RECT 36.455 4.44 36.63 4.77 ;
      RECT 36.245 3.83 36.52 4.24 ;
      RECT 36.125 3.83 36.52 4.04 ;
      RECT 34.59 4.44 34.765 4.8 ;
      RECT 34.59 4.52 35.935 4.69 ;
      RECT 35.765 4.35 35.935 4.69 ;
      RECT 34.495 10.05 34.67 10.6 ;
      RECT 34.495 7.31 34.665 10.6 ;
      RECT 34.495 7.31 34.67 8.45 ;
      RECT 34.325 3.87 34.495 4.24 ;
      RECT 33.845 3.87 34.495 4.14 ;
      RECT 33.765 3.87 34.575 4.04 ;
      RECT 33.125 3.11 33.295 3.4 ;
      RECT 33.125 3.11 34.365 3.28 ;
      RECT 34.065 7.31 34.235 9.52 ;
      RECT 34.065 7.31 34.24 8.57 ;
      RECT 33.845 3.45 34.015 3.66 ;
      RECT 33.485 3.45 34.015 3.62 ;
      RECT 33.11 10.11 33.285 10.6 ;
      RECT 33.11 7.31 33.28 10.6 ;
      RECT 33.11 9.61 33.52 9.94 ;
      RECT 33.11 8.77 33.52 9.1 ;
      RECT 33.11 7.31 33.285 8.57 ;
      RECT 32.885 4.52 33.375 4.69 ;
      RECT 32.885 4.35 33.055 4.69 ;
      RECT 32.165 4.52 32.335 5.08 ;
      RECT 32.06 4.52 32.39 4.69 ;
      RECT 32.125 3.13 32.295 3.4 ;
      RECT 32.165 3.05 32.335 3.38 ;
      RECT 32.03 3.13 32.335 3.35 ;
      RECT 30.605 4.52 30.895 5.08 ;
      RECT 30.725 4.44 30.895 5.08 ;
      RECT 26.55 7.31 26.72 9.52 ;
      RECT 26.55 7.31 26.725 8.57 ;
      RECT 26.12 10.15 26.29 10.6 ;
      RECT 26.18 8.37 26.35 10.32 ;
      RECT 26.12 7.31 26.29 8.54 ;
      RECT 25.595 10.11 25.77 10.6 ;
      RECT 25.595 7.31 25.765 10.6 ;
      RECT 25.595 9.61 26.005 9.94 ;
      RECT 25.595 8.77 26.005 9.1 ;
      RECT 25.595 7.31 25.77 8.57 ;
      RECT 103.5 10.09 103.675 10.6 ;
      RECT 102.51 1.865 102.685 2.375 ;
      RECT 102.51 10.09 102.685 10.6 ;
      RECT 100.72 1.865 100.895 2.375 ;
      RECT 100.72 10.09 100.895 10.6 ;
      RECT 97.045 3.05 97.215 3.4 ;
      RECT 96.805 3.79 96.975 4.12 ;
      RECT 96.325 3.79 96.495 4.24 ;
      RECT 96.085 3.05 96.255 3.4 ;
      RECT 95.845 3.79 96.015 4.12 ;
      RECT 95.105 10.09 95.28 10.6 ;
      RECT 95.1 4.78 95.27 5.11 ;
      RECT 94.405 3.79 94.575 4.24 ;
      RECT 93.925 3.79 94.095 4.12 ;
      RECT 93.445 3.79 93.615 4.12 ;
      RECT 92.965 3.79 93.135 4.24 ;
      RECT 92.725 4.78 92.895 5.11 ;
      RECT 92.485 3.79 92.655 4.52 ;
      RECT 92.005 3.79 92.175 4.12 ;
      RECT 91.765 3.05 91.935 3.4 ;
      RECT 91.285 4.35 91.455 4.77 ;
      RECT 91.045 3.79 91.215 4.12 ;
      RECT 90.805 4.44 90.975 4.8 ;
      RECT 90.565 3.79 90.735 4.24 ;
      RECT 89.87 3.05 90.04 3.4 ;
      RECT 89.87 4.44 90.04 4.8 ;
      RECT 88.24 10.09 88.415 10.6 ;
      RECT 87.25 1.865 87.425 2.375 ;
      RECT 87.25 10.09 87.425 10.6 ;
      RECT 85.46 1.865 85.635 2.375 ;
      RECT 85.46 10.09 85.635 10.6 ;
      RECT 81.785 3.05 81.955 3.4 ;
      RECT 81.545 3.79 81.715 4.12 ;
      RECT 81.065 3.79 81.235 4.24 ;
      RECT 80.825 3.05 80.995 3.4 ;
      RECT 80.585 3.79 80.755 4.12 ;
      RECT 79.845 10.09 80.02 10.6 ;
      RECT 79.84 4.78 80.01 5.11 ;
      RECT 79.145 3.79 79.315 4.24 ;
      RECT 78.665 3.79 78.835 4.12 ;
      RECT 78.185 3.79 78.355 4.12 ;
      RECT 77.705 3.79 77.875 4.24 ;
      RECT 77.465 4.78 77.635 5.11 ;
      RECT 77.225 3.79 77.395 4.52 ;
      RECT 76.745 3.79 76.915 4.12 ;
      RECT 76.505 3.05 76.675 3.4 ;
      RECT 76.025 4.35 76.195 4.77 ;
      RECT 75.785 3.79 75.955 4.12 ;
      RECT 75.545 4.44 75.715 4.8 ;
      RECT 75.305 3.79 75.475 4.24 ;
      RECT 74.61 3.05 74.78 3.4 ;
      RECT 74.61 4.44 74.78 4.8 ;
      RECT 72.98 10.09 73.155 10.6 ;
      RECT 71.99 1.865 72.165 2.375 ;
      RECT 71.99 10.09 72.165 10.6 ;
      RECT 70.2 1.865 70.375 2.375 ;
      RECT 70.2 10.09 70.375 10.6 ;
      RECT 66.525 3.05 66.695 3.4 ;
      RECT 66.285 3.79 66.455 4.12 ;
      RECT 65.805 3.79 65.975 4.24 ;
      RECT 65.565 3.05 65.735 3.4 ;
      RECT 65.325 3.79 65.495 4.12 ;
      RECT 64.585 10.09 64.76 10.6 ;
      RECT 64.58 4.78 64.75 5.11 ;
      RECT 63.885 3.79 64.055 4.24 ;
      RECT 63.405 3.79 63.575 4.12 ;
      RECT 62.925 3.79 63.095 4.12 ;
      RECT 62.445 3.79 62.615 4.24 ;
      RECT 62.205 4.78 62.375 5.11 ;
      RECT 61.965 3.79 62.135 4.52 ;
      RECT 61.485 3.79 61.655 4.12 ;
      RECT 61.245 3.05 61.415 3.4 ;
      RECT 60.765 4.35 60.935 4.77 ;
      RECT 60.525 3.79 60.695 4.12 ;
      RECT 60.285 4.44 60.455 4.8 ;
      RECT 60.045 3.79 60.215 4.24 ;
      RECT 59.35 3.05 59.52 3.4 ;
      RECT 59.35 4.44 59.52 4.8 ;
      RECT 57.72 10.09 57.895 10.6 ;
      RECT 56.73 1.865 56.905 2.375 ;
      RECT 56.73 10.09 56.905 10.6 ;
      RECT 54.94 1.865 55.115 2.375 ;
      RECT 54.94 10.09 55.115 10.6 ;
      RECT 51.265 3.05 51.435 3.4 ;
      RECT 51.025 3.79 51.195 4.12 ;
      RECT 50.545 3.79 50.715 4.24 ;
      RECT 50.305 3.05 50.475 3.4 ;
      RECT 50.065 3.79 50.235 4.12 ;
      RECT 49.325 10.09 49.5 10.6 ;
      RECT 49.32 4.78 49.49 5.11 ;
      RECT 48.625 3.79 48.795 4.24 ;
      RECT 48.145 3.79 48.315 4.12 ;
      RECT 47.665 3.79 47.835 4.12 ;
      RECT 47.185 3.79 47.355 4.24 ;
      RECT 46.945 4.78 47.115 5.11 ;
      RECT 46.705 3.79 46.875 4.52 ;
      RECT 46.225 3.79 46.395 4.12 ;
      RECT 45.985 3.05 46.155 3.4 ;
      RECT 45.505 4.35 45.675 4.77 ;
      RECT 45.265 3.79 45.435 4.12 ;
      RECT 45.025 4.44 45.195 4.8 ;
      RECT 44.785 3.79 44.955 4.24 ;
      RECT 44.09 3.05 44.26 3.4 ;
      RECT 44.09 4.44 44.26 4.8 ;
      RECT 42.46 10.09 42.635 10.6 ;
      RECT 41.47 1.865 41.645 2.375 ;
      RECT 41.47 10.09 41.645 10.6 ;
      RECT 39.68 1.865 39.855 2.375 ;
      RECT 39.68 10.09 39.855 10.6 ;
      RECT 36.005 3.05 36.175 3.4 ;
      RECT 35.765 3.79 35.935 4.12 ;
      RECT 35.285 3.79 35.455 4.24 ;
      RECT 35.045 3.05 35.215 3.4 ;
      RECT 34.805 3.79 34.975 4.12 ;
      RECT 34.065 10.09 34.24 10.6 ;
      RECT 34.06 4.78 34.23 5.11 ;
      RECT 33.365 3.79 33.535 4.24 ;
      RECT 32.885 3.79 33.055 4.12 ;
      RECT 32.405 3.79 32.575 4.12 ;
      RECT 31.925 3.79 32.095 4.24 ;
      RECT 31.685 4.78 31.855 5.11 ;
      RECT 31.445 3.79 31.615 4.52 ;
      RECT 30.965 3.79 31.135 4.12 ;
      RECT 30.725 3.05 30.895 3.4 ;
      RECT 30.245 4.35 30.415 4.77 ;
      RECT 30.005 3.79 30.175 4.12 ;
      RECT 29.765 4.44 29.935 4.8 ;
      RECT 29.525 3.79 29.695 4.24 ;
      RECT 28.83 3.05 29 3.4 ;
      RECT 28.83 4.44 29 4.8 ;
      RECT 26.55 10.09 26.725 10.6 ;
  END
END sky130_osu_ring_oscillator_mpr2xa_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2xa_8_b0r2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2xa_8_b0r2 ;
  SIZE 104.095 BY 12.465 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 42.405 0 42.785 5.26 ;
      LAYER met2 ;
        RECT 42.405 4.88 42.785 5.26 ;
      LAYER li1 ;
        RECT 42.505 1.865 42.68 2.375 ;
        RECT 42.505 3.895 42.68 5.155 ;
        RECT 42.505 3.685 42.675 5.155 ;
      LAYER met1 ;
        RECT 42.42 4.925 42.77 5.215 ;
        RECT 42.445 2.175 42.74 2.405 ;
        RECT 42.445 3.655 42.735 3.885 ;
        RECT 42.505 2.175 42.675 3.885 ;
      LAYER via1 ;
        RECT 42.52 4.995 42.67 5.145 ;
      LAYER via2 ;
        RECT 42.495 4.97 42.695 5.17 ;
      LAYER mcon ;
        RECT 42.505 3.685 42.675 3.855 ;
        RECT 42.505 2.205 42.675 2.375 ;
        RECT 42.51 4.985 42.68 5.155 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 57.665 0 58.045 5.26 ;
      LAYER met2 ;
        RECT 57.665 4.88 58.045 5.26 ;
      LAYER li1 ;
        RECT 57.765 1.865 57.94 2.375 ;
        RECT 57.765 3.895 57.94 5.155 ;
        RECT 57.765 3.685 57.935 5.155 ;
      LAYER met1 ;
        RECT 57.68 4.925 58.03 5.215 ;
        RECT 57.705 2.175 58 2.405 ;
        RECT 57.705 3.655 57.995 3.885 ;
        RECT 57.765 2.175 57.935 3.885 ;
      LAYER via1 ;
        RECT 57.78 4.995 57.93 5.145 ;
      LAYER via2 ;
        RECT 57.755 4.97 57.955 5.17 ;
      LAYER mcon ;
        RECT 57.765 3.685 57.935 3.855 ;
        RECT 57.765 2.205 57.935 2.375 ;
        RECT 57.77 4.985 57.94 5.155 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 72.925 0 73.305 5.26 ;
      LAYER met2 ;
        RECT 72.925 4.88 73.305 5.26 ;
      LAYER li1 ;
        RECT 73.025 1.865 73.2 2.375 ;
        RECT 73.025 3.895 73.2 5.155 ;
        RECT 73.025 3.685 73.195 5.155 ;
      LAYER met1 ;
        RECT 72.94 4.925 73.29 5.215 ;
        RECT 72.965 2.175 73.26 2.405 ;
        RECT 72.965 3.655 73.255 3.885 ;
        RECT 73.025 2.175 73.195 3.885 ;
      LAYER via1 ;
        RECT 73.04 4.995 73.19 5.145 ;
      LAYER via2 ;
        RECT 73.015 4.97 73.215 5.17 ;
      LAYER mcon ;
        RECT 73.025 3.685 73.195 3.855 ;
        RECT 73.025 2.205 73.195 2.375 ;
        RECT 73.03 4.985 73.2 5.155 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 88.185 0 88.565 5.26 ;
      LAYER met2 ;
        RECT 88.185 4.88 88.565 5.26 ;
      LAYER li1 ;
        RECT 88.285 1.865 88.46 2.375 ;
        RECT 88.285 3.895 88.46 5.155 ;
        RECT 88.285 3.685 88.455 5.155 ;
      LAYER met1 ;
        RECT 88.2 4.925 88.55 5.215 ;
        RECT 88.225 2.175 88.52 2.405 ;
        RECT 88.225 3.655 88.515 3.885 ;
        RECT 88.285 2.175 88.455 3.885 ;
      LAYER via1 ;
        RECT 88.3 4.995 88.45 5.145 ;
      LAYER via2 ;
        RECT 88.275 4.97 88.475 5.17 ;
      LAYER mcon ;
        RECT 88.285 3.685 88.455 3.855 ;
        RECT 88.285 2.205 88.455 2.375 ;
        RECT 88.29 4.985 88.46 5.155 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 103.445 0 103.825 5.26 ;
      LAYER met2 ;
        RECT 103.445 4.88 103.825 5.26 ;
      LAYER li1 ;
        RECT 103.545 1.865 103.72 2.375 ;
        RECT 103.545 3.895 103.72 5.155 ;
        RECT 103.545 3.685 103.715 5.155 ;
      LAYER met1 ;
        RECT 103.46 4.925 103.81 5.215 ;
        RECT 103.485 2.175 103.78 2.405 ;
        RECT 103.485 3.655 103.775 3.885 ;
        RECT 103.545 2.175 103.715 3.885 ;
      LAYER via1 ;
        RECT 103.56 4.995 103.71 5.145 ;
      LAYER via2 ;
        RECT 103.535 4.97 103.735 5.17 ;
      LAYER mcon ;
        RECT 103.545 3.685 103.715 3.855 ;
        RECT 103.545 2.205 103.715 2.375 ;
        RECT 103.55 4.985 103.72 5.155 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 38.28 8.15 38.62 8.5 ;
        RECT 38.28 4 38.62 4.35 ;
        RECT 38.36 4 38.53 8.5 ;
      LAYER li1 ;
        RECT 38.355 2.955 38.525 4.225 ;
        RECT 38.355 8.24 38.525 9.51 ;
        RECT 32.74 8.24 32.91 9.51 ;
      LAYER met1 ;
        RECT 38.28 4.055 38.755 4.225 ;
        RECT 38.28 4 38.62 4.35 ;
        RECT 38.28 8.24 38.755 8.41 ;
        RECT 38.28 8.15 38.62 8.5 ;
        RECT 32.68 8.235 38.62 8.405 ;
        RECT 32.68 8.235 33.14 8.41 ;
        RECT 32.68 8.21 32.97 8.44 ;
      LAYER via1 ;
        RECT 38.38 8.25 38.53 8.4 ;
        RECT 38.38 4.1 38.53 4.25 ;
      LAYER mcon ;
        RECT 32.74 8.24 32.91 8.41 ;
        RECT 38.355 8.24 38.525 8.41 ;
        RECT 38.355 4.055 38.525 4.225 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 53.54 8.15 53.88 8.5 ;
        RECT 53.54 4 53.88 4.35 ;
        RECT 53.62 4 53.79 8.5 ;
      LAYER li1 ;
        RECT 53.615 2.955 53.785 4.225 ;
        RECT 53.615 8.24 53.785 9.51 ;
        RECT 48 8.24 48.17 9.51 ;
      LAYER met1 ;
        RECT 53.54 4.055 54.015 4.225 ;
        RECT 53.54 4 53.88 4.35 ;
        RECT 53.54 8.24 54.015 8.41 ;
        RECT 53.54 8.15 53.88 8.5 ;
        RECT 47.94 8.235 53.88 8.405 ;
        RECT 47.94 8.235 48.4 8.41 ;
        RECT 47.94 8.21 48.23 8.44 ;
      LAYER via1 ;
        RECT 53.64 8.25 53.79 8.4 ;
        RECT 53.64 4.1 53.79 4.25 ;
      LAYER mcon ;
        RECT 48 8.24 48.17 8.41 ;
        RECT 53.615 8.24 53.785 8.41 ;
        RECT 53.615 4.055 53.785 4.225 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 68.8 8.15 69.14 8.5 ;
        RECT 68.8 4 69.14 4.35 ;
        RECT 68.88 4 69.05 8.5 ;
      LAYER li1 ;
        RECT 68.875 2.955 69.045 4.225 ;
        RECT 68.875 8.24 69.045 9.51 ;
        RECT 63.26 8.24 63.43 9.51 ;
      LAYER met1 ;
        RECT 68.8 4.055 69.275 4.225 ;
        RECT 68.8 4 69.14 4.35 ;
        RECT 68.8 8.24 69.275 8.41 ;
        RECT 68.8 8.15 69.14 8.5 ;
        RECT 63.2 8.235 69.14 8.405 ;
        RECT 63.2 8.235 63.66 8.41 ;
        RECT 63.2 8.21 63.49 8.44 ;
      LAYER via1 ;
        RECT 68.9 8.25 69.05 8.4 ;
        RECT 68.9 4.1 69.05 4.25 ;
      LAYER mcon ;
        RECT 63.26 8.24 63.43 8.41 ;
        RECT 68.875 8.24 69.045 8.41 ;
        RECT 68.875 4.055 69.045 4.225 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 84.06 8.15 84.4 8.5 ;
        RECT 84.06 4 84.4 4.35 ;
        RECT 84.14 4 84.31 8.5 ;
      LAYER li1 ;
        RECT 84.135 2.955 84.305 4.225 ;
        RECT 84.135 8.24 84.305 9.51 ;
        RECT 78.52 8.24 78.69 9.51 ;
      LAYER met1 ;
        RECT 84.06 4.055 84.535 4.225 ;
        RECT 84.06 4 84.4 4.35 ;
        RECT 84.06 8.24 84.535 8.41 ;
        RECT 84.06 8.15 84.4 8.5 ;
        RECT 78.46 8.235 84.4 8.405 ;
        RECT 78.46 8.235 78.92 8.41 ;
        RECT 78.46 8.21 78.75 8.44 ;
      LAYER via1 ;
        RECT 84.16 8.25 84.31 8.4 ;
        RECT 84.16 4.1 84.31 4.25 ;
      LAYER mcon ;
        RECT 78.52 8.24 78.69 8.41 ;
        RECT 84.135 8.24 84.305 8.41 ;
        RECT 84.135 4.055 84.305 4.225 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 99.32 8.15 99.66 8.5 ;
        RECT 99.32 4 99.66 4.35 ;
        RECT 99.4 4 99.57 8.5 ;
      LAYER li1 ;
        RECT 99.395 2.955 99.565 4.225 ;
        RECT 99.395 8.24 99.565 9.51 ;
        RECT 93.78 8.24 93.95 9.51 ;
      LAYER met1 ;
        RECT 99.32 4.055 99.795 4.225 ;
        RECT 99.32 4 99.66 4.35 ;
        RECT 99.32 8.24 99.795 8.41 ;
        RECT 99.32 8.15 99.66 8.5 ;
        RECT 93.72 8.235 99.66 8.405 ;
        RECT 93.72 8.235 94.18 8.41 ;
        RECT 93.72 8.21 94.01 8.44 ;
      LAYER via1 ;
        RECT 99.42 8.25 99.57 8.4 ;
        RECT 99.42 4.1 99.57 4.25 ;
      LAYER mcon ;
        RECT 93.78 8.24 93.95 8.41 ;
        RECT 99.395 8.24 99.565 8.41 ;
        RECT 99.395 4.055 99.565 4.225 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 25.225 8.24 25.395 9.51 ;
      LAYER met1 ;
        RECT 25.165 8.24 25.625 8.41 ;
        RECT 25.17 8.205 25.46 8.435 ;
        RECT 25.165 8.21 25.455 8.44 ;
      LAYER mcon ;
        RECT 25.225 8.24 25.395 8.41 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 5.435 104.095 7.035 ;
        RECT 89.585 5.43 104.095 7.035 ;
        RECT 99.215 5.43 103.94 7.04 ;
        RECT 99.215 5.425 103.935 7.04 ;
        RECT 103.12 5.425 103.29 7.77 ;
        RECT 103.115 4.695 103.285 7.04 ;
        RECT 102.13 4.695 102.3 7.77 ;
        RECT 99.385 4.695 99.555 7.77 ;
        RECT 96.615 4.93 96.785 7.035 ;
        RECT 93.6 5.43 96.35 7.04 ;
        RECT 94.695 4.93 94.865 7.04 ;
        RECT 93.77 5.43 93.94 7.77 ;
        RECT 93.755 4.93 93.925 7.04 ;
        RECT 92.295 4.93 92.465 7.035 ;
        RECT 90.375 4.93 90.545 7.035 ;
        RECT 74.325 5.43 88.835 7.035 ;
        RECT 83.955 5.43 88.68 7.04 ;
        RECT 83.955 5.425 88.675 7.04 ;
        RECT 87.86 5.425 88.03 7.77 ;
        RECT 87.855 4.695 88.025 7.04 ;
        RECT 86.87 4.695 87.04 7.77 ;
        RECT 84.125 4.695 84.295 7.77 ;
        RECT 81.355 4.93 81.525 7.035 ;
        RECT 78.34 5.43 81.09 7.04 ;
        RECT 79.435 4.93 79.605 7.04 ;
        RECT 78.51 5.43 78.68 7.77 ;
        RECT 78.495 4.93 78.665 7.04 ;
        RECT 77.035 4.93 77.205 7.035 ;
        RECT 75.115 4.93 75.285 7.035 ;
        RECT 59.065 5.43 73.575 7.035 ;
        RECT 68.695 5.43 73.42 7.04 ;
        RECT 68.695 5.425 73.415 7.04 ;
        RECT 72.6 5.425 72.77 7.77 ;
        RECT 72.595 4.695 72.765 7.04 ;
        RECT 71.61 4.695 71.78 7.77 ;
        RECT 68.865 4.695 69.035 7.77 ;
        RECT 66.095 4.93 66.265 7.035 ;
        RECT 63.08 5.43 65.83 7.04 ;
        RECT 64.175 4.93 64.345 7.04 ;
        RECT 63.25 5.43 63.42 7.77 ;
        RECT 63.235 4.93 63.405 7.04 ;
        RECT 61.775 4.93 61.945 7.035 ;
        RECT 59.855 4.93 60.025 7.035 ;
        RECT 43.805 5.43 58.315 7.035 ;
        RECT 53.435 5.43 58.16 7.04 ;
        RECT 53.435 5.425 58.155 7.04 ;
        RECT 57.34 5.425 57.51 7.77 ;
        RECT 57.335 4.695 57.505 7.04 ;
        RECT 56.35 4.695 56.52 7.77 ;
        RECT 53.605 4.695 53.775 7.77 ;
        RECT 50.835 4.93 51.005 7.035 ;
        RECT 47.82 5.43 50.57 7.04 ;
        RECT 48.915 4.93 49.085 7.04 ;
        RECT 47.99 5.43 48.16 7.77 ;
        RECT 47.975 4.93 48.145 7.04 ;
        RECT 46.515 4.93 46.685 7.035 ;
        RECT 44.595 4.93 44.765 7.035 ;
        RECT 28.545 5.43 43.055 7.035 ;
        RECT 38.175 5.43 42.9 7.04 ;
        RECT 38.175 5.425 42.895 7.04 ;
        RECT 42.08 5.425 42.25 7.77 ;
        RECT 42.075 4.695 42.245 7.04 ;
        RECT 41.09 4.695 41.26 7.77 ;
        RECT 38.345 4.695 38.515 7.77 ;
        RECT 35.575 4.93 35.745 7.035 ;
        RECT 32.56 5.43 35.31 7.04 ;
        RECT 33.655 4.93 33.825 7.04 ;
        RECT 32.73 5.43 32.9 7.77 ;
        RECT 32.715 4.93 32.885 7.04 ;
        RECT 31.255 4.93 31.425 7.035 ;
        RECT 29.335 4.93 29.505 7.035 ;
        RECT 25.045 5.435 27.795 7.04 ;
        RECT 27.03 10.05 27.205 10.6 ;
        RECT 27.03 7.31 27.205 8.45 ;
        RECT 27.03 5.435 27.2 10.6 ;
        RECT 25.215 5.435 25.385 7.77 ;
      LAYER met1 ;
        RECT 0 5.435 104.095 7.035 ;
        RECT 89.585 5.43 104.095 7.035 ;
        RECT 99.215 5.43 103.94 7.04 ;
        RECT 99.215 5.425 103.935 7.04 ;
        RECT 89.585 5.4 98.325 7.035 ;
        RECT 93.6 5.4 96.35 7.04 ;
        RECT 74.325 5.43 88.835 7.035 ;
        RECT 83.955 5.43 88.68 7.04 ;
        RECT 83.955 5.425 88.675 7.04 ;
        RECT 74.325 5.4 83.065 7.035 ;
        RECT 78.34 5.4 81.09 7.04 ;
        RECT 59.065 5.43 73.575 7.035 ;
        RECT 68.695 5.43 73.42 7.04 ;
        RECT 68.695 5.425 73.415 7.04 ;
        RECT 59.065 5.4 67.805 7.035 ;
        RECT 63.08 5.4 65.83 7.04 ;
        RECT 43.805 5.43 58.315 7.035 ;
        RECT 53.435 5.43 58.16 7.04 ;
        RECT 53.435 5.425 58.155 7.04 ;
        RECT 43.805 5.4 52.545 7.035 ;
        RECT 47.82 5.4 50.57 7.04 ;
        RECT 28.545 5.43 43.055 7.035 ;
        RECT 38.175 5.43 42.9 7.04 ;
        RECT 38.175 5.425 42.895 7.04 ;
        RECT 28.545 5.4 37.285 7.035 ;
        RECT 32.56 5.4 35.31 7.04 ;
        RECT 25.045 5.435 27.795 7.04 ;
        RECT 26.97 8.95 27.26 9.18 ;
        RECT 26.8 8.98 27.26 9.15 ;
      LAYER mcon ;
        RECT 27.03 8.98 27.2 9.15 ;
        RECT 27.335 6.84 27.505 7.01 ;
        RECT 28.69 5.43 28.86 5.6 ;
        RECT 29.15 5.43 29.32 5.6 ;
        RECT 29.61 5.43 29.78 5.6 ;
        RECT 30.07 5.43 30.24 5.6 ;
        RECT 30.53 5.43 30.7 5.6 ;
        RECT 30.99 5.43 31.16 5.6 ;
        RECT 31.45 5.43 31.62 5.6 ;
        RECT 31.91 5.43 32.08 5.6 ;
        RECT 32.37 5.43 32.54 5.6 ;
        RECT 32.83 5.43 33 5.6 ;
        RECT 33.29 5.43 33.46 5.6 ;
        RECT 33.75 5.43 33.92 5.6 ;
        RECT 34.21 5.43 34.38 5.6 ;
        RECT 34.67 5.43 34.84 5.6 ;
        RECT 34.85 6.84 35.02 7.01 ;
        RECT 35.13 5.43 35.3 5.6 ;
        RECT 35.59 5.43 35.76 5.6 ;
        RECT 36.05 5.43 36.22 5.6 ;
        RECT 36.51 5.43 36.68 5.6 ;
        RECT 36.97 5.43 37.14 5.6 ;
        RECT 40.465 6.84 40.635 7.01 ;
        RECT 40.465 5.455 40.635 5.625 ;
        RECT 41.17 6.84 41.34 7.01 ;
        RECT 41.17 5.455 41.34 5.625 ;
        RECT 42.155 5.455 42.325 5.625 ;
        RECT 42.16 6.84 42.33 7.01 ;
        RECT 43.95 5.43 44.12 5.6 ;
        RECT 44.41 5.43 44.58 5.6 ;
        RECT 44.87 5.43 45.04 5.6 ;
        RECT 45.33 5.43 45.5 5.6 ;
        RECT 45.79 5.43 45.96 5.6 ;
        RECT 46.25 5.43 46.42 5.6 ;
        RECT 46.71 5.43 46.88 5.6 ;
        RECT 47.17 5.43 47.34 5.6 ;
        RECT 47.63 5.43 47.8 5.6 ;
        RECT 48.09 5.43 48.26 5.6 ;
        RECT 48.55 5.43 48.72 5.6 ;
        RECT 49.01 5.43 49.18 5.6 ;
        RECT 49.47 5.43 49.64 5.6 ;
        RECT 49.93 5.43 50.1 5.6 ;
        RECT 50.11 6.84 50.28 7.01 ;
        RECT 50.39 5.43 50.56 5.6 ;
        RECT 50.85 5.43 51.02 5.6 ;
        RECT 51.31 5.43 51.48 5.6 ;
        RECT 51.77 5.43 51.94 5.6 ;
        RECT 52.23 5.43 52.4 5.6 ;
        RECT 55.725 6.84 55.895 7.01 ;
        RECT 55.725 5.455 55.895 5.625 ;
        RECT 56.43 6.84 56.6 7.01 ;
        RECT 56.43 5.455 56.6 5.625 ;
        RECT 57.415 5.455 57.585 5.625 ;
        RECT 57.42 6.84 57.59 7.01 ;
        RECT 59.21 5.43 59.38 5.6 ;
        RECT 59.67 5.43 59.84 5.6 ;
        RECT 60.13 5.43 60.3 5.6 ;
        RECT 60.59 5.43 60.76 5.6 ;
        RECT 61.05 5.43 61.22 5.6 ;
        RECT 61.51 5.43 61.68 5.6 ;
        RECT 61.97 5.43 62.14 5.6 ;
        RECT 62.43 5.43 62.6 5.6 ;
        RECT 62.89 5.43 63.06 5.6 ;
        RECT 63.35 5.43 63.52 5.6 ;
        RECT 63.81 5.43 63.98 5.6 ;
        RECT 64.27 5.43 64.44 5.6 ;
        RECT 64.73 5.43 64.9 5.6 ;
        RECT 65.19 5.43 65.36 5.6 ;
        RECT 65.37 6.84 65.54 7.01 ;
        RECT 65.65 5.43 65.82 5.6 ;
        RECT 66.11 5.43 66.28 5.6 ;
        RECT 66.57 5.43 66.74 5.6 ;
        RECT 67.03 5.43 67.2 5.6 ;
        RECT 67.49 5.43 67.66 5.6 ;
        RECT 70.985 6.84 71.155 7.01 ;
        RECT 70.985 5.455 71.155 5.625 ;
        RECT 71.69 6.84 71.86 7.01 ;
        RECT 71.69 5.455 71.86 5.625 ;
        RECT 72.675 5.455 72.845 5.625 ;
        RECT 72.68 6.84 72.85 7.01 ;
        RECT 74.47 5.43 74.64 5.6 ;
        RECT 74.93 5.43 75.1 5.6 ;
        RECT 75.39 5.43 75.56 5.6 ;
        RECT 75.85 5.43 76.02 5.6 ;
        RECT 76.31 5.43 76.48 5.6 ;
        RECT 76.77 5.43 76.94 5.6 ;
        RECT 77.23 5.43 77.4 5.6 ;
        RECT 77.69 5.43 77.86 5.6 ;
        RECT 78.15 5.43 78.32 5.6 ;
        RECT 78.61 5.43 78.78 5.6 ;
        RECT 79.07 5.43 79.24 5.6 ;
        RECT 79.53 5.43 79.7 5.6 ;
        RECT 79.99 5.43 80.16 5.6 ;
        RECT 80.45 5.43 80.62 5.6 ;
        RECT 80.63 6.84 80.8 7.01 ;
        RECT 80.91 5.43 81.08 5.6 ;
        RECT 81.37 5.43 81.54 5.6 ;
        RECT 81.83 5.43 82 5.6 ;
        RECT 82.29 5.43 82.46 5.6 ;
        RECT 82.75 5.43 82.92 5.6 ;
        RECT 86.245 6.84 86.415 7.01 ;
        RECT 86.245 5.455 86.415 5.625 ;
        RECT 86.95 6.84 87.12 7.01 ;
        RECT 86.95 5.455 87.12 5.625 ;
        RECT 87.935 5.455 88.105 5.625 ;
        RECT 87.94 6.84 88.11 7.01 ;
        RECT 89.73 5.43 89.9 5.6 ;
        RECT 90.19 5.43 90.36 5.6 ;
        RECT 90.65 5.43 90.82 5.6 ;
        RECT 91.11 5.43 91.28 5.6 ;
        RECT 91.57 5.43 91.74 5.6 ;
        RECT 92.03 5.43 92.2 5.6 ;
        RECT 92.49 5.43 92.66 5.6 ;
        RECT 92.95 5.43 93.12 5.6 ;
        RECT 93.41 5.43 93.58 5.6 ;
        RECT 93.87 5.43 94.04 5.6 ;
        RECT 94.33 5.43 94.5 5.6 ;
        RECT 94.79 5.43 94.96 5.6 ;
        RECT 95.25 5.43 95.42 5.6 ;
        RECT 95.71 5.43 95.88 5.6 ;
        RECT 95.89 6.84 96.06 7.01 ;
        RECT 96.17 5.43 96.34 5.6 ;
        RECT 96.63 5.43 96.8 5.6 ;
        RECT 97.09 5.43 97.26 5.6 ;
        RECT 97.55 5.43 97.72 5.6 ;
        RECT 98.01 5.43 98.18 5.6 ;
        RECT 101.505 6.84 101.675 7.01 ;
        RECT 101.505 5.455 101.675 5.625 ;
        RECT 102.21 6.84 102.38 7.01 ;
        RECT 102.21 5.455 102.38 5.625 ;
        RECT 103.195 5.455 103.365 5.625 ;
        RECT 103.2 6.84 103.37 7.01 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 90.415 3.15 91.145 3.48 ;
        RECT 75.155 3.15 75.885 3.48 ;
        RECT 59.895 3.15 60.625 3.48 ;
        RECT 44.635 3.15 45.365 3.48 ;
        RECT 29.375 3.15 30.105 3.48 ;
      LAYER met2 ;
        RECT 90.56 3.155 90.95 3.475 ;
        RECT 90.56 3.13 90.84 3.5 ;
        RECT 75.3 3.155 75.69 3.475 ;
        RECT 75.3 3.13 75.58 3.5 ;
        RECT 60.04 3.155 60.43 3.475 ;
        RECT 60.04 3.13 60.32 3.5 ;
        RECT 44.78 3.155 45.17 3.475 ;
        RECT 44.78 3.13 45.06 3.5 ;
        RECT 29.52 3.155 29.91 3.475 ;
        RECT 29.52 3.13 29.8 3.5 ;
      LAYER li1 ;
        RECT 0 0 104.095 1.6 ;
        RECT 103.115 0 103.285 2.225 ;
        RECT 102.13 0 102.3 2.225 ;
        RECT 99.385 0 99.555 2.225 ;
        RECT 89.585 0 98.325 2.88 ;
        RECT 97.555 0 97.725 3.38 ;
        RECT 96.615 0 96.785 3.38 ;
        RECT 95.655 0 95.825 3.38 ;
        RECT 94.61 0 94.805 2.89 ;
        RECT 93.735 0 93.905 3.38 ;
        RECT 92.775 0 92.945 3.38 ;
        RECT 90.855 0 91.13 2.89 ;
        RECT 90.855 0 91.025 3.38 ;
        RECT 87.855 0 88.025 2.225 ;
        RECT 86.87 0 87.04 2.225 ;
        RECT 84.125 0 84.295 2.225 ;
        RECT 74.325 0 83.065 2.88 ;
        RECT 82.295 0 82.465 3.38 ;
        RECT 81.355 0 81.525 3.38 ;
        RECT 80.395 0 80.565 3.38 ;
        RECT 79.35 0 79.545 2.89 ;
        RECT 78.475 0 78.645 3.38 ;
        RECT 77.515 0 77.685 3.38 ;
        RECT 75.595 0 75.87 2.89 ;
        RECT 75.595 0 75.765 3.38 ;
        RECT 72.595 0 72.765 2.225 ;
        RECT 71.61 0 71.78 2.225 ;
        RECT 68.865 0 69.035 2.225 ;
        RECT 59.065 0 67.805 2.88 ;
        RECT 67.035 0 67.205 3.38 ;
        RECT 66.095 0 66.265 3.38 ;
        RECT 65.135 0 65.305 3.38 ;
        RECT 64.09 0 64.285 2.89 ;
        RECT 63.215 0 63.385 3.38 ;
        RECT 62.255 0 62.425 3.38 ;
        RECT 60.335 0 60.61 2.89 ;
        RECT 60.335 0 60.505 3.38 ;
        RECT 57.335 0 57.505 2.225 ;
        RECT 56.35 0 56.52 2.225 ;
        RECT 53.605 0 53.775 2.225 ;
        RECT 43.805 0 52.545 2.88 ;
        RECT 51.775 0 51.945 3.38 ;
        RECT 50.835 0 51.005 3.38 ;
        RECT 49.875 0 50.045 3.38 ;
        RECT 48.83 0 49.025 2.89 ;
        RECT 47.955 0 48.125 3.38 ;
        RECT 46.995 0 47.165 3.38 ;
        RECT 45.075 0 45.35 2.89 ;
        RECT 45.075 0 45.245 3.38 ;
        RECT 42.075 0 42.245 2.225 ;
        RECT 41.09 0 41.26 2.225 ;
        RECT 38.345 0 38.515 2.225 ;
        RECT 28.545 0 37.285 2.88 ;
        RECT 36.515 0 36.685 3.38 ;
        RECT 35.575 0 35.745 3.38 ;
        RECT 34.615 0 34.785 3.38 ;
        RECT 33.57 0 33.765 2.89 ;
        RECT 32.695 0 32.865 3.38 ;
        RECT 31.735 0 31.905 3.38 ;
        RECT 29.815 0 30.09 2.89 ;
        RECT 29.815 0 29.985 3.38 ;
        RECT 0 10.865 104.095 12.465 ;
        RECT 103.12 10.24 103.29 12.465 ;
        RECT 102.13 10.24 102.3 12.465 ;
        RECT 99.385 10.24 99.555 12.465 ;
        RECT 93.77 10.24 93.94 12.465 ;
        RECT 87.86 10.24 88.03 12.465 ;
        RECT 86.87 10.24 87.04 12.465 ;
        RECT 84.125 10.24 84.295 12.465 ;
        RECT 78.51 10.24 78.68 12.465 ;
        RECT 72.6 10.24 72.77 12.465 ;
        RECT 71.61 10.24 71.78 12.465 ;
        RECT 68.865 10.24 69.035 12.465 ;
        RECT 63.25 10.24 63.42 12.465 ;
        RECT 57.34 10.24 57.51 12.465 ;
        RECT 56.35 10.24 56.52 12.465 ;
        RECT 53.605 10.24 53.775 12.465 ;
        RECT 47.99 10.24 48.16 12.465 ;
        RECT 42.08 10.24 42.25 12.465 ;
        RECT 41.09 10.24 41.26 12.465 ;
        RECT 38.345 10.24 38.515 12.465 ;
        RECT 32.73 10.24 32.9 12.465 ;
        RECT 25.215 10.24 25.385 12.465 ;
        RECT 94.785 8.37 94.955 10.32 ;
        RECT 94.725 10.15 94.895 10.6 ;
        RECT 94.725 7.31 94.895 8.54 ;
        RECT 91.455 3.87 91.825 4.04 ;
        RECT 91.455 3.23 91.625 4.04 ;
        RECT 91.335 3.23 91.625 3.4 ;
        RECT 90.135 3.79 90.305 4.24 ;
        RECT 79.525 8.37 79.695 10.32 ;
        RECT 79.465 10.15 79.635 10.6 ;
        RECT 79.465 7.31 79.635 8.54 ;
        RECT 76.195 3.87 76.565 4.04 ;
        RECT 76.195 3.23 76.365 4.04 ;
        RECT 76.075 3.23 76.365 3.4 ;
        RECT 74.875 3.79 75.045 4.24 ;
        RECT 64.265 8.37 64.435 10.32 ;
        RECT 64.205 10.15 64.375 10.6 ;
        RECT 64.205 7.31 64.375 8.54 ;
        RECT 60.935 3.87 61.305 4.04 ;
        RECT 60.935 3.23 61.105 4.04 ;
        RECT 60.815 3.23 61.105 3.4 ;
        RECT 59.615 3.79 59.785 4.24 ;
        RECT 49.005 8.37 49.175 10.32 ;
        RECT 48.945 10.15 49.115 10.6 ;
        RECT 48.945 7.31 49.115 8.54 ;
        RECT 45.675 3.87 46.045 4.04 ;
        RECT 45.675 3.23 45.845 4.04 ;
        RECT 45.555 3.23 45.845 3.4 ;
        RECT 44.355 3.79 44.525 4.24 ;
        RECT 33.745 8.37 33.915 10.32 ;
        RECT 33.685 10.15 33.855 10.6 ;
        RECT 33.685 7.31 33.855 8.54 ;
        RECT 30.415 3.87 30.785 4.04 ;
        RECT 30.415 3.23 30.585 4.04 ;
        RECT 30.295 3.23 30.585 3.4 ;
        RECT 29.095 3.79 29.265 4.24 ;
      LAYER met1 ;
        RECT 0 0 104.095 1.6 ;
        RECT 89.585 0 98.325 2.915 ;
        RECT 91.275 3.2 91.565 3.43 ;
        RECT 90.39 3.245 91.565 3.385 ;
        RECT 90.57 3.185 90.98 3.445 ;
        RECT 90.57 0 90.86 3.445 ;
        RECT 90.15 3.665 90.77 3.805 ;
        RECT 90.63 0 90.77 3.805 ;
        RECT 90.39 3.245 90.77 3.505 ;
        RECT 90.075 4.04 90.365 4.27 ;
        RECT 90.15 3.665 90.29 4.27 ;
        RECT 74.325 0 83.065 2.915 ;
        RECT 76.015 3.2 76.305 3.43 ;
        RECT 75.13 3.245 76.305 3.385 ;
        RECT 75.31 3.185 75.72 3.445 ;
        RECT 75.31 0 75.6 3.445 ;
        RECT 74.89 3.665 75.51 3.805 ;
        RECT 75.37 0 75.51 3.805 ;
        RECT 75.13 3.245 75.51 3.505 ;
        RECT 74.815 4.04 75.105 4.27 ;
        RECT 74.89 3.665 75.03 4.27 ;
        RECT 59.065 0 67.805 2.915 ;
        RECT 60.755 3.2 61.045 3.43 ;
        RECT 59.87 3.245 61.045 3.385 ;
        RECT 60.05 3.185 60.46 3.445 ;
        RECT 60.05 0 60.34 3.445 ;
        RECT 59.63 3.665 60.25 3.805 ;
        RECT 60.11 0 60.25 3.805 ;
        RECT 59.87 3.245 60.25 3.505 ;
        RECT 59.555 4.04 59.845 4.27 ;
        RECT 59.63 3.665 59.77 4.27 ;
        RECT 43.805 0 52.545 2.915 ;
        RECT 45.495 3.2 45.785 3.43 ;
        RECT 44.61 3.245 45.785 3.385 ;
        RECT 44.79 3.185 45.2 3.445 ;
        RECT 44.79 0 45.08 3.445 ;
        RECT 44.37 3.665 44.99 3.805 ;
        RECT 44.85 0 44.99 3.805 ;
        RECT 44.61 3.245 44.99 3.505 ;
        RECT 44.295 4.04 44.585 4.27 ;
        RECT 44.37 3.665 44.51 4.27 ;
        RECT 28.545 0 37.285 2.915 ;
        RECT 30.235 3.2 30.525 3.43 ;
        RECT 29.35 3.245 30.525 3.385 ;
        RECT 29.53 3.185 29.94 3.445 ;
        RECT 29.53 0 29.82 3.445 ;
        RECT 29.11 3.665 29.73 3.805 ;
        RECT 29.59 0 29.73 3.805 ;
        RECT 29.35 3.245 29.73 3.505 ;
        RECT 29.035 4.04 29.325 4.27 ;
        RECT 29.11 3.665 29.25 4.27 ;
        RECT 0 10.865 104.095 12.465 ;
        RECT 94.725 8.58 95.015 8.81 ;
        RECT 94.555 8.605 94.725 12.465 ;
        RECT 94.55 8.61 95.015 8.78 ;
        RECT 79.465 8.58 79.755 8.81 ;
        RECT 79.295 8.605 79.465 12.465 ;
        RECT 79.29 8.61 79.755 8.78 ;
        RECT 64.205 8.58 64.495 8.81 ;
        RECT 64.035 8.605 64.205 12.465 ;
        RECT 64.03 8.61 64.495 8.78 ;
        RECT 48.945 8.58 49.235 8.81 ;
        RECT 48.775 8.605 48.945 12.465 ;
        RECT 48.77 8.61 49.235 8.78 ;
        RECT 33.685 8.58 33.975 8.81 ;
        RECT 33.515 8.605 33.685 12.465 ;
        RECT 33.51 8.61 33.975 8.78 ;
      LAYER via1 ;
        RECT 29.705 3.24 29.855 3.39 ;
        RECT 44.965 3.24 45.115 3.39 ;
        RECT 60.225 3.24 60.375 3.39 ;
        RECT 75.485 3.24 75.635 3.39 ;
        RECT 90.745 3.24 90.895 3.39 ;
      LAYER via2 ;
        RECT 29.56 3.215 29.76 3.415 ;
        RECT 44.82 3.215 45.02 3.415 ;
        RECT 60.08 3.215 60.28 3.415 ;
        RECT 75.34 3.215 75.54 3.415 ;
        RECT 90.6 3.215 90.8 3.415 ;
      LAYER mcon ;
        RECT 25.295 10.9 25.465 11.07 ;
        RECT 25.975 10.9 26.145 11.07 ;
        RECT 26.655 10.9 26.825 11.07 ;
        RECT 27.335 10.9 27.505 11.07 ;
        RECT 28.69 2.71 28.86 2.88 ;
        RECT 29.095 4.07 29.265 4.24 ;
        RECT 29.15 2.71 29.32 2.88 ;
        RECT 29.61 2.71 29.78 2.88 ;
        RECT 30.07 2.71 30.24 2.88 ;
        RECT 30.295 3.23 30.465 3.4 ;
        RECT 30.53 2.71 30.7 2.88 ;
        RECT 30.99 2.71 31.16 2.88 ;
        RECT 31.45 2.71 31.62 2.88 ;
        RECT 31.91 2.71 32.08 2.88 ;
        RECT 32.37 2.71 32.54 2.88 ;
        RECT 32.81 10.9 32.98 11.07 ;
        RECT 32.83 2.71 33 2.88 ;
        RECT 33.29 2.71 33.46 2.88 ;
        RECT 33.49 10.9 33.66 11.07 ;
        RECT 33.745 8.61 33.915 8.78 ;
        RECT 33.75 2.71 33.92 2.88 ;
        RECT 34.17 10.9 34.34 11.07 ;
        RECT 34.21 2.71 34.38 2.88 ;
        RECT 34.67 2.71 34.84 2.88 ;
        RECT 34.85 10.9 35.02 11.07 ;
        RECT 35.13 2.71 35.3 2.88 ;
        RECT 35.59 2.71 35.76 2.88 ;
        RECT 36.05 2.71 36.22 2.88 ;
        RECT 36.51 2.71 36.68 2.88 ;
        RECT 36.97 2.71 37.14 2.88 ;
        RECT 38.425 10.9 38.595 11.07 ;
        RECT 38.425 1.395 38.595 1.565 ;
        RECT 39.105 10.9 39.275 11.07 ;
        RECT 39.105 1.395 39.275 1.565 ;
        RECT 39.785 10.9 39.955 11.07 ;
        RECT 39.785 1.395 39.955 1.565 ;
        RECT 40.465 10.9 40.635 11.07 ;
        RECT 40.465 1.395 40.635 1.565 ;
        RECT 41.17 10.9 41.34 11.07 ;
        RECT 41.17 1.395 41.34 1.565 ;
        RECT 42.155 1.395 42.325 1.565 ;
        RECT 42.16 10.9 42.33 11.07 ;
        RECT 43.95 2.71 44.12 2.88 ;
        RECT 44.355 4.07 44.525 4.24 ;
        RECT 44.41 2.71 44.58 2.88 ;
        RECT 44.87 2.71 45.04 2.88 ;
        RECT 45.33 2.71 45.5 2.88 ;
        RECT 45.555 3.23 45.725 3.4 ;
        RECT 45.79 2.71 45.96 2.88 ;
        RECT 46.25 2.71 46.42 2.88 ;
        RECT 46.71 2.71 46.88 2.88 ;
        RECT 47.17 2.71 47.34 2.88 ;
        RECT 47.63 2.71 47.8 2.88 ;
        RECT 48.07 10.9 48.24 11.07 ;
        RECT 48.09 2.71 48.26 2.88 ;
        RECT 48.55 2.71 48.72 2.88 ;
        RECT 48.75 10.9 48.92 11.07 ;
        RECT 49.005 8.61 49.175 8.78 ;
        RECT 49.01 2.71 49.18 2.88 ;
        RECT 49.43 10.9 49.6 11.07 ;
        RECT 49.47 2.71 49.64 2.88 ;
        RECT 49.93 2.71 50.1 2.88 ;
        RECT 50.11 10.9 50.28 11.07 ;
        RECT 50.39 2.71 50.56 2.88 ;
        RECT 50.85 2.71 51.02 2.88 ;
        RECT 51.31 2.71 51.48 2.88 ;
        RECT 51.77 2.71 51.94 2.88 ;
        RECT 52.23 2.71 52.4 2.88 ;
        RECT 53.685 10.9 53.855 11.07 ;
        RECT 53.685 1.395 53.855 1.565 ;
        RECT 54.365 10.9 54.535 11.07 ;
        RECT 54.365 1.395 54.535 1.565 ;
        RECT 55.045 10.9 55.215 11.07 ;
        RECT 55.045 1.395 55.215 1.565 ;
        RECT 55.725 10.9 55.895 11.07 ;
        RECT 55.725 1.395 55.895 1.565 ;
        RECT 56.43 10.9 56.6 11.07 ;
        RECT 56.43 1.395 56.6 1.565 ;
        RECT 57.415 1.395 57.585 1.565 ;
        RECT 57.42 10.9 57.59 11.07 ;
        RECT 59.21 2.71 59.38 2.88 ;
        RECT 59.615 4.07 59.785 4.24 ;
        RECT 59.67 2.71 59.84 2.88 ;
        RECT 60.13 2.71 60.3 2.88 ;
        RECT 60.59 2.71 60.76 2.88 ;
        RECT 60.815 3.23 60.985 3.4 ;
        RECT 61.05 2.71 61.22 2.88 ;
        RECT 61.51 2.71 61.68 2.88 ;
        RECT 61.97 2.71 62.14 2.88 ;
        RECT 62.43 2.71 62.6 2.88 ;
        RECT 62.89 2.71 63.06 2.88 ;
        RECT 63.33 10.9 63.5 11.07 ;
        RECT 63.35 2.71 63.52 2.88 ;
        RECT 63.81 2.71 63.98 2.88 ;
        RECT 64.01 10.9 64.18 11.07 ;
        RECT 64.265 8.61 64.435 8.78 ;
        RECT 64.27 2.71 64.44 2.88 ;
        RECT 64.69 10.9 64.86 11.07 ;
        RECT 64.73 2.71 64.9 2.88 ;
        RECT 65.19 2.71 65.36 2.88 ;
        RECT 65.37 10.9 65.54 11.07 ;
        RECT 65.65 2.71 65.82 2.88 ;
        RECT 66.11 2.71 66.28 2.88 ;
        RECT 66.57 2.71 66.74 2.88 ;
        RECT 67.03 2.71 67.2 2.88 ;
        RECT 67.49 2.71 67.66 2.88 ;
        RECT 68.945 10.9 69.115 11.07 ;
        RECT 68.945 1.395 69.115 1.565 ;
        RECT 69.625 10.9 69.795 11.07 ;
        RECT 69.625 1.395 69.795 1.565 ;
        RECT 70.305 10.9 70.475 11.07 ;
        RECT 70.305 1.395 70.475 1.565 ;
        RECT 70.985 10.9 71.155 11.07 ;
        RECT 70.985 1.395 71.155 1.565 ;
        RECT 71.69 10.9 71.86 11.07 ;
        RECT 71.69 1.395 71.86 1.565 ;
        RECT 72.675 1.395 72.845 1.565 ;
        RECT 72.68 10.9 72.85 11.07 ;
        RECT 74.47 2.71 74.64 2.88 ;
        RECT 74.875 4.07 75.045 4.24 ;
        RECT 74.93 2.71 75.1 2.88 ;
        RECT 75.39 2.71 75.56 2.88 ;
        RECT 75.85 2.71 76.02 2.88 ;
        RECT 76.075 3.23 76.245 3.4 ;
        RECT 76.31 2.71 76.48 2.88 ;
        RECT 76.77 2.71 76.94 2.88 ;
        RECT 77.23 2.71 77.4 2.88 ;
        RECT 77.69 2.71 77.86 2.88 ;
        RECT 78.15 2.71 78.32 2.88 ;
        RECT 78.59 10.9 78.76 11.07 ;
        RECT 78.61 2.71 78.78 2.88 ;
        RECT 79.07 2.71 79.24 2.88 ;
        RECT 79.27 10.9 79.44 11.07 ;
        RECT 79.525 8.61 79.695 8.78 ;
        RECT 79.53 2.71 79.7 2.88 ;
        RECT 79.95 10.9 80.12 11.07 ;
        RECT 79.99 2.71 80.16 2.88 ;
        RECT 80.45 2.71 80.62 2.88 ;
        RECT 80.63 10.9 80.8 11.07 ;
        RECT 80.91 2.71 81.08 2.88 ;
        RECT 81.37 2.71 81.54 2.88 ;
        RECT 81.83 2.71 82 2.88 ;
        RECT 82.29 2.71 82.46 2.88 ;
        RECT 82.75 2.71 82.92 2.88 ;
        RECT 84.205 10.9 84.375 11.07 ;
        RECT 84.205 1.395 84.375 1.565 ;
        RECT 84.885 10.9 85.055 11.07 ;
        RECT 84.885 1.395 85.055 1.565 ;
        RECT 85.565 10.9 85.735 11.07 ;
        RECT 85.565 1.395 85.735 1.565 ;
        RECT 86.245 10.9 86.415 11.07 ;
        RECT 86.245 1.395 86.415 1.565 ;
        RECT 86.95 10.9 87.12 11.07 ;
        RECT 86.95 1.395 87.12 1.565 ;
        RECT 87.935 1.395 88.105 1.565 ;
        RECT 87.94 10.9 88.11 11.07 ;
        RECT 89.73 2.71 89.9 2.88 ;
        RECT 90.135 4.07 90.305 4.24 ;
        RECT 90.19 2.71 90.36 2.88 ;
        RECT 90.65 2.71 90.82 2.88 ;
        RECT 91.11 2.71 91.28 2.88 ;
        RECT 91.335 3.23 91.505 3.4 ;
        RECT 91.57 2.71 91.74 2.88 ;
        RECT 92.03 2.71 92.2 2.88 ;
        RECT 92.49 2.71 92.66 2.88 ;
        RECT 92.95 2.71 93.12 2.88 ;
        RECT 93.41 2.71 93.58 2.88 ;
        RECT 93.85 10.9 94.02 11.07 ;
        RECT 93.87 2.71 94.04 2.88 ;
        RECT 94.33 2.71 94.5 2.88 ;
        RECT 94.53 10.9 94.7 11.07 ;
        RECT 94.785 8.61 94.955 8.78 ;
        RECT 94.79 2.71 94.96 2.88 ;
        RECT 95.21 10.9 95.38 11.07 ;
        RECT 95.25 2.71 95.42 2.88 ;
        RECT 95.71 2.71 95.88 2.88 ;
        RECT 95.89 10.9 96.06 11.07 ;
        RECT 96.17 2.71 96.34 2.88 ;
        RECT 96.63 2.71 96.8 2.88 ;
        RECT 97.09 2.71 97.26 2.88 ;
        RECT 97.55 2.71 97.72 2.88 ;
        RECT 98.01 2.71 98.18 2.88 ;
        RECT 99.465 10.9 99.635 11.07 ;
        RECT 99.465 1.395 99.635 1.565 ;
        RECT 100.145 10.9 100.315 11.07 ;
        RECT 100.145 1.395 100.315 1.565 ;
        RECT 100.825 10.9 100.995 11.07 ;
        RECT 100.825 1.395 100.995 1.565 ;
        RECT 101.505 10.9 101.675 11.07 ;
        RECT 101.505 1.395 101.675 1.565 ;
        RECT 102.21 10.9 102.38 11.07 ;
        RECT 102.21 1.395 102.38 1.565 ;
        RECT 103.195 1.395 103.365 1.565 ;
        RECT 103.2 10.9 103.37 11.07 ;
    END
  END vssd1
  OBS
    LAYER met4 ;
      RECT 91.735 4.27 92.065 4.6 ;
      RECT 91.75 3.795 92.065 4.6 ;
      RECT 93.895 3.78 94.225 4.135 ;
      RECT 91.75 3.795 94.225 4.095 ;
      RECT 76.475 4.27 76.805 4.6 ;
      RECT 76.49 3.795 76.805 4.6 ;
      RECT 78.635 3.78 78.965 4.135 ;
      RECT 76.49 3.795 78.965 4.095 ;
      RECT 61.215 4.27 61.545 4.6 ;
      RECT 61.23 3.795 61.545 4.6 ;
      RECT 63.375 3.78 63.705 4.135 ;
      RECT 61.23 3.795 63.705 4.095 ;
      RECT 45.955 4.27 46.285 4.6 ;
      RECT 45.97 3.795 46.285 4.6 ;
      RECT 48.115 3.78 48.445 4.135 ;
      RECT 45.97 3.795 48.445 4.095 ;
      RECT 30.695 4.27 31.025 4.6 ;
      RECT 30.71 3.795 31.025 4.6 ;
      RECT 32.855 3.78 33.185 4.135 ;
      RECT 30.71 3.795 33.185 4.095 ;
    LAYER via3 ;
      RECT 93.96 3.87 94.16 4.07 ;
      RECT 91.8 4.335 92 4.535 ;
      RECT 78.7 3.87 78.9 4.07 ;
      RECT 76.54 4.335 76.74 4.535 ;
      RECT 63.44 3.87 63.64 4.07 ;
      RECT 61.28 4.335 61.48 4.535 ;
      RECT 48.18 3.87 48.38 4.07 ;
      RECT 46.02 4.335 46.22 4.535 ;
      RECT 32.92 3.87 33.12 4.07 ;
      RECT 30.76 4.335 30.96 4.535 ;
    LAYER met3 ;
      RECT 98.76 3.94 99.12 4.365 ;
      RECT 98.76 2.4 99.1 4.365 ;
      RECT 93.02 3.175 93.75 3.505 ;
      RECT 93.17 2.4 93.47 3.505 ;
      RECT 93.17 2.4 99.1 2.7 ;
      RECT 95.055 9.345 95.425 9.715 ;
      RECT 95.09 5.77 95.39 9.715 ;
      RECT 93.65 5.77 95.39 7.065 ;
      RECT 90.855 5.55 93.95 6.845 ;
      RECT 93.65 3.81 93.95 7.065 ;
      RECT 90.855 4.27 91.155 6.845 ;
      RECT 94.375 4.805 94.705 5.16 ;
      RECT 92.47 4.845 94.705 5.145 ;
      RECT 92.47 3.71 92.77 5.145 ;
      RECT 90.55 4.27 91.28 4.6 ;
      RECT 93.445 3.815 94.225 4.16 ;
      RECT 93.9 3.78 94.225 4.16 ;
      RECT 92.455 3.71 92.785 4.04 ;
      RECT 91.74 3.71 92.06 4.625 ;
      RECT 91.74 3.71 92.07 4.245 ;
      RECT 83.5 3.94 83.86 4.365 ;
      RECT 83.5 2.4 83.84 4.365 ;
      RECT 77.76 3.175 78.49 3.505 ;
      RECT 77.91 2.4 78.21 3.505 ;
      RECT 77.91 2.4 83.84 2.7 ;
      RECT 79.795 9.345 80.165 9.715 ;
      RECT 79.83 5.77 80.13 9.715 ;
      RECT 78.39 5.77 80.13 7.065 ;
      RECT 75.595 5.55 78.69 6.845 ;
      RECT 78.39 3.81 78.69 7.065 ;
      RECT 75.595 4.27 75.895 6.845 ;
      RECT 79.115 4.805 79.445 5.16 ;
      RECT 77.21 4.845 79.445 5.145 ;
      RECT 77.21 3.71 77.51 5.145 ;
      RECT 75.29 4.27 76.02 4.6 ;
      RECT 78.185 3.815 78.965 4.16 ;
      RECT 78.64 3.78 78.965 4.16 ;
      RECT 77.195 3.71 77.525 4.04 ;
      RECT 76.48 3.71 76.8 4.625 ;
      RECT 76.48 3.71 76.81 4.245 ;
      RECT 68.24 3.94 68.6 4.365 ;
      RECT 68.24 2.4 68.58 4.365 ;
      RECT 62.5 3.175 63.23 3.505 ;
      RECT 62.65 2.4 62.95 3.505 ;
      RECT 62.65 2.4 68.58 2.7 ;
      RECT 64.535 9.345 64.905 9.715 ;
      RECT 64.57 5.77 64.87 9.715 ;
      RECT 63.13 5.77 64.87 7.065 ;
      RECT 60.335 5.55 63.43 6.845 ;
      RECT 63.13 3.81 63.43 7.065 ;
      RECT 60.335 4.27 60.635 6.845 ;
      RECT 63.855 4.805 64.185 5.16 ;
      RECT 61.95 4.845 64.185 5.145 ;
      RECT 61.95 3.71 62.25 5.145 ;
      RECT 60.03 4.27 60.76 4.6 ;
      RECT 62.925 3.815 63.705 4.16 ;
      RECT 63.38 3.78 63.705 4.16 ;
      RECT 61.935 3.71 62.265 4.04 ;
      RECT 61.22 3.71 61.54 4.625 ;
      RECT 61.22 3.71 61.55 4.245 ;
      RECT 52.98 3.94 53.34 4.365 ;
      RECT 52.98 2.4 53.32 4.365 ;
      RECT 47.24 3.175 47.97 3.505 ;
      RECT 47.39 2.4 47.69 3.505 ;
      RECT 47.39 2.4 53.32 2.7 ;
      RECT 49.275 9.345 49.645 9.715 ;
      RECT 49.31 5.77 49.61 9.715 ;
      RECT 47.87 5.77 49.61 7.065 ;
      RECT 45.075 5.55 48.17 6.845 ;
      RECT 47.87 3.81 48.17 7.065 ;
      RECT 45.075 4.27 45.375 6.845 ;
      RECT 48.595 4.805 48.925 5.16 ;
      RECT 46.69 4.845 48.925 5.145 ;
      RECT 46.69 3.71 46.99 5.145 ;
      RECT 44.77 4.27 45.5 4.6 ;
      RECT 47.665 3.815 48.445 4.16 ;
      RECT 48.12 3.78 48.445 4.16 ;
      RECT 46.675 3.71 47.005 4.04 ;
      RECT 45.96 3.71 46.28 4.625 ;
      RECT 45.96 3.71 46.29 4.245 ;
      RECT 37.72 3.94 38.08 4.365 ;
      RECT 37.72 2.4 38.06 4.365 ;
      RECT 31.98 3.175 32.71 3.505 ;
      RECT 32.13 2.4 32.43 3.505 ;
      RECT 32.13 2.4 38.06 2.7 ;
      RECT 34.015 9.345 34.385 9.715 ;
      RECT 34.05 5.77 34.35 9.715 ;
      RECT 32.61 5.77 34.35 7.065 ;
      RECT 29.815 5.55 32.91 6.845 ;
      RECT 32.61 3.81 32.91 7.065 ;
      RECT 29.815 4.27 30.115 6.845 ;
      RECT 33.335 4.805 33.665 5.16 ;
      RECT 31.43 4.845 33.665 5.145 ;
      RECT 31.43 3.71 31.73 5.145 ;
      RECT 29.51 4.27 30.24 4.6 ;
      RECT 32.405 3.815 33.185 4.16 ;
      RECT 32.86 3.78 33.185 4.16 ;
      RECT 31.415 3.71 31.745 4.04 ;
      RECT 30.7 3.71 31.02 4.625 ;
      RECT 30.7 3.71 31.03 4.245 ;
      RECT 103.45 7.205 103.83 12.465 ;
      RECT 97.295 3.15 98.025 3.48 ;
      RECT 95.605 3.165 96.335 3.495 ;
      RECT 94.57 3.15 95.3 3.5 ;
      RECT 88.19 7.205 88.57 12.465 ;
      RECT 82.035 3.15 82.765 3.48 ;
      RECT 80.345 3.165 81.075 3.495 ;
      RECT 79.31 3.15 80.04 3.5 ;
      RECT 72.93 7.205 73.31 12.465 ;
      RECT 66.775 3.15 67.505 3.48 ;
      RECT 65.085 3.165 65.815 3.495 ;
      RECT 64.05 3.15 64.78 3.5 ;
      RECT 57.67 7.205 58.05 12.465 ;
      RECT 51.515 3.15 52.245 3.48 ;
      RECT 49.825 3.165 50.555 3.495 ;
      RECT 48.79 3.15 49.52 3.5 ;
      RECT 42.41 7.205 42.79 12.465 ;
      RECT 36.255 3.15 36.985 3.48 ;
      RECT 34.565 3.165 35.295 3.495 ;
      RECT 33.53 3.15 34.26 3.5 ;
    LAYER via2 ;
      RECT 103.54 7.295 103.74 7.495 ;
      RECT 98.835 4.07 99.035 4.27 ;
      RECT 97.53 3.215 97.73 3.415 ;
      RECT 95.67 3.23 95.87 3.43 ;
      RECT 95.14 9.43 95.34 9.63 ;
      RECT 94.65 3.235 94.85 3.435 ;
      RECT 94.44 4.87 94.64 5.07 ;
      RECT 93.96 3.87 94.16 4.07 ;
      RECT 93.21 3.24 93.41 3.44 ;
      RECT 92.52 3.775 92.72 3.975 ;
      RECT 91.805 3.775 92.005 3.975 ;
      RECT 90.84 4.335 91.04 4.535 ;
      RECT 88.28 7.295 88.48 7.495 ;
      RECT 83.575 4.07 83.775 4.27 ;
      RECT 82.27 3.215 82.47 3.415 ;
      RECT 80.41 3.23 80.61 3.43 ;
      RECT 79.88 9.43 80.08 9.63 ;
      RECT 79.39 3.235 79.59 3.435 ;
      RECT 79.18 4.87 79.38 5.07 ;
      RECT 78.7 3.87 78.9 4.07 ;
      RECT 77.95 3.24 78.15 3.44 ;
      RECT 77.26 3.775 77.46 3.975 ;
      RECT 76.545 3.775 76.745 3.975 ;
      RECT 75.58 4.335 75.78 4.535 ;
      RECT 73.02 7.295 73.22 7.495 ;
      RECT 68.315 4.07 68.515 4.27 ;
      RECT 67.01 3.215 67.21 3.415 ;
      RECT 65.15 3.23 65.35 3.43 ;
      RECT 64.62 9.43 64.82 9.63 ;
      RECT 64.13 3.235 64.33 3.435 ;
      RECT 63.92 4.87 64.12 5.07 ;
      RECT 63.44 3.87 63.64 4.07 ;
      RECT 62.69 3.24 62.89 3.44 ;
      RECT 62 3.775 62.2 3.975 ;
      RECT 61.285 3.775 61.485 3.975 ;
      RECT 60.32 4.335 60.52 4.535 ;
      RECT 57.76 7.295 57.96 7.495 ;
      RECT 53.055 4.07 53.255 4.27 ;
      RECT 51.75 3.215 51.95 3.415 ;
      RECT 49.89 3.23 50.09 3.43 ;
      RECT 49.36 9.43 49.56 9.63 ;
      RECT 48.87 3.235 49.07 3.435 ;
      RECT 48.66 4.87 48.86 5.07 ;
      RECT 48.18 3.87 48.38 4.07 ;
      RECT 47.43 3.24 47.63 3.44 ;
      RECT 46.74 3.775 46.94 3.975 ;
      RECT 46.025 3.775 46.225 3.975 ;
      RECT 45.06 4.335 45.26 4.535 ;
      RECT 42.5 7.295 42.7 7.495 ;
      RECT 37.795 4.07 37.995 4.27 ;
      RECT 36.49 3.215 36.69 3.415 ;
      RECT 34.63 3.23 34.83 3.43 ;
      RECT 34.1 9.43 34.3 9.63 ;
      RECT 33.61 3.235 33.81 3.435 ;
      RECT 33.4 4.87 33.6 5.07 ;
      RECT 32.92 3.87 33.12 4.07 ;
      RECT 32.17 3.24 32.37 3.44 ;
      RECT 31.48 3.775 31.68 3.975 ;
      RECT 30.765 3.775 30.965 3.975 ;
      RECT 29.8 4.335 30 4.535 ;
    LAYER met2 ;
      RECT 26.23 10.69 103.725 10.86 ;
      RECT 103.555 9.565 103.725 10.86 ;
      RECT 26.23 8.545 26.4 10.86 ;
      RECT 103.525 9.565 103.875 9.915 ;
      RECT 26.165 8.545 26.455 8.895 ;
      RECT 100.365 8.51 100.685 8.835 ;
      RECT 100.395 7.985 100.565 8.835 ;
      RECT 100.395 7.985 100.57 8.335 ;
      RECT 100.395 7.985 101.37 8.16 ;
      RECT 101.195 3.26 101.37 8.16 ;
      RECT 101.14 3.26 101.49 3.61 ;
      RECT 101.165 8.945 101.49 9.27 ;
      RECT 100.05 9.035 101.49 9.205 ;
      RECT 100.05 3.69 100.21 9.205 ;
      RECT 100.365 3.66 100.685 3.98 ;
      RECT 100.05 3.69 100.685 3.86 ;
      RECT 98.79 3.98 99.08 4.36 ;
      RECT 98.76 3.995 99.1 4.345 ;
      RECT 97.5 4.835 97.76 5.155 ;
      RECT 97.56 3.13 97.7 5.155 ;
      RECT 97.385 3.69 97.7 4.06 ;
      RECT 97.455 3.245 97.7 4.06 ;
      RECT 97.49 3.13 97.77 3.5 ;
      RECT 96.81 3.715 97.07 4.035 ;
      RECT 96.15 3.805 97.07 3.945 ;
      RECT 96.15 2.865 96.29 3.945 ;
      RECT 92.61 3.155 92.87 3.475 ;
      RECT 92.79 2.865 92.93 3.385 ;
      RECT 92.79 2.865 96.29 3.005 ;
      RECT 88.24 8.95 88.59 9.3 ;
      RECT 95.725 8.905 96.075 9.255 ;
      RECT 88.24 8.98 96.075 9.18 ;
      RECT 95.64 4.555 95.9 4.875 ;
      RECT 95.7 3.145 95.84 4.875 ;
      RECT 95.63 3.145 95.91 3.515 ;
      RECT 93.03 5.305 95.465 5.445 ;
      RECT 95.325 3.995 95.465 5.445 ;
      RECT 93.03 4.925 93.17 5.445 ;
      RECT 92.73 4.925 93.17 5.155 ;
      RECT 90.39 4.925 93.17 5.065 ;
      RECT 92.73 4.835 92.99 5.155 ;
      RECT 90.39 4.645 90.53 5.065 ;
      RECT 89.88 4.555 90.14 4.875 ;
      RECT 89.88 4.645 90.53 4.785 ;
      RECT 89.935 4.435 90.08 4.875 ;
      RECT 89.94 3.155 90.08 4.875 ;
      RECT 95.265 3.995 95.525 4.315 ;
      RECT 89.935 3.155 90.08 3.615 ;
      RECT 89.875 3.155 90.14 3.475 ;
      RECT 94.89 4.835 95.155 5.155 ;
      RECT 94.95 3.245 95.09 5.155 ;
      RECT 94.61 3.245 95.09 3.52 ;
      RECT 94.41 3.15 94.89 3.495 ;
      RECT 94.4 4.785 94.68 5.155 ;
      RECT 94.47 3.69 94.61 5.155 ;
      RECT 94.41 3.69 94.67 4.315 ;
      RECT 94.4 3.69 94.68 4.06 ;
      RECT 93.33 4.835 93.59 5.155 ;
      RECT 93.33 4.645 93.53 5.155 ;
      RECT 93.135 4.645 93.53 4.785 ;
      RECT 93.135 3.155 93.275 4.785 ;
      RECT 93.135 3.155 93.45 3.525 ;
      RECT 93.075 3.155 93.45 3.475 ;
      RECT 90.8 4.25 91.08 4.62 ;
      RECT 92.25 4.275 92.51 4.595 ;
      RECT 90.63 4.365 92.51 4.505 ;
      RECT 90.63 4.25 91.08 4.505 ;
      RECT 90.57 3.69 90.83 4.315 ;
      RECT 90.56 3.69 90.84 4.06 ;
      RECT 91.64 3.69 92.05 4.06 ;
      RECT 91.05 3.715 91.31 4.035 ;
      RECT 91.05 3.805 92.05 3.945 ;
      RECT 85.105 8.51 85.425 8.835 ;
      RECT 85.135 7.985 85.305 8.835 ;
      RECT 85.135 7.985 85.31 8.335 ;
      RECT 85.135 7.985 86.11 8.16 ;
      RECT 85.935 3.26 86.11 8.16 ;
      RECT 85.88 3.26 86.23 3.61 ;
      RECT 85.905 8.945 86.23 9.27 ;
      RECT 84.79 9.035 86.23 9.205 ;
      RECT 84.79 3.69 84.95 9.205 ;
      RECT 85.105 3.66 85.425 3.98 ;
      RECT 84.79 3.69 85.425 3.86 ;
      RECT 83.53 3.98 83.82 4.36 ;
      RECT 83.5 3.995 83.84 4.345 ;
      RECT 82.24 4.835 82.5 5.155 ;
      RECT 82.3 3.13 82.44 5.155 ;
      RECT 82.125 3.69 82.44 4.06 ;
      RECT 82.195 3.245 82.44 4.06 ;
      RECT 82.23 3.13 82.51 3.5 ;
      RECT 81.55 3.715 81.81 4.035 ;
      RECT 80.89 3.805 81.81 3.945 ;
      RECT 80.89 2.865 81.03 3.945 ;
      RECT 77.35 3.155 77.61 3.475 ;
      RECT 77.53 2.865 77.67 3.385 ;
      RECT 77.53 2.865 81.03 3.005 ;
      RECT 72.98 8.95 73.33 9.3 ;
      RECT 80.47 8.905 80.82 9.255 ;
      RECT 72.98 8.98 80.82 9.18 ;
      RECT 80.38 4.555 80.64 4.875 ;
      RECT 80.44 3.145 80.58 4.875 ;
      RECT 80.37 3.145 80.65 3.515 ;
      RECT 77.77 5.305 80.205 5.445 ;
      RECT 80.065 3.995 80.205 5.445 ;
      RECT 77.77 4.925 77.91 5.445 ;
      RECT 77.47 4.925 77.91 5.155 ;
      RECT 75.13 4.925 77.91 5.065 ;
      RECT 77.47 4.835 77.73 5.155 ;
      RECT 75.13 4.645 75.27 5.065 ;
      RECT 74.62 4.555 74.88 4.875 ;
      RECT 74.62 4.645 75.27 4.785 ;
      RECT 74.675 4.435 74.82 4.875 ;
      RECT 74.68 3.155 74.82 4.875 ;
      RECT 80.005 3.995 80.265 4.315 ;
      RECT 74.675 3.155 74.82 3.615 ;
      RECT 74.615 3.155 74.88 3.475 ;
      RECT 79.63 4.835 79.895 5.155 ;
      RECT 79.69 3.245 79.83 5.155 ;
      RECT 79.35 3.245 79.83 3.52 ;
      RECT 79.15 3.15 79.63 3.495 ;
      RECT 79.14 4.785 79.42 5.155 ;
      RECT 79.21 3.69 79.35 5.155 ;
      RECT 79.15 3.69 79.41 4.315 ;
      RECT 79.14 3.69 79.42 4.06 ;
      RECT 78.07 4.835 78.33 5.155 ;
      RECT 78.07 4.645 78.27 5.155 ;
      RECT 77.875 4.645 78.27 4.785 ;
      RECT 77.875 3.155 78.015 4.785 ;
      RECT 77.875 3.155 78.19 3.525 ;
      RECT 77.815 3.155 78.19 3.475 ;
      RECT 75.54 4.25 75.82 4.62 ;
      RECT 76.99 4.275 77.25 4.595 ;
      RECT 75.37 4.365 77.25 4.505 ;
      RECT 75.37 4.25 75.82 4.505 ;
      RECT 75.31 3.69 75.57 4.315 ;
      RECT 75.3 3.69 75.58 4.06 ;
      RECT 76.38 3.69 76.79 4.06 ;
      RECT 75.79 3.715 76.05 4.035 ;
      RECT 75.79 3.805 76.79 3.945 ;
      RECT 69.845 8.51 70.165 8.835 ;
      RECT 69.875 7.985 70.045 8.835 ;
      RECT 69.875 7.985 70.05 8.335 ;
      RECT 69.875 7.985 70.85 8.16 ;
      RECT 70.675 3.26 70.85 8.16 ;
      RECT 70.62 3.26 70.97 3.61 ;
      RECT 70.645 8.945 70.97 9.27 ;
      RECT 69.53 9.035 70.97 9.205 ;
      RECT 69.53 3.69 69.69 9.205 ;
      RECT 69.845 3.66 70.165 3.98 ;
      RECT 69.53 3.69 70.165 3.86 ;
      RECT 68.27 3.98 68.56 4.36 ;
      RECT 68.24 3.995 68.58 4.345 ;
      RECT 66.98 4.835 67.24 5.155 ;
      RECT 67.04 3.13 67.18 5.155 ;
      RECT 66.865 3.69 67.18 4.06 ;
      RECT 66.935 3.245 67.18 4.06 ;
      RECT 66.97 3.13 67.25 3.5 ;
      RECT 66.29 3.715 66.55 4.035 ;
      RECT 65.63 3.805 66.55 3.945 ;
      RECT 65.63 2.865 65.77 3.945 ;
      RECT 62.09 3.155 62.35 3.475 ;
      RECT 62.27 2.865 62.41 3.385 ;
      RECT 62.27 2.865 65.77 3.005 ;
      RECT 57.765 8.95 58.115 9.3 ;
      RECT 65.205 8.905 65.555 9.255 ;
      RECT 57.765 8.98 65.555 9.18 ;
      RECT 65.12 4.555 65.38 4.875 ;
      RECT 65.18 3.145 65.32 4.875 ;
      RECT 65.11 3.145 65.39 3.515 ;
      RECT 62.51 5.305 64.945 5.445 ;
      RECT 64.805 3.995 64.945 5.445 ;
      RECT 62.51 4.925 62.65 5.445 ;
      RECT 62.21 4.925 62.65 5.155 ;
      RECT 59.87 4.925 62.65 5.065 ;
      RECT 62.21 4.835 62.47 5.155 ;
      RECT 59.87 4.645 60.01 5.065 ;
      RECT 59.36 4.555 59.62 4.875 ;
      RECT 59.36 4.645 60.01 4.785 ;
      RECT 59.415 4.435 59.56 4.875 ;
      RECT 59.42 3.155 59.56 4.875 ;
      RECT 64.745 3.995 65.005 4.315 ;
      RECT 59.415 3.155 59.56 3.615 ;
      RECT 59.355 3.155 59.62 3.475 ;
      RECT 64.37 4.835 64.635 5.155 ;
      RECT 64.43 3.245 64.57 5.155 ;
      RECT 64.09 3.245 64.57 3.52 ;
      RECT 63.89 3.15 64.37 3.495 ;
      RECT 63.88 4.785 64.16 5.155 ;
      RECT 63.95 3.69 64.09 5.155 ;
      RECT 63.89 3.69 64.15 4.315 ;
      RECT 63.88 3.69 64.16 4.06 ;
      RECT 62.81 4.835 63.07 5.155 ;
      RECT 62.81 4.645 63.01 5.155 ;
      RECT 62.615 4.645 63.01 4.785 ;
      RECT 62.615 3.155 62.755 4.785 ;
      RECT 62.615 3.155 62.93 3.525 ;
      RECT 62.555 3.155 62.93 3.475 ;
      RECT 60.28 4.25 60.56 4.62 ;
      RECT 61.73 4.275 61.99 4.595 ;
      RECT 60.11 4.365 61.99 4.505 ;
      RECT 60.11 4.25 60.56 4.505 ;
      RECT 60.05 3.69 60.31 4.315 ;
      RECT 60.04 3.69 60.32 4.06 ;
      RECT 61.12 3.69 61.53 4.06 ;
      RECT 60.53 3.715 60.79 4.035 ;
      RECT 60.53 3.805 61.53 3.945 ;
      RECT 54.585 8.51 54.905 8.835 ;
      RECT 54.615 7.985 54.785 8.835 ;
      RECT 54.615 7.985 54.79 8.335 ;
      RECT 54.615 7.985 55.59 8.16 ;
      RECT 55.415 3.26 55.59 8.16 ;
      RECT 55.36 3.26 55.71 3.61 ;
      RECT 55.385 8.945 55.71 9.27 ;
      RECT 54.27 9.035 55.71 9.205 ;
      RECT 54.27 3.69 54.43 9.205 ;
      RECT 54.585 3.66 54.905 3.98 ;
      RECT 54.27 3.69 54.905 3.86 ;
      RECT 53.01 3.98 53.3 4.36 ;
      RECT 52.98 3.995 53.32 4.345 ;
      RECT 51.72 4.835 51.98 5.155 ;
      RECT 51.78 3.13 51.92 5.155 ;
      RECT 51.605 3.69 51.92 4.06 ;
      RECT 51.675 3.245 51.92 4.06 ;
      RECT 51.71 3.13 51.99 3.5 ;
      RECT 51.03 3.715 51.29 4.035 ;
      RECT 50.37 3.805 51.29 3.945 ;
      RECT 50.37 2.865 50.51 3.945 ;
      RECT 46.83 3.155 47.09 3.475 ;
      RECT 47.01 2.865 47.15 3.385 ;
      RECT 47.01 2.865 50.51 3.005 ;
      RECT 42.505 8.95 42.855 9.3 ;
      RECT 49.945 8.905 50.295 9.255 ;
      RECT 42.505 8.98 50.295 9.18 ;
      RECT 49.86 4.555 50.12 4.875 ;
      RECT 49.92 3.145 50.06 4.875 ;
      RECT 49.85 3.145 50.13 3.515 ;
      RECT 47.25 5.305 49.685 5.445 ;
      RECT 49.545 3.995 49.685 5.445 ;
      RECT 47.25 4.925 47.39 5.445 ;
      RECT 46.95 4.925 47.39 5.155 ;
      RECT 44.61 4.925 47.39 5.065 ;
      RECT 46.95 4.835 47.21 5.155 ;
      RECT 44.61 4.645 44.75 5.065 ;
      RECT 44.1 4.555 44.36 4.875 ;
      RECT 44.1 4.645 44.75 4.785 ;
      RECT 44.155 4.435 44.3 4.875 ;
      RECT 44.16 3.155 44.3 4.875 ;
      RECT 49.485 3.995 49.745 4.315 ;
      RECT 44.155 3.155 44.3 3.615 ;
      RECT 44.095 3.155 44.36 3.475 ;
      RECT 49.11 4.835 49.375 5.155 ;
      RECT 49.17 3.245 49.31 5.155 ;
      RECT 48.83 3.245 49.31 3.52 ;
      RECT 48.63 3.15 49.11 3.495 ;
      RECT 48.62 4.785 48.9 5.155 ;
      RECT 48.69 3.69 48.83 5.155 ;
      RECT 48.63 3.69 48.89 4.315 ;
      RECT 48.62 3.69 48.9 4.06 ;
      RECT 47.55 4.835 47.81 5.155 ;
      RECT 47.55 4.645 47.75 5.155 ;
      RECT 47.355 4.645 47.75 4.785 ;
      RECT 47.355 3.155 47.495 4.785 ;
      RECT 47.355 3.155 47.67 3.525 ;
      RECT 47.295 3.155 47.67 3.475 ;
      RECT 45.02 4.25 45.3 4.62 ;
      RECT 46.47 4.275 46.73 4.595 ;
      RECT 44.85 4.365 46.73 4.505 ;
      RECT 44.85 4.25 45.3 4.505 ;
      RECT 44.79 3.69 45.05 4.315 ;
      RECT 44.78 3.69 45.06 4.06 ;
      RECT 45.86 3.69 46.27 4.06 ;
      RECT 45.27 3.715 45.53 4.035 ;
      RECT 45.27 3.805 46.27 3.945 ;
      RECT 39.325 8.51 39.645 8.835 ;
      RECT 39.355 7.985 39.525 8.835 ;
      RECT 39.355 7.985 39.53 8.335 ;
      RECT 39.355 7.985 40.33 8.16 ;
      RECT 40.155 3.26 40.33 8.16 ;
      RECT 40.1 3.26 40.45 3.61 ;
      RECT 40.125 8.945 40.45 9.27 ;
      RECT 39.01 9.035 40.45 9.205 ;
      RECT 39.01 3.69 39.17 9.205 ;
      RECT 39.325 3.66 39.645 3.98 ;
      RECT 39.01 3.69 39.645 3.86 ;
      RECT 37.75 3.98 38.04 4.36 ;
      RECT 37.72 3.995 38.06 4.345 ;
      RECT 36.46 4.835 36.72 5.155 ;
      RECT 36.52 3.13 36.66 5.155 ;
      RECT 36.345 3.69 36.66 4.06 ;
      RECT 36.415 3.245 36.66 4.06 ;
      RECT 36.45 3.13 36.73 3.5 ;
      RECT 35.77 3.715 36.03 4.035 ;
      RECT 35.11 3.805 36.03 3.945 ;
      RECT 35.11 2.865 35.25 3.945 ;
      RECT 31.57 3.155 31.83 3.475 ;
      RECT 31.75 2.865 31.89 3.385 ;
      RECT 31.75 2.865 35.25 3.005 ;
      RECT 26.54 9.285 26.83 9.635 ;
      RECT 26.54 9.34 27.795 9.51 ;
      RECT 27.625 8.975 27.795 9.51 ;
      RECT 34.685 8.895 35.035 9.245 ;
      RECT 27.625 8.975 35.035 9.145 ;
      RECT 34.6 4.555 34.86 4.875 ;
      RECT 34.66 3.145 34.8 4.875 ;
      RECT 34.59 3.145 34.87 3.515 ;
      RECT 31.99 5.305 34.425 5.445 ;
      RECT 34.285 3.995 34.425 5.445 ;
      RECT 31.99 4.925 32.13 5.445 ;
      RECT 31.69 4.925 32.13 5.155 ;
      RECT 29.35 4.925 32.13 5.065 ;
      RECT 31.69 4.835 31.95 5.155 ;
      RECT 29.35 4.645 29.49 5.065 ;
      RECT 28.84 4.555 29.1 4.875 ;
      RECT 28.84 4.645 29.49 4.785 ;
      RECT 28.895 4.435 29.04 4.875 ;
      RECT 28.9 3.155 29.04 4.875 ;
      RECT 34.225 3.995 34.485 4.315 ;
      RECT 28.895 3.155 29.04 3.615 ;
      RECT 28.835 3.155 29.1 3.475 ;
      RECT 33.85 4.835 34.115 5.155 ;
      RECT 33.91 3.245 34.05 5.155 ;
      RECT 33.57 3.245 34.05 3.52 ;
      RECT 33.37 3.15 33.85 3.495 ;
      RECT 33.36 4.785 33.64 5.155 ;
      RECT 33.43 3.69 33.57 5.155 ;
      RECT 33.37 3.69 33.63 4.315 ;
      RECT 33.36 3.69 33.64 4.06 ;
      RECT 32.29 4.835 32.55 5.155 ;
      RECT 32.29 4.645 32.49 5.155 ;
      RECT 32.095 4.645 32.49 4.785 ;
      RECT 32.095 3.155 32.235 4.785 ;
      RECT 32.095 3.155 32.41 3.525 ;
      RECT 32.035 3.155 32.41 3.475 ;
      RECT 29.76 4.25 30.04 4.62 ;
      RECT 31.21 4.275 31.47 4.595 ;
      RECT 29.59 4.365 31.47 4.505 ;
      RECT 29.59 4.25 30.04 4.505 ;
      RECT 29.53 3.69 29.79 4.315 ;
      RECT 29.52 3.69 29.8 4.06 ;
      RECT 30.6 3.69 31.01 4.06 ;
      RECT 30.01 3.715 30.27 4.035 ;
      RECT 30.01 3.805 31.01 3.945 ;
      RECT 103.45 7.205 103.83 7.585 ;
      RECT 95.055 9.345 95.425 9.715 ;
      RECT 93.92 3.69 94.2 4.155 ;
      RECT 93.68 3.155 93.96 3.5 ;
      RECT 92.48 3.69 92.76 4.06 ;
      RECT 88.19 7.205 88.57 7.585 ;
      RECT 79.795 9.345 80.165 9.715 ;
      RECT 78.66 3.69 78.94 4.155 ;
      RECT 78.42 3.155 78.7 3.5 ;
      RECT 77.22 3.69 77.5 4.06 ;
      RECT 72.93 7.205 73.31 7.585 ;
      RECT 64.535 9.345 64.905 9.715 ;
      RECT 63.4 3.69 63.68 4.155 ;
      RECT 63.16 3.155 63.44 3.5 ;
      RECT 61.96 3.69 62.24 4.06 ;
      RECT 57.67 7.205 58.05 7.585 ;
      RECT 49.275 9.345 49.645 9.715 ;
      RECT 48.14 3.69 48.42 4.155 ;
      RECT 47.9 3.155 48.18 3.5 ;
      RECT 46.7 3.69 46.98 4.06 ;
      RECT 42.41 7.205 42.79 7.585 ;
      RECT 34.015 9.345 34.385 9.715 ;
      RECT 32.88 3.69 33.16 4.155 ;
      RECT 32.64 3.155 32.92 3.5 ;
      RECT 31.44 3.69 31.72 4.06 ;
    LAYER via1 ;
      RECT 103.625 9.665 103.775 9.815 ;
      RECT 103.565 7.32 103.715 7.47 ;
      RECT 101.255 9.03 101.405 9.18 ;
      RECT 101.24 3.36 101.39 3.51 ;
      RECT 100.45 3.745 100.6 3.895 ;
      RECT 100.45 8.615 100.6 8.765 ;
      RECT 98.86 4.095 99.01 4.245 ;
      RECT 97.555 3.24 97.705 3.39 ;
      RECT 97.555 4.92 97.705 5.07 ;
      RECT 96.865 3.8 97.015 3.95 ;
      RECT 95.825 9.005 95.975 9.155 ;
      RECT 95.695 3.24 95.845 3.39 ;
      RECT 95.695 4.64 95.845 4.79 ;
      RECT 95.32 4.08 95.47 4.23 ;
      RECT 95.165 9.455 95.315 9.605 ;
      RECT 94.945 4.92 95.095 5.07 ;
      RECT 94.465 3.24 94.615 3.39 ;
      RECT 94.465 4.08 94.615 4.23 ;
      RECT 93.985 3.8 94.135 3.95 ;
      RECT 93.745 3.24 93.895 3.39 ;
      RECT 93.385 4.92 93.535 5.07 ;
      RECT 93.13 3.24 93.28 3.39 ;
      RECT 92.785 4.92 92.935 5.07 ;
      RECT 92.665 3.24 92.815 3.39 ;
      RECT 92.545 3.8 92.695 3.95 ;
      RECT 92.305 4.36 92.455 4.51 ;
      RECT 91.105 3.8 91.255 3.95 ;
      RECT 90.625 4.08 90.775 4.23 ;
      RECT 89.935 4.64 90.085 4.79 ;
      RECT 89.93 3.24 90.08 3.39 ;
      RECT 88.34 9.05 88.49 9.2 ;
      RECT 88.305 7.32 88.455 7.47 ;
      RECT 85.995 9.03 86.145 9.18 ;
      RECT 85.98 3.36 86.13 3.51 ;
      RECT 85.19 3.745 85.34 3.895 ;
      RECT 85.19 8.615 85.34 8.765 ;
      RECT 83.6 4.095 83.75 4.245 ;
      RECT 82.295 3.24 82.445 3.39 ;
      RECT 82.295 4.92 82.445 5.07 ;
      RECT 81.605 3.8 81.755 3.95 ;
      RECT 80.57 9.005 80.72 9.155 ;
      RECT 80.435 3.24 80.585 3.39 ;
      RECT 80.435 4.64 80.585 4.79 ;
      RECT 80.06 4.08 80.21 4.23 ;
      RECT 79.905 9.455 80.055 9.605 ;
      RECT 79.685 4.92 79.835 5.07 ;
      RECT 79.205 3.24 79.355 3.39 ;
      RECT 79.205 4.08 79.355 4.23 ;
      RECT 78.725 3.8 78.875 3.95 ;
      RECT 78.485 3.24 78.635 3.39 ;
      RECT 78.125 4.92 78.275 5.07 ;
      RECT 77.87 3.24 78.02 3.39 ;
      RECT 77.525 4.92 77.675 5.07 ;
      RECT 77.405 3.24 77.555 3.39 ;
      RECT 77.285 3.8 77.435 3.95 ;
      RECT 77.045 4.36 77.195 4.51 ;
      RECT 75.845 3.8 75.995 3.95 ;
      RECT 75.365 4.08 75.515 4.23 ;
      RECT 74.675 4.64 74.825 4.79 ;
      RECT 74.67 3.24 74.82 3.39 ;
      RECT 73.08 9.05 73.23 9.2 ;
      RECT 73.045 7.32 73.195 7.47 ;
      RECT 70.735 9.03 70.885 9.18 ;
      RECT 70.72 3.36 70.87 3.51 ;
      RECT 69.93 3.745 70.08 3.895 ;
      RECT 69.93 8.615 70.08 8.765 ;
      RECT 68.34 4.095 68.49 4.245 ;
      RECT 67.035 3.24 67.185 3.39 ;
      RECT 67.035 4.92 67.185 5.07 ;
      RECT 66.345 3.8 66.495 3.95 ;
      RECT 65.305 9.005 65.455 9.155 ;
      RECT 65.175 3.24 65.325 3.39 ;
      RECT 65.175 4.64 65.325 4.79 ;
      RECT 64.8 4.08 64.95 4.23 ;
      RECT 64.645 9.455 64.795 9.605 ;
      RECT 64.425 4.92 64.575 5.07 ;
      RECT 63.945 3.24 64.095 3.39 ;
      RECT 63.945 4.08 64.095 4.23 ;
      RECT 63.465 3.8 63.615 3.95 ;
      RECT 63.225 3.24 63.375 3.39 ;
      RECT 62.865 4.92 63.015 5.07 ;
      RECT 62.61 3.24 62.76 3.39 ;
      RECT 62.265 4.92 62.415 5.07 ;
      RECT 62.145 3.24 62.295 3.39 ;
      RECT 62.025 3.8 62.175 3.95 ;
      RECT 61.785 4.36 61.935 4.51 ;
      RECT 60.585 3.8 60.735 3.95 ;
      RECT 60.105 4.08 60.255 4.23 ;
      RECT 59.415 4.64 59.565 4.79 ;
      RECT 59.41 3.24 59.56 3.39 ;
      RECT 57.865 9.05 58.015 9.2 ;
      RECT 57.785 7.32 57.935 7.47 ;
      RECT 55.475 9.03 55.625 9.18 ;
      RECT 55.46 3.36 55.61 3.51 ;
      RECT 54.67 3.745 54.82 3.895 ;
      RECT 54.67 8.615 54.82 8.765 ;
      RECT 53.08 4.095 53.23 4.245 ;
      RECT 51.775 3.24 51.925 3.39 ;
      RECT 51.775 4.92 51.925 5.07 ;
      RECT 51.085 3.8 51.235 3.95 ;
      RECT 50.045 9.005 50.195 9.155 ;
      RECT 49.915 3.24 50.065 3.39 ;
      RECT 49.915 4.64 50.065 4.79 ;
      RECT 49.54 4.08 49.69 4.23 ;
      RECT 49.385 9.455 49.535 9.605 ;
      RECT 49.165 4.92 49.315 5.07 ;
      RECT 48.685 3.24 48.835 3.39 ;
      RECT 48.685 4.08 48.835 4.23 ;
      RECT 48.205 3.8 48.355 3.95 ;
      RECT 47.965 3.24 48.115 3.39 ;
      RECT 47.605 4.92 47.755 5.07 ;
      RECT 47.35 3.24 47.5 3.39 ;
      RECT 47.005 4.92 47.155 5.07 ;
      RECT 46.885 3.24 47.035 3.39 ;
      RECT 46.765 3.8 46.915 3.95 ;
      RECT 46.525 4.36 46.675 4.51 ;
      RECT 45.325 3.8 45.475 3.95 ;
      RECT 44.845 4.08 44.995 4.23 ;
      RECT 44.155 4.64 44.305 4.79 ;
      RECT 44.15 3.24 44.3 3.39 ;
      RECT 42.605 9.05 42.755 9.2 ;
      RECT 42.525 7.32 42.675 7.47 ;
      RECT 40.215 9.03 40.365 9.18 ;
      RECT 40.2 3.36 40.35 3.51 ;
      RECT 39.41 3.745 39.56 3.895 ;
      RECT 39.41 8.615 39.56 8.765 ;
      RECT 37.82 4.095 37.97 4.245 ;
      RECT 36.515 3.24 36.665 3.39 ;
      RECT 36.515 4.92 36.665 5.07 ;
      RECT 35.825 3.8 35.975 3.95 ;
      RECT 34.785 8.995 34.935 9.145 ;
      RECT 34.655 3.24 34.805 3.39 ;
      RECT 34.655 4.64 34.805 4.79 ;
      RECT 34.28 4.08 34.43 4.23 ;
      RECT 34.125 9.455 34.275 9.605 ;
      RECT 33.905 4.92 34.055 5.07 ;
      RECT 33.425 3.24 33.575 3.39 ;
      RECT 33.425 4.08 33.575 4.23 ;
      RECT 32.945 3.8 33.095 3.95 ;
      RECT 32.705 3.24 32.855 3.39 ;
      RECT 32.345 4.92 32.495 5.07 ;
      RECT 32.09 3.24 32.24 3.39 ;
      RECT 31.745 4.92 31.895 5.07 ;
      RECT 31.625 3.24 31.775 3.39 ;
      RECT 31.505 3.8 31.655 3.95 ;
      RECT 31.265 4.36 31.415 4.51 ;
      RECT 30.065 3.8 30.215 3.95 ;
      RECT 29.585 4.08 29.735 4.23 ;
      RECT 28.895 4.64 29.045 4.79 ;
      RECT 28.89 3.24 29.04 3.39 ;
      RECT 26.61 9.385 26.76 9.535 ;
      RECT 26.235 8.645 26.385 8.795 ;
    LAYER met1 ;
      RECT 103.49 10.06 103.785 10.29 ;
      RECT 103.55 9.565 103.725 10.29 ;
      RECT 103.525 9.565 103.875 9.915 ;
      RECT 103.55 8.58 103.72 10.29 ;
      RECT 103.49 8.58 103.78 8.81 ;
      RECT 102.5 10.06 102.795 10.29 ;
      RECT 102.56 8.58 102.73 10.29 ;
      RECT 102.5 8.58 102.79 8.81 ;
      RECT 102.5 8.615 103.35 8.775 ;
      RECT 103.185 8.21 103.35 8.775 ;
      RECT 102.5 8.61 102.895 8.775 ;
      RECT 103.12 8.21 103.41 8.44 ;
      RECT 103.12 8.24 103.58 8.41 ;
      RECT 103.085 4.025 103.405 4.26 ;
      RECT 103.085 4.055 103.575 4.225 ;
      RECT 103.085 3.69 103.275 4.26 ;
      RECT 102.5 3.655 102.79 3.885 ;
      RECT 102.5 3.69 103.275 3.86 ;
      RECT 102.56 2.175 102.73 3.885 ;
      RECT 102.5 2.175 102.795 2.405 ;
      RECT 102.13 4.025 102.42 4.255 ;
      RECT 102.13 4.055 102.59 4.225 ;
      RECT 102.195 2.95 102.36 4.255 ;
      RECT 100.71 2.915 101 3.145 ;
      RECT 100.71 2.95 102.36 3.12 ;
      RECT 100.77 2.175 100.94 3.145 ;
      RECT 100.71 2.175 101 2.405 ;
      RECT 100.71 10.06 101 10.29 ;
      RECT 100.77 9.32 100.94 10.29 ;
      RECT 100.77 9.41 102.36 9.58 ;
      RECT 102.19 8.21 102.36 9.58 ;
      RECT 100.71 9.32 101 9.55 ;
      RECT 102.13 8.21 102.42 8.44 ;
      RECT 102.13 8.24 102.59 8.41 ;
      RECT 98.76 3.995 99.1 4.345 ;
      RECT 98.85 3.32 99.02 4.345 ;
      RECT 101.14 3.26 101.49 3.61 ;
      RECT 98.85 3.32 101.49 3.49 ;
      RECT 100.97 3.315 101.49 3.49 ;
      RECT 101.165 8.945 101.49 9.27 ;
      RECT 95.725 8.905 96.075 9.255 ;
      RECT 101.14 8.95 101.49 9.18 ;
      RECT 95.525 8.95 96.075 9.18 ;
      RECT 100.97 8.975 101.49 9.15 ;
      RECT 95.355 8.98 96.075 9.15 ;
      RECT 95.415 8.975 101.49 9.145 ;
      RECT 100.365 3.66 100.685 3.98 ;
      RECT 100.34 3.655 100.63 3.885 ;
      RECT 100.33 3.685 100.685 3.86 ;
      RECT 100.165 3.685 100.685 3.855 ;
      RECT 100.365 8.545 100.685 8.835 ;
      RECT 100.34 8.58 100.685 8.81 ;
      RECT 100.165 8.61 100.685 8.78 ;
      RECT 97.47 3.185 97.79 3.445 ;
      RECT 97.035 3.2 97.325 3.43 ;
      RECT 97.035 3.245 97.79 3.385 ;
      RECT 97.47 4.865 97.79 5.125 ;
      RECT 97.035 4.88 97.325 5.11 ;
      RECT 97.035 4.925 97.79 5.065 ;
      RECT 96.795 4.32 97.085 4.55 ;
      RECT 96.795 4.365 97.37 4.505 ;
      RECT 97.23 4.225 97.49 4.365 ;
      RECT 97.275 4.04 97.565 4.27 ;
      RECT 95.43 4.225 96.53 4.365 ;
      RECT 95.235 4.025 95.555 4.285 ;
      RECT 96.315 4.04 96.605 4.27 ;
      RECT 95.235 4.04 95.645 4.285 ;
      RECT 95.61 3.185 95.93 3.445 ;
      RECT 96.075 3.2 96.365 3.43 ;
      RECT 95.61 3.245 96.365 3.385 ;
      RECT 93.225 4.365 93.4 4.69 ;
      RECT 92.91 4.45 95.09 4.59 ;
      RECT 94.95 3.46 95.09 4.59 ;
      RECT 92.91 4.365 94.205 4.59 ;
      RECT 93.915 4.32 94.205 4.59 ;
      RECT 92.91 4.085 93.245 4.59 ;
      RECT 92.955 4.04 93.245 4.59 ;
      RECT 95.835 3.76 96.125 3.99 ;
      RECT 94.95 3.665 96.05 3.805 ;
      RECT 94.875 3.46 95.165 3.71 ;
      RECT 95.095 10.06 95.385 10.29 ;
      RECT 95.155 9.32 95.325 10.29 ;
      RECT 95.055 9.345 95.425 9.715 ;
      RECT 95.095 9.32 95.385 9.715 ;
      RECT 94.86 4.865 95.185 5.125 ;
      RECT 94.86 4.88 95.38 5.11 ;
      RECT 93.435 3.76 93.725 3.99 ;
      RECT 93.585 3.365 93.725 3.99 ;
      RECT 93.585 3.365 93.89 3.505 ;
      RECT 94.38 3.185 94.7 3.445 ;
      RECT 93.66 3.185 93.98 3.445 ;
      RECT 94.155 3.2 94.7 3.43 ;
      RECT 93.66 3.245 94.7 3.385 ;
      RECT 93.3 4.865 93.62 5.125 ;
      RECT 93.195 4.88 93.62 5.11 ;
      RECT 91.275 4.32 91.565 4.55 ;
      RECT 91.275 4.32 91.73 4.505 ;
      RECT 91.59 3.845 91.73 4.505 ;
      RECT 91.71 3.245 91.85 3.985 ;
      RECT 92.58 3.185 92.9 3.445 ;
      RECT 91.755 3.2 92.045 3.43 ;
      RECT 91.71 3.245 92.9 3.385 ;
      RECT 92.46 3.745 92.78 4.005 ;
      RECT 91.995 3.76 92.285 3.99 ;
      RECT 91.995 3.805 92.78 3.945 ;
      RECT 92.22 4.305 92.54 4.565 ;
      RECT 92.22 4.32 92.765 4.55 ;
      RECT 91.755 4.88 92.045 5.11 ;
      RECT 90.87 4.76 91.97 4.9 ;
      RECT 90.795 4.6 91.085 4.83 ;
      RECT 88.23 10.06 88.525 10.29 ;
      RECT 88.29 8.58 88.46 10.29 ;
      RECT 88.24 8.95 88.59 9.3 ;
      RECT 88.23 8.58 88.52 8.81 ;
      RECT 87.24 10.06 87.535 10.29 ;
      RECT 87.3 8.58 87.47 10.29 ;
      RECT 87.24 8.58 87.53 8.81 ;
      RECT 87.24 8.615 88.09 8.775 ;
      RECT 87.925 8.21 88.09 8.775 ;
      RECT 87.24 8.61 87.635 8.775 ;
      RECT 87.86 8.21 88.15 8.44 ;
      RECT 87.86 8.24 88.32 8.41 ;
      RECT 87.825 4.025 88.145 4.26 ;
      RECT 87.825 4.055 88.315 4.225 ;
      RECT 87.825 3.69 88.015 4.26 ;
      RECT 87.24 3.655 87.53 3.885 ;
      RECT 87.24 3.69 88.015 3.86 ;
      RECT 87.3 2.175 87.47 3.885 ;
      RECT 87.24 2.175 87.535 2.405 ;
      RECT 86.87 4.025 87.16 4.255 ;
      RECT 86.87 4.055 87.33 4.225 ;
      RECT 86.935 2.95 87.1 4.255 ;
      RECT 85.45 2.915 85.74 3.145 ;
      RECT 85.45 2.95 87.1 3.12 ;
      RECT 85.51 2.175 85.68 3.145 ;
      RECT 85.45 2.175 85.74 2.405 ;
      RECT 85.45 10.06 85.74 10.29 ;
      RECT 85.51 9.32 85.68 10.29 ;
      RECT 85.51 9.41 87.1 9.58 ;
      RECT 86.93 8.21 87.1 9.58 ;
      RECT 85.45 9.32 85.74 9.55 ;
      RECT 86.87 8.21 87.16 8.44 ;
      RECT 86.87 8.24 87.33 8.41 ;
      RECT 83.5 3.995 83.84 4.345 ;
      RECT 83.59 3.32 83.76 4.345 ;
      RECT 85.88 3.26 86.23 3.61 ;
      RECT 83.59 3.32 86.23 3.49 ;
      RECT 85.71 3.315 86.23 3.49 ;
      RECT 85.905 8.945 86.23 9.27 ;
      RECT 80.47 8.905 80.82 9.255 ;
      RECT 85.88 8.95 86.23 9.18 ;
      RECT 80.265 8.95 80.82 9.18 ;
      RECT 85.71 8.975 86.23 9.15 ;
      RECT 80.095 8.98 80.82 9.15 ;
      RECT 80.155 8.975 86.23 9.145 ;
      RECT 85.105 3.66 85.425 3.98 ;
      RECT 85.08 3.655 85.37 3.885 ;
      RECT 85.07 3.685 85.425 3.86 ;
      RECT 84.905 3.685 85.425 3.855 ;
      RECT 85.105 8.545 85.425 8.835 ;
      RECT 85.08 8.58 85.425 8.81 ;
      RECT 84.905 8.61 85.425 8.78 ;
      RECT 82.21 3.185 82.53 3.445 ;
      RECT 81.775 3.2 82.065 3.43 ;
      RECT 81.775 3.245 82.53 3.385 ;
      RECT 82.21 4.865 82.53 5.125 ;
      RECT 81.775 4.88 82.065 5.11 ;
      RECT 81.775 4.925 82.53 5.065 ;
      RECT 81.535 4.32 81.825 4.55 ;
      RECT 81.535 4.365 82.11 4.505 ;
      RECT 81.97 4.225 82.23 4.365 ;
      RECT 82.015 4.04 82.305 4.27 ;
      RECT 80.17 4.225 81.27 4.365 ;
      RECT 79.975 4.025 80.295 4.285 ;
      RECT 81.055 4.04 81.345 4.27 ;
      RECT 79.975 4.04 80.385 4.285 ;
      RECT 80.35 3.185 80.67 3.445 ;
      RECT 80.815 3.2 81.105 3.43 ;
      RECT 80.35 3.245 81.105 3.385 ;
      RECT 77.965 4.365 78.14 4.69 ;
      RECT 77.65 4.45 79.83 4.59 ;
      RECT 79.69 3.46 79.83 4.59 ;
      RECT 77.65 4.365 78.945 4.59 ;
      RECT 78.655 4.32 78.945 4.59 ;
      RECT 77.65 4.085 77.985 4.59 ;
      RECT 77.695 4.04 77.985 4.59 ;
      RECT 80.575 3.76 80.865 3.99 ;
      RECT 79.69 3.665 80.79 3.805 ;
      RECT 79.615 3.46 79.905 3.71 ;
      RECT 79.835 10.06 80.125 10.29 ;
      RECT 79.895 9.32 80.065 10.29 ;
      RECT 79.795 9.345 80.165 9.715 ;
      RECT 79.835 9.32 80.125 9.715 ;
      RECT 79.6 4.865 79.925 5.125 ;
      RECT 79.6 4.88 80.12 5.11 ;
      RECT 78.175 3.76 78.465 3.99 ;
      RECT 78.325 3.365 78.465 3.99 ;
      RECT 78.325 3.365 78.63 3.505 ;
      RECT 79.12 3.185 79.44 3.445 ;
      RECT 78.4 3.185 78.72 3.445 ;
      RECT 78.895 3.2 79.44 3.43 ;
      RECT 78.4 3.245 79.44 3.385 ;
      RECT 78.04 4.865 78.36 5.125 ;
      RECT 77.935 4.88 78.36 5.11 ;
      RECT 76.015 4.32 76.305 4.55 ;
      RECT 76.015 4.32 76.47 4.505 ;
      RECT 76.33 3.845 76.47 4.505 ;
      RECT 76.45 3.245 76.59 3.985 ;
      RECT 77.32 3.185 77.64 3.445 ;
      RECT 76.495 3.2 76.785 3.43 ;
      RECT 76.45 3.245 77.64 3.385 ;
      RECT 77.2 3.745 77.52 4.005 ;
      RECT 76.735 3.76 77.025 3.99 ;
      RECT 76.735 3.805 77.52 3.945 ;
      RECT 76.96 4.305 77.28 4.565 ;
      RECT 76.96 4.32 77.505 4.55 ;
      RECT 76.495 4.88 76.785 5.11 ;
      RECT 75.61 4.76 76.71 4.9 ;
      RECT 75.535 4.6 75.825 4.83 ;
      RECT 72.97 10.06 73.265 10.29 ;
      RECT 73.03 8.58 73.2 10.29 ;
      RECT 72.98 8.95 73.33 9.3 ;
      RECT 72.97 8.58 73.26 8.81 ;
      RECT 71.98 10.06 72.275 10.29 ;
      RECT 72.04 8.58 72.21 10.29 ;
      RECT 71.98 8.58 72.27 8.81 ;
      RECT 71.98 8.615 72.83 8.775 ;
      RECT 72.665 8.21 72.83 8.775 ;
      RECT 71.98 8.61 72.375 8.775 ;
      RECT 72.6 8.21 72.89 8.44 ;
      RECT 72.6 8.24 73.06 8.41 ;
      RECT 72.565 4.025 72.885 4.26 ;
      RECT 72.565 4.055 73.055 4.225 ;
      RECT 72.565 3.69 72.755 4.26 ;
      RECT 71.98 3.655 72.27 3.885 ;
      RECT 71.98 3.69 72.755 3.86 ;
      RECT 72.04 2.175 72.21 3.885 ;
      RECT 71.98 2.175 72.275 2.405 ;
      RECT 71.61 4.025 71.9 4.255 ;
      RECT 71.61 4.055 72.07 4.225 ;
      RECT 71.675 2.95 71.84 4.255 ;
      RECT 70.19 2.915 70.48 3.145 ;
      RECT 70.19 2.95 71.84 3.12 ;
      RECT 70.25 2.175 70.42 3.145 ;
      RECT 70.19 2.175 70.48 2.405 ;
      RECT 70.19 10.06 70.48 10.29 ;
      RECT 70.25 9.32 70.42 10.29 ;
      RECT 70.25 9.41 71.84 9.58 ;
      RECT 71.67 8.21 71.84 9.58 ;
      RECT 70.19 9.32 70.48 9.55 ;
      RECT 71.61 8.21 71.9 8.44 ;
      RECT 71.61 8.24 72.07 8.41 ;
      RECT 68.24 3.995 68.58 4.345 ;
      RECT 68.33 3.32 68.5 4.345 ;
      RECT 70.62 3.26 70.97 3.61 ;
      RECT 68.33 3.32 70.97 3.49 ;
      RECT 70.45 3.315 70.97 3.49 ;
      RECT 70.645 8.945 70.97 9.27 ;
      RECT 65.205 8.905 65.555 9.255 ;
      RECT 70.62 8.95 70.97 9.18 ;
      RECT 65.005 8.95 65.555 9.18 ;
      RECT 70.45 8.975 70.97 9.15 ;
      RECT 64.835 8.98 65.555 9.15 ;
      RECT 64.895 8.975 70.97 9.145 ;
      RECT 69.845 3.66 70.165 3.98 ;
      RECT 69.82 3.655 70.11 3.885 ;
      RECT 69.81 3.685 70.165 3.86 ;
      RECT 69.645 3.685 70.165 3.855 ;
      RECT 69.845 8.545 70.165 8.835 ;
      RECT 69.82 8.58 70.165 8.81 ;
      RECT 69.645 8.61 70.165 8.78 ;
      RECT 66.95 3.185 67.27 3.445 ;
      RECT 66.515 3.2 66.805 3.43 ;
      RECT 66.515 3.245 67.27 3.385 ;
      RECT 66.95 4.865 67.27 5.125 ;
      RECT 66.515 4.88 66.805 5.11 ;
      RECT 66.515 4.925 67.27 5.065 ;
      RECT 66.275 4.32 66.565 4.55 ;
      RECT 66.275 4.365 66.85 4.505 ;
      RECT 66.71 4.225 66.97 4.365 ;
      RECT 66.755 4.04 67.045 4.27 ;
      RECT 64.91 4.225 66.01 4.365 ;
      RECT 64.715 4.025 65.035 4.285 ;
      RECT 65.795 4.04 66.085 4.27 ;
      RECT 64.715 4.04 65.125 4.285 ;
      RECT 65.09 3.185 65.41 3.445 ;
      RECT 65.555 3.2 65.845 3.43 ;
      RECT 65.09 3.245 65.845 3.385 ;
      RECT 62.705 4.365 62.88 4.69 ;
      RECT 62.39 4.45 64.57 4.59 ;
      RECT 64.43 3.46 64.57 4.59 ;
      RECT 62.39 4.365 63.685 4.59 ;
      RECT 63.395 4.32 63.685 4.59 ;
      RECT 62.39 4.085 62.725 4.59 ;
      RECT 62.435 4.04 62.725 4.59 ;
      RECT 65.315 3.76 65.605 3.99 ;
      RECT 64.43 3.665 65.53 3.805 ;
      RECT 64.355 3.46 64.645 3.71 ;
      RECT 64.575 10.06 64.865 10.29 ;
      RECT 64.635 9.32 64.805 10.29 ;
      RECT 64.535 9.345 64.905 9.715 ;
      RECT 64.575 9.32 64.865 9.715 ;
      RECT 64.34 4.865 64.665 5.125 ;
      RECT 64.34 4.88 64.86 5.11 ;
      RECT 62.915 3.76 63.205 3.99 ;
      RECT 63.065 3.365 63.205 3.99 ;
      RECT 63.065 3.365 63.37 3.505 ;
      RECT 63.86 3.185 64.18 3.445 ;
      RECT 63.14 3.185 63.46 3.445 ;
      RECT 63.635 3.2 64.18 3.43 ;
      RECT 63.14 3.245 64.18 3.385 ;
      RECT 62.78 4.865 63.1 5.125 ;
      RECT 62.675 4.88 63.1 5.11 ;
      RECT 60.755 4.32 61.045 4.55 ;
      RECT 60.755 4.32 61.21 4.505 ;
      RECT 61.07 3.845 61.21 4.505 ;
      RECT 61.19 3.245 61.33 3.985 ;
      RECT 62.06 3.185 62.38 3.445 ;
      RECT 61.235 3.2 61.525 3.43 ;
      RECT 61.19 3.245 62.38 3.385 ;
      RECT 61.94 3.745 62.26 4.005 ;
      RECT 61.475 3.76 61.765 3.99 ;
      RECT 61.475 3.805 62.26 3.945 ;
      RECT 61.7 4.305 62.02 4.565 ;
      RECT 61.7 4.32 62.245 4.55 ;
      RECT 61.235 4.88 61.525 5.11 ;
      RECT 60.35 4.76 61.45 4.9 ;
      RECT 60.275 4.6 60.565 4.83 ;
      RECT 57.71 10.06 58.005 10.29 ;
      RECT 57.77 8.58 57.94 10.29 ;
      RECT 57.76 8.95 58.115 9.305 ;
      RECT 57.71 8.58 58 8.81 ;
      RECT 56.72 10.06 57.015 10.29 ;
      RECT 56.78 8.58 56.95 10.29 ;
      RECT 56.72 8.58 57.01 8.81 ;
      RECT 56.72 8.615 57.57 8.775 ;
      RECT 57.405 8.21 57.57 8.775 ;
      RECT 56.72 8.61 57.115 8.775 ;
      RECT 57.34 8.21 57.63 8.44 ;
      RECT 57.34 8.24 57.8 8.41 ;
      RECT 57.305 4.025 57.625 4.26 ;
      RECT 57.305 4.055 57.795 4.225 ;
      RECT 57.305 3.69 57.495 4.26 ;
      RECT 56.72 3.655 57.01 3.885 ;
      RECT 56.72 3.69 57.495 3.86 ;
      RECT 56.78 2.175 56.95 3.885 ;
      RECT 56.72 2.175 57.015 2.405 ;
      RECT 56.35 4.025 56.64 4.255 ;
      RECT 56.35 4.055 56.81 4.225 ;
      RECT 56.415 2.95 56.58 4.255 ;
      RECT 54.93 2.915 55.22 3.145 ;
      RECT 54.93 2.95 56.58 3.12 ;
      RECT 54.99 2.175 55.16 3.145 ;
      RECT 54.93 2.175 55.22 2.405 ;
      RECT 54.93 10.06 55.22 10.29 ;
      RECT 54.99 9.32 55.16 10.29 ;
      RECT 54.99 9.41 56.58 9.58 ;
      RECT 56.41 8.21 56.58 9.58 ;
      RECT 54.93 9.32 55.22 9.55 ;
      RECT 56.35 8.21 56.64 8.44 ;
      RECT 56.35 8.24 56.81 8.41 ;
      RECT 52.98 3.995 53.32 4.345 ;
      RECT 53.07 3.32 53.24 4.345 ;
      RECT 55.36 3.26 55.71 3.61 ;
      RECT 53.07 3.32 55.71 3.49 ;
      RECT 55.19 3.315 55.71 3.49 ;
      RECT 55.385 8.945 55.71 9.27 ;
      RECT 49.945 8.905 50.295 9.255 ;
      RECT 55.36 8.95 55.71 9.18 ;
      RECT 49.745 8.95 50.295 9.18 ;
      RECT 55.19 8.975 55.71 9.15 ;
      RECT 49.575 8.98 50.295 9.15 ;
      RECT 49.635 8.975 55.71 9.145 ;
      RECT 54.585 3.66 54.905 3.98 ;
      RECT 54.56 3.655 54.85 3.885 ;
      RECT 54.55 3.685 54.905 3.86 ;
      RECT 54.385 3.685 54.905 3.855 ;
      RECT 54.585 8.545 54.905 8.835 ;
      RECT 54.56 8.58 54.905 8.81 ;
      RECT 54.385 8.61 54.905 8.78 ;
      RECT 51.69 3.185 52.01 3.445 ;
      RECT 51.255 3.2 51.545 3.43 ;
      RECT 51.255 3.245 52.01 3.385 ;
      RECT 51.69 4.865 52.01 5.125 ;
      RECT 51.255 4.88 51.545 5.11 ;
      RECT 51.255 4.925 52.01 5.065 ;
      RECT 51.015 4.32 51.305 4.55 ;
      RECT 51.015 4.365 51.59 4.505 ;
      RECT 51.45 4.225 51.71 4.365 ;
      RECT 51.495 4.04 51.785 4.27 ;
      RECT 49.65 4.225 50.75 4.365 ;
      RECT 49.455 4.025 49.775 4.285 ;
      RECT 50.535 4.04 50.825 4.27 ;
      RECT 49.455 4.04 49.865 4.285 ;
      RECT 49.83 3.185 50.15 3.445 ;
      RECT 50.295 3.2 50.585 3.43 ;
      RECT 49.83 3.245 50.585 3.385 ;
      RECT 47.445 4.365 47.62 4.69 ;
      RECT 47.13 4.45 49.31 4.59 ;
      RECT 49.17 3.46 49.31 4.59 ;
      RECT 47.13 4.365 48.425 4.59 ;
      RECT 48.135 4.32 48.425 4.59 ;
      RECT 47.13 4.085 47.465 4.59 ;
      RECT 47.175 4.04 47.465 4.59 ;
      RECT 50.055 3.76 50.345 3.99 ;
      RECT 49.17 3.665 50.27 3.805 ;
      RECT 49.095 3.46 49.385 3.71 ;
      RECT 49.315 10.06 49.605 10.29 ;
      RECT 49.375 9.32 49.545 10.29 ;
      RECT 49.275 9.345 49.645 9.715 ;
      RECT 49.315 9.32 49.605 9.715 ;
      RECT 49.08 4.865 49.405 5.125 ;
      RECT 49.08 4.88 49.6 5.11 ;
      RECT 47.655 3.76 47.945 3.99 ;
      RECT 47.805 3.365 47.945 3.99 ;
      RECT 47.805 3.365 48.11 3.505 ;
      RECT 48.6 3.185 48.92 3.445 ;
      RECT 47.88 3.185 48.2 3.445 ;
      RECT 48.375 3.2 48.92 3.43 ;
      RECT 47.88 3.245 48.92 3.385 ;
      RECT 47.52 4.865 47.84 5.125 ;
      RECT 47.415 4.88 47.84 5.11 ;
      RECT 45.495 4.32 45.785 4.55 ;
      RECT 45.495 4.32 45.95 4.505 ;
      RECT 45.81 3.845 45.95 4.505 ;
      RECT 45.93 3.245 46.07 3.985 ;
      RECT 46.8 3.185 47.12 3.445 ;
      RECT 45.975 3.2 46.265 3.43 ;
      RECT 45.93 3.245 47.12 3.385 ;
      RECT 46.68 3.745 47 4.005 ;
      RECT 46.215 3.76 46.505 3.99 ;
      RECT 46.215 3.805 47 3.945 ;
      RECT 46.44 4.305 46.76 4.565 ;
      RECT 46.44 4.32 46.985 4.55 ;
      RECT 45.975 4.88 46.265 5.11 ;
      RECT 45.09 4.76 46.19 4.9 ;
      RECT 45.015 4.6 45.305 4.83 ;
      RECT 42.45 10.06 42.745 10.29 ;
      RECT 42.51 8.58 42.68 10.29 ;
      RECT 42.505 8.95 42.855 9.3 ;
      RECT 42.45 8.58 42.74 8.81 ;
      RECT 41.46 10.06 41.755 10.29 ;
      RECT 41.52 8.58 41.69 10.29 ;
      RECT 41.46 8.58 41.75 8.81 ;
      RECT 41.46 8.615 42.31 8.775 ;
      RECT 42.145 8.21 42.31 8.775 ;
      RECT 41.46 8.61 41.855 8.775 ;
      RECT 42.08 8.21 42.37 8.44 ;
      RECT 42.08 8.24 42.54 8.41 ;
      RECT 42.045 4.025 42.365 4.26 ;
      RECT 42.045 4.055 42.535 4.225 ;
      RECT 42.045 3.69 42.235 4.26 ;
      RECT 41.46 3.655 41.75 3.885 ;
      RECT 41.46 3.69 42.235 3.86 ;
      RECT 41.52 2.175 41.69 3.885 ;
      RECT 41.46 2.175 41.755 2.405 ;
      RECT 41.09 4.025 41.38 4.255 ;
      RECT 41.09 4.055 41.55 4.225 ;
      RECT 41.155 2.95 41.32 4.255 ;
      RECT 39.67 2.915 39.96 3.145 ;
      RECT 39.67 2.95 41.32 3.12 ;
      RECT 39.73 2.175 39.9 3.145 ;
      RECT 39.67 2.175 39.96 2.405 ;
      RECT 39.67 10.06 39.96 10.29 ;
      RECT 39.73 9.32 39.9 10.29 ;
      RECT 39.73 9.41 41.32 9.58 ;
      RECT 41.15 8.21 41.32 9.58 ;
      RECT 39.67 9.32 39.96 9.55 ;
      RECT 41.09 8.21 41.38 8.44 ;
      RECT 41.09 8.24 41.55 8.41 ;
      RECT 37.72 3.995 38.06 4.345 ;
      RECT 37.81 3.32 37.98 4.345 ;
      RECT 40.1 3.26 40.45 3.61 ;
      RECT 37.81 3.32 40.45 3.49 ;
      RECT 39.93 3.315 40.45 3.49 ;
      RECT 40.125 8.945 40.45 9.27 ;
      RECT 34.685 8.895 35.035 9.245 ;
      RECT 40.1 8.95 40.45 9.18 ;
      RECT 34.485 8.95 35.035 9.18 ;
      RECT 39.93 8.975 40.45 9.15 ;
      RECT 34.315 8.98 35.035 9.15 ;
      RECT 34.375 8.975 40.45 9.145 ;
      RECT 39.325 3.66 39.645 3.98 ;
      RECT 39.3 3.655 39.59 3.885 ;
      RECT 39.29 3.685 39.645 3.86 ;
      RECT 39.125 3.685 39.645 3.855 ;
      RECT 39.325 8.545 39.645 8.835 ;
      RECT 39.3 8.58 39.645 8.81 ;
      RECT 39.125 8.61 39.645 8.78 ;
      RECT 36.43 3.185 36.75 3.445 ;
      RECT 35.995 3.2 36.285 3.43 ;
      RECT 35.995 3.245 36.75 3.385 ;
      RECT 36.43 4.865 36.75 5.125 ;
      RECT 35.995 4.88 36.285 5.11 ;
      RECT 35.995 4.925 36.75 5.065 ;
      RECT 35.755 4.32 36.045 4.55 ;
      RECT 35.755 4.365 36.33 4.505 ;
      RECT 36.19 4.225 36.45 4.365 ;
      RECT 36.235 4.04 36.525 4.27 ;
      RECT 34.39 4.225 35.49 4.365 ;
      RECT 34.195 4.025 34.515 4.285 ;
      RECT 35.275 4.04 35.565 4.27 ;
      RECT 34.195 4.04 34.605 4.285 ;
      RECT 34.57 3.185 34.89 3.445 ;
      RECT 35.035 3.2 35.325 3.43 ;
      RECT 34.57 3.245 35.325 3.385 ;
      RECT 32.185 4.365 32.36 4.69 ;
      RECT 31.87 4.45 34.05 4.59 ;
      RECT 33.91 3.46 34.05 4.59 ;
      RECT 31.87 4.365 33.165 4.59 ;
      RECT 32.875 4.32 33.165 4.59 ;
      RECT 31.87 4.085 32.205 4.59 ;
      RECT 31.915 4.04 32.205 4.59 ;
      RECT 34.795 3.76 35.085 3.99 ;
      RECT 33.91 3.665 35.01 3.805 ;
      RECT 33.835 3.46 34.125 3.71 ;
      RECT 34.055 10.06 34.345 10.29 ;
      RECT 34.115 9.32 34.285 10.29 ;
      RECT 34.015 9.345 34.385 9.715 ;
      RECT 34.055 9.32 34.345 9.715 ;
      RECT 33.82 4.865 34.145 5.125 ;
      RECT 33.82 4.88 34.34 5.11 ;
      RECT 32.395 3.76 32.685 3.99 ;
      RECT 32.545 3.365 32.685 3.99 ;
      RECT 32.545 3.365 32.85 3.505 ;
      RECT 33.34 3.185 33.66 3.445 ;
      RECT 32.62 3.185 32.94 3.445 ;
      RECT 33.115 3.2 33.66 3.43 ;
      RECT 32.62 3.245 33.66 3.385 ;
      RECT 32.26 4.865 32.58 5.125 ;
      RECT 32.155 4.88 32.58 5.11 ;
      RECT 30.235 4.32 30.525 4.55 ;
      RECT 30.235 4.32 30.69 4.505 ;
      RECT 30.55 3.845 30.69 4.505 ;
      RECT 30.67 3.245 30.81 3.985 ;
      RECT 31.54 3.185 31.86 3.445 ;
      RECT 30.715 3.2 31.005 3.43 ;
      RECT 30.67 3.245 31.86 3.385 ;
      RECT 31.42 3.745 31.74 4.005 ;
      RECT 30.955 3.76 31.245 3.99 ;
      RECT 30.955 3.805 31.74 3.945 ;
      RECT 31.18 4.305 31.5 4.565 ;
      RECT 31.18 4.32 31.725 4.55 ;
      RECT 30.715 4.88 31.005 5.11 ;
      RECT 29.83 4.76 30.93 4.9 ;
      RECT 29.755 4.6 30.045 4.83 ;
      RECT 26.54 10.06 26.83 10.29 ;
      RECT 26.6 9.315 26.77 10.29 ;
      RECT 26.51 9.315 26.86 9.605 ;
      RECT 26.135 8.575 26.485 8.865 ;
      RECT 25.995 8.61 26.485 8.78 ;
      RECT 103.465 7.25 103.815 7.54 ;
      RECT 96.78 3.745 97.1 4.005 ;
      RECT 95.61 4.585 95.93 4.845 ;
      RECT 94.38 4.025 94.7 4.285 ;
      RECT 93.9 3.745 94.22 4.005 ;
      RECT 93.045 3.185 93.445 3.445 ;
      RECT 92.7 4.865 93.02 5.125 ;
      RECT 91.02 3.745 91.34 4.005 ;
      RECT 90.54 4.025 90.86 4.285 ;
      RECT 89.845 3.185 90.17 3.445 ;
      RECT 89.85 4.585 90.17 4.845 ;
      RECT 88.205 7.25 88.555 7.54 ;
      RECT 81.52 3.745 81.84 4.005 ;
      RECT 80.35 4.585 80.67 4.845 ;
      RECT 79.12 4.025 79.44 4.285 ;
      RECT 78.64 3.745 78.96 4.005 ;
      RECT 77.785 3.185 78.185 3.445 ;
      RECT 77.44 4.865 77.76 5.125 ;
      RECT 75.76 3.745 76.08 4.005 ;
      RECT 75.28 4.025 75.6 4.285 ;
      RECT 74.585 3.185 74.91 3.445 ;
      RECT 74.59 4.585 74.91 4.845 ;
      RECT 72.945 7.25 73.295 7.54 ;
      RECT 66.26 3.745 66.58 4.005 ;
      RECT 65.09 4.585 65.41 4.845 ;
      RECT 63.86 4.025 64.18 4.285 ;
      RECT 63.38 3.745 63.7 4.005 ;
      RECT 62.525 3.185 62.925 3.445 ;
      RECT 62.18 4.865 62.5 5.125 ;
      RECT 60.5 3.745 60.82 4.005 ;
      RECT 60.02 4.025 60.34 4.285 ;
      RECT 59.325 3.185 59.65 3.445 ;
      RECT 59.33 4.585 59.65 4.845 ;
      RECT 57.685 7.25 58.035 7.54 ;
      RECT 51 3.745 51.32 4.005 ;
      RECT 49.83 4.585 50.15 4.845 ;
      RECT 48.6 4.025 48.92 4.285 ;
      RECT 48.12 3.745 48.44 4.005 ;
      RECT 47.265 3.185 47.665 3.445 ;
      RECT 46.92 4.865 47.24 5.125 ;
      RECT 45.24 3.745 45.56 4.005 ;
      RECT 44.76 4.025 45.08 4.285 ;
      RECT 44.065 3.185 44.39 3.445 ;
      RECT 44.07 4.585 44.39 4.845 ;
      RECT 42.425 7.25 42.775 7.54 ;
      RECT 35.74 3.745 36.06 4.005 ;
      RECT 34.57 4.585 34.89 4.845 ;
      RECT 33.34 4.025 33.66 4.285 ;
      RECT 32.86 3.745 33.18 4.005 ;
      RECT 32.005 3.185 32.405 3.445 ;
      RECT 31.66 4.865 31.98 5.125 ;
      RECT 29.98 3.745 30.3 4.005 ;
      RECT 29.5 4.025 29.82 4.285 ;
      RECT 28.805 3.185 29.13 3.445 ;
      RECT 28.81 4.585 29.13 4.845 ;
    LAYER mcon ;
      RECT 103.555 7.31 103.725 7.48 ;
      RECT 103.55 8.61 103.72 8.78 ;
      RECT 103.55 10.09 103.72 10.26 ;
      RECT 103.18 8.24 103.35 8.41 ;
      RECT 103.175 4.055 103.345 4.225 ;
      RECT 102.56 2.205 102.73 2.375 ;
      RECT 102.56 3.685 102.73 3.855 ;
      RECT 102.56 8.61 102.73 8.78 ;
      RECT 102.56 10.09 102.73 10.26 ;
      RECT 102.19 4.055 102.36 4.225 ;
      RECT 102.19 8.24 102.36 8.41 ;
      RECT 101.2 3.315 101.37 3.485 ;
      RECT 101.2 8.98 101.37 9.15 ;
      RECT 100.77 2.205 100.94 2.375 ;
      RECT 100.77 2.945 100.94 3.115 ;
      RECT 100.77 9.35 100.94 9.52 ;
      RECT 100.77 10.09 100.94 10.26 ;
      RECT 100.4 3.685 100.57 3.855 ;
      RECT 100.4 8.61 100.57 8.78 ;
      RECT 97.335 4.07 97.505 4.24 ;
      RECT 97.095 3.23 97.265 3.4 ;
      RECT 97.095 4.91 97.265 5.08 ;
      RECT 96.855 3.79 97.025 3.96 ;
      RECT 96.855 4.35 97.025 4.52 ;
      RECT 96.375 4.07 96.545 4.24 ;
      RECT 96.135 3.23 96.305 3.4 ;
      RECT 95.895 3.79 96.065 3.96 ;
      RECT 95.685 4.63 95.855 4.8 ;
      RECT 95.585 8.98 95.755 9.15 ;
      RECT 95.415 4.07 95.585 4.24 ;
      RECT 95.155 9.35 95.325 9.52 ;
      RECT 95.155 10.09 95.325 10.26 ;
      RECT 95.15 4.91 95.32 5.08 ;
      RECT 94.935 3.49 95.105 3.66 ;
      RECT 94.455 4.07 94.625 4.24 ;
      RECT 94.215 3.23 94.385 3.4 ;
      RECT 93.975 3.79 94.145 3.96 ;
      RECT 93.975 4.35 94.145 4.52 ;
      RECT 93.495 3.79 93.665 3.96 ;
      RECT 93.255 4.91 93.425 5.08 ;
      RECT 93.215 3.23 93.385 3.4 ;
      RECT 93.015 4.07 93.185 4.24 ;
      RECT 92.775 4.91 92.945 5.08 ;
      RECT 92.535 4.35 92.705 4.52 ;
      RECT 92.055 3.79 92.225 3.96 ;
      RECT 91.815 3.23 91.985 3.4 ;
      RECT 91.815 4.91 91.985 5.08 ;
      RECT 91.335 4.35 91.505 4.52 ;
      RECT 91.095 3.79 91.265 3.96 ;
      RECT 90.855 4.63 91.025 4.8 ;
      RECT 90.615 4.07 90.785 4.24 ;
      RECT 89.92 3.23 90.09 3.4 ;
      RECT 89.92 4.63 90.09 4.8 ;
      RECT 88.295 7.31 88.465 7.48 ;
      RECT 88.29 8.61 88.46 8.78 ;
      RECT 88.29 10.09 88.46 10.26 ;
      RECT 87.92 8.24 88.09 8.41 ;
      RECT 87.915 4.055 88.085 4.225 ;
      RECT 87.3 2.205 87.47 2.375 ;
      RECT 87.3 3.685 87.47 3.855 ;
      RECT 87.3 8.61 87.47 8.78 ;
      RECT 87.3 10.09 87.47 10.26 ;
      RECT 86.93 4.055 87.1 4.225 ;
      RECT 86.93 8.24 87.1 8.41 ;
      RECT 85.94 3.315 86.11 3.485 ;
      RECT 85.94 8.98 86.11 9.15 ;
      RECT 85.51 2.205 85.68 2.375 ;
      RECT 85.51 2.945 85.68 3.115 ;
      RECT 85.51 9.35 85.68 9.52 ;
      RECT 85.51 10.09 85.68 10.26 ;
      RECT 85.14 3.685 85.31 3.855 ;
      RECT 85.14 8.61 85.31 8.78 ;
      RECT 82.075 4.07 82.245 4.24 ;
      RECT 81.835 3.23 82.005 3.4 ;
      RECT 81.835 4.91 82.005 5.08 ;
      RECT 81.595 3.79 81.765 3.96 ;
      RECT 81.595 4.35 81.765 4.52 ;
      RECT 81.115 4.07 81.285 4.24 ;
      RECT 80.875 3.23 81.045 3.4 ;
      RECT 80.635 3.79 80.805 3.96 ;
      RECT 80.425 4.63 80.595 4.8 ;
      RECT 80.325 8.98 80.495 9.15 ;
      RECT 80.155 4.07 80.325 4.24 ;
      RECT 79.895 9.35 80.065 9.52 ;
      RECT 79.895 10.09 80.065 10.26 ;
      RECT 79.89 4.91 80.06 5.08 ;
      RECT 79.675 3.49 79.845 3.66 ;
      RECT 79.195 4.07 79.365 4.24 ;
      RECT 78.955 3.23 79.125 3.4 ;
      RECT 78.715 3.79 78.885 3.96 ;
      RECT 78.715 4.35 78.885 4.52 ;
      RECT 78.235 3.79 78.405 3.96 ;
      RECT 77.995 4.91 78.165 5.08 ;
      RECT 77.955 3.23 78.125 3.4 ;
      RECT 77.755 4.07 77.925 4.24 ;
      RECT 77.515 4.91 77.685 5.08 ;
      RECT 77.275 4.35 77.445 4.52 ;
      RECT 76.795 3.79 76.965 3.96 ;
      RECT 76.555 3.23 76.725 3.4 ;
      RECT 76.555 4.91 76.725 5.08 ;
      RECT 76.075 4.35 76.245 4.52 ;
      RECT 75.835 3.79 76.005 3.96 ;
      RECT 75.595 4.63 75.765 4.8 ;
      RECT 75.355 4.07 75.525 4.24 ;
      RECT 74.66 3.23 74.83 3.4 ;
      RECT 74.66 4.63 74.83 4.8 ;
      RECT 73.035 7.31 73.205 7.48 ;
      RECT 73.03 8.61 73.2 8.78 ;
      RECT 73.03 10.09 73.2 10.26 ;
      RECT 72.66 8.24 72.83 8.41 ;
      RECT 72.655 4.055 72.825 4.225 ;
      RECT 72.04 2.205 72.21 2.375 ;
      RECT 72.04 3.685 72.21 3.855 ;
      RECT 72.04 8.61 72.21 8.78 ;
      RECT 72.04 10.09 72.21 10.26 ;
      RECT 71.67 4.055 71.84 4.225 ;
      RECT 71.67 8.24 71.84 8.41 ;
      RECT 70.68 3.315 70.85 3.485 ;
      RECT 70.68 8.98 70.85 9.15 ;
      RECT 70.25 2.205 70.42 2.375 ;
      RECT 70.25 2.945 70.42 3.115 ;
      RECT 70.25 9.35 70.42 9.52 ;
      RECT 70.25 10.09 70.42 10.26 ;
      RECT 69.88 3.685 70.05 3.855 ;
      RECT 69.88 8.61 70.05 8.78 ;
      RECT 66.815 4.07 66.985 4.24 ;
      RECT 66.575 3.23 66.745 3.4 ;
      RECT 66.575 4.91 66.745 5.08 ;
      RECT 66.335 3.79 66.505 3.96 ;
      RECT 66.335 4.35 66.505 4.52 ;
      RECT 65.855 4.07 66.025 4.24 ;
      RECT 65.615 3.23 65.785 3.4 ;
      RECT 65.375 3.79 65.545 3.96 ;
      RECT 65.165 4.63 65.335 4.8 ;
      RECT 65.065 8.98 65.235 9.15 ;
      RECT 64.895 4.07 65.065 4.24 ;
      RECT 64.635 9.35 64.805 9.52 ;
      RECT 64.635 10.09 64.805 10.26 ;
      RECT 64.63 4.91 64.8 5.08 ;
      RECT 64.415 3.49 64.585 3.66 ;
      RECT 63.935 4.07 64.105 4.24 ;
      RECT 63.695 3.23 63.865 3.4 ;
      RECT 63.455 3.79 63.625 3.96 ;
      RECT 63.455 4.35 63.625 4.52 ;
      RECT 62.975 3.79 63.145 3.96 ;
      RECT 62.735 4.91 62.905 5.08 ;
      RECT 62.695 3.23 62.865 3.4 ;
      RECT 62.495 4.07 62.665 4.24 ;
      RECT 62.255 4.91 62.425 5.08 ;
      RECT 62.015 4.35 62.185 4.52 ;
      RECT 61.535 3.79 61.705 3.96 ;
      RECT 61.295 3.23 61.465 3.4 ;
      RECT 61.295 4.91 61.465 5.08 ;
      RECT 60.815 4.35 60.985 4.52 ;
      RECT 60.575 3.79 60.745 3.96 ;
      RECT 60.335 4.63 60.505 4.8 ;
      RECT 60.095 4.07 60.265 4.24 ;
      RECT 59.4 3.23 59.57 3.4 ;
      RECT 59.4 4.63 59.57 4.8 ;
      RECT 57.775 7.31 57.945 7.48 ;
      RECT 57.77 8.61 57.94 8.78 ;
      RECT 57.77 10.09 57.94 10.26 ;
      RECT 57.4 8.24 57.57 8.41 ;
      RECT 57.395 4.055 57.565 4.225 ;
      RECT 56.78 2.205 56.95 2.375 ;
      RECT 56.78 3.685 56.95 3.855 ;
      RECT 56.78 8.61 56.95 8.78 ;
      RECT 56.78 10.09 56.95 10.26 ;
      RECT 56.41 4.055 56.58 4.225 ;
      RECT 56.41 8.24 56.58 8.41 ;
      RECT 55.42 3.315 55.59 3.485 ;
      RECT 55.42 8.98 55.59 9.15 ;
      RECT 54.99 2.205 55.16 2.375 ;
      RECT 54.99 2.945 55.16 3.115 ;
      RECT 54.99 9.35 55.16 9.52 ;
      RECT 54.99 10.09 55.16 10.26 ;
      RECT 54.62 3.685 54.79 3.855 ;
      RECT 54.62 8.61 54.79 8.78 ;
      RECT 51.555 4.07 51.725 4.24 ;
      RECT 51.315 3.23 51.485 3.4 ;
      RECT 51.315 4.91 51.485 5.08 ;
      RECT 51.075 3.79 51.245 3.96 ;
      RECT 51.075 4.35 51.245 4.52 ;
      RECT 50.595 4.07 50.765 4.24 ;
      RECT 50.355 3.23 50.525 3.4 ;
      RECT 50.115 3.79 50.285 3.96 ;
      RECT 49.905 4.63 50.075 4.8 ;
      RECT 49.805 8.98 49.975 9.15 ;
      RECT 49.635 4.07 49.805 4.24 ;
      RECT 49.375 9.35 49.545 9.52 ;
      RECT 49.375 10.09 49.545 10.26 ;
      RECT 49.37 4.91 49.54 5.08 ;
      RECT 49.155 3.49 49.325 3.66 ;
      RECT 48.675 4.07 48.845 4.24 ;
      RECT 48.435 3.23 48.605 3.4 ;
      RECT 48.195 3.79 48.365 3.96 ;
      RECT 48.195 4.35 48.365 4.52 ;
      RECT 47.715 3.79 47.885 3.96 ;
      RECT 47.475 4.91 47.645 5.08 ;
      RECT 47.435 3.23 47.605 3.4 ;
      RECT 47.235 4.07 47.405 4.24 ;
      RECT 46.995 4.91 47.165 5.08 ;
      RECT 46.755 4.35 46.925 4.52 ;
      RECT 46.275 3.79 46.445 3.96 ;
      RECT 46.035 3.23 46.205 3.4 ;
      RECT 46.035 4.91 46.205 5.08 ;
      RECT 45.555 4.35 45.725 4.52 ;
      RECT 45.315 3.79 45.485 3.96 ;
      RECT 45.075 4.63 45.245 4.8 ;
      RECT 44.835 4.07 45.005 4.24 ;
      RECT 44.14 3.23 44.31 3.4 ;
      RECT 44.14 4.63 44.31 4.8 ;
      RECT 42.515 7.31 42.685 7.48 ;
      RECT 42.51 8.61 42.68 8.78 ;
      RECT 42.51 10.09 42.68 10.26 ;
      RECT 42.14 8.24 42.31 8.41 ;
      RECT 42.135 4.055 42.305 4.225 ;
      RECT 41.52 2.205 41.69 2.375 ;
      RECT 41.52 3.685 41.69 3.855 ;
      RECT 41.52 8.61 41.69 8.78 ;
      RECT 41.52 10.09 41.69 10.26 ;
      RECT 41.15 4.055 41.32 4.225 ;
      RECT 41.15 8.24 41.32 8.41 ;
      RECT 40.16 3.315 40.33 3.485 ;
      RECT 40.16 8.98 40.33 9.15 ;
      RECT 39.73 2.205 39.9 2.375 ;
      RECT 39.73 2.945 39.9 3.115 ;
      RECT 39.73 9.35 39.9 9.52 ;
      RECT 39.73 10.09 39.9 10.26 ;
      RECT 39.36 3.685 39.53 3.855 ;
      RECT 39.36 8.61 39.53 8.78 ;
      RECT 36.295 4.07 36.465 4.24 ;
      RECT 36.055 3.23 36.225 3.4 ;
      RECT 36.055 4.91 36.225 5.08 ;
      RECT 35.815 3.79 35.985 3.96 ;
      RECT 35.815 4.35 35.985 4.52 ;
      RECT 35.335 4.07 35.505 4.24 ;
      RECT 35.095 3.23 35.265 3.4 ;
      RECT 34.855 3.79 35.025 3.96 ;
      RECT 34.645 4.63 34.815 4.8 ;
      RECT 34.545 8.98 34.715 9.15 ;
      RECT 34.375 4.07 34.545 4.24 ;
      RECT 34.115 9.35 34.285 9.52 ;
      RECT 34.115 10.09 34.285 10.26 ;
      RECT 34.11 4.91 34.28 5.08 ;
      RECT 33.895 3.49 34.065 3.66 ;
      RECT 33.415 4.07 33.585 4.24 ;
      RECT 33.175 3.23 33.345 3.4 ;
      RECT 32.935 3.79 33.105 3.96 ;
      RECT 32.935 4.35 33.105 4.52 ;
      RECT 32.455 3.79 32.625 3.96 ;
      RECT 32.215 4.91 32.385 5.08 ;
      RECT 32.175 3.23 32.345 3.4 ;
      RECT 31.975 4.07 32.145 4.24 ;
      RECT 31.735 4.91 31.905 5.08 ;
      RECT 31.495 4.35 31.665 4.52 ;
      RECT 31.015 3.79 31.185 3.96 ;
      RECT 30.775 3.23 30.945 3.4 ;
      RECT 30.775 4.91 30.945 5.08 ;
      RECT 30.295 4.35 30.465 4.52 ;
      RECT 30.055 3.79 30.225 3.96 ;
      RECT 29.815 4.63 29.985 4.8 ;
      RECT 29.575 4.07 29.745 4.24 ;
      RECT 28.88 3.23 29.05 3.4 ;
      RECT 28.88 4.63 29.05 4.8 ;
      RECT 26.6 9.35 26.77 9.52 ;
      RECT 26.6 10.09 26.77 10.26 ;
      RECT 26.23 8.61 26.4 8.78 ;
    LAYER li1 ;
      RECT 103.55 7.31 103.72 8.78 ;
      RECT 103.55 7.31 103.725 8.57 ;
      RECT 103.18 9.26 103.65 9.43 ;
      RECT 103.18 8.24 103.35 9.43 ;
      RECT 103.175 3.035 103.345 4.225 ;
      RECT 103.175 3.035 103.645 3.205 ;
      RECT 102.56 3.895 102.735 5.155 ;
      RECT 102.56 3.685 102.73 5.155 ;
      RECT 102.56 7.31 102.73 8.78 ;
      RECT 102.56 7.31 102.735 8.57 ;
      RECT 102.19 3.035 102.36 4.225 ;
      RECT 102.19 3.035 102.66 3.205 ;
      RECT 102.19 9.26 102.66 9.43 ;
      RECT 102.19 8.24 102.36 9.43 ;
      RECT 101.2 4.015 101.375 5.155 ;
      RECT 101.2 1.865 101.37 5.155 ;
      RECT 101.2 1.865 101.375 2.415 ;
      RECT 101.2 10.05 101.375 10.6 ;
      RECT 101.2 7.31 101.37 10.6 ;
      RECT 101.2 7.31 101.375 8.45 ;
      RECT 100.77 3.895 100.945 5.155 ;
      RECT 100.77 2.945 100.94 5.155 ;
      RECT 100.77 7.31 100.94 9.52 ;
      RECT 100.77 7.31 100.945 8.57 ;
      RECT 100.34 3.925 100.51 5.155 ;
      RECT 100.4 2.145 100.57 4.095 ;
      RECT 100.34 1.865 100.51 2.315 ;
      RECT 100.34 10.15 100.51 10.6 ;
      RECT 100.4 8.37 100.57 10.32 ;
      RECT 100.34 7.31 100.51 8.54 ;
      RECT 99.815 3.895 99.99 5.155 ;
      RECT 99.815 1.865 99.985 5.155 ;
      RECT 99.815 3.365 100.225 3.695 ;
      RECT 99.815 2.525 100.225 2.855 ;
      RECT 99.815 1.865 99.99 2.355 ;
      RECT 99.815 10.11 99.99 10.6 ;
      RECT 99.815 7.31 99.985 10.6 ;
      RECT 99.815 9.61 100.225 9.94 ;
      RECT 99.815 8.77 100.225 9.1 ;
      RECT 99.815 7.31 99.99 8.57 ;
      RECT 97.095 4.91 97.61 5.08 ;
      RECT 97.44 4.52 97.61 5.08 ;
      RECT 97.545 4.44 97.72 4.77 ;
      RECT 97.335 3.83 97.61 4.24 ;
      RECT 97.215 3.83 97.61 4.04 ;
      RECT 95.68 4.44 95.855 4.8 ;
      RECT 95.68 4.52 97.025 4.69 ;
      RECT 96.855 4.35 97.025 4.69 ;
      RECT 95.585 10.05 95.76 10.6 ;
      RECT 95.585 7.31 95.755 10.6 ;
      RECT 95.585 7.31 95.76 8.45 ;
      RECT 95.415 3.87 95.585 4.24 ;
      RECT 94.935 3.87 95.585 4.14 ;
      RECT 94.855 3.87 95.665 4.04 ;
      RECT 94.215 3.11 94.385 3.4 ;
      RECT 94.215 3.11 95.455 3.28 ;
      RECT 95.155 7.31 95.325 9.52 ;
      RECT 95.155 7.31 95.33 8.57 ;
      RECT 94.935 3.45 95.105 3.66 ;
      RECT 94.575 3.45 95.105 3.62 ;
      RECT 94.2 10.11 94.375 10.6 ;
      RECT 94.2 7.31 94.37 10.6 ;
      RECT 94.2 9.61 94.61 9.94 ;
      RECT 94.2 8.77 94.61 9.1 ;
      RECT 94.2 7.31 94.375 8.57 ;
      RECT 93.975 4.52 94.465 4.69 ;
      RECT 93.975 4.35 94.145 4.69 ;
      RECT 93.255 4.52 93.425 5.08 ;
      RECT 93.15 4.52 93.48 4.69 ;
      RECT 93.215 3.13 93.385 3.4 ;
      RECT 93.255 3.05 93.425 3.38 ;
      RECT 93.12 3.13 93.425 3.35 ;
      RECT 91.695 4.52 91.985 5.08 ;
      RECT 91.815 4.44 91.985 5.08 ;
      RECT 88.29 7.31 88.46 8.78 ;
      RECT 88.29 7.31 88.465 8.57 ;
      RECT 87.92 9.26 88.39 9.43 ;
      RECT 87.92 8.24 88.09 9.43 ;
      RECT 87.915 3.035 88.085 4.225 ;
      RECT 87.915 3.035 88.385 3.205 ;
      RECT 87.3 3.895 87.475 5.155 ;
      RECT 87.3 3.685 87.47 5.155 ;
      RECT 87.3 7.31 87.47 8.78 ;
      RECT 87.3 7.31 87.475 8.57 ;
      RECT 86.93 3.035 87.1 4.225 ;
      RECT 86.93 3.035 87.4 3.205 ;
      RECT 86.93 9.26 87.4 9.43 ;
      RECT 86.93 8.24 87.1 9.43 ;
      RECT 85.94 4.015 86.115 5.155 ;
      RECT 85.94 1.865 86.11 5.155 ;
      RECT 85.94 1.865 86.115 2.415 ;
      RECT 85.94 10.05 86.115 10.6 ;
      RECT 85.94 7.31 86.11 10.6 ;
      RECT 85.94 7.31 86.115 8.45 ;
      RECT 85.51 3.895 85.685 5.155 ;
      RECT 85.51 2.945 85.68 5.155 ;
      RECT 85.51 7.31 85.68 9.52 ;
      RECT 85.51 7.31 85.685 8.57 ;
      RECT 85.08 3.925 85.25 5.155 ;
      RECT 85.14 2.145 85.31 4.095 ;
      RECT 85.08 1.865 85.25 2.315 ;
      RECT 85.08 10.15 85.25 10.6 ;
      RECT 85.14 8.37 85.31 10.32 ;
      RECT 85.08 7.31 85.25 8.54 ;
      RECT 84.555 3.895 84.73 5.155 ;
      RECT 84.555 1.865 84.725 5.155 ;
      RECT 84.555 3.365 84.965 3.695 ;
      RECT 84.555 2.525 84.965 2.855 ;
      RECT 84.555 1.865 84.73 2.355 ;
      RECT 84.555 10.11 84.73 10.6 ;
      RECT 84.555 7.31 84.725 10.6 ;
      RECT 84.555 9.61 84.965 9.94 ;
      RECT 84.555 8.77 84.965 9.1 ;
      RECT 84.555 7.31 84.73 8.57 ;
      RECT 81.835 4.91 82.35 5.08 ;
      RECT 82.18 4.52 82.35 5.08 ;
      RECT 82.285 4.44 82.46 4.77 ;
      RECT 82.075 3.83 82.35 4.24 ;
      RECT 81.955 3.83 82.35 4.04 ;
      RECT 80.42 4.44 80.595 4.8 ;
      RECT 80.42 4.52 81.765 4.69 ;
      RECT 81.595 4.35 81.765 4.69 ;
      RECT 80.325 10.05 80.5 10.6 ;
      RECT 80.325 7.31 80.495 10.6 ;
      RECT 80.325 7.31 80.5 8.45 ;
      RECT 80.155 3.87 80.325 4.24 ;
      RECT 79.675 3.87 80.325 4.14 ;
      RECT 79.595 3.87 80.405 4.04 ;
      RECT 78.955 3.11 79.125 3.4 ;
      RECT 78.955 3.11 80.195 3.28 ;
      RECT 79.895 7.31 80.065 9.52 ;
      RECT 79.895 7.31 80.07 8.57 ;
      RECT 79.675 3.45 79.845 3.66 ;
      RECT 79.315 3.45 79.845 3.62 ;
      RECT 78.94 10.11 79.115 10.6 ;
      RECT 78.94 7.31 79.11 10.6 ;
      RECT 78.94 9.61 79.35 9.94 ;
      RECT 78.94 8.77 79.35 9.1 ;
      RECT 78.94 7.31 79.115 8.57 ;
      RECT 78.715 4.52 79.205 4.69 ;
      RECT 78.715 4.35 78.885 4.69 ;
      RECT 77.995 4.52 78.165 5.08 ;
      RECT 77.89 4.52 78.22 4.69 ;
      RECT 77.955 3.13 78.125 3.4 ;
      RECT 77.995 3.05 78.165 3.38 ;
      RECT 77.86 3.13 78.165 3.35 ;
      RECT 76.435 4.52 76.725 5.08 ;
      RECT 76.555 4.44 76.725 5.08 ;
      RECT 73.03 7.31 73.2 8.78 ;
      RECT 73.03 7.31 73.205 8.57 ;
      RECT 72.66 9.26 73.13 9.43 ;
      RECT 72.66 8.24 72.83 9.43 ;
      RECT 72.655 3.035 72.825 4.225 ;
      RECT 72.655 3.035 73.125 3.205 ;
      RECT 72.04 3.895 72.215 5.155 ;
      RECT 72.04 3.685 72.21 5.155 ;
      RECT 72.04 7.31 72.21 8.78 ;
      RECT 72.04 7.31 72.215 8.57 ;
      RECT 71.67 3.035 71.84 4.225 ;
      RECT 71.67 3.035 72.14 3.205 ;
      RECT 71.67 9.26 72.14 9.43 ;
      RECT 71.67 8.24 71.84 9.43 ;
      RECT 70.68 4.015 70.855 5.155 ;
      RECT 70.68 1.865 70.85 5.155 ;
      RECT 70.68 1.865 70.855 2.415 ;
      RECT 70.68 10.05 70.855 10.6 ;
      RECT 70.68 7.31 70.85 10.6 ;
      RECT 70.68 7.31 70.855 8.45 ;
      RECT 70.25 3.895 70.425 5.155 ;
      RECT 70.25 2.945 70.42 5.155 ;
      RECT 70.25 7.31 70.42 9.52 ;
      RECT 70.25 7.31 70.425 8.57 ;
      RECT 69.82 3.925 69.99 5.155 ;
      RECT 69.88 2.145 70.05 4.095 ;
      RECT 69.82 1.865 69.99 2.315 ;
      RECT 69.82 10.15 69.99 10.6 ;
      RECT 69.88 8.37 70.05 10.32 ;
      RECT 69.82 7.31 69.99 8.54 ;
      RECT 69.295 3.895 69.47 5.155 ;
      RECT 69.295 1.865 69.465 5.155 ;
      RECT 69.295 3.365 69.705 3.695 ;
      RECT 69.295 2.525 69.705 2.855 ;
      RECT 69.295 1.865 69.47 2.355 ;
      RECT 69.295 10.11 69.47 10.6 ;
      RECT 69.295 7.31 69.465 10.6 ;
      RECT 69.295 9.61 69.705 9.94 ;
      RECT 69.295 8.77 69.705 9.1 ;
      RECT 69.295 7.31 69.47 8.57 ;
      RECT 66.575 4.91 67.09 5.08 ;
      RECT 66.92 4.52 67.09 5.08 ;
      RECT 67.025 4.44 67.2 4.77 ;
      RECT 66.815 3.83 67.09 4.24 ;
      RECT 66.695 3.83 67.09 4.04 ;
      RECT 65.16 4.44 65.335 4.8 ;
      RECT 65.16 4.52 66.505 4.69 ;
      RECT 66.335 4.35 66.505 4.69 ;
      RECT 65.065 10.05 65.24 10.6 ;
      RECT 65.065 7.31 65.235 10.6 ;
      RECT 65.065 7.31 65.24 8.45 ;
      RECT 64.895 3.87 65.065 4.24 ;
      RECT 64.415 3.87 65.065 4.14 ;
      RECT 64.335 3.87 65.145 4.04 ;
      RECT 63.695 3.11 63.865 3.4 ;
      RECT 63.695 3.11 64.935 3.28 ;
      RECT 64.635 7.31 64.805 9.52 ;
      RECT 64.635 7.31 64.81 8.57 ;
      RECT 64.415 3.45 64.585 3.66 ;
      RECT 64.055 3.45 64.585 3.62 ;
      RECT 63.68 10.11 63.855 10.6 ;
      RECT 63.68 7.31 63.85 10.6 ;
      RECT 63.68 9.61 64.09 9.94 ;
      RECT 63.68 8.77 64.09 9.1 ;
      RECT 63.68 7.31 63.855 8.57 ;
      RECT 63.455 4.52 63.945 4.69 ;
      RECT 63.455 4.35 63.625 4.69 ;
      RECT 62.735 4.52 62.905 5.08 ;
      RECT 62.63 4.52 62.96 4.69 ;
      RECT 62.695 3.13 62.865 3.4 ;
      RECT 62.735 3.05 62.905 3.38 ;
      RECT 62.6 3.13 62.905 3.35 ;
      RECT 61.175 4.52 61.465 5.08 ;
      RECT 61.295 4.44 61.465 5.08 ;
      RECT 57.77 7.31 57.94 8.78 ;
      RECT 57.77 7.31 57.945 8.57 ;
      RECT 57.4 9.26 57.87 9.43 ;
      RECT 57.4 8.24 57.57 9.43 ;
      RECT 57.395 3.035 57.565 4.225 ;
      RECT 57.395 3.035 57.865 3.205 ;
      RECT 56.78 3.895 56.955 5.155 ;
      RECT 56.78 3.685 56.95 5.155 ;
      RECT 56.78 7.31 56.95 8.78 ;
      RECT 56.78 7.31 56.955 8.57 ;
      RECT 56.41 3.035 56.58 4.225 ;
      RECT 56.41 3.035 56.88 3.205 ;
      RECT 56.41 9.26 56.88 9.43 ;
      RECT 56.41 8.24 56.58 9.43 ;
      RECT 55.42 4.015 55.595 5.155 ;
      RECT 55.42 1.865 55.59 5.155 ;
      RECT 55.42 1.865 55.595 2.415 ;
      RECT 55.42 10.05 55.595 10.6 ;
      RECT 55.42 7.31 55.59 10.6 ;
      RECT 55.42 7.31 55.595 8.45 ;
      RECT 54.99 3.895 55.165 5.155 ;
      RECT 54.99 2.945 55.16 5.155 ;
      RECT 54.99 7.31 55.16 9.52 ;
      RECT 54.99 7.31 55.165 8.57 ;
      RECT 54.56 3.925 54.73 5.155 ;
      RECT 54.62 2.145 54.79 4.095 ;
      RECT 54.56 1.865 54.73 2.315 ;
      RECT 54.56 10.15 54.73 10.6 ;
      RECT 54.62 8.37 54.79 10.32 ;
      RECT 54.56 7.31 54.73 8.54 ;
      RECT 54.035 3.895 54.21 5.155 ;
      RECT 54.035 1.865 54.205 5.155 ;
      RECT 54.035 3.365 54.445 3.695 ;
      RECT 54.035 2.525 54.445 2.855 ;
      RECT 54.035 1.865 54.21 2.355 ;
      RECT 54.035 10.11 54.21 10.6 ;
      RECT 54.035 7.31 54.205 10.6 ;
      RECT 54.035 9.61 54.445 9.94 ;
      RECT 54.035 8.77 54.445 9.1 ;
      RECT 54.035 7.31 54.21 8.57 ;
      RECT 51.315 4.91 51.83 5.08 ;
      RECT 51.66 4.52 51.83 5.08 ;
      RECT 51.765 4.44 51.94 4.77 ;
      RECT 51.555 3.83 51.83 4.24 ;
      RECT 51.435 3.83 51.83 4.04 ;
      RECT 49.9 4.44 50.075 4.8 ;
      RECT 49.9 4.52 51.245 4.69 ;
      RECT 51.075 4.35 51.245 4.69 ;
      RECT 49.805 10.05 49.98 10.6 ;
      RECT 49.805 7.31 49.975 10.6 ;
      RECT 49.805 7.31 49.98 8.45 ;
      RECT 49.635 3.87 49.805 4.24 ;
      RECT 49.155 3.87 49.805 4.14 ;
      RECT 49.075 3.87 49.885 4.04 ;
      RECT 48.435 3.11 48.605 3.4 ;
      RECT 48.435 3.11 49.675 3.28 ;
      RECT 49.375 7.31 49.545 9.52 ;
      RECT 49.375 7.31 49.55 8.57 ;
      RECT 49.155 3.45 49.325 3.66 ;
      RECT 48.795 3.45 49.325 3.62 ;
      RECT 48.42 10.11 48.595 10.6 ;
      RECT 48.42 7.31 48.59 10.6 ;
      RECT 48.42 9.61 48.83 9.94 ;
      RECT 48.42 8.77 48.83 9.1 ;
      RECT 48.42 7.31 48.595 8.57 ;
      RECT 48.195 4.52 48.685 4.69 ;
      RECT 48.195 4.35 48.365 4.69 ;
      RECT 47.475 4.52 47.645 5.08 ;
      RECT 47.37 4.52 47.7 4.69 ;
      RECT 47.435 3.13 47.605 3.4 ;
      RECT 47.475 3.05 47.645 3.38 ;
      RECT 47.34 3.13 47.645 3.35 ;
      RECT 45.915 4.52 46.205 5.08 ;
      RECT 46.035 4.44 46.205 5.08 ;
      RECT 42.51 7.31 42.68 8.78 ;
      RECT 42.51 7.31 42.685 8.57 ;
      RECT 42.14 9.26 42.61 9.43 ;
      RECT 42.14 8.24 42.31 9.43 ;
      RECT 42.135 3.035 42.305 4.225 ;
      RECT 42.135 3.035 42.605 3.205 ;
      RECT 41.52 3.895 41.695 5.155 ;
      RECT 41.52 3.685 41.69 5.155 ;
      RECT 41.52 7.31 41.69 8.78 ;
      RECT 41.52 7.31 41.695 8.57 ;
      RECT 41.15 3.035 41.32 4.225 ;
      RECT 41.15 3.035 41.62 3.205 ;
      RECT 41.15 9.26 41.62 9.43 ;
      RECT 41.15 8.24 41.32 9.43 ;
      RECT 40.16 4.015 40.335 5.155 ;
      RECT 40.16 1.865 40.33 5.155 ;
      RECT 40.16 1.865 40.335 2.415 ;
      RECT 40.16 10.05 40.335 10.6 ;
      RECT 40.16 7.31 40.33 10.6 ;
      RECT 40.16 7.31 40.335 8.45 ;
      RECT 39.73 3.895 39.905 5.155 ;
      RECT 39.73 2.945 39.9 5.155 ;
      RECT 39.73 7.31 39.9 9.52 ;
      RECT 39.73 7.31 39.905 8.57 ;
      RECT 39.3 3.925 39.47 5.155 ;
      RECT 39.36 2.145 39.53 4.095 ;
      RECT 39.3 1.865 39.47 2.315 ;
      RECT 39.3 10.15 39.47 10.6 ;
      RECT 39.36 8.37 39.53 10.32 ;
      RECT 39.3 7.31 39.47 8.54 ;
      RECT 38.775 3.895 38.95 5.155 ;
      RECT 38.775 1.865 38.945 5.155 ;
      RECT 38.775 3.365 39.185 3.695 ;
      RECT 38.775 2.525 39.185 2.855 ;
      RECT 38.775 1.865 38.95 2.355 ;
      RECT 38.775 10.11 38.95 10.6 ;
      RECT 38.775 7.31 38.945 10.6 ;
      RECT 38.775 9.61 39.185 9.94 ;
      RECT 38.775 8.77 39.185 9.1 ;
      RECT 38.775 7.31 38.95 8.57 ;
      RECT 36.055 4.91 36.57 5.08 ;
      RECT 36.4 4.52 36.57 5.08 ;
      RECT 36.505 4.44 36.68 4.77 ;
      RECT 36.295 3.83 36.57 4.24 ;
      RECT 36.175 3.83 36.57 4.04 ;
      RECT 34.64 4.44 34.815 4.8 ;
      RECT 34.64 4.52 35.985 4.69 ;
      RECT 35.815 4.35 35.985 4.69 ;
      RECT 34.545 10.05 34.72 10.6 ;
      RECT 34.545 7.31 34.715 10.6 ;
      RECT 34.545 7.31 34.72 8.45 ;
      RECT 34.375 3.87 34.545 4.24 ;
      RECT 33.895 3.87 34.545 4.14 ;
      RECT 33.815 3.87 34.625 4.04 ;
      RECT 33.175 3.11 33.345 3.4 ;
      RECT 33.175 3.11 34.415 3.28 ;
      RECT 34.115 7.31 34.285 9.52 ;
      RECT 34.115 7.31 34.29 8.57 ;
      RECT 33.895 3.45 34.065 3.66 ;
      RECT 33.535 3.45 34.065 3.62 ;
      RECT 33.16 10.11 33.335 10.6 ;
      RECT 33.16 7.31 33.33 10.6 ;
      RECT 33.16 9.61 33.57 9.94 ;
      RECT 33.16 8.77 33.57 9.1 ;
      RECT 33.16 7.31 33.335 8.57 ;
      RECT 32.935 4.52 33.425 4.69 ;
      RECT 32.935 4.35 33.105 4.69 ;
      RECT 32.215 4.52 32.385 5.08 ;
      RECT 32.11 4.52 32.44 4.69 ;
      RECT 32.175 3.13 32.345 3.4 ;
      RECT 32.215 3.05 32.385 3.38 ;
      RECT 32.08 3.13 32.385 3.35 ;
      RECT 30.655 4.52 30.945 5.08 ;
      RECT 30.775 4.44 30.945 5.08 ;
      RECT 26.6 7.31 26.77 9.52 ;
      RECT 26.6 7.31 26.775 8.57 ;
      RECT 26.17 10.15 26.34 10.6 ;
      RECT 26.23 8.37 26.4 10.32 ;
      RECT 26.17 7.31 26.34 8.54 ;
      RECT 25.645 10.11 25.82 10.6 ;
      RECT 25.645 7.31 25.815 10.6 ;
      RECT 25.645 9.61 26.055 9.94 ;
      RECT 25.645 8.77 26.055 9.1 ;
      RECT 25.645 7.31 25.82 8.57 ;
      RECT 103.55 10.09 103.725 10.6 ;
      RECT 102.56 1.865 102.735 2.375 ;
      RECT 102.56 10.09 102.735 10.6 ;
      RECT 100.77 1.865 100.945 2.375 ;
      RECT 100.77 10.09 100.945 10.6 ;
      RECT 97.095 3.05 97.265 3.4 ;
      RECT 96.855 3.79 97.025 4.12 ;
      RECT 96.375 3.79 96.545 4.24 ;
      RECT 96.135 3.05 96.305 3.4 ;
      RECT 95.895 3.79 96.065 4.12 ;
      RECT 95.155 10.09 95.33 10.6 ;
      RECT 95.15 4.78 95.32 5.11 ;
      RECT 94.455 3.79 94.625 4.24 ;
      RECT 93.975 3.79 94.145 4.12 ;
      RECT 93.495 3.79 93.665 4.12 ;
      RECT 93.015 3.79 93.185 4.24 ;
      RECT 92.775 4.78 92.945 5.11 ;
      RECT 92.535 3.79 92.705 4.52 ;
      RECT 92.055 3.79 92.225 4.12 ;
      RECT 91.815 3.05 91.985 3.4 ;
      RECT 91.335 4.35 91.505 4.77 ;
      RECT 91.095 3.79 91.265 4.12 ;
      RECT 90.855 4.44 91.025 4.8 ;
      RECT 90.615 3.79 90.785 4.24 ;
      RECT 89.92 3.05 90.09 3.4 ;
      RECT 89.92 4.44 90.09 4.8 ;
      RECT 88.29 10.09 88.465 10.6 ;
      RECT 87.3 1.865 87.475 2.375 ;
      RECT 87.3 10.09 87.475 10.6 ;
      RECT 85.51 1.865 85.685 2.375 ;
      RECT 85.51 10.09 85.685 10.6 ;
      RECT 81.835 3.05 82.005 3.4 ;
      RECT 81.595 3.79 81.765 4.12 ;
      RECT 81.115 3.79 81.285 4.24 ;
      RECT 80.875 3.05 81.045 3.4 ;
      RECT 80.635 3.79 80.805 4.12 ;
      RECT 79.895 10.09 80.07 10.6 ;
      RECT 79.89 4.78 80.06 5.11 ;
      RECT 79.195 3.79 79.365 4.24 ;
      RECT 78.715 3.79 78.885 4.12 ;
      RECT 78.235 3.79 78.405 4.12 ;
      RECT 77.755 3.79 77.925 4.24 ;
      RECT 77.515 4.78 77.685 5.11 ;
      RECT 77.275 3.79 77.445 4.52 ;
      RECT 76.795 3.79 76.965 4.12 ;
      RECT 76.555 3.05 76.725 3.4 ;
      RECT 76.075 4.35 76.245 4.77 ;
      RECT 75.835 3.79 76.005 4.12 ;
      RECT 75.595 4.44 75.765 4.8 ;
      RECT 75.355 3.79 75.525 4.24 ;
      RECT 74.66 3.05 74.83 3.4 ;
      RECT 74.66 4.44 74.83 4.8 ;
      RECT 73.03 10.09 73.205 10.6 ;
      RECT 72.04 1.865 72.215 2.375 ;
      RECT 72.04 10.09 72.215 10.6 ;
      RECT 70.25 1.865 70.425 2.375 ;
      RECT 70.25 10.09 70.425 10.6 ;
      RECT 66.575 3.05 66.745 3.4 ;
      RECT 66.335 3.79 66.505 4.12 ;
      RECT 65.855 3.79 66.025 4.24 ;
      RECT 65.615 3.05 65.785 3.4 ;
      RECT 65.375 3.79 65.545 4.12 ;
      RECT 64.635 10.09 64.81 10.6 ;
      RECT 64.63 4.78 64.8 5.11 ;
      RECT 63.935 3.79 64.105 4.24 ;
      RECT 63.455 3.79 63.625 4.12 ;
      RECT 62.975 3.79 63.145 4.12 ;
      RECT 62.495 3.79 62.665 4.24 ;
      RECT 62.255 4.78 62.425 5.11 ;
      RECT 62.015 3.79 62.185 4.52 ;
      RECT 61.535 3.79 61.705 4.12 ;
      RECT 61.295 3.05 61.465 3.4 ;
      RECT 60.815 4.35 60.985 4.77 ;
      RECT 60.575 3.79 60.745 4.12 ;
      RECT 60.335 4.44 60.505 4.8 ;
      RECT 60.095 3.79 60.265 4.24 ;
      RECT 59.4 3.05 59.57 3.4 ;
      RECT 59.4 4.44 59.57 4.8 ;
      RECT 57.77 10.09 57.945 10.6 ;
      RECT 56.78 1.865 56.955 2.375 ;
      RECT 56.78 10.09 56.955 10.6 ;
      RECT 54.99 1.865 55.165 2.375 ;
      RECT 54.99 10.09 55.165 10.6 ;
      RECT 51.315 3.05 51.485 3.4 ;
      RECT 51.075 3.79 51.245 4.12 ;
      RECT 50.595 3.79 50.765 4.24 ;
      RECT 50.355 3.05 50.525 3.4 ;
      RECT 50.115 3.79 50.285 4.12 ;
      RECT 49.375 10.09 49.55 10.6 ;
      RECT 49.37 4.78 49.54 5.11 ;
      RECT 48.675 3.79 48.845 4.24 ;
      RECT 48.195 3.79 48.365 4.12 ;
      RECT 47.715 3.79 47.885 4.12 ;
      RECT 47.235 3.79 47.405 4.24 ;
      RECT 46.995 4.78 47.165 5.11 ;
      RECT 46.755 3.79 46.925 4.52 ;
      RECT 46.275 3.79 46.445 4.12 ;
      RECT 46.035 3.05 46.205 3.4 ;
      RECT 45.555 4.35 45.725 4.77 ;
      RECT 45.315 3.79 45.485 4.12 ;
      RECT 45.075 4.44 45.245 4.8 ;
      RECT 44.835 3.79 45.005 4.24 ;
      RECT 44.14 3.05 44.31 3.4 ;
      RECT 44.14 4.44 44.31 4.8 ;
      RECT 42.51 10.09 42.685 10.6 ;
      RECT 41.52 1.865 41.695 2.375 ;
      RECT 41.52 10.09 41.695 10.6 ;
      RECT 39.73 1.865 39.905 2.375 ;
      RECT 39.73 10.09 39.905 10.6 ;
      RECT 36.055 3.05 36.225 3.4 ;
      RECT 35.815 3.79 35.985 4.12 ;
      RECT 35.335 3.79 35.505 4.24 ;
      RECT 35.095 3.05 35.265 3.4 ;
      RECT 34.855 3.79 35.025 4.12 ;
      RECT 34.115 10.09 34.29 10.6 ;
      RECT 34.11 4.78 34.28 5.11 ;
      RECT 33.415 3.79 33.585 4.24 ;
      RECT 32.935 3.79 33.105 4.12 ;
      RECT 32.455 3.79 32.625 4.12 ;
      RECT 31.975 3.79 32.145 4.24 ;
      RECT 31.735 4.78 31.905 5.11 ;
      RECT 31.495 3.79 31.665 4.52 ;
      RECT 31.015 3.79 31.185 4.12 ;
      RECT 30.775 3.05 30.945 3.4 ;
      RECT 30.295 4.35 30.465 4.77 ;
      RECT 30.055 3.79 30.225 4.12 ;
      RECT 29.815 4.44 29.985 4.8 ;
      RECT 29.575 3.79 29.745 4.24 ;
      RECT 28.88 3.05 29.05 3.4 ;
      RECT 28.88 4.44 29.05 4.8 ;
      RECT 26.6 10.09 26.775 10.6 ;
  END
END sky130_osu_ring_oscillator_mpr2xa_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2ya_8_b0r1
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ya_8_b0r1 ;
  SIZE 94.1 BY 12.465 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 32.405 0 32.785 5.265 ;
      LAYER met2 ;
        RECT 32.405 4.885 32.785 5.265 ;
      LAYER li1 ;
        RECT 32.51 1.865 32.685 2.375 ;
        RECT 32.51 3.895 32.685 5.155 ;
        RECT 32.51 3.685 32.68 5.155 ;
      LAYER met1 ;
        RECT 32.42 4.93 32.77 5.22 ;
        RECT 32.45 2.175 32.745 2.405 ;
        RECT 32.45 3.655 32.74 3.885 ;
        RECT 32.51 2.175 32.68 3.885 ;
      LAYER via1 ;
        RECT 32.52 5 32.67 5.15 ;
      LAYER via2 ;
        RECT 32.495 4.975 32.695 5.175 ;
      LAYER mcon ;
        RECT 32.51 3.685 32.68 3.855 ;
        RECT 32.515 4.985 32.685 5.155 ;
        RECT 32.51 2.205 32.685 2.375 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 47.665 0 48.045 5.265 ;
      LAYER met2 ;
        RECT 47.665 4.885 48.045 5.265 ;
      LAYER li1 ;
        RECT 47.77 1.865 47.945 2.375 ;
        RECT 47.77 3.895 47.945 5.155 ;
        RECT 47.77 3.685 47.94 5.155 ;
      LAYER met1 ;
        RECT 47.68 4.93 48.03 5.22 ;
        RECT 47.71 2.175 48.005 2.405 ;
        RECT 47.71 3.655 48 3.885 ;
        RECT 47.77 2.175 47.94 3.885 ;
      LAYER via1 ;
        RECT 47.78 5 47.93 5.15 ;
      LAYER via2 ;
        RECT 47.755 4.975 47.955 5.175 ;
      LAYER mcon ;
        RECT 47.77 3.685 47.94 3.855 ;
        RECT 47.775 4.985 47.945 5.155 ;
        RECT 47.77 2.205 47.945 2.375 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 62.925 0 63.305 5.265 ;
      LAYER met2 ;
        RECT 62.925 4.885 63.305 5.265 ;
      LAYER li1 ;
        RECT 63.03 1.865 63.205 2.375 ;
        RECT 63.03 3.895 63.205 5.155 ;
        RECT 63.03 3.685 63.2 5.155 ;
      LAYER met1 ;
        RECT 62.94 4.93 63.29 5.22 ;
        RECT 62.97 2.175 63.265 2.405 ;
        RECT 62.97 3.655 63.26 3.885 ;
        RECT 63.03 2.175 63.2 3.885 ;
      LAYER via1 ;
        RECT 63.04 5 63.19 5.15 ;
      LAYER via2 ;
        RECT 63.015 4.975 63.215 5.175 ;
      LAYER mcon ;
        RECT 63.03 3.685 63.2 3.855 ;
        RECT 63.035 4.985 63.205 5.155 ;
        RECT 63.03 2.205 63.205 2.375 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 78.185 0 78.565 5.265 ;
      LAYER met2 ;
        RECT 78.185 4.885 78.565 5.265 ;
      LAYER li1 ;
        RECT 78.29 1.865 78.465 2.375 ;
        RECT 78.29 3.895 78.465 5.155 ;
        RECT 78.29 3.685 78.46 5.155 ;
      LAYER met1 ;
        RECT 78.2 4.93 78.55 5.22 ;
        RECT 78.23 2.175 78.525 2.405 ;
        RECT 78.23 3.655 78.52 3.885 ;
        RECT 78.29 2.175 78.46 3.885 ;
      LAYER via1 ;
        RECT 78.3 5 78.45 5.15 ;
      LAYER via2 ;
        RECT 78.275 4.975 78.475 5.175 ;
      LAYER mcon ;
        RECT 78.29 3.685 78.46 3.855 ;
        RECT 78.295 4.985 78.465 5.155 ;
        RECT 78.29 2.205 78.465 2.375 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 93.445 0 93.825 5.265 ;
      LAYER met2 ;
        RECT 93.445 4.885 93.825 5.265 ;
      LAYER li1 ;
        RECT 93.55 1.865 93.725 2.375 ;
        RECT 93.55 3.895 93.725 5.155 ;
        RECT 93.55 3.685 93.72 5.155 ;
      LAYER met1 ;
        RECT 93.46 4.93 93.81 5.22 ;
        RECT 93.49 2.175 93.785 2.405 ;
        RECT 93.49 3.655 93.78 3.885 ;
        RECT 93.55 2.175 93.72 3.885 ;
      LAYER via1 ;
        RECT 93.56 5 93.71 5.15 ;
      LAYER via2 ;
        RECT 93.535 4.975 93.735 5.175 ;
      LAYER mcon ;
        RECT 93.55 3.685 93.72 3.855 ;
        RECT 93.555 4.985 93.725 5.155 ;
        RECT 93.55 2.205 93.725 2.375 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 28.285 4 28.625 4.35 ;
        RECT 28.28 8.15 28.62 8.5 ;
        RECT 28.36 4 28.535 8.5 ;
      LAYER li1 ;
        RECT 28.36 2.955 28.53 4.225 ;
        RECT 28.36 8.24 28.53 9.51 ;
        RECT 22.725 8.24 22.895 9.51 ;
      LAYER met1 ;
        RECT 28.285 4.055 28.76 4.225 ;
        RECT 28.285 4 28.625 4.35 ;
        RECT 28.28 8.24 28.76 8.41 ;
        RECT 28.28 8.15 28.62 8.5 ;
        RECT 22.665 8.235 28.62 8.405 ;
        RECT 22.665 8.235 23.125 8.41 ;
        RECT 22.665 8.21 22.955 8.44 ;
      LAYER via1 ;
        RECT 28.38 8.25 28.53 8.4 ;
        RECT 28.385 4.1 28.535 4.25 ;
      LAYER mcon ;
        RECT 22.725 8.24 22.895 8.41 ;
        RECT 28.36 8.24 28.53 8.41 ;
        RECT 28.36 4.055 28.53 4.225 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 43.545 4 43.885 4.35 ;
        RECT 43.54 8.15 43.88 8.5 ;
        RECT 43.62 4 43.795 8.5 ;
      LAYER li1 ;
        RECT 43.62 2.955 43.79 4.225 ;
        RECT 43.62 8.24 43.79 9.51 ;
        RECT 37.985 8.24 38.155 9.51 ;
      LAYER met1 ;
        RECT 43.545 4.055 44.02 4.225 ;
        RECT 43.545 4 43.885 4.35 ;
        RECT 43.54 8.24 44.02 8.41 ;
        RECT 43.54 8.15 43.88 8.5 ;
        RECT 37.925 8.235 43.88 8.405 ;
        RECT 37.925 8.235 38.385 8.41 ;
        RECT 37.925 8.21 38.215 8.44 ;
      LAYER via1 ;
        RECT 43.64 8.25 43.79 8.4 ;
        RECT 43.645 4.1 43.795 4.25 ;
      LAYER mcon ;
        RECT 37.985 8.24 38.155 8.41 ;
        RECT 43.62 8.24 43.79 8.41 ;
        RECT 43.62 4.055 43.79 4.225 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 58.805 4 59.145 4.35 ;
        RECT 58.8 8.15 59.14 8.5 ;
        RECT 58.88 4 59.055 8.5 ;
      LAYER li1 ;
        RECT 58.88 2.955 59.05 4.225 ;
        RECT 58.88 8.24 59.05 9.51 ;
        RECT 53.245 8.24 53.415 9.51 ;
      LAYER met1 ;
        RECT 58.805 4.055 59.28 4.225 ;
        RECT 58.805 4 59.145 4.35 ;
        RECT 58.8 8.24 59.28 8.41 ;
        RECT 58.8 8.15 59.14 8.5 ;
        RECT 53.185 8.235 59.14 8.405 ;
        RECT 53.185 8.235 53.645 8.41 ;
        RECT 53.185 8.21 53.475 8.44 ;
      LAYER via1 ;
        RECT 58.9 8.25 59.05 8.4 ;
        RECT 58.905 4.1 59.055 4.25 ;
      LAYER mcon ;
        RECT 53.245 8.24 53.415 8.41 ;
        RECT 58.88 8.24 59.05 8.41 ;
        RECT 58.88 4.055 59.05 4.225 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 74.065 4 74.405 4.35 ;
        RECT 74.06 8.15 74.4 8.5 ;
        RECT 74.14 4 74.315 8.5 ;
      LAYER li1 ;
        RECT 74.14 2.955 74.31 4.225 ;
        RECT 74.14 8.24 74.31 9.51 ;
        RECT 68.505 8.24 68.675 9.51 ;
      LAYER met1 ;
        RECT 74.065 4.055 74.54 4.225 ;
        RECT 74.065 4 74.405 4.35 ;
        RECT 74.06 8.24 74.54 8.41 ;
        RECT 74.06 8.15 74.4 8.5 ;
        RECT 68.445 8.235 74.4 8.405 ;
        RECT 68.445 8.235 68.905 8.41 ;
        RECT 68.445 8.21 68.735 8.44 ;
      LAYER via1 ;
        RECT 74.16 8.25 74.31 8.4 ;
        RECT 74.165 4.1 74.315 4.25 ;
      LAYER mcon ;
        RECT 68.505 8.24 68.675 8.41 ;
        RECT 74.14 8.24 74.31 8.41 ;
        RECT 74.14 4.055 74.31 4.225 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 89.325 4 89.665 4.35 ;
        RECT 89.32 8.15 89.66 8.5 ;
        RECT 89.4 4 89.575 8.5 ;
      LAYER li1 ;
        RECT 89.4 2.955 89.57 4.225 ;
        RECT 89.4 8.24 89.57 9.51 ;
        RECT 83.765 8.24 83.935 9.51 ;
      LAYER met1 ;
        RECT 89.325 4.055 89.8 4.225 ;
        RECT 89.325 4 89.665 4.35 ;
        RECT 89.32 8.24 89.8 8.41 ;
        RECT 89.32 8.15 89.66 8.5 ;
        RECT 83.705 8.235 89.66 8.405 ;
        RECT 83.705 8.235 84.165 8.41 ;
        RECT 83.705 8.21 83.995 8.44 ;
      LAYER via1 ;
        RECT 89.42 8.25 89.57 8.4 ;
        RECT 89.425 4.1 89.575 4.25 ;
      LAYER mcon ;
        RECT 83.765 8.24 83.935 8.41 ;
        RECT 89.4 8.24 89.57 8.41 ;
        RECT 89.4 4.055 89.57 4.225 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 15.23 8.24 15.4 9.51 ;
      LAYER met1 ;
        RECT 15.17 8.24 15.63 8.41 ;
        RECT 15.175 8.205 15.465 8.435 ;
        RECT 15.17 8.21 15.46 8.44 ;
      LAYER mcon ;
        RECT 15.23 8.24 15.4 8.41 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 5.435 94.1 7.035 ;
        RECT 79.59 5.43 94.1 7.035 ;
        RECT 89.22 5.43 93.945 7.04 ;
        RECT 89.22 5.425 93.94 7.04 ;
        RECT 93.125 5.425 93.295 7.77 ;
        RECT 93.12 4.695 93.29 7.04 ;
        RECT 92.135 4.695 92.305 7.77 ;
        RECT 89.39 4.695 89.56 7.77 ;
        RECT 86.62 4.93 86.79 7.035 ;
        RECT 83.585 5.43 86.335 7.04 ;
        RECT 84.7 4.93 84.87 7.04 ;
        RECT 83.76 4.93 83.93 7.04 ;
        RECT 83.755 5.43 83.925 7.77 ;
        RECT 82.3 4.93 82.47 7.035 ;
        RECT 80.38 4.93 80.55 7.035 ;
        RECT 64.33 5.43 78.84 7.035 ;
        RECT 73.96 5.43 78.685 7.04 ;
        RECT 73.96 5.425 78.68 7.04 ;
        RECT 77.865 5.425 78.035 7.77 ;
        RECT 77.86 4.695 78.03 7.04 ;
        RECT 76.875 4.695 77.045 7.77 ;
        RECT 74.13 4.695 74.3 7.77 ;
        RECT 71.36 4.93 71.53 7.035 ;
        RECT 68.325 5.43 71.075 7.04 ;
        RECT 69.44 4.93 69.61 7.04 ;
        RECT 68.5 4.93 68.67 7.04 ;
        RECT 68.495 5.43 68.665 7.77 ;
        RECT 67.04 4.93 67.21 7.035 ;
        RECT 65.12 4.93 65.29 7.035 ;
        RECT 49.07 5.43 63.58 7.035 ;
        RECT 58.7 5.43 63.425 7.04 ;
        RECT 58.7 5.425 63.42 7.04 ;
        RECT 62.605 5.425 62.775 7.77 ;
        RECT 62.6 4.695 62.77 7.04 ;
        RECT 61.615 4.695 61.785 7.77 ;
        RECT 58.87 4.695 59.04 7.77 ;
        RECT 56.1 4.93 56.27 7.035 ;
        RECT 53.065 5.43 55.815 7.04 ;
        RECT 54.18 4.93 54.35 7.04 ;
        RECT 53.24 4.93 53.41 7.04 ;
        RECT 53.235 5.43 53.405 7.77 ;
        RECT 51.78 4.93 51.95 7.035 ;
        RECT 49.86 4.93 50.03 7.035 ;
        RECT 33.81 5.43 48.32 7.035 ;
        RECT 43.44 5.43 48.165 7.04 ;
        RECT 43.44 5.425 48.16 7.04 ;
        RECT 47.345 5.425 47.515 7.77 ;
        RECT 47.34 4.695 47.51 7.04 ;
        RECT 46.355 4.695 46.525 7.77 ;
        RECT 43.61 4.695 43.78 7.77 ;
        RECT 40.84 4.93 41.01 7.035 ;
        RECT 37.805 5.43 40.555 7.04 ;
        RECT 38.92 4.93 39.09 7.04 ;
        RECT 37.98 4.93 38.15 7.04 ;
        RECT 37.975 5.43 38.145 7.77 ;
        RECT 36.52 4.93 36.69 7.035 ;
        RECT 34.6 4.93 34.77 7.035 ;
        RECT 18.55 5.43 33.06 7.035 ;
        RECT 28.18 5.43 32.905 7.04 ;
        RECT 28.18 5.425 32.9 7.04 ;
        RECT 32.085 5.425 32.255 7.77 ;
        RECT 32.08 4.695 32.25 7.04 ;
        RECT 31.095 4.695 31.265 7.77 ;
        RECT 28.35 4.695 28.52 7.77 ;
        RECT 25.58 4.93 25.75 7.035 ;
        RECT 22.545 5.43 25.295 7.04 ;
        RECT 23.66 4.93 23.83 7.04 ;
        RECT 22.72 4.93 22.89 7.04 ;
        RECT 22.715 5.43 22.885 7.77 ;
        RECT 21.26 4.93 21.43 7.035 ;
        RECT 19.34 4.93 19.51 7.035 ;
        RECT 15.05 5.435 17.8 7.04 ;
        RECT 17.035 10.05 17.21 10.6 ;
        RECT 17.035 7.31 17.21 8.45 ;
        RECT 17.035 5.435 17.205 10.6 ;
        RECT 15.22 5.435 15.39 7.77 ;
      LAYER met1 ;
        RECT 0 5.435 94.1 7.035 ;
        RECT 79.59 5.43 94.1 7.035 ;
        RECT 89.22 5.43 93.945 7.04 ;
        RECT 89.22 5.425 93.94 7.04 ;
        RECT 79.59 5.275 88.33 7.035 ;
        RECT 83.585 5.275 86.335 7.04 ;
        RECT 64.33 5.43 78.84 7.035 ;
        RECT 73.96 5.43 78.685 7.04 ;
        RECT 73.96 5.425 78.68 7.04 ;
        RECT 64.33 5.275 73.07 7.035 ;
        RECT 68.325 5.275 71.075 7.04 ;
        RECT 49.07 5.43 63.58 7.035 ;
        RECT 58.7 5.43 63.425 7.04 ;
        RECT 58.7 5.425 63.42 7.04 ;
        RECT 49.07 5.275 57.81 7.035 ;
        RECT 53.065 5.275 55.815 7.04 ;
        RECT 33.81 5.43 48.32 7.035 ;
        RECT 43.44 5.43 48.165 7.04 ;
        RECT 43.44 5.425 48.16 7.04 ;
        RECT 33.81 5.275 42.55 7.035 ;
        RECT 37.805 5.275 40.555 7.04 ;
        RECT 18.55 5.43 33.06 7.035 ;
        RECT 28.18 5.43 32.905 7.04 ;
        RECT 28.18 5.425 32.9 7.04 ;
        RECT 18.55 5.275 27.29 7.035 ;
        RECT 22.545 5.275 25.295 7.04 ;
        RECT 15.05 5.435 17.8 7.04 ;
        RECT 16.975 8.95 17.265 9.18 ;
        RECT 16.805 8.98 17.265 9.15 ;
      LAYER mcon ;
        RECT 17.035 8.98 17.205 9.15 ;
        RECT 17.34 6.84 17.51 7.01 ;
        RECT 18.695 5.43 18.865 5.6 ;
        RECT 19.155 5.43 19.325 5.6 ;
        RECT 19.615 5.43 19.785 5.6 ;
        RECT 20.075 5.43 20.245 5.6 ;
        RECT 20.535 5.43 20.705 5.6 ;
        RECT 20.995 5.43 21.165 5.6 ;
        RECT 21.455 5.43 21.625 5.6 ;
        RECT 21.915 5.43 22.085 5.6 ;
        RECT 22.375 5.43 22.545 5.6 ;
        RECT 22.835 5.43 23.005 5.6 ;
        RECT 23.295 5.43 23.465 5.6 ;
        RECT 23.755 5.43 23.925 5.6 ;
        RECT 24.215 5.43 24.385 5.6 ;
        RECT 24.675 5.43 24.845 5.6 ;
        RECT 24.835 6.84 25.005 7.01 ;
        RECT 25.135 5.43 25.305 5.6 ;
        RECT 25.595 5.43 25.765 5.6 ;
        RECT 26.055 5.43 26.225 5.6 ;
        RECT 26.515 5.43 26.685 5.6 ;
        RECT 26.975 5.43 27.145 5.6 ;
        RECT 30.47 6.84 30.64 7.01 ;
        RECT 30.47 5.455 30.64 5.625 ;
        RECT 31.175 6.84 31.345 7.01 ;
        RECT 31.175 5.455 31.345 5.625 ;
        RECT 32.16 5.455 32.33 5.625 ;
        RECT 32.165 6.84 32.335 7.01 ;
        RECT 33.955 5.43 34.125 5.6 ;
        RECT 34.415 5.43 34.585 5.6 ;
        RECT 34.875 5.43 35.045 5.6 ;
        RECT 35.335 5.43 35.505 5.6 ;
        RECT 35.795 5.43 35.965 5.6 ;
        RECT 36.255 5.43 36.425 5.6 ;
        RECT 36.715 5.43 36.885 5.6 ;
        RECT 37.175 5.43 37.345 5.6 ;
        RECT 37.635 5.43 37.805 5.6 ;
        RECT 38.095 5.43 38.265 5.6 ;
        RECT 38.555 5.43 38.725 5.6 ;
        RECT 39.015 5.43 39.185 5.6 ;
        RECT 39.475 5.43 39.645 5.6 ;
        RECT 39.935 5.43 40.105 5.6 ;
        RECT 40.095 6.84 40.265 7.01 ;
        RECT 40.395 5.43 40.565 5.6 ;
        RECT 40.855 5.43 41.025 5.6 ;
        RECT 41.315 5.43 41.485 5.6 ;
        RECT 41.775 5.43 41.945 5.6 ;
        RECT 42.235 5.43 42.405 5.6 ;
        RECT 45.73 6.84 45.9 7.01 ;
        RECT 45.73 5.455 45.9 5.625 ;
        RECT 46.435 6.84 46.605 7.01 ;
        RECT 46.435 5.455 46.605 5.625 ;
        RECT 47.42 5.455 47.59 5.625 ;
        RECT 47.425 6.84 47.595 7.01 ;
        RECT 49.215 5.43 49.385 5.6 ;
        RECT 49.675 5.43 49.845 5.6 ;
        RECT 50.135 5.43 50.305 5.6 ;
        RECT 50.595 5.43 50.765 5.6 ;
        RECT 51.055 5.43 51.225 5.6 ;
        RECT 51.515 5.43 51.685 5.6 ;
        RECT 51.975 5.43 52.145 5.6 ;
        RECT 52.435 5.43 52.605 5.6 ;
        RECT 52.895 5.43 53.065 5.6 ;
        RECT 53.355 5.43 53.525 5.6 ;
        RECT 53.815 5.43 53.985 5.6 ;
        RECT 54.275 5.43 54.445 5.6 ;
        RECT 54.735 5.43 54.905 5.6 ;
        RECT 55.195 5.43 55.365 5.6 ;
        RECT 55.355 6.84 55.525 7.01 ;
        RECT 55.655 5.43 55.825 5.6 ;
        RECT 56.115 5.43 56.285 5.6 ;
        RECT 56.575 5.43 56.745 5.6 ;
        RECT 57.035 5.43 57.205 5.6 ;
        RECT 57.495 5.43 57.665 5.6 ;
        RECT 60.99 6.84 61.16 7.01 ;
        RECT 60.99 5.455 61.16 5.625 ;
        RECT 61.695 6.84 61.865 7.01 ;
        RECT 61.695 5.455 61.865 5.625 ;
        RECT 62.68 5.455 62.85 5.625 ;
        RECT 62.685 6.84 62.855 7.01 ;
        RECT 64.475 5.43 64.645 5.6 ;
        RECT 64.935 5.43 65.105 5.6 ;
        RECT 65.395 5.43 65.565 5.6 ;
        RECT 65.855 5.43 66.025 5.6 ;
        RECT 66.315 5.43 66.485 5.6 ;
        RECT 66.775 5.43 66.945 5.6 ;
        RECT 67.235 5.43 67.405 5.6 ;
        RECT 67.695 5.43 67.865 5.6 ;
        RECT 68.155 5.43 68.325 5.6 ;
        RECT 68.615 5.43 68.785 5.6 ;
        RECT 69.075 5.43 69.245 5.6 ;
        RECT 69.535 5.43 69.705 5.6 ;
        RECT 69.995 5.43 70.165 5.6 ;
        RECT 70.455 5.43 70.625 5.6 ;
        RECT 70.615 6.84 70.785 7.01 ;
        RECT 70.915 5.43 71.085 5.6 ;
        RECT 71.375 5.43 71.545 5.6 ;
        RECT 71.835 5.43 72.005 5.6 ;
        RECT 72.295 5.43 72.465 5.6 ;
        RECT 72.755 5.43 72.925 5.6 ;
        RECT 76.25 6.84 76.42 7.01 ;
        RECT 76.25 5.455 76.42 5.625 ;
        RECT 76.955 6.84 77.125 7.01 ;
        RECT 76.955 5.455 77.125 5.625 ;
        RECT 77.94 5.455 78.11 5.625 ;
        RECT 77.945 6.84 78.115 7.01 ;
        RECT 79.735 5.43 79.905 5.6 ;
        RECT 80.195 5.43 80.365 5.6 ;
        RECT 80.655 5.43 80.825 5.6 ;
        RECT 81.115 5.43 81.285 5.6 ;
        RECT 81.575 5.43 81.745 5.6 ;
        RECT 82.035 5.43 82.205 5.6 ;
        RECT 82.495 5.43 82.665 5.6 ;
        RECT 82.955 5.43 83.125 5.6 ;
        RECT 83.415 5.43 83.585 5.6 ;
        RECT 83.875 5.43 84.045 5.6 ;
        RECT 84.335 5.43 84.505 5.6 ;
        RECT 84.795 5.43 84.965 5.6 ;
        RECT 85.255 5.43 85.425 5.6 ;
        RECT 85.715 5.43 85.885 5.6 ;
        RECT 85.875 6.84 86.045 7.01 ;
        RECT 86.175 5.43 86.345 5.6 ;
        RECT 86.635 5.43 86.805 5.6 ;
        RECT 87.095 5.43 87.265 5.6 ;
        RECT 87.555 5.43 87.725 5.6 ;
        RECT 88.015 5.43 88.185 5.6 ;
        RECT 91.51 6.84 91.68 7.01 ;
        RECT 91.51 5.455 91.68 5.625 ;
        RECT 92.215 6.84 92.385 7.01 ;
        RECT 92.215 5.455 92.385 5.625 ;
        RECT 93.2 5.455 93.37 5.625 ;
        RECT 93.205 6.84 93.375 7.01 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 81.5 3.31 81.83 4.04 ;
        RECT 66.24 3.31 66.57 4.04 ;
        RECT 50.98 3.31 51.31 4.04 ;
        RECT 35.72 3.31 36.05 4.04 ;
        RECT 20.46 3.31 20.79 4.04 ;
      LAYER met2 ;
        RECT 81.605 2.24 81.975 2.61 ;
        RECT 81.615 3.625 81.875 3.885 ;
        RECT 81.705 2.24 81.87 3.885 ;
        RECT 81.525 3.735 81.825 3.935 ;
        RECT 81.525 3.735 81.805 4.015 ;
        RECT 81.58 3.72 81.875 3.885 ;
        RECT 66.345 2.24 66.715 2.61 ;
        RECT 66.355 3.625 66.615 3.885 ;
        RECT 66.445 2.24 66.61 3.885 ;
        RECT 66.265 3.735 66.565 3.935 ;
        RECT 66.265 3.735 66.545 4.015 ;
        RECT 66.32 3.72 66.615 3.885 ;
        RECT 51.085 2.24 51.455 2.61 ;
        RECT 51.095 3.625 51.355 3.885 ;
        RECT 51.185 2.24 51.35 3.885 ;
        RECT 51.005 3.735 51.305 3.935 ;
        RECT 51.005 3.735 51.285 4.015 ;
        RECT 51.06 3.72 51.355 3.885 ;
        RECT 35.825 2.24 36.195 2.61 ;
        RECT 35.835 3.625 36.095 3.885 ;
        RECT 35.925 2.24 36.09 3.885 ;
        RECT 35.745 3.735 36.045 3.935 ;
        RECT 35.745 3.735 36.025 4.015 ;
        RECT 35.8 3.72 36.095 3.885 ;
        RECT 20.565 2.24 20.935 2.61 ;
        RECT 20.575 3.625 20.835 3.885 ;
        RECT 20.665 2.24 20.83 3.885 ;
        RECT 20.485 3.735 20.785 3.935 ;
        RECT 20.485 3.735 20.765 4.015 ;
        RECT 20.54 3.72 20.835 3.885 ;
      LAYER li1 ;
        RECT 0.005 0 94.1 1.6 ;
        RECT 93.12 0 93.29 2.225 ;
        RECT 92.135 0 92.305 2.225 ;
        RECT 89.39 0 89.56 2.225 ;
        RECT 79.59 0 88.33 2.88 ;
        RECT 87.56 0 87.73 3.38 ;
        RECT 86.62 0 86.79 3.38 ;
        RECT 85.66 0 85.83 3.38 ;
        RECT 84.615 0 84.81 2.89 ;
        RECT 83.74 0 83.91 3.38 ;
        RECT 82.78 0 82.95 3.38 ;
        RECT 80.86 0 81.135 2.89 ;
        RECT 80.86 0 81.03 3.38 ;
        RECT 77.86 0 78.03 2.225 ;
        RECT 76.875 0 77.045 2.225 ;
        RECT 74.13 0 74.3 2.225 ;
        RECT 64.33 0 73.07 2.88 ;
        RECT 72.3 0 72.47 3.38 ;
        RECT 71.36 0 71.53 3.38 ;
        RECT 70.4 0 70.57 3.38 ;
        RECT 69.355 0 69.55 2.89 ;
        RECT 68.48 0 68.65 3.38 ;
        RECT 67.52 0 67.69 3.38 ;
        RECT 65.6 0 65.875 2.89 ;
        RECT 65.6 0 65.77 3.38 ;
        RECT 62.6 0 62.77 2.225 ;
        RECT 61.615 0 61.785 2.225 ;
        RECT 58.87 0 59.04 2.225 ;
        RECT 49.07 0 57.81 2.88 ;
        RECT 57.04 0 57.21 3.38 ;
        RECT 56.1 0 56.27 3.38 ;
        RECT 55.14 0 55.31 3.38 ;
        RECT 54.095 0 54.29 2.89 ;
        RECT 53.22 0 53.39 3.38 ;
        RECT 52.26 0 52.43 3.38 ;
        RECT 50.34 0 50.615 2.89 ;
        RECT 50.34 0 50.51 3.38 ;
        RECT 47.34 0 47.51 2.225 ;
        RECT 46.355 0 46.525 2.225 ;
        RECT 43.61 0 43.78 2.225 ;
        RECT 33.81 0 42.55 2.88 ;
        RECT 41.78 0 41.95 3.38 ;
        RECT 40.84 0 41.01 3.38 ;
        RECT 39.88 0 40.05 3.38 ;
        RECT 38.835 0 39.03 2.89 ;
        RECT 37.96 0 38.13 3.38 ;
        RECT 37 0 37.17 3.38 ;
        RECT 35.08 0 35.355 2.89 ;
        RECT 35.08 0 35.25 3.38 ;
        RECT 32.08 0 32.25 2.225 ;
        RECT 31.095 0 31.265 2.225 ;
        RECT 28.35 0 28.52 2.225 ;
        RECT 18.55 0 27.29 2.88 ;
        RECT 26.52 0 26.69 3.38 ;
        RECT 25.58 0 25.75 3.38 ;
        RECT 24.62 0 24.79 3.38 ;
        RECT 23.575 0 23.77 2.89 ;
        RECT 22.7 0 22.87 3.38 ;
        RECT 21.74 0 21.91 3.38 ;
        RECT 19.82 0 20.095 2.89 ;
        RECT 19.82 0 19.99 3.38 ;
        RECT 0.01 10.865 94.1 12.465 ;
        RECT 93.125 10.24 93.295 12.465 ;
        RECT 92.135 10.24 92.305 12.465 ;
        RECT 89.39 10.24 89.56 12.465 ;
        RECT 83.755 10.24 83.925 12.465 ;
        RECT 77.865 10.24 78.035 12.465 ;
        RECT 76.875 10.24 77.045 12.465 ;
        RECT 74.13 10.24 74.3 12.465 ;
        RECT 68.495 10.24 68.665 12.465 ;
        RECT 62.605 10.24 62.775 12.465 ;
        RECT 61.615 10.24 61.785 12.465 ;
        RECT 58.87 10.24 59.04 12.465 ;
        RECT 53.235 10.24 53.405 12.465 ;
        RECT 47.345 10.24 47.515 12.465 ;
        RECT 46.355 10.24 46.525 12.465 ;
        RECT 43.61 10.24 43.78 12.465 ;
        RECT 37.975 10.24 38.145 12.465 ;
        RECT 32.085 10.24 32.255 12.465 ;
        RECT 31.095 10.24 31.265 12.465 ;
        RECT 28.35 10.24 28.52 12.465 ;
        RECT 22.715 10.24 22.885 12.465 ;
        RECT 15.22 10.24 15.39 12.465 ;
        RECT 84.77 8.37 84.94 10.32 ;
        RECT 84.71 10.15 84.88 10.6 ;
        RECT 84.71 7.31 84.88 8.54 ;
        RECT 81.475 3.62 81.825 4.04 ;
        RECT 81.455 3.62 81.825 3.91 ;
        RECT 81.45 3.62 81.825 3.875 ;
        RECT 81.44 3.62 81.825 3.87 ;
        RECT 81.41 3.62 81.825 3.855 ;
        RECT 80.115 3.585 81.435 3.765 ;
        RECT 81.385 3.62 81.825 3.815 ;
        RECT 81.355 3.62 81.825 3.785 ;
        RECT 80.115 3.58 81.23 3.765 ;
        RECT 80.115 3.575 81.225 3.765 ;
        RECT 80.115 3.57 81.185 3.765 ;
        RECT 80.115 3.565 81.18 3.765 ;
        RECT 80.115 3.56 81.155 3.765 ;
        RECT 80.115 3.555 81.145 3.765 ;
        RECT 80.115 3.535 81.105 3.765 ;
        RECT 80.115 3.535 80.47 3.77 ;
        RECT 80.115 3.535 80.445 3.865 ;
        RECT 80.115 3.535 80.405 3.88 ;
        RECT 80.115 3.535 80.395 4.055 ;
        RECT 69.51 8.37 69.68 10.32 ;
        RECT 69.45 10.15 69.62 10.6 ;
        RECT 69.45 7.31 69.62 8.54 ;
        RECT 66.215 3.62 66.565 4.04 ;
        RECT 66.195 3.62 66.565 3.91 ;
        RECT 66.19 3.62 66.565 3.875 ;
        RECT 66.18 3.62 66.565 3.87 ;
        RECT 66.15 3.62 66.565 3.855 ;
        RECT 64.855 3.585 66.175 3.765 ;
        RECT 66.125 3.62 66.565 3.815 ;
        RECT 66.095 3.62 66.565 3.785 ;
        RECT 64.855 3.58 65.97 3.765 ;
        RECT 64.855 3.575 65.965 3.765 ;
        RECT 64.855 3.57 65.925 3.765 ;
        RECT 64.855 3.565 65.92 3.765 ;
        RECT 64.855 3.56 65.895 3.765 ;
        RECT 64.855 3.555 65.885 3.765 ;
        RECT 64.855 3.535 65.845 3.765 ;
        RECT 64.855 3.535 65.21 3.77 ;
        RECT 64.855 3.535 65.185 3.865 ;
        RECT 64.855 3.535 65.145 3.88 ;
        RECT 64.855 3.535 65.135 4.055 ;
        RECT 54.25 8.37 54.42 10.32 ;
        RECT 54.19 10.15 54.36 10.6 ;
        RECT 54.19 7.31 54.36 8.54 ;
        RECT 50.955 3.62 51.305 4.04 ;
        RECT 50.935 3.62 51.305 3.91 ;
        RECT 50.93 3.62 51.305 3.875 ;
        RECT 50.92 3.62 51.305 3.87 ;
        RECT 50.89 3.62 51.305 3.855 ;
        RECT 49.595 3.585 50.915 3.765 ;
        RECT 50.865 3.62 51.305 3.815 ;
        RECT 50.835 3.62 51.305 3.785 ;
        RECT 49.595 3.58 50.71 3.765 ;
        RECT 49.595 3.575 50.705 3.765 ;
        RECT 49.595 3.57 50.665 3.765 ;
        RECT 49.595 3.565 50.66 3.765 ;
        RECT 49.595 3.56 50.635 3.765 ;
        RECT 49.595 3.555 50.625 3.765 ;
        RECT 49.595 3.535 50.585 3.765 ;
        RECT 49.595 3.535 49.95 3.77 ;
        RECT 49.595 3.535 49.925 3.865 ;
        RECT 49.595 3.535 49.885 3.88 ;
        RECT 49.595 3.535 49.875 4.055 ;
        RECT 38.99 8.37 39.16 10.32 ;
        RECT 38.93 10.15 39.1 10.6 ;
        RECT 38.93 7.31 39.1 8.54 ;
        RECT 35.695 3.62 36.045 4.04 ;
        RECT 35.675 3.62 36.045 3.91 ;
        RECT 35.67 3.62 36.045 3.875 ;
        RECT 35.66 3.62 36.045 3.87 ;
        RECT 35.63 3.62 36.045 3.855 ;
        RECT 34.335 3.585 35.655 3.765 ;
        RECT 35.605 3.62 36.045 3.815 ;
        RECT 35.575 3.62 36.045 3.785 ;
        RECT 34.335 3.58 35.45 3.765 ;
        RECT 34.335 3.575 35.445 3.765 ;
        RECT 34.335 3.57 35.405 3.765 ;
        RECT 34.335 3.565 35.4 3.765 ;
        RECT 34.335 3.56 35.375 3.765 ;
        RECT 34.335 3.555 35.365 3.765 ;
        RECT 34.335 3.535 35.325 3.765 ;
        RECT 34.335 3.535 34.69 3.77 ;
        RECT 34.335 3.535 34.665 3.865 ;
        RECT 34.335 3.535 34.625 3.88 ;
        RECT 34.335 3.535 34.615 4.055 ;
        RECT 23.73 8.37 23.9 10.32 ;
        RECT 23.67 10.15 23.84 10.6 ;
        RECT 23.67 7.31 23.84 8.54 ;
        RECT 20.435 3.62 20.785 4.04 ;
        RECT 20.415 3.62 20.785 3.91 ;
        RECT 20.41 3.62 20.785 3.875 ;
        RECT 20.4 3.62 20.785 3.87 ;
        RECT 20.37 3.62 20.785 3.855 ;
        RECT 19.075 3.585 20.395 3.765 ;
        RECT 20.345 3.62 20.785 3.815 ;
        RECT 20.315 3.62 20.785 3.785 ;
        RECT 19.075 3.58 20.19 3.765 ;
        RECT 19.075 3.575 20.185 3.765 ;
        RECT 19.075 3.57 20.145 3.765 ;
        RECT 19.075 3.565 20.14 3.765 ;
        RECT 19.075 3.56 20.115 3.765 ;
        RECT 19.075 3.555 20.105 3.765 ;
        RECT 19.075 3.535 20.065 3.765 ;
        RECT 19.075 3.535 19.43 3.77 ;
        RECT 19.075 3.535 19.405 3.865 ;
        RECT 19.075 3.535 19.365 3.88 ;
        RECT 19.075 3.535 19.355 4.055 ;
      LAYER met1 ;
        RECT 0.005 0 94.1 1.6 ;
        RECT 79.59 0 88.33 3.035 ;
        RECT 64.33 0 73.07 3.035 ;
        RECT 49.07 0 57.81 3.035 ;
        RECT 33.81 0 42.55 3.035 ;
        RECT 18.55 0 27.29 3.035 ;
        RECT 0.01 10.865 94.1 12.465 ;
        RECT 84.71 8.58 85 8.81 ;
        RECT 84.535 8.61 85 8.78 ;
        RECT 84.535 8.605 84.705 12.465 ;
        RECT 69.45 8.58 69.74 8.81 ;
        RECT 69.275 8.61 69.74 8.78 ;
        RECT 69.275 8.605 69.445 12.465 ;
        RECT 54.19 8.58 54.48 8.81 ;
        RECT 54.015 8.61 54.48 8.78 ;
        RECT 54.015 8.605 54.185 12.465 ;
        RECT 38.93 8.58 39.22 8.81 ;
        RECT 38.755 8.61 39.22 8.78 ;
        RECT 38.755 8.605 38.925 12.465 ;
        RECT 23.67 8.58 23.96 8.81 ;
        RECT 23.495 8.61 23.96 8.78 ;
        RECT 23.495 8.605 23.665 12.465 ;
        RECT 81.455 3.625 81.875 3.885 ;
        RECT 81.455 3.62 81.825 3.91 ;
        RECT 81.475 3.62 81.82 3.93 ;
        RECT 66.195 3.625 66.615 3.885 ;
        RECT 66.195 3.62 66.565 3.91 ;
        RECT 66.215 3.62 66.56 3.93 ;
        RECT 50.935 3.625 51.355 3.885 ;
        RECT 50.935 3.62 51.305 3.91 ;
        RECT 50.955 3.62 51.3 3.93 ;
        RECT 35.675 3.625 36.095 3.885 ;
        RECT 35.675 3.62 36.045 3.91 ;
        RECT 35.695 3.62 36.04 3.93 ;
        RECT 20.415 3.625 20.835 3.885 ;
        RECT 20.415 3.62 20.785 3.91 ;
        RECT 20.435 3.62 20.78 3.93 ;
      LAYER via1 ;
        RECT 20.63 3.68 20.78 3.83 ;
        RECT 20.675 2.35 20.825 2.5 ;
        RECT 35.89 3.68 36.04 3.83 ;
        RECT 35.935 2.35 36.085 2.5 ;
        RECT 51.15 3.68 51.3 3.83 ;
        RECT 51.195 2.35 51.345 2.5 ;
        RECT 66.41 3.68 66.56 3.83 ;
        RECT 66.455 2.35 66.605 2.5 ;
        RECT 81.67 3.68 81.82 3.83 ;
        RECT 81.715 2.35 81.865 2.5 ;
      LAYER via2 ;
        RECT 20.525 3.775 20.725 3.975 ;
        RECT 35.785 3.775 35.985 3.975 ;
        RECT 51.045 3.775 51.245 3.975 ;
        RECT 66.305 3.775 66.505 3.975 ;
        RECT 81.565 3.775 81.765 3.975 ;
      LAYER mcon ;
        RECT 15.3 10.9 15.47 11.07 ;
        RECT 15.98 10.9 16.15 11.07 ;
        RECT 16.66 10.9 16.83 11.07 ;
        RECT 17.34 10.9 17.51 11.07 ;
        RECT 18.695 2.71 18.865 2.88 ;
        RECT 19.155 2.71 19.325 2.88 ;
        RECT 19.615 2.71 19.785 2.88 ;
        RECT 20.075 2.71 20.245 2.88 ;
        RECT 20.525 3.71 20.695 3.88 ;
        RECT 20.535 2.71 20.705 2.88 ;
        RECT 20.995 2.71 21.165 2.88 ;
        RECT 21.455 2.71 21.625 2.88 ;
        RECT 21.915 2.71 22.085 2.88 ;
        RECT 22.375 2.71 22.545 2.88 ;
        RECT 22.795 10.9 22.965 11.07 ;
        RECT 22.835 2.71 23.005 2.88 ;
        RECT 23.295 2.71 23.465 2.88 ;
        RECT 23.475 10.9 23.645 11.07 ;
        RECT 23.73 8.61 23.9 8.78 ;
        RECT 23.755 2.71 23.925 2.88 ;
        RECT 24.155 10.9 24.325 11.07 ;
        RECT 24.215 2.71 24.385 2.88 ;
        RECT 24.675 2.71 24.845 2.88 ;
        RECT 24.835 10.9 25.005 11.07 ;
        RECT 25.135 2.71 25.305 2.88 ;
        RECT 25.595 2.71 25.765 2.88 ;
        RECT 26.055 2.71 26.225 2.88 ;
        RECT 26.515 2.71 26.685 2.88 ;
        RECT 26.975 2.71 27.145 2.88 ;
        RECT 28.43 10.9 28.6 11.07 ;
        RECT 28.43 1.395 28.6 1.565 ;
        RECT 29.11 10.9 29.28 11.07 ;
        RECT 29.11 1.395 29.28 1.565 ;
        RECT 29.79 10.9 29.96 11.07 ;
        RECT 29.79 1.395 29.96 1.565 ;
        RECT 30.47 10.9 30.64 11.07 ;
        RECT 30.47 1.395 30.64 1.565 ;
        RECT 31.175 10.9 31.345 11.07 ;
        RECT 31.175 1.395 31.345 1.565 ;
        RECT 32.16 1.395 32.33 1.565 ;
        RECT 32.165 10.9 32.335 11.07 ;
        RECT 33.955 2.71 34.125 2.88 ;
        RECT 34.415 2.71 34.585 2.88 ;
        RECT 34.875 2.71 35.045 2.88 ;
        RECT 35.335 2.71 35.505 2.88 ;
        RECT 35.785 3.71 35.955 3.88 ;
        RECT 35.795 2.71 35.965 2.88 ;
        RECT 36.255 2.71 36.425 2.88 ;
        RECT 36.715 2.71 36.885 2.88 ;
        RECT 37.175 2.71 37.345 2.88 ;
        RECT 37.635 2.71 37.805 2.88 ;
        RECT 38.055 10.9 38.225 11.07 ;
        RECT 38.095 2.71 38.265 2.88 ;
        RECT 38.555 2.71 38.725 2.88 ;
        RECT 38.735 10.9 38.905 11.07 ;
        RECT 38.99 8.61 39.16 8.78 ;
        RECT 39.015 2.71 39.185 2.88 ;
        RECT 39.415 10.9 39.585 11.07 ;
        RECT 39.475 2.71 39.645 2.88 ;
        RECT 39.935 2.71 40.105 2.88 ;
        RECT 40.095 10.9 40.265 11.07 ;
        RECT 40.395 2.71 40.565 2.88 ;
        RECT 40.855 2.71 41.025 2.88 ;
        RECT 41.315 2.71 41.485 2.88 ;
        RECT 41.775 2.71 41.945 2.88 ;
        RECT 42.235 2.71 42.405 2.88 ;
        RECT 43.69 10.9 43.86 11.07 ;
        RECT 43.69 1.395 43.86 1.565 ;
        RECT 44.37 10.9 44.54 11.07 ;
        RECT 44.37 1.395 44.54 1.565 ;
        RECT 45.05 10.9 45.22 11.07 ;
        RECT 45.05 1.395 45.22 1.565 ;
        RECT 45.73 10.9 45.9 11.07 ;
        RECT 45.73 1.395 45.9 1.565 ;
        RECT 46.435 10.9 46.605 11.07 ;
        RECT 46.435 1.395 46.605 1.565 ;
        RECT 47.42 1.395 47.59 1.565 ;
        RECT 47.425 10.9 47.595 11.07 ;
        RECT 49.215 2.71 49.385 2.88 ;
        RECT 49.675 2.71 49.845 2.88 ;
        RECT 50.135 2.71 50.305 2.88 ;
        RECT 50.595 2.71 50.765 2.88 ;
        RECT 51.045 3.71 51.215 3.88 ;
        RECT 51.055 2.71 51.225 2.88 ;
        RECT 51.515 2.71 51.685 2.88 ;
        RECT 51.975 2.71 52.145 2.88 ;
        RECT 52.435 2.71 52.605 2.88 ;
        RECT 52.895 2.71 53.065 2.88 ;
        RECT 53.315 10.9 53.485 11.07 ;
        RECT 53.355 2.71 53.525 2.88 ;
        RECT 53.815 2.71 53.985 2.88 ;
        RECT 53.995 10.9 54.165 11.07 ;
        RECT 54.25 8.61 54.42 8.78 ;
        RECT 54.275 2.71 54.445 2.88 ;
        RECT 54.675 10.9 54.845 11.07 ;
        RECT 54.735 2.71 54.905 2.88 ;
        RECT 55.195 2.71 55.365 2.88 ;
        RECT 55.355 10.9 55.525 11.07 ;
        RECT 55.655 2.71 55.825 2.88 ;
        RECT 56.115 2.71 56.285 2.88 ;
        RECT 56.575 2.71 56.745 2.88 ;
        RECT 57.035 2.71 57.205 2.88 ;
        RECT 57.495 2.71 57.665 2.88 ;
        RECT 58.95 10.9 59.12 11.07 ;
        RECT 58.95 1.395 59.12 1.565 ;
        RECT 59.63 10.9 59.8 11.07 ;
        RECT 59.63 1.395 59.8 1.565 ;
        RECT 60.31 10.9 60.48 11.07 ;
        RECT 60.31 1.395 60.48 1.565 ;
        RECT 60.99 10.9 61.16 11.07 ;
        RECT 60.99 1.395 61.16 1.565 ;
        RECT 61.695 10.9 61.865 11.07 ;
        RECT 61.695 1.395 61.865 1.565 ;
        RECT 62.68 1.395 62.85 1.565 ;
        RECT 62.685 10.9 62.855 11.07 ;
        RECT 64.475 2.71 64.645 2.88 ;
        RECT 64.935 2.71 65.105 2.88 ;
        RECT 65.395 2.71 65.565 2.88 ;
        RECT 65.855 2.71 66.025 2.88 ;
        RECT 66.305 3.71 66.475 3.88 ;
        RECT 66.315 2.71 66.485 2.88 ;
        RECT 66.775 2.71 66.945 2.88 ;
        RECT 67.235 2.71 67.405 2.88 ;
        RECT 67.695 2.71 67.865 2.88 ;
        RECT 68.155 2.71 68.325 2.88 ;
        RECT 68.575 10.9 68.745 11.07 ;
        RECT 68.615 2.71 68.785 2.88 ;
        RECT 69.075 2.71 69.245 2.88 ;
        RECT 69.255 10.9 69.425 11.07 ;
        RECT 69.51 8.61 69.68 8.78 ;
        RECT 69.535 2.71 69.705 2.88 ;
        RECT 69.935 10.9 70.105 11.07 ;
        RECT 69.995 2.71 70.165 2.88 ;
        RECT 70.455 2.71 70.625 2.88 ;
        RECT 70.615 10.9 70.785 11.07 ;
        RECT 70.915 2.71 71.085 2.88 ;
        RECT 71.375 2.71 71.545 2.88 ;
        RECT 71.835 2.71 72.005 2.88 ;
        RECT 72.295 2.71 72.465 2.88 ;
        RECT 72.755 2.71 72.925 2.88 ;
        RECT 74.21 10.9 74.38 11.07 ;
        RECT 74.21 1.395 74.38 1.565 ;
        RECT 74.89 10.9 75.06 11.07 ;
        RECT 74.89 1.395 75.06 1.565 ;
        RECT 75.57 10.9 75.74 11.07 ;
        RECT 75.57 1.395 75.74 1.565 ;
        RECT 76.25 10.9 76.42 11.07 ;
        RECT 76.25 1.395 76.42 1.565 ;
        RECT 76.955 10.9 77.125 11.07 ;
        RECT 76.955 1.395 77.125 1.565 ;
        RECT 77.94 1.395 78.11 1.565 ;
        RECT 77.945 10.9 78.115 11.07 ;
        RECT 79.735 2.71 79.905 2.88 ;
        RECT 80.195 2.71 80.365 2.88 ;
        RECT 80.655 2.71 80.825 2.88 ;
        RECT 81.115 2.71 81.285 2.88 ;
        RECT 81.565 3.71 81.735 3.88 ;
        RECT 81.575 2.71 81.745 2.88 ;
        RECT 82.035 2.71 82.205 2.88 ;
        RECT 82.495 2.71 82.665 2.88 ;
        RECT 82.955 2.71 83.125 2.88 ;
        RECT 83.415 2.71 83.585 2.88 ;
        RECT 83.835 10.9 84.005 11.07 ;
        RECT 83.875 2.71 84.045 2.88 ;
        RECT 84.335 2.71 84.505 2.88 ;
        RECT 84.515 10.9 84.685 11.07 ;
        RECT 84.77 8.61 84.94 8.78 ;
        RECT 84.795 2.71 84.965 2.88 ;
        RECT 85.195 10.9 85.365 11.07 ;
        RECT 85.255 2.71 85.425 2.88 ;
        RECT 85.715 2.71 85.885 2.88 ;
        RECT 85.875 10.9 86.045 11.07 ;
        RECT 86.175 2.71 86.345 2.88 ;
        RECT 86.635 2.71 86.805 2.88 ;
        RECT 87.095 2.71 87.265 2.88 ;
        RECT 87.555 2.71 87.725 2.88 ;
        RECT 88.015 2.71 88.185 2.88 ;
        RECT 89.47 10.9 89.64 11.07 ;
        RECT 89.47 1.395 89.64 1.565 ;
        RECT 90.15 10.9 90.32 11.07 ;
        RECT 90.15 1.395 90.32 1.565 ;
        RECT 90.83 10.9 91 11.07 ;
        RECT 90.83 1.395 91 1.565 ;
        RECT 91.51 10.9 91.68 11.07 ;
        RECT 91.51 1.395 91.68 1.565 ;
        RECT 92.215 10.9 92.385 11.07 ;
        RECT 92.215 1.395 92.385 1.565 ;
        RECT 93.2 1.395 93.37 1.565 ;
        RECT 93.205 10.9 93.375 11.07 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 85.04 9.345 85.41 9.715 ;
      RECT 85.075 5.565 85.375 9.715 ;
      RECT 80.885 5.565 85.375 6.86 ;
      RECT 84.065 3.15 84.365 6.86 ;
      RECT 80.885 3.73 81.185 6.86 ;
      RECT 84.02 4.055 84.365 4.785 ;
      RECT 80.78 3.31 81.11 4.04 ;
      RECT 83.66 3.15 84.39 3.48 ;
      RECT 69.78 9.345 70.15 9.715 ;
      RECT 69.815 5.565 70.115 9.715 ;
      RECT 65.625 5.565 70.115 6.86 ;
      RECT 68.805 3.15 69.105 6.86 ;
      RECT 65.625 3.73 65.925 6.86 ;
      RECT 68.76 4.055 69.105 4.785 ;
      RECT 65.52 3.31 65.85 4.04 ;
      RECT 68.4 3.15 69.13 3.48 ;
      RECT 54.52 9.345 54.89 9.715 ;
      RECT 54.555 5.565 54.855 9.715 ;
      RECT 50.365 5.565 54.855 6.86 ;
      RECT 53.545 3.15 53.845 6.86 ;
      RECT 50.365 3.73 50.665 6.86 ;
      RECT 53.5 4.055 53.845 4.785 ;
      RECT 50.26 3.31 50.59 4.04 ;
      RECT 53.14 3.15 53.87 3.48 ;
      RECT 39.26 9.345 39.63 9.715 ;
      RECT 39.295 5.565 39.595 9.715 ;
      RECT 35.105 5.565 39.595 6.86 ;
      RECT 38.285 3.15 38.585 6.86 ;
      RECT 35.105 3.73 35.405 6.86 ;
      RECT 38.24 4.055 38.585 4.785 ;
      RECT 35 3.31 35.33 4.04 ;
      RECT 37.88 3.15 38.61 3.48 ;
      RECT 24 9.345 24.37 9.715 ;
      RECT 24.035 5.565 24.335 9.715 ;
      RECT 19.845 5.565 24.335 6.86 ;
      RECT 23.025 3.15 23.325 6.86 ;
      RECT 19.845 3.73 20.145 6.86 ;
      RECT 22.98 4.055 23.325 4.785 ;
      RECT 19.74 3.31 20.07 4.04 ;
      RECT 22.62 3.15 23.35 3.48 ;
      RECT 93.455 7.205 93.835 12.465 ;
      RECT 87.14 3.31 87.47 4.04 ;
      RECT 85.94 4.175 86.27 4.905 ;
      RECT 85.1 3.15 85.83 3.48 ;
      RECT 82.7 3.15 83.03 3.88 ;
      RECT 78.195 7.205 78.575 12.465 ;
      RECT 71.88 3.31 72.21 4.04 ;
      RECT 70.68 4.175 71.01 4.905 ;
      RECT 69.84 3.15 70.57 3.48 ;
      RECT 67.44 3.15 67.77 3.88 ;
      RECT 62.935 7.205 63.315 12.465 ;
      RECT 56.62 3.31 56.95 4.04 ;
      RECT 55.42 4.175 55.75 4.905 ;
      RECT 54.58 3.15 55.31 3.48 ;
      RECT 52.18 3.15 52.51 3.88 ;
      RECT 47.675 7.205 48.055 12.465 ;
      RECT 41.36 3.31 41.69 4.04 ;
      RECT 40.16 4.175 40.49 4.905 ;
      RECT 39.32 3.15 40.05 3.48 ;
      RECT 36.92 3.15 37.25 3.88 ;
      RECT 32.415 7.205 32.795 12.465 ;
      RECT 26.1 3.31 26.43 4.04 ;
      RECT 24.9 4.175 25.23 4.905 ;
      RECT 24.06 3.15 24.79 3.48 ;
      RECT 21.66 3.15 21.99 3.88 ;
    LAYER via2 ;
      RECT 93.545 7.295 93.745 7.495 ;
      RECT 87.205 3.775 87.405 3.975 ;
      RECT 86.005 4.335 86.205 4.535 ;
      RECT 85.165 3.215 85.365 3.415 ;
      RECT 85.125 9.43 85.325 9.63 ;
      RECT 84.085 4.12 84.285 4.32 ;
      RECT 83.725 3.215 83.925 3.415 ;
      RECT 82.765 3.215 82.965 3.415 ;
      RECT 80.845 3.775 81.045 3.975 ;
      RECT 78.285 7.295 78.485 7.495 ;
      RECT 71.945 3.775 72.145 3.975 ;
      RECT 70.745 4.335 70.945 4.535 ;
      RECT 69.905 3.215 70.105 3.415 ;
      RECT 69.865 9.43 70.065 9.63 ;
      RECT 68.825 4.12 69.025 4.32 ;
      RECT 68.465 3.215 68.665 3.415 ;
      RECT 67.505 3.215 67.705 3.415 ;
      RECT 65.585 3.775 65.785 3.975 ;
      RECT 63.025 7.295 63.225 7.495 ;
      RECT 56.685 3.775 56.885 3.975 ;
      RECT 55.485 4.335 55.685 4.535 ;
      RECT 54.645 3.215 54.845 3.415 ;
      RECT 54.605 9.43 54.805 9.63 ;
      RECT 53.565 4.12 53.765 4.32 ;
      RECT 53.205 3.215 53.405 3.415 ;
      RECT 52.245 3.215 52.445 3.415 ;
      RECT 50.325 3.775 50.525 3.975 ;
      RECT 47.765 7.295 47.965 7.495 ;
      RECT 41.425 3.775 41.625 3.975 ;
      RECT 40.225 4.335 40.425 4.535 ;
      RECT 39.385 3.215 39.585 3.415 ;
      RECT 39.345 9.43 39.545 9.63 ;
      RECT 38.305 4.12 38.505 4.32 ;
      RECT 37.945 3.215 38.145 3.415 ;
      RECT 36.985 3.215 37.185 3.415 ;
      RECT 35.065 3.775 35.265 3.975 ;
      RECT 32.505 7.295 32.705 7.495 ;
      RECT 26.165 3.775 26.365 3.975 ;
      RECT 24.965 4.335 25.165 4.535 ;
      RECT 24.125 3.215 24.325 3.415 ;
      RECT 24.085 9.43 24.285 9.63 ;
      RECT 23.045 4.12 23.245 4.32 ;
      RECT 22.685 3.215 22.885 3.415 ;
      RECT 21.725 3.215 21.925 3.415 ;
      RECT 19.805 3.775 20.005 3.975 ;
    LAYER met2 ;
      RECT 16.235 10.69 93.73 10.86 ;
      RECT 93.56 9.565 93.73 10.86 ;
      RECT 16.235 8.545 16.405 10.86 ;
      RECT 93.53 9.565 93.88 9.915 ;
      RECT 16.17 8.545 16.46 8.895 ;
      RECT 90.37 8.51 90.69 8.835 ;
      RECT 90.4 7.985 90.57 8.835 ;
      RECT 90.4 7.985 90.575 8.335 ;
      RECT 90.4 7.985 91.375 8.16 ;
      RECT 91.2 3.26 91.375 8.16 ;
      RECT 91.145 3.26 91.495 3.61 ;
      RECT 91.17 8.945 91.495 9.27 ;
      RECT 90.055 9.035 91.495 9.205 ;
      RECT 90.055 3.69 90.215 9.205 ;
      RECT 90.37 3.66 90.69 3.98 ;
      RECT 90.055 3.69 90.69 3.86 ;
      RECT 88.765 4 89.105 4.35 ;
      RECT 88.16 4.065 89.105 4.265 ;
      RECT 88.16 4.06 88.375 4.265 ;
      RECT 88.175 3.635 88.375 4.265 ;
      RECT 87.165 3.635 87.445 4.015 ;
      RECT 88.855 3.995 89.025 4.35 ;
      RECT 87.16 3.635 87.445 3.968 ;
      RECT 87.14 3.635 87.445 3.945 ;
      RECT 87.13 3.635 87.445 3.925 ;
      RECT 87.12 3.635 87.445 3.91 ;
      RECT 87.095 3.635 87.445 3.883 ;
      RECT 87.085 3.635 87.445 3.858 ;
      RECT 87.04 3.59 87.32 3.85 ;
      RECT 87.04 3.635 88.375 3.835 ;
      RECT 87.04 3.63 87.365 3.85 ;
      RECT 87.04 3.622 87.36 3.85 ;
      RECT 87.04 3.612 87.355 3.85 ;
      RECT 87.04 3.6 87.35 3.85 ;
      RECT 85.965 4.295 86.245 4.575 ;
      RECT 85.965 4.295 86.28 4.555 ;
      RECT 78.245 8.95 78.595 9.3 ;
      RECT 85.71 8.905 86.06 9.255 ;
      RECT 78.245 8.98 86.06 9.18 ;
      RECT 86 3.715 86.05 3.975 ;
      RECT 85.79 3.715 85.795 3.975 ;
      RECT 84.985 3.27 85.015 3.53 ;
      RECT 84.755 3.27 84.83 3.53 ;
      RECT 85.975 3.665 86 3.975 ;
      RECT 85.97 3.622 85.975 3.975 ;
      RECT 85.965 3.605 85.97 3.975 ;
      RECT 85.96 3.592 85.965 3.975 ;
      RECT 85.885 3.475 85.96 3.975 ;
      RECT 85.84 3.292 85.885 3.975 ;
      RECT 85.835 3.22 85.84 3.975 ;
      RECT 85.82 3.195 85.835 3.975 ;
      RECT 85.795 3.157 85.82 3.975 ;
      RECT 85.785 3.137 85.795 3.697 ;
      RECT 85.77 3.129 85.785 3.652 ;
      RECT 85.765 3.121 85.77 3.623 ;
      RECT 85.76 3.118 85.765 3.603 ;
      RECT 85.755 3.115 85.76 3.583 ;
      RECT 85.75 3.112 85.755 3.563 ;
      RECT 85.72 3.101 85.75 3.5 ;
      RECT 85.7 3.086 85.72 3.415 ;
      RECT 85.695 3.078 85.7 3.378 ;
      RECT 85.685 3.072 85.695 3.345 ;
      RECT 85.67 3.064 85.685 3.305 ;
      RECT 85.665 3.057 85.67 3.265 ;
      RECT 85.66 3.054 85.665 3.243 ;
      RECT 85.655 3.051 85.66 3.23 ;
      RECT 85.65 3.05 85.655 3.22 ;
      RECT 85.635 3.044 85.65 3.21 ;
      RECT 85.61 3.031 85.635 3.195 ;
      RECT 85.56 3.006 85.61 3.166 ;
      RECT 85.545 2.985 85.56 3.141 ;
      RECT 85.535 2.978 85.545 3.13 ;
      RECT 85.48 2.959 85.535 3.103 ;
      RECT 85.455 2.937 85.48 3.076 ;
      RECT 85.45 2.93 85.455 3.071 ;
      RECT 85.435 2.93 85.45 3.069 ;
      RECT 85.41 2.922 85.435 3.065 ;
      RECT 85.395 2.92 85.41 3.061 ;
      RECT 85.365 2.92 85.395 3.058 ;
      RECT 85.355 2.92 85.365 3.053 ;
      RECT 85.31 2.92 85.355 3.051 ;
      RECT 85.281 2.92 85.31 3.052 ;
      RECT 85.195 2.92 85.281 3.054 ;
      RECT 85.181 2.921 85.195 3.056 ;
      RECT 85.095 2.922 85.181 3.058 ;
      RECT 85.08 2.923 85.095 3.068 ;
      RECT 85.075 2.924 85.08 3.077 ;
      RECT 85.055 2.927 85.075 3.087 ;
      RECT 85.04 2.935 85.055 3.102 ;
      RECT 85.02 2.953 85.04 3.117 ;
      RECT 85.01 2.965 85.02 3.14 ;
      RECT 85 2.974 85.01 3.17 ;
      RECT 84.985 2.986 85 3.215 ;
      RECT 84.93 3.019 84.985 3.53 ;
      RECT 84.925 3.047 84.93 3.53 ;
      RECT 84.905 3.062 84.925 3.53 ;
      RECT 84.87 3.122 84.905 3.53 ;
      RECT 84.868 3.172 84.87 3.53 ;
      RECT 84.865 3.18 84.868 3.53 ;
      RECT 84.855 3.195 84.865 3.53 ;
      RECT 84.85 3.207 84.855 3.53 ;
      RECT 84.84 3.232 84.85 3.53 ;
      RECT 84.83 3.26 84.84 3.53 ;
      RECT 82.735 4.765 82.785 5.025 ;
      RECT 85.645 4.315 85.705 4.575 ;
      RECT 85.63 4.315 85.645 4.585 ;
      RECT 85.611 4.315 85.63 4.618 ;
      RECT 85.525 4.315 85.611 4.743 ;
      RECT 85.445 4.315 85.525 4.925 ;
      RECT 85.44 4.552 85.445 5.01 ;
      RECT 85.415 4.622 85.44 5.038 ;
      RECT 85.41 4.692 85.415 5.065 ;
      RECT 85.39 4.764 85.41 5.087 ;
      RECT 85.385 4.831 85.39 5.11 ;
      RECT 85.375 4.86 85.385 5.125 ;
      RECT 85.365 4.882 85.375 5.142 ;
      RECT 85.36 4.892 85.365 5.153 ;
      RECT 85.355 4.9 85.36 5.161 ;
      RECT 85.345 4.908 85.355 5.173 ;
      RECT 85.34 4.92 85.345 5.183 ;
      RECT 85.335 4.928 85.34 5.188 ;
      RECT 85.315 4.946 85.335 5.198 ;
      RECT 85.31 4.963 85.315 5.205 ;
      RECT 85.305 4.971 85.31 5.206 ;
      RECT 85.3 4.982 85.305 5.208 ;
      RECT 85.26 5.02 85.3 5.218 ;
      RECT 85.255 5.055 85.26 5.229 ;
      RECT 85.25 5.06 85.255 5.232 ;
      RECT 85.225 5.07 85.25 5.239 ;
      RECT 85.215 5.084 85.225 5.248 ;
      RECT 85.195 5.096 85.215 5.251 ;
      RECT 85.145 5.115 85.195 5.255 ;
      RECT 85.1 5.13 85.145 5.26 ;
      RECT 85.035 5.133 85.1 5.266 ;
      RECT 85.02 5.131 85.035 5.273 ;
      RECT 84.99 5.13 85.02 5.273 ;
      RECT 84.951 5.129 84.99 5.269 ;
      RECT 84.865 5.126 84.951 5.265 ;
      RECT 84.848 5.124 84.865 5.262 ;
      RECT 84.762 5.122 84.848 5.259 ;
      RECT 84.676 5.119 84.762 5.253 ;
      RECT 84.59 5.115 84.676 5.248 ;
      RECT 84.512 5.112 84.59 5.244 ;
      RECT 84.426 5.109 84.512 5.242 ;
      RECT 84.34 5.106 84.426 5.239 ;
      RECT 84.282 5.104 84.34 5.236 ;
      RECT 84.196 5.101 84.282 5.234 ;
      RECT 84.11 5.097 84.196 5.232 ;
      RECT 84.024 5.094 84.11 5.229 ;
      RECT 83.938 5.09 84.024 5.227 ;
      RECT 83.852 5.086 83.938 5.224 ;
      RECT 83.766 5.083 83.852 5.222 ;
      RECT 83.68 5.079 83.766 5.219 ;
      RECT 83.594 5.076 83.68 5.217 ;
      RECT 83.508 5.072 83.594 5.214 ;
      RECT 83.422 5.069 83.508 5.212 ;
      RECT 83.336 5.065 83.422 5.209 ;
      RECT 83.25 5.062 83.336 5.207 ;
      RECT 83.24 5.06 83.25 5.203 ;
      RECT 83.235 5.06 83.24 5.201 ;
      RECT 83.195 5.055 83.235 5.195 ;
      RECT 83.181 5.046 83.195 5.188 ;
      RECT 83.095 5.016 83.181 5.173 ;
      RECT 83.075 4.982 83.095 5.158 ;
      RECT 83.005 4.951 83.075 5.145 ;
      RECT 83 4.926 83.005 5.134 ;
      RECT 82.995 4.92 83 5.132 ;
      RECT 82.926 4.765 82.995 5.12 ;
      RECT 82.84 4.765 82.926 5.094 ;
      RECT 82.815 4.765 82.84 5.073 ;
      RECT 82.81 4.765 82.815 5.063 ;
      RECT 82.805 4.765 82.81 5.055 ;
      RECT 82.785 4.765 82.805 5.038 ;
      RECT 85.205 3.335 85.465 3.595 ;
      RECT 85.19 3.335 85.465 3.498 ;
      RECT 85.16 3.335 85.465 3.473 ;
      RECT 85.125 3.175 85.405 3.455 ;
      RECT 85.095 4.665 85.155 4.925 ;
      RECT 84.12 3.355 84.175 3.615 ;
      RECT 85.055 4.622 85.095 4.925 ;
      RECT 85.026 4.543 85.055 4.925 ;
      RECT 84.94 4.415 85.026 4.925 ;
      RECT 84.92 4.295 84.94 4.925 ;
      RECT 84.895 4.246 84.92 4.925 ;
      RECT 84.89 4.211 84.895 4.775 ;
      RECT 84.86 4.171 84.89 4.713 ;
      RECT 84.835 4.108 84.86 4.628 ;
      RECT 84.825 4.07 84.835 4.565 ;
      RECT 84.81 4.045 84.825 4.526 ;
      RECT 84.767 4.003 84.81 4.432 ;
      RECT 84.765 3.976 84.767 4.359 ;
      RECT 84.76 3.971 84.765 4.35 ;
      RECT 84.755 3.964 84.76 4.325 ;
      RECT 84.75 3.958 84.755 4.31 ;
      RECT 84.745 3.952 84.75 4.298 ;
      RECT 84.735 3.943 84.745 4.28 ;
      RECT 84.73 3.934 84.735 4.258 ;
      RECT 84.705 3.915 84.73 4.208 ;
      RECT 84.7 3.896 84.705 4.158 ;
      RECT 84.685 3.882 84.7 4.118 ;
      RECT 84.68 3.868 84.685 4.085 ;
      RECT 84.675 3.861 84.68 4.078 ;
      RECT 84.66 3.848 84.675 4.07 ;
      RECT 84.615 3.81 84.66 4.043 ;
      RECT 84.585 3.763 84.615 4.008 ;
      RECT 84.565 3.732 84.585 3.985 ;
      RECT 84.485 3.665 84.565 3.938 ;
      RECT 84.455 3.595 84.485 3.885 ;
      RECT 84.45 3.572 84.455 3.868 ;
      RECT 84.42 3.55 84.45 3.853 ;
      RECT 84.39 3.509 84.42 3.825 ;
      RECT 84.385 3.484 84.39 3.81 ;
      RECT 84.38 3.478 84.385 3.803 ;
      RECT 84.37 3.355 84.38 3.795 ;
      RECT 84.36 3.355 84.37 3.788 ;
      RECT 84.355 3.355 84.36 3.78 ;
      RECT 84.335 3.355 84.355 3.768 ;
      RECT 84.285 3.355 84.335 3.738 ;
      RECT 84.23 3.355 84.285 3.688 ;
      RECT 84.2 3.355 84.23 3.648 ;
      RECT 84.175 3.355 84.2 3.625 ;
      RECT 84.045 4.08 84.325 4.36 ;
      RECT 84.01 3.995 84.27 4.255 ;
      RECT 84.01 4.077 84.28 4.255 ;
      RECT 82.21 3.45 82.215 3.935 ;
      RECT 82.1 3.635 82.105 3.935 ;
      RECT 82.01 3.675 82.075 3.935 ;
      RECT 83.685 3.175 83.775 3.805 ;
      RECT 83.65 3.225 83.655 3.805 ;
      RECT 83.595 3.25 83.605 3.805 ;
      RECT 83.55 3.25 83.56 3.805 ;
      RECT 83.92 3.175 83.965 3.455 ;
      RECT 82.77 2.905 82.97 3.045 ;
      RECT 83.886 3.175 83.92 3.467 ;
      RECT 83.8 3.175 83.886 3.507 ;
      RECT 83.785 3.175 83.8 3.548 ;
      RECT 83.78 3.175 83.785 3.568 ;
      RECT 83.775 3.175 83.78 3.588 ;
      RECT 83.655 3.217 83.685 3.805 ;
      RECT 83.605 3.237 83.65 3.805 ;
      RECT 83.59 3.252 83.595 3.805 ;
      RECT 83.56 3.252 83.59 3.805 ;
      RECT 83.515 3.237 83.55 3.805 ;
      RECT 83.51 3.225 83.515 3.585 ;
      RECT 83.505 3.222 83.51 3.565 ;
      RECT 83.49 3.212 83.505 3.518 ;
      RECT 83.485 3.205 83.49 3.481 ;
      RECT 83.48 3.202 83.485 3.464 ;
      RECT 83.465 3.192 83.48 3.42 ;
      RECT 83.46 3.183 83.465 3.38 ;
      RECT 83.455 3.179 83.46 3.365 ;
      RECT 83.445 3.173 83.455 3.348 ;
      RECT 83.405 3.154 83.445 3.323 ;
      RECT 83.4 3.136 83.405 3.303 ;
      RECT 83.39 3.13 83.4 3.298 ;
      RECT 83.36 3.114 83.39 3.285 ;
      RECT 83.345 3.096 83.36 3.268 ;
      RECT 83.33 3.084 83.345 3.255 ;
      RECT 83.325 3.076 83.33 3.248 ;
      RECT 83.295 3.062 83.325 3.235 ;
      RECT 83.29 3.047 83.295 3.223 ;
      RECT 83.28 3.041 83.29 3.215 ;
      RECT 83.26 3.029 83.28 3.203 ;
      RECT 83.25 3.017 83.26 3.19 ;
      RECT 83.22 3.001 83.25 3.175 ;
      RECT 83.2 2.981 83.22 3.158 ;
      RECT 83.195 2.971 83.2 3.148 ;
      RECT 83.17 2.959 83.195 3.135 ;
      RECT 83.165 2.947 83.17 3.123 ;
      RECT 83.16 2.942 83.165 3.119 ;
      RECT 83.145 2.935 83.16 3.111 ;
      RECT 83.135 2.922 83.145 3.101 ;
      RECT 83.13 2.92 83.135 3.095 ;
      RECT 83.105 2.913 83.13 3.084 ;
      RECT 83.1 2.906 83.105 3.073 ;
      RECT 83.075 2.905 83.1 3.06 ;
      RECT 83.056 2.905 83.075 3.05 ;
      RECT 82.97 2.905 83.056 3.047 ;
      RECT 82.74 2.905 82.77 3.05 ;
      RECT 82.7 2.912 82.74 3.063 ;
      RECT 82.675 2.922 82.7 3.076 ;
      RECT 82.66 2.931 82.675 3.086 ;
      RECT 82.63 2.936 82.66 3.105 ;
      RECT 82.625 2.942 82.63 3.123 ;
      RECT 82.605 2.952 82.625 3.138 ;
      RECT 82.595 2.965 82.605 3.158 ;
      RECT 82.58 2.977 82.595 3.175 ;
      RECT 82.575 2.987 82.58 3.185 ;
      RECT 82.57 2.992 82.575 3.19 ;
      RECT 82.56 3 82.57 3.203 ;
      RECT 82.51 3.032 82.56 3.24 ;
      RECT 82.495 3.067 82.51 3.281 ;
      RECT 82.49 3.077 82.495 3.296 ;
      RECT 82.485 3.082 82.49 3.303 ;
      RECT 82.46 3.098 82.485 3.323 ;
      RECT 82.445 3.119 82.46 3.348 ;
      RECT 82.42 3.14 82.445 3.373 ;
      RECT 82.41 3.159 82.42 3.396 ;
      RECT 82.385 3.177 82.41 3.419 ;
      RECT 82.37 3.197 82.385 3.443 ;
      RECT 82.365 3.207 82.37 3.455 ;
      RECT 82.35 3.219 82.365 3.475 ;
      RECT 82.34 3.234 82.35 3.515 ;
      RECT 82.335 3.242 82.34 3.543 ;
      RECT 82.325 3.252 82.335 3.563 ;
      RECT 82.32 3.265 82.325 3.588 ;
      RECT 82.315 3.278 82.32 3.608 ;
      RECT 82.31 3.284 82.315 3.63 ;
      RECT 82.3 3.293 82.31 3.65 ;
      RECT 82.295 3.313 82.3 3.673 ;
      RECT 82.29 3.319 82.295 3.693 ;
      RECT 82.285 3.326 82.29 3.715 ;
      RECT 82.28 3.337 82.285 3.728 ;
      RECT 82.27 3.347 82.28 3.753 ;
      RECT 82.25 3.372 82.27 3.935 ;
      RECT 82.22 3.412 82.25 3.935 ;
      RECT 82.215 3.442 82.22 3.935 ;
      RECT 82.19 3.47 82.21 3.935 ;
      RECT 82.16 3.515 82.19 3.935 ;
      RECT 82.155 3.542 82.16 3.935 ;
      RECT 82.135 3.56 82.155 3.935 ;
      RECT 82.125 3.585 82.135 3.935 ;
      RECT 82.12 3.597 82.125 3.935 ;
      RECT 82.105 3.62 82.12 3.935 ;
      RECT 82.085 3.647 82.1 3.935 ;
      RECT 82.075 3.67 82.085 3.935 ;
      RECT 83.865 4.555 83.945 4.815 ;
      RECT 83.1 3.775 83.17 4.035 ;
      RECT 83.831 4.522 83.865 4.815 ;
      RECT 83.745 4.425 83.831 4.815 ;
      RECT 83.725 4.337 83.745 4.815 ;
      RECT 83.715 4.307 83.725 4.815 ;
      RECT 83.705 4.287 83.715 4.815 ;
      RECT 83.685 4.274 83.705 4.815 ;
      RECT 83.67 4.264 83.685 4.643 ;
      RECT 83.665 4.257 83.67 4.598 ;
      RECT 83.655 4.251 83.665 4.588 ;
      RECT 83.645 4.243 83.655 4.57 ;
      RECT 83.64 4.237 83.645 4.558 ;
      RECT 83.63 4.232 83.64 4.545 ;
      RECT 83.61 4.222 83.63 4.518 ;
      RECT 83.57 4.201 83.61 4.47 ;
      RECT 83.555 4.182 83.57 4.428 ;
      RECT 83.53 4.168 83.555 4.398 ;
      RECT 83.52 4.156 83.53 4.365 ;
      RECT 83.515 4.151 83.52 4.355 ;
      RECT 83.485 4.137 83.515 4.335 ;
      RECT 83.475 4.121 83.485 4.308 ;
      RECT 83.47 4.116 83.475 4.298 ;
      RECT 83.445 4.107 83.47 4.278 ;
      RECT 83.435 4.095 83.445 4.258 ;
      RECT 83.365 4.063 83.435 4.233 ;
      RECT 83.36 4.032 83.365 4.21 ;
      RECT 83.311 3.775 83.36 4.193 ;
      RECT 83.225 3.775 83.311 4.152 ;
      RECT 83.17 3.775 83.225 4.08 ;
      RECT 83.26 4.56 83.42 4.82 ;
      RECT 82.785 3.175 82.835 3.86 ;
      RECT 82.575 3.6 82.61 3.86 ;
      RECT 82.89 3.175 82.895 3.635 ;
      RECT 82.98 3.175 83.005 3.455 ;
      RECT 83.255 4.557 83.26 4.82 ;
      RECT 83.22 4.545 83.255 4.82 ;
      RECT 83.16 4.518 83.22 4.82 ;
      RECT 83.155 4.501 83.16 4.674 ;
      RECT 83.15 4.498 83.155 4.661 ;
      RECT 83.13 4.491 83.15 4.648 ;
      RECT 83.095 4.474 83.13 4.63 ;
      RECT 83.055 4.453 83.095 4.61 ;
      RECT 83.05 4.441 83.055 4.598 ;
      RECT 83.01 4.427 83.05 4.584 ;
      RECT 82.99 4.41 83.01 4.566 ;
      RECT 82.98 4.402 82.99 4.558 ;
      RECT 82.965 3.175 82.98 3.473 ;
      RECT 82.95 4.392 82.98 4.545 ;
      RECT 82.935 3.175 82.965 3.518 ;
      RECT 82.94 4.382 82.95 4.532 ;
      RECT 82.91 4.367 82.94 4.519 ;
      RECT 82.895 3.175 82.935 3.585 ;
      RECT 82.895 4.335 82.91 4.505 ;
      RECT 82.89 4.307 82.895 4.499 ;
      RECT 82.885 3.175 82.89 3.64 ;
      RECT 82.875 4.277 82.89 4.493 ;
      RECT 82.88 3.175 82.885 3.653 ;
      RECT 82.87 3.175 82.88 3.673 ;
      RECT 82.835 4.19 82.875 4.478 ;
      RECT 82.835 3.175 82.87 3.713 ;
      RECT 82.83 4.122 82.835 4.466 ;
      RECT 82.815 4.077 82.83 4.461 ;
      RECT 82.81 4.015 82.815 4.456 ;
      RECT 82.785 3.922 82.81 4.449 ;
      RECT 82.78 3.175 82.785 4.441 ;
      RECT 82.765 3.175 82.78 4.428 ;
      RECT 82.745 3.175 82.765 4.385 ;
      RECT 82.735 3.175 82.745 4.335 ;
      RECT 82.73 3.175 82.735 4.308 ;
      RECT 82.725 3.175 82.73 4.286 ;
      RECT 82.72 3.401 82.725 4.269 ;
      RECT 82.715 3.423 82.72 4.247 ;
      RECT 82.71 3.465 82.715 4.23 ;
      RECT 82.68 3.515 82.71 4.174 ;
      RECT 82.675 3.542 82.68 4.116 ;
      RECT 82.66 3.56 82.675 4.08 ;
      RECT 82.655 3.578 82.66 4.044 ;
      RECT 82.649 3.585 82.655 4.025 ;
      RECT 82.645 3.592 82.649 4.008 ;
      RECT 82.64 3.597 82.645 3.977 ;
      RECT 82.63 3.6 82.64 3.952 ;
      RECT 82.62 3.6 82.63 3.918 ;
      RECT 82.615 3.6 82.62 3.895 ;
      RECT 82.61 3.6 82.615 3.875 ;
      RECT 81.23 4.765 81.49 5.025 ;
      RECT 81.25 4.692 81.43 5.025 ;
      RECT 81.25 4.435 81.425 5.025 ;
      RECT 81.25 4.227 81.415 5.025 ;
      RECT 81.255 4.145 81.415 5.025 ;
      RECT 81.255 3.91 81.405 5.025 ;
      RECT 81.255 3.757 81.4 5.025 ;
      RECT 81.26 3.742 81.4 5.025 ;
      RECT 81.31 3.457 81.4 5.025 ;
      RECT 81.265 3.692 81.4 5.025 ;
      RECT 81.295 3.51 81.4 5.025 ;
      RECT 81.28 3.622 81.4 5.025 ;
      RECT 81.285 3.58 81.4 5.025 ;
      RECT 81.28 3.622 81.415 3.685 ;
      RECT 81.315 3.21 81.42 3.63 ;
      RECT 81.315 3.21 81.435 3.613 ;
      RECT 81.315 3.21 81.47 3.575 ;
      RECT 81.31 3.457 81.52 3.508 ;
      RECT 81.315 3.21 81.575 3.47 ;
      RECT 80.575 3.915 80.835 4.175 ;
      RECT 80.575 3.915 80.845 4.133 ;
      RECT 80.575 3.915 80.931 4.104 ;
      RECT 80.575 3.915 81 4.056 ;
      RECT 80.575 3.915 81.035 4.025 ;
      RECT 80.805 3.735 81.085 4.015 ;
      RECT 80.64 3.9 81.085 4.015 ;
      RECT 80.73 3.777 80.835 4.175 ;
      RECT 80.66 3.84 81.085 4.015 ;
      RECT 75.11 8.51 75.43 8.835 ;
      RECT 75.14 7.985 75.31 8.835 ;
      RECT 75.14 7.985 75.315 8.335 ;
      RECT 75.14 7.985 76.115 8.16 ;
      RECT 75.94 3.26 76.115 8.16 ;
      RECT 75.885 3.26 76.235 3.61 ;
      RECT 75.91 8.945 76.235 9.27 ;
      RECT 74.795 9.035 76.235 9.205 ;
      RECT 74.795 3.69 74.955 9.205 ;
      RECT 75.11 3.66 75.43 3.98 ;
      RECT 74.795 3.69 75.43 3.86 ;
      RECT 73.505 4 73.845 4.35 ;
      RECT 72.9 4.065 73.845 4.265 ;
      RECT 72.9 4.06 73.115 4.265 ;
      RECT 72.915 3.635 73.115 4.265 ;
      RECT 71.905 3.635 72.185 4.015 ;
      RECT 73.595 3.995 73.765 4.35 ;
      RECT 71.9 3.635 72.185 3.968 ;
      RECT 71.88 3.635 72.185 3.945 ;
      RECT 71.87 3.635 72.185 3.925 ;
      RECT 71.86 3.635 72.185 3.91 ;
      RECT 71.835 3.635 72.185 3.883 ;
      RECT 71.825 3.635 72.185 3.858 ;
      RECT 71.78 3.59 72.06 3.85 ;
      RECT 71.78 3.635 73.115 3.835 ;
      RECT 71.78 3.63 72.105 3.85 ;
      RECT 71.78 3.622 72.1 3.85 ;
      RECT 71.78 3.612 72.095 3.85 ;
      RECT 71.78 3.6 72.09 3.85 ;
      RECT 70.705 4.295 70.985 4.575 ;
      RECT 70.705 4.295 71.02 4.555 ;
      RECT 62.985 8.95 63.335 9.3 ;
      RECT 70.45 8.905 70.8 9.255 ;
      RECT 62.985 8.98 70.8 9.18 ;
      RECT 70.74 3.715 70.79 3.975 ;
      RECT 70.53 3.715 70.535 3.975 ;
      RECT 69.725 3.27 69.755 3.53 ;
      RECT 69.495 3.27 69.57 3.53 ;
      RECT 70.715 3.665 70.74 3.975 ;
      RECT 70.71 3.622 70.715 3.975 ;
      RECT 70.705 3.605 70.71 3.975 ;
      RECT 70.7 3.592 70.705 3.975 ;
      RECT 70.625 3.475 70.7 3.975 ;
      RECT 70.58 3.292 70.625 3.975 ;
      RECT 70.575 3.22 70.58 3.975 ;
      RECT 70.56 3.195 70.575 3.975 ;
      RECT 70.535 3.157 70.56 3.975 ;
      RECT 70.525 3.137 70.535 3.697 ;
      RECT 70.51 3.129 70.525 3.652 ;
      RECT 70.505 3.121 70.51 3.623 ;
      RECT 70.5 3.118 70.505 3.603 ;
      RECT 70.495 3.115 70.5 3.583 ;
      RECT 70.49 3.112 70.495 3.563 ;
      RECT 70.46 3.101 70.49 3.5 ;
      RECT 70.44 3.086 70.46 3.415 ;
      RECT 70.435 3.078 70.44 3.378 ;
      RECT 70.425 3.072 70.435 3.345 ;
      RECT 70.41 3.064 70.425 3.305 ;
      RECT 70.405 3.057 70.41 3.265 ;
      RECT 70.4 3.054 70.405 3.243 ;
      RECT 70.395 3.051 70.4 3.23 ;
      RECT 70.39 3.05 70.395 3.22 ;
      RECT 70.375 3.044 70.39 3.21 ;
      RECT 70.35 3.031 70.375 3.195 ;
      RECT 70.3 3.006 70.35 3.166 ;
      RECT 70.285 2.985 70.3 3.141 ;
      RECT 70.275 2.978 70.285 3.13 ;
      RECT 70.22 2.959 70.275 3.103 ;
      RECT 70.195 2.937 70.22 3.076 ;
      RECT 70.19 2.93 70.195 3.071 ;
      RECT 70.175 2.93 70.19 3.069 ;
      RECT 70.15 2.922 70.175 3.065 ;
      RECT 70.135 2.92 70.15 3.061 ;
      RECT 70.105 2.92 70.135 3.058 ;
      RECT 70.095 2.92 70.105 3.053 ;
      RECT 70.05 2.92 70.095 3.051 ;
      RECT 70.021 2.92 70.05 3.052 ;
      RECT 69.935 2.92 70.021 3.054 ;
      RECT 69.921 2.921 69.935 3.056 ;
      RECT 69.835 2.922 69.921 3.058 ;
      RECT 69.82 2.923 69.835 3.068 ;
      RECT 69.815 2.924 69.82 3.077 ;
      RECT 69.795 2.927 69.815 3.087 ;
      RECT 69.78 2.935 69.795 3.102 ;
      RECT 69.76 2.953 69.78 3.117 ;
      RECT 69.75 2.965 69.76 3.14 ;
      RECT 69.74 2.974 69.75 3.17 ;
      RECT 69.725 2.986 69.74 3.215 ;
      RECT 69.67 3.019 69.725 3.53 ;
      RECT 69.665 3.047 69.67 3.53 ;
      RECT 69.645 3.062 69.665 3.53 ;
      RECT 69.61 3.122 69.645 3.53 ;
      RECT 69.608 3.172 69.61 3.53 ;
      RECT 69.605 3.18 69.608 3.53 ;
      RECT 69.595 3.195 69.605 3.53 ;
      RECT 69.59 3.207 69.595 3.53 ;
      RECT 69.58 3.232 69.59 3.53 ;
      RECT 69.57 3.26 69.58 3.53 ;
      RECT 67.475 4.765 67.525 5.025 ;
      RECT 70.385 4.315 70.445 4.575 ;
      RECT 70.37 4.315 70.385 4.585 ;
      RECT 70.351 4.315 70.37 4.618 ;
      RECT 70.265 4.315 70.351 4.743 ;
      RECT 70.185 4.315 70.265 4.925 ;
      RECT 70.18 4.552 70.185 5.01 ;
      RECT 70.155 4.622 70.18 5.038 ;
      RECT 70.15 4.692 70.155 5.065 ;
      RECT 70.13 4.764 70.15 5.087 ;
      RECT 70.125 4.831 70.13 5.11 ;
      RECT 70.115 4.86 70.125 5.125 ;
      RECT 70.105 4.882 70.115 5.142 ;
      RECT 70.1 4.892 70.105 5.153 ;
      RECT 70.095 4.9 70.1 5.161 ;
      RECT 70.085 4.908 70.095 5.173 ;
      RECT 70.08 4.92 70.085 5.183 ;
      RECT 70.075 4.928 70.08 5.188 ;
      RECT 70.055 4.946 70.075 5.198 ;
      RECT 70.05 4.963 70.055 5.205 ;
      RECT 70.045 4.971 70.05 5.206 ;
      RECT 70.04 4.982 70.045 5.208 ;
      RECT 70 5.02 70.04 5.218 ;
      RECT 69.995 5.055 70 5.229 ;
      RECT 69.99 5.06 69.995 5.232 ;
      RECT 69.965 5.07 69.99 5.239 ;
      RECT 69.955 5.084 69.965 5.248 ;
      RECT 69.935 5.096 69.955 5.251 ;
      RECT 69.885 5.115 69.935 5.255 ;
      RECT 69.84 5.13 69.885 5.26 ;
      RECT 69.775 5.133 69.84 5.266 ;
      RECT 69.76 5.131 69.775 5.273 ;
      RECT 69.73 5.13 69.76 5.273 ;
      RECT 69.691 5.129 69.73 5.269 ;
      RECT 69.605 5.126 69.691 5.265 ;
      RECT 69.588 5.124 69.605 5.262 ;
      RECT 69.502 5.122 69.588 5.259 ;
      RECT 69.416 5.119 69.502 5.253 ;
      RECT 69.33 5.115 69.416 5.248 ;
      RECT 69.252 5.112 69.33 5.244 ;
      RECT 69.166 5.109 69.252 5.242 ;
      RECT 69.08 5.106 69.166 5.239 ;
      RECT 69.022 5.104 69.08 5.236 ;
      RECT 68.936 5.101 69.022 5.234 ;
      RECT 68.85 5.097 68.936 5.232 ;
      RECT 68.764 5.094 68.85 5.229 ;
      RECT 68.678 5.09 68.764 5.227 ;
      RECT 68.592 5.086 68.678 5.224 ;
      RECT 68.506 5.083 68.592 5.222 ;
      RECT 68.42 5.079 68.506 5.219 ;
      RECT 68.334 5.076 68.42 5.217 ;
      RECT 68.248 5.072 68.334 5.214 ;
      RECT 68.162 5.069 68.248 5.212 ;
      RECT 68.076 5.065 68.162 5.209 ;
      RECT 67.99 5.062 68.076 5.207 ;
      RECT 67.98 5.06 67.99 5.203 ;
      RECT 67.975 5.06 67.98 5.201 ;
      RECT 67.935 5.055 67.975 5.195 ;
      RECT 67.921 5.046 67.935 5.188 ;
      RECT 67.835 5.016 67.921 5.173 ;
      RECT 67.815 4.982 67.835 5.158 ;
      RECT 67.745 4.951 67.815 5.145 ;
      RECT 67.74 4.926 67.745 5.134 ;
      RECT 67.735 4.92 67.74 5.132 ;
      RECT 67.666 4.765 67.735 5.12 ;
      RECT 67.58 4.765 67.666 5.094 ;
      RECT 67.555 4.765 67.58 5.073 ;
      RECT 67.55 4.765 67.555 5.063 ;
      RECT 67.545 4.765 67.55 5.055 ;
      RECT 67.525 4.765 67.545 5.038 ;
      RECT 69.945 3.335 70.205 3.595 ;
      RECT 69.93 3.335 70.205 3.498 ;
      RECT 69.9 3.335 70.205 3.473 ;
      RECT 69.865 3.175 70.145 3.455 ;
      RECT 69.835 4.665 69.895 4.925 ;
      RECT 68.86 3.355 68.915 3.615 ;
      RECT 69.795 4.622 69.835 4.925 ;
      RECT 69.766 4.543 69.795 4.925 ;
      RECT 69.68 4.415 69.766 4.925 ;
      RECT 69.66 4.295 69.68 4.925 ;
      RECT 69.635 4.246 69.66 4.925 ;
      RECT 69.63 4.211 69.635 4.775 ;
      RECT 69.6 4.171 69.63 4.713 ;
      RECT 69.575 4.108 69.6 4.628 ;
      RECT 69.565 4.07 69.575 4.565 ;
      RECT 69.55 4.045 69.565 4.526 ;
      RECT 69.507 4.003 69.55 4.432 ;
      RECT 69.505 3.976 69.507 4.359 ;
      RECT 69.5 3.971 69.505 4.35 ;
      RECT 69.495 3.964 69.5 4.325 ;
      RECT 69.49 3.958 69.495 4.31 ;
      RECT 69.485 3.952 69.49 4.298 ;
      RECT 69.475 3.943 69.485 4.28 ;
      RECT 69.47 3.934 69.475 4.258 ;
      RECT 69.445 3.915 69.47 4.208 ;
      RECT 69.44 3.896 69.445 4.158 ;
      RECT 69.425 3.882 69.44 4.118 ;
      RECT 69.42 3.868 69.425 4.085 ;
      RECT 69.415 3.861 69.42 4.078 ;
      RECT 69.4 3.848 69.415 4.07 ;
      RECT 69.355 3.81 69.4 4.043 ;
      RECT 69.325 3.763 69.355 4.008 ;
      RECT 69.305 3.732 69.325 3.985 ;
      RECT 69.225 3.665 69.305 3.938 ;
      RECT 69.195 3.595 69.225 3.885 ;
      RECT 69.19 3.572 69.195 3.868 ;
      RECT 69.16 3.55 69.19 3.853 ;
      RECT 69.13 3.509 69.16 3.825 ;
      RECT 69.125 3.484 69.13 3.81 ;
      RECT 69.12 3.478 69.125 3.803 ;
      RECT 69.11 3.355 69.12 3.795 ;
      RECT 69.1 3.355 69.11 3.788 ;
      RECT 69.095 3.355 69.1 3.78 ;
      RECT 69.075 3.355 69.095 3.768 ;
      RECT 69.025 3.355 69.075 3.738 ;
      RECT 68.97 3.355 69.025 3.688 ;
      RECT 68.94 3.355 68.97 3.648 ;
      RECT 68.915 3.355 68.94 3.625 ;
      RECT 68.785 4.08 69.065 4.36 ;
      RECT 68.75 3.995 69.01 4.255 ;
      RECT 68.75 4.077 69.02 4.255 ;
      RECT 66.95 3.45 66.955 3.935 ;
      RECT 66.84 3.635 66.845 3.935 ;
      RECT 66.75 3.675 66.815 3.935 ;
      RECT 68.425 3.175 68.515 3.805 ;
      RECT 68.39 3.225 68.395 3.805 ;
      RECT 68.335 3.25 68.345 3.805 ;
      RECT 68.29 3.25 68.3 3.805 ;
      RECT 68.66 3.175 68.705 3.455 ;
      RECT 67.51 2.905 67.71 3.045 ;
      RECT 68.626 3.175 68.66 3.467 ;
      RECT 68.54 3.175 68.626 3.507 ;
      RECT 68.525 3.175 68.54 3.548 ;
      RECT 68.52 3.175 68.525 3.568 ;
      RECT 68.515 3.175 68.52 3.588 ;
      RECT 68.395 3.217 68.425 3.805 ;
      RECT 68.345 3.237 68.39 3.805 ;
      RECT 68.33 3.252 68.335 3.805 ;
      RECT 68.3 3.252 68.33 3.805 ;
      RECT 68.255 3.237 68.29 3.805 ;
      RECT 68.25 3.225 68.255 3.585 ;
      RECT 68.245 3.222 68.25 3.565 ;
      RECT 68.23 3.212 68.245 3.518 ;
      RECT 68.225 3.205 68.23 3.481 ;
      RECT 68.22 3.202 68.225 3.464 ;
      RECT 68.205 3.192 68.22 3.42 ;
      RECT 68.2 3.183 68.205 3.38 ;
      RECT 68.195 3.179 68.2 3.365 ;
      RECT 68.185 3.173 68.195 3.348 ;
      RECT 68.145 3.154 68.185 3.323 ;
      RECT 68.14 3.136 68.145 3.303 ;
      RECT 68.13 3.13 68.14 3.298 ;
      RECT 68.1 3.114 68.13 3.285 ;
      RECT 68.085 3.096 68.1 3.268 ;
      RECT 68.07 3.084 68.085 3.255 ;
      RECT 68.065 3.076 68.07 3.248 ;
      RECT 68.035 3.062 68.065 3.235 ;
      RECT 68.03 3.047 68.035 3.223 ;
      RECT 68.02 3.041 68.03 3.215 ;
      RECT 68 3.029 68.02 3.203 ;
      RECT 67.99 3.017 68 3.19 ;
      RECT 67.96 3.001 67.99 3.175 ;
      RECT 67.94 2.981 67.96 3.158 ;
      RECT 67.935 2.971 67.94 3.148 ;
      RECT 67.91 2.959 67.935 3.135 ;
      RECT 67.905 2.947 67.91 3.123 ;
      RECT 67.9 2.942 67.905 3.119 ;
      RECT 67.885 2.935 67.9 3.111 ;
      RECT 67.875 2.922 67.885 3.101 ;
      RECT 67.87 2.92 67.875 3.095 ;
      RECT 67.845 2.913 67.87 3.084 ;
      RECT 67.84 2.906 67.845 3.073 ;
      RECT 67.815 2.905 67.84 3.06 ;
      RECT 67.796 2.905 67.815 3.05 ;
      RECT 67.71 2.905 67.796 3.047 ;
      RECT 67.48 2.905 67.51 3.05 ;
      RECT 67.44 2.912 67.48 3.063 ;
      RECT 67.415 2.922 67.44 3.076 ;
      RECT 67.4 2.931 67.415 3.086 ;
      RECT 67.37 2.936 67.4 3.105 ;
      RECT 67.365 2.942 67.37 3.123 ;
      RECT 67.345 2.952 67.365 3.138 ;
      RECT 67.335 2.965 67.345 3.158 ;
      RECT 67.32 2.977 67.335 3.175 ;
      RECT 67.315 2.987 67.32 3.185 ;
      RECT 67.31 2.992 67.315 3.19 ;
      RECT 67.3 3 67.31 3.203 ;
      RECT 67.25 3.032 67.3 3.24 ;
      RECT 67.235 3.067 67.25 3.281 ;
      RECT 67.23 3.077 67.235 3.296 ;
      RECT 67.225 3.082 67.23 3.303 ;
      RECT 67.2 3.098 67.225 3.323 ;
      RECT 67.185 3.119 67.2 3.348 ;
      RECT 67.16 3.14 67.185 3.373 ;
      RECT 67.15 3.159 67.16 3.396 ;
      RECT 67.125 3.177 67.15 3.419 ;
      RECT 67.11 3.197 67.125 3.443 ;
      RECT 67.105 3.207 67.11 3.455 ;
      RECT 67.09 3.219 67.105 3.475 ;
      RECT 67.08 3.234 67.09 3.515 ;
      RECT 67.075 3.242 67.08 3.543 ;
      RECT 67.065 3.252 67.075 3.563 ;
      RECT 67.06 3.265 67.065 3.588 ;
      RECT 67.055 3.278 67.06 3.608 ;
      RECT 67.05 3.284 67.055 3.63 ;
      RECT 67.04 3.293 67.05 3.65 ;
      RECT 67.035 3.313 67.04 3.673 ;
      RECT 67.03 3.319 67.035 3.693 ;
      RECT 67.025 3.326 67.03 3.715 ;
      RECT 67.02 3.337 67.025 3.728 ;
      RECT 67.01 3.347 67.02 3.753 ;
      RECT 66.99 3.372 67.01 3.935 ;
      RECT 66.96 3.412 66.99 3.935 ;
      RECT 66.955 3.442 66.96 3.935 ;
      RECT 66.93 3.47 66.95 3.935 ;
      RECT 66.9 3.515 66.93 3.935 ;
      RECT 66.895 3.542 66.9 3.935 ;
      RECT 66.875 3.56 66.895 3.935 ;
      RECT 66.865 3.585 66.875 3.935 ;
      RECT 66.86 3.597 66.865 3.935 ;
      RECT 66.845 3.62 66.86 3.935 ;
      RECT 66.825 3.647 66.84 3.935 ;
      RECT 66.815 3.67 66.825 3.935 ;
      RECT 68.605 4.555 68.685 4.815 ;
      RECT 67.84 3.775 67.91 4.035 ;
      RECT 68.571 4.522 68.605 4.815 ;
      RECT 68.485 4.425 68.571 4.815 ;
      RECT 68.465 4.337 68.485 4.815 ;
      RECT 68.455 4.307 68.465 4.815 ;
      RECT 68.445 4.287 68.455 4.815 ;
      RECT 68.425 4.274 68.445 4.815 ;
      RECT 68.41 4.264 68.425 4.643 ;
      RECT 68.405 4.257 68.41 4.598 ;
      RECT 68.395 4.251 68.405 4.588 ;
      RECT 68.385 4.243 68.395 4.57 ;
      RECT 68.38 4.237 68.385 4.558 ;
      RECT 68.37 4.232 68.38 4.545 ;
      RECT 68.35 4.222 68.37 4.518 ;
      RECT 68.31 4.201 68.35 4.47 ;
      RECT 68.295 4.182 68.31 4.428 ;
      RECT 68.27 4.168 68.295 4.398 ;
      RECT 68.26 4.156 68.27 4.365 ;
      RECT 68.255 4.151 68.26 4.355 ;
      RECT 68.225 4.137 68.255 4.335 ;
      RECT 68.215 4.121 68.225 4.308 ;
      RECT 68.21 4.116 68.215 4.298 ;
      RECT 68.185 4.107 68.21 4.278 ;
      RECT 68.175 4.095 68.185 4.258 ;
      RECT 68.105 4.063 68.175 4.233 ;
      RECT 68.1 4.032 68.105 4.21 ;
      RECT 68.051 3.775 68.1 4.193 ;
      RECT 67.965 3.775 68.051 4.152 ;
      RECT 67.91 3.775 67.965 4.08 ;
      RECT 68 4.56 68.16 4.82 ;
      RECT 67.525 3.175 67.575 3.86 ;
      RECT 67.315 3.6 67.35 3.86 ;
      RECT 67.63 3.175 67.635 3.635 ;
      RECT 67.72 3.175 67.745 3.455 ;
      RECT 67.995 4.557 68 4.82 ;
      RECT 67.96 4.545 67.995 4.82 ;
      RECT 67.9 4.518 67.96 4.82 ;
      RECT 67.895 4.501 67.9 4.674 ;
      RECT 67.89 4.498 67.895 4.661 ;
      RECT 67.87 4.491 67.89 4.648 ;
      RECT 67.835 4.474 67.87 4.63 ;
      RECT 67.795 4.453 67.835 4.61 ;
      RECT 67.79 4.441 67.795 4.598 ;
      RECT 67.75 4.427 67.79 4.584 ;
      RECT 67.73 4.41 67.75 4.566 ;
      RECT 67.72 4.402 67.73 4.558 ;
      RECT 67.705 3.175 67.72 3.473 ;
      RECT 67.69 4.392 67.72 4.545 ;
      RECT 67.675 3.175 67.705 3.518 ;
      RECT 67.68 4.382 67.69 4.532 ;
      RECT 67.65 4.367 67.68 4.519 ;
      RECT 67.635 3.175 67.675 3.585 ;
      RECT 67.635 4.335 67.65 4.505 ;
      RECT 67.63 4.307 67.635 4.499 ;
      RECT 67.625 3.175 67.63 3.64 ;
      RECT 67.615 4.277 67.63 4.493 ;
      RECT 67.62 3.175 67.625 3.653 ;
      RECT 67.61 3.175 67.62 3.673 ;
      RECT 67.575 4.19 67.615 4.478 ;
      RECT 67.575 3.175 67.61 3.713 ;
      RECT 67.57 4.122 67.575 4.466 ;
      RECT 67.555 4.077 67.57 4.461 ;
      RECT 67.55 4.015 67.555 4.456 ;
      RECT 67.525 3.922 67.55 4.449 ;
      RECT 67.52 3.175 67.525 4.441 ;
      RECT 67.505 3.175 67.52 4.428 ;
      RECT 67.485 3.175 67.505 4.385 ;
      RECT 67.475 3.175 67.485 4.335 ;
      RECT 67.47 3.175 67.475 4.308 ;
      RECT 67.465 3.175 67.47 4.286 ;
      RECT 67.46 3.401 67.465 4.269 ;
      RECT 67.455 3.423 67.46 4.247 ;
      RECT 67.45 3.465 67.455 4.23 ;
      RECT 67.42 3.515 67.45 4.174 ;
      RECT 67.415 3.542 67.42 4.116 ;
      RECT 67.4 3.56 67.415 4.08 ;
      RECT 67.395 3.578 67.4 4.044 ;
      RECT 67.389 3.585 67.395 4.025 ;
      RECT 67.385 3.592 67.389 4.008 ;
      RECT 67.38 3.597 67.385 3.977 ;
      RECT 67.37 3.6 67.38 3.952 ;
      RECT 67.36 3.6 67.37 3.918 ;
      RECT 67.355 3.6 67.36 3.895 ;
      RECT 67.35 3.6 67.355 3.875 ;
      RECT 65.97 4.765 66.23 5.025 ;
      RECT 65.99 4.692 66.17 5.025 ;
      RECT 65.99 4.435 66.165 5.025 ;
      RECT 65.99 4.227 66.155 5.025 ;
      RECT 65.995 4.145 66.155 5.025 ;
      RECT 65.995 3.91 66.145 5.025 ;
      RECT 65.995 3.757 66.14 5.025 ;
      RECT 66 3.742 66.14 5.025 ;
      RECT 66.05 3.457 66.14 5.025 ;
      RECT 66.005 3.692 66.14 5.025 ;
      RECT 66.035 3.51 66.14 5.025 ;
      RECT 66.02 3.622 66.14 5.025 ;
      RECT 66.025 3.58 66.14 5.025 ;
      RECT 66.02 3.622 66.155 3.685 ;
      RECT 66.055 3.21 66.16 3.63 ;
      RECT 66.055 3.21 66.175 3.613 ;
      RECT 66.055 3.21 66.21 3.575 ;
      RECT 66.05 3.457 66.26 3.508 ;
      RECT 66.055 3.21 66.315 3.47 ;
      RECT 65.315 3.915 65.575 4.175 ;
      RECT 65.315 3.915 65.585 4.133 ;
      RECT 65.315 3.915 65.671 4.104 ;
      RECT 65.315 3.915 65.74 4.056 ;
      RECT 65.315 3.915 65.775 4.025 ;
      RECT 65.545 3.735 65.825 4.015 ;
      RECT 65.38 3.9 65.825 4.015 ;
      RECT 65.47 3.777 65.575 4.175 ;
      RECT 65.4 3.84 65.825 4.015 ;
      RECT 59.85 8.51 60.17 8.835 ;
      RECT 59.88 7.985 60.05 8.835 ;
      RECT 59.88 7.985 60.055 8.335 ;
      RECT 59.88 7.985 60.855 8.16 ;
      RECT 60.68 3.26 60.855 8.16 ;
      RECT 60.625 3.26 60.975 3.61 ;
      RECT 60.65 8.945 60.975 9.27 ;
      RECT 59.535 9.035 60.975 9.205 ;
      RECT 59.535 3.69 59.695 9.205 ;
      RECT 59.85 3.66 60.17 3.98 ;
      RECT 59.535 3.69 60.17 3.86 ;
      RECT 58.245 4 58.585 4.35 ;
      RECT 57.64 4.065 58.585 4.265 ;
      RECT 57.64 4.06 57.855 4.265 ;
      RECT 57.655 3.635 57.855 4.265 ;
      RECT 56.645 3.635 56.925 4.015 ;
      RECT 58.335 3.995 58.505 4.35 ;
      RECT 56.64 3.635 56.925 3.968 ;
      RECT 56.62 3.635 56.925 3.945 ;
      RECT 56.61 3.635 56.925 3.925 ;
      RECT 56.6 3.635 56.925 3.91 ;
      RECT 56.575 3.635 56.925 3.883 ;
      RECT 56.565 3.635 56.925 3.858 ;
      RECT 56.52 3.59 56.8 3.85 ;
      RECT 56.52 3.635 57.855 3.835 ;
      RECT 56.52 3.63 56.845 3.85 ;
      RECT 56.52 3.622 56.84 3.85 ;
      RECT 56.52 3.612 56.835 3.85 ;
      RECT 56.52 3.6 56.83 3.85 ;
      RECT 55.445 4.295 55.725 4.575 ;
      RECT 55.445 4.295 55.76 4.555 ;
      RECT 47.77 8.95 48.12 9.3 ;
      RECT 55.19 8.905 55.54 9.255 ;
      RECT 47.77 8.98 55.54 9.18 ;
      RECT 55.48 3.715 55.53 3.975 ;
      RECT 55.27 3.715 55.275 3.975 ;
      RECT 54.465 3.27 54.495 3.53 ;
      RECT 54.235 3.27 54.31 3.53 ;
      RECT 55.455 3.665 55.48 3.975 ;
      RECT 55.45 3.622 55.455 3.975 ;
      RECT 55.445 3.605 55.45 3.975 ;
      RECT 55.44 3.592 55.445 3.975 ;
      RECT 55.365 3.475 55.44 3.975 ;
      RECT 55.32 3.292 55.365 3.975 ;
      RECT 55.315 3.22 55.32 3.975 ;
      RECT 55.3 3.195 55.315 3.975 ;
      RECT 55.275 3.157 55.3 3.975 ;
      RECT 55.265 3.137 55.275 3.697 ;
      RECT 55.25 3.129 55.265 3.652 ;
      RECT 55.245 3.121 55.25 3.623 ;
      RECT 55.24 3.118 55.245 3.603 ;
      RECT 55.235 3.115 55.24 3.583 ;
      RECT 55.23 3.112 55.235 3.563 ;
      RECT 55.2 3.101 55.23 3.5 ;
      RECT 55.18 3.086 55.2 3.415 ;
      RECT 55.175 3.078 55.18 3.378 ;
      RECT 55.165 3.072 55.175 3.345 ;
      RECT 55.15 3.064 55.165 3.305 ;
      RECT 55.145 3.057 55.15 3.265 ;
      RECT 55.14 3.054 55.145 3.243 ;
      RECT 55.135 3.051 55.14 3.23 ;
      RECT 55.13 3.05 55.135 3.22 ;
      RECT 55.115 3.044 55.13 3.21 ;
      RECT 55.09 3.031 55.115 3.195 ;
      RECT 55.04 3.006 55.09 3.166 ;
      RECT 55.025 2.985 55.04 3.141 ;
      RECT 55.015 2.978 55.025 3.13 ;
      RECT 54.96 2.959 55.015 3.103 ;
      RECT 54.935 2.937 54.96 3.076 ;
      RECT 54.93 2.93 54.935 3.071 ;
      RECT 54.915 2.93 54.93 3.069 ;
      RECT 54.89 2.922 54.915 3.065 ;
      RECT 54.875 2.92 54.89 3.061 ;
      RECT 54.845 2.92 54.875 3.058 ;
      RECT 54.835 2.92 54.845 3.053 ;
      RECT 54.79 2.92 54.835 3.051 ;
      RECT 54.761 2.92 54.79 3.052 ;
      RECT 54.675 2.92 54.761 3.054 ;
      RECT 54.661 2.921 54.675 3.056 ;
      RECT 54.575 2.922 54.661 3.058 ;
      RECT 54.56 2.923 54.575 3.068 ;
      RECT 54.555 2.924 54.56 3.077 ;
      RECT 54.535 2.927 54.555 3.087 ;
      RECT 54.52 2.935 54.535 3.102 ;
      RECT 54.5 2.953 54.52 3.117 ;
      RECT 54.49 2.965 54.5 3.14 ;
      RECT 54.48 2.974 54.49 3.17 ;
      RECT 54.465 2.986 54.48 3.215 ;
      RECT 54.41 3.019 54.465 3.53 ;
      RECT 54.405 3.047 54.41 3.53 ;
      RECT 54.385 3.062 54.405 3.53 ;
      RECT 54.35 3.122 54.385 3.53 ;
      RECT 54.348 3.172 54.35 3.53 ;
      RECT 54.345 3.18 54.348 3.53 ;
      RECT 54.335 3.195 54.345 3.53 ;
      RECT 54.33 3.207 54.335 3.53 ;
      RECT 54.32 3.232 54.33 3.53 ;
      RECT 54.31 3.26 54.32 3.53 ;
      RECT 52.215 4.765 52.265 5.025 ;
      RECT 55.125 4.315 55.185 4.575 ;
      RECT 55.11 4.315 55.125 4.585 ;
      RECT 55.091 4.315 55.11 4.618 ;
      RECT 55.005 4.315 55.091 4.743 ;
      RECT 54.925 4.315 55.005 4.925 ;
      RECT 54.92 4.552 54.925 5.01 ;
      RECT 54.895 4.622 54.92 5.038 ;
      RECT 54.89 4.692 54.895 5.065 ;
      RECT 54.87 4.764 54.89 5.087 ;
      RECT 54.865 4.831 54.87 5.11 ;
      RECT 54.855 4.86 54.865 5.125 ;
      RECT 54.845 4.882 54.855 5.142 ;
      RECT 54.84 4.892 54.845 5.153 ;
      RECT 54.835 4.9 54.84 5.161 ;
      RECT 54.825 4.908 54.835 5.173 ;
      RECT 54.82 4.92 54.825 5.183 ;
      RECT 54.815 4.928 54.82 5.188 ;
      RECT 54.795 4.946 54.815 5.198 ;
      RECT 54.79 4.963 54.795 5.205 ;
      RECT 54.785 4.971 54.79 5.206 ;
      RECT 54.78 4.982 54.785 5.208 ;
      RECT 54.74 5.02 54.78 5.218 ;
      RECT 54.735 5.055 54.74 5.229 ;
      RECT 54.73 5.06 54.735 5.232 ;
      RECT 54.705 5.07 54.73 5.239 ;
      RECT 54.695 5.084 54.705 5.248 ;
      RECT 54.675 5.096 54.695 5.251 ;
      RECT 54.625 5.115 54.675 5.255 ;
      RECT 54.58 5.13 54.625 5.26 ;
      RECT 54.515 5.133 54.58 5.266 ;
      RECT 54.5 5.131 54.515 5.273 ;
      RECT 54.47 5.13 54.5 5.273 ;
      RECT 54.431 5.129 54.47 5.269 ;
      RECT 54.345 5.126 54.431 5.265 ;
      RECT 54.328 5.124 54.345 5.262 ;
      RECT 54.242 5.122 54.328 5.259 ;
      RECT 54.156 5.119 54.242 5.253 ;
      RECT 54.07 5.115 54.156 5.248 ;
      RECT 53.992 5.112 54.07 5.244 ;
      RECT 53.906 5.109 53.992 5.242 ;
      RECT 53.82 5.106 53.906 5.239 ;
      RECT 53.762 5.104 53.82 5.236 ;
      RECT 53.676 5.101 53.762 5.234 ;
      RECT 53.59 5.097 53.676 5.232 ;
      RECT 53.504 5.094 53.59 5.229 ;
      RECT 53.418 5.09 53.504 5.227 ;
      RECT 53.332 5.086 53.418 5.224 ;
      RECT 53.246 5.083 53.332 5.222 ;
      RECT 53.16 5.079 53.246 5.219 ;
      RECT 53.074 5.076 53.16 5.217 ;
      RECT 52.988 5.072 53.074 5.214 ;
      RECT 52.902 5.069 52.988 5.212 ;
      RECT 52.816 5.065 52.902 5.209 ;
      RECT 52.73 5.062 52.816 5.207 ;
      RECT 52.72 5.06 52.73 5.203 ;
      RECT 52.715 5.06 52.72 5.201 ;
      RECT 52.675 5.055 52.715 5.195 ;
      RECT 52.661 5.046 52.675 5.188 ;
      RECT 52.575 5.016 52.661 5.173 ;
      RECT 52.555 4.982 52.575 5.158 ;
      RECT 52.485 4.951 52.555 5.145 ;
      RECT 52.48 4.926 52.485 5.134 ;
      RECT 52.475 4.92 52.48 5.132 ;
      RECT 52.406 4.765 52.475 5.12 ;
      RECT 52.32 4.765 52.406 5.094 ;
      RECT 52.295 4.765 52.32 5.073 ;
      RECT 52.29 4.765 52.295 5.063 ;
      RECT 52.285 4.765 52.29 5.055 ;
      RECT 52.265 4.765 52.285 5.038 ;
      RECT 54.685 3.335 54.945 3.595 ;
      RECT 54.67 3.335 54.945 3.498 ;
      RECT 54.64 3.335 54.945 3.473 ;
      RECT 54.605 3.175 54.885 3.455 ;
      RECT 54.575 4.665 54.635 4.925 ;
      RECT 53.6 3.355 53.655 3.615 ;
      RECT 54.535 4.622 54.575 4.925 ;
      RECT 54.506 4.543 54.535 4.925 ;
      RECT 54.42 4.415 54.506 4.925 ;
      RECT 54.4 4.295 54.42 4.925 ;
      RECT 54.375 4.246 54.4 4.925 ;
      RECT 54.37 4.211 54.375 4.775 ;
      RECT 54.34 4.171 54.37 4.713 ;
      RECT 54.315 4.108 54.34 4.628 ;
      RECT 54.305 4.07 54.315 4.565 ;
      RECT 54.29 4.045 54.305 4.526 ;
      RECT 54.247 4.003 54.29 4.432 ;
      RECT 54.245 3.976 54.247 4.359 ;
      RECT 54.24 3.971 54.245 4.35 ;
      RECT 54.235 3.964 54.24 4.325 ;
      RECT 54.23 3.958 54.235 4.31 ;
      RECT 54.225 3.952 54.23 4.298 ;
      RECT 54.215 3.943 54.225 4.28 ;
      RECT 54.21 3.934 54.215 4.258 ;
      RECT 54.185 3.915 54.21 4.208 ;
      RECT 54.18 3.896 54.185 4.158 ;
      RECT 54.165 3.882 54.18 4.118 ;
      RECT 54.16 3.868 54.165 4.085 ;
      RECT 54.155 3.861 54.16 4.078 ;
      RECT 54.14 3.848 54.155 4.07 ;
      RECT 54.095 3.81 54.14 4.043 ;
      RECT 54.065 3.763 54.095 4.008 ;
      RECT 54.045 3.732 54.065 3.985 ;
      RECT 53.965 3.665 54.045 3.938 ;
      RECT 53.935 3.595 53.965 3.885 ;
      RECT 53.93 3.572 53.935 3.868 ;
      RECT 53.9 3.55 53.93 3.853 ;
      RECT 53.87 3.509 53.9 3.825 ;
      RECT 53.865 3.484 53.87 3.81 ;
      RECT 53.86 3.478 53.865 3.803 ;
      RECT 53.85 3.355 53.86 3.795 ;
      RECT 53.84 3.355 53.85 3.788 ;
      RECT 53.835 3.355 53.84 3.78 ;
      RECT 53.815 3.355 53.835 3.768 ;
      RECT 53.765 3.355 53.815 3.738 ;
      RECT 53.71 3.355 53.765 3.688 ;
      RECT 53.68 3.355 53.71 3.648 ;
      RECT 53.655 3.355 53.68 3.625 ;
      RECT 53.525 4.08 53.805 4.36 ;
      RECT 53.49 3.995 53.75 4.255 ;
      RECT 53.49 4.077 53.76 4.255 ;
      RECT 51.69 3.45 51.695 3.935 ;
      RECT 51.58 3.635 51.585 3.935 ;
      RECT 51.49 3.675 51.555 3.935 ;
      RECT 53.165 3.175 53.255 3.805 ;
      RECT 53.13 3.225 53.135 3.805 ;
      RECT 53.075 3.25 53.085 3.805 ;
      RECT 53.03 3.25 53.04 3.805 ;
      RECT 53.4 3.175 53.445 3.455 ;
      RECT 52.25 2.905 52.45 3.045 ;
      RECT 53.366 3.175 53.4 3.467 ;
      RECT 53.28 3.175 53.366 3.507 ;
      RECT 53.265 3.175 53.28 3.548 ;
      RECT 53.26 3.175 53.265 3.568 ;
      RECT 53.255 3.175 53.26 3.588 ;
      RECT 53.135 3.217 53.165 3.805 ;
      RECT 53.085 3.237 53.13 3.805 ;
      RECT 53.07 3.252 53.075 3.805 ;
      RECT 53.04 3.252 53.07 3.805 ;
      RECT 52.995 3.237 53.03 3.805 ;
      RECT 52.99 3.225 52.995 3.585 ;
      RECT 52.985 3.222 52.99 3.565 ;
      RECT 52.97 3.212 52.985 3.518 ;
      RECT 52.965 3.205 52.97 3.481 ;
      RECT 52.96 3.202 52.965 3.464 ;
      RECT 52.945 3.192 52.96 3.42 ;
      RECT 52.94 3.183 52.945 3.38 ;
      RECT 52.935 3.179 52.94 3.365 ;
      RECT 52.925 3.173 52.935 3.348 ;
      RECT 52.885 3.154 52.925 3.323 ;
      RECT 52.88 3.136 52.885 3.303 ;
      RECT 52.87 3.13 52.88 3.298 ;
      RECT 52.84 3.114 52.87 3.285 ;
      RECT 52.825 3.096 52.84 3.268 ;
      RECT 52.81 3.084 52.825 3.255 ;
      RECT 52.805 3.076 52.81 3.248 ;
      RECT 52.775 3.062 52.805 3.235 ;
      RECT 52.77 3.047 52.775 3.223 ;
      RECT 52.76 3.041 52.77 3.215 ;
      RECT 52.74 3.029 52.76 3.203 ;
      RECT 52.73 3.017 52.74 3.19 ;
      RECT 52.7 3.001 52.73 3.175 ;
      RECT 52.68 2.981 52.7 3.158 ;
      RECT 52.675 2.971 52.68 3.148 ;
      RECT 52.65 2.959 52.675 3.135 ;
      RECT 52.645 2.947 52.65 3.123 ;
      RECT 52.64 2.942 52.645 3.119 ;
      RECT 52.625 2.935 52.64 3.111 ;
      RECT 52.615 2.922 52.625 3.101 ;
      RECT 52.61 2.92 52.615 3.095 ;
      RECT 52.585 2.913 52.61 3.084 ;
      RECT 52.58 2.906 52.585 3.073 ;
      RECT 52.555 2.905 52.58 3.06 ;
      RECT 52.536 2.905 52.555 3.05 ;
      RECT 52.45 2.905 52.536 3.047 ;
      RECT 52.22 2.905 52.25 3.05 ;
      RECT 52.18 2.912 52.22 3.063 ;
      RECT 52.155 2.922 52.18 3.076 ;
      RECT 52.14 2.931 52.155 3.086 ;
      RECT 52.11 2.936 52.14 3.105 ;
      RECT 52.105 2.942 52.11 3.123 ;
      RECT 52.085 2.952 52.105 3.138 ;
      RECT 52.075 2.965 52.085 3.158 ;
      RECT 52.06 2.977 52.075 3.175 ;
      RECT 52.055 2.987 52.06 3.185 ;
      RECT 52.05 2.992 52.055 3.19 ;
      RECT 52.04 3 52.05 3.203 ;
      RECT 51.99 3.032 52.04 3.24 ;
      RECT 51.975 3.067 51.99 3.281 ;
      RECT 51.97 3.077 51.975 3.296 ;
      RECT 51.965 3.082 51.97 3.303 ;
      RECT 51.94 3.098 51.965 3.323 ;
      RECT 51.925 3.119 51.94 3.348 ;
      RECT 51.9 3.14 51.925 3.373 ;
      RECT 51.89 3.159 51.9 3.396 ;
      RECT 51.865 3.177 51.89 3.419 ;
      RECT 51.85 3.197 51.865 3.443 ;
      RECT 51.845 3.207 51.85 3.455 ;
      RECT 51.83 3.219 51.845 3.475 ;
      RECT 51.82 3.234 51.83 3.515 ;
      RECT 51.815 3.242 51.82 3.543 ;
      RECT 51.805 3.252 51.815 3.563 ;
      RECT 51.8 3.265 51.805 3.588 ;
      RECT 51.795 3.278 51.8 3.608 ;
      RECT 51.79 3.284 51.795 3.63 ;
      RECT 51.78 3.293 51.79 3.65 ;
      RECT 51.775 3.313 51.78 3.673 ;
      RECT 51.77 3.319 51.775 3.693 ;
      RECT 51.765 3.326 51.77 3.715 ;
      RECT 51.76 3.337 51.765 3.728 ;
      RECT 51.75 3.347 51.76 3.753 ;
      RECT 51.73 3.372 51.75 3.935 ;
      RECT 51.7 3.412 51.73 3.935 ;
      RECT 51.695 3.442 51.7 3.935 ;
      RECT 51.67 3.47 51.69 3.935 ;
      RECT 51.64 3.515 51.67 3.935 ;
      RECT 51.635 3.542 51.64 3.935 ;
      RECT 51.615 3.56 51.635 3.935 ;
      RECT 51.605 3.585 51.615 3.935 ;
      RECT 51.6 3.597 51.605 3.935 ;
      RECT 51.585 3.62 51.6 3.935 ;
      RECT 51.565 3.647 51.58 3.935 ;
      RECT 51.555 3.67 51.565 3.935 ;
      RECT 53.345 4.555 53.425 4.815 ;
      RECT 52.58 3.775 52.65 4.035 ;
      RECT 53.311 4.522 53.345 4.815 ;
      RECT 53.225 4.425 53.311 4.815 ;
      RECT 53.205 4.337 53.225 4.815 ;
      RECT 53.195 4.307 53.205 4.815 ;
      RECT 53.185 4.287 53.195 4.815 ;
      RECT 53.165 4.274 53.185 4.815 ;
      RECT 53.15 4.264 53.165 4.643 ;
      RECT 53.145 4.257 53.15 4.598 ;
      RECT 53.135 4.251 53.145 4.588 ;
      RECT 53.125 4.243 53.135 4.57 ;
      RECT 53.12 4.237 53.125 4.558 ;
      RECT 53.11 4.232 53.12 4.545 ;
      RECT 53.09 4.222 53.11 4.518 ;
      RECT 53.05 4.201 53.09 4.47 ;
      RECT 53.035 4.182 53.05 4.428 ;
      RECT 53.01 4.168 53.035 4.398 ;
      RECT 53 4.156 53.01 4.365 ;
      RECT 52.995 4.151 53 4.355 ;
      RECT 52.965 4.137 52.995 4.335 ;
      RECT 52.955 4.121 52.965 4.308 ;
      RECT 52.95 4.116 52.955 4.298 ;
      RECT 52.925 4.107 52.95 4.278 ;
      RECT 52.915 4.095 52.925 4.258 ;
      RECT 52.845 4.063 52.915 4.233 ;
      RECT 52.84 4.032 52.845 4.21 ;
      RECT 52.791 3.775 52.84 4.193 ;
      RECT 52.705 3.775 52.791 4.152 ;
      RECT 52.65 3.775 52.705 4.08 ;
      RECT 52.74 4.56 52.9 4.82 ;
      RECT 52.265 3.175 52.315 3.86 ;
      RECT 52.055 3.6 52.09 3.86 ;
      RECT 52.37 3.175 52.375 3.635 ;
      RECT 52.46 3.175 52.485 3.455 ;
      RECT 52.735 4.557 52.74 4.82 ;
      RECT 52.7 4.545 52.735 4.82 ;
      RECT 52.64 4.518 52.7 4.82 ;
      RECT 52.635 4.501 52.64 4.674 ;
      RECT 52.63 4.498 52.635 4.661 ;
      RECT 52.61 4.491 52.63 4.648 ;
      RECT 52.575 4.474 52.61 4.63 ;
      RECT 52.535 4.453 52.575 4.61 ;
      RECT 52.53 4.441 52.535 4.598 ;
      RECT 52.49 4.427 52.53 4.584 ;
      RECT 52.47 4.41 52.49 4.566 ;
      RECT 52.46 4.402 52.47 4.558 ;
      RECT 52.445 3.175 52.46 3.473 ;
      RECT 52.43 4.392 52.46 4.545 ;
      RECT 52.415 3.175 52.445 3.518 ;
      RECT 52.42 4.382 52.43 4.532 ;
      RECT 52.39 4.367 52.42 4.519 ;
      RECT 52.375 3.175 52.415 3.585 ;
      RECT 52.375 4.335 52.39 4.505 ;
      RECT 52.37 4.307 52.375 4.499 ;
      RECT 52.365 3.175 52.37 3.64 ;
      RECT 52.355 4.277 52.37 4.493 ;
      RECT 52.36 3.175 52.365 3.653 ;
      RECT 52.35 3.175 52.36 3.673 ;
      RECT 52.315 4.19 52.355 4.478 ;
      RECT 52.315 3.175 52.35 3.713 ;
      RECT 52.31 4.122 52.315 4.466 ;
      RECT 52.295 4.077 52.31 4.461 ;
      RECT 52.29 4.015 52.295 4.456 ;
      RECT 52.265 3.922 52.29 4.449 ;
      RECT 52.26 3.175 52.265 4.441 ;
      RECT 52.245 3.175 52.26 4.428 ;
      RECT 52.225 3.175 52.245 4.385 ;
      RECT 52.215 3.175 52.225 4.335 ;
      RECT 52.21 3.175 52.215 4.308 ;
      RECT 52.205 3.175 52.21 4.286 ;
      RECT 52.2 3.401 52.205 4.269 ;
      RECT 52.195 3.423 52.2 4.247 ;
      RECT 52.19 3.465 52.195 4.23 ;
      RECT 52.16 3.515 52.19 4.174 ;
      RECT 52.155 3.542 52.16 4.116 ;
      RECT 52.14 3.56 52.155 4.08 ;
      RECT 52.135 3.578 52.14 4.044 ;
      RECT 52.129 3.585 52.135 4.025 ;
      RECT 52.125 3.592 52.129 4.008 ;
      RECT 52.12 3.597 52.125 3.977 ;
      RECT 52.11 3.6 52.12 3.952 ;
      RECT 52.1 3.6 52.11 3.918 ;
      RECT 52.095 3.6 52.1 3.895 ;
      RECT 52.09 3.6 52.095 3.875 ;
      RECT 50.71 4.765 50.97 5.025 ;
      RECT 50.73 4.692 50.91 5.025 ;
      RECT 50.73 4.435 50.905 5.025 ;
      RECT 50.73 4.227 50.895 5.025 ;
      RECT 50.735 4.145 50.895 5.025 ;
      RECT 50.735 3.91 50.885 5.025 ;
      RECT 50.735 3.757 50.88 5.025 ;
      RECT 50.74 3.742 50.88 5.025 ;
      RECT 50.79 3.457 50.88 5.025 ;
      RECT 50.745 3.692 50.88 5.025 ;
      RECT 50.775 3.51 50.88 5.025 ;
      RECT 50.76 3.622 50.88 5.025 ;
      RECT 50.765 3.58 50.88 5.025 ;
      RECT 50.76 3.622 50.895 3.685 ;
      RECT 50.795 3.21 50.9 3.63 ;
      RECT 50.795 3.21 50.915 3.613 ;
      RECT 50.795 3.21 50.95 3.575 ;
      RECT 50.79 3.457 51 3.508 ;
      RECT 50.795 3.21 51.055 3.47 ;
      RECT 50.055 3.915 50.315 4.175 ;
      RECT 50.055 3.915 50.325 4.133 ;
      RECT 50.055 3.915 50.411 4.104 ;
      RECT 50.055 3.915 50.48 4.056 ;
      RECT 50.055 3.915 50.515 4.025 ;
      RECT 50.285 3.735 50.565 4.015 ;
      RECT 50.12 3.9 50.565 4.015 ;
      RECT 50.21 3.777 50.315 4.175 ;
      RECT 50.14 3.84 50.565 4.015 ;
      RECT 44.59 8.51 44.91 8.835 ;
      RECT 44.62 7.985 44.79 8.835 ;
      RECT 44.62 7.985 44.795 8.335 ;
      RECT 44.62 7.985 45.595 8.16 ;
      RECT 45.42 3.26 45.595 8.16 ;
      RECT 45.365 3.26 45.715 3.61 ;
      RECT 45.39 8.945 45.715 9.27 ;
      RECT 44.275 9.035 45.715 9.205 ;
      RECT 44.275 3.69 44.435 9.205 ;
      RECT 44.59 3.66 44.91 3.98 ;
      RECT 44.275 3.69 44.91 3.86 ;
      RECT 42.985 4 43.325 4.35 ;
      RECT 42.38 4.065 43.325 4.265 ;
      RECT 42.38 4.06 42.595 4.265 ;
      RECT 42.395 3.635 42.595 4.265 ;
      RECT 41.385 3.635 41.665 4.015 ;
      RECT 43.075 3.995 43.245 4.35 ;
      RECT 41.38 3.635 41.665 3.968 ;
      RECT 41.36 3.635 41.665 3.945 ;
      RECT 41.35 3.635 41.665 3.925 ;
      RECT 41.34 3.635 41.665 3.91 ;
      RECT 41.315 3.635 41.665 3.883 ;
      RECT 41.305 3.635 41.665 3.858 ;
      RECT 41.26 3.59 41.54 3.85 ;
      RECT 41.26 3.635 42.595 3.835 ;
      RECT 41.26 3.63 41.585 3.85 ;
      RECT 41.26 3.622 41.58 3.85 ;
      RECT 41.26 3.612 41.575 3.85 ;
      RECT 41.26 3.6 41.57 3.85 ;
      RECT 40.185 4.295 40.465 4.575 ;
      RECT 40.185 4.295 40.5 4.555 ;
      RECT 32.51 8.95 32.86 9.3 ;
      RECT 39.93 8.905 40.28 9.255 ;
      RECT 32.51 8.98 40.28 9.18 ;
      RECT 40.22 3.715 40.27 3.975 ;
      RECT 40.01 3.715 40.015 3.975 ;
      RECT 39.205 3.27 39.235 3.53 ;
      RECT 38.975 3.27 39.05 3.53 ;
      RECT 40.195 3.665 40.22 3.975 ;
      RECT 40.19 3.622 40.195 3.975 ;
      RECT 40.185 3.605 40.19 3.975 ;
      RECT 40.18 3.592 40.185 3.975 ;
      RECT 40.105 3.475 40.18 3.975 ;
      RECT 40.06 3.292 40.105 3.975 ;
      RECT 40.055 3.22 40.06 3.975 ;
      RECT 40.04 3.195 40.055 3.975 ;
      RECT 40.015 3.157 40.04 3.975 ;
      RECT 40.005 3.137 40.015 3.697 ;
      RECT 39.99 3.129 40.005 3.652 ;
      RECT 39.985 3.121 39.99 3.623 ;
      RECT 39.98 3.118 39.985 3.603 ;
      RECT 39.975 3.115 39.98 3.583 ;
      RECT 39.97 3.112 39.975 3.563 ;
      RECT 39.94 3.101 39.97 3.5 ;
      RECT 39.92 3.086 39.94 3.415 ;
      RECT 39.915 3.078 39.92 3.378 ;
      RECT 39.905 3.072 39.915 3.345 ;
      RECT 39.89 3.064 39.905 3.305 ;
      RECT 39.885 3.057 39.89 3.265 ;
      RECT 39.88 3.054 39.885 3.243 ;
      RECT 39.875 3.051 39.88 3.23 ;
      RECT 39.87 3.05 39.875 3.22 ;
      RECT 39.855 3.044 39.87 3.21 ;
      RECT 39.83 3.031 39.855 3.195 ;
      RECT 39.78 3.006 39.83 3.166 ;
      RECT 39.765 2.985 39.78 3.141 ;
      RECT 39.755 2.978 39.765 3.13 ;
      RECT 39.7 2.959 39.755 3.103 ;
      RECT 39.675 2.937 39.7 3.076 ;
      RECT 39.67 2.93 39.675 3.071 ;
      RECT 39.655 2.93 39.67 3.069 ;
      RECT 39.63 2.922 39.655 3.065 ;
      RECT 39.615 2.92 39.63 3.061 ;
      RECT 39.585 2.92 39.615 3.058 ;
      RECT 39.575 2.92 39.585 3.053 ;
      RECT 39.53 2.92 39.575 3.051 ;
      RECT 39.501 2.92 39.53 3.052 ;
      RECT 39.415 2.92 39.501 3.054 ;
      RECT 39.401 2.921 39.415 3.056 ;
      RECT 39.315 2.922 39.401 3.058 ;
      RECT 39.3 2.923 39.315 3.068 ;
      RECT 39.295 2.924 39.3 3.077 ;
      RECT 39.275 2.927 39.295 3.087 ;
      RECT 39.26 2.935 39.275 3.102 ;
      RECT 39.24 2.953 39.26 3.117 ;
      RECT 39.23 2.965 39.24 3.14 ;
      RECT 39.22 2.974 39.23 3.17 ;
      RECT 39.205 2.986 39.22 3.215 ;
      RECT 39.15 3.019 39.205 3.53 ;
      RECT 39.145 3.047 39.15 3.53 ;
      RECT 39.125 3.062 39.145 3.53 ;
      RECT 39.09 3.122 39.125 3.53 ;
      RECT 39.088 3.172 39.09 3.53 ;
      RECT 39.085 3.18 39.088 3.53 ;
      RECT 39.075 3.195 39.085 3.53 ;
      RECT 39.07 3.207 39.075 3.53 ;
      RECT 39.06 3.232 39.07 3.53 ;
      RECT 39.05 3.26 39.06 3.53 ;
      RECT 36.955 4.765 37.005 5.025 ;
      RECT 39.865 4.315 39.925 4.575 ;
      RECT 39.85 4.315 39.865 4.585 ;
      RECT 39.831 4.315 39.85 4.618 ;
      RECT 39.745 4.315 39.831 4.743 ;
      RECT 39.665 4.315 39.745 4.925 ;
      RECT 39.66 4.552 39.665 5.01 ;
      RECT 39.635 4.622 39.66 5.038 ;
      RECT 39.63 4.692 39.635 5.065 ;
      RECT 39.61 4.764 39.63 5.087 ;
      RECT 39.605 4.831 39.61 5.11 ;
      RECT 39.595 4.86 39.605 5.125 ;
      RECT 39.585 4.882 39.595 5.142 ;
      RECT 39.58 4.892 39.585 5.153 ;
      RECT 39.575 4.9 39.58 5.161 ;
      RECT 39.565 4.908 39.575 5.173 ;
      RECT 39.56 4.92 39.565 5.183 ;
      RECT 39.555 4.928 39.56 5.188 ;
      RECT 39.535 4.946 39.555 5.198 ;
      RECT 39.53 4.963 39.535 5.205 ;
      RECT 39.525 4.971 39.53 5.206 ;
      RECT 39.52 4.982 39.525 5.208 ;
      RECT 39.48 5.02 39.52 5.218 ;
      RECT 39.475 5.055 39.48 5.229 ;
      RECT 39.47 5.06 39.475 5.232 ;
      RECT 39.445 5.07 39.47 5.239 ;
      RECT 39.435 5.084 39.445 5.248 ;
      RECT 39.415 5.096 39.435 5.251 ;
      RECT 39.365 5.115 39.415 5.255 ;
      RECT 39.32 5.13 39.365 5.26 ;
      RECT 39.255 5.133 39.32 5.266 ;
      RECT 39.24 5.131 39.255 5.273 ;
      RECT 39.21 5.13 39.24 5.273 ;
      RECT 39.171 5.129 39.21 5.269 ;
      RECT 39.085 5.126 39.171 5.265 ;
      RECT 39.068 5.124 39.085 5.262 ;
      RECT 38.982 5.122 39.068 5.259 ;
      RECT 38.896 5.119 38.982 5.253 ;
      RECT 38.81 5.115 38.896 5.248 ;
      RECT 38.732 5.112 38.81 5.244 ;
      RECT 38.646 5.109 38.732 5.242 ;
      RECT 38.56 5.106 38.646 5.239 ;
      RECT 38.502 5.104 38.56 5.236 ;
      RECT 38.416 5.101 38.502 5.234 ;
      RECT 38.33 5.097 38.416 5.232 ;
      RECT 38.244 5.094 38.33 5.229 ;
      RECT 38.158 5.09 38.244 5.227 ;
      RECT 38.072 5.086 38.158 5.224 ;
      RECT 37.986 5.083 38.072 5.222 ;
      RECT 37.9 5.079 37.986 5.219 ;
      RECT 37.814 5.076 37.9 5.217 ;
      RECT 37.728 5.072 37.814 5.214 ;
      RECT 37.642 5.069 37.728 5.212 ;
      RECT 37.556 5.065 37.642 5.209 ;
      RECT 37.47 5.062 37.556 5.207 ;
      RECT 37.46 5.06 37.47 5.203 ;
      RECT 37.455 5.06 37.46 5.201 ;
      RECT 37.415 5.055 37.455 5.195 ;
      RECT 37.401 5.046 37.415 5.188 ;
      RECT 37.315 5.016 37.401 5.173 ;
      RECT 37.295 4.982 37.315 5.158 ;
      RECT 37.225 4.951 37.295 5.145 ;
      RECT 37.22 4.926 37.225 5.134 ;
      RECT 37.215 4.92 37.22 5.132 ;
      RECT 37.146 4.765 37.215 5.12 ;
      RECT 37.06 4.765 37.146 5.094 ;
      RECT 37.035 4.765 37.06 5.073 ;
      RECT 37.03 4.765 37.035 5.063 ;
      RECT 37.025 4.765 37.03 5.055 ;
      RECT 37.005 4.765 37.025 5.038 ;
      RECT 39.425 3.335 39.685 3.595 ;
      RECT 39.41 3.335 39.685 3.498 ;
      RECT 39.38 3.335 39.685 3.473 ;
      RECT 39.345 3.175 39.625 3.455 ;
      RECT 39.315 4.665 39.375 4.925 ;
      RECT 38.34 3.355 38.395 3.615 ;
      RECT 39.275 4.622 39.315 4.925 ;
      RECT 39.246 4.543 39.275 4.925 ;
      RECT 39.16 4.415 39.246 4.925 ;
      RECT 39.14 4.295 39.16 4.925 ;
      RECT 39.115 4.246 39.14 4.925 ;
      RECT 39.11 4.211 39.115 4.775 ;
      RECT 39.08 4.171 39.11 4.713 ;
      RECT 39.055 4.108 39.08 4.628 ;
      RECT 39.045 4.07 39.055 4.565 ;
      RECT 39.03 4.045 39.045 4.526 ;
      RECT 38.987 4.003 39.03 4.432 ;
      RECT 38.985 3.976 38.987 4.359 ;
      RECT 38.98 3.971 38.985 4.35 ;
      RECT 38.975 3.964 38.98 4.325 ;
      RECT 38.97 3.958 38.975 4.31 ;
      RECT 38.965 3.952 38.97 4.298 ;
      RECT 38.955 3.943 38.965 4.28 ;
      RECT 38.95 3.934 38.955 4.258 ;
      RECT 38.925 3.915 38.95 4.208 ;
      RECT 38.92 3.896 38.925 4.158 ;
      RECT 38.905 3.882 38.92 4.118 ;
      RECT 38.9 3.868 38.905 4.085 ;
      RECT 38.895 3.861 38.9 4.078 ;
      RECT 38.88 3.848 38.895 4.07 ;
      RECT 38.835 3.81 38.88 4.043 ;
      RECT 38.805 3.763 38.835 4.008 ;
      RECT 38.785 3.732 38.805 3.985 ;
      RECT 38.705 3.665 38.785 3.938 ;
      RECT 38.675 3.595 38.705 3.885 ;
      RECT 38.67 3.572 38.675 3.868 ;
      RECT 38.64 3.55 38.67 3.853 ;
      RECT 38.61 3.509 38.64 3.825 ;
      RECT 38.605 3.484 38.61 3.81 ;
      RECT 38.6 3.478 38.605 3.803 ;
      RECT 38.59 3.355 38.6 3.795 ;
      RECT 38.58 3.355 38.59 3.788 ;
      RECT 38.575 3.355 38.58 3.78 ;
      RECT 38.555 3.355 38.575 3.768 ;
      RECT 38.505 3.355 38.555 3.738 ;
      RECT 38.45 3.355 38.505 3.688 ;
      RECT 38.42 3.355 38.45 3.648 ;
      RECT 38.395 3.355 38.42 3.625 ;
      RECT 38.265 4.08 38.545 4.36 ;
      RECT 38.23 3.995 38.49 4.255 ;
      RECT 38.23 4.077 38.5 4.255 ;
      RECT 36.43 3.45 36.435 3.935 ;
      RECT 36.32 3.635 36.325 3.935 ;
      RECT 36.23 3.675 36.295 3.935 ;
      RECT 37.905 3.175 37.995 3.805 ;
      RECT 37.87 3.225 37.875 3.805 ;
      RECT 37.815 3.25 37.825 3.805 ;
      RECT 37.77 3.25 37.78 3.805 ;
      RECT 38.14 3.175 38.185 3.455 ;
      RECT 36.99 2.905 37.19 3.045 ;
      RECT 38.106 3.175 38.14 3.467 ;
      RECT 38.02 3.175 38.106 3.507 ;
      RECT 38.005 3.175 38.02 3.548 ;
      RECT 38 3.175 38.005 3.568 ;
      RECT 37.995 3.175 38 3.588 ;
      RECT 37.875 3.217 37.905 3.805 ;
      RECT 37.825 3.237 37.87 3.805 ;
      RECT 37.81 3.252 37.815 3.805 ;
      RECT 37.78 3.252 37.81 3.805 ;
      RECT 37.735 3.237 37.77 3.805 ;
      RECT 37.73 3.225 37.735 3.585 ;
      RECT 37.725 3.222 37.73 3.565 ;
      RECT 37.71 3.212 37.725 3.518 ;
      RECT 37.705 3.205 37.71 3.481 ;
      RECT 37.7 3.202 37.705 3.464 ;
      RECT 37.685 3.192 37.7 3.42 ;
      RECT 37.68 3.183 37.685 3.38 ;
      RECT 37.675 3.179 37.68 3.365 ;
      RECT 37.665 3.173 37.675 3.348 ;
      RECT 37.625 3.154 37.665 3.323 ;
      RECT 37.62 3.136 37.625 3.303 ;
      RECT 37.61 3.13 37.62 3.298 ;
      RECT 37.58 3.114 37.61 3.285 ;
      RECT 37.565 3.096 37.58 3.268 ;
      RECT 37.55 3.084 37.565 3.255 ;
      RECT 37.545 3.076 37.55 3.248 ;
      RECT 37.515 3.062 37.545 3.235 ;
      RECT 37.51 3.047 37.515 3.223 ;
      RECT 37.5 3.041 37.51 3.215 ;
      RECT 37.48 3.029 37.5 3.203 ;
      RECT 37.47 3.017 37.48 3.19 ;
      RECT 37.44 3.001 37.47 3.175 ;
      RECT 37.42 2.981 37.44 3.158 ;
      RECT 37.415 2.971 37.42 3.148 ;
      RECT 37.39 2.959 37.415 3.135 ;
      RECT 37.385 2.947 37.39 3.123 ;
      RECT 37.38 2.942 37.385 3.119 ;
      RECT 37.365 2.935 37.38 3.111 ;
      RECT 37.355 2.922 37.365 3.101 ;
      RECT 37.35 2.92 37.355 3.095 ;
      RECT 37.325 2.913 37.35 3.084 ;
      RECT 37.32 2.906 37.325 3.073 ;
      RECT 37.295 2.905 37.32 3.06 ;
      RECT 37.276 2.905 37.295 3.05 ;
      RECT 37.19 2.905 37.276 3.047 ;
      RECT 36.96 2.905 36.99 3.05 ;
      RECT 36.92 2.912 36.96 3.063 ;
      RECT 36.895 2.922 36.92 3.076 ;
      RECT 36.88 2.931 36.895 3.086 ;
      RECT 36.85 2.936 36.88 3.105 ;
      RECT 36.845 2.942 36.85 3.123 ;
      RECT 36.825 2.952 36.845 3.138 ;
      RECT 36.815 2.965 36.825 3.158 ;
      RECT 36.8 2.977 36.815 3.175 ;
      RECT 36.795 2.987 36.8 3.185 ;
      RECT 36.79 2.992 36.795 3.19 ;
      RECT 36.78 3 36.79 3.203 ;
      RECT 36.73 3.032 36.78 3.24 ;
      RECT 36.715 3.067 36.73 3.281 ;
      RECT 36.71 3.077 36.715 3.296 ;
      RECT 36.705 3.082 36.71 3.303 ;
      RECT 36.68 3.098 36.705 3.323 ;
      RECT 36.665 3.119 36.68 3.348 ;
      RECT 36.64 3.14 36.665 3.373 ;
      RECT 36.63 3.159 36.64 3.396 ;
      RECT 36.605 3.177 36.63 3.419 ;
      RECT 36.59 3.197 36.605 3.443 ;
      RECT 36.585 3.207 36.59 3.455 ;
      RECT 36.57 3.219 36.585 3.475 ;
      RECT 36.56 3.234 36.57 3.515 ;
      RECT 36.555 3.242 36.56 3.543 ;
      RECT 36.545 3.252 36.555 3.563 ;
      RECT 36.54 3.265 36.545 3.588 ;
      RECT 36.535 3.278 36.54 3.608 ;
      RECT 36.53 3.284 36.535 3.63 ;
      RECT 36.52 3.293 36.53 3.65 ;
      RECT 36.515 3.313 36.52 3.673 ;
      RECT 36.51 3.319 36.515 3.693 ;
      RECT 36.505 3.326 36.51 3.715 ;
      RECT 36.5 3.337 36.505 3.728 ;
      RECT 36.49 3.347 36.5 3.753 ;
      RECT 36.47 3.372 36.49 3.935 ;
      RECT 36.44 3.412 36.47 3.935 ;
      RECT 36.435 3.442 36.44 3.935 ;
      RECT 36.41 3.47 36.43 3.935 ;
      RECT 36.38 3.515 36.41 3.935 ;
      RECT 36.375 3.542 36.38 3.935 ;
      RECT 36.355 3.56 36.375 3.935 ;
      RECT 36.345 3.585 36.355 3.935 ;
      RECT 36.34 3.597 36.345 3.935 ;
      RECT 36.325 3.62 36.34 3.935 ;
      RECT 36.305 3.647 36.32 3.935 ;
      RECT 36.295 3.67 36.305 3.935 ;
      RECT 38.085 4.555 38.165 4.815 ;
      RECT 37.32 3.775 37.39 4.035 ;
      RECT 38.051 4.522 38.085 4.815 ;
      RECT 37.965 4.425 38.051 4.815 ;
      RECT 37.945 4.337 37.965 4.815 ;
      RECT 37.935 4.307 37.945 4.815 ;
      RECT 37.925 4.287 37.935 4.815 ;
      RECT 37.905 4.274 37.925 4.815 ;
      RECT 37.89 4.264 37.905 4.643 ;
      RECT 37.885 4.257 37.89 4.598 ;
      RECT 37.875 4.251 37.885 4.588 ;
      RECT 37.865 4.243 37.875 4.57 ;
      RECT 37.86 4.237 37.865 4.558 ;
      RECT 37.85 4.232 37.86 4.545 ;
      RECT 37.83 4.222 37.85 4.518 ;
      RECT 37.79 4.201 37.83 4.47 ;
      RECT 37.775 4.182 37.79 4.428 ;
      RECT 37.75 4.168 37.775 4.398 ;
      RECT 37.74 4.156 37.75 4.365 ;
      RECT 37.735 4.151 37.74 4.355 ;
      RECT 37.705 4.137 37.735 4.335 ;
      RECT 37.695 4.121 37.705 4.308 ;
      RECT 37.69 4.116 37.695 4.298 ;
      RECT 37.665 4.107 37.69 4.278 ;
      RECT 37.655 4.095 37.665 4.258 ;
      RECT 37.585 4.063 37.655 4.233 ;
      RECT 37.58 4.032 37.585 4.21 ;
      RECT 37.531 3.775 37.58 4.193 ;
      RECT 37.445 3.775 37.531 4.152 ;
      RECT 37.39 3.775 37.445 4.08 ;
      RECT 37.48 4.56 37.64 4.82 ;
      RECT 37.005 3.175 37.055 3.86 ;
      RECT 36.795 3.6 36.83 3.86 ;
      RECT 37.11 3.175 37.115 3.635 ;
      RECT 37.2 3.175 37.225 3.455 ;
      RECT 37.475 4.557 37.48 4.82 ;
      RECT 37.44 4.545 37.475 4.82 ;
      RECT 37.38 4.518 37.44 4.82 ;
      RECT 37.375 4.501 37.38 4.674 ;
      RECT 37.37 4.498 37.375 4.661 ;
      RECT 37.35 4.491 37.37 4.648 ;
      RECT 37.315 4.474 37.35 4.63 ;
      RECT 37.275 4.453 37.315 4.61 ;
      RECT 37.27 4.441 37.275 4.598 ;
      RECT 37.23 4.427 37.27 4.584 ;
      RECT 37.21 4.41 37.23 4.566 ;
      RECT 37.2 4.402 37.21 4.558 ;
      RECT 37.185 3.175 37.2 3.473 ;
      RECT 37.17 4.392 37.2 4.545 ;
      RECT 37.155 3.175 37.185 3.518 ;
      RECT 37.16 4.382 37.17 4.532 ;
      RECT 37.13 4.367 37.16 4.519 ;
      RECT 37.115 3.175 37.155 3.585 ;
      RECT 37.115 4.335 37.13 4.505 ;
      RECT 37.11 4.307 37.115 4.499 ;
      RECT 37.105 3.175 37.11 3.64 ;
      RECT 37.095 4.277 37.11 4.493 ;
      RECT 37.1 3.175 37.105 3.653 ;
      RECT 37.09 3.175 37.1 3.673 ;
      RECT 37.055 4.19 37.095 4.478 ;
      RECT 37.055 3.175 37.09 3.713 ;
      RECT 37.05 4.122 37.055 4.466 ;
      RECT 37.035 4.077 37.05 4.461 ;
      RECT 37.03 4.015 37.035 4.456 ;
      RECT 37.005 3.922 37.03 4.449 ;
      RECT 37 3.175 37.005 4.441 ;
      RECT 36.985 3.175 37 4.428 ;
      RECT 36.965 3.175 36.985 4.385 ;
      RECT 36.955 3.175 36.965 4.335 ;
      RECT 36.95 3.175 36.955 4.308 ;
      RECT 36.945 3.175 36.95 4.286 ;
      RECT 36.94 3.401 36.945 4.269 ;
      RECT 36.935 3.423 36.94 4.247 ;
      RECT 36.93 3.465 36.935 4.23 ;
      RECT 36.9 3.515 36.93 4.174 ;
      RECT 36.895 3.542 36.9 4.116 ;
      RECT 36.88 3.56 36.895 4.08 ;
      RECT 36.875 3.578 36.88 4.044 ;
      RECT 36.869 3.585 36.875 4.025 ;
      RECT 36.865 3.592 36.869 4.008 ;
      RECT 36.86 3.597 36.865 3.977 ;
      RECT 36.85 3.6 36.86 3.952 ;
      RECT 36.84 3.6 36.85 3.918 ;
      RECT 36.835 3.6 36.84 3.895 ;
      RECT 36.83 3.6 36.835 3.875 ;
      RECT 35.45 4.765 35.71 5.025 ;
      RECT 35.47 4.692 35.65 5.025 ;
      RECT 35.47 4.435 35.645 5.025 ;
      RECT 35.47 4.227 35.635 5.025 ;
      RECT 35.475 4.145 35.635 5.025 ;
      RECT 35.475 3.91 35.625 5.025 ;
      RECT 35.475 3.757 35.62 5.025 ;
      RECT 35.48 3.742 35.62 5.025 ;
      RECT 35.53 3.457 35.62 5.025 ;
      RECT 35.485 3.692 35.62 5.025 ;
      RECT 35.515 3.51 35.62 5.025 ;
      RECT 35.5 3.622 35.62 5.025 ;
      RECT 35.505 3.58 35.62 5.025 ;
      RECT 35.5 3.622 35.635 3.685 ;
      RECT 35.535 3.21 35.64 3.63 ;
      RECT 35.535 3.21 35.655 3.613 ;
      RECT 35.535 3.21 35.69 3.575 ;
      RECT 35.53 3.457 35.74 3.508 ;
      RECT 35.535 3.21 35.795 3.47 ;
      RECT 34.795 3.915 35.055 4.175 ;
      RECT 34.795 3.915 35.065 4.133 ;
      RECT 34.795 3.915 35.151 4.104 ;
      RECT 34.795 3.915 35.22 4.056 ;
      RECT 34.795 3.915 35.255 4.025 ;
      RECT 35.025 3.735 35.305 4.015 ;
      RECT 34.86 3.9 35.305 4.015 ;
      RECT 34.95 3.777 35.055 4.175 ;
      RECT 34.88 3.84 35.305 4.015 ;
      RECT 29.33 8.51 29.65 8.835 ;
      RECT 29.36 7.985 29.53 8.835 ;
      RECT 29.36 7.985 29.535 8.335 ;
      RECT 29.36 7.985 30.335 8.16 ;
      RECT 30.16 3.26 30.335 8.16 ;
      RECT 30.105 3.26 30.455 3.61 ;
      RECT 30.13 8.945 30.455 9.27 ;
      RECT 29.015 9.035 30.455 9.205 ;
      RECT 29.015 3.69 29.175 9.205 ;
      RECT 29.33 3.66 29.65 3.98 ;
      RECT 29.015 3.69 29.65 3.86 ;
      RECT 27.725 4 28.065 4.35 ;
      RECT 27.12 4.065 28.065 4.265 ;
      RECT 27.12 4.06 27.335 4.265 ;
      RECT 27.135 3.635 27.335 4.265 ;
      RECT 26.125 3.635 26.405 4.015 ;
      RECT 27.815 3.995 27.985 4.35 ;
      RECT 26.12 3.635 26.405 3.968 ;
      RECT 26.1 3.635 26.405 3.945 ;
      RECT 26.09 3.635 26.405 3.925 ;
      RECT 26.08 3.635 26.405 3.91 ;
      RECT 26.055 3.635 26.405 3.883 ;
      RECT 26.045 3.635 26.405 3.858 ;
      RECT 26 3.59 26.28 3.85 ;
      RECT 26 3.635 27.335 3.835 ;
      RECT 26 3.63 26.325 3.85 ;
      RECT 26 3.622 26.32 3.85 ;
      RECT 26 3.612 26.315 3.85 ;
      RECT 26 3.6 26.31 3.85 ;
      RECT 24.925 4.295 25.205 4.575 ;
      RECT 24.925 4.295 25.24 4.555 ;
      RECT 16.545 9.285 16.835 9.635 ;
      RECT 16.545 9.345 17.875 9.515 ;
      RECT 17.705 8.975 17.875 9.515 ;
      RECT 24.67 8.895 25.02 9.245 ;
      RECT 17.705 8.975 25.02 9.145 ;
      RECT 24.96 3.715 25.01 3.975 ;
      RECT 24.75 3.715 24.755 3.975 ;
      RECT 23.945 3.27 23.975 3.53 ;
      RECT 23.715 3.27 23.79 3.53 ;
      RECT 24.935 3.665 24.96 3.975 ;
      RECT 24.93 3.622 24.935 3.975 ;
      RECT 24.925 3.605 24.93 3.975 ;
      RECT 24.92 3.592 24.925 3.975 ;
      RECT 24.845 3.475 24.92 3.975 ;
      RECT 24.8 3.292 24.845 3.975 ;
      RECT 24.795 3.22 24.8 3.975 ;
      RECT 24.78 3.195 24.795 3.975 ;
      RECT 24.755 3.157 24.78 3.975 ;
      RECT 24.745 3.137 24.755 3.697 ;
      RECT 24.73 3.129 24.745 3.652 ;
      RECT 24.725 3.121 24.73 3.623 ;
      RECT 24.72 3.118 24.725 3.603 ;
      RECT 24.715 3.115 24.72 3.583 ;
      RECT 24.71 3.112 24.715 3.563 ;
      RECT 24.68 3.101 24.71 3.5 ;
      RECT 24.66 3.086 24.68 3.415 ;
      RECT 24.655 3.078 24.66 3.378 ;
      RECT 24.645 3.072 24.655 3.345 ;
      RECT 24.63 3.064 24.645 3.305 ;
      RECT 24.625 3.057 24.63 3.265 ;
      RECT 24.62 3.054 24.625 3.243 ;
      RECT 24.615 3.051 24.62 3.23 ;
      RECT 24.61 3.05 24.615 3.22 ;
      RECT 24.595 3.044 24.61 3.21 ;
      RECT 24.57 3.031 24.595 3.195 ;
      RECT 24.52 3.006 24.57 3.166 ;
      RECT 24.505 2.985 24.52 3.141 ;
      RECT 24.495 2.978 24.505 3.13 ;
      RECT 24.44 2.959 24.495 3.103 ;
      RECT 24.415 2.937 24.44 3.076 ;
      RECT 24.41 2.93 24.415 3.071 ;
      RECT 24.395 2.93 24.41 3.069 ;
      RECT 24.37 2.922 24.395 3.065 ;
      RECT 24.355 2.92 24.37 3.061 ;
      RECT 24.325 2.92 24.355 3.058 ;
      RECT 24.315 2.92 24.325 3.053 ;
      RECT 24.27 2.92 24.315 3.051 ;
      RECT 24.241 2.92 24.27 3.052 ;
      RECT 24.155 2.92 24.241 3.054 ;
      RECT 24.141 2.921 24.155 3.056 ;
      RECT 24.055 2.922 24.141 3.058 ;
      RECT 24.04 2.923 24.055 3.068 ;
      RECT 24.035 2.924 24.04 3.077 ;
      RECT 24.015 2.927 24.035 3.087 ;
      RECT 24 2.935 24.015 3.102 ;
      RECT 23.98 2.953 24 3.117 ;
      RECT 23.97 2.965 23.98 3.14 ;
      RECT 23.96 2.974 23.97 3.17 ;
      RECT 23.945 2.986 23.96 3.215 ;
      RECT 23.89 3.019 23.945 3.53 ;
      RECT 23.885 3.047 23.89 3.53 ;
      RECT 23.865 3.062 23.885 3.53 ;
      RECT 23.83 3.122 23.865 3.53 ;
      RECT 23.828 3.172 23.83 3.53 ;
      RECT 23.825 3.18 23.828 3.53 ;
      RECT 23.815 3.195 23.825 3.53 ;
      RECT 23.81 3.207 23.815 3.53 ;
      RECT 23.8 3.232 23.81 3.53 ;
      RECT 23.79 3.26 23.8 3.53 ;
      RECT 21.695 4.765 21.745 5.025 ;
      RECT 24.605 4.315 24.665 4.575 ;
      RECT 24.59 4.315 24.605 4.585 ;
      RECT 24.571 4.315 24.59 4.618 ;
      RECT 24.485 4.315 24.571 4.743 ;
      RECT 24.405 4.315 24.485 4.925 ;
      RECT 24.4 4.552 24.405 5.01 ;
      RECT 24.375 4.622 24.4 5.038 ;
      RECT 24.37 4.692 24.375 5.065 ;
      RECT 24.35 4.764 24.37 5.087 ;
      RECT 24.345 4.831 24.35 5.11 ;
      RECT 24.335 4.86 24.345 5.125 ;
      RECT 24.325 4.882 24.335 5.142 ;
      RECT 24.32 4.892 24.325 5.153 ;
      RECT 24.315 4.9 24.32 5.161 ;
      RECT 24.305 4.908 24.315 5.173 ;
      RECT 24.3 4.92 24.305 5.183 ;
      RECT 24.295 4.928 24.3 5.188 ;
      RECT 24.275 4.946 24.295 5.198 ;
      RECT 24.27 4.963 24.275 5.205 ;
      RECT 24.265 4.971 24.27 5.206 ;
      RECT 24.26 4.982 24.265 5.208 ;
      RECT 24.22 5.02 24.26 5.218 ;
      RECT 24.215 5.055 24.22 5.229 ;
      RECT 24.21 5.06 24.215 5.232 ;
      RECT 24.185 5.07 24.21 5.239 ;
      RECT 24.175 5.084 24.185 5.248 ;
      RECT 24.155 5.096 24.175 5.251 ;
      RECT 24.105 5.115 24.155 5.255 ;
      RECT 24.06 5.13 24.105 5.26 ;
      RECT 23.995 5.133 24.06 5.266 ;
      RECT 23.98 5.131 23.995 5.273 ;
      RECT 23.95 5.13 23.98 5.273 ;
      RECT 23.911 5.129 23.95 5.269 ;
      RECT 23.825 5.126 23.911 5.265 ;
      RECT 23.808 5.124 23.825 5.262 ;
      RECT 23.722 5.122 23.808 5.259 ;
      RECT 23.636 5.119 23.722 5.253 ;
      RECT 23.55 5.115 23.636 5.248 ;
      RECT 23.472 5.112 23.55 5.244 ;
      RECT 23.386 5.109 23.472 5.242 ;
      RECT 23.3 5.106 23.386 5.239 ;
      RECT 23.242 5.104 23.3 5.236 ;
      RECT 23.156 5.101 23.242 5.234 ;
      RECT 23.07 5.097 23.156 5.232 ;
      RECT 22.984 5.094 23.07 5.229 ;
      RECT 22.898 5.09 22.984 5.227 ;
      RECT 22.812 5.086 22.898 5.224 ;
      RECT 22.726 5.083 22.812 5.222 ;
      RECT 22.64 5.079 22.726 5.219 ;
      RECT 22.554 5.076 22.64 5.217 ;
      RECT 22.468 5.072 22.554 5.214 ;
      RECT 22.382 5.069 22.468 5.212 ;
      RECT 22.296 5.065 22.382 5.209 ;
      RECT 22.21 5.062 22.296 5.207 ;
      RECT 22.2 5.06 22.21 5.203 ;
      RECT 22.195 5.06 22.2 5.201 ;
      RECT 22.155 5.055 22.195 5.195 ;
      RECT 22.141 5.046 22.155 5.188 ;
      RECT 22.055 5.016 22.141 5.173 ;
      RECT 22.035 4.982 22.055 5.158 ;
      RECT 21.965 4.951 22.035 5.145 ;
      RECT 21.96 4.926 21.965 5.134 ;
      RECT 21.955 4.92 21.96 5.132 ;
      RECT 21.886 4.765 21.955 5.12 ;
      RECT 21.8 4.765 21.886 5.094 ;
      RECT 21.775 4.765 21.8 5.073 ;
      RECT 21.77 4.765 21.775 5.063 ;
      RECT 21.765 4.765 21.77 5.055 ;
      RECT 21.745 4.765 21.765 5.038 ;
      RECT 24.165 3.335 24.425 3.595 ;
      RECT 24.15 3.335 24.425 3.498 ;
      RECT 24.12 3.335 24.425 3.473 ;
      RECT 24.085 3.175 24.365 3.455 ;
      RECT 24.055 4.665 24.115 4.925 ;
      RECT 23.08 3.355 23.135 3.615 ;
      RECT 24.015 4.622 24.055 4.925 ;
      RECT 23.986 4.543 24.015 4.925 ;
      RECT 23.9 4.415 23.986 4.925 ;
      RECT 23.88 4.295 23.9 4.925 ;
      RECT 23.855 4.246 23.88 4.925 ;
      RECT 23.85 4.211 23.855 4.775 ;
      RECT 23.82 4.171 23.85 4.713 ;
      RECT 23.795 4.108 23.82 4.628 ;
      RECT 23.785 4.07 23.795 4.565 ;
      RECT 23.77 4.045 23.785 4.526 ;
      RECT 23.727 4.003 23.77 4.432 ;
      RECT 23.725 3.976 23.727 4.359 ;
      RECT 23.72 3.971 23.725 4.35 ;
      RECT 23.715 3.964 23.72 4.325 ;
      RECT 23.71 3.958 23.715 4.31 ;
      RECT 23.705 3.952 23.71 4.298 ;
      RECT 23.695 3.943 23.705 4.28 ;
      RECT 23.69 3.934 23.695 4.258 ;
      RECT 23.665 3.915 23.69 4.208 ;
      RECT 23.66 3.896 23.665 4.158 ;
      RECT 23.645 3.882 23.66 4.118 ;
      RECT 23.64 3.868 23.645 4.085 ;
      RECT 23.635 3.861 23.64 4.078 ;
      RECT 23.62 3.848 23.635 4.07 ;
      RECT 23.575 3.81 23.62 4.043 ;
      RECT 23.545 3.763 23.575 4.008 ;
      RECT 23.525 3.732 23.545 3.985 ;
      RECT 23.445 3.665 23.525 3.938 ;
      RECT 23.415 3.595 23.445 3.885 ;
      RECT 23.41 3.572 23.415 3.868 ;
      RECT 23.38 3.55 23.41 3.853 ;
      RECT 23.35 3.509 23.38 3.825 ;
      RECT 23.345 3.484 23.35 3.81 ;
      RECT 23.34 3.478 23.345 3.803 ;
      RECT 23.33 3.355 23.34 3.795 ;
      RECT 23.32 3.355 23.33 3.788 ;
      RECT 23.315 3.355 23.32 3.78 ;
      RECT 23.295 3.355 23.315 3.768 ;
      RECT 23.245 3.355 23.295 3.738 ;
      RECT 23.19 3.355 23.245 3.688 ;
      RECT 23.16 3.355 23.19 3.648 ;
      RECT 23.135 3.355 23.16 3.625 ;
      RECT 23.005 4.08 23.285 4.36 ;
      RECT 22.97 3.995 23.23 4.255 ;
      RECT 22.97 4.077 23.24 4.255 ;
      RECT 21.17 3.45 21.175 3.935 ;
      RECT 21.06 3.635 21.065 3.935 ;
      RECT 20.97 3.675 21.035 3.935 ;
      RECT 22.645 3.175 22.735 3.805 ;
      RECT 22.61 3.225 22.615 3.805 ;
      RECT 22.555 3.25 22.565 3.805 ;
      RECT 22.51 3.25 22.52 3.805 ;
      RECT 22.88 3.175 22.925 3.455 ;
      RECT 21.73 2.905 21.93 3.045 ;
      RECT 22.846 3.175 22.88 3.467 ;
      RECT 22.76 3.175 22.846 3.507 ;
      RECT 22.745 3.175 22.76 3.548 ;
      RECT 22.74 3.175 22.745 3.568 ;
      RECT 22.735 3.175 22.74 3.588 ;
      RECT 22.615 3.217 22.645 3.805 ;
      RECT 22.565 3.237 22.61 3.805 ;
      RECT 22.55 3.252 22.555 3.805 ;
      RECT 22.52 3.252 22.55 3.805 ;
      RECT 22.475 3.237 22.51 3.805 ;
      RECT 22.47 3.225 22.475 3.585 ;
      RECT 22.465 3.222 22.47 3.565 ;
      RECT 22.45 3.212 22.465 3.518 ;
      RECT 22.445 3.205 22.45 3.481 ;
      RECT 22.44 3.202 22.445 3.464 ;
      RECT 22.425 3.192 22.44 3.42 ;
      RECT 22.42 3.183 22.425 3.38 ;
      RECT 22.415 3.179 22.42 3.365 ;
      RECT 22.405 3.173 22.415 3.348 ;
      RECT 22.365 3.154 22.405 3.323 ;
      RECT 22.36 3.136 22.365 3.303 ;
      RECT 22.35 3.13 22.36 3.298 ;
      RECT 22.32 3.114 22.35 3.285 ;
      RECT 22.305 3.096 22.32 3.268 ;
      RECT 22.29 3.084 22.305 3.255 ;
      RECT 22.285 3.076 22.29 3.248 ;
      RECT 22.255 3.062 22.285 3.235 ;
      RECT 22.25 3.047 22.255 3.223 ;
      RECT 22.24 3.041 22.25 3.215 ;
      RECT 22.22 3.029 22.24 3.203 ;
      RECT 22.21 3.017 22.22 3.19 ;
      RECT 22.18 3.001 22.21 3.175 ;
      RECT 22.16 2.981 22.18 3.158 ;
      RECT 22.155 2.971 22.16 3.148 ;
      RECT 22.13 2.959 22.155 3.135 ;
      RECT 22.125 2.947 22.13 3.123 ;
      RECT 22.12 2.942 22.125 3.119 ;
      RECT 22.105 2.935 22.12 3.111 ;
      RECT 22.095 2.922 22.105 3.101 ;
      RECT 22.09 2.92 22.095 3.095 ;
      RECT 22.065 2.913 22.09 3.084 ;
      RECT 22.06 2.906 22.065 3.073 ;
      RECT 22.035 2.905 22.06 3.06 ;
      RECT 22.016 2.905 22.035 3.05 ;
      RECT 21.93 2.905 22.016 3.047 ;
      RECT 21.7 2.905 21.73 3.05 ;
      RECT 21.66 2.912 21.7 3.063 ;
      RECT 21.635 2.922 21.66 3.076 ;
      RECT 21.62 2.931 21.635 3.086 ;
      RECT 21.59 2.936 21.62 3.105 ;
      RECT 21.585 2.942 21.59 3.123 ;
      RECT 21.565 2.952 21.585 3.138 ;
      RECT 21.555 2.965 21.565 3.158 ;
      RECT 21.54 2.977 21.555 3.175 ;
      RECT 21.535 2.987 21.54 3.185 ;
      RECT 21.53 2.992 21.535 3.19 ;
      RECT 21.52 3 21.53 3.203 ;
      RECT 21.47 3.032 21.52 3.24 ;
      RECT 21.455 3.067 21.47 3.281 ;
      RECT 21.45 3.077 21.455 3.296 ;
      RECT 21.445 3.082 21.45 3.303 ;
      RECT 21.42 3.098 21.445 3.323 ;
      RECT 21.405 3.119 21.42 3.348 ;
      RECT 21.38 3.14 21.405 3.373 ;
      RECT 21.37 3.159 21.38 3.396 ;
      RECT 21.345 3.177 21.37 3.419 ;
      RECT 21.33 3.197 21.345 3.443 ;
      RECT 21.325 3.207 21.33 3.455 ;
      RECT 21.31 3.219 21.325 3.475 ;
      RECT 21.3 3.234 21.31 3.515 ;
      RECT 21.295 3.242 21.3 3.543 ;
      RECT 21.285 3.252 21.295 3.563 ;
      RECT 21.28 3.265 21.285 3.588 ;
      RECT 21.275 3.278 21.28 3.608 ;
      RECT 21.27 3.284 21.275 3.63 ;
      RECT 21.26 3.293 21.27 3.65 ;
      RECT 21.255 3.313 21.26 3.673 ;
      RECT 21.25 3.319 21.255 3.693 ;
      RECT 21.245 3.326 21.25 3.715 ;
      RECT 21.24 3.337 21.245 3.728 ;
      RECT 21.23 3.347 21.24 3.753 ;
      RECT 21.21 3.372 21.23 3.935 ;
      RECT 21.18 3.412 21.21 3.935 ;
      RECT 21.175 3.442 21.18 3.935 ;
      RECT 21.15 3.47 21.17 3.935 ;
      RECT 21.12 3.515 21.15 3.935 ;
      RECT 21.115 3.542 21.12 3.935 ;
      RECT 21.095 3.56 21.115 3.935 ;
      RECT 21.085 3.585 21.095 3.935 ;
      RECT 21.08 3.597 21.085 3.935 ;
      RECT 21.065 3.62 21.08 3.935 ;
      RECT 21.045 3.647 21.06 3.935 ;
      RECT 21.035 3.67 21.045 3.935 ;
      RECT 22.825 4.555 22.905 4.815 ;
      RECT 22.06 3.775 22.13 4.035 ;
      RECT 22.791 4.522 22.825 4.815 ;
      RECT 22.705 4.425 22.791 4.815 ;
      RECT 22.685 4.337 22.705 4.815 ;
      RECT 22.675 4.307 22.685 4.815 ;
      RECT 22.665 4.287 22.675 4.815 ;
      RECT 22.645 4.274 22.665 4.815 ;
      RECT 22.63 4.264 22.645 4.643 ;
      RECT 22.625 4.257 22.63 4.598 ;
      RECT 22.615 4.251 22.625 4.588 ;
      RECT 22.605 4.243 22.615 4.57 ;
      RECT 22.6 4.237 22.605 4.558 ;
      RECT 22.59 4.232 22.6 4.545 ;
      RECT 22.57 4.222 22.59 4.518 ;
      RECT 22.53 4.201 22.57 4.47 ;
      RECT 22.515 4.182 22.53 4.428 ;
      RECT 22.49 4.168 22.515 4.398 ;
      RECT 22.48 4.156 22.49 4.365 ;
      RECT 22.475 4.151 22.48 4.355 ;
      RECT 22.445 4.137 22.475 4.335 ;
      RECT 22.435 4.121 22.445 4.308 ;
      RECT 22.43 4.116 22.435 4.298 ;
      RECT 22.405 4.107 22.43 4.278 ;
      RECT 22.395 4.095 22.405 4.258 ;
      RECT 22.325 4.063 22.395 4.233 ;
      RECT 22.32 4.032 22.325 4.21 ;
      RECT 22.271 3.775 22.32 4.193 ;
      RECT 22.185 3.775 22.271 4.152 ;
      RECT 22.13 3.775 22.185 4.08 ;
      RECT 22.22 4.56 22.38 4.82 ;
      RECT 21.745 3.175 21.795 3.86 ;
      RECT 21.535 3.6 21.57 3.86 ;
      RECT 21.85 3.175 21.855 3.635 ;
      RECT 21.94 3.175 21.965 3.455 ;
      RECT 22.215 4.557 22.22 4.82 ;
      RECT 22.18 4.545 22.215 4.82 ;
      RECT 22.12 4.518 22.18 4.82 ;
      RECT 22.115 4.501 22.12 4.674 ;
      RECT 22.11 4.498 22.115 4.661 ;
      RECT 22.09 4.491 22.11 4.648 ;
      RECT 22.055 4.474 22.09 4.63 ;
      RECT 22.015 4.453 22.055 4.61 ;
      RECT 22.01 4.441 22.015 4.598 ;
      RECT 21.97 4.427 22.01 4.584 ;
      RECT 21.95 4.41 21.97 4.566 ;
      RECT 21.94 4.402 21.95 4.558 ;
      RECT 21.925 3.175 21.94 3.473 ;
      RECT 21.91 4.392 21.94 4.545 ;
      RECT 21.895 3.175 21.925 3.518 ;
      RECT 21.9 4.382 21.91 4.532 ;
      RECT 21.87 4.367 21.9 4.519 ;
      RECT 21.855 3.175 21.895 3.585 ;
      RECT 21.855 4.335 21.87 4.505 ;
      RECT 21.85 4.307 21.855 4.499 ;
      RECT 21.845 3.175 21.85 3.64 ;
      RECT 21.835 4.277 21.85 4.493 ;
      RECT 21.84 3.175 21.845 3.653 ;
      RECT 21.83 3.175 21.84 3.673 ;
      RECT 21.795 4.19 21.835 4.478 ;
      RECT 21.795 3.175 21.83 3.713 ;
      RECT 21.79 4.122 21.795 4.466 ;
      RECT 21.775 4.077 21.79 4.461 ;
      RECT 21.77 4.015 21.775 4.456 ;
      RECT 21.745 3.922 21.77 4.449 ;
      RECT 21.74 3.175 21.745 4.441 ;
      RECT 21.725 3.175 21.74 4.428 ;
      RECT 21.705 3.175 21.725 4.385 ;
      RECT 21.695 3.175 21.705 4.335 ;
      RECT 21.69 3.175 21.695 4.308 ;
      RECT 21.685 3.175 21.69 4.286 ;
      RECT 21.68 3.401 21.685 4.269 ;
      RECT 21.675 3.423 21.68 4.247 ;
      RECT 21.67 3.465 21.675 4.23 ;
      RECT 21.64 3.515 21.67 4.174 ;
      RECT 21.635 3.542 21.64 4.116 ;
      RECT 21.62 3.56 21.635 4.08 ;
      RECT 21.615 3.578 21.62 4.044 ;
      RECT 21.609 3.585 21.615 4.025 ;
      RECT 21.605 3.592 21.609 4.008 ;
      RECT 21.6 3.597 21.605 3.977 ;
      RECT 21.59 3.6 21.6 3.952 ;
      RECT 21.58 3.6 21.59 3.918 ;
      RECT 21.575 3.6 21.58 3.895 ;
      RECT 21.57 3.6 21.575 3.875 ;
      RECT 20.19 4.765 20.45 5.025 ;
      RECT 20.21 4.692 20.39 5.025 ;
      RECT 20.21 4.435 20.385 5.025 ;
      RECT 20.21 4.227 20.375 5.025 ;
      RECT 20.215 4.145 20.375 5.025 ;
      RECT 20.215 3.91 20.365 5.025 ;
      RECT 20.215 3.757 20.36 5.025 ;
      RECT 20.22 3.742 20.36 5.025 ;
      RECT 20.27 3.457 20.36 5.025 ;
      RECT 20.225 3.692 20.36 5.025 ;
      RECT 20.255 3.51 20.36 5.025 ;
      RECT 20.24 3.622 20.36 5.025 ;
      RECT 20.245 3.58 20.36 5.025 ;
      RECT 20.24 3.622 20.375 3.685 ;
      RECT 20.275 3.21 20.38 3.63 ;
      RECT 20.275 3.21 20.395 3.613 ;
      RECT 20.275 3.21 20.43 3.575 ;
      RECT 20.27 3.457 20.48 3.508 ;
      RECT 20.275 3.21 20.535 3.47 ;
      RECT 19.535 3.915 19.795 4.175 ;
      RECT 19.535 3.915 19.805 4.133 ;
      RECT 19.535 3.915 19.891 4.104 ;
      RECT 19.535 3.915 19.96 4.056 ;
      RECT 19.535 3.915 19.995 4.025 ;
      RECT 19.765 3.735 20.045 4.015 ;
      RECT 19.6 3.9 20.045 4.015 ;
      RECT 19.69 3.777 19.795 4.175 ;
      RECT 19.62 3.84 20.045 4.015 ;
      RECT 93.455 7.205 93.835 7.585 ;
      RECT 85.04 9.345 85.41 9.715 ;
      RECT 78.195 7.205 78.575 7.585 ;
      RECT 69.78 9.345 70.15 9.715 ;
      RECT 62.935 7.205 63.315 7.585 ;
      RECT 54.52 9.345 54.89 9.715 ;
      RECT 47.675 7.205 48.055 7.585 ;
      RECT 39.26 9.345 39.63 9.715 ;
      RECT 32.415 7.205 32.795 7.585 ;
      RECT 24 9.345 24.37 9.715 ;
    LAYER via1 ;
      RECT 93.63 9.665 93.78 9.815 ;
      RECT 93.57 7.32 93.72 7.47 ;
      RECT 91.26 9.03 91.41 9.18 ;
      RECT 91.245 3.36 91.395 3.51 ;
      RECT 90.455 3.745 90.605 3.895 ;
      RECT 90.455 8.615 90.605 8.765 ;
      RECT 88.865 4.1 89.015 4.25 ;
      RECT 87.095 3.645 87.245 3.795 ;
      RECT 86.075 4.35 86.225 4.5 ;
      RECT 85.845 3.77 85.995 3.92 ;
      RECT 85.81 9.005 85.96 9.155 ;
      RECT 85.5 4.37 85.65 4.52 ;
      RECT 85.26 3.39 85.41 3.54 ;
      RECT 85.15 9.455 85.3 9.605 ;
      RECT 84.95 4.72 85.1 4.87 ;
      RECT 84.81 3.325 84.96 3.475 ;
      RECT 84.175 3.41 84.325 3.56 ;
      RECT 84.065 4.05 84.215 4.2 ;
      RECT 83.74 4.61 83.89 4.76 ;
      RECT 83.57 3.6 83.72 3.75 ;
      RECT 83.215 4.615 83.365 4.765 ;
      RECT 83.155 3.83 83.305 3.98 ;
      RECT 82.79 4.82 82.94 4.97 ;
      RECT 82.63 3.655 82.78 3.805 ;
      RECT 82.065 3.73 82.215 3.88 ;
      RECT 81.37 3.265 81.52 3.415 ;
      RECT 81.285 4.82 81.435 4.97 ;
      RECT 80.63 3.97 80.78 4.12 ;
      RECT 78.345 9.05 78.495 9.2 ;
      RECT 78.31 7.32 78.46 7.47 ;
      RECT 76 9.03 76.15 9.18 ;
      RECT 75.985 3.36 76.135 3.51 ;
      RECT 75.195 3.745 75.345 3.895 ;
      RECT 75.195 8.615 75.345 8.765 ;
      RECT 73.605 4.1 73.755 4.25 ;
      RECT 71.835 3.645 71.985 3.795 ;
      RECT 70.815 4.35 70.965 4.5 ;
      RECT 70.585 3.77 70.735 3.92 ;
      RECT 70.55 9.005 70.7 9.155 ;
      RECT 70.24 4.37 70.39 4.52 ;
      RECT 70 3.39 70.15 3.54 ;
      RECT 69.89 9.455 70.04 9.605 ;
      RECT 69.69 4.72 69.84 4.87 ;
      RECT 69.55 3.325 69.7 3.475 ;
      RECT 68.915 3.41 69.065 3.56 ;
      RECT 68.805 4.05 68.955 4.2 ;
      RECT 68.48 4.61 68.63 4.76 ;
      RECT 68.31 3.6 68.46 3.75 ;
      RECT 67.955 4.615 68.105 4.765 ;
      RECT 67.895 3.83 68.045 3.98 ;
      RECT 67.53 4.82 67.68 4.97 ;
      RECT 67.37 3.655 67.52 3.805 ;
      RECT 66.805 3.73 66.955 3.88 ;
      RECT 66.11 3.265 66.26 3.415 ;
      RECT 66.025 4.82 66.175 4.97 ;
      RECT 65.37 3.97 65.52 4.12 ;
      RECT 63.085 9.05 63.235 9.2 ;
      RECT 63.05 7.32 63.2 7.47 ;
      RECT 60.74 9.03 60.89 9.18 ;
      RECT 60.725 3.36 60.875 3.51 ;
      RECT 59.935 3.745 60.085 3.895 ;
      RECT 59.935 8.615 60.085 8.765 ;
      RECT 58.345 4.1 58.495 4.25 ;
      RECT 56.575 3.645 56.725 3.795 ;
      RECT 55.555 4.35 55.705 4.5 ;
      RECT 55.325 3.77 55.475 3.92 ;
      RECT 55.29 9.005 55.44 9.155 ;
      RECT 54.98 4.37 55.13 4.52 ;
      RECT 54.74 3.39 54.89 3.54 ;
      RECT 54.63 9.455 54.78 9.605 ;
      RECT 54.43 4.72 54.58 4.87 ;
      RECT 54.29 3.325 54.44 3.475 ;
      RECT 53.655 3.41 53.805 3.56 ;
      RECT 53.545 4.05 53.695 4.2 ;
      RECT 53.22 4.61 53.37 4.76 ;
      RECT 53.05 3.6 53.2 3.75 ;
      RECT 52.695 4.615 52.845 4.765 ;
      RECT 52.635 3.83 52.785 3.98 ;
      RECT 52.27 4.82 52.42 4.97 ;
      RECT 52.11 3.655 52.26 3.805 ;
      RECT 51.545 3.73 51.695 3.88 ;
      RECT 50.85 3.265 51 3.415 ;
      RECT 50.765 4.82 50.915 4.97 ;
      RECT 50.11 3.97 50.26 4.12 ;
      RECT 47.87 9.05 48.02 9.2 ;
      RECT 47.79 7.32 47.94 7.47 ;
      RECT 45.48 9.03 45.63 9.18 ;
      RECT 45.465 3.36 45.615 3.51 ;
      RECT 44.675 3.745 44.825 3.895 ;
      RECT 44.675 8.615 44.825 8.765 ;
      RECT 43.085 4.1 43.235 4.25 ;
      RECT 41.315 3.645 41.465 3.795 ;
      RECT 40.295 4.35 40.445 4.5 ;
      RECT 40.065 3.77 40.215 3.92 ;
      RECT 40.03 9.005 40.18 9.155 ;
      RECT 39.72 4.37 39.87 4.52 ;
      RECT 39.48 3.39 39.63 3.54 ;
      RECT 39.37 9.455 39.52 9.605 ;
      RECT 39.17 4.72 39.32 4.87 ;
      RECT 39.03 3.325 39.18 3.475 ;
      RECT 38.395 3.41 38.545 3.56 ;
      RECT 38.285 4.05 38.435 4.2 ;
      RECT 37.96 4.61 38.11 4.76 ;
      RECT 37.79 3.6 37.94 3.75 ;
      RECT 37.435 4.615 37.585 4.765 ;
      RECT 37.375 3.83 37.525 3.98 ;
      RECT 37.01 4.82 37.16 4.97 ;
      RECT 36.85 3.655 37 3.805 ;
      RECT 36.285 3.73 36.435 3.88 ;
      RECT 35.59 3.265 35.74 3.415 ;
      RECT 35.505 4.82 35.655 4.97 ;
      RECT 34.85 3.97 35 4.12 ;
      RECT 32.61 9.05 32.76 9.2 ;
      RECT 32.53 7.32 32.68 7.47 ;
      RECT 30.22 9.03 30.37 9.18 ;
      RECT 30.205 3.36 30.355 3.51 ;
      RECT 29.415 3.745 29.565 3.895 ;
      RECT 29.415 8.615 29.565 8.765 ;
      RECT 27.825 4.1 27.975 4.25 ;
      RECT 26.055 3.645 26.205 3.795 ;
      RECT 25.035 4.35 25.185 4.5 ;
      RECT 24.805 3.77 24.955 3.92 ;
      RECT 24.77 8.995 24.92 9.145 ;
      RECT 24.46 4.37 24.61 4.52 ;
      RECT 24.22 3.39 24.37 3.54 ;
      RECT 24.11 9.455 24.26 9.605 ;
      RECT 23.91 4.72 24.06 4.87 ;
      RECT 23.77 3.325 23.92 3.475 ;
      RECT 23.135 3.41 23.285 3.56 ;
      RECT 23.025 4.05 23.175 4.2 ;
      RECT 22.7 4.61 22.85 4.76 ;
      RECT 22.53 3.6 22.68 3.75 ;
      RECT 22.175 4.615 22.325 4.765 ;
      RECT 22.115 3.83 22.265 3.98 ;
      RECT 21.75 4.82 21.9 4.97 ;
      RECT 21.59 3.655 21.74 3.805 ;
      RECT 21.025 3.73 21.175 3.88 ;
      RECT 20.33 3.265 20.48 3.415 ;
      RECT 20.245 4.82 20.395 4.97 ;
      RECT 19.59 3.97 19.74 4.12 ;
      RECT 16.615 9.385 16.765 9.535 ;
      RECT 16.24 8.645 16.39 8.795 ;
    LAYER met1 ;
      RECT 93.495 10.06 93.79 10.29 ;
      RECT 93.555 9.565 93.73 10.29 ;
      RECT 93.53 9.565 93.88 9.915 ;
      RECT 93.555 8.58 93.725 10.29 ;
      RECT 93.495 8.58 93.785 8.81 ;
      RECT 92.505 10.06 92.8 10.29 ;
      RECT 92.565 8.58 92.735 10.29 ;
      RECT 92.505 8.58 92.795 8.81 ;
      RECT 92.505 8.615 93.355 8.775 ;
      RECT 93.19 8.21 93.355 8.775 ;
      RECT 92.505 8.61 92.9 8.775 ;
      RECT 93.125 8.21 93.415 8.44 ;
      RECT 93.125 8.24 93.585 8.41 ;
      RECT 93.09 4.025 93.41 4.26 ;
      RECT 93.09 4.055 93.58 4.225 ;
      RECT 93.09 3.69 93.28 4.26 ;
      RECT 92.505 3.655 92.795 3.885 ;
      RECT 92.505 3.69 93.28 3.86 ;
      RECT 92.565 2.175 92.735 3.885 ;
      RECT 92.505 2.175 92.8 2.405 ;
      RECT 92.135 4.025 92.425 4.255 ;
      RECT 92.135 4.055 92.595 4.225 ;
      RECT 92.2 2.95 92.365 4.255 ;
      RECT 90.715 2.915 91.005 3.145 ;
      RECT 90.715 2.95 92.365 3.12 ;
      RECT 90.775 2.175 90.945 3.145 ;
      RECT 90.715 2.175 91.005 2.405 ;
      RECT 90.715 10.06 91.005 10.29 ;
      RECT 90.775 9.32 90.945 10.29 ;
      RECT 90.775 9.41 92.365 9.58 ;
      RECT 92.195 8.21 92.365 9.58 ;
      RECT 90.715 9.32 91.005 9.55 ;
      RECT 92.135 8.21 92.425 8.44 ;
      RECT 92.135 8.24 92.595 8.41 ;
      RECT 88.765 4 89.105 4.35 ;
      RECT 88.855 3.32 89.025 4.35 ;
      RECT 91.145 3.26 91.495 3.61 ;
      RECT 88.855 3.32 91.495 3.49 ;
      RECT 90.975 3.315 91.495 3.49 ;
      RECT 91.17 8.945 91.495 9.27 ;
      RECT 85.71 8.905 86.06 9.255 ;
      RECT 91.145 8.95 91.495 9.18 ;
      RECT 85.51 8.95 86.06 9.18 ;
      RECT 90.975 8.975 91.495 9.15 ;
      RECT 85.34 8.98 86.06 9.15 ;
      RECT 85.39 8.975 91.495 9.145 ;
      RECT 90.37 3.66 90.69 3.98 ;
      RECT 90.345 3.655 90.635 3.885 ;
      RECT 90.34 3.685 90.69 3.86 ;
      RECT 90.17 3.685 90.69 3.855 ;
      RECT 90.37 8.545 90.69 8.835 ;
      RECT 90.345 8.58 90.69 8.81 ;
      RECT 90.17 8.61 90.69 8.78 ;
      RECT 86.06 4.28 86.21 4.555 ;
      RECT 86.6 3.36 86.605 3.58 ;
      RECT 87.75 3.56 87.765 3.758 ;
      RECT 87.715 3.552 87.75 3.765 ;
      RECT 87.685 3.545 87.715 3.765 ;
      RECT 87.63 3.51 87.685 3.765 ;
      RECT 87.565 3.447 87.63 3.765 ;
      RECT 87.56 3.412 87.565 3.763 ;
      RECT 87.555 3.407 87.56 3.755 ;
      RECT 87.55 3.402 87.555 3.741 ;
      RECT 87.545 3.399 87.55 3.734 ;
      RECT 87.5 3.389 87.545 3.685 ;
      RECT 87.48 3.376 87.5 3.62 ;
      RECT 87.475 3.371 87.48 3.593 ;
      RECT 87.47 3.37 87.475 3.586 ;
      RECT 87.465 3.369 87.47 3.579 ;
      RECT 87.38 3.354 87.465 3.525 ;
      RECT 87.35 3.335 87.38 3.475 ;
      RECT 87.27 3.318 87.35 3.46 ;
      RECT 87.235 3.305 87.27 3.445 ;
      RECT 87.227 3.305 87.235 3.44 ;
      RECT 87.141 3.306 87.227 3.44 ;
      RECT 87.055 3.308 87.141 3.44 ;
      RECT 87.03 3.309 87.055 3.444 ;
      RECT 86.955 3.315 87.03 3.459 ;
      RECT 86.872 3.327 86.955 3.483 ;
      RECT 86.786 3.34 86.872 3.509 ;
      RECT 86.7 3.353 86.786 3.535 ;
      RECT 86.665 3.362 86.7 3.554 ;
      RECT 86.615 3.362 86.665 3.567 ;
      RECT 86.605 3.36 86.615 3.578 ;
      RECT 86.59 3.357 86.6 3.58 ;
      RECT 86.575 3.349 86.59 3.588 ;
      RECT 86.56 3.341 86.575 3.608 ;
      RECT 86.555 3.336 86.56 3.665 ;
      RECT 86.54 3.331 86.555 3.738 ;
      RECT 86.535 3.326 86.54 3.78 ;
      RECT 86.53 3.324 86.535 3.808 ;
      RECT 86.525 3.322 86.53 3.83 ;
      RECT 86.515 3.318 86.525 3.873 ;
      RECT 86.51 3.315 86.515 3.898 ;
      RECT 86.505 3.313 86.51 3.918 ;
      RECT 86.5 3.311 86.505 3.942 ;
      RECT 86.495 3.307 86.5 3.965 ;
      RECT 86.49 3.303 86.495 3.988 ;
      RECT 86.455 3.293 86.49 4.095 ;
      RECT 86.45 3.283 86.455 4.193 ;
      RECT 86.445 3.281 86.45 4.22 ;
      RECT 86.44 3.28 86.445 4.24 ;
      RECT 86.435 3.272 86.44 4.26 ;
      RECT 86.43 3.267 86.435 4.295 ;
      RECT 86.425 3.265 86.43 4.313 ;
      RECT 86.42 3.265 86.425 4.338 ;
      RECT 86.415 3.265 86.42 4.36 ;
      RECT 86.38 3.265 86.415 4.403 ;
      RECT 86.355 3.265 86.38 4.432 ;
      RECT 86.345 3.265 86.355 3.618 ;
      RECT 86.348 3.675 86.355 4.442 ;
      RECT 86.345 3.732 86.348 4.445 ;
      RECT 86.34 3.265 86.345 3.59 ;
      RECT 86.34 3.782 86.345 4.448 ;
      RECT 86.33 3.265 86.34 3.58 ;
      RECT 86.335 3.835 86.34 4.451 ;
      RECT 86.33 3.92 86.335 4.455 ;
      RECT 86.32 3.265 86.33 3.568 ;
      RECT 86.325 3.967 86.33 4.459 ;
      RECT 86.32 4.042 86.325 4.463 ;
      RECT 86.285 3.265 86.32 3.543 ;
      RECT 86.31 4.125 86.32 4.468 ;
      RECT 86.3 4.192 86.31 4.475 ;
      RECT 86.295 4.22 86.3 4.48 ;
      RECT 86.285 4.233 86.295 4.486 ;
      RECT 86.24 3.265 86.285 3.5 ;
      RECT 86.28 4.238 86.285 4.493 ;
      RECT 86.24 4.255 86.28 4.555 ;
      RECT 86.235 3.267 86.24 3.473 ;
      RECT 86.21 4.275 86.24 4.555 ;
      RECT 86.23 3.272 86.235 3.445 ;
      RECT 86.02 4.284 86.06 4.555 ;
      RECT 85.995 4.292 86.02 4.525 ;
      RECT 85.95 4.3 85.995 4.525 ;
      RECT 85.935 4.305 85.95 4.52 ;
      RECT 85.925 4.305 85.935 4.514 ;
      RECT 85.915 4.312 85.925 4.511 ;
      RECT 85.91 4.35 85.915 4.5 ;
      RECT 85.905 4.412 85.91 4.478 ;
      RECT 87.175 4.287 87.36 4.51 ;
      RECT 87.175 4.302 87.365 4.506 ;
      RECT 87.165 3.575 87.25 4.505 ;
      RECT 87.165 4.302 87.37 4.499 ;
      RECT 87.16 4.31 87.37 4.498 ;
      RECT 87.365 4.03 87.685 4.35 ;
      RECT 87.16 4.202 87.33 4.293 ;
      RECT 87.155 4.202 87.33 4.275 ;
      RECT 87.145 4.01 87.28 4.25 ;
      RECT 87.14 4.01 87.28 4.195 ;
      RECT 87.1 3.59 87.27 4.095 ;
      RECT 87.085 3.59 87.27 3.965 ;
      RECT 87.08 3.59 87.27 3.918 ;
      RECT 87.075 3.59 87.27 3.898 ;
      RECT 87.07 3.59 87.27 3.873 ;
      RECT 87.04 3.59 87.3 3.85 ;
      RECT 87.05 3.587 87.26 3.85 ;
      RECT 87.175 3.582 87.26 4.51 ;
      RECT 87.06 3.575 87.25 3.85 ;
      RECT 87.055 3.58 87.25 3.85 ;
      RECT 85.885 3.792 86.07 4.005 ;
      RECT 85.885 3.8 86.08 3.998 ;
      RECT 85.865 3.8 86.08 3.995 ;
      RECT 85.86 3.8 86.08 3.98 ;
      RECT 85.79 3.715 86.05 3.975 ;
      RECT 85.79 3.86 86.085 3.888 ;
      RECT 85.445 4.315 85.705 4.575 ;
      RECT 85.47 4.26 85.665 4.575 ;
      RECT 85.465 4.009 85.645 4.303 ;
      RECT 85.465 4.015 85.655 4.303 ;
      RECT 85.445 4.017 85.655 4.248 ;
      RECT 85.44 4.027 85.655 4.115 ;
      RECT 85.47 4.007 85.645 4.575 ;
      RECT 85.556 4.005 85.645 4.575 ;
      RECT 85.415 3.225 85.45 3.595 ;
      RECT 85.205 3.335 85.21 3.595 ;
      RECT 85.45 3.232 85.465 3.595 ;
      RECT 85.34 3.225 85.415 3.673 ;
      RECT 85.33 3.225 85.34 3.758 ;
      RECT 85.305 3.225 85.33 3.793 ;
      RECT 85.265 3.225 85.305 3.861 ;
      RECT 85.255 3.232 85.265 3.913 ;
      RECT 85.225 3.335 85.255 3.954 ;
      RECT 85.22 3.335 85.225 3.993 ;
      RECT 85.21 3.335 85.22 4.013 ;
      RECT 85.205 3.63 85.21 4.05 ;
      RECT 85.2 3.647 85.205 4.07 ;
      RECT 85.185 3.71 85.2 4.11 ;
      RECT 85.18 3.753 85.185 4.145 ;
      RECT 85.175 3.761 85.18 4.158 ;
      RECT 85.165 3.775 85.175 4.18 ;
      RECT 85.14 3.81 85.165 4.245 ;
      RECT 85.13 3.845 85.14 4.308 ;
      RECT 85.11 3.875 85.13 4.369 ;
      RECT 85.095 3.911 85.11 4.436 ;
      RECT 85.085 3.939 85.095 4.475 ;
      RECT 85.075 3.961 85.085 4.495 ;
      RECT 85.07 3.971 85.075 4.506 ;
      RECT 85.065 3.98 85.07 4.509 ;
      RECT 85.055 3.998 85.065 4.513 ;
      RECT 85.045 4.016 85.055 4.514 ;
      RECT 85.02 4.055 85.045 4.511 ;
      RECT 85 4.097 85.02 4.508 ;
      RECT 84.985 4.135 85 4.507 ;
      RECT 84.95 4.17 84.985 4.504 ;
      RECT 84.945 4.192 84.95 4.502 ;
      RECT 84.88 4.232 84.945 4.499 ;
      RECT 84.875 4.272 84.88 4.495 ;
      RECT 84.86 4.282 84.875 4.486 ;
      RECT 84.85 4.402 84.86 4.471 ;
      RECT 85.33 4.815 85.34 5.075 ;
      RECT 85.33 4.818 85.35 5.074 ;
      RECT 85.32 4.808 85.33 5.073 ;
      RECT 85.31 4.823 85.39 5.069 ;
      RECT 85.295 4.802 85.31 5.067 ;
      RECT 85.27 4.827 85.395 5.063 ;
      RECT 85.255 4.787 85.27 5.058 ;
      RECT 85.255 4.829 85.405 5.057 ;
      RECT 85.255 4.837 85.42 5.05 ;
      RECT 85.195 4.774 85.255 5.04 ;
      RECT 85.185 4.761 85.195 5.022 ;
      RECT 85.16 4.751 85.185 5.012 ;
      RECT 85.155 4.741 85.16 5.004 ;
      RECT 85.09 4.837 85.42 4.986 ;
      RECT 85.005 4.837 85.42 4.948 ;
      RECT 84.895 4.665 85.155 4.925 ;
      RECT 85.27 4.795 85.295 5.063 ;
      RECT 85.31 4.805 85.32 5.069 ;
      RECT 84.895 4.813 85.335 4.925 ;
      RECT 85.08 10.06 85.37 10.29 ;
      RECT 85.14 9.32 85.31 10.29 ;
      RECT 85.04 9.345 85.41 9.715 ;
      RECT 85.08 9.32 85.37 9.715 ;
      RECT 84.11 4.57 84.14 4.87 ;
      RECT 83.885 4.555 83.89 4.83 ;
      RECT 83.685 4.555 83.84 4.815 ;
      RECT 84.985 3.27 85.015 3.53 ;
      RECT 84.975 3.27 84.985 3.638 ;
      RECT 84.955 3.27 84.975 3.648 ;
      RECT 84.94 3.27 84.955 3.66 ;
      RECT 84.885 3.27 84.94 3.71 ;
      RECT 84.87 3.27 84.885 3.758 ;
      RECT 84.84 3.27 84.87 3.793 ;
      RECT 84.785 3.27 84.84 3.855 ;
      RECT 84.765 3.27 84.785 3.923 ;
      RECT 84.76 3.27 84.765 3.953 ;
      RECT 84.755 3.27 84.76 3.965 ;
      RECT 84.75 3.387 84.755 3.983 ;
      RECT 84.73 3.405 84.75 4.008 ;
      RECT 84.71 3.432 84.73 4.058 ;
      RECT 84.705 3.452 84.71 4.089 ;
      RECT 84.7 3.46 84.705 4.106 ;
      RECT 84.685 3.486 84.7 4.135 ;
      RECT 84.67 3.528 84.685 4.17 ;
      RECT 84.665 3.557 84.67 4.193 ;
      RECT 84.66 3.572 84.665 4.206 ;
      RECT 84.655 3.595 84.66 4.217 ;
      RECT 84.645 3.615 84.655 4.235 ;
      RECT 84.635 3.645 84.645 4.258 ;
      RECT 84.63 3.667 84.635 4.278 ;
      RECT 84.625 3.682 84.63 4.293 ;
      RECT 84.61 3.712 84.625 4.32 ;
      RECT 84.605 3.742 84.61 4.346 ;
      RECT 84.6 3.76 84.605 4.358 ;
      RECT 84.59 3.79 84.6 4.377 ;
      RECT 84.58 3.815 84.59 4.402 ;
      RECT 84.575 3.835 84.58 4.421 ;
      RECT 84.57 3.852 84.575 4.434 ;
      RECT 84.56 3.878 84.57 4.453 ;
      RECT 84.55 3.916 84.56 4.48 ;
      RECT 84.545 3.942 84.55 4.5 ;
      RECT 84.54 3.952 84.545 4.51 ;
      RECT 84.535 3.965 84.54 4.525 ;
      RECT 84.53 3.98 84.535 4.535 ;
      RECT 84.525 4.002 84.53 4.55 ;
      RECT 84.52 4.02 84.525 4.561 ;
      RECT 84.515 4.03 84.52 4.572 ;
      RECT 84.51 4.038 84.515 4.584 ;
      RECT 84.505 4.046 84.51 4.595 ;
      RECT 84.5 4.072 84.505 4.608 ;
      RECT 84.49 4.1 84.5 4.621 ;
      RECT 84.485 4.13 84.49 4.63 ;
      RECT 84.48 4.145 84.485 4.637 ;
      RECT 84.465 4.17 84.48 4.644 ;
      RECT 84.46 4.192 84.465 4.65 ;
      RECT 84.455 4.217 84.46 4.653 ;
      RECT 84.446 4.245 84.455 4.657 ;
      RECT 84.44 4.262 84.446 4.662 ;
      RECT 84.435 4.28 84.44 4.666 ;
      RECT 84.43 4.292 84.435 4.669 ;
      RECT 84.425 4.313 84.43 4.673 ;
      RECT 84.42 4.331 84.425 4.676 ;
      RECT 84.415 4.345 84.42 4.679 ;
      RECT 84.41 4.362 84.415 4.682 ;
      RECT 84.405 4.375 84.41 4.685 ;
      RECT 84.38 4.412 84.405 4.693 ;
      RECT 84.375 4.457 84.38 4.702 ;
      RECT 84.37 4.485 84.375 4.705 ;
      RECT 84.36 4.505 84.37 4.709 ;
      RECT 84.355 4.525 84.36 4.714 ;
      RECT 84.35 4.54 84.355 4.717 ;
      RECT 84.33 4.55 84.35 4.724 ;
      RECT 84.265 4.557 84.33 4.75 ;
      RECT 84.23 4.56 84.265 4.778 ;
      RECT 84.215 4.563 84.23 4.793 ;
      RECT 84.205 4.564 84.215 4.808 ;
      RECT 84.195 4.565 84.205 4.825 ;
      RECT 84.19 4.565 84.195 4.84 ;
      RECT 84.185 4.565 84.19 4.848 ;
      RECT 84.17 4.566 84.185 4.863 ;
      RECT 84.14 4.568 84.17 4.87 ;
      RECT 84.03 4.575 84.11 4.87 ;
      RECT 83.985 4.58 84.03 4.87 ;
      RECT 83.975 4.581 83.985 4.86 ;
      RECT 83.965 4.582 83.975 4.853 ;
      RECT 83.945 4.584 83.965 4.848 ;
      RECT 83.935 4.555 83.945 4.843 ;
      RECT 83.89 4.555 83.935 4.835 ;
      RECT 83.86 4.555 83.885 4.825 ;
      RECT 83.84 4.555 83.86 4.818 ;
      RECT 84.12 3.355 84.38 3.615 ;
      RECT 84 3.37 84.01 3.535 ;
      RECT 83.985 3.37 83.99 3.53 ;
      RECT 81.35 3.21 81.535 3.5 ;
      RECT 83.165 3.335 83.18 3.49 ;
      RECT 81.315 3.21 81.34 3.47 ;
      RECT 83.73 3.26 83.735 3.402 ;
      RECT 83.645 3.255 83.67 3.395 ;
      RECT 84.045 3.372 84.12 3.565 ;
      RECT 84.03 3.37 84.045 3.548 ;
      RECT 84.01 3.37 84.03 3.54 ;
      RECT 83.99 3.37 84 3.533 ;
      RECT 83.945 3.365 83.985 3.523 ;
      RECT 83.905 3.34 83.945 3.508 ;
      RECT 83.89 3.315 83.905 3.498 ;
      RECT 83.885 3.309 83.89 3.496 ;
      RECT 83.85 3.301 83.885 3.479 ;
      RECT 83.845 3.294 83.85 3.467 ;
      RECT 83.825 3.289 83.845 3.455 ;
      RECT 83.815 3.283 83.825 3.44 ;
      RECT 83.795 3.278 83.815 3.425 ;
      RECT 83.785 3.273 83.795 3.418 ;
      RECT 83.78 3.271 83.785 3.413 ;
      RECT 83.775 3.27 83.78 3.41 ;
      RECT 83.735 3.265 83.775 3.406 ;
      RECT 83.715 3.259 83.73 3.401 ;
      RECT 83.68 3.256 83.715 3.398 ;
      RECT 83.67 3.255 83.68 3.396 ;
      RECT 83.61 3.255 83.645 3.393 ;
      RECT 83.565 3.255 83.61 3.393 ;
      RECT 83.515 3.255 83.565 3.396 ;
      RECT 83.5 3.257 83.515 3.398 ;
      RECT 83.485 3.26 83.5 3.399 ;
      RECT 83.475 3.265 83.485 3.4 ;
      RECT 83.445 3.27 83.475 3.405 ;
      RECT 83.435 3.276 83.445 3.413 ;
      RECT 83.425 3.278 83.435 3.417 ;
      RECT 83.415 3.282 83.425 3.421 ;
      RECT 83.39 3.288 83.415 3.429 ;
      RECT 83.38 3.293 83.39 3.437 ;
      RECT 83.365 3.297 83.38 3.441 ;
      RECT 83.33 3.303 83.365 3.449 ;
      RECT 83.31 3.308 83.33 3.459 ;
      RECT 83.28 3.315 83.31 3.468 ;
      RECT 83.235 3.324 83.28 3.482 ;
      RECT 83.23 3.329 83.235 3.493 ;
      RECT 83.21 3.332 83.23 3.494 ;
      RECT 83.18 3.335 83.21 3.492 ;
      RECT 83.145 3.335 83.165 3.488 ;
      RECT 83.075 3.335 83.145 3.479 ;
      RECT 83.06 3.332 83.075 3.471 ;
      RECT 83.02 3.325 83.06 3.466 ;
      RECT 82.995 3.315 83.02 3.459 ;
      RECT 82.99 3.309 82.995 3.456 ;
      RECT 82.95 3.303 82.99 3.453 ;
      RECT 82.935 3.296 82.95 3.448 ;
      RECT 82.915 3.292 82.935 3.443 ;
      RECT 82.9 3.287 82.915 3.439 ;
      RECT 82.885 3.282 82.9 3.437 ;
      RECT 82.87 3.278 82.885 3.436 ;
      RECT 82.855 3.276 82.87 3.432 ;
      RECT 82.845 3.274 82.855 3.427 ;
      RECT 82.83 3.271 82.845 3.423 ;
      RECT 82.82 3.269 82.83 3.418 ;
      RECT 82.8 3.266 82.82 3.414 ;
      RECT 82.755 3.265 82.8 3.412 ;
      RECT 82.695 3.267 82.755 3.413 ;
      RECT 82.675 3.269 82.695 3.415 ;
      RECT 82.645 3.272 82.675 3.416 ;
      RECT 82.595 3.277 82.645 3.418 ;
      RECT 82.59 3.28 82.595 3.42 ;
      RECT 82.58 3.282 82.59 3.423 ;
      RECT 82.575 3.284 82.58 3.426 ;
      RECT 82.525 3.287 82.575 3.433 ;
      RECT 82.505 3.291 82.525 3.445 ;
      RECT 82.495 3.294 82.505 3.451 ;
      RECT 82.485 3.295 82.495 3.454 ;
      RECT 82.446 3.298 82.485 3.456 ;
      RECT 82.36 3.305 82.446 3.459 ;
      RECT 82.286 3.315 82.36 3.463 ;
      RECT 82.2 3.326 82.286 3.468 ;
      RECT 82.185 3.333 82.2 3.47 ;
      RECT 82.13 3.337 82.185 3.471 ;
      RECT 82.116 3.34 82.13 3.473 ;
      RECT 82.03 3.34 82.116 3.475 ;
      RECT 81.99 3.337 82.03 3.478 ;
      RECT 81.966 3.333 81.99 3.48 ;
      RECT 81.88 3.323 81.966 3.483 ;
      RECT 81.85 3.312 81.88 3.484 ;
      RECT 81.831 3.308 81.85 3.483 ;
      RECT 81.745 3.301 81.831 3.48 ;
      RECT 81.685 3.29 81.745 3.477 ;
      RECT 81.665 3.282 81.685 3.475 ;
      RECT 81.63 3.277 81.665 3.474 ;
      RECT 81.605 3.272 81.63 3.473 ;
      RECT 81.575 3.267 81.605 3.472 ;
      RECT 81.55 3.21 81.575 3.471 ;
      RECT 81.535 3.21 81.55 3.495 ;
      RECT 81.34 3.21 81.35 3.495 ;
      RECT 83.115 4.23 83.12 4.37 ;
      RECT 82.775 4.23 82.81 4.368 ;
      RECT 82.35 4.215 82.365 4.36 ;
      RECT 84.18 3.995 84.27 4.255 ;
      RECT 84.01 3.86 84.11 4.255 ;
      RECT 81.045 3.835 81.125 4.045 ;
      RECT 84.135 3.972 84.18 4.255 ;
      RECT 84.125 3.942 84.135 4.255 ;
      RECT 84.11 3.865 84.125 4.255 ;
      RECT 83.925 3.86 84.01 4.22 ;
      RECT 83.92 3.862 83.925 4.215 ;
      RECT 83.915 3.867 83.92 4.215 ;
      RECT 83.88 3.967 83.915 4.215 ;
      RECT 83.87 3.995 83.88 4.215 ;
      RECT 83.86 4.01 83.87 4.215 ;
      RECT 83.85 4.022 83.86 4.215 ;
      RECT 83.845 4.032 83.85 4.215 ;
      RECT 83.83 4.042 83.845 4.217 ;
      RECT 83.825 4.057 83.83 4.219 ;
      RECT 83.81 4.07 83.825 4.221 ;
      RECT 83.805 4.085 83.81 4.224 ;
      RECT 83.785 4.095 83.805 4.228 ;
      RECT 83.77 4.105 83.785 4.231 ;
      RECT 83.735 4.112 83.77 4.236 ;
      RECT 83.691 4.119 83.735 4.244 ;
      RECT 83.605 4.131 83.691 4.257 ;
      RECT 83.58 4.142 83.605 4.268 ;
      RECT 83.55 4.147 83.58 4.273 ;
      RECT 83.515 4.152 83.55 4.281 ;
      RECT 83.485 4.157 83.515 4.288 ;
      RECT 83.46 4.162 83.485 4.293 ;
      RECT 83.395 4.169 83.46 4.302 ;
      RECT 83.325 4.182 83.395 4.318 ;
      RECT 83.295 4.192 83.325 4.33 ;
      RECT 83.27 4.197 83.295 4.337 ;
      RECT 83.215 4.204 83.27 4.345 ;
      RECT 83.21 4.211 83.215 4.35 ;
      RECT 83.205 4.213 83.21 4.351 ;
      RECT 83.19 4.215 83.205 4.353 ;
      RECT 83.185 4.215 83.19 4.356 ;
      RECT 83.12 4.222 83.185 4.363 ;
      RECT 83.085 4.232 83.115 4.373 ;
      RECT 83.068 4.235 83.085 4.375 ;
      RECT 82.982 4.234 83.068 4.374 ;
      RECT 82.896 4.232 82.982 4.371 ;
      RECT 82.81 4.231 82.896 4.369 ;
      RECT 82.709 4.229 82.775 4.368 ;
      RECT 82.623 4.226 82.709 4.366 ;
      RECT 82.537 4.222 82.623 4.364 ;
      RECT 82.451 4.219 82.537 4.363 ;
      RECT 82.365 4.216 82.451 4.361 ;
      RECT 82.265 4.215 82.35 4.358 ;
      RECT 82.215 4.213 82.265 4.356 ;
      RECT 82.195 4.21 82.215 4.354 ;
      RECT 82.175 4.208 82.195 4.351 ;
      RECT 82.15 4.204 82.175 4.348 ;
      RECT 82.105 4.198 82.15 4.343 ;
      RECT 82.065 4.192 82.105 4.335 ;
      RECT 82.04 4.187 82.065 4.328 ;
      RECT 81.985 4.18 82.04 4.32 ;
      RECT 81.961 4.173 81.985 4.313 ;
      RECT 81.875 4.164 81.961 4.303 ;
      RECT 81.845 4.156 81.875 4.293 ;
      RECT 81.815 4.152 81.845 4.288 ;
      RECT 81.81 4.149 81.815 4.285 ;
      RECT 81.805 4.148 81.81 4.285 ;
      RECT 81.73 4.141 81.805 4.278 ;
      RECT 81.691 4.132 81.73 4.267 ;
      RECT 81.605 4.122 81.691 4.255 ;
      RECT 81.565 4.112 81.605 4.243 ;
      RECT 81.526 4.107 81.565 4.236 ;
      RECT 81.44 4.097 81.526 4.225 ;
      RECT 81.4 4.085 81.44 4.214 ;
      RECT 81.365 4.07 81.4 4.207 ;
      RECT 81.355 4.06 81.365 4.204 ;
      RECT 81.335 4.045 81.355 4.202 ;
      RECT 81.305 4.015 81.335 4.198 ;
      RECT 81.295 3.995 81.305 4.193 ;
      RECT 81.29 3.987 81.295 4.19 ;
      RECT 81.285 3.98 81.29 4.188 ;
      RECT 81.27 3.967 81.285 4.181 ;
      RECT 81.265 3.957 81.27 4.173 ;
      RECT 81.26 3.95 81.265 4.168 ;
      RECT 81.255 3.945 81.26 4.164 ;
      RECT 81.24 3.932 81.255 4.156 ;
      RECT 81.235 3.842 81.24 4.145 ;
      RECT 81.23 3.837 81.235 4.138 ;
      RECT 81.155 3.835 81.23 4.098 ;
      RECT 81.125 3.835 81.155 4.053 ;
      RECT 81.03 3.84 81.045 4.04 ;
      RECT 83.515 3.545 83.775 3.805 ;
      RECT 83.5 3.533 83.68 3.77 ;
      RECT 83.495 3.534 83.68 3.768 ;
      RECT 83.48 3.538 83.69 3.758 ;
      RECT 83.475 3.543 83.695 3.728 ;
      RECT 83.48 3.54 83.695 3.758 ;
      RECT 83.495 3.535 83.69 3.768 ;
      RECT 83.515 3.532 83.68 3.805 ;
      RECT 83.515 3.531 83.67 3.805 ;
      RECT 83.54 3.53 83.67 3.805 ;
      RECT 83.1 3.775 83.36 4.035 ;
      RECT 82.975 3.82 83.36 4.03 ;
      RECT 82.965 3.825 83.36 4.025 ;
      RECT 82.98 4.765 82.995 5.075 ;
      RECT 81.575 4.535 81.585 4.665 ;
      RECT 81.355 4.53 81.46 4.665 ;
      RECT 81.27 4.535 81.32 4.665 ;
      RECT 79.82 3.27 79.825 4.375 ;
      RECT 83.075 4.857 83.08 4.993 ;
      RECT 83.07 4.852 83.075 5.053 ;
      RECT 83.065 4.85 83.07 5.066 ;
      RECT 83.05 4.847 83.065 5.068 ;
      RECT 83.045 4.842 83.05 5.07 ;
      RECT 83.04 4.838 83.045 5.073 ;
      RECT 83.025 4.833 83.04 5.075 ;
      RECT 82.995 4.825 83.025 5.075 ;
      RECT 82.956 4.765 82.98 5.075 ;
      RECT 82.87 4.765 82.956 5.072 ;
      RECT 82.84 4.765 82.87 5.065 ;
      RECT 82.815 4.765 82.84 5.058 ;
      RECT 82.79 4.765 82.815 5.05 ;
      RECT 82.775 4.765 82.79 5.043 ;
      RECT 82.75 4.765 82.775 5.035 ;
      RECT 82.735 4.765 82.75 5.028 ;
      RECT 82.695 4.775 82.735 5.017 ;
      RECT 82.685 4.77 82.695 5.007 ;
      RECT 82.681 4.769 82.685 5.004 ;
      RECT 82.595 4.761 82.681 4.987 ;
      RECT 82.562 4.75 82.595 4.964 ;
      RECT 82.476 4.739 82.562 4.942 ;
      RECT 82.39 4.723 82.476 4.911 ;
      RECT 82.32 4.708 82.39 4.883 ;
      RECT 82.31 4.701 82.32 4.87 ;
      RECT 82.28 4.698 82.31 4.86 ;
      RECT 82.255 4.694 82.28 4.853 ;
      RECT 82.24 4.691 82.255 4.848 ;
      RECT 82.235 4.69 82.24 4.843 ;
      RECT 82.205 4.685 82.235 4.836 ;
      RECT 82.2 4.68 82.205 4.831 ;
      RECT 82.185 4.677 82.2 4.826 ;
      RECT 82.18 4.672 82.185 4.821 ;
      RECT 82.16 4.667 82.18 4.818 ;
      RECT 82.145 4.662 82.16 4.81 ;
      RECT 82.13 4.656 82.145 4.805 ;
      RECT 82.1 4.647 82.13 4.798 ;
      RECT 82.095 4.64 82.1 4.79 ;
      RECT 82.09 4.638 82.095 4.788 ;
      RECT 82.085 4.637 82.09 4.785 ;
      RECT 82.045 4.63 82.085 4.778 ;
      RECT 82.031 4.62 82.045 4.768 ;
      RECT 81.98 4.609 82.031 4.756 ;
      RECT 81.955 4.595 81.98 4.742 ;
      RECT 81.93 4.584 81.955 4.734 ;
      RECT 81.91 4.573 81.93 4.728 ;
      RECT 81.9 4.567 81.91 4.723 ;
      RECT 81.895 4.565 81.9 4.719 ;
      RECT 81.875 4.56 81.895 4.714 ;
      RECT 81.845 4.55 81.875 4.704 ;
      RECT 81.84 4.542 81.845 4.697 ;
      RECT 81.825 4.54 81.84 4.693 ;
      RECT 81.805 4.54 81.825 4.688 ;
      RECT 81.8 4.539 81.805 4.686 ;
      RECT 81.795 4.539 81.8 4.683 ;
      RECT 81.755 4.538 81.795 4.678 ;
      RECT 81.73 4.537 81.755 4.673 ;
      RECT 81.67 4.536 81.73 4.67 ;
      RECT 81.585 4.535 81.67 4.668 ;
      RECT 81.546 4.534 81.575 4.665 ;
      RECT 81.46 4.532 81.546 4.665 ;
      RECT 81.32 4.532 81.355 4.665 ;
      RECT 81.23 4.536 81.27 4.668 ;
      RECT 81.215 4.539 81.23 4.675 ;
      RECT 81.205 4.54 81.215 4.682 ;
      RECT 81.18 4.543 81.205 4.687 ;
      RECT 81.175 4.545 81.18 4.69 ;
      RECT 81.125 4.547 81.175 4.691 ;
      RECT 81.086 4.551 81.125 4.693 ;
      RECT 81 4.553 81.086 4.696 ;
      RECT 80.982 4.555 81 4.698 ;
      RECT 80.896 4.558 80.982 4.7 ;
      RECT 80.81 4.562 80.896 4.703 ;
      RECT 80.773 4.566 80.81 4.706 ;
      RECT 80.687 4.569 80.773 4.709 ;
      RECT 80.601 4.573 80.687 4.712 ;
      RECT 80.515 4.578 80.601 4.716 ;
      RECT 80.495 4.58 80.515 4.719 ;
      RECT 80.475 4.579 80.495 4.72 ;
      RECT 80.426 4.576 80.475 4.721 ;
      RECT 80.34 4.571 80.426 4.724 ;
      RECT 80.29 4.566 80.34 4.726 ;
      RECT 80.266 4.564 80.29 4.727 ;
      RECT 80.18 4.559 80.266 4.729 ;
      RECT 80.155 4.555 80.18 4.728 ;
      RECT 80.145 4.552 80.155 4.726 ;
      RECT 80.135 4.545 80.145 4.723 ;
      RECT 80.13 4.525 80.135 4.718 ;
      RECT 80.12 4.495 80.13 4.713 ;
      RECT 80.105 4.365 80.12 4.704 ;
      RECT 80.1 4.357 80.105 4.697 ;
      RECT 80.08 4.35 80.1 4.689 ;
      RECT 80.075 4.332 80.08 4.681 ;
      RECT 80.065 4.312 80.075 4.676 ;
      RECT 80.06 4.285 80.065 4.672 ;
      RECT 80.055 4.262 80.06 4.669 ;
      RECT 80.035 4.22 80.055 4.661 ;
      RECT 80 4.135 80.035 4.645 ;
      RECT 79.995 4.067 80 4.633 ;
      RECT 79.98 4.037 79.995 4.627 ;
      RECT 79.975 3.282 79.98 3.528 ;
      RECT 79.965 4.007 79.98 4.618 ;
      RECT 79.97 3.277 79.975 3.56 ;
      RECT 79.965 3.272 79.97 3.603 ;
      RECT 79.96 3.27 79.965 3.638 ;
      RECT 79.945 3.97 79.965 4.608 ;
      RECT 79.955 3.27 79.96 3.675 ;
      RECT 79.94 3.27 79.955 3.773 ;
      RECT 79.94 3.943 79.945 4.601 ;
      RECT 79.935 3.27 79.94 3.848 ;
      RECT 79.935 3.931 79.94 4.598 ;
      RECT 79.93 3.27 79.935 3.88 ;
      RECT 79.93 3.91 79.935 4.595 ;
      RECT 79.925 3.27 79.93 4.592 ;
      RECT 79.89 3.27 79.925 4.578 ;
      RECT 79.875 3.27 79.89 4.56 ;
      RECT 79.855 3.27 79.875 4.55 ;
      RECT 79.83 3.27 79.855 4.533 ;
      RECT 79.825 3.27 79.83 4.483 ;
      RECT 79.815 3.27 79.82 4.313 ;
      RECT 79.81 3.27 79.815 4.22 ;
      RECT 79.805 3.27 79.81 4.133 ;
      RECT 79.8 3.27 79.805 4.065 ;
      RECT 79.795 3.27 79.8 4.008 ;
      RECT 79.785 3.27 79.795 3.903 ;
      RECT 79.78 3.27 79.785 3.775 ;
      RECT 79.775 3.27 79.78 3.693 ;
      RECT 79.77 3.272 79.775 3.61 ;
      RECT 79.765 3.277 79.77 3.543 ;
      RECT 79.76 3.282 79.765 3.47 ;
      RECT 82.575 3.6 82.835 3.86 ;
      RECT 82.595 3.567 82.805 3.86 ;
      RECT 82.595 3.565 82.795 3.86 ;
      RECT 82.605 3.552 82.795 3.86 ;
      RECT 82.605 3.55 82.72 3.86 ;
      RECT 82.08 3.675 82.255 3.955 ;
      RECT 82.075 3.675 82.255 3.953 ;
      RECT 82.075 3.675 82.27 3.95 ;
      RECT 82.065 3.675 82.27 3.948 ;
      RECT 82.01 3.675 82.27 3.935 ;
      RECT 82.01 3.75 82.275 3.913 ;
      RECT 81.54 4.873 81.545 5.08 ;
      RECT 81.49 4.867 81.54 5.079 ;
      RECT 81.457 4.881 81.55 5.078 ;
      RECT 81.371 4.881 81.55 5.077 ;
      RECT 81.285 4.881 81.55 5.076 ;
      RECT 81.285 4.98 81.555 5.073 ;
      RECT 81.28 4.98 81.555 5.068 ;
      RECT 81.275 4.98 81.555 5.05 ;
      RECT 81.27 4.98 81.555 5.033 ;
      RECT 81.23 4.765 81.49 5.025 ;
      RECT 80.69 3.915 80.776 4.329 ;
      RECT 80.69 3.915 80.815 4.326 ;
      RECT 80.69 3.915 80.835 4.316 ;
      RECT 80.645 3.915 80.835 4.313 ;
      RECT 80.645 4.067 80.845 4.303 ;
      RECT 80.645 4.088 80.85 4.297 ;
      RECT 80.645 4.106 80.855 4.293 ;
      RECT 80.645 4.126 80.865 4.288 ;
      RECT 80.62 4.126 80.865 4.285 ;
      RECT 80.61 4.126 80.865 4.263 ;
      RECT 80.61 4.142 80.87 4.233 ;
      RECT 80.575 3.915 80.835 4.22 ;
      RECT 80.575 4.154 80.875 4.175 ;
      RECT 78.235 10.06 78.53 10.29 ;
      RECT 78.295 8.58 78.465 10.29 ;
      RECT 78.245 8.95 78.595 9.3 ;
      RECT 78.235 8.58 78.525 8.81 ;
      RECT 77.245 10.06 77.54 10.29 ;
      RECT 77.305 8.58 77.475 10.29 ;
      RECT 77.245 8.58 77.535 8.81 ;
      RECT 77.245 8.615 78.095 8.775 ;
      RECT 77.93 8.21 78.095 8.775 ;
      RECT 77.245 8.61 77.64 8.775 ;
      RECT 77.865 8.21 78.155 8.44 ;
      RECT 77.865 8.24 78.325 8.41 ;
      RECT 77.83 4.025 78.15 4.26 ;
      RECT 77.83 4.055 78.32 4.225 ;
      RECT 77.83 3.69 78.02 4.26 ;
      RECT 77.245 3.655 77.535 3.885 ;
      RECT 77.245 3.69 78.02 3.86 ;
      RECT 77.305 2.175 77.475 3.885 ;
      RECT 77.245 2.175 77.54 2.405 ;
      RECT 76.875 4.025 77.165 4.255 ;
      RECT 76.875 4.055 77.335 4.225 ;
      RECT 76.94 2.95 77.105 4.255 ;
      RECT 75.455 2.915 75.745 3.145 ;
      RECT 75.455 2.95 77.105 3.12 ;
      RECT 75.515 2.175 75.685 3.145 ;
      RECT 75.455 2.175 75.745 2.405 ;
      RECT 75.455 10.06 75.745 10.29 ;
      RECT 75.515 9.32 75.685 10.29 ;
      RECT 75.515 9.41 77.105 9.58 ;
      RECT 76.935 8.21 77.105 9.58 ;
      RECT 75.455 9.32 75.745 9.55 ;
      RECT 76.875 8.21 77.165 8.44 ;
      RECT 76.875 8.24 77.335 8.41 ;
      RECT 73.505 4 73.845 4.35 ;
      RECT 73.595 3.32 73.765 4.35 ;
      RECT 75.885 3.26 76.235 3.61 ;
      RECT 73.595 3.32 76.235 3.49 ;
      RECT 75.715 3.315 76.235 3.49 ;
      RECT 75.91 8.945 76.235 9.27 ;
      RECT 70.45 8.905 70.8 9.255 ;
      RECT 75.885 8.95 76.235 9.18 ;
      RECT 70.25 8.95 70.8 9.18 ;
      RECT 75.715 8.975 76.235 9.15 ;
      RECT 70.08 8.98 70.8 9.15 ;
      RECT 70.13 8.975 76.235 9.145 ;
      RECT 75.11 3.66 75.43 3.98 ;
      RECT 75.085 3.655 75.375 3.885 ;
      RECT 75.08 3.685 75.43 3.86 ;
      RECT 74.91 3.685 75.43 3.855 ;
      RECT 75.11 8.545 75.43 8.835 ;
      RECT 75.085 8.58 75.43 8.81 ;
      RECT 74.91 8.61 75.43 8.78 ;
      RECT 70.8 4.28 70.95 4.555 ;
      RECT 71.34 3.36 71.345 3.58 ;
      RECT 72.49 3.56 72.505 3.758 ;
      RECT 72.455 3.552 72.49 3.765 ;
      RECT 72.425 3.545 72.455 3.765 ;
      RECT 72.37 3.51 72.425 3.765 ;
      RECT 72.305 3.447 72.37 3.765 ;
      RECT 72.3 3.412 72.305 3.763 ;
      RECT 72.295 3.407 72.3 3.755 ;
      RECT 72.29 3.402 72.295 3.741 ;
      RECT 72.285 3.399 72.29 3.734 ;
      RECT 72.24 3.389 72.285 3.685 ;
      RECT 72.22 3.376 72.24 3.62 ;
      RECT 72.215 3.371 72.22 3.593 ;
      RECT 72.21 3.37 72.215 3.586 ;
      RECT 72.205 3.369 72.21 3.579 ;
      RECT 72.12 3.354 72.205 3.525 ;
      RECT 72.09 3.335 72.12 3.475 ;
      RECT 72.01 3.318 72.09 3.46 ;
      RECT 71.975 3.305 72.01 3.445 ;
      RECT 71.967 3.305 71.975 3.44 ;
      RECT 71.881 3.306 71.967 3.44 ;
      RECT 71.795 3.308 71.881 3.44 ;
      RECT 71.77 3.309 71.795 3.444 ;
      RECT 71.695 3.315 71.77 3.459 ;
      RECT 71.612 3.327 71.695 3.483 ;
      RECT 71.526 3.34 71.612 3.509 ;
      RECT 71.44 3.353 71.526 3.535 ;
      RECT 71.405 3.362 71.44 3.554 ;
      RECT 71.355 3.362 71.405 3.567 ;
      RECT 71.345 3.36 71.355 3.578 ;
      RECT 71.33 3.357 71.34 3.58 ;
      RECT 71.315 3.349 71.33 3.588 ;
      RECT 71.3 3.341 71.315 3.608 ;
      RECT 71.295 3.336 71.3 3.665 ;
      RECT 71.28 3.331 71.295 3.738 ;
      RECT 71.275 3.326 71.28 3.78 ;
      RECT 71.27 3.324 71.275 3.808 ;
      RECT 71.265 3.322 71.27 3.83 ;
      RECT 71.255 3.318 71.265 3.873 ;
      RECT 71.25 3.315 71.255 3.898 ;
      RECT 71.245 3.313 71.25 3.918 ;
      RECT 71.24 3.311 71.245 3.942 ;
      RECT 71.235 3.307 71.24 3.965 ;
      RECT 71.23 3.303 71.235 3.988 ;
      RECT 71.195 3.293 71.23 4.095 ;
      RECT 71.19 3.283 71.195 4.193 ;
      RECT 71.185 3.281 71.19 4.22 ;
      RECT 71.18 3.28 71.185 4.24 ;
      RECT 71.175 3.272 71.18 4.26 ;
      RECT 71.17 3.267 71.175 4.295 ;
      RECT 71.165 3.265 71.17 4.313 ;
      RECT 71.16 3.265 71.165 4.338 ;
      RECT 71.155 3.265 71.16 4.36 ;
      RECT 71.12 3.265 71.155 4.403 ;
      RECT 71.095 3.265 71.12 4.432 ;
      RECT 71.085 3.265 71.095 3.618 ;
      RECT 71.088 3.675 71.095 4.442 ;
      RECT 71.085 3.732 71.088 4.445 ;
      RECT 71.08 3.265 71.085 3.59 ;
      RECT 71.08 3.782 71.085 4.448 ;
      RECT 71.07 3.265 71.08 3.58 ;
      RECT 71.075 3.835 71.08 4.451 ;
      RECT 71.07 3.92 71.075 4.455 ;
      RECT 71.06 3.265 71.07 3.568 ;
      RECT 71.065 3.967 71.07 4.459 ;
      RECT 71.06 4.042 71.065 4.463 ;
      RECT 71.025 3.265 71.06 3.543 ;
      RECT 71.05 4.125 71.06 4.468 ;
      RECT 71.04 4.192 71.05 4.475 ;
      RECT 71.035 4.22 71.04 4.48 ;
      RECT 71.025 4.233 71.035 4.486 ;
      RECT 70.98 3.265 71.025 3.5 ;
      RECT 71.02 4.238 71.025 4.493 ;
      RECT 70.98 4.255 71.02 4.555 ;
      RECT 70.975 3.267 70.98 3.473 ;
      RECT 70.95 4.275 70.98 4.555 ;
      RECT 70.97 3.272 70.975 3.445 ;
      RECT 70.76 4.284 70.8 4.555 ;
      RECT 70.735 4.292 70.76 4.525 ;
      RECT 70.69 4.3 70.735 4.525 ;
      RECT 70.675 4.305 70.69 4.52 ;
      RECT 70.665 4.305 70.675 4.514 ;
      RECT 70.655 4.312 70.665 4.511 ;
      RECT 70.65 4.35 70.655 4.5 ;
      RECT 70.645 4.412 70.65 4.478 ;
      RECT 71.915 4.287 72.1 4.51 ;
      RECT 71.915 4.302 72.105 4.506 ;
      RECT 71.905 3.575 71.99 4.505 ;
      RECT 71.905 4.302 72.11 4.499 ;
      RECT 71.9 4.31 72.11 4.498 ;
      RECT 72.105 4.03 72.425 4.35 ;
      RECT 71.9 4.202 72.07 4.293 ;
      RECT 71.895 4.202 72.07 4.275 ;
      RECT 71.885 4.01 72.02 4.25 ;
      RECT 71.88 4.01 72.02 4.195 ;
      RECT 71.84 3.59 72.01 4.095 ;
      RECT 71.825 3.59 72.01 3.965 ;
      RECT 71.82 3.59 72.01 3.918 ;
      RECT 71.815 3.59 72.01 3.898 ;
      RECT 71.81 3.59 72.01 3.873 ;
      RECT 71.78 3.59 72.04 3.85 ;
      RECT 71.79 3.587 72 3.85 ;
      RECT 71.915 3.582 72 4.51 ;
      RECT 71.8 3.575 71.99 3.85 ;
      RECT 71.795 3.58 71.99 3.85 ;
      RECT 70.625 3.792 70.81 4.005 ;
      RECT 70.625 3.8 70.82 3.998 ;
      RECT 70.605 3.8 70.82 3.995 ;
      RECT 70.6 3.8 70.82 3.98 ;
      RECT 70.53 3.715 70.79 3.975 ;
      RECT 70.53 3.86 70.825 3.888 ;
      RECT 70.185 4.315 70.445 4.575 ;
      RECT 70.21 4.26 70.405 4.575 ;
      RECT 70.205 4.009 70.385 4.303 ;
      RECT 70.205 4.015 70.395 4.303 ;
      RECT 70.185 4.017 70.395 4.248 ;
      RECT 70.18 4.027 70.395 4.115 ;
      RECT 70.21 4.007 70.385 4.575 ;
      RECT 70.296 4.005 70.385 4.575 ;
      RECT 70.155 3.225 70.19 3.595 ;
      RECT 69.945 3.335 69.95 3.595 ;
      RECT 70.19 3.232 70.205 3.595 ;
      RECT 70.08 3.225 70.155 3.673 ;
      RECT 70.07 3.225 70.08 3.758 ;
      RECT 70.045 3.225 70.07 3.793 ;
      RECT 70.005 3.225 70.045 3.861 ;
      RECT 69.995 3.232 70.005 3.913 ;
      RECT 69.965 3.335 69.995 3.954 ;
      RECT 69.96 3.335 69.965 3.993 ;
      RECT 69.95 3.335 69.96 4.013 ;
      RECT 69.945 3.63 69.95 4.05 ;
      RECT 69.94 3.647 69.945 4.07 ;
      RECT 69.925 3.71 69.94 4.11 ;
      RECT 69.92 3.753 69.925 4.145 ;
      RECT 69.915 3.761 69.92 4.158 ;
      RECT 69.905 3.775 69.915 4.18 ;
      RECT 69.88 3.81 69.905 4.245 ;
      RECT 69.87 3.845 69.88 4.308 ;
      RECT 69.85 3.875 69.87 4.369 ;
      RECT 69.835 3.911 69.85 4.436 ;
      RECT 69.825 3.939 69.835 4.475 ;
      RECT 69.815 3.961 69.825 4.495 ;
      RECT 69.81 3.971 69.815 4.506 ;
      RECT 69.805 3.98 69.81 4.509 ;
      RECT 69.795 3.998 69.805 4.513 ;
      RECT 69.785 4.016 69.795 4.514 ;
      RECT 69.76 4.055 69.785 4.511 ;
      RECT 69.74 4.097 69.76 4.508 ;
      RECT 69.725 4.135 69.74 4.507 ;
      RECT 69.69 4.17 69.725 4.504 ;
      RECT 69.685 4.192 69.69 4.502 ;
      RECT 69.62 4.232 69.685 4.499 ;
      RECT 69.615 4.272 69.62 4.495 ;
      RECT 69.6 4.282 69.615 4.486 ;
      RECT 69.59 4.402 69.6 4.471 ;
      RECT 70.07 4.815 70.08 5.075 ;
      RECT 70.07 4.818 70.09 5.074 ;
      RECT 70.06 4.808 70.07 5.073 ;
      RECT 70.05 4.823 70.13 5.069 ;
      RECT 70.035 4.802 70.05 5.067 ;
      RECT 70.01 4.827 70.135 5.063 ;
      RECT 69.995 4.787 70.01 5.058 ;
      RECT 69.995 4.829 70.145 5.057 ;
      RECT 69.995 4.837 70.16 5.05 ;
      RECT 69.935 4.774 69.995 5.04 ;
      RECT 69.925 4.761 69.935 5.022 ;
      RECT 69.9 4.751 69.925 5.012 ;
      RECT 69.895 4.741 69.9 5.004 ;
      RECT 69.83 4.837 70.16 4.986 ;
      RECT 69.745 4.837 70.16 4.948 ;
      RECT 69.635 4.665 69.895 4.925 ;
      RECT 70.01 4.795 70.035 5.063 ;
      RECT 70.05 4.805 70.06 5.069 ;
      RECT 69.635 4.813 70.075 4.925 ;
      RECT 69.82 10.06 70.11 10.29 ;
      RECT 69.88 9.32 70.05 10.29 ;
      RECT 69.78 9.345 70.15 9.715 ;
      RECT 69.82 9.32 70.11 9.715 ;
      RECT 68.85 4.57 68.88 4.87 ;
      RECT 68.625 4.555 68.63 4.83 ;
      RECT 68.425 4.555 68.58 4.815 ;
      RECT 69.725 3.27 69.755 3.53 ;
      RECT 69.715 3.27 69.725 3.638 ;
      RECT 69.695 3.27 69.715 3.648 ;
      RECT 69.68 3.27 69.695 3.66 ;
      RECT 69.625 3.27 69.68 3.71 ;
      RECT 69.61 3.27 69.625 3.758 ;
      RECT 69.58 3.27 69.61 3.793 ;
      RECT 69.525 3.27 69.58 3.855 ;
      RECT 69.505 3.27 69.525 3.923 ;
      RECT 69.5 3.27 69.505 3.953 ;
      RECT 69.495 3.27 69.5 3.965 ;
      RECT 69.49 3.387 69.495 3.983 ;
      RECT 69.47 3.405 69.49 4.008 ;
      RECT 69.45 3.432 69.47 4.058 ;
      RECT 69.445 3.452 69.45 4.089 ;
      RECT 69.44 3.46 69.445 4.106 ;
      RECT 69.425 3.486 69.44 4.135 ;
      RECT 69.41 3.528 69.425 4.17 ;
      RECT 69.405 3.557 69.41 4.193 ;
      RECT 69.4 3.572 69.405 4.206 ;
      RECT 69.395 3.595 69.4 4.217 ;
      RECT 69.385 3.615 69.395 4.235 ;
      RECT 69.375 3.645 69.385 4.258 ;
      RECT 69.37 3.667 69.375 4.278 ;
      RECT 69.365 3.682 69.37 4.293 ;
      RECT 69.35 3.712 69.365 4.32 ;
      RECT 69.345 3.742 69.35 4.346 ;
      RECT 69.34 3.76 69.345 4.358 ;
      RECT 69.33 3.79 69.34 4.377 ;
      RECT 69.32 3.815 69.33 4.402 ;
      RECT 69.315 3.835 69.32 4.421 ;
      RECT 69.31 3.852 69.315 4.434 ;
      RECT 69.3 3.878 69.31 4.453 ;
      RECT 69.29 3.916 69.3 4.48 ;
      RECT 69.285 3.942 69.29 4.5 ;
      RECT 69.28 3.952 69.285 4.51 ;
      RECT 69.275 3.965 69.28 4.525 ;
      RECT 69.27 3.98 69.275 4.535 ;
      RECT 69.265 4.002 69.27 4.55 ;
      RECT 69.26 4.02 69.265 4.561 ;
      RECT 69.255 4.03 69.26 4.572 ;
      RECT 69.25 4.038 69.255 4.584 ;
      RECT 69.245 4.046 69.25 4.595 ;
      RECT 69.24 4.072 69.245 4.608 ;
      RECT 69.23 4.1 69.24 4.621 ;
      RECT 69.225 4.13 69.23 4.63 ;
      RECT 69.22 4.145 69.225 4.637 ;
      RECT 69.205 4.17 69.22 4.644 ;
      RECT 69.2 4.192 69.205 4.65 ;
      RECT 69.195 4.217 69.2 4.653 ;
      RECT 69.186 4.245 69.195 4.657 ;
      RECT 69.18 4.262 69.186 4.662 ;
      RECT 69.175 4.28 69.18 4.666 ;
      RECT 69.17 4.292 69.175 4.669 ;
      RECT 69.165 4.313 69.17 4.673 ;
      RECT 69.16 4.331 69.165 4.676 ;
      RECT 69.155 4.345 69.16 4.679 ;
      RECT 69.15 4.362 69.155 4.682 ;
      RECT 69.145 4.375 69.15 4.685 ;
      RECT 69.12 4.412 69.145 4.693 ;
      RECT 69.115 4.457 69.12 4.702 ;
      RECT 69.11 4.485 69.115 4.705 ;
      RECT 69.1 4.505 69.11 4.709 ;
      RECT 69.095 4.525 69.1 4.714 ;
      RECT 69.09 4.54 69.095 4.717 ;
      RECT 69.07 4.55 69.09 4.724 ;
      RECT 69.005 4.557 69.07 4.75 ;
      RECT 68.97 4.56 69.005 4.778 ;
      RECT 68.955 4.563 68.97 4.793 ;
      RECT 68.945 4.564 68.955 4.808 ;
      RECT 68.935 4.565 68.945 4.825 ;
      RECT 68.93 4.565 68.935 4.84 ;
      RECT 68.925 4.565 68.93 4.848 ;
      RECT 68.91 4.566 68.925 4.863 ;
      RECT 68.88 4.568 68.91 4.87 ;
      RECT 68.77 4.575 68.85 4.87 ;
      RECT 68.725 4.58 68.77 4.87 ;
      RECT 68.715 4.581 68.725 4.86 ;
      RECT 68.705 4.582 68.715 4.853 ;
      RECT 68.685 4.584 68.705 4.848 ;
      RECT 68.675 4.555 68.685 4.843 ;
      RECT 68.63 4.555 68.675 4.835 ;
      RECT 68.6 4.555 68.625 4.825 ;
      RECT 68.58 4.555 68.6 4.818 ;
      RECT 68.86 3.355 69.12 3.615 ;
      RECT 68.74 3.37 68.75 3.535 ;
      RECT 68.725 3.37 68.73 3.53 ;
      RECT 66.09 3.21 66.275 3.5 ;
      RECT 67.905 3.335 67.92 3.49 ;
      RECT 66.055 3.21 66.08 3.47 ;
      RECT 68.47 3.26 68.475 3.402 ;
      RECT 68.385 3.255 68.41 3.395 ;
      RECT 68.785 3.372 68.86 3.565 ;
      RECT 68.77 3.37 68.785 3.548 ;
      RECT 68.75 3.37 68.77 3.54 ;
      RECT 68.73 3.37 68.74 3.533 ;
      RECT 68.685 3.365 68.725 3.523 ;
      RECT 68.645 3.34 68.685 3.508 ;
      RECT 68.63 3.315 68.645 3.498 ;
      RECT 68.625 3.309 68.63 3.496 ;
      RECT 68.59 3.301 68.625 3.479 ;
      RECT 68.585 3.294 68.59 3.467 ;
      RECT 68.565 3.289 68.585 3.455 ;
      RECT 68.555 3.283 68.565 3.44 ;
      RECT 68.535 3.278 68.555 3.425 ;
      RECT 68.525 3.273 68.535 3.418 ;
      RECT 68.52 3.271 68.525 3.413 ;
      RECT 68.515 3.27 68.52 3.41 ;
      RECT 68.475 3.265 68.515 3.406 ;
      RECT 68.455 3.259 68.47 3.401 ;
      RECT 68.42 3.256 68.455 3.398 ;
      RECT 68.41 3.255 68.42 3.396 ;
      RECT 68.35 3.255 68.385 3.393 ;
      RECT 68.305 3.255 68.35 3.393 ;
      RECT 68.255 3.255 68.305 3.396 ;
      RECT 68.24 3.257 68.255 3.398 ;
      RECT 68.225 3.26 68.24 3.399 ;
      RECT 68.215 3.265 68.225 3.4 ;
      RECT 68.185 3.27 68.215 3.405 ;
      RECT 68.175 3.276 68.185 3.413 ;
      RECT 68.165 3.278 68.175 3.417 ;
      RECT 68.155 3.282 68.165 3.421 ;
      RECT 68.13 3.288 68.155 3.429 ;
      RECT 68.12 3.293 68.13 3.437 ;
      RECT 68.105 3.297 68.12 3.441 ;
      RECT 68.07 3.303 68.105 3.449 ;
      RECT 68.05 3.308 68.07 3.459 ;
      RECT 68.02 3.315 68.05 3.468 ;
      RECT 67.975 3.324 68.02 3.482 ;
      RECT 67.97 3.329 67.975 3.493 ;
      RECT 67.95 3.332 67.97 3.494 ;
      RECT 67.92 3.335 67.95 3.492 ;
      RECT 67.885 3.335 67.905 3.488 ;
      RECT 67.815 3.335 67.885 3.479 ;
      RECT 67.8 3.332 67.815 3.471 ;
      RECT 67.76 3.325 67.8 3.466 ;
      RECT 67.735 3.315 67.76 3.459 ;
      RECT 67.73 3.309 67.735 3.456 ;
      RECT 67.69 3.303 67.73 3.453 ;
      RECT 67.675 3.296 67.69 3.448 ;
      RECT 67.655 3.292 67.675 3.443 ;
      RECT 67.64 3.287 67.655 3.439 ;
      RECT 67.625 3.282 67.64 3.437 ;
      RECT 67.61 3.278 67.625 3.436 ;
      RECT 67.595 3.276 67.61 3.432 ;
      RECT 67.585 3.274 67.595 3.427 ;
      RECT 67.57 3.271 67.585 3.423 ;
      RECT 67.56 3.269 67.57 3.418 ;
      RECT 67.54 3.266 67.56 3.414 ;
      RECT 67.495 3.265 67.54 3.412 ;
      RECT 67.435 3.267 67.495 3.413 ;
      RECT 67.415 3.269 67.435 3.415 ;
      RECT 67.385 3.272 67.415 3.416 ;
      RECT 67.335 3.277 67.385 3.418 ;
      RECT 67.33 3.28 67.335 3.42 ;
      RECT 67.32 3.282 67.33 3.423 ;
      RECT 67.315 3.284 67.32 3.426 ;
      RECT 67.265 3.287 67.315 3.433 ;
      RECT 67.245 3.291 67.265 3.445 ;
      RECT 67.235 3.294 67.245 3.451 ;
      RECT 67.225 3.295 67.235 3.454 ;
      RECT 67.186 3.298 67.225 3.456 ;
      RECT 67.1 3.305 67.186 3.459 ;
      RECT 67.026 3.315 67.1 3.463 ;
      RECT 66.94 3.326 67.026 3.468 ;
      RECT 66.925 3.333 66.94 3.47 ;
      RECT 66.87 3.337 66.925 3.471 ;
      RECT 66.856 3.34 66.87 3.473 ;
      RECT 66.77 3.34 66.856 3.475 ;
      RECT 66.73 3.337 66.77 3.478 ;
      RECT 66.706 3.333 66.73 3.48 ;
      RECT 66.62 3.323 66.706 3.483 ;
      RECT 66.59 3.312 66.62 3.484 ;
      RECT 66.571 3.308 66.59 3.483 ;
      RECT 66.485 3.301 66.571 3.48 ;
      RECT 66.425 3.29 66.485 3.477 ;
      RECT 66.405 3.282 66.425 3.475 ;
      RECT 66.37 3.277 66.405 3.474 ;
      RECT 66.345 3.272 66.37 3.473 ;
      RECT 66.315 3.267 66.345 3.472 ;
      RECT 66.29 3.21 66.315 3.471 ;
      RECT 66.275 3.21 66.29 3.495 ;
      RECT 66.08 3.21 66.09 3.495 ;
      RECT 67.855 4.23 67.86 4.37 ;
      RECT 67.515 4.23 67.55 4.368 ;
      RECT 67.09 4.215 67.105 4.36 ;
      RECT 68.92 3.995 69.01 4.255 ;
      RECT 68.75 3.86 68.85 4.255 ;
      RECT 65.785 3.835 65.865 4.045 ;
      RECT 68.875 3.972 68.92 4.255 ;
      RECT 68.865 3.942 68.875 4.255 ;
      RECT 68.85 3.865 68.865 4.255 ;
      RECT 68.665 3.86 68.75 4.22 ;
      RECT 68.66 3.862 68.665 4.215 ;
      RECT 68.655 3.867 68.66 4.215 ;
      RECT 68.62 3.967 68.655 4.215 ;
      RECT 68.61 3.995 68.62 4.215 ;
      RECT 68.6 4.01 68.61 4.215 ;
      RECT 68.59 4.022 68.6 4.215 ;
      RECT 68.585 4.032 68.59 4.215 ;
      RECT 68.57 4.042 68.585 4.217 ;
      RECT 68.565 4.057 68.57 4.219 ;
      RECT 68.55 4.07 68.565 4.221 ;
      RECT 68.545 4.085 68.55 4.224 ;
      RECT 68.525 4.095 68.545 4.228 ;
      RECT 68.51 4.105 68.525 4.231 ;
      RECT 68.475 4.112 68.51 4.236 ;
      RECT 68.431 4.119 68.475 4.244 ;
      RECT 68.345 4.131 68.431 4.257 ;
      RECT 68.32 4.142 68.345 4.268 ;
      RECT 68.29 4.147 68.32 4.273 ;
      RECT 68.255 4.152 68.29 4.281 ;
      RECT 68.225 4.157 68.255 4.288 ;
      RECT 68.2 4.162 68.225 4.293 ;
      RECT 68.135 4.169 68.2 4.302 ;
      RECT 68.065 4.182 68.135 4.318 ;
      RECT 68.035 4.192 68.065 4.33 ;
      RECT 68.01 4.197 68.035 4.337 ;
      RECT 67.955 4.204 68.01 4.345 ;
      RECT 67.95 4.211 67.955 4.35 ;
      RECT 67.945 4.213 67.95 4.351 ;
      RECT 67.93 4.215 67.945 4.353 ;
      RECT 67.925 4.215 67.93 4.356 ;
      RECT 67.86 4.222 67.925 4.363 ;
      RECT 67.825 4.232 67.855 4.373 ;
      RECT 67.808 4.235 67.825 4.375 ;
      RECT 67.722 4.234 67.808 4.374 ;
      RECT 67.636 4.232 67.722 4.371 ;
      RECT 67.55 4.231 67.636 4.369 ;
      RECT 67.449 4.229 67.515 4.368 ;
      RECT 67.363 4.226 67.449 4.366 ;
      RECT 67.277 4.222 67.363 4.364 ;
      RECT 67.191 4.219 67.277 4.363 ;
      RECT 67.105 4.216 67.191 4.361 ;
      RECT 67.005 4.215 67.09 4.358 ;
      RECT 66.955 4.213 67.005 4.356 ;
      RECT 66.935 4.21 66.955 4.354 ;
      RECT 66.915 4.208 66.935 4.351 ;
      RECT 66.89 4.204 66.915 4.348 ;
      RECT 66.845 4.198 66.89 4.343 ;
      RECT 66.805 4.192 66.845 4.335 ;
      RECT 66.78 4.187 66.805 4.328 ;
      RECT 66.725 4.18 66.78 4.32 ;
      RECT 66.701 4.173 66.725 4.313 ;
      RECT 66.615 4.164 66.701 4.303 ;
      RECT 66.585 4.156 66.615 4.293 ;
      RECT 66.555 4.152 66.585 4.288 ;
      RECT 66.55 4.149 66.555 4.285 ;
      RECT 66.545 4.148 66.55 4.285 ;
      RECT 66.47 4.141 66.545 4.278 ;
      RECT 66.431 4.132 66.47 4.267 ;
      RECT 66.345 4.122 66.431 4.255 ;
      RECT 66.305 4.112 66.345 4.243 ;
      RECT 66.266 4.107 66.305 4.236 ;
      RECT 66.18 4.097 66.266 4.225 ;
      RECT 66.14 4.085 66.18 4.214 ;
      RECT 66.105 4.07 66.14 4.207 ;
      RECT 66.095 4.06 66.105 4.204 ;
      RECT 66.075 4.045 66.095 4.202 ;
      RECT 66.045 4.015 66.075 4.198 ;
      RECT 66.035 3.995 66.045 4.193 ;
      RECT 66.03 3.987 66.035 4.19 ;
      RECT 66.025 3.98 66.03 4.188 ;
      RECT 66.01 3.967 66.025 4.181 ;
      RECT 66.005 3.957 66.01 4.173 ;
      RECT 66 3.95 66.005 4.168 ;
      RECT 65.995 3.945 66 4.164 ;
      RECT 65.98 3.932 65.995 4.156 ;
      RECT 65.975 3.842 65.98 4.145 ;
      RECT 65.97 3.837 65.975 4.138 ;
      RECT 65.895 3.835 65.97 4.098 ;
      RECT 65.865 3.835 65.895 4.053 ;
      RECT 65.77 3.84 65.785 4.04 ;
      RECT 68.255 3.545 68.515 3.805 ;
      RECT 68.24 3.533 68.42 3.77 ;
      RECT 68.235 3.534 68.42 3.768 ;
      RECT 68.22 3.538 68.43 3.758 ;
      RECT 68.215 3.543 68.435 3.728 ;
      RECT 68.22 3.54 68.435 3.758 ;
      RECT 68.235 3.535 68.43 3.768 ;
      RECT 68.255 3.532 68.42 3.805 ;
      RECT 68.255 3.531 68.41 3.805 ;
      RECT 68.28 3.53 68.41 3.805 ;
      RECT 67.84 3.775 68.1 4.035 ;
      RECT 67.715 3.82 68.1 4.03 ;
      RECT 67.705 3.825 68.1 4.025 ;
      RECT 67.72 4.765 67.735 5.075 ;
      RECT 66.315 4.535 66.325 4.665 ;
      RECT 66.095 4.53 66.2 4.665 ;
      RECT 66.01 4.535 66.06 4.665 ;
      RECT 64.56 3.27 64.565 4.375 ;
      RECT 67.815 4.857 67.82 4.993 ;
      RECT 67.81 4.852 67.815 5.053 ;
      RECT 67.805 4.85 67.81 5.066 ;
      RECT 67.79 4.847 67.805 5.068 ;
      RECT 67.785 4.842 67.79 5.07 ;
      RECT 67.78 4.838 67.785 5.073 ;
      RECT 67.765 4.833 67.78 5.075 ;
      RECT 67.735 4.825 67.765 5.075 ;
      RECT 67.696 4.765 67.72 5.075 ;
      RECT 67.61 4.765 67.696 5.072 ;
      RECT 67.58 4.765 67.61 5.065 ;
      RECT 67.555 4.765 67.58 5.058 ;
      RECT 67.53 4.765 67.555 5.05 ;
      RECT 67.515 4.765 67.53 5.043 ;
      RECT 67.49 4.765 67.515 5.035 ;
      RECT 67.475 4.765 67.49 5.028 ;
      RECT 67.435 4.775 67.475 5.017 ;
      RECT 67.425 4.77 67.435 5.007 ;
      RECT 67.421 4.769 67.425 5.004 ;
      RECT 67.335 4.761 67.421 4.987 ;
      RECT 67.302 4.75 67.335 4.964 ;
      RECT 67.216 4.739 67.302 4.942 ;
      RECT 67.13 4.723 67.216 4.911 ;
      RECT 67.06 4.708 67.13 4.883 ;
      RECT 67.05 4.701 67.06 4.87 ;
      RECT 67.02 4.698 67.05 4.86 ;
      RECT 66.995 4.694 67.02 4.853 ;
      RECT 66.98 4.691 66.995 4.848 ;
      RECT 66.975 4.69 66.98 4.843 ;
      RECT 66.945 4.685 66.975 4.836 ;
      RECT 66.94 4.68 66.945 4.831 ;
      RECT 66.925 4.677 66.94 4.826 ;
      RECT 66.92 4.672 66.925 4.821 ;
      RECT 66.9 4.667 66.92 4.818 ;
      RECT 66.885 4.662 66.9 4.81 ;
      RECT 66.87 4.656 66.885 4.805 ;
      RECT 66.84 4.647 66.87 4.798 ;
      RECT 66.835 4.64 66.84 4.79 ;
      RECT 66.83 4.638 66.835 4.788 ;
      RECT 66.825 4.637 66.83 4.785 ;
      RECT 66.785 4.63 66.825 4.778 ;
      RECT 66.771 4.62 66.785 4.768 ;
      RECT 66.72 4.609 66.771 4.756 ;
      RECT 66.695 4.595 66.72 4.742 ;
      RECT 66.67 4.584 66.695 4.734 ;
      RECT 66.65 4.573 66.67 4.728 ;
      RECT 66.64 4.567 66.65 4.723 ;
      RECT 66.635 4.565 66.64 4.719 ;
      RECT 66.615 4.56 66.635 4.714 ;
      RECT 66.585 4.55 66.615 4.704 ;
      RECT 66.58 4.542 66.585 4.697 ;
      RECT 66.565 4.54 66.58 4.693 ;
      RECT 66.545 4.54 66.565 4.688 ;
      RECT 66.54 4.539 66.545 4.686 ;
      RECT 66.535 4.539 66.54 4.683 ;
      RECT 66.495 4.538 66.535 4.678 ;
      RECT 66.47 4.537 66.495 4.673 ;
      RECT 66.41 4.536 66.47 4.67 ;
      RECT 66.325 4.535 66.41 4.668 ;
      RECT 66.286 4.534 66.315 4.665 ;
      RECT 66.2 4.532 66.286 4.665 ;
      RECT 66.06 4.532 66.095 4.665 ;
      RECT 65.97 4.536 66.01 4.668 ;
      RECT 65.955 4.539 65.97 4.675 ;
      RECT 65.945 4.54 65.955 4.682 ;
      RECT 65.92 4.543 65.945 4.687 ;
      RECT 65.915 4.545 65.92 4.69 ;
      RECT 65.865 4.547 65.915 4.691 ;
      RECT 65.826 4.551 65.865 4.693 ;
      RECT 65.74 4.553 65.826 4.696 ;
      RECT 65.722 4.555 65.74 4.698 ;
      RECT 65.636 4.558 65.722 4.7 ;
      RECT 65.55 4.562 65.636 4.703 ;
      RECT 65.513 4.566 65.55 4.706 ;
      RECT 65.427 4.569 65.513 4.709 ;
      RECT 65.341 4.573 65.427 4.712 ;
      RECT 65.255 4.578 65.341 4.716 ;
      RECT 65.235 4.58 65.255 4.719 ;
      RECT 65.215 4.579 65.235 4.72 ;
      RECT 65.166 4.576 65.215 4.721 ;
      RECT 65.08 4.571 65.166 4.724 ;
      RECT 65.03 4.566 65.08 4.726 ;
      RECT 65.006 4.564 65.03 4.727 ;
      RECT 64.92 4.559 65.006 4.729 ;
      RECT 64.895 4.555 64.92 4.728 ;
      RECT 64.885 4.552 64.895 4.726 ;
      RECT 64.875 4.545 64.885 4.723 ;
      RECT 64.87 4.525 64.875 4.718 ;
      RECT 64.86 4.495 64.87 4.713 ;
      RECT 64.845 4.365 64.86 4.704 ;
      RECT 64.84 4.357 64.845 4.697 ;
      RECT 64.82 4.35 64.84 4.689 ;
      RECT 64.815 4.332 64.82 4.681 ;
      RECT 64.805 4.312 64.815 4.676 ;
      RECT 64.8 4.285 64.805 4.672 ;
      RECT 64.795 4.262 64.8 4.669 ;
      RECT 64.775 4.22 64.795 4.661 ;
      RECT 64.74 4.135 64.775 4.645 ;
      RECT 64.735 4.067 64.74 4.633 ;
      RECT 64.72 4.037 64.735 4.627 ;
      RECT 64.715 3.282 64.72 3.528 ;
      RECT 64.705 4.007 64.72 4.618 ;
      RECT 64.71 3.277 64.715 3.56 ;
      RECT 64.705 3.272 64.71 3.603 ;
      RECT 64.7 3.27 64.705 3.638 ;
      RECT 64.685 3.97 64.705 4.608 ;
      RECT 64.695 3.27 64.7 3.675 ;
      RECT 64.68 3.27 64.695 3.773 ;
      RECT 64.68 3.943 64.685 4.601 ;
      RECT 64.675 3.27 64.68 3.848 ;
      RECT 64.675 3.931 64.68 4.598 ;
      RECT 64.67 3.27 64.675 3.88 ;
      RECT 64.67 3.91 64.675 4.595 ;
      RECT 64.665 3.27 64.67 4.592 ;
      RECT 64.63 3.27 64.665 4.578 ;
      RECT 64.615 3.27 64.63 4.56 ;
      RECT 64.595 3.27 64.615 4.55 ;
      RECT 64.57 3.27 64.595 4.533 ;
      RECT 64.565 3.27 64.57 4.483 ;
      RECT 64.555 3.27 64.56 4.313 ;
      RECT 64.55 3.27 64.555 4.22 ;
      RECT 64.545 3.27 64.55 4.133 ;
      RECT 64.54 3.27 64.545 4.065 ;
      RECT 64.535 3.27 64.54 4.008 ;
      RECT 64.525 3.27 64.535 3.903 ;
      RECT 64.52 3.27 64.525 3.775 ;
      RECT 64.515 3.27 64.52 3.693 ;
      RECT 64.51 3.272 64.515 3.61 ;
      RECT 64.505 3.277 64.51 3.543 ;
      RECT 64.5 3.282 64.505 3.47 ;
      RECT 67.315 3.6 67.575 3.86 ;
      RECT 67.335 3.567 67.545 3.86 ;
      RECT 67.335 3.565 67.535 3.86 ;
      RECT 67.345 3.552 67.535 3.86 ;
      RECT 67.345 3.55 67.46 3.86 ;
      RECT 66.82 3.675 66.995 3.955 ;
      RECT 66.815 3.675 66.995 3.953 ;
      RECT 66.815 3.675 67.01 3.95 ;
      RECT 66.805 3.675 67.01 3.948 ;
      RECT 66.75 3.675 67.01 3.935 ;
      RECT 66.75 3.75 67.015 3.913 ;
      RECT 66.28 4.873 66.285 5.08 ;
      RECT 66.23 4.867 66.28 5.079 ;
      RECT 66.197 4.881 66.29 5.078 ;
      RECT 66.111 4.881 66.29 5.077 ;
      RECT 66.025 4.881 66.29 5.076 ;
      RECT 66.025 4.98 66.295 5.073 ;
      RECT 66.02 4.98 66.295 5.068 ;
      RECT 66.015 4.98 66.295 5.05 ;
      RECT 66.01 4.98 66.295 5.033 ;
      RECT 65.97 4.765 66.23 5.025 ;
      RECT 65.43 3.915 65.516 4.329 ;
      RECT 65.43 3.915 65.555 4.326 ;
      RECT 65.43 3.915 65.575 4.316 ;
      RECT 65.385 3.915 65.575 4.313 ;
      RECT 65.385 4.067 65.585 4.303 ;
      RECT 65.385 4.088 65.59 4.297 ;
      RECT 65.385 4.106 65.595 4.293 ;
      RECT 65.385 4.126 65.605 4.288 ;
      RECT 65.36 4.126 65.605 4.285 ;
      RECT 65.35 4.126 65.605 4.263 ;
      RECT 65.35 4.142 65.61 4.233 ;
      RECT 65.315 3.915 65.575 4.22 ;
      RECT 65.315 4.154 65.615 4.175 ;
      RECT 62.975 10.06 63.27 10.29 ;
      RECT 63.035 8.58 63.205 10.29 ;
      RECT 62.985 8.95 63.335 9.3 ;
      RECT 62.975 8.58 63.265 8.81 ;
      RECT 61.985 10.06 62.28 10.29 ;
      RECT 62.045 8.58 62.215 10.29 ;
      RECT 61.985 8.58 62.275 8.81 ;
      RECT 61.985 8.615 62.835 8.775 ;
      RECT 62.67 8.21 62.835 8.775 ;
      RECT 61.985 8.61 62.38 8.775 ;
      RECT 62.605 8.21 62.895 8.44 ;
      RECT 62.605 8.24 63.065 8.41 ;
      RECT 62.57 4.025 62.89 4.26 ;
      RECT 62.57 4.055 63.06 4.225 ;
      RECT 62.57 3.69 62.76 4.26 ;
      RECT 61.985 3.655 62.275 3.885 ;
      RECT 61.985 3.69 62.76 3.86 ;
      RECT 62.045 2.175 62.215 3.885 ;
      RECT 61.985 2.175 62.28 2.405 ;
      RECT 61.615 4.025 61.905 4.255 ;
      RECT 61.615 4.055 62.075 4.225 ;
      RECT 61.68 2.95 61.845 4.255 ;
      RECT 60.195 2.915 60.485 3.145 ;
      RECT 60.195 2.95 61.845 3.12 ;
      RECT 60.255 2.175 60.425 3.145 ;
      RECT 60.195 2.175 60.485 2.405 ;
      RECT 60.195 10.06 60.485 10.29 ;
      RECT 60.255 9.32 60.425 10.29 ;
      RECT 60.255 9.41 61.845 9.58 ;
      RECT 61.675 8.21 61.845 9.58 ;
      RECT 60.195 9.32 60.485 9.55 ;
      RECT 61.615 8.21 61.905 8.44 ;
      RECT 61.615 8.24 62.075 8.41 ;
      RECT 58.245 4 58.585 4.35 ;
      RECT 58.335 3.32 58.505 4.35 ;
      RECT 60.625 3.26 60.975 3.61 ;
      RECT 58.335 3.32 60.975 3.49 ;
      RECT 60.455 3.315 60.975 3.49 ;
      RECT 60.65 8.945 60.975 9.27 ;
      RECT 55.19 8.905 55.54 9.255 ;
      RECT 60.625 8.95 60.975 9.18 ;
      RECT 54.99 8.95 55.54 9.18 ;
      RECT 60.455 8.975 60.975 9.15 ;
      RECT 54.82 8.98 55.54 9.15 ;
      RECT 54.87 8.975 60.975 9.145 ;
      RECT 59.85 3.66 60.17 3.98 ;
      RECT 59.825 3.655 60.115 3.885 ;
      RECT 59.82 3.685 60.17 3.86 ;
      RECT 59.65 3.685 60.17 3.855 ;
      RECT 59.85 8.545 60.17 8.835 ;
      RECT 59.825 8.58 60.17 8.81 ;
      RECT 59.65 8.61 60.17 8.78 ;
      RECT 55.54 4.28 55.69 4.555 ;
      RECT 56.08 3.36 56.085 3.58 ;
      RECT 57.23 3.56 57.245 3.758 ;
      RECT 57.195 3.552 57.23 3.765 ;
      RECT 57.165 3.545 57.195 3.765 ;
      RECT 57.11 3.51 57.165 3.765 ;
      RECT 57.045 3.447 57.11 3.765 ;
      RECT 57.04 3.412 57.045 3.763 ;
      RECT 57.035 3.407 57.04 3.755 ;
      RECT 57.03 3.402 57.035 3.741 ;
      RECT 57.025 3.399 57.03 3.734 ;
      RECT 56.98 3.389 57.025 3.685 ;
      RECT 56.96 3.376 56.98 3.62 ;
      RECT 56.955 3.371 56.96 3.593 ;
      RECT 56.95 3.37 56.955 3.586 ;
      RECT 56.945 3.369 56.95 3.579 ;
      RECT 56.86 3.354 56.945 3.525 ;
      RECT 56.83 3.335 56.86 3.475 ;
      RECT 56.75 3.318 56.83 3.46 ;
      RECT 56.715 3.305 56.75 3.445 ;
      RECT 56.707 3.305 56.715 3.44 ;
      RECT 56.621 3.306 56.707 3.44 ;
      RECT 56.535 3.308 56.621 3.44 ;
      RECT 56.51 3.309 56.535 3.444 ;
      RECT 56.435 3.315 56.51 3.459 ;
      RECT 56.352 3.327 56.435 3.483 ;
      RECT 56.266 3.34 56.352 3.509 ;
      RECT 56.18 3.353 56.266 3.535 ;
      RECT 56.145 3.362 56.18 3.554 ;
      RECT 56.095 3.362 56.145 3.567 ;
      RECT 56.085 3.36 56.095 3.578 ;
      RECT 56.07 3.357 56.08 3.58 ;
      RECT 56.055 3.349 56.07 3.588 ;
      RECT 56.04 3.341 56.055 3.608 ;
      RECT 56.035 3.336 56.04 3.665 ;
      RECT 56.02 3.331 56.035 3.738 ;
      RECT 56.015 3.326 56.02 3.78 ;
      RECT 56.01 3.324 56.015 3.808 ;
      RECT 56.005 3.322 56.01 3.83 ;
      RECT 55.995 3.318 56.005 3.873 ;
      RECT 55.99 3.315 55.995 3.898 ;
      RECT 55.985 3.313 55.99 3.918 ;
      RECT 55.98 3.311 55.985 3.942 ;
      RECT 55.975 3.307 55.98 3.965 ;
      RECT 55.97 3.303 55.975 3.988 ;
      RECT 55.935 3.293 55.97 4.095 ;
      RECT 55.93 3.283 55.935 4.193 ;
      RECT 55.925 3.281 55.93 4.22 ;
      RECT 55.92 3.28 55.925 4.24 ;
      RECT 55.915 3.272 55.92 4.26 ;
      RECT 55.91 3.267 55.915 4.295 ;
      RECT 55.905 3.265 55.91 4.313 ;
      RECT 55.9 3.265 55.905 4.338 ;
      RECT 55.895 3.265 55.9 4.36 ;
      RECT 55.86 3.265 55.895 4.403 ;
      RECT 55.835 3.265 55.86 4.432 ;
      RECT 55.825 3.265 55.835 3.618 ;
      RECT 55.828 3.675 55.835 4.442 ;
      RECT 55.825 3.732 55.828 4.445 ;
      RECT 55.82 3.265 55.825 3.59 ;
      RECT 55.82 3.782 55.825 4.448 ;
      RECT 55.81 3.265 55.82 3.58 ;
      RECT 55.815 3.835 55.82 4.451 ;
      RECT 55.81 3.92 55.815 4.455 ;
      RECT 55.8 3.265 55.81 3.568 ;
      RECT 55.805 3.967 55.81 4.459 ;
      RECT 55.8 4.042 55.805 4.463 ;
      RECT 55.765 3.265 55.8 3.543 ;
      RECT 55.79 4.125 55.8 4.468 ;
      RECT 55.78 4.192 55.79 4.475 ;
      RECT 55.775 4.22 55.78 4.48 ;
      RECT 55.765 4.233 55.775 4.486 ;
      RECT 55.72 3.265 55.765 3.5 ;
      RECT 55.76 4.238 55.765 4.493 ;
      RECT 55.72 4.255 55.76 4.555 ;
      RECT 55.715 3.267 55.72 3.473 ;
      RECT 55.69 4.275 55.72 4.555 ;
      RECT 55.71 3.272 55.715 3.445 ;
      RECT 55.5 4.284 55.54 4.555 ;
      RECT 55.475 4.292 55.5 4.525 ;
      RECT 55.43 4.3 55.475 4.525 ;
      RECT 55.415 4.305 55.43 4.52 ;
      RECT 55.405 4.305 55.415 4.514 ;
      RECT 55.395 4.312 55.405 4.511 ;
      RECT 55.39 4.35 55.395 4.5 ;
      RECT 55.385 4.412 55.39 4.478 ;
      RECT 56.655 4.287 56.84 4.51 ;
      RECT 56.655 4.302 56.845 4.506 ;
      RECT 56.645 3.575 56.73 4.505 ;
      RECT 56.645 4.302 56.85 4.499 ;
      RECT 56.64 4.31 56.85 4.498 ;
      RECT 56.845 4.03 57.165 4.35 ;
      RECT 56.64 4.202 56.81 4.293 ;
      RECT 56.635 4.202 56.81 4.275 ;
      RECT 56.625 4.01 56.76 4.25 ;
      RECT 56.62 4.01 56.76 4.195 ;
      RECT 56.58 3.59 56.75 4.095 ;
      RECT 56.565 3.59 56.75 3.965 ;
      RECT 56.56 3.59 56.75 3.918 ;
      RECT 56.555 3.59 56.75 3.898 ;
      RECT 56.55 3.59 56.75 3.873 ;
      RECT 56.52 3.59 56.78 3.85 ;
      RECT 56.53 3.587 56.74 3.85 ;
      RECT 56.655 3.582 56.74 4.51 ;
      RECT 56.54 3.575 56.73 3.85 ;
      RECT 56.535 3.58 56.73 3.85 ;
      RECT 55.365 3.792 55.55 4.005 ;
      RECT 55.365 3.8 55.56 3.998 ;
      RECT 55.345 3.8 55.56 3.995 ;
      RECT 55.34 3.8 55.56 3.98 ;
      RECT 55.27 3.715 55.53 3.975 ;
      RECT 55.27 3.86 55.565 3.888 ;
      RECT 54.925 4.315 55.185 4.575 ;
      RECT 54.95 4.26 55.145 4.575 ;
      RECT 54.945 4.009 55.125 4.303 ;
      RECT 54.945 4.015 55.135 4.303 ;
      RECT 54.925 4.017 55.135 4.248 ;
      RECT 54.92 4.027 55.135 4.115 ;
      RECT 54.95 4.007 55.125 4.575 ;
      RECT 55.036 4.005 55.125 4.575 ;
      RECT 54.895 3.225 54.93 3.595 ;
      RECT 54.685 3.335 54.69 3.595 ;
      RECT 54.93 3.232 54.945 3.595 ;
      RECT 54.82 3.225 54.895 3.673 ;
      RECT 54.81 3.225 54.82 3.758 ;
      RECT 54.785 3.225 54.81 3.793 ;
      RECT 54.745 3.225 54.785 3.861 ;
      RECT 54.735 3.232 54.745 3.913 ;
      RECT 54.705 3.335 54.735 3.954 ;
      RECT 54.7 3.335 54.705 3.993 ;
      RECT 54.69 3.335 54.7 4.013 ;
      RECT 54.685 3.63 54.69 4.05 ;
      RECT 54.68 3.647 54.685 4.07 ;
      RECT 54.665 3.71 54.68 4.11 ;
      RECT 54.66 3.753 54.665 4.145 ;
      RECT 54.655 3.761 54.66 4.158 ;
      RECT 54.645 3.775 54.655 4.18 ;
      RECT 54.62 3.81 54.645 4.245 ;
      RECT 54.61 3.845 54.62 4.308 ;
      RECT 54.59 3.875 54.61 4.369 ;
      RECT 54.575 3.911 54.59 4.436 ;
      RECT 54.565 3.939 54.575 4.475 ;
      RECT 54.555 3.961 54.565 4.495 ;
      RECT 54.55 3.971 54.555 4.506 ;
      RECT 54.545 3.98 54.55 4.509 ;
      RECT 54.535 3.998 54.545 4.513 ;
      RECT 54.525 4.016 54.535 4.514 ;
      RECT 54.5 4.055 54.525 4.511 ;
      RECT 54.48 4.097 54.5 4.508 ;
      RECT 54.465 4.135 54.48 4.507 ;
      RECT 54.43 4.17 54.465 4.504 ;
      RECT 54.425 4.192 54.43 4.502 ;
      RECT 54.36 4.232 54.425 4.499 ;
      RECT 54.355 4.272 54.36 4.495 ;
      RECT 54.34 4.282 54.355 4.486 ;
      RECT 54.33 4.402 54.34 4.471 ;
      RECT 54.81 4.815 54.82 5.075 ;
      RECT 54.81 4.818 54.83 5.074 ;
      RECT 54.8 4.808 54.81 5.073 ;
      RECT 54.79 4.823 54.87 5.069 ;
      RECT 54.775 4.802 54.79 5.067 ;
      RECT 54.75 4.827 54.875 5.063 ;
      RECT 54.735 4.787 54.75 5.058 ;
      RECT 54.735 4.829 54.885 5.057 ;
      RECT 54.735 4.837 54.9 5.05 ;
      RECT 54.675 4.774 54.735 5.04 ;
      RECT 54.665 4.761 54.675 5.022 ;
      RECT 54.64 4.751 54.665 5.012 ;
      RECT 54.635 4.741 54.64 5.004 ;
      RECT 54.57 4.837 54.9 4.986 ;
      RECT 54.485 4.837 54.9 4.948 ;
      RECT 54.375 4.665 54.635 4.925 ;
      RECT 54.75 4.795 54.775 5.063 ;
      RECT 54.79 4.805 54.8 5.069 ;
      RECT 54.375 4.813 54.815 4.925 ;
      RECT 54.56 10.06 54.85 10.29 ;
      RECT 54.62 9.32 54.79 10.29 ;
      RECT 54.52 9.345 54.89 9.715 ;
      RECT 54.56 9.32 54.85 9.715 ;
      RECT 53.59 4.57 53.62 4.87 ;
      RECT 53.365 4.555 53.37 4.83 ;
      RECT 53.165 4.555 53.32 4.815 ;
      RECT 54.465 3.27 54.495 3.53 ;
      RECT 54.455 3.27 54.465 3.638 ;
      RECT 54.435 3.27 54.455 3.648 ;
      RECT 54.42 3.27 54.435 3.66 ;
      RECT 54.365 3.27 54.42 3.71 ;
      RECT 54.35 3.27 54.365 3.758 ;
      RECT 54.32 3.27 54.35 3.793 ;
      RECT 54.265 3.27 54.32 3.855 ;
      RECT 54.245 3.27 54.265 3.923 ;
      RECT 54.24 3.27 54.245 3.953 ;
      RECT 54.235 3.27 54.24 3.965 ;
      RECT 54.23 3.387 54.235 3.983 ;
      RECT 54.21 3.405 54.23 4.008 ;
      RECT 54.19 3.432 54.21 4.058 ;
      RECT 54.185 3.452 54.19 4.089 ;
      RECT 54.18 3.46 54.185 4.106 ;
      RECT 54.165 3.486 54.18 4.135 ;
      RECT 54.15 3.528 54.165 4.17 ;
      RECT 54.145 3.557 54.15 4.193 ;
      RECT 54.14 3.572 54.145 4.206 ;
      RECT 54.135 3.595 54.14 4.217 ;
      RECT 54.125 3.615 54.135 4.235 ;
      RECT 54.115 3.645 54.125 4.258 ;
      RECT 54.11 3.667 54.115 4.278 ;
      RECT 54.105 3.682 54.11 4.293 ;
      RECT 54.09 3.712 54.105 4.32 ;
      RECT 54.085 3.742 54.09 4.346 ;
      RECT 54.08 3.76 54.085 4.358 ;
      RECT 54.07 3.79 54.08 4.377 ;
      RECT 54.06 3.815 54.07 4.402 ;
      RECT 54.055 3.835 54.06 4.421 ;
      RECT 54.05 3.852 54.055 4.434 ;
      RECT 54.04 3.878 54.05 4.453 ;
      RECT 54.03 3.916 54.04 4.48 ;
      RECT 54.025 3.942 54.03 4.5 ;
      RECT 54.02 3.952 54.025 4.51 ;
      RECT 54.015 3.965 54.02 4.525 ;
      RECT 54.01 3.98 54.015 4.535 ;
      RECT 54.005 4.002 54.01 4.55 ;
      RECT 54 4.02 54.005 4.561 ;
      RECT 53.995 4.03 54 4.572 ;
      RECT 53.99 4.038 53.995 4.584 ;
      RECT 53.985 4.046 53.99 4.595 ;
      RECT 53.98 4.072 53.985 4.608 ;
      RECT 53.97 4.1 53.98 4.621 ;
      RECT 53.965 4.13 53.97 4.63 ;
      RECT 53.96 4.145 53.965 4.637 ;
      RECT 53.945 4.17 53.96 4.644 ;
      RECT 53.94 4.192 53.945 4.65 ;
      RECT 53.935 4.217 53.94 4.653 ;
      RECT 53.926 4.245 53.935 4.657 ;
      RECT 53.92 4.262 53.926 4.662 ;
      RECT 53.915 4.28 53.92 4.666 ;
      RECT 53.91 4.292 53.915 4.669 ;
      RECT 53.905 4.313 53.91 4.673 ;
      RECT 53.9 4.331 53.905 4.676 ;
      RECT 53.895 4.345 53.9 4.679 ;
      RECT 53.89 4.362 53.895 4.682 ;
      RECT 53.885 4.375 53.89 4.685 ;
      RECT 53.86 4.412 53.885 4.693 ;
      RECT 53.855 4.457 53.86 4.702 ;
      RECT 53.85 4.485 53.855 4.705 ;
      RECT 53.84 4.505 53.85 4.709 ;
      RECT 53.835 4.525 53.84 4.714 ;
      RECT 53.83 4.54 53.835 4.717 ;
      RECT 53.81 4.55 53.83 4.724 ;
      RECT 53.745 4.557 53.81 4.75 ;
      RECT 53.71 4.56 53.745 4.778 ;
      RECT 53.695 4.563 53.71 4.793 ;
      RECT 53.685 4.564 53.695 4.808 ;
      RECT 53.675 4.565 53.685 4.825 ;
      RECT 53.67 4.565 53.675 4.84 ;
      RECT 53.665 4.565 53.67 4.848 ;
      RECT 53.65 4.566 53.665 4.863 ;
      RECT 53.62 4.568 53.65 4.87 ;
      RECT 53.51 4.575 53.59 4.87 ;
      RECT 53.465 4.58 53.51 4.87 ;
      RECT 53.455 4.581 53.465 4.86 ;
      RECT 53.445 4.582 53.455 4.853 ;
      RECT 53.425 4.584 53.445 4.848 ;
      RECT 53.415 4.555 53.425 4.843 ;
      RECT 53.37 4.555 53.415 4.835 ;
      RECT 53.34 4.555 53.365 4.825 ;
      RECT 53.32 4.555 53.34 4.818 ;
      RECT 53.6 3.355 53.86 3.615 ;
      RECT 53.48 3.37 53.49 3.535 ;
      RECT 53.465 3.37 53.47 3.53 ;
      RECT 50.83 3.21 51.015 3.5 ;
      RECT 52.645 3.335 52.66 3.49 ;
      RECT 50.795 3.21 50.82 3.47 ;
      RECT 53.21 3.26 53.215 3.402 ;
      RECT 53.125 3.255 53.15 3.395 ;
      RECT 53.525 3.372 53.6 3.565 ;
      RECT 53.51 3.37 53.525 3.548 ;
      RECT 53.49 3.37 53.51 3.54 ;
      RECT 53.47 3.37 53.48 3.533 ;
      RECT 53.425 3.365 53.465 3.523 ;
      RECT 53.385 3.34 53.425 3.508 ;
      RECT 53.37 3.315 53.385 3.498 ;
      RECT 53.365 3.309 53.37 3.496 ;
      RECT 53.33 3.301 53.365 3.479 ;
      RECT 53.325 3.294 53.33 3.467 ;
      RECT 53.305 3.289 53.325 3.455 ;
      RECT 53.295 3.283 53.305 3.44 ;
      RECT 53.275 3.278 53.295 3.425 ;
      RECT 53.265 3.273 53.275 3.418 ;
      RECT 53.26 3.271 53.265 3.413 ;
      RECT 53.255 3.27 53.26 3.41 ;
      RECT 53.215 3.265 53.255 3.406 ;
      RECT 53.195 3.259 53.21 3.401 ;
      RECT 53.16 3.256 53.195 3.398 ;
      RECT 53.15 3.255 53.16 3.396 ;
      RECT 53.09 3.255 53.125 3.393 ;
      RECT 53.045 3.255 53.09 3.393 ;
      RECT 52.995 3.255 53.045 3.396 ;
      RECT 52.98 3.257 52.995 3.398 ;
      RECT 52.965 3.26 52.98 3.399 ;
      RECT 52.955 3.265 52.965 3.4 ;
      RECT 52.925 3.27 52.955 3.405 ;
      RECT 52.915 3.276 52.925 3.413 ;
      RECT 52.905 3.278 52.915 3.417 ;
      RECT 52.895 3.282 52.905 3.421 ;
      RECT 52.87 3.288 52.895 3.429 ;
      RECT 52.86 3.293 52.87 3.437 ;
      RECT 52.845 3.297 52.86 3.441 ;
      RECT 52.81 3.303 52.845 3.449 ;
      RECT 52.79 3.308 52.81 3.459 ;
      RECT 52.76 3.315 52.79 3.468 ;
      RECT 52.715 3.324 52.76 3.482 ;
      RECT 52.71 3.329 52.715 3.493 ;
      RECT 52.69 3.332 52.71 3.494 ;
      RECT 52.66 3.335 52.69 3.492 ;
      RECT 52.625 3.335 52.645 3.488 ;
      RECT 52.555 3.335 52.625 3.479 ;
      RECT 52.54 3.332 52.555 3.471 ;
      RECT 52.5 3.325 52.54 3.466 ;
      RECT 52.475 3.315 52.5 3.459 ;
      RECT 52.47 3.309 52.475 3.456 ;
      RECT 52.43 3.303 52.47 3.453 ;
      RECT 52.415 3.296 52.43 3.448 ;
      RECT 52.395 3.292 52.415 3.443 ;
      RECT 52.38 3.287 52.395 3.439 ;
      RECT 52.365 3.282 52.38 3.437 ;
      RECT 52.35 3.278 52.365 3.436 ;
      RECT 52.335 3.276 52.35 3.432 ;
      RECT 52.325 3.274 52.335 3.427 ;
      RECT 52.31 3.271 52.325 3.423 ;
      RECT 52.3 3.269 52.31 3.418 ;
      RECT 52.28 3.266 52.3 3.414 ;
      RECT 52.235 3.265 52.28 3.412 ;
      RECT 52.175 3.267 52.235 3.413 ;
      RECT 52.155 3.269 52.175 3.415 ;
      RECT 52.125 3.272 52.155 3.416 ;
      RECT 52.075 3.277 52.125 3.418 ;
      RECT 52.07 3.28 52.075 3.42 ;
      RECT 52.06 3.282 52.07 3.423 ;
      RECT 52.055 3.284 52.06 3.426 ;
      RECT 52.005 3.287 52.055 3.433 ;
      RECT 51.985 3.291 52.005 3.445 ;
      RECT 51.975 3.294 51.985 3.451 ;
      RECT 51.965 3.295 51.975 3.454 ;
      RECT 51.926 3.298 51.965 3.456 ;
      RECT 51.84 3.305 51.926 3.459 ;
      RECT 51.766 3.315 51.84 3.463 ;
      RECT 51.68 3.326 51.766 3.468 ;
      RECT 51.665 3.333 51.68 3.47 ;
      RECT 51.61 3.337 51.665 3.471 ;
      RECT 51.596 3.34 51.61 3.473 ;
      RECT 51.51 3.34 51.596 3.475 ;
      RECT 51.47 3.337 51.51 3.478 ;
      RECT 51.446 3.333 51.47 3.48 ;
      RECT 51.36 3.323 51.446 3.483 ;
      RECT 51.33 3.312 51.36 3.484 ;
      RECT 51.311 3.308 51.33 3.483 ;
      RECT 51.225 3.301 51.311 3.48 ;
      RECT 51.165 3.29 51.225 3.477 ;
      RECT 51.145 3.282 51.165 3.475 ;
      RECT 51.11 3.277 51.145 3.474 ;
      RECT 51.085 3.272 51.11 3.473 ;
      RECT 51.055 3.267 51.085 3.472 ;
      RECT 51.03 3.21 51.055 3.471 ;
      RECT 51.015 3.21 51.03 3.495 ;
      RECT 50.82 3.21 50.83 3.495 ;
      RECT 52.595 4.23 52.6 4.37 ;
      RECT 52.255 4.23 52.29 4.368 ;
      RECT 51.83 4.215 51.845 4.36 ;
      RECT 53.66 3.995 53.75 4.255 ;
      RECT 53.49 3.86 53.59 4.255 ;
      RECT 50.525 3.835 50.605 4.045 ;
      RECT 53.615 3.972 53.66 4.255 ;
      RECT 53.605 3.942 53.615 4.255 ;
      RECT 53.59 3.865 53.605 4.255 ;
      RECT 53.405 3.86 53.49 4.22 ;
      RECT 53.4 3.862 53.405 4.215 ;
      RECT 53.395 3.867 53.4 4.215 ;
      RECT 53.36 3.967 53.395 4.215 ;
      RECT 53.35 3.995 53.36 4.215 ;
      RECT 53.34 4.01 53.35 4.215 ;
      RECT 53.33 4.022 53.34 4.215 ;
      RECT 53.325 4.032 53.33 4.215 ;
      RECT 53.31 4.042 53.325 4.217 ;
      RECT 53.305 4.057 53.31 4.219 ;
      RECT 53.29 4.07 53.305 4.221 ;
      RECT 53.285 4.085 53.29 4.224 ;
      RECT 53.265 4.095 53.285 4.228 ;
      RECT 53.25 4.105 53.265 4.231 ;
      RECT 53.215 4.112 53.25 4.236 ;
      RECT 53.171 4.119 53.215 4.244 ;
      RECT 53.085 4.131 53.171 4.257 ;
      RECT 53.06 4.142 53.085 4.268 ;
      RECT 53.03 4.147 53.06 4.273 ;
      RECT 52.995 4.152 53.03 4.281 ;
      RECT 52.965 4.157 52.995 4.288 ;
      RECT 52.94 4.162 52.965 4.293 ;
      RECT 52.875 4.169 52.94 4.302 ;
      RECT 52.805 4.182 52.875 4.318 ;
      RECT 52.775 4.192 52.805 4.33 ;
      RECT 52.75 4.197 52.775 4.337 ;
      RECT 52.695 4.204 52.75 4.345 ;
      RECT 52.69 4.211 52.695 4.35 ;
      RECT 52.685 4.213 52.69 4.351 ;
      RECT 52.67 4.215 52.685 4.353 ;
      RECT 52.665 4.215 52.67 4.356 ;
      RECT 52.6 4.222 52.665 4.363 ;
      RECT 52.565 4.232 52.595 4.373 ;
      RECT 52.548 4.235 52.565 4.375 ;
      RECT 52.462 4.234 52.548 4.374 ;
      RECT 52.376 4.232 52.462 4.371 ;
      RECT 52.29 4.231 52.376 4.369 ;
      RECT 52.189 4.229 52.255 4.368 ;
      RECT 52.103 4.226 52.189 4.366 ;
      RECT 52.017 4.222 52.103 4.364 ;
      RECT 51.931 4.219 52.017 4.363 ;
      RECT 51.845 4.216 51.931 4.361 ;
      RECT 51.745 4.215 51.83 4.358 ;
      RECT 51.695 4.213 51.745 4.356 ;
      RECT 51.675 4.21 51.695 4.354 ;
      RECT 51.655 4.208 51.675 4.351 ;
      RECT 51.63 4.204 51.655 4.348 ;
      RECT 51.585 4.198 51.63 4.343 ;
      RECT 51.545 4.192 51.585 4.335 ;
      RECT 51.52 4.187 51.545 4.328 ;
      RECT 51.465 4.18 51.52 4.32 ;
      RECT 51.441 4.173 51.465 4.313 ;
      RECT 51.355 4.164 51.441 4.303 ;
      RECT 51.325 4.156 51.355 4.293 ;
      RECT 51.295 4.152 51.325 4.288 ;
      RECT 51.29 4.149 51.295 4.285 ;
      RECT 51.285 4.148 51.29 4.285 ;
      RECT 51.21 4.141 51.285 4.278 ;
      RECT 51.171 4.132 51.21 4.267 ;
      RECT 51.085 4.122 51.171 4.255 ;
      RECT 51.045 4.112 51.085 4.243 ;
      RECT 51.006 4.107 51.045 4.236 ;
      RECT 50.92 4.097 51.006 4.225 ;
      RECT 50.88 4.085 50.92 4.214 ;
      RECT 50.845 4.07 50.88 4.207 ;
      RECT 50.835 4.06 50.845 4.204 ;
      RECT 50.815 4.045 50.835 4.202 ;
      RECT 50.785 4.015 50.815 4.198 ;
      RECT 50.775 3.995 50.785 4.193 ;
      RECT 50.77 3.987 50.775 4.19 ;
      RECT 50.765 3.98 50.77 4.188 ;
      RECT 50.75 3.967 50.765 4.181 ;
      RECT 50.745 3.957 50.75 4.173 ;
      RECT 50.74 3.95 50.745 4.168 ;
      RECT 50.735 3.945 50.74 4.164 ;
      RECT 50.72 3.932 50.735 4.156 ;
      RECT 50.715 3.842 50.72 4.145 ;
      RECT 50.71 3.837 50.715 4.138 ;
      RECT 50.635 3.835 50.71 4.098 ;
      RECT 50.605 3.835 50.635 4.053 ;
      RECT 50.51 3.84 50.525 4.04 ;
      RECT 52.995 3.545 53.255 3.805 ;
      RECT 52.98 3.533 53.16 3.77 ;
      RECT 52.975 3.534 53.16 3.768 ;
      RECT 52.96 3.538 53.17 3.758 ;
      RECT 52.955 3.543 53.175 3.728 ;
      RECT 52.96 3.54 53.175 3.758 ;
      RECT 52.975 3.535 53.17 3.768 ;
      RECT 52.995 3.532 53.16 3.805 ;
      RECT 52.995 3.531 53.15 3.805 ;
      RECT 53.02 3.53 53.15 3.805 ;
      RECT 52.58 3.775 52.84 4.035 ;
      RECT 52.455 3.82 52.84 4.03 ;
      RECT 52.445 3.825 52.84 4.025 ;
      RECT 52.46 4.765 52.475 5.075 ;
      RECT 51.055 4.535 51.065 4.665 ;
      RECT 50.835 4.53 50.94 4.665 ;
      RECT 50.75 4.535 50.8 4.665 ;
      RECT 49.3 3.27 49.305 4.375 ;
      RECT 52.555 4.857 52.56 4.993 ;
      RECT 52.55 4.852 52.555 5.053 ;
      RECT 52.545 4.85 52.55 5.066 ;
      RECT 52.53 4.847 52.545 5.068 ;
      RECT 52.525 4.842 52.53 5.07 ;
      RECT 52.52 4.838 52.525 5.073 ;
      RECT 52.505 4.833 52.52 5.075 ;
      RECT 52.475 4.825 52.505 5.075 ;
      RECT 52.436 4.765 52.46 5.075 ;
      RECT 52.35 4.765 52.436 5.072 ;
      RECT 52.32 4.765 52.35 5.065 ;
      RECT 52.295 4.765 52.32 5.058 ;
      RECT 52.27 4.765 52.295 5.05 ;
      RECT 52.255 4.765 52.27 5.043 ;
      RECT 52.23 4.765 52.255 5.035 ;
      RECT 52.215 4.765 52.23 5.028 ;
      RECT 52.175 4.775 52.215 5.017 ;
      RECT 52.165 4.77 52.175 5.007 ;
      RECT 52.161 4.769 52.165 5.004 ;
      RECT 52.075 4.761 52.161 4.987 ;
      RECT 52.042 4.75 52.075 4.964 ;
      RECT 51.956 4.739 52.042 4.942 ;
      RECT 51.87 4.723 51.956 4.911 ;
      RECT 51.8 4.708 51.87 4.883 ;
      RECT 51.79 4.701 51.8 4.87 ;
      RECT 51.76 4.698 51.79 4.86 ;
      RECT 51.735 4.694 51.76 4.853 ;
      RECT 51.72 4.691 51.735 4.848 ;
      RECT 51.715 4.69 51.72 4.843 ;
      RECT 51.685 4.685 51.715 4.836 ;
      RECT 51.68 4.68 51.685 4.831 ;
      RECT 51.665 4.677 51.68 4.826 ;
      RECT 51.66 4.672 51.665 4.821 ;
      RECT 51.64 4.667 51.66 4.818 ;
      RECT 51.625 4.662 51.64 4.81 ;
      RECT 51.61 4.656 51.625 4.805 ;
      RECT 51.58 4.647 51.61 4.798 ;
      RECT 51.575 4.64 51.58 4.79 ;
      RECT 51.57 4.638 51.575 4.788 ;
      RECT 51.565 4.637 51.57 4.785 ;
      RECT 51.525 4.63 51.565 4.778 ;
      RECT 51.511 4.62 51.525 4.768 ;
      RECT 51.46 4.609 51.511 4.756 ;
      RECT 51.435 4.595 51.46 4.742 ;
      RECT 51.41 4.584 51.435 4.734 ;
      RECT 51.39 4.573 51.41 4.728 ;
      RECT 51.38 4.567 51.39 4.723 ;
      RECT 51.375 4.565 51.38 4.719 ;
      RECT 51.355 4.56 51.375 4.714 ;
      RECT 51.325 4.55 51.355 4.704 ;
      RECT 51.32 4.542 51.325 4.697 ;
      RECT 51.305 4.54 51.32 4.693 ;
      RECT 51.285 4.54 51.305 4.688 ;
      RECT 51.28 4.539 51.285 4.686 ;
      RECT 51.275 4.539 51.28 4.683 ;
      RECT 51.235 4.538 51.275 4.678 ;
      RECT 51.21 4.537 51.235 4.673 ;
      RECT 51.15 4.536 51.21 4.67 ;
      RECT 51.065 4.535 51.15 4.668 ;
      RECT 51.026 4.534 51.055 4.665 ;
      RECT 50.94 4.532 51.026 4.665 ;
      RECT 50.8 4.532 50.835 4.665 ;
      RECT 50.71 4.536 50.75 4.668 ;
      RECT 50.695 4.539 50.71 4.675 ;
      RECT 50.685 4.54 50.695 4.682 ;
      RECT 50.66 4.543 50.685 4.687 ;
      RECT 50.655 4.545 50.66 4.69 ;
      RECT 50.605 4.547 50.655 4.691 ;
      RECT 50.566 4.551 50.605 4.693 ;
      RECT 50.48 4.553 50.566 4.696 ;
      RECT 50.462 4.555 50.48 4.698 ;
      RECT 50.376 4.558 50.462 4.7 ;
      RECT 50.29 4.562 50.376 4.703 ;
      RECT 50.253 4.566 50.29 4.706 ;
      RECT 50.167 4.569 50.253 4.709 ;
      RECT 50.081 4.573 50.167 4.712 ;
      RECT 49.995 4.578 50.081 4.716 ;
      RECT 49.975 4.58 49.995 4.719 ;
      RECT 49.955 4.579 49.975 4.72 ;
      RECT 49.906 4.576 49.955 4.721 ;
      RECT 49.82 4.571 49.906 4.724 ;
      RECT 49.77 4.566 49.82 4.726 ;
      RECT 49.746 4.564 49.77 4.727 ;
      RECT 49.66 4.559 49.746 4.729 ;
      RECT 49.635 4.555 49.66 4.728 ;
      RECT 49.625 4.552 49.635 4.726 ;
      RECT 49.615 4.545 49.625 4.723 ;
      RECT 49.61 4.525 49.615 4.718 ;
      RECT 49.6 4.495 49.61 4.713 ;
      RECT 49.585 4.365 49.6 4.704 ;
      RECT 49.58 4.357 49.585 4.697 ;
      RECT 49.56 4.35 49.58 4.689 ;
      RECT 49.555 4.332 49.56 4.681 ;
      RECT 49.545 4.312 49.555 4.676 ;
      RECT 49.54 4.285 49.545 4.672 ;
      RECT 49.535 4.262 49.54 4.669 ;
      RECT 49.515 4.22 49.535 4.661 ;
      RECT 49.48 4.135 49.515 4.645 ;
      RECT 49.475 4.067 49.48 4.633 ;
      RECT 49.46 4.037 49.475 4.627 ;
      RECT 49.455 3.282 49.46 3.528 ;
      RECT 49.445 4.007 49.46 4.618 ;
      RECT 49.45 3.277 49.455 3.56 ;
      RECT 49.445 3.272 49.45 3.603 ;
      RECT 49.44 3.27 49.445 3.638 ;
      RECT 49.425 3.97 49.445 4.608 ;
      RECT 49.435 3.27 49.44 3.675 ;
      RECT 49.42 3.27 49.435 3.773 ;
      RECT 49.42 3.943 49.425 4.601 ;
      RECT 49.415 3.27 49.42 3.848 ;
      RECT 49.415 3.931 49.42 4.598 ;
      RECT 49.41 3.27 49.415 3.88 ;
      RECT 49.41 3.91 49.415 4.595 ;
      RECT 49.405 3.27 49.41 4.592 ;
      RECT 49.37 3.27 49.405 4.578 ;
      RECT 49.355 3.27 49.37 4.56 ;
      RECT 49.335 3.27 49.355 4.55 ;
      RECT 49.31 3.27 49.335 4.533 ;
      RECT 49.305 3.27 49.31 4.483 ;
      RECT 49.295 3.27 49.3 4.313 ;
      RECT 49.29 3.27 49.295 4.22 ;
      RECT 49.285 3.27 49.29 4.133 ;
      RECT 49.28 3.27 49.285 4.065 ;
      RECT 49.275 3.27 49.28 4.008 ;
      RECT 49.265 3.27 49.275 3.903 ;
      RECT 49.26 3.27 49.265 3.775 ;
      RECT 49.255 3.27 49.26 3.693 ;
      RECT 49.25 3.272 49.255 3.61 ;
      RECT 49.245 3.277 49.25 3.543 ;
      RECT 49.24 3.282 49.245 3.47 ;
      RECT 52.055 3.6 52.315 3.86 ;
      RECT 52.075 3.567 52.285 3.86 ;
      RECT 52.075 3.565 52.275 3.86 ;
      RECT 52.085 3.552 52.275 3.86 ;
      RECT 52.085 3.55 52.2 3.86 ;
      RECT 51.56 3.675 51.735 3.955 ;
      RECT 51.555 3.675 51.735 3.953 ;
      RECT 51.555 3.675 51.75 3.95 ;
      RECT 51.545 3.675 51.75 3.948 ;
      RECT 51.49 3.675 51.75 3.935 ;
      RECT 51.49 3.75 51.755 3.913 ;
      RECT 51.02 4.873 51.025 5.08 ;
      RECT 50.97 4.867 51.02 5.079 ;
      RECT 50.937 4.881 51.03 5.078 ;
      RECT 50.851 4.881 51.03 5.077 ;
      RECT 50.765 4.881 51.03 5.076 ;
      RECT 50.765 4.98 51.035 5.073 ;
      RECT 50.76 4.98 51.035 5.068 ;
      RECT 50.755 4.98 51.035 5.05 ;
      RECT 50.75 4.98 51.035 5.033 ;
      RECT 50.71 4.765 50.97 5.025 ;
      RECT 50.17 3.915 50.256 4.329 ;
      RECT 50.17 3.915 50.295 4.326 ;
      RECT 50.17 3.915 50.315 4.316 ;
      RECT 50.125 3.915 50.315 4.313 ;
      RECT 50.125 4.067 50.325 4.303 ;
      RECT 50.125 4.088 50.33 4.297 ;
      RECT 50.125 4.106 50.335 4.293 ;
      RECT 50.125 4.126 50.345 4.288 ;
      RECT 50.1 4.126 50.345 4.285 ;
      RECT 50.09 4.126 50.345 4.263 ;
      RECT 50.09 4.142 50.35 4.233 ;
      RECT 50.055 3.915 50.315 4.22 ;
      RECT 50.055 4.154 50.355 4.175 ;
      RECT 47.715 10.06 48.01 10.29 ;
      RECT 47.775 8.58 47.945 10.29 ;
      RECT 47.765 8.95 48.12 9.305 ;
      RECT 47.715 8.58 48.005 8.81 ;
      RECT 46.725 10.06 47.02 10.29 ;
      RECT 46.785 8.58 46.955 10.29 ;
      RECT 46.725 8.58 47.015 8.81 ;
      RECT 46.725 8.615 47.575 8.775 ;
      RECT 47.41 8.21 47.575 8.775 ;
      RECT 46.725 8.61 47.12 8.775 ;
      RECT 47.345 8.21 47.635 8.44 ;
      RECT 47.345 8.24 47.805 8.41 ;
      RECT 47.31 4.025 47.63 4.26 ;
      RECT 47.31 4.055 47.8 4.225 ;
      RECT 47.31 3.69 47.5 4.26 ;
      RECT 46.725 3.655 47.015 3.885 ;
      RECT 46.725 3.69 47.5 3.86 ;
      RECT 46.785 2.175 46.955 3.885 ;
      RECT 46.725 2.175 47.02 2.405 ;
      RECT 46.355 4.025 46.645 4.255 ;
      RECT 46.355 4.055 46.815 4.225 ;
      RECT 46.42 2.95 46.585 4.255 ;
      RECT 44.935 2.915 45.225 3.145 ;
      RECT 44.935 2.95 46.585 3.12 ;
      RECT 44.995 2.175 45.165 3.145 ;
      RECT 44.935 2.175 45.225 2.405 ;
      RECT 44.935 10.06 45.225 10.29 ;
      RECT 44.995 9.32 45.165 10.29 ;
      RECT 44.995 9.41 46.585 9.58 ;
      RECT 46.415 8.21 46.585 9.58 ;
      RECT 44.935 9.32 45.225 9.55 ;
      RECT 46.355 8.21 46.645 8.44 ;
      RECT 46.355 8.24 46.815 8.41 ;
      RECT 42.985 4 43.325 4.35 ;
      RECT 43.075 3.32 43.245 4.35 ;
      RECT 45.365 3.26 45.715 3.61 ;
      RECT 43.075 3.32 45.715 3.49 ;
      RECT 45.195 3.315 45.715 3.49 ;
      RECT 45.39 8.945 45.715 9.27 ;
      RECT 39.93 8.905 40.28 9.255 ;
      RECT 45.365 8.95 45.715 9.18 ;
      RECT 39.73 8.95 40.28 9.18 ;
      RECT 45.195 8.975 45.715 9.15 ;
      RECT 39.56 8.98 40.28 9.15 ;
      RECT 39.61 8.975 45.715 9.145 ;
      RECT 44.59 3.66 44.91 3.98 ;
      RECT 44.565 3.655 44.855 3.885 ;
      RECT 44.56 3.685 44.91 3.86 ;
      RECT 44.39 3.685 44.91 3.855 ;
      RECT 44.59 8.545 44.91 8.835 ;
      RECT 44.565 8.58 44.91 8.81 ;
      RECT 44.39 8.61 44.91 8.78 ;
      RECT 40.28 4.28 40.43 4.555 ;
      RECT 40.82 3.36 40.825 3.58 ;
      RECT 41.97 3.56 41.985 3.758 ;
      RECT 41.935 3.552 41.97 3.765 ;
      RECT 41.905 3.545 41.935 3.765 ;
      RECT 41.85 3.51 41.905 3.765 ;
      RECT 41.785 3.447 41.85 3.765 ;
      RECT 41.78 3.412 41.785 3.763 ;
      RECT 41.775 3.407 41.78 3.755 ;
      RECT 41.77 3.402 41.775 3.741 ;
      RECT 41.765 3.399 41.77 3.734 ;
      RECT 41.72 3.389 41.765 3.685 ;
      RECT 41.7 3.376 41.72 3.62 ;
      RECT 41.695 3.371 41.7 3.593 ;
      RECT 41.69 3.37 41.695 3.586 ;
      RECT 41.685 3.369 41.69 3.579 ;
      RECT 41.6 3.354 41.685 3.525 ;
      RECT 41.57 3.335 41.6 3.475 ;
      RECT 41.49 3.318 41.57 3.46 ;
      RECT 41.455 3.305 41.49 3.445 ;
      RECT 41.447 3.305 41.455 3.44 ;
      RECT 41.361 3.306 41.447 3.44 ;
      RECT 41.275 3.308 41.361 3.44 ;
      RECT 41.25 3.309 41.275 3.444 ;
      RECT 41.175 3.315 41.25 3.459 ;
      RECT 41.092 3.327 41.175 3.483 ;
      RECT 41.006 3.34 41.092 3.509 ;
      RECT 40.92 3.353 41.006 3.535 ;
      RECT 40.885 3.362 40.92 3.554 ;
      RECT 40.835 3.362 40.885 3.567 ;
      RECT 40.825 3.36 40.835 3.578 ;
      RECT 40.81 3.357 40.82 3.58 ;
      RECT 40.795 3.349 40.81 3.588 ;
      RECT 40.78 3.341 40.795 3.608 ;
      RECT 40.775 3.336 40.78 3.665 ;
      RECT 40.76 3.331 40.775 3.738 ;
      RECT 40.755 3.326 40.76 3.78 ;
      RECT 40.75 3.324 40.755 3.808 ;
      RECT 40.745 3.322 40.75 3.83 ;
      RECT 40.735 3.318 40.745 3.873 ;
      RECT 40.73 3.315 40.735 3.898 ;
      RECT 40.725 3.313 40.73 3.918 ;
      RECT 40.72 3.311 40.725 3.942 ;
      RECT 40.715 3.307 40.72 3.965 ;
      RECT 40.71 3.303 40.715 3.988 ;
      RECT 40.675 3.293 40.71 4.095 ;
      RECT 40.67 3.283 40.675 4.193 ;
      RECT 40.665 3.281 40.67 4.22 ;
      RECT 40.66 3.28 40.665 4.24 ;
      RECT 40.655 3.272 40.66 4.26 ;
      RECT 40.65 3.267 40.655 4.295 ;
      RECT 40.645 3.265 40.65 4.313 ;
      RECT 40.64 3.265 40.645 4.338 ;
      RECT 40.635 3.265 40.64 4.36 ;
      RECT 40.6 3.265 40.635 4.403 ;
      RECT 40.575 3.265 40.6 4.432 ;
      RECT 40.565 3.265 40.575 3.618 ;
      RECT 40.568 3.675 40.575 4.442 ;
      RECT 40.565 3.732 40.568 4.445 ;
      RECT 40.56 3.265 40.565 3.59 ;
      RECT 40.56 3.782 40.565 4.448 ;
      RECT 40.55 3.265 40.56 3.58 ;
      RECT 40.555 3.835 40.56 4.451 ;
      RECT 40.55 3.92 40.555 4.455 ;
      RECT 40.54 3.265 40.55 3.568 ;
      RECT 40.545 3.967 40.55 4.459 ;
      RECT 40.54 4.042 40.545 4.463 ;
      RECT 40.505 3.265 40.54 3.543 ;
      RECT 40.53 4.125 40.54 4.468 ;
      RECT 40.52 4.192 40.53 4.475 ;
      RECT 40.515 4.22 40.52 4.48 ;
      RECT 40.505 4.233 40.515 4.486 ;
      RECT 40.46 3.265 40.505 3.5 ;
      RECT 40.5 4.238 40.505 4.493 ;
      RECT 40.46 4.255 40.5 4.555 ;
      RECT 40.455 3.267 40.46 3.473 ;
      RECT 40.43 4.275 40.46 4.555 ;
      RECT 40.45 3.272 40.455 3.445 ;
      RECT 40.24 4.284 40.28 4.555 ;
      RECT 40.215 4.292 40.24 4.525 ;
      RECT 40.17 4.3 40.215 4.525 ;
      RECT 40.155 4.305 40.17 4.52 ;
      RECT 40.145 4.305 40.155 4.514 ;
      RECT 40.135 4.312 40.145 4.511 ;
      RECT 40.13 4.35 40.135 4.5 ;
      RECT 40.125 4.412 40.13 4.478 ;
      RECT 41.395 4.287 41.58 4.51 ;
      RECT 41.395 4.302 41.585 4.506 ;
      RECT 41.385 3.575 41.47 4.505 ;
      RECT 41.385 4.302 41.59 4.499 ;
      RECT 41.38 4.31 41.59 4.498 ;
      RECT 41.585 4.03 41.905 4.35 ;
      RECT 41.38 4.202 41.55 4.293 ;
      RECT 41.375 4.202 41.55 4.275 ;
      RECT 41.365 4.01 41.5 4.25 ;
      RECT 41.36 4.01 41.5 4.195 ;
      RECT 41.32 3.59 41.49 4.095 ;
      RECT 41.305 3.59 41.49 3.965 ;
      RECT 41.3 3.59 41.49 3.918 ;
      RECT 41.295 3.59 41.49 3.898 ;
      RECT 41.29 3.59 41.49 3.873 ;
      RECT 41.26 3.59 41.52 3.85 ;
      RECT 41.27 3.587 41.48 3.85 ;
      RECT 41.395 3.582 41.48 4.51 ;
      RECT 41.28 3.575 41.47 3.85 ;
      RECT 41.275 3.58 41.47 3.85 ;
      RECT 40.105 3.792 40.29 4.005 ;
      RECT 40.105 3.8 40.3 3.998 ;
      RECT 40.085 3.8 40.3 3.995 ;
      RECT 40.08 3.8 40.3 3.98 ;
      RECT 40.01 3.715 40.27 3.975 ;
      RECT 40.01 3.86 40.305 3.888 ;
      RECT 39.665 4.315 39.925 4.575 ;
      RECT 39.69 4.26 39.885 4.575 ;
      RECT 39.685 4.009 39.865 4.303 ;
      RECT 39.685 4.015 39.875 4.303 ;
      RECT 39.665 4.017 39.875 4.248 ;
      RECT 39.66 4.027 39.875 4.115 ;
      RECT 39.69 4.007 39.865 4.575 ;
      RECT 39.776 4.005 39.865 4.575 ;
      RECT 39.635 3.225 39.67 3.595 ;
      RECT 39.425 3.335 39.43 3.595 ;
      RECT 39.67 3.232 39.685 3.595 ;
      RECT 39.56 3.225 39.635 3.673 ;
      RECT 39.55 3.225 39.56 3.758 ;
      RECT 39.525 3.225 39.55 3.793 ;
      RECT 39.485 3.225 39.525 3.861 ;
      RECT 39.475 3.232 39.485 3.913 ;
      RECT 39.445 3.335 39.475 3.954 ;
      RECT 39.44 3.335 39.445 3.993 ;
      RECT 39.43 3.335 39.44 4.013 ;
      RECT 39.425 3.63 39.43 4.05 ;
      RECT 39.42 3.647 39.425 4.07 ;
      RECT 39.405 3.71 39.42 4.11 ;
      RECT 39.4 3.753 39.405 4.145 ;
      RECT 39.395 3.761 39.4 4.158 ;
      RECT 39.385 3.775 39.395 4.18 ;
      RECT 39.36 3.81 39.385 4.245 ;
      RECT 39.35 3.845 39.36 4.308 ;
      RECT 39.33 3.875 39.35 4.369 ;
      RECT 39.315 3.911 39.33 4.436 ;
      RECT 39.305 3.939 39.315 4.475 ;
      RECT 39.295 3.961 39.305 4.495 ;
      RECT 39.29 3.971 39.295 4.506 ;
      RECT 39.285 3.98 39.29 4.509 ;
      RECT 39.275 3.998 39.285 4.513 ;
      RECT 39.265 4.016 39.275 4.514 ;
      RECT 39.24 4.055 39.265 4.511 ;
      RECT 39.22 4.097 39.24 4.508 ;
      RECT 39.205 4.135 39.22 4.507 ;
      RECT 39.17 4.17 39.205 4.504 ;
      RECT 39.165 4.192 39.17 4.502 ;
      RECT 39.1 4.232 39.165 4.499 ;
      RECT 39.095 4.272 39.1 4.495 ;
      RECT 39.08 4.282 39.095 4.486 ;
      RECT 39.07 4.402 39.08 4.471 ;
      RECT 39.55 4.815 39.56 5.075 ;
      RECT 39.55 4.818 39.57 5.074 ;
      RECT 39.54 4.808 39.55 5.073 ;
      RECT 39.53 4.823 39.61 5.069 ;
      RECT 39.515 4.802 39.53 5.067 ;
      RECT 39.49 4.827 39.615 5.063 ;
      RECT 39.475 4.787 39.49 5.058 ;
      RECT 39.475 4.829 39.625 5.057 ;
      RECT 39.475 4.837 39.64 5.05 ;
      RECT 39.415 4.774 39.475 5.04 ;
      RECT 39.405 4.761 39.415 5.022 ;
      RECT 39.38 4.751 39.405 5.012 ;
      RECT 39.375 4.741 39.38 5.004 ;
      RECT 39.31 4.837 39.64 4.986 ;
      RECT 39.225 4.837 39.64 4.948 ;
      RECT 39.115 4.665 39.375 4.925 ;
      RECT 39.49 4.795 39.515 5.063 ;
      RECT 39.53 4.805 39.54 5.069 ;
      RECT 39.115 4.813 39.555 4.925 ;
      RECT 39.3 10.06 39.59 10.29 ;
      RECT 39.36 9.32 39.53 10.29 ;
      RECT 39.26 9.345 39.63 9.715 ;
      RECT 39.3 9.32 39.59 9.715 ;
      RECT 38.33 4.57 38.36 4.87 ;
      RECT 38.105 4.555 38.11 4.83 ;
      RECT 37.905 4.555 38.06 4.815 ;
      RECT 39.205 3.27 39.235 3.53 ;
      RECT 39.195 3.27 39.205 3.638 ;
      RECT 39.175 3.27 39.195 3.648 ;
      RECT 39.16 3.27 39.175 3.66 ;
      RECT 39.105 3.27 39.16 3.71 ;
      RECT 39.09 3.27 39.105 3.758 ;
      RECT 39.06 3.27 39.09 3.793 ;
      RECT 39.005 3.27 39.06 3.855 ;
      RECT 38.985 3.27 39.005 3.923 ;
      RECT 38.98 3.27 38.985 3.953 ;
      RECT 38.975 3.27 38.98 3.965 ;
      RECT 38.97 3.387 38.975 3.983 ;
      RECT 38.95 3.405 38.97 4.008 ;
      RECT 38.93 3.432 38.95 4.058 ;
      RECT 38.925 3.452 38.93 4.089 ;
      RECT 38.92 3.46 38.925 4.106 ;
      RECT 38.905 3.486 38.92 4.135 ;
      RECT 38.89 3.528 38.905 4.17 ;
      RECT 38.885 3.557 38.89 4.193 ;
      RECT 38.88 3.572 38.885 4.206 ;
      RECT 38.875 3.595 38.88 4.217 ;
      RECT 38.865 3.615 38.875 4.235 ;
      RECT 38.855 3.645 38.865 4.258 ;
      RECT 38.85 3.667 38.855 4.278 ;
      RECT 38.845 3.682 38.85 4.293 ;
      RECT 38.83 3.712 38.845 4.32 ;
      RECT 38.825 3.742 38.83 4.346 ;
      RECT 38.82 3.76 38.825 4.358 ;
      RECT 38.81 3.79 38.82 4.377 ;
      RECT 38.8 3.815 38.81 4.402 ;
      RECT 38.795 3.835 38.8 4.421 ;
      RECT 38.79 3.852 38.795 4.434 ;
      RECT 38.78 3.878 38.79 4.453 ;
      RECT 38.77 3.916 38.78 4.48 ;
      RECT 38.765 3.942 38.77 4.5 ;
      RECT 38.76 3.952 38.765 4.51 ;
      RECT 38.755 3.965 38.76 4.525 ;
      RECT 38.75 3.98 38.755 4.535 ;
      RECT 38.745 4.002 38.75 4.55 ;
      RECT 38.74 4.02 38.745 4.561 ;
      RECT 38.735 4.03 38.74 4.572 ;
      RECT 38.73 4.038 38.735 4.584 ;
      RECT 38.725 4.046 38.73 4.595 ;
      RECT 38.72 4.072 38.725 4.608 ;
      RECT 38.71 4.1 38.72 4.621 ;
      RECT 38.705 4.13 38.71 4.63 ;
      RECT 38.7 4.145 38.705 4.637 ;
      RECT 38.685 4.17 38.7 4.644 ;
      RECT 38.68 4.192 38.685 4.65 ;
      RECT 38.675 4.217 38.68 4.653 ;
      RECT 38.666 4.245 38.675 4.657 ;
      RECT 38.66 4.262 38.666 4.662 ;
      RECT 38.655 4.28 38.66 4.666 ;
      RECT 38.65 4.292 38.655 4.669 ;
      RECT 38.645 4.313 38.65 4.673 ;
      RECT 38.64 4.331 38.645 4.676 ;
      RECT 38.635 4.345 38.64 4.679 ;
      RECT 38.63 4.362 38.635 4.682 ;
      RECT 38.625 4.375 38.63 4.685 ;
      RECT 38.6 4.412 38.625 4.693 ;
      RECT 38.595 4.457 38.6 4.702 ;
      RECT 38.59 4.485 38.595 4.705 ;
      RECT 38.58 4.505 38.59 4.709 ;
      RECT 38.575 4.525 38.58 4.714 ;
      RECT 38.57 4.54 38.575 4.717 ;
      RECT 38.55 4.55 38.57 4.724 ;
      RECT 38.485 4.557 38.55 4.75 ;
      RECT 38.45 4.56 38.485 4.778 ;
      RECT 38.435 4.563 38.45 4.793 ;
      RECT 38.425 4.564 38.435 4.808 ;
      RECT 38.415 4.565 38.425 4.825 ;
      RECT 38.41 4.565 38.415 4.84 ;
      RECT 38.405 4.565 38.41 4.848 ;
      RECT 38.39 4.566 38.405 4.863 ;
      RECT 38.36 4.568 38.39 4.87 ;
      RECT 38.25 4.575 38.33 4.87 ;
      RECT 38.205 4.58 38.25 4.87 ;
      RECT 38.195 4.581 38.205 4.86 ;
      RECT 38.185 4.582 38.195 4.853 ;
      RECT 38.165 4.584 38.185 4.848 ;
      RECT 38.155 4.555 38.165 4.843 ;
      RECT 38.11 4.555 38.155 4.835 ;
      RECT 38.08 4.555 38.105 4.825 ;
      RECT 38.06 4.555 38.08 4.818 ;
      RECT 38.34 3.355 38.6 3.615 ;
      RECT 38.22 3.37 38.23 3.535 ;
      RECT 38.205 3.37 38.21 3.53 ;
      RECT 35.57 3.21 35.755 3.5 ;
      RECT 37.385 3.335 37.4 3.49 ;
      RECT 35.535 3.21 35.56 3.47 ;
      RECT 37.95 3.26 37.955 3.402 ;
      RECT 37.865 3.255 37.89 3.395 ;
      RECT 38.265 3.372 38.34 3.565 ;
      RECT 38.25 3.37 38.265 3.548 ;
      RECT 38.23 3.37 38.25 3.54 ;
      RECT 38.21 3.37 38.22 3.533 ;
      RECT 38.165 3.365 38.205 3.523 ;
      RECT 38.125 3.34 38.165 3.508 ;
      RECT 38.11 3.315 38.125 3.498 ;
      RECT 38.105 3.309 38.11 3.496 ;
      RECT 38.07 3.301 38.105 3.479 ;
      RECT 38.065 3.294 38.07 3.467 ;
      RECT 38.045 3.289 38.065 3.455 ;
      RECT 38.035 3.283 38.045 3.44 ;
      RECT 38.015 3.278 38.035 3.425 ;
      RECT 38.005 3.273 38.015 3.418 ;
      RECT 38 3.271 38.005 3.413 ;
      RECT 37.995 3.27 38 3.41 ;
      RECT 37.955 3.265 37.995 3.406 ;
      RECT 37.935 3.259 37.95 3.401 ;
      RECT 37.9 3.256 37.935 3.398 ;
      RECT 37.89 3.255 37.9 3.396 ;
      RECT 37.83 3.255 37.865 3.393 ;
      RECT 37.785 3.255 37.83 3.393 ;
      RECT 37.735 3.255 37.785 3.396 ;
      RECT 37.72 3.257 37.735 3.398 ;
      RECT 37.705 3.26 37.72 3.399 ;
      RECT 37.695 3.265 37.705 3.4 ;
      RECT 37.665 3.27 37.695 3.405 ;
      RECT 37.655 3.276 37.665 3.413 ;
      RECT 37.645 3.278 37.655 3.417 ;
      RECT 37.635 3.282 37.645 3.421 ;
      RECT 37.61 3.288 37.635 3.429 ;
      RECT 37.6 3.293 37.61 3.437 ;
      RECT 37.585 3.297 37.6 3.441 ;
      RECT 37.55 3.303 37.585 3.449 ;
      RECT 37.53 3.308 37.55 3.459 ;
      RECT 37.5 3.315 37.53 3.468 ;
      RECT 37.455 3.324 37.5 3.482 ;
      RECT 37.45 3.329 37.455 3.493 ;
      RECT 37.43 3.332 37.45 3.494 ;
      RECT 37.4 3.335 37.43 3.492 ;
      RECT 37.365 3.335 37.385 3.488 ;
      RECT 37.295 3.335 37.365 3.479 ;
      RECT 37.28 3.332 37.295 3.471 ;
      RECT 37.24 3.325 37.28 3.466 ;
      RECT 37.215 3.315 37.24 3.459 ;
      RECT 37.21 3.309 37.215 3.456 ;
      RECT 37.17 3.303 37.21 3.453 ;
      RECT 37.155 3.296 37.17 3.448 ;
      RECT 37.135 3.292 37.155 3.443 ;
      RECT 37.12 3.287 37.135 3.439 ;
      RECT 37.105 3.282 37.12 3.437 ;
      RECT 37.09 3.278 37.105 3.436 ;
      RECT 37.075 3.276 37.09 3.432 ;
      RECT 37.065 3.274 37.075 3.427 ;
      RECT 37.05 3.271 37.065 3.423 ;
      RECT 37.04 3.269 37.05 3.418 ;
      RECT 37.02 3.266 37.04 3.414 ;
      RECT 36.975 3.265 37.02 3.412 ;
      RECT 36.915 3.267 36.975 3.413 ;
      RECT 36.895 3.269 36.915 3.415 ;
      RECT 36.865 3.272 36.895 3.416 ;
      RECT 36.815 3.277 36.865 3.418 ;
      RECT 36.81 3.28 36.815 3.42 ;
      RECT 36.8 3.282 36.81 3.423 ;
      RECT 36.795 3.284 36.8 3.426 ;
      RECT 36.745 3.287 36.795 3.433 ;
      RECT 36.725 3.291 36.745 3.445 ;
      RECT 36.715 3.294 36.725 3.451 ;
      RECT 36.705 3.295 36.715 3.454 ;
      RECT 36.666 3.298 36.705 3.456 ;
      RECT 36.58 3.305 36.666 3.459 ;
      RECT 36.506 3.315 36.58 3.463 ;
      RECT 36.42 3.326 36.506 3.468 ;
      RECT 36.405 3.333 36.42 3.47 ;
      RECT 36.35 3.337 36.405 3.471 ;
      RECT 36.336 3.34 36.35 3.473 ;
      RECT 36.25 3.34 36.336 3.475 ;
      RECT 36.21 3.337 36.25 3.478 ;
      RECT 36.186 3.333 36.21 3.48 ;
      RECT 36.1 3.323 36.186 3.483 ;
      RECT 36.07 3.312 36.1 3.484 ;
      RECT 36.051 3.308 36.07 3.483 ;
      RECT 35.965 3.301 36.051 3.48 ;
      RECT 35.905 3.29 35.965 3.477 ;
      RECT 35.885 3.282 35.905 3.475 ;
      RECT 35.85 3.277 35.885 3.474 ;
      RECT 35.825 3.272 35.85 3.473 ;
      RECT 35.795 3.267 35.825 3.472 ;
      RECT 35.77 3.21 35.795 3.471 ;
      RECT 35.755 3.21 35.77 3.495 ;
      RECT 35.56 3.21 35.57 3.495 ;
      RECT 37.335 4.23 37.34 4.37 ;
      RECT 36.995 4.23 37.03 4.368 ;
      RECT 36.57 4.215 36.585 4.36 ;
      RECT 38.4 3.995 38.49 4.255 ;
      RECT 38.23 3.86 38.33 4.255 ;
      RECT 35.265 3.835 35.345 4.045 ;
      RECT 38.355 3.972 38.4 4.255 ;
      RECT 38.345 3.942 38.355 4.255 ;
      RECT 38.33 3.865 38.345 4.255 ;
      RECT 38.145 3.86 38.23 4.22 ;
      RECT 38.14 3.862 38.145 4.215 ;
      RECT 38.135 3.867 38.14 4.215 ;
      RECT 38.1 3.967 38.135 4.215 ;
      RECT 38.09 3.995 38.1 4.215 ;
      RECT 38.08 4.01 38.09 4.215 ;
      RECT 38.07 4.022 38.08 4.215 ;
      RECT 38.065 4.032 38.07 4.215 ;
      RECT 38.05 4.042 38.065 4.217 ;
      RECT 38.045 4.057 38.05 4.219 ;
      RECT 38.03 4.07 38.045 4.221 ;
      RECT 38.025 4.085 38.03 4.224 ;
      RECT 38.005 4.095 38.025 4.228 ;
      RECT 37.99 4.105 38.005 4.231 ;
      RECT 37.955 4.112 37.99 4.236 ;
      RECT 37.911 4.119 37.955 4.244 ;
      RECT 37.825 4.131 37.911 4.257 ;
      RECT 37.8 4.142 37.825 4.268 ;
      RECT 37.77 4.147 37.8 4.273 ;
      RECT 37.735 4.152 37.77 4.281 ;
      RECT 37.705 4.157 37.735 4.288 ;
      RECT 37.68 4.162 37.705 4.293 ;
      RECT 37.615 4.169 37.68 4.302 ;
      RECT 37.545 4.182 37.615 4.318 ;
      RECT 37.515 4.192 37.545 4.33 ;
      RECT 37.49 4.197 37.515 4.337 ;
      RECT 37.435 4.204 37.49 4.345 ;
      RECT 37.43 4.211 37.435 4.35 ;
      RECT 37.425 4.213 37.43 4.351 ;
      RECT 37.41 4.215 37.425 4.353 ;
      RECT 37.405 4.215 37.41 4.356 ;
      RECT 37.34 4.222 37.405 4.363 ;
      RECT 37.305 4.232 37.335 4.373 ;
      RECT 37.288 4.235 37.305 4.375 ;
      RECT 37.202 4.234 37.288 4.374 ;
      RECT 37.116 4.232 37.202 4.371 ;
      RECT 37.03 4.231 37.116 4.369 ;
      RECT 36.929 4.229 36.995 4.368 ;
      RECT 36.843 4.226 36.929 4.366 ;
      RECT 36.757 4.222 36.843 4.364 ;
      RECT 36.671 4.219 36.757 4.363 ;
      RECT 36.585 4.216 36.671 4.361 ;
      RECT 36.485 4.215 36.57 4.358 ;
      RECT 36.435 4.213 36.485 4.356 ;
      RECT 36.415 4.21 36.435 4.354 ;
      RECT 36.395 4.208 36.415 4.351 ;
      RECT 36.37 4.204 36.395 4.348 ;
      RECT 36.325 4.198 36.37 4.343 ;
      RECT 36.285 4.192 36.325 4.335 ;
      RECT 36.26 4.187 36.285 4.328 ;
      RECT 36.205 4.18 36.26 4.32 ;
      RECT 36.181 4.173 36.205 4.313 ;
      RECT 36.095 4.164 36.181 4.303 ;
      RECT 36.065 4.156 36.095 4.293 ;
      RECT 36.035 4.152 36.065 4.288 ;
      RECT 36.03 4.149 36.035 4.285 ;
      RECT 36.025 4.148 36.03 4.285 ;
      RECT 35.95 4.141 36.025 4.278 ;
      RECT 35.911 4.132 35.95 4.267 ;
      RECT 35.825 4.122 35.911 4.255 ;
      RECT 35.785 4.112 35.825 4.243 ;
      RECT 35.746 4.107 35.785 4.236 ;
      RECT 35.66 4.097 35.746 4.225 ;
      RECT 35.62 4.085 35.66 4.214 ;
      RECT 35.585 4.07 35.62 4.207 ;
      RECT 35.575 4.06 35.585 4.204 ;
      RECT 35.555 4.045 35.575 4.202 ;
      RECT 35.525 4.015 35.555 4.198 ;
      RECT 35.515 3.995 35.525 4.193 ;
      RECT 35.51 3.987 35.515 4.19 ;
      RECT 35.505 3.98 35.51 4.188 ;
      RECT 35.49 3.967 35.505 4.181 ;
      RECT 35.485 3.957 35.49 4.173 ;
      RECT 35.48 3.95 35.485 4.168 ;
      RECT 35.475 3.945 35.48 4.164 ;
      RECT 35.46 3.932 35.475 4.156 ;
      RECT 35.455 3.842 35.46 4.145 ;
      RECT 35.45 3.837 35.455 4.138 ;
      RECT 35.375 3.835 35.45 4.098 ;
      RECT 35.345 3.835 35.375 4.053 ;
      RECT 35.25 3.84 35.265 4.04 ;
      RECT 37.735 3.545 37.995 3.805 ;
      RECT 37.72 3.533 37.9 3.77 ;
      RECT 37.715 3.534 37.9 3.768 ;
      RECT 37.7 3.538 37.91 3.758 ;
      RECT 37.695 3.543 37.915 3.728 ;
      RECT 37.7 3.54 37.915 3.758 ;
      RECT 37.715 3.535 37.91 3.768 ;
      RECT 37.735 3.532 37.9 3.805 ;
      RECT 37.735 3.531 37.89 3.805 ;
      RECT 37.76 3.53 37.89 3.805 ;
      RECT 37.32 3.775 37.58 4.035 ;
      RECT 37.195 3.82 37.58 4.03 ;
      RECT 37.185 3.825 37.58 4.025 ;
      RECT 37.2 4.765 37.215 5.075 ;
      RECT 35.795 4.535 35.805 4.665 ;
      RECT 35.575 4.53 35.68 4.665 ;
      RECT 35.49 4.535 35.54 4.665 ;
      RECT 34.04 3.27 34.045 4.375 ;
      RECT 37.295 4.857 37.3 4.993 ;
      RECT 37.29 4.852 37.295 5.053 ;
      RECT 37.285 4.85 37.29 5.066 ;
      RECT 37.27 4.847 37.285 5.068 ;
      RECT 37.265 4.842 37.27 5.07 ;
      RECT 37.26 4.838 37.265 5.073 ;
      RECT 37.245 4.833 37.26 5.075 ;
      RECT 37.215 4.825 37.245 5.075 ;
      RECT 37.176 4.765 37.2 5.075 ;
      RECT 37.09 4.765 37.176 5.072 ;
      RECT 37.06 4.765 37.09 5.065 ;
      RECT 37.035 4.765 37.06 5.058 ;
      RECT 37.01 4.765 37.035 5.05 ;
      RECT 36.995 4.765 37.01 5.043 ;
      RECT 36.97 4.765 36.995 5.035 ;
      RECT 36.955 4.765 36.97 5.028 ;
      RECT 36.915 4.775 36.955 5.017 ;
      RECT 36.905 4.77 36.915 5.007 ;
      RECT 36.901 4.769 36.905 5.004 ;
      RECT 36.815 4.761 36.901 4.987 ;
      RECT 36.782 4.75 36.815 4.964 ;
      RECT 36.696 4.739 36.782 4.942 ;
      RECT 36.61 4.723 36.696 4.911 ;
      RECT 36.54 4.708 36.61 4.883 ;
      RECT 36.53 4.701 36.54 4.87 ;
      RECT 36.5 4.698 36.53 4.86 ;
      RECT 36.475 4.694 36.5 4.853 ;
      RECT 36.46 4.691 36.475 4.848 ;
      RECT 36.455 4.69 36.46 4.843 ;
      RECT 36.425 4.685 36.455 4.836 ;
      RECT 36.42 4.68 36.425 4.831 ;
      RECT 36.405 4.677 36.42 4.826 ;
      RECT 36.4 4.672 36.405 4.821 ;
      RECT 36.38 4.667 36.4 4.818 ;
      RECT 36.365 4.662 36.38 4.81 ;
      RECT 36.35 4.656 36.365 4.805 ;
      RECT 36.32 4.647 36.35 4.798 ;
      RECT 36.315 4.64 36.32 4.79 ;
      RECT 36.31 4.638 36.315 4.788 ;
      RECT 36.305 4.637 36.31 4.785 ;
      RECT 36.265 4.63 36.305 4.778 ;
      RECT 36.251 4.62 36.265 4.768 ;
      RECT 36.2 4.609 36.251 4.756 ;
      RECT 36.175 4.595 36.2 4.742 ;
      RECT 36.15 4.584 36.175 4.734 ;
      RECT 36.13 4.573 36.15 4.728 ;
      RECT 36.12 4.567 36.13 4.723 ;
      RECT 36.115 4.565 36.12 4.719 ;
      RECT 36.095 4.56 36.115 4.714 ;
      RECT 36.065 4.55 36.095 4.704 ;
      RECT 36.06 4.542 36.065 4.697 ;
      RECT 36.045 4.54 36.06 4.693 ;
      RECT 36.025 4.54 36.045 4.688 ;
      RECT 36.02 4.539 36.025 4.686 ;
      RECT 36.015 4.539 36.02 4.683 ;
      RECT 35.975 4.538 36.015 4.678 ;
      RECT 35.95 4.537 35.975 4.673 ;
      RECT 35.89 4.536 35.95 4.67 ;
      RECT 35.805 4.535 35.89 4.668 ;
      RECT 35.766 4.534 35.795 4.665 ;
      RECT 35.68 4.532 35.766 4.665 ;
      RECT 35.54 4.532 35.575 4.665 ;
      RECT 35.45 4.536 35.49 4.668 ;
      RECT 35.435 4.539 35.45 4.675 ;
      RECT 35.425 4.54 35.435 4.682 ;
      RECT 35.4 4.543 35.425 4.687 ;
      RECT 35.395 4.545 35.4 4.69 ;
      RECT 35.345 4.547 35.395 4.691 ;
      RECT 35.306 4.551 35.345 4.693 ;
      RECT 35.22 4.553 35.306 4.696 ;
      RECT 35.202 4.555 35.22 4.698 ;
      RECT 35.116 4.558 35.202 4.7 ;
      RECT 35.03 4.562 35.116 4.703 ;
      RECT 34.993 4.566 35.03 4.706 ;
      RECT 34.907 4.569 34.993 4.709 ;
      RECT 34.821 4.573 34.907 4.712 ;
      RECT 34.735 4.578 34.821 4.716 ;
      RECT 34.715 4.58 34.735 4.719 ;
      RECT 34.695 4.579 34.715 4.72 ;
      RECT 34.646 4.576 34.695 4.721 ;
      RECT 34.56 4.571 34.646 4.724 ;
      RECT 34.51 4.566 34.56 4.726 ;
      RECT 34.486 4.564 34.51 4.727 ;
      RECT 34.4 4.559 34.486 4.729 ;
      RECT 34.375 4.555 34.4 4.728 ;
      RECT 34.365 4.552 34.375 4.726 ;
      RECT 34.355 4.545 34.365 4.723 ;
      RECT 34.35 4.525 34.355 4.718 ;
      RECT 34.34 4.495 34.35 4.713 ;
      RECT 34.325 4.365 34.34 4.704 ;
      RECT 34.32 4.357 34.325 4.697 ;
      RECT 34.3 4.35 34.32 4.689 ;
      RECT 34.295 4.332 34.3 4.681 ;
      RECT 34.285 4.312 34.295 4.676 ;
      RECT 34.28 4.285 34.285 4.672 ;
      RECT 34.275 4.262 34.28 4.669 ;
      RECT 34.255 4.22 34.275 4.661 ;
      RECT 34.22 4.135 34.255 4.645 ;
      RECT 34.215 4.067 34.22 4.633 ;
      RECT 34.2 4.037 34.215 4.627 ;
      RECT 34.195 3.282 34.2 3.528 ;
      RECT 34.185 4.007 34.2 4.618 ;
      RECT 34.19 3.277 34.195 3.56 ;
      RECT 34.185 3.272 34.19 3.603 ;
      RECT 34.18 3.27 34.185 3.638 ;
      RECT 34.165 3.97 34.185 4.608 ;
      RECT 34.175 3.27 34.18 3.675 ;
      RECT 34.16 3.27 34.175 3.773 ;
      RECT 34.16 3.943 34.165 4.601 ;
      RECT 34.155 3.27 34.16 3.848 ;
      RECT 34.155 3.931 34.16 4.598 ;
      RECT 34.15 3.27 34.155 3.88 ;
      RECT 34.15 3.91 34.155 4.595 ;
      RECT 34.145 3.27 34.15 4.592 ;
      RECT 34.11 3.27 34.145 4.578 ;
      RECT 34.095 3.27 34.11 4.56 ;
      RECT 34.075 3.27 34.095 4.55 ;
      RECT 34.05 3.27 34.075 4.533 ;
      RECT 34.045 3.27 34.05 4.483 ;
      RECT 34.035 3.27 34.04 4.313 ;
      RECT 34.03 3.27 34.035 4.22 ;
      RECT 34.025 3.27 34.03 4.133 ;
      RECT 34.02 3.27 34.025 4.065 ;
      RECT 34.015 3.27 34.02 4.008 ;
      RECT 34.005 3.27 34.015 3.903 ;
      RECT 34 3.27 34.005 3.775 ;
      RECT 33.995 3.27 34 3.693 ;
      RECT 33.99 3.272 33.995 3.61 ;
      RECT 33.985 3.277 33.99 3.543 ;
      RECT 33.98 3.282 33.985 3.47 ;
      RECT 36.795 3.6 37.055 3.86 ;
      RECT 36.815 3.567 37.025 3.86 ;
      RECT 36.815 3.565 37.015 3.86 ;
      RECT 36.825 3.552 37.015 3.86 ;
      RECT 36.825 3.55 36.94 3.86 ;
      RECT 36.3 3.675 36.475 3.955 ;
      RECT 36.295 3.675 36.475 3.953 ;
      RECT 36.295 3.675 36.49 3.95 ;
      RECT 36.285 3.675 36.49 3.948 ;
      RECT 36.23 3.675 36.49 3.935 ;
      RECT 36.23 3.75 36.495 3.913 ;
      RECT 35.76 4.873 35.765 5.08 ;
      RECT 35.71 4.867 35.76 5.079 ;
      RECT 35.677 4.881 35.77 5.078 ;
      RECT 35.591 4.881 35.77 5.077 ;
      RECT 35.505 4.881 35.77 5.076 ;
      RECT 35.505 4.98 35.775 5.073 ;
      RECT 35.5 4.98 35.775 5.068 ;
      RECT 35.495 4.98 35.775 5.05 ;
      RECT 35.49 4.98 35.775 5.033 ;
      RECT 35.45 4.765 35.71 5.025 ;
      RECT 34.91 3.915 34.996 4.329 ;
      RECT 34.91 3.915 35.035 4.326 ;
      RECT 34.91 3.915 35.055 4.316 ;
      RECT 34.865 3.915 35.055 4.313 ;
      RECT 34.865 4.067 35.065 4.303 ;
      RECT 34.865 4.088 35.07 4.297 ;
      RECT 34.865 4.106 35.075 4.293 ;
      RECT 34.865 4.126 35.085 4.288 ;
      RECT 34.84 4.126 35.085 4.285 ;
      RECT 34.83 4.126 35.085 4.263 ;
      RECT 34.83 4.142 35.09 4.233 ;
      RECT 34.795 3.915 35.055 4.22 ;
      RECT 34.795 4.154 35.095 4.175 ;
      RECT 32.455 10.06 32.75 10.29 ;
      RECT 32.515 8.58 32.685 10.29 ;
      RECT 32.51 8.95 32.86 9.3 ;
      RECT 32.455 8.58 32.745 8.81 ;
      RECT 31.465 10.06 31.76 10.29 ;
      RECT 31.525 8.58 31.695 10.29 ;
      RECT 31.465 8.58 31.755 8.81 ;
      RECT 31.465 8.615 32.315 8.775 ;
      RECT 32.15 8.21 32.315 8.775 ;
      RECT 31.465 8.61 31.86 8.775 ;
      RECT 32.085 8.21 32.375 8.44 ;
      RECT 32.085 8.24 32.545 8.41 ;
      RECT 32.05 4.025 32.37 4.26 ;
      RECT 32.05 4.055 32.54 4.225 ;
      RECT 32.05 3.69 32.24 4.26 ;
      RECT 31.465 3.655 31.755 3.885 ;
      RECT 31.465 3.69 32.24 3.86 ;
      RECT 31.525 2.175 31.695 3.885 ;
      RECT 31.465 2.175 31.76 2.405 ;
      RECT 31.095 4.025 31.385 4.255 ;
      RECT 31.095 4.055 31.555 4.225 ;
      RECT 31.16 2.95 31.325 4.255 ;
      RECT 29.675 2.915 29.965 3.145 ;
      RECT 29.675 2.95 31.325 3.12 ;
      RECT 29.735 2.175 29.905 3.145 ;
      RECT 29.675 2.175 29.965 2.405 ;
      RECT 29.675 10.06 29.965 10.29 ;
      RECT 29.735 9.32 29.905 10.29 ;
      RECT 29.735 9.41 31.325 9.58 ;
      RECT 31.155 8.21 31.325 9.58 ;
      RECT 29.675 9.32 29.965 9.55 ;
      RECT 31.095 8.21 31.385 8.44 ;
      RECT 31.095 8.24 31.555 8.41 ;
      RECT 27.725 4 28.065 4.35 ;
      RECT 27.815 3.32 27.985 4.35 ;
      RECT 30.105 3.26 30.455 3.61 ;
      RECT 27.815 3.32 30.455 3.49 ;
      RECT 29.935 3.315 30.455 3.49 ;
      RECT 30.13 8.945 30.455 9.27 ;
      RECT 24.67 8.895 25.02 9.245 ;
      RECT 30.105 8.95 30.455 9.18 ;
      RECT 24.47 8.95 25.02 9.18 ;
      RECT 29.935 8.975 30.455 9.15 ;
      RECT 24.3 8.98 25.02 9.15 ;
      RECT 24.35 8.975 30.455 9.145 ;
      RECT 29.33 3.66 29.65 3.98 ;
      RECT 29.305 3.655 29.595 3.885 ;
      RECT 29.3 3.685 29.65 3.86 ;
      RECT 29.13 3.685 29.65 3.855 ;
      RECT 29.33 8.545 29.65 8.835 ;
      RECT 29.305 8.58 29.65 8.81 ;
      RECT 29.13 8.61 29.65 8.78 ;
      RECT 25.02 4.28 25.17 4.555 ;
      RECT 25.56 3.36 25.565 3.58 ;
      RECT 26.71 3.56 26.725 3.758 ;
      RECT 26.675 3.552 26.71 3.765 ;
      RECT 26.645 3.545 26.675 3.765 ;
      RECT 26.59 3.51 26.645 3.765 ;
      RECT 26.525 3.447 26.59 3.765 ;
      RECT 26.52 3.412 26.525 3.763 ;
      RECT 26.515 3.407 26.52 3.755 ;
      RECT 26.51 3.402 26.515 3.741 ;
      RECT 26.505 3.399 26.51 3.734 ;
      RECT 26.46 3.389 26.505 3.685 ;
      RECT 26.44 3.376 26.46 3.62 ;
      RECT 26.435 3.371 26.44 3.593 ;
      RECT 26.43 3.37 26.435 3.586 ;
      RECT 26.425 3.369 26.43 3.579 ;
      RECT 26.34 3.354 26.425 3.525 ;
      RECT 26.31 3.335 26.34 3.475 ;
      RECT 26.23 3.318 26.31 3.46 ;
      RECT 26.195 3.305 26.23 3.445 ;
      RECT 26.187 3.305 26.195 3.44 ;
      RECT 26.101 3.306 26.187 3.44 ;
      RECT 26.015 3.308 26.101 3.44 ;
      RECT 25.99 3.309 26.015 3.444 ;
      RECT 25.915 3.315 25.99 3.459 ;
      RECT 25.832 3.327 25.915 3.483 ;
      RECT 25.746 3.34 25.832 3.509 ;
      RECT 25.66 3.353 25.746 3.535 ;
      RECT 25.625 3.362 25.66 3.554 ;
      RECT 25.575 3.362 25.625 3.567 ;
      RECT 25.565 3.36 25.575 3.578 ;
      RECT 25.55 3.357 25.56 3.58 ;
      RECT 25.535 3.349 25.55 3.588 ;
      RECT 25.52 3.341 25.535 3.608 ;
      RECT 25.515 3.336 25.52 3.665 ;
      RECT 25.5 3.331 25.515 3.738 ;
      RECT 25.495 3.326 25.5 3.78 ;
      RECT 25.49 3.324 25.495 3.808 ;
      RECT 25.485 3.322 25.49 3.83 ;
      RECT 25.475 3.318 25.485 3.873 ;
      RECT 25.47 3.315 25.475 3.898 ;
      RECT 25.465 3.313 25.47 3.918 ;
      RECT 25.46 3.311 25.465 3.942 ;
      RECT 25.455 3.307 25.46 3.965 ;
      RECT 25.45 3.303 25.455 3.988 ;
      RECT 25.415 3.293 25.45 4.095 ;
      RECT 25.41 3.283 25.415 4.193 ;
      RECT 25.405 3.281 25.41 4.22 ;
      RECT 25.4 3.28 25.405 4.24 ;
      RECT 25.395 3.272 25.4 4.26 ;
      RECT 25.39 3.267 25.395 4.295 ;
      RECT 25.385 3.265 25.39 4.313 ;
      RECT 25.38 3.265 25.385 4.338 ;
      RECT 25.375 3.265 25.38 4.36 ;
      RECT 25.34 3.265 25.375 4.403 ;
      RECT 25.315 3.265 25.34 4.432 ;
      RECT 25.305 3.265 25.315 3.618 ;
      RECT 25.308 3.675 25.315 4.442 ;
      RECT 25.305 3.732 25.308 4.445 ;
      RECT 25.3 3.265 25.305 3.59 ;
      RECT 25.3 3.782 25.305 4.448 ;
      RECT 25.29 3.265 25.3 3.58 ;
      RECT 25.295 3.835 25.3 4.451 ;
      RECT 25.29 3.92 25.295 4.455 ;
      RECT 25.28 3.265 25.29 3.568 ;
      RECT 25.285 3.967 25.29 4.459 ;
      RECT 25.28 4.042 25.285 4.463 ;
      RECT 25.245 3.265 25.28 3.543 ;
      RECT 25.27 4.125 25.28 4.468 ;
      RECT 25.26 4.192 25.27 4.475 ;
      RECT 25.255 4.22 25.26 4.48 ;
      RECT 25.245 4.233 25.255 4.486 ;
      RECT 25.2 3.265 25.245 3.5 ;
      RECT 25.24 4.238 25.245 4.493 ;
      RECT 25.2 4.255 25.24 4.555 ;
      RECT 25.195 3.267 25.2 3.473 ;
      RECT 25.17 4.275 25.2 4.555 ;
      RECT 25.19 3.272 25.195 3.445 ;
      RECT 24.98 4.284 25.02 4.555 ;
      RECT 24.955 4.292 24.98 4.525 ;
      RECT 24.91 4.3 24.955 4.525 ;
      RECT 24.895 4.305 24.91 4.52 ;
      RECT 24.885 4.305 24.895 4.514 ;
      RECT 24.875 4.312 24.885 4.511 ;
      RECT 24.87 4.35 24.875 4.5 ;
      RECT 24.865 4.412 24.87 4.478 ;
      RECT 26.135 4.287 26.32 4.51 ;
      RECT 26.135 4.302 26.325 4.506 ;
      RECT 26.125 3.575 26.21 4.505 ;
      RECT 26.125 4.302 26.33 4.499 ;
      RECT 26.12 4.31 26.33 4.498 ;
      RECT 26.325 4.03 26.645 4.35 ;
      RECT 26.12 4.202 26.29 4.293 ;
      RECT 26.115 4.202 26.29 4.275 ;
      RECT 26.105 4.01 26.24 4.25 ;
      RECT 26.1 4.01 26.24 4.195 ;
      RECT 26.06 3.59 26.23 4.095 ;
      RECT 26.045 3.59 26.23 3.965 ;
      RECT 26.04 3.59 26.23 3.918 ;
      RECT 26.035 3.59 26.23 3.898 ;
      RECT 26.03 3.59 26.23 3.873 ;
      RECT 26 3.59 26.26 3.85 ;
      RECT 26.01 3.587 26.22 3.85 ;
      RECT 26.135 3.582 26.22 4.51 ;
      RECT 26.02 3.575 26.21 3.85 ;
      RECT 26.015 3.58 26.21 3.85 ;
      RECT 24.845 3.792 25.03 4.005 ;
      RECT 24.845 3.8 25.04 3.998 ;
      RECT 24.825 3.8 25.04 3.995 ;
      RECT 24.82 3.8 25.04 3.98 ;
      RECT 24.75 3.715 25.01 3.975 ;
      RECT 24.75 3.86 25.045 3.888 ;
      RECT 24.405 4.315 24.665 4.575 ;
      RECT 24.43 4.26 24.625 4.575 ;
      RECT 24.425 4.009 24.605 4.303 ;
      RECT 24.425 4.015 24.615 4.303 ;
      RECT 24.405 4.017 24.615 4.248 ;
      RECT 24.4 4.027 24.615 4.115 ;
      RECT 24.43 4.007 24.605 4.575 ;
      RECT 24.516 4.005 24.605 4.575 ;
      RECT 24.375 3.225 24.41 3.595 ;
      RECT 24.165 3.335 24.17 3.595 ;
      RECT 24.41 3.232 24.425 3.595 ;
      RECT 24.3 3.225 24.375 3.673 ;
      RECT 24.29 3.225 24.3 3.758 ;
      RECT 24.265 3.225 24.29 3.793 ;
      RECT 24.225 3.225 24.265 3.861 ;
      RECT 24.215 3.232 24.225 3.913 ;
      RECT 24.185 3.335 24.215 3.954 ;
      RECT 24.18 3.335 24.185 3.993 ;
      RECT 24.17 3.335 24.18 4.013 ;
      RECT 24.165 3.63 24.17 4.05 ;
      RECT 24.16 3.647 24.165 4.07 ;
      RECT 24.145 3.71 24.16 4.11 ;
      RECT 24.14 3.753 24.145 4.145 ;
      RECT 24.135 3.761 24.14 4.158 ;
      RECT 24.125 3.775 24.135 4.18 ;
      RECT 24.1 3.81 24.125 4.245 ;
      RECT 24.09 3.845 24.1 4.308 ;
      RECT 24.07 3.875 24.09 4.369 ;
      RECT 24.055 3.911 24.07 4.436 ;
      RECT 24.045 3.939 24.055 4.475 ;
      RECT 24.035 3.961 24.045 4.495 ;
      RECT 24.03 3.971 24.035 4.506 ;
      RECT 24.025 3.98 24.03 4.509 ;
      RECT 24.015 3.998 24.025 4.513 ;
      RECT 24.005 4.016 24.015 4.514 ;
      RECT 23.98 4.055 24.005 4.511 ;
      RECT 23.96 4.097 23.98 4.508 ;
      RECT 23.945 4.135 23.96 4.507 ;
      RECT 23.91 4.17 23.945 4.504 ;
      RECT 23.905 4.192 23.91 4.502 ;
      RECT 23.84 4.232 23.905 4.499 ;
      RECT 23.835 4.272 23.84 4.495 ;
      RECT 23.82 4.282 23.835 4.486 ;
      RECT 23.81 4.402 23.82 4.471 ;
      RECT 24.29 4.815 24.3 5.075 ;
      RECT 24.29 4.818 24.31 5.074 ;
      RECT 24.28 4.808 24.29 5.073 ;
      RECT 24.27 4.823 24.35 5.069 ;
      RECT 24.255 4.802 24.27 5.067 ;
      RECT 24.23 4.827 24.355 5.063 ;
      RECT 24.215 4.787 24.23 5.058 ;
      RECT 24.215 4.829 24.365 5.057 ;
      RECT 24.215 4.837 24.38 5.05 ;
      RECT 24.155 4.774 24.215 5.04 ;
      RECT 24.145 4.761 24.155 5.022 ;
      RECT 24.12 4.751 24.145 5.012 ;
      RECT 24.115 4.741 24.12 5.004 ;
      RECT 24.05 4.837 24.38 4.986 ;
      RECT 23.965 4.837 24.38 4.948 ;
      RECT 23.855 4.665 24.115 4.925 ;
      RECT 24.23 4.795 24.255 5.063 ;
      RECT 24.27 4.805 24.28 5.069 ;
      RECT 23.855 4.813 24.295 4.925 ;
      RECT 24.04 10.06 24.33 10.29 ;
      RECT 24.1 9.32 24.27 10.29 ;
      RECT 24 9.345 24.37 9.715 ;
      RECT 24.04 9.32 24.33 9.715 ;
      RECT 23.07 4.57 23.1 4.87 ;
      RECT 22.845 4.555 22.85 4.83 ;
      RECT 22.645 4.555 22.8 4.815 ;
      RECT 23.945 3.27 23.975 3.53 ;
      RECT 23.935 3.27 23.945 3.638 ;
      RECT 23.915 3.27 23.935 3.648 ;
      RECT 23.9 3.27 23.915 3.66 ;
      RECT 23.845 3.27 23.9 3.71 ;
      RECT 23.83 3.27 23.845 3.758 ;
      RECT 23.8 3.27 23.83 3.793 ;
      RECT 23.745 3.27 23.8 3.855 ;
      RECT 23.725 3.27 23.745 3.923 ;
      RECT 23.72 3.27 23.725 3.953 ;
      RECT 23.715 3.27 23.72 3.965 ;
      RECT 23.71 3.387 23.715 3.983 ;
      RECT 23.69 3.405 23.71 4.008 ;
      RECT 23.67 3.432 23.69 4.058 ;
      RECT 23.665 3.452 23.67 4.089 ;
      RECT 23.66 3.46 23.665 4.106 ;
      RECT 23.645 3.486 23.66 4.135 ;
      RECT 23.63 3.528 23.645 4.17 ;
      RECT 23.625 3.557 23.63 4.193 ;
      RECT 23.62 3.572 23.625 4.206 ;
      RECT 23.615 3.595 23.62 4.217 ;
      RECT 23.605 3.615 23.615 4.235 ;
      RECT 23.595 3.645 23.605 4.258 ;
      RECT 23.59 3.667 23.595 4.278 ;
      RECT 23.585 3.682 23.59 4.293 ;
      RECT 23.57 3.712 23.585 4.32 ;
      RECT 23.565 3.742 23.57 4.346 ;
      RECT 23.56 3.76 23.565 4.358 ;
      RECT 23.55 3.79 23.56 4.377 ;
      RECT 23.54 3.815 23.55 4.402 ;
      RECT 23.535 3.835 23.54 4.421 ;
      RECT 23.53 3.852 23.535 4.434 ;
      RECT 23.52 3.878 23.53 4.453 ;
      RECT 23.51 3.916 23.52 4.48 ;
      RECT 23.505 3.942 23.51 4.5 ;
      RECT 23.5 3.952 23.505 4.51 ;
      RECT 23.495 3.965 23.5 4.525 ;
      RECT 23.49 3.98 23.495 4.535 ;
      RECT 23.485 4.002 23.49 4.55 ;
      RECT 23.48 4.02 23.485 4.561 ;
      RECT 23.475 4.03 23.48 4.572 ;
      RECT 23.47 4.038 23.475 4.584 ;
      RECT 23.465 4.046 23.47 4.595 ;
      RECT 23.46 4.072 23.465 4.608 ;
      RECT 23.45 4.1 23.46 4.621 ;
      RECT 23.445 4.13 23.45 4.63 ;
      RECT 23.44 4.145 23.445 4.637 ;
      RECT 23.425 4.17 23.44 4.644 ;
      RECT 23.42 4.192 23.425 4.65 ;
      RECT 23.415 4.217 23.42 4.653 ;
      RECT 23.406 4.245 23.415 4.657 ;
      RECT 23.4 4.262 23.406 4.662 ;
      RECT 23.395 4.28 23.4 4.666 ;
      RECT 23.39 4.292 23.395 4.669 ;
      RECT 23.385 4.313 23.39 4.673 ;
      RECT 23.38 4.331 23.385 4.676 ;
      RECT 23.375 4.345 23.38 4.679 ;
      RECT 23.37 4.362 23.375 4.682 ;
      RECT 23.365 4.375 23.37 4.685 ;
      RECT 23.34 4.412 23.365 4.693 ;
      RECT 23.335 4.457 23.34 4.702 ;
      RECT 23.33 4.485 23.335 4.705 ;
      RECT 23.32 4.505 23.33 4.709 ;
      RECT 23.315 4.525 23.32 4.714 ;
      RECT 23.31 4.54 23.315 4.717 ;
      RECT 23.29 4.55 23.31 4.724 ;
      RECT 23.225 4.557 23.29 4.75 ;
      RECT 23.19 4.56 23.225 4.778 ;
      RECT 23.175 4.563 23.19 4.793 ;
      RECT 23.165 4.564 23.175 4.808 ;
      RECT 23.155 4.565 23.165 4.825 ;
      RECT 23.15 4.565 23.155 4.84 ;
      RECT 23.145 4.565 23.15 4.848 ;
      RECT 23.13 4.566 23.145 4.863 ;
      RECT 23.1 4.568 23.13 4.87 ;
      RECT 22.99 4.575 23.07 4.87 ;
      RECT 22.945 4.58 22.99 4.87 ;
      RECT 22.935 4.581 22.945 4.86 ;
      RECT 22.925 4.582 22.935 4.853 ;
      RECT 22.905 4.584 22.925 4.848 ;
      RECT 22.895 4.555 22.905 4.843 ;
      RECT 22.85 4.555 22.895 4.835 ;
      RECT 22.82 4.555 22.845 4.825 ;
      RECT 22.8 4.555 22.82 4.818 ;
      RECT 23.08 3.355 23.34 3.615 ;
      RECT 22.96 3.37 22.97 3.535 ;
      RECT 22.945 3.37 22.95 3.53 ;
      RECT 20.31 3.21 20.495 3.5 ;
      RECT 22.125 3.335 22.14 3.49 ;
      RECT 20.275 3.21 20.3 3.47 ;
      RECT 22.69 3.26 22.695 3.402 ;
      RECT 22.605 3.255 22.63 3.395 ;
      RECT 23.005 3.372 23.08 3.565 ;
      RECT 22.99 3.37 23.005 3.548 ;
      RECT 22.97 3.37 22.99 3.54 ;
      RECT 22.95 3.37 22.96 3.533 ;
      RECT 22.905 3.365 22.945 3.523 ;
      RECT 22.865 3.34 22.905 3.508 ;
      RECT 22.85 3.315 22.865 3.498 ;
      RECT 22.845 3.309 22.85 3.496 ;
      RECT 22.81 3.301 22.845 3.479 ;
      RECT 22.805 3.294 22.81 3.467 ;
      RECT 22.785 3.289 22.805 3.455 ;
      RECT 22.775 3.283 22.785 3.44 ;
      RECT 22.755 3.278 22.775 3.425 ;
      RECT 22.745 3.273 22.755 3.418 ;
      RECT 22.74 3.271 22.745 3.413 ;
      RECT 22.735 3.27 22.74 3.41 ;
      RECT 22.695 3.265 22.735 3.406 ;
      RECT 22.675 3.259 22.69 3.401 ;
      RECT 22.64 3.256 22.675 3.398 ;
      RECT 22.63 3.255 22.64 3.396 ;
      RECT 22.57 3.255 22.605 3.393 ;
      RECT 22.525 3.255 22.57 3.393 ;
      RECT 22.475 3.255 22.525 3.396 ;
      RECT 22.46 3.257 22.475 3.398 ;
      RECT 22.445 3.26 22.46 3.399 ;
      RECT 22.435 3.265 22.445 3.4 ;
      RECT 22.405 3.27 22.435 3.405 ;
      RECT 22.395 3.276 22.405 3.413 ;
      RECT 22.385 3.278 22.395 3.417 ;
      RECT 22.375 3.282 22.385 3.421 ;
      RECT 22.35 3.288 22.375 3.429 ;
      RECT 22.34 3.293 22.35 3.437 ;
      RECT 22.325 3.297 22.34 3.441 ;
      RECT 22.29 3.303 22.325 3.449 ;
      RECT 22.27 3.308 22.29 3.459 ;
      RECT 22.24 3.315 22.27 3.468 ;
      RECT 22.195 3.324 22.24 3.482 ;
      RECT 22.19 3.329 22.195 3.493 ;
      RECT 22.17 3.332 22.19 3.494 ;
      RECT 22.14 3.335 22.17 3.492 ;
      RECT 22.105 3.335 22.125 3.488 ;
      RECT 22.035 3.335 22.105 3.479 ;
      RECT 22.02 3.332 22.035 3.471 ;
      RECT 21.98 3.325 22.02 3.466 ;
      RECT 21.955 3.315 21.98 3.459 ;
      RECT 21.95 3.309 21.955 3.456 ;
      RECT 21.91 3.303 21.95 3.453 ;
      RECT 21.895 3.296 21.91 3.448 ;
      RECT 21.875 3.292 21.895 3.443 ;
      RECT 21.86 3.287 21.875 3.439 ;
      RECT 21.845 3.282 21.86 3.437 ;
      RECT 21.83 3.278 21.845 3.436 ;
      RECT 21.815 3.276 21.83 3.432 ;
      RECT 21.805 3.274 21.815 3.427 ;
      RECT 21.79 3.271 21.805 3.423 ;
      RECT 21.78 3.269 21.79 3.418 ;
      RECT 21.76 3.266 21.78 3.414 ;
      RECT 21.715 3.265 21.76 3.412 ;
      RECT 21.655 3.267 21.715 3.413 ;
      RECT 21.635 3.269 21.655 3.415 ;
      RECT 21.605 3.272 21.635 3.416 ;
      RECT 21.555 3.277 21.605 3.418 ;
      RECT 21.55 3.28 21.555 3.42 ;
      RECT 21.54 3.282 21.55 3.423 ;
      RECT 21.535 3.284 21.54 3.426 ;
      RECT 21.485 3.287 21.535 3.433 ;
      RECT 21.465 3.291 21.485 3.445 ;
      RECT 21.455 3.294 21.465 3.451 ;
      RECT 21.445 3.295 21.455 3.454 ;
      RECT 21.406 3.298 21.445 3.456 ;
      RECT 21.32 3.305 21.406 3.459 ;
      RECT 21.246 3.315 21.32 3.463 ;
      RECT 21.16 3.326 21.246 3.468 ;
      RECT 21.145 3.333 21.16 3.47 ;
      RECT 21.09 3.337 21.145 3.471 ;
      RECT 21.076 3.34 21.09 3.473 ;
      RECT 20.99 3.34 21.076 3.475 ;
      RECT 20.95 3.337 20.99 3.478 ;
      RECT 20.926 3.333 20.95 3.48 ;
      RECT 20.84 3.323 20.926 3.483 ;
      RECT 20.81 3.312 20.84 3.484 ;
      RECT 20.791 3.308 20.81 3.483 ;
      RECT 20.705 3.301 20.791 3.48 ;
      RECT 20.645 3.29 20.705 3.477 ;
      RECT 20.625 3.282 20.645 3.475 ;
      RECT 20.59 3.277 20.625 3.474 ;
      RECT 20.565 3.272 20.59 3.473 ;
      RECT 20.535 3.267 20.565 3.472 ;
      RECT 20.51 3.21 20.535 3.471 ;
      RECT 20.495 3.21 20.51 3.495 ;
      RECT 20.3 3.21 20.31 3.495 ;
      RECT 22.075 4.23 22.08 4.37 ;
      RECT 21.735 4.23 21.77 4.368 ;
      RECT 21.31 4.215 21.325 4.36 ;
      RECT 23.14 3.995 23.23 4.255 ;
      RECT 22.97 3.86 23.07 4.255 ;
      RECT 20.005 3.835 20.085 4.045 ;
      RECT 23.095 3.972 23.14 4.255 ;
      RECT 23.085 3.942 23.095 4.255 ;
      RECT 23.07 3.865 23.085 4.255 ;
      RECT 22.885 3.86 22.97 4.22 ;
      RECT 22.88 3.862 22.885 4.215 ;
      RECT 22.875 3.867 22.88 4.215 ;
      RECT 22.84 3.967 22.875 4.215 ;
      RECT 22.83 3.995 22.84 4.215 ;
      RECT 22.82 4.01 22.83 4.215 ;
      RECT 22.81 4.022 22.82 4.215 ;
      RECT 22.805 4.032 22.81 4.215 ;
      RECT 22.79 4.042 22.805 4.217 ;
      RECT 22.785 4.057 22.79 4.219 ;
      RECT 22.77 4.07 22.785 4.221 ;
      RECT 22.765 4.085 22.77 4.224 ;
      RECT 22.745 4.095 22.765 4.228 ;
      RECT 22.73 4.105 22.745 4.231 ;
      RECT 22.695 4.112 22.73 4.236 ;
      RECT 22.651 4.119 22.695 4.244 ;
      RECT 22.565 4.131 22.651 4.257 ;
      RECT 22.54 4.142 22.565 4.268 ;
      RECT 22.51 4.147 22.54 4.273 ;
      RECT 22.475 4.152 22.51 4.281 ;
      RECT 22.445 4.157 22.475 4.288 ;
      RECT 22.42 4.162 22.445 4.293 ;
      RECT 22.355 4.169 22.42 4.302 ;
      RECT 22.285 4.182 22.355 4.318 ;
      RECT 22.255 4.192 22.285 4.33 ;
      RECT 22.23 4.197 22.255 4.337 ;
      RECT 22.175 4.204 22.23 4.345 ;
      RECT 22.17 4.211 22.175 4.35 ;
      RECT 22.165 4.213 22.17 4.351 ;
      RECT 22.15 4.215 22.165 4.353 ;
      RECT 22.145 4.215 22.15 4.356 ;
      RECT 22.08 4.222 22.145 4.363 ;
      RECT 22.045 4.232 22.075 4.373 ;
      RECT 22.028 4.235 22.045 4.375 ;
      RECT 21.942 4.234 22.028 4.374 ;
      RECT 21.856 4.232 21.942 4.371 ;
      RECT 21.77 4.231 21.856 4.369 ;
      RECT 21.669 4.229 21.735 4.368 ;
      RECT 21.583 4.226 21.669 4.366 ;
      RECT 21.497 4.222 21.583 4.364 ;
      RECT 21.411 4.219 21.497 4.363 ;
      RECT 21.325 4.216 21.411 4.361 ;
      RECT 21.225 4.215 21.31 4.358 ;
      RECT 21.175 4.213 21.225 4.356 ;
      RECT 21.155 4.21 21.175 4.354 ;
      RECT 21.135 4.208 21.155 4.351 ;
      RECT 21.11 4.204 21.135 4.348 ;
      RECT 21.065 4.198 21.11 4.343 ;
      RECT 21.025 4.192 21.065 4.335 ;
      RECT 21 4.187 21.025 4.328 ;
      RECT 20.945 4.18 21 4.32 ;
      RECT 20.921 4.173 20.945 4.313 ;
      RECT 20.835 4.164 20.921 4.303 ;
      RECT 20.805 4.156 20.835 4.293 ;
      RECT 20.775 4.152 20.805 4.288 ;
      RECT 20.77 4.149 20.775 4.285 ;
      RECT 20.765 4.148 20.77 4.285 ;
      RECT 20.69 4.141 20.765 4.278 ;
      RECT 20.651 4.132 20.69 4.267 ;
      RECT 20.565 4.122 20.651 4.255 ;
      RECT 20.525 4.112 20.565 4.243 ;
      RECT 20.486 4.107 20.525 4.236 ;
      RECT 20.4 4.097 20.486 4.225 ;
      RECT 20.36 4.085 20.4 4.214 ;
      RECT 20.325 4.07 20.36 4.207 ;
      RECT 20.315 4.06 20.325 4.204 ;
      RECT 20.295 4.045 20.315 4.202 ;
      RECT 20.265 4.015 20.295 4.198 ;
      RECT 20.255 3.995 20.265 4.193 ;
      RECT 20.25 3.987 20.255 4.19 ;
      RECT 20.245 3.98 20.25 4.188 ;
      RECT 20.23 3.967 20.245 4.181 ;
      RECT 20.225 3.957 20.23 4.173 ;
      RECT 20.22 3.95 20.225 4.168 ;
      RECT 20.215 3.945 20.22 4.164 ;
      RECT 20.2 3.932 20.215 4.156 ;
      RECT 20.195 3.842 20.2 4.145 ;
      RECT 20.19 3.837 20.195 4.138 ;
      RECT 20.115 3.835 20.19 4.098 ;
      RECT 20.085 3.835 20.115 4.053 ;
      RECT 19.99 3.84 20.005 4.04 ;
      RECT 22.475 3.545 22.735 3.805 ;
      RECT 22.46 3.533 22.64 3.77 ;
      RECT 22.455 3.534 22.64 3.768 ;
      RECT 22.44 3.538 22.65 3.758 ;
      RECT 22.435 3.543 22.655 3.728 ;
      RECT 22.44 3.54 22.655 3.758 ;
      RECT 22.455 3.535 22.65 3.768 ;
      RECT 22.475 3.532 22.64 3.805 ;
      RECT 22.475 3.531 22.63 3.805 ;
      RECT 22.5 3.53 22.63 3.805 ;
      RECT 22.06 3.775 22.32 4.035 ;
      RECT 21.935 3.82 22.32 4.03 ;
      RECT 21.925 3.825 22.32 4.025 ;
      RECT 21.94 4.765 21.955 5.075 ;
      RECT 20.535 4.535 20.545 4.665 ;
      RECT 20.315 4.53 20.42 4.665 ;
      RECT 20.23 4.535 20.28 4.665 ;
      RECT 18.78 3.27 18.785 4.375 ;
      RECT 22.035 4.857 22.04 4.993 ;
      RECT 22.03 4.852 22.035 5.053 ;
      RECT 22.025 4.85 22.03 5.066 ;
      RECT 22.01 4.847 22.025 5.068 ;
      RECT 22.005 4.842 22.01 5.07 ;
      RECT 22 4.838 22.005 5.073 ;
      RECT 21.985 4.833 22 5.075 ;
      RECT 21.955 4.825 21.985 5.075 ;
      RECT 21.916 4.765 21.94 5.075 ;
      RECT 21.83 4.765 21.916 5.072 ;
      RECT 21.8 4.765 21.83 5.065 ;
      RECT 21.775 4.765 21.8 5.058 ;
      RECT 21.75 4.765 21.775 5.05 ;
      RECT 21.735 4.765 21.75 5.043 ;
      RECT 21.71 4.765 21.735 5.035 ;
      RECT 21.695 4.765 21.71 5.028 ;
      RECT 21.655 4.775 21.695 5.017 ;
      RECT 21.645 4.77 21.655 5.007 ;
      RECT 21.641 4.769 21.645 5.004 ;
      RECT 21.555 4.761 21.641 4.987 ;
      RECT 21.522 4.75 21.555 4.964 ;
      RECT 21.436 4.739 21.522 4.942 ;
      RECT 21.35 4.723 21.436 4.911 ;
      RECT 21.28 4.708 21.35 4.883 ;
      RECT 21.27 4.701 21.28 4.87 ;
      RECT 21.24 4.698 21.27 4.86 ;
      RECT 21.215 4.694 21.24 4.853 ;
      RECT 21.2 4.691 21.215 4.848 ;
      RECT 21.195 4.69 21.2 4.843 ;
      RECT 21.165 4.685 21.195 4.836 ;
      RECT 21.16 4.68 21.165 4.831 ;
      RECT 21.145 4.677 21.16 4.826 ;
      RECT 21.14 4.672 21.145 4.821 ;
      RECT 21.12 4.667 21.14 4.818 ;
      RECT 21.105 4.662 21.12 4.81 ;
      RECT 21.09 4.656 21.105 4.805 ;
      RECT 21.06 4.647 21.09 4.798 ;
      RECT 21.055 4.64 21.06 4.79 ;
      RECT 21.05 4.638 21.055 4.788 ;
      RECT 21.045 4.637 21.05 4.785 ;
      RECT 21.005 4.63 21.045 4.778 ;
      RECT 20.991 4.62 21.005 4.768 ;
      RECT 20.94 4.609 20.991 4.756 ;
      RECT 20.915 4.595 20.94 4.742 ;
      RECT 20.89 4.584 20.915 4.734 ;
      RECT 20.87 4.573 20.89 4.728 ;
      RECT 20.86 4.567 20.87 4.723 ;
      RECT 20.855 4.565 20.86 4.719 ;
      RECT 20.835 4.56 20.855 4.714 ;
      RECT 20.805 4.55 20.835 4.704 ;
      RECT 20.8 4.542 20.805 4.697 ;
      RECT 20.785 4.54 20.8 4.693 ;
      RECT 20.765 4.54 20.785 4.688 ;
      RECT 20.76 4.539 20.765 4.686 ;
      RECT 20.755 4.539 20.76 4.683 ;
      RECT 20.715 4.538 20.755 4.678 ;
      RECT 20.69 4.537 20.715 4.673 ;
      RECT 20.63 4.536 20.69 4.67 ;
      RECT 20.545 4.535 20.63 4.668 ;
      RECT 20.506 4.534 20.535 4.665 ;
      RECT 20.42 4.532 20.506 4.665 ;
      RECT 20.28 4.532 20.315 4.665 ;
      RECT 20.19 4.536 20.23 4.668 ;
      RECT 20.175 4.539 20.19 4.675 ;
      RECT 20.165 4.54 20.175 4.682 ;
      RECT 20.14 4.543 20.165 4.687 ;
      RECT 20.135 4.545 20.14 4.69 ;
      RECT 20.085 4.547 20.135 4.691 ;
      RECT 20.046 4.551 20.085 4.693 ;
      RECT 19.96 4.553 20.046 4.696 ;
      RECT 19.942 4.555 19.96 4.698 ;
      RECT 19.856 4.558 19.942 4.7 ;
      RECT 19.77 4.562 19.856 4.703 ;
      RECT 19.733 4.566 19.77 4.706 ;
      RECT 19.647 4.569 19.733 4.709 ;
      RECT 19.561 4.573 19.647 4.712 ;
      RECT 19.475 4.578 19.561 4.716 ;
      RECT 19.455 4.58 19.475 4.719 ;
      RECT 19.435 4.579 19.455 4.72 ;
      RECT 19.386 4.576 19.435 4.721 ;
      RECT 19.3 4.571 19.386 4.724 ;
      RECT 19.25 4.566 19.3 4.726 ;
      RECT 19.226 4.564 19.25 4.727 ;
      RECT 19.14 4.559 19.226 4.729 ;
      RECT 19.115 4.555 19.14 4.728 ;
      RECT 19.105 4.552 19.115 4.726 ;
      RECT 19.095 4.545 19.105 4.723 ;
      RECT 19.09 4.525 19.095 4.718 ;
      RECT 19.08 4.495 19.09 4.713 ;
      RECT 19.065 4.365 19.08 4.704 ;
      RECT 19.06 4.357 19.065 4.697 ;
      RECT 19.04 4.35 19.06 4.689 ;
      RECT 19.035 4.332 19.04 4.681 ;
      RECT 19.025 4.312 19.035 4.676 ;
      RECT 19.02 4.285 19.025 4.672 ;
      RECT 19.015 4.262 19.02 4.669 ;
      RECT 18.995 4.22 19.015 4.661 ;
      RECT 18.96 4.135 18.995 4.645 ;
      RECT 18.955 4.067 18.96 4.633 ;
      RECT 18.94 4.037 18.955 4.627 ;
      RECT 18.935 3.282 18.94 3.528 ;
      RECT 18.925 4.007 18.94 4.618 ;
      RECT 18.93 3.277 18.935 3.56 ;
      RECT 18.925 3.272 18.93 3.603 ;
      RECT 18.92 3.27 18.925 3.638 ;
      RECT 18.905 3.97 18.925 4.608 ;
      RECT 18.915 3.27 18.92 3.675 ;
      RECT 18.9 3.27 18.915 3.773 ;
      RECT 18.9 3.943 18.905 4.601 ;
      RECT 18.895 3.27 18.9 3.848 ;
      RECT 18.895 3.931 18.9 4.598 ;
      RECT 18.89 3.27 18.895 3.88 ;
      RECT 18.89 3.91 18.895 4.595 ;
      RECT 18.885 3.27 18.89 4.592 ;
      RECT 18.85 3.27 18.885 4.578 ;
      RECT 18.835 3.27 18.85 4.56 ;
      RECT 18.815 3.27 18.835 4.55 ;
      RECT 18.79 3.27 18.815 4.533 ;
      RECT 18.785 3.27 18.79 4.483 ;
      RECT 18.775 3.27 18.78 4.313 ;
      RECT 18.77 3.27 18.775 4.22 ;
      RECT 18.765 3.27 18.77 4.133 ;
      RECT 18.76 3.27 18.765 4.065 ;
      RECT 18.755 3.27 18.76 4.008 ;
      RECT 18.745 3.27 18.755 3.903 ;
      RECT 18.74 3.27 18.745 3.775 ;
      RECT 18.735 3.27 18.74 3.693 ;
      RECT 18.73 3.272 18.735 3.61 ;
      RECT 18.725 3.277 18.73 3.543 ;
      RECT 18.72 3.282 18.725 3.47 ;
      RECT 21.535 3.6 21.795 3.86 ;
      RECT 21.555 3.567 21.765 3.86 ;
      RECT 21.555 3.565 21.755 3.86 ;
      RECT 21.565 3.552 21.755 3.86 ;
      RECT 21.565 3.55 21.68 3.86 ;
      RECT 21.04 3.675 21.215 3.955 ;
      RECT 21.035 3.675 21.215 3.953 ;
      RECT 21.035 3.675 21.23 3.95 ;
      RECT 21.025 3.675 21.23 3.948 ;
      RECT 20.97 3.675 21.23 3.935 ;
      RECT 20.97 3.75 21.235 3.913 ;
      RECT 20.5 4.873 20.505 5.08 ;
      RECT 20.45 4.867 20.5 5.079 ;
      RECT 20.417 4.881 20.51 5.078 ;
      RECT 20.331 4.881 20.51 5.077 ;
      RECT 20.245 4.881 20.51 5.076 ;
      RECT 20.245 4.98 20.515 5.073 ;
      RECT 20.24 4.98 20.515 5.068 ;
      RECT 20.235 4.98 20.515 5.05 ;
      RECT 20.23 4.98 20.515 5.033 ;
      RECT 20.19 4.765 20.45 5.025 ;
      RECT 19.65 3.915 19.736 4.329 ;
      RECT 19.65 3.915 19.775 4.326 ;
      RECT 19.65 3.915 19.795 4.316 ;
      RECT 19.605 3.915 19.795 4.313 ;
      RECT 19.605 4.067 19.805 4.303 ;
      RECT 19.605 4.088 19.81 4.297 ;
      RECT 19.605 4.106 19.815 4.293 ;
      RECT 19.605 4.126 19.825 4.288 ;
      RECT 19.58 4.126 19.825 4.285 ;
      RECT 19.57 4.126 19.825 4.263 ;
      RECT 19.57 4.142 19.83 4.233 ;
      RECT 19.535 3.915 19.795 4.22 ;
      RECT 19.535 4.154 19.835 4.175 ;
      RECT 16.545 10.06 16.835 10.29 ;
      RECT 16.605 9.315 16.775 10.29 ;
      RECT 16.515 9.315 16.865 9.605 ;
      RECT 16.14 8.575 16.49 8.865 ;
      RECT 16 8.61 16.49 8.78 ;
      RECT 93.47 7.25 93.82 7.54 ;
      RECT 83.16 4.56 83.42 4.82 ;
      RECT 78.21 7.25 78.56 7.54 ;
      RECT 67.9 4.56 68.16 4.82 ;
      RECT 62.95 7.25 63.3 7.54 ;
      RECT 52.64 4.56 52.9 4.82 ;
      RECT 47.69 7.25 48.04 7.54 ;
      RECT 37.38 4.56 37.64 4.82 ;
      RECT 32.43 7.25 32.78 7.54 ;
      RECT 22.12 4.56 22.38 4.82 ;
    LAYER mcon ;
      RECT 93.56 7.31 93.73 7.48 ;
      RECT 93.555 8.61 93.725 8.78 ;
      RECT 93.555 10.09 93.725 10.26 ;
      RECT 93.185 8.24 93.355 8.41 ;
      RECT 93.18 4.055 93.35 4.225 ;
      RECT 92.565 2.205 92.735 2.375 ;
      RECT 92.565 3.685 92.735 3.855 ;
      RECT 92.565 8.61 92.735 8.78 ;
      RECT 92.565 10.09 92.735 10.26 ;
      RECT 92.195 4.055 92.365 4.225 ;
      RECT 92.195 8.24 92.365 8.41 ;
      RECT 91.205 3.315 91.375 3.485 ;
      RECT 91.205 8.98 91.375 9.15 ;
      RECT 90.775 2.205 90.945 2.375 ;
      RECT 90.775 2.945 90.945 3.115 ;
      RECT 90.775 9.35 90.945 9.52 ;
      RECT 90.775 10.09 90.945 10.26 ;
      RECT 90.405 3.685 90.575 3.855 ;
      RECT 90.405 8.61 90.575 8.78 ;
      RECT 87.575 3.575 87.745 3.745 ;
      RECT 87.18 4.32 87.35 4.49 ;
      RECT 87.07 3.595 87.24 3.765 ;
      RECT 86.25 3.285 86.42 3.455 ;
      RECT 85.935 4.325 86.105 4.495 ;
      RECT 85.89 3.815 86.06 3.985 ;
      RECT 85.57 8.98 85.74 9.15 ;
      RECT 85.465 4.025 85.635 4.195 ;
      RECT 85.275 3.245 85.445 3.415 ;
      RECT 85.225 4.855 85.395 5.025 ;
      RECT 85.14 9.35 85.31 9.52 ;
      RECT 85.14 10.09 85.31 10.26 ;
      RECT 84.89 4.295 85.06 4.465 ;
      RECT 84.795 3.455 84.965 3.625 ;
      RECT 83.995 4.68 84.165 4.85 ;
      RECT 83.935 3.88 84.105 4.05 ;
      RECT 83.495 3.55 83.665 3.72 ;
      RECT 83.23 4.6 83.4 4.77 ;
      RECT 82.985 3.84 83.155 4.01 ;
      RECT 82.89 4.87 83.06 5.04 ;
      RECT 82.615 3.565 82.785 3.735 ;
      RECT 82.085 3.765 82.255 3.935 ;
      RECT 81.36 3.31 81.53 3.48 ;
      RECT 81.36 4.89 81.53 5.06 ;
      RECT 81.05 3.855 81.22 4.025 ;
      RECT 80.64 4.08 80.81 4.25 ;
      RECT 79.93 4.38 80.1 4.55 ;
      RECT 79.785 3.29 79.955 3.46 ;
      RECT 78.3 7.31 78.47 7.48 ;
      RECT 78.295 8.61 78.465 8.78 ;
      RECT 78.295 10.09 78.465 10.26 ;
      RECT 77.925 8.24 78.095 8.41 ;
      RECT 77.92 4.055 78.09 4.225 ;
      RECT 77.305 2.205 77.475 2.375 ;
      RECT 77.305 3.685 77.475 3.855 ;
      RECT 77.305 8.61 77.475 8.78 ;
      RECT 77.305 10.09 77.475 10.26 ;
      RECT 76.935 4.055 77.105 4.225 ;
      RECT 76.935 8.24 77.105 8.41 ;
      RECT 75.945 3.315 76.115 3.485 ;
      RECT 75.945 8.98 76.115 9.15 ;
      RECT 75.515 2.205 75.685 2.375 ;
      RECT 75.515 2.945 75.685 3.115 ;
      RECT 75.515 9.35 75.685 9.52 ;
      RECT 75.515 10.09 75.685 10.26 ;
      RECT 75.145 3.685 75.315 3.855 ;
      RECT 75.145 8.61 75.315 8.78 ;
      RECT 72.315 3.575 72.485 3.745 ;
      RECT 71.92 4.32 72.09 4.49 ;
      RECT 71.81 3.595 71.98 3.765 ;
      RECT 70.99 3.285 71.16 3.455 ;
      RECT 70.675 4.325 70.845 4.495 ;
      RECT 70.63 3.815 70.8 3.985 ;
      RECT 70.31 8.98 70.48 9.15 ;
      RECT 70.205 4.025 70.375 4.195 ;
      RECT 70.015 3.245 70.185 3.415 ;
      RECT 69.965 4.855 70.135 5.025 ;
      RECT 69.88 9.35 70.05 9.52 ;
      RECT 69.88 10.09 70.05 10.26 ;
      RECT 69.63 4.295 69.8 4.465 ;
      RECT 69.535 3.455 69.705 3.625 ;
      RECT 68.735 4.68 68.905 4.85 ;
      RECT 68.675 3.88 68.845 4.05 ;
      RECT 68.235 3.55 68.405 3.72 ;
      RECT 67.97 4.6 68.14 4.77 ;
      RECT 67.725 3.84 67.895 4.01 ;
      RECT 67.63 4.87 67.8 5.04 ;
      RECT 67.355 3.565 67.525 3.735 ;
      RECT 66.825 3.765 66.995 3.935 ;
      RECT 66.1 3.31 66.27 3.48 ;
      RECT 66.1 4.89 66.27 5.06 ;
      RECT 65.79 3.855 65.96 4.025 ;
      RECT 65.38 4.08 65.55 4.25 ;
      RECT 64.67 4.38 64.84 4.55 ;
      RECT 64.525 3.29 64.695 3.46 ;
      RECT 63.04 7.31 63.21 7.48 ;
      RECT 63.035 8.61 63.205 8.78 ;
      RECT 63.035 10.09 63.205 10.26 ;
      RECT 62.665 8.24 62.835 8.41 ;
      RECT 62.66 4.055 62.83 4.225 ;
      RECT 62.045 2.205 62.215 2.375 ;
      RECT 62.045 3.685 62.215 3.855 ;
      RECT 62.045 8.61 62.215 8.78 ;
      RECT 62.045 10.09 62.215 10.26 ;
      RECT 61.675 4.055 61.845 4.225 ;
      RECT 61.675 8.24 61.845 8.41 ;
      RECT 60.685 3.315 60.855 3.485 ;
      RECT 60.685 8.98 60.855 9.15 ;
      RECT 60.255 2.205 60.425 2.375 ;
      RECT 60.255 2.945 60.425 3.115 ;
      RECT 60.255 9.35 60.425 9.52 ;
      RECT 60.255 10.09 60.425 10.26 ;
      RECT 59.885 3.685 60.055 3.855 ;
      RECT 59.885 8.61 60.055 8.78 ;
      RECT 57.055 3.575 57.225 3.745 ;
      RECT 56.66 4.32 56.83 4.49 ;
      RECT 56.55 3.595 56.72 3.765 ;
      RECT 55.73 3.285 55.9 3.455 ;
      RECT 55.415 4.325 55.585 4.495 ;
      RECT 55.37 3.815 55.54 3.985 ;
      RECT 55.05 8.98 55.22 9.15 ;
      RECT 54.945 4.025 55.115 4.195 ;
      RECT 54.755 3.245 54.925 3.415 ;
      RECT 54.705 4.855 54.875 5.025 ;
      RECT 54.62 9.35 54.79 9.52 ;
      RECT 54.62 10.09 54.79 10.26 ;
      RECT 54.37 4.295 54.54 4.465 ;
      RECT 54.275 3.455 54.445 3.625 ;
      RECT 53.475 4.68 53.645 4.85 ;
      RECT 53.415 3.88 53.585 4.05 ;
      RECT 52.975 3.55 53.145 3.72 ;
      RECT 52.71 4.6 52.88 4.77 ;
      RECT 52.465 3.84 52.635 4.01 ;
      RECT 52.37 4.87 52.54 5.04 ;
      RECT 52.095 3.565 52.265 3.735 ;
      RECT 51.565 3.765 51.735 3.935 ;
      RECT 50.84 3.31 51.01 3.48 ;
      RECT 50.84 4.89 51.01 5.06 ;
      RECT 50.53 3.855 50.7 4.025 ;
      RECT 50.12 4.08 50.29 4.25 ;
      RECT 49.41 4.38 49.58 4.55 ;
      RECT 49.265 3.29 49.435 3.46 ;
      RECT 47.78 7.31 47.95 7.48 ;
      RECT 47.775 8.61 47.945 8.78 ;
      RECT 47.775 10.09 47.945 10.26 ;
      RECT 47.405 8.24 47.575 8.41 ;
      RECT 47.4 4.055 47.57 4.225 ;
      RECT 46.785 2.205 46.955 2.375 ;
      RECT 46.785 3.685 46.955 3.855 ;
      RECT 46.785 8.61 46.955 8.78 ;
      RECT 46.785 10.09 46.955 10.26 ;
      RECT 46.415 4.055 46.585 4.225 ;
      RECT 46.415 8.24 46.585 8.41 ;
      RECT 45.425 3.315 45.595 3.485 ;
      RECT 45.425 8.98 45.595 9.15 ;
      RECT 44.995 2.205 45.165 2.375 ;
      RECT 44.995 2.945 45.165 3.115 ;
      RECT 44.995 9.35 45.165 9.52 ;
      RECT 44.995 10.09 45.165 10.26 ;
      RECT 44.625 3.685 44.795 3.855 ;
      RECT 44.625 8.61 44.795 8.78 ;
      RECT 41.795 3.575 41.965 3.745 ;
      RECT 41.4 4.32 41.57 4.49 ;
      RECT 41.29 3.595 41.46 3.765 ;
      RECT 40.47 3.285 40.64 3.455 ;
      RECT 40.155 4.325 40.325 4.495 ;
      RECT 40.11 3.815 40.28 3.985 ;
      RECT 39.79 8.98 39.96 9.15 ;
      RECT 39.685 4.025 39.855 4.195 ;
      RECT 39.495 3.245 39.665 3.415 ;
      RECT 39.445 4.855 39.615 5.025 ;
      RECT 39.36 9.35 39.53 9.52 ;
      RECT 39.36 10.09 39.53 10.26 ;
      RECT 39.11 4.295 39.28 4.465 ;
      RECT 39.015 3.455 39.185 3.625 ;
      RECT 38.215 4.68 38.385 4.85 ;
      RECT 38.155 3.88 38.325 4.05 ;
      RECT 37.715 3.55 37.885 3.72 ;
      RECT 37.45 4.6 37.62 4.77 ;
      RECT 37.205 3.84 37.375 4.01 ;
      RECT 37.11 4.87 37.28 5.04 ;
      RECT 36.835 3.565 37.005 3.735 ;
      RECT 36.305 3.765 36.475 3.935 ;
      RECT 35.58 3.31 35.75 3.48 ;
      RECT 35.58 4.89 35.75 5.06 ;
      RECT 35.27 3.855 35.44 4.025 ;
      RECT 34.86 4.08 35.03 4.25 ;
      RECT 34.15 4.38 34.32 4.55 ;
      RECT 34.005 3.29 34.175 3.46 ;
      RECT 32.52 7.31 32.69 7.48 ;
      RECT 32.515 8.61 32.685 8.78 ;
      RECT 32.515 10.09 32.685 10.26 ;
      RECT 32.145 8.24 32.315 8.41 ;
      RECT 32.14 4.055 32.31 4.225 ;
      RECT 31.525 2.205 31.695 2.375 ;
      RECT 31.525 3.685 31.695 3.855 ;
      RECT 31.525 8.61 31.695 8.78 ;
      RECT 31.525 10.09 31.695 10.26 ;
      RECT 31.155 4.055 31.325 4.225 ;
      RECT 31.155 8.24 31.325 8.41 ;
      RECT 30.165 3.315 30.335 3.485 ;
      RECT 30.165 8.98 30.335 9.15 ;
      RECT 29.735 2.205 29.905 2.375 ;
      RECT 29.735 2.945 29.905 3.115 ;
      RECT 29.735 9.35 29.905 9.52 ;
      RECT 29.735 10.09 29.905 10.26 ;
      RECT 29.365 3.685 29.535 3.855 ;
      RECT 29.365 8.61 29.535 8.78 ;
      RECT 26.535 3.575 26.705 3.745 ;
      RECT 26.14 4.32 26.31 4.49 ;
      RECT 26.03 3.595 26.2 3.765 ;
      RECT 25.21 3.285 25.38 3.455 ;
      RECT 24.895 4.325 25.065 4.495 ;
      RECT 24.85 3.815 25.02 3.985 ;
      RECT 24.53 8.98 24.7 9.15 ;
      RECT 24.425 4.025 24.595 4.195 ;
      RECT 24.235 3.245 24.405 3.415 ;
      RECT 24.185 4.855 24.355 5.025 ;
      RECT 24.1 9.35 24.27 9.52 ;
      RECT 24.1 10.09 24.27 10.26 ;
      RECT 23.85 4.295 24.02 4.465 ;
      RECT 23.755 3.455 23.925 3.625 ;
      RECT 22.955 4.68 23.125 4.85 ;
      RECT 22.895 3.88 23.065 4.05 ;
      RECT 22.455 3.55 22.625 3.72 ;
      RECT 22.19 4.6 22.36 4.77 ;
      RECT 21.945 3.84 22.115 4.01 ;
      RECT 21.85 4.87 22.02 5.04 ;
      RECT 21.575 3.565 21.745 3.735 ;
      RECT 21.045 3.765 21.215 3.935 ;
      RECT 20.32 3.31 20.49 3.48 ;
      RECT 20.32 4.89 20.49 5.06 ;
      RECT 20.01 3.855 20.18 4.025 ;
      RECT 19.6 4.08 19.77 4.25 ;
      RECT 18.89 4.38 19.06 4.55 ;
      RECT 18.745 3.29 18.915 3.46 ;
      RECT 16.605 9.35 16.775 9.52 ;
      RECT 16.605 10.09 16.775 10.26 ;
      RECT 16.235 8.61 16.405 8.78 ;
    LAYER li1 ;
      RECT 93.555 7.31 93.725 8.78 ;
      RECT 93.555 7.31 93.73 8.57 ;
      RECT 93.185 9.26 93.655 9.43 ;
      RECT 93.185 8.24 93.355 9.43 ;
      RECT 93.18 3.035 93.35 4.225 ;
      RECT 93.18 3.035 93.65 3.205 ;
      RECT 92.565 3.895 92.74 5.155 ;
      RECT 92.565 3.685 92.735 5.155 ;
      RECT 92.565 7.31 92.735 8.78 ;
      RECT 92.565 7.31 92.74 8.57 ;
      RECT 92.195 3.035 92.365 4.225 ;
      RECT 92.195 3.035 92.665 3.205 ;
      RECT 92.195 9.26 92.665 9.43 ;
      RECT 92.195 8.24 92.365 9.43 ;
      RECT 91.205 4.015 91.38 5.155 ;
      RECT 91.205 1.865 91.375 5.155 ;
      RECT 91.205 1.865 91.38 2.415 ;
      RECT 91.205 10.05 91.38 10.6 ;
      RECT 91.205 7.31 91.375 10.6 ;
      RECT 91.205 7.31 91.38 8.45 ;
      RECT 90.775 3.895 90.95 5.155 ;
      RECT 90.775 2.945 90.945 5.155 ;
      RECT 90.775 7.31 90.945 9.52 ;
      RECT 90.775 7.31 90.95 8.57 ;
      RECT 90.345 3.925 90.515 5.155 ;
      RECT 90.405 2.145 90.575 4.095 ;
      RECT 90.345 1.865 90.515 2.315 ;
      RECT 90.345 10.15 90.515 10.6 ;
      RECT 90.405 8.37 90.575 10.32 ;
      RECT 90.345 7.31 90.515 8.54 ;
      RECT 89.82 3.895 89.995 5.155 ;
      RECT 89.82 1.865 89.99 5.155 ;
      RECT 89.82 3.365 90.23 3.695 ;
      RECT 89.82 2.525 90.23 2.855 ;
      RECT 89.82 1.865 89.995 2.355 ;
      RECT 89.82 10.11 89.995 10.6 ;
      RECT 89.82 7.31 89.99 10.6 ;
      RECT 89.82 9.61 90.23 9.94 ;
      RECT 89.82 8.77 90.23 9.1 ;
      RECT 89.82 7.31 89.995 8.57 ;
      RECT 87.75 4.421 87.755 4.593 ;
      RECT 87.745 4.414 87.75 4.683 ;
      RECT 87.74 4.408 87.745 4.702 ;
      RECT 87.72 4.402 87.74 4.712 ;
      RECT 87.705 4.397 87.72 4.72 ;
      RECT 87.668 4.391 87.705 4.718 ;
      RECT 87.582 4.377 87.668 4.714 ;
      RECT 87.496 4.359 87.582 4.709 ;
      RECT 87.41 4.34 87.496 4.703 ;
      RECT 87.38 4.328 87.41 4.699 ;
      RECT 87.36 4.322 87.38 4.698 ;
      RECT 87.295 4.32 87.36 4.696 ;
      RECT 87.28 4.32 87.295 4.688 ;
      RECT 87.265 4.32 87.28 4.675 ;
      RECT 87.26 4.32 87.265 4.665 ;
      RECT 87.245 4.32 87.26 4.643 ;
      RECT 87.23 4.32 87.245 4.61 ;
      RECT 87.225 4.32 87.23 4.588 ;
      RECT 87.215 4.32 87.225 4.57 ;
      RECT 87.2 4.32 87.215 4.548 ;
      RECT 87.18 4.32 87.2 4.51 ;
      RECT 87.53 3.605 87.565 4.044 ;
      RECT 87.53 3.605 87.57 4.043 ;
      RECT 87.475 3.665 87.57 4.042 ;
      RECT 87.34 3.837 87.57 4.041 ;
      RECT 87.45 3.715 87.57 4.041 ;
      RECT 87.34 3.837 87.595 4.031 ;
      RECT 87.395 3.782 87.675 3.948 ;
      RECT 87.57 3.576 87.575 4.039 ;
      RECT 87.425 3.752 87.715 3.825 ;
      RECT 87.44 3.735 87.57 4.041 ;
      RECT 87.575 3.575 87.745 3.763 ;
      RECT 87.565 3.578 87.745 3.763 ;
      RECT 87.07 3.455 87.24 3.765 ;
      RECT 87.07 3.455 87.245 3.738 ;
      RECT 87.07 3.455 87.25 3.715 ;
      RECT 87.07 3.455 87.26 3.665 ;
      RECT 87.065 3.56 87.26 3.635 ;
      RECT 87.1 3.13 87.27 3.608 ;
      RECT 87.1 3.13 87.285 3.529 ;
      RECT 87.09 3.34 87.285 3.529 ;
      RECT 87.1 3.14 87.295 3.444 ;
      RECT 87.03 3.882 87.035 4.085 ;
      RECT 87.02 3.87 87.03 4.195 ;
      RECT 86.995 3.87 87.02 4.235 ;
      RECT 86.915 3.87 86.995 4.32 ;
      RECT 86.905 3.87 86.915 4.39 ;
      RECT 86.88 3.87 86.905 4.413 ;
      RECT 86.86 3.87 86.88 4.448 ;
      RECT 86.815 3.88 86.86 4.491 ;
      RECT 86.805 3.892 86.815 4.528 ;
      RECT 86.785 3.906 86.805 4.548 ;
      RECT 86.775 3.924 86.785 4.564 ;
      RECT 86.76 3.95 86.775 4.574 ;
      RECT 86.745 3.991 86.76 4.588 ;
      RECT 86.735 4.026 86.745 4.598 ;
      RECT 86.73 4.042 86.735 4.603 ;
      RECT 86.72 4.057 86.73 4.608 ;
      RECT 86.7 4.1 86.72 4.618 ;
      RECT 86.68 4.137 86.7 4.631 ;
      RECT 86.645 4.16 86.68 4.649 ;
      RECT 86.635 4.174 86.645 4.665 ;
      RECT 86.615 4.184 86.635 4.675 ;
      RECT 86.61 4.193 86.615 4.683 ;
      RECT 86.6 4.2 86.61 4.69 ;
      RECT 86.59 4.207 86.6 4.698 ;
      RECT 86.575 4.217 86.59 4.706 ;
      RECT 86.565 4.231 86.575 4.716 ;
      RECT 86.555 4.243 86.565 4.728 ;
      RECT 86.54 4.265 86.555 4.741 ;
      RECT 86.53 4.287 86.54 4.752 ;
      RECT 86.52 4.307 86.53 4.761 ;
      RECT 86.515 4.322 86.52 4.768 ;
      RECT 86.485 4.355 86.515 4.782 ;
      RECT 86.475 4.39 86.485 4.797 ;
      RECT 86.47 4.397 86.475 4.803 ;
      RECT 86.45 4.412 86.47 4.81 ;
      RECT 86.445 4.427 86.45 4.818 ;
      RECT 86.44 4.436 86.445 4.823 ;
      RECT 86.425 4.442 86.44 4.83 ;
      RECT 86.42 4.448 86.425 4.838 ;
      RECT 86.415 4.452 86.42 4.845 ;
      RECT 86.41 4.456 86.415 4.855 ;
      RECT 86.4 4.461 86.41 4.865 ;
      RECT 86.38 4.472 86.4 4.893 ;
      RECT 86.365 4.484 86.38 4.92 ;
      RECT 86.345 4.497 86.365 4.945 ;
      RECT 86.325 4.512 86.345 4.969 ;
      RECT 86.31 4.527 86.325 4.984 ;
      RECT 86.305 4.538 86.31 4.993 ;
      RECT 86.24 4.583 86.305 5.003 ;
      RECT 86.205 4.642 86.24 5.016 ;
      RECT 86.2 4.665 86.205 5.022 ;
      RECT 86.195 4.672 86.2 5.024 ;
      RECT 86.18 4.682 86.195 5.027 ;
      RECT 86.15 4.707 86.18 5.031 ;
      RECT 86.145 4.725 86.15 5.035 ;
      RECT 86.14 4.732 86.145 5.036 ;
      RECT 86.12 4.74 86.14 5.04 ;
      RECT 86.11 4.747 86.12 5.044 ;
      RECT 86.066 4.758 86.11 5.051 ;
      RECT 85.98 4.786 86.066 5.067 ;
      RECT 85.92 4.81 85.98 5.085 ;
      RECT 85.875 4.82 85.92 5.099 ;
      RECT 85.816 4.828 85.875 5.113 ;
      RECT 85.73 4.835 85.816 5.132 ;
      RECT 85.705 4.84 85.73 5.147 ;
      RECT 85.625 4.843 85.705 5.15 ;
      RECT 85.545 4.847 85.625 5.137 ;
      RECT 85.536 4.85 85.545 5.122 ;
      RECT 85.45 4.85 85.536 5.107 ;
      RECT 85.39 4.852 85.45 5.084 ;
      RECT 85.386 4.855 85.39 5.074 ;
      RECT 85.3 4.855 85.386 5.059 ;
      RECT 85.225 4.855 85.3 5.035 ;
      RECT 86.54 3.864 86.55 4.04 ;
      RECT 86.495 3.831 86.54 4.04 ;
      RECT 86.45 3.782 86.495 4.04 ;
      RECT 86.42 3.752 86.45 4.041 ;
      RECT 86.415 3.735 86.42 4.042 ;
      RECT 86.39 3.715 86.415 4.043 ;
      RECT 86.375 3.69 86.39 4.044 ;
      RECT 86.37 3.677 86.375 4.045 ;
      RECT 86.365 3.671 86.37 4.043 ;
      RECT 86.36 3.663 86.365 4.037 ;
      RECT 86.335 3.655 86.36 4.017 ;
      RECT 86.315 3.644 86.335 3.988 ;
      RECT 86.285 3.629 86.315 3.959 ;
      RECT 86.265 3.615 86.285 3.931 ;
      RECT 86.255 3.609 86.265 3.91 ;
      RECT 86.25 3.606 86.255 3.893 ;
      RECT 86.245 3.603 86.25 3.878 ;
      RECT 86.23 3.598 86.245 3.843 ;
      RECT 86.225 3.594 86.23 3.81 ;
      RECT 86.205 3.589 86.225 3.786 ;
      RECT 86.175 3.581 86.205 3.751 ;
      RECT 86.16 3.575 86.175 3.728 ;
      RECT 86.12 3.568 86.16 3.713 ;
      RECT 86.095 3.56 86.12 3.693 ;
      RECT 86.075 3.555 86.095 3.683 ;
      RECT 86.04 3.549 86.075 3.678 ;
      RECT 85.995 3.54 86.04 3.677 ;
      RECT 85.965 3.536 85.995 3.679 ;
      RECT 85.88 3.544 85.965 3.683 ;
      RECT 85.81 3.555 85.88 3.705 ;
      RECT 85.797 3.561 85.81 3.728 ;
      RECT 85.711 3.568 85.797 3.75 ;
      RECT 85.625 3.58 85.711 3.787 ;
      RECT 85.625 3.957 85.635 4.195 ;
      RECT 85.62 3.586 85.625 3.81 ;
      RECT 85.615 3.842 85.625 4.195 ;
      RECT 85.615 3.587 85.62 3.815 ;
      RECT 85.61 3.588 85.615 4.195 ;
      RECT 85.586 3.59 85.61 4.196 ;
      RECT 85.5 3.598 85.586 4.198 ;
      RECT 85.48 3.612 85.5 4.201 ;
      RECT 85.475 3.64 85.48 4.202 ;
      RECT 85.47 3.652 85.475 4.203 ;
      RECT 85.465 3.667 85.47 4.204 ;
      RECT 85.455 3.697 85.465 4.205 ;
      RECT 85.45 3.735 85.455 4.203 ;
      RECT 85.445 3.755 85.45 4.198 ;
      RECT 85.43 3.79 85.445 4.183 ;
      RECT 85.42 3.842 85.43 4.163 ;
      RECT 85.415 3.872 85.42 4.151 ;
      RECT 85.4 3.885 85.415 4.134 ;
      RECT 85.375 3.889 85.4 4.101 ;
      RECT 85.36 3.887 85.375 4.078 ;
      RECT 85.345 3.886 85.36 4.075 ;
      RECT 85.285 3.884 85.345 4.073 ;
      RECT 85.275 3.882 85.285 4.068 ;
      RECT 85.235 3.881 85.275 4.065 ;
      RECT 85.165 3.878 85.235 4.063 ;
      RECT 85.11 3.876 85.165 4.058 ;
      RECT 85.04 3.87 85.11 4.053 ;
      RECT 85.031 3.87 85.04 4.05 ;
      RECT 84.945 3.87 85.031 4.045 ;
      RECT 84.94 3.87 84.945 4.04 ;
      RECT 86.245 3.105 86.42 3.455 ;
      RECT 86.245 3.12 86.43 3.453 ;
      RECT 86.22 3.07 86.365 3.45 ;
      RECT 86.2 3.071 86.365 3.443 ;
      RECT 86.19 3.072 86.375 3.438 ;
      RECT 86.16 3.073 86.375 3.425 ;
      RECT 86.11 3.074 86.375 3.401 ;
      RECT 86.105 3.076 86.375 3.386 ;
      RECT 86.105 3.142 86.435 3.38 ;
      RECT 86.085 3.083 86.39 3.36 ;
      RECT 86.075 3.092 86.4 3.215 ;
      RECT 86.085 3.087 86.4 3.36 ;
      RECT 86.105 3.077 86.39 3.386 ;
      RECT 85.69 4.402 85.86 4.69 ;
      RECT 85.685 4.42 85.87 4.685 ;
      RECT 85.65 4.428 85.935 4.605 ;
      RECT 85.65 4.428 86.021 4.595 ;
      RECT 85.65 4.428 86.075 4.541 ;
      RECT 85.935 4.325 86.105 4.509 ;
      RECT 85.65 4.48 86.11 4.497 ;
      RECT 85.635 4.45 86.105 4.493 ;
      RECT 85.895 4.332 85.935 4.644 ;
      RECT 85.775 4.369 86.105 4.509 ;
      RECT 85.87 4.344 85.895 4.67 ;
      RECT 85.86 4.351 86.105 4.509 ;
      RECT 85.991 3.815 86.06 4.074 ;
      RECT 85.991 3.87 86.065 4.073 ;
      RECT 85.905 3.87 86.065 4.072 ;
      RECT 85.9 3.87 86.07 4.065 ;
      RECT 85.89 3.815 86.06 4.06 ;
      RECT 85.57 10.05 85.745 10.6 ;
      RECT 85.57 7.31 85.74 10.6 ;
      RECT 85.57 7.31 85.745 8.45 ;
      RECT 85.27 3.114 85.445 3.415 ;
      RECT 85.255 3.102 85.27 3.4 ;
      RECT 85.225 3.101 85.255 3.353 ;
      RECT 85.225 3.119 85.45 3.348 ;
      RECT 85.21 3.103 85.27 3.313 ;
      RECT 85.205 3.125 85.46 3.213 ;
      RECT 85.205 3.108 85.356 3.213 ;
      RECT 85.205 3.11 85.36 3.213 ;
      RECT 85.21 3.106 85.356 3.313 ;
      RECT 85.315 4.342 85.32 4.69 ;
      RECT 85.305 4.332 85.315 4.696 ;
      RECT 85.27 4.322 85.305 4.698 ;
      RECT 85.232 4.317 85.27 4.702 ;
      RECT 85.146 4.31 85.232 4.709 ;
      RECT 85.06 4.3 85.146 4.719 ;
      RECT 85.015 4.295 85.06 4.727 ;
      RECT 85.011 4.295 85.015 4.731 ;
      RECT 84.925 4.295 85.011 4.738 ;
      RECT 84.91 4.295 84.925 4.738 ;
      RECT 84.9 4.293 84.91 4.71 ;
      RECT 84.89 4.289 84.9 4.653 ;
      RECT 84.87 4.283 84.89 4.585 ;
      RECT 84.865 4.279 84.87 4.533 ;
      RECT 84.855 4.278 84.865 4.5 ;
      RECT 84.805 4.276 84.855 4.485 ;
      RECT 84.78 4.274 84.805 4.48 ;
      RECT 84.737 4.272 84.78 4.476 ;
      RECT 84.651 4.268 84.737 4.464 ;
      RECT 84.565 4.263 84.651 4.448 ;
      RECT 84.535 4.26 84.565 4.435 ;
      RECT 84.51 4.259 84.535 4.423 ;
      RECT 84.505 4.259 84.51 4.413 ;
      RECT 84.465 4.258 84.505 4.405 ;
      RECT 84.45 4.257 84.465 4.398 ;
      RECT 84.4 4.256 84.45 4.39 ;
      RECT 84.398 4.255 84.4 4.385 ;
      RECT 84.312 4.253 84.398 4.385 ;
      RECT 84.226 4.248 84.312 4.385 ;
      RECT 84.14 4.244 84.226 4.385 ;
      RECT 84.091 4.24 84.14 4.383 ;
      RECT 84.005 4.237 84.091 4.378 ;
      RECT 83.982 4.234 84.005 4.374 ;
      RECT 83.896 4.231 83.982 4.369 ;
      RECT 83.81 4.227 83.896 4.36 ;
      RECT 83.785 4.22 83.81 4.355 ;
      RECT 83.725 4.185 83.785 4.352 ;
      RECT 83.705 4.11 83.725 4.349 ;
      RECT 83.7 4.052 83.705 4.348 ;
      RECT 83.675 3.992 83.7 4.347 ;
      RECT 83.6 3.87 83.675 4.343 ;
      RECT 83.59 3.87 83.6 4.335 ;
      RECT 83.575 3.87 83.59 4.325 ;
      RECT 83.56 3.87 83.575 4.295 ;
      RECT 83.545 3.87 83.56 4.24 ;
      RECT 83.53 3.87 83.545 4.178 ;
      RECT 83.505 3.87 83.53 4.103 ;
      RECT 83.5 3.87 83.505 4.053 ;
      RECT 85.14 7.31 85.31 9.52 ;
      RECT 85.14 7.31 85.315 8.57 ;
      RECT 84.845 3.415 84.865 3.724 ;
      RECT 84.831 3.417 84.88 3.721 ;
      RECT 84.831 3.422 84.9 3.712 ;
      RECT 84.745 3.42 84.88 3.706 ;
      RECT 84.745 3.428 84.935 3.689 ;
      RECT 84.71 3.43 84.935 3.688 ;
      RECT 84.68 3.438 84.935 3.679 ;
      RECT 84.67 3.443 84.955 3.665 ;
      RECT 84.71 3.433 84.955 3.665 ;
      RECT 84.71 3.436 84.965 3.653 ;
      RECT 84.68 3.438 84.975 3.64 ;
      RECT 84.68 3.442 84.985 3.583 ;
      RECT 84.67 3.447 84.99 3.498 ;
      RECT 84.831 3.415 84.865 3.721 ;
      RECT 84.27 3.518 84.275 3.73 ;
      RECT 84.145 3.515 84.16 3.73 ;
      RECT 83.61 3.545 83.68 3.73 ;
      RECT 83.495 3.545 83.53 3.725 ;
      RECT 84.616 3.847 84.635 4.041 ;
      RECT 84.53 3.802 84.616 4.042 ;
      RECT 84.52 3.755 84.53 4.044 ;
      RECT 84.515 3.735 84.52 4.045 ;
      RECT 84.495 3.7 84.515 4.046 ;
      RECT 84.48 3.65 84.495 4.047 ;
      RECT 84.46 3.587 84.48 4.048 ;
      RECT 84.45 3.55 84.46 4.049 ;
      RECT 84.435 3.539 84.45 4.05 ;
      RECT 84.43 3.531 84.435 4.048 ;
      RECT 84.42 3.53 84.43 4.04 ;
      RECT 84.39 3.527 84.42 4.019 ;
      RECT 84.315 3.522 84.39 3.964 ;
      RECT 84.3 3.518 84.315 3.91 ;
      RECT 84.29 3.518 84.3 3.805 ;
      RECT 84.275 3.518 84.29 3.738 ;
      RECT 84.26 3.518 84.27 3.728 ;
      RECT 84.205 3.517 84.26 3.725 ;
      RECT 84.16 3.515 84.205 3.728 ;
      RECT 84.132 3.515 84.145 3.731 ;
      RECT 84.046 3.519 84.132 3.733 ;
      RECT 83.96 3.525 84.046 3.738 ;
      RECT 83.94 3.529 83.96 3.74 ;
      RECT 83.938 3.53 83.94 3.739 ;
      RECT 83.852 3.532 83.938 3.738 ;
      RECT 83.766 3.537 83.852 3.735 ;
      RECT 83.68 3.542 83.766 3.732 ;
      RECT 83.53 3.545 83.61 3.728 ;
      RECT 84.185 10.11 84.36 10.6 ;
      RECT 84.185 7.31 84.355 10.6 ;
      RECT 84.185 9.61 84.595 9.94 ;
      RECT 84.185 8.77 84.595 9.1 ;
      RECT 84.185 7.31 84.36 8.57 ;
      RECT 84.306 4.52 84.355 4.854 ;
      RECT 84.306 4.52 84.36 4.853 ;
      RECT 84.22 4.52 84.36 4.852 ;
      RECT 83.995 4.628 84.365 4.85 ;
      RECT 84.22 4.52 84.39 4.843 ;
      RECT 84.19 4.532 84.395 4.834 ;
      RECT 84.175 4.55 84.4 4.831 ;
      RECT 83.99 4.634 84.4 4.758 ;
      RECT 83.985 4.641 84.4 4.718 ;
      RECT 84 4.607 84.4 4.831 ;
      RECT 84.161 4.553 84.365 4.85 ;
      RECT 84.075 4.573 84.4 4.831 ;
      RECT 84.175 4.547 84.395 4.834 ;
      RECT 83.945 3.871 84.135 4.065 ;
      RECT 83.94 3.873 84.135 4.064 ;
      RECT 83.935 3.877 84.15 4.061 ;
      RECT 83.95 3.87 84.15 4.061 ;
      RECT 83.935 3.98 84.155 4.056 ;
      RECT 83.23 4.48 83.321 4.778 ;
      RECT 83.225 4.482 83.4 4.773 ;
      RECT 83.23 4.48 83.4 4.773 ;
      RECT 83.225 4.486 83.42 4.771 ;
      RECT 83.225 4.541 83.46 4.77 ;
      RECT 83.225 4.576 83.475 4.764 ;
      RECT 83.225 4.61 83.485 4.754 ;
      RECT 83.215 4.49 83.42 4.605 ;
      RECT 83.215 4.51 83.435 4.605 ;
      RECT 83.215 4.493 83.425 4.605 ;
      RECT 83.44 3.261 83.445 3.323 ;
      RECT 83.435 3.183 83.44 3.346 ;
      RECT 83.43 3.14 83.435 3.357 ;
      RECT 83.425 3.13 83.43 3.369 ;
      RECT 83.42 3.13 83.425 3.378 ;
      RECT 83.395 3.13 83.42 3.41 ;
      RECT 83.39 3.13 83.395 3.443 ;
      RECT 83.375 3.13 83.39 3.468 ;
      RECT 83.365 3.13 83.375 3.495 ;
      RECT 83.36 3.13 83.365 3.508 ;
      RECT 83.355 3.13 83.36 3.523 ;
      RECT 83.345 3.13 83.355 3.538 ;
      RECT 83.34 3.13 83.345 3.558 ;
      RECT 83.315 3.13 83.34 3.593 ;
      RECT 83.27 3.13 83.315 3.638 ;
      RECT 83.26 3.13 83.27 3.651 ;
      RECT 83.175 3.215 83.26 3.658 ;
      RECT 83.14 3.337 83.175 3.667 ;
      RECT 83.135 3.377 83.14 3.671 ;
      RECT 83.115 3.4 83.135 3.673 ;
      RECT 83.11 3.43 83.115 3.676 ;
      RECT 83.1 3.442 83.11 3.677 ;
      RECT 83.055 3.465 83.1 3.682 ;
      RECT 83.015 3.495 83.055 3.69 ;
      RECT 82.98 3.507 83.015 3.696 ;
      RECT 82.975 3.512 82.98 3.7 ;
      RECT 82.905 3.522 82.975 3.707 ;
      RECT 82.865 3.532 82.905 3.717 ;
      RECT 82.845 3.537 82.865 3.723 ;
      RECT 82.835 3.541 82.845 3.728 ;
      RECT 82.83 3.544 82.835 3.731 ;
      RECT 82.82 3.545 82.83 3.732 ;
      RECT 82.795 3.547 82.82 3.736 ;
      RECT 82.785 3.552 82.795 3.739 ;
      RECT 82.74 3.56 82.785 3.74 ;
      RECT 82.615 3.565 82.74 3.74 ;
      RECT 83.17 3.862 83.19 4.044 ;
      RECT 83.121 3.847 83.17 4.043 ;
      RECT 83.035 3.862 83.19 4.041 ;
      RECT 83.02 3.862 83.19 4.04 ;
      RECT 82.985 3.84 83.155 4.025 ;
      RECT 83.055 4.86 83.07 5.069 ;
      RECT 83.055 4.868 83.075 5.068 ;
      RECT 83 4.868 83.075 5.067 ;
      RECT 82.98 4.872 83.08 5.065 ;
      RECT 82.96 4.822 83 5.064 ;
      RECT 82.905 4.88 83.085 5.062 ;
      RECT 82.87 4.837 83 5.06 ;
      RECT 82.866 4.84 83.055 5.059 ;
      RECT 82.78 4.848 83.055 5.057 ;
      RECT 82.78 4.892 83.09 5.05 ;
      RECT 82.77 4.985 83.09 5.048 ;
      RECT 82.78 4.904 83.095 5.033 ;
      RECT 82.78 4.925 83.11 5.003 ;
      RECT 82.78 4.952 83.115 4.973 ;
      RECT 82.905 4.83 83 5.062 ;
      RECT 82.535 3.875 82.54 4.413 ;
      RECT 82.34 4.205 82.345 4.4 ;
      RECT 80.64 3.87 80.655 4.25 ;
      RECT 82.705 3.87 82.71 4.04 ;
      RECT 82.7 3.87 82.705 4.05 ;
      RECT 82.695 3.87 82.7 4.063 ;
      RECT 82.67 3.87 82.695 4.105 ;
      RECT 82.645 3.87 82.67 4.178 ;
      RECT 82.63 3.87 82.645 4.23 ;
      RECT 82.625 3.87 82.63 4.26 ;
      RECT 82.6 3.87 82.625 4.3 ;
      RECT 82.585 3.87 82.6 4.355 ;
      RECT 82.58 3.87 82.585 4.388 ;
      RECT 82.555 3.87 82.58 4.408 ;
      RECT 82.54 3.87 82.555 4.414 ;
      RECT 82.47 3.905 82.535 4.41 ;
      RECT 82.42 3.96 82.47 4.405 ;
      RECT 82.41 3.992 82.42 4.403 ;
      RECT 82.405 4.017 82.41 4.403 ;
      RECT 82.385 4.09 82.405 4.403 ;
      RECT 82.375 4.17 82.385 4.402 ;
      RECT 82.36 4.2 82.375 4.402 ;
      RECT 82.345 4.205 82.36 4.401 ;
      RECT 82.285 4.207 82.34 4.398 ;
      RECT 82.255 4.212 82.285 4.394 ;
      RECT 82.253 4.215 82.255 4.393 ;
      RECT 82.167 4.217 82.253 4.39 ;
      RECT 82.081 4.223 82.167 4.384 ;
      RECT 81.995 4.228 82.081 4.378 ;
      RECT 81.922 4.233 81.995 4.379 ;
      RECT 81.836 4.239 81.922 4.387 ;
      RECT 81.75 4.245 81.836 4.396 ;
      RECT 81.73 4.249 81.75 4.401 ;
      RECT 81.683 4.251 81.73 4.404 ;
      RECT 81.597 4.256 81.683 4.41 ;
      RECT 81.511 4.261 81.597 4.419 ;
      RECT 81.425 4.267 81.511 4.427 ;
      RECT 81.34 4.265 81.425 4.436 ;
      RECT 81.336 4.26 81.34 4.44 ;
      RECT 81.25 4.255 81.336 4.432 ;
      RECT 81.186 4.246 81.25 4.42 ;
      RECT 81.1 4.237 81.186 4.407 ;
      RECT 81.076 4.23 81.1 4.398 ;
      RECT 80.99 4.224 81.076 4.385 ;
      RECT 80.95 4.217 80.99 4.371 ;
      RECT 80.945 4.207 80.95 4.367 ;
      RECT 80.935 4.195 80.945 4.366 ;
      RECT 80.915 4.165 80.935 4.363 ;
      RECT 80.86 4.085 80.915 4.357 ;
      RECT 80.84 4.004 80.86 4.352 ;
      RECT 80.82 3.962 80.84 4.348 ;
      RECT 80.795 3.915 80.82 4.342 ;
      RECT 80.79 3.89 80.795 4.339 ;
      RECT 80.755 3.87 80.79 4.334 ;
      RECT 80.746 3.87 80.755 4.327 ;
      RECT 80.66 3.87 80.746 4.297 ;
      RECT 80.655 3.87 80.66 4.26 ;
      RECT 80.62 3.87 80.64 4.182 ;
      RECT 80.615 3.912 80.62 4.147 ;
      RECT 80.61 3.987 80.615 4.103 ;
      RECT 82.06 3.792 82.235 4.04 ;
      RECT 82.06 3.792 82.24 4.038 ;
      RECT 82.055 3.824 82.24 3.998 ;
      RECT 82.085 3.765 82.255 3.985 ;
      RECT 82.05 3.842 82.255 3.918 ;
      RECT 81.36 3.305 81.53 3.48 ;
      RECT 81.36 3.305 81.702 3.472 ;
      RECT 81.36 3.305 81.785 3.466 ;
      RECT 81.36 3.305 81.82 3.462 ;
      RECT 81.36 3.305 81.84 3.461 ;
      RECT 81.36 3.305 81.926 3.457 ;
      RECT 81.82 3.13 81.99 3.452 ;
      RECT 81.395 3.237 82.02 3.45 ;
      RECT 81.385 3.292 82.025 3.448 ;
      RECT 81.36 3.328 82.035 3.443 ;
      RECT 81.36 3.355 82.04 3.373 ;
      RECT 81.425 3.18 82 3.45 ;
      RECT 81.616 3.165 82 3.45 ;
      RECT 81.45 3.168 82 3.45 ;
      RECT 81.53 3.166 81.616 3.477 ;
      RECT 81.616 3.163 81.995 3.45 ;
      RECT 81.8 3.14 81.995 3.45 ;
      RECT 81.702 3.161 81.995 3.45 ;
      RECT 81.785 3.155 81.8 3.463 ;
      RECT 81.935 4.52 81.94 4.72 ;
      RECT 81.4 4.585 81.445 4.72 ;
      RECT 81.97 4.52 81.99 4.693 ;
      RECT 81.94 4.52 81.97 4.708 ;
      RECT 81.875 4.52 81.935 4.745 ;
      RECT 81.86 4.52 81.875 4.775 ;
      RECT 81.845 4.52 81.86 4.788 ;
      RECT 81.825 4.52 81.845 4.803 ;
      RECT 81.82 4.52 81.825 4.812 ;
      RECT 81.81 4.524 81.82 4.817 ;
      RECT 81.795 4.534 81.81 4.828 ;
      RECT 81.77 4.55 81.795 4.838 ;
      RECT 81.76 4.564 81.77 4.84 ;
      RECT 81.74 4.576 81.76 4.837 ;
      RECT 81.71 4.597 81.74 4.831 ;
      RECT 81.7 4.609 81.71 4.826 ;
      RECT 81.69 4.607 81.7 4.823 ;
      RECT 81.675 4.606 81.69 4.818 ;
      RECT 81.67 4.605 81.675 4.813 ;
      RECT 81.635 4.603 81.67 4.803 ;
      RECT 81.615 4.6 81.635 4.785 ;
      RECT 81.605 4.598 81.615 4.78 ;
      RECT 81.595 4.597 81.605 4.775 ;
      RECT 81.56 4.595 81.595 4.763 ;
      RECT 81.505 4.591 81.56 4.743 ;
      RECT 81.495 4.589 81.505 4.728 ;
      RECT 81.49 4.589 81.495 4.723 ;
      RECT 81.445 4.587 81.49 4.72 ;
      RECT 81.35 4.585 81.4 4.724 ;
      RECT 81.34 4.586 81.35 4.729 ;
      RECT 81.28 4.593 81.34 4.743 ;
      RECT 81.255 4.601 81.28 4.763 ;
      RECT 81.245 4.605 81.255 4.775 ;
      RECT 81.24 4.606 81.245 4.78 ;
      RECT 81.225 4.608 81.24 4.783 ;
      RECT 81.21 4.61 81.225 4.788 ;
      RECT 81.205 4.61 81.21 4.791 ;
      RECT 81.16 4.615 81.205 4.802 ;
      RECT 81.155 4.619 81.16 4.814 ;
      RECT 81.13 4.615 81.155 4.818 ;
      RECT 81.12 4.611 81.13 4.822 ;
      RECT 81.11 4.61 81.12 4.826 ;
      RECT 81.095 4.6 81.11 4.832 ;
      RECT 81.09 4.588 81.095 4.836 ;
      RECT 81.085 4.585 81.09 4.837 ;
      RECT 81.08 4.582 81.085 4.839 ;
      RECT 81.065 4.57 81.08 4.838 ;
      RECT 81.05 4.552 81.065 4.835 ;
      RECT 81.03 4.531 81.05 4.828 ;
      RECT 80.965 4.52 81.03 4.8 ;
      RECT 80.961 4.52 80.965 4.779 ;
      RECT 80.875 4.52 80.961 4.749 ;
      RECT 80.86 4.52 80.875 4.705 ;
      RECT 81.51 4.871 81.525 5.13 ;
      RECT 81.51 4.886 81.53 5.129 ;
      RECT 81.426 4.886 81.53 5.127 ;
      RECT 81.426 4.9 81.535 5.126 ;
      RECT 81.34 4.942 81.54 5.123 ;
      RECT 81.335 4.885 81.525 5.118 ;
      RECT 81.335 4.956 81.545 5.115 ;
      RECT 81.33 4.987 81.545 5.113 ;
      RECT 81.335 4.984 81.56 5.103 ;
      RECT 81.33 5.03 81.575 5.088 ;
      RECT 81.33 5.058 81.58 5.073 ;
      RECT 81.34 4.86 81.51 5.123 ;
      RECT 81.1 3.87 81.27 4.04 ;
      RECT 81.065 3.87 81.27 4.035 ;
      RECT 81.055 3.87 81.27 4.028 ;
      RECT 81.05 3.855 81.22 4.025 ;
      RECT 79.88 4.392 80.145 4.835 ;
      RECT 79.875 4.363 80.09 4.833 ;
      RECT 79.87 4.517 80.15 4.828 ;
      RECT 79.875 4.412 80.15 4.828 ;
      RECT 79.875 4.423 80.16 4.815 ;
      RECT 79.875 4.37 80.12 4.833 ;
      RECT 79.88 4.357 80.09 4.835 ;
      RECT 79.88 4.355 80.04 4.835 ;
      RECT 79.981 4.347 80.04 4.835 ;
      RECT 79.895 4.348 80.04 4.835 ;
      RECT 79.981 4.346 80.03 4.835 ;
      RECT 79.785 3.161 79.96 3.46 ;
      RECT 79.835 3.123 79.96 3.46 ;
      RECT 79.82 3.125 80.046 3.452 ;
      RECT 79.82 3.128 80.085 3.439 ;
      RECT 79.82 3.129 80.095 3.425 ;
      RECT 79.775 3.18 80.095 3.415 ;
      RECT 79.82 3.13 80.1 3.41 ;
      RECT 79.775 3.34 80.105 3.4 ;
      RECT 79.76 3.2 80.1 3.34 ;
      RECT 79.755 3.216 80.1 3.28 ;
      RECT 79.8 3.14 80.1 3.41 ;
      RECT 79.835 3.121 79.921 3.46 ;
      RECT 78.295 7.31 78.465 8.78 ;
      RECT 78.295 7.31 78.47 8.57 ;
      RECT 77.925 9.26 78.395 9.43 ;
      RECT 77.925 8.24 78.095 9.43 ;
      RECT 77.92 3.035 78.09 4.225 ;
      RECT 77.92 3.035 78.39 3.205 ;
      RECT 77.305 3.895 77.48 5.155 ;
      RECT 77.305 3.685 77.475 5.155 ;
      RECT 77.305 7.31 77.475 8.78 ;
      RECT 77.305 7.31 77.48 8.57 ;
      RECT 76.935 3.035 77.105 4.225 ;
      RECT 76.935 3.035 77.405 3.205 ;
      RECT 76.935 9.26 77.405 9.43 ;
      RECT 76.935 8.24 77.105 9.43 ;
      RECT 75.945 4.015 76.12 5.155 ;
      RECT 75.945 1.865 76.115 5.155 ;
      RECT 75.945 1.865 76.12 2.415 ;
      RECT 75.945 10.05 76.12 10.6 ;
      RECT 75.945 7.31 76.115 10.6 ;
      RECT 75.945 7.31 76.12 8.45 ;
      RECT 75.515 3.895 75.69 5.155 ;
      RECT 75.515 2.945 75.685 5.155 ;
      RECT 75.515 7.31 75.685 9.52 ;
      RECT 75.515 7.31 75.69 8.57 ;
      RECT 75.085 3.925 75.255 5.155 ;
      RECT 75.145 2.145 75.315 4.095 ;
      RECT 75.085 1.865 75.255 2.315 ;
      RECT 75.085 10.15 75.255 10.6 ;
      RECT 75.145 8.37 75.315 10.32 ;
      RECT 75.085 7.31 75.255 8.54 ;
      RECT 74.56 3.895 74.735 5.155 ;
      RECT 74.56 1.865 74.73 5.155 ;
      RECT 74.56 3.365 74.97 3.695 ;
      RECT 74.56 2.525 74.97 2.855 ;
      RECT 74.56 1.865 74.735 2.355 ;
      RECT 74.56 10.11 74.735 10.6 ;
      RECT 74.56 7.31 74.73 10.6 ;
      RECT 74.56 9.61 74.97 9.94 ;
      RECT 74.56 8.77 74.97 9.1 ;
      RECT 74.56 7.31 74.735 8.57 ;
      RECT 72.49 4.421 72.495 4.593 ;
      RECT 72.485 4.414 72.49 4.683 ;
      RECT 72.48 4.408 72.485 4.702 ;
      RECT 72.46 4.402 72.48 4.712 ;
      RECT 72.445 4.397 72.46 4.72 ;
      RECT 72.408 4.391 72.445 4.718 ;
      RECT 72.322 4.377 72.408 4.714 ;
      RECT 72.236 4.359 72.322 4.709 ;
      RECT 72.15 4.34 72.236 4.703 ;
      RECT 72.12 4.328 72.15 4.699 ;
      RECT 72.1 4.322 72.12 4.698 ;
      RECT 72.035 4.32 72.1 4.696 ;
      RECT 72.02 4.32 72.035 4.688 ;
      RECT 72.005 4.32 72.02 4.675 ;
      RECT 72 4.32 72.005 4.665 ;
      RECT 71.985 4.32 72 4.643 ;
      RECT 71.97 4.32 71.985 4.61 ;
      RECT 71.965 4.32 71.97 4.588 ;
      RECT 71.955 4.32 71.965 4.57 ;
      RECT 71.94 4.32 71.955 4.548 ;
      RECT 71.92 4.32 71.94 4.51 ;
      RECT 72.27 3.605 72.305 4.044 ;
      RECT 72.27 3.605 72.31 4.043 ;
      RECT 72.215 3.665 72.31 4.042 ;
      RECT 72.08 3.837 72.31 4.041 ;
      RECT 72.19 3.715 72.31 4.041 ;
      RECT 72.08 3.837 72.335 4.031 ;
      RECT 72.135 3.782 72.415 3.948 ;
      RECT 72.31 3.576 72.315 4.039 ;
      RECT 72.165 3.752 72.455 3.825 ;
      RECT 72.18 3.735 72.31 4.041 ;
      RECT 72.315 3.575 72.485 3.763 ;
      RECT 72.305 3.578 72.485 3.763 ;
      RECT 71.81 3.455 71.98 3.765 ;
      RECT 71.81 3.455 71.985 3.738 ;
      RECT 71.81 3.455 71.99 3.715 ;
      RECT 71.81 3.455 72 3.665 ;
      RECT 71.805 3.56 72 3.635 ;
      RECT 71.84 3.13 72.01 3.608 ;
      RECT 71.84 3.13 72.025 3.529 ;
      RECT 71.83 3.34 72.025 3.529 ;
      RECT 71.84 3.14 72.035 3.444 ;
      RECT 71.77 3.882 71.775 4.085 ;
      RECT 71.76 3.87 71.77 4.195 ;
      RECT 71.735 3.87 71.76 4.235 ;
      RECT 71.655 3.87 71.735 4.32 ;
      RECT 71.645 3.87 71.655 4.39 ;
      RECT 71.62 3.87 71.645 4.413 ;
      RECT 71.6 3.87 71.62 4.448 ;
      RECT 71.555 3.88 71.6 4.491 ;
      RECT 71.545 3.892 71.555 4.528 ;
      RECT 71.525 3.906 71.545 4.548 ;
      RECT 71.515 3.924 71.525 4.564 ;
      RECT 71.5 3.95 71.515 4.574 ;
      RECT 71.485 3.991 71.5 4.588 ;
      RECT 71.475 4.026 71.485 4.598 ;
      RECT 71.47 4.042 71.475 4.603 ;
      RECT 71.46 4.057 71.47 4.608 ;
      RECT 71.44 4.1 71.46 4.618 ;
      RECT 71.42 4.137 71.44 4.631 ;
      RECT 71.385 4.16 71.42 4.649 ;
      RECT 71.375 4.174 71.385 4.665 ;
      RECT 71.355 4.184 71.375 4.675 ;
      RECT 71.35 4.193 71.355 4.683 ;
      RECT 71.34 4.2 71.35 4.69 ;
      RECT 71.33 4.207 71.34 4.698 ;
      RECT 71.315 4.217 71.33 4.706 ;
      RECT 71.305 4.231 71.315 4.716 ;
      RECT 71.295 4.243 71.305 4.728 ;
      RECT 71.28 4.265 71.295 4.741 ;
      RECT 71.27 4.287 71.28 4.752 ;
      RECT 71.26 4.307 71.27 4.761 ;
      RECT 71.255 4.322 71.26 4.768 ;
      RECT 71.225 4.355 71.255 4.782 ;
      RECT 71.215 4.39 71.225 4.797 ;
      RECT 71.21 4.397 71.215 4.803 ;
      RECT 71.19 4.412 71.21 4.81 ;
      RECT 71.185 4.427 71.19 4.818 ;
      RECT 71.18 4.436 71.185 4.823 ;
      RECT 71.165 4.442 71.18 4.83 ;
      RECT 71.16 4.448 71.165 4.838 ;
      RECT 71.155 4.452 71.16 4.845 ;
      RECT 71.15 4.456 71.155 4.855 ;
      RECT 71.14 4.461 71.15 4.865 ;
      RECT 71.12 4.472 71.14 4.893 ;
      RECT 71.105 4.484 71.12 4.92 ;
      RECT 71.085 4.497 71.105 4.945 ;
      RECT 71.065 4.512 71.085 4.969 ;
      RECT 71.05 4.527 71.065 4.984 ;
      RECT 71.045 4.538 71.05 4.993 ;
      RECT 70.98 4.583 71.045 5.003 ;
      RECT 70.945 4.642 70.98 5.016 ;
      RECT 70.94 4.665 70.945 5.022 ;
      RECT 70.935 4.672 70.94 5.024 ;
      RECT 70.92 4.682 70.935 5.027 ;
      RECT 70.89 4.707 70.92 5.031 ;
      RECT 70.885 4.725 70.89 5.035 ;
      RECT 70.88 4.732 70.885 5.036 ;
      RECT 70.86 4.74 70.88 5.04 ;
      RECT 70.85 4.747 70.86 5.044 ;
      RECT 70.806 4.758 70.85 5.051 ;
      RECT 70.72 4.786 70.806 5.067 ;
      RECT 70.66 4.81 70.72 5.085 ;
      RECT 70.615 4.82 70.66 5.099 ;
      RECT 70.556 4.828 70.615 5.113 ;
      RECT 70.47 4.835 70.556 5.132 ;
      RECT 70.445 4.84 70.47 5.147 ;
      RECT 70.365 4.843 70.445 5.15 ;
      RECT 70.285 4.847 70.365 5.137 ;
      RECT 70.276 4.85 70.285 5.122 ;
      RECT 70.19 4.85 70.276 5.107 ;
      RECT 70.13 4.852 70.19 5.084 ;
      RECT 70.126 4.855 70.13 5.074 ;
      RECT 70.04 4.855 70.126 5.059 ;
      RECT 69.965 4.855 70.04 5.035 ;
      RECT 71.28 3.864 71.29 4.04 ;
      RECT 71.235 3.831 71.28 4.04 ;
      RECT 71.19 3.782 71.235 4.04 ;
      RECT 71.16 3.752 71.19 4.041 ;
      RECT 71.155 3.735 71.16 4.042 ;
      RECT 71.13 3.715 71.155 4.043 ;
      RECT 71.115 3.69 71.13 4.044 ;
      RECT 71.11 3.677 71.115 4.045 ;
      RECT 71.105 3.671 71.11 4.043 ;
      RECT 71.1 3.663 71.105 4.037 ;
      RECT 71.075 3.655 71.1 4.017 ;
      RECT 71.055 3.644 71.075 3.988 ;
      RECT 71.025 3.629 71.055 3.959 ;
      RECT 71.005 3.615 71.025 3.931 ;
      RECT 70.995 3.609 71.005 3.91 ;
      RECT 70.99 3.606 70.995 3.893 ;
      RECT 70.985 3.603 70.99 3.878 ;
      RECT 70.97 3.598 70.985 3.843 ;
      RECT 70.965 3.594 70.97 3.81 ;
      RECT 70.945 3.589 70.965 3.786 ;
      RECT 70.915 3.581 70.945 3.751 ;
      RECT 70.9 3.575 70.915 3.728 ;
      RECT 70.86 3.568 70.9 3.713 ;
      RECT 70.835 3.56 70.86 3.693 ;
      RECT 70.815 3.555 70.835 3.683 ;
      RECT 70.78 3.549 70.815 3.678 ;
      RECT 70.735 3.54 70.78 3.677 ;
      RECT 70.705 3.536 70.735 3.679 ;
      RECT 70.62 3.544 70.705 3.683 ;
      RECT 70.55 3.555 70.62 3.705 ;
      RECT 70.537 3.561 70.55 3.728 ;
      RECT 70.451 3.568 70.537 3.75 ;
      RECT 70.365 3.58 70.451 3.787 ;
      RECT 70.365 3.957 70.375 4.195 ;
      RECT 70.36 3.586 70.365 3.81 ;
      RECT 70.355 3.842 70.365 4.195 ;
      RECT 70.355 3.587 70.36 3.815 ;
      RECT 70.35 3.588 70.355 4.195 ;
      RECT 70.326 3.59 70.35 4.196 ;
      RECT 70.24 3.598 70.326 4.198 ;
      RECT 70.22 3.612 70.24 4.201 ;
      RECT 70.215 3.64 70.22 4.202 ;
      RECT 70.21 3.652 70.215 4.203 ;
      RECT 70.205 3.667 70.21 4.204 ;
      RECT 70.195 3.697 70.205 4.205 ;
      RECT 70.19 3.735 70.195 4.203 ;
      RECT 70.185 3.755 70.19 4.198 ;
      RECT 70.17 3.79 70.185 4.183 ;
      RECT 70.16 3.842 70.17 4.163 ;
      RECT 70.155 3.872 70.16 4.151 ;
      RECT 70.14 3.885 70.155 4.134 ;
      RECT 70.115 3.889 70.14 4.101 ;
      RECT 70.1 3.887 70.115 4.078 ;
      RECT 70.085 3.886 70.1 4.075 ;
      RECT 70.025 3.884 70.085 4.073 ;
      RECT 70.015 3.882 70.025 4.068 ;
      RECT 69.975 3.881 70.015 4.065 ;
      RECT 69.905 3.878 69.975 4.063 ;
      RECT 69.85 3.876 69.905 4.058 ;
      RECT 69.78 3.87 69.85 4.053 ;
      RECT 69.771 3.87 69.78 4.05 ;
      RECT 69.685 3.87 69.771 4.045 ;
      RECT 69.68 3.87 69.685 4.04 ;
      RECT 70.985 3.105 71.16 3.455 ;
      RECT 70.985 3.12 71.17 3.453 ;
      RECT 70.96 3.07 71.105 3.45 ;
      RECT 70.94 3.071 71.105 3.443 ;
      RECT 70.93 3.072 71.115 3.438 ;
      RECT 70.9 3.073 71.115 3.425 ;
      RECT 70.85 3.074 71.115 3.401 ;
      RECT 70.845 3.076 71.115 3.386 ;
      RECT 70.845 3.142 71.175 3.38 ;
      RECT 70.825 3.083 71.13 3.36 ;
      RECT 70.815 3.092 71.14 3.215 ;
      RECT 70.825 3.087 71.14 3.36 ;
      RECT 70.845 3.077 71.13 3.386 ;
      RECT 70.43 4.402 70.6 4.69 ;
      RECT 70.425 4.42 70.61 4.685 ;
      RECT 70.39 4.428 70.675 4.605 ;
      RECT 70.39 4.428 70.761 4.595 ;
      RECT 70.39 4.428 70.815 4.541 ;
      RECT 70.675 4.325 70.845 4.509 ;
      RECT 70.39 4.48 70.85 4.497 ;
      RECT 70.375 4.45 70.845 4.493 ;
      RECT 70.635 4.332 70.675 4.644 ;
      RECT 70.515 4.369 70.845 4.509 ;
      RECT 70.61 4.344 70.635 4.67 ;
      RECT 70.6 4.351 70.845 4.509 ;
      RECT 70.731 3.815 70.8 4.074 ;
      RECT 70.731 3.87 70.805 4.073 ;
      RECT 70.645 3.87 70.805 4.072 ;
      RECT 70.64 3.87 70.81 4.065 ;
      RECT 70.63 3.815 70.8 4.06 ;
      RECT 70.31 10.05 70.485 10.6 ;
      RECT 70.31 7.31 70.48 10.6 ;
      RECT 70.31 7.31 70.485 8.45 ;
      RECT 70.01 3.114 70.185 3.415 ;
      RECT 69.995 3.102 70.01 3.4 ;
      RECT 69.965 3.101 69.995 3.353 ;
      RECT 69.965 3.119 70.19 3.348 ;
      RECT 69.95 3.103 70.01 3.313 ;
      RECT 69.945 3.125 70.2 3.213 ;
      RECT 69.945 3.108 70.096 3.213 ;
      RECT 69.945 3.11 70.1 3.213 ;
      RECT 69.95 3.106 70.096 3.313 ;
      RECT 70.055 4.342 70.06 4.69 ;
      RECT 70.045 4.332 70.055 4.696 ;
      RECT 70.01 4.322 70.045 4.698 ;
      RECT 69.972 4.317 70.01 4.702 ;
      RECT 69.886 4.31 69.972 4.709 ;
      RECT 69.8 4.3 69.886 4.719 ;
      RECT 69.755 4.295 69.8 4.727 ;
      RECT 69.751 4.295 69.755 4.731 ;
      RECT 69.665 4.295 69.751 4.738 ;
      RECT 69.65 4.295 69.665 4.738 ;
      RECT 69.64 4.293 69.65 4.71 ;
      RECT 69.63 4.289 69.64 4.653 ;
      RECT 69.61 4.283 69.63 4.585 ;
      RECT 69.605 4.279 69.61 4.533 ;
      RECT 69.595 4.278 69.605 4.5 ;
      RECT 69.545 4.276 69.595 4.485 ;
      RECT 69.52 4.274 69.545 4.48 ;
      RECT 69.477 4.272 69.52 4.476 ;
      RECT 69.391 4.268 69.477 4.464 ;
      RECT 69.305 4.263 69.391 4.448 ;
      RECT 69.275 4.26 69.305 4.435 ;
      RECT 69.25 4.259 69.275 4.423 ;
      RECT 69.245 4.259 69.25 4.413 ;
      RECT 69.205 4.258 69.245 4.405 ;
      RECT 69.19 4.257 69.205 4.398 ;
      RECT 69.14 4.256 69.19 4.39 ;
      RECT 69.138 4.255 69.14 4.385 ;
      RECT 69.052 4.253 69.138 4.385 ;
      RECT 68.966 4.248 69.052 4.385 ;
      RECT 68.88 4.244 68.966 4.385 ;
      RECT 68.831 4.24 68.88 4.383 ;
      RECT 68.745 4.237 68.831 4.378 ;
      RECT 68.722 4.234 68.745 4.374 ;
      RECT 68.636 4.231 68.722 4.369 ;
      RECT 68.55 4.227 68.636 4.36 ;
      RECT 68.525 4.22 68.55 4.355 ;
      RECT 68.465 4.185 68.525 4.352 ;
      RECT 68.445 4.11 68.465 4.349 ;
      RECT 68.44 4.052 68.445 4.348 ;
      RECT 68.415 3.992 68.44 4.347 ;
      RECT 68.34 3.87 68.415 4.343 ;
      RECT 68.33 3.87 68.34 4.335 ;
      RECT 68.315 3.87 68.33 4.325 ;
      RECT 68.3 3.87 68.315 4.295 ;
      RECT 68.285 3.87 68.3 4.24 ;
      RECT 68.27 3.87 68.285 4.178 ;
      RECT 68.245 3.87 68.27 4.103 ;
      RECT 68.24 3.87 68.245 4.053 ;
      RECT 69.88 7.31 70.05 9.52 ;
      RECT 69.88 7.31 70.055 8.57 ;
      RECT 69.585 3.415 69.605 3.724 ;
      RECT 69.571 3.417 69.62 3.721 ;
      RECT 69.571 3.422 69.64 3.712 ;
      RECT 69.485 3.42 69.62 3.706 ;
      RECT 69.485 3.428 69.675 3.689 ;
      RECT 69.45 3.43 69.675 3.688 ;
      RECT 69.42 3.438 69.675 3.679 ;
      RECT 69.41 3.443 69.695 3.665 ;
      RECT 69.45 3.433 69.695 3.665 ;
      RECT 69.45 3.436 69.705 3.653 ;
      RECT 69.42 3.438 69.715 3.64 ;
      RECT 69.42 3.442 69.725 3.583 ;
      RECT 69.41 3.447 69.73 3.498 ;
      RECT 69.571 3.415 69.605 3.721 ;
      RECT 69.01 3.518 69.015 3.73 ;
      RECT 68.885 3.515 68.9 3.73 ;
      RECT 68.35 3.545 68.42 3.73 ;
      RECT 68.235 3.545 68.27 3.725 ;
      RECT 69.356 3.847 69.375 4.041 ;
      RECT 69.27 3.802 69.356 4.042 ;
      RECT 69.26 3.755 69.27 4.044 ;
      RECT 69.255 3.735 69.26 4.045 ;
      RECT 69.235 3.7 69.255 4.046 ;
      RECT 69.22 3.65 69.235 4.047 ;
      RECT 69.2 3.587 69.22 4.048 ;
      RECT 69.19 3.55 69.2 4.049 ;
      RECT 69.175 3.539 69.19 4.05 ;
      RECT 69.17 3.531 69.175 4.048 ;
      RECT 69.16 3.53 69.17 4.04 ;
      RECT 69.13 3.527 69.16 4.019 ;
      RECT 69.055 3.522 69.13 3.964 ;
      RECT 69.04 3.518 69.055 3.91 ;
      RECT 69.03 3.518 69.04 3.805 ;
      RECT 69.015 3.518 69.03 3.738 ;
      RECT 69 3.518 69.01 3.728 ;
      RECT 68.945 3.517 69 3.725 ;
      RECT 68.9 3.515 68.945 3.728 ;
      RECT 68.872 3.515 68.885 3.731 ;
      RECT 68.786 3.519 68.872 3.733 ;
      RECT 68.7 3.525 68.786 3.738 ;
      RECT 68.68 3.529 68.7 3.74 ;
      RECT 68.678 3.53 68.68 3.739 ;
      RECT 68.592 3.532 68.678 3.738 ;
      RECT 68.506 3.537 68.592 3.735 ;
      RECT 68.42 3.542 68.506 3.732 ;
      RECT 68.27 3.545 68.35 3.728 ;
      RECT 68.925 10.11 69.1 10.6 ;
      RECT 68.925 7.31 69.095 10.6 ;
      RECT 68.925 9.61 69.335 9.94 ;
      RECT 68.925 8.77 69.335 9.1 ;
      RECT 68.925 7.31 69.1 8.57 ;
      RECT 69.046 4.52 69.095 4.854 ;
      RECT 69.046 4.52 69.1 4.853 ;
      RECT 68.96 4.52 69.1 4.852 ;
      RECT 68.735 4.628 69.105 4.85 ;
      RECT 68.96 4.52 69.13 4.843 ;
      RECT 68.93 4.532 69.135 4.834 ;
      RECT 68.915 4.55 69.14 4.831 ;
      RECT 68.73 4.634 69.14 4.758 ;
      RECT 68.725 4.641 69.14 4.718 ;
      RECT 68.74 4.607 69.14 4.831 ;
      RECT 68.901 4.553 69.105 4.85 ;
      RECT 68.815 4.573 69.14 4.831 ;
      RECT 68.915 4.547 69.135 4.834 ;
      RECT 68.685 3.871 68.875 4.065 ;
      RECT 68.68 3.873 68.875 4.064 ;
      RECT 68.675 3.877 68.89 4.061 ;
      RECT 68.69 3.87 68.89 4.061 ;
      RECT 68.675 3.98 68.895 4.056 ;
      RECT 67.97 4.48 68.061 4.778 ;
      RECT 67.965 4.482 68.14 4.773 ;
      RECT 67.97 4.48 68.14 4.773 ;
      RECT 67.965 4.486 68.16 4.771 ;
      RECT 67.965 4.541 68.2 4.77 ;
      RECT 67.965 4.576 68.215 4.764 ;
      RECT 67.965 4.61 68.225 4.754 ;
      RECT 67.955 4.49 68.16 4.605 ;
      RECT 67.955 4.51 68.175 4.605 ;
      RECT 67.955 4.493 68.165 4.605 ;
      RECT 68.18 3.261 68.185 3.323 ;
      RECT 68.175 3.183 68.18 3.346 ;
      RECT 68.17 3.14 68.175 3.357 ;
      RECT 68.165 3.13 68.17 3.369 ;
      RECT 68.16 3.13 68.165 3.378 ;
      RECT 68.135 3.13 68.16 3.41 ;
      RECT 68.13 3.13 68.135 3.443 ;
      RECT 68.115 3.13 68.13 3.468 ;
      RECT 68.105 3.13 68.115 3.495 ;
      RECT 68.1 3.13 68.105 3.508 ;
      RECT 68.095 3.13 68.1 3.523 ;
      RECT 68.085 3.13 68.095 3.538 ;
      RECT 68.08 3.13 68.085 3.558 ;
      RECT 68.055 3.13 68.08 3.593 ;
      RECT 68.01 3.13 68.055 3.638 ;
      RECT 68 3.13 68.01 3.651 ;
      RECT 67.915 3.215 68 3.658 ;
      RECT 67.88 3.337 67.915 3.667 ;
      RECT 67.875 3.377 67.88 3.671 ;
      RECT 67.855 3.4 67.875 3.673 ;
      RECT 67.85 3.43 67.855 3.676 ;
      RECT 67.84 3.442 67.85 3.677 ;
      RECT 67.795 3.465 67.84 3.682 ;
      RECT 67.755 3.495 67.795 3.69 ;
      RECT 67.72 3.507 67.755 3.696 ;
      RECT 67.715 3.512 67.72 3.7 ;
      RECT 67.645 3.522 67.715 3.707 ;
      RECT 67.605 3.532 67.645 3.717 ;
      RECT 67.585 3.537 67.605 3.723 ;
      RECT 67.575 3.541 67.585 3.728 ;
      RECT 67.57 3.544 67.575 3.731 ;
      RECT 67.56 3.545 67.57 3.732 ;
      RECT 67.535 3.547 67.56 3.736 ;
      RECT 67.525 3.552 67.535 3.739 ;
      RECT 67.48 3.56 67.525 3.74 ;
      RECT 67.355 3.565 67.48 3.74 ;
      RECT 67.91 3.862 67.93 4.044 ;
      RECT 67.861 3.847 67.91 4.043 ;
      RECT 67.775 3.862 67.93 4.041 ;
      RECT 67.76 3.862 67.93 4.04 ;
      RECT 67.725 3.84 67.895 4.025 ;
      RECT 67.795 4.86 67.81 5.069 ;
      RECT 67.795 4.868 67.815 5.068 ;
      RECT 67.74 4.868 67.815 5.067 ;
      RECT 67.72 4.872 67.82 5.065 ;
      RECT 67.7 4.822 67.74 5.064 ;
      RECT 67.645 4.88 67.825 5.062 ;
      RECT 67.61 4.837 67.74 5.06 ;
      RECT 67.606 4.84 67.795 5.059 ;
      RECT 67.52 4.848 67.795 5.057 ;
      RECT 67.52 4.892 67.83 5.05 ;
      RECT 67.51 4.985 67.83 5.048 ;
      RECT 67.52 4.904 67.835 5.033 ;
      RECT 67.52 4.925 67.85 5.003 ;
      RECT 67.52 4.952 67.855 4.973 ;
      RECT 67.645 4.83 67.74 5.062 ;
      RECT 67.275 3.875 67.28 4.413 ;
      RECT 67.08 4.205 67.085 4.4 ;
      RECT 65.38 3.87 65.395 4.25 ;
      RECT 67.445 3.87 67.45 4.04 ;
      RECT 67.44 3.87 67.445 4.05 ;
      RECT 67.435 3.87 67.44 4.063 ;
      RECT 67.41 3.87 67.435 4.105 ;
      RECT 67.385 3.87 67.41 4.178 ;
      RECT 67.37 3.87 67.385 4.23 ;
      RECT 67.365 3.87 67.37 4.26 ;
      RECT 67.34 3.87 67.365 4.3 ;
      RECT 67.325 3.87 67.34 4.355 ;
      RECT 67.32 3.87 67.325 4.388 ;
      RECT 67.295 3.87 67.32 4.408 ;
      RECT 67.28 3.87 67.295 4.414 ;
      RECT 67.21 3.905 67.275 4.41 ;
      RECT 67.16 3.96 67.21 4.405 ;
      RECT 67.15 3.992 67.16 4.403 ;
      RECT 67.145 4.017 67.15 4.403 ;
      RECT 67.125 4.09 67.145 4.403 ;
      RECT 67.115 4.17 67.125 4.402 ;
      RECT 67.1 4.2 67.115 4.402 ;
      RECT 67.085 4.205 67.1 4.401 ;
      RECT 67.025 4.207 67.08 4.398 ;
      RECT 66.995 4.212 67.025 4.394 ;
      RECT 66.993 4.215 66.995 4.393 ;
      RECT 66.907 4.217 66.993 4.39 ;
      RECT 66.821 4.223 66.907 4.384 ;
      RECT 66.735 4.228 66.821 4.378 ;
      RECT 66.662 4.233 66.735 4.379 ;
      RECT 66.576 4.239 66.662 4.387 ;
      RECT 66.49 4.245 66.576 4.396 ;
      RECT 66.47 4.249 66.49 4.401 ;
      RECT 66.423 4.251 66.47 4.404 ;
      RECT 66.337 4.256 66.423 4.41 ;
      RECT 66.251 4.261 66.337 4.419 ;
      RECT 66.165 4.267 66.251 4.427 ;
      RECT 66.08 4.265 66.165 4.436 ;
      RECT 66.076 4.26 66.08 4.44 ;
      RECT 65.99 4.255 66.076 4.432 ;
      RECT 65.926 4.246 65.99 4.42 ;
      RECT 65.84 4.237 65.926 4.407 ;
      RECT 65.816 4.23 65.84 4.398 ;
      RECT 65.73 4.224 65.816 4.385 ;
      RECT 65.69 4.217 65.73 4.371 ;
      RECT 65.685 4.207 65.69 4.367 ;
      RECT 65.675 4.195 65.685 4.366 ;
      RECT 65.655 4.165 65.675 4.363 ;
      RECT 65.6 4.085 65.655 4.357 ;
      RECT 65.58 4.004 65.6 4.352 ;
      RECT 65.56 3.962 65.58 4.348 ;
      RECT 65.535 3.915 65.56 4.342 ;
      RECT 65.53 3.89 65.535 4.339 ;
      RECT 65.495 3.87 65.53 4.334 ;
      RECT 65.486 3.87 65.495 4.327 ;
      RECT 65.4 3.87 65.486 4.297 ;
      RECT 65.395 3.87 65.4 4.26 ;
      RECT 65.36 3.87 65.38 4.182 ;
      RECT 65.355 3.912 65.36 4.147 ;
      RECT 65.35 3.987 65.355 4.103 ;
      RECT 66.8 3.792 66.975 4.04 ;
      RECT 66.8 3.792 66.98 4.038 ;
      RECT 66.795 3.824 66.98 3.998 ;
      RECT 66.825 3.765 66.995 3.985 ;
      RECT 66.79 3.842 66.995 3.918 ;
      RECT 66.1 3.305 66.27 3.48 ;
      RECT 66.1 3.305 66.442 3.472 ;
      RECT 66.1 3.305 66.525 3.466 ;
      RECT 66.1 3.305 66.56 3.462 ;
      RECT 66.1 3.305 66.58 3.461 ;
      RECT 66.1 3.305 66.666 3.457 ;
      RECT 66.56 3.13 66.73 3.452 ;
      RECT 66.135 3.237 66.76 3.45 ;
      RECT 66.125 3.292 66.765 3.448 ;
      RECT 66.1 3.328 66.775 3.443 ;
      RECT 66.1 3.355 66.78 3.373 ;
      RECT 66.165 3.18 66.74 3.45 ;
      RECT 66.356 3.165 66.74 3.45 ;
      RECT 66.19 3.168 66.74 3.45 ;
      RECT 66.27 3.166 66.356 3.477 ;
      RECT 66.356 3.163 66.735 3.45 ;
      RECT 66.54 3.14 66.735 3.45 ;
      RECT 66.442 3.161 66.735 3.45 ;
      RECT 66.525 3.155 66.54 3.463 ;
      RECT 66.675 4.52 66.68 4.72 ;
      RECT 66.14 4.585 66.185 4.72 ;
      RECT 66.71 4.52 66.73 4.693 ;
      RECT 66.68 4.52 66.71 4.708 ;
      RECT 66.615 4.52 66.675 4.745 ;
      RECT 66.6 4.52 66.615 4.775 ;
      RECT 66.585 4.52 66.6 4.788 ;
      RECT 66.565 4.52 66.585 4.803 ;
      RECT 66.56 4.52 66.565 4.812 ;
      RECT 66.55 4.524 66.56 4.817 ;
      RECT 66.535 4.534 66.55 4.828 ;
      RECT 66.51 4.55 66.535 4.838 ;
      RECT 66.5 4.564 66.51 4.84 ;
      RECT 66.48 4.576 66.5 4.837 ;
      RECT 66.45 4.597 66.48 4.831 ;
      RECT 66.44 4.609 66.45 4.826 ;
      RECT 66.43 4.607 66.44 4.823 ;
      RECT 66.415 4.606 66.43 4.818 ;
      RECT 66.41 4.605 66.415 4.813 ;
      RECT 66.375 4.603 66.41 4.803 ;
      RECT 66.355 4.6 66.375 4.785 ;
      RECT 66.345 4.598 66.355 4.78 ;
      RECT 66.335 4.597 66.345 4.775 ;
      RECT 66.3 4.595 66.335 4.763 ;
      RECT 66.245 4.591 66.3 4.743 ;
      RECT 66.235 4.589 66.245 4.728 ;
      RECT 66.23 4.589 66.235 4.723 ;
      RECT 66.185 4.587 66.23 4.72 ;
      RECT 66.09 4.585 66.14 4.724 ;
      RECT 66.08 4.586 66.09 4.729 ;
      RECT 66.02 4.593 66.08 4.743 ;
      RECT 65.995 4.601 66.02 4.763 ;
      RECT 65.985 4.605 65.995 4.775 ;
      RECT 65.98 4.606 65.985 4.78 ;
      RECT 65.965 4.608 65.98 4.783 ;
      RECT 65.95 4.61 65.965 4.788 ;
      RECT 65.945 4.61 65.95 4.791 ;
      RECT 65.9 4.615 65.945 4.802 ;
      RECT 65.895 4.619 65.9 4.814 ;
      RECT 65.87 4.615 65.895 4.818 ;
      RECT 65.86 4.611 65.87 4.822 ;
      RECT 65.85 4.61 65.86 4.826 ;
      RECT 65.835 4.6 65.85 4.832 ;
      RECT 65.83 4.588 65.835 4.836 ;
      RECT 65.825 4.585 65.83 4.837 ;
      RECT 65.82 4.582 65.825 4.839 ;
      RECT 65.805 4.57 65.82 4.838 ;
      RECT 65.79 4.552 65.805 4.835 ;
      RECT 65.77 4.531 65.79 4.828 ;
      RECT 65.705 4.52 65.77 4.8 ;
      RECT 65.701 4.52 65.705 4.779 ;
      RECT 65.615 4.52 65.701 4.749 ;
      RECT 65.6 4.52 65.615 4.705 ;
      RECT 66.25 4.871 66.265 5.13 ;
      RECT 66.25 4.886 66.27 5.129 ;
      RECT 66.166 4.886 66.27 5.127 ;
      RECT 66.166 4.9 66.275 5.126 ;
      RECT 66.08 4.942 66.28 5.123 ;
      RECT 66.075 4.885 66.265 5.118 ;
      RECT 66.075 4.956 66.285 5.115 ;
      RECT 66.07 4.987 66.285 5.113 ;
      RECT 66.075 4.984 66.3 5.103 ;
      RECT 66.07 5.03 66.315 5.088 ;
      RECT 66.07 5.058 66.32 5.073 ;
      RECT 66.08 4.86 66.25 5.123 ;
      RECT 65.84 3.87 66.01 4.04 ;
      RECT 65.805 3.87 66.01 4.035 ;
      RECT 65.795 3.87 66.01 4.028 ;
      RECT 65.79 3.855 65.96 4.025 ;
      RECT 64.62 4.392 64.885 4.835 ;
      RECT 64.615 4.363 64.83 4.833 ;
      RECT 64.61 4.517 64.89 4.828 ;
      RECT 64.615 4.412 64.89 4.828 ;
      RECT 64.615 4.423 64.9 4.815 ;
      RECT 64.615 4.37 64.86 4.833 ;
      RECT 64.62 4.357 64.83 4.835 ;
      RECT 64.62 4.355 64.78 4.835 ;
      RECT 64.721 4.347 64.78 4.835 ;
      RECT 64.635 4.348 64.78 4.835 ;
      RECT 64.721 4.346 64.77 4.835 ;
      RECT 64.525 3.161 64.7 3.46 ;
      RECT 64.575 3.123 64.7 3.46 ;
      RECT 64.56 3.125 64.786 3.452 ;
      RECT 64.56 3.128 64.825 3.439 ;
      RECT 64.56 3.129 64.835 3.425 ;
      RECT 64.515 3.18 64.835 3.415 ;
      RECT 64.56 3.13 64.84 3.41 ;
      RECT 64.515 3.34 64.845 3.4 ;
      RECT 64.5 3.2 64.84 3.34 ;
      RECT 64.495 3.216 64.84 3.28 ;
      RECT 64.54 3.14 64.84 3.41 ;
      RECT 64.575 3.121 64.661 3.46 ;
      RECT 63.035 7.31 63.205 8.78 ;
      RECT 63.035 7.31 63.21 8.57 ;
      RECT 62.665 9.26 63.135 9.43 ;
      RECT 62.665 8.24 62.835 9.43 ;
      RECT 62.66 3.035 62.83 4.225 ;
      RECT 62.66 3.035 63.13 3.205 ;
      RECT 62.045 3.895 62.22 5.155 ;
      RECT 62.045 3.685 62.215 5.155 ;
      RECT 62.045 7.31 62.215 8.78 ;
      RECT 62.045 7.31 62.22 8.57 ;
      RECT 61.675 3.035 61.845 4.225 ;
      RECT 61.675 3.035 62.145 3.205 ;
      RECT 61.675 9.26 62.145 9.43 ;
      RECT 61.675 8.24 61.845 9.43 ;
      RECT 60.685 4.015 60.86 5.155 ;
      RECT 60.685 1.865 60.855 5.155 ;
      RECT 60.685 1.865 60.86 2.415 ;
      RECT 60.685 10.05 60.86 10.6 ;
      RECT 60.685 7.31 60.855 10.6 ;
      RECT 60.685 7.31 60.86 8.45 ;
      RECT 60.255 3.895 60.43 5.155 ;
      RECT 60.255 2.945 60.425 5.155 ;
      RECT 60.255 7.31 60.425 9.52 ;
      RECT 60.255 7.31 60.43 8.57 ;
      RECT 59.825 3.925 59.995 5.155 ;
      RECT 59.885 2.145 60.055 4.095 ;
      RECT 59.825 1.865 59.995 2.315 ;
      RECT 59.825 10.15 59.995 10.6 ;
      RECT 59.885 8.37 60.055 10.32 ;
      RECT 59.825 7.31 59.995 8.54 ;
      RECT 59.3 3.895 59.475 5.155 ;
      RECT 59.3 1.865 59.47 5.155 ;
      RECT 59.3 3.365 59.71 3.695 ;
      RECT 59.3 2.525 59.71 2.855 ;
      RECT 59.3 1.865 59.475 2.355 ;
      RECT 59.3 10.11 59.475 10.6 ;
      RECT 59.3 7.31 59.47 10.6 ;
      RECT 59.3 9.61 59.71 9.94 ;
      RECT 59.3 8.77 59.71 9.1 ;
      RECT 59.3 7.31 59.475 8.57 ;
      RECT 57.23 4.421 57.235 4.593 ;
      RECT 57.225 4.414 57.23 4.683 ;
      RECT 57.22 4.408 57.225 4.702 ;
      RECT 57.2 4.402 57.22 4.712 ;
      RECT 57.185 4.397 57.2 4.72 ;
      RECT 57.148 4.391 57.185 4.718 ;
      RECT 57.062 4.377 57.148 4.714 ;
      RECT 56.976 4.359 57.062 4.709 ;
      RECT 56.89 4.34 56.976 4.703 ;
      RECT 56.86 4.328 56.89 4.699 ;
      RECT 56.84 4.322 56.86 4.698 ;
      RECT 56.775 4.32 56.84 4.696 ;
      RECT 56.76 4.32 56.775 4.688 ;
      RECT 56.745 4.32 56.76 4.675 ;
      RECT 56.74 4.32 56.745 4.665 ;
      RECT 56.725 4.32 56.74 4.643 ;
      RECT 56.71 4.32 56.725 4.61 ;
      RECT 56.705 4.32 56.71 4.588 ;
      RECT 56.695 4.32 56.705 4.57 ;
      RECT 56.68 4.32 56.695 4.548 ;
      RECT 56.66 4.32 56.68 4.51 ;
      RECT 57.01 3.605 57.045 4.044 ;
      RECT 57.01 3.605 57.05 4.043 ;
      RECT 56.955 3.665 57.05 4.042 ;
      RECT 56.82 3.837 57.05 4.041 ;
      RECT 56.93 3.715 57.05 4.041 ;
      RECT 56.82 3.837 57.075 4.031 ;
      RECT 56.875 3.782 57.155 3.948 ;
      RECT 57.05 3.576 57.055 4.039 ;
      RECT 56.905 3.752 57.195 3.825 ;
      RECT 56.92 3.735 57.05 4.041 ;
      RECT 57.055 3.575 57.225 3.763 ;
      RECT 57.045 3.578 57.225 3.763 ;
      RECT 56.55 3.455 56.72 3.765 ;
      RECT 56.55 3.455 56.725 3.738 ;
      RECT 56.55 3.455 56.73 3.715 ;
      RECT 56.55 3.455 56.74 3.665 ;
      RECT 56.545 3.56 56.74 3.635 ;
      RECT 56.58 3.13 56.75 3.608 ;
      RECT 56.58 3.13 56.765 3.529 ;
      RECT 56.57 3.34 56.765 3.529 ;
      RECT 56.58 3.14 56.775 3.444 ;
      RECT 56.51 3.882 56.515 4.085 ;
      RECT 56.5 3.87 56.51 4.195 ;
      RECT 56.475 3.87 56.5 4.235 ;
      RECT 56.395 3.87 56.475 4.32 ;
      RECT 56.385 3.87 56.395 4.39 ;
      RECT 56.36 3.87 56.385 4.413 ;
      RECT 56.34 3.87 56.36 4.448 ;
      RECT 56.295 3.88 56.34 4.491 ;
      RECT 56.285 3.892 56.295 4.528 ;
      RECT 56.265 3.906 56.285 4.548 ;
      RECT 56.255 3.924 56.265 4.564 ;
      RECT 56.24 3.95 56.255 4.574 ;
      RECT 56.225 3.991 56.24 4.588 ;
      RECT 56.215 4.026 56.225 4.598 ;
      RECT 56.21 4.042 56.215 4.603 ;
      RECT 56.2 4.057 56.21 4.608 ;
      RECT 56.18 4.1 56.2 4.618 ;
      RECT 56.16 4.137 56.18 4.631 ;
      RECT 56.125 4.16 56.16 4.649 ;
      RECT 56.115 4.174 56.125 4.665 ;
      RECT 56.095 4.184 56.115 4.675 ;
      RECT 56.09 4.193 56.095 4.683 ;
      RECT 56.08 4.2 56.09 4.69 ;
      RECT 56.07 4.207 56.08 4.698 ;
      RECT 56.055 4.217 56.07 4.706 ;
      RECT 56.045 4.231 56.055 4.716 ;
      RECT 56.035 4.243 56.045 4.728 ;
      RECT 56.02 4.265 56.035 4.741 ;
      RECT 56.01 4.287 56.02 4.752 ;
      RECT 56 4.307 56.01 4.761 ;
      RECT 55.995 4.322 56 4.768 ;
      RECT 55.965 4.355 55.995 4.782 ;
      RECT 55.955 4.39 55.965 4.797 ;
      RECT 55.95 4.397 55.955 4.803 ;
      RECT 55.93 4.412 55.95 4.81 ;
      RECT 55.925 4.427 55.93 4.818 ;
      RECT 55.92 4.436 55.925 4.823 ;
      RECT 55.905 4.442 55.92 4.83 ;
      RECT 55.9 4.448 55.905 4.838 ;
      RECT 55.895 4.452 55.9 4.845 ;
      RECT 55.89 4.456 55.895 4.855 ;
      RECT 55.88 4.461 55.89 4.865 ;
      RECT 55.86 4.472 55.88 4.893 ;
      RECT 55.845 4.484 55.86 4.92 ;
      RECT 55.825 4.497 55.845 4.945 ;
      RECT 55.805 4.512 55.825 4.969 ;
      RECT 55.79 4.527 55.805 4.984 ;
      RECT 55.785 4.538 55.79 4.993 ;
      RECT 55.72 4.583 55.785 5.003 ;
      RECT 55.685 4.642 55.72 5.016 ;
      RECT 55.68 4.665 55.685 5.022 ;
      RECT 55.675 4.672 55.68 5.024 ;
      RECT 55.66 4.682 55.675 5.027 ;
      RECT 55.63 4.707 55.66 5.031 ;
      RECT 55.625 4.725 55.63 5.035 ;
      RECT 55.62 4.732 55.625 5.036 ;
      RECT 55.6 4.74 55.62 5.04 ;
      RECT 55.59 4.747 55.6 5.044 ;
      RECT 55.546 4.758 55.59 5.051 ;
      RECT 55.46 4.786 55.546 5.067 ;
      RECT 55.4 4.81 55.46 5.085 ;
      RECT 55.355 4.82 55.4 5.099 ;
      RECT 55.296 4.828 55.355 5.113 ;
      RECT 55.21 4.835 55.296 5.132 ;
      RECT 55.185 4.84 55.21 5.147 ;
      RECT 55.105 4.843 55.185 5.15 ;
      RECT 55.025 4.847 55.105 5.137 ;
      RECT 55.016 4.85 55.025 5.122 ;
      RECT 54.93 4.85 55.016 5.107 ;
      RECT 54.87 4.852 54.93 5.084 ;
      RECT 54.866 4.855 54.87 5.074 ;
      RECT 54.78 4.855 54.866 5.059 ;
      RECT 54.705 4.855 54.78 5.035 ;
      RECT 56.02 3.864 56.03 4.04 ;
      RECT 55.975 3.831 56.02 4.04 ;
      RECT 55.93 3.782 55.975 4.04 ;
      RECT 55.9 3.752 55.93 4.041 ;
      RECT 55.895 3.735 55.9 4.042 ;
      RECT 55.87 3.715 55.895 4.043 ;
      RECT 55.855 3.69 55.87 4.044 ;
      RECT 55.85 3.677 55.855 4.045 ;
      RECT 55.845 3.671 55.85 4.043 ;
      RECT 55.84 3.663 55.845 4.037 ;
      RECT 55.815 3.655 55.84 4.017 ;
      RECT 55.795 3.644 55.815 3.988 ;
      RECT 55.765 3.629 55.795 3.959 ;
      RECT 55.745 3.615 55.765 3.931 ;
      RECT 55.735 3.609 55.745 3.91 ;
      RECT 55.73 3.606 55.735 3.893 ;
      RECT 55.725 3.603 55.73 3.878 ;
      RECT 55.71 3.598 55.725 3.843 ;
      RECT 55.705 3.594 55.71 3.81 ;
      RECT 55.685 3.589 55.705 3.786 ;
      RECT 55.655 3.581 55.685 3.751 ;
      RECT 55.64 3.575 55.655 3.728 ;
      RECT 55.6 3.568 55.64 3.713 ;
      RECT 55.575 3.56 55.6 3.693 ;
      RECT 55.555 3.555 55.575 3.683 ;
      RECT 55.52 3.549 55.555 3.678 ;
      RECT 55.475 3.54 55.52 3.677 ;
      RECT 55.445 3.536 55.475 3.679 ;
      RECT 55.36 3.544 55.445 3.683 ;
      RECT 55.29 3.555 55.36 3.705 ;
      RECT 55.277 3.561 55.29 3.728 ;
      RECT 55.191 3.568 55.277 3.75 ;
      RECT 55.105 3.58 55.191 3.787 ;
      RECT 55.105 3.957 55.115 4.195 ;
      RECT 55.1 3.586 55.105 3.81 ;
      RECT 55.095 3.842 55.105 4.195 ;
      RECT 55.095 3.587 55.1 3.815 ;
      RECT 55.09 3.588 55.095 4.195 ;
      RECT 55.066 3.59 55.09 4.196 ;
      RECT 54.98 3.598 55.066 4.198 ;
      RECT 54.96 3.612 54.98 4.201 ;
      RECT 54.955 3.64 54.96 4.202 ;
      RECT 54.95 3.652 54.955 4.203 ;
      RECT 54.945 3.667 54.95 4.204 ;
      RECT 54.935 3.697 54.945 4.205 ;
      RECT 54.93 3.735 54.935 4.203 ;
      RECT 54.925 3.755 54.93 4.198 ;
      RECT 54.91 3.79 54.925 4.183 ;
      RECT 54.9 3.842 54.91 4.163 ;
      RECT 54.895 3.872 54.9 4.151 ;
      RECT 54.88 3.885 54.895 4.134 ;
      RECT 54.855 3.889 54.88 4.101 ;
      RECT 54.84 3.887 54.855 4.078 ;
      RECT 54.825 3.886 54.84 4.075 ;
      RECT 54.765 3.884 54.825 4.073 ;
      RECT 54.755 3.882 54.765 4.068 ;
      RECT 54.715 3.881 54.755 4.065 ;
      RECT 54.645 3.878 54.715 4.063 ;
      RECT 54.59 3.876 54.645 4.058 ;
      RECT 54.52 3.87 54.59 4.053 ;
      RECT 54.511 3.87 54.52 4.05 ;
      RECT 54.425 3.87 54.511 4.045 ;
      RECT 54.42 3.87 54.425 4.04 ;
      RECT 55.725 3.105 55.9 3.455 ;
      RECT 55.725 3.12 55.91 3.453 ;
      RECT 55.7 3.07 55.845 3.45 ;
      RECT 55.68 3.071 55.845 3.443 ;
      RECT 55.67 3.072 55.855 3.438 ;
      RECT 55.64 3.073 55.855 3.425 ;
      RECT 55.59 3.074 55.855 3.401 ;
      RECT 55.585 3.076 55.855 3.386 ;
      RECT 55.585 3.142 55.915 3.38 ;
      RECT 55.565 3.083 55.87 3.36 ;
      RECT 55.555 3.092 55.88 3.215 ;
      RECT 55.565 3.087 55.88 3.36 ;
      RECT 55.585 3.077 55.87 3.386 ;
      RECT 55.17 4.402 55.34 4.69 ;
      RECT 55.165 4.42 55.35 4.685 ;
      RECT 55.13 4.428 55.415 4.605 ;
      RECT 55.13 4.428 55.501 4.595 ;
      RECT 55.13 4.428 55.555 4.541 ;
      RECT 55.415 4.325 55.585 4.509 ;
      RECT 55.13 4.48 55.59 4.497 ;
      RECT 55.115 4.45 55.585 4.493 ;
      RECT 55.375 4.332 55.415 4.644 ;
      RECT 55.255 4.369 55.585 4.509 ;
      RECT 55.35 4.344 55.375 4.67 ;
      RECT 55.34 4.351 55.585 4.509 ;
      RECT 55.471 3.815 55.54 4.074 ;
      RECT 55.471 3.87 55.545 4.073 ;
      RECT 55.385 3.87 55.545 4.072 ;
      RECT 55.38 3.87 55.55 4.065 ;
      RECT 55.37 3.815 55.54 4.06 ;
      RECT 55.05 10.05 55.225 10.6 ;
      RECT 55.05 7.31 55.22 10.6 ;
      RECT 55.05 7.31 55.225 8.45 ;
      RECT 54.75 3.114 54.925 3.415 ;
      RECT 54.735 3.102 54.75 3.4 ;
      RECT 54.705 3.101 54.735 3.353 ;
      RECT 54.705 3.119 54.93 3.348 ;
      RECT 54.69 3.103 54.75 3.313 ;
      RECT 54.685 3.125 54.94 3.213 ;
      RECT 54.685 3.108 54.836 3.213 ;
      RECT 54.685 3.11 54.84 3.213 ;
      RECT 54.69 3.106 54.836 3.313 ;
      RECT 54.795 4.342 54.8 4.69 ;
      RECT 54.785 4.332 54.795 4.696 ;
      RECT 54.75 4.322 54.785 4.698 ;
      RECT 54.712 4.317 54.75 4.702 ;
      RECT 54.626 4.31 54.712 4.709 ;
      RECT 54.54 4.3 54.626 4.719 ;
      RECT 54.495 4.295 54.54 4.727 ;
      RECT 54.491 4.295 54.495 4.731 ;
      RECT 54.405 4.295 54.491 4.738 ;
      RECT 54.39 4.295 54.405 4.738 ;
      RECT 54.38 4.293 54.39 4.71 ;
      RECT 54.37 4.289 54.38 4.653 ;
      RECT 54.35 4.283 54.37 4.585 ;
      RECT 54.345 4.279 54.35 4.533 ;
      RECT 54.335 4.278 54.345 4.5 ;
      RECT 54.285 4.276 54.335 4.485 ;
      RECT 54.26 4.274 54.285 4.48 ;
      RECT 54.217 4.272 54.26 4.476 ;
      RECT 54.131 4.268 54.217 4.464 ;
      RECT 54.045 4.263 54.131 4.448 ;
      RECT 54.015 4.26 54.045 4.435 ;
      RECT 53.99 4.259 54.015 4.423 ;
      RECT 53.985 4.259 53.99 4.413 ;
      RECT 53.945 4.258 53.985 4.405 ;
      RECT 53.93 4.257 53.945 4.398 ;
      RECT 53.88 4.256 53.93 4.39 ;
      RECT 53.878 4.255 53.88 4.385 ;
      RECT 53.792 4.253 53.878 4.385 ;
      RECT 53.706 4.248 53.792 4.385 ;
      RECT 53.62 4.244 53.706 4.385 ;
      RECT 53.571 4.24 53.62 4.383 ;
      RECT 53.485 4.237 53.571 4.378 ;
      RECT 53.462 4.234 53.485 4.374 ;
      RECT 53.376 4.231 53.462 4.369 ;
      RECT 53.29 4.227 53.376 4.36 ;
      RECT 53.265 4.22 53.29 4.355 ;
      RECT 53.205 4.185 53.265 4.352 ;
      RECT 53.185 4.11 53.205 4.349 ;
      RECT 53.18 4.052 53.185 4.348 ;
      RECT 53.155 3.992 53.18 4.347 ;
      RECT 53.08 3.87 53.155 4.343 ;
      RECT 53.07 3.87 53.08 4.335 ;
      RECT 53.055 3.87 53.07 4.325 ;
      RECT 53.04 3.87 53.055 4.295 ;
      RECT 53.025 3.87 53.04 4.24 ;
      RECT 53.01 3.87 53.025 4.178 ;
      RECT 52.985 3.87 53.01 4.103 ;
      RECT 52.98 3.87 52.985 4.053 ;
      RECT 54.62 7.31 54.79 9.52 ;
      RECT 54.62 7.31 54.795 8.57 ;
      RECT 54.325 3.415 54.345 3.724 ;
      RECT 54.311 3.417 54.36 3.721 ;
      RECT 54.311 3.422 54.38 3.712 ;
      RECT 54.225 3.42 54.36 3.706 ;
      RECT 54.225 3.428 54.415 3.689 ;
      RECT 54.19 3.43 54.415 3.688 ;
      RECT 54.16 3.438 54.415 3.679 ;
      RECT 54.15 3.443 54.435 3.665 ;
      RECT 54.19 3.433 54.435 3.665 ;
      RECT 54.19 3.436 54.445 3.653 ;
      RECT 54.16 3.438 54.455 3.64 ;
      RECT 54.16 3.442 54.465 3.583 ;
      RECT 54.15 3.447 54.47 3.498 ;
      RECT 54.311 3.415 54.345 3.721 ;
      RECT 53.75 3.518 53.755 3.73 ;
      RECT 53.625 3.515 53.64 3.73 ;
      RECT 53.09 3.545 53.16 3.73 ;
      RECT 52.975 3.545 53.01 3.725 ;
      RECT 54.096 3.847 54.115 4.041 ;
      RECT 54.01 3.802 54.096 4.042 ;
      RECT 54 3.755 54.01 4.044 ;
      RECT 53.995 3.735 54 4.045 ;
      RECT 53.975 3.7 53.995 4.046 ;
      RECT 53.96 3.65 53.975 4.047 ;
      RECT 53.94 3.587 53.96 4.048 ;
      RECT 53.93 3.55 53.94 4.049 ;
      RECT 53.915 3.539 53.93 4.05 ;
      RECT 53.91 3.531 53.915 4.048 ;
      RECT 53.9 3.53 53.91 4.04 ;
      RECT 53.87 3.527 53.9 4.019 ;
      RECT 53.795 3.522 53.87 3.964 ;
      RECT 53.78 3.518 53.795 3.91 ;
      RECT 53.77 3.518 53.78 3.805 ;
      RECT 53.755 3.518 53.77 3.738 ;
      RECT 53.74 3.518 53.75 3.728 ;
      RECT 53.685 3.517 53.74 3.725 ;
      RECT 53.64 3.515 53.685 3.728 ;
      RECT 53.612 3.515 53.625 3.731 ;
      RECT 53.526 3.519 53.612 3.733 ;
      RECT 53.44 3.525 53.526 3.738 ;
      RECT 53.42 3.529 53.44 3.74 ;
      RECT 53.418 3.53 53.42 3.739 ;
      RECT 53.332 3.532 53.418 3.738 ;
      RECT 53.246 3.537 53.332 3.735 ;
      RECT 53.16 3.542 53.246 3.732 ;
      RECT 53.01 3.545 53.09 3.728 ;
      RECT 53.665 10.11 53.84 10.6 ;
      RECT 53.665 7.31 53.835 10.6 ;
      RECT 53.665 9.61 54.075 9.94 ;
      RECT 53.665 8.77 54.075 9.1 ;
      RECT 53.665 7.31 53.84 8.57 ;
      RECT 53.786 4.52 53.835 4.854 ;
      RECT 53.786 4.52 53.84 4.853 ;
      RECT 53.7 4.52 53.84 4.852 ;
      RECT 53.475 4.628 53.845 4.85 ;
      RECT 53.7 4.52 53.87 4.843 ;
      RECT 53.67 4.532 53.875 4.834 ;
      RECT 53.655 4.55 53.88 4.831 ;
      RECT 53.47 4.634 53.88 4.758 ;
      RECT 53.465 4.641 53.88 4.718 ;
      RECT 53.48 4.607 53.88 4.831 ;
      RECT 53.641 4.553 53.845 4.85 ;
      RECT 53.555 4.573 53.88 4.831 ;
      RECT 53.655 4.547 53.875 4.834 ;
      RECT 53.425 3.871 53.615 4.065 ;
      RECT 53.42 3.873 53.615 4.064 ;
      RECT 53.415 3.877 53.63 4.061 ;
      RECT 53.43 3.87 53.63 4.061 ;
      RECT 53.415 3.98 53.635 4.056 ;
      RECT 52.71 4.48 52.801 4.778 ;
      RECT 52.705 4.482 52.88 4.773 ;
      RECT 52.71 4.48 52.88 4.773 ;
      RECT 52.705 4.486 52.9 4.771 ;
      RECT 52.705 4.541 52.94 4.77 ;
      RECT 52.705 4.576 52.955 4.764 ;
      RECT 52.705 4.61 52.965 4.754 ;
      RECT 52.695 4.49 52.9 4.605 ;
      RECT 52.695 4.51 52.915 4.605 ;
      RECT 52.695 4.493 52.905 4.605 ;
      RECT 52.92 3.261 52.925 3.323 ;
      RECT 52.915 3.183 52.92 3.346 ;
      RECT 52.91 3.14 52.915 3.357 ;
      RECT 52.905 3.13 52.91 3.369 ;
      RECT 52.9 3.13 52.905 3.378 ;
      RECT 52.875 3.13 52.9 3.41 ;
      RECT 52.87 3.13 52.875 3.443 ;
      RECT 52.855 3.13 52.87 3.468 ;
      RECT 52.845 3.13 52.855 3.495 ;
      RECT 52.84 3.13 52.845 3.508 ;
      RECT 52.835 3.13 52.84 3.523 ;
      RECT 52.825 3.13 52.835 3.538 ;
      RECT 52.82 3.13 52.825 3.558 ;
      RECT 52.795 3.13 52.82 3.593 ;
      RECT 52.75 3.13 52.795 3.638 ;
      RECT 52.74 3.13 52.75 3.651 ;
      RECT 52.655 3.215 52.74 3.658 ;
      RECT 52.62 3.337 52.655 3.667 ;
      RECT 52.615 3.377 52.62 3.671 ;
      RECT 52.595 3.4 52.615 3.673 ;
      RECT 52.59 3.43 52.595 3.676 ;
      RECT 52.58 3.442 52.59 3.677 ;
      RECT 52.535 3.465 52.58 3.682 ;
      RECT 52.495 3.495 52.535 3.69 ;
      RECT 52.46 3.507 52.495 3.696 ;
      RECT 52.455 3.512 52.46 3.7 ;
      RECT 52.385 3.522 52.455 3.707 ;
      RECT 52.345 3.532 52.385 3.717 ;
      RECT 52.325 3.537 52.345 3.723 ;
      RECT 52.315 3.541 52.325 3.728 ;
      RECT 52.31 3.544 52.315 3.731 ;
      RECT 52.3 3.545 52.31 3.732 ;
      RECT 52.275 3.547 52.3 3.736 ;
      RECT 52.265 3.552 52.275 3.739 ;
      RECT 52.22 3.56 52.265 3.74 ;
      RECT 52.095 3.565 52.22 3.74 ;
      RECT 52.65 3.862 52.67 4.044 ;
      RECT 52.601 3.847 52.65 4.043 ;
      RECT 52.515 3.862 52.67 4.041 ;
      RECT 52.5 3.862 52.67 4.04 ;
      RECT 52.465 3.84 52.635 4.025 ;
      RECT 52.535 4.86 52.55 5.069 ;
      RECT 52.535 4.868 52.555 5.068 ;
      RECT 52.48 4.868 52.555 5.067 ;
      RECT 52.46 4.872 52.56 5.065 ;
      RECT 52.44 4.822 52.48 5.064 ;
      RECT 52.385 4.88 52.565 5.062 ;
      RECT 52.35 4.837 52.48 5.06 ;
      RECT 52.346 4.84 52.535 5.059 ;
      RECT 52.26 4.848 52.535 5.057 ;
      RECT 52.26 4.892 52.57 5.05 ;
      RECT 52.25 4.985 52.57 5.048 ;
      RECT 52.26 4.904 52.575 5.033 ;
      RECT 52.26 4.925 52.59 5.003 ;
      RECT 52.26 4.952 52.595 4.973 ;
      RECT 52.385 4.83 52.48 5.062 ;
      RECT 52.015 3.875 52.02 4.413 ;
      RECT 51.82 4.205 51.825 4.4 ;
      RECT 50.12 3.87 50.135 4.25 ;
      RECT 52.185 3.87 52.19 4.04 ;
      RECT 52.18 3.87 52.185 4.05 ;
      RECT 52.175 3.87 52.18 4.063 ;
      RECT 52.15 3.87 52.175 4.105 ;
      RECT 52.125 3.87 52.15 4.178 ;
      RECT 52.11 3.87 52.125 4.23 ;
      RECT 52.105 3.87 52.11 4.26 ;
      RECT 52.08 3.87 52.105 4.3 ;
      RECT 52.065 3.87 52.08 4.355 ;
      RECT 52.06 3.87 52.065 4.388 ;
      RECT 52.035 3.87 52.06 4.408 ;
      RECT 52.02 3.87 52.035 4.414 ;
      RECT 51.95 3.905 52.015 4.41 ;
      RECT 51.9 3.96 51.95 4.405 ;
      RECT 51.89 3.992 51.9 4.403 ;
      RECT 51.885 4.017 51.89 4.403 ;
      RECT 51.865 4.09 51.885 4.403 ;
      RECT 51.855 4.17 51.865 4.402 ;
      RECT 51.84 4.2 51.855 4.402 ;
      RECT 51.825 4.205 51.84 4.401 ;
      RECT 51.765 4.207 51.82 4.398 ;
      RECT 51.735 4.212 51.765 4.394 ;
      RECT 51.733 4.215 51.735 4.393 ;
      RECT 51.647 4.217 51.733 4.39 ;
      RECT 51.561 4.223 51.647 4.384 ;
      RECT 51.475 4.228 51.561 4.378 ;
      RECT 51.402 4.233 51.475 4.379 ;
      RECT 51.316 4.239 51.402 4.387 ;
      RECT 51.23 4.245 51.316 4.396 ;
      RECT 51.21 4.249 51.23 4.401 ;
      RECT 51.163 4.251 51.21 4.404 ;
      RECT 51.077 4.256 51.163 4.41 ;
      RECT 50.991 4.261 51.077 4.419 ;
      RECT 50.905 4.267 50.991 4.427 ;
      RECT 50.82 4.265 50.905 4.436 ;
      RECT 50.816 4.26 50.82 4.44 ;
      RECT 50.73 4.255 50.816 4.432 ;
      RECT 50.666 4.246 50.73 4.42 ;
      RECT 50.58 4.237 50.666 4.407 ;
      RECT 50.556 4.23 50.58 4.398 ;
      RECT 50.47 4.224 50.556 4.385 ;
      RECT 50.43 4.217 50.47 4.371 ;
      RECT 50.425 4.207 50.43 4.367 ;
      RECT 50.415 4.195 50.425 4.366 ;
      RECT 50.395 4.165 50.415 4.363 ;
      RECT 50.34 4.085 50.395 4.357 ;
      RECT 50.32 4.004 50.34 4.352 ;
      RECT 50.3 3.962 50.32 4.348 ;
      RECT 50.275 3.915 50.3 4.342 ;
      RECT 50.27 3.89 50.275 4.339 ;
      RECT 50.235 3.87 50.27 4.334 ;
      RECT 50.226 3.87 50.235 4.327 ;
      RECT 50.14 3.87 50.226 4.297 ;
      RECT 50.135 3.87 50.14 4.26 ;
      RECT 50.1 3.87 50.12 4.182 ;
      RECT 50.095 3.912 50.1 4.147 ;
      RECT 50.09 3.987 50.095 4.103 ;
      RECT 51.54 3.792 51.715 4.04 ;
      RECT 51.54 3.792 51.72 4.038 ;
      RECT 51.535 3.824 51.72 3.998 ;
      RECT 51.565 3.765 51.735 3.985 ;
      RECT 51.53 3.842 51.735 3.918 ;
      RECT 50.84 3.305 51.01 3.48 ;
      RECT 50.84 3.305 51.182 3.472 ;
      RECT 50.84 3.305 51.265 3.466 ;
      RECT 50.84 3.305 51.3 3.462 ;
      RECT 50.84 3.305 51.32 3.461 ;
      RECT 50.84 3.305 51.406 3.457 ;
      RECT 51.3 3.13 51.47 3.452 ;
      RECT 50.875 3.237 51.5 3.45 ;
      RECT 50.865 3.292 51.505 3.448 ;
      RECT 50.84 3.328 51.515 3.443 ;
      RECT 50.84 3.355 51.52 3.373 ;
      RECT 50.905 3.18 51.48 3.45 ;
      RECT 51.096 3.165 51.48 3.45 ;
      RECT 50.93 3.168 51.48 3.45 ;
      RECT 51.01 3.166 51.096 3.477 ;
      RECT 51.096 3.163 51.475 3.45 ;
      RECT 51.28 3.14 51.475 3.45 ;
      RECT 51.182 3.161 51.475 3.45 ;
      RECT 51.265 3.155 51.28 3.463 ;
      RECT 51.415 4.52 51.42 4.72 ;
      RECT 50.88 4.585 50.925 4.72 ;
      RECT 51.45 4.52 51.47 4.693 ;
      RECT 51.42 4.52 51.45 4.708 ;
      RECT 51.355 4.52 51.415 4.745 ;
      RECT 51.34 4.52 51.355 4.775 ;
      RECT 51.325 4.52 51.34 4.788 ;
      RECT 51.305 4.52 51.325 4.803 ;
      RECT 51.3 4.52 51.305 4.812 ;
      RECT 51.29 4.524 51.3 4.817 ;
      RECT 51.275 4.534 51.29 4.828 ;
      RECT 51.25 4.55 51.275 4.838 ;
      RECT 51.24 4.564 51.25 4.84 ;
      RECT 51.22 4.576 51.24 4.837 ;
      RECT 51.19 4.597 51.22 4.831 ;
      RECT 51.18 4.609 51.19 4.826 ;
      RECT 51.17 4.607 51.18 4.823 ;
      RECT 51.155 4.606 51.17 4.818 ;
      RECT 51.15 4.605 51.155 4.813 ;
      RECT 51.115 4.603 51.15 4.803 ;
      RECT 51.095 4.6 51.115 4.785 ;
      RECT 51.085 4.598 51.095 4.78 ;
      RECT 51.075 4.597 51.085 4.775 ;
      RECT 51.04 4.595 51.075 4.763 ;
      RECT 50.985 4.591 51.04 4.743 ;
      RECT 50.975 4.589 50.985 4.728 ;
      RECT 50.97 4.589 50.975 4.723 ;
      RECT 50.925 4.587 50.97 4.72 ;
      RECT 50.83 4.585 50.88 4.724 ;
      RECT 50.82 4.586 50.83 4.729 ;
      RECT 50.76 4.593 50.82 4.743 ;
      RECT 50.735 4.601 50.76 4.763 ;
      RECT 50.725 4.605 50.735 4.775 ;
      RECT 50.72 4.606 50.725 4.78 ;
      RECT 50.705 4.608 50.72 4.783 ;
      RECT 50.69 4.61 50.705 4.788 ;
      RECT 50.685 4.61 50.69 4.791 ;
      RECT 50.64 4.615 50.685 4.802 ;
      RECT 50.635 4.619 50.64 4.814 ;
      RECT 50.61 4.615 50.635 4.818 ;
      RECT 50.6 4.611 50.61 4.822 ;
      RECT 50.59 4.61 50.6 4.826 ;
      RECT 50.575 4.6 50.59 4.832 ;
      RECT 50.57 4.588 50.575 4.836 ;
      RECT 50.565 4.585 50.57 4.837 ;
      RECT 50.56 4.582 50.565 4.839 ;
      RECT 50.545 4.57 50.56 4.838 ;
      RECT 50.53 4.552 50.545 4.835 ;
      RECT 50.51 4.531 50.53 4.828 ;
      RECT 50.445 4.52 50.51 4.8 ;
      RECT 50.441 4.52 50.445 4.779 ;
      RECT 50.355 4.52 50.441 4.749 ;
      RECT 50.34 4.52 50.355 4.705 ;
      RECT 50.99 4.871 51.005 5.13 ;
      RECT 50.99 4.886 51.01 5.129 ;
      RECT 50.906 4.886 51.01 5.127 ;
      RECT 50.906 4.9 51.015 5.126 ;
      RECT 50.82 4.942 51.02 5.123 ;
      RECT 50.815 4.885 51.005 5.118 ;
      RECT 50.815 4.956 51.025 5.115 ;
      RECT 50.81 4.987 51.025 5.113 ;
      RECT 50.815 4.984 51.04 5.103 ;
      RECT 50.81 5.03 51.055 5.088 ;
      RECT 50.81 5.058 51.06 5.073 ;
      RECT 50.82 4.86 50.99 5.123 ;
      RECT 50.58 3.87 50.75 4.04 ;
      RECT 50.545 3.87 50.75 4.035 ;
      RECT 50.535 3.87 50.75 4.028 ;
      RECT 50.53 3.855 50.7 4.025 ;
      RECT 49.36 4.392 49.625 4.835 ;
      RECT 49.355 4.363 49.57 4.833 ;
      RECT 49.35 4.517 49.63 4.828 ;
      RECT 49.355 4.412 49.63 4.828 ;
      RECT 49.355 4.423 49.64 4.815 ;
      RECT 49.355 4.37 49.6 4.833 ;
      RECT 49.36 4.357 49.57 4.835 ;
      RECT 49.36 4.355 49.52 4.835 ;
      RECT 49.461 4.347 49.52 4.835 ;
      RECT 49.375 4.348 49.52 4.835 ;
      RECT 49.461 4.346 49.51 4.835 ;
      RECT 49.265 3.161 49.44 3.46 ;
      RECT 49.315 3.123 49.44 3.46 ;
      RECT 49.3 3.125 49.526 3.452 ;
      RECT 49.3 3.128 49.565 3.439 ;
      RECT 49.3 3.129 49.575 3.425 ;
      RECT 49.255 3.18 49.575 3.415 ;
      RECT 49.3 3.13 49.58 3.41 ;
      RECT 49.255 3.34 49.585 3.4 ;
      RECT 49.24 3.2 49.58 3.34 ;
      RECT 49.235 3.216 49.58 3.28 ;
      RECT 49.28 3.14 49.58 3.41 ;
      RECT 49.315 3.121 49.401 3.46 ;
      RECT 47.775 7.31 47.945 8.78 ;
      RECT 47.775 7.31 47.95 8.57 ;
      RECT 47.405 9.26 47.875 9.43 ;
      RECT 47.405 8.24 47.575 9.43 ;
      RECT 47.4 3.035 47.57 4.225 ;
      RECT 47.4 3.035 47.87 3.205 ;
      RECT 46.785 3.895 46.96 5.155 ;
      RECT 46.785 3.685 46.955 5.155 ;
      RECT 46.785 7.31 46.955 8.78 ;
      RECT 46.785 7.31 46.96 8.57 ;
      RECT 46.415 3.035 46.585 4.225 ;
      RECT 46.415 3.035 46.885 3.205 ;
      RECT 46.415 9.26 46.885 9.43 ;
      RECT 46.415 8.24 46.585 9.43 ;
      RECT 45.425 4.015 45.6 5.155 ;
      RECT 45.425 1.865 45.595 5.155 ;
      RECT 45.425 1.865 45.6 2.415 ;
      RECT 45.425 10.05 45.6 10.6 ;
      RECT 45.425 7.31 45.595 10.6 ;
      RECT 45.425 7.31 45.6 8.45 ;
      RECT 44.995 3.895 45.17 5.155 ;
      RECT 44.995 2.945 45.165 5.155 ;
      RECT 44.995 7.31 45.165 9.52 ;
      RECT 44.995 7.31 45.17 8.57 ;
      RECT 44.565 3.925 44.735 5.155 ;
      RECT 44.625 2.145 44.795 4.095 ;
      RECT 44.565 1.865 44.735 2.315 ;
      RECT 44.565 10.15 44.735 10.6 ;
      RECT 44.625 8.37 44.795 10.32 ;
      RECT 44.565 7.31 44.735 8.54 ;
      RECT 44.04 3.895 44.215 5.155 ;
      RECT 44.04 1.865 44.21 5.155 ;
      RECT 44.04 3.365 44.45 3.695 ;
      RECT 44.04 2.525 44.45 2.855 ;
      RECT 44.04 1.865 44.215 2.355 ;
      RECT 44.04 10.11 44.215 10.6 ;
      RECT 44.04 7.31 44.21 10.6 ;
      RECT 44.04 9.61 44.45 9.94 ;
      RECT 44.04 8.77 44.45 9.1 ;
      RECT 44.04 7.31 44.215 8.57 ;
      RECT 41.97 4.421 41.975 4.593 ;
      RECT 41.965 4.414 41.97 4.683 ;
      RECT 41.96 4.408 41.965 4.702 ;
      RECT 41.94 4.402 41.96 4.712 ;
      RECT 41.925 4.397 41.94 4.72 ;
      RECT 41.888 4.391 41.925 4.718 ;
      RECT 41.802 4.377 41.888 4.714 ;
      RECT 41.716 4.359 41.802 4.709 ;
      RECT 41.63 4.34 41.716 4.703 ;
      RECT 41.6 4.328 41.63 4.699 ;
      RECT 41.58 4.322 41.6 4.698 ;
      RECT 41.515 4.32 41.58 4.696 ;
      RECT 41.5 4.32 41.515 4.688 ;
      RECT 41.485 4.32 41.5 4.675 ;
      RECT 41.48 4.32 41.485 4.665 ;
      RECT 41.465 4.32 41.48 4.643 ;
      RECT 41.45 4.32 41.465 4.61 ;
      RECT 41.445 4.32 41.45 4.588 ;
      RECT 41.435 4.32 41.445 4.57 ;
      RECT 41.42 4.32 41.435 4.548 ;
      RECT 41.4 4.32 41.42 4.51 ;
      RECT 41.75 3.605 41.785 4.044 ;
      RECT 41.75 3.605 41.79 4.043 ;
      RECT 41.695 3.665 41.79 4.042 ;
      RECT 41.56 3.837 41.79 4.041 ;
      RECT 41.67 3.715 41.79 4.041 ;
      RECT 41.56 3.837 41.815 4.031 ;
      RECT 41.615 3.782 41.895 3.948 ;
      RECT 41.79 3.576 41.795 4.039 ;
      RECT 41.645 3.752 41.935 3.825 ;
      RECT 41.66 3.735 41.79 4.041 ;
      RECT 41.795 3.575 41.965 3.763 ;
      RECT 41.785 3.578 41.965 3.763 ;
      RECT 41.29 3.455 41.46 3.765 ;
      RECT 41.29 3.455 41.465 3.738 ;
      RECT 41.29 3.455 41.47 3.715 ;
      RECT 41.29 3.455 41.48 3.665 ;
      RECT 41.285 3.56 41.48 3.635 ;
      RECT 41.32 3.13 41.49 3.608 ;
      RECT 41.32 3.13 41.505 3.529 ;
      RECT 41.31 3.34 41.505 3.529 ;
      RECT 41.32 3.14 41.515 3.444 ;
      RECT 41.25 3.882 41.255 4.085 ;
      RECT 41.24 3.87 41.25 4.195 ;
      RECT 41.215 3.87 41.24 4.235 ;
      RECT 41.135 3.87 41.215 4.32 ;
      RECT 41.125 3.87 41.135 4.39 ;
      RECT 41.1 3.87 41.125 4.413 ;
      RECT 41.08 3.87 41.1 4.448 ;
      RECT 41.035 3.88 41.08 4.491 ;
      RECT 41.025 3.892 41.035 4.528 ;
      RECT 41.005 3.906 41.025 4.548 ;
      RECT 40.995 3.924 41.005 4.564 ;
      RECT 40.98 3.95 40.995 4.574 ;
      RECT 40.965 3.991 40.98 4.588 ;
      RECT 40.955 4.026 40.965 4.598 ;
      RECT 40.95 4.042 40.955 4.603 ;
      RECT 40.94 4.057 40.95 4.608 ;
      RECT 40.92 4.1 40.94 4.618 ;
      RECT 40.9 4.137 40.92 4.631 ;
      RECT 40.865 4.16 40.9 4.649 ;
      RECT 40.855 4.174 40.865 4.665 ;
      RECT 40.835 4.184 40.855 4.675 ;
      RECT 40.83 4.193 40.835 4.683 ;
      RECT 40.82 4.2 40.83 4.69 ;
      RECT 40.81 4.207 40.82 4.698 ;
      RECT 40.795 4.217 40.81 4.706 ;
      RECT 40.785 4.231 40.795 4.716 ;
      RECT 40.775 4.243 40.785 4.728 ;
      RECT 40.76 4.265 40.775 4.741 ;
      RECT 40.75 4.287 40.76 4.752 ;
      RECT 40.74 4.307 40.75 4.761 ;
      RECT 40.735 4.322 40.74 4.768 ;
      RECT 40.705 4.355 40.735 4.782 ;
      RECT 40.695 4.39 40.705 4.797 ;
      RECT 40.69 4.397 40.695 4.803 ;
      RECT 40.67 4.412 40.69 4.81 ;
      RECT 40.665 4.427 40.67 4.818 ;
      RECT 40.66 4.436 40.665 4.823 ;
      RECT 40.645 4.442 40.66 4.83 ;
      RECT 40.64 4.448 40.645 4.838 ;
      RECT 40.635 4.452 40.64 4.845 ;
      RECT 40.63 4.456 40.635 4.855 ;
      RECT 40.62 4.461 40.63 4.865 ;
      RECT 40.6 4.472 40.62 4.893 ;
      RECT 40.585 4.484 40.6 4.92 ;
      RECT 40.565 4.497 40.585 4.945 ;
      RECT 40.545 4.512 40.565 4.969 ;
      RECT 40.53 4.527 40.545 4.984 ;
      RECT 40.525 4.538 40.53 4.993 ;
      RECT 40.46 4.583 40.525 5.003 ;
      RECT 40.425 4.642 40.46 5.016 ;
      RECT 40.42 4.665 40.425 5.022 ;
      RECT 40.415 4.672 40.42 5.024 ;
      RECT 40.4 4.682 40.415 5.027 ;
      RECT 40.37 4.707 40.4 5.031 ;
      RECT 40.365 4.725 40.37 5.035 ;
      RECT 40.36 4.732 40.365 5.036 ;
      RECT 40.34 4.74 40.36 5.04 ;
      RECT 40.33 4.747 40.34 5.044 ;
      RECT 40.286 4.758 40.33 5.051 ;
      RECT 40.2 4.786 40.286 5.067 ;
      RECT 40.14 4.81 40.2 5.085 ;
      RECT 40.095 4.82 40.14 5.099 ;
      RECT 40.036 4.828 40.095 5.113 ;
      RECT 39.95 4.835 40.036 5.132 ;
      RECT 39.925 4.84 39.95 5.147 ;
      RECT 39.845 4.843 39.925 5.15 ;
      RECT 39.765 4.847 39.845 5.137 ;
      RECT 39.756 4.85 39.765 5.122 ;
      RECT 39.67 4.85 39.756 5.107 ;
      RECT 39.61 4.852 39.67 5.084 ;
      RECT 39.606 4.855 39.61 5.074 ;
      RECT 39.52 4.855 39.606 5.059 ;
      RECT 39.445 4.855 39.52 5.035 ;
      RECT 40.76 3.864 40.77 4.04 ;
      RECT 40.715 3.831 40.76 4.04 ;
      RECT 40.67 3.782 40.715 4.04 ;
      RECT 40.64 3.752 40.67 4.041 ;
      RECT 40.635 3.735 40.64 4.042 ;
      RECT 40.61 3.715 40.635 4.043 ;
      RECT 40.595 3.69 40.61 4.044 ;
      RECT 40.59 3.677 40.595 4.045 ;
      RECT 40.585 3.671 40.59 4.043 ;
      RECT 40.58 3.663 40.585 4.037 ;
      RECT 40.555 3.655 40.58 4.017 ;
      RECT 40.535 3.644 40.555 3.988 ;
      RECT 40.505 3.629 40.535 3.959 ;
      RECT 40.485 3.615 40.505 3.931 ;
      RECT 40.475 3.609 40.485 3.91 ;
      RECT 40.47 3.606 40.475 3.893 ;
      RECT 40.465 3.603 40.47 3.878 ;
      RECT 40.45 3.598 40.465 3.843 ;
      RECT 40.445 3.594 40.45 3.81 ;
      RECT 40.425 3.589 40.445 3.786 ;
      RECT 40.395 3.581 40.425 3.751 ;
      RECT 40.38 3.575 40.395 3.728 ;
      RECT 40.34 3.568 40.38 3.713 ;
      RECT 40.315 3.56 40.34 3.693 ;
      RECT 40.295 3.555 40.315 3.683 ;
      RECT 40.26 3.549 40.295 3.678 ;
      RECT 40.215 3.54 40.26 3.677 ;
      RECT 40.185 3.536 40.215 3.679 ;
      RECT 40.1 3.544 40.185 3.683 ;
      RECT 40.03 3.555 40.1 3.705 ;
      RECT 40.017 3.561 40.03 3.728 ;
      RECT 39.931 3.568 40.017 3.75 ;
      RECT 39.845 3.58 39.931 3.787 ;
      RECT 39.845 3.957 39.855 4.195 ;
      RECT 39.84 3.586 39.845 3.81 ;
      RECT 39.835 3.842 39.845 4.195 ;
      RECT 39.835 3.587 39.84 3.815 ;
      RECT 39.83 3.588 39.835 4.195 ;
      RECT 39.806 3.59 39.83 4.196 ;
      RECT 39.72 3.598 39.806 4.198 ;
      RECT 39.7 3.612 39.72 4.201 ;
      RECT 39.695 3.64 39.7 4.202 ;
      RECT 39.69 3.652 39.695 4.203 ;
      RECT 39.685 3.667 39.69 4.204 ;
      RECT 39.675 3.697 39.685 4.205 ;
      RECT 39.67 3.735 39.675 4.203 ;
      RECT 39.665 3.755 39.67 4.198 ;
      RECT 39.65 3.79 39.665 4.183 ;
      RECT 39.64 3.842 39.65 4.163 ;
      RECT 39.635 3.872 39.64 4.151 ;
      RECT 39.62 3.885 39.635 4.134 ;
      RECT 39.595 3.889 39.62 4.101 ;
      RECT 39.58 3.887 39.595 4.078 ;
      RECT 39.565 3.886 39.58 4.075 ;
      RECT 39.505 3.884 39.565 4.073 ;
      RECT 39.495 3.882 39.505 4.068 ;
      RECT 39.455 3.881 39.495 4.065 ;
      RECT 39.385 3.878 39.455 4.063 ;
      RECT 39.33 3.876 39.385 4.058 ;
      RECT 39.26 3.87 39.33 4.053 ;
      RECT 39.251 3.87 39.26 4.05 ;
      RECT 39.165 3.87 39.251 4.045 ;
      RECT 39.16 3.87 39.165 4.04 ;
      RECT 40.465 3.105 40.64 3.455 ;
      RECT 40.465 3.12 40.65 3.453 ;
      RECT 40.44 3.07 40.585 3.45 ;
      RECT 40.42 3.071 40.585 3.443 ;
      RECT 40.41 3.072 40.595 3.438 ;
      RECT 40.38 3.073 40.595 3.425 ;
      RECT 40.33 3.074 40.595 3.401 ;
      RECT 40.325 3.076 40.595 3.386 ;
      RECT 40.325 3.142 40.655 3.38 ;
      RECT 40.305 3.083 40.61 3.36 ;
      RECT 40.295 3.092 40.62 3.215 ;
      RECT 40.305 3.087 40.62 3.36 ;
      RECT 40.325 3.077 40.61 3.386 ;
      RECT 39.91 4.402 40.08 4.69 ;
      RECT 39.905 4.42 40.09 4.685 ;
      RECT 39.87 4.428 40.155 4.605 ;
      RECT 39.87 4.428 40.241 4.595 ;
      RECT 39.87 4.428 40.295 4.541 ;
      RECT 40.155 4.325 40.325 4.509 ;
      RECT 39.87 4.48 40.33 4.497 ;
      RECT 39.855 4.45 40.325 4.493 ;
      RECT 40.115 4.332 40.155 4.644 ;
      RECT 39.995 4.369 40.325 4.509 ;
      RECT 40.09 4.344 40.115 4.67 ;
      RECT 40.08 4.351 40.325 4.509 ;
      RECT 40.211 3.815 40.28 4.074 ;
      RECT 40.211 3.87 40.285 4.073 ;
      RECT 40.125 3.87 40.285 4.072 ;
      RECT 40.12 3.87 40.29 4.065 ;
      RECT 40.11 3.815 40.28 4.06 ;
      RECT 39.79 10.05 39.965 10.6 ;
      RECT 39.79 7.31 39.96 10.6 ;
      RECT 39.79 7.31 39.965 8.45 ;
      RECT 39.49 3.114 39.665 3.415 ;
      RECT 39.475 3.102 39.49 3.4 ;
      RECT 39.445 3.101 39.475 3.353 ;
      RECT 39.445 3.119 39.67 3.348 ;
      RECT 39.43 3.103 39.49 3.313 ;
      RECT 39.425 3.125 39.68 3.213 ;
      RECT 39.425 3.108 39.576 3.213 ;
      RECT 39.425 3.11 39.58 3.213 ;
      RECT 39.43 3.106 39.576 3.313 ;
      RECT 39.535 4.342 39.54 4.69 ;
      RECT 39.525 4.332 39.535 4.696 ;
      RECT 39.49 4.322 39.525 4.698 ;
      RECT 39.452 4.317 39.49 4.702 ;
      RECT 39.366 4.31 39.452 4.709 ;
      RECT 39.28 4.3 39.366 4.719 ;
      RECT 39.235 4.295 39.28 4.727 ;
      RECT 39.231 4.295 39.235 4.731 ;
      RECT 39.145 4.295 39.231 4.738 ;
      RECT 39.13 4.295 39.145 4.738 ;
      RECT 39.12 4.293 39.13 4.71 ;
      RECT 39.11 4.289 39.12 4.653 ;
      RECT 39.09 4.283 39.11 4.585 ;
      RECT 39.085 4.279 39.09 4.533 ;
      RECT 39.075 4.278 39.085 4.5 ;
      RECT 39.025 4.276 39.075 4.485 ;
      RECT 39 4.274 39.025 4.48 ;
      RECT 38.957 4.272 39 4.476 ;
      RECT 38.871 4.268 38.957 4.464 ;
      RECT 38.785 4.263 38.871 4.448 ;
      RECT 38.755 4.26 38.785 4.435 ;
      RECT 38.73 4.259 38.755 4.423 ;
      RECT 38.725 4.259 38.73 4.413 ;
      RECT 38.685 4.258 38.725 4.405 ;
      RECT 38.67 4.257 38.685 4.398 ;
      RECT 38.62 4.256 38.67 4.39 ;
      RECT 38.618 4.255 38.62 4.385 ;
      RECT 38.532 4.253 38.618 4.385 ;
      RECT 38.446 4.248 38.532 4.385 ;
      RECT 38.36 4.244 38.446 4.385 ;
      RECT 38.311 4.24 38.36 4.383 ;
      RECT 38.225 4.237 38.311 4.378 ;
      RECT 38.202 4.234 38.225 4.374 ;
      RECT 38.116 4.231 38.202 4.369 ;
      RECT 38.03 4.227 38.116 4.36 ;
      RECT 38.005 4.22 38.03 4.355 ;
      RECT 37.945 4.185 38.005 4.352 ;
      RECT 37.925 4.11 37.945 4.349 ;
      RECT 37.92 4.052 37.925 4.348 ;
      RECT 37.895 3.992 37.92 4.347 ;
      RECT 37.82 3.87 37.895 4.343 ;
      RECT 37.81 3.87 37.82 4.335 ;
      RECT 37.795 3.87 37.81 4.325 ;
      RECT 37.78 3.87 37.795 4.295 ;
      RECT 37.765 3.87 37.78 4.24 ;
      RECT 37.75 3.87 37.765 4.178 ;
      RECT 37.725 3.87 37.75 4.103 ;
      RECT 37.72 3.87 37.725 4.053 ;
      RECT 39.36 7.31 39.53 9.52 ;
      RECT 39.36 7.31 39.535 8.57 ;
      RECT 39.065 3.415 39.085 3.724 ;
      RECT 39.051 3.417 39.1 3.721 ;
      RECT 39.051 3.422 39.12 3.712 ;
      RECT 38.965 3.42 39.1 3.706 ;
      RECT 38.965 3.428 39.155 3.689 ;
      RECT 38.93 3.43 39.155 3.688 ;
      RECT 38.9 3.438 39.155 3.679 ;
      RECT 38.89 3.443 39.175 3.665 ;
      RECT 38.93 3.433 39.175 3.665 ;
      RECT 38.93 3.436 39.185 3.653 ;
      RECT 38.9 3.438 39.195 3.64 ;
      RECT 38.9 3.442 39.205 3.583 ;
      RECT 38.89 3.447 39.21 3.498 ;
      RECT 39.051 3.415 39.085 3.721 ;
      RECT 38.49 3.518 38.495 3.73 ;
      RECT 38.365 3.515 38.38 3.73 ;
      RECT 37.83 3.545 37.9 3.73 ;
      RECT 37.715 3.545 37.75 3.725 ;
      RECT 38.836 3.847 38.855 4.041 ;
      RECT 38.75 3.802 38.836 4.042 ;
      RECT 38.74 3.755 38.75 4.044 ;
      RECT 38.735 3.735 38.74 4.045 ;
      RECT 38.715 3.7 38.735 4.046 ;
      RECT 38.7 3.65 38.715 4.047 ;
      RECT 38.68 3.587 38.7 4.048 ;
      RECT 38.67 3.55 38.68 4.049 ;
      RECT 38.655 3.539 38.67 4.05 ;
      RECT 38.65 3.531 38.655 4.048 ;
      RECT 38.64 3.53 38.65 4.04 ;
      RECT 38.61 3.527 38.64 4.019 ;
      RECT 38.535 3.522 38.61 3.964 ;
      RECT 38.52 3.518 38.535 3.91 ;
      RECT 38.51 3.518 38.52 3.805 ;
      RECT 38.495 3.518 38.51 3.738 ;
      RECT 38.48 3.518 38.49 3.728 ;
      RECT 38.425 3.517 38.48 3.725 ;
      RECT 38.38 3.515 38.425 3.728 ;
      RECT 38.352 3.515 38.365 3.731 ;
      RECT 38.266 3.519 38.352 3.733 ;
      RECT 38.18 3.525 38.266 3.738 ;
      RECT 38.16 3.529 38.18 3.74 ;
      RECT 38.158 3.53 38.16 3.739 ;
      RECT 38.072 3.532 38.158 3.738 ;
      RECT 37.986 3.537 38.072 3.735 ;
      RECT 37.9 3.542 37.986 3.732 ;
      RECT 37.75 3.545 37.83 3.728 ;
      RECT 38.405 10.11 38.58 10.6 ;
      RECT 38.405 7.31 38.575 10.6 ;
      RECT 38.405 9.61 38.815 9.94 ;
      RECT 38.405 8.77 38.815 9.1 ;
      RECT 38.405 7.31 38.58 8.57 ;
      RECT 38.526 4.52 38.575 4.854 ;
      RECT 38.526 4.52 38.58 4.853 ;
      RECT 38.44 4.52 38.58 4.852 ;
      RECT 38.215 4.628 38.585 4.85 ;
      RECT 38.44 4.52 38.61 4.843 ;
      RECT 38.41 4.532 38.615 4.834 ;
      RECT 38.395 4.55 38.62 4.831 ;
      RECT 38.21 4.634 38.62 4.758 ;
      RECT 38.205 4.641 38.62 4.718 ;
      RECT 38.22 4.607 38.62 4.831 ;
      RECT 38.381 4.553 38.585 4.85 ;
      RECT 38.295 4.573 38.62 4.831 ;
      RECT 38.395 4.547 38.615 4.834 ;
      RECT 38.165 3.871 38.355 4.065 ;
      RECT 38.16 3.873 38.355 4.064 ;
      RECT 38.155 3.877 38.37 4.061 ;
      RECT 38.17 3.87 38.37 4.061 ;
      RECT 38.155 3.98 38.375 4.056 ;
      RECT 37.45 4.48 37.541 4.778 ;
      RECT 37.445 4.482 37.62 4.773 ;
      RECT 37.45 4.48 37.62 4.773 ;
      RECT 37.445 4.486 37.64 4.771 ;
      RECT 37.445 4.541 37.68 4.77 ;
      RECT 37.445 4.576 37.695 4.764 ;
      RECT 37.445 4.61 37.705 4.754 ;
      RECT 37.435 4.49 37.64 4.605 ;
      RECT 37.435 4.51 37.655 4.605 ;
      RECT 37.435 4.493 37.645 4.605 ;
      RECT 37.66 3.261 37.665 3.323 ;
      RECT 37.655 3.183 37.66 3.346 ;
      RECT 37.65 3.14 37.655 3.357 ;
      RECT 37.645 3.13 37.65 3.369 ;
      RECT 37.64 3.13 37.645 3.378 ;
      RECT 37.615 3.13 37.64 3.41 ;
      RECT 37.61 3.13 37.615 3.443 ;
      RECT 37.595 3.13 37.61 3.468 ;
      RECT 37.585 3.13 37.595 3.495 ;
      RECT 37.58 3.13 37.585 3.508 ;
      RECT 37.575 3.13 37.58 3.523 ;
      RECT 37.565 3.13 37.575 3.538 ;
      RECT 37.56 3.13 37.565 3.558 ;
      RECT 37.535 3.13 37.56 3.593 ;
      RECT 37.49 3.13 37.535 3.638 ;
      RECT 37.48 3.13 37.49 3.651 ;
      RECT 37.395 3.215 37.48 3.658 ;
      RECT 37.36 3.337 37.395 3.667 ;
      RECT 37.355 3.377 37.36 3.671 ;
      RECT 37.335 3.4 37.355 3.673 ;
      RECT 37.33 3.43 37.335 3.676 ;
      RECT 37.32 3.442 37.33 3.677 ;
      RECT 37.275 3.465 37.32 3.682 ;
      RECT 37.235 3.495 37.275 3.69 ;
      RECT 37.2 3.507 37.235 3.696 ;
      RECT 37.195 3.512 37.2 3.7 ;
      RECT 37.125 3.522 37.195 3.707 ;
      RECT 37.085 3.532 37.125 3.717 ;
      RECT 37.065 3.537 37.085 3.723 ;
      RECT 37.055 3.541 37.065 3.728 ;
      RECT 37.05 3.544 37.055 3.731 ;
      RECT 37.04 3.545 37.05 3.732 ;
      RECT 37.015 3.547 37.04 3.736 ;
      RECT 37.005 3.552 37.015 3.739 ;
      RECT 36.96 3.56 37.005 3.74 ;
      RECT 36.835 3.565 36.96 3.74 ;
      RECT 37.39 3.862 37.41 4.044 ;
      RECT 37.341 3.847 37.39 4.043 ;
      RECT 37.255 3.862 37.41 4.041 ;
      RECT 37.24 3.862 37.41 4.04 ;
      RECT 37.205 3.84 37.375 4.025 ;
      RECT 37.275 4.86 37.29 5.069 ;
      RECT 37.275 4.868 37.295 5.068 ;
      RECT 37.22 4.868 37.295 5.067 ;
      RECT 37.2 4.872 37.3 5.065 ;
      RECT 37.18 4.822 37.22 5.064 ;
      RECT 37.125 4.88 37.305 5.062 ;
      RECT 37.09 4.837 37.22 5.06 ;
      RECT 37.086 4.84 37.275 5.059 ;
      RECT 37 4.848 37.275 5.057 ;
      RECT 37 4.892 37.31 5.05 ;
      RECT 36.99 4.985 37.31 5.048 ;
      RECT 37 4.904 37.315 5.033 ;
      RECT 37 4.925 37.33 5.003 ;
      RECT 37 4.952 37.335 4.973 ;
      RECT 37.125 4.83 37.22 5.062 ;
      RECT 36.755 3.875 36.76 4.413 ;
      RECT 36.56 4.205 36.565 4.4 ;
      RECT 34.86 3.87 34.875 4.25 ;
      RECT 36.925 3.87 36.93 4.04 ;
      RECT 36.92 3.87 36.925 4.05 ;
      RECT 36.915 3.87 36.92 4.063 ;
      RECT 36.89 3.87 36.915 4.105 ;
      RECT 36.865 3.87 36.89 4.178 ;
      RECT 36.85 3.87 36.865 4.23 ;
      RECT 36.845 3.87 36.85 4.26 ;
      RECT 36.82 3.87 36.845 4.3 ;
      RECT 36.805 3.87 36.82 4.355 ;
      RECT 36.8 3.87 36.805 4.388 ;
      RECT 36.775 3.87 36.8 4.408 ;
      RECT 36.76 3.87 36.775 4.414 ;
      RECT 36.69 3.905 36.755 4.41 ;
      RECT 36.64 3.96 36.69 4.405 ;
      RECT 36.63 3.992 36.64 4.403 ;
      RECT 36.625 4.017 36.63 4.403 ;
      RECT 36.605 4.09 36.625 4.403 ;
      RECT 36.595 4.17 36.605 4.402 ;
      RECT 36.58 4.2 36.595 4.402 ;
      RECT 36.565 4.205 36.58 4.401 ;
      RECT 36.505 4.207 36.56 4.398 ;
      RECT 36.475 4.212 36.505 4.394 ;
      RECT 36.473 4.215 36.475 4.393 ;
      RECT 36.387 4.217 36.473 4.39 ;
      RECT 36.301 4.223 36.387 4.384 ;
      RECT 36.215 4.228 36.301 4.378 ;
      RECT 36.142 4.233 36.215 4.379 ;
      RECT 36.056 4.239 36.142 4.387 ;
      RECT 35.97 4.245 36.056 4.396 ;
      RECT 35.95 4.249 35.97 4.401 ;
      RECT 35.903 4.251 35.95 4.404 ;
      RECT 35.817 4.256 35.903 4.41 ;
      RECT 35.731 4.261 35.817 4.419 ;
      RECT 35.645 4.267 35.731 4.427 ;
      RECT 35.56 4.265 35.645 4.436 ;
      RECT 35.556 4.26 35.56 4.44 ;
      RECT 35.47 4.255 35.556 4.432 ;
      RECT 35.406 4.246 35.47 4.42 ;
      RECT 35.32 4.237 35.406 4.407 ;
      RECT 35.296 4.23 35.32 4.398 ;
      RECT 35.21 4.224 35.296 4.385 ;
      RECT 35.17 4.217 35.21 4.371 ;
      RECT 35.165 4.207 35.17 4.367 ;
      RECT 35.155 4.195 35.165 4.366 ;
      RECT 35.135 4.165 35.155 4.363 ;
      RECT 35.08 4.085 35.135 4.357 ;
      RECT 35.06 4.004 35.08 4.352 ;
      RECT 35.04 3.962 35.06 4.348 ;
      RECT 35.015 3.915 35.04 4.342 ;
      RECT 35.01 3.89 35.015 4.339 ;
      RECT 34.975 3.87 35.01 4.334 ;
      RECT 34.966 3.87 34.975 4.327 ;
      RECT 34.88 3.87 34.966 4.297 ;
      RECT 34.875 3.87 34.88 4.26 ;
      RECT 34.84 3.87 34.86 4.182 ;
      RECT 34.835 3.912 34.84 4.147 ;
      RECT 34.83 3.987 34.835 4.103 ;
      RECT 36.28 3.792 36.455 4.04 ;
      RECT 36.28 3.792 36.46 4.038 ;
      RECT 36.275 3.824 36.46 3.998 ;
      RECT 36.305 3.765 36.475 3.985 ;
      RECT 36.27 3.842 36.475 3.918 ;
      RECT 35.58 3.305 35.75 3.48 ;
      RECT 35.58 3.305 35.922 3.472 ;
      RECT 35.58 3.305 36.005 3.466 ;
      RECT 35.58 3.305 36.04 3.462 ;
      RECT 35.58 3.305 36.06 3.461 ;
      RECT 35.58 3.305 36.146 3.457 ;
      RECT 36.04 3.13 36.21 3.452 ;
      RECT 35.615 3.237 36.24 3.45 ;
      RECT 35.605 3.292 36.245 3.448 ;
      RECT 35.58 3.328 36.255 3.443 ;
      RECT 35.58 3.355 36.26 3.373 ;
      RECT 35.645 3.18 36.22 3.45 ;
      RECT 35.836 3.165 36.22 3.45 ;
      RECT 35.67 3.168 36.22 3.45 ;
      RECT 35.75 3.166 35.836 3.477 ;
      RECT 35.836 3.163 36.215 3.45 ;
      RECT 36.02 3.14 36.215 3.45 ;
      RECT 35.922 3.161 36.215 3.45 ;
      RECT 36.005 3.155 36.02 3.463 ;
      RECT 36.155 4.52 36.16 4.72 ;
      RECT 35.62 4.585 35.665 4.72 ;
      RECT 36.19 4.52 36.21 4.693 ;
      RECT 36.16 4.52 36.19 4.708 ;
      RECT 36.095 4.52 36.155 4.745 ;
      RECT 36.08 4.52 36.095 4.775 ;
      RECT 36.065 4.52 36.08 4.788 ;
      RECT 36.045 4.52 36.065 4.803 ;
      RECT 36.04 4.52 36.045 4.812 ;
      RECT 36.03 4.524 36.04 4.817 ;
      RECT 36.015 4.534 36.03 4.828 ;
      RECT 35.99 4.55 36.015 4.838 ;
      RECT 35.98 4.564 35.99 4.84 ;
      RECT 35.96 4.576 35.98 4.837 ;
      RECT 35.93 4.597 35.96 4.831 ;
      RECT 35.92 4.609 35.93 4.826 ;
      RECT 35.91 4.607 35.92 4.823 ;
      RECT 35.895 4.606 35.91 4.818 ;
      RECT 35.89 4.605 35.895 4.813 ;
      RECT 35.855 4.603 35.89 4.803 ;
      RECT 35.835 4.6 35.855 4.785 ;
      RECT 35.825 4.598 35.835 4.78 ;
      RECT 35.815 4.597 35.825 4.775 ;
      RECT 35.78 4.595 35.815 4.763 ;
      RECT 35.725 4.591 35.78 4.743 ;
      RECT 35.715 4.589 35.725 4.728 ;
      RECT 35.71 4.589 35.715 4.723 ;
      RECT 35.665 4.587 35.71 4.72 ;
      RECT 35.57 4.585 35.62 4.724 ;
      RECT 35.56 4.586 35.57 4.729 ;
      RECT 35.5 4.593 35.56 4.743 ;
      RECT 35.475 4.601 35.5 4.763 ;
      RECT 35.465 4.605 35.475 4.775 ;
      RECT 35.46 4.606 35.465 4.78 ;
      RECT 35.445 4.608 35.46 4.783 ;
      RECT 35.43 4.61 35.445 4.788 ;
      RECT 35.425 4.61 35.43 4.791 ;
      RECT 35.38 4.615 35.425 4.802 ;
      RECT 35.375 4.619 35.38 4.814 ;
      RECT 35.35 4.615 35.375 4.818 ;
      RECT 35.34 4.611 35.35 4.822 ;
      RECT 35.33 4.61 35.34 4.826 ;
      RECT 35.315 4.6 35.33 4.832 ;
      RECT 35.31 4.588 35.315 4.836 ;
      RECT 35.305 4.585 35.31 4.837 ;
      RECT 35.3 4.582 35.305 4.839 ;
      RECT 35.285 4.57 35.3 4.838 ;
      RECT 35.27 4.552 35.285 4.835 ;
      RECT 35.25 4.531 35.27 4.828 ;
      RECT 35.185 4.52 35.25 4.8 ;
      RECT 35.181 4.52 35.185 4.779 ;
      RECT 35.095 4.52 35.181 4.749 ;
      RECT 35.08 4.52 35.095 4.705 ;
      RECT 35.73 4.871 35.745 5.13 ;
      RECT 35.73 4.886 35.75 5.129 ;
      RECT 35.646 4.886 35.75 5.127 ;
      RECT 35.646 4.9 35.755 5.126 ;
      RECT 35.56 4.942 35.76 5.123 ;
      RECT 35.555 4.885 35.745 5.118 ;
      RECT 35.555 4.956 35.765 5.115 ;
      RECT 35.55 4.987 35.765 5.113 ;
      RECT 35.555 4.984 35.78 5.103 ;
      RECT 35.55 5.03 35.795 5.088 ;
      RECT 35.55 5.058 35.8 5.073 ;
      RECT 35.56 4.86 35.73 5.123 ;
      RECT 35.32 3.87 35.49 4.04 ;
      RECT 35.285 3.87 35.49 4.035 ;
      RECT 35.275 3.87 35.49 4.028 ;
      RECT 35.27 3.855 35.44 4.025 ;
      RECT 34.1 4.392 34.365 4.835 ;
      RECT 34.095 4.363 34.31 4.833 ;
      RECT 34.09 4.517 34.37 4.828 ;
      RECT 34.095 4.412 34.37 4.828 ;
      RECT 34.095 4.423 34.38 4.815 ;
      RECT 34.095 4.37 34.34 4.833 ;
      RECT 34.1 4.357 34.31 4.835 ;
      RECT 34.1 4.355 34.26 4.835 ;
      RECT 34.201 4.347 34.26 4.835 ;
      RECT 34.115 4.348 34.26 4.835 ;
      RECT 34.201 4.346 34.25 4.835 ;
      RECT 34.005 3.161 34.18 3.46 ;
      RECT 34.055 3.123 34.18 3.46 ;
      RECT 34.04 3.125 34.266 3.452 ;
      RECT 34.04 3.128 34.305 3.439 ;
      RECT 34.04 3.129 34.315 3.425 ;
      RECT 33.995 3.18 34.315 3.415 ;
      RECT 34.04 3.13 34.32 3.41 ;
      RECT 33.995 3.34 34.325 3.4 ;
      RECT 33.98 3.2 34.32 3.34 ;
      RECT 33.975 3.216 34.32 3.28 ;
      RECT 34.02 3.14 34.32 3.41 ;
      RECT 34.055 3.121 34.141 3.46 ;
      RECT 32.515 7.31 32.685 8.78 ;
      RECT 32.515 7.31 32.69 8.57 ;
      RECT 32.145 9.26 32.615 9.43 ;
      RECT 32.145 8.24 32.315 9.43 ;
      RECT 32.14 3.035 32.31 4.225 ;
      RECT 32.14 3.035 32.61 3.205 ;
      RECT 31.525 3.895 31.7 5.155 ;
      RECT 31.525 3.685 31.695 5.155 ;
      RECT 31.525 7.31 31.695 8.78 ;
      RECT 31.525 7.31 31.7 8.57 ;
      RECT 31.155 3.035 31.325 4.225 ;
      RECT 31.155 3.035 31.625 3.205 ;
      RECT 31.155 9.26 31.625 9.43 ;
      RECT 31.155 8.24 31.325 9.43 ;
      RECT 30.165 4.015 30.34 5.155 ;
      RECT 30.165 1.865 30.335 5.155 ;
      RECT 30.165 1.865 30.34 2.415 ;
      RECT 30.165 10.05 30.34 10.6 ;
      RECT 30.165 7.31 30.335 10.6 ;
      RECT 30.165 7.31 30.34 8.45 ;
      RECT 29.735 3.895 29.91 5.155 ;
      RECT 29.735 2.945 29.905 5.155 ;
      RECT 29.735 7.31 29.905 9.52 ;
      RECT 29.735 7.31 29.91 8.57 ;
      RECT 29.305 3.925 29.475 5.155 ;
      RECT 29.365 2.145 29.535 4.095 ;
      RECT 29.305 1.865 29.475 2.315 ;
      RECT 29.305 10.15 29.475 10.6 ;
      RECT 29.365 8.37 29.535 10.32 ;
      RECT 29.305 7.31 29.475 8.54 ;
      RECT 28.78 3.895 28.955 5.155 ;
      RECT 28.78 1.865 28.95 5.155 ;
      RECT 28.78 3.365 29.19 3.695 ;
      RECT 28.78 2.525 29.19 2.855 ;
      RECT 28.78 1.865 28.955 2.355 ;
      RECT 28.78 10.11 28.955 10.6 ;
      RECT 28.78 7.31 28.95 10.6 ;
      RECT 28.78 9.61 29.19 9.94 ;
      RECT 28.78 8.77 29.19 9.1 ;
      RECT 28.78 7.31 28.955 8.57 ;
      RECT 26.71 4.421 26.715 4.593 ;
      RECT 26.705 4.414 26.71 4.683 ;
      RECT 26.7 4.408 26.705 4.702 ;
      RECT 26.68 4.402 26.7 4.712 ;
      RECT 26.665 4.397 26.68 4.72 ;
      RECT 26.628 4.391 26.665 4.718 ;
      RECT 26.542 4.377 26.628 4.714 ;
      RECT 26.456 4.359 26.542 4.709 ;
      RECT 26.37 4.34 26.456 4.703 ;
      RECT 26.34 4.328 26.37 4.699 ;
      RECT 26.32 4.322 26.34 4.698 ;
      RECT 26.255 4.32 26.32 4.696 ;
      RECT 26.24 4.32 26.255 4.688 ;
      RECT 26.225 4.32 26.24 4.675 ;
      RECT 26.22 4.32 26.225 4.665 ;
      RECT 26.205 4.32 26.22 4.643 ;
      RECT 26.19 4.32 26.205 4.61 ;
      RECT 26.185 4.32 26.19 4.588 ;
      RECT 26.175 4.32 26.185 4.57 ;
      RECT 26.16 4.32 26.175 4.548 ;
      RECT 26.14 4.32 26.16 4.51 ;
      RECT 26.49 3.605 26.525 4.044 ;
      RECT 26.49 3.605 26.53 4.043 ;
      RECT 26.435 3.665 26.53 4.042 ;
      RECT 26.3 3.837 26.53 4.041 ;
      RECT 26.41 3.715 26.53 4.041 ;
      RECT 26.3 3.837 26.555 4.031 ;
      RECT 26.355 3.782 26.635 3.948 ;
      RECT 26.53 3.576 26.535 4.039 ;
      RECT 26.385 3.752 26.675 3.825 ;
      RECT 26.4 3.735 26.53 4.041 ;
      RECT 26.535 3.575 26.705 3.763 ;
      RECT 26.525 3.578 26.705 3.763 ;
      RECT 26.03 3.455 26.2 3.765 ;
      RECT 26.03 3.455 26.205 3.738 ;
      RECT 26.03 3.455 26.21 3.715 ;
      RECT 26.03 3.455 26.22 3.665 ;
      RECT 26.025 3.56 26.22 3.635 ;
      RECT 26.06 3.13 26.23 3.608 ;
      RECT 26.06 3.13 26.245 3.529 ;
      RECT 26.05 3.34 26.245 3.529 ;
      RECT 26.06 3.14 26.255 3.444 ;
      RECT 25.99 3.882 25.995 4.085 ;
      RECT 25.98 3.87 25.99 4.195 ;
      RECT 25.955 3.87 25.98 4.235 ;
      RECT 25.875 3.87 25.955 4.32 ;
      RECT 25.865 3.87 25.875 4.39 ;
      RECT 25.84 3.87 25.865 4.413 ;
      RECT 25.82 3.87 25.84 4.448 ;
      RECT 25.775 3.88 25.82 4.491 ;
      RECT 25.765 3.892 25.775 4.528 ;
      RECT 25.745 3.906 25.765 4.548 ;
      RECT 25.735 3.924 25.745 4.564 ;
      RECT 25.72 3.95 25.735 4.574 ;
      RECT 25.705 3.991 25.72 4.588 ;
      RECT 25.695 4.026 25.705 4.598 ;
      RECT 25.69 4.042 25.695 4.603 ;
      RECT 25.68 4.057 25.69 4.608 ;
      RECT 25.66 4.1 25.68 4.618 ;
      RECT 25.64 4.137 25.66 4.631 ;
      RECT 25.605 4.16 25.64 4.649 ;
      RECT 25.595 4.174 25.605 4.665 ;
      RECT 25.575 4.184 25.595 4.675 ;
      RECT 25.57 4.193 25.575 4.683 ;
      RECT 25.56 4.2 25.57 4.69 ;
      RECT 25.55 4.207 25.56 4.698 ;
      RECT 25.535 4.217 25.55 4.706 ;
      RECT 25.525 4.231 25.535 4.716 ;
      RECT 25.515 4.243 25.525 4.728 ;
      RECT 25.5 4.265 25.515 4.741 ;
      RECT 25.49 4.287 25.5 4.752 ;
      RECT 25.48 4.307 25.49 4.761 ;
      RECT 25.475 4.322 25.48 4.768 ;
      RECT 25.445 4.355 25.475 4.782 ;
      RECT 25.435 4.39 25.445 4.797 ;
      RECT 25.43 4.397 25.435 4.803 ;
      RECT 25.41 4.412 25.43 4.81 ;
      RECT 25.405 4.427 25.41 4.818 ;
      RECT 25.4 4.436 25.405 4.823 ;
      RECT 25.385 4.442 25.4 4.83 ;
      RECT 25.38 4.448 25.385 4.838 ;
      RECT 25.375 4.452 25.38 4.845 ;
      RECT 25.37 4.456 25.375 4.855 ;
      RECT 25.36 4.461 25.37 4.865 ;
      RECT 25.34 4.472 25.36 4.893 ;
      RECT 25.325 4.484 25.34 4.92 ;
      RECT 25.305 4.497 25.325 4.945 ;
      RECT 25.285 4.512 25.305 4.969 ;
      RECT 25.27 4.527 25.285 4.984 ;
      RECT 25.265 4.538 25.27 4.993 ;
      RECT 25.2 4.583 25.265 5.003 ;
      RECT 25.165 4.642 25.2 5.016 ;
      RECT 25.16 4.665 25.165 5.022 ;
      RECT 25.155 4.672 25.16 5.024 ;
      RECT 25.14 4.682 25.155 5.027 ;
      RECT 25.11 4.707 25.14 5.031 ;
      RECT 25.105 4.725 25.11 5.035 ;
      RECT 25.1 4.732 25.105 5.036 ;
      RECT 25.08 4.74 25.1 5.04 ;
      RECT 25.07 4.747 25.08 5.044 ;
      RECT 25.026 4.758 25.07 5.051 ;
      RECT 24.94 4.786 25.026 5.067 ;
      RECT 24.88 4.81 24.94 5.085 ;
      RECT 24.835 4.82 24.88 5.099 ;
      RECT 24.776 4.828 24.835 5.113 ;
      RECT 24.69 4.835 24.776 5.132 ;
      RECT 24.665 4.84 24.69 5.147 ;
      RECT 24.585 4.843 24.665 5.15 ;
      RECT 24.505 4.847 24.585 5.137 ;
      RECT 24.496 4.85 24.505 5.122 ;
      RECT 24.41 4.85 24.496 5.107 ;
      RECT 24.35 4.852 24.41 5.084 ;
      RECT 24.346 4.855 24.35 5.074 ;
      RECT 24.26 4.855 24.346 5.059 ;
      RECT 24.185 4.855 24.26 5.035 ;
      RECT 25.5 3.864 25.51 4.04 ;
      RECT 25.455 3.831 25.5 4.04 ;
      RECT 25.41 3.782 25.455 4.04 ;
      RECT 25.38 3.752 25.41 4.041 ;
      RECT 25.375 3.735 25.38 4.042 ;
      RECT 25.35 3.715 25.375 4.043 ;
      RECT 25.335 3.69 25.35 4.044 ;
      RECT 25.33 3.677 25.335 4.045 ;
      RECT 25.325 3.671 25.33 4.043 ;
      RECT 25.32 3.663 25.325 4.037 ;
      RECT 25.295 3.655 25.32 4.017 ;
      RECT 25.275 3.644 25.295 3.988 ;
      RECT 25.245 3.629 25.275 3.959 ;
      RECT 25.225 3.615 25.245 3.931 ;
      RECT 25.215 3.609 25.225 3.91 ;
      RECT 25.21 3.606 25.215 3.893 ;
      RECT 25.205 3.603 25.21 3.878 ;
      RECT 25.19 3.598 25.205 3.843 ;
      RECT 25.185 3.594 25.19 3.81 ;
      RECT 25.165 3.589 25.185 3.786 ;
      RECT 25.135 3.581 25.165 3.751 ;
      RECT 25.12 3.575 25.135 3.728 ;
      RECT 25.08 3.568 25.12 3.713 ;
      RECT 25.055 3.56 25.08 3.693 ;
      RECT 25.035 3.555 25.055 3.683 ;
      RECT 25 3.549 25.035 3.678 ;
      RECT 24.955 3.54 25 3.677 ;
      RECT 24.925 3.536 24.955 3.679 ;
      RECT 24.84 3.544 24.925 3.683 ;
      RECT 24.77 3.555 24.84 3.705 ;
      RECT 24.757 3.561 24.77 3.728 ;
      RECT 24.671 3.568 24.757 3.75 ;
      RECT 24.585 3.58 24.671 3.787 ;
      RECT 24.585 3.957 24.595 4.195 ;
      RECT 24.58 3.586 24.585 3.81 ;
      RECT 24.575 3.842 24.585 4.195 ;
      RECT 24.575 3.587 24.58 3.815 ;
      RECT 24.57 3.588 24.575 4.195 ;
      RECT 24.546 3.59 24.57 4.196 ;
      RECT 24.46 3.598 24.546 4.198 ;
      RECT 24.44 3.612 24.46 4.201 ;
      RECT 24.435 3.64 24.44 4.202 ;
      RECT 24.43 3.652 24.435 4.203 ;
      RECT 24.425 3.667 24.43 4.204 ;
      RECT 24.415 3.697 24.425 4.205 ;
      RECT 24.41 3.735 24.415 4.203 ;
      RECT 24.405 3.755 24.41 4.198 ;
      RECT 24.39 3.79 24.405 4.183 ;
      RECT 24.38 3.842 24.39 4.163 ;
      RECT 24.375 3.872 24.38 4.151 ;
      RECT 24.36 3.885 24.375 4.134 ;
      RECT 24.335 3.889 24.36 4.101 ;
      RECT 24.32 3.887 24.335 4.078 ;
      RECT 24.305 3.886 24.32 4.075 ;
      RECT 24.245 3.884 24.305 4.073 ;
      RECT 24.235 3.882 24.245 4.068 ;
      RECT 24.195 3.881 24.235 4.065 ;
      RECT 24.125 3.878 24.195 4.063 ;
      RECT 24.07 3.876 24.125 4.058 ;
      RECT 24 3.87 24.07 4.053 ;
      RECT 23.991 3.87 24 4.05 ;
      RECT 23.905 3.87 23.991 4.045 ;
      RECT 23.9 3.87 23.905 4.04 ;
      RECT 25.205 3.105 25.38 3.455 ;
      RECT 25.205 3.12 25.39 3.453 ;
      RECT 25.18 3.07 25.325 3.45 ;
      RECT 25.16 3.071 25.325 3.443 ;
      RECT 25.15 3.072 25.335 3.438 ;
      RECT 25.12 3.073 25.335 3.425 ;
      RECT 25.07 3.074 25.335 3.401 ;
      RECT 25.065 3.076 25.335 3.386 ;
      RECT 25.065 3.142 25.395 3.38 ;
      RECT 25.045 3.083 25.35 3.36 ;
      RECT 25.035 3.092 25.36 3.215 ;
      RECT 25.045 3.087 25.36 3.36 ;
      RECT 25.065 3.077 25.35 3.386 ;
      RECT 24.65 4.402 24.82 4.69 ;
      RECT 24.645 4.42 24.83 4.685 ;
      RECT 24.61 4.428 24.895 4.605 ;
      RECT 24.61 4.428 24.981 4.595 ;
      RECT 24.61 4.428 25.035 4.541 ;
      RECT 24.895 4.325 25.065 4.509 ;
      RECT 24.61 4.48 25.07 4.497 ;
      RECT 24.595 4.45 25.065 4.493 ;
      RECT 24.855 4.332 24.895 4.644 ;
      RECT 24.735 4.369 25.065 4.509 ;
      RECT 24.83 4.344 24.855 4.67 ;
      RECT 24.82 4.351 25.065 4.509 ;
      RECT 24.951 3.815 25.02 4.074 ;
      RECT 24.951 3.87 25.025 4.073 ;
      RECT 24.865 3.87 25.025 4.072 ;
      RECT 24.86 3.87 25.03 4.065 ;
      RECT 24.85 3.815 25.02 4.06 ;
      RECT 24.53 10.05 24.705 10.6 ;
      RECT 24.53 7.31 24.7 10.6 ;
      RECT 24.53 7.31 24.705 8.45 ;
      RECT 24.23 3.114 24.405 3.415 ;
      RECT 24.215 3.102 24.23 3.4 ;
      RECT 24.185 3.101 24.215 3.353 ;
      RECT 24.185 3.119 24.41 3.348 ;
      RECT 24.17 3.103 24.23 3.313 ;
      RECT 24.165 3.125 24.42 3.213 ;
      RECT 24.165 3.108 24.316 3.213 ;
      RECT 24.165 3.11 24.32 3.213 ;
      RECT 24.17 3.106 24.316 3.313 ;
      RECT 24.275 4.342 24.28 4.69 ;
      RECT 24.265 4.332 24.275 4.696 ;
      RECT 24.23 4.322 24.265 4.698 ;
      RECT 24.192 4.317 24.23 4.702 ;
      RECT 24.106 4.31 24.192 4.709 ;
      RECT 24.02 4.3 24.106 4.719 ;
      RECT 23.975 4.295 24.02 4.727 ;
      RECT 23.971 4.295 23.975 4.731 ;
      RECT 23.885 4.295 23.971 4.738 ;
      RECT 23.87 4.295 23.885 4.738 ;
      RECT 23.86 4.293 23.87 4.71 ;
      RECT 23.85 4.289 23.86 4.653 ;
      RECT 23.83 4.283 23.85 4.585 ;
      RECT 23.825 4.279 23.83 4.533 ;
      RECT 23.815 4.278 23.825 4.5 ;
      RECT 23.765 4.276 23.815 4.485 ;
      RECT 23.74 4.274 23.765 4.48 ;
      RECT 23.697 4.272 23.74 4.476 ;
      RECT 23.611 4.268 23.697 4.464 ;
      RECT 23.525 4.263 23.611 4.448 ;
      RECT 23.495 4.26 23.525 4.435 ;
      RECT 23.47 4.259 23.495 4.423 ;
      RECT 23.465 4.259 23.47 4.413 ;
      RECT 23.425 4.258 23.465 4.405 ;
      RECT 23.41 4.257 23.425 4.398 ;
      RECT 23.36 4.256 23.41 4.39 ;
      RECT 23.358 4.255 23.36 4.385 ;
      RECT 23.272 4.253 23.358 4.385 ;
      RECT 23.186 4.248 23.272 4.385 ;
      RECT 23.1 4.244 23.186 4.385 ;
      RECT 23.051 4.24 23.1 4.383 ;
      RECT 22.965 4.237 23.051 4.378 ;
      RECT 22.942 4.234 22.965 4.374 ;
      RECT 22.856 4.231 22.942 4.369 ;
      RECT 22.77 4.227 22.856 4.36 ;
      RECT 22.745 4.22 22.77 4.355 ;
      RECT 22.685 4.185 22.745 4.352 ;
      RECT 22.665 4.11 22.685 4.349 ;
      RECT 22.66 4.052 22.665 4.348 ;
      RECT 22.635 3.992 22.66 4.347 ;
      RECT 22.56 3.87 22.635 4.343 ;
      RECT 22.55 3.87 22.56 4.335 ;
      RECT 22.535 3.87 22.55 4.325 ;
      RECT 22.52 3.87 22.535 4.295 ;
      RECT 22.505 3.87 22.52 4.24 ;
      RECT 22.49 3.87 22.505 4.178 ;
      RECT 22.465 3.87 22.49 4.103 ;
      RECT 22.46 3.87 22.465 4.053 ;
      RECT 24.1 7.31 24.27 9.52 ;
      RECT 24.1 7.31 24.275 8.57 ;
      RECT 23.805 3.415 23.825 3.724 ;
      RECT 23.791 3.417 23.84 3.721 ;
      RECT 23.791 3.422 23.86 3.712 ;
      RECT 23.705 3.42 23.84 3.706 ;
      RECT 23.705 3.428 23.895 3.689 ;
      RECT 23.67 3.43 23.895 3.688 ;
      RECT 23.64 3.438 23.895 3.679 ;
      RECT 23.63 3.443 23.915 3.665 ;
      RECT 23.67 3.433 23.915 3.665 ;
      RECT 23.67 3.436 23.925 3.653 ;
      RECT 23.64 3.438 23.935 3.64 ;
      RECT 23.64 3.442 23.945 3.583 ;
      RECT 23.63 3.447 23.95 3.498 ;
      RECT 23.791 3.415 23.825 3.721 ;
      RECT 23.23 3.518 23.235 3.73 ;
      RECT 23.105 3.515 23.12 3.73 ;
      RECT 22.57 3.545 22.64 3.73 ;
      RECT 22.455 3.545 22.49 3.725 ;
      RECT 23.576 3.847 23.595 4.041 ;
      RECT 23.49 3.802 23.576 4.042 ;
      RECT 23.48 3.755 23.49 4.044 ;
      RECT 23.475 3.735 23.48 4.045 ;
      RECT 23.455 3.7 23.475 4.046 ;
      RECT 23.44 3.65 23.455 4.047 ;
      RECT 23.42 3.587 23.44 4.048 ;
      RECT 23.41 3.55 23.42 4.049 ;
      RECT 23.395 3.539 23.41 4.05 ;
      RECT 23.39 3.531 23.395 4.048 ;
      RECT 23.38 3.53 23.39 4.04 ;
      RECT 23.35 3.527 23.38 4.019 ;
      RECT 23.275 3.522 23.35 3.964 ;
      RECT 23.26 3.518 23.275 3.91 ;
      RECT 23.25 3.518 23.26 3.805 ;
      RECT 23.235 3.518 23.25 3.738 ;
      RECT 23.22 3.518 23.23 3.728 ;
      RECT 23.165 3.517 23.22 3.725 ;
      RECT 23.12 3.515 23.165 3.728 ;
      RECT 23.092 3.515 23.105 3.731 ;
      RECT 23.006 3.519 23.092 3.733 ;
      RECT 22.92 3.525 23.006 3.738 ;
      RECT 22.9 3.529 22.92 3.74 ;
      RECT 22.898 3.53 22.9 3.739 ;
      RECT 22.812 3.532 22.898 3.738 ;
      RECT 22.726 3.537 22.812 3.735 ;
      RECT 22.64 3.542 22.726 3.732 ;
      RECT 22.49 3.545 22.57 3.728 ;
      RECT 23.145 10.11 23.32 10.6 ;
      RECT 23.145 7.31 23.315 10.6 ;
      RECT 23.145 9.61 23.555 9.94 ;
      RECT 23.145 8.77 23.555 9.1 ;
      RECT 23.145 7.31 23.32 8.57 ;
      RECT 23.266 4.52 23.315 4.854 ;
      RECT 23.266 4.52 23.32 4.853 ;
      RECT 23.18 4.52 23.32 4.852 ;
      RECT 22.955 4.628 23.325 4.85 ;
      RECT 23.18 4.52 23.35 4.843 ;
      RECT 23.15 4.532 23.355 4.834 ;
      RECT 23.135 4.55 23.36 4.831 ;
      RECT 22.95 4.634 23.36 4.758 ;
      RECT 22.945 4.641 23.36 4.718 ;
      RECT 22.96 4.607 23.36 4.831 ;
      RECT 23.121 4.553 23.325 4.85 ;
      RECT 23.035 4.573 23.36 4.831 ;
      RECT 23.135 4.547 23.355 4.834 ;
      RECT 22.905 3.871 23.095 4.065 ;
      RECT 22.9 3.873 23.095 4.064 ;
      RECT 22.895 3.877 23.11 4.061 ;
      RECT 22.91 3.87 23.11 4.061 ;
      RECT 22.895 3.98 23.115 4.056 ;
      RECT 22.19 4.48 22.281 4.778 ;
      RECT 22.185 4.482 22.36 4.773 ;
      RECT 22.19 4.48 22.36 4.773 ;
      RECT 22.185 4.486 22.38 4.771 ;
      RECT 22.185 4.541 22.42 4.77 ;
      RECT 22.185 4.576 22.435 4.764 ;
      RECT 22.185 4.61 22.445 4.754 ;
      RECT 22.175 4.49 22.38 4.605 ;
      RECT 22.175 4.51 22.395 4.605 ;
      RECT 22.175 4.493 22.385 4.605 ;
      RECT 22.4 3.261 22.405 3.323 ;
      RECT 22.395 3.183 22.4 3.346 ;
      RECT 22.39 3.14 22.395 3.357 ;
      RECT 22.385 3.13 22.39 3.369 ;
      RECT 22.38 3.13 22.385 3.378 ;
      RECT 22.355 3.13 22.38 3.41 ;
      RECT 22.35 3.13 22.355 3.443 ;
      RECT 22.335 3.13 22.35 3.468 ;
      RECT 22.325 3.13 22.335 3.495 ;
      RECT 22.32 3.13 22.325 3.508 ;
      RECT 22.315 3.13 22.32 3.523 ;
      RECT 22.305 3.13 22.315 3.538 ;
      RECT 22.3 3.13 22.305 3.558 ;
      RECT 22.275 3.13 22.3 3.593 ;
      RECT 22.23 3.13 22.275 3.638 ;
      RECT 22.22 3.13 22.23 3.651 ;
      RECT 22.135 3.215 22.22 3.658 ;
      RECT 22.1 3.337 22.135 3.667 ;
      RECT 22.095 3.377 22.1 3.671 ;
      RECT 22.075 3.4 22.095 3.673 ;
      RECT 22.07 3.43 22.075 3.676 ;
      RECT 22.06 3.442 22.07 3.677 ;
      RECT 22.015 3.465 22.06 3.682 ;
      RECT 21.975 3.495 22.015 3.69 ;
      RECT 21.94 3.507 21.975 3.696 ;
      RECT 21.935 3.512 21.94 3.7 ;
      RECT 21.865 3.522 21.935 3.707 ;
      RECT 21.825 3.532 21.865 3.717 ;
      RECT 21.805 3.537 21.825 3.723 ;
      RECT 21.795 3.541 21.805 3.728 ;
      RECT 21.79 3.544 21.795 3.731 ;
      RECT 21.78 3.545 21.79 3.732 ;
      RECT 21.755 3.547 21.78 3.736 ;
      RECT 21.745 3.552 21.755 3.739 ;
      RECT 21.7 3.56 21.745 3.74 ;
      RECT 21.575 3.565 21.7 3.74 ;
      RECT 22.13 3.862 22.15 4.044 ;
      RECT 22.081 3.847 22.13 4.043 ;
      RECT 21.995 3.862 22.15 4.041 ;
      RECT 21.98 3.862 22.15 4.04 ;
      RECT 21.945 3.84 22.115 4.025 ;
      RECT 22.015 4.86 22.03 5.069 ;
      RECT 22.015 4.868 22.035 5.068 ;
      RECT 21.96 4.868 22.035 5.067 ;
      RECT 21.94 4.872 22.04 5.065 ;
      RECT 21.92 4.822 21.96 5.064 ;
      RECT 21.865 4.88 22.045 5.062 ;
      RECT 21.83 4.837 21.96 5.06 ;
      RECT 21.826 4.84 22.015 5.059 ;
      RECT 21.74 4.848 22.015 5.057 ;
      RECT 21.74 4.892 22.05 5.05 ;
      RECT 21.73 4.985 22.05 5.048 ;
      RECT 21.74 4.904 22.055 5.033 ;
      RECT 21.74 4.925 22.07 5.003 ;
      RECT 21.74 4.952 22.075 4.973 ;
      RECT 21.865 4.83 21.96 5.062 ;
      RECT 21.495 3.875 21.5 4.413 ;
      RECT 21.3 4.205 21.305 4.4 ;
      RECT 19.6 3.87 19.615 4.25 ;
      RECT 21.665 3.87 21.67 4.04 ;
      RECT 21.66 3.87 21.665 4.05 ;
      RECT 21.655 3.87 21.66 4.063 ;
      RECT 21.63 3.87 21.655 4.105 ;
      RECT 21.605 3.87 21.63 4.178 ;
      RECT 21.59 3.87 21.605 4.23 ;
      RECT 21.585 3.87 21.59 4.26 ;
      RECT 21.56 3.87 21.585 4.3 ;
      RECT 21.545 3.87 21.56 4.355 ;
      RECT 21.54 3.87 21.545 4.388 ;
      RECT 21.515 3.87 21.54 4.408 ;
      RECT 21.5 3.87 21.515 4.414 ;
      RECT 21.43 3.905 21.495 4.41 ;
      RECT 21.38 3.96 21.43 4.405 ;
      RECT 21.37 3.992 21.38 4.403 ;
      RECT 21.365 4.017 21.37 4.403 ;
      RECT 21.345 4.09 21.365 4.403 ;
      RECT 21.335 4.17 21.345 4.402 ;
      RECT 21.32 4.2 21.335 4.402 ;
      RECT 21.305 4.205 21.32 4.401 ;
      RECT 21.245 4.207 21.3 4.398 ;
      RECT 21.215 4.212 21.245 4.394 ;
      RECT 21.213 4.215 21.215 4.393 ;
      RECT 21.127 4.217 21.213 4.39 ;
      RECT 21.041 4.223 21.127 4.384 ;
      RECT 20.955 4.228 21.041 4.378 ;
      RECT 20.882 4.233 20.955 4.379 ;
      RECT 20.796 4.239 20.882 4.387 ;
      RECT 20.71 4.245 20.796 4.396 ;
      RECT 20.69 4.249 20.71 4.401 ;
      RECT 20.643 4.251 20.69 4.404 ;
      RECT 20.557 4.256 20.643 4.41 ;
      RECT 20.471 4.261 20.557 4.419 ;
      RECT 20.385 4.267 20.471 4.427 ;
      RECT 20.3 4.265 20.385 4.436 ;
      RECT 20.296 4.26 20.3 4.44 ;
      RECT 20.21 4.255 20.296 4.432 ;
      RECT 20.146 4.246 20.21 4.42 ;
      RECT 20.06 4.237 20.146 4.407 ;
      RECT 20.036 4.23 20.06 4.398 ;
      RECT 19.95 4.224 20.036 4.385 ;
      RECT 19.91 4.217 19.95 4.371 ;
      RECT 19.905 4.207 19.91 4.367 ;
      RECT 19.895 4.195 19.905 4.366 ;
      RECT 19.875 4.165 19.895 4.363 ;
      RECT 19.82 4.085 19.875 4.357 ;
      RECT 19.8 4.004 19.82 4.352 ;
      RECT 19.78 3.962 19.8 4.348 ;
      RECT 19.755 3.915 19.78 4.342 ;
      RECT 19.75 3.89 19.755 4.339 ;
      RECT 19.715 3.87 19.75 4.334 ;
      RECT 19.706 3.87 19.715 4.327 ;
      RECT 19.62 3.87 19.706 4.297 ;
      RECT 19.615 3.87 19.62 4.26 ;
      RECT 19.58 3.87 19.6 4.182 ;
      RECT 19.575 3.912 19.58 4.147 ;
      RECT 19.57 3.987 19.575 4.103 ;
      RECT 21.02 3.792 21.195 4.04 ;
      RECT 21.02 3.792 21.2 4.038 ;
      RECT 21.015 3.824 21.2 3.998 ;
      RECT 21.045 3.765 21.215 3.985 ;
      RECT 21.01 3.842 21.215 3.918 ;
      RECT 20.32 3.305 20.49 3.48 ;
      RECT 20.32 3.305 20.662 3.472 ;
      RECT 20.32 3.305 20.745 3.466 ;
      RECT 20.32 3.305 20.78 3.462 ;
      RECT 20.32 3.305 20.8 3.461 ;
      RECT 20.32 3.305 20.886 3.457 ;
      RECT 20.78 3.13 20.95 3.452 ;
      RECT 20.355 3.237 20.98 3.45 ;
      RECT 20.345 3.292 20.985 3.448 ;
      RECT 20.32 3.328 20.995 3.443 ;
      RECT 20.32 3.355 21 3.373 ;
      RECT 20.385 3.18 20.96 3.45 ;
      RECT 20.576 3.165 20.96 3.45 ;
      RECT 20.41 3.168 20.96 3.45 ;
      RECT 20.49 3.166 20.576 3.477 ;
      RECT 20.576 3.163 20.955 3.45 ;
      RECT 20.76 3.14 20.955 3.45 ;
      RECT 20.662 3.161 20.955 3.45 ;
      RECT 20.745 3.155 20.76 3.463 ;
      RECT 20.895 4.52 20.9 4.72 ;
      RECT 20.36 4.585 20.405 4.72 ;
      RECT 20.93 4.52 20.95 4.693 ;
      RECT 20.9 4.52 20.93 4.708 ;
      RECT 20.835 4.52 20.895 4.745 ;
      RECT 20.82 4.52 20.835 4.775 ;
      RECT 20.805 4.52 20.82 4.788 ;
      RECT 20.785 4.52 20.805 4.803 ;
      RECT 20.78 4.52 20.785 4.812 ;
      RECT 20.77 4.524 20.78 4.817 ;
      RECT 20.755 4.534 20.77 4.828 ;
      RECT 20.73 4.55 20.755 4.838 ;
      RECT 20.72 4.564 20.73 4.84 ;
      RECT 20.7 4.576 20.72 4.837 ;
      RECT 20.67 4.597 20.7 4.831 ;
      RECT 20.66 4.609 20.67 4.826 ;
      RECT 20.65 4.607 20.66 4.823 ;
      RECT 20.635 4.606 20.65 4.818 ;
      RECT 20.63 4.605 20.635 4.813 ;
      RECT 20.595 4.603 20.63 4.803 ;
      RECT 20.575 4.6 20.595 4.785 ;
      RECT 20.565 4.598 20.575 4.78 ;
      RECT 20.555 4.597 20.565 4.775 ;
      RECT 20.52 4.595 20.555 4.763 ;
      RECT 20.465 4.591 20.52 4.743 ;
      RECT 20.455 4.589 20.465 4.728 ;
      RECT 20.45 4.589 20.455 4.723 ;
      RECT 20.405 4.587 20.45 4.72 ;
      RECT 20.31 4.585 20.36 4.724 ;
      RECT 20.3 4.586 20.31 4.729 ;
      RECT 20.24 4.593 20.3 4.743 ;
      RECT 20.215 4.601 20.24 4.763 ;
      RECT 20.205 4.605 20.215 4.775 ;
      RECT 20.2 4.606 20.205 4.78 ;
      RECT 20.185 4.608 20.2 4.783 ;
      RECT 20.17 4.61 20.185 4.788 ;
      RECT 20.165 4.61 20.17 4.791 ;
      RECT 20.12 4.615 20.165 4.802 ;
      RECT 20.115 4.619 20.12 4.814 ;
      RECT 20.09 4.615 20.115 4.818 ;
      RECT 20.08 4.611 20.09 4.822 ;
      RECT 20.07 4.61 20.08 4.826 ;
      RECT 20.055 4.6 20.07 4.832 ;
      RECT 20.05 4.588 20.055 4.836 ;
      RECT 20.045 4.585 20.05 4.837 ;
      RECT 20.04 4.582 20.045 4.839 ;
      RECT 20.025 4.57 20.04 4.838 ;
      RECT 20.01 4.552 20.025 4.835 ;
      RECT 19.99 4.531 20.01 4.828 ;
      RECT 19.925 4.52 19.99 4.8 ;
      RECT 19.921 4.52 19.925 4.779 ;
      RECT 19.835 4.52 19.921 4.749 ;
      RECT 19.82 4.52 19.835 4.705 ;
      RECT 20.47 4.871 20.485 5.13 ;
      RECT 20.47 4.886 20.49 5.129 ;
      RECT 20.386 4.886 20.49 5.127 ;
      RECT 20.386 4.9 20.495 5.126 ;
      RECT 20.3 4.942 20.5 5.123 ;
      RECT 20.295 4.885 20.485 5.118 ;
      RECT 20.295 4.956 20.505 5.115 ;
      RECT 20.29 4.987 20.505 5.113 ;
      RECT 20.295 4.984 20.52 5.103 ;
      RECT 20.29 5.03 20.535 5.088 ;
      RECT 20.29 5.058 20.54 5.073 ;
      RECT 20.3 4.86 20.47 5.123 ;
      RECT 20.06 3.87 20.23 4.04 ;
      RECT 20.025 3.87 20.23 4.035 ;
      RECT 20.015 3.87 20.23 4.028 ;
      RECT 20.01 3.855 20.18 4.025 ;
      RECT 18.84 4.392 19.105 4.835 ;
      RECT 18.835 4.363 19.05 4.833 ;
      RECT 18.83 4.517 19.11 4.828 ;
      RECT 18.835 4.412 19.11 4.828 ;
      RECT 18.835 4.423 19.12 4.815 ;
      RECT 18.835 4.37 19.08 4.833 ;
      RECT 18.84 4.357 19.05 4.835 ;
      RECT 18.84 4.355 19 4.835 ;
      RECT 18.941 4.347 19 4.835 ;
      RECT 18.855 4.348 19 4.835 ;
      RECT 18.941 4.346 18.99 4.835 ;
      RECT 18.745 3.161 18.92 3.46 ;
      RECT 18.795 3.123 18.92 3.46 ;
      RECT 18.78 3.125 19.006 3.452 ;
      RECT 18.78 3.128 19.045 3.439 ;
      RECT 18.78 3.129 19.055 3.425 ;
      RECT 18.735 3.18 19.055 3.415 ;
      RECT 18.78 3.13 19.06 3.41 ;
      RECT 18.735 3.34 19.065 3.4 ;
      RECT 18.72 3.2 19.06 3.34 ;
      RECT 18.715 3.216 19.06 3.28 ;
      RECT 18.76 3.14 19.06 3.41 ;
      RECT 18.795 3.121 18.881 3.46 ;
      RECT 16.605 7.31 16.775 9.52 ;
      RECT 16.605 7.31 16.78 8.57 ;
      RECT 16.175 10.15 16.345 10.6 ;
      RECT 16.235 8.37 16.405 10.32 ;
      RECT 16.175 7.31 16.345 8.54 ;
      RECT 15.65 10.11 15.825 10.6 ;
      RECT 15.65 7.31 15.82 10.6 ;
      RECT 15.65 9.61 16.06 9.94 ;
      RECT 15.65 8.77 16.06 9.1 ;
      RECT 15.65 7.31 15.825 8.57 ;
      RECT 93.555 10.09 93.73 10.6 ;
      RECT 92.565 1.865 92.74 2.375 ;
      RECT 92.565 10.09 92.74 10.6 ;
      RECT 90.775 1.865 90.95 2.375 ;
      RECT 90.775 10.09 90.95 10.6 ;
      RECT 85.14 10.09 85.315 10.6 ;
      RECT 78.295 10.09 78.47 10.6 ;
      RECT 77.305 1.865 77.48 2.375 ;
      RECT 77.305 10.09 77.48 10.6 ;
      RECT 75.515 1.865 75.69 2.375 ;
      RECT 75.515 10.09 75.69 10.6 ;
      RECT 69.88 10.09 70.055 10.6 ;
      RECT 63.035 10.09 63.21 10.6 ;
      RECT 62.045 1.865 62.22 2.375 ;
      RECT 62.045 10.09 62.22 10.6 ;
      RECT 60.255 1.865 60.43 2.375 ;
      RECT 60.255 10.09 60.43 10.6 ;
      RECT 54.62 10.09 54.795 10.6 ;
      RECT 47.775 10.09 47.95 10.6 ;
      RECT 46.785 1.865 46.96 2.375 ;
      RECT 46.785 10.09 46.96 10.6 ;
      RECT 44.995 1.865 45.17 2.375 ;
      RECT 44.995 10.09 45.17 10.6 ;
      RECT 39.36 10.09 39.535 10.6 ;
      RECT 32.515 10.09 32.69 10.6 ;
      RECT 31.525 1.865 31.7 2.375 ;
      RECT 31.525 10.09 31.7 10.6 ;
      RECT 29.735 1.865 29.91 2.375 ;
      RECT 29.735 10.09 29.91 10.6 ;
      RECT 24.1 10.09 24.275 10.6 ;
      RECT 16.605 10.09 16.78 10.6 ;
  END
END sky130_osu_ring_oscillator_mpr2ya_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2ya_8_b0r2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ya_8_b0r2 ;
  SIZE 94.105 BY 12.465 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 32.41 0 32.79 5.26 ;
      LAYER met2 ;
        RECT 32.41 4.88 32.79 5.26 ;
      LAYER li1 ;
        RECT 32.51 1.865 32.685 2.375 ;
        RECT 32.51 3.895 32.685 5.155 ;
        RECT 32.51 3.685 32.68 5.155 ;
      LAYER met1 ;
        RECT 32.425 4.925 32.775 5.215 ;
        RECT 32.45 2.175 32.745 2.405 ;
        RECT 32.45 3.655 32.74 3.885 ;
        RECT 32.51 2.175 32.68 3.885 ;
      LAYER via1 ;
        RECT 32.525 4.995 32.675 5.145 ;
      LAYER via2 ;
        RECT 32.5 4.97 32.7 5.17 ;
      LAYER mcon ;
        RECT 32.51 3.685 32.68 3.855 ;
        RECT 32.515 4.985 32.685 5.155 ;
        RECT 32.51 2.205 32.685 2.375 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 47.67 0 48.05 5.26 ;
      LAYER met2 ;
        RECT 47.67 4.88 48.05 5.26 ;
      LAYER li1 ;
        RECT 47.77 1.865 47.945 2.375 ;
        RECT 47.77 3.895 47.945 5.155 ;
        RECT 47.77 3.685 47.94 5.155 ;
      LAYER met1 ;
        RECT 47.685 4.925 48.035 5.215 ;
        RECT 47.71 2.175 48.005 2.405 ;
        RECT 47.71 3.655 48 3.885 ;
        RECT 47.77 2.175 47.94 3.885 ;
      LAYER via1 ;
        RECT 47.785 4.995 47.935 5.145 ;
      LAYER via2 ;
        RECT 47.76 4.97 47.96 5.17 ;
      LAYER mcon ;
        RECT 47.77 3.685 47.94 3.855 ;
        RECT 47.775 4.985 47.945 5.155 ;
        RECT 47.77 2.205 47.945 2.375 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 62.93 0 63.31 5.26 ;
      LAYER met2 ;
        RECT 62.93 4.88 63.31 5.26 ;
      LAYER li1 ;
        RECT 63.03 1.865 63.205 2.375 ;
        RECT 63.03 3.895 63.205 5.155 ;
        RECT 63.03 3.685 63.2 5.155 ;
      LAYER met1 ;
        RECT 62.945 4.925 63.295 5.215 ;
        RECT 62.97 2.175 63.265 2.405 ;
        RECT 62.97 3.655 63.26 3.885 ;
        RECT 63.03 2.175 63.2 3.885 ;
      LAYER via1 ;
        RECT 63.045 4.995 63.195 5.145 ;
      LAYER via2 ;
        RECT 63.02 4.97 63.22 5.17 ;
      LAYER mcon ;
        RECT 63.03 3.685 63.2 3.855 ;
        RECT 63.035 4.985 63.205 5.155 ;
        RECT 63.03 2.205 63.205 2.375 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 78.19 0 78.57 5.26 ;
      LAYER met2 ;
        RECT 78.19 4.88 78.57 5.26 ;
      LAYER li1 ;
        RECT 78.29 1.865 78.465 2.375 ;
        RECT 78.29 3.895 78.465 5.155 ;
        RECT 78.29 3.685 78.46 5.155 ;
      LAYER met1 ;
        RECT 78.205 4.925 78.555 5.215 ;
        RECT 78.23 2.175 78.525 2.405 ;
        RECT 78.23 3.655 78.52 3.885 ;
        RECT 78.29 2.175 78.46 3.885 ;
      LAYER via1 ;
        RECT 78.305 4.995 78.455 5.145 ;
      LAYER via2 ;
        RECT 78.28 4.97 78.48 5.17 ;
      LAYER mcon ;
        RECT 78.29 3.685 78.46 3.855 ;
        RECT 78.295 4.985 78.465 5.155 ;
        RECT 78.29 2.205 78.465 2.375 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.14575 ;
    PORT
      LAYER met3 ;
        RECT 93.45 0 93.83 5.26 ;
      LAYER met2 ;
        RECT 93.45 4.88 93.83 5.26 ;
      LAYER li1 ;
        RECT 93.55 1.865 93.725 2.375 ;
        RECT 93.55 3.895 93.725 5.155 ;
        RECT 93.55 3.685 93.72 5.155 ;
      LAYER met1 ;
        RECT 93.465 4.925 93.815 5.215 ;
        RECT 93.49 2.175 93.785 2.405 ;
        RECT 93.49 3.655 93.78 3.885 ;
        RECT 93.55 2.175 93.72 3.885 ;
      LAYER via1 ;
        RECT 93.565 4.995 93.715 5.145 ;
      LAYER via2 ;
        RECT 93.54 4.97 93.74 5.17 ;
      LAYER mcon ;
        RECT 93.55 3.685 93.72 3.855 ;
        RECT 93.555 4.985 93.725 5.155 ;
        RECT 93.55 2.205 93.725 2.375 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 28.285 4 28.625 4.35 ;
        RECT 28.28 8.15 28.62 8.5 ;
        RECT 28.36 4 28.535 8.5 ;
      LAYER li1 ;
        RECT 28.36 2.955 28.53 4.225 ;
        RECT 28.36 8.24 28.53 9.51 ;
        RECT 22.725 8.24 22.895 9.51 ;
      LAYER met1 ;
        RECT 28.285 4.055 28.76 4.225 ;
        RECT 28.285 4 28.625 4.35 ;
        RECT 28.28 8.24 28.76 8.41 ;
        RECT 28.28 8.15 28.62 8.5 ;
        RECT 22.665 8.235 28.62 8.405 ;
        RECT 22.665 8.235 23.125 8.41 ;
        RECT 22.665 8.21 22.955 8.44 ;
      LAYER via1 ;
        RECT 28.38 8.25 28.53 8.4 ;
        RECT 28.385 4.1 28.535 4.25 ;
      LAYER mcon ;
        RECT 22.725 8.24 22.895 8.41 ;
        RECT 28.36 8.24 28.53 8.41 ;
        RECT 28.36 4.055 28.53 4.225 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 43.545 4 43.885 4.35 ;
        RECT 43.54 8.15 43.88 8.5 ;
        RECT 43.62 4 43.795 8.5 ;
      LAYER li1 ;
        RECT 43.62 2.955 43.79 4.225 ;
        RECT 43.62 8.24 43.79 9.51 ;
        RECT 37.985 8.24 38.155 9.51 ;
      LAYER met1 ;
        RECT 43.545 4.055 44.02 4.225 ;
        RECT 43.545 4 43.885 4.35 ;
        RECT 43.54 8.24 44.02 8.41 ;
        RECT 43.54 8.15 43.88 8.5 ;
        RECT 37.925 8.235 43.88 8.405 ;
        RECT 37.925 8.235 38.385 8.41 ;
        RECT 37.925 8.21 38.215 8.44 ;
      LAYER via1 ;
        RECT 43.64 8.25 43.79 8.4 ;
        RECT 43.645 4.1 43.795 4.25 ;
      LAYER mcon ;
        RECT 37.985 8.24 38.155 8.41 ;
        RECT 43.62 8.24 43.79 8.41 ;
        RECT 43.62 4.055 43.79 4.225 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 58.805 4 59.145 4.35 ;
        RECT 58.8 8.15 59.14 8.5 ;
        RECT 58.88 4 59.055 8.5 ;
      LAYER li1 ;
        RECT 58.88 2.955 59.05 4.225 ;
        RECT 58.88 8.24 59.05 9.51 ;
        RECT 53.245 8.24 53.415 9.51 ;
      LAYER met1 ;
        RECT 58.805 4.055 59.28 4.225 ;
        RECT 58.805 4 59.145 4.35 ;
        RECT 58.8 8.24 59.28 8.41 ;
        RECT 58.8 8.15 59.14 8.5 ;
        RECT 53.185 8.235 59.14 8.405 ;
        RECT 53.185 8.235 53.645 8.41 ;
        RECT 53.185 8.21 53.475 8.44 ;
      LAYER via1 ;
        RECT 58.9 8.25 59.05 8.4 ;
        RECT 58.905 4.1 59.055 4.25 ;
      LAYER mcon ;
        RECT 53.245 8.24 53.415 8.41 ;
        RECT 58.88 8.24 59.05 8.41 ;
        RECT 58.88 4.055 59.05 4.225 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 74.065 4 74.405 4.35 ;
        RECT 74.06 8.15 74.4 8.5 ;
        RECT 74.14 4 74.315 8.5 ;
      LAYER li1 ;
        RECT 74.14 2.955 74.31 4.225 ;
        RECT 74.14 8.24 74.31 9.51 ;
        RECT 68.505 8.24 68.675 9.51 ;
      LAYER met1 ;
        RECT 74.065 4.055 74.54 4.225 ;
        RECT 74.065 4 74.405 4.35 ;
        RECT 74.06 8.24 74.54 8.41 ;
        RECT 74.06 8.15 74.4 8.5 ;
        RECT 68.445 8.235 74.4 8.405 ;
        RECT 68.445 8.235 68.905 8.41 ;
        RECT 68.445 8.21 68.735 8.44 ;
      LAYER via1 ;
        RECT 74.16 8.25 74.31 8.4 ;
        RECT 74.165 4.1 74.315 4.25 ;
      LAYER mcon ;
        RECT 68.505 8.24 68.675 8.41 ;
        RECT 74.14 8.24 74.31 8.41 ;
        RECT 74.14 4.055 74.31 4.225 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER met2 ;
        RECT 89.325 4 89.665 4.35 ;
        RECT 89.32 8.15 89.66 8.5 ;
        RECT 89.4 4 89.575 8.5 ;
      LAYER li1 ;
        RECT 89.4 2.955 89.57 4.225 ;
        RECT 89.4 8.24 89.57 9.51 ;
        RECT 83.765 8.24 83.935 9.51 ;
      LAYER met1 ;
        RECT 89.325 4.055 89.8 4.225 ;
        RECT 89.325 4 89.665 4.35 ;
        RECT 89.32 8.24 89.8 8.41 ;
        RECT 89.32 8.15 89.66 8.5 ;
        RECT 83.705 8.235 89.66 8.405 ;
        RECT 83.705 8.235 84.165 8.41 ;
        RECT 83.705 8.21 83.995 8.44 ;
      LAYER via1 ;
        RECT 89.42 8.25 89.57 8.4 ;
        RECT 89.425 4.1 89.575 4.25 ;
      LAYER mcon ;
        RECT 83.765 8.24 83.935 8.41 ;
        RECT 89.4 8.24 89.57 8.41 ;
        RECT 89.4 4.055 89.57 4.225 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 15.23 8.24 15.4 9.51 ;
      LAYER met1 ;
        RECT 15.17 8.24 15.63 8.41 ;
        RECT 15.175 8.205 15.465 8.435 ;
        RECT 15.17 8.21 15.46 8.44 ;
      LAYER mcon ;
        RECT 15.23 8.24 15.4 8.41 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 5.435 94.1 7.035 ;
        RECT 79.59 5.43 94.1 7.035 ;
        RECT 89.22 5.43 93.945 7.04 ;
        RECT 89.22 5.425 93.94 7.04 ;
        RECT 93.125 5.425 93.295 7.77 ;
        RECT 93.12 4.695 93.29 7.04 ;
        RECT 92.135 4.695 92.305 7.77 ;
        RECT 89.39 4.695 89.56 7.77 ;
        RECT 86.62 4.93 86.79 7.035 ;
        RECT 83.585 5.43 86.335 7.04 ;
        RECT 84.7 4.93 84.87 7.04 ;
        RECT 83.76 4.93 83.93 7.04 ;
        RECT 83.755 5.43 83.925 7.77 ;
        RECT 82.3 4.93 82.47 7.035 ;
        RECT 80.38 4.93 80.55 7.035 ;
        RECT 64.33 5.43 78.84 7.035 ;
        RECT 73.96 5.43 78.685 7.04 ;
        RECT 73.96 5.425 78.68 7.04 ;
        RECT 77.865 5.425 78.035 7.77 ;
        RECT 77.86 4.695 78.03 7.04 ;
        RECT 76.875 4.695 77.045 7.77 ;
        RECT 74.13 4.695 74.3 7.77 ;
        RECT 71.36 4.93 71.53 7.035 ;
        RECT 68.325 5.43 71.075 7.04 ;
        RECT 69.44 4.93 69.61 7.04 ;
        RECT 68.5 4.93 68.67 7.04 ;
        RECT 68.495 5.43 68.665 7.77 ;
        RECT 67.04 4.93 67.21 7.035 ;
        RECT 65.12 4.93 65.29 7.035 ;
        RECT 49.07 5.43 63.58 7.035 ;
        RECT 58.7 5.43 63.425 7.04 ;
        RECT 58.7 5.425 63.42 7.04 ;
        RECT 62.605 5.425 62.775 7.77 ;
        RECT 62.6 4.695 62.77 7.04 ;
        RECT 61.615 4.695 61.785 7.77 ;
        RECT 58.87 4.695 59.04 7.77 ;
        RECT 56.1 4.93 56.27 7.035 ;
        RECT 53.065 5.43 55.815 7.04 ;
        RECT 54.18 4.93 54.35 7.04 ;
        RECT 53.24 4.93 53.41 7.04 ;
        RECT 53.235 5.43 53.405 7.77 ;
        RECT 51.78 4.93 51.95 7.035 ;
        RECT 49.86 4.93 50.03 7.035 ;
        RECT 33.81 5.43 48.32 7.035 ;
        RECT 43.44 5.43 48.165 7.04 ;
        RECT 43.44 5.425 48.16 7.04 ;
        RECT 47.345 5.425 47.515 7.77 ;
        RECT 47.34 4.695 47.51 7.04 ;
        RECT 46.355 4.695 46.525 7.77 ;
        RECT 43.61 4.695 43.78 7.77 ;
        RECT 40.84 4.93 41.01 7.035 ;
        RECT 37.805 5.43 40.555 7.04 ;
        RECT 38.92 4.93 39.09 7.04 ;
        RECT 37.98 4.93 38.15 7.04 ;
        RECT 37.975 5.43 38.145 7.77 ;
        RECT 36.52 4.93 36.69 7.035 ;
        RECT 34.6 4.93 34.77 7.035 ;
        RECT 18.55 5.43 33.06 7.035 ;
        RECT 28.18 5.43 32.905 7.04 ;
        RECT 28.18 5.425 32.9 7.04 ;
        RECT 32.085 5.425 32.255 7.77 ;
        RECT 32.08 4.695 32.25 7.04 ;
        RECT 31.095 4.695 31.265 7.77 ;
        RECT 28.35 4.695 28.52 7.77 ;
        RECT 25.58 4.93 25.75 7.035 ;
        RECT 22.545 5.43 25.295 7.04 ;
        RECT 23.66 4.93 23.83 7.04 ;
        RECT 22.72 4.93 22.89 7.04 ;
        RECT 22.715 5.43 22.885 7.77 ;
        RECT 21.26 4.93 21.43 7.035 ;
        RECT 19.34 4.93 19.51 7.035 ;
        RECT 15.05 5.435 17.8 7.04 ;
        RECT 17.035 10.05 17.21 10.6 ;
        RECT 17.035 7.31 17.21 8.45 ;
        RECT 17.035 5.435 17.205 10.6 ;
        RECT 15.22 5.435 15.39 7.77 ;
      LAYER met1 ;
        RECT 17.805 5.43 94.105 7.03 ;
        RECT 0 5.435 94.1 7.035 ;
        RECT 89.22 5.43 93.945 7.04 ;
        RECT 89.22 5.425 93.94 7.04 ;
        RECT 79.59 5.275 88.33 7.035 ;
        RECT 83.585 5.275 86.335 7.04 ;
        RECT 73.96 5.43 78.685 7.04 ;
        RECT 73.96 5.425 78.68 7.04 ;
        RECT 64.33 5.275 73.07 7.035 ;
        RECT 68.325 5.275 71.075 7.04 ;
        RECT 58.7 5.43 63.425 7.04 ;
        RECT 58.7 5.425 63.42 7.04 ;
        RECT 49.07 5.275 57.81 7.035 ;
        RECT 53.065 5.275 55.815 7.04 ;
        RECT 43.44 5.43 48.165 7.04 ;
        RECT 43.44 5.425 48.16 7.04 ;
        RECT 33.81 5.275 42.55 7.035 ;
        RECT 37.805 5.275 40.555 7.04 ;
        RECT 28.18 5.43 32.905 7.04 ;
        RECT 28.18 5.425 32.9 7.04 ;
        RECT 18.55 5.275 27.29 7.035 ;
        RECT 22.545 5.275 25.295 7.04 ;
        RECT 15.05 5.435 17.8 7.04 ;
        RECT 16.975 8.95 17.265 9.18 ;
        RECT 16.805 8.98 17.265 9.15 ;
      LAYER mcon ;
        RECT 17.035 8.98 17.205 9.15 ;
        RECT 17.34 6.84 17.51 7.01 ;
        RECT 18.695 5.43 18.865 5.6 ;
        RECT 19.155 5.43 19.325 5.6 ;
        RECT 19.615 5.43 19.785 5.6 ;
        RECT 20.075 5.43 20.245 5.6 ;
        RECT 20.535 5.43 20.705 5.6 ;
        RECT 20.995 5.43 21.165 5.6 ;
        RECT 21.455 5.43 21.625 5.6 ;
        RECT 21.915 5.43 22.085 5.6 ;
        RECT 22.375 5.43 22.545 5.6 ;
        RECT 22.835 5.43 23.005 5.6 ;
        RECT 23.295 5.43 23.465 5.6 ;
        RECT 23.755 5.43 23.925 5.6 ;
        RECT 24.215 5.43 24.385 5.6 ;
        RECT 24.675 5.43 24.845 5.6 ;
        RECT 24.835 6.84 25.005 7.01 ;
        RECT 25.135 5.43 25.305 5.6 ;
        RECT 25.595 5.43 25.765 5.6 ;
        RECT 26.055 5.43 26.225 5.6 ;
        RECT 26.515 5.43 26.685 5.6 ;
        RECT 26.975 5.43 27.145 5.6 ;
        RECT 30.47 6.84 30.64 7.01 ;
        RECT 30.47 5.455 30.64 5.625 ;
        RECT 31.175 6.84 31.345 7.01 ;
        RECT 31.175 5.455 31.345 5.625 ;
        RECT 32.16 5.455 32.33 5.625 ;
        RECT 32.165 6.84 32.335 7.01 ;
        RECT 33.955 5.43 34.125 5.6 ;
        RECT 34.415 5.43 34.585 5.6 ;
        RECT 34.875 5.43 35.045 5.6 ;
        RECT 35.335 5.43 35.505 5.6 ;
        RECT 35.795 5.43 35.965 5.6 ;
        RECT 36.255 5.43 36.425 5.6 ;
        RECT 36.715 5.43 36.885 5.6 ;
        RECT 37.175 5.43 37.345 5.6 ;
        RECT 37.635 5.43 37.805 5.6 ;
        RECT 38.095 5.43 38.265 5.6 ;
        RECT 38.555 5.43 38.725 5.6 ;
        RECT 39.015 5.43 39.185 5.6 ;
        RECT 39.475 5.43 39.645 5.6 ;
        RECT 39.935 5.43 40.105 5.6 ;
        RECT 40.095 6.84 40.265 7.01 ;
        RECT 40.395 5.43 40.565 5.6 ;
        RECT 40.855 5.43 41.025 5.6 ;
        RECT 41.315 5.43 41.485 5.6 ;
        RECT 41.775 5.43 41.945 5.6 ;
        RECT 42.235 5.43 42.405 5.6 ;
        RECT 45.73 6.84 45.9 7.01 ;
        RECT 45.73 5.455 45.9 5.625 ;
        RECT 46.435 6.84 46.605 7.01 ;
        RECT 46.435 5.455 46.605 5.625 ;
        RECT 47.42 5.455 47.59 5.625 ;
        RECT 47.425 6.84 47.595 7.01 ;
        RECT 49.215 5.43 49.385 5.6 ;
        RECT 49.675 5.43 49.845 5.6 ;
        RECT 50.135 5.43 50.305 5.6 ;
        RECT 50.595 5.43 50.765 5.6 ;
        RECT 51.055 5.43 51.225 5.6 ;
        RECT 51.515 5.43 51.685 5.6 ;
        RECT 51.975 5.43 52.145 5.6 ;
        RECT 52.435 5.43 52.605 5.6 ;
        RECT 52.895 5.43 53.065 5.6 ;
        RECT 53.355 5.43 53.525 5.6 ;
        RECT 53.815 5.43 53.985 5.6 ;
        RECT 54.275 5.43 54.445 5.6 ;
        RECT 54.735 5.43 54.905 5.6 ;
        RECT 55.195 5.43 55.365 5.6 ;
        RECT 55.355 6.84 55.525 7.01 ;
        RECT 55.655 5.43 55.825 5.6 ;
        RECT 56.115 5.43 56.285 5.6 ;
        RECT 56.575 5.43 56.745 5.6 ;
        RECT 57.035 5.43 57.205 5.6 ;
        RECT 57.495 5.43 57.665 5.6 ;
        RECT 60.99 6.84 61.16 7.01 ;
        RECT 60.99 5.455 61.16 5.625 ;
        RECT 61.695 6.84 61.865 7.01 ;
        RECT 61.695 5.455 61.865 5.625 ;
        RECT 62.68 5.455 62.85 5.625 ;
        RECT 62.685 6.84 62.855 7.01 ;
        RECT 64.475 5.43 64.645 5.6 ;
        RECT 64.935 5.43 65.105 5.6 ;
        RECT 65.395 5.43 65.565 5.6 ;
        RECT 65.855 5.43 66.025 5.6 ;
        RECT 66.315 5.43 66.485 5.6 ;
        RECT 66.775 5.43 66.945 5.6 ;
        RECT 67.235 5.43 67.405 5.6 ;
        RECT 67.695 5.43 67.865 5.6 ;
        RECT 68.155 5.43 68.325 5.6 ;
        RECT 68.615 5.43 68.785 5.6 ;
        RECT 69.075 5.43 69.245 5.6 ;
        RECT 69.535 5.43 69.705 5.6 ;
        RECT 69.995 5.43 70.165 5.6 ;
        RECT 70.455 5.43 70.625 5.6 ;
        RECT 70.615 6.84 70.785 7.01 ;
        RECT 70.915 5.43 71.085 5.6 ;
        RECT 71.375 5.43 71.545 5.6 ;
        RECT 71.835 5.43 72.005 5.6 ;
        RECT 72.295 5.43 72.465 5.6 ;
        RECT 72.755 5.43 72.925 5.6 ;
        RECT 76.25 6.84 76.42 7.01 ;
        RECT 76.25 5.455 76.42 5.625 ;
        RECT 76.955 6.84 77.125 7.01 ;
        RECT 76.955 5.455 77.125 5.625 ;
        RECT 77.94 5.455 78.11 5.625 ;
        RECT 77.945 6.84 78.115 7.01 ;
        RECT 79.735 5.43 79.905 5.6 ;
        RECT 80.195 5.43 80.365 5.6 ;
        RECT 80.655 5.43 80.825 5.6 ;
        RECT 81.115 5.43 81.285 5.6 ;
        RECT 81.575 5.43 81.745 5.6 ;
        RECT 82.035 5.43 82.205 5.6 ;
        RECT 82.495 5.43 82.665 5.6 ;
        RECT 82.955 5.43 83.125 5.6 ;
        RECT 83.415 5.43 83.585 5.6 ;
        RECT 83.875 5.43 84.045 5.6 ;
        RECT 84.335 5.43 84.505 5.6 ;
        RECT 84.795 5.43 84.965 5.6 ;
        RECT 85.255 5.43 85.425 5.6 ;
        RECT 85.715 5.43 85.885 5.6 ;
        RECT 85.875 6.84 86.045 7.01 ;
        RECT 86.175 5.43 86.345 5.6 ;
        RECT 86.635 5.43 86.805 5.6 ;
        RECT 87.095 5.43 87.265 5.6 ;
        RECT 87.555 5.43 87.725 5.6 ;
        RECT 88.015 5.43 88.185 5.6 ;
        RECT 91.51 6.84 91.68 7.01 ;
        RECT 91.51 5.455 91.68 5.625 ;
        RECT 92.215 6.84 92.385 7.01 ;
        RECT 92.215 5.455 92.385 5.625 ;
        RECT 93.2 5.455 93.37 5.625 ;
        RECT 93.205 6.84 93.375 7.01 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 81.5 3.31 81.83 4.04 ;
        RECT 66.24 3.31 66.57 4.04 ;
        RECT 50.98 3.31 51.31 4.04 ;
        RECT 35.72 3.31 36.05 4.04 ;
        RECT 20.46 3.31 20.79 4.04 ;
      LAYER met2 ;
        RECT 81.605 2.24 81.975 2.61 ;
        RECT 81.615 3.625 81.875 3.885 ;
        RECT 81.705 2.24 81.87 3.885 ;
        RECT 81.525 3.735 81.83 3.945 ;
        RECT 81.525 3.735 81.805 4.015 ;
        RECT 81.58 3.72 81.875 3.885 ;
        RECT 66.345 2.24 66.715 2.61 ;
        RECT 66.355 3.625 66.615 3.885 ;
        RECT 66.445 2.24 66.61 3.885 ;
        RECT 66.265 3.735 66.57 3.945 ;
        RECT 66.265 3.735 66.545 4.015 ;
        RECT 66.32 3.72 66.615 3.885 ;
        RECT 51.085 2.24 51.455 2.61 ;
        RECT 51.095 3.625 51.355 3.885 ;
        RECT 51.185 2.24 51.35 3.885 ;
        RECT 51.005 3.735 51.31 3.945 ;
        RECT 51.005 3.735 51.285 4.015 ;
        RECT 51.06 3.72 51.355 3.885 ;
        RECT 35.825 2.24 36.195 2.61 ;
        RECT 35.835 3.625 36.095 3.885 ;
        RECT 35.925 2.24 36.09 3.885 ;
        RECT 35.745 3.735 36.05 3.945 ;
        RECT 35.745 3.735 36.025 4.015 ;
        RECT 35.8 3.72 36.095 3.885 ;
        RECT 20.565 2.24 20.935 2.61 ;
        RECT 20.575 3.625 20.835 3.885 ;
        RECT 20.665 2.24 20.83 3.885 ;
        RECT 20.485 3.735 20.79 3.945 ;
        RECT 20.485 3.735 20.765 4.015 ;
        RECT 20.54 3.72 20.835 3.885 ;
      LAYER li1 ;
        RECT 0.005 0 94.1 1.6 ;
        RECT 93.12 0 93.29 2.225 ;
        RECT 92.135 0 92.305 2.225 ;
        RECT 89.39 0 89.56 2.225 ;
        RECT 79.59 0 88.33 2.88 ;
        RECT 87.56 0 87.73 3.38 ;
        RECT 86.62 0 86.79 3.38 ;
        RECT 85.66 0 85.83 3.38 ;
        RECT 84.615 0 84.81 2.89 ;
        RECT 83.74 0 83.91 3.38 ;
        RECT 82.78 0 82.95 3.38 ;
        RECT 80.86 0 81.135 2.89 ;
        RECT 80.86 0 81.03 3.38 ;
        RECT 77.86 0 78.03 2.225 ;
        RECT 76.875 0 77.045 2.225 ;
        RECT 74.13 0 74.3 2.225 ;
        RECT 64.33 0 73.07 2.88 ;
        RECT 72.3 0 72.47 3.38 ;
        RECT 71.36 0 71.53 3.38 ;
        RECT 70.4 0 70.57 3.38 ;
        RECT 69.355 0 69.55 2.89 ;
        RECT 68.48 0 68.65 3.38 ;
        RECT 67.52 0 67.69 3.38 ;
        RECT 65.6 0 65.875 2.89 ;
        RECT 65.6 0 65.77 3.38 ;
        RECT 62.6 0 62.77 2.225 ;
        RECT 61.615 0 61.785 2.225 ;
        RECT 58.87 0 59.04 2.225 ;
        RECT 49.07 0 57.81 2.88 ;
        RECT 57.04 0 57.21 3.38 ;
        RECT 56.1 0 56.27 3.38 ;
        RECT 55.14 0 55.31 3.38 ;
        RECT 54.095 0 54.29 2.89 ;
        RECT 53.22 0 53.39 3.38 ;
        RECT 52.26 0 52.43 3.38 ;
        RECT 50.34 0 50.615 2.89 ;
        RECT 50.34 0 50.51 3.38 ;
        RECT 47.34 0 47.51 2.225 ;
        RECT 46.355 0 46.525 2.225 ;
        RECT 43.61 0 43.78 2.225 ;
        RECT 33.81 0 42.55 2.88 ;
        RECT 41.78 0 41.95 3.38 ;
        RECT 40.84 0 41.01 3.38 ;
        RECT 39.88 0 40.05 3.38 ;
        RECT 38.835 0 39.03 2.89 ;
        RECT 37.96 0 38.13 3.38 ;
        RECT 37 0 37.17 3.38 ;
        RECT 35.08 0 35.355 2.89 ;
        RECT 35.08 0 35.25 3.38 ;
        RECT 32.08 0 32.25 2.225 ;
        RECT 31.095 0 31.265 2.225 ;
        RECT 28.35 0 28.52 2.225 ;
        RECT 18.55 0 27.29 2.88 ;
        RECT 26.52 0 26.69 3.38 ;
        RECT 25.58 0 25.75 3.38 ;
        RECT 24.62 0 24.79 3.38 ;
        RECT 23.575 0 23.77 2.89 ;
        RECT 22.7 0 22.87 3.38 ;
        RECT 21.74 0 21.91 3.38 ;
        RECT 19.82 0 20.095 2.89 ;
        RECT 19.82 0 19.99 3.38 ;
        RECT 0.005 10.865 94.1 12.465 ;
        RECT 93.125 10.24 93.295 12.465 ;
        RECT 92.135 10.24 92.305 12.465 ;
        RECT 89.39 10.24 89.56 12.465 ;
        RECT 83.755 10.24 83.925 12.465 ;
        RECT 77.865 10.24 78.035 12.465 ;
        RECT 76.875 10.24 77.045 12.465 ;
        RECT 74.13 10.24 74.3 12.465 ;
        RECT 68.495 10.24 68.665 12.465 ;
        RECT 62.605 10.24 62.775 12.465 ;
        RECT 61.615 10.24 61.785 12.465 ;
        RECT 58.87 10.24 59.04 12.465 ;
        RECT 53.235 10.24 53.405 12.465 ;
        RECT 47.345 10.24 47.515 12.465 ;
        RECT 46.355 10.24 46.525 12.465 ;
        RECT 43.61 10.24 43.78 12.465 ;
        RECT 37.975 10.24 38.145 12.465 ;
        RECT 32.085 10.24 32.255 12.465 ;
        RECT 31.095 10.24 31.265 12.465 ;
        RECT 28.35 10.24 28.52 12.465 ;
        RECT 22.715 10.24 22.885 12.465 ;
        RECT 15.22 10.24 15.39 12.465 ;
        RECT 84.77 8.37 84.94 10.32 ;
        RECT 84.71 10.15 84.88 10.6 ;
        RECT 84.71 7.31 84.88 8.54 ;
        RECT 81.455 3.63 81.78 3.88 ;
        RECT 81.505 3.63 81.775 4.04 ;
        RECT 81.5 3.63 81.775 3.98 ;
        RECT 81.475 3.63 81.775 3.945 ;
        RECT 80.125 3.62 81.49 3.715 ;
        RECT 81.455 3.63 81.775 3.91 ;
        RECT 81.45 3.63 81.78 3.875 ;
        RECT 81.44 3.63 81.78 3.87 ;
        RECT 81.435 3.63 81.78 3.855 ;
        RECT 80.125 3.585 81.435 3.715 ;
        RECT 81.42 3.63 81.78 3.85 ;
        RECT 81.405 3.63 81.78 3.83 ;
        RECT 81.385 3.63 81.78 3.815 ;
        RECT 81.37 3.63 81.78 3.785 ;
        RECT 81.35 3.63 81.78 3.775 ;
        RECT 81.335 3.63 81.78 3.76 ;
        RECT 81.3 3.63 81.78 3.745 ;
        RECT 81.205 3.63 81.78 3.735 ;
        RECT 80.125 3.565 81.235 3.715 ;
        RECT 80.91 3.63 81.78 3.725 ;
        RECT 80.125 3.555 81.145 3.715 ;
        RECT 80.125 3.55 81.105 3.715 ;
        RECT 80.125 3.545 81.09 3.715 ;
        RECT 80.125 3.535 81.065 3.715 ;
        RECT 80.125 3.535 80.755 3.72 ;
        RECT 80.125 3.535 80.72 3.73 ;
        RECT 80.125 3.535 80.68 3.74 ;
        RECT 80.125 3.535 80.565 3.745 ;
        RECT 80.125 3.535 80.55 3.765 ;
        RECT 80.125 3.535 80.47 3.77 ;
        RECT 80.125 3.535 80.445 3.795 ;
        RECT 80.125 3.535 80.42 3.815 ;
        RECT 80.125 3.535 80.415 3.83 ;
        RECT 80.125 3.535 80.41 3.85 ;
        RECT 80.125 3.535 80.405 3.855 ;
        RECT 80.125 3.535 80.4 3.87 ;
        RECT 80.115 3.95 80.395 4.05 ;
        RECT 80.125 3.535 80.395 4.05 ;
        RECT 69.51 8.37 69.68 10.32 ;
        RECT 69.45 10.15 69.62 10.6 ;
        RECT 69.45 7.31 69.62 8.54 ;
        RECT 66.195 3.63 66.52 3.88 ;
        RECT 66.245 3.63 66.515 4.04 ;
        RECT 66.24 3.63 66.515 3.98 ;
        RECT 66.215 3.63 66.515 3.945 ;
        RECT 64.865 3.62 66.23 3.715 ;
        RECT 66.195 3.63 66.515 3.91 ;
        RECT 66.19 3.63 66.52 3.875 ;
        RECT 66.18 3.63 66.52 3.87 ;
        RECT 66.175 3.63 66.52 3.855 ;
        RECT 64.865 3.585 66.175 3.715 ;
        RECT 66.16 3.63 66.52 3.85 ;
        RECT 66.145 3.63 66.52 3.83 ;
        RECT 66.125 3.63 66.52 3.815 ;
        RECT 66.11 3.63 66.52 3.785 ;
        RECT 66.09 3.63 66.52 3.775 ;
        RECT 66.075 3.63 66.52 3.76 ;
        RECT 66.04 3.63 66.52 3.745 ;
        RECT 65.945 3.63 66.52 3.735 ;
        RECT 64.865 3.565 65.975 3.715 ;
        RECT 65.65 3.63 66.52 3.725 ;
        RECT 64.865 3.555 65.885 3.715 ;
        RECT 64.865 3.55 65.845 3.715 ;
        RECT 64.865 3.545 65.83 3.715 ;
        RECT 64.865 3.535 65.805 3.715 ;
        RECT 64.865 3.535 65.495 3.72 ;
        RECT 64.865 3.535 65.46 3.73 ;
        RECT 64.865 3.535 65.42 3.74 ;
        RECT 64.865 3.535 65.305 3.745 ;
        RECT 64.865 3.535 65.29 3.765 ;
        RECT 64.865 3.535 65.21 3.77 ;
        RECT 64.865 3.535 65.185 3.795 ;
        RECT 64.865 3.535 65.16 3.815 ;
        RECT 64.865 3.535 65.155 3.83 ;
        RECT 64.865 3.535 65.15 3.85 ;
        RECT 64.865 3.535 65.145 3.855 ;
        RECT 64.865 3.535 65.14 3.87 ;
        RECT 64.855 3.95 65.135 4.05 ;
        RECT 64.865 3.535 65.135 4.05 ;
        RECT 54.25 8.37 54.42 10.32 ;
        RECT 54.19 10.15 54.36 10.6 ;
        RECT 54.19 7.31 54.36 8.54 ;
        RECT 50.935 3.63 51.26 3.88 ;
        RECT 50.985 3.63 51.255 4.04 ;
        RECT 50.98 3.63 51.255 3.98 ;
        RECT 50.955 3.63 51.255 3.945 ;
        RECT 49.605 3.62 50.97 3.715 ;
        RECT 50.935 3.63 51.255 3.91 ;
        RECT 50.93 3.63 51.26 3.875 ;
        RECT 50.92 3.63 51.26 3.87 ;
        RECT 50.915 3.63 51.26 3.855 ;
        RECT 49.605 3.585 50.915 3.715 ;
        RECT 50.9 3.63 51.26 3.85 ;
        RECT 50.885 3.63 51.26 3.83 ;
        RECT 50.865 3.63 51.26 3.815 ;
        RECT 50.85 3.63 51.26 3.785 ;
        RECT 50.83 3.63 51.26 3.775 ;
        RECT 50.815 3.63 51.26 3.76 ;
        RECT 50.78 3.63 51.26 3.745 ;
        RECT 50.685 3.63 51.26 3.735 ;
        RECT 49.605 3.565 50.715 3.715 ;
        RECT 50.39 3.63 51.26 3.725 ;
        RECT 49.605 3.555 50.625 3.715 ;
        RECT 49.605 3.55 50.585 3.715 ;
        RECT 49.605 3.545 50.57 3.715 ;
        RECT 49.605 3.535 50.545 3.715 ;
        RECT 49.605 3.535 50.235 3.72 ;
        RECT 49.605 3.535 50.2 3.73 ;
        RECT 49.605 3.535 50.16 3.74 ;
        RECT 49.605 3.535 50.045 3.745 ;
        RECT 49.605 3.535 50.03 3.765 ;
        RECT 49.605 3.535 49.95 3.77 ;
        RECT 49.605 3.535 49.925 3.795 ;
        RECT 49.605 3.535 49.9 3.815 ;
        RECT 49.605 3.535 49.895 3.83 ;
        RECT 49.605 3.535 49.89 3.85 ;
        RECT 49.605 3.535 49.885 3.855 ;
        RECT 49.605 3.535 49.88 3.87 ;
        RECT 49.595 3.95 49.875 4.05 ;
        RECT 49.605 3.535 49.875 4.05 ;
        RECT 38.99 8.37 39.16 10.32 ;
        RECT 38.93 10.15 39.1 10.6 ;
        RECT 38.93 7.31 39.1 8.54 ;
        RECT 35.675 3.63 36 3.88 ;
        RECT 35.725 3.63 35.995 4.04 ;
        RECT 35.72 3.63 35.995 3.98 ;
        RECT 35.695 3.63 35.995 3.945 ;
        RECT 34.345 3.62 35.71 3.715 ;
        RECT 35.675 3.63 35.995 3.91 ;
        RECT 35.67 3.63 36 3.875 ;
        RECT 35.66 3.63 36 3.87 ;
        RECT 35.655 3.63 36 3.855 ;
        RECT 34.345 3.585 35.655 3.715 ;
        RECT 35.64 3.63 36 3.85 ;
        RECT 35.625 3.63 36 3.83 ;
        RECT 35.605 3.63 36 3.815 ;
        RECT 35.59 3.63 36 3.785 ;
        RECT 35.57 3.63 36 3.775 ;
        RECT 35.555 3.63 36 3.76 ;
        RECT 35.52 3.63 36 3.745 ;
        RECT 35.425 3.63 36 3.735 ;
        RECT 34.345 3.565 35.455 3.715 ;
        RECT 35.13 3.63 36 3.725 ;
        RECT 34.345 3.555 35.365 3.715 ;
        RECT 34.345 3.55 35.325 3.715 ;
        RECT 34.345 3.545 35.31 3.715 ;
        RECT 34.345 3.535 35.285 3.715 ;
        RECT 34.345 3.535 34.975 3.72 ;
        RECT 34.345 3.535 34.94 3.73 ;
        RECT 34.345 3.535 34.9 3.74 ;
        RECT 34.345 3.535 34.785 3.745 ;
        RECT 34.345 3.535 34.77 3.765 ;
        RECT 34.345 3.535 34.69 3.77 ;
        RECT 34.345 3.535 34.665 3.795 ;
        RECT 34.345 3.535 34.64 3.815 ;
        RECT 34.345 3.535 34.635 3.83 ;
        RECT 34.345 3.535 34.63 3.85 ;
        RECT 34.345 3.535 34.625 3.855 ;
        RECT 34.345 3.535 34.62 3.87 ;
        RECT 34.335 3.95 34.615 4.05 ;
        RECT 34.345 3.535 34.615 4.05 ;
        RECT 23.73 8.37 23.9 10.32 ;
        RECT 23.67 10.15 23.84 10.6 ;
        RECT 23.67 7.31 23.84 8.54 ;
        RECT 20.415 3.63 20.74 3.88 ;
        RECT 20.465 3.63 20.735 4.04 ;
        RECT 20.46 3.63 20.735 3.98 ;
        RECT 20.435 3.63 20.735 3.945 ;
        RECT 19.085 3.62 20.45 3.715 ;
        RECT 20.415 3.63 20.735 3.91 ;
        RECT 20.41 3.63 20.74 3.875 ;
        RECT 20.4 3.63 20.74 3.87 ;
        RECT 20.395 3.63 20.74 3.855 ;
        RECT 19.085 3.585 20.395 3.715 ;
        RECT 20.38 3.63 20.74 3.85 ;
        RECT 20.365 3.63 20.74 3.83 ;
        RECT 20.345 3.63 20.74 3.815 ;
        RECT 20.33 3.63 20.74 3.785 ;
        RECT 20.31 3.63 20.74 3.775 ;
        RECT 20.295 3.63 20.74 3.76 ;
        RECT 20.26 3.63 20.74 3.745 ;
        RECT 20.165 3.63 20.74 3.735 ;
        RECT 19.085 3.565 20.195 3.715 ;
        RECT 19.87 3.63 20.74 3.725 ;
        RECT 19.085 3.555 20.105 3.715 ;
        RECT 19.085 3.55 20.065 3.715 ;
        RECT 19.085 3.545 20.05 3.715 ;
        RECT 19.085 3.535 20.025 3.715 ;
        RECT 19.085 3.535 19.715 3.72 ;
        RECT 19.085 3.535 19.68 3.73 ;
        RECT 19.085 3.535 19.64 3.74 ;
        RECT 19.085 3.535 19.525 3.745 ;
        RECT 19.085 3.535 19.51 3.765 ;
        RECT 19.085 3.535 19.43 3.77 ;
        RECT 19.085 3.535 19.405 3.795 ;
        RECT 19.085 3.535 19.38 3.815 ;
        RECT 19.085 3.535 19.375 3.83 ;
        RECT 19.085 3.535 19.37 3.85 ;
        RECT 19.085 3.535 19.365 3.855 ;
        RECT 19.085 3.535 19.36 3.87 ;
        RECT 19.075 3.95 19.355 4.05 ;
        RECT 19.085 3.535 19.355 4.05 ;
      LAYER met1 ;
        RECT 0.005 0 94.1 1.6 ;
        RECT 79.59 0 88.33 3.035 ;
        RECT 64.33 0 73.07 3.035 ;
        RECT 49.07 0 57.81 3.035 ;
        RECT 33.81 0 42.55 3.035 ;
        RECT 18.55 0 27.29 3.035 ;
        RECT 0.005 10.865 94.1 12.465 ;
        RECT 84.71 8.58 85 8.81 ;
        RECT 84.535 8.61 85 8.78 ;
        RECT 84.535 8.605 84.705 12.465 ;
        RECT 69.45 8.58 69.74 8.81 ;
        RECT 69.275 8.61 69.74 8.78 ;
        RECT 69.275 8.605 69.445 12.465 ;
        RECT 54.19 8.58 54.48 8.81 ;
        RECT 54.015 8.61 54.48 8.78 ;
        RECT 54.015 8.605 54.185 12.465 ;
        RECT 38.93 8.58 39.22 8.81 ;
        RECT 38.755 8.61 39.22 8.78 ;
        RECT 38.755 8.605 38.925 12.465 ;
        RECT 23.67 8.58 23.96 8.81 ;
        RECT 23.495 8.61 23.96 8.78 ;
        RECT 23.495 8.605 23.665 12.465 ;
        RECT 81.615 3.625 81.875 3.885 ;
        RECT 81.475 3.63 81.82 3.93 ;
        RECT 81.475 3.63 81.775 3.945 ;
        RECT 81.455 3.63 81.82 3.91 ;
        RECT 66.355 3.625 66.615 3.885 ;
        RECT 66.215 3.63 66.56 3.93 ;
        RECT 66.215 3.63 66.515 3.945 ;
        RECT 66.195 3.63 66.56 3.91 ;
        RECT 51.095 3.625 51.355 3.885 ;
        RECT 50.955 3.63 51.3 3.93 ;
        RECT 50.955 3.63 51.255 3.945 ;
        RECT 50.935 3.63 51.3 3.91 ;
        RECT 35.835 3.625 36.095 3.885 ;
        RECT 35.695 3.63 36.04 3.93 ;
        RECT 35.695 3.63 35.995 3.945 ;
        RECT 35.675 3.63 36.04 3.91 ;
        RECT 20.575 3.625 20.835 3.885 ;
        RECT 20.435 3.63 20.78 3.93 ;
        RECT 20.435 3.63 20.735 3.945 ;
        RECT 20.415 3.63 20.78 3.91 ;
      LAYER via1 ;
        RECT 20.63 3.68 20.78 3.83 ;
        RECT 20.675 2.35 20.825 2.5 ;
        RECT 35.89 3.68 36.04 3.83 ;
        RECT 35.935 2.35 36.085 2.5 ;
        RECT 51.15 3.68 51.3 3.83 ;
        RECT 51.195 2.35 51.345 2.5 ;
        RECT 66.41 3.68 66.56 3.83 ;
        RECT 66.455 2.35 66.605 2.5 ;
        RECT 81.67 3.68 81.82 3.83 ;
        RECT 81.715 2.35 81.865 2.5 ;
      LAYER via2 ;
        RECT 20.525 3.775 20.725 3.975 ;
        RECT 35.785 3.775 35.985 3.975 ;
        RECT 51.045 3.775 51.245 3.975 ;
        RECT 66.305 3.775 66.505 3.975 ;
        RECT 81.565 3.775 81.765 3.975 ;
      LAYER mcon ;
        RECT 15.3 10.9 15.47 11.07 ;
        RECT 15.98 10.9 16.15 11.07 ;
        RECT 16.66 10.9 16.83 11.07 ;
        RECT 17.34 10.9 17.51 11.07 ;
        RECT 18.695 2.71 18.865 2.88 ;
        RECT 19.155 2.71 19.325 2.88 ;
        RECT 19.615 2.71 19.785 2.88 ;
        RECT 20.075 2.71 20.245 2.88 ;
        RECT 20.525 3.71 20.695 3.88 ;
        RECT 20.535 2.71 20.705 2.88 ;
        RECT 20.995 2.71 21.165 2.88 ;
        RECT 21.455 2.71 21.625 2.88 ;
        RECT 21.915 2.71 22.085 2.88 ;
        RECT 22.375 2.71 22.545 2.88 ;
        RECT 22.795 10.9 22.965 11.07 ;
        RECT 22.835 2.71 23.005 2.88 ;
        RECT 23.295 2.71 23.465 2.88 ;
        RECT 23.475 10.9 23.645 11.07 ;
        RECT 23.73 8.61 23.9 8.78 ;
        RECT 23.755 2.71 23.925 2.88 ;
        RECT 24.155 10.9 24.325 11.07 ;
        RECT 24.215 2.71 24.385 2.88 ;
        RECT 24.675 2.71 24.845 2.88 ;
        RECT 24.835 10.9 25.005 11.07 ;
        RECT 25.135 2.71 25.305 2.88 ;
        RECT 25.595 2.71 25.765 2.88 ;
        RECT 26.055 2.71 26.225 2.88 ;
        RECT 26.515 2.71 26.685 2.88 ;
        RECT 26.975 2.71 27.145 2.88 ;
        RECT 28.43 10.9 28.6 11.07 ;
        RECT 28.43 1.395 28.6 1.565 ;
        RECT 29.11 10.9 29.28 11.07 ;
        RECT 29.11 1.395 29.28 1.565 ;
        RECT 29.79 10.9 29.96 11.07 ;
        RECT 29.79 1.395 29.96 1.565 ;
        RECT 30.47 10.9 30.64 11.07 ;
        RECT 30.47 1.395 30.64 1.565 ;
        RECT 31.175 10.9 31.345 11.07 ;
        RECT 31.175 1.395 31.345 1.565 ;
        RECT 32.16 1.395 32.33 1.565 ;
        RECT 32.165 10.9 32.335 11.07 ;
        RECT 33.955 2.71 34.125 2.88 ;
        RECT 34.415 2.71 34.585 2.88 ;
        RECT 34.875 2.71 35.045 2.88 ;
        RECT 35.335 2.71 35.505 2.88 ;
        RECT 35.785 3.71 35.955 3.88 ;
        RECT 35.795 2.71 35.965 2.88 ;
        RECT 36.255 2.71 36.425 2.88 ;
        RECT 36.715 2.71 36.885 2.88 ;
        RECT 37.175 2.71 37.345 2.88 ;
        RECT 37.635 2.71 37.805 2.88 ;
        RECT 38.055 10.9 38.225 11.07 ;
        RECT 38.095 2.71 38.265 2.88 ;
        RECT 38.555 2.71 38.725 2.88 ;
        RECT 38.735 10.9 38.905 11.07 ;
        RECT 38.99 8.61 39.16 8.78 ;
        RECT 39.015 2.71 39.185 2.88 ;
        RECT 39.415 10.9 39.585 11.07 ;
        RECT 39.475 2.71 39.645 2.88 ;
        RECT 39.935 2.71 40.105 2.88 ;
        RECT 40.095 10.9 40.265 11.07 ;
        RECT 40.395 2.71 40.565 2.88 ;
        RECT 40.855 2.71 41.025 2.88 ;
        RECT 41.315 2.71 41.485 2.88 ;
        RECT 41.775 2.71 41.945 2.88 ;
        RECT 42.235 2.71 42.405 2.88 ;
        RECT 43.69 10.9 43.86 11.07 ;
        RECT 43.69 1.395 43.86 1.565 ;
        RECT 44.37 10.9 44.54 11.07 ;
        RECT 44.37 1.395 44.54 1.565 ;
        RECT 45.05 10.9 45.22 11.07 ;
        RECT 45.05 1.395 45.22 1.565 ;
        RECT 45.73 10.9 45.9 11.07 ;
        RECT 45.73 1.395 45.9 1.565 ;
        RECT 46.435 10.9 46.605 11.07 ;
        RECT 46.435 1.395 46.605 1.565 ;
        RECT 47.42 1.395 47.59 1.565 ;
        RECT 47.425 10.9 47.595 11.07 ;
        RECT 49.215 2.71 49.385 2.88 ;
        RECT 49.675 2.71 49.845 2.88 ;
        RECT 50.135 2.71 50.305 2.88 ;
        RECT 50.595 2.71 50.765 2.88 ;
        RECT 51.045 3.71 51.215 3.88 ;
        RECT 51.055 2.71 51.225 2.88 ;
        RECT 51.515 2.71 51.685 2.88 ;
        RECT 51.975 2.71 52.145 2.88 ;
        RECT 52.435 2.71 52.605 2.88 ;
        RECT 52.895 2.71 53.065 2.88 ;
        RECT 53.315 10.9 53.485 11.07 ;
        RECT 53.355 2.71 53.525 2.88 ;
        RECT 53.815 2.71 53.985 2.88 ;
        RECT 53.995 10.9 54.165 11.07 ;
        RECT 54.25 8.61 54.42 8.78 ;
        RECT 54.275 2.71 54.445 2.88 ;
        RECT 54.675 10.9 54.845 11.07 ;
        RECT 54.735 2.71 54.905 2.88 ;
        RECT 55.195 2.71 55.365 2.88 ;
        RECT 55.355 10.9 55.525 11.07 ;
        RECT 55.655 2.71 55.825 2.88 ;
        RECT 56.115 2.71 56.285 2.88 ;
        RECT 56.575 2.71 56.745 2.88 ;
        RECT 57.035 2.71 57.205 2.88 ;
        RECT 57.495 2.71 57.665 2.88 ;
        RECT 58.95 10.9 59.12 11.07 ;
        RECT 58.95 1.395 59.12 1.565 ;
        RECT 59.63 10.9 59.8 11.07 ;
        RECT 59.63 1.395 59.8 1.565 ;
        RECT 60.31 10.9 60.48 11.07 ;
        RECT 60.31 1.395 60.48 1.565 ;
        RECT 60.99 10.9 61.16 11.07 ;
        RECT 60.99 1.395 61.16 1.565 ;
        RECT 61.695 10.9 61.865 11.07 ;
        RECT 61.695 1.395 61.865 1.565 ;
        RECT 62.68 1.395 62.85 1.565 ;
        RECT 62.685 10.9 62.855 11.07 ;
        RECT 64.475 2.71 64.645 2.88 ;
        RECT 64.935 2.71 65.105 2.88 ;
        RECT 65.395 2.71 65.565 2.88 ;
        RECT 65.855 2.71 66.025 2.88 ;
        RECT 66.305 3.71 66.475 3.88 ;
        RECT 66.315 2.71 66.485 2.88 ;
        RECT 66.775 2.71 66.945 2.88 ;
        RECT 67.235 2.71 67.405 2.88 ;
        RECT 67.695 2.71 67.865 2.88 ;
        RECT 68.155 2.71 68.325 2.88 ;
        RECT 68.575 10.9 68.745 11.07 ;
        RECT 68.615 2.71 68.785 2.88 ;
        RECT 69.075 2.71 69.245 2.88 ;
        RECT 69.255 10.9 69.425 11.07 ;
        RECT 69.51 8.61 69.68 8.78 ;
        RECT 69.535 2.71 69.705 2.88 ;
        RECT 69.935 10.9 70.105 11.07 ;
        RECT 69.995 2.71 70.165 2.88 ;
        RECT 70.455 2.71 70.625 2.88 ;
        RECT 70.615 10.9 70.785 11.07 ;
        RECT 70.915 2.71 71.085 2.88 ;
        RECT 71.375 2.71 71.545 2.88 ;
        RECT 71.835 2.71 72.005 2.88 ;
        RECT 72.295 2.71 72.465 2.88 ;
        RECT 72.755 2.71 72.925 2.88 ;
        RECT 74.21 10.9 74.38 11.07 ;
        RECT 74.21 1.395 74.38 1.565 ;
        RECT 74.89 10.9 75.06 11.07 ;
        RECT 74.89 1.395 75.06 1.565 ;
        RECT 75.57 10.9 75.74 11.07 ;
        RECT 75.57 1.395 75.74 1.565 ;
        RECT 76.25 10.9 76.42 11.07 ;
        RECT 76.25 1.395 76.42 1.565 ;
        RECT 76.955 10.9 77.125 11.07 ;
        RECT 76.955 1.395 77.125 1.565 ;
        RECT 77.94 1.395 78.11 1.565 ;
        RECT 77.945 10.9 78.115 11.07 ;
        RECT 79.735 2.71 79.905 2.88 ;
        RECT 80.195 2.71 80.365 2.88 ;
        RECT 80.655 2.71 80.825 2.88 ;
        RECT 81.115 2.71 81.285 2.88 ;
        RECT 81.565 3.71 81.735 3.88 ;
        RECT 81.575 2.71 81.745 2.88 ;
        RECT 82.035 2.71 82.205 2.88 ;
        RECT 82.495 2.71 82.665 2.88 ;
        RECT 82.955 2.71 83.125 2.88 ;
        RECT 83.415 2.71 83.585 2.88 ;
        RECT 83.835 10.9 84.005 11.07 ;
        RECT 83.875 2.71 84.045 2.88 ;
        RECT 84.335 2.71 84.505 2.88 ;
        RECT 84.515 10.9 84.685 11.07 ;
        RECT 84.77 8.61 84.94 8.78 ;
        RECT 84.795 2.71 84.965 2.88 ;
        RECT 85.195 10.9 85.365 11.07 ;
        RECT 85.255 2.71 85.425 2.88 ;
        RECT 85.715 2.71 85.885 2.88 ;
        RECT 85.875 10.9 86.045 11.07 ;
        RECT 86.175 2.71 86.345 2.88 ;
        RECT 86.635 2.71 86.805 2.88 ;
        RECT 87.095 2.71 87.265 2.88 ;
        RECT 87.555 2.71 87.725 2.88 ;
        RECT 88.015 2.71 88.185 2.88 ;
        RECT 89.47 10.9 89.64 11.07 ;
        RECT 89.47 1.395 89.64 1.565 ;
        RECT 90.15 10.9 90.32 11.07 ;
        RECT 90.15 1.395 90.32 1.565 ;
        RECT 90.83 10.9 91 11.07 ;
        RECT 90.83 1.395 91 1.565 ;
        RECT 91.51 10.9 91.68 11.07 ;
        RECT 91.51 1.395 91.68 1.565 ;
        RECT 92.215 10.9 92.385 11.07 ;
        RECT 92.215 1.395 92.385 1.565 ;
        RECT 93.2 1.395 93.37 1.565 ;
        RECT 93.205 10.9 93.375 11.07 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 88.705 3.97 89.105 4.355 ;
      RECT 88.71 2.245 89.04 4.355 ;
      RECT 82.7 2.245 83.03 3.88 ;
      RECT 82.7 2.245 89.04 2.575 ;
      RECT 85.04 9.345 85.41 9.715 ;
      RECT 85.075 5.565 85.375 9.715 ;
      RECT 80.885 6.525 85.375 6.86 ;
      RECT 84.025 5.565 85.375 6.86 ;
      RECT 80.885 5.435 81.19 6.86 ;
      RECT 84.065 3.15 84.365 6.86 ;
      RECT 80.885 3.73 81.185 6.86 ;
      RECT 84.02 4.055 84.365 4.785 ;
      RECT 80.78 3.31 81.11 4.04 ;
      RECT 83.66 3.15 84.39 3.48 ;
      RECT 73.445 3.97 73.845 4.355 ;
      RECT 73.45 2.245 73.78 4.355 ;
      RECT 67.44 2.245 67.77 3.88 ;
      RECT 67.44 2.245 73.78 2.575 ;
      RECT 69.78 9.345 70.15 9.715 ;
      RECT 69.815 5.565 70.115 9.715 ;
      RECT 65.625 6.525 70.115 6.86 ;
      RECT 68.765 5.565 70.115 6.86 ;
      RECT 65.625 5.435 65.93 6.86 ;
      RECT 68.805 3.15 69.105 6.86 ;
      RECT 65.625 3.73 65.925 6.86 ;
      RECT 68.76 4.055 69.105 4.785 ;
      RECT 65.52 3.31 65.85 4.04 ;
      RECT 68.4 3.15 69.13 3.48 ;
      RECT 58.185 3.97 58.585 4.355 ;
      RECT 58.19 2.245 58.52 4.355 ;
      RECT 52.18 2.245 52.51 3.88 ;
      RECT 52.18 2.245 58.52 2.575 ;
      RECT 54.52 9.345 54.89 9.715 ;
      RECT 54.555 5.565 54.855 9.715 ;
      RECT 50.365 6.525 54.855 6.86 ;
      RECT 53.505 5.565 54.855 6.86 ;
      RECT 50.365 5.435 50.67 6.86 ;
      RECT 53.545 3.15 53.845 6.86 ;
      RECT 50.365 3.73 50.665 6.86 ;
      RECT 53.5 4.055 53.845 4.785 ;
      RECT 50.26 3.31 50.59 4.04 ;
      RECT 53.14 3.15 53.87 3.48 ;
      RECT 42.925 3.97 43.325 4.355 ;
      RECT 42.93 2.245 43.26 4.355 ;
      RECT 36.92 2.245 37.25 3.88 ;
      RECT 36.92 2.245 43.26 2.575 ;
      RECT 39.26 9.345 39.63 9.715 ;
      RECT 39.295 5.565 39.595 9.715 ;
      RECT 35.105 6.525 39.595 6.86 ;
      RECT 38.245 5.565 39.595 6.86 ;
      RECT 35.105 5.435 35.41 6.86 ;
      RECT 38.285 3.15 38.585 6.86 ;
      RECT 35.105 3.73 35.405 6.86 ;
      RECT 38.24 4.055 38.585 4.785 ;
      RECT 35 3.31 35.33 4.04 ;
      RECT 37.88 3.15 38.61 3.48 ;
      RECT 27.665 3.97 28.065 4.355 ;
      RECT 27.67 2.245 28 4.355 ;
      RECT 21.66 2.245 21.99 3.88 ;
      RECT 21.66 2.245 28 2.575 ;
      RECT 24 9.345 24.37 9.715 ;
      RECT 24.035 5.565 24.335 9.715 ;
      RECT 19.845 6.525 24.335 6.86 ;
      RECT 22.985 5.565 24.335 6.86 ;
      RECT 19.845 5.435 20.15 6.86 ;
      RECT 23.025 3.15 23.325 6.86 ;
      RECT 19.845 3.73 20.145 6.86 ;
      RECT 22.98 4.055 23.325 4.785 ;
      RECT 19.74 3.31 20.07 4.04 ;
      RECT 22.62 3.15 23.35 3.48 ;
      RECT 93.455 7.205 93.835 12.465 ;
      RECT 87.14 3.31 87.47 4.04 ;
      RECT 85.94 4.175 86.27 4.905 ;
      RECT 85.1 3.15 85.83 3.48 ;
      RECT 78.195 7.205 78.575 12.465 ;
      RECT 71.88 3.31 72.21 4.04 ;
      RECT 70.68 4.175 71.01 4.905 ;
      RECT 69.84 3.15 70.57 3.48 ;
      RECT 62.935 7.205 63.315 12.465 ;
      RECT 56.62 3.31 56.95 4.04 ;
      RECT 55.42 4.175 55.75 4.905 ;
      RECT 54.58 3.15 55.31 3.48 ;
      RECT 47.675 7.205 48.055 12.465 ;
      RECT 41.36 3.31 41.69 4.04 ;
      RECT 40.16 4.175 40.49 4.905 ;
      RECT 39.32 3.15 40.05 3.48 ;
      RECT 32.415 7.205 32.795 12.465 ;
      RECT 26.1 3.31 26.43 4.04 ;
      RECT 24.9 4.175 25.23 4.905 ;
      RECT 24.06 3.15 24.79 3.48 ;
    LAYER via2 ;
      RECT 93.545 7.295 93.745 7.495 ;
      RECT 88.81 4.075 89.01 4.275 ;
      RECT 87.205 3.775 87.405 3.975 ;
      RECT 86.005 4.335 86.205 4.535 ;
      RECT 85.165 3.215 85.365 3.415 ;
      RECT 85.125 9.43 85.325 9.63 ;
      RECT 84.085 4.12 84.285 4.32 ;
      RECT 83.725 3.215 83.925 3.415 ;
      RECT 82.765 3.215 82.965 3.415 ;
      RECT 80.845 3.775 81.045 3.975 ;
      RECT 78.285 7.295 78.485 7.495 ;
      RECT 73.55 4.075 73.75 4.275 ;
      RECT 71.945 3.775 72.145 3.975 ;
      RECT 70.745 4.335 70.945 4.535 ;
      RECT 69.905 3.215 70.105 3.415 ;
      RECT 69.865 9.43 70.065 9.63 ;
      RECT 68.825 4.12 69.025 4.32 ;
      RECT 68.465 3.215 68.665 3.415 ;
      RECT 67.505 3.215 67.705 3.415 ;
      RECT 65.585 3.775 65.785 3.975 ;
      RECT 63.025 7.295 63.225 7.495 ;
      RECT 58.29 4.075 58.49 4.275 ;
      RECT 56.685 3.775 56.885 3.975 ;
      RECT 55.485 4.335 55.685 4.535 ;
      RECT 54.645 3.215 54.845 3.415 ;
      RECT 54.605 9.43 54.805 9.63 ;
      RECT 53.565 4.12 53.765 4.32 ;
      RECT 53.205 3.215 53.405 3.415 ;
      RECT 52.245 3.215 52.445 3.415 ;
      RECT 50.325 3.775 50.525 3.975 ;
      RECT 47.765 7.295 47.965 7.495 ;
      RECT 43.03 4.075 43.23 4.275 ;
      RECT 41.425 3.775 41.625 3.975 ;
      RECT 40.225 4.335 40.425 4.535 ;
      RECT 39.385 3.215 39.585 3.415 ;
      RECT 39.345 9.43 39.545 9.63 ;
      RECT 38.305 4.12 38.505 4.32 ;
      RECT 37.945 3.215 38.145 3.415 ;
      RECT 36.985 3.215 37.185 3.415 ;
      RECT 35.065 3.775 35.265 3.975 ;
      RECT 32.505 7.295 32.705 7.495 ;
      RECT 27.77 4.075 27.97 4.275 ;
      RECT 26.165 3.775 26.365 3.975 ;
      RECT 24.965 4.335 25.165 4.535 ;
      RECT 24.125 3.215 24.325 3.415 ;
      RECT 24.085 9.43 24.285 9.63 ;
      RECT 23.045 4.12 23.245 4.32 ;
      RECT 22.685 3.215 22.885 3.415 ;
      RECT 21.725 3.215 21.925 3.415 ;
      RECT 19.805 3.775 20.005 3.975 ;
    LAYER met2 ;
      RECT 16.23 10.69 93.73 10.86 ;
      RECT 93.56 9.565 93.73 10.86 ;
      RECT 16.23 8.545 16.4 10.86 ;
      RECT 93.53 9.565 93.88 9.915 ;
      RECT 16.17 8.545 16.46 8.895 ;
      RECT 90.37 8.51 90.69 8.835 ;
      RECT 90.4 7.985 90.57 8.835 ;
      RECT 90.4 7.985 90.575 8.335 ;
      RECT 90.4 7.985 91.375 8.16 ;
      RECT 91.2 3.26 91.375 8.16 ;
      RECT 91.145 3.26 91.495 3.61 ;
      RECT 91.17 8.945 91.495 9.27 ;
      RECT 90.055 9.035 91.495 9.205 ;
      RECT 90.055 3.69 90.215 9.205 ;
      RECT 90.37 3.66 90.69 3.98 ;
      RECT 90.055 3.69 90.69 3.86 ;
      RECT 88.72 4 89.105 4.35 ;
      RECT 88.71 4.065 89.105 4.265 ;
      RECT 88.855 3.995 89.025 4.35 ;
      RECT 87.165 3.735 87.445 4.015 ;
      RECT 87.16 3.735 87.445 3.968 ;
      RECT 87.14 3.735 87.445 3.945 ;
      RECT 87.13 3.735 87.445 3.925 ;
      RECT 87.12 3.735 87.445 3.91 ;
      RECT 87.095 3.735 87.445 3.883 ;
      RECT 87.085 3.735 87.445 3.858 ;
      RECT 87.04 3.59 87.32 3.85 ;
      RECT 87.04 3.685 87.42 3.85 ;
      RECT 87.04 3.63 87.365 3.85 ;
      RECT 87.04 3.622 87.36 3.85 ;
      RECT 87.04 3.612 87.355 3.85 ;
      RECT 87.04 3.6 87.35 3.85 ;
      RECT 85.965 4.295 86.245 4.575 ;
      RECT 85.965 4.295 86.28 4.555 ;
      RECT 78.245 8.95 78.595 9.3 ;
      RECT 85.71 8.905 86.06 9.255 ;
      RECT 78.245 8.98 86.06 9.18 ;
      RECT 86 3.715 86.05 3.975 ;
      RECT 85.79 3.715 85.795 3.975 ;
      RECT 84.985 3.27 85.015 3.53 ;
      RECT 84.755 3.27 84.83 3.53 ;
      RECT 85.975 3.665 86 3.975 ;
      RECT 85.97 3.622 85.975 3.975 ;
      RECT 85.965 3.605 85.97 3.975 ;
      RECT 85.96 3.592 85.965 3.975 ;
      RECT 85.885 3.475 85.96 3.975 ;
      RECT 85.84 3.292 85.885 3.975 ;
      RECT 85.835 3.22 85.84 3.975 ;
      RECT 85.82 3.195 85.835 3.975 ;
      RECT 85.795 3.157 85.82 3.975 ;
      RECT 85.785 3.137 85.795 3.697 ;
      RECT 85.77 3.129 85.785 3.652 ;
      RECT 85.765 3.121 85.77 3.623 ;
      RECT 85.76 3.118 85.765 3.603 ;
      RECT 85.755 3.115 85.76 3.583 ;
      RECT 85.75 3.112 85.755 3.563 ;
      RECT 85.72 3.101 85.75 3.5 ;
      RECT 85.7 3.086 85.72 3.415 ;
      RECT 85.695 3.078 85.7 3.378 ;
      RECT 85.685 3.072 85.695 3.345 ;
      RECT 85.67 3.064 85.685 3.305 ;
      RECT 85.665 3.057 85.67 3.265 ;
      RECT 85.66 3.054 85.665 3.243 ;
      RECT 85.655 3.051 85.66 3.23 ;
      RECT 85.65 3.05 85.655 3.22 ;
      RECT 85.635 3.044 85.65 3.21 ;
      RECT 85.61 3.031 85.635 3.195 ;
      RECT 85.56 3.006 85.61 3.166 ;
      RECT 85.545 2.985 85.56 3.141 ;
      RECT 85.535 2.978 85.545 3.13 ;
      RECT 85.48 2.959 85.535 3.103 ;
      RECT 85.455 2.937 85.48 3.076 ;
      RECT 85.45 2.93 85.455 3.071 ;
      RECT 85.435 2.93 85.45 3.069 ;
      RECT 85.41 2.922 85.435 3.065 ;
      RECT 85.395 2.92 85.41 3.061 ;
      RECT 85.365 2.92 85.395 3.058 ;
      RECT 85.355 2.92 85.365 3.053 ;
      RECT 85.31 2.92 85.355 3.051 ;
      RECT 85.281 2.92 85.31 3.052 ;
      RECT 85.195 2.92 85.281 3.054 ;
      RECT 85.181 2.921 85.195 3.056 ;
      RECT 85.095 2.922 85.181 3.058 ;
      RECT 85.08 2.923 85.095 3.068 ;
      RECT 85.075 2.924 85.08 3.077 ;
      RECT 85.055 2.927 85.075 3.087 ;
      RECT 85.04 2.935 85.055 3.102 ;
      RECT 85.02 2.953 85.04 3.117 ;
      RECT 85.01 2.965 85.02 3.14 ;
      RECT 85 2.974 85.01 3.17 ;
      RECT 84.985 2.986 85 3.215 ;
      RECT 84.93 3.019 84.985 3.53 ;
      RECT 84.925 3.047 84.93 3.53 ;
      RECT 84.905 3.062 84.925 3.53 ;
      RECT 84.87 3.122 84.905 3.53 ;
      RECT 84.868 3.172 84.87 3.53 ;
      RECT 84.865 3.18 84.868 3.53 ;
      RECT 84.855 3.195 84.865 3.53 ;
      RECT 84.85 3.207 84.855 3.53 ;
      RECT 84.84 3.232 84.85 3.53 ;
      RECT 84.83 3.26 84.84 3.53 ;
      RECT 82.735 4.765 82.785 5.025 ;
      RECT 85.645 4.315 85.705 4.575 ;
      RECT 85.63 4.315 85.645 4.585 ;
      RECT 85.611 4.315 85.63 4.618 ;
      RECT 85.525 4.315 85.611 4.743 ;
      RECT 85.445 4.315 85.525 4.925 ;
      RECT 85.44 4.552 85.445 5.01 ;
      RECT 85.415 4.622 85.44 5.038 ;
      RECT 85.41 4.692 85.415 5.065 ;
      RECT 85.39 4.764 85.41 5.087 ;
      RECT 85.385 4.831 85.39 5.11 ;
      RECT 85.375 4.86 85.385 5.125 ;
      RECT 85.365 4.882 85.375 5.142 ;
      RECT 85.36 4.892 85.365 5.153 ;
      RECT 85.355 4.9 85.36 5.161 ;
      RECT 85.345 4.908 85.355 5.173 ;
      RECT 85.34 4.92 85.345 5.183 ;
      RECT 85.335 4.928 85.34 5.188 ;
      RECT 85.315 4.946 85.335 5.198 ;
      RECT 85.31 4.963 85.315 5.205 ;
      RECT 85.305 4.971 85.31 5.206 ;
      RECT 85.3 4.982 85.305 5.208 ;
      RECT 85.26 5.02 85.3 5.218 ;
      RECT 85.255 5.055 85.26 5.229 ;
      RECT 85.25 5.06 85.255 5.232 ;
      RECT 85.225 5.07 85.25 5.239 ;
      RECT 85.215 5.084 85.225 5.248 ;
      RECT 85.195 5.096 85.215 5.251 ;
      RECT 85.145 5.115 85.195 5.255 ;
      RECT 85.1 5.13 85.145 5.26 ;
      RECT 85.035 5.133 85.1 5.266 ;
      RECT 85.02 5.131 85.035 5.273 ;
      RECT 84.99 5.13 85.02 5.273 ;
      RECT 84.951 5.129 84.99 5.269 ;
      RECT 84.865 5.126 84.951 5.265 ;
      RECT 84.848 5.124 84.865 5.262 ;
      RECT 84.762 5.122 84.848 5.259 ;
      RECT 84.676 5.119 84.762 5.253 ;
      RECT 84.59 5.115 84.676 5.248 ;
      RECT 84.512 5.112 84.59 5.244 ;
      RECT 84.426 5.109 84.512 5.242 ;
      RECT 84.34 5.106 84.426 5.239 ;
      RECT 84.282 5.104 84.34 5.236 ;
      RECT 84.196 5.101 84.282 5.234 ;
      RECT 84.11 5.097 84.196 5.232 ;
      RECT 84.024 5.094 84.11 5.229 ;
      RECT 83.938 5.09 84.024 5.227 ;
      RECT 83.852 5.086 83.938 5.224 ;
      RECT 83.766 5.083 83.852 5.222 ;
      RECT 83.68 5.079 83.766 5.219 ;
      RECT 83.594 5.076 83.68 5.217 ;
      RECT 83.508 5.072 83.594 5.214 ;
      RECT 83.422 5.069 83.508 5.212 ;
      RECT 83.336 5.065 83.422 5.209 ;
      RECT 83.25 5.062 83.336 5.207 ;
      RECT 83.24 5.06 83.25 5.203 ;
      RECT 83.235 5.06 83.24 5.201 ;
      RECT 83.195 5.055 83.235 5.195 ;
      RECT 83.181 5.046 83.195 5.188 ;
      RECT 83.095 5.016 83.181 5.173 ;
      RECT 83.075 4.982 83.095 5.158 ;
      RECT 83.005 4.951 83.075 5.145 ;
      RECT 83 4.926 83.005 5.134 ;
      RECT 82.995 4.92 83 5.132 ;
      RECT 82.926 4.765 82.995 5.12 ;
      RECT 82.84 4.765 82.926 5.094 ;
      RECT 82.815 4.765 82.84 5.073 ;
      RECT 82.81 4.765 82.815 5.063 ;
      RECT 82.805 4.765 82.81 5.055 ;
      RECT 82.785 4.765 82.805 5.038 ;
      RECT 85.205 3.335 85.465 3.595 ;
      RECT 85.19 3.335 85.465 3.498 ;
      RECT 85.16 3.335 85.465 3.473 ;
      RECT 85.125 3.175 85.405 3.455 ;
      RECT 85.095 4.665 85.155 4.925 ;
      RECT 84.12 3.355 84.175 3.615 ;
      RECT 85.055 4.622 85.095 4.925 ;
      RECT 85.026 4.543 85.055 4.925 ;
      RECT 84.94 4.415 85.026 4.925 ;
      RECT 84.92 4.295 84.94 4.925 ;
      RECT 84.895 4.246 84.92 4.925 ;
      RECT 84.89 4.211 84.895 4.775 ;
      RECT 84.86 4.171 84.89 4.713 ;
      RECT 84.835 4.108 84.86 4.628 ;
      RECT 84.825 4.07 84.835 4.565 ;
      RECT 84.81 4.045 84.825 4.526 ;
      RECT 84.767 4.003 84.81 4.432 ;
      RECT 84.765 3.976 84.767 4.359 ;
      RECT 84.76 3.971 84.765 4.35 ;
      RECT 84.755 3.964 84.76 4.325 ;
      RECT 84.75 3.958 84.755 4.31 ;
      RECT 84.745 3.952 84.75 4.298 ;
      RECT 84.735 3.943 84.745 4.28 ;
      RECT 84.73 3.934 84.735 4.258 ;
      RECT 84.705 3.915 84.73 4.208 ;
      RECT 84.7 3.896 84.705 4.158 ;
      RECT 84.685 3.882 84.7 4.118 ;
      RECT 84.68 3.868 84.685 4.085 ;
      RECT 84.675 3.861 84.68 4.078 ;
      RECT 84.66 3.848 84.675 4.07 ;
      RECT 84.615 3.81 84.66 4.043 ;
      RECT 84.585 3.763 84.615 4.008 ;
      RECT 84.565 3.732 84.585 3.985 ;
      RECT 84.485 3.665 84.565 3.938 ;
      RECT 84.455 3.595 84.485 3.885 ;
      RECT 84.45 3.572 84.455 3.868 ;
      RECT 84.42 3.55 84.45 3.853 ;
      RECT 84.39 3.509 84.42 3.825 ;
      RECT 84.385 3.484 84.39 3.81 ;
      RECT 84.38 3.478 84.385 3.803 ;
      RECT 84.37 3.355 84.38 3.795 ;
      RECT 84.36 3.355 84.37 3.788 ;
      RECT 84.355 3.355 84.36 3.78 ;
      RECT 84.335 3.355 84.355 3.768 ;
      RECT 84.285 3.355 84.335 3.738 ;
      RECT 84.23 3.355 84.285 3.688 ;
      RECT 84.2 3.355 84.23 3.648 ;
      RECT 84.175 3.355 84.2 3.625 ;
      RECT 84.045 4.08 84.325 4.36 ;
      RECT 84.01 3.995 84.27 4.255 ;
      RECT 84.01 4.077 84.28 4.255 ;
      RECT 82.21 3.45 82.215 3.935 ;
      RECT 82.1 3.635 82.105 3.935 ;
      RECT 82.01 3.675 82.075 3.935 ;
      RECT 83.685 3.175 83.775 3.805 ;
      RECT 83.65 3.225 83.655 3.805 ;
      RECT 83.595 3.25 83.605 3.805 ;
      RECT 83.55 3.25 83.56 3.805 ;
      RECT 83.92 3.175 83.965 3.455 ;
      RECT 82.77 2.905 82.97 3.045 ;
      RECT 83.886 3.175 83.92 3.467 ;
      RECT 83.8 3.175 83.886 3.507 ;
      RECT 83.785 3.175 83.8 3.548 ;
      RECT 83.78 3.175 83.785 3.568 ;
      RECT 83.775 3.175 83.78 3.588 ;
      RECT 83.655 3.217 83.685 3.805 ;
      RECT 83.605 3.237 83.65 3.805 ;
      RECT 83.59 3.252 83.595 3.805 ;
      RECT 83.56 3.252 83.59 3.805 ;
      RECT 83.515 3.237 83.55 3.805 ;
      RECT 83.51 3.225 83.515 3.585 ;
      RECT 83.505 3.222 83.51 3.565 ;
      RECT 83.49 3.212 83.505 3.518 ;
      RECT 83.485 3.205 83.49 3.481 ;
      RECT 83.48 3.202 83.485 3.464 ;
      RECT 83.465 3.192 83.48 3.42 ;
      RECT 83.46 3.183 83.465 3.38 ;
      RECT 83.455 3.179 83.46 3.365 ;
      RECT 83.445 3.173 83.455 3.348 ;
      RECT 83.405 3.154 83.445 3.323 ;
      RECT 83.4 3.136 83.405 3.303 ;
      RECT 83.39 3.13 83.4 3.298 ;
      RECT 83.36 3.114 83.39 3.285 ;
      RECT 83.345 3.096 83.36 3.268 ;
      RECT 83.33 3.084 83.345 3.255 ;
      RECT 83.325 3.076 83.33 3.248 ;
      RECT 83.295 3.062 83.325 3.235 ;
      RECT 83.29 3.047 83.295 3.223 ;
      RECT 83.28 3.041 83.29 3.215 ;
      RECT 83.26 3.029 83.28 3.203 ;
      RECT 83.25 3.017 83.26 3.19 ;
      RECT 83.22 3.001 83.25 3.175 ;
      RECT 83.2 2.981 83.22 3.158 ;
      RECT 83.195 2.971 83.2 3.148 ;
      RECT 83.17 2.959 83.195 3.135 ;
      RECT 83.165 2.947 83.17 3.123 ;
      RECT 83.16 2.942 83.165 3.119 ;
      RECT 83.145 2.935 83.16 3.111 ;
      RECT 83.135 2.922 83.145 3.101 ;
      RECT 83.13 2.92 83.135 3.095 ;
      RECT 83.105 2.913 83.13 3.084 ;
      RECT 83.1 2.906 83.105 3.073 ;
      RECT 83.075 2.905 83.1 3.06 ;
      RECT 83.056 2.905 83.075 3.05 ;
      RECT 82.97 2.905 83.056 3.047 ;
      RECT 82.74 2.905 82.77 3.05 ;
      RECT 82.7 2.912 82.74 3.063 ;
      RECT 82.675 2.922 82.7 3.076 ;
      RECT 82.66 2.931 82.675 3.086 ;
      RECT 82.63 2.936 82.66 3.105 ;
      RECT 82.625 2.942 82.63 3.123 ;
      RECT 82.605 2.952 82.625 3.138 ;
      RECT 82.595 2.965 82.605 3.158 ;
      RECT 82.58 2.977 82.595 3.175 ;
      RECT 82.575 2.987 82.58 3.185 ;
      RECT 82.57 2.992 82.575 3.19 ;
      RECT 82.56 3 82.57 3.203 ;
      RECT 82.51 3.032 82.56 3.24 ;
      RECT 82.495 3.067 82.51 3.281 ;
      RECT 82.49 3.077 82.495 3.296 ;
      RECT 82.485 3.082 82.49 3.303 ;
      RECT 82.46 3.098 82.485 3.323 ;
      RECT 82.445 3.119 82.46 3.348 ;
      RECT 82.42 3.14 82.445 3.373 ;
      RECT 82.41 3.159 82.42 3.396 ;
      RECT 82.385 3.177 82.41 3.419 ;
      RECT 82.37 3.197 82.385 3.443 ;
      RECT 82.365 3.207 82.37 3.455 ;
      RECT 82.35 3.219 82.365 3.475 ;
      RECT 82.34 3.234 82.35 3.515 ;
      RECT 82.335 3.242 82.34 3.543 ;
      RECT 82.325 3.252 82.335 3.563 ;
      RECT 82.32 3.265 82.325 3.588 ;
      RECT 82.315 3.278 82.32 3.608 ;
      RECT 82.31 3.284 82.315 3.63 ;
      RECT 82.3 3.293 82.31 3.65 ;
      RECT 82.295 3.313 82.3 3.673 ;
      RECT 82.29 3.319 82.295 3.693 ;
      RECT 82.285 3.326 82.29 3.715 ;
      RECT 82.28 3.337 82.285 3.728 ;
      RECT 82.27 3.347 82.28 3.753 ;
      RECT 82.25 3.372 82.27 3.935 ;
      RECT 82.22 3.412 82.25 3.935 ;
      RECT 82.215 3.442 82.22 3.935 ;
      RECT 82.19 3.47 82.21 3.935 ;
      RECT 82.16 3.515 82.19 3.935 ;
      RECT 82.155 3.542 82.16 3.935 ;
      RECT 82.135 3.56 82.155 3.935 ;
      RECT 82.125 3.585 82.135 3.935 ;
      RECT 82.12 3.597 82.125 3.935 ;
      RECT 82.105 3.62 82.12 3.935 ;
      RECT 82.085 3.647 82.1 3.935 ;
      RECT 82.075 3.67 82.085 3.935 ;
      RECT 83.865 4.555 83.945 4.815 ;
      RECT 83.1 3.775 83.17 4.035 ;
      RECT 83.831 4.522 83.865 4.815 ;
      RECT 83.745 4.425 83.831 4.815 ;
      RECT 83.725 4.337 83.745 4.815 ;
      RECT 83.715 4.307 83.725 4.815 ;
      RECT 83.705 4.287 83.715 4.815 ;
      RECT 83.685 4.274 83.705 4.815 ;
      RECT 83.67 4.264 83.685 4.643 ;
      RECT 83.665 4.257 83.67 4.598 ;
      RECT 83.655 4.251 83.665 4.588 ;
      RECT 83.645 4.243 83.655 4.57 ;
      RECT 83.64 4.237 83.645 4.558 ;
      RECT 83.63 4.232 83.64 4.545 ;
      RECT 83.61 4.222 83.63 4.518 ;
      RECT 83.57 4.201 83.61 4.47 ;
      RECT 83.555 4.182 83.57 4.428 ;
      RECT 83.53 4.168 83.555 4.398 ;
      RECT 83.52 4.156 83.53 4.365 ;
      RECT 83.515 4.151 83.52 4.355 ;
      RECT 83.485 4.137 83.515 4.335 ;
      RECT 83.475 4.121 83.485 4.308 ;
      RECT 83.47 4.116 83.475 4.298 ;
      RECT 83.445 4.107 83.47 4.278 ;
      RECT 83.435 4.095 83.445 4.258 ;
      RECT 83.365 4.063 83.435 4.233 ;
      RECT 83.36 4.032 83.365 4.21 ;
      RECT 83.311 3.775 83.36 4.193 ;
      RECT 83.225 3.775 83.311 4.152 ;
      RECT 83.17 3.775 83.225 4.08 ;
      RECT 83.26 4.56 83.42 4.82 ;
      RECT 82.785 3.175 82.835 3.86 ;
      RECT 82.575 3.6 82.61 3.86 ;
      RECT 82.89 3.175 82.895 3.635 ;
      RECT 82.98 3.175 83.005 3.455 ;
      RECT 83.255 4.557 83.26 4.82 ;
      RECT 83.22 4.545 83.255 4.82 ;
      RECT 83.16 4.518 83.22 4.82 ;
      RECT 83.155 4.501 83.16 4.674 ;
      RECT 83.15 4.498 83.155 4.661 ;
      RECT 83.13 4.491 83.15 4.648 ;
      RECT 83.095 4.474 83.13 4.63 ;
      RECT 83.055 4.453 83.095 4.61 ;
      RECT 83.05 4.441 83.055 4.598 ;
      RECT 83.01 4.427 83.05 4.584 ;
      RECT 82.99 4.41 83.01 4.566 ;
      RECT 82.98 4.402 82.99 4.558 ;
      RECT 82.965 3.175 82.98 3.473 ;
      RECT 82.95 4.392 82.98 4.545 ;
      RECT 82.935 3.175 82.965 3.518 ;
      RECT 82.94 4.382 82.95 4.532 ;
      RECT 82.91 4.367 82.94 4.519 ;
      RECT 82.895 3.175 82.935 3.585 ;
      RECT 82.895 4.335 82.91 4.505 ;
      RECT 82.89 4.307 82.895 4.499 ;
      RECT 82.885 3.175 82.89 3.64 ;
      RECT 82.875 4.277 82.89 4.493 ;
      RECT 82.88 3.175 82.885 3.653 ;
      RECT 82.87 3.175 82.88 3.673 ;
      RECT 82.835 4.19 82.875 4.478 ;
      RECT 82.835 3.175 82.87 3.713 ;
      RECT 82.83 4.122 82.835 4.466 ;
      RECT 82.815 4.077 82.83 4.461 ;
      RECT 82.81 4.015 82.815 4.456 ;
      RECT 82.785 3.922 82.81 4.449 ;
      RECT 82.78 3.175 82.785 4.441 ;
      RECT 82.765 3.175 82.78 4.428 ;
      RECT 82.745 3.175 82.765 4.385 ;
      RECT 82.735 3.175 82.745 4.335 ;
      RECT 82.73 3.175 82.735 4.308 ;
      RECT 82.725 3.175 82.73 4.286 ;
      RECT 82.72 3.401 82.725 4.269 ;
      RECT 82.715 3.423 82.72 4.247 ;
      RECT 82.71 3.465 82.715 4.23 ;
      RECT 82.68 3.515 82.71 4.174 ;
      RECT 82.675 3.542 82.68 4.116 ;
      RECT 82.66 3.56 82.675 4.08 ;
      RECT 82.655 3.578 82.66 4.044 ;
      RECT 82.649 3.585 82.655 4.025 ;
      RECT 82.645 3.592 82.649 4.008 ;
      RECT 82.64 3.597 82.645 3.977 ;
      RECT 82.63 3.6 82.64 3.952 ;
      RECT 82.62 3.6 82.63 3.918 ;
      RECT 82.615 3.6 82.62 3.895 ;
      RECT 82.61 3.6 82.615 3.875 ;
      RECT 81.23 4.765 81.49 5.025 ;
      RECT 81.25 4.692 81.43 5.025 ;
      RECT 81.25 4.435 81.425 5.025 ;
      RECT 81.25 4.227 81.415 5.025 ;
      RECT 81.255 4.145 81.415 5.025 ;
      RECT 81.255 3.91 81.405 5.025 ;
      RECT 81.255 3.757 81.4 5.025 ;
      RECT 81.26 3.742 81.4 5.025 ;
      RECT 81.31 3.457 81.4 5.025 ;
      RECT 81.265 3.692 81.4 5.025 ;
      RECT 81.295 3.51 81.4 5.025 ;
      RECT 81.28 3.622 81.4 5.025 ;
      RECT 81.285 3.58 81.4 5.025 ;
      RECT 81.28 3.622 81.415 3.685 ;
      RECT 81.315 3.21 81.42 3.63 ;
      RECT 81.315 3.21 81.435 3.613 ;
      RECT 81.315 3.21 81.47 3.575 ;
      RECT 81.31 3.457 81.52 3.508 ;
      RECT 81.315 3.21 81.575 3.47 ;
      RECT 80.575 3.915 80.835 4.175 ;
      RECT 80.575 3.915 80.845 4.133 ;
      RECT 80.575 3.915 80.931 4.104 ;
      RECT 80.575 3.915 81 4.056 ;
      RECT 80.575 3.915 81.035 4.025 ;
      RECT 80.805 3.735 81.085 4.015 ;
      RECT 80.64 3.9 81.085 4.015 ;
      RECT 80.73 3.777 80.835 4.175 ;
      RECT 80.66 3.84 81.085 4.015 ;
      RECT 75.11 8.51 75.43 8.835 ;
      RECT 75.14 7.985 75.31 8.835 ;
      RECT 75.14 7.985 75.315 8.335 ;
      RECT 75.14 7.985 76.115 8.16 ;
      RECT 75.94 3.26 76.115 8.16 ;
      RECT 75.885 3.26 76.235 3.61 ;
      RECT 75.91 8.945 76.235 9.27 ;
      RECT 74.795 9.035 76.235 9.205 ;
      RECT 74.795 3.69 74.955 9.205 ;
      RECT 75.11 3.66 75.43 3.98 ;
      RECT 74.795 3.69 75.43 3.86 ;
      RECT 73.46 4 73.845 4.35 ;
      RECT 73.45 4.065 73.845 4.265 ;
      RECT 73.595 3.995 73.765 4.35 ;
      RECT 71.905 3.735 72.185 4.015 ;
      RECT 71.9 3.735 72.185 3.968 ;
      RECT 71.88 3.735 72.185 3.945 ;
      RECT 71.87 3.735 72.185 3.925 ;
      RECT 71.86 3.735 72.185 3.91 ;
      RECT 71.835 3.735 72.185 3.883 ;
      RECT 71.825 3.735 72.185 3.858 ;
      RECT 71.78 3.59 72.06 3.85 ;
      RECT 71.78 3.685 72.16 3.85 ;
      RECT 71.78 3.63 72.105 3.85 ;
      RECT 71.78 3.622 72.1 3.85 ;
      RECT 71.78 3.612 72.095 3.85 ;
      RECT 71.78 3.6 72.09 3.85 ;
      RECT 70.705 4.295 70.985 4.575 ;
      RECT 70.705 4.295 71.02 4.555 ;
      RECT 62.985 8.95 63.335 9.3 ;
      RECT 70.45 8.905 70.8 9.255 ;
      RECT 62.985 8.98 70.8 9.18 ;
      RECT 70.74 3.715 70.79 3.975 ;
      RECT 70.53 3.715 70.535 3.975 ;
      RECT 69.725 3.27 69.755 3.53 ;
      RECT 69.495 3.27 69.57 3.53 ;
      RECT 70.715 3.665 70.74 3.975 ;
      RECT 70.71 3.622 70.715 3.975 ;
      RECT 70.705 3.605 70.71 3.975 ;
      RECT 70.7 3.592 70.705 3.975 ;
      RECT 70.625 3.475 70.7 3.975 ;
      RECT 70.58 3.292 70.625 3.975 ;
      RECT 70.575 3.22 70.58 3.975 ;
      RECT 70.56 3.195 70.575 3.975 ;
      RECT 70.535 3.157 70.56 3.975 ;
      RECT 70.525 3.137 70.535 3.697 ;
      RECT 70.51 3.129 70.525 3.652 ;
      RECT 70.505 3.121 70.51 3.623 ;
      RECT 70.5 3.118 70.505 3.603 ;
      RECT 70.495 3.115 70.5 3.583 ;
      RECT 70.49 3.112 70.495 3.563 ;
      RECT 70.46 3.101 70.49 3.5 ;
      RECT 70.44 3.086 70.46 3.415 ;
      RECT 70.435 3.078 70.44 3.378 ;
      RECT 70.425 3.072 70.435 3.345 ;
      RECT 70.41 3.064 70.425 3.305 ;
      RECT 70.405 3.057 70.41 3.265 ;
      RECT 70.4 3.054 70.405 3.243 ;
      RECT 70.395 3.051 70.4 3.23 ;
      RECT 70.39 3.05 70.395 3.22 ;
      RECT 70.375 3.044 70.39 3.21 ;
      RECT 70.35 3.031 70.375 3.195 ;
      RECT 70.3 3.006 70.35 3.166 ;
      RECT 70.285 2.985 70.3 3.141 ;
      RECT 70.275 2.978 70.285 3.13 ;
      RECT 70.22 2.959 70.275 3.103 ;
      RECT 70.195 2.937 70.22 3.076 ;
      RECT 70.19 2.93 70.195 3.071 ;
      RECT 70.175 2.93 70.19 3.069 ;
      RECT 70.15 2.922 70.175 3.065 ;
      RECT 70.135 2.92 70.15 3.061 ;
      RECT 70.105 2.92 70.135 3.058 ;
      RECT 70.095 2.92 70.105 3.053 ;
      RECT 70.05 2.92 70.095 3.051 ;
      RECT 70.021 2.92 70.05 3.052 ;
      RECT 69.935 2.92 70.021 3.054 ;
      RECT 69.921 2.921 69.935 3.056 ;
      RECT 69.835 2.922 69.921 3.058 ;
      RECT 69.82 2.923 69.835 3.068 ;
      RECT 69.815 2.924 69.82 3.077 ;
      RECT 69.795 2.927 69.815 3.087 ;
      RECT 69.78 2.935 69.795 3.102 ;
      RECT 69.76 2.953 69.78 3.117 ;
      RECT 69.75 2.965 69.76 3.14 ;
      RECT 69.74 2.974 69.75 3.17 ;
      RECT 69.725 2.986 69.74 3.215 ;
      RECT 69.67 3.019 69.725 3.53 ;
      RECT 69.665 3.047 69.67 3.53 ;
      RECT 69.645 3.062 69.665 3.53 ;
      RECT 69.61 3.122 69.645 3.53 ;
      RECT 69.608 3.172 69.61 3.53 ;
      RECT 69.605 3.18 69.608 3.53 ;
      RECT 69.595 3.195 69.605 3.53 ;
      RECT 69.59 3.207 69.595 3.53 ;
      RECT 69.58 3.232 69.59 3.53 ;
      RECT 69.57 3.26 69.58 3.53 ;
      RECT 67.475 4.765 67.525 5.025 ;
      RECT 70.385 4.315 70.445 4.575 ;
      RECT 70.37 4.315 70.385 4.585 ;
      RECT 70.351 4.315 70.37 4.618 ;
      RECT 70.265 4.315 70.351 4.743 ;
      RECT 70.185 4.315 70.265 4.925 ;
      RECT 70.18 4.552 70.185 5.01 ;
      RECT 70.155 4.622 70.18 5.038 ;
      RECT 70.15 4.692 70.155 5.065 ;
      RECT 70.13 4.764 70.15 5.087 ;
      RECT 70.125 4.831 70.13 5.11 ;
      RECT 70.115 4.86 70.125 5.125 ;
      RECT 70.105 4.882 70.115 5.142 ;
      RECT 70.1 4.892 70.105 5.153 ;
      RECT 70.095 4.9 70.1 5.161 ;
      RECT 70.085 4.908 70.095 5.173 ;
      RECT 70.08 4.92 70.085 5.183 ;
      RECT 70.075 4.928 70.08 5.188 ;
      RECT 70.055 4.946 70.075 5.198 ;
      RECT 70.05 4.963 70.055 5.205 ;
      RECT 70.045 4.971 70.05 5.206 ;
      RECT 70.04 4.982 70.045 5.208 ;
      RECT 70 5.02 70.04 5.218 ;
      RECT 69.995 5.055 70 5.229 ;
      RECT 69.99 5.06 69.995 5.232 ;
      RECT 69.965 5.07 69.99 5.239 ;
      RECT 69.955 5.084 69.965 5.248 ;
      RECT 69.935 5.096 69.955 5.251 ;
      RECT 69.885 5.115 69.935 5.255 ;
      RECT 69.84 5.13 69.885 5.26 ;
      RECT 69.775 5.133 69.84 5.266 ;
      RECT 69.76 5.131 69.775 5.273 ;
      RECT 69.73 5.13 69.76 5.273 ;
      RECT 69.691 5.129 69.73 5.269 ;
      RECT 69.605 5.126 69.691 5.265 ;
      RECT 69.588 5.124 69.605 5.262 ;
      RECT 69.502 5.122 69.588 5.259 ;
      RECT 69.416 5.119 69.502 5.253 ;
      RECT 69.33 5.115 69.416 5.248 ;
      RECT 69.252 5.112 69.33 5.244 ;
      RECT 69.166 5.109 69.252 5.242 ;
      RECT 69.08 5.106 69.166 5.239 ;
      RECT 69.022 5.104 69.08 5.236 ;
      RECT 68.936 5.101 69.022 5.234 ;
      RECT 68.85 5.097 68.936 5.232 ;
      RECT 68.764 5.094 68.85 5.229 ;
      RECT 68.678 5.09 68.764 5.227 ;
      RECT 68.592 5.086 68.678 5.224 ;
      RECT 68.506 5.083 68.592 5.222 ;
      RECT 68.42 5.079 68.506 5.219 ;
      RECT 68.334 5.076 68.42 5.217 ;
      RECT 68.248 5.072 68.334 5.214 ;
      RECT 68.162 5.069 68.248 5.212 ;
      RECT 68.076 5.065 68.162 5.209 ;
      RECT 67.99 5.062 68.076 5.207 ;
      RECT 67.98 5.06 67.99 5.203 ;
      RECT 67.975 5.06 67.98 5.201 ;
      RECT 67.935 5.055 67.975 5.195 ;
      RECT 67.921 5.046 67.935 5.188 ;
      RECT 67.835 5.016 67.921 5.173 ;
      RECT 67.815 4.982 67.835 5.158 ;
      RECT 67.745 4.951 67.815 5.145 ;
      RECT 67.74 4.926 67.745 5.134 ;
      RECT 67.735 4.92 67.74 5.132 ;
      RECT 67.666 4.765 67.735 5.12 ;
      RECT 67.58 4.765 67.666 5.094 ;
      RECT 67.555 4.765 67.58 5.073 ;
      RECT 67.55 4.765 67.555 5.063 ;
      RECT 67.545 4.765 67.55 5.055 ;
      RECT 67.525 4.765 67.545 5.038 ;
      RECT 69.945 3.335 70.205 3.595 ;
      RECT 69.93 3.335 70.205 3.498 ;
      RECT 69.9 3.335 70.205 3.473 ;
      RECT 69.865 3.175 70.145 3.455 ;
      RECT 69.835 4.665 69.895 4.925 ;
      RECT 68.86 3.355 68.915 3.615 ;
      RECT 69.795 4.622 69.835 4.925 ;
      RECT 69.766 4.543 69.795 4.925 ;
      RECT 69.68 4.415 69.766 4.925 ;
      RECT 69.66 4.295 69.68 4.925 ;
      RECT 69.635 4.246 69.66 4.925 ;
      RECT 69.63 4.211 69.635 4.775 ;
      RECT 69.6 4.171 69.63 4.713 ;
      RECT 69.575 4.108 69.6 4.628 ;
      RECT 69.565 4.07 69.575 4.565 ;
      RECT 69.55 4.045 69.565 4.526 ;
      RECT 69.507 4.003 69.55 4.432 ;
      RECT 69.505 3.976 69.507 4.359 ;
      RECT 69.5 3.971 69.505 4.35 ;
      RECT 69.495 3.964 69.5 4.325 ;
      RECT 69.49 3.958 69.495 4.31 ;
      RECT 69.485 3.952 69.49 4.298 ;
      RECT 69.475 3.943 69.485 4.28 ;
      RECT 69.47 3.934 69.475 4.258 ;
      RECT 69.445 3.915 69.47 4.208 ;
      RECT 69.44 3.896 69.445 4.158 ;
      RECT 69.425 3.882 69.44 4.118 ;
      RECT 69.42 3.868 69.425 4.085 ;
      RECT 69.415 3.861 69.42 4.078 ;
      RECT 69.4 3.848 69.415 4.07 ;
      RECT 69.355 3.81 69.4 4.043 ;
      RECT 69.325 3.763 69.355 4.008 ;
      RECT 69.305 3.732 69.325 3.985 ;
      RECT 69.225 3.665 69.305 3.938 ;
      RECT 69.195 3.595 69.225 3.885 ;
      RECT 69.19 3.572 69.195 3.868 ;
      RECT 69.16 3.55 69.19 3.853 ;
      RECT 69.13 3.509 69.16 3.825 ;
      RECT 69.125 3.484 69.13 3.81 ;
      RECT 69.12 3.478 69.125 3.803 ;
      RECT 69.11 3.355 69.12 3.795 ;
      RECT 69.1 3.355 69.11 3.788 ;
      RECT 69.095 3.355 69.1 3.78 ;
      RECT 69.075 3.355 69.095 3.768 ;
      RECT 69.025 3.355 69.075 3.738 ;
      RECT 68.97 3.355 69.025 3.688 ;
      RECT 68.94 3.355 68.97 3.648 ;
      RECT 68.915 3.355 68.94 3.625 ;
      RECT 68.785 4.08 69.065 4.36 ;
      RECT 68.75 3.995 69.01 4.255 ;
      RECT 68.75 4.077 69.02 4.255 ;
      RECT 66.95 3.45 66.955 3.935 ;
      RECT 66.84 3.635 66.845 3.935 ;
      RECT 66.75 3.675 66.815 3.935 ;
      RECT 68.425 3.175 68.515 3.805 ;
      RECT 68.39 3.225 68.395 3.805 ;
      RECT 68.335 3.25 68.345 3.805 ;
      RECT 68.29 3.25 68.3 3.805 ;
      RECT 68.66 3.175 68.705 3.455 ;
      RECT 67.51 2.905 67.71 3.045 ;
      RECT 68.626 3.175 68.66 3.467 ;
      RECT 68.54 3.175 68.626 3.507 ;
      RECT 68.525 3.175 68.54 3.548 ;
      RECT 68.52 3.175 68.525 3.568 ;
      RECT 68.515 3.175 68.52 3.588 ;
      RECT 68.395 3.217 68.425 3.805 ;
      RECT 68.345 3.237 68.39 3.805 ;
      RECT 68.33 3.252 68.335 3.805 ;
      RECT 68.3 3.252 68.33 3.805 ;
      RECT 68.255 3.237 68.29 3.805 ;
      RECT 68.25 3.225 68.255 3.585 ;
      RECT 68.245 3.222 68.25 3.565 ;
      RECT 68.23 3.212 68.245 3.518 ;
      RECT 68.225 3.205 68.23 3.481 ;
      RECT 68.22 3.202 68.225 3.464 ;
      RECT 68.205 3.192 68.22 3.42 ;
      RECT 68.2 3.183 68.205 3.38 ;
      RECT 68.195 3.179 68.2 3.365 ;
      RECT 68.185 3.173 68.195 3.348 ;
      RECT 68.145 3.154 68.185 3.323 ;
      RECT 68.14 3.136 68.145 3.303 ;
      RECT 68.13 3.13 68.14 3.298 ;
      RECT 68.1 3.114 68.13 3.285 ;
      RECT 68.085 3.096 68.1 3.268 ;
      RECT 68.07 3.084 68.085 3.255 ;
      RECT 68.065 3.076 68.07 3.248 ;
      RECT 68.035 3.062 68.065 3.235 ;
      RECT 68.03 3.047 68.035 3.223 ;
      RECT 68.02 3.041 68.03 3.215 ;
      RECT 68 3.029 68.02 3.203 ;
      RECT 67.99 3.017 68 3.19 ;
      RECT 67.96 3.001 67.99 3.175 ;
      RECT 67.94 2.981 67.96 3.158 ;
      RECT 67.935 2.971 67.94 3.148 ;
      RECT 67.91 2.959 67.935 3.135 ;
      RECT 67.905 2.947 67.91 3.123 ;
      RECT 67.9 2.942 67.905 3.119 ;
      RECT 67.885 2.935 67.9 3.111 ;
      RECT 67.875 2.922 67.885 3.101 ;
      RECT 67.87 2.92 67.875 3.095 ;
      RECT 67.845 2.913 67.87 3.084 ;
      RECT 67.84 2.906 67.845 3.073 ;
      RECT 67.815 2.905 67.84 3.06 ;
      RECT 67.796 2.905 67.815 3.05 ;
      RECT 67.71 2.905 67.796 3.047 ;
      RECT 67.48 2.905 67.51 3.05 ;
      RECT 67.44 2.912 67.48 3.063 ;
      RECT 67.415 2.922 67.44 3.076 ;
      RECT 67.4 2.931 67.415 3.086 ;
      RECT 67.37 2.936 67.4 3.105 ;
      RECT 67.365 2.942 67.37 3.123 ;
      RECT 67.345 2.952 67.365 3.138 ;
      RECT 67.335 2.965 67.345 3.158 ;
      RECT 67.32 2.977 67.335 3.175 ;
      RECT 67.315 2.987 67.32 3.185 ;
      RECT 67.31 2.992 67.315 3.19 ;
      RECT 67.3 3 67.31 3.203 ;
      RECT 67.25 3.032 67.3 3.24 ;
      RECT 67.235 3.067 67.25 3.281 ;
      RECT 67.23 3.077 67.235 3.296 ;
      RECT 67.225 3.082 67.23 3.303 ;
      RECT 67.2 3.098 67.225 3.323 ;
      RECT 67.185 3.119 67.2 3.348 ;
      RECT 67.16 3.14 67.185 3.373 ;
      RECT 67.15 3.159 67.16 3.396 ;
      RECT 67.125 3.177 67.15 3.419 ;
      RECT 67.11 3.197 67.125 3.443 ;
      RECT 67.105 3.207 67.11 3.455 ;
      RECT 67.09 3.219 67.105 3.475 ;
      RECT 67.08 3.234 67.09 3.515 ;
      RECT 67.075 3.242 67.08 3.543 ;
      RECT 67.065 3.252 67.075 3.563 ;
      RECT 67.06 3.265 67.065 3.588 ;
      RECT 67.055 3.278 67.06 3.608 ;
      RECT 67.05 3.284 67.055 3.63 ;
      RECT 67.04 3.293 67.05 3.65 ;
      RECT 67.035 3.313 67.04 3.673 ;
      RECT 67.03 3.319 67.035 3.693 ;
      RECT 67.025 3.326 67.03 3.715 ;
      RECT 67.02 3.337 67.025 3.728 ;
      RECT 67.01 3.347 67.02 3.753 ;
      RECT 66.99 3.372 67.01 3.935 ;
      RECT 66.96 3.412 66.99 3.935 ;
      RECT 66.955 3.442 66.96 3.935 ;
      RECT 66.93 3.47 66.95 3.935 ;
      RECT 66.9 3.515 66.93 3.935 ;
      RECT 66.895 3.542 66.9 3.935 ;
      RECT 66.875 3.56 66.895 3.935 ;
      RECT 66.865 3.585 66.875 3.935 ;
      RECT 66.86 3.597 66.865 3.935 ;
      RECT 66.845 3.62 66.86 3.935 ;
      RECT 66.825 3.647 66.84 3.935 ;
      RECT 66.815 3.67 66.825 3.935 ;
      RECT 68.605 4.555 68.685 4.815 ;
      RECT 67.84 3.775 67.91 4.035 ;
      RECT 68.571 4.522 68.605 4.815 ;
      RECT 68.485 4.425 68.571 4.815 ;
      RECT 68.465 4.337 68.485 4.815 ;
      RECT 68.455 4.307 68.465 4.815 ;
      RECT 68.445 4.287 68.455 4.815 ;
      RECT 68.425 4.274 68.445 4.815 ;
      RECT 68.41 4.264 68.425 4.643 ;
      RECT 68.405 4.257 68.41 4.598 ;
      RECT 68.395 4.251 68.405 4.588 ;
      RECT 68.385 4.243 68.395 4.57 ;
      RECT 68.38 4.237 68.385 4.558 ;
      RECT 68.37 4.232 68.38 4.545 ;
      RECT 68.35 4.222 68.37 4.518 ;
      RECT 68.31 4.201 68.35 4.47 ;
      RECT 68.295 4.182 68.31 4.428 ;
      RECT 68.27 4.168 68.295 4.398 ;
      RECT 68.26 4.156 68.27 4.365 ;
      RECT 68.255 4.151 68.26 4.355 ;
      RECT 68.225 4.137 68.255 4.335 ;
      RECT 68.215 4.121 68.225 4.308 ;
      RECT 68.21 4.116 68.215 4.298 ;
      RECT 68.185 4.107 68.21 4.278 ;
      RECT 68.175 4.095 68.185 4.258 ;
      RECT 68.105 4.063 68.175 4.233 ;
      RECT 68.1 4.032 68.105 4.21 ;
      RECT 68.051 3.775 68.1 4.193 ;
      RECT 67.965 3.775 68.051 4.152 ;
      RECT 67.91 3.775 67.965 4.08 ;
      RECT 68 4.56 68.16 4.82 ;
      RECT 67.525 3.175 67.575 3.86 ;
      RECT 67.315 3.6 67.35 3.86 ;
      RECT 67.63 3.175 67.635 3.635 ;
      RECT 67.72 3.175 67.745 3.455 ;
      RECT 67.995 4.557 68 4.82 ;
      RECT 67.96 4.545 67.995 4.82 ;
      RECT 67.9 4.518 67.96 4.82 ;
      RECT 67.895 4.501 67.9 4.674 ;
      RECT 67.89 4.498 67.895 4.661 ;
      RECT 67.87 4.491 67.89 4.648 ;
      RECT 67.835 4.474 67.87 4.63 ;
      RECT 67.795 4.453 67.835 4.61 ;
      RECT 67.79 4.441 67.795 4.598 ;
      RECT 67.75 4.427 67.79 4.584 ;
      RECT 67.73 4.41 67.75 4.566 ;
      RECT 67.72 4.402 67.73 4.558 ;
      RECT 67.705 3.175 67.72 3.473 ;
      RECT 67.69 4.392 67.72 4.545 ;
      RECT 67.675 3.175 67.705 3.518 ;
      RECT 67.68 4.382 67.69 4.532 ;
      RECT 67.65 4.367 67.68 4.519 ;
      RECT 67.635 3.175 67.675 3.585 ;
      RECT 67.635 4.335 67.65 4.505 ;
      RECT 67.63 4.307 67.635 4.499 ;
      RECT 67.625 3.175 67.63 3.64 ;
      RECT 67.615 4.277 67.63 4.493 ;
      RECT 67.62 3.175 67.625 3.653 ;
      RECT 67.61 3.175 67.62 3.673 ;
      RECT 67.575 4.19 67.615 4.478 ;
      RECT 67.575 3.175 67.61 3.713 ;
      RECT 67.57 4.122 67.575 4.466 ;
      RECT 67.555 4.077 67.57 4.461 ;
      RECT 67.55 4.015 67.555 4.456 ;
      RECT 67.525 3.922 67.55 4.449 ;
      RECT 67.52 3.175 67.525 4.441 ;
      RECT 67.505 3.175 67.52 4.428 ;
      RECT 67.485 3.175 67.505 4.385 ;
      RECT 67.475 3.175 67.485 4.335 ;
      RECT 67.47 3.175 67.475 4.308 ;
      RECT 67.465 3.175 67.47 4.286 ;
      RECT 67.46 3.401 67.465 4.269 ;
      RECT 67.455 3.423 67.46 4.247 ;
      RECT 67.45 3.465 67.455 4.23 ;
      RECT 67.42 3.515 67.45 4.174 ;
      RECT 67.415 3.542 67.42 4.116 ;
      RECT 67.4 3.56 67.415 4.08 ;
      RECT 67.395 3.578 67.4 4.044 ;
      RECT 67.389 3.585 67.395 4.025 ;
      RECT 67.385 3.592 67.389 4.008 ;
      RECT 67.38 3.597 67.385 3.977 ;
      RECT 67.37 3.6 67.38 3.952 ;
      RECT 67.36 3.6 67.37 3.918 ;
      RECT 67.355 3.6 67.36 3.895 ;
      RECT 67.35 3.6 67.355 3.875 ;
      RECT 65.97 4.765 66.23 5.025 ;
      RECT 65.99 4.692 66.17 5.025 ;
      RECT 65.99 4.435 66.165 5.025 ;
      RECT 65.99 4.227 66.155 5.025 ;
      RECT 65.995 4.145 66.155 5.025 ;
      RECT 65.995 3.91 66.145 5.025 ;
      RECT 65.995 3.757 66.14 5.025 ;
      RECT 66 3.742 66.14 5.025 ;
      RECT 66.05 3.457 66.14 5.025 ;
      RECT 66.005 3.692 66.14 5.025 ;
      RECT 66.035 3.51 66.14 5.025 ;
      RECT 66.02 3.622 66.14 5.025 ;
      RECT 66.025 3.58 66.14 5.025 ;
      RECT 66.02 3.622 66.155 3.685 ;
      RECT 66.055 3.21 66.16 3.63 ;
      RECT 66.055 3.21 66.175 3.613 ;
      RECT 66.055 3.21 66.21 3.575 ;
      RECT 66.05 3.457 66.26 3.508 ;
      RECT 66.055 3.21 66.315 3.47 ;
      RECT 65.315 3.915 65.575 4.175 ;
      RECT 65.315 3.915 65.585 4.133 ;
      RECT 65.315 3.915 65.671 4.104 ;
      RECT 65.315 3.915 65.74 4.056 ;
      RECT 65.315 3.915 65.775 4.025 ;
      RECT 65.545 3.735 65.825 4.015 ;
      RECT 65.38 3.9 65.825 4.015 ;
      RECT 65.47 3.777 65.575 4.175 ;
      RECT 65.4 3.84 65.825 4.015 ;
      RECT 59.85 8.51 60.17 8.835 ;
      RECT 59.88 7.985 60.05 8.835 ;
      RECT 59.88 7.985 60.055 8.335 ;
      RECT 59.88 7.985 60.855 8.16 ;
      RECT 60.68 3.26 60.855 8.16 ;
      RECT 60.625 3.26 60.975 3.61 ;
      RECT 60.65 8.945 60.975 9.27 ;
      RECT 59.535 9.035 60.975 9.205 ;
      RECT 59.535 3.69 59.695 9.205 ;
      RECT 59.85 3.66 60.17 3.98 ;
      RECT 59.535 3.69 60.17 3.86 ;
      RECT 58.2 4 58.585 4.35 ;
      RECT 58.19 4.065 58.585 4.265 ;
      RECT 58.335 3.995 58.505 4.35 ;
      RECT 56.645 3.735 56.925 4.015 ;
      RECT 56.64 3.735 56.925 3.968 ;
      RECT 56.62 3.735 56.925 3.945 ;
      RECT 56.61 3.735 56.925 3.925 ;
      RECT 56.6 3.735 56.925 3.91 ;
      RECT 56.575 3.735 56.925 3.883 ;
      RECT 56.565 3.735 56.925 3.858 ;
      RECT 56.52 3.59 56.8 3.85 ;
      RECT 56.52 3.685 56.9 3.85 ;
      RECT 56.52 3.63 56.845 3.85 ;
      RECT 56.52 3.622 56.84 3.85 ;
      RECT 56.52 3.612 56.835 3.85 ;
      RECT 56.52 3.6 56.83 3.85 ;
      RECT 55.445 4.295 55.725 4.575 ;
      RECT 55.445 4.295 55.76 4.555 ;
      RECT 47.77 8.95 48.12 9.3 ;
      RECT 55.19 8.905 55.54 9.255 ;
      RECT 47.77 8.98 55.54 9.18 ;
      RECT 55.48 3.715 55.53 3.975 ;
      RECT 55.27 3.715 55.275 3.975 ;
      RECT 54.465 3.27 54.495 3.53 ;
      RECT 54.235 3.27 54.31 3.53 ;
      RECT 55.455 3.665 55.48 3.975 ;
      RECT 55.45 3.622 55.455 3.975 ;
      RECT 55.445 3.605 55.45 3.975 ;
      RECT 55.44 3.592 55.445 3.975 ;
      RECT 55.365 3.475 55.44 3.975 ;
      RECT 55.32 3.292 55.365 3.975 ;
      RECT 55.315 3.22 55.32 3.975 ;
      RECT 55.3 3.195 55.315 3.975 ;
      RECT 55.275 3.157 55.3 3.975 ;
      RECT 55.265 3.137 55.275 3.697 ;
      RECT 55.25 3.129 55.265 3.652 ;
      RECT 55.245 3.121 55.25 3.623 ;
      RECT 55.24 3.118 55.245 3.603 ;
      RECT 55.235 3.115 55.24 3.583 ;
      RECT 55.23 3.112 55.235 3.563 ;
      RECT 55.2 3.101 55.23 3.5 ;
      RECT 55.18 3.086 55.2 3.415 ;
      RECT 55.175 3.078 55.18 3.378 ;
      RECT 55.165 3.072 55.175 3.345 ;
      RECT 55.15 3.064 55.165 3.305 ;
      RECT 55.145 3.057 55.15 3.265 ;
      RECT 55.14 3.054 55.145 3.243 ;
      RECT 55.135 3.051 55.14 3.23 ;
      RECT 55.13 3.05 55.135 3.22 ;
      RECT 55.115 3.044 55.13 3.21 ;
      RECT 55.09 3.031 55.115 3.195 ;
      RECT 55.04 3.006 55.09 3.166 ;
      RECT 55.025 2.985 55.04 3.141 ;
      RECT 55.015 2.978 55.025 3.13 ;
      RECT 54.96 2.959 55.015 3.103 ;
      RECT 54.935 2.937 54.96 3.076 ;
      RECT 54.93 2.93 54.935 3.071 ;
      RECT 54.915 2.93 54.93 3.069 ;
      RECT 54.89 2.922 54.915 3.065 ;
      RECT 54.875 2.92 54.89 3.061 ;
      RECT 54.845 2.92 54.875 3.058 ;
      RECT 54.835 2.92 54.845 3.053 ;
      RECT 54.79 2.92 54.835 3.051 ;
      RECT 54.761 2.92 54.79 3.052 ;
      RECT 54.675 2.92 54.761 3.054 ;
      RECT 54.661 2.921 54.675 3.056 ;
      RECT 54.575 2.922 54.661 3.058 ;
      RECT 54.56 2.923 54.575 3.068 ;
      RECT 54.555 2.924 54.56 3.077 ;
      RECT 54.535 2.927 54.555 3.087 ;
      RECT 54.52 2.935 54.535 3.102 ;
      RECT 54.5 2.953 54.52 3.117 ;
      RECT 54.49 2.965 54.5 3.14 ;
      RECT 54.48 2.974 54.49 3.17 ;
      RECT 54.465 2.986 54.48 3.215 ;
      RECT 54.41 3.019 54.465 3.53 ;
      RECT 54.405 3.047 54.41 3.53 ;
      RECT 54.385 3.062 54.405 3.53 ;
      RECT 54.35 3.122 54.385 3.53 ;
      RECT 54.348 3.172 54.35 3.53 ;
      RECT 54.345 3.18 54.348 3.53 ;
      RECT 54.335 3.195 54.345 3.53 ;
      RECT 54.33 3.207 54.335 3.53 ;
      RECT 54.32 3.232 54.33 3.53 ;
      RECT 54.31 3.26 54.32 3.53 ;
      RECT 52.215 4.765 52.265 5.025 ;
      RECT 55.125 4.315 55.185 4.575 ;
      RECT 55.11 4.315 55.125 4.585 ;
      RECT 55.091 4.315 55.11 4.618 ;
      RECT 55.005 4.315 55.091 4.743 ;
      RECT 54.925 4.315 55.005 4.925 ;
      RECT 54.92 4.552 54.925 5.01 ;
      RECT 54.895 4.622 54.92 5.038 ;
      RECT 54.89 4.692 54.895 5.065 ;
      RECT 54.87 4.764 54.89 5.087 ;
      RECT 54.865 4.831 54.87 5.11 ;
      RECT 54.855 4.86 54.865 5.125 ;
      RECT 54.845 4.882 54.855 5.142 ;
      RECT 54.84 4.892 54.845 5.153 ;
      RECT 54.835 4.9 54.84 5.161 ;
      RECT 54.825 4.908 54.835 5.173 ;
      RECT 54.82 4.92 54.825 5.183 ;
      RECT 54.815 4.928 54.82 5.188 ;
      RECT 54.795 4.946 54.815 5.198 ;
      RECT 54.79 4.963 54.795 5.205 ;
      RECT 54.785 4.971 54.79 5.206 ;
      RECT 54.78 4.982 54.785 5.208 ;
      RECT 54.74 5.02 54.78 5.218 ;
      RECT 54.735 5.055 54.74 5.229 ;
      RECT 54.73 5.06 54.735 5.232 ;
      RECT 54.705 5.07 54.73 5.239 ;
      RECT 54.695 5.084 54.705 5.248 ;
      RECT 54.675 5.096 54.695 5.251 ;
      RECT 54.625 5.115 54.675 5.255 ;
      RECT 54.58 5.13 54.625 5.26 ;
      RECT 54.515 5.133 54.58 5.266 ;
      RECT 54.5 5.131 54.515 5.273 ;
      RECT 54.47 5.13 54.5 5.273 ;
      RECT 54.431 5.129 54.47 5.269 ;
      RECT 54.345 5.126 54.431 5.265 ;
      RECT 54.328 5.124 54.345 5.262 ;
      RECT 54.242 5.122 54.328 5.259 ;
      RECT 54.156 5.119 54.242 5.253 ;
      RECT 54.07 5.115 54.156 5.248 ;
      RECT 53.992 5.112 54.07 5.244 ;
      RECT 53.906 5.109 53.992 5.242 ;
      RECT 53.82 5.106 53.906 5.239 ;
      RECT 53.762 5.104 53.82 5.236 ;
      RECT 53.676 5.101 53.762 5.234 ;
      RECT 53.59 5.097 53.676 5.232 ;
      RECT 53.504 5.094 53.59 5.229 ;
      RECT 53.418 5.09 53.504 5.227 ;
      RECT 53.332 5.086 53.418 5.224 ;
      RECT 53.246 5.083 53.332 5.222 ;
      RECT 53.16 5.079 53.246 5.219 ;
      RECT 53.074 5.076 53.16 5.217 ;
      RECT 52.988 5.072 53.074 5.214 ;
      RECT 52.902 5.069 52.988 5.212 ;
      RECT 52.816 5.065 52.902 5.209 ;
      RECT 52.73 5.062 52.816 5.207 ;
      RECT 52.72 5.06 52.73 5.203 ;
      RECT 52.715 5.06 52.72 5.201 ;
      RECT 52.675 5.055 52.715 5.195 ;
      RECT 52.661 5.046 52.675 5.188 ;
      RECT 52.575 5.016 52.661 5.173 ;
      RECT 52.555 4.982 52.575 5.158 ;
      RECT 52.485 4.951 52.555 5.145 ;
      RECT 52.48 4.926 52.485 5.134 ;
      RECT 52.475 4.92 52.48 5.132 ;
      RECT 52.406 4.765 52.475 5.12 ;
      RECT 52.32 4.765 52.406 5.094 ;
      RECT 52.295 4.765 52.32 5.073 ;
      RECT 52.29 4.765 52.295 5.063 ;
      RECT 52.285 4.765 52.29 5.055 ;
      RECT 52.265 4.765 52.285 5.038 ;
      RECT 54.685 3.335 54.945 3.595 ;
      RECT 54.67 3.335 54.945 3.498 ;
      RECT 54.64 3.335 54.945 3.473 ;
      RECT 54.605 3.175 54.885 3.455 ;
      RECT 54.575 4.665 54.635 4.925 ;
      RECT 53.6 3.355 53.655 3.615 ;
      RECT 54.535 4.622 54.575 4.925 ;
      RECT 54.506 4.543 54.535 4.925 ;
      RECT 54.42 4.415 54.506 4.925 ;
      RECT 54.4 4.295 54.42 4.925 ;
      RECT 54.375 4.246 54.4 4.925 ;
      RECT 54.37 4.211 54.375 4.775 ;
      RECT 54.34 4.171 54.37 4.713 ;
      RECT 54.315 4.108 54.34 4.628 ;
      RECT 54.305 4.07 54.315 4.565 ;
      RECT 54.29 4.045 54.305 4.526 ;
      RECT 54.247 4.003 54.29 4.432 ;
      RECT 54.245 3.976 54.247 4.359 ;
      RECT 54.24 3.971 54.245 4.35 ;
      RECT 54.235 3.964 54.24 4.325 ;
      RECT 54.23 3.958 54.235 4.31 ;
      RECT 54.225 3.952 54.23 4.298 ;
      RECT 54.215 3.943 54.225 4.28 ;
      RECT 54.21 3.934 54.215 4.258 ;
      RECT 54.185 3.915 54.21 4.208 ;
      RECT 54.18 3.896 54.185 4.158 ;
      RECT 54.165 3.882 54.18 4.118 ;
      RECT 54.16 3.868 54.165 4.085 ;
      RECT 54.155 3.861 54.16 4.078 ;
      RECT 54.14 3.848 54.155 4.07 ;
      RECT 54.095 3.81 54.14 4.043 ;
      RECT 54.065 3.763 54.095 4.008 ;
      RECT 54.045 3.732 54.065 3.985 ;
      RECT 53.965 3.665 54.045 3.938 ;
      RECT 53.935 3.595 53.965 3.885 ;
      RECT 53.93 3.572 53.935 3.868 ;
      RECT 53.9 3.55 53.93 3.853 ;
      RECT 53.87 3.509 53.9 3.825 ;
      RECT 53.865 3.484 53.87 3.81 ;
      RECT 53.86 3.478 53.865 3.803 ;
      RECT 53.85 3.355 53.86 3.795 ;
      RECT 53.84 3.355 53.85 3.788 ;
      RECT 53.835 3.355 53.84 3.78 ;
      RECT 53.815 3.355 53.835 3.768 ;
      RECT 53.765 3.355 53.815 3.738 ;
      RECT 53.71 3.355 53.765 3.688 ;
      RECT 53.68 3.355 53.71 3.648 ;
      RECT 53.655 3.355 53.68 3.625 ;
      RECT 53.525 4.08 53.805 4.36 ;
      RECT 53.49 3.995 53.75 4.255 ;
      RECT 53.49 4.077 53.76 4.255 ;
      RECT 51.69 3.45 51.695 3.935 ;
      RECT 51.58 3.635 51.585 3.935 ;
      RECT 51.49 3.675 51.555 3.935 ;
      RECT 53.165 3.175 53.255 3.805 ;
      RECT 53.13 3.225 53.135 3.805 ;
      RECT 53.075 3.25 53.085 3.805 ;
      RECT 53.03 3.25 53.04 3.805 ;
      RECT 53.4 3.175 53.445 3.455 ;
      RECT 52.25 2.905 52.45 3.045 ;
      RECT 53.366 3.175 53.4 3.467 ;
      RECT 53.28 3.175 53.366 3.507 ;
      RECT 53.265 3.175 53.28 3.548 ;
      RECT 53.26 3.175 53.265 3.568 ;
      RECT 53.255 3.175 53.26 3.588 ;
      RECT 53.135 3.217 53.165 3.805 ;
      RECT 53.085 3.237 53.13 3.805 ;
      RECT 53.07 3.252 53.075 3.805 ;
      RECT 53.04 3.252 53.07 3.805 ;
      RECT 52.995 3.237 53.03 3.805 ;
      RECT 52.99 3.225 52.995 3.585 ;
      RECT 52.985 3.222 52.99 3.565 ;
      RECT 52.97 3.212 52.985 3.518 ;
      RECT 52.965 3.205 52.97 3.481 ;
      RECT 52.96 3.202 52.965 3.464 ;
      RECT 52.945 3.192 52.96 3.42 ;
      RECT 52.94 3.183 52.945 3.38 ;
      RECT 52.935 3.179 52.94 3.365 ;
      RECT 52.925 3.173 52.935 3.348 ;
      RECT 52.885 3.154 52.925 3.323 ;
      RECT 52.88 3.136 52.885 3.303 ;
      RECT 52.87 3.13 52.88 3.298 ;
      RECT 52.84 3.114 52.87 3.285 ;
      RECT 52.825 3.096 52.84 3.268 ;
      RECT 52.81 3.084 52.825 3.255 ;
      RECT 52.805 3.076 52.81 3.248 ;
      RECT 52.775 3.062 52.805 3.235 ;
      RECT 52.77 3.047 52.775 3.223 ;
      RECT 52.76 3.041 52.77 3.215 ;
      RECT 52.74 3.029 52.76 3.203 ;
      RECT 52.73 3.017 52.74 3.19 ;
      RECT 52.7 3.001 52.73 3.175 ;
      RECT 52.68 2.981 52.7 3.158 ;
      RECT 52.675 2.971 52.68 3.148 ;
      RECT 52.65 2.959 52.675 3.135 ;
      RECT 52.645 2.947 52.65 3.123 ;
      RECT 52.64 2.942 52.645 3.119 ;
      RECT 52.625 2.935 52.64 3.111 ;
      RECT 52.615 2.922 52.625 3.101 ;
      RECT 52.61 2.92 52.615 3.095 ;
      RECT 52.585 2.913 52.61 3.084 ;
      RECT 52.58 2.906 52.585 3.073 ;
      RECT 52.555 2.905 52.58 3.06 ;
      RECT 52.536 2.905 52.555 3.05 ;
      RECT 52.45 2.905 52.536 3.047 ;
      RECT 52.22 2.905 52.25 3.05 ;
      RECT 52.18 2.912 52.22 3.063 ;
      RECT 52.155 2.922 52.18 3.076 ;
      RECT 52.14 2.931 52.155 3.086 ;
      RECT 52.11 2.936 52.14 3.105 ;
      RECT 52.105 2.942 52.11 3.123 ;
      RECT 52.085 2.952 52.105 3.138 ;
      RECT 52.075 2.965 52.085 3.158 ;
      RECT 52.06 2.977 52.075 3.175 ;
      RECT 52.055 2.987 52.06 3.185 ;
      RECT 52.05 2.992 52.055 3.19 ;
      RECT 52.04 3 52.05 3.203 ;
      RECT 51.99 3.032 52.04 3.24 ;
      RECT 51.975 3.067 51.99 3.281 ;
      RECT 51.97 3.077 51.975 3.296 ;
      RECT 51.965 3.082 51.97 3.303 ;
      RECT 51.94 3.098 51.965 3.323 ;
      RECT 51.925 3.119 51.94 3.348 ;
      RECT 51.9 3.14 51.925 3.373 ;
      RECT 51.89 3.159 51.9 3.396 ;
      RECT 51.865 3.177 51.89 3.419 ;
      RECT 51.85 3.197 51.865 3.443 ;
      RECT 51.845 3.207 51.85 3.455 ;
      RECT 51.83 3.219 51.845 3.475 ;
      RECT 51.82 3.234 51.83 3.515 ;
      RECT 51.815 3.242 51.82 3.543 ;
      RECT 51.805 3.252 51.815 3.563 ;
      RECT 51.8 3.265 51.805 3.588 ;
      RECT 51.795 3.278 51.8 3.608 ;
      RECT 51.79 3.284 51.795 3.63 ;
      RECT 51.78 3.293 51.79 3.65 ;
      RECT 51.775 3.313 51.78 3.673 ;
      RECT 51.77 3.319 51.775 3.693 ;
      RECT 51.765 3.326 51.77 3.715 ;
      RECT 51.76 3.337 51.765 3.728 ;
      RECT 51.75 3.347 51.76 3.753 ;
      RECT 51.73 3.372 51.75 3.935 ;
      RECT 51.7 3.412 51.73 3.935 ;
      RECT 51.695 3.442 51.7 3.935 ;
      RECT 51.67 3.47 51.69 3.935 ;
      RECT 51.64 3.515 51.67 3.935 ;
      RECT 51.635 3.542 51.64 3.935 ;
      RECT 51.615 3.56 51.635 3.935 ;
      RECT 51.605 3.585 51.615 3.935 ;
      RECT 51.6 3.597 51.605 3.935 ;
      RECT 51.585 3.62 51.6 3.935 ;
      RECT 51.565 3.647 51.58 3.935 ;
      RECT 51.555 3.67 51.565 3.935 ;
      RECT 53.345 4.555 53.425 4.815 ;
      RECT 52.58 3.775 52.65 4.035 ;
      RECT 53.311 4.522 53.345 4.815 ;
      RECT 53.225 4.425 53.311 4.815 ;
      RECT 53.205 4.337 53.225 4.815 ;
      RECT 53.195 4.307 53.205 4.815 ;
      RECT 53.185 4.287 53.195 4.815 ;
      RECT 53.165 4.274 53.185 4.815 ;
      RECT 53.15 4.264 53.165 4.643 ;
      RECT 53.145 4.257 53.15 4.598 ;
      RECT 53.135 4.251 53.145 4.588 ;
      RECT 53.125 4.243 53.135 4.57 ;
      RECT 53.12 4.237 53.125 4.558 ;
      RECT 53.11 4.232 53.12 4.545 ;
      RECT 53.09 4.222 53.11 4.518 ;
      RECT 53.05 4.201 53.09 4.47 ;
      RECT 53.035 4.182 53.05 4.428 ;
      RECT 53.01 4.168 53.035 4.398 ;
      RECT 53 4.156 53.01 4.365 ;
      RECT 52.995 4.151 53 4.355 ;
      RECT 52.965 4.137 52.995 4.335 ;
      RECT 52.955 4.121 52.965 4.308 ;
      RECT 52.95 4.116 52.955 4.298 ;
      RECT 52.925 4.107 52.95 4.278 ;
      RECT 52.915 4.095 52.925 4.258 ;
      RECT 52.845 4.063 52.915 4.233 ;
      RECT 52.84 4.032 52.845 4.21 ;
      RECT 52.791 3.775 52.84 4.193 ;
      RECT 52.705 3.775 52.791 4.152 ;
      RECT 52.65 3.775 52.705 4.08 ;
      RECT 52.74 4.56 52.9 4.82 ;
      RECT 52.265 3.175 52.315 3.86 ;
      RECT 52.055 3.6 52.09 3.86 ;
      RECT 52.37 3.175 52.375 3.635 ;
      RECT 52.46 3.175 52.485 3.455 ;
      RECT 52.735 4.557 52.74 4.82 ;
      RECT 52.7 4.545 52.735 4.82 ;
      RECT 52.64 4.518 52.7 4.82 ;
      RECT 52.635 4.501 52.64 4.674 ;
      RECT 52.63 4.498 52.635 4.661 ;
      RECT 52.61 4.491 52.63 4.648 ;
      RECT 52.575 4.474 52.61 4.63 ;
      RECT 52.535 4.453 52.575 4.61 ;
      RECT 52.53 4.441 52.535 4.598 ;
      RECT 52.49 4.427 52.53 4.584 ;
      RECT 52.47 4.41 52.49 4.566 ;
      RECT 52.46 4.402 52.47 4.558 ;
      RECT 52.445 3.175 52.46 3.473 ;
      RECT 52.43 4.392 52.46 4.545 ;
      RECT 52.415 3.175 52.445 3.518 ;
      RECT 52.42 4.382 52.43 4.532 ;
      RECT 52.39 4.367 52.42 4.519 ;
      RECT 52.375 3.175 52.415 3.585 ;
      RECT 52.375 4.335 52.39 4.505 ;
      RECT 52.37 4.307 52.375 4.499 ;
      RECT 52.365 3.175 52.37 3.64 ;
      RECT 52.355 4.277 52.37 4.493 ;
      RECT 52.36 3.175 52.365 3.653 ;
      RECT 52.35 3.175 52.36 3.673 ;
      RECT 52.315 4.19 52.355 4.478 ;
      RECT 52.315 3.175 52.35 3.713 ;
      RECT 52.31 4.122 52.315 4.466 ;
      RECT 52.295 4.077 52.31 4.461 ;
      RECT 52.29 4.015 52.295 4.456 ;
      RECT 52.265 3.922 52.29 4.449 ;
      RECT 52.26 3.175 52.265 4.441 ;
      RECT 52.245 3.175 52.26 4.428 ;
      RECT 52.225 3.175 52.245 4.385 ;
      RECT 52.215 3.175 52.225 4.335 ;
      RECT 52.21 3.175 52.215 4.308 ;
      RECT 52.205 3.175 52.21 4.286 ;
      RECT 52.2 3.401 52.205 4.269 ;
      RECT 52.195 3.423 52.2 4.247 ;
      RECT 52.19 3.465 52.195 4.23 ;
      RECT 52.16 3.515 52.19 4.174 ;
      RECT 52.155 3.542 52.16 4.116 ;
      RECT 52.14 3.56 52.155 4.08 ;
      RECT 52.135 3.578 52.14 4.044 ;
      RECT 52.129 3.585 52.135 4.025 ;
      RECT 52.125 3.592 52.129 4.008 ;
      RECT 52.12 3.597 52.125 3.977 ;
      RECT 52.11 3.6 52.12 3.952 ;
      RECT 52.1 3.6 52.11 3.918 ;
      RECT 52.095 3.6 52.1 3.895 ;
      RECT 52.09 3.6 52.095 3.875 ;
      RECT 50.71 4.765 50.97 5.025 ;
      RECT 50.73 4.692 50.91 5.025 ;
      RECT 50.73 4.435 50.905 5.025 ;
      RECT 50.73 4.227 50.895 5.025 ;
      RECT 50.735 4.145 50.895 5.025 ;
      RECT 50.735 3.91 50.885 5.025 ;
      RECT 50.735 3.757 50.88 5.025 ;
      RECT 50.74 3.742 50.88 5.025 ;
      RECT 50.79 3.457 50.88 5.025 ;
      RECT 50.745 3.692 50.88 5.025 ;
      RECT 50.775 3.51 50.88 5.025 ;
      RECT 50.76 3.622 50.88 5.025 ;
      RECT 50.765 3.58 50.88 5.025 ;
      RECT 50.76 3.622 50.895 3.685 ;
      RECT 50.795 3.21 50.9 3.63 ;
      RECT 50.795 3.21 50.915 3.613 ;
      RECT 50.795 3.21 50.95 3.575 ;
      RECT 50.79 3.457 51 3.508 ;
      RECT 50.795 3.21 51.055 3.47 ;
      RECT 50.055 3.915 50.315 4.175 ;
      RECT 50.055 3.915 50.325 4.133 ;
      RECT 50.055 3.915 50.411 4.104 ;
      RECT 50.055 3.915 50.48 4.056 ;
      RECT 50.055 3.915 50.515 4.025 ;
      RECT 50.285 3.735 50.565 4.015 ;
      RECT 50.12 3.9 50.565 4.015 ;
      RECT 50.21 3.777 50.315 4.175 ;
      RECT 50.14 3.84 50.565 4.015 ;
      RECT 44.59 8.51 44.91 8.835 ;
      RECT 44.62 7.985 44.79 8.835 ;
      RECT 44.62 7.985 44.795 8.335 ;
      RECT 44.62 7.985 45.595 8.16 ;
      RECT 45.42 3.26 45.595 8.16 ;
      RECT 45.365 3.26 45.715 3.61 ;
      RECT 45.39 8.945 45.715 9.27 ;
      RECT 44.275 9.035 45.715 9.205 ;
      RECT 44.275 3.69 44.435 9.205 ;
      RECT 44.59 3.66 44.91 3.98 ;
      RECT 44.275 3.69 44.91 3.86 ;
      RECT 42.94 4 43.325 4.35 ;
      RECT 42.93 4.065 43.325 4.265 ;
      RECT 43.075 3.995 43.245 4.35 ;
      RECT 41.385 3.735 41.665 4.015 ;
      RECT 41.38 3.735 41.665 3.968 ;
      RECT 41.36 3.735 41.665 3.945 ;
      RECT 41.35 3.735 41.665 3.925 ;
      RECT 41.34 3.735 41.665 3.91 ;
      RECT 41.315 3.735 41.665 3.883 ;
      RECT 41.305 3.735 41.665 3.858 ;
      RECT 41.26 3.59 41.54 3.85 ;
      RECT 41.26 3.685 41.64 3.85 ;
      RECT 41.26 3.63 41.585 3.85 ;
      RECT 41.26 3.622 41.58 3.85 ;
      RECT 41.26 3.612 41.575 3.85 ;
      RECT 41.26 3.6 41.57 3.85 ;
      RECT 40.185 4.295 40.465 4.575 ;
      RECT 40.185 4.295 40.5 4.555 ;
      RECT 32.51 8.95 32.86 9.3 ;
      RECT 39.93 8.905 40.28 9.255 ;
      RECT 32.51 8.98 40.28 9.18 ;
      RECT 40.22 3.715 40.27 3.975 ;
      RECT 40.01 3.715 40.015 3.975 ;
      RECT 39.205 3.27 39.235 3.53 ;
      RECT 38.975 3.27 39.05 3.53 ;
      RECT 40.195 3.665 40.22 3.975 ;
      RECT 40.19 3.622 40.195 3.975 ;
      RECT 40.185 3.605 40.19 3.975 ;
      RECT 40.18 3.592 40.185 3.975 ;
      RECT 40.105 3.475 40.18 3.975 ;
      RECT 40.06 3.292 40.105 3.975 ;
      RECT 40.055 3.22 40.06 3.975 ;
      RECT 40.04 3.195 40.055 3.975 ;
      RECT 40.015 3.157 40.04 3.975 ;
      RECT 40.005 3.137 40.015 3.697 ;
      RECT 39.99 3.129 40.005 3.652 ;
      RECT 39.985 3.121 39.99 3.623 ;
      RECT 39.98 3.118 39.985 3.603 ;
      RECT 39.975 3.115 39.98 3.583 ;
      RECT 39.97 3.112 39.975 3.563 ;
      RECT 39.94 3.101 39.97 3.5 ;
      RECT 39.92 3.086 39.94 3.415 ;
      RECT 39.915 3.078 39.92 3.378 ;
      RECT 39.905 3.072 39.915 3.345 ;
      RECT 39.89 3.064 39.905 3.305 ;
      RECT 39.885 3.057 39.89 3.265 ;
      RECT 39.88 3.054 39.885 3.243 ;
      RECT 39.875 3.051 39.88 3.23 ;
      RECT 39.87 3.05 39.875 3.22 ;
      RECT 39.855 3.044 39.87 3.21 ;
      RECT 39.83 3.031 39.855 3.195 ;
      RECT 39.78 3.006 39.83 3.166 ;
      RECT 39.765 2.985 39.78 3.141 ;
      RECT 39.755 2.978 39.765 3.13 ;
      RECT 39.7 2.959 39.755 3.103 ;
      RECT 39.675 2.937 39.7 3.076 ;
      RECT 39.67 2.93 39.675 3.071 ;
      RECT 39.655 2.93 39.67 3.069 ;
      RECT 39.63 2.922 39.655 3.065 ;
      RECT 39.615 2.92 39.63 3.061 ;
      RECT 39.585 2.92 39.615 3.058 ;
      RECT 39.575 2.92 39.585 3.053 ;
      RECT 39.53 2.92 39.575 3.051 ;
      RECT 39.501 2.92 39.53 3.052 ;
      RECT 39.415 2.92 39.501 3.054 ;
      RECT 39.401 2.921 39.415 3.056 ;
      RECT 39.315 2.922 39.401 3.058 ;
      RECT 39.3 2.923 39.315 3.068 ;
      RECT 39.295 2.924 39.3 3.077 ;
      RECT 39.275 2.927 39.295 3.087 ;
      RECT 39.26 2.935 39.275 3.102 ;
      RECT 39.24 2.953 39.26 3.117 ;
      RECT 39.23 2.965 39.24 3.14 ;
      RECT 39.22 2.974 39.23 3.17 ;
      RECT 39.205 2.986 39.22 3.215 ;
      RECT 39.15 3.019 39.205 3.53 ;
      RECT 39.145 3.047 39.15 3.53 ;
      RECT 39.125 3.062 39.145 3.53 ;
      RECT 39.09 3.122 39.125 3.53 ;
      RECT 39.088 3.172 39.09 3.53 ;
      RECT 39.085 3.18 39.088 3.53 ;
      RECT 39.075 3.195 39.085 3.53 ;
      RECT 39.07 3.207 39.075 3.53 ;
      RECT 39.06 3.232 39.07 3.53 ;
      RECT 39.05 3.26 39.06 3.53 ;
      RECT 36.955 4.765 37.005 5.025 ;
      RECT 39.865 4.315 39.925 4.575 ;
      RECT 39.85 4.315 39.865 4.585 ;
      RECT 39.831 4.315 39.85 4.618 ;
      RECT 39.745 4.315 39.831 4.743 ;
      RECT 39.665 4.315 39.745 4.925 ;
      RECT 39.66 4.552 39.665 5.01 ;
      RECT 39.635 4.622 39.66 5.038 ;
      RECT 39.63 4.692 39.635 5.065 ;
      RECT 39.61 4.764 39.63 5.087 ;
      RECT 39.605 4.831 39.61 5.11 ;
      RECT 39.595 4.86 39.605 5.125 ;
      RECT 39.585 4.882 39.595 5.142 ;
      RECT 39.58 4.892 39.585 5.153 ;
      RECT 39.575 4.9 39.58 5.161 ;
      RECT 39.565 4.908 39.575 5.173 ;
      RECT 39.56 4.92 39.565 5.183 ;
      RECT 39.555 4.928 39.56 5.188 ;
      RECT 39.535 4.946 39.555 5.198 ;
      RECT 39.53 4.963 39.535 5.205 ;
      RECT 39.525 4.971 39.53 5.206 ;
      RECT 39.52 4.982 39.525 5.208 ;
      RECT 39.48 5.02 39.52 5.218 ;
      RECT 39.475 5.055 39.48 5.229 ;
      RECT 39.47 5.06 39.475 5.232 ;
      RECT 39.445 5.07 39.47 5.239 ;
      RECT 39.435 5.084 39.445 5.248 ;
      RECT 39.415 5.096 39.435 5.251 ;
      RECT 39.365 5.115 39.415 5.255 ;
      RECT 39.32 5.13 39.365 5.26 ;
      RECT 39.255 5.133 39.32 5.266 ;
      RECT 39.24 5.131 39.255 5.273 ;
      RECT 39.21 5.13 39.24 5.273 ;
      RECT 39.171 5.129 39.21 5.269 ;
      RECT 39.085 5.126 39.171 5.265 ;
      RECT 39.068 5.124 39.085 5.262 ;
      RECT 38.982 5.122 39.068 5.259 ;
      RECT 38.896 5.119 38.982 5.253 ;
      RECT 38.81 5.115 38.896 5.248 ;
      RECT 38.732 5.112 38.81 5.244 ;
      RECT 38.646 5.109 38.732 5.242 ;
      RECT 38.56 5.106 38.646 5.239 ;
      RECT 38.502 5.104 38.56 5.236 ;
      RECT 38.416 5.101 38.502 5.234 ;
      RECT 38.33 5.097 38.416 5.232 ;
      RECT 38.244 5.094 38.33 5.229 ;
      RECT 38.158 5.09 38.244 5.227 ;
      RECT 38.072 5.086 38.158 5.224 ;
      RECT 37.986 5.083 38.072 5.222 ;
      RECT 37.9 5.079 37.986 5.219 ;
      RECT 37.814 5.076 37.9 5.217 ;
      RECT 37.728 5.072 37.814 5.214 ;
      RECT 37.642 5.069 37.728 5.212 ;
      RECT 37.556 5.065 37.642 5.209 ;
      RECT 37.47 5.062 37.556 5.207 ;
      RECT 37.46 5.06 37.47 5.203 ;
      RECT 37.455 5.06 37.46 5.201 ;
      RECT 37.415 5.055 37.455 5.195 ;
      RECT 37.401 5.046 37.415 5.188 ;
      RECT 37.315 5.016 37.401 5.173 ;
      RECT 37.295 4.982 37.315 5.158 ;
      RECT 37.225 4.951 37.295 5.145 ;
      RECT 37.22 4.926 37.225 5.134 ;
      RECT 37.215 4.92 37.22 5.132 ;
      RECT 37.146 4.765 37.215 5.12 ;
      RECT 37.06 4.765 37.146 5.094 ;
      RECT 37.035 4.765 37.06 5.073 ;
      RECT 37.03 4.765 37.035 5.063 ;
      RECT 37.025 4.765 37.03 5.055 ;
      RECT 37.005 4.765 37.025 5.038 ;
      RECT 39.425 3.335 39.685 3.595 ;
      RECT 39.41 3.335 39.685 3.498 ;
      RECT 39.38 3.335 39.685 3.473 ;
      RECT 39.345 3.175 39.625 3.455 ;
      RECT 39.315 4.665 39.375 4.925 ;
      RECT 38.34 3.355 38.395 3.615 ;
      RECT 39.275 4.622 39.315 4.925 ;
      RECT 39.246 4.543 39.275 4.925 ;
      RECT 39.16 4.415 39.246 4.925 ;
      RECT 39.14 4.295 39.16 4.925 ;
      RECT 39.115 4.246 39.14 4.925 ;
      RECT 39.11 4.211 39.115 4.775 ;
      RECT 39.08 4.171 39.11 4.713 ;
      RECT 39.055 4.108 39.08 4.628 ;
      RECT 39.045 4.07 39.055 4.565 ;
      RECT 39.03 4.045 39.045 4.526 ;
      RECT 38.987 4.003 39.03 4.432 ;
      RECT 38.985 3.976 38.987 4.359 ;
      RECT 38.98 3.971 38.985 4.35 ;
      RECT 38.975 3.964 38.98 4.325 ;
      RECT 38.97 3.958 38.975 4.31 ;
      RECT 38.965 3.952 38.97 4.298 ;
      RECT 38.955 3.943 38.965 4.28 ;
      RECT 38.95 3.934 38.955 4.258 ;
      RECT 38.925 3.915 38.95 4.208 ;
      RECT 38.92 3.896 38.925 4.158 ;
      RECT 38.905 3.882 38.92 4.118 ;
      RECT 38.9 3.868 38.905 4.085 ;
      RECT 38.895 3.861 38.9 4.078 ;
      RECT 38.88 3.848 38.895 4.07 ;
      RECT 38.835 3.81 38.88 4.043 ;
      RECT 38.805 3.763 38.835 4.008 ;
      RECT 38.785 3.732 38.805 3.985 ;
      RECT 38.705 3.665 38.785 3.938 ;
      RECT 38.675 3.595 38.705 3.885 ;
      RECT 38.67 3.572 38.675 3.868 ;
      RECT 38.64 3.55 38.67 3.853 ;
      RECT 38.61 3.509 38.64 3.825 ;
      RECT 38.605 3.484 38.61 3.81 ;
      RECT 38.6 3.478 38.605 3.803 ;
      RECT 38.59 3.355 38.6 3.795 ;
      RECT 38.58 3.355 38.59 3.788 ;
      RECT 38.575 3.355 38.58 3.78 ;
      RECT 38.555 3.355 38.575 3.768 ;
      RECT 38.505 3.355 38.555 3.738 ;
      RECT 38.45 3.355 38.505 3.688 ;
      RECT 38.42 3.355 38.45 3.648 ;
      RECT 38.395 3.355 38.42 3.625 ;
      RECT 38.265 4.08 38.545 4.36 ;
      RECT 38.23 3.995 38.49 4.255 ;
      RECT 38.23 4.077 38.5 4.255 ;
      RECT 36.43 3.45 36.435 3.935 ;
      RECT 36.32 3.635 36.325 3.935 ;
      RECT 36.23 3.675 36.295 3.935 ;
      RECT 37.905 3.175 37.995 3.805 ;
      RECT 37.87 3.225 37.875 3.805 ;
      RECT 37.815 3.25 37.825 3.805 ;
      RECT 37.77 3.25 37.78 3.805 ;
      RECT 38.14 3.175 38.185 3.455 ;
      RECT 36.99 2.905 37.19 3.045 ;
      RECT 38.106 3.175 38.14 3.467 ;
      RECT 38.02 3.175 38.106 3.507 ;
      RECT 38.005 3.175 38.02 3.548 ;
      RECT 38 3.175 38.005 3.568 ;
      RECT 37.995 3.175 38 3.588 ;
      RECT 37.875 3.217 37.905 3.805 ;
      RECT 37.825 3.237 37.87 3.805 ;
      RECT 37.81 3.252 37.815 3.805 ;
      RECT 37.78 3.252 37.81 3.805 ;
      RECT 37.735 3.237 37.77 3.805 ;
      RECT 37.73 3.225 37.735 3.585 ;
      RECT 37.725 3.222 37.73 3.565 ;
      RECT 37.71 3.212 37.725 3.518 ;
      RECT 37.705 3.205 37.71 3.481 ;
      RECT 37.7 3.202 37.705 3.464 ;
      RECT 37.685 3.192 37.7 3.42 ;
      RECT 37.68 3.183 37.685 3.38 ;
      RECT 37.675 3.179 37.68 3.365 ;
      RECT 37.665 3.173 37.675 3.348 ;
      RECT 37.625 3.154 37.665 3.323 ;
      RECT 37.62 3.136 37.625 3.303 ;
      RECT 37.61 3.13 37.62 3.298 ;
      RECT 37.58 3.114 37.61 3.285 ;
      RECT 37.565 3.096 37.58 3.268 ;
      RECT 37.55 3.084 37.565 3.255 ;
      RECT 37.545 3.076 37.55 3.248 ;
      RECT 37.515 3.062 37.545 3.235 ;
      RECT 37.51 3.047 37.515 3.223 ;
      RECT 37.5 3.041 37.51 3.215 ;
      RECT 37.48 3.029 37.5 3.203 ;
      RECT 37.47 3.017 37.48 3.19 ;
      RECT 37.44 3.001 37.47 3.175 ;
      RECT 37.42 2.981 37.44 3.158 ;
      RECT 37.415 2.971 37.42 3.148 ;
      RECT 37.39 2.959 37.415 3.135 ;
      RECT 37.385 2.947 37.39 3.123 ;
      RECT 37.38 2.942 37.385 3.119 ;
      RECT 37.365 2.935 37.38 3.111 ;
      RECT 37.355 2.922 37.365 3.101 ;
      RECT 37.35 2.92 37.355 3.095 ;
      RECT 37.325 2.913 37.35 3.084 ;
      RECT 37.32 2.906 37.325 3.073 ;
      RECT 37.295 2.905 37.32 3.06 ;
      RECT 37.276 2.905 37.295 3.05 ;
      RECT 37.19 2.905 37.276 3.047 ;
      RECT 36.96 2.905 36.99 3.05 ;
      RECT 36.92 2.912 36.96 3.063 ;
      RECT 36.895 2.922 36.92 3.076 ;
      RECT 36.88 2.931 36.895 3.086 ;
      RECT 36.85 2.936 36.88 3.105 ;
      RECT 36.845 2.942 36.85 3.123 ;
      RECT 36.825 2.952 36.845 3.138 ;
      RECT 36.815 2.965 36.825 3.158 ;
      RECT 36.8 2.977 36.815 3.175 ;
      RECT 36.795 2.987 36.8 3.185 ;
      RECT 36.79 2.992 36.795 3.19 ;
      RECT 36.78 3 36.79 3.203 ;
      RECT 36.73 3.032 36.78 3.24 ;
      RECT 36.715 3.067 36.73 3.281 ;
      RECT 36.71 3.077 36.715 3.296 ;
      RECT 36.705 3.082 36.71 3.303 ;
      RECT 36.68 3.098 36.705 3.323 ;
      RECT 36.665 3.119 36.68 3.348 ;
      RECT 36.64 3.14 36.665 3.373 ;
      RECT 36.63 3.159 36.64 3.396 ;
      RECT 36.605 3.177 36.63 3.419 ;
      RECT 36.59 3.197 36.605 3.443 ;
      RECT 36.585 3.207 36.59 3.455 ;
      RECT 36.57 3.219 36.585 3.475 ;
      RECT 36.56 3.234 36.57 3.515 ;
      RECT 36.555 3.242 36.56 3.543 ;
      RECT 36.545 3.252 36.555 3.563 ;
      RECT 36.54 3.265 36.545 3.588 ;
      RECT 36.535 3.278 36.54 3.608 ;
      RECT 36.53 3.284 36.535 3.63 ;
      RECT 36.52 3.293 36.53 3.65 ;
      RECT 36.515 3.313 36.52 3.673 ;
      RECT 36.51 3.319 36.515 3.693 ;
      RECT 36.505 3.326 36.51 3.715 ;
      RECT 36.5 3.337 36.505 3.728 ;
      RECT 36.49 3.347 36.5 3.753 ;
      RECT 36.47 3.372 36.49 3.935 ;
      RECT 36.44 3.412 36.47 3.935 ;
      RECT 36.435 3.442 36.44 3.935 ;
      RECT 36.41 3.47 36.43 3.935 ;
      RECT 36.38 3.515 36.41 3.935 ;
      RECT 36.375 3.542 36.38 3.935 ;
      RECT 36.355 3.56 36.375 3.935 ;
      RECT 36.345 3.585 36.355 3.935 ;
      RECT 36.34 3.597 36.345 3.935 ;
      RECT 36.325 3.62 36.34 3.935 ;
      RECT 36.305 3.647 36.32 3.935 ;
      RECT 36.295 3.67 36.305 3.935 ;
      RECT 38.085 4.555 38.165 4.815 ;
      RECT 37.32 3.775 37.39 4.035 ;
      RECT 38.051 4.522 38.085 4.815 ;
      RECT 37.965 4.425 38.051 4.815 ;
      RECT 37.945 4.337 37.965 4.815 ;
      RECT 37.935 4.307 37.945 4.815 ;
      RECT 37.925 4.287 37.935 4.815 ;
      RECT 37.905 4.274 37.925 4.815 ;
      RECT 37.89 4.264 37.905 4.643 ;
      RECT 37.885 4.257 37.89 4.598 ;
      RECT 37.875 4.251 37.885 4.588 ;
      RECT 37.865 4.243 37.875 4.57 ;
      RECT 37.86 4.237 37.865 4.558 ;
      RECT 37.85 4.232 37.86 4.545 ;
      RECT 37.83 4.222 37.85 4.518 ;
      RECT 37.79 4.201 37.83 4.47 ;
      RECT 37.775 4.182 37.79 4.428 ;
      RECT 37.75 4.168 37.775 4.398 ;
      RECT 37.74 4.156 37.75 4.365 ;
      RECT 37.735 4.151 37.74 4.355 ;
      RECT 37.705 4.137 37.735 4.335 ;
      RECT 37.695 4.121 37.705 4.308 ;
      RECT 37.69 4.116 37.695 4.298 ;
      RECT 37.665 4.107 37.69 4.278 ;
      RECT 37.655 4.095 37.665 4.258 ;
      RECT 37.585 4.063 37.655 4.233 ;
      RECT 37.58 4.032 37.585 4.21 ;
      RECT 37.531 3.775 37.58 4.193 ;
      RECT 37.445 3.775 37.531 4.152 ;
      RECT 37.39 3.775 37.445 4.08 ;
      RECT 37.48 4.56 37.64 4.82 ;
      RECT 37.005 3.175 37.055 3.86 ;
      RECT 36.795 3.6 36.83 3.86 ;
      RECT 37.11 3.175 37.115 3.635 ;
      RECT 37.2 3.175 37.225 3.455 ;
      RECT 37.475 4.557 37.48 4.82 ;
      RECT 37.44 4.545 37.475 4.82 ;
      RECT 37.38 4.518 37.44 4.82 ;
      RECT 37.375 4.501 37.38 4.674 ;
      RECT 37.37 4.498 37.375 4.661 ;
      RECT 37.35 4.491 37.37 4.648 ;
      RECT 37.315 4.474 37.35 4.63 ;
      RECT 37.275 4.453 37.315 4.61 ;
      RECT 37.27 4.441 37.275 4.598 ;
      RECT 37.23 4.427 37.27 4.584 ;
      RECT 37.21 4.41 37.23 4.566 ;
      RECT 37.2 4.402 37.21 4.558 ;
      RECT 37.185 3.175 37.2 3.473 ;
      RECT 37.17 4.392 37.2 4.545 ;
      RECT 37.155 3.175 37.185 3.518 ;
      RECT 37.16 4.382 37.17 4.532 ;
      RECT 37.13 4.367 37.16 4.519 ;
      RECT 37.115 3.175 37.155 3.585 ;
      RECT 37.115 4.335 37.13 4.505 ;
      RECT 37.11 4.307 37.115 4.499 ;
      RECT 37.105 3.175 37.11 3.64 ;
      RECT 37.095 4.277 37.11 4.493 ;
      RECT 37.1 3.175 37.105 3.653 ;
      RECT 37.09 3.175 37.1 3.673 ;
      RECT 37.055 4.19 37.095 4.478 ;
      RECT 37.055 3.175 37.09 3.713 ;
      RECT 37.05 4.122 37.055 4.466 ;
      RECT 37.035 4.077 37.05 4.461 ;
      RECT 37.03 4.015 37.035 4.456 ;
      RECT 37.005 3.922 37.03 4.449 ;
      RECT 37 3.175 37.005 4.441 ;
      RECT 36.985 3.175 37 4.428 ;
      RECT 36.965 3.175 36.985 4.385 ;
      RECT 36.955 3.175 36.965 4.335 ;
      RECT 36.95 3.175 36.955 4.308 ;
      RECT 36.945 3.175 36.95 4.286 ;
      RECT 36.94 3.401 36.945 4.269 ;
      RECT 36.935 3.423 36.94 4.247 ;
      RECT 36.93 3.465 36.935 4.23 ;
      RECT 36.9 3.515 36.93 4.174 ;
      RECT 36.895 3.542 36.9 4.116 ;
      RECT 36.88 3.56 36.895 4.08 ;
      RECT 36.875 3.578 36.88 4.044 ;
      RECT 36.869 3.585 36.875 4.025 ;
      RECT 36.865 3.592 36.869 4.008 ;
      RECT 36.86 3.597 36.865 3.977 ;
      RECT 36.85 3.6 36.86 3.952 ;
      RECT 36.84 3.6 36.85 3.918 ;
      RECT 36.835 3.6 36.84 3.895 ;
      RECT 36.83 3.6 36.835 3.875 ;
      RECT 35.45 4.765 35.71 5.025 ;
      RECT 35.47 4.692 35.65 5.025 ;
      RECT 35.47 4.435 35.645 5.025 ;
      RECT 35.47 4.227 35.635 5.025 ;
      RECT 35.475 4.145 35.635 5.025 ;
      RECT 35.475 3.91 35.625 5.025 ;
      RECT 35.475 3.757 35.62 5.025 ;
      RECT 35.48 3.742 35.62 5.025 ;
      RECT 35.53 3.457 35.62 5.025 ;
      RECT 35.485 3.692 35.62 5.025 ;
      RECT 35.515 3.51 35.62 5.025 ;
      RECT 35.5 3.622 35.62 5.025 ;
      RECT 35.505 3.58 35.62 5.025 ;
      RECT 35.5 3.622 35.635 3.685 ;
      RECT 35.535 3.21 35.64 3.63 ;
      RECT 35.535 3.21 35.655 3.613 ;
      RECT 35.535 3.21 35.69 3.575 ;
      RECT 35.53 3.457 35.74 3.508 ;
      RECT 35.535 3.21 35.795 3.47 ;
      RECT 34.795 3.915 35.055 4.175 ;
      RECT 34.795 3.915 35.065 4.133 ;
      RECT 34.795 3.915 35.151 4.104 ;
      RECT 34.795 3.915 35.22 4.056 ;
      RECT 34.795 3.915 35.255 4.025 ;
      RECT 35.025 3.735 35.305 4.015 ;
      RECT 34.86 3.9 35.305 4.015 ;
      RECT 34.95 3.777 35.055 4.175 ;
      RECT 34.88 3.84 35.305 4.015 ;
      RECT 29.33 8.51 29.65 8.835 ;
      RECT 29.36 7.985 29.53 8.835 ;
      RECT 29.36 7.985 29.535 8.335 ;
      RECT 29.36 7.985 30.335 8.16 ;
      RECT 30.16 3.26 30.335 8.16 ;
      RECT 30.105 3.26 30.455 3.61 ;
      RECT 30.13 8.945 30.455 9.27 ;
      RECT 29.015 9.035 30.455 9.205 ;
      RECT 29.015 3.69 29.175 9.205 ;
      RECT 29.33 3.66 29.65 3.98 ;
      RECT 29.015 3.69 29.65 3.86 ;
      RECT 27.68 4 28.065 4.35 ;
      RECT 27.67 4.065 28.065 4.265 ;
      RECT 27.815 3.995 27.985 4.35 ;
      RECT 26.125 3.735 26.405 4.015 ;
      RECT 26.12 3.735 26.405 3.968 ;
      RECT 26.1 3.735 26.405 3.945 ;
      RECT 26.09 3.735 26.405 3.925 ;
      RECT 26.08 3.735 26.405 3.91 ;
      RECT 26.055 3.735 26.405 3.883 ;
      RECT 26.045 3.735 26.405 3.858 ;
      RECT 26 3.59 26.28 3.85 ;
      RECT 26 3.685 26.38 3.85 ;
      RECT 26 3.63 26.325 3.85 ;
      RECT 26 3.622 26.32 3.85 ;
      RECT 26 3.612 26.315 3.85 ;
      RECT 26 3.6 26.31 3.85 ;
      RECT 24.925 4.295 25.205 4.575 ;
      RECT 24.925 4.295 25.24 4.555 ;
      RECT 16.545 9.285 16.835 9.635 ;
      RECT 16.545 9.36 17.91 9.53 ;
      RECT 17.74 8.975 17.91 9.53 ;
      RECT 24.67 8.895 25.02 9.245 ;
      RECT 17.74 8.975 25.02 9.145 ;
      RECT 24.96 3.715 25.01 3.975 ;
      RECT 24.75 3.715 24.755 3.975 ;
      RECT 23.945 3.27 23.975 3.53 ;
      RECT 23.715 3.27 23.79 3.53 ;
      RECT 24.935 3.665 24.96 3.975 ;
      RECT 24.93 3.622 24.935 3.975 ;
      RECT 24.925 3.605 24.93 3.975 ;
      RECT 24.92 3.592 24.925 3.975 ;
      RECT 24.845 3.475 24.92 3.975 ;
      RECT 24.8 3.292 24.845 3.975 ;
      RECT 24.795 3.22 24.8 3.975 ;
      RECT 24.78 3.195 24.795 3.975 ;
      RECT 24.755 3.157 24.78 3.975 ;
      RECT 24.745 3.137 24.755 3.697 ;
      RECT 24.73 3.129 24.745 3.652 ;
      RECT 24.725 3.121 24.73 3.623 ;
      RECT 24.72 3.118 24.725 3.603 ;
      RECT 24.715 3.115 24.72 3.583 ;
      RECT 24.71 3.112 24.715 3.563 ;
      RECT 24.68 3.101 24.71 3.5 ;
      RECT 24.66 3.086 24.68 3.415 ;
      RECT 24.655 3.078 24.66 3.378 ;
      RECT 24.645 3.072 24.655 3.345 ;
      RECT 24.63 3.064 24.645 3.305 ;
      RECT 24.625 3.057 24.63 3.265 ;
      RECT 24.62 3.054 24.625 3.243 ;
      RECT 24.615 3.051 24.62 3.23 ;
      RECT 24.61 3.05 24.615 3.22 ;
      RECT 24.595 3.044 24.61 3.21 ;
      RECT 24.57 3.031 24.595 3.195 ;
      RECT 24.52 3.006 24.57 3.166 ;
      RECT 24.505 2.985 24.52 3.141 ;
      RECT 24.495 2.978 24.505 3.13 ;
      RECT 24.44 2.959 24.495 3.103 ;
      RECT 24.415 2.937 24.44 3.076 ;
      RECT 24.41 2.93 24.415 3.071 ;
      RECT 24.395 2.93 24.41 3.069 ;
      RECT 24.37 2.922 24.395 3.065 ;
      RECT 24.355 2.92 24.37 3.061 ;
      RECT 24.325 2.92 24.355 3.058 ;
      RECT 24.315 2.92 24.325 3.053 ;
      RECT 24.27 2.92 24.315 3.051 ;
      RECT 24.241 2.92 24.27 3.052 ;
      RECT 24.155 2.92 24.241 3.054 ;
      RECT 24.141 2.921 24.155 3.056 ;
      RECT 24.055 2.922 24.141 3.058 ;
      RECT 24.04 2.923 24.055 3.068 ;
      RECT 24.035 2.924 24.04 3.077 ;
      RECT 24.015 2.927 24.035 3.087 ;
      RECT 24 2.935 24.015 3.102 ;
      RECT 23.98 2.953 24 3.117 ;
      RECT 23.97 2.965 23.98 3.14 ;
      RECT 23.96 2.974 23.97 3.17 ;
      RECT 23.945 2.986 23.96 3.215 ;
      RECT 23.89 3.019 23.945 3.53 ;
      RECT 23.885 3.047 23.89 3.53 ;
      RECT 23.865 3.062 23.885 3.53 ;
      RECT 23.83 3.122 23.865 3.53 ;
      RECT 23.828 3.172 23.83 3.53 ;
      RECT 23.825 3.18 23.828 3.53 ;
      RECT 23.815 3.195 23.825 3.53 ;
      RECT 23.81 3.207 23.815 3.53 ;
      RECT 23.8 3.232 23.81 3.53 ;
      RECT 23.79 3.26 23.8 3.53 ;
      RECT 21.695 4.765 21.745 5.025 ;
      RECT 24.605 4.315 24.665 4.575 ;
      RECT 24.59 4.315 24.605 4.585 ;
      RECT 24.571 4.315 24.59 4.618 ;
      RECT 24.485 4.315 24.571 4.743 ;
      RECT 24.405 4.315 24.485 4.925 ;
      RECT 24.4 4.552 24.405 5.01 ;
      RECT 24.375 4.622 24.4 5.038 ;
      RECT 24.37 4.692 24.375 5.065 ;
      RECT 24.35 4.764 24.37 5.087 ;
      RECT 24.345 4.831 24.35 5.11 ;
      RECT 24.335 4.86 24.345 5.125 ;
      RECT 24.325 4.882 24.335 5.142 ;
      RECT 24.32 4.892 24.325 5.153 ;
      RECT 24.315 4.9 24.32 5.161 ;
      RECT 24.305 4.908 24.315 5.173 ;
      RECT 24.3 4.92 24.305 5.183 ;
      RECT 24.295 4.928 24.3 5.188 ;
      RECT 24.275 4.946 24.295 5.198 ;
      RECT 24.27 4.963 24.275 5.205 ;
      RECT 24.265 4.971 24.27 5.206 ;
      RECT 24.26 4.982 24.265 5.208 ;
      RECT 24.22 5.02 24.26 5.218 ;
      RECT 24.215 5.055 24.22 5.229 ;
      RECT 24.21 5.06 24.215 5.232 ;
      RECT 24.185 5.07 24.21 5.239 ;
      RECT 24.175 5.084 24.185 5.248 ;
      RECT 24.155 5.096 24.175 5.251 ;
      RECT 24.105 5.115 24.155 5.255 ;
      RECT 24.06 5.13 24.105 5.26 ;
      RECT 23.995 5.133 24.06 5.266 ;
      RECT 23.98 5.131 23.995 5.273 ;
      RECT 23.95 5.13 23.98 5.273 ;
      RECT 23.911 5.129 23.95 5.269 ;
      RECT 23.825 5.126 23.911 5.265 ;
      RECT 23.808 5.124 23.825 5.262 ;
      RECT 23.722 5.122 23.808 5.259 ;
      RECT 23.636 5.119 23.722 5.253 ;
      RECT 23.55 5.115 23.636 5.248 ;
      RECT 23.472 5.112 23.55 5.244 ;
      RECT 23.386 5.109 23.472 5.242 ;
      RECT 23.3 5.106 23.386 5.239 ;
      RECT 23.242 5.104 23.3 5.236 ;
      RECT 23.156 5.101 23.242 5.234 ;
      RECT 23.07 5.097 23.156 5.232 ;
      RECT 22.984 5.094 23.07 5.229 ;
      RECT 22.898 5.09 22.984 5.227 ;
      RECT 22.812 5.086 22.898 5.224 ;
      RECT 22.726 5.083 22.812 5.222 ;
      RECT 22.64 5.079 22.726 5.219 ;
      RECT 22.554 5.076 22.64 5.217 ;
      RECT 22.468 5.072 22.554 5.214 ;
      RECT 22.382 5.069 22.468 5.212 ;
      RECT 22.296 5.065 22.382 5.209 ;
      RECT 22.21 5.062 22.296 5.207 ;
      RECT 22.2 5.06 22.21 5.203 ;
      RECT 22.195 5.06 22.2 5.201 ;
      RECT 22.155 5.055 22.195 5.195 ;
      RECT 22.141 5.046 22.155 5.188 ;
      RECT 22.055 5.016 22.141 5.173 ;
      RECT 22.035 4.982 22.055 5.158 ;
      RECT 21.965 4.951 22.035 5.145 ;
      RECT 21.96 4.926 21.965 5.134 ;
      RECT 21.955 4.92 21.96 5.132 ;
      RECT 21.886 4.765 21.955 5.12 ;
      RECT 21.8 4.765 21.886 5.094 ;
      RECT 21.775 4.765 21.8 5.073 ;
      RECT 21.77 4.765 21.775 5.063 ;
      RECT 21.765 4.765 21.77 5.055 ;
      RECT 21.745 4.765 21.765 5.038 ;
      RECT 24.165 3.335 24.425 3.595 ;
      RECT 24.15 3.335 24.425 3.498 ;
      RECT 24.12 3.335 24.425 3.473 ;
      RECT 24.085 3.175 24.365 3.455 ;
      RECT 24.055 4.665 24.115 4.925 ;
      RECT 23.08 3.355 23.135 3.615 ;
      RECT 24.015 4.622 24.055 4.925 ;
      RECT 23.986 4.543 24.015 4.925 ;
      RECT 23.9 4.415 23.986 4.925 ;
      RECT 23.88 4.295 23.9 4.925 ;
      RECT 23.855 4.246 23.88 4.925 ;
      RECT 23.85 4.211 23.855 4.775 ;
      RECT 23.82 4.171 23.85 4.713 ;
      RECT 23.795 4.108 23.82 4.628 ;
      RECT 23.785 4.07 23.795 4.565 ;
      RECT 23.77 4.045 23.785 4.526 ;
      RECT 23.727 4.003 23.77 4.432 ;
      RECT 23.725 3.976 23.727 4.359 ;
      RECT 23.72 3.971 23.725 4.35 ;
      RECT 23.715 3.964 23.72 4.325 ;
      RECT 23.71 3.958 23.715 4.31 ;
      RECT 23.705 3.952 23.71 4.298 ;
      RECT 23.695 3.943 23.705 4.28 ;
      RECT 23.69 3.934 23.695 4.258 ;
      RECT 23.665 3.915 23.69 4.208 ;
      RECT 23.66 3.896 23.665 4.158 ;
      RECT 23.645 3.882 23.66 4.118 ;
      RECT 23.64 3.868 23.645 4.085 ;
      RECT 23.635 3.861 23.64 4.078 ;
      RECT 23.62 3.848 23.635 4.07 ;
      RECT 23.575 3.81 23.62 4.043 ;
      RECT 23.545 3.763 23.575 4.008 ;
      RECT 23.525 3.732 23.545 3.985 ;
      RECT 23.445 3.665 23.525 3.938 ;
      RECT 23.415 3.595 23.445 3.885 ;
      RECT 23.41 3.572 23.415 3.868 ;
      RECT 23.38 3.55 23.41 3.853 ;
      RECT 23.35 3.509 23.38 3.825 ;
      RECT 23.345 3.484 23.35 3.81 ;
      RECT 23.34 3.478 23.345 3.803 ;
      RECT 23.33 3.355 23.34 3.795 ;
      RECT 23.32 3.355 23.33 3.788 ;
      RECT 23.315 3.355 23.32 3.78 ;
      RECT 23.295 3.355 23.315 3.768 ;
      RECT 23.245 3.355 23.295 3.738 ;
      RECT 23.19 3.355 23.245 3.688 ;
      RECT 23.16 3.355 23.19 3.648 ;
      RECT 23.135 3.355 23.16 3.625 ;
      RECT 23.005 4.08 23.285 4.36 ;
      RECT 22.97 3.995 23.23 4.255 ;
      RECT 22.97 4.077 23.24 4.255 ;
      RECT 21.17 3.45 21.175 3.935 ;
      RECT 21.06 3.635 21.065 3.935 ;
      RECT 20.97 3.675 21.035 3.935 ;
      RECT 22.645 3.175 22.735 3.805 ;
      RECT 22.61 3.225 22.615 3.805 ;
      RECT 22.555 3.25 22.565 3.805 ;
      RECT 22.51 3.25 22.52 3.805 ;
      RECT 22.88 3.175 22.925 3.455 ;
      RECT 21.73 2.905 21.93 3.045 ;
      RECT 22.846 3.175 22.88 3.467 ;
      RECT 22.76 3.175 22.846 3.507 ;
      RECT 22.745 3.175 22.76 3.548 ;
      RECT 22.74 3.175 22.745 3.568 ;
      RECT 22.735 3.175 22.74 3.588 ;
      RECT 22.615 3.217 22.645 3.805 ;
      RECT 22.565 3.237 22.61 3.805 ;
      RECT 22.55 3.252 22.555 3.805 ;
      RECT 22.52 3.252 22.55 3.805 ;
      RECT 22.475 3.237 22.51 3.805 ;
      RECT 22.47 3.225 22.475 3.585 ;
      RECT 22.465 3.222 22.47 3.565 ;
      RECT 22.45 3.212 22.465 3.518 ;
      RECT 22.445 3.205 22.45 3.481 ;
      RECT 22.44 3.202 22.445 3.464 ;
      RECT 22.425 3.192 22.44 3.42 ;
      RECT 22.42 3.183 22.425 3.38 ;
      RECT 22.415 3.179 22.42 3.365 ;
      RECT 22.405 3.173 22.415 3.348 ;
      RECT 22.365 3.154 22.405 3.323 ;
      RECT 22.36 3.136 22.365 3.303 ;
      RECT 22.35 3.13 22.36 3.298 ;
      RECT 22.32 3.114 22.35 3.285 ;
      RECT 22.305 3.096 22.32 3.268 ;
      RECT 22.29 3.084 22.305 3.255 ;
      RECT 22.285 3.076 22.29 3.248 ;
      RECT 22.255 3.062 22.285 3.235 ;
      RECT 22.25 3.047 22.255 3.223 ;
      RECT 22.24 3.041 22.25 3.215 ;
      RECT 22.22 3.029 22.24 3.203 ;
      RECT 22.21 3.017 22.22 3.19 ;
      RECT 22.18 3.001 22.21 3.175 ;
      RECT 22.16 2.981 22.18 3.158 ;
      RECT 22.155 2.971 22.16 3.148 ;
      RECT 22.13 2.959 22.155 3.135 ;
      RECT 22.125 2.947 22.13 3.123 ;
      RECT 22.12 2.942 22.125 3.119 ;
      RECT 22.105 2.935 22.12 3.111 ;
      RECT 22.095 2.922 22.105 3.101 ;
      RECT 22.09 2.92 22.095 3.095 ;
      RECT 22.065 2.913 22.09 3.084 ;
      RECT 22.06 2.906 22.065 3.073 ;
      RECT 22.035 2.905 22.06 3.06 ;
      RECT 22.016 2.905 22.035 3.05 ;
      RECT 21.93 2.905 22.016 3.047 ;
      RECT 21.7 2.905 21.73 3.05 ;
      RECT 21.66 2.912 21.7 3.063 ;
      RECT 21.635 2.922 21.66 3.076 ;
      RECT 21.62 2.931 21.635 3.086 ;
      RECT 21.59 2.936 21.62 3.105 ;
      RECT 21.585 2.942 21.59 3.123 ;
      RECT 21.565 2.952 21.585 3.138 ;
      RECT 21.555 2.965 21.565 3.158 ;
      RECT 21.54 2.977 21.555 3.175 ;
      RECT 21.535 2.987 21.54 3.185 ;
      RECT 21.53 2.992 21.535 3.19 ;
      RECT 21.52 3 21.53 3.203 ;
      RECT 21.47 3.032 21.52 3.24 ;
      RECT 21.455 3.067 21.47 3.281 ;
      RECT 21.45 3.077 21.455 3.296 ;
      RECT 21.445 3.082 21.45 3.303 ;
      RECT 21.42 3.098 21.445 3.323 ;
      RECT 21.405 3.119 21.42 3.348 ;
      RECT 21.38 3.14 21.405 3.373 ;
      RECT 21.37 3.159 21.38 3.396 ;
      RECT 21.345 3.177 21.37 3.419 ;
      RECT 21.33 3.197 21.345 3.443 ;
      RECT 21.325 3.207 21.33 3.455 ;
      RECT 21.31 3.219 21.325 3.475 ;
      RECT 21.3 3.234 21.31 3.515 ;
      RECT 21.295 3.242 21.3 3.543 ;
      RECT 21.285 3.252 21.295 3.563 ;
      RECT 21.28 3.265 21.285 3.588 ;
      RECT 21.275 3.278 21.28 3.608 ;
      RECT 21.27 3.284 21.275 3.63 ;
      RECT 21.26 3.293 21.27 3.65 ;
      RECT 21.255 3.313 21.26 3.673 ;
      RECT 21.25 3.319 21.255 3.693 ;
      RECT 21.245 3.326 21.25 3.715 ;
      RECT 21.24 3.337 21.245 3.728 ;
      RECT 21.23 3.347 21.24 3.753 ;
      RECT 21.21 3.372 21.23 3.935 ;
      RECT 21.18 3.412 21.21 3.935 ;
      RECT 21.175 3.442 21.18 3.935 ;
      RECT 21.15 3.47 21.17 3.935 ;
      RECT 21.12 3.515 21.15 3.935 ;
      RECT 21.115 3.542 21.12 3.935 ;
      RECT 21.095 3.56 21.115 3.935 ;
      RECT 21.085 3.585 21.095 3.935 ;
      RECT 21.08 3.597 21.085 3.935 ;
      RECT 21.065 3.62 21.08 3.935 ;
      RECT 21.045 3.647 21.06 3.935 ;
      RECT 21.035 3.67 21.045 3.935 ;
      RECT 22.825 4.555 22.905 4.815 ;
      RECT 22.06 3.775 22.13 4.035 ;
      RECT 22.791 4.522 22.825 4.815 ;
      RECT 22.705 4.425 22.791 4.815 ;
      RECT 22.685 4.337 22.705 4.815 ;
      RECT 22.675 4.307 22.685 4.815 ;
      RECT 22.665 4.287 22.675 4.815 ;
      RECT 22.645 4.274 22.665 4.815 ;
      RECT 22.63 4.264 22.645 4.643 ;
      RECT 22.625 4.257 22.63 4.598 ;
      RECT 22.615 4.251 22.625 4.588 ;
      RECT 22.605 4.243 22.615 4.57 ;
      RECT 22.6 4.237 22.605 4.558 ;
      RECT 22.59 4.232 22.6 4.545 ;
      RECT 22.57 4.222 22.59 4.518 ;
      RECT 22.53 4.201 22.57 4.47 ;
      RECT 22.515 4.182 22.53 4.428 ;
      RECT 22.49 4.168 22.515 4.398 ;
      RECT 22.48 4.156 22.49 4.365 ;
      RECT 22.475 4.151 22.48 4.355 ;
      RECT 22.445 4.137 22.475 4.335 ;
      RECT 22.435 4.121 22.445 4.308 ;
      RECT 22.43 4.116 22.435 4.298 ;
      RECT 22.405 4.107 22.43 4.278 ;
      RECT 22.395 4.095 22.405 4.258 ;
      RECT 22.325 4.063 22.395 4.233 ;
      RECT 22.32 4.032 22.325 4.21 ;
      RECT 22.271 3.775 22.32 4.193 ;
      RECT 22.185 3.775 22.271 4.152 ;
      RECT 22.13 3.775 22.185 4.08 ;
      RECT 22.22 4.56 22.38 4.82 ;
      RECT 21.745 3.175 21.795 3.86 ;
      RECT 21.535 3.6 21.57 3.86 ;
      RECT 21.85 3.175 21.855 3.635 ;
      RECT 21.94 3.175 21.965 3.455 ;
      RECT 22.215 4.557 22.22 4.82 ;
      RECT 22.18 4.545 22.215 4.82 ;
      RECT 22.12 4.518 22.18 4.82 ;
      RECT 22.115 4.501 22.12 4.674 ;
      RECT 22.11 4.498 22.115 4.661 ;
      RECT 22.09 4.491 22.11 4.648 ;
      RECT 22.055 4.474 22.09 4.63 ;
      RECT 22.015 4.453 22.055 4.61 ;
      RECT 22.01 4.441 22.015 4.598 ;
      RECT 21.97 4.427 22.01 4.584 ;
      RECT 21.95 4.41 21.97 4.566 ;
      RECT 21.94 4.402 21.95 4.558 ;
      RECT 21.925 3.175 21.94 3.473 ;
      RECT 21.91 4.392 21.94 4.545 ;
      RECT 21.895 3.175 21.925 3.518 ;
      RECT 21.9 4.382 21.91 4.532 ;
      RECT 21.87 4.367 21.9 4.519 ;
      RECT 21.855 3.175 21.895 3.585 ;
      RECT 21.855 4.335 21.87 4.505 ;
      RECT 21.85 4.307 21.855 4.499 ;
      RECT 21.845 3.175 21.85 3.64 ;
      RECT 21.835 4.277 21.85 4.493 ;
      RECT 21.84 3.175 21.845 3.653 ;
      RECT 21.83 3.175 21.84 3.673 ;
      RECT 21.795 4.19 21.835 4.478 ;
      RECT 21.795 3.175 21.83 3.713 ;
      RECT 21.79 4.122 21.795 4.466 ;
      RECT 21.775 4.077 21.79 4.461 ;
      RECT 21.77 4.015 21.775 4.456 ;
      RECT 21.745 3.922 21.77 4.449 ;
      RECT 21.74 3.175 21.745 4.441 ;
      RECT 21.725 3.175 21.74 4.428 ;
      RECT 21.705 3.175 21.725 4.385 ;
      RECT 21.695 3.175 21.705 4.335 ;
      RECT 21.69 3.175 21.695 4.308 ;
      RECT 21.685 3.175 21.69 4.286 ;
      RECT 21.68 3.401 21.685 4.269 ;
      RECT 21.675 3.423 21.68 4.247 ;
      RECT 21.67 3.465 21.675 4.23 ;
      RECT 21.64 3.515 21.67 4.174 ;
      RECT 21.635 3.542 21.64 4.116 ;
      RECT 21.62 3.56 21.635 4.08 ;
      RECT 21.615 3.578 21.62 4.044 ;
      RECT 21.609 3.585 21.615 4.025 ;
      RECT 21.605 3.592 21.609 4.008 ;
      RECT 21.6 3.597 21.605 3.977 ;
      RECT 21.59 3.6 21.6 3.952 ;
      RECT 21.58 3.6 21.59 3.918 ;
      RECT 21.575 3.6 21.58 3.895 ;
      RECT 21.57 3.6 21.575 3.875 ;
      RECT 20.19 4.765 20.45 5.025 ;
      RECT 20.21 4.692 20.39 5.025 ;
      RECT 20.21 4.435 20.385 5.025 ;
      RECT 20.21 4.227 20.375 5.025 ;
      RECT 20.215 4.145 20.375 5.025 ;
      RECT 20.215 3.91 20.365 5.025 ;
      RECT 20.215 3.757 20.36 5.025 ;
      RECT 20.22 3.742 20.36 5.025 ;
      RECT 20.27 3.457 20.36 5.025 ;
      RECT 20.225 3.692 20.36 5.025 ;
      RECT 20.255 3.51 20.36 5.025 ;
      RECT 20.24 3.622 20.36 5.025 ;
      RECT 20.245 3.58 20.36 5.025 ;
      RECT 20.24 3.622 20.375 3.685 ;
      RECT 20.275 3.21 20.38 3.63 ;
      RECT 20.275 3.21 20.395 3.613 ;
      RECT 20.275 3.21 20.43 3.575 ;
      RECT 20.27 3.457 20.48 3.508 ;
      RECT 20.275 3.21 20.535 3.47 ;
      RECT 19.535 3.915 19.795 4.175 ;
      RECT 19.535 3.915 19.805 4.133 ;
      RECT 19.535 3.915 19.891 4.104 ;
      RECT 19.535 3.915 19.96 4.056 ;
      RECT 19.535 3.915 19.995 4.025 ;
      RECT 19.765 3.735 20.045 4.015 ;
      RECT 19.6 3.9 20.045 4.015 ;
      RECT 19.69 3.777 19.795 4.175 ;
      RECT 19.62 3.84 20.045 4.015 ;
      RECT 93.455 7.205 93.835 7.585 ;
      RECT 85.04 9.345 85.41 9.715 ;
      RECT 78.195 7.205 78.575 7.585 ;
      RECT 69.78 9.345 70.15 9.715 ;
      RECT 62.935 7.205 63.315 7.585 ;
      RECT 54.52 9.345 54.89 9.715 ;
      RECT 47.675 7.205 48.055 7.585 ;
      RECT 39.26 9.345 39.63 9.715 ;
      RECT 32.415 7.205 32.795 7.585 ;
      RECT 24 9.345 24.37 9.715 ;
    LAYER via1 ;
      RECT 93.63 9.665 93.78 9.815 ;
      RECT 93.57 7.32 93.72 7.47 ;
      RECT 91.26 9.03 91.41 9.18 ;
      RECT 91.245 3.36 91.395 3.51 ;
      RECT 90.455 3.745 90.605 3.895 ;
      RECT 90.455 8.615 90.605 8.765 ;
      RECT 88.865 4.1 89.015 4.25 ;
      RECT 87.095 3.645 87.245 3.795 ;
      RECT 86.075 4.35 86.225 4.5 ;
      RECT 85.845 3.77 85.995 3.92 ;
      RECT 85.81 9.005 85.96 9.155 ;
      RECT 85.5 4.37 85.65 4.52 ;
      RECT 85.26 3.39 85.41 3.54 ;
      RECT 85.15 9.455 85.3 9.605 ;
      RECT 84.95 4.72 85.1 4.87 ;
      RECT 84.81 3.325 84.96 3.475 ;
      RECT 84.175 3.41 84.325 3.56 ;
      RECT 84.065 4.05 84.215 4.2 ;
      RECT 83.74 4.61 83.89 4.76 ;
      RECT 83.57 3.6 83.72 3.75 ;
      RECT 83.215 4.615 83.365 4.765 ;
      RECT 83.155 3.83 83.305 3.98 ;
      RECT 82.79 4.82 82.94 4.97 ;
      RECT 82.63 3.655 82.78 3.805 ;
      RECT 82.065 3.73 82.215 3.88 ;
      RECT 81.37 3.265 81.52 3.415 ;
      RECT 81.285 4.82 81.435 4.97 ;
      RECT 80.63 3.97 80.78 4.12 ;
      RECT 78.345 9.05 78.495 9.2 ;
      RECT 78.31 7.32 78.46 7.47 ;
      RECT 76 9.03 76.15 9.18 ;
      RECT 75.985 3.36 76.135 3.51 ;
      RECT 75.195 3.745 75.345 3.895 ;
      RECT 75.195 8.615 75.345 8.765 ;
      RECT 73.605 4.1 73.755 4.25 ;
      RECT 71.835 3.645 71.985 3.795 ;
      RECT 70.815 4.35 70.965 4.5 ;
      RECT 70.585 3.77 70.735 3.92 ;
      RECT 70.55 9.005 70.7 9.155 ;
      RECT 70.24 4.37 70.39 4.52 ;
      RECT 70 3.39 70.15 3.54 ;
      RECT 69.89 9.455 70.04 9.605 ;
      RECT 69.69 4.72 69.84 4.87 ;
      RECT 69.55 3.325 69.7 3.475 ;
      RECT 68.915 3.41 69.065 3.56 ;
      RECT 68.805 4.05 68.955 4.2 ;
      RECT 68.48 4.61 68.63 4.76 ;
      RECT 68.31 3.6 68.46 3.75 ;
      RECT 67.955 4.615 68.105 4.765 ;
      RECT 67.895 3.83 68.045 3.98 ;
      RECT 67.53 4.82 67.68 4.97 ;
      RECT 67.37 3.655 67.52 3.805 ;
      RECT 66.805 3.73 66.955 3.88 ;
      RECT 66.11 3.265 66.26 3.415 ;
      RECT 66.025 4.82 66.175 4.97 ;
      RECT 65.37 3.97 65.52 4.12 ;
      RECT 63.085 9.05 63.235 9.2 ;
      RECT 63.05 7.32 63.2 7.47 ;
      RECT 60.74 9.03 60.89 9.18 ;
      RECT 60.725 3.36 60.875 3.51 ;
      RECT 59.935 3.745 60.085 3.895 ;
      RECT 59.935 8.615 60.085 8.765 ;
      RECT 58.345 4.1 58.495 4.25 ;
      RECT 56.575 3.645 56.725 3.795 ;
      RECT 55.555 4.35 55.705 4.5 ;
      RECT 55.325 3.77 55.475 3.92 ;
      RECT 55.29 9.005 55.44 9.155 ;
      RECT 54.98 4.37 55.13 4.52 ;
      RECT 54.74 3.39 54.89 3.54 ;
      RECT 54.63 9.455 54.78 9.605 ;
      RECT 54.43 4.72 54.58 4.87 ;
      RECT 54.29 3.325 54.44 3.475 ;
      RECT 53.655 3.41 53.805 3.56 ;
      RECT 53.545 4.05 53.695 4.2 ;
      RECT 53.22 4.61 53.37 4.76 ;
      RECT 53.05 3.6 53.2 3.75 ;
      RECT 52.695 4.615 52.845 4.765 ;
      RECT 52.635 3.83 52.785 3.98 ;
      RECT 52.27 4.82 52.42 4.97 ;
      RECT 52.11 3.655 52.26 3.805 ;
      RECT 51.545 3.73 51.695 3.88 ;
      RECT 50.85 3.265 51 3.415 ;
      RECT 50.765 4.82 50.915 4.97 ;
      RECT 50.11 3.97 50.26 4.12 ;
      RECT 47.87 9.05 48.02 9.2 ;
      RECT 47.79 7.32 47.94 7.47 ;
      RECT 45.48 9.03 45.63 9.18 ;
      RECT 45.465 3.36 45.615 3.51 ;
      RECT 44.675 3.745 44.825 3.895 ;
      RECT 44.675 8.615 44.825 8.765 ;
      RECT 43.085 4.1 43.235 4.25 ;
      RECT 41.315 3.645 41.465 3.795 ;
      RECT 40.295 4.35 40.445 4.5 ;
      RECT 40.065 3.77 40.215 3.92 ;
      RECT 40.03 9.005 40.18 9.155 ;
      RECT 39.72 4.37 39.87 4.52 ;
      RECT 39.48 3.39 39.63 3.54 ;
      RECT 39.37 9.455 39.52 9.605 ;
      RECT 39.17 4.72 39.32 4.87 ;
      RECT 39.03 3.325 39.18 3.475 ;
      RECT 38.395 3.41 38.545 3.56 ;
      RECT 38.285 4.05 38.435 4.2 ;
      RECT 37.96 4.61 38.11 4.76 ;
      RECT 37.79 3.6 37.94 3.75 ;
      RECT 37.435 4.615 37.585 4.765 ;
      RECT 37.375 3.83 37.525 3.98 ;
      RECT 37.01 4.82 37.16 4.97 ;
      RECT 36.85 3.655 37 3.805 ;
      RECT 36.285 3.73 36.435 3.88 ;
      RECT 35.59 3.265 35.74 3.415 ;
      RECT 35.505 4.82 35.655 4.97 ;
      RECT 34.85 3.97 35 4.12 ;
      RECT 32.61 9.05 32.76 9.2 ;
      RECT 32.53 7.32 32.68 7.47 ;
      RECT 30.22 9.03 30.37 9.18 ;
      RECT 30.205 3.36 30.355 3.51 ;
      RECT 29.415 3.745 29.565 3.895 ;
      RECT 29.415 8.615 29.565 8.765 ;
      RECT 27.825 4.1 27.975 4.25 ;
      RECT 26.055 3.645 26.205 3.795 ;
      RECT 25.035 4.35 25.185 4.5 ;
      RECT 24.805 3.77 24.955 3.92 ;
      RECT 24.77 8.995 24.92 9.145 ;
      RECT 24.46 4.37 24.61 4.52 ;
      RECT 24.22 3.39 24.37 3.54 ;
      RECT 24.11 9.455 24.26 9.605 ;
      RECT 23.91 4.72 24.06 4.87 ;
      RECT 23.77 3.325 23.92 3.475 ;
      RECT 23.135 3.41 23.285 3.56 ;
      RECT 23.025 4.05 23.175 4.2 ;
      RECT 22.7 4.61 22.85 4.76 ;
      RECT 22.53 3.6 22.68 3.75 ;
      RECT 22.175 4.615 22.325 4.765 ;
      RECT 22.115 3.83 22.265 3.98 ;
      RECT 21.75 4.82 21.9 4.97 ;
      RECT 21.59 3.655 21.74 3.805 ;
      RECT 21.025 3.73 21.175 3.88 ;
      RECT 20.33 3.265 20.48 3.415 ;
      RECT 20.245 4.82 20.395 4.97 ;
      RECT 19.59 3.97 19.74 4.12 ;
      RECT 16.615 9.385 16.765 9.535 ;
      RECT 16.24 8.645 16.39 8.795 ;
    LAYER met1 ;
      RECT 93.495 10.06 93.79 10.29 ;
      RECT 93.555 9.565 93.73 10.29 ;
      RECT 93.53 9.565 93.88 9.915 ;
      RECT 93.555 8.58 93.725 10.29 ;
      RECT 93.495 8.58 93.785 8.81 ;
      RECT 92.505 10.06 92.8 10.29 ;
      RECT 92.565 8.58 92.735 10.29 ;
      RECT 92.505 8.58 92.795 8.81 ;
      RECT 92.505 8.615 93.355 8.775 ;
      RECT 93.19 8.21 93.355 8.775 ;
      RECT 92.505 8.61 92.9 8.775 ;
      RECT 93.125 8.21 93.415 8.44 ;
      RECT 93.125 8.24 93.585 8.41 ;
      RECT 93.09 4.005 93.41 4.26 ;
      RECT 93.09 4.055 93.58 4.225 ;
      RECT 93.09 3.69 93.28 4.26 ;
      RECT 92.505 3.655 92.795 3.885 ;
      RECT 92.505 3.69 93.28 3.86 ;
      RECT 92.565 2.175 92.735 3.885 ;
      RECT 92.505 2.175 92.8 2.405 ;
      RECT 92.135 4.025 92.425 4.255 ;
      RECT 92.135 4.055 92.595 4.225 ;
      RECT 92.2 2.95 92.365 4.255 ;
      RECT 90.715 2.915 91.005 3.145 ;
      RECT 90.715 2.95 92.365 3.12 ;
      RECT 90.775 2.175 90.945 3.145 ;
      RECT 90.715 2.175 91.005 2.405 ;
      RECT 90.715 10.06 91.005 10.29 ;
      RECT 90.775 9.32 90.945 10.29 ;
      RECT 90.775 9.41 92.365 9.58 ;
      RECT 92.195 8.21 92.365 9.58 ;
      RECT 90.715 9.32 91.005 9.55 ;
      RECT 92.135 8.21 92.425 8.44 ;
      RECT 92.135 8.24 92.595 8.41 ;
      RECT 88.765 4 89.105 4.35 ;
      RECT 88.855 3.32 89.025 4.35 ;
      RECT 91.145 3.26 91.495 3.61 ;
      RECT 88.855 3.32 91.495 3.49 ;
      RECT 90.975 3.315 91.495 3.49 ;
      RECT 91.17 8.945 91.495 9.27 ;
      RECT 85.71 8.905 86.06 9.255 ;
      RECT 91.145 8.95 91.495 9.18 ;
      RECT 85.51 8.95 86.06 9.18 ;
      RECT 90.975 8.975 91.495 9.15 ;
      RECT 85.34 8.98 86.06 9.15 ;
      RECT 85.39 8.975 91.495 9.145 ;
      RECT 90.37 3.66 90.69 3.98 ;
      RECT 90.345 3.655 90.635 3.885 ;
      RECT 90.34 3.685 90.69 3.86 ;
      RECT 90.17 3.685 90.69 3.855 ;
      RECT 90.37 8.545 90.69 8.835 ;
      RECT 90.345 8.58 90.69 8.81 ;
      RECT 90.17 8.61 90.69 8.78 ;
      RECT 86.06 4.28 86.21 4.555 ;
      RECT 86.6 3.36 86.605 3.58 ;
      RECT 87.75 3.56 87.765 3.758 ;
      RECT 87.715 3.552 87.75 3.765 ;
      RECT 87.685 3.545 87.715 3.765 ;
      RECT 87.63 3.51 87.685 3.765 ;
      RECT 87.565 3.447 87.63 3.765 ;
      RECT 87.56 3.412 87.565 3.763 ;
      RECT 87.555 3.407 87.56 3.755 ;
      RECT 87.55 3.402 87.555 3.741 ;
      RECT 87.545 3.399 87.55 3.734 ;
      RECT 87.5 3.389 87.545 3.685 ;
      RECT 87.48 3.376 87.5 3.62 ;
      RECT 87.475 3.371 87.48 3.593 ;
      RECT 87.47 3.37 87.475 3.586 ;
      RECT 87.465 3.369 87.47 3.579 ;
      RECT 87.38 3.354 87.465 3.525 ;
      RECT 87.35 3.335 87.38 3.475 ;
      RECT 87.27 3.318 87.35 3.46 ;
      RECT 87.235 3.305 87.27 3.445 ;
      RECT 87.227 3.305 87.235 3.44 ;
      RECT 87.141 3.306 87.227 3.44 ;
      RECT 87.055 3.308 87.141 3.44 ;
      RECT 87.03 3.309 87.055 3.444 ;
      RECT 86.955 3.315 87.03 3.459 ;
      RECT 86.872 3.327 86.955 3.483 ;
      RECT 86.786 3.34 86.872 3.509 ;
      RECT 86.7 3.353 86.786 3.535 ;
      RECT 86.665 3.362 86.7 3.554 ;
      RECT 86.615 3.362 86.665 3.567 ;
      RECT 86.605 3.36 86.615 3.578 ;
      RECT 86.59 3.357 86.6 3.58 ;
      RECT 86.575 3.349 86.59 3.588 ;
      RECT 86.56 3.341 86.575 3.608 ;
      RECT 86.555 3.336 86.56 3.665 ;
      RECT 86.54 3.331 86.555 3.738 ;
      RECT 86.535 3.326 86.54 3.78 ;
      RECT 86.53 3.324 86.535 3.808 ;
      RECT 86.525 3.322 86.53 3.83 ;
      RECT 86.515 3.318 86.525 3.873 ;
      RECT 86.51 3.315 86.515 3.898 ;
      RECT 86.505 3.313 86.51 3.918 ;
      RECT 86.5 3.311 86.505 3.942 ;
      RECT 86.495 3.307 86.5 3.965 ;
      RECT 86.49 3.303 86.495 3.988 ;
      RECT 86.455 3.293 86.49 4.095 ;
      RECT 86.45 3.283 86.455 4.193 ;
      RECT 86.445 3.281 86.45 4.22 ;
      RECT 86.44 3.28 86.445 4.24 ;
      RECT 86.435 3.272 86.44 4.26 ;
      RECT 86.43 3.267 86.435 4.295 ;
      RECT 86.425 3.265 86.43 4.313 ;
      RECT 86.42 3.265 86.425 4.338 ;
      RECT 86.415 3.265 86.42 4.36 ;
      RECT 86.38 3.265 86.415 4.403 ;
      RECT 86.355 3.265 86.38 4.432 ;
      RECT 86.345 3.265 86.355 3.618 ;
      RECT 86.348 3.675 86.355 4.442 ;
      RECT 86.345 3.732 86.348 4.445 ;
      RECT 86.34 3.265 86.345 3.59 ;
      RECT 86.34 3.782 86.345 4.448 ;
      RECT 86.33 3.265 86.34 3.58 ;
      RECT 86.335 3.835 86.34 4.451 ;
      RECT 86.33 3.92 86.335 4.455 ;
      RECT 86.32 3.265 86.33 3.568 ;
      RECT 86.325 3.967 86.33 4.459 ;
      RECT 86.32 4.042 86.325 4.463 ;
      RECT 86.285 3.265 86.32 3.543 ;
      RECT 86.31 4.125 86.32 4.468 ;
      RECT 86.3 4.192 86.31 4.475 ;
      RECT 86.295 4.22 86.3 4.48 ;
      RECT 86.285 4.233 86.295 4.486 ;
      RECT 86.24 3.265 86.285 3.5 ;
      RECT 86.28 4.238 86.285 4.493 ;
      RECT 86.24 4.255 86.28 4.555 ;
      RECT 86.235 3.267 86.24 3.473 ;
      RECT 86.21 4.275 86.24 4.555 ;
      RECT 86.23 3.272 86.235 3.445 ;
      RECT 86.02 4.284 86.06 4.555 ;
      RECT 85.995 4.292 86.02 4.525 ;
      RECT 85.95 4.3 85.995 4.525 ;
      RECT 85.935 4.305 85.95 4.52 ;
      RECT 85.925 4.305 85.935 4.514 ;
      RECT 85.915 4.312 85.925 4.511 ;
      RECT 85.91 4.35 85.915 4.5 ;
      RECT 85.905 4.412 85.91 4.478 ;
      RECT 87.175 4.287 87.36 4.51 ;
      RECT 87.175 4.302 87.365 4.506 ;
      RECT 87.165 3.575 87.25 4.505 ;
      RECT 87.165 4.302 87.37 4.499 ;
      RECT 87.16 4.31 87.37 4.498 ;
      RECT 87.365 4.03 87.685 4.35 ;
      RECT 87.16 4.202 87.33 4.293 ;
      RECT 87.155 4.202 87.33 4.275 ;
      RECT 87.145 4.01 87.28 4.25 ;
      RECT 87.14 4.01 87.28 4.195 ;
      RECT 87.1 3.59 87.27 4.095 ;
      RECT 87.085 3.59 87.27 3.965 ;
      RECT 87.08 3.59 87.27 3.918 ;
      RECT 87.075 3.59 87.27 3.898 ;
      RECT 87.07 3.59 87.27 3.873 ;
      RECT 87.04 3.59 87.3 3.85 ;
      RECT 87.05 3.587 87.26 3.85 ;
      RECT 87.175 3.582 87.26 4.51 ;
      RECT 87.06 3.575 87.25 3.85 ;
      RECT 87.055 3.58 87.25 3.85 ;
      RECT 85.885 3.792 86.07 4.005 ;
      RECT 85.885 3.8 86.08 3.998 ;
      RECT 85.865 3.8 86.08 3.995 ;
      RECT 85.86 3.8 86.08 3.98 ;
      RECT 85.79 3.715 86.05 3.975 ;
      RECT 85.79 3.86 86.085 3.888 ;
      RECT 85.445 4.315 85.705 4.575 ;
      RECT 85.47 4.26 85.665 4.575 ;
      RECT 85.465 4.009 85.645 4.303 ;
      RECT 85.465 4.015 85.655 4.303 ;
      RECT 85.445 4.017 85.655 4.248 ;
      RECT 85.44 4.027 85.655 4.115 ;
      RECT 85.47 4.007 85.645 4.575 ;
      RECT 85.556 4.005 85.645 4.575 ;
      RECT 85.415 3.225 85.45 3.595 ;
      RECT 85.205 3.335 85.21 3.595 ;
      RECT 85.45 3.232 85.465 3.595 ;
      RECT 85.34 3.225 85.415 3.673 ;
      RECT 85.33 3.225 85.34 3.758 ;
      RECT 85.305 3.225 85.33 3.793 ;
      RECT 85.265 3.225 85.305 3.861 ;
      RECT 85.255 3.232 85.265 3.913 ;
      RECT 85.225 3.335 85.255 3.954 ;
      RECT 85.22 3.335 85.225 3.993 ;
      RECT 85.21 3.335 85.22 4.013 ;
      RECT 85.205 3.63 85.21 4.05 ;
      RECT 85.2 3.647 85.205 4.07 ;
      RECT 85.185 3.71 85.2 4.11 ;
      RECT 85.18 3.753 85.185 4.145 ;
      RECT 85.175 3.761 85.18 4.158 ;
      RECT 85.165 3.775 85.175 4.18 ;
      RECT 85.14 3.81 85.165 4.245 ;
      RECT 85.13 3.845 85.14 4.308 ;
      RECT 85.11 3.875 85.13 4.369 ;
      RECT 85.095 3.911 85.11 4.436 ;
      RECT 85.085 3.939 85.095 4.475 ;
      RECT 85.075 3.961 85.085 4.495 ;
      RECT 85.07 3.971 85.075 4.506 ;
      RECT 85.065 3.98 85.07 4.509 ;
      RECT 85.055 3.998 85.065 4.513 ;
      RECT 85.045 4.016 85.055 4.514 ;
      RECT 85.02 4.055 85.045 4.511 ;
      RECT 85 4.097 85.02 4.508 ;
      RECT 84.985 4.135 85 4.507 ;
      RECT 84.95 4.17 84.985 4.504 ;
      RECT 84.945 4.192 84.95 4.502 ;
      RECT 84.88 4.232 84.945 4.499 ;
      RECT 84.875 4.272 84.88 4.495 ;
      RECT 84.86 4.282 84.875 4.486 ;
      RECT 84.85 4.402 84.86 4.471 ;
      RECT 85.33 4.815 85.34 5.075 ;
      RECT 85.33 4.818 85.35 5.074 ;
      RECT 85.32 4.808 85.33 5.073 ;
      RECT 85.31 4.823 85.39 5.069 ;
      RECT 85.295 4.802 85.31 5.067 ;
      RECT 85.27 4.827 85.395 5.063 ;
      RECT 85.255 4.787 85.27 5.058 ;
      RECT 85.255 4.829 85.405 5.057 ;
      RECT 85.255 4.837 85.42 5.05 ;
      RECT 85.195 4.774 85.255 5.04 ;
      RECT 85.185 4.761 85.195 5.022 ;
      RECT 85.16 4.751 85.185 5.012 ;
      RECT 85.155 4.741 85.16 5.004 ;
      RECT 85.09 4.837 85.42 4.986 ;
      RECT 85.005 4.837 85.42 4.948 ;
      RECT 84.895 4.665 85.155 4.925 ;
      RECT 85.27 4.795 85.295 5.063 ;
      RECT 85.31 4.805 85.32 5.069 ;
      RECT 84.895 4.813 85.335 4.925 ;
      RECT 85.08 10.06 85.37 10.29 ;
      RECT 85.14 9.32 85.31 10.29 ;
      RECT 85.04 9.345 85.41 9.715 ;
      RECT 85.08 9.32 85.37 9.715 ;
      RECT 84.11 4.57 84.14 4.87 ;
      RECT 83.885 4.555 83.89 4.83 ;
      RECT 83.685 4.555 83.84 4.815 ;
      RECT 84.985 3.27 85.015 3.53 ;
      RECT 84.975 3.27 84.985 3.638 ;
      RECT 84.955 3.27 84.975 3.648 ;
      RECT 84.94 3.27 84.955 3.66 ;
      RECT 84.885 3.27 84.94 3.71 ;
      RECT 84.87 3.27 84.885 3.758 ;
      RECT 84.84 3.27 84.87 3.793 ;
      RECT 84.785 3.27 84.84 3.855 ;
      RECT 84.765 3.27 84.785 3.923 ;
      RECT 84.76 3.27 84.765 3.953 ;
      RECT 84.755 3.27 84.76 3.965 ;
      RECT 84.75 3.387 84.755 3.983 ;
      RECT 84.73 3.405 84.75 4.008 ;
      RECT 84.71 3.432 84.73 4.058 ;
      RECT 84.705 3.452 84.71 4.089 ;
      RECT 84.7 3.46 84.705 4.106 ;
      RECT 84.685 3.486 84.7 4.135 ;
      RECT 84.67 3.528 84.685 4.17 ;
      RECT 84.665 3.557 84.67 4.193 ;
      RECT 84.66 3.572 84.665 4.206 ;
      RECT 84.655 3.595 84.66 4.217 ;
      RECT 84.645 3.615 84.655 4.235 ;
      RECT 84.635 3.645 84.645 4.258 ;
      RECT 84.63 3.667 84.635 4.278 ;
      RECT 84.625 3.682 84.63 4.293 ;
      RECT 84.61 3.712 84.625 4.32 ;
      RECT 84.605 3.742 84.61 4.346 ;
      RECT 84.6 3.76 84.605 4.358 ;
      RECT 84.59 3.79 84.6 4.377 ;
      RECT 84.58 3.815 84.59 4.402 ;
      RECT 84.575 3.835 84.58 4.421 ;
      RECT 84.57 3.852 84.575 4.434 ;
      RECT 84.56 3.878 84.57 4.453 ;
      RECT 84.55 3.916 84.56 4.48 ;
      RECT 84.545 3.942 84.55 4.5 ;
      RECT 84.54 3.952 84.545 4.51 ;
      RECT 84.535 3.965 84.54 4.525 ;
      RECT 84.53 3.98 84.535 4.535 ;
      RECT 84.525 4.002 84.53 4.55 ;
      RECT 84.52 4.02 84.525 4.561 ;
      RECT 84.515 4.03 84.52 4.572 ;
      RECT 84.51 4.038 84.515 4.584 ;
      RECT 84.505 4.046 84.51 4.595 ;
      RECT 84.5 4.072 84.505 4.608 ;
      RECT 84.49 4.1 84.5 4.621 ;
      RECT 84.485 4.13 84.49 4.63 ;
      RECT 84.48 4.145 84.485 4.637 ;
      RECT 84.465 4.17 84.48 4.644 ;
      RECT 84.46 4.192 84.465 4.65 ;
      RECT 84.455 4.217 84.46 4.653 ;
      RECT 84.446 4.245 84.455 4.657 ;
      RECT 84.44 4.262 84.446 4.662 ;
      RECT 84.435 4.28 84.44 4.666 ;
      RECT 84.43 4.292 84.435 4.669 ;
      RECT 84.425 4.313 84.43 4.673 ;
      RECT 84.42 4.331 84.425 4.676 ;
      RECT 84.415 4.345 84.42 4.679 ;
      RECT 84.41 4.362 84.415 4.682 ;
      RECT 84.405 4.375 84.41 4.685 ;
      RECT 84.38 4.412 84.405 4.693 ;
      RECT 84.375 4.457 84.38 4.702 ;
      RECT 84.37 4.485 84.375 4.705 ;
      RECT 84.36 4.505 84.37 4.709 ;
      RECT 84.355 4.525 84.36 4.714 ;
      RECT 84.35 4.54 84.355 4.717 ;
      RECT 84.33 4.55 84.35 4.724 ;
      RECT 84.265 4.557 84.33 4.75 ;
      RECT 84.23 4.56 84.265 4.778 ;
      RECT 84.215 4.563 84.23 4.793 ;
      RECT 84.205 4.564 84.215 4.808 ;
      RECT 84.195 4.565 84.205 4.825 ;
      RECT 84.19 4.565 84.195 4.84 ;
      RECT 84.185 4.565 84.19 4.848 ;
      RECT 84.17 4.566 84.185 4.863 ;
      RECT 84.14 4.568 84.17 4.87 ;
      RECT 84.03 4.575 84.11 4.87 ;
      RECT 83.985 4.58 84.03 4.87 ;
      RECT 83.975 4.581 83.985 4.86 ;
      RECT 83.965 4.582 83.975 4.853 ;
      RECT 83.945 4.584 83.965 4.848 ;
      RECT 83.935 4.555 83.945 4.843 ;
      RECT 83.89 4.555 83.935 4.835 ;
      RECT 83.86 4.555 83.885 4.825 ;
      RECT 83.84 4.555 83.86 4.818 ;
      RECT 84.12 3.355 84.38 3.615 ;
      RECT 84 3.37 84.01 3.535 ;
      RECT 83.985 3.37 83.99 3.53 ;
      RECT 81.35 3.21 81.535 3.5 ;
      RECT 83.165 3.335 83.18 3.49 ;
      RECT 81.315 3.21 81.34 3.47 ;
      RECT 83.73 3.26 83.735 3.402 ;
      RECT 83.645 3.255 83.67 3.395 ;
      RECT 84.045 3.372 84.12 3.565 ;
      RECT 84.03 3.37 84.045 3.548 ;
      RECT 84.01 3.37 84.03 3.54 ;
      RECT 83.99 3.37 84 3.533 ;
      RECT 83.945 3.365 83.985 3.523 ;
      RECT 83.905 3.34 83.945 3.508 ;
      RECT 83.89 3.315 83.905 3.498 ;
      RECT 83.885 3.309 83.89 3.496 ;
      RECT 83.85 3.301 83.885 3.479 ;
      RECT 83.845 3.294 83.85 3.467 ;
      RECT 83.825 3.289 83.845 3.455 ;
      RECT 83.815 3.283 83.825 3.44 ;
      RECT 83.795 3.278 83.815 3.425 ;
      RECT 83.785 3.273 83.795 3.418 ;
      RECT 83.78 3.271 83.785 3.413 ;
      RECT 83.775 3.27 83.78 3.41 ;
      RECT 83.735 3.265 83.775 3.406 ;
      RECT 83.715 3.259 83.73 3.401 ;
      RECT 83.68 3.256 83.715 3.398 ;
      RECT 83.67 3.255 83.68 3.396 ;
      RECT 83.61 3.255 83.645 3.393 ;
      RECT 83.565 3.255 83.61 3.393 ;
      RECT 83.515 3.255 83.565 3.396 ;
      RECT 83.5 3.257 83.515 3.398 ;
      RECT 83.485 3.26 83.5 3.399 ;
      RECT 83.475 3.265 83.485 3.4 ;
      RECT 83.445 3.27 83.475 3.405 ;
      RECT 83.435 3.276 83.445 3.413 ;
      RECT 83.425 3.278 83.435 3.417 ;
      RECT 83.415 3.282 83.425 3.421 ;
      RECT 83.39 3.288 83.415 3.429 ;
      RECT 83.38 3.293 83.39 3.437 ;
      RECT 83.365 3.297 83.38 3.441 ;
      RECT 83.33 3.303 83.365 3.449 ;
      RECT 83.31 3.308 83.33 3.459 ;
      RECT 83.28 3.315 83.31 3.468 ;
      RECT 83.235 3.324 83.28 3.482 ;
      RECT 83.23 3.329 83.235 3.493 ;
      RECT 83.21 3.332 83.23 3.494 ;
      RECT 83.18 3.335 83.21 3.492 ;
      RECT 83.145 3.335 83.165 3.488 ;
      RECT 83.075 3.335 83.145 3.479 ;
      RECT 83.06 3.332 83.075 3.471 ;
      RECT 83.02 3.325 83.06 3.466 ;
      RECT 82.995 3.315 83.02 3.459 ;
      RECT 82.99 3.309 82.995 3.456 ;
      RECT 82.95 3.303 82.99 3.453 ;
      RECT 82.935 3.296 82.95 3.448 ;
      RECT 82.915 3.292 82.935 3.443 ;
      RECT 82.9 3.287 82.915 3.439 ;
      RECT 82.885 3.282 82.9 3.437 ;
      RECT 82.87 3.278 82.885 3.436 ;
      RECT 82.855 3.276 82.87 3.432 ;
      RECT 82.845 3.274 82.855 3.427 ;
      RECT 82.83 3.271 82.845 3.423 ;
      RECT 82.82 3.269 82.83 3.418 ;
      RECT 82.8 3.266 82.82 3.414 ;
      RECT 82.755 3.265 82.8 3.412 ;
      RECT 82.695 3.267 82.755 3.413 ;
      RECT 82.675 3.269 82.695 3.415 ;
      RECT 82.645 3.272 82.675 3.416 ;
      RECT 82.595 3.277 82.645 3.418 ;
      RECT 82.59 3.28 82.595 3.42 ;
      RECT 82.58 3.282 82.59 3.423 ;
      RECT 82.575 3.284 82.58 3.426 ;
      RECT 82.525 3.287 82.575 3.433 ;
      RECT 82.505 3.291 82.525 3.445 ;
      RECT 82.495 3.294 82.505 3.451 ;
      RECT 82.485 3.295 82.495 3.454 ;
      RECT 82.446 3.298 82.485 3.456 ;
      RECT 82.36 3.305 82.446 3.459 ;
      RECT 82.286 3.315 82.36 3.463 ;
      RECT 82.2 3.326 82.286 3.468 ;
      RECT 82.185 3.333 82.2 3.47 ;
      RECT 82.13 3.337 82.185 3.471 ;
      RECT 82.116 3.34 82.13 3.473 ;
      RECT 82.03 3.34 82.116 3.475 ;
      RECT 81.99 3.337 82.03 3.478 ;
      RECT 81.966 3.333 81.99 3.48 ;
      RECT 81.88 3.323 81.966 3.483 ;
      RECT 81.85 3.312 81.88 3.484 ;
      RECT 81.831 3.308 81.85 3.483 ;
      RECT 81.745 3.301 81.831 3.48 ;
      RECT 81.685 3.29 81.745 3.477 ;
      RECT 81.665 3.282 81.685 3.475 ;
      RECT 81.63 3.277 81.665 3.474 ;
      RECT 81.605 3.272 81.63 3.473 ;
      RECT 81.575 3.267 81.605 3.472 ;
      RECT 81.55 3.21 81.575 3.471 ;
      RECT 81.535 3.21 81.55 3.495 ;
      RECT 81.34 3.21 81.35 3.495 ;
      RECT 83.115 4.23 83.12 4.37 ;
      RECT 82.775 4.23 82.81 4.368 ;
      RECT 82.35 4.215 82.365 4.36 ;
      RECT 84.18 3.995 84.27 4.255 ;
      RECT 84.01 3.86 84.11 4.255 ;
      RECT 81.045 3.835 81.125 4.045 ;
      RECT 84.135 3.972 84.18 4.255 ;
      RECT 84.125 3.942 84.135 4.255 ;
      RECT 84.11 3.865 84.125 4.255 ;
      RECT 83.925 3.86 84.01 4.22 ;
      RECT 83.92 3.862 83.925 4.215 ;
      RECT 83.915 3.867 83.92 4.215 ;
      RECT 83.88 3.967 83.915 4.215 ;
      RECT 83.87 3.995 83.88 4.215 ;
      RECT 83.86 4.01 83.87 4.215 ;
      RECT 83.85 4.022 83.86 4.215 ;
      RECT 83.845 4.032 83.85 4.215 ;
      RECT 83.83 4.042 83.845 4.217 ;
      RECT 83.825 4.057 83.83 4.219 ;
      RECT 83.81 4.07 83.825 4.221 ;
      RECT 83.805 4.085 83.81 4.224 ;
      RECT 83.785 4.095 83.805 4.228 ;
      RECT 83.77 4.105 83.785 4.231 ;
      RECT 83.735 4.112 83.77 4.236 ;
      RECT 83.691 4.119 83.735 4.244 ;
      RECT 83.605 4.131 83.691 4.257 ;
      RECT 83.58 4.142 83.605 4.268 ;
      RECT 83.55 4.147 83.58 4.273 ;
      RECT 83.515 4.152 83.55 4.281 ;
      RECT 83.485 4.157 83.515 4.288 ;
      RECT 83.46 4.162 83.485 4.293 ;
      RECT 83.395 4.169 83.46 4.302 ;
      RECT 83.325 4.182 83.395 4.318 ;
      RECT 83.295 4.192 83.325 4.33 ;
      RECT 83.27 4.197 83.295 4.337 ;
      RECT 83.215 4.204 83.27 4.345 ;
      RECT 83.21 4.211 83.215 4.35 ;
      RECT 83.205 4.213 83.21 4.351 ;
      RECT 83.19 4.215 83.205 4.353 ;
      RECT 83.185 4.215 83.19 4.356 ;
      RECT 83.12 4.222 83.185 4.363 ;
      RECT 83.085 4.232 83.115 4.373 ;
      RECT 83.068 4.235 83.085 4.375 ;
      RECT 82.982 4.234 83.068 4.374 ;
      RECT 82.896 4.232 82.982 4.371 ;
      RECT 82.81 4.231 82.896 4.369 ;
      RECT 82.709 4.229 82.775 4.368 ;
      RECT 82.623 4.226 82.709 4.366 ;
      RECT 82.537 4.222 82.623 4.364 ;
      RECT 82.451 4.219 82.537 4.363 ;
      RECT 82.365 4.216 82.451 4.361 ;
      RECT 82.265 4.215 82.35 4.358 ;
      RECT 82.215 4.213 82.265 4.356 ;
      RECT 82.195 4.21 82.215 4.354 ;
      RECT 82.175 4.208 82.195 4.351 ;
      RECT 82.15 4.204 82.175 4.348 ;
      RECT 82.105 4.198 82.15 4.343 ;
      RECT 82.065 4.192 82.105 4.335 ;
      RECT 82.04 4.187 82.065 4.328 ;
      RECT 81.985 4.18 82.04 4.32 ;
      RECT 81.961 4.173 81.985 4.313 ;
      RECT 81.875 4.164 81.961 4.303 ;
      RECT 81.845 4.156 81.875 4.293 ;
      RECT 81.815 4.152 81.845 4.288 ;
      RECT 81.81 4.149 81.815 4.285 ;
      RECT 81.805 4.148 81.81 4.285 ;
      RECT 81.73 4.141 81.805 4.278 ;
      RECT 81.691 4.132 81.73 4.267 ;
      RECT 81.605 4.122 81.691 4.255 ;
      RECT 81.565 4.112 81.605 4.243 ;
      RECT 81.526 4.107 81.565 4.236 ;
      RECT 81.44 4.097 81.526 4.225 ;
      RECT 81.4 4.085 81.44 4.214 ;
      RECT 81.365 4.07 81.4 4.207 ;
      RECT 81.355 4.06 81.365 4.204 ;
      RECT 81.335 4.045 81.355 4.202 ;
      RECT 81.305 4.015 81.335 4.198 ;
      RECT 81.295 3.995 81.305 4.193 ;
      RECT 81.29 3.987 81.295 4.19 ;
      RECT 81.285 3.98 81.29 4.188 ;
      RECT 81.27 3.967 81.285 4.181 ;
      RECT 81.265 3.957 81.27 4.173 ;
      RECT 81.26 3.95 81.265 4.168 ;
      RECT 81.255 3.945 81.26 4.164 ;
      RECT 81.24 3.932 81.255 4.156 ;
      RECT 81.235 3.842 81.24 4.145 ;
      RECT 81.23 3.837 81.235 4.138 ;
      RECT 81.155 3.835 81.23 4.098 ;
      RECT 81.125 3.835 81.155 4.053 ;
      RECT 81.03 3.84 81.045 4.04 ;
      RECT 83.515 3.545 83.775 3.805 ;
      RECT 83.5 3.533 83.68 3.77 ;
      RECT 83.495 3.534 83.68 3.768 ;
      RECT 83.48 3.538 83.69 3.758 ;
      RECT 83.475 3.543 83.695 3.728 ;
      RECT 83.48 3.54 83.695 3.758 ;
      RECT 83.495 3.535 83.69 3.768 ;
      RECT 83.515 3.532 83.68 3.805 ;
      RECT 83.515 3.531 83.67 3.805 ;
      RECT 83.54 3.53 83.67 3.805 ;
      RECT 83.1 3.775 83.36 4.035 ;
      RECT 82.975 3.82 83.36 4.03 ;
      RECT 82.965 3.825 83.36 4.025 ;
      RECT 82.98 4.765 82.995 5.075 ;
      RECT 81.575 4.535 81.585 4.665 ;
      RECT 81.355 4.53 81.46 4.665 ;
      RECT 81.27 4.535 81.32 4.665 ;
      RECT 79.82 3.27 79.825 4.375 ;
      RECT 83.075 4.857 83.08 4.993 ;
      RECT 83.07 4.852 83.075 5.053 ;
      RECT 83.065 4.85 83.07 5.066 ;
      RECT 83.05 4.847 83.065 5.068 ;
      RECT 83.045 4.842 83.05 5.07 ;
      RECT 83.04 4.838 83.045 5.073 ;
      RECT 83.025 4.833 83.04 5.075 ;
      RECT 82.995 4.825 83.025 5.075 ;
      RECT 82.956 4.765 82.98 5.075 ;
      RECT 82.87 4.765 82.956 5.072 ;
      RECT 82.84 4.765 82.87 5.065 ;
      RECT 82.815 4.765 82.84 5.058 ;
      RECT 82.79 4.765 82.815 5.05 ;
      RECT 82.775 4.765 82.79 5.043 ;
      RECT 82.75 4.765 82.775 5.035 ;
      RECT 82.735 4.765 82.75 5.028 ;
      RECT 82.695 4.775 82.735 5.017 ;
      RECT 82.685 4.77 82.695 5.007 ;
      RECT 82.681 4.769 82.685 5.004 ;
      RECT 82.595 4.761 82.681 4.987 ;
      RECT 82.562 4.75 82.595 4.964 ;
      RECT 82.476 4.739 82.562 4.942 ;
      RECT 82.39 4.723 82.476 4.911 ;
      RECT 82.32 4.708 82.39 4.883 ;
      RECT 82.31 4.701 82.32 4.87 ;
      RECT 82.28 4.698 82.31 4.86 ;
      RECT 82.255 4.694 82.28 4.853 ;
      RECT 82.24 4.691 82.255 4.848 ;
      RECT 82.235 4.69 82.24 4.843 ;
      RECT 82.205 4.685 82.235 4.836 ;
      RECT 82.2 4.68 82.205 4.831 ;
      RECT 82.185 4.677 82.2 4.826 ;
      RECT 82.18 4.672 82.185 4.821 ;
      RECT 82.16 4.667 82.18 4.818 ;
      RECT 82.145 4.662 82.16 4.81 ;
      RECT 82.13 4.656 82.145 4.805 ;
      RECT 82.1 4.647 82.13 4.798 ;
      RECT 82.095 4.64 82.1 4.79 ;
      RECT 82.09 4.638 82.095 4.788 ;
      RECT 82.085 4.637 82.09 4.785 ;
      RECT 82.045 4.63 82.085 4.778 ;
      RECT 82.031 4.62 82.045 4.768 ;
      RECT 81.98 4.609 82.031 4.756 ;
      RECT 81.955 4.595 81.98 4.742 ;
      RECT 81.93 4.584 81.955 4.734 ;
      RECT 81.91 4.573 81.93 4.728 ;
      RECT 81.9 4.567 81.91 4.723 ;
      RECT 81.895 4.565 81.9 4.719 ;
      RECT 81.875 4.56 81.895 4.714 ;
      RECT 81.845 4.55 81.875 4.704 ;
      RECT 81.84 4.542 81.845 4.697 ;
      RECT 81.825 4.54 81.84 4.693 ;
      RECT 81.805 4.54 81.825 4.688 ;
      RECT 81.8 4.539 81.805 4.686 ;
      RECT 81.795 4.539 81.8 4.683 ;
      RECT 81.755 4.538 81.795 4.678 ;
      RECT 81.73 4.537 81.755 4.673 ;
      RECT 81.67 4.536 81.73 4.67 ;
      RECT 81.585 4.535 81.67 4.668 ;
      RECT 81.546 4.534 81.575 4.665 ;
      RECT 81.46 4.532 81.546 4.665 ;
      RECT 81.32 4.532 81.355 4.665 ;
      RECT 81.23 4.536 81.27 4.668 ;
      RECT 81.215 4.539 81.23 4.675 ;
      RECT 81.205 4.54 81.215 4.682 ;
      RECT 81.18 4.543 81.205 4.687 ;
      RECT 81.175 4.545 81.18 4.69 ;
      RECT 81.125 4.547 81.175 4.691 ;
      RECT 81.086 4.551 81.125 4.693 ;
      RECT 81 4.553 81.086 4.696 ;
      RECT 80.982 4.555 81 4.698 ;
      RECT 80.896 4.558 80.982 4.7 ;
      RECT 80.81 4.562 80.896 4.703 ;
      RECT 80.773 4.566 80.81 4.706 ;
      RECT 80.687 4.569 80.773 4.709 ;
      RECT 80.601 4.573 80.687 4.712 ;
      RECT 80.515 4.578 80.601 4.716 ;
      RECT 80.495 4.58 80.515 4.719 ;
      RECT 80.475 4.579 80.495 4.72 ;
      RECT 80.426 4.576 80.475 4.721 ;
      RECT 80.34 4.571 80.426 4.724 ;
      RECT 80.29 4.566 80.34 4.726 ;
      RECT 80.266 4.564 80.29 4.727 ;
      RECT 80.18 4.559 80.266 4.729 ;
      RECT 80.155 4.555 80.18 4.728 ;
      RECT 80.145 4.552 80.155 4.726 ;
      RECT 80.135 4.545 80.145 4.723 ;
      RECT 80.13 4.525 80.135 4.718 ;
      RECT 80.12 4.495 80.13 4.713 ;
      RECT 80.105 4.365 80.12 4.704 ;
      RECT 80.1 4.357 80.105 4.697 ;
      RECT 80.08 4.35 80.1 4.689 ;
      RECT 80.075 4.332 80.08 4.681 ;
      RECT 80.065 4.312 80.075 4.676 ;
      RECT 80.06 4.285 80.065 4.672 ;
      RECT 80.055 4.262 80.06 4.669 ;
      RECT 80.035 4.22 80.055 4.661 ;
      RECT 80 4.135 80.035 4.645 ;
      RECT 79.995 4.067 80 4.633 ;
      RECT 79.98 4.037 79.995 4.627 ;
      RECT 79.975 3.282 79.98 3.528 ;
      RECT 79.965 4.007 79.98 4.618 ;
      RECT 79.97 3.277 79.975 3.56 ;
      RECT 79.965 3.272 79.97 3.603 ;
      RECT 79.96 3.27 79.965 3.638 ;
      RECT 79.945 3.97 79.965 4.608 ;
      RECT 79.955 3.27 79.96 3.675 ;
      RECT 79.94 3.27 79.955 3.773 ;
      RECT 79.94 3.943 79.945 4.601 ;
      RECT 79.935 3.27 79.94 3.848 ;
      RECT 79.935 3.931 79.94 4.598 ;
      RECT 79.93 3.27 79.935 3.88 ;
      RECT 79.93 3.91 79.935 4.595 ;
      RECT 79.925 3.27 79.93 4.592 ;
      RECT 79.89 3.27 79.925 4.578 ;
      RECT 79.875 3.27 79.89 4.56 ;
      RECT 79.855 3.27 79.875 4.55 ;
      RECT 79.83 3.27 79.855 4.533 ;
      RECT 79.825 3.27 79.83 4.483 ;
      RECT 79.815 3.27 79.82 4.313 ;
      RECT 79.81 3.27 79.815 4.22 ;
      RECT 79.805 3.27 79.81 4.133 ;
      RECT 79.8 3.27 79.805 4.065 ;
      RECT 79.795 3.27 79.8 4.008 ;
      RECT 79.785 3.27 79.795 3.903 ;
      RECT 79.78 3.27 79.785 3.775 ;
      RECT 79.775 3.27 79.78 3.693 ;
      RECT 79.77 3.272 79.775 3.61 ;
      RECT 79.765 3.277 79.77 3.543 ;
      RECT 79.76 3.282 79.765 3.47 ;
      RECT 82.575 3.6 82.835 3.86 ;
      RECT 82.595 3.567 82.805 3.86 ;
      RECT 82.595 3.565 82.795 3.86 ;
      RECT 82.605 3.552 82.795 3.86 ;
      RECT 82.605 3.55 82.72 3.86 ;
      RECT 82.08 3.675 82.255 3.955 ;
      RECT 82.075 3.675 82.255 3.953 ;
      RECT 82.075 3.675 82.27 3.95 ;
      RECT 82.065 3.675 82.27 3.948 ;
      RECT 82.01 3.675 82.27 3.935 ;
      RECT 82.01 3.75 82.275 3.913 ;
      RECT 81.54 4.873 81.545 5.08 ;
      RECT 81.49 4.867 81.54 5.079 ;
      RECT 81.457 4.881 81.55 5.078 ;
      RECT 81.371 4.881 81.55 5.077 ;
      RECT 81.285 4.881 81.55 5.076 ;
      RECT 81.285 4.98 81.555 5.073 ;
      RECT 81.28 4.98 81.555 5.068 ;
      RECT 81.275 4.98 81.555 5.05 ;
      RECT 81.27 4.98 81.555 5.033 ;
      RECT 81.23 4.765 81.49 5.025 ;
      RECT 80.69 3.915 80.776 4.329 ;
      RECT 80.69 3.915 80.815 4.326 ;
      RECT 80.69 3.915 80.835 4.316 ;
      RECT 80.645 3.915 80.835 4.313 ;
      RECT 80.645 4.067 80.845 4.303 ;
      RECT 80.645 4.088 80.85 4.297 ;
      RECT 80.645 4.106 80.855 4.293 ;
      RECT 80.645 4.126 80.865 4.288 ;
      RECT 80.62 4.126 80.865 4.285 ;
      RECT 80.61 4.126 80.865 4.263 ;
      RECT 80.61 4.142 80.87 4.233 ;
      RECT 80.575 3.915 80.835 4.22 ;
      RECT 80.575 4.154 80.875 4.175 ;
      RECT 78.235 10.06 78.53 10.29 ;
      RECT 78.295 8.58 78.465 10.29 ;
      RECT 78.245 8.95 78.595 9.3 ;
      RECT 78.235 8.58 78.525 8.81 ;
      RECT 77.245 10.06 77.54 10.29 ;
      RECT 77.305 8.58 77.475 10.29 ;
      RECT 77.245 8.58 77.535 8.81 ;
      RECT 77.245 8.615 78.095 8.775 ;
      RECT 77.93 8.21 78.095 8.775 ;
      RECT 77.245 8.61 77.64 8.775 ;
      RECT 77.865 8.21 78.155 8.44 ;
      RECT 77.865 8.24 78.325 8.41 ;
      RECT 77.83 4.005 78.15 4.26 ;
      RECT 77.83 4.055 78.32 4.225 ;
      RECT 77.83 3.69 78.02 4.26 ;
      RECT 77.245 3.655 77.535 3.885 ;
      RECT 77.245 3.69 78.02 3.86 ;
      RECT 77.305 2.175 77.475 3.885 ;
      RECT 77.245 2.175 77.54 2.405 ;
      RECT 76.875 4.025 77.165 4.255 ;
      RECT 76.875 4.055 77.335 4.225 ;
      RECT 76.94 2.95 77.105 4.255 ;
      RECT 75.455 2.915 75.745 3.145 ;
      RECT 75.455 2.95 77.105 3.12 ;
      RECT 75.515 2.175 75.685 3.145 ;
      RECT 75.455 2.175 75.745 2.405 ;
      RECT 75.455 10.06 75.745 10.29 ;
      RECT 75.515 9.32 75.685 10.29 ;
      RECT 75.515 9.41 77.105 9.58 ;
      RECT 76.935 8.21 77.105 9.58 ;
      RECT 75.455 9.32 75.745 9.55 ;
      RECT 76.875 8.21 77.165 8.44 ;
      RECT 76.875 8.24 77.335 8.41 ;
      RECT 73.505 4 73.845 4.35 ;
      RECT 73.595 3.32 73.765 4.35 ;
      RECT 75.885 3.26 76.235 3.61 ;
      RECT 73.595 3.32 76.235 3.49 ;
      RECT 75.715 3.315 76.235 3.49 ;
      RECT 75.91 8.945 76.235 9.27 ;
      RECT 70.45 8.905 70.8 9.255 ;
      RECT 75.885 8.95 76.235 9.18 ;
      RECT 70.25 8.95 70.8 9.18 ;
      RECT 75.715 8.975 76.235 9.15 ;
      RECT 70.08 8.98 70.8 9.15 ;
      RECT 70.13 8.975 76.235 9.145 ;
      RECT 75.11 3.66 75.43 3.98 ;
      RECT 75.085 3.655 75.375 3.885 ;
      RECT 75.08 3.685 75.43 3.86 ;
      RECT 74.91 3.685 75.43 3.855 ;
      RECT 75.11 8.545 75.43 8.835 ;
      RECT 75.085 8.58 75.43 8.81 ;
      RECT 74.91 8.61 75.43 8.78 ;
      RECT 70.8 4.28 70.95 4.555 ;
      RECT 71.34 3.36 71.345 3.58 ;
      RECT 72.49 3.56 72.505 3.758 ;
      RECT 72.455 3.552 72.49 3.765 ;
      RECT 72.425 3.545 72.455 3.765 ;
      RECT 72.37 3.51 72.425 3.765 ;
      RECT 72.305 3.447 72.37 3.765 ;
      RECT 72.3 3.412 72.305 3.763 ;
      RECT 72.295 3.407 72.3 3.755 ;
      RECT 72.29 3.402 72.295 3.741 ;
      RECT 72.285 3.399 72.29 3.734 ;
      RECT 72.24 3.389 72.285 3.685 ;
      RECT 72.22 3.376 72.24 3.62 ;
      RECT 72.215 3.371 72.22 3.593 ;
      RECT 72.21 3.37 72.215 3.586 ;
      RECT 72.205 3.369 72.21 3.579 ;
      RECT 72.12 3.354 72.205 3.525 ;
      RECT 72.09 3.335 72.12 3.475 ;
      RECT 72.01 3.318 72.09 3.46 ;
      RECT 71.975 3.305 72.01 3.445 ;
      RECT 71.967 3.305 71.975 3.44 ;
      RECT 71.881 3.306 71.967 3.44 ;
      RECT 71.795 3.308 71.881 3.44 ;
      RECT 71.77 3.309 71.795 3.444 ;
      RECT 71.695 3.315 71.77 3.459 ;
      RECT 71.612 3.327 71.695 3.483 ;
      RECT 71.526 3.34 71.612 3.509 ;
      RECT 71.44 3.353 71.526 3.535 ;
      RECT 71.405 3.362 71.44 3.554 ;
      RECT 71.355 3.362 71.405 3.567 ;
      RECT 71.345 3.36 71.355 3.578 ;
      RECT 71.33 3.357 71.34 3.58 ;
      RECT 71.315 3.349 71.33 3.588 ;
      RECT 71.3 3.341 71.315 3.608 ;
      RECT 71.295 3.336 71.3 3.665 ;
      RECT 71.28 3.331 71.295 3.738 ;
      RECT 71.275 3.326 71.28 3.78 ;
      RECT 71.27 3.324 71.275 3.808 ;
      RECT 71.265 3.322 71.27 3.83 ;
      RECT 71.255 3.318 71.265 3.873 ;
      RECT 71.25 3.315 71.255 3.898 ;
      RECT 71.245 3.313 71.25 3.918 ;
      RECT 71.24 3.311 71.245 3.942 ;
      RECT 71.235 3.307 71.24 3.965 ;
      RECT 71.23 3.303 71.235 3.988 ;
      RECT 71.195 3.293 71.23 4.095 ;
      RECT 71.19 3.283 71.195 4.193 ;
      RECT 71.185 3.281 71.19 4.22 ;
      RECT 71.18 3.28 71.185 4.24 ;
      RECT 71.175 3.272 71.18 4.26 ;
      RECT 71.17 3.267 71.175 4.295 ;
      RECT 71.165 3.265 71.17 4.313 ;
      RECT 71.16 3.265 71.165 4.338 ;
      RECT 71.155 3.265 71.16 4.36 ;
      RECT 71.12 3.265 71.155 4.403 ;
      RECT 71.095 3.265 71.12 4.432 ;
      RECT 71.085 3.265 71.095 3.618 ;
      RECT 71.088 3.675 71.095 4.442 ;
      RECT 71.085 3.732 71.088 4.445 ;
      RECT 71.08 3.265 71.085 3.59 ;
      RECT 71.08 3.782 71.085 4.448 ;
      RECT 71.07 3.265 71.08 3.58 ;
      RECT 71.075 3.835 71.08 4.451 ;
      RECT 71.07 3.92 71.075 4.455 ;
      RECT 71.06 3.265 71.07 3.568 ;
      RECT 71.065 3.967 71.07 4.459 ;
      RECT 71.06 4.042 71.065 4.463 ;
      RECT 71.025 3.265 71.06 3.543 ;
      RECT 71.05 4.125 71.06 4.468 ;
      RECT 71.04 4.192 71.05 4.475 ;
      RECT 71.035 4.22 71.04 4.48 ;
      RECT 71.025 4.233 71.035 4.486 ;
      RECT 70.98 3.265 71.025 3.5 ;
      RECT 71.02 4.238 71.025 4.493 ;
      RECT 70.98 4.255 71.02 4.555 ;
      RECT 70.975 3.267 70.98 3.473 ;
      RECT 70.95 4.275 70.98 4.555 ;
      RECT 70.97 3.272 70.975 3.445 ;
      RECT 70.76 4.284 70.8 4.555 ;
      RECT 70.735 4.292 70.76 4.525 ;
      RECT 70.69 4.3 70.735 4.525 ;
      RECT 70.675 4.305 70.69 4.52 ;
      RECT 70.665 4.305 70.675 4.514 ;
      RECT 70.655 4.312 70.665 4.511 ;
      RECT 70.65 4.35 70.655 4.5 ;
      RECT 70.645 4.412 70.65 4.478 ;
      RECT 71.915 4.287 72.1 4.51 ;
      RECT 71.915 4.302 72.105 4.506 ;
      RECT 71.905 3.575 71.99 4.505 ;
      RECT 71.905 4.302 72.11 4.499 ;
      RECT 71.9 4.31 72.11 4.498 ;
      RECT 72.105 4.03 72.425 4.35 ;
      RECT 71.9 4.202 72.07 4.293 ;
      RECT 71.895 4.202 72.07 4.275 ;
      RECT 71.885 4.01 72.02 4.25 ;
      RECT 71.88 4.01 72.02 4.195 ;
      RECT 71.84 3.59 72.01 4.095 ;
      RECT 71.825 3.59 72.01 3.965 ;
      RECT 71.82 3.59 72.01 3.918 ;
      RECT 71.815 3.59 72.01 3.898 ;
      RECT 71.81 3.59 72.01 3.873 ;
      RECT 71.78 3.59 72.04 3.85 ;
      RECT 71.79 3.587 72 3.85 ;
      RECT 71.915 3.582 72 4.51 ;
      RECT 71.8 3.575 71.99 3.85 ;
      RECT 71.795 3.58 71.99 3.85 ;
      RECT 70.625 3.792 70.81 4.005 ;
      RECT 70.625 3.8 70.82 3.998 ;
      RECT 70.605 3.8 70.82 3.995 ;
      RECT 70.6 3.8 70.82 3.98 ;
      RECT 70.53 3.715 70.79 3.975 ;
      RECT 70.53 3.86 70.825 3.888 ;
      RECT 70.185 4.315 70.445 4.575 ;
      RECT 70.21 4.26 70.405 4.575 ;
      RECT 70.205 4.009 70.385 4.303 ;
      RECT 70.205 4.015 70.395 4.303 ;
      RECT 70.185 4.017 70.395 4.248 ;
      RECT 70.18 4.027 70.395 4.115 ;
      RECT 70.21 4.007 70.385 4.575 ;
      RECT 70.296 4.005 70.385 4.575 ;
      RECT 70.155 3.225 70.19 3.595 ;
      RECT 69.945 3.335 69.95 3.595 ;
      RECT 70.19 3.232 70.205 3.595 ;
      RECT 70.08 3.225 70.155 3.673 ;
      RECT 70.07 3.225 70.08 3.758 ;
      RECT 70.045 3.225 70.07 3.793 ;
      RECT 70.005 3.225 70.045 3.861 ;
      RECT 69.995 3.232 70.005 3.913 ;
      RECT 69.965 3.335 69.995 3.954 ;
      RECT 69.96 3.335 69.965 3.993 ;
      RECT 69.95 3.335 69.96 4.013 ;
      RECT 69.945 3.63 69.95 4.05 ;
      RECT 69.94 3.647 69.945 4.07 ;
      RECT 69.925 3.71 69.94 4.11 ;
      RECT 69.92 3.753 69.925 4.145 ;
      RECT 69.915 3.761 69.92 4.158 ;
      RECT 69.905 3.775 69.915 4.18 ;
      RECT 69.88 3.81 69.905 4.245 ;
      RECT 69.87 3.845 69.88 4.308 ;
      RECT 69.85 3.875 69.87 4.369 ;
      RECT 69.835 3.911 69.85 4.436 ;
      RECT 69.825 3.939 69.835 4.475 ;
      RECT 69.815 3.961 69.825 4.495 ;
      RECT 69.81 3.971 69.815 4.506 ;
      RECT 69.805 3.98 69.81 4.509 ;
      RECT 69.795 3.998 69.805 4.513 ;
      RECT 69.785 4.016 69.795 4.514 ;
      RECT 69.76 4.055 69.785 4.511 ;
      RECT 69.74 4.097 69.76 4.508 ;
      RECT 69.725 4.135 69.74 4.507 ;
      RECT 69.69 4.17 69.725 4.504 ;
      RECT 69.685 4.192 69.69 4.502 ;
      RECT 69.62 4.232 69.685 4.499 ;
      RECT 69.615 4.272 69.62 4.495 ;
      RECT 69.6 4.282 69.615 4.486 ;
      RECT 69.59 4.402 69.6 4.471 ;
      RECT 70.07 4.815 70.08 5.075 ;
      RECT 70.07 4.818 70.09 5.074 ;
      RECT 70.06 4.808 70.07 5.073 ;
      RECT 70.05 4.823 70.13 5.069 ;
      RECT 70.035 4.802 70.05 5.067 ;
      RECT 70.01 4.827 70.135 5.063 ;
      RECT 69.995 4.787 70.01 5.058 ;
      RECT 69.995 4.829 70.145 5.057 ;
      RECT 69.995 4.837 70.16 5.05 ;
      RECT 69.935 4.774 69.995 5.04 ;
      RECT 69.925 4.761 69.935 5.022 ;
      RECT 69.9 4.751 69.925 5.012 ;
      RECT 69.895 4.741 69.9 5.004 ;
      RECT 69.83 4.837 70.16 4.986 ;
      RECT 69.745 4.837 70.16 4.948 ;
      RECT 69.635 4.665 69.895 4.925 ;
      RECT 70.01 4.795 70.035 5.063 ;
      RECT 70.05 4.805 70.06 5.069 ;
      RECT 69.635 4.813 70.075 4.925 ;
      RECT 69.82 10.06 70.11 10.29 ;
      RECT 69.88 9.32 70.05 10.29 ;
      RECT 69.78 9.345 70.15 9.715 ;
      RECT 69.82 9.32 70.11 9.715 ;
      RECT 68.85 4.57 68.88 4.87 ;
      RECT 68.625 4.555 68.63 4.83 ;
      RECT 68.425 4.555 68.58 4.815 ;
      RECT 69.725 3.27 69.755 3.53 ;
      RECT 69.715 3.27 69.725 3.638 ;
      RECT 69.695 3.27 69.715 3.648 ;
      RECT 69.68 3.27 69.695 3.66 ;
      RECT 69.625 3.27 69.68 3.71 ;
      RECT 69.61 3.27 69.625 3.758 ;
      RECT 69.58 3.27 69.61 3.793 ;
      RECT 69.525 3.27 69.58 3.855 ;
      RECT 69.505 3.27 69.525 3.923 ;
      RECT 69.5 3.27 69.505 3.953 ;
      RECT 69.495 3.27 69.5 3.965 ;
      RECT 69.49 3.387 69.495 3.983 ;
      RECT 69.47 3.405 69.49 4.008 ;
      RECT 69.45 3.432 69.47 4.058 ;
      RECT 69.445 3.452 69.45 4.089 ;
      RECT 69.44 3.46 69.445 4.106 ;
      RECT 69.425 3.486 69.44 4.135 ;
      RECT 69.41 3.528 69.425 4.17 ;
      RECT 69.405 3.557 69.41 4.193 ;
      RECT 69.4 3.572 69.405 4.206 ;
      RECT 69.395 3.595 69.4 4.217 ;
      RECT 69.385 3.615 69.395 4.235 ;
      RECT 69.375 3.645 69.385 4.258 ;
      RECT 69.37 3.667 69.375 4.278 ;
      RECT 69.365 3.682 69.37 4.293 ;
      RECT 69.35 3.712 69.365 4.32 ;
      RECT 69.345 3.742 69.35 4.346 ;
      RECT 69.34 3.76 69.345 4.358 ;
      RECT 69.33 3.79 69.34 4.377 ;
      RECT 69.32 3.815 69.33 4.402 ;
      RECT 69.315 3.835 69.32 4.421 ;
      RECT 69.31 3.852 69.315 4.434 ;
      RECT 69.3 3.878 69.31 4.453 ;
      RECT 69.29 3.916 69.3 4.48 ;
      RECT 69.285 3.942 69.29 4.5 ;
      RECT 69.28 3.952 69.285 4.51 ;
      RECT 69.275 3.965 69.28 4.525 ;
      RECT 69.27 3.98 69.275 4.535 ;
      RECT 69.265 4.002 69.27 4.55 ;
      RECT 69.26 4.02 69.265 4.561 ;
      RECT 69.255 4.03 69.26 4.572 ;
      RECT 69.25 4.038 69.255 4.584 ;
      RECT 69.245 4.046 69.25 4.595 ;
      RECT 69.24 4.072 69.245 4.608 ;
      RECT 69.23 4.1 69.24 4.621 ;
      RECT 69.225 4.13 69.23 4.63 ;
      RECT 69.22 4.145 69.225 4.637 ;
      RECT 69.205 4.17 69.22 4.644 ;
      RECT 69.2 4.192 69.205 4.65 ;
      RECT 69.195 4.217 69.2 4.653 ;
      RECT 69.186 4.245 69.195 4.657 ;
      RECT 69.18 4.262 69.186 4.662 ;
      RECT 69.175 4.28 69.18 4.666 ;
      RECT 69.17 4.292 69.175 4.669 ;
      RECT 69.165 4.313 69.17 4.673 ;
      RECT 69.16 4.331 69.165 4.676 ;
      RECT 69.155 4.345 69.16 4.679 ;
      RECT 69.15 4.362 69.155 4.682 ;
      RECT 69.145 4.375 69.15 4.685 ;
      RECT 69.12 4.412 69.145 4.693 ;
      RECT 69.115 4.457 69.12 4.702 ;
      RECT 69.11 4.485 69.115 4.705 ;
      RECT 69.1 4.505 69.11 4.709 ;
      RECT 69.095 4.525 69.1 4.714 ;
      RECT 69.09 4.54 69.095 4.717 ;
      RECT 69.07 4.55 69.09 4.724 ;
      RECT 69.005 4.557 69.07 4.75 ;
      RECT 68.97 4.56 69.005 4.778 ;
      RECT 68.955 4.563 68.97 4.793 ;
      RECT 68.945 4.564 68.955 4.808 ;
      RECT 68.935 4.565 68.945 4.825 ;
      RECT 68.93 4.565 68.935 4.84 ;
      RECT 68.925 4.565 68.93 4.848 ;
      RECT 68.91 4.566 68.925 4.863 ;
      RECT 68.88 4.568 68.91 4.87 ;
      RECT 68.77 4.575 68.85 4.87 ;
      RECT 68.725 4.58 68.77 4.87 ;
      RECT 68.715 4.581 68.725 4.86 ;
      RECT 68.705 4.582 68.715 4.853 ;
      RECT 68.685 4.584 68.705 4.848 ;
      RECT 68.675 4.555 68.685 4.843 ;
      RECT 68.63 4.555 68.675 4.835 ;
      RECT 68.6 4.555 68.625 4.825 ;
      RECT 68.58 4.555 68.6 4.818 ;
      RECT 68.86 3.355 69.12 3.615 ;
      RECT 68.74 3.37 68.75 3.535 ;
      RECT 68.725 3.37 68.73 3.53 ;
      RECT 66.09 3.21 66.275 3.5 ;
      RECT 67.905 3.335 67.92 3.49 ;
      RECT 66.055 3.21 66.08 3.47 ;
      RECT 68.47 3.26 68.475 3.402 ;
      RECT 68.385 3.255 68.41 3.395 ;
      RECT 68.785 3.372 68.86 3.565 ;
      RECT 68.77 3.37 68.785 3.548 ;
      RECT 68.75 3.37 68.77 3.54 ;
      RECT 68.73 3.37 68.74 3.533 ;
      RECT 68.685 3.365 68.725 3.523 ;
      RECT 68.645 3.34 68.685 3.508 ;
      RECT 68.63 3.315 68.645 3.498 ;
      RECT 68.625 3.309 68.63 3.496 ;
      RECT 68.59 3.301 68.625 3.479 ;
      RECT 68.585 3.294 68.59 3.467 ;
      RECT 68.565 3.289 68.585 3.455 ;
      RECT 68.555 3.283 68.565 3.44 ;
      RECT 68.535 3.278 68.555 3.425 ;
      RECT 68.525 3.273 68.535 3.418 ;
      RECT 68.52 3.271 68.525 3.413 ;
      RECT 68.515 3.27 68.52 3.41 ;
      RECT 68.475 3.265 68.515 3.406 ;
      RECT 68.455 3.259 68.47 3.401 ;
      RECT 68.42 3.256 68.455 3.398 ;
      RECT 68.41 3.255 68.42 3.396 ;
      RECT 68.35 3.255 68.385 3.393 ;
      RECT 68.305 3.255 68.35 3.393 ;
      RECT 68.255 3.255 68.305 3.396 ;
      RECT 68.24 3.257 68.255 3.398 ;
      RECT 68.225 3.26 68.24 3.399 ;
      RECT 68.215 3.265 68.225 3.4 ;
      RECT 68.185 3.27 68.215 3.405 ;
      RECT 68.175 3.276 68.185 3.413 ;
      RECT 68.165 3.278 68.175 3.417 ;
      RECT 68.155 3.282 68.165 3.421 ;
      RECT 68.13 3.288 68.155 3.429 ;
      RECT 68.12 3.293 68.13 3.437 ;
      RECT 68.105 3.297 68.12 3.441 ;
      RECT 68.07 3.303 68.105 3.449 ;
      RECT 68.05 3.308 68.07 3.459 ;
      RECT 68.02 3.315 68.05 3.468 ;
      RECT 67.975 3.324 68.02 3.482 ;
      RECT 67.97 3.329 67.975 3.493 ;
      RECT 67.95 3.332 67.97 3.494 ;
      RECT 67.92 3.335 67.95 3.492 ;
      RECT 67.885 3.335 67.905 3.488 ;
      RECT 67.815 3.335 67.885 3.479 ;
      RECT 67.8 3.332 67.815 3.471 ;
      RECT 67.76 3.325 67.8 3.466 ;
      RECT 67.735 3.315 67.76 3.459 ;
      RECT 67.73 3.309 67.735 3.456 ;
      RECT 67.69 3.303 67.73 3.453 ;
      RECT 67.675 3.296 67.69 3.448 ;
      RECT 67.655 3.292 67.675 3.443 ;
      RECT 67.64 3.287 67.655 3.439 ;
      RECT 67.625 3.282 67.64 3.437 ;
      RECT 67.61 3.278 67.625 3.436 ;
      RECT 67.595 3.276 67.61 3.432 ;
      RECT 67.585 3.274 67.595 3.427 ;
      RECT 67.57 3.271 67.585 3.423 ;
      RECT 67.56 3.269 67.57 3.418 ;
      RECT 67.54 3.266 67.56 3.414 ;
      RECT 67.495 3.265 67.54 3.412 ;
      RECT 67.435 3.267 67.495 3.413 ;
      RECT 67.415 3.269 67.435 3.415 ;
      RECT 67.385 3.272 67.415 3.416 ;
      RECT 67.335 3.277 67.385 3.418 ;
      RECT 67.33 3.28 67.335 3.42 ;
      RECT 67.32 3.282 67.33 3.423 ;
      RECT 67.315 3.284 67.32 3.426 ;
      RECT 67.265 3.287 67.315 3.433 ;
      RECT 67.245 3.291 67.265 3.445 ;
      RECT 67.235 3.294 67.245 3.451 ;
      RECT 67.225 3.295 67.235 3.454 ;
      RECT 67.186 3.298 67.225 3.456 ;
      RECT 67.1 3.305 67.186 3.459 ;
      RECT 67.026 3.315 67.1 3.463 ;
      RECT 66.94 3.326 67.026 3.468 ;
      RECT 66.925 3.333 66.94 3.47 ;
      RECT 66.87 3.337 66.925 3.471 ;
      RECT 66.856 3.34 66.87 3.473 ;
      RECT 66.77 3.34 66.856 3.475 ;
      RECT 66.73 3.337 66.77 3.478 ;
      RECT 66.706 3.333 66.73 3.48 ;
      RECT 66.62 3.323 66.706 3.483 ;
      RECT 66.59 3.312 66.62 3.484 ;
      RECT 66.571 3.308 66.59 3.483 ;
      RECT 66.485 3.301 66.571 3.48 ;
      RECT 66.425 3.29 66.485 3.477 ;
      RECT 66.405 3.282 66.425 3.475 ;
      RECT 66.37 3.277 66.405 3.474 ;
      RECT 66.345 3.272 66.37 3.473 ;
      RECT 66.315 3.267 66.345 3.472 ;
      RECT 66.29 3.21 66.315 3.471 ;
      RECT 66.275 3.21 66.29 3.495 ;
      RECT 66.08 3.21 66.09 3.495 ;
      RECT 67.855 4.23 67.86 4.37 ;
      RECT 67.515 4.23 67.55 4.368 ;
      RECT 67.09 4.215 67.105 4.36 ;
      RECT 68.92 3.995 69.01 4.255 ;
      RECT 68.75 3.86 68.85 4.255 ;
      RECT 65.785 3.835 65.865 4.045 ;
      RECT 68.875 3.972 68.92 4.255 ;
      RECT 68.865 3.942 68.875 4.255 ;
      RECT 68.85 3.865 68.865 4.255 ;
      RECT 68.665 3.86 68.75 4.22 ;
      RECT 68.66 3.862 68.665 4.215 ;
      RECT 68.655 3.867 68.66 4.215 ;
      RECT 68.62 3.967 68.655 4.215 ;
      RECT 68.61 3.995 68.62 4.215 ;
      RECT 68.6 4.01 68.61 4.215 ;
      RECT 68.59 4.022 68.6 4.215 ;
      RECT 68.585 4.032 68.59 4.215 ;
      RECT 68.57 4.042 68.585 4.217 ;
      RECT 68.565 4.057 68.57 4.219 ;
      RECT 68.55 4.07 68.565 4.221 ;
      RECT 68.545 4.085 68.55 4.224 ;
      RECT 68.525 4.095 68.545 4.228 ;
      RECT 68.51 4.105 68.525 4.231 ;
      RECT 68.475 4.112 68.51 4.236 ;
      RECT 68.431 4.119 68.475 4.244 ;
      RECT 68.345 4.131 68.431 4.257 ;
      RECT 68.32 4.142 68.345 4.268 ;
      RECT 68.29 4.147 68.32 4.273 ;
      RECT 68.255 4.152 68.29 4.281 ;
      RECT 68.225 4.157 68.255 4.288 ;
      RECT 68.2 4.162 68.225 4.293 ;
      RECT 68.135 4.169 68.2 4.302 ;
      RECT 68.065 4.182 68.135 4.318 ;
      RECT 68.035 4.192 68.065 4.33 ;
      RECT 68.01 4.197 68.035 4.337 ;
      RECT 67.955 4.204 68.01 4.345 ;
      RECT 67.95 4.211 67.955 4.35 ;
      RECT 67.945 4.213 67.95 4.351 ;
      RECT 67.93 4.215 67.945 4.353 ;
      RECT 67.925 4.215 67.93 4.356 ;
      RECT 67.86 4.222 67.925 4.363 ;
      RECT 67.825 4.232 67.855 4.373 ;
      RECT 67.808 4.235 67.825 4.375 ;
      RECT 67.722 4.234 67.808 4.374 ;
      RECT 67.636 4.232 67.722 4.371 ;
      RECT 67.55 4.231 67.636 4.369 ;
      RECT 67.449 4.229 67.515 4.368 ;
      RECT 67.363 4.226 67.449 4.366 ;
      RECT 67.277 4.222 67.363 4.364 ;
      RECT 67.191 4.219 67.277 4.363 ;
      RECT 67.105 4.216 67.191 4.361 ;
      RECT 67.005 4.215 67.09 4.358 ;
      RECT 66.955 4.213 67.005 4.356 ;
      RECT 66.935 4.21 66.955 4.354 ;
      RECT 66.915 4.208 66.935 4.351 ;
      RECT 66.89 4.204 66.915 4.348 ;
      RECT 66.845 4.198 66.89 4.343 ;
      RECT 66.805 4.192 66.845 4.335 ;
      RECT 66.78 4.187 66.805 4.328 ;
      RECT 66.725 4.18 66.78 4.32 ;
      RECT 66.701 4.173 66.725 4.313 ;
      RECT 66.615 4.164 66.701 4.303 ;
      RECT 66.585 4.156 66.615 4.293 ;
      RECT 66.555 4.152 66.585 4.288 ;
      RECT 66.55 4.149 66.555 4.285 ;
      RECT 66.545 4.148 66.55 4.285 ;
      RECT 66.47 4.141 66.545 4.278 ;
      RECT 66.431 4.132 66.47 4.267 ;
      RECT 66.345 4.122 66.431 4.255 ;
      RECT 66.305 4.112 66.345 4.243 ;
      RECT 66.266 4.107 66.305 4.236 ;
      RECT 66.18 4.097 66.266 4.225 ;
      RECT 66.14 4.085 66.18 4.214 ;
      RECT 66.105 4.07 66.14 4.207 ;
      RECT 66.095 4.06 66.105 4.204 ;
      RECT 66.075 4.045 66.095 4.202 ;
      RECT 66.045 4.015 66.075 4.198 ;
      RECT 66.035 3.995 66.045 4.193 ;
      RECT 66.03 3.987 66.035 4.19 ;
      RECT 66.025 3.98 66.03 4.188 ;
      RECT 66.01 3.967 66.025 4.181 ;
      RECT 66.005 3.957 66.01 4.173 ;
      RECT 66 3.95 66.005 4.168 ;
      RECT 65.995 3.945 66 4.164 ;
      RECT 65.98 3.932 65.995 4.156 ;
      RECT 65.975 3.842 65.98 4.145 ;
      RECT 65.97 3.837 65.975 4.138 ;
      RECT 65.895 3.835 65.97 4.098 ;
      RECT 65.865 3.835 65.895 4.053 ;
      RECT 65.77 3.84 65.785 4.04 ;
      RECT 68.255 3.545 68.515 3.805 ;
      RECT 68.24 3.533 68.42 3.77 ;
      RECT 68.235 3.534 68.42 3.768 ;
      RECT 68.22 3.538 68.43 3.758 ;
      RECT 68.215 3.543 68.435 3.728 ;
      RECT 68.22 3.54 68.435 3.758 ;
      RECT 68.235 3.535 68.43 3.768 ;
      RECT 68.255 3.532 68.42 3.805 ;
      RECT 68.255 3.531 68.41 3.805 ;
      RECT 68.28 3.53 68.41 3.805 ;
      RECT 67.84 3.775 68.1 4.035 ;
      RECT 67.715 3.82 68.1 4.03 ;
      RECT 67.705 3.825 68.1 4.025 ;
      RECT 67.72 4.765 67.735 5.075 ;
      RECT 66.315 4.535 66.325 4.665 ;
      RECT 66.095 4.53 66.2 4.665 ;
      RECT 66.01 4.535 66.06 4.665 ;
      RECT 64.56 3.27 64.565 4.375 ;
      RECT 67.815 4.857 67.82 4.993 ;
      RECT 67.81 4.852 67.815 5.053 ;
      RECT 67.805 4.85 67.81 5.066 ;
      RECT 67.79 4.847 67.805 5.068 ;
      RECT 67.785 4.842 67.79 5.07 ;
      RECT 67.78 4.838 67.785 5.073 ;
      RECT 67.765 4.833 67.78 5.075 ;
      RECT 67.735 4.825 67.765 5.075 ;
      RECT 67.696 4.765 67.72 5.075 ;
      RECT 67.61 4.765 67.696 5.072 ;
      RECT 67.58 4.765 67.61 5.065 ;
      RECT 67.555 4.765 67.58 5.058 ;
      RECT 67.53 4.765 67.555 5.05 ;
      RECT 67.515 4.765 67.53 5.043 ;
      RECT 67.49 4.765 67.515 5.035 ;
      RECT 67.475 4.765 67.49 5.028 ;
      RECT 67.435 4.775 67.475 5.017 ;
      RECT 67.425 4.77 67.435 5.007 ;
      RECT 67.421 4.769 67.425 5.004 ;
      RECT 67.335 4.761 67.421 4.987 ;
      RECT 67.302 4.75 67.335 4.964 ;
      RECT 67.216 4.739 67.302 4.942 ;
      RECT 67.13 4.723 67.216 4.911 ;
      RECT 67.06 4.708 67.13 4.883 ;
      RECT 67.05 4.701 67.06 4.87 ;
      RECT 67.02 4.698 67.05 4.86 ;
      RECT 66.995 4.694 67.02 4.853 ;
      RECT 66.98 4.691 66.995 4.848 ;
      RECT 66.975 4.69 66.98 4.843 ;
      RECT 66.945 4.685 66.975 4.836 ;
      RECT 66.94 4.68 66.945 4.831 ;
      RECT 66.925 4.677 66.94 4.826 ;
      RECT 66.92 4.672 66.925 4.821 ;
      RECT 66.9 4.667 66.92 4.818 ;
      RECT 66.885 4.662 66.9 4.81 ;
      RECT 66.87 4.656 66.885 4.805 ;
      RECT 66.84 4.647 66.87 4.798 ;
      RECT 66.835 4.64 66.84 4.79 ;
      RECT 66.83 4.638 66.835 4.788 ;
      RECT 66.825 4.637 66.83 4.785 ;
      RECT 66.785 4.63 66.825 4.778 ;
      RECT 66.771 4.62 66.785 4.768 ;
      RECT 66.72 4.609 66.771 4.756 ;
      RECT 66.695 4.595 66.72 4.742 ;
      RECT 66.67 4.584 66.695 4.734 ;
      RECT 66.65 4.573 66.67 4.728 ;
      RECT 66.64 4.567 66.65 4.723 ;
      RECT 66.635 4.565 66.64 4.719 ;
      RECT 66.615 4.56 66.635 4.714 ;
      RECT 66.585 4.55 66.615 4.704 ;
      RECT 66.58 4.542 66.585 4.697 ;
      RECT 66.565 4.54 66.58 4.693 ;
      RECT 66.545 4.54 66.565 4.688 ;
      RECT 66.54 4.539 66.545 4.686 ;
      RECT 66.535 4.539 66.54 4.683 ;
      RECT 66.495 4.538 66.535 4.678 ;
      RECT 66.47 4.537 66.495 4.673 ;
      RECT 66.41 4.536 66.47 4.67 ;
      RECT 66.325 4.535 66.41 4.668 ;
      RECT 66.286 4.534 66.315 4.665 ;
      RECT 66.2 4.532 66.286 4.665 ;
      RECT 66.06 4.532 66.095 4.665 ;
      RECT 65.97 4.536 66.01 4.668 ;
      RECT 65.955 4.539 65.97 4.675 ;
      RECT 65.945 4.54 65.955 4.682 ;
      RECT 65.92 4.543 65.945 4.687 ;
      RECT 65.915 4.545 65.92 4.69 ;
      RECT 65.865 4.547 65.915 4.691 ;
      RECT 65.826 4.551 65.865 4.693 ;
      RECT 65.74 4.553 65.826 4.696 ;
      RECT 65.722 4.555 65.74 4.698 ;
      RECT 65.636 4.558 65.722 4.7 ;
      RECT 65.55 4.562 65.636 4.703 ;
      RECT 65.513 4.566 65.55 4.706 ;
      RECT 65.427 4.569 65.513 4.709 ;
      RECT 65.341 4.573 65.427 4.712 ;
      RECT 65.255 4.578 65.341 4.716 ;
      RECT 65.235 4.58 65.255 4.719 ;
      RECT 65.215 4.579 65.235 4.72 ;
      RECT 65.166 4.576 65.215 4.721 ;
      RECT 65.08 4.571 65.166 4.724 ;
      RECT 65.03 4.566 65.08 4.726 ;
      RECT 65.006 4.564 65.03 4.727 ;
      RECT 64.92 4.559 65.006 4.729 ;
      RECT 64.895 4.555 64.92 4.728 ;
      RECT 64.885 4.552 64.895 4.726 ;
      RECT 64.875 4.545 64.885 4.723 ;
      RECT 64.87 4.525 64.875 4.718 ;
      RECT 64.86 4.495 64.87 4.713 ;
      RECT 64.845 4.365 64.86 4.704 ;
      RECT 64.84 4.357 64.845 4.697 ;
      RECT 64.82 4.35 64.84 4.689 ;
      RECT 64.815 4.332 64.82 4.681 ;
      RECT 64.805 4.312 64.815 4.676 ;
      RECT 64.8 4.285 64.805 4.672 ;
      RECT 64.795 4.262 64.8 4.669 ;
      RECT 64.775 4.22 64.795 4.661 ;
      RECT 64.74 4.135 64.775 4.645 ;
      RECT 64.735 4.067 64.74 4.633 ;
      RECT 64.72 4.037 64.735 4.627 ;
      RECT 64.715 3.282 64.72 3.528 ;
      RECT 64.705 4.007 64.72 4.618 ;
      RECT 64.71 3.277 64.715 3.56 ;
      RECT 64.705 3.272 64.71 3.603 ;
      RECT 64.7 3.27 64.705 3.638 ;
      RECT 64.685 3.97 64.705 4.608 ;
      RECT 64.695 3.27 64.7 3.675 ;
      RECT 64.68 3.27 64.695 3.773 ;
      RECT 64.68 3.943 64.685 4.601 ;
      RECT 64.675 3.27 64.68 3.848 ;
      RECT 64.675 3.931 64.68 4.598 ;
      RECT 64.67 3.27 64.675 3.88 ;
      RECT 64.67 3.91 64.675 4.595 ;
      RECT 64.665 3.27 64.67 4.592 ;
      RECT 64.63 3.27 64.665 4.578 ;
      RECT 64.615 3.27 64.63 4.56 ;
      RECT 64.595 3.27 64.615 4.55 ;
      RECT 64.57 3.27 64.595 4.533 ;
      RECT 64.565 3.27 64.57 4.483 ;
      RECT 64.555 3.27 64.56 4.313 ;
      RECT 64.55 3.27 64.555 4.22 ;
      RECT 64.545 3.27 64.55 4.133 ;
      RECT 64.54 3.27 64.545 4.065 ;
      RECT 64.535 3.27 64.54 4.008 ;
      RECT 64.525 3.27 64.535 3.903 ;
      RECT 64.52 3.27 64.525 3.775 ;
      RECT 64.515 3.27 64.52 3.693 ;
      RECT 64.51 3.272 64.515 3.61 ;
      RECT 64.505 3.277 64.51 3.543 ;
      RECT 64.5 3.282 64.505 3.47 ;
      RECT 67.315 3.6 67.575 3.86 ;
      RECT 67.335 3.567 67.545 3.86 ;
      RECT 67.335 3.565 67.535 3.86 ;
      RECT 67.345 3.552 67.535 3.86 ;
      RECT 67.345 3.55 67.46 3.86 ;
      RECT 66.82 3.675 66.995 3.955 ;
      RECT 66.815 3.675 66.995 3.953 ;
      RECT 66.815 3.675 67.01 3.95 ;
      RECT 66.805 3.675 67.01 3.948 ;
      RECT 66.75 3.675 67.01 3.935 ;
      RECT 66.75 3.75 67.015 3.913 ;
      RECT 66.28 4.873 66.285 5.08 ;
      RECT 66.23 4.867 66.28 5.079 ;
      RECT 66.197 4.881 66.29 5.078 ;
      RECT 66.111 4.881 66.29 5.077 ;
      RECT 66.025 4.881 66.29 5.076 ;
      RECT 66.025 4.98 66.295 5.073 ;
      RECT 66.02 4.98 66.295 5.068 ;
      RECT 66.015 4.98 66.295 5.05 ;
      RECT 66.01 4.98 66.295 5.033 ;
      RECT 65.97 4.765 66.23 5.025 ;
      RECT 65.43 3.915 65.516 4.329 ;
      RECT 65.43 3.915 65.555 4.326 ;
      RECT 65.43 3.915 65.575 4.316 ;
      RECT 65.385 3.915 65.575 4.313 ;
      RECT 65.385 4.067 65.585 4.303 ;
      RECT 65.385 4.088 65.59 4.297 ;
      RECT 65.385 4.106 65.595 4.293 ;
      RECT 65.385 4.126 65.605 4.288 ;
      RECT 65.36 4.126 65.605 4.285 ;
      RECT 65.35 4.126 65.605 4.263 ;
      RECT 65.35 4.142 65.61 4.233 ;
      RECT 65.315 3.915 65.575 4.22 ;
      RECT 65.315 4.154 65.615 4.175 ;
      RECT 62.975 10.06 63.27 10.29 ;
      RECT 63.035 8.58 63.205 10.29 ;
      RECT 62.985 8.95 63.335 9.3 ;
      RECT 62.975 8.58 63.265 8.81 ;
      RECT 61.985 10.06 62.28 10.29 ;
      RECT 62.045 8.58 62.215 10.29 ;
      RECT 61.985 8.58 62.275 8.81 ;
      RECT 61.985 8.615 62.835 8.775 ;
      RECT 62.67 8.21 62.835 8.775 ;
      RECT 61.985 8.61 62.38 8.775 ;
      RECT 62.605 8.21 62.895 8.44 ;
      RECT 62.605 8.24 63.065 8.41 ;
      RECT 62.57 4.005 62.89 4.26 ;
      RECT 62.57 4.055 63.06 4.225 ;
      RECT 62.57 3.69 62.76 4.26 ;
      RECT 61.985 3.655 62.275 3.885 ;
      RECT 61.985 3.69 62.76 3.86 ;
      RECT 62.045 2.175 62.215 3.885 ;
      RECT 61.985 2.175 62.28 2.405 ;
      RECT 61.615 4.025 61.905 4.255 ;
      RECT 61.615 4.055 62.075 4.225 ;
      RECT 61.68 2.95 61.845 4.255 ;
      RECT 60.195 2.915 60.485 3.145 ;
      RECT 60.195 2.95 61.845 3.12 ;
      RECT 60.255 2.175 60.425 3.145 ;
      RECT 60.195 2.175 60.485 2.405 ;
      RECT 60.195 10.06 60.485 10.29 ;
      RECT 60.255 9.32 60.425 10.29 ;
      RECT 60.255 9.41 61.845 9.58 ;
      RECT 61.675 8.21 61.845 9.58 ;
      RECT 60.195 9.32 60.485 9.55 ;
      RECT 61.615 8.21 61.905 8.44 ;
      RECT 61.615 8.24 62.075 8.41 ;
      RECT 58.245 4 58.585 4.35 ;
      RECT 58.335 3.32 58.505 4.35 ;
      RECT 60.625 3.26 60.975 3.61 ;
      RECT 58.335 3.32 60.975 3.49 ;
      RECT 60.455 3.315 60.975 3.49 ;
      RECT 60.65 8.945 60.975 9.27 ;
      RECT 55.19 8.905 55.54 9.255 ;
      RECT 60.625 8.95 60.975 9.18 ;
      RECT 54.99 8.95 55.54 9.18 ;
      RECT 60.455 8.975 60.975 9.15 ;
      RECT 54.82 8.98 55.54 9.15 ;
      RECT 54.87 8.975 60.975 9.145 ;
      RECT 59.85 3.66 60.17 3.98 ;
      RECT 59.825 3.655 60.115 3.885 ;
      RECT 59.82 3.685 60.17 3.86 ;
      RECT 59.65 3.685 60.17 3.855 ;
      RECT 59.85 8.545 60.17 8.835 ;
      RECT 59.825 8.58 60.17 8.81 ;
      RECT 59.65 8.61 60.17 8.78 ;
      RECT 55.54 4.28 55.69 4.555 ;
      RECT 56.08 3.36 56.085 3.58 ;
      RECT 57.23 3.56 57.245 3.758 ;
      RECT 57.195 3.552 57.23 3.765 ;
      RECT 57.165 3.545 57.195 3.765 ;
      RECT 57.11 3.51 57.165 3.765 ;
      RECT 57.045 3.447 57.11 3.765 ;
      RECT 57.04 3.412 57.045 3.763 ;
      RECT 57.035 3.407 57.04 3.755 ;
      RECT 57.03 3.402 57.035 3.741 ;
      RECT 57.025 3.399 57.03 3.734 ;
      RECT 56.98 3.389 57.025 3.685 ;
      RECT 56.96 3.376 56.98 3.62 ;
      RECT 56.955 3.371 56.96 3.593 ;
      RECT 56.95 3.37 56.955 3.586 ;
      RECT 56.945 3.369 56.95 3.579 ;
      RECT 56.86 3.354 56.945 3.525 ;
      RECT 56.83 3.335 56.86 3.475 ;
      RECT 56.75 3.318 56.83 3.46 ;
      RECT 56.715 3.305 56.75 3.445 ;
      RECT 56.707 3.305 56.715 3.44 ;
      RECT 56.621 3.306 56.707 3.44 ;
      RECT 56.535 3.308 56.621 3.44 ;
      RECT 56.51 3.309 56.535 3.444 ;
      RECT 56.435 3.315 56.51 3.459 ;
      RECT 56.352 3.327 56.435 3.483 ;
      RECT 56.266 3.34 56.352 3.509 ;
      RECT 56.18 3.353 56.266 3.535 ;
      RECT 56.145 3.362 56.18 3.554 ;
      RECT 56.095 3.362 56.145 3.567 ;
      RECT 56.085 3.36 56.095 3.578 ;
      RECT 56.07 3.357 56.08 3.58 ;
      RECT 56.055 3.349 56.07 3.588 ;
      RECT 56.04 3.341 56.055 3.608 ;
      RECT 56.035 3.336 56.04 3.665 ;
      RECT 56.02 3.331 56.035 3.738 ;
      RECT 56.015 3.326 56.02 3.78 ;
      RECT 56.01 3.324 56.015 3.808 ;
      RECT 56.005 3.322 56.01 3.83 ;
      RECT 55.995 3.318 56.005 3.873 ;
      RECT 55.99 3.315 55.995 3.898 ;
      RECT 55.985 3.313 55.99 3.918 ;
      RECT 55.98 3.311 55.985 3.942 ;
      RECT 55.975 3.307 55.98 3.965 ;
      RECT 55.97 3.303 55.975 3.988 ;
      RECT 55.935 3.293 55.97 4.095 ;
      RECT 55.93 3.283 55.935 4.193 ;
      RECT 55.925 3.281 55.93 4.22 ;
      RECT 55.92 3.28 55.925 4.24 ;
      RECT 55.915 3.272 55.92 4.26 ;
      RECT 55.91 3.267 55.915 4.295 ;
      RECT 55.905 3.265 55.91 4.313 ;
      RECT 55.9 3.265 55.905 4.338 ;
      RECT 55.895 3.265 55.9 4.36 ;
      RECT 55.86 3.265 55.895 4.403 ;
      RECT 55.835 3.265 55.86 4.432 ;
      RECT 55.825 3.265 55.835 3.618 ;
      RECT 55.828 3.675 55.835 4.442 ;
      RECT 55.825 3.732 55.828 4.445 ;
      RECT 55.82 3.265 55.825 3.59 ;
      RECT 55.82 3.782 55.825 4.448 ;
      RECT 55.81 3.265 55.82 3.58 ;
      RECT 55.815 3.835 55.82 4.451 ;
      RECT 55.81 3.92 55.815 4.455 ;
      RECT 55.8 3.265 55.81 3.568 ;
      RECT 55.805 3.967 55.81 4.459 ;
      RECT 55.8 4.042 55.805 4.463 ;
      RECT 55.765 3.265 55.8 3.543 ;
      RECT 55.79 4.125 55.8 4.468 ;
      RECT 55.78 4.192 55.79 4.475 ;
      RECT 55.775 4.22 55.78 4.48 ;
      RECT 55.765 4.233 55.775 4.486 ;
      RECT 55.72 3.265 55.765 3.5 ;
      RECT 55.76 4.238 55.765 4.493 ;
      RECT 55.72 4.255 55.76 4.555 ;
      RECT 55.715 3.267 55.72 3.473 ;
      RECT 55.69 4.275 55.72 4.555 ;
      RECT 55.71 3.272 55.715 3.445 ;
      RECT 55.5 4.284 55.54 4.555 ;
      RECT 55.475 4.292 55.5 4.525 ;
      RECT 55.43 4.3 55.475 4.525 ;
      RECT 55.415 4.305 55.43 4.52 ;
      RECT 55.405 4.305 55.415 4.514 ;
      RECT 55.395 4.312 55.405 4.511 ;
      RECT 55.39 4.35 55.395 4.5 ;
      RECT 55.385 4.412 55.39 4.478 ;
      RECT 56.655 4.287 56.84 4.51 ;
      RECT 56.655 4.302 56.845 4.506 ;
      RECT 56.645 3.575 56.73 4.505 ;
      RECT 56.645 4.302 56.85 4.499 ;
      RECT 56.64 4.31 56.85 4.498 ;
      RECT 56.845 4.03 57.165 4.35 ;
      RECT 56.64 4.202 56.81 4.293 ;
      RECT 56.635 4.202 56.81 4.275 ;
      RECT 56.625 4.01 56.76 4.25 ;
      RECT 56.62 4.01 56.76 4.195 ;
      RECT 56.58 3.59 56.75 4.095 ;
      RECT 56.565 3.59 56.75 3.965 ;
      RECT 56.56 3.59 56.75 3.918 ;
      RECT 56.555 3.59 56.75 3.898 ;
      RECT 56.55 3.59 56.75 3.873 ;
      RECT 56.52 3.59 56.78 3.85 ;
      RECT 56.53 3.587 56.74 3.85 ;
      RECT 56.655 3.582 56.74 4.51 ;
      RECT 56.54 3.575 56.73 3.85 ;
      RECT 56.535 3.58 56.73 3.85 ;
      RECT 55.365 3.792 55.55 4.005 ;
      RECT 55.365 3.8 55.56 3.998 ;
      RECT 55.345 3.8 55.56 3.995 ;
      RECT 55.34 3.8 55.56 3.98 ;
      RECT 55.27 3.715 55.53 3.975 ;
      RECT 55.27 3.86 55.565 3.888 ;
      RECT 54.925 4.315 55.185 4.575 ;
      RECT 54.95 4.26 55.145 4.575 ;
      RECT 54.945 4.009 55.125 4.303 ;
      RECT 54.945 4.015 55.135 4.303 ;
      RECT 54.925 4.017 55.135 4.248 ;
      RECT 54.92 4.027 55.135 4.115 ;
      RECT 54.95 4.007 55.125 4.575 ;
      RECT 55.036 4.005 55.125 4.575 ;
      RECT 54.895 3.225 54.93 3.595 ;
      RECT 54.685 3.335 54.69 3.595 ;
      RECT 54.93 3.232 54.945 3.595 ;
      RECT 54.82 3.225 54.895 3.673 ;
      RECT 54.81 3.225 54.82 3.758 ;
      RECT 54.785 3.225 54.81 3.793 ;
      RECT 54.745 3.225 54.785 3.861 ;
      RECT 54.735 3.232 54.745 3.913 ;
      RECT 54.705 3.335 54.735 3.954 ;
      RECT 54.7 3.335 54.705 3.993 ;
      RECT 54.69 3.335 54.7 4.013 ;
      RECT 54.685 3.63 54.69 4.05 ;
      RECT 54.68 3.647 54.685 4.07 ;
      RECT 54.665 3.71 54.68 4.11 ;
      RECT 54.66 3.753 54.665 4.145 ;
      RECT 54.655 3.761 54.66 4.158 ;
      RECT 54.645 3.775 54.655 4.18 ;
      RECT 54.62 3.81 54.645 4.245 ;
      RECT 54.61 3.845 54.62 4.308 ;
      RECT 54.59 3.875 54.61 4.369 ;
      RECT 54.575 3.911 54.59 4.436 ;
      RECT 54.565 3.939 54.575 4.475 ;
      RECT 54.555 3.961 54.565 4.495 ;
      RECT 54.55 3.971 54.555 4.506 ;
      RECT 54.545 3.98 54.55 4.509 ;
      RECT 54.535 3.998 54.545 4.513 ;
      RECT 54.525 4.016 54.535 4.514 ;
      RECT 54.5 4.055 54.525 4.511 ;
      RECT 54.48 4.097 54.5 4.508 ;
      RECT 54.465 4.135 54.48 4.507 ;
      RECT 54.43 4.17 54.465 4.504 ;
      RECT 54.425 4.192 54.43 4.502 ;
      RECT 54.36 4.232 54.425 4.499 ;
      RECT 54.355 4.272 54.36 4.495 ;
      RECT 54.34 4.282 54.355 4.486 ;
      RECT 54.33 4.402 54.34 4.471 ;
      RECT 54.81 4.815 54.82 5.075 ;
      RECT 54.81 4.818 54.83 5.074 ;
      RECT 54.8 4.808 54.81 5.073 ;
      RECT 54.79 4.823 54.87 5.069 ;
      RECT 54.775 4.802 54.79 5.067 ;
      RECT 54.75 4.827 54.875 5.063 ;
      RECT 54.735 4.787 54.75 5.058 ;
      RECT 54.735 4.829 54.885 5.057 ;
      RECT 54.735 4.837 54.9 5.05 ;
      RECT 54.675 4.774 54.735 5.04 ;
      RECT 54.665 4.761 54.675 5.022 ;
      RECT 54.64 4.751 54.665 5.012 ;
      RECT 54.635 4.741 54.64 5.004 ;
      RECT 54.57 4.837 54.9 4.986 ;
      RECT 54.485 4.837 54.9 4.948 ;
      RECT 54.375 4.665 54.635 4.925 ;
      RECT 54.75 4.795 54.775 5.063 ;
      RECT 54.79 4.805 54.8 5.069 ;
      RECT 54.375 4.813 54.815 4.925 ;
      RECT 54.56 10.06 54.85 10.29 ;
      RECT 54.62 9.32 54.79 10.29 ;
      RECT 54.52 9.345 54.89 9.715 ;
      RECT 54.56 9.32 54.85 9.715 ;
      RECT 53.59 4.57 53.62 4.87 ;
      RECT 53.365 4.555 53.37 4.83 ;
      RECT 53.165 4.555 53.32 4.815 ;
      RECT 54.465 3.27 54.495 3.53 ;
      RECT 54.455 3.27 54.465 3.638 ;
      RECT 54.435 3.27 54.455 3.648 ;
      RECT 54.42 3.27 54.435 3.66 ;
      RECT 54.365 3.27 54.42 3.71 ;
      RECT 54.35 3.27 54.365 3.758 ;
      RECT 54.32 3.27 54.35 3.793 ;
      RECT 54.265 3.27 54.32 3.855 ;
      RECT 54.245 3.27 54.265 3.923 ;
      RECT 54.24 3.27 54.245 3.953 ;
      RECT 54.235 3.27 54.24 3.965 ;
      RECT 54.23 3.387 54.235 3.983 ;
      RECT 54.21 3.405 54.23 4.008 ;
      RECT 54.19 3.432 54.21 4.058 ;
      RECT 54.185 3.452 54.19 4.089 ;
      RECT 54.18 3.46 54.185 4.106 ;
      RECT 54.165 3.486 54.18 4.135 ;
      RECT 54.15 3.528 54.165 4.17 ;
      RECT 54.145 3.557 54.15 4.193 ;
      RECT 54.14 3.572 54.145 4.206 ;
      RECT 54.135 3.595 54.14 4.217 ;
      RECT 54.125 3.615 54.135 4.235 ;
      RECT 54.115 3.645 54.125 4.258 ;
      RECT 54.11 3.667 54.115 4.278 ;
      RECT 54.105 3.682 54.11 4.293 ;
      RECT 54.09 3.712 54.105 4.32 ;
      RECT 54.085 3.742 54.09 4.346 ;
      RECT 54.08 3.76 54.085 4.358 ;
      RECT 54.07 3.79 54.08 4.377 ;
      RECT 54.06 3.815 54.07 4.402 ;
      RECT 54.055 3.835 54.06 4.421 ;
      RECT 54.05 3.852 54.055 4.434 ;
      RECT 54.04 3.878 54.05 4.453 ;
      RECT 54.03 3.916 54.04 4.48 ;
      RECT 54.025 3.942 54.03 4.5 ;
      RECT 54.02 3.952 54.025 4.51 ;
      RECT 54.015 3.965 54.02 4.525 ;
      RECT 54.01 3.98 54.015 4.535 ;
      RECT 54.005 4.002 54.01 4.55 ;
      RECT 54 4.02 54.005 4.561 ;
      RECT 53.995 4.03 54 4.572 ;
      RECT 53.99 4.038 53.995 4.584 ;
      RECT 53.985 4.046 53.99 4.595 ;
      RECT 53.98 4.072 53.985 4.608 ;
      RECT 53.97 4.1 53.98 4.621 ;
      RECT 53.965 4.13 53.97 4.63 ;
      RECT 53.96 4.145 53.965 4.637 ;
      RECT 53.945 4.17 53.96 4.644 ;
      RECT 53.94 4.192 53.945 4.65 ;
      RECT 53.935 4.217 53.94 4.653 ;
      RECT 53.926 4.245 53.935 4.657 ;
      RECT 53.92 4.262 53.926 4.662 ;
      RECT 53.915 4.28 53.92 4.666 ;
      RECT 53.91 4.292 53.915 4.669 ;
      RECT 53.905 4.313 53.91 4.673 ;
      RECT 53.9 4.331 53.905 4.676 ;
      RECT 53.895 4.345 53.9 4.679 ;
      RECT 53.89 4.362 53.895 4.682 ;
      RECT 53.885 4.375 53.89 4.685 ;
      RECT 53.86 4.412 53.885 4.693 ;
      RECT 53.855 4.457 53.86 4.702 ;
      RECT 53.85 4.485 53.855 4.705 ;
      RECT 53.84 4.505 53.85 4.709 ;
      RECT 53.835 4.525 53.84 4.714 ;
      RECT 53.83 4.54 53.835 4.717 ;
      RECT 53.81 4.55 53.83 4.724 ;
      RECT 53.745 4.557 53.81 4.75 ;
      RECT 53.71 4.56 53.745 4.778 ;
      RECT 53.695 4.563 53.71 4.793 ;
      RECT 53.685 4.564 53.695 4.808 ;
      RECT 53.675 4.565 53.685 4.825 ;
      RECT 53.67 4.565 53.675 4.84 ;
      RECT 53.665 4.565 53.67 4.848 ;
      RECT 53.65 4.566 53.665 4.863 ;
      RECT 53.62 4.568 53.65 4.87 ;
      RECT 53.51 4.575 53.59 4.87 ;
      RECT 53.465 4.58 53.51 4.87 ;
      RECT 53.455 4.581 53.465 4.86 ;
      RECT 53.445 4.582 53.455 4.853 ;
      RECT 53.425 4.584 53.445 4.848 ;
      RECT 53.415 4.555 53.425 4.843 ;
      RECT 53.37 4.555 53.415 4.835 ;
      RECT 53.34 4.555 53.365 4.825 ;
      RECT 53.32 4.555 53.34 4.818 ;
      RECT 53.6 3.355 53.86 3.615 ;
      RECT 53.48 3.37 53.49 3.535 ;
      RECT 53.465 3.37 53.47 3.53 ;
      RECT 50.83 3.21 51.015 3.5 ;
      RECT 52.645 3.335 52.66 3.49 ;
      RECT 50.795 3.21 50.82 3.47 ;
      RECT 53.21 3.26 53.215 3.402 ;
      RECT 53.125 3.255 53.15 3.395 ;
      RECT 53.525 3.372 53.6 3.565 ;
      RECT 53.51 3.37 53.525 3.548 ;
      RECT 53.49 3.37 53.51 3.54 ;
      RECT 53.47 3.37 53.48 3.533 ;
      RECT 53.425 3.365 53.465 3.523 ;
      RECT 53.385 3.34 53.425 3.508 ;
      RECT 53.37 3.315 53.385 3.498 ;
      RECT 53.365 3.309 53.37 3.496 ;
      RECT 53.33 3.301 53.365 3.479 ;
      RECT 53.325 3.294 53.33 3.467 ;
      RECT 53.305 3.289 53.325 3.455 ;
      RECT 53.295 3.283 53.305 3.44 ;
      RECT 53.275 3.278 53.295 3.425 ;
      RECT 53.265 3.273 53.275 3.418 ;
      RECT 53.26 3.271 53.265 3.413 ;
      RECT 53.255 3.27 53.26 3.41 ;
      RECT 53.215 3.265 53.255 3.406 ;
      RECT 53.195 3.259 53.21 3.401 ;
      RECT 53.16 3.256 53.195 3.398 ;
      RECT 53.15 3.255 53.16 3.396 ;
      RECT 53.09 3.255 53.125 3.393 ;
      RECT 53.045 3.255 53.09 3.393 ;
      RECT 52.995 3.255 53.045 3.396 ;
      RECT 52.98 3.257 52.995 3.398 ;
      RECT 52.965 3.26 52.98 3.399 ;
      RECT 52.955 3.265 52.965 3.4 ;
      RECT 52.925 3.27 52.955 3.405 ;
      RECT 52.915 3.276 52.925 3.413 ;
      RECT 52.905 3.278 52.915 3.417 ;
      RECT 52.895 3.282 52.905 3.421 ;
      RECT 52.87 3.288 52.895 3.429 ;
      RECT 52.86 3.293 52.87 3.437 ;
      RECT 52.845 3.297 52.86 3.441 ;
      RECT 52.81 3.303 52.845 3.449 ;
      RECT 52.79 3.308 52.81 3.459 ;
      RECT 52.76 3.315 52.79 3.468 ;
      RECT 52.715 3.324 52.76 3.482 ;
      RECT 52.71 3.329 52.715 3.493 ;
      RECT 52.69 3.332 52.71 3.494 ;
      RECT 52.66 3.335 52.69 3.492 ;
      RECT 52.625 3.335 52.645 3.488 ;
      RECT 52.555 3.335 52.625 3.479 ;
      RECT 52.54 3.332 52.555 3.471 ;
      RECT 52.5 3.325 52.54 3.466 ;
      RECT 52.475 3.315 52.5 3.459 ;
      RECT 52.47 3.309 52.475 3.456 ;
      RECT 52.43 3.303 52.47 3.453 ;
      RECT 52.415 3.296 52.43 3.448 ;
      RECT 52.395 3.292 52.415 3.443 ;
      RECT 52.38 3.287 52.395 3.439 ;
      RECT 52.365 3.282 52.38 3.437 ;
      RECT 52.35 3.278 52.365 3.436 ;
      RECT 52.335 3.276 52.35 3.432 ;
      RECT 52.325 3.274 52.335 3.427 ;
      RECT 52.31 3.271 52.325 3.423 ;
      RECT 52.3 3.269 52.31 3.418 ;
      RECT 52.28 3.266 52.3 3.414 ;
      RECT 52.235 3.265 52.28 3.412 ;
      RECT 52.175 3.267 52.235 3.413 ;
      RECT 52.155 3.269 52.175 3.415 ;
      RECT 52.125 3.272 52.155 3.416 ;
      RECT 52.075 3.277 52.125 3.418 ;
      RECT 52.07 3.28 52.075 3.42 ;
      RECT 52.06 3.282 52.07 3.423 ;
      RECT 52.055 3.284 52.06 3.426 ;
      RECT 52.005 3.287 52.055 3.433 ;
      RECT 51.985 3.291 52.005 3.445 ;
      RECT 51.975 3.294 51.985 3.451 ;
      RECT 51.965 3.295 51.975 3.454 ;
      RECT 51.926 3.298 51.965 3.456 ;
      RECT 51.84 3.305 51.926 3.459 ;
      RECT 51.766 3.315 51.84 3.463 ;
      RECT 51.68 3.326 51.766 3.468 ;
      RECT 51.665 3.333 51.68 3.47 ;
      RECT 51.61 3.337 51.665 3.471 ;
      RECT 51.596 3.34 51.61 3.473 ;
      RECT 51.51 3.34 51.596 3.475 ;
      RECT 51.47 3.337 51.51 3.478 ;
      RECT 51.446 3.333 51.47 3.48 ;
      RECT 51.36 3.323 51.446 3.483 ;
      RECT 51.33 3.312 51.36 3.484 ;
      RECT 51.311 3.308 51.33 3.483 ;
      RECT 51.225 3.301 51.311 3.48 ;
      RECT 51.165 3.29 51.225 3.477 ;
      RECT 51.145 3.282 51.165 3.475 ;
      RECT 51.11 3.277 51.145 3.474 ;
      RECT 51.085 3.272 51.11 3.473 ;
      RECT 51.055 3.267 51.085 3.472 ;
      RECT 51.03 3.21 51.055 3.471 ;
      RECT 51.015 3.21 51.03 3.495 ;
      RECT 50.82 3.21 50.83 3.495 ;
      RECT 52.595 4.23 52.6 4.37 ;
      RECT 52.255 4.23 52.29 4.368 ;
      RECT 51.83 4.215 51.845 4.36 ;
      RECT 53.66 3.995 53.75 4.255 ;
      RECT 53.49 3.86 53.59 4.255 ;
      RECT 50.525 3.835 50.605 4.045 ;
      RECT 53.615 3.972 53.66 4.255 ;
      RECT 53.605 3.942 53.615 4.255 ;
      RECT 53.59 3.865 53.605 4.255 ;
      RECT 53.405 3.86 53.49 4.22 ;
      RECT 53.4 3.862 53.405 4.215 ;
      RECT 53.395 3.867 53.4 4.215 ;
      RECT 53.36 3.967 53.395 4.215 ;
      RECT 53.35 3.995 53.36 4.215 ;
      RECT 53.34 4.01 53.35 4.215 ;
      RECT 53.33 4.022 53.34 4.215 ;
      RECT 53.325 4.032 53.33 4.215 ;
      RECT 53.31 4.042 53.325 4.217 ;
      RECT 53.305 4.057 53.31 4.219 ;
      RECT 53.29 4.07 53.305 4.221 ;
      RECT 53.285 4.085 53.29 4.224 ;
      RECT 53.265 4.095 53.285 4.228 ;
      RECT 53.25 4.105 53.265 4.231 ;
      RECT 53.215 4.112 53.25 4.236 ;
      RECT 53.171 4.119 53.215 4.244 ;
      RECT 53.085 4.131 53.171 4.257 ;
      RECT 53.06 4.142 53.085 4.268 ;
      RECT 53.03 4.147 53.06 4.273 ;
      RECT 52.995 4.152 53.03 4.281 ;
      RECT 52.965 4.157 52.995 4.288 ;
      RECT 52.94 4.162 52.965 4.293 ;
      RECT 52.875 4.169 52.94 4.302 ;
      RECT 52.805 4.182 52.875 4.318 ;
      RECT 52.775 4.192 52.805 4.33 ;
      RECT 52.75 4.197 52.775 4.337 ;
      RECT 52.695 4.204 52.75 4.345 ;
      RECT 52.69 4.211 52.695 4.35 ;
      RECT 52.685 4.213 52.69 4.351 ;
      RECT 52.67 4.215 52.685 4.353 ;
      RECT 52.665 4.215 52.67 4.356 ;
      RECT 52.6 4.222 52.665 4.363 ;
      RECT 52.565 4.232 52.595 4.373 ;
      RECT 52.548 4.235 52.565 4.375 ;
      RECT 52.462 4.234 52.548 4.374 ;
      RECT 52.376 4.232 52.462 4.371 ;
      RECT 52.29 4.231 52.376 4.369 ;
      RECT 52.189 4.229 52.255 4.368 ;
      RECT 52.103 4.226 52.189 4.366 ;
      RECT 52.017 4.222 52.103 4.364 ;
      RECT 51.931 4.219 52.017 4.363 ;
      RECT 51.845 4.216 51.931 4.361 ;
      RECT 51.745 4.215 51.83 4.358 ;
      RECT 51.695 4.213 51.745 4.356 ;
      RECT 51.675 4.21 51.695 4.354 ;
      RECT 51.655 4.208 51.675 4.351 ;
      RECT 51.63 4.204 51.655 4.348 ;
      RECT 51.585 4.198 51.63 4.343 ;
      RECT 51.545 4.192 51.585 4.335 ;
      RECT 51.52 4.187 51.545 4.328 ;
      RECT 51.465 4.18 51.52 4.32 ;
      RECT 51.441 4.173 51.465 4.313 ;
      RECT 51.355 4.164 51.441 4.303 ;
      RECT 51.325 4.156 51.355 4.293 ;
      RECT 51.295 4.152 51.325 4.288 ;
      RECT 51.29 4.149 51.295 4.285 ;
      RECT 51.285 4.148 51.29 4.285 ;
      RECT 51.21 4.141 51.285 4.278 ;
      RECT 51.171 4.132 51.21 4.267 ;
      RECT 51.085 4.122 51.171 4.255 ;
      RECT 51.045 4.112 51.085 4.243 ;
      RECT 51.006 4.107 51.045 4.236 ;
      RECT 50.92 4.097 51.006 4.225 ;
      RECT 50.88 4.085 50.92 4.214 ;
      RECT 50.845 4.07 50.88 4.207 ;
      RECT 50.835 4.06 50.845 4.204 ;
      RECT 50.815 4.045 50.835 4.202 ;
      RECT 50.785 4.015 50.815 4.198 ;
      RECT 50.775 3.995 50.785 4.193 ;
      RECT 50.77 3.987 50.775 4.19 ;
      RECT 50.765 3.98 50.77 4.188 ;
      RECT 50.75 3.967 50.765 4.181 ;
      RECT 50.745 3.957 50.75 4.173 ;
      RECT 50.74 3.95 50.745 4.168 ;
      RECT 50.735 3.945 50.74 4.164 ;
      RECT 50.72 3.932 50.735 4.156 ;
      RECT 50.715 3.842 50.72 4.145 ;
      RECT 50.71 3.837 50.715 4.138 ;
      RECT 50.635 3.835 50.71 4.098 ;
      RECT 50.605 3.835 50.635 4.053 ;
      RECT 50.51 3.84 50.525 4.04 ;
      RECT 52.995 3.545 53.255 3.805 ;
      RECT 52.98 3.533 53.16 3.77 ;
      RECT 52.975 3.534 53.16 3.768 ;
      RECT 52.96 3.538 53.17 3.758 ;
      RECT 52.955 3.543 53.175 3.728 ;
      RECT 52.96 3.54 53.175 3.758 ;
      RECT 52.975 3.535 53.17 3.768 ;
      RECT 52.995 3.532 53.16 3.805 ;
      RECT 52.995 3.531 53.15 3.805 ;
      RECT 53.02 3.53 53.15 3.805 ;
      RECT 52.58 3.775 52.84 4.035 ;
      RECT 52.455 3.82 52.84 4.03 ;
      RECT 52.445 3.825 52.84 4.025 ;
      RECT 52.46 4.765 52.475 5.075 ;
      RECT 51.055 4.535 51.065 4.665 ;
      RECT 50.835 4.53 50.94 4.665 ;
      RECT 50.75 4.535 50.8 4.665 ;
      RECT 49.3 3.27 49.305 4.375 ;
      RECT 52.555 4.857 52.56 4.993 ;
      RECT 52.55 4.852 52.555 5.053 ;
      RECT 52.545 4.85 52.55 5.066 ;
      RECT 52.53 4.847 52.545 5.068 ;
      RECT 52.525 4.842 52.53 5.07 ;
      RECT 52.52 4.838 52.525 5.073 ;
      RECT 52.505 4.833 52.52 5.075 ;
      RECT 52.475 4.825 52.505 5.075 ;
      RECT 52.436 4.765 52.46 5.075 ;
      RECT 52.35 4.765 52.436 5.072 ;
      RECT 52.32 4.765 52.35 5.065 ;
      RECT 52.295 4.765 52.32 5.058 ;
      RECT 52.27 4.765 52.295 5.05 ;
      RECT 52.255 4.765 52.27 5.043 ;
      RECT 52.23 4.765 52.255 5.035 ;
      RECT 52.215 4.765 52.23 5.028 ;
      RECT 52.175 4.775 52.215 5.017 ;
      RECT 52.165 4.77 52.175 5.007 ;
      RECT 52.161 4.769 52.165 5.004 ;
      RECT 52.075 4.761 52.161 4.987 ;
      RECT 52.042 4.75 52.075 4.964 ;
      RECT 51.956 4.739 52.042 4.942 ;
      RECT 51.87 4.723 51.956 4.911 ;
      RECT 51.8 4.708 51.87 4.883 ;
      RECT 51.79 4.701 51.8 4.87 ;
      RECT 51.76 4.698 51.79 4.86 ;
      RECT 51.735 4.694 51.76 4.853 ;
      RECT 51.72 4.691 51.735 4.848 ;
      RECT 51.715 4.69 51.72 4.843 ;
      RECT 51.685 4.685 51.715 4.836 ;
      RECT 51.68 4.68 51.685 4.831 ;
      RECT 51.665 4.677 51.68 4.826 ;
      RECT 51.66 4.672 51.665 4.821 ;
      RECT 51.64 4.667 51.66 4.818 ;
      RECT 51.625 4.662 51.64 4.81 ;
      RECT 51.61 4.656 51.625 4.805 ;
      RECT 51.58 4.647 51.61 4.798 ;
      RECT 51.575 4.64 51.58 4.79 ;
      RECT 51.57 4.638 51.575 4.788 ;
      RECT 51.565 4.637 51.57 4.785 ;
      RECT 51.525 4.63 51.565 4.778 ;
      RECT 51.511 4.62 51.525 4.768 ;
      RECT 51.46 4.609 51.511 4.756 ;
      RECT 51.435 4.595 51.46 4.742 ;
      RECT 51.41 4.584 51.435 4.734 ;
      RECT 51.39 4.573 51.41 4.728 ;
      RECT 51.38 4.567 51.39 4.723 ;
      RECT 51.375 4.565 51.38 4.719 ;
      RECT 51.355 4.56 51.375 4.714 ;
      RECT 51.325 4.55 51.355 4.704 ;
      RECT 51.32 4.542 51.325 4.697 ;
      RECT 51.305 4.54 51.32 4.693 ;
      RECT 51.285 4.54 51.305 4.688 ;
      RECT 51.28 4.539 51.285 4.686 ;
      RECT 51.275 4.539 51.28 4.683 ;
      RECT 51.235 4.538 51.275 4.678 ;
      RECT 51.21 4.537 51.235 4.673 ;
      RECT 51.15 4.536 51.21 4.67 ;
      RECT 51.065 4.535 51.15 4.668 ;
      RECT 51.026 4.534 51.055 4.665 ;
      RECT 50.94 4.532 51.026 4.665 ;
      RECT 50.8 4.532 50.835 4.665 ;
      RECT 50.71 4.536 50.75 4.668 ;
      RECT 50.695 4.539 50.71 4.675 ;
      RECT 50.685 4.54 50.695 4.682 ;
      RECT 50.66 4.543 50.685 4.687 ;
      RECT 50.655 4.545 50.66 4.69 ;
      RECT 50.605 4.547 50.655 4.691 ;
      RECT 50.566 4.551 50.605 4.693 ;
      RECT 50.48 4.553 50.566 4.696 ;
      RECT 50.462 4.555 50.48 4.698 ;
      RECT 50.376 4.558 50.462 4.7 ;
      RECT 50.29 4.562 50.376 4.703 ;
      RECT 50.253 4.566 50.29 4.706 ;
      RECT 50.167 4.569 50.253 4.709 ;
      RECT 50.081 4.573 50.167 4.712 ;
      RECT 49.995 4.578 50.081 4.716 ;
      RECT 49.975 4.58 49.995 4.719 ;
      RECT 49.955 4.579 49.975 4.72 ;
      RECT 49.906 4.576 49.955 4.721 ;
      RECT 49.82 4.571 49.906 4.724 ;
      RECT 49.77 4.566 49.82 4.726 ;
      RECT 49.746 4.564 49.77 4.727 ;
      RECT 49.66 4.559 49.746 4.729 ;
      RECT 49.635 4.555 49.66 4.728 ;
      RECT 49.625 4.552 49.635 4.726 ;
      RECT 49.615 4.545 49.625 4.723 ;
      RECT 49.61 4.525 49.615 4.718 ;
      RECT 49.6 4.495 49.61 4.713 ;
      RECT 49.585 4.365 49.6 4.704 ;
      RECT 49.58 4.357 49.585 4.697 ;
      RECT 49.56 4.35 49.58 4.689 ;
      RECT 49.555 4.332 49.56 4.681 ;
      RECT 49.545 4.312 49.555 4.676 ;
      RECT 49.54 4.285 49.545 4.672 ;
      RECT 49.535 4.262 49.54 4.669 ;
      RECT 49.515 4.22 49.535 4.661 ;
      RECT 49.48 4.135 49.515 4.645 ;
      RECT 49.475 4.067 49.48 4.633 ;
      RECT 49.46 4.037 49.475 4.627 ;
      RECT 49.455 3.282 49.46 3.528 ;
      RECT 49.445 4.007 49.46 4.618 ;
      RECT 49.45 3.277 49.455 3.56 ;
      RECT 49.445 3.272 49.45 3.603 ;
      RECT 49.44 3.27 49.445 3.638 ;
      RECT 49.425 3.97 49.445 4.608 ;
      RECT 49.435 3.27 49.44 3.675 ;
      RECT 49.42 3.27 49.435 3.773 ;
      RECT 49.42 3.943 49.425 4.601 ;
      RECT 49.415 3.27 49.42 3.848 ;
      RECT 49.415 3.931 49.42 4.598 ;
      RECT 49.41 3.27 49.415 3.88 ;
      RECT 49.41 3.91 49.415 4.595 ;
      RECT 49.405 3.27 49.41 4.592 ;
      RECT 49.37 3.27 49.405 4.578 ;
      RECT 49.355 3.27 49.37 4.56 ;
      RECT 49.335 3.27 49.355 4.55 ;
      RECT 49.31 3.27 49.335 4.533 ;
      RECT 49.305 3.27 49.31 4.483 ;
      RECT 49.295 3.27 49.3 4.313 ;
      RECT 49.29 3.27 49.295 4.22 ;
      RECT 49.285 3.27 49.29 4.133 ;
      RECT 49.28 3.27 49.285 4.065 ;
      RECT 49.275 3.27 49.28 4.008 ;
      RECT 49.265 3.27 49.275 3.903 ;
      RECT 49.26 3.27 49.265 3.775 ;
      RECT 49.255 3.27 49.26 3.693 ;
      RECT 49.25 3.272 49.255 3.61 ;
      RECT 49.245 3.277 49.25 3.543 ;
      RECT 49.24 3.282 49.245 3.47 ;
      RECT 52.055 3.6 52.315 3.86 ;
      RECT 52.075 3.567 52.285 3.86 ;
      RECT 52.075 3.565 52.275 3.86 ;
      RECT 52.085 3.552 52.275 3.86 ;
      RECT 52.085 3.55 52.2 3.86 ;
      RECT 51.56 3.675 51.735 3.955 ;
      RECT 51.555 3.675 51.735 3.953 ;
      RECT 51.555 3.675 51.75 3.95 ;
      RECT 51.545 3.675 51.75 3.948 ;
      RECT 51.49 3.675 51.75 3.935 ;
      RECT 51.49 3.75 51.755 3.913 ;
      RECT 51.02 4.873 51.025 5.08 ;
      RECT 50.97 4.867 51.02 5.079 ;
      RECT 50.937 4.881 51.03 5.078 ;
      RECT 50.851 4.881 51.03 5.077 ;
      RECT 50.765 4.881 51.03 5.076 ;
      RECT 50.765 4.98 51.035 5.073 ;
      RECT 50.76 4.98 51.035 5.068 ;
      RECT 50.755 4.98 51.035 5.05 ;
      RECT 50.75 4.98 51.035 5.033 ;
      RECT 50.71 4.765 50.97 5.025 ;
      RECT 50.17 3.915 50.256 4.329 ;
      RECT 50.17 3.915 50.295 4.326 ;
      RECT 50.17 3.915 50.315 4.316 ;
      RECT 50.125 3.915 50.315 4.313 ;
      RECT 50.125 4.067 50.325 4.303 ;
      RECT 50.125 4.088 50.33 4.297 ;
      RECT 50.125 4.106 50.335 4.293 ;
      RECT 50.125 4.126 50.345 4.288 ;
      RECT 50.1 4.126 50.345 4.285 ;
      RECT 50.09 4.126 50.345 4.263 ;
      RECT 50.09 4.142 50.35 4.233 ;
      RECT 50.055 3.915 50.315 4.22 ;
      RECT 50.055 4.154 50.355 4.175 ;
      RECT 47.715 10.06 48.01 10.29 ;
      RECT 47.775 8.58 47.945 10.29 ;
      RECT 47.765 8.95 48.12 9.305 ;
      RECT 47.715 8.58 48.005 8.81 ;
      RECT 46.725 10.06 47.02 10.29 ;
      RECT 46.785 8.58 46.955 10.29 ;
      RECT 46.725 8.58 47.015 8.81 ;
      RECT 46.725 8.615 47.575 8.775 ;
      RECT 47.41 8.21 47.575 8.775 ;
      RECT 46.725 8.61 47.12 8.775 ;
      RECT 47.345 8.21 47.635 8.44 ;
      RECT 47.345 8.24 47.805 8.41 ;
      RECT 47.31 4.005 47.63 4.26 ;
      RECT 47.31 4.055 47.8 4.225 ;
      RECT 47.31 3.69 47.5 4.26 ;
      RECT 46.725 3.655 47.015 3.885 ;
      RECT 46.725 3.69 47.5 3.86 ;
      RECT 46.785 2.175 46.955 3.885 ;
      RECT 46.725 2.175 47.02 2.405 ;
      RECT 46.355 4.025 46.645 4.255 ;
      RECT 46.355 4.055 46.815 4.225 ;
      RECT 46.42 2.95 46.585 4.255 ;
      RECT 44.935 2.915 45.225 3.145 ;
      RECT 44.935 2.95 46.585 3.12 ;
      RECT 44.995 2.175 45.165 3.145 ;
      RECT 44.935 2.175 45.225 2.405 ;
      RECT 44.935 10.06 45.225 10.29 ;
      RECT 44.995 9.32 45.165 10.29 ;
      RECT 44.995 9.41 46.585 9.58 ;
      RECT 46.415 8.21 46.585 9.58 ;
      RECT 44.935 9.32 45.225 9.55 ;
      RECT 46.355 8.21 46.645 8.44 ;
      RECT 46.355 8.24 46.815 8.41 ;
      RECT 42.985 4 43.325 4.35 ;
      RECT 43.075 3.32 43.245 4.35 ;
      RECT 45.365 3.26 45.715 3.61 ;
      RECT 43.075 3.32 45.715 3.49 ;
      RECT 45.195 3.315 45.715 3.49 ;
      RECT 45.39 8.945 45.715 9.27 ;
      RECT 39.93 8.905 40.28 9.255 ;
      RECT 45.365 8.95 45.715 9.18 ;
      RECT 39.73 8.95 40.28 9.18 ;
      RECT 45.195 8.975 45.715 9.15 ;
      RECT 39.56 8.98 40.28 9.15 ;
      RECT 39.61 8.975 45.715 9.145 ;
      RECT 44.59 3.66 44.91 3.98 ;
      RECT 44.565 3.655 44.855 3.885 ;
      RECT 44.56 3.685 44.91 3.86 ;
      RECT 44.39 3.685 44.91 3.855 ;
      RECT 44.59 8.545 44.91 8.835 ;
      RECT 44.565 8.58 44.91 8.81 ;
      RECT 44.39 8.61 44.91 8.78 ;
      RECT 40.28 4.28 40.43 4.555 ;
      RECT 40.82 3.36 40.825 3.58 ;
      RECT 41.97 3.56 41.985 3.758 ;
      RECT 41.935 3.552 41.97 3.765 ;
      RECT 41.905 3.545 41.935 3.765 ;
      RECT 41.85 3.51 41.905 3.765 ;
      RECT 41.785 3.447 41.85 3.765 ;
      RECT 41.78 3.412 41.785 3.763 ;
      RECT 41.775 3.407 41.78 3.755 ;
      RECT 41.77 3.402 41.775 3.741 ;
      RECT 41.765 3.399 41.77 3.734 ;
      RECT 41.72 3.389 41.765 3.685 ;
      RECT 41.7 3.376 41.72 3.62 ;
      RECT 41.695 3.371 41.7 3.593 ;
      RECT 41.69 3.37 41.695 3.586 ;
      RECT 41.685 3.369 41.69 3.579 ;
      RECT 41.6 3.354 41.685 3.525 ;
      RECT 41.57 3.335 41.6 3.475 ;
      RECT 41.49 3.318 41.57 3.46 ;
      RECT 41.455 3.305 41.49 3.445 ;
      RECT 41.447 3.305 41.455 3.44 ;
      RECT 41.361 3.306 41.447 3.44 ;
      RECT 41.275 3.308 41.361 3.44 ;
      RECT 41.25 3.309 41.275 3.444 ;
      RECT 41.175 3.315 41.25 3.459 ;
      RECT 41.092 3.327 41.175 3.483 ;
      RECT 41.006 3.34 41.092 3.509 ;
      RECT 40.92 3.353 41.006 3.535 ;
      RECT 40.885 3.362 40.92 3.554 ;
      RECT 40.835 3.362 40.885 3.567 ;
      RECT 40.825 3.36 40.835 3.578 ;
      RECT 40.81 3.357 40.82 3.58 ;
      RECT 40.795 3.349 40.81 3.588 ;
      RECT 40.78 3.341 40.795 3.608 ;
      RECT 40.775 3.336 40.78 3.665 ;
      RECT 40.76 3.331 40.775 3.738 ;
      RECT 40.755 3.326 40.76 3.78 ;
      RECT 40.75 3.324 40.755 3.808 ;
      RECT 40.745 3.322 40.75 3.83 ;
      RECT 40.735 3.318 40.745 3.873 ;
      RECT 40.73 3.315 40.735 3.898 ;
      RECT 40.725 3.313 40.73 3.918 ;
      RECT 40.72 3.311 40.725 3.942 ;
      RECT 40.715 3.307 40.72 3.965 ;
      RECT 40.71 3.303 40.715 3.988 ;
      RECT 40.675 3.293 40.71 4.095 ;
      RECT 40.67 3.283 40.675 4.193 ;
      RECT 40.665 3.281 40.67 4.22 ;
      RECT 40.66 3.28 40.665 4.24 ;
      RECT 40.655 3.272 40.66 4.26 ;
      RECT 40.65 3.267 40.655 4.295 ;
      RECT 40.645 3.265 40.65 4.313 ;
      RECT 40.64 3.265 40.645 4.338 ;
      RECT 40.635 3.265 40.64 4.36 ;
      RECT 40.6 3.265 40.635 4.403 ;
      RECT 40.575 3.265 40.6 4.432 ;
      RECT 40.565 3.265 40.575 3.618 ;
      RECT 40.568 3.675 40.575 4.442 ;
      RECT 40.565 3.732 40.568 4.445 ;
      RECT 40.56 3.265 40.565 3.59 ;
      RECT 40.56 3.782 40.565 4.448 ;
      RECT 40.55 3.265 40.56 3.58 ;
      RECT 40.555 3.835 40.56 4.451 ;
      RECT 40.55 3.92 40.555 4.455 ;
      RECT 40.54 3.265 40.55 3.568 ;
      RECT 40.545 3.967 40.55 4.459 ;
      RECT 40.54 4.042 40.545 4.463 ;
      RECT 40.505 3.265 40.54 3.543 ;
      RECT 40.53 4.125 40.54 4.468 ;
      RECT 40.52 4.192 40.53 4.475 ;
      RECT 40.515 4.22 40.52 4.48 ;
      RECT 40.505 4.233 40.515 4.486 ;
      RECT 40.46 3.265 40.505 3.5 ;
      RECT 40.5 4.238 40.505 4.493 ;
      RECT 40.46 4.255 40.5 4.555 ;
      RECT 40.455 3.267 40.46 3.473 ;
      RECT 40.43 4.275 40.46 4.555 ;
      RECT 40.45 3.272 40.455 3.445 ;
      RECT 40.24 4.284 40.28 4.555 ;
      RECT 40.215 4.292 40.24 4.525 ;
      RECT 40.17 4.3 40.215 4.525 ;
      RECT 40.155 4.305 40.17 4.52 ;
      RECT 40.145 4.305 40.155 4.514 ;
      RECT 40.135 4.312 40.145 4.511 ;
      RECT 40.13 4.35 40.135 4.5 ;
      RECT 40.125 4.412 40.13 4.478 ;
      RECT 41.395 4.287 41.58 4.51 ;
      RECT 41.395 4.302 41.585 4.506 ;
      RECT 41.385 3.575 41.47 4.505 ;
      RECT 41.385 4.302 41.59 4.499 ;
      RECT 41.38 4.31 41.59 4.498 ;
      RECT 41.585 4.03 41.905 4.35 ;
      RECT 41.38 4.202 41.55 4.293 ;
      RECT 41.375 4.202 41.55 4.275 ;
      RECT 41.365 4.01 41.5 4.25 ;
      RECT 41.36 4.01 41.5 4.195 ;
      RECT 41.32 3.59 41.49 4.095 ;
      RECT 41.305 3.59 41.49 3.965 ;
      RECT 41.3 3.59 41.49 3.918 ;
      RECT 41.295 3.59 41.49 3.898 ;
      RECT 41.29 3.59 41.49 3.873 ;
      RECT 41.26 3.59 41.52 3.85 ;
      RECT 41.27 3.587 41.48 3.85 ;
      RECT 41.395 3.582 41.48 4.51 ;
      RECT 41.28 3.575 41.47 3.85 ;
      RECT 41.275 3.58 41.47 3.85 ;
      RECT 40.105 3.792 40.29 4.005 ;
      RECT 40.105 3.8 40.3 3.998 ;
      RECT 40.085 3.8 40.3 3.995 ;
      RECT 40.08 3.8 40.3 3.98 ;
      RECT 40.01 3.715 40.27 3.975 ;
      RECT 40.01 3.86 40.305 3.888 ;
      RECT 39.665 4.315 39.925 4.575 ;
      RECT 39.69 4.26 39.885 4.575 ;
      RECT 39.685 4.009 39.865 4.303 ;
      RECT 39.685 4.015 39.875 4.303 ;
      RECT 39.665 4.017 39.875 4.248 ;
      RECT 39.66 4.027 39.875 4.115 ;
      RECT 39.69 4.007 39.865 4.575 ;
      RECT 39.776 4.005 39.865 4.575 ;
      RECT 39.635 3.225 39.67 3.595 ;
      RECT 39.425 3.335 39.43 3.595 ;
      RECT 39.67 3.232 39.685 3.595 ;
      RECT 39.56 3.225 39.635 3.673 ;
      RECT 39.55 3.225 39.56 3.758 ;
      RECT 39.525 3.225 39.55 3.793 ;
      RECT 39.485 3.225 39.525 3.861 ;
      RECT 39.475 3.232 39.485 3.913 ;
      RECT 39.445 3.335 39.475 3.954 ;
      RECT 39.44 3.335 39.445 3.993 ;
      RECT 39.43 3.335 39.44 4.013 ;
      RECT 39.425 3.63 39.43 4.05 ;
      RECT 39.42 3.647 39.425 4.07 ;
      RECT 39.405 3.71 39.42 4.11 ;
      RECT 39.4 3.753 39.405 4.145 ;
      RECT 39.395 3.761 39.4 4.158 ;
      RECT 39.385 3.775 39.395 4.18 ;
      RECT 39.36 3.81 39.385 4.245 ;
      RECT 39.35 3.845 39.36 4.308 ;
      RECT 39.33 3.875 39.35 4.369 ;
      RECT 39.315 3.911 39.33 4.436 ;
      RECT 39.305 3.939 39.315 4.475 ;
      RECT 39.295 3.961 39.305 4.495 ;
      RECT 39.29 3.971 39.295 4.506 ;
      RECT 39.285 3.98 39.29 4.509 ;
      RECT 39.275 3.998 39.285 4.513 ;
      RECT 39.265 4.016 39.275 4.514 ;
      RECT 39.24 4.055 39.265 4.511 ;
      RECT 39.22 4.097 39.24 4.508 ;
      RECT 39.205 4.135 39.22 4.507 ;
      RECT 39.17 4.17 39.205 4.504 ;
      RECT 39.165 4.192 39.17 4.502 ;
      RECT 39.1 4.232 39.165 4.499 ;
      RECT 39.095 4.272 39.1 4.495 ;
      RECT 39.08 4.282 39.095 4.486 ;
      RECT 39.07 4.402 39.08 4.471 ;
      RECT 39.55 4.815 39.56 5.075 ;
      RECT 39.55 4.818 39.57 5.074 ;
      RECT 39.54 4.808 39.55 5.073 ;
      RECT 39.53 4.823 39.61 5.069 ;
      RECT 39.515 4.802 39.53 5.067 ;
      RECT 39.49 4.827 39.615 5.063 ;
      RECT 39.475 4.787 39.49 5.058 ;
      RECT 39.475 4.829 39.625 5.057 ;
      RECT 39.475 4.837 39.64 5.05 ;
      RECT 39.415 4.774 39.475 5.04 ;
      RECT 39.405 4.761 39.415 5.022 ;
      RECT 39.38 4.751 39.405 5.012 ;
      RECT 39.375 4.741 39.38 5.004 ;
      RECT 39.31 4.837 39.64 4.986 ;
      RECT 39.225 4.837 39.64 4.948 ;
      RECT 39.115 4.665 39.375 4.925 ;
      RECT 39.49 4.795 39.515 5.063 ;
      RECT 39.53 4.805 39.54 5.069 ;
      RECT 39.115 4.813 39.555 4.925 ;
      RECT 39.3 10.06 39.59 10.29 ;
      RECT 39.36 9.32 39.53 10.29 ;
      RECT 39.26 9.345 39.63 9.715 ;
      RECT 39.3 9.32 39.59 9.715 ;
      RECT 38.33 4.57 38.36 4.87 ;
      RECT 38.105 4.555 38.11 4.83 ;
      RECT 37.905 4.555 38.06 4.815 ;
      RECT 39.205 3.27 39.235 3.53 ;
      RECT 39.195 3.27 39.205 3.638 ;
      RECT 39.175 3.27 39.195 3.648 ;
      RECT 39.16 3.27 39.175 3.66 ;
      RECT 39.105 3.27 39.16 3.71 ;
      RECT 39.09 3.27 39.105 3.758 ;
      RECT 39.06 3.27 39.09 3.793 ;
      RECT 39.005 3.27 39.06 3.855 ;
      RECT 38.985 3.27 39.005 3.923 ;
      RECT 38.98 3.27 38.985 3.953 ;
      RECT 38.975 3.27 38.98 3.965 ;
      RECT 38.97 3.387 38.975 3.983 ;
      RECT 38.95 3.405 38.97 4.008 ;
      RECT 38.93 3.432 38.95 4.058 ;
      RECT 38.925 3.452 38.93 4.089 ;
      RECT 38.92 3.46 38.925 4.106 ;
      RECT 38.905 3.486 38.92 4.135 ;
      RECT 38.89 3.528 38.905 4.17 ;
      RECT 38.885 3.557 38.89 4.193 ;
      RECT 38.88 3.572 38.885 4.206 ;
      RECT 38.875 3.595 38.88 4.217 ;
      RECT 38.865 3.615 38.875 4.235 ;
      RECT 38.855 3.645 38.865 4.258 ;
      RECT 38.85 3.667 38.855 4.278 ;
      RECT 38.845 3.682 38.85 4.293 ;
      RECT 38.83 3.712 38.845 4.32 ;
      RECT 38.825 3.742 38.83 4.346 ;
      RECT 38.82 3.76 38.825 4.358 ;
      RECT 38.81 3.79 38.82 4.377 ;
      RECT 38.8 3.815 38.81 4.402 ;
      RECT 38.795 3.835 38.8 4.421 ;
      RECT 38.79 3.852 38.795 4.434 ;
      RECT 38.78 3.878 38.79 4.453 ;
      RECT 38.77 3.916 38.78 4.48 ;
      RECT 38.765 3.942 38.77 4.5 ;
      RECT 38.76 3.952 38.765 4.51 ;
      RECT 38.755 3.965 38.76 4.525 ;
      RECT 38.75 3.98 38.755 4.535 ;
      RECT 38.745 4.002 38.75 4.55 ;
      RECT 38.74 4.02 38.745 4.561 ;
      RECT 38.735 4.03 38.74 4.572 ;
      RECT 38.73 4.038 38.735 4.584 ;
      RECT 38.725 4.046 38.73 4.595 ;
      RECT 38.72 4.072 38.725 4.608 ;
      RECT 38.71 4.1 38.72 4.621 ;
      RECT 38.705 4.13 38.71 4.63 ;
      RECT 38.7 4.145 38.705 4.637 ;
      RECT 38.685 4.17 38.7 4.644 ;
      RECT 38.68 4.192 38.685 4.65 ;
      RECT 38.675 4.217 38.68 4.653 ;
      RECT 38.666 4.245 38.675 4.657 ;
      RECT 38.66 4.262 38.666 4.662 ;
      RECT 38.655 4.28 38.66 4.666 ;
      RECT 38.65 4.292 38.655 4.669 ;
      RECT 38.645 4.313 38.65 4.673 ;
      RECT 38.64 4.331 38.645 4.676 ;
      RECT 38.635 4.345 38.64 4.679 ;
      RECT 38.63 4.362 38.635 4.682 ;
      RECT 38.625 4.375 38.63 4.685 ;
      RECT 38.6 4.412 38.625 4.693 ;
      RECT 38.595 4.457 38.6 4.702 ;
      RECT 38.59 4.485 38.595 4.705 ;
      RECT 38.58 4.505 38.59 4.709 ;
      RECT 38.575 4.525 38.58 4.714 ;
      RECT 38.57 4.54 38.575 4.717 ;
      RECT 38.55 4.55 38.57 4.724 ;
      RECT 38.485 4.557 38.55 4.75 ;
      RECT 38.45 4.56 38.485 4.778 ;
      RECT 38.435 4.563 38.45 4.793 ;
      RECT 38.425 4.564 38.435 4.808 ;
      RECT 38.415 4.565 38.425 4.825 ;
      RECT 38.41 4.565 38.415 4.84 ;
      RECT 38.405 4.565 38.41 4.848 ;
      RECT 38.39 4.566 38.405 4.863 ;
      RECT 38.36 4.568 38.39 4.87 ;
      RECT 38.25 4.575 38.33 4.87 ;
      RECT 38.205 4.58 38.25 4.87 ;
      RECT 38.195 4.581 38.205 4.86 ;
      RECT 38.185 4.582 38.195 4.853 ;
      RECT 38.165 4.584 38.185 4.848 ;
      RECT 38.155 4.555 38.165 4.843 ;
      RECT 38.11 4.555 38.155 4.835 ;
      RECT 38.08 4.555 38.105 4.825 ;
      RECT 38.06 4.555 38.08 4.818 ;
      RECT 38.34 3.355 38.6 3.615 ;
      RECT 38.22 3.37 38.23 3.535 ;
      RECT 38.205 3.37 38.21 3.53 ;
      RECT 35.57 3.21 35.755 3.5 ;
      RECT 37.385 3.335 37.4 3.49 ;
      RECT 35.535 3.21 35.56 3.47 ;
      RECT 37.95 3.26 37.955 3.402 ;
      RECT 37.865 3.255 37.89 3.395 ;
      RECT 38.265 3.372 38.34 3.565 ;
      RECT 38.25 3.37 38.265 3.548 ;
      RECT 38.23 3.37 38.25 3.54 ;
      RECT 38.21 3.37 38.22 3.533 ;
      RECT 38.165 3.365 38.205 3.523 ;
      RECT 38.125 3.34 38.165 3.508 ;
      RECT 38.11 3.315 38.125 3.498 ;
      RECT 38.105 3.309 38.11 3.496 ;
      RECT 38.07 3.301 38.105 3.479 ;
      RECT 38.065 3.294 38.07 3.467 ;
      RECT 38.045 3.289 38.065 3.455 ;
      RECT 38.035 3.283 38.045 3.44 ;
      RECT 38.015 3.278 38.035 3.425 ;
      RECT 38.005 3.273 38.015 3.418 ;
      RECT 38 3.271 38.005 3.413 ;
      RECT 37.995 3.27 38 3.41 ;
      RECT 37.955 3.265 37.995 3.406 ;
      RECT 37.935 3.259 37.95 3.401 ;
      RECT 37.9 3.256 37.935 3.398 ;
      RECT 37.89 3.255 37.9 3.396 ;
      RECT 37.83 3.255 37.865 3.393 ;
      RECT 37.785 3.255 37.83 3.393 ;
      RECT 37.735 3.255 37.785 3.396 ;
      RECT 37.72 3.257 37.735 3.398 ;
      RECT 37.705 3.26 37.72 3.399 ;
      RECT 37.695 3.265 37.705 3.4 ;
      RECT 37.665 3.27 37.695 3.405 ;
      RECT 37.655 3.276 37.665 3.413 ;
      RECT 37.645 3.278 37.655 3.417 ;
      RECT 37.635 3.282 37.645 3.421 ;
      RECT 37.61 3.288 37.635 3.429 ;
      RECT 37.6 3.293 37.61 3.437 ;
      RECT 37.585 3.297 37.6 3.441 ;
      RECT 37.55 3.303 37.585 3.449 ;
      RECT 37.53 3.308 37.55 3.459 ;
      RECT 37.5 3.315 37.53 3.468 ;
      RECT 37.455 3.324 37.5 3.482 ;
      RECT 37.45 3.329 37.455 3.493 ;
      RECT 37.43 3.332 37.45 3.494 ;
      RECT 37.4 3.335 37.43 3.492 ;
      RECT 37.365 3.335 37.385 3.488 ;
      RECT 37.295 3.335 37.365 3.479 ;
      RECT 37.28 3.332 37.295 3.471 ;
      RECT 37.24 3.325 37.28 3.466 ;
      RECT 37.215 3.315 37.24 3.459 ;
      RECT 37.21 3.309 37.215 3.456 ;
      RECT 37.17 3.303 37.21 3.453 ;
      RECT 37.155 3.296 37.17 3.448 ;
      RECT 37.135 3.292 37.155 3.443 ;
      RECT 37.12 3.287 37.135 3.439 ;
      RECT 37.105 3.282 37.12 3.437 ;
      RECT 37.09 3.278 37.105 3.436 ;
      RECT 37.075 3.276 37.09 3.432 ;
      RECT 37.065 3.274 37.075 3.427 ;
      RECT 37.05 3.271 37.065 3.423 ;
      RECT 37.04 3.269 37.05 3.418 ;
      RECT 37.02 3.266 37.04 3.414 ;
      RECT 36.975 3.265 37.02 3.412 ;
      RECT 36.915 3.267 36.975 3.413 ;
      RECT 36.895 3.269 36.915 3.415 ;
      RECT 36.865 3.272 36.895 3.416 ;
      RECT 36.815 3.277 36.865 3.418 ;
      RECT 36.81 3.28 36.815 3.42 ;
      RECT 36.8 3.282 36.81 3.423 ;
      RECT 36.795 3.284 36.8 3.426 ;
      RECT 36.745 3.287 36.795 3.433 ;
      RECT 36.725 3.291 36.745 3.445 ;
      RECT 36.715 3.294 36.725 3.451 ;
      RECT 36.705 3.295 36.715 3.454 ;
      RECT 36.666 3.298 36.705 3.456 ;
      RECT 36.58 3.305 36.666 3.459 ;
      RECT 36.506 3.315 36.58 3.463 ;
      RECT 36.42 3.326 36.506 3.468 ;
      RECT 36.405 3.333 36.42 3.47 ;
      RECT 36.35 3.337 36.405 3.471 ;
      RECT 36.336 3.34 36.35 3.473 ;
      RECT 36.25 3.34 36.336 3.475 ;
      RECT 36.21 3.337 36.25 3.478 ;
      RECT 36.186 3.333 36.21 3.48 ;
      RECT 36.1 3.323 36.186 3.483 ;
      RECT 36.07 3.312 36.1 3.484 ;
      RECT 36.051 3.308 36.07 3.483 ;
      RECT 35.965 3.301 36.051 3.48 ;
      RECT 35.905 3.29 35.965 3.477 ;
      RECT 35.885 3.282 35.905 3.475 ;
      RECT 35.85 3.277 35.885 3.474 ;
      RECT 35.825 3.272 35.85 3.473 ;
      RECT 35.795 3.267 35.825 3.472 ;
      RECT 35.77 3.21 35.795 3.471 ;
      RECT 35.755 3.21 35.77 3.495 ;
      RECT 35.56 3.21 35.57 3.495 ;
      RECT 37.335 4.23 37.34 4.37 ;
      RECT 36.995 4.23 37.03 4.368 ;
      RECT 36.57 4.215 36.585 4.36 ;
      RECT 38.4 3.995 38.49 4.255 ;
      RECT 38.23 3.86 38.33 4.255 ;
      RECT 35.265 3.835 35.345 4.045 ;
      RECT 38.355 3.972 38.4 4.255 ;
      RECT 38.345 3.942 38.355 4.255 ;
      RECT 38.33 3.865 38.345 4.255 ;
      RECT 38.145 3.86 38.23 4.22 ;
      RECT 38.14 3.862 38.145 4.215 ;
      RECT 38.135 3.867 38.14 4.215 ;
      RECT 38.1 3.967 38.135 4.215 ;
      RECT 38.09 3.995 38.1 4.215 ;
      RECT 38.08 4.01 38.09 4.215 ;
      RECT 38.07 4.022 38.08 4.215 ;
      RECT 38.065 4.032 38.07 4.215 ;
      RECT 38.05 4.042 38.065 4.217 ;
      RECT 38.045 4.057 38.05 4.219 ;
      RECT 38.03 4.07 38.045 4.221 ;
      RECT 38.025 4.085 38.03 4.224 ;
      RECT 38.005 4.095 38.025 4.228 ;
      RECT 37.99 4.105 38.005 4.231 ;
      RECT 37.955 4.112 37.99 4.236 ;
      RECT 37.911 4.119 37.955 4.244 ;
      RECT 37.825 4.131 37.911 4.257 ;
      RECT 37.8 4.142 37.825 4.268 ;
      RECT 37.77 4.147 37.8 4.273 ;
      RECT 37.735 4.152 37.77 4.281 ;
      RECT 37.705 4.157 37.735 4.288 ;
      RECT 37.68 4.162 37.705 4.293 ;
      RECT 37.615 4.169 37.68 4.302 ;
      RECT 37.545 4.182 37.615 4.318 ;
      RECT 37.515 4.192 37.545 4.33 ;
      RECT 37.49 4.197 37.515 4.337 ;
      RECT 37.435 4.204 37.49 4.345 ;
      RECT 37.43 4.211 37.435 4.35 ;
      RECT 37.425 4.213 37.43 4.351 ;
      RECT 37.41 4.215 37.425 4.353 ;
      RECT 37.405 4.215 37.41 4.356 ;
      RECT 37.34 4.222 37.405 4.363 ;
      RECT 37.305 4.232 37.335 4.373 ;
      RECT 37.288 4.235 37.305 4.375 ;
      RECT 37.202 4.234 37.288 4.374 ;
      RECT 37.116 4.232 37.202 4.371 ;
      RECT 37.03 4.231 37.116 4.369 ;
      RECT 36.929 4.229 36.995 4.368 ;
      RECT 36.843 4.226 36.929 4.366 ;
      RECT 36.757 4.222 36.843 4.364 ;
      RECT 36.671 4.219 36.757 4.363 ;
      RECT 36.585 4.216 36.671 4.361 ;
      RECT 36.485 4.215 36.57 4.358 ;
      RECT 36.435 4.213 36.485 4.356 ;
      RECT 36.415 4.21 36.435 4.354 ;
      RECT 36.395 4.208 36.415 4.351 ;
      RECT 36.37 4.204 36.395 4.348 ;
      RECT 36.325 4.198 36.37 4.343 ;
      RECT 36.285 4.192 36.325 4.335 ;
      RECT 36.26 4.187 36.285 4.328 ;
      RECT 36.205 4.18 36.26 4.32 ;
      RECT 36.181 4.173 36.205 4.313 ;
      RECT 36.095 4.164 36.181 4.303 ;
      RECT 36.065 4.156 36.095 4.293 ;
      RECT 36.035 4.152 36.065 4.288 ;
      RECT 36.03 4.149 36.035 4.285 ;
      RECT 36.025 4.148 36.03 4.285 ;
      RECT 35.95 4.141 36.025 4.278 ;
      RECT 35.911 4.132 35.95 4.267 ;
      RECT 35.825 4.122 35.911 4.255 ;
      RECT 35.785 4.112 35.825 4.243 ;
      RECT 35.746 4.107 35.785 4.236 ;
      RECT 35.66 4.097 35.746 4.225 ;
      RECT 35.62 4.085 35.66 4.214 ;
      RECT 35.585 4.07 35.62 4.207 ;
      RECT 35.575 4.06 35.585 4.204 ;
      RECT 35.555 4.045 35.575 4.202 ;
      RECT 35.525 4.015 35.555 4.198 ;
      RECT 35.515 3.995 35.525 4.193 ;
      RECT 35.51 3.987 35.515 4.19 ;
      RECT 35.505 3.98 35.51 4.188 ;
      RECT 35.49 3.967 35.505 4.181 ;
      RECT 35.485 3.957 35.49 4.173 ;
      RECT 35.48 3.95 35.485 4.168 ;
      RECT 35.475 3.945 35.48 4.164 ;
      RECT 35.46 3.932 35.475 4.156 ;
      RECT 35.455 3.842 35.46 4.145 ;
      RECT 35.45 3.837 35.455 4.138 ;
      RECT 35.375 3.835 35.45 4.098 ;
      RECT 35.345 3.835 35.375 4.053 ;
      RECT 35.25 3.84 35.265 4.04 ;
      RECT 37.735 3.545 37.995 3.805 ;
      RECT 37.72 3.533 37.9 3.77 ;
      RECT 37.715 3.534 37.9 3.768 ;
      RECT 37.7 3.538 37.91 3.758 ;
      RECT 37.695 3.543 37.915 3.728 ;
      RECT 37.7 3.54 37.915 3.758 ;
      RECT 37.715 3.535 37.91 3.768 ;
      RECT 37.735 3.532 37.9 3.805 ;
      RECT 37.735 3.531 37.89 3.805 ;
      RECT 37.76 3.53 37.89 3.805 ;
      RECT 37.32 3.775 37.58 4.035 ;
      RECT 37.195 3.82 37.58 4.03 ;
      RECT 37.185 3.825 37.58 4.025 ;
      RECT 37.2 4.765 37.215 5.075 ;
      RECT 35.795 4.535 35.805 4.665 ;
      RECT 35.575 4.53 35.68 4.665 ;
      RECT 35.49 4.535 35.54 4.665 ;
      RECT 34.04 3.27 34.045 4.375 ;
      RECT 37.295 4.857 37.3 4.993 ;
      RECT 37.29 4.852 37.295 5.053 ;
      RECT 37.285 4.85 37.29 5.066 ;
      RECT 37.27 4.847 37.285 5.068 ;
      RECT 37.265 4.842 37.27 5.07 ;
      RECT 37.26 4.838 37.265 5.073 ;
      RECT 37.245 4.833 37.26 5.075 ;
      RECT 37.215 4.825 37.245 5.075 ;
      RECT 37.176 4.765 37.2 5.075 ;
      RECT 37.09 4.765 37.176 5.072 ;
      RECT 37.06 4.765 37.09 5.065 ;
      RECT 37.035 4.765 37.06 5.058 ;
      RECT 37.01 4.765 37.035 5.05 ;
      RECT 36.995 4.765 37.01 5.043 ;
      RECT 36.97 4.765 36.995 5.035 ;
      RECT 36.955 4.765 36.97 5.028 ;
      RECT 36.915 4.775 36.955 5.017 ;
      RECT 36.905 4.77 36.915 5.007 ;
      RECT 36.901 4.769 36.905 5.004 ;
      RECT 36.815 4.761 36.901 4.987 ;
      RECT 36.782 4.75 36.815 4.964 ;
      RECT 36.696 4.739 36.782 4.942 ;
      RECT 36.61 4.723 36.696 4.911 ;
      RECT 36.54 4.708 36.61 4.883 ;
      RECT 36.53 4.701 36.54 4.87 ;
      RECT 36.5 4.698 36.53 4.86 ;
      RECT 36.475 4.694 36.5 4.853 ;
      RECT 36.46 4.691 36.475 4.848 ;
      RECT 36.455 4.69 36.46 4.843 ;
      RECT 36.425 4.685 36.455 4.836 ;
      RECT 36.42 4.68 36.425 4.831 ;
      RECT 36.405 4.677 36.42 4.826 ;
      RECT 36.4 4.672 36.405 4.821 ;
      RECT 36.38 4.667 36.4 4.818 ;
      RECT 36.365 4.662 36.38 4.81 ;
      RECT 36.35 4.656 36.365 4.805 ;
      RECT 36.32 4.647 36.35 4.798 ;
      RECT 36.315 4.64 36.32 4.79 ;
      RECT 36.31 4.638 36.315 4.788 ;
      RECT 36.305 4.637 36.31 4.785 ;
      RECT 36.265 4.63 36.305 4.778 ;
      RECT 36.251 4.62 36.265 4.768 ;
      RECT 36.2 4.609 36.251 4.756 ;
      RECT 36.175 4.595 36.2 4.742 ;
      RECT 36.15 4.584 36.175 4.734 ;
      RECT 36.13 4.573 36.15 4.728 ;
      RECT 36.12 4.567 36.13 4.723 ;
      RECT 36.115 4.565 36.12 4.719 ;
      RECT 36.095 4.56 36.115 4.714 ;
      RECT 36.065 4.55 36.095 4.704 ;
      RECT 36.06 4.542 36.065 4.697 ;
      RECT 36.045 4.54 36.06 4.693 ;
      RECT 36.025 4.54 36.045 4.688 ;
      RECT 36.02 4.539 36.025 4.686 ;
      RECT 36.015 4.539 36.02 4.683 ;
      RECT 35.975 4.538 36.015 4.678 ;
      RECT 35.95 4.537 35.975 4.673 ;
      RECT 35.89 4.536 35.95 4.67 ;
      RECT 35.805 4.535 35.89 4.668 ;
      RECT 35.766 4.534 35.795 4.665 ;
      RECT 35.68 4.532 35.766 4.665 ;
      RECT 35.54 4.532 35.575 4.665 ;
      RECT 35.45 4.536 35.49 4.668 ;
      RECT 35.435 4.539 35.45 4.675 ;
      RECT 35.425 4.54 35.435 4.682 ;
      RECT 35.4 4.543 35.425 4.687 ;
      RECT 35.395 4.545 35.4 4.69 ;
      RECT 35.345 4.547 35.395 4.691 ;
      RECT 35.306 4.551 35.345 4.693 ;
      RECT 35.22 4.553 35.306 4.696 ;
      RECT 35.202 4.555 35.22 4.698 ;
      RECT 35.116 4.558 35.202 4.7 ;
      RECT 35.03 4.562 35.116 4.703 ;
      RECT 34.993 4.566 35.03 4.706 ;
      RECT 34.907 4.569 34.993 4.709 ;
      RECT 34.821 4.573 34.907 4.712 ;
      RECT 34.735 4.578 34.821 4.716 ;
      RECT 34.715 4.58 34.735 4.719 ;
      RECT 34.695 4.579 34.715 4.72 ;
      RECT 34.646 4.576 34.695 4.721 ;
      RECT 34.56 4.571 34.646 4.724 ;
      RECT 34.51 4.566 34.56 4.726 ;
      RECT 34.486 4.564 34.51 4.727 ;
      RECT 34.4 4.559 34.486 4.729 ;
      RECT 34.375 4.555 34.4 4.728 ;
      RECT 34.365 4.552 34.375 4.726 ;
      RECT 34.355 4.545 34.365 4.723 ;
      RECT 34.35 4.525 34.355 4.718 ;
      RECT 34.34 4.495 34.35 4.713 ;
      RECT 34.325 4.365 34.34 4.704 ;
      RECT 34.32 4.357 34.325 4.697 ;
      RECT 34.3 4.35 34.32 4.689 ;
      RECT 34.295 4.332 34.3 4.681 ;
      RECT 34.285 4.312 34.295 4.676 ;
      RECT 34.28 4.285 34.285 4.672 ;
      RECT 34.275 4.262 34.28 4.669 ;
      RECT 34.255 4.22 34.275 4.661 ;
      RECT 34.22 4.135 34.255 4.645 ;
      RECT 34.215 4.067 34.22 4.633 ;
      RECT 34.2 4.037 34.215 4.627 ;
      RECT 34.195 3.282 34.2 3.528 ;
      RECT 34.185 4.007 34.2 4.618 ;
      RECT 34.19 3.277 34.195 3.56 ;
      RECT 34.185 3.272 34.19 3.603 ;
      RECT 34.18 3.27 34.185 3.638 ;
      RECT 34.165 3.97 34.185 4.608 ;
      RECT 34.175 3.27 34.18 3.675 ;
      RECT 34.16 3.27 34.175 3.773 ;
      RECT 34.16 3.943 34.165 4.601 ;
      RECT 34.155 3.27 34.16 3.848 ;
      RECT 34.155 3.931 34.16 4.598 ;
      RECT 34.15 3.27 34.155 3.88 ;
      RECT 34.15 3.91 34.155 4.595 ;
      RECT 34.145 3.27 34.15 4.592 ;
      RECT 34.11 3.27 34.145 4.578 ;
      RECT 34.095 3.27 34.11 4.56 ;
      RECT 34.075 3.27 34.095 4.55 ;
      RECT 34.05 3.27 34.075 4.533 ;
      RECT 34.045 3.27 34.05 4.483 ;
      RECT 34.035 3.27 34.04 4.313 ;
      RECT 34.03 3.27 34.035 4.22 ;
      RECT 34.025 3.27 34.03 4.133 ;
      RECT 34.02 3.27 34.025 4.065 ;
      RECT 34.015 3.27 34.02 4.008 ;
      RECT 34.005 3.27 34.015 3.903 ;
      RECT 34 3.27 34.005 3.775 ;
      RECT 33.995 3.27 34 3.693 ;
      RECT 33.99 3.272 33.995 3.61 ;
      RECT 33.985 3.277 33.99 3.543 ;
      RECT 33.98 3.282 33.985 3.47 ;
      RECT 36.795 3.6 37.055 3.86 ;
      RECT 36.815 3.567 37.025 3.86 ;
      RECT 36.815 3.565 37.015 3.86 ;
      RECT 36.825 3.552 37.015 3.86 ;
      RECT 36.825 3.55 36.94 3.86 ;
      RECT 36.3 3.675 36.475 3.955 ;
      RECT 36.295 3.675 36.475 3.953 ;
      RECT 36.295 3.675 36.49 3.95 ;
      RECT 36.285 3.675 36.49 3.948 ;
      RECT 36.23 3.675 36.49 3.935 ;
      RECT 36.23 3.75 36.495 3.913 ;
      RECT 35.76 4.873 35.765 5.08 ;
      RECT 35.71 4.867 35.76 5.079 ;
      RECT 35.677 4.881 35.77 5.078 ;
      RECT 35.591 4.881 35.77 5.077 ;
      RECT 35.505 4.881 35.77 5.076 ;
      RECT 35.505 4.98 35.775 5.073 ;
      RECT 35.5 4.98 35.775 5.068 ;
      RECT 35.495 4.98 35.775 5.05 ;
      RECT 35.49 4.98 35.775 5.033 ;
      RECT 35.45 4.765 35.71 5.025 ;
      RECT 34.91 3.915 34.996 4.329 ;
      RECT 34.91 3.915 35.035 4.326 ;
      RECT 34.91 3.915 35.055 4.316 ;
      RECT 34.865 3.915 35.055 4.313 ;
      RECT 34.865 4.067 35.065 4.303 ;
      RECT 34.865 4.088 35.07 4.297 ;
      RECT 34.865 4.106 35.075 4.293 ;
      RECT 34.865 4.126 35.085 4.288 ;
      RECT 34.84 4.126 35.085 4.285 ;
      RECT 34.83 4.126 35.085 4.263 ;
      RECT 34.83 4.142 35.09 4.233 ;
      RECT 34.795 3.915 35.055 4.22 ;
      RECT 34.795 4.154 35.095 4.175 ;
      RECT 32.455 10.06 32.75 10.29 ;
      RECT 32.515 8.58 32.685 10.29 ;
      RECT 32.51 8.95 32.86 9.3 ;
      RECT 32.455 8.58 32.745 8.81 ;
      RECT 31.465 10.06 31.76 10.29 ;
      RECT 31.525 8.58 31.695 10.29 ;
      RECT 31.465 8.58 31.755 8.81 ;
      RECT 31.465 8.615 32.315 8.775 ;
      RECT 32.15 8.21 32.315 8.775 ;
      RECT 31.465 8.61 31.86 8.775 ;
      RECT 32.085 8.21 32.375 8.44 ;
      RECT 32.085 8.24 32.545 8.41 ;
      RECT 32.05 4.005 32.37 4.26 ;
      RECT 32.05 4.055 32.54 4.225 ;
      RECT 32.05 3.69 32.24 4.26 ;
      RECT 31.465 3.655 31.755 3.885 ;
      RECT 31.465 3.69 32.24 3.86 ;
      RECT 31.525 2.175 31.695 3.885 ;
      RECT 31.465 2.175 31.76 2.405 ;
      RECT 31.095 4.025 31.385 4.255 ;
      RECT 31.095 4.055 31.555 4.225 ;
      RECT 31.16 2.95 31.325 4.255 ;
      RECT 29.675 2.915 29.965 3.145 ;
      RECT 29.675 2.95 31.325 3.12 ;
      RECT 29.735 2.175 29.905 3.145 ;
      RECT 29.675 2.175 29.965 2.405 ;
      RECT 29.675 10.06 29.965 10.29 ;
      RECT 29.735 9.32 29.905 10.29 ;
      RECT 29.735 9.41 31.325 9.58 ;
      RECT 31.155 8.21 31.325 9.58 ;
      RECT 29.675 9.32 29.965 9.55 ;
      RECT 31.095 8.21 31.385 8.44 ;
      RECT 31.095 8.24 31.555 8.41 ;
      RECT 27.725 4 28.065 4.35 ;
      RECT 27.815 3.32 27.985 4.35 ;
      RECT 30.105 3.26 30.455 3.61 ;
      RECT 27.815 3.32 30.455 3.49 ;
      RECT 29.935 3.315 30.455 3.49 ;
      RECT 30.13 8.945 30.455 9.27 ;
      RECT 24.67 8.895 25.02 9.245 ;
      RECT 30.105 8.95 30.455 9.18 ;
      RECT 24.47 8.95 25.02 9.18 ;
      RECT 29.935 8.975 30.455 9.15 ;
      RECT 24.3 8.98 25.02 9.15 ;
      RECT 24.35 8.975 30.455 9.145 ;
      RECT 29.33 3.66 29.65 3.98 ;
      RECT 29.305 3.655 29.595 3.885 ;
      RECT 29.3 3.685 29.65 3.86 ;
      RECT 29.13 3.685 29.65 3.855 ;
      RECT 29.33 8.545 29.65 8.835 ;
      RECT 29.305 8.58 29.65 8.81 ;
      RECT 29.13 8.61 29.65 8.78 ;
      RECT 25.02 4.28 25.17 4.555 ;
      RECT 25.56 3.36 25.565 3.58 ;
      RECT 26.71 3.56 26.725 3.758 ;
      RECT 26.675 3.552 26.71 3.765 ;
      RECT 26.645 3.545 26.675 3.765 ;
      RECT 26.59 3.51 26.645 3.765 ;
      RECT 26.525 3.447 26.59 3.765 ;
      RECT 26.52 3.412 26.525 3.763 ;
      RECT 26.515 3.407 26.52 3.755 ;
      RECT 26.51 3.402 26.515 3.741 ;
      RECT 26.505 3.399 26.51 3.734 ;
      RECT 26.46 3.389 26.505 3.685 ;
      RECT 26.44 3.376 26.46 3.62 ;
      RECT 26.435 3.371 26.44 3.593 ;
      RECT 26.43 3.37 26.435 3.586 ;
      RECT 26.425 3.369 26.43 3.579 ;
      RECT 26.34 3.354 26.425 3.525 ;
      RECT 26.31 3.335 26.34 3.475 ;
      RECT 26.23 3.318 26.31 3.46 ;
      RECT 26.195 3.305 26.23 3.445 ;
      RECT 26.187 3.305 26.195 3.44 ;
      RECT 26.101 3.306 26.187 3.44 ;
      RECT 26.015 3.308 26.101 3.44 ;
      RECT 25.99 3.309 26.015 3.444 ;
      RECT 25.915 3.315 25.99 3.459 ;
      RECT 25.832 3.327 25.915 3.483 ;
      RECT 25.746 3.34 25.832 3.509 ;
      RECT 25.66 3.353 25.746 3.535 ;
      RECT 25.625 3.362 25.66 3.554 ;
      RECT 25.575 3.362 25.625 3.567 ;
      RECT 25.565 3.36 25.575 3.578 ;
      RECT 25.55 3.357 25.56 3.58 ;
      RECT 25.535 3.349 25.55 3.588 ;
      RECT 25.52 3.341 25.535 3.608 ;
      RECT 25.515 3.336 25.52 3.665 ;
      RECT 25.5 3.331 25.515 3.738 ;
      RECT 25.495 3.326 25.5 3.78 ;
      RECT 25.49 3.324 25.495 3.808 ;
      RECT 25.485 3.322 25.49 3.83 ;
      RECT 25.475 3.318 25.485 3.873 ;
      RECT 25.47 3.315 25.475 3.898 ;
      RECT 25.465 3.313 25.47 3.918 ;
      RECT 25.46 3.311 25.465 3.942 ;
      RECT 25.455 3.307 25.46 3.965 ;
      RECT 25.45 3.303 25.455 3.988 ;
      RECT 25.415 3.293 25.45 4.095 ;
      RECT 25.41 3.283 25.415 4.193 ;
      RECT 25.405 3.281 25.41 4.22 ;
      RECT 25.4 3.28 25.405 4.24 ;
      RECT 25.395 3.272 25.4 4.26 ;
      RECT 25.39 3.267 25.395 4.295 ;
      RECT 25.385 3.265 25.39 4.313 ;
      RECT 25.38 3.265 25.385 4.338 ;
      RECT 25.375 3.265 25.38 4.36 ;
      RECT 25.34 3.265 25.375 4.403 ;
      RECT 25.315 3.265 25.34 4.432 ;
      RECT 25.305 3.265 25.315 3.618 ;
      RECT 25.308 3.675 25.315 4.442 ;
      RECT 25.305 3.732 25.308 4.445 ;
      RECT 25.3 3.265 25.305 3.59 ;
      RECT 25.3 3.782 25.305 4.448 ;
      RECT 25.29 3.265 25.3 3.58 ;
      RECT 25.295 3.835 25.3 4.451 ;
      RECT 25.29 3.92 25.295 4.455 ;
      RECT 25.28 3.265 25.29 3.568 ;
      RECT 25.285 3.967 25.29 4.459 ;
      RECT 25.28 4.042 25.285 4.463 ;
      RECT 25.245 3.265 25.28 3.543 ;
      RECT 25.27 4.125 25.28 4.468 ;
      RECT 25.26 4.192 25.27 4.475 ;
      RECT 25.255 4.22 25.26 4.48 ;
      RECT 25.245 4.233 25.255 4.486 ;
      RECT 25.2 3.265 25.245 3.5 ;
      RECT 25.24 4.238 25.245 4.493 ;
      RECT 25.2 4.255 25.24 4.555 ;
      RECT 25.195 3.267 25.2 3.473 ;
      RECT 25.17 4.275 25.2 4.555 ;
      RECT 25.19 3.272 25.195 3.445 ;
      RECT 24.98 4.284 25.02 4.555 ;
      RECT 24.955 4.292 24.98 4.525 ;
      RECT 24.91 4.3 24.955 4.525 ;
      RECT 24.895 4.305 24.91 4.52 ;
      RECT 24.885 4.305 24.895 4.514 ;
      RECT 24.875 4.312 24.885 4.511 ;
      RECT 24.87 4.35 24.875 4.5 ;
      RECT 24.865 4.412 24.87 4.478 ;
      RECT 26.135 4.287 26.32 4.51 ;
      RECT 26.135 4.302 26.325 4.506 ;
      RECT 26.125 3.575 26.21 4.505 ;
      RECT 26.125 4.302 26.33 4.499 ;
      RECT 26.12 4.31 26.33 4.498 ;
      RECT 26.325 4.03 26.645 4.35 ;
      RECT 26.12 4.202 26.29 4.293 ;
      RECT 26.115 4.202 26.29 4.275 ;
      RECT 26.105 4.01 26.24 4.25 ;
      RECT 26.1 4.01 26.24 4.195 ;
      RECT 26.06 3.59 26.23 4.095 ;
      RECT 26.045 3.59 26.23 3.965 ;
      RECT 26.04 3.59 26.23 3.918 ;
      RECT 26.035 3.59 26.23 3.898 ;
      RECT 26.03 3.59 26.23 3.873 ;
      RECT 26 3.59 26.26 3.85 ;
      RECT 26.01 3.587 26.22 3.85 ;
      RECT 26.135 3.582 26.22 4.51 ;
      RECT 26.02 3.575 26.21 3.85 ;
      RECT 26.015 3.58 26.21 3.85 ;
      RECT 24.845 3.792 25.03 4.005 ;
      RECT 24.845 3.8 25.04 3.998 ;
      RECT 24.825 3.8 25.04 3.995 ;
      RECT 24.82 3.8 25.04 3.98 ;
      RECT 24.75 3.715 25.01 3.975 ;
      RECT 24.75 3.86 25.045 3.888 ;
      RECT 24.405 4.315 24.665 4.575 ;
      RECT 24.43 4.26 24.625 4.575 ;
      RECT 24.425 4.009 24.605 4.303 ;
      RECT 24.425 4.015 24.615 4.303 ;
      RECT 24.405 4.017 24.615 4.248 ;
      RECT 24.4 4.027 24.615 4.115 ;
      RECT 24.43 4.007 24.605 4.575 ;
      RECT 24.516 4.005 24.605 4.575 ;
      RECT 24.375 3.225 24.41 3.595 ;
      RECT 24.165 3.335 24.17 3.595 ;
      RECT 24.41 3.232 24.425 3.595 ;
      RECT 24.3 3.225 24.375 3.673 ;
      RECT 24.29 3.225 24.3 3.758 ;
      RECT 24.265 3.225 24.29 3.793 ;
      RECT 24.225 3.225 24.265 3.861 ;
      RECT 24.215 3.232 24.225 3.913 ;
      RECT 24.185 3.335 24.215 3.954 ;
      RECT 24.18 3.335 24.185 3.993 ;
      RECT 24.17 3.335 24.18 4.013 ;
      RECT 24.165 3.63 24.17 4.05 ;
      RECT 24.16 3.647 24.165 4.07 ;
      RECT 24.145 3.71 24.16 4.11 ;
      RECT 24.14 3.753 24.145 4.145 ;
      RECT 24.135 3.761 24.14 4.158 ;
      RECT 24.125 3.775 24.135 4.18 ;
      RECT 24.1 3.81 24.125 4.245 ;
      RECT 24.09 3.845 24.1 4.308 ;
      RECT 24.07 3.875 24.09 4.369 ;
      RECT 24.055 3.911 24.07 4.436 ;
      RECT 24.045 3.939 24.055 4.475 ;
      RECT 24.035 3.961 24.045 4.495 ;
      RECT 24.03 3.971 24.035 4.506 ;
      RECT 24.025 3.98 24.03 4.509 ;
      RECT 24.015 3.998 24.025 4.513 ;
      RECT 24.005 4.016 24.015 4.514 ;
      RECT 23.98 4.055 24.005 4.511 ;
      RECT 23.96 4.097 23.98 4.508 ;
      RECT 23.945 4.135 23.96 4.507 ;
      RECT 23.91 4.17 23.945 4.504 ;
      RECT 23.905 4.192 23.91 4.502 ;
      RECT 23.84 4.232 23.905 4.499 ;
      RECT 23.835 4.272 23.84 4.495 ;
      RECT 23.82 4.282 23.835 4.486 ;
      RECT 23.81 4.402 23.82 4.471 ;
      RECT 24.29 4.815 24.3 5.075 ;
      RECT 24.29 4.818 24.31 5.074 ;
      RECT 24.28 4.808 24.29 5.073 ;
      RECT 24.27 4.823 24.35 5.069 ;
      RECT 24.255 4.802 24.27 5.067 ;
      RECT 24.23 4.827 24.355 5.063 ;
      RECT 24.215 4.787 24.23 5.058 ;
      RECT 24.215 4.829 24.365 5.057 ;
      RECT 24.215 4.837 24.38 5.05 ;
      RECT 24.155 4.774 24.215 5.04 ;
      RECT 24.145 4.761 24.155 5.022 ;
      RECT 24.12 4.751 24.145 5.012 ;
      RECT 24.115 4.741 24.12 5.004 ;
      RECT 24.05 4.837 24.38 4.986 ;
      RECT 23.965 4.837 24.38 4.948 ;
      RECT 23.855 4.665 24.115 4.925 ;
      RECT 24.23 4.795 24.255 5.063 ;
      RECT 24.27 4.805 24.28 5.069 ;
      RECT 23.855 4.813 24.295 4.925 ;
      RECT 24.04 10.06 24.33 10.29 ;
      RECT 24.1 9.32 24.27 10.29 ;
      RECT 24 9.345 24.37 9.715 ;
      RECT 24.04 9.32 24.33 9.715 ;
      RECT 23.07 4.57 23.1 4.87 ;
      RECT 22.845 4.555 22.85 4.83 ;
      RECT 22.645 4.555 22.8 4.815 ;
      RECT 23.945 3.27 23.975 3.53 ;
      RECT 23.935 3.27 23.945 3.638 ;
      RECT 23.915 3.27 23.935 3.648 ;
      RECT 23.9 3.27 23.915 3.66 ;
      RECT 23.845 3.27 23.9 3.71 ;
      RECT 23.83 3.27 23.845 3.758 ;
      RECT 23.8 3.27 23.83 3.793 ;
      RECT 23.745 3.27 23.8 3.855 ;
      RECT 23.725 3.27 23.745 3.923 ;
      RECT 23.72 3.27 23.725 3.953 ;
      RECT 23.715 3.27 23.72 3.965 ;
      RECT 23.71 3.387 23.715 3.983 ;
      RECT 23.69 3.405 23.71 4.008 ;
      RECT 23.67 3.432 23.69 4.058 ;
      RECT 23.665 3.452 23.67 4.089 ;
      RECT 23.66 3.46 23.665 4.106 ;
      RECT 23.645 3.486 23.66 4.135 ;
      RECT 23.63 3.528 23.645 4.17 ;
      RECT 23.625 3.557 23.63 4.193 ;
      RECT 23.62 3.572 23.625 4.206 ;
      RECT 23.615 3.595 23.62 4.217 ;
      RECT 23.605 3.615 23.615 4.235 ;
      RECT 23.595 3.645 23.605 4.258 ;
      RECT 23.59 3.667 23.595 4.278 ;
      RECT 23.585 3.682 23.59 4.293 ;
      RECT 23.57 3.712 23.585 4.32 ;
      RECT 23.565 3.742 23.57 4.346 ;
      RECT 23.56 3.76 23.565 4.358 ;
      RECT 23.55 3.79 23.56 4.377 ;
      RECT 23.54 3.815 23.55 4.402 ;
      RECT 23.535 3.835 23.54 4.421 ;
      RECT 23.53 3.852 23.535 4.434 ;
      RECT 23.52 3.878 23.53 4.453 ;
      RECT 23.51 3.916 23.52 4.48 ;
      RECT 23.505 3.942 23.51 4.5 ;
      RECT 23.5 3.952 23.505 4.51 ;
      RECT 23.495 3.965 23.5 4.525 ;
      RECT 23.49 3.98 23.495 4.535 ;
      RECT 23.485 4.002 23.49 4.55 ;
      RECT 23.48 4.02 23.485 4.561 ;
      RECT 23.475 4.03 23.48 4.572 ;
      RECT 23.47 4.038 23.475 4.584 ;
      RECT 23.465 4.046 23.47 4.595 ;
      RECT 23.46 4.072 23.465 4.608 ;
      RECT 23.45 4.1 23.46 4.621 ;
      RECT 23.445 4.13 23.45 4.63 ;
      RECT 23.44 4.145 23.445 4.637 ;
      RECT 23.425 4.17 23.44 4.644 ;
      RECT 23.42 4.192 23.425 4.65 ;
      RECT 23.415 4.217 23.42 4.653 ;
      RECT 23.406 4.245 23.415 4.657 ;
      RECT 23.4 4.262 23.406 4.662 ;
      RECT 23.395 4.28 23.4 4.666 ;
      RECT 23.39 4.292 23.395 4.669 ;
      RECT 23.385 4.313 23.39 4.673 ;
      RECT 23.38 4.331 23.385 4.676 ;
      RECT 23.375 4.345 23.38 4.679 ;
      RECT 23.37 4.362 23.375 4.682 ;
      RECT 23.365 4.375 23.37 4.685 ;
      RECT 23.34 4.412 23.365 4.693 ;
      RECT 23.335 4.457 23.34 4.702 ;
      RECT 23.33 4.485 23.335 4.705 ;
      RECT 23.32 4.505 23.33 4.709 ;
      RECT 23.315 4.525 23.32 4.714 ;
      RECT 23.31 4.54 23.315 4.717 ;
      RECT 23.29 4.55 23.31 4.724 ;
      RECT 23.225 4.557 23.29 4.75 ;
      RECT 23.19 4.56 23.225 4.778 ;
      RECT 23.175 4.563 23.19 4.793 ;
      RECT 23.165 4.564 23.175 4.808 ;
      RECT 23.155 4.565 23.165 4.825 ;
      RECT 23.15 4.565 23.155 4.84 ;
      RECT 23.145 4.565 23.15 4.848 ;
      RECT 23.13 4.566 23.145 4.863 ;
      RECT 23.1 4.568 23.13 4.87 ;
      RECT 22.99 4.575 23.07 4.87 ;
      RECT 22.945 4.58 22.99 4.87 ;
      RECT 22.935 4.581 22.945 4.86 ;
      RECT 22.925 4.582 22.935 4.853 ;
      RECT 22.905 4.584 22.925 4.848 ;
      RECT 22.895 4.555 22.905 4.843 ;
      RECT 22.85 4.555 22.895 4.835 ;
      RECT 22.82 4.555 22.845 4.825 ;
      RECT 22.8 4.555 22.82 4.818 ;
      RECT 23.08 3.355 23.34 3.615 ;
      RECT 22.96 3.37 22.97 3.535 ;
      RECT 22.945 3.37 22.95 3.53 ;
      RECT 20.31 3.21 20.495 3.5 ;
      RECT 22.125 3.335 22.14 3.49 ;
      RECT 20.275 3.21 20.3 3.47 ;
      RECT 22.69 3.26 22.695 3.402 ;
      RECT 22.605 3.255 22.63 3.395 ;
      RECT 23.005 3.372 23.08 3.565 ;
      RECT 22.99 3.37 23.005 3.548 ;
      RECT 22.97 3.37 22.99 3.54 ;
      RECT 22.95 3.37 22.96 3.533 ;
      RECT 22.905 3.365 22.945 3.523 ;
      RECT 22.865 3.34 22.905 3.508 ;
      RECT 22.85 3.315 22.865 3.498 ;
      RECT 22.845 3.309 22.85 3.496 ;
      RECT 22.81 3.301 22.845 3.479 ;
      RECT 22.805 3.294 22.81 3.467 ;
      RECT 22.785 3.289 22.805 3.455 ;
      RECT 22.775 3.283 22.785 3.44 ;
      RECT 22.755 3.278 22.775 3.425 ;
      RECT 22.745 3.273 22.755 3.418 ;
      RECT 22.74 3.271 22.745 3.413 ;
      RECT 22.735 3.27 22.74 3.41 ;
      RECT 22.695 3.265 22.735 3.406 ;
      RECT 22.675 3.259 22.69 3.401 ;
      RECT 22.64 3.256 22.675 3.398 ;
      RECT 22.63 3.255 22.64 3.396 ;
      RECT 22.57 3.255 22.605 3.393 ;
      RECT 22.525 3.255 22.57 3.393 ;
      RECT 22.475 3.255 22.525 3.396 ;
      RECT 22.46 3.257 22.475 3.398 ;
      RECT 22.445 3.26 22.46 3.399 ;
      RECT 22.435 3.265 22.445 3.4 ;
      RECT 22.405 3.27 22.435 3.405 ;
      RECT 22.395 3.276 22.405 3.413 ;
      RECT 22.385 3.278 22.395 3.417 ;
      RECT 22.375 3.282 22.385 3.421 ;
      RECT 22.35 3.288 22.375 3.429 ;
      RECT 22.34 3.293 22.35 3.437 ;
      RECT 22.325 3.297 22.34 3.441 ;
      RECT 22.29 3.303 22.325 3.449 ;
      RECT 22.27 3.308 22.29 3.459 ;
      RECT 22.24 3.315 22.27 3.468 ;
      RECT 22.195 3.324 22.24 3.482 ;
      RECT 22.19 3.329 22.195 3.493 ;
      RECT 22.17 3.332 22.19 3.494 ;
      RECT 22.14 3.335 22.17 3.492 ;
      RECT 22.105 3.335 22.125 3.488 ;
      RECT 22.035 3.335 22.105 3.479 ;
      RECT 22.02 3.332 22.035 3.471 ;
      RECT 21.98 3.325 22.02 3.466 ;
      RECT 21.955 3.315 21.98 3.459 ;
      RECT 21.95 3.309 21.955 3.456 ;
      RECT 21.91 3.303 21.95 3.453 ;
      RECT 21.895 3.296 21.91 3.448 ;
      RECT 21.875 3.292 21.895 3.443 ;
      RECT 21.86 3.287 21.875 3.439 ;
      RECT 21.845 3.282 21.86 3.437 ;
      RECT 21.83 3.278 21.845 3.436 ;
      RECT 21.815 3.276 21.83 3.432 ;
      RECT 21.805 3.274 21.815 3.427 ;
      RECT 21.79 3.271 21.805 3.423 ;
      RECT 21.78 3.269 21.79 3.418 ;
      RECT 21.76 3.266 21.78 3.414 ;
      RECT 21.715 3.265 21.76 3.412 ;
      RECT 21.655 3.267 21.715 3.413 ;
      RECT 21.635 3.269 21.655 3.415 ;
      RECT 21.605 3.272 21.635 3.416 ;
      RECT 21.555 3.277 21.605 3.418 ;
      RECT 21.55 3.28 21.555 3.42 ;
      RECT 21.54 3.282 21.55 3.423 ;
      RECT 21.535 3.284 21.54 3.426 ;
      RECT 21.485 3.287 21.535 3.433 ;
      RECT 21.465 3.291 21.485 3.445 ;
      RECT 21.455 3.294 21.465 3.451 ;
      RECT 21.445 3.295 21.455 3.454 ;
      RECT 21.406 3.298 21.445 3.456 ;
      RECT 21.32 3.305 21.406 3.459 ;
      RECT 21.246 3.315 21.32 3.463 ;
      RECT 21.16 3.326 21.246 3.468 ;
      RECT 21.145 3.333 21.16 3.47 ;
      RECT 21.09 3.337 21.145 3.471 ;
      RECT 21.076 3.34 21.09 3.473 ;
      RECT 20.99 3.34 21.076 3.475 ;
      RECT 20.95 3.337 20.99 3.478 ;
      RECT 20.926 3.333 20.95 3.48 ;
      RECT 20.84 3.323 20.926 3.483 ;
      RECT 20.81 3.312 20.84 3.484 ;
      RECT 20.791 3.308 20.81 3.483 ;
      RECT 20.705 3.301 20.791 3.48 ;
      RECT 20.645 3.29 20.705 3.477 ;
      RECT 20.625 3.282 20.645 3.475 ;
      RECT 20.59 3.277 20.625 3.474 ;
      RECT 20.565 3.272 20.59 3.473 ;
      RECT 20.535 3.267 20.565 3.472 ;
      RECT 20.51 3.21 20.535 3.471 ;
      RECT 20.495 3.21 20.51 3.495 ;
      RECT 20.3 3.21 20.31 3.495 ;
      RECT 22.075 4.23 22.08 4.37 ;
      RECT 21.735 4.23 21.77 4.368 ;
      RECT 21.31 4.215 21.325 4.36 ;
      RECT 23.14 3.995 23.23 4.255 ;
      RECT 22.97 3.86 23.07 4.255 ;
      RECT 20.005 3.835 20.085 4.045 ;
      RECT 23.095 3.972 23.14 4.255 ;
      RECT 23.085 3.942 23.095 4.255 ;
      RECT 23.07 3.865 23.085 4.255 ;
      RECT 22.885 3.86 22.97 4.22 ;
      RECT 22.88 3.862 22.885 4.215 ;
      RECT 22.875 3.867 22.88 4.215 ;
      RECT 22.84 3.967 22.875 4.215 ;
      RECT 22.83 3.995 22.84 4.215 ;
      RECT 22.82 4.01 22.83 4.215 ;
      RECT 22.81 4.022 22.82 4.215 ;
      RECT 22.805 4.032 22.81 4.215 ;
      RECT 22.79 4.042 22.805 4.217 ;
      RECT 22.785 4.057 22.79 4.219 ;
      RECT 22.77 4.07 22.785 4.221 ;
      RECT 22.765 4.085 22.77 4.224 ;
      RECT 22.745 4.095 22.765 4.228 ;
      RECT 22.73 4.105 22.745 4.231 ;
      RECT 22.695 4.112 22.73 4.236 ;
      RECT 22.651 4.119 22.695 4.244 ;
      RECT 22.565 4.131 22.651 4.257 ;
      RECT 22.54 4.142 22.565 4.268 ;
      RECT 22.51 4.147 22.54 4.273 ;
      RECT 22.475 4.152 22.51 4.281 ;
      RECT 22.445 4.157 22.475 4.288 ;
      RECT 22.42 4.162 22.445 4.293 ;
      RECT 22.355 4.169 22.42 4.302 ;
      RECT 22.285 4.182 22.355 4.318 ;
      RECT 22.255 4.192 22.285 4.33 ;
      RECT 22.23 4.197 22.255 4.337 ;
      RECT 22.175 4.204 22.23 4.345 ;
      RECT 22.17 4.211 22.175 4.35 ;
      RECT 22.165 4.213 22.17 4.351 ;
      RECT 22.15 4.215 22.165 4.353 ;
      RECT 22.145 4.215 22.15 4.356 ;
      RECT 22.08 4.222 22.145 4.363 ;
      RECT 22.045 4.232 22.075 4.373 ;
      RECT 22.028 4.235 22.045 4.375 ;
      RECT 21.942 4.234 22.028 4.374 ;
      RECT 21.856 4.232 21.942 4.371 ;
      RECT 21.77 4.231 21.856 4.369 ;
      RECT 21.669 4.229 21.735 4.368 ;
      RECT 21.583 4.226 21.669 4.366 ;
      RECT 21.497 4.222 21.583 4.364 ;
      RECT 21.411 4.219 21.497 4.363 ;
      RECT 21.325 4.216 21.411 4.361 ;
      RECT 21.225 4.215 21.31 4.358 ;
      RECT 21.175 4.213 21.225 4.356 ;
      RECT 21.155 4.21 21.175 4.354 ;
      RECT 21.135 4.208 21.155 4.351 ;
      RECT 21.11 4.204 21.135 4.348 ;
      RECT 21.065 4.198 21.11 4.343 ;
      RECT 21.025 4.192 21.065 4.335 ;
      RECT 21 4.187 21.025 4.328 ;
      RECT 20.945 4.18 21 4.32 ;
      RECT 20.921 4.173 20.945 4.313 ;
      RECT 20.835 4.164 20.921 4.303 ;
      RECT 20.805 4.156 20.835 4.293 ;
      RECT 20.775 4.152 20.805 4.288 ;
      RECT 20.77 4.149 20.775 4.285 ;
      RECT 20.765 4.148 20.77 4.285 ;
      RECT 20.69 4.141 20.765 4.278 ;
      RECT 20.651 4.132 20.69 4.267 ;
      RECT 20.565 4.122 20.651 4.255 ;
      RECT 20.525 4.112 20.565 4.243 ;
      RECT 20.486 4.107 20.525 4.236 ;
      RECT 20.4 4.097 20.486 4.225 ;
      RECT 20.36 4.085 20.4 4.214 ;
      RECT 20.325 4.07 20.36 4.207 ;
      RECT 20.315 4.06 20.325 4.204 ;
      RECT 20.295 4.045 20.315 4.202 ;
      RECT 20.265 4.015 20.295 4.198 ;
      RECT 20.255 3.995 20.265 4.193 ;
      RECT 20.25 3.987 20.255 4.19 ;
      RECT 20.245 3.98 20.25 4.188 ;
      RECT 20.23 3.967 20.245 4.181 ;
      RECT 20.225 3.957 20.23 4.173 ;
      RECT 20.22 3.95 20.225 4.168 ;
      RECT 20.215 3.945 20.22 4.164 ;
      RECT 20.2 3.932 20.215 4.156 ;
      RECT 20.195 3.842 20.2 4.145 ;
      RECT 20.19 3.837 20.195 4.138 ;
      RECT 20.115 3.835 20.19 4.098 ;
      RECT 20.085 3.835 20.115 4.053 ;
      RECT 19.99 3.84 20.005 4.04 ;
      RECT 22.475 3.545 22.735 3.805 ;
      RECT 22.46 3.533 22.64 3.77 ;
      RECT 22.455 3.534 22.64 3.768 ;
      RECT 22.44 3.538 22.65 3.758 ;
      RECT 22.435 3.543 22.655 3.728 ;
      RECT 22.44 3.54 22.655 3.758 ;
      RECT 22.455 3.535 22.65 3.768 ;
      RECT 22.475 3.532 22.64 3.805 ;
      RECT 22.475 3.531 22.63 3.805 ;
      RECT 22.5 3.53 22.63 3.805 ;
      RECT 22.06 3.775 22.32 4.035 ;
      RECT 21.935 3.82 22.32 4.03 ;
      RECT 21.925 3.825 22.32 4.025 ;
      RECT 21.94 4.765 21.955 5.075 ;
      RECT 20.535 4.535 20.545 4.665 ;
      RECT 20.315 4.53 20.42 4.665 ;
      RECT 20.23 4.535 20.28 4.665 ;
      RECT 18.78 3.27 18.785 4.375 ;
      RECT 22.035 4.857 22.04 4.993 ;
      RECT 22.03 4.852 22.035 5.053 ;
      RECT 22.025 4.85 22.03 5.066 ;
      RECT 22.01 4.847 22.025 5.068 ;
      RECT 22.005 4.842 22.01 5.07 ;
      RECT 22 4.838 22.005 5.073 ;
      RECT 21.985 4.833 22 5.075 ;
      RECT 21.955 4.825 21.985 5.075 ;
      RECT 21.916 4.765 21.94 5.075 ;
      RECT 21.83 4.765 21.916 5.072 ;
      RECT 21.8 4.765 21.83 5.065 ;
      RECT 21.775 4.765 21.8 5.058 ;
      RECT 21.75 4.765 21.775 5.05 ;
      RECT 21.735 4.765 21.75 5.043 ;
      RECT 21.71 4.765 21.735 5.035 ;
      RECT 21.695 4.765 21.71 5.028 ;
      RECT 21.655 4.775 21.695 5.017 ;
      RECT 21.645 4.77 21.655 5.007 ;
      RECT 21.641 4.769 21.645 5.004 ;
      RECT 21.555 4.761 21.641 4.987 ;
      RECT 21.522 4.75 21.555 4.964 ;
      RECT 21.436 4.739 21.522 4.942 ;
      RECT 21.35 4.723 21.436 4.911 ;
      RECT 21.28 4.708 21.35 4.883 ;
      RECT 21.27 4.701 21.28 4.87 ;
      RECT 21.24 4.698 21.27 4.86 ;
      RECT 21.215 4.694 21.24 4.853 ;
      RECT 21.2 4.691 21.215 4.848 ;
      RECT 21.195 4.69 21.2 4.843 ;
      RECT 21.165 4.685 21.195 4.836 ;
      RECT 21.16 4.68 21.165 4.831 ;
      RECT 21.145 4.677 21.16 4.826 ;
      RECT 21.14 4.672 21.145 4.821 ;
      RECT 21.12 4.667 21.14 4.818 ;
      RECT 21.105 4.662 21.12 4.81 ;
      RECT 21.09 4.656 21.105 4.805 ;
      RECT 21.06 4.647 21.09 4.798 ;
      RECT 21.055 4.64 21.06 4.79 ;
      RECT 21.05 4.638 21.055 4.788 ;
      RECT 21.045 4.637 21.05 4.785 ;
      RECT 21.005 4.63 21.045 4.778 ;
      RECT 20.991 4.62 21.005 4.768 ;
      RECT 20.94 4.609 20.991 4.756 ;
      RECT 20.915 4.595 20.94 4.742 ;
      RECT 20.89 4.584 20.915 4.734 ;
      RECT 20.87 4.573 20.89 4.728 ;
      RECT 20.86 4.567 20.87 4.723 ;
      RECT 20.855 4.565 20.86 4.719 ;
      RECT 20.835 4.56 20.855 4.714 ;
      RECT 20.805 4.55 20.835 4.704 ;
      RECT 20.8 4.542 20.805 4.697 ;
      RECT 20.785 4.54 20.8 4.693 ;
      RECT 20.765 4.54 20.785 4.688 ;
      RECT 20.76 4.539 20.765 4.686 ;
      RECT 20.755 4.539 20.76 4.683 ;
      RECT 20.715 4.538 20.755 4.678 ;
      RECT 20.69 4.537 20.715 4.673 ;
      RECT 20.63 4.536 20.69 4.67 ;
      RECT 20.545 4.535 20.63 4.668 ;
      RECT 20.506 4.534 20.535 4.665 ;
      RECT 20.42 4.532 20.506 4.665 ;
      RECT 20.28 4.532 20.315 4.665 ;
      RECT 20.19 4.536 20.23 4.668 ;
      RECT 20.175 4.539 20.19 4.675 ;
      RECT 20.165 4.54 20.175 4.682 ;
      RECT 20.14 4.543 20.165 4.687 ;
      RECT 20.135 4.545 20.14 4.69 ;
      RECT 20.085 4.547 20.135 4.691 ;
      RECT 20.046 4.551 20.085 4.693 ;
      RECT 19.96 4.553 20.046 4.696 ;
      RECT 19.942 4.555 19.96 4.698 ;
      RECT 19.856 4.558 19.942 4.7 ;
      RECT 19.77 4.562 19.856 4.703 ;
      RECT 19.733 4.566 19.77 4.706 ;
      RECT 19.647 4.569 19.733 4.709 ;
      RECT 19.561 4.573 19.647 4.712 ;
      RECT 19.475 4.578 19.561 4.716 ;
      RECT 19.455 4.58 19.475 4.719 ;
      RECT 19.435 4.579 19.455 4.72 ;
      RECT 19.386 4.576 19.435 4.721 ;
      RECT 19.3 4.571 19.386 4.724 ;
      RECT 19.25 4.566 19.3 4.726 ;
      RECT 19.226 4.564 19.25 4.727 ;
      RECT 19.14 4.559 19.226 4.729 ;
      RECT 19.115 4.555 19.14 4.728 ;
      RECT 19.105 4.552 19.115 4.726 ;
      RECT 19.095 4.545 19.105 4.723 ;
      RECT 19.09 4.525 19.095 4.718 ;
      RECT 19.08 4.495 19.09 4.713 ;
      RECT 19.065 4.365 19.08 4.704 ;
      RECT 19.06 4.357 19.065 4.697 ;
      RECT 19.04 4.35 19.06 4.689 ;
      RECT 19.035 4.332 19.04 4.681 ;
      RECT 19.025 4.312 19.035 4.676 ;
      RECT 19.02 4.285 19.025 4.672 ;
      RECT 19.015 4.262 19.02 4.669 ;
      RECT 18.995 4.22 19.015 4.661 ;
      RECT 18.96 4.135 18.995 4.645 ;
      RECT 18.955 4.067 18.96 4.633 ;
      RECT 18.94 4.037 18.955 4.627 ;
      RECT 18.935 3.282 18.94 3.528 ;
      RECT 18.925 4.007 18.94 4.618 ;
      RECT 18.93 3.277 18.935 3.56 ;
      RECT 18.925 3.272 18.93 3.603 ;
      RECT 18.92 3.27 18.925 3.638 ;
      RECT 18.905 3.97 18.925 4.608 ;
      RECT 18.915 3.27 18.92 3.675 ;
      RECT 18.9 3.27 18.915 3.773 ;
      RECT 18.9 3.943 18.905 4.601 ;
      RECT 18.895 3.27 18.9 3.848 ;
      RECT 18.895 3.931 18.9 4.598 ;
      RECT 18.89 3.27 18.895 3.88 ;
      RECT 18.89 3.91 18.895 4.595 ;
      RECT 18.885 3.27 18.89 4.592 ;
      RECT 18.85 3.27 18.885 4.578 ;
      RECT 18.835 3.27 18.85 4.56 ;
      RECT 18.815 3.27 18.835 4.55 ;
      RECT 18.79 3.27 18.815 4.533 ;
      RECT 18.785 3.27 18.79 4.483 ;
      RECT 18.775 3.27 18.78 4.313 ;
      RECT 18.77 3.27 18.775 4.22 ;
      RECT 18.765 3.27 18.77 4.133 ;
      RECT 18.76 3.27 18.765 4.065 ;
      RECT 18.755 3.27 18.76 4.008 ;
      RECT 18.745 3.27 18.755 3.903 ;
      RECT 18.74 3.27 18.745 3.775 ;
      RECT 18.735 3.27 18.74 3.693 ;
      RECT 18.73 3.272 18.735 3.61 ;
      RECT 18.725 3.277 18.73 3.543 ;
      RECT 18.72 3.282 18.725 3.47 ;
      RECT 21.535 3.6 21.795 3.86 ;
      RECT 21.555 3.567 21.765 3.86 ;
      RECT 21.555 3.565 21.755 3.86 ;
      RECT 21.565 3.552 21.755 3.86 ;
      RECT 21.565 3.55 21.68 3.86 ;
      RECT 21.04 3.675 21.215 3.955 ;
      RECT 21.035 3.675 21.215 3.953 ;
      RECT 21.035 3.675 21.23 3.95 ;
      RECT 21.025 3.675 21.23 3.948 ;
      RECT 20.97 3.675 21.23 3.935 ;
      RECT 20.97 3.75 21.235 3.913 ;
      RECT 20.5 4.873 20.505 5.08 ;
      RECT 20.45 4.867 20.5 5.079 ;
      RECT 20.417 4.881 20.51 5.078 ;
      RECT 20.331 4.881 20.51 5.077 ;
      RECT 20.245 4.881 20.51 5.076 ;
      RECT 20.245 4.98 20.515 5.073 ;
      RECT 20.24 4.98 20.515 5.068 ;
      RECT 20.235 4.98 20.515 5.05 ;
      RECT 20.23 4.98 20.515 5.033 ;
      RECT 20.19 4.765 20.45 5.025 ;
      RECT 19.65 3.915 19.736 4.329 ;
      RECT 19.65 3.915 19.775 4.326 ;
      RECT 19.65 3.915 19.795 4.316 ;
      RECT 19.605 3.915 19.795 4.313 ;
      RECT 19.605 4.067 19.805 4.303 ;
      RECT 19.605 4.088 19.81 4.297 ;
      RECT 19.605 4.106 19.815 4.293 ;
      RECT 19.605 4.126 19.825 4.288 ;
      RECT 19.58 4.126 19.825 4.285 ;
      RECT 19.57 4.126 19.825 4.263 ;
      RECT 19.57 4.142 19.83 4.233 ;
      RECT 19.535 3.915 19.795 4.22 ;
      RECT 19.535 4.154 19.835 4.175 ;
      RECT 16.545 10.06 16.835 10.29 ;
      RECT 16.605 9.315 16.775 10.29 ;
      RECT 16.515 9.315 16.865 9.605 ;
      RECT 16.14 8.575 16.49 8.865 ;
      RECT 16 8.61 16.49 8.78 ;
      RECT 93.47 7.25 93.82 7.54 ;
      RECT 83.16 4.56 83.42 4.82 ;
      RECT 78.21 7.25 78.56 7.54 ;
      RECT 67.9 4.56 68.16 4.82 ;
      RECT 62.95 7.25 63.3 7.54 ;
      RECT 52.64 4.56 52.9 4.82 ;
      RECT 47.69 7.25 48.04 7.54 ;
      RECT 37.38 4.56 37.64 4.82 ;
      RECT 32.43 7.25 32.78 7.54 ;
      RECT 22.12 4.56 22.38 4.82 ;
    LAYER mcon ;
      RECT 93.56 7.31 93.73 7.48 ;
      RECT 93.555 8.61 93.725 8.78 ;
      RECT 93.555 10.09 93.725 10.26 ;
      RECT 93.185 8.24 93.355 8.41 ;
      RECT 93.18 4.055 93.35 4.225 ;
      RECT 92.565 2.205 92.735 2.375 ;
      RECT 92.565 3.685 92.735 3.855 ;
      RECT 92.565 8.61 92.735 8.78 ;
      RECT 92.565 10.09 92.735 10.26 ;
      RECT 92.195 4.055 92.365 4.225 ;
      RECT 92.195 8.24 92.365 8.41 ;
      RECT 91.205 3.315 91.375 3.485 ;
      RECT 91.205 8.98 91.375 9.15 ;
      RECT 90.775 2.205 90.945 2.375 ;
      RECT 90.775 2.945 90.945 3.115 ;
      RECT 90.775 9.35 90.945 9.52 ;
      RECT 90.775 10.09 90.945 10.26 ;
      RECT 90.405 3.685 90.575 3.855 ;
      RECT 90.405 8.61 90.575 8.78 ;
      RECT 87.575 3.575 87.745 3.745 ;
      RECT 87.18 4.32 87.35 4.49 ;
      RECT 87.07 3.595 87.24 3.765 ;
      RECT 86.25 3.285 86.42 3.455 ;
      RECT 85.935 4.325 86.105 4.495 ;
      RECT 85.89 3.815 86.06 3.985 ;
      RECT 85.57 8.98 85.74 9.15 ;
      RECT 85.465 4.025 85.635 4.195 ;
      RECT 85.275 3.245 85.445 3.415 ;
      RECT 85.225 4.855 85.395 5.025 ;
      RECT 85.14 9.35 85.31 9.52 ;
      RECT 85.14 10.09 85.31 10.26 ;
      RECT 84.89 4.295 85.06 4.465 ;
      RECT 84.795 3.455 84.965 3.625 ;
      RECT 83.995 4.68 84.165 4.85 ;
      RECT 83.935 3.88 84.105 4.05 ;
      RECT 83.495 3.55 83.665 3.72 ;
      RECT 83.23 4.6 83.4 4.77 ;
      RECT 82.985 3.84 83.155 4.01 ;
      RECT 82.89 4.87 83.06 5.04 ;
      RECT 82.615 3.565 82.785 3.735 ;
      RECT 82.085 3.765 82.255 3.935 ;
      RECT 81.36 3.31 81.53 3.48 ;
      RECT 81.36 4.89 81.53 5.06 ;
      RECT 81.05 3.855 81.22 4.025 ;
      RECT 80.64 4.08 80.81 4.25 ;
      RECT 79.93 4.38 80.1 4.55 ;
      RECT 79.785 3.29 79.955 3.46 ;
      RECT 78.3 7.31 78.47 7.48 ;
      RECT 78.295 8.61 78.465 8.78 ;
      RECT 78.295 10.09 78.465 10.26 ;
      RECT 77.925 8.24 78.095 8.41 ;
      RECT 77.92 4.055 78.09 4.225 ;
      RECT 77.305 2.205 77.475 2.375 ;
      RECT 77.305 3.685 77.475 3.855 ;
      RECT 77.305 8.61 77.475 8.78 ;
      RECT 77.305 10.09 77.475 10.26 ;
      RECT 76.935 4.055 77.105 4.225 ;
      RECT 76.935 8.24 77.105 8.41 ;
      RECT 75.945 3.315 76.115 3.485 ;
      RECT 75.945 8.98 76.115 9.15 ;
      RECT 75.515 2.205 75.685 2.375 ;
      RECT 75.515 2.945 75.685 3.115 ;
      RECT 75.515 9.35 75.685 9.52 ;
      RECT 75.515 10.09 75.685 10.26 ;
      RECT 75.145 3.685 75.315 3.855 ;
      RECT 75.145 8.61 75.315 8.78 ;
      RECT 72.315 3.575 72.485 3.745 ;
      RECT 71.92 4.32 72.09 4.49 ;
      RECT 71.81 3.595 71.98 3.765 ;
      RECT 70.99 3.285 71.16 3.455 ;
      RECT 70.675 4.325 70.845 4.495 ;
      RECT 70.63 3.815 70.8 3.985 ;
      RECT 70.31 8.98 70.48 9.15 ;
      RECT 70.205 4.025 70.375 4.195 ;
      RECT 70.015 3.245 70.185 3.415 ;
      RECT 69.965 4.855 70.135 5.025 ;
      RECT 69.88 9.35 70.05 9.52 ;
      RECT 69.88 10.09 70.05 10.26 ;
      RECT 69.63 4.295 69.8 4.465 ;
      RECT 69.535 3.455 69.705 3.625 ;
      RECT 68.735 4.68 68.905 4.85 ;
      RECT 68.675 3.88 68.845 4.05 ;
      RECT 68.235 3.55 68.405 3.72 ;
      RECT 67.97 4.6 68.14 4.77 ;
      RECT 67.725 3.84 67.895 4.01 ;
      RECT 67.63 4.87 67.8 5.04 ;
      RECT 67.355 3.565 67.525 3.735 ;
      RECT 66.825 3.765 66.995 3.935 ;
      RECT 66.1 3.31 66.27 3.48 ;
      RECT 66.1 4.89 66.27 5.06 ;
      RECT 65.79 3.855 65.96 4.025 ;
      RECT 65.38 4.08 65.55 4.25 ;
      RECT 64.67 4.38 64.84 4.55 ;
      RECT 64.525 3.29 64.695 3.46 ;
      RECT 63.04 7.31 63.21 7.48 ;
      RECT 63.035 8.61 63.205 8.78 ;
      RECT 63.035 10.09 63.205 10.26 ;
      RECT 62.665 8.24 62.835 8.41 ;
      RECT 62.66 4.055 62.83 4.225 ;
      RECT 62.045 2.205 62.215 2.375 ;
      RECT 62.045 3.685 62.215 3.855 ;
      RECT 62.045 8.61 62.215 8.78 ;
      RECT 62.045 10.09 62.215 10.26 ;
      RECT 61.675 4.055 61.845 4.225 ;
      RECT 61.675 8.24 61.845 8.41 ;
      RECT 60.685 3.315 60.855 3.485 ;
      RECT 60.685 8.98 60.855 9.15 ;
      RECT 60.255 2.205 60.425 2.375 ;
      RECT 60.255 2.945 60.425 3.115 ;
      RECT 60.255 9.35 60.425 9.52 ;
      RECT 60.255 10.09 60.425 10.26 ;
      RECT 59.885 3.685 60.055 3.855 ;
      RECT 59.885 8.61 60.055 8.78 ;
      RECT 57.055 3.575 57.225 3.745 ;
      RECT 56.66 4.32 56.83 4.49 ;
      RECT 56.55 3.595 56.72 3.765 ;
      RECT 55.73 3.285 55.9 3.455 ;
      RECT 55.415 4.325 55.585 4.495 ;
      RECT 55.37 3.815 55.54 3.985 ;
      RECT 55.05 8.98 55.22 9.15 ;
      RECT 54.945 4.025 55.115 4.195 ;
      RECT 54.755 3.245 54.925 3.415 ;
      RECT 54.705 4.855 54.875 5.025 ;
      RECT 54.62 9.35 54.79 9.52 ;
      RECT 54.62 10.09 54.79 10.26 ;
      RECT 54.37 4.295 54.54 4.465 ;
      RECT 54.275 3.455 54.445 3.625 ;
      RECT 53.475 4.68 53.645 4.85 ;
      RECT 53.415 3.88 53.585 4.05 ;
      RECT 52.975 3.55 53.145 3.72 ;
      RECT 52.71 4.6 52.88 4.77 ;
      RECT 52.465 3.84 52.635 4.01 ;
      RECT 52.37 4.87 52.54 5.04 ;
      RECT 52.095 3.565 52.265 3.735 ;
      RECT 51.565 3.765 51.735 3.935 ;
      RECT 50.84 3.31 51.01 3.48 ;
      RECT 50.84 4.89 51.01 5.06 ;
      RECT 50.53 3.855 50.7 4.025 ;
      RECT 50.12 4.08 50.29 4.25 ;
      RECT 49.41 4.38 49.58 4.55 ;
      RECT 49.265 3.29 49.435 3.46 ;
      RECT 47.78 7.31 47.95 7.48 ;
      RECT 47.775 8.61 47.945 8.78 ;
      RECT 47.775 10.09 47.945 10.26 ;
      RECT 47.405 8.24 47.575 8.41 ;
      RECT 47.4 4.055 47.57 4.225 ;
      RECT 46.785 2.205 46.955 2.375 ;
      RECT 46.785 3.685 46.955 3.855 ;
      RECT 46.785 8.61 46.955 8.78 ;
      RECT 46.785 10.09 46.955 10.26 ;
      RECT 46.415 4.055 46.585 4.225 ;
      RECT 46.415 8.24 46.585 8.41 ;
      RECT 45.425 3.315 45.595 3.485 ;
      RECT 45.425 8.98 45.595 9.15 ;
      RECT 44.995 2.205 45.165 2.375 ;
      RECT 44.995 2.945 45.165 3.115 ;
      RECT 44.995 9.35 45.165 9.52 ;
      RECT 44.995 10.09 45.165 10.26 ;
      RECT 44.625 3.685 44.795 3.855 ;
      RECT 44.625 8.61 44.795 8.78 ;
      RECT 41.795 3.575 41.965 3.745 ;
      RECT 41.4 4.32 41.57 4.49 ;
      RECT 41.29 3.595 41.46 3.765 ;
      RECT 40.47 3.285 40.64 3.455 ;
      RECT 40.155 4.325 40.325 4.495 ;
      RECT 40.11 3.815 40.28 3.985 ;
      RECT 39.79 8.98 39.96 9.15 ;
      RECT 39.685 4.025 39.855 4.195 ;
      RECT 39.495 3.245 39.665 3.415 ;
      RECT 39.445 4.855 39.615 5.025 ;
      RECT 39.36 9.35 39.53 9.52 ;
      RECT 39.36 10.09 39.53 10.26 ;
      RECT 39.11 4.295 39.28 4.465 ;
      RECT 39.015 3.455 39.185 3.625 ;
      RECT 38.215 4.68 38.385 4.85 ;
      RECT 38.155 3.88 38.325 4.05 ;
      RECT 37.715 3.55 37.885 3.72 ;
      RECT 37.45 4.6 37.62 4.77 ;
      RECT 37.205 3.84 37.375 4.01 ;
      RECT 37.11 4.87 37.28 5.04 ;
      RECT 36.835 3.565 37.005 3.735 ;
      RECT 36.305 3.765 36.475 3.935 ;
      RECT 35.58 3.31 35.75 3.48 ;
      RECT 35.58 4.89 35.75 5.06 ;
      RECT 35.27 3.855 35.44 4.025 ;
      RECT 34.86 4.08 35.03 4.25 ;
      RECT 34.15 4.38 34.32 4.55 ;
      RECT 34.005 3.29 34.175 3.46 ;
      RECT 32.52 7.31 32.69 7.48 ;
      RECT 32.515 8.61 32.685 8.78 ;
      RECT 32.515 10.09 32.685 10.26 ;
      RECT 32.145 8.24 32.315 8.41 ;
      RECT 32.14 4.055 32.31 4.225 ;
      RECT 31.525 2.205 31.695 2.375 ;
      RECT 31.525 3.685 31.695 3.855 ;
      RECT 31.525 8.61 31.695 8.78 ;
      RECT 31.525 10.09 31.695 10.26 ;
      RECT 31.155 4.055 31.325 4.225 ;
      RECT 31.155 8.24 31.325 8.41 ;
      RECT 30.165 3.315 30.335 3.485 ;
      RECT 30.165 8.98 30.335 9.15 ;
      RECT 29.735 2.205 29.905 2.375 ;
      RECT 29.735 2.945 29.905 3.115 ;
      RECT 29.735 9.35 29.905 9.52 ;
      RECT 29.735 10.09 29.905 10.26 ;
      RECT 29.365 3.685 29.535 3.855 ;
      RECT 29.365 8.61 29.535 8.78 ;
      RECT 26.535 3.575 26.705 3.745 ;
      RECT 26.14 4.32 26.31 4.49 ;
      RECT 26.03 3.595 26.2 3.765 ;
      RECT 25.21 3.285 25.38 3.455 ;
      RECT 24.895 4.325 25.065 4.495 ;
      RECT 24.85 3.815 25.02 3.985 ;
      RECT 24.53 8.98 24.7 9.15 ;
      RECT 24.425 4.025 24.595 4.195 ;
      RECT 24.235 3.245 24.405 3.415 ;
      RECT 24.185 4.855 24.355 5.025 ;
      RECT 24.1 9.35 24.27 9.52 ;
      RECT 24.1 10.09 24.27 10.26 ;
      RECT 23.85 4.295 24.02 4.465 ;
      RECT 23.755 3.455 23.925 3.625 ;
      RECT 22.955 4.68 23.125 4.85 ;
      RECT 22.895 3.88 23.065 4.05 ;
      RECT 22.455 3.55 22.625 3.72 ;
      RECT 22.19 4.6 22.36 4.77 ;
      RECT 21.945 3.84 22.115 4.01 ;
      RECT 21.85 4.87 22.02 5.04 ;
      RECT 21.575 3.565 21.745 3.735 ;
      RECT 21.045 3.765 21.215 3.935 ;
      RECT 20.32 3.31 20.49 3.48 ;
      RECT 20.32 4.89 20.49 5.06 ;
      RECT 20.01 3.855 20.18 4.025 ;
      RECT 19.6 4.08 19.77 4.25 ;
      RECT 18.89 4.38 19.06 4.55 ;
      RECT 18.745 3.29 18.915 3.46 ;
      RECT 16.605 9.35 16.775 9.52 ;
      RECT 16.605 10.09 16.775 10.26 ;
      RECT 16.235 8.61 16.405 8.78 ;
    LAYER li1 ;
      RECT 93.555 7.31 93.725 8.78 ;
      RECT 93.555 7.31 93.73 8.57 ;
      RECT 93.185 9.26 93.655 9.43 ;
      RECT 93.185 8.24 93.355 9.43 ;
      RECT 93.18 3.035 93.35 4.225 ;
      RECT 93.18 3.035 93.65 3.205 ;
      RECT 92.565 3.895 92.74 5.155 ;
      RECT 92.565 3.685 92.735 5.155 ;
      RECT 92.565 7.31 92.735 8.78 ;
      RECT 92.565 7.31 92.74 8.57 ;
      RECT 92.195 3.035 92.365 4.225 ;
      RECT 92.195 3.035 92.665 3.205 ;
      RECT 92.195 9.26 92.665 9.43 ;
      RECT 92.195 8.24 92.365 9.43 ;
      RECT 91.205 4.015 91.38 5.155 ;
      RECT 91.205 1.865 91.375 5.155 ;
      RECT 91.205 1.865 91.38 2.415 ;
      RECT 91.205 10.05 91.38 10.6 ;
      RECT 91.205 7.31 91.375 10.6 ;
      RECT 91.205 7.31 91.38 8.45 ;
      RECT 90.775 3.895 90.95 5.155 ;
      RECT 90.775 2.945 90.945 5.155 ;
      RECT 90.775 7.31 90.945 9.52 ;
      RECT 90.775 7.31 90.95 8.57 ;
      RECT 90.345 3.925 90.515 5.155 ;
      RECT 90.405 2.145 90.575 4.095 ;
      RECT 90.345 1.865 90.515 2.315 ;
      RECT 90.345 10.15 90.515 10.6 ;
      RECT 90.405 8.37 90.575 10.32 ;
      RECT 90.345 7.31 90.515 8.54 ;
      RECT 89.82 3.895 89.995 5.155 ;
      RECT 89.82 1.865 89.99 5.155 ;
      RECT 89.82 3.365 90.23 3.695 ;
      RECT 89.82 2.525 90.23 2.855 ;
      RECT 89.82 1.865 89.995 2.355 ;
      RECT 89.82 10.11 89.995 10.6 ;
      RECT 89.82 7.31 89.99 10.6 ;
      RECT 89.82 9.61 90.23 9.94 ;
      RECT 89.82 8.77 90.23 9.1 ;
      RECT 89.82 7.31 89.995 8.57 ;
      RECT 87.75 4.421 87.755 4.593 ;
      RECT 87.745 4.414 87.75 4.683 ;
      RECT 87.74 4.408 87.745 4.702 ;
      RECT 87.72 4.402 87.74 4.712 ;
      RECT 87.705 4.397 87.72 4.72 ;
      RECT 87.668 4.391 87.705 4.718 ;
      RECT 87.582 4.377 87.668 4.714 ;
      RECT 87.496 4.359 87.582 4.709 ;
      RECT 87.41 4.34 87.496 4.703 ;
      RECT 87.38 4.328 87.41 4.699 ;
      RECT 87.36 4.322 87.38 4.698 ;
      RECT 87.295 4.32 87.36 4.696 ;
      RECT 87.28 4.32 87.295 4.688 ;
      RECT 87.265 4.32 87.28 4.675 ;
      RECT 87.26 4.32 87.265 4.665 ;
      RECT 87.245 4.32 87.26 4.643 ;
      RECT 87.23 4.32 87.245 4.61 ;
      RECT 87.225 4.32 87.23 4.588 ;
      RECT 87.215 4.32 87.225 4.57 ;
      RECT 87.2 4.32 87.215 4.548 ;
      RECT 87.18 4.32 87.2 4.51 ;
      RECT 87.53 3.605 87.565 4.044 ;
      RECT 87.53 3.605 87.57 4.043 ;
      RECT 87.475 3.665 87.57 4.042 ;
      RECT 87.34 3.837 87.57 4.041 ;
      RECT 87.45 3.715 87.57 4.041 ;
      RECT 87.34 3.837 87.595 4.031 ;
      RECT 87.395 3.782 87.675 3.948 ;
      RECT 87.57 3.576 87.575 4.039 ;
      RECT 87.425 3.752 87.715 3.825 ;
      RECT 87.44 3.735 87.57 4.041 ;
      RECT 87.575 3.575 87.745 3.763 ;
      RECT 87.565 3.578 87.745 3.763 ;
      RECT 87.07 3.455 87.24 3.765 ;
      RECT 87.07 3.455 87.245 3.738 ;
      RECT 87.07 3.455 87.25 3.715 ;
      RECT 87.07 3.455 87.26 3.665 ;
      RECT 87.065 3.56 87.26 3.635 ;
      RECT 87.1 3.13 87.27 3.608 ;
      RECT 87.1 3.13 87.285 3.529 ;
      RECT 87.09 3.34 87.285 3.529 ;
      RECT 87.1 3.14 87.295 3.444 ;
      RECT 87.03 3.882 87.035 4.085 ;
      RECT 87.02 3.87 87.03 4.195 ;
      RECT 86.995 3.87 87.02 4.235 ;
      RECT 86.915 3.87 86.995 4.32 ;
      RECT 86.905 3.87 86.915 4.39 ;
      RECT 86.88 3.87 86.905 4.413 ;
      RECT 86.86 3.87 86.88 4.448 ;
      RECT 86.815 3.88 86.86 4.491 ;
      RECT 86.805 3.892 86.815 4.528 ;
      RECT 86.785 3.906 86.805 4.548 ;
      RECT 86.775 3.924 86.785 4.564 ;
      RECT 86.76 3.95 86.775 4.574 ;
      RECT 86.745 3.991 86.76 4.588 ;
      RECT 86.735 4.026 86.745 4.598 ;
      RECT 86.73 4.042 86.735 4.603 ;
      RECT 86.72 4.057 86.73 4.608 ;
      RECT 86.7 4.1 86.72 4.618 ;
      RECT 86.68 4.137 86.7 4.631 ;
      RECT 86.645 4.16 86.68 4.649 ;
      RECT 86.635 4.174 86.645 4.665 ;
      RECT 86.615 4.184 86.635 4.675 ;
      RECT 86.61 4.193 86.615 4.683 ;
      RECT 86.6 4.2 86.61 4.69 ;
      RECT 86.59 4.207 86.6 4.698 ;
      RECT 86.575 4.217 86.59 4.706 ;
      RECT 86.565 4.231 86.575 4.716 ;
      RECT 86.555 4.243 86.565 4.728 ;
      RECT 86.54 4.265 86.555 4.741 ;
      RECT 86.53 4.287 86.54 4.752 ;
      RECT 86.52 4.307 86.53 4.761 ;
      RECT 86.515 4.322 86.52 4.768 ;
      RECT 86.485 4.355 86.515 4.782 ;
      RECT 86.475 4.39 86.485 4.797 ;
      RECT 86.47 4.397 86.475 4.803 ;
      RECT 86.45 4.412 86.47 4.81 ;
      RECT 86.445 4.427 86.45 4.818 ;
      RECT 86.44 4.436 86.445 4.823 ;
      RECT 86.425 4.442 86.44 4.83 ;
      RECT 86.42 4.448 86.425 4.838 ;
      RECT 86.415 4.452 86.42 4.845 ;
      RECT 86.41 4.456 86.415 4.855 ;
      RECT 86.4 4.461 86.41 4.865 ;
      RECT 86.38 4.472 86.4 4.893 ;
      RECT 86.365 4.484 86.38 4.92 ;
      RECT 86.345 4.497 86.365 4.945 ;
      RECT 86.325 4.512 86.345 4.969 ;
      RECT 86.31 4.527 86.325 4.984 ;
      RECT 86.305 4.538 86.31 4.993 ;
      RECT 86.24 4.583 86.305 5.003 ;
      RECT 86.205 4.642 86.24 5.016 ;
      RECT 86.2 4.665 86.205 5.022 ;
      RECT 86.195 4.672 86.2 5.024 ;
      RECT 86.18 4.682 86.195 5.027 ;
      RECT 86.15 4.707 86.18 5.031 ;
      RECT 86.145 4.725 86.15 5.035 ;
      RECT 86.14 4.732 86.145 5.036 ;
      RECT 86.12 4.74 86.14 5.04 ;
      RECT 86.11 4.747 86.12 5.044 ;
      RECT 86.066 4.758 86.11 5.051 ;
      RECT 85.98 4.786 86.066 5.067 ;
      RECT 85.92 4.81 85.98 5.085 ;
      RECT 85.875 4.82 85.92 5.099 ;
      RECT 85.816 4.828 85.875 5.113 ;
      RECT 85.73 4.835 85.816 5.132 ;
      RECT 85.705 4.84 85.73 5.147 ;
      RECT 85.625 4.843 85.705 5.15 ;
      RECT 85.545 4.847 85.625 5.137 ;
      RECT 85.536 4.85 85.545 5.122 ;
      RECT 85.45 4.85 85.536 5.107 ;
      RECT 85.39 4.852 85.45 5.084 ;
      RECT 85.386 4.855 85.39 5.074 ;
      RECT 85.3 4.855 85.386 5.059 ;
      RECT 85.225 4.855 85.3 5.035 ;
      RECT 86.54 3.864 86.55 4.04 ;
      RECT 86.495 3.831 86.54 4.04 ;
      RECT 86.45 3.782 86.495 4.04 ;
      RECT 86.42 3.752 86.45 4.041 ;
      RECT 86.415 3.735 86.42 4.042 ;
      RECT 86.39 3.715 86.415 4.043 ;
      RECT 86.375 3.69 86.39 4.044 ;
      RECT 86.37 3.677 86.375 4.045 ;
      RECT 86.365 3.671 86.37 4.043 ;
      RECT 86.36 3.663 86.365 4.037 ;
      RECT 86.335 3.655 86.36 4.017 ;
      RECT 86.315 3.644 86.335 3.988 ;
      RECT 86.285 3.629 86.315 3.959 ;
      RECT 86.265 3.615 86.285 3.931 ;
      RECT 86.255 3.609 86.265 3.91 ;
      RECT 86.25 3.606 86.255 3.893 ;
      RECT 86.245 3.603 86.25 3.878 ;
      RECT 86.23 3.598 86.245 3.843 ;
      RECT 86.225 3.594 86.23 3.81 ;
      RECT 86.205 3.589 86.225 3.786 ;
      RECT 86.175 3.581 86.205 3.751 ;
      RECT 86.16 3.575 86.175 3.728 ;
      RECT 86.12 3.568 86.16 3.713 ;
      RECT 86.095 3.56 86.12 3.693 ;
      RECT 86.075 3.555 86.095 3.683 ;
      RECT 86.04 3.549 86.075 3.678 ;
      RECT 85.995 3.54 86.04 3.677 ;
      RECT 85.965 3.536 85.995 3.679 ;
      RECT 85.88 3.544 85.965 3.683 ;
      RECT 85.81 3.555 85.88 3.705 ;
      RECT 85.797 3.561 85.81 3.728 ;
      RECT 85.711 3.568 85.797 3.75 ;
      RECT 85.625 3.58 85.711 3.787 ;
      RECT 85.625 3.957 85.635 4.195 ;
      RECT 85.62 3.586 85.625 3.81 ;
      RECT 85.615 3.842 85.625 4.195 ;
      RECT 85.615 3.587 85.62 3.815 ;
      RECT 85.61 3.588 85.615 4.195 ;
      RECT 85.586 3.59 85.61 4.196 ;
      RECT 85.5 3.598 85.586 4.198 ;
      RECT 85.48 3.612 85.5 4.201 ;
      RECT 85.475 3.64 85.48 4.202 ;
      RECT 85.47 3.652 85.475 4.203 ;
      RECT 85.465 3.667 85.47 4.204 ;
      RECT 85.455 3.697 85.465 4.205 ;
      RECT 85.45 3.735 85.455 4.203 ;
      RECT 85.445 3.755 85.45 4.198 ;
      RECT 85.43 3.79 85.445 4.183 ;
      RECT 85.42 3.842 85.43 4.163 ;
      RECT 85.415 3.872 85.42 4.151 ;
      RECT 85.4 3.885 85.415 4.134 ;
      RECT 85.375 3.889 85.4 4.101 ;
      RECT 85.36 3.887 85.375 4.078 ;
      RECT 85.345 3.886 85.36 4.075 ;
      RECT 85.285 3.884 85.345 4.073 ;
      RECT 85.275 3.882 85.285 4.068 ;
      RECT 85.235 3.881 85.275 4.065 ;
      RECT 85.165 3.878 85.235 4.063 ;
      RECT 85.11 3.876 85.165 4.058 ;
      RECT 85.04 3.87 85.11 4.053 ;
      RECT 85.031 3.87 85.04 4.05 ;
      RECT 84.945 3.87 85.031 4.045 ;
      RECT 84.94 3.87 84.945 4.04 ;
      RECT 86.245 3.105 86.42 3.455 ;
      RECT 86.245 3.12 86.43 3.453 ;
      RECT 86.22 3.07 86.365 3.45 ;
      RECT 86.2 3.071 86.365 3.443 ;
      RECT 86.19 3.072 86.375 3.438 ;
      RECT 86.16 3.073 86.375 3.425 ;
      RECT 86.11 3.074 86.375 3.401 ;
      RECT 86.105 3.076 86.375 3.386 ;
      RECT 86.105 3.142 86.435 3.38 ;
      RECT 86.085 3.083 86.39 3.36 ;
      RECT 86.075 3.092 86.4 3.215 ;
      RECT 86.085 3.087 86.4 3.36 ;
      RECT 86.105 3.077 86.39 3.386 ;
      RECT 85.69 4.402 85.86 4.69 ;
      RECT 85.685 4.42 85.87 4.685 ;
      RECT 85.65 4.428 85.935 4.605 ;
      RECT 85.65 4.428 86.021 4.595 ;
      RECT 85.65 4.428 86.075 4.541 ;
      RECT 85.935 4.325 86.105 4.509 ;
      RECT 85.65 4.48 86.11 4.497 ;
      RECT 85.635 4.45 86.105 4.493 ;
      RECT 85.895 4.332 85.935 4.644 ;
      RECT 85.775 4.369 86.105 4.509 ;
      RECT 85.87 4.344 85.895 4.67 ;
      RECT 85.86 4.351 86.105 4.509 ;
      RECT 85.991 3.815 86.06 4.074 ;
      RECT 85.991 3.87 86.065 4.073 ;
      RECT 85.905 3.87 86.065 4.072 ;
      RECT 85.9 3.87 86.07 4.065 ;
      RECT 85.89 3.815 86.06 4.06 ;
      RECT 85.57 10.05 85.745 10.6 ;
      RECT 85.57 7.31 85.74 10.6 ;
      RECT 85.57 7.31 85.745 8.45 ;
      RECT 85.27 3.114 85.445 3.415 ;
      RECT 85.255 3.102 85.27 3.4 ;
      RECT 85.225 3.101 85.255 3.353 ;
      RECT 85.225 3.119 85.45 3.348 ;
      RECT 85.21 3.103 85.27 3.313 ;
      RECT 85.205 3.125 85.46 3.213 ;
      RECT 85.205 3.108 85.356 3.213 ;
      RECT 85.205 3.11 85.36 3.213 ;
      RECT 85.21 3.106 85.356 3.313 ;
      RECT 85.315 4.342 85.32 4.69 ;
      RECT 85.305 4.332 85.315 4.696 ;
      RECT 85.27 4.322 85.305 4.698 ;
      RECT 85.232 4.317 85.27 4.702 ;
      RECT 85.146 4.31 85.232 4.709 ;
      RECT 85.06 4.3 85.146 4.719 ;
      RECT 85.015 4.295 85.06 4.727 ;
      RECT 85.011 4.295 85.015 4.731 ;
      RECT 84.925 4.295 85.011 4.738 ;
      RECT 84.91 4.295 84.925 4.738 ;
      RECT 84.9 4.293 84.91 4.71 ;
      RECT 84.89 4.289 84.9 4.653 ;
      RECT 84.87 4.283 84.89 4.585 ;
      RECT 84.865 4.279 84.87 4.533 ;
      RECT 84.855 4.278 84.865 4.5 ;
      RECT 84.805 4.276 84.855 4.485 ;
      RECT 84.78 4.274 84.805 4.48 ;
      RECT 84.737 4.272 84.78 4.476 ;
      RECT 84.651 4.268 84.737 4.464 ;
      RECT 84.565 4.263 84.651 4.448 ;
      RECT 84.535 4.26 84.565 4.435 ;
      RECT 84.51 4.259 84.535 4.423 ;
      RECT 84.505 4.259 84.51 4.413 ;
      RECT 84.465 4.258 84.505 4.405 ;
      RECT 84.45 4.257 84.465 4.398 ;
      RECT 84.4 4.256 84.45 4.39 ;
      RECT 84.398 4.255 84.4 4.385 ;
      RECT 84.312 4.253 84.398 4.385 ;
      RECT 84.226 4.248 84.312 4.385 ;
      RECT 84.14 4.244 84.226 4.385 ;
      RECT 84.091 4.24 84.14 4.383 ;
      RECT 84.005 4.237 84.091 4.378 ;
      RECT 83.982 4.234 84.005 4.374 ;
      RECT 83.896 4.231 83.982 4.369 ;
      RECT 83.81 4.227 83.896 4.36 ;
      RECT 83.785 4.22 83.81 4.355 ;
      RECT 83.725 4.185 83.785 4.352 ;
      RECT 83.705 4.11 83.725 4.349 ;
      RECT 83.7 4.052 83.705 4.348 ;
      RECT 83.675 3.992 83.7 4.347 ;
      RECT 83.6 3.87 83.675 4.343 ;
      RECT 83.59 3.87 83.6 4.335 ;
      RECT 83.575 3.87 83.59 4.325 ;
      RECT 83.56 3.87 83.575 4.295 ;
      RECT 83.545 3.87 83.56 4.24 ;
      RECT 83.53 3.87 83.545 4.178 ;
      RECT 83.505 3.87 83.53 4.103 ;
      RECT 83.5 3.87 83.505 4.053 ;
      RECT 85.14 7.31 85.31 9.52 ;
      RECT 85.14 7.31 85.315 8.57 ;
      RECT 84.845 3.415 84.865 3.724 ;
      RECT 84.831 3.417 84.88 3.721 ;
      RECT 84.831 3.422 84.9 3.712 ;
      RECT 84.745 3.42 84.88 3.706 ;
      RECT 84.745 3.428 84.935 3.689 ;
      RECT 84.71 3.43 84.935 3.688 ;
      RECT 84.68 3.438 84.935 3.679 ;
      RECT 84.67 3.443 84.955 3.665 ;
      RECT 84.71 3.433 84.955 3.665 ;
      RECT 84.71 3.436 84.965 3.653 ;
      RECT 84.68 3.438 84.975 3.64 ;
      RECT 84.68 3.442 84.985 3.583 ;
      RECT 84.67 3.447 84.99 3.498 ;
      RECT 84.831 3.415 84.865 3.721 ;
      RECT 84.27 3.518 84.275 3.73 ;
      RECT 84.145 3.515 84.16 3.73 ;
      RECT 83.61 3.545 83.68 3.73 ;
      RECT 83.495 3.545 83.53 3.725 ;
      RECT 84.616 3.847 84.635 4.041 ;
      RECT 84.53 3.802 84.616 4.042 ;
      RECT 84.52 3.755 84.53 4.044 ;
      RECT 84.515 3.735 84.52 4.045 ;
      RECT 84.495 3.7 84.515 4.046 ;
      RECT 84.48 3.65 84.495 4.047 ;
      RECT 84.46 3.587 84.48 4.048 ;
      RECT 84.45 3.55 84.46 4.049 ;
      RECT 84.435 3.539 84.45 4.05 ;
      RECT 84.43 3.531 84.435 4.048 ;
      RECT 84.42 3.53 84.43 4.04 ;
      RECT 84.39 3.527 84.42 4.019 ;
      RECT 84.315 3.522 84.39 3.964 ;
      RECT 84.3 3.518 84.315 3.91 ;
      RECT 84.29 3.518 84.3 3.805 ;
      RECT 84.275 3.518 84.29 3.738 ;
      RECT 84.26 3.518 84.27 3.728 ;
      RECT 84.205 3.517 84.26 3.725 ;
      RECT 84.16 3.515 84.205 3.728 ;
      RECT 84.132 3.515 84.145 3.731 ;
      RECT 84.046 3.519 84.132 3.733 ;
      RECT 83.96 3.525 84.046 3.738 ;
      RECT 83.94 3.529 83.96 3.74 ;
      RECT 83.938 3.53 83.94 3.739 ;
      RECT 83.852 3.532 83.938 3.738 ;
      RECT 83.766 3.537 83.852 3.735 ;
      RECT 83.68 3.542 83.766 3.732 ;
      RECT 83.53 3.545 83.61 3.728 ;
      RECT 84.185 10.11 84.36 10.6 ;
      RECT 84.185 7.31 84.355 10.6 ;
      RECT 84.185 9.61 84.595 9.94 ;
      RECT 84.185 8.77 84.595 9.1 ;
      RECT 84.185 7.31 84.36 8.57 ;
      RECT 84.306 4.52 84.355 4.854 ;
      RECT 84.306 4.52 84.36 4.853 ;
      RECT 84.22 4.52 84.36 4.852 ;
      RECT 83.995 4.628 84.365 4.85 ;
      RECT 84.22 4.52 84.39 4.843 ;
      RECT 84.19 4.532 84.395 4.834 ;
      RECT 84.175 4.55 84.4 4.831 ;
      RECT 83.99 4.634 84.4 4.758 ;
      RECT 83.985 4.641 84.4 4.718 ;
      RECT 84 4.607 84.4 4.831 ;
      RECT 84.161 4.553 84.365 4.85 ;
      RECT 84.075 4.573 84.4 4.831 ;
      RECT 84.175 4.547 84.395 4.834 ;
      RECT 83.945 3.871 84.135 4.065 ;
      RECT 83.94 3.873 84.135 4.064 ;
      RECT 83.935 3.877 84.15 4.061 ;
      RECT 83.95 3.87 84.15 4.061 ;
      RECT 83.935 3.98 84.155 4.056 ;
      RECT 83.23 4.48 83.321 4.778 ;
      RECT 83.225 4.482 83.4 4.773 ;
      RECT 83.23 4.48 83.4 4.773 ;
      RECT 83.225 4.486 83.42 4.771 ;
      RECT 83.225 4.541 83.46 4.77 ;
      RECT 83.225 4.576 83.475 4.764 ;
      RECT 83.225 4.61 83.485 4.754 ;
      RECT 83.215 4.49 83.42 4.605 ;
      RECT 83.215 4.51 83.435 4.605 ;
      RECT 83.215 4.493 83.425 4.605 ;
      RECT 83.44 3.261 83.445 3.323 ;
      RECT 83.435 3.183 83.44 3.346 ;
      RECT 83.43 3.14 83.435 3.357 ;
      RECT 83.425 3.13 83.43 3.369 ;
      RECT 83.42 3.13 83.425 3.378 ;
      RECT 83.395 3.13 83.42 3.41 ;
      RECT 83.39 3.13 83.395 3.443 ;
      RECT 83.375 3.13 83.39 3.468 ;
      RECT 83.365 3.13 83.375 3.495 ;
      RECT 83.36 3.13 83.365 3.508 ;
      RECT 83.355 3.13 83.36 3.523 ;
      RECT 83.345 3.13 83.355 3.538 ;
      RECT 83.34 3.13 83.345 3.558 ;
      RECT 83.315 3.13 83.34 3.593 ;
      RECT 83.27 3.13 83.315 3.638 ;
      RECT 83.26 3.13 83.27 3.651 ;
      RECT 83.175 3.215 83.26 3.658 ;
      RECT 83.14 3.337 83.175 3.667 ;
      RECT 83.135 3.377 83.14 3.671 ;
      RECT 83.115 3.4 83.135 3.673 ;
      RECT 83.11 3.43 83.115 3.676 ;
      RECT 83.1 3.442 83.11 3.677 ;
      RECT 83.055 3.465 83.1 3.682 ;
      RECT 83.015 3.495 83.055 3.69 ;
      RECT 82.98 3.507 83.015 3.696 ;
      RECT 82.975 3.512 82.98 3.7 ;
      RECT 82.905 3.522 82.975 3.707 ;
      RECT 82.865 3.532 82.905 3.717 ;
      RECT 82.845 3.537 82.865 3.723 ;
      RECT 82.835 3.541 82.845 3.728 ;
      RECT 82.83 3.544 82.835 3.731 ;
      RECT 82.82 3.545 82.83 3.732 ;
      RECT 82.795 3.547 82.82 3.736 ;
      RECT 82.785 3.552 82.795 3.739 ;
      RECT 82.74 3.56 82.785 3.74 ;
      RECT 82.615 3.565 82.74 3.74 ;
      RECT 83.17 3.862 83.19 4.044 ;
      RECT 83.121 3.847 83.17 4.043 ;
      RECT 83.035 3.862 83.19 4.041 ;
      RECT 83.02 3.862 83.19 4.04 ;
      RECT 82.985 3.84 83.155 4.025 ;
      RECT 83.055 4.86 83.07 5.069 ;
      RECT 83.055 4.868 83.075 5.068 ;
      RECT 83 4.868 83.075 5.067 ;
      RECT 82.98 4.872 83.08 5.065 ;
      RECT 82.96 4.822 83 5.064 ;
      RECT 82.905 4.88 83.085 5.062 ;
      RECT 82.87 4.837 83 5.06 ;
      RECT 82.866 4.84 83.055 5.059 ;
      RECT 82.78 4.848 83.055 5.057 ;
      RECT 82.78 4.892 83.09 5.05 ;
      RECT 82.77 4.985 83.09 5.048 ;
      RECT 82.78 4.904 83.095 5.033 ;
      RECT 82.78 4.925 83.11 5.003 ;
      RECT 82.78 4.952 83.115 4.973 ;
      RECT 82.905 4.83 83 5.062 ;
      RECT 82.535 3.875 82.54 4.413 ;
      RECT 82.34 4.205 82.345 4.4 ;
      RECT 80.64 3.87 80.655 4.25 ;
      RECT 82.705 3.87 82.71 4.04 ;
      RECT 82.7 3.87 82.705 4.05 ;
      RECT 82.695 3.87 82.7 4.063 ;
      RECT 82.67 3.87 82.695 4.105 ;
      RECT 82.645 3.87 82.67 4.178 ;
      RECT 82.63 3.87 82.645 4.23 ;
      RECT 82.625 3.87 82.63 4.26 ;
      RECT 82.6 3.87 82.625 4.3 ;
      RECT 82.585 3.87 82.6 4.355 ;
      RECT 82.58 3.87 82.585 4.388 ;
      RECT 82.555 3.87 82.58 4.408 ;
      RECT 82.54 3.87 82.555 4.414 ;
      RECT 82.47 3.905 82.535 4.41 ;
      RECT 82.42 3.96 82.47 4.405 ;
      RECT 82.41 3.992 82.42 4.403 ;
      RECT 82.405 4.017 82.41 4.403 ;
      RECT 82.385 4.09 82.405 4.403 ;
      RECT 82.375 4.17 82.385 4.402 ;
      RECT 82.36 4.2 82.375 4.402 ;
      RECT 82.345 4.205 82.36 4.401 ;
      RECT 82.285 4.207 82.34 4.398 ;
      RECT 82.255 4.212 82.285 4.394 ;
      RECT 82.253 4.215 82.255 4.393 ;
      RECT 82.167 4.217 82.253 4.39 ;
      RECT 82.081 4.223 82.167 4.384 ;
      RECT 81.995 4.228 82.081 4.378 ;
      RECT 81.922 4.233 81.995 4.379 ;
      RECT 81.836 4.239 81.922 4.387 ;
      RECT 81.75 4.245 81.836 4.396 ;
      RECT 81.73 4.249 81.75 4.401 ;
      RECT 81.683 4.251 81.73 4.404 ;
      RECT 81.597 4.256 81.683 4.41 ;
      RECT 81.511 4.261 81.597 4.419 ;
      RECT 81.425 4.267 81.511 4.427 ;
      RECT 81.34 4.265 81.425 4.436 ;
      RECT 81.336 4.26 81.34 4.44 ;
      RECT 81.25 4.255 81.336 4.432 ;
      RECT 81.186 4.246 81.25 4.42 ;
      RECT 81.1 4.237 81.186 4.407 ;
      RECT 81.076 4.23 81.1 4.398 ;
      RECT 80.99 4.224 81.076 4.385 ;
      RECT 80.95 4.217 80.99 4.371 ;
      RECT 80.945 4.207 80.95 4.367 ;
      RECT 80.935 4.195 80.945 4.366 ;
      RECT 80.915 4.165 80.935 4.363 ;
      RECT 80.86 4.085 80.915 4.357 ;
      RECT 80.84 4.004 80.86 4.352 ;
      RECT 80.82 3.962 80.84 4.348 ;
      RECT 80.795 3.915 80.82 4.342 ;
      RECT 80.79 3.89 80.795 4.339 ;
      RECT 80.755 3.87 80.79 4.334 ;
      RECT 80.746 3.87 80.755 4.327 ;
      RECT 80.66 3.87 80.746 4.297 ;
      RECT 80.655 3.87 80.66 4.26 ;
      RECT 80.62 3.87 80.64 4.182 ;
      RECT 80.615 3.912 80.62 4.147 ;
      RECT 80.61 3.987 80.615 4.103 ;
      RECT 82.06 3.792 82.235 4.04 ;
      RECT 82.06 3.792 82.24 4.038 ;
      RECT 82.055 3.824 82.24 3.998 ;
      RECT 82.085 3.765 82.255 3.985 ;
      RECT 82.05 3.842 82.255 3.918 ;
      RECT 81.36 3.305 81.53 3.48 ;
      RECT 81.36 3.305 81.702 3.472 ;
      RECT 81.36 3.305 81.785 3.466 ;
      RECT 81.36 3.305 81.82 3.462 ;
      RECT 81.36 3.305 81.84 3.461 ;
      RECT 81.36 3.305 81.926 3.457 ;
      RECT 81.82 3.13 81.99 3.452 ;
      RECT 81.395 3.237 82.02 3.45 ;
      RECT 81.385 3.292 82.025 3.448 ;
      RECT 81.36 3.328 82.035 3.443 ;
      RECT 81.36 3.355 82.04 3.373 ;
      RECT 81.425 3.18 82 3.45 ;
      RECT 81.616 3.165 82 3.45 ;
      RECT 81.45 3.168 82 3.45 ;
      RECT 81.53 3.166 81.616 3.477 ;
      RECT 81.616 3.163 81.995 3.45 ;
      RECT 81.8 3.14 81.995 3.45 ;
      RECT 81.702 3.161 81.995 3.45 ;
      RECT 81.785 3.155 81.8 3.463 ;
      RECT 81.935 4.52 81.94 4.72 ;
      RECT 81.4 4.585 81.445 4.72 ;
      RECT 81.97 4.52 81.99 4.693 ;
      RECT 81.94 4.52 81.97 4.708 ;
      RECT 81.875 4.52 81.935 4.745 ;
      RECT 81.86 4.52 81.875 4.775 ;
      RECT 81.845 4.52 81.86 4.788 ;
      RECT 81.825 4.52 81.845 4.803 ;
      RECT 81.82 4.52 81.825 4.812 ;
      RECT 81.81 4.524 81.82 4.817 ;
      RECT 81.795 4.534 81.81 4.828 ;
      RECT 81.77 4.55 81.795 4.838 ;
      RECT 81.76 4.564 81.77 4.84 ;
      RECT 81.74 4.576 81.76 4.837 ;
      RECT 81.71 4.597 81.74 4.831 ;
      RECT 81.7 4.609 81.71 4.826 ;
      RECT 81.69 4.607 81.7 4.823 ;
      RECT 81.675 4.606 81.69 4.818 ;
      RECT 81.67 4.605 81.675 4.813 ;
      RECT 81.635 4.603 81.67 4.803 ;
      RECT 81.615 4.6 81.635 4.785 ;
      RECT 81.605 4.598 81.615 4.78 ;
      RECT 81.595 4.597 81.605 4.775 ;
      RECT 81.56 4.595 81.595 4.763 ;
      RECT 81.505 4.591 81.56 4.743 ;
      RECT 81.495 4.589 81.505 4.728 ;
      RECT 81.49 4.589 81.495 4.723 ;
      RECT 81.445 4.587 81.49 4.72 ;
      RECT 81.35 4.585 81.4 4.724 ;
      RECT 81.34 4.586 81.35 4.729 ;
      RECT 81.28 4.593 81.34 4.743 ;
      RECT 81.255 4.601 81.28 4.763 ;
      RECT 81.245 4.605 81.255 4.775 ;
      RECT 81.24 4.606 81.245 4.78 ;
      RECT 81.225 4.608 81.24 4.783 ;
      RECT 81.21 4.61 81.225 4.788 ;
      RECT 81.205 4.61 81.21 4.791 ;
      RECT 81.16 4.615 81.205 4.802 ;
      RECT 81.155 4.619 81.16 4.814 ;
      RECT 81.13 4.615 81.155 4.818 ;
      RECT 81.12 4.611 81.13 4.822 ;
      RECT 81.11 4.61 81.12 4.826 ;
      RECT 81.095 4.6 81.11 4.832 ;
      RECT 81.09 4.588 81.095 4.836 ;
      RECT 81.085 4.585 81.09 4.837 ;
      RECT 81.08 4.582 81.085 4.839 ;
      RECT 81.065 4.57 81.08 4.838 ;
      RECT 81.05 4.552 81.065 4.835 ;
      RECT 81.03 4.531 81.05 4.828 ;
      RECT 80.965 4.52 81.03 4.8 ;
      RECT 80.961 4.52 80.965 4.779 ;
      RECT 80.875 4.52 80.961 4.749 ;
      RECT 80.86 4.52 80.875 4.705 ;
      RECT 81.51 4.871 81.525 5.13 ;
      RECT 81.51 4.886 81.53 5.129 ;
      RECT 81.426 4.886 81.53 5.127 ;
      RECT 81.426 4.9 81.535 5.126 ;
      RECT 81.34 4.942 81.54 5.123 ;
      RECT 81.335 4.885 81.525 5.118 ;
      RECT 81.335 4.956 81.545 5.115 ;
      RECT 81.33 4.987 81.545 5.113 ;
      RECT 81.335 4.984 81.56 5.103 ;
      RECT 81.33 5.03 81.575 5.088 ;
      RECT 81.33 5.058 81.58 5.073 ;
      RECT 81.34 4.86 81.51 5.123 ;
      RECT 81.1 3.87 81.27 4.04 ;
      RECT 81.065 3.87 81.27 4.035 ;
      RECT 81.055 3.87 81.27 4.028 ;
      RECT 81.05 3.855 81.22 4.025 ;
      RECT 79.88 4.392 80.145 4.835 ;
      RECT 79.875 4.363 80.09 4.833 ;
      RECT 79.87 4.517 80.15 4.828 ;
      RECT 79.875 4.412 80.15 4.828 ;
      RECT 79.875 4.423 80.16 4.815 ;
      RECT 79.875 4.37 80.12 4.833 ;
      RECT 79.88 4.357 80.09 4.835 ;
      RECT 79.88 4.355 80.04 4.835 ;
      RECT 79.981 4.347 80.04 4.835 ;
      RECT 79.895 4.348 80.04 4.835 ;
      RECT 79.981 4.346 80.03 4.835 ;
      RECT 79.785 3.161 79.96 3.46 ;
      RECT 79.835 3.123 79.96 3.46 ;
      RECT 79.82 3.125 80.046 3.452 ;
      RECT 79.82 3.128 80.085 3.439 ;
      RECT 79.82 3.129 80.095 3.425 ;
      RECT 79.775 3.18 80.095 3.415 ;
      RECT 79.82 3.13 80.1 3.41 ;
      RECT 79.775 3.34 80.105 3.4 ;
      RECT 79.76 3.2 80.1 3.34 ;
      RECT 79.755 3.216 80.1 3.28 ;
      RECT 79.8 3.14 80.1 3.41 ;
      RECT 79.835 3.121 79.921 3.46 ;
      RECT 78.295 7.31 78.465 8.78 ;
      RECT 78.295 7.31 78.47 8.57 ;
      RECT 77.925 9.26 78.395 9.43 ;
      RECT 77.925 8.24 78.095 9.43 ;
      RECT 77.92 3.035 78.09 4.225 ;
      RECT 77.92 3.035 78.39 3.205 ;
      RECT 77.305 3.895 77.48 5.155 ;
      RECT 77.305 3.685 77.475 5.155 ;
      RECT 77.305 7.31 77.475 8.78 ;
      RECT 77.305 7.31 77.48 8.57 ;
      RECT 76.935 3.035 77.105 4.225 ;
      RECT 76.935 3.035 77.405 3.205 ;
      RECT 76.935 9.26 77.405 9.43 ;
      RECT 76.935 8.24 77.105 9.43 ;
      RECT 75.945 4.015 76.12 5.155 ;
      RECT 75.945 1.865 76.115 5.155 ;
      RECT 75.945 1.865 76.12 2.415 ;
      RECT 75.945 10.05 76.12 10.6 ;
      RECT 75.945 7.31 76.115 10.6 ;
      RECT 75.945 7.31 76.12 8.45 ;
      RECT 75.515 3.895 75.69 5.155 ;
      RECT 75.515 2.945 75.685 5.155 ;
      RECT 75.515 7.31 75.685 9.52 ;
      RECT 75.515 7.31 75.69 8.57 ;
      RECT 75.085 3.925 75.255 5.155 ;
      RECT 75.145 2.145 75.315 4.095 ;
      RECT 75.085 1.865 75.255 2.315 ;
      RECT 75.085 10.15 75.255 10.6 ;
      RECT 75.145 8.37 75.315 10.32 ;
      RECT 75.085 7.31 75.255 8.54 ;
      RECT 74.56 3.895 74.735 5.155 ;
      RECT 74.56 1.865 74.73 5.155 ;
      RECT 74.56 3.365 74.97 3.695 ;
      RECT 74.56 2.525 74.97 2.855 ;
      RECT 74.56 1.865 74.735 2.355 ;
      RECT 74.56 10.11 74.735 10.6 ;
      RECT 74.56 7.31 74.73 10.6 ;
      RECT 74.56 9.61 74.97 9.94 ;
      RECT 74.56 8.77 74.97 9.1 ;
      RECT 74.56 7.31 74.735 8.57 ;
      RECT 72.49 4.421 72.495 4.593 ;
      RECT 72.485 4.414 72.49 4.683 ;
      RECT 72.48 4.408 72.485 4.702 ;
      RECT 72.46 4.402 72.48 4.712 ;
      RECT 72.445 4.397 72.46 4.72 ;
      RECT 72.408 4.391 72.445 4.718 ;
      RECT 72.322 4.377 72.408 4.714 ;
      RECT 72.236 4.359 72.322 4.709 ;
      RECT 72.15 4.34 72.236 4.703 ;
      RECT 72.12 4.328 72.15 4.699 ;
      RECT 72.1 4.322 72.12 4.698 ;
      RECT 72.035 4.32 72.1 4.696 ;
      RECT 72.02 4.32 72.035 4.688 ;
      RECT 72.005 4.32 72.02 4.675 ;
      RECT 72 4.32 72.005 4.665 ;
      RECT 71.985 4.32 72 4.643 ;
      RECT 71.97 4.32 71.985 4.61 ;
      RECT 71.965 4.32 71.97 4.588 ;
      RECT 71.955 4.32 71.965 4.57 ;
      RECT 71.94 4.32 71.955 4.548 ;
      RECT 71.92 4.32 71.94 4.51 ;
      RECT 72.27 3.605 72.305 4.044 ;
      RECT 72.27 3.605 72.31 4.043 ;
      RECT 72.215 3.665 72.31 4.042 ;
      RECT 72.08 3.837 72.31 4.041 ;
      RECT 72.19 3.715 72.31 4.041 ;
      RECT 72.08 3.837 72.335 4.031 ;
      RECT 72.135 3.782 72.415 3.948 ;
      RECT 72.31 3.576 72.315 4.039 ;
      RECT 72.165 3.752 72.455 3.825 ;
      RECT 72.18 3.735 72.31 4.041 ;
      RECT 72.315 3.575 72.485 3.763 ;
      RECT 72.305 3.578 72.485 3.763 ;
      RECT 71.81 3.455 71.98 3.765 ;
      RECT 71.81 3.455 71.985 3.738 ;
      RECT 71.81 3.455 71.99 3.715 ;
      RECT 71.81 3.455 72 3.665 ;
      RECT 71.805 3.56 72 3.635 ;
      RECT 71.84 3.13 72.01 3.608 ;
      RECT 71.84 3.13 72.025 3.529 ;
      RECT 71.83 3.34 72.025 3.529 ;
      RECT 71.84 3.14 72.035 3.444 ;
      RECT 71.77 3.882 71.775 4.085 ;
      RECT 71.76 3.87 71.77 4.195 ;
      RECT 71.735 3.87 71.76 4.235 ;
      RECT 71.655 3.87 71.735 4.32 ;
      RECT 71.645 3.87 71.655 4.39 ;
      RECT 71.62 3.87 71.645 4.413 ;
      RECT 71.6 3.87 71.62 4.448 ;
      RECT 71.555 3.88 71.6 4.491 ;
      RECT 71.545 3.892 71.555 4.528 ;
      RECT 71.525 3.906 71.545 4.548 ;
      RECT 71.515 3.924 71.525 4.564 ;
      RECT 71.5 3.95 71.515 4.574 ;
      RECT 71.485 3.991 71.5 4.588 ;
      RECT 71.475 4.026 71.485 4.598 ;
      RECT 71.47 4.042 71.475 4.603 ;
      RECT 71.46 4.057 71.47 4.608 ;
      RECT 71.44 4.1 71.46 4.618 ;
      RECT 71.42 4.137 71.44 4.631 ;
      RECT 71.385 4.16 71.42 4.649 ;
      RECT 71.375 4.174 71.385 4.665 ;
      RECT 71.355 4.184 71.375 4.675 ;
      RECT 71.35 4.193 71.355 4.683 ;
      RECT 71.34 4.2 71.35 4.69 ;
      RECT 71.33 4.207 71.34 4.698 ;
      RECT 71.315 4.217 71.33 4.706 ;
      RECT 71.305 4.231 71.315 4.716 ;
      RECT 71.295 4.243 71.305 4.728 ;
      RECT 71.28 4.265 71.295 4.741 ;
      RECT 71.27 4.287 71.28 4.752 ;
      RECT 71.26 4.307 71.27 4.761 ;
      RECT 71.255 4.322 71.26 4.768 ;
      RECT 71.225 4.355 71.255 4.782 ;
      RECT 71.215 4.39 71.225 4.797 ;
      RECT 71.21 4.397 71.215 4.803 ;
      RECT 71.19 4.412 71.21 4.81 ;
      RECT 71.185 4.427 71.19 4.818 ;
      RECT 71.18 4.436 71.185 4.823 ;
      RECT 71.165 4.442 71.18 4.83 ;
      RECT 71.16 4.448 71.165 4.838 ;
      RECT 71.155 4.452 71.16 4.845 ;
      RECT 71.15 4.456 71.155 4.855 ;
      RECT 71.14 4.461 71.15 4.865 ;
      RECT 71.12 4.472 71.14 4.893 ;
      RECT 71.105 4.484 71.12 4.92 ;
      RECT 71.085 4.497 71.105 4.945 ;
      RECT 71.065 4.512 71.085 4.969 ;
      RECT 71.05 4.527 71.065 4.984 ;
      RECT 71.045 4.538 71.05 4.993 ;
      RECT 70.98 4.583 71.045 5.003 ;
      RECT 70.945 4.642 70.98 5.016 ;
      RECT 70.94 4.665 70.945 5.022 ;
      RECT 70.935 4.672 70.94 5.024 ;
      RECT 70.92 4.682 70.935 5.027 ;
      RECT 70.89 4.707 70.92 5.031 ;
      RECT 70.885 4.725 70.89 5.035 ;
      RECT 70.88 4.732 70.885 5.036 ;
      RECT 70.86 4.74 70.88 5.04 ;
      RECT 70.85 4.747 70.86 5.044 ;
      RECT 70.806 4.758 70.85 5.051 ;
      RECT 70.72 4.786 70.806 5.067 ;
      RECT 70.66 4.81 70.72 5.085 ;
      RECT 70.615 4.82 70.66 5.099 ;
      RECT 70.556 4.828 70.615 5.113 ;
      RECT 70.47 4.835 70.556 5.132 ;
      RECT 70.445 4.84 70.47 5.147 ;
      RECT 70.365 4.843 70.445 5.15 ;
      RECT 70.285 4.847 70.365 5.137 ;
      RECT 70.276 4.85 70.285 5.122 ;
      RECT 70.19 4.85 70.276 5.107 ;
      RECT 70.13 4.852 70.19 5.084 ;
      RECT 70.126 4.855 70.13 5.074 ;
      RECT 70.04 4.855 70.126 5.059 ;
      RECT 69.965 4.855 70.04 5.035 ;
      RECT 71.28 3.864 71.29 4.04 ;
      RECT 71.235 3.831 71.28 4.04 ;
      RECT 71.19 3.782 71.235 4.04 ;
      RECT 71.16 3.752 71.19 4.041 ;
      RECT 71.155 3.735 71.16 4.042 ;
      RECT 71.13 3.715 71.155 4.043 ;
      RECT 71.115 3.69 71.13 4.044 ;
      RECT 71.11 3.677 71.115 4.045 ;
      RECT 71.105 3.671 71.11 4.043 ;
      RECT 71.1 3.663 71.105 4.037 ;
      RECT 71.075 3.655 71.1 4.017 ;
      RECT 71.055 3.644 71.075 3.988 ;
      RECT 71.025 3.629 71.055 3.959 ;
      RECT 71.005 3.615 71.025 3.931 ;
      RECT 70.995 3.609 71.005 3.91 ;
      RECT 70.99 3.606 70.995 3.893 ;
      RECT 70.985 3.603 70.99 3.878 ;
      RECT 70.97 3.598 70.985 3.843 ;
      RECT 70.965 3.594 70.97 3.81 ;
      RECT 70.945 3.589 70.965 3.786 ;
      RECT 70.915 3.581 70.945 3.751 ;
      RECT 70.9 3.575 70.915 3.728 ;
      RECT 70.86 3.568 70.9 3.713 ;
      RECT 70.835 3.56 70.86 3.693 ;
      RECT 70.815 3.555 70.835 3.683 ;
      RECT 70.78 3.549 70.815 3.678 ;
      RECT 70.735 3.54 70.78 3.677 ;
      RECT 70.705 3.536 70.735 3.679 ;
      RECT 70.62 3.544 70.705 3.683 ;
      RECT 70.55 3.555 70.62 3.705 ;
      RECT 70.537 3.561 70.55 3.728 ;
      RECT 70.451 3.568 70.537 3.75 ;
      RECT 70.365 3.58 70.451 3.787 ;
      RECT 70.365 3.957 70.375 4.195 ;
      RECT 70.36 3.586 70.365 3.81 ;
      RECT 70.355 3.842 70.365 4.195 ;
      RECT 70.355 3.587 70.36 3.815 ;
      RECT 70.35 3.588 70.355 4.195 ;
      RECT 70.326 3.59 70.35 4.196 ;
      RECT 70.24 3.598 70.326 4.198 ;
      RECT 70.22 3.612 70.24 4.201 ;
      RECT 70.215 3.64 70.22 4.202 ;
      RECT 70.21 3.652 70.215 4.203 ;
      RECT 70.205 3.667 70.21 4.204 ;
      RECT 70.195 3.697 70.205 4.205 ;
      RECT 70.19 3.735 70.195 4.203 ;
      RECT 70.185 3.755 70.19 4.198 ;
      RECT 70.17 3.79 70.185 4.183 ;
      RECT 70.16 3.842 70.17 4.163 ;
      RECT 70.155 3.872 70.16 4.151 ;
      RECT 70.14 3.885 70.155 4.134 ;
      RECT 70.115 3.889 70.14 4.101 ;
      RECT 70.1 3.887 70.115 4.078 ;
      RECT 70.085 3.886 70.1 4.075 ;
      RECT 70.025 3.884 70.085 4.073 ;
      RECT 70.015 3.882 70.025 4.068 ;
      RECT 69.975 3.881 70.015 4.065 ;
      RECT 69.905 3.878 69.975 4.063 ;
      RECT 69.85 3.876 69.905 4.058 ;
      RECT 69.78 3.87 69.85 4.053 ;
      RECT 69.771 3.87 69.78 4.05 ;
      RECT 69.685 3.87 69.771 4.045 ;
      RECT 69.68 3.87 69.685 4.04 ;
      RECT 70.985 3.105 71.16 3.455 ;
      RECT 70.985 3.12 71.17 3.453 ;
      RECT 70.96 3.07 71.105 3.45 ;
      RECT 70.94 3.071 71.105 3.443 ;
      RECT 70.93 3.072 71.115 3.438 ;
      RECT 70.9 3.073 71.115 3.425 ;
      RECT 70.85 3.074 71.115 3.401 ;
      RECT 70.845 3.076 71.115 3.386 ;
      RECT 70.845 3.142 71.175 3.38 ;
      RECT 70.825 3.083 71.13 3.36 ;
      RECT 70.815 3.092 71.14 3.215 ;
      RECT 70.825 3.087 71.14 3.36 ;
      RECT 70.845 3.077 71.13 3.386 ;
      RECT 70.43 4.402 70.6 4.69 ;
      RECT 70.425 4.42 70.61 4.685 ;
      RECT 70.39 4.428 70.675 4.605 ;
      RECT 70.39 4.428 70.761 4.595 ;
      RECT 70.39 4.428 70.815 4.541 ;
      RECT 70.675 4.325 70.845 4.509 ;
      RECT 70.39 4.48 70.85 4.497 ;
      RECT 70.375 4.45 70.845 4.493 ;
      RECT 70.635 4.332 70.675 4.644 ;
      RECT 70.515 4.369 70.845 4.509 ;
      RECT 70.61 4.344 70.635 4.67 ;
      RECT 70.6 4.351 70.845 4.509 ;
      RECT 70.731 3.815 70.8 4.074 ;
      RECT 70.731 3.87 70.805 4.073 ;
      RECT 70.645 3.87 70.805 4.072 ;
      RECT 70.64 3.87 70.81 4.065 ;
      RECT 70.63 3.815 70.8 4.06 ;
      RECT 70.31 10.05 70.485 10.6 ;
      RECT 70.31 7.31 70.48 10.6 ;
      RECT 70.31 7.31 70.485 8.45 ;
      RECT 70.01 3.114 70.185 3.415 ;
      RECT 69.995 3.102 70.01 3.4 ;
      RECT 69.965 3.101 69.995 3.353 ;
      RECT 69.965 3.119 70.19 3.348 ;
      RECT 69.95 3.103 70.01 3.313 ;
      RECT 69.945 3.125 70.2 3.213 ;
      RECT 69.945 3.108 70.096 3.213 ;
      RECT 69.945 3.11 70.1 3.213 ;
      RECT 69.95 3.106 70.096 3.313 ;
      RECT 70.055 4.342 70.06 4.69 ;
      RECT 70.045 4.332 70.055 4.696 ;
      RECT 70.01 4.322 70.045 4.698 ;
      RECT 69.972 4.317 70.01 4.702 ;
      RECT 69.886 4.31 69.972 4.709 ;
      RECT 69.8 4.3 69.886 4.719 ;
      RECT 69.755 4.295 69.8 4.727 ;
      RECT 69.751 4.295 69.755 4.731 ;
      RECT 69.665 4.295 69.751 4.738 ;
      RECT 69.65 4.295 69.665 4.738 ;
      RECT 69.64 4.293 69.65 4.71 ;
      RECT 69.63 4.289 69.64 4.653 ;
      RECT 69.61 4.283 69.63 4.585 ;
      RECT 69.605 4.279 69.61 4.533 ;
      RECT 69.595 4.278 69.605 4.5 ;
      RECT 69.545 4.276 69.595 4.485 ;
      RECT 69.52 4.274 69.545 4.48 ;
      RECT 69.477 4.272 69.52 4.476 ;
      RECT 69.391 4.268 69.477 4.464 ;
      RECT 69.305 4.263 69.391 4.448 ;
      RECT 69.275 4.26 69.305 4.435 ;
      RECT 69.25 4.259 69.275 4.423 ;
      RECT 69.245 4.259 69.25 4.413 ;
      RECT 69.205 4.258 69.245 4.405 ;
      RECT 69.19 4.257 69.205 4.398 ;
      RECT 69.14 4.256 69.19 4.39 ;
      RECT 69.138 4.255 69.14 4.385 ;
      RECT 69.052 4.253 69.138 4.385 ;
      RECT 68.966 4.248 69.052 4.385 ;
      RECT 68.88 4.244 68.966 4.385 ;
      RECT 68.831 4.24 68.88 4.383 ;
      RECT 68.745 4.237 68.831 4.378 ;
      RECT 68.722 4.234 68.745 4.374 ;
      RECT 68.636 4.231 68.722 4.369 ;
      RECT 68.55 4.227 68.636 4.36 ;
      RECT 68.525 4.22 68.55 4.355 ;
      RECT 68.465 4.185 68.525 4.352 ;
      RECT 68.445 4.11 68.465 4.349 ;
      RECT 68.44 4.052 68.445 4.348 ;
      RECT 68.415 3.992 68.44 4.347 ;
      RECT 68.34 3.87 68.415 4.343 ;
      RECT 68.33 3.87 68.34 4.335 ;
      RECT 68.315 3.87 68.33 4.325 ;
      RECT 68.3 3.87 68.315 4.295 ;
      RECT 68.285 3.87 68.3 4.24 ;
      RECT 68.27 3.87 68.285 4.178 ;
      RECT 68.245 3.87 68.27 4.103 ;
      RECT 68.24 3.87 68.245 4.053 ;
      RECT 69.88 7.31 70.05 9.52 ;
      RECT 69.88 7.31 70.055 8.57 ;
      RECT 69.585 3.415 69.605 3.724 ;
      RECT 69.571 3.417 69.62 3.721 ;
      RECT 69.571 3.422 69.64 3.712 ;
      RECT 69.485 3.42 69.62 3.706 ;
      RECT 69.485 3.428 69.675 3.689 ;
      RECT 69.45 3.43 69.675 3.688 ;
      RECT 69.42 3.438 69.675 3.679 ;
      RECT 69.41 3.443 69.695 3.665 ;
      RECT 69.45 3.433 69.695 3.665 ;
      RECT 69.45 3.436 69.705 3.653 ;
      RECT 69.42 3.438 69.715 3.64 ;
      RECT 69.42 3.442 69.725 3.583 ;
      RECT 69.41 3.447 69.73 3.498 ;
      RECT 69.571 3.415 69.605 3.721 ;
      RECT 69.01 3.518 69.015 3.73 ;
      RECT 68.885 3.515 68.9 3.73 ;
      RECT 68.35 3.545 68.42 3.73 ;
      RECT 68.235 3.545 68.27 3.725 ;
      RECT 69.356 3.847 69.375 4.041 ;
      RECT 69.27 3.802 69.356 4.042 ;
      RECT 69.26 3.755 69.27 4.044 ;
      RECT 69.255 3.735 69.26 4.045 ;
      RECT 69.235 3.7 69.255 4.046 ;
      RECT 69.22 3.65 69.235 4.047 ;
      RECT 69.2 3.587 69.22 4.048 ;
      RECT 69.19 3.55 69.2 4.049 ;
      RECT 69.175 3.539 69.19 4.05 ;
      RECT 69.17 3.531 69.175 4.048 ;
      RECT 69.16 3.53 69.17 4.04 ;
      RECT 69.13 3.527 69.16 4.019 ;
      RECT 69.055 3.522 69.13 3.964 ;
      RECT 69.04 3.518 69.055 3.91 ;
      RECT 69.03 3.518 69.04 3.805 ;
      RECT 69.015 3.518 69.03 3.738 ;
      RECT 69 3.518 69.01 3.728 ;
      RECT 68.945 3.517 69 3.725 ;
      RECT 68.9 3.515 68.945 3.728 ;
      RECT 68.872 3.515 68.885 3.731 ;
      RECT 68.786 3.519 68.872 3.733 ;
      RECT 68.7 3.525 68.786 3.738 ;
      RECT 68.68 3.529 68.7 3.74 ;
      RECT 68.678 3.53 68.68 3.739 ;
      RECT 68.592 3.532 68.678 3.738 ;
      RECT 68.506 3.537 68.592 3.735 ;
      RECT 68.42 3.542 68.506 3.732 ;
      RECT 68.27 3.545 68.35 3.728 ;
      RECT 68.925 10.11 69.1 10.6 ;
      RECT 68.925 7.31 69.095 10.6 ;
      RECT 68.925 9.61 69.335 9.94 ;
      RECT 68.925 8.77 69.335 9.1 ;
      RECT 68.925 7.31 69.1 8.57 ;
      RECT 69.046 4.52 69.095 4.854 ;
      RECT 69.046 4.52 69.1 4.853 ;
      RECT 68.96 4.52 69.1 4.852 ;
      RECT 68.735 4.628 69.105 4.85 ;
      RECT 68.96 4.52 69.13 4.843 ;
      RECT 68.93 4.532 69.135 4.834 ;
      RECT 68.915 4.55 69.14 4.831 ;
      RECT 68.73 4.634 69.14 4.758 ;
      RECT 68.725 4.641 69.14 4.718 ;
      RECT 68.74 4.607 69.14 4.831 ;
      RECT 68.901 4.553 69.105 4.85 ;
      RECT 68.815 4.573 69.14 4.831 ;
      RECT 68.915 4.547 69.135 4.834 ;
      RECT 68.685 3.871 68.875 4.065 ;
      RECT 68.68 3.873 68.875 4.064 ;
      RECT 68.675 3.877 68.89 4.061 ;
      RECT 68.69 3.87 68.89 4.061 ;
      RECT 68.675 3.98 68.895 4.056 ;
      RECT 67.97 4.48 68.061 4.778 ;
      RECT 67.965 4.482 68.14 4.773 ;
      RECT 67.97 4.48 68.14 4.773 ;
      RECT 67.965 4.486 68.16 4.771 ;
      RECT 67.965 4.541 68.2 4.77 ;
      RECT 67.965 4.576 68.215 4.764 ;
      RECT 67.965 4.61 68.225 4.754 ;
      RECT 67.955 4.49 68.16 4.605 ;
      RECT 67.955 4.51 68.175 4.605 ;
      RECT 67.955 4.493 68.165 4.605 ;
      RECT 68.18 3.261 68.185 3.323 ;
      RECT 68.175 3.183 68.18 3.346 ;
      RECT 68.17 3.14 68.175 3.357 ;
      RECT 68.165 3.13 68.17 3.369 ;
      RECT 68.16 3.13 68.165 3.378 ;
      RECT 68.135 3.13 68.16 3.41 ;
      RECT 68.13 3.13 68.135 3.443 ;
      RECT 68.115 3.13 68.13 3.468 ;
      RECT 68.105 3.13 68.115 3.495 ;
      RECT 68.1 3.13 68.105 3.508 ;
      RECT 68.095 3.13 68.1 3.523 ;
      RECT 68.085 3.13 68.095 3.538 ;
      RECT 68.08 3.13 68.085 3.558 ;
      RECT 68.055 3.13 68.08 3.593 ;
      RECT 68.01 3.13 68.055 3.638 ;
      RECT 68 3.13 68.01 3.651 ;
      RECT 67.915 3.215 68 3.658 ;
      RECT 67.88 3.337 67.915 3.667 ;
      RECT 67.875 3.377 67.88 3.671 ;
      RECT 67.855 3.4 67.875 3.673 ;
      RECT 67.85 3.43 67.855 3.676 ;
      RECT 67.84 3.442 67.85 3.677 ;
      RECT 67.795 3.465 67.84 3.682 ;
      RECT 67.755 3.495 67.795 3.69 ;
      RECT 67.72 3.507 67.755 3.696 ;
      RECT 67.715 3.512 67.72 3.7 ;
      RECT 67.645 3.522 67.715 3.707 ;
      RECT 67.605 3.532 67.645 3.717 ;
      RECT 67.585 3.537 67.605 3.723 ;
      RECT 67.575 3.541 67.585 3.728 ;
      RECT 67.57 3.544 67.575 3.731 ;
      RECT 67.56 3.545 67.57 3.732 ;
      RECT 67.535 3.547 67.56 3.736 ;
      RECT 67.525 3.552 67.535 3.739 ;
      RECT 67.48 3.56 67.525 3.74 ;
      RECT 67.355 3.565 67.48 3.74 ;
      RECT 67.91 3.862 67.93 4.044 ;
      RECT 67.861 3.847 67.91 4.043 ;
      RECT 67.775 3.862 67.93 4.041 ;
      RECT 67.76 3.862 67.93 4.04 ;
      RECT 67.725 3.84 67.895 4.025 ;
      RECT 67.795 4.86 67.81 5.069 ;
      RECT 67.795 4.868 67.815 5.068 ;
      RECT 67.74 4.868 67.815 5.067 ;
      RECT 67.72 4.872 67.82 5.065 ;
      RECT 67.7 4.822 67.74 5.064 ;
      RECT 67.645 4.88 67.825 5.062 ;
      RECT 67.61 4.837 67.74 5.06 ;
      RECT 67.606 4.84 67.795 5.059 ;
      RECT 67.52 4.848 67.795 5.057 ;
      RECT 67.52 4.892 67.83 5.05 ;
      RECT 67.51 4.985 67.83 5.048 ;
      RECT 67.52 4.904 67.835 5.033 ;
      RECT 67.52 4.925 67.85 5.003 ;
      RECT 67.52 4.952 67.855 4.973 ;
      RECT 67.645 4.83 67.74 5.062 ;
      RECT 67.275 3.875 67.28 4.413 ;
      RECT 67.08 4.205 67.085 4.4 ;
      RECT 65.38 3.87 65.395 4.25 ;
      RECT 67.445 3.87 67.45 4.04 ;
      RECT 67.44 3.87 67.445 4.05 ;
      RECT 67.435 3.87 67.44 4.063 ;
      RECT 67.41 3.87 67.435 4.105 ;
      RECT 67.385 3.87 67.41 4.178 ;
      RECT 67.37 3.87 67.385 4.23 ;
      RECT 67.365 3.87 67.37 4.26 ;
      RECT 67.34 3.87 67.365 4.3 ;
      RECT 67.325 3.87 67.34 4.355 ;
      RECT 67.32 3.87 67.325 4.388 ;
      RECT 67.295 3.87 67.32 4.408 ;
      RECT 67.28 3.87 67.295 4.414 ;
      RECT 67.21 3.905 67.275 4.41 ;
      RECT 67.16 3.96 67.21 4.405 ;
      RECT 67.15 3.992 67.16 4.403 ;
      RECT 67.145 4.017 67.15 4.403 ;
      RECT 67.125 4.09 67.145 4.403 ;
      RECT 67.115 4.17 67.125 4.402 ;
      RECT 67.1 4.2 67.115 4.402 ;
      RECT 67.085 4.205 67.1 4.401 ;
      RECT 67.025 4.207 67.08 4.398 ;
      RECT 66.995 4.212 67.025 4.394 ;
      RECT 66.993 4.215 66.995 4.393 ;
      RECT 66.907 4.217 66.993 4.39 ;
      RECT 66.821 4.223 66.907 4.384 ;
      RECT 66.735 4.228 66.821 4.378 ;
      RECT 66.662 4.233 66.735 4.379 ;
      RECT 66.576 4.239 66.662 4.387 ;
      RECT 66.49 4.245 66.576 4.396 ;
      RECT 66.47 4.249 66.49 4.401 ;
      RECT 66.423 4.251 66.47 4.404 ;
      RECT 66.337 4.256 66.423 4.41 ;
      RECT 66.251 4.261 66.337 4.419 ;
      RECT 66.165 4.267 66.251 4.427 ;
      RECT 66.08 4.265 66.165 4.436 ;
      RECT 66.076 4.26 66.08 4.44 ;
      RECT 65.99 4.255 66.076 4.432 ;
      RECT 65.926 4.246 65.99 4.42 ;
      RECT 65.84 4.237 65.926 4.407 ;
      RECT 65.816 4.23 65.84 4.398 ;
      RECT 65.73 4.224 65.816 4.385 ;
      RECT 65.69 4.217 65.73 4.371 ;
      RECT 65.685 4.207 65.69 4.367 ;
      RECT 65.675 4.195 65.685 4.366 ;
      RECT 65.655 4.165 65.675 4.363 ;
      RECT 65.6 4.085 65.655 4.357 ;
      RECT 65.58 4.004 65.6 4.352 ;
      RECT 65.56 3.962 65.58 4.348 ;
      RECT 65.535 3.915 65.56 4.342 ;
      RECT 65.53 3.89 65.535 4.339 ;
      RECT 65.495 3.87 65.53 4.334 ;
      RECT 65.486 3.87 65.495 4.327 ;
      RECT 65.4 3.87 65.486 4.297 ;
      RECT 65.395 3.87 65.4 4.26 ;
      RECT 65.36 3.87 65.38 4.182 ;
      RECT 65.355 3.912 65.36 4.147 ;
      RECT 65.35 3.987 65.355 4.103 ;
      RECT 66.8 3.792 66.975 4.04 ;
      RECT 66.8 3.792 66.98 4.038 ;
      RECT 66.795 3.824 66.98 3.998 ;
      RECT 66.825 3.765 66.995 3.985 ;
      RECT 66.79 3.842 66.995 3.918 ;
      RECT 66.1 3.305 66.27 3.48 ;
      RECT 66.1 3.305 66.442 3.472 ;
      RECT 66.1 3.305 66.525 3.466 ;
      RECT 66.1 3.305 66.56 3.462 ;
      RECT 66.1 3.305 66.58 3.461 ;
      RECT 66.1 3.305 66.666 3.457 ;
      RECT 66.56 3.13 66.73 3.452 ;
      RECT 66.135 3.237 66.76 3.45 ;
      RECT 66.125 3.292 66.765 3.448 ;
      RECT 66.1 3.328 66.775 3.443 ;
      RECT 66.1 3.355 66.78 3.373 ;
      RECT 66.165 3.18 66.74 3.45 ;
      RECT 66.356 3.165 66.74 3.45 ;
      RECT 66.19 3.168 66.74 3.45 ;
      RECT 66.27 3.166 66.356 3.477 ;
      RECT 66.356 3.163 66.735 3.45 ;
      RECT 66.54 3.14 66.735 3.45 ;
      RECT 66.442 3.161 66.735 3.45 ;
      RECT 66.525 3.155 66.54 3.463 ;
      RECT 66.675 4.52 66.68 4.72 ;
      RECT 66.14 4.585 66.185 4.72 ;
      RECT 66.71 4.52 66.73 4.693 ;
      RECT 66.68 4.52 66.71 4.708 ;
      RECT 66.615 4.52 66.675 4.745 ;
      RECT 66.6 4.52 66.615 4.775 ;
      RECT 66.585 4.52 66.6 4.788 ;
      RECT 66.565 4.52 66.585 4.803 ;
      RECT 66.56 4.52 66.565 4.812 ;
      RECT 66.55 4.524 66.56 4.817 ;
      RECT 66.535 4.534 66.55 4.828 ;
      RECT 66.51 4.55 66.535 4.838 ;
      RECT 66.5 4.564 66.51 4.84 ;
      RECT 66.48 4.576 66.5 4.837 ;
      RECT 66.45 4.597 66.48 4.831 ;
      RECT 66.44 4.609 66.45 4.826 ;
      RECT 66.43 4.607 66.44 4.823 ;
      RECT 66.415 4.606 66.43 4.818 ;
      RECT 66.41 4.605 66.415 4.813 ;
      RECT 66.375 4.603 66.41 4.803 ;
      RECT 66.355 4.6 66.375 4.785 ;
      RECT 66.345 4.598 66.355 4.78 ;
      RECT 66.335 4.597 66.345 4.775 ;
      RECT 66.3 4.595 66.335 4.763 ;
      RECT 66.245 4.591 66.3 4.743 ;
      RECT 66.235 4.589 66.245 4.728 ;
      RECT 66.23 4.589 66.235 4.723 ;
      RECT 66.185 4.587 66.23 4.72 ;
      RECT 66.09 4.585 66.14 4.724 ;
      RECT 66.08 4.586 66.09 4.729 ;
      RECT 66.02 4.593 66.08 4.743 ;
      RECT 65.995 4.601 66.02 4.763 ;
      RECT 65.985 4.605 65.995 4.775 ;
      RECT 65.98 4.606 65.985 4.78 ;
      RECT 65.965 4.608 65.98 4.783 ;
      RECT 65.95 4.61 65.965 4.788 ;
      RECT 65.945 4.61 65.95 4.791 ;
      RECT 65.9 4.615 65.945 4.802 ;
      RECT 65.895 4.619 65.9 4.814 ;
      RECT 65.87 4.615 65.895 4.818 ;
      RECT 65.86 4.611 65.87 4.822 ;
      RECT 65.85 4.61 65.86 4.826 ;
      RECT 65.835 4.6 65.85 4.832 ;
      RECT 65.83 4.588 65.835 4.836 ;
      RECT 65.825 4.585 65.83 4.837 ;
      RECT 65.82 4.582 65.825 4.839 ;
      RECT 65.805 4.57 65.82 4.838 ;
      RECT 65.79 4.552 65.805 4.835 ;
      RECT 65.77 4.531 65.79 4.828 ;
      RECT 65.705 4.52 65.77 4.8 ;
      RECT 65.701 4.52 65.705 4.779 ;
      RECT 65.615 4.52 65.701 4.749 ;
      RECT 65.6 4.52 65.615 4.705 ;
      RECT 66.25 4.871 66.265 5.13 ;
      RECT 66.25 4.886 66.27 5.129 ;
      RECT 66.166 4.886 66.27 5.127 ;
      RECT 66.166 4.9 66.275 5.126 ;
      RECT 66.08 4.942 66.28 5.123 ;
      RECT 66.075 4.885 66.265 5.118 ;
      RECT 66.075 4.956 66.285 5.115 ;
      RECT 66.07 4.987 66.285 5.113 ;
      RECT 66.075 4.984 66.3 5.103 ;
      RECT 66.07 5.03 66.315 5.088 ;
      RECT 66.07 5.058 66.32 5.073 ;
      RECT 66.08 4.86 66.25 5.123 ;
      RECT 65.84 3.87 66.01 4.04 ;
      RECT 65.805 3.87 66.01 4.035 ;
      RECT 65.795 3.87 66.01 4.028 ;
      RECT 65.79 3.855 65.96 4.025 ;
      RECT 64.62 4.392 64.885 4.835 ;
      RECT 64.615 4.363 64.83 4.833 ;
      RECT 64.61 4.517 64.89 4.828 ;
      RECT 64.615 4.412 64.89 4.828 ;
      RECT 64.615 4.423 64.9 4.815 ;
      RECT 64.615 4.37 64.86 4.833 ;
      RECT 64.62 4.357 64.83 4.835 ;
      RECT 64.62 4.355 64.78 4.835 ;
      RECT 64.721 4.347 64.78 4.835 ;
      RECT 64.635 4.348 64.78 4.835 ;
      RECT 64.721 4.346 64.77 4.835 ;
      RECT 64.525 3.161 64.7 3.46 ;
      RECT 64.575 3.123 64.7 3.46 ;
      RECT 64.56 3.125 64.786 3.452 ;
      RECT 64.56 3.128 64.825 3.439 ;
      RECT 64.56 3.129 64.835 3.425 ;
      RECT 64.515 3.18 64.835 3.415 ;
      RECT 64.56 3.13 64.84 3.41 ;
      RECT 64.515 3.34 64.845 3.4 ;
      RECT 64.5 3.2 64.84 3.34 ;
      RECT 64.495 3.216 64.84 3.28 ;
      RECT 64.54 3.14 64.84 3.41 ;
      RECT 64.575 3.121 64.661 3.46 ;
      RECT 63.035 7.31 63.205 8.78 ;
      RECT 63.035 7.31 63.21 8.57 ;
      RECT 62.665 9.26 63.135 9.43 ;
      RECT 62.665 8.24 62.835 9.43 ;
      RECT 62.66 3.035 62.83 4.225 ;
      RECT 62.66 3.035 63.13 3.205 ;
      RECT 62.045 3.895 62.22 5.155 ;
      RECT 62.045 3.685 62.215 5.155 ;
      RECT 62.045 7.31 62.215 8.78 ;
      RECT 62.045 7.31 62.22 8.57 ;
      RECT 61.675 3.035 61.845 4.225 ;
      RECT 61.675 3.035 62.145 3.205 ;
      RECT 61.675 9.26 62.145 9.43 ;
      RECT 61.675 8.24 61.845 9.43 ;
      RECT 60.685 4.015 60.86 5.155 ;
      RECT 60.685 1.865 60.855 5.155 ;
      RECT 60.685 1.865 60.86 2.415 ;
      RECT 60.685 10.05 60.86 10.6 ;
      RECT 60.685 7.31 60.855 10.6 ;
      RECT 60.685 7.31 60.86 8.45 ;
      RECT 60.255 3.895 60.43 5.155 ;
      RECT 60.255 2.945 60.425 5.155 ;
      RECT 60.255 7.31 60.425 9.52 ;
      RECT 60.255 7.31 60.43 8.57 ;
      RECT 59.825 3.925 59.995 5.155 ;
      RECT 59.885 2.145 60.055 4.095 ;
      RECT 59.825 1.865 59.995 2.315 ;
      RECT 59.825 10.15 59.995 10.6 ;
      RECT 59.885 8.37 60.055 10.32 ;
      RECT 59.825 7.31 59.995 8.54 ;
      RECT 59.3 3.895 59.475 5.155 ;
      RECT 59.3 1.865 59.47 5.155 ;
      RECT 59.3 3.365 59.71 3.695 ;
      RECT 59.3 2.525 59.71 2.855 ;
      RECT 59.3 1.865 59.475 2.355 ;
      RECT 59.3 10.11 59.475 10.6 ;
      RECT 59.3 7.31 59.47 10.6 ;
      RECT 59.3 9.61 59.71 9.94 ;
      RECT 59.3 8.77 59.71 9.1 ;
      RECT 59.3 7.31 59.475 8.57 ;
      RECT 57.23 4.421 57.235 4.593 ;
      RECT 57.225 4.414 57.23 4.683 ;
      RECT 57.22 4.408 57.225 4.702 ;
      RECT 57.2 4.402 57.22 4.712 ;
      RECT 57.185 4.397 57.2 4.72 ;
      RECT 57.148 4.391 57.185 4.718 ;
      RECT 57.062 4.377 57.148 4.714 ;
      RECT 56.976 4.359 57.062 4.709 ;
      RECT 56.89 4.34 56.976 4.703 ;
      RECT 56.86 4.328 56.89 4.699 ;
      RECT 56.84 4.322 56.86 4.698 ;
      RECT 56.775 4.32 56.84 4.696 ;
      RECT 56.76 4.32 56.775 4.688 ;
      RECT 56.745 4.32 56.76 4.675 ;
      RECT 56.74 4.32 56.745 4.665 ;
      RECT 56.725 4.32 56.74 4.643 ;
      RECT 56.71 4.32 56.725 4.61 ;
      RECT 56.705 4.32 56.71 4.588 ;
      RECT 56.695 4.32 56.705 4.57 ;
      RECT 56.68 4.32 56.695 4.548 ;
      RECT 56.66 4.32 56.68 4.51 ;
      RECT 57.01 3.605 57.045 4.044 ;
      RECT 57.01 3.605 57.05 4.043 ;
      RECT 56.955 3.665 57.05 4.042 ;
      RECT 56.82 3.837 57.05 4.041 ;
      RECT 56.93 3.715 57.05 4.041 ;
      RECT 56.82 3.837 57.075 4.031 ;
      RECT 56.875 3.782 57.155 3.948 ;
      RECT 57.05 3.576 57.055 4.039 ;
      RECT 56.905 3.752 57.195 3.825 ;
      RECT 56.92 3.735 57.05 4.041 ;
      RECT 57.055 3.575 57.225 3.763 ;
      RECT 57.045 3.578 57.225 3.763 ;
      RECT 56.55 3.455 56.72 3.765 ;
      RECT 56.55 3.455 56.725 3.738 ;
      RECT 56.55 3.455 56.73 3.715 ;
      RECT 56.55 3.455 56.74 3.665 ;
      RECT 56.545 3.56 56.74 3.635 ;
      RECT 56.58 3.13 56.75 3.608 ;
      RECT 56.58 3.13 56.765 3.529 ;
      RECT 56.57 3.34 56.765 3.529 ;
      RECT 56.58 3.14 56.775 3.444 ;
      RECT 56.51 3.882 56.515 4.085 ;
      RECT 56.5 3.87 56.51 4.195 ;
      RECT 56.475 3.87 56.5 4.235 ;
      RECT 56.395 3.87 56.475 4.32 ;
      RECT 56.385 3.87 56.395 4.39 ;
      RECT 56.36 3.87 56.385 4.413 ;
      RECT 56.34 3.87 56.36 4.448 ;
      RECT 56.295 3.88 56.34 4.491 ;
      RECT 56.285 3.892 56.295 4.528 ;
      RECT 56.265 3.906 56.285 4.548 ;
      RECT 56.255 3.924 56.265 4.564 ;
      RECT 56.24 3.95 56.255 4.574 ;
      RECT 56.225 3.991 56.24 4.588 ;
      RECT 56.215 4.026 56.225 4.598 ;
      RECT 56.21 4.042 56.215 4.603 ;
      RECT 56.2 4.057 56.21 4.608 ;
      RECT 56.18 4.1 56.2 4.618 ;
      RECT 56.16 4.137 56.18 4.631 ;
      RECT 56.125 4.16 56.16 4.649 ;
      RECT 56.115 4.174 56.125 4.665 ;
      RECT 56.095 4.184 56.115 4.675 ;
      RECT 56.09 4.193 56.095 4.683 ;
      RECT 56.08 4.2 56.09 4.69 ;
      RECT 56.07 4.207 56.08 4.698 ;
      RECT 56.055 4.217 56.07 4.706 ;
      RECT 56.045 4.231 56.055 4.716 ;
      RECT 56.035 4.243 56.045 4.728 ;
      RECT 56.02 4.265 56.035 4.741 ;
      RECT 56.01 4.287 56.02 4.752 ;
      RECT 56 4.307 56.01 4.761 ;
      RECT 55.995 4.322 56 4.768 ;
      RECT 55.965 4.355 55.995 4.782 ;
      RECT 55.955 4.39 55.965 4.797 ;
      RECT 55.95 4.397 55.955 4.803 ;
      RECT 55.93 4.412 55.95 4.81 ;
      RECT 55.925 4.427 55.93 4.818 ;
      RECT 55.92 4.436 55.925 4.823 ;
      RECT 55.905 4.442 55.92 4.83 ;
      RECT 55.9 4.448 55.905 4.838 ;
      RECT 55.895 4.452 55.9 4.845 ;
      RECT 55.89 4.456 55.895 4.855 ;
      RECT 55.88 4.461 55.89 4.865 ;
      RECT 55.86 4.472 55.88 4.893 ;
      RECT 55.845 4.484 55.86 4.92 ;
      RECT 55.825 4.497 55.845 4.945 ;
      RECT 55.805 4.512 55.825 4.969 ;
      RECT 55.79 4.527 55.805 4.984 ;
      RECT 55.785 4.538 55.79 4.993 ;
      RECT 55.72 4.583 55.785 5.003 ;
      RECT 55.685 4.642 55.72 5.016 ;
      RECT 55.68 4.665 55.685 5.022 ;
      RECT 55.675 4.672 55.68 5.024 ;
      RECT 55.66 4.682 55.675 5.027 ;
      RECT 55.63 4.707 55.66 5.031 ;
      RECT 55.625 4.725 55.63 5.035 ;
      RECT 55.62 4.732 55.625 5.036 ;
      RECT 55.6 4.74 55.62 5.04 ;
      RECT 55.59 4.747 55.6 5.044 ;
      RECT 55.546 4.758 55.59 5.051 ;
      RECT 55.46 4.786 55.546 5.067 ;
      RECT 55.4 4.81 55.46 5.085 ;
      RECT 55.355 4.82 55.4 5.099 ;
      RECT 55.296 4.828 55.355 5.113 ;
      RECT 55.21 4.835 55.296 5.132 ;
      RECT 55.185 4.84 55.21 5.147 ;
      RECT 55.105 4.843 55.185 5.15 ;
      RECT 55.025 4.847 55.105 5.137 ;
      RECT 55.016 4.85 55.025 5.122 ;
      RECT 54.93 4.85 55.016 5.107 ;
      RECT 54.87 4.852 54.93 5.084 ;
      RECT 54.866 4.855 54.87 5.074 ;
      RECT 54.78 4.855 54.866 5.059 ;
      RECT 54.705 4.855 54.78 5.035 ;
      RECT 56.02 3.864 56.03 4.04 ;
      RECT 55.975 3.831 56.02 4.04 ;
      RECT 55.93 3.782 55.975 4.04 ;
      RECT 55.9 3.752 55.93 4.041 ;
      RECT 55.895 3.735 55.9 4.042 ;
      RECT 55.87 3.715 55.895 4.043 ;
      RECT 55.855 3.69 55.87 4.044 ;
      RECT 55.85 3.677 55.855 4.045 ;
      RECT 55.845 3.671 55.85 4.043 ;
      RECT 55.84 3.663 55.845 4.037 ;
      RECT 55.815 3.655 55.84 4.017 ;
      RECT 55.795 3.644 55.815 3.988 ;
      RECT 55.765 3.629 55.795 3.959 ;
      RECT 55.745 3.615 55.765 3.931 ;
      RECT 55.735 3.609 55.745 3.91 ;
      RECT 55.73 3.606 55.735 3.893 ;
      RECT 55.725 3.603 55.73 3.878 ;
      RECT 55.71 3.598 55.725 3.843 ;
      RECT 55.705 3.594 55.71 3.81 ;
      RECT 55.685 3.589 55.705 3.786 ;
      RECT 55.655 3.581 55.685 3.751 ;
      RECT 55.64 3.575 55.655 3.728 ;
      RECT 55.6 3.568 55.64 3.713 ;
      RECT 55.575 3.56 55.6 3.693 ;
      RECT 55.555 3.555 55.575 3.683 ;
      RECT 55.52 3.549 55.555 3.678 ;
      RECT 55.475 3.54 55.52 3.677 ;
      RECT 55.445 3.536 55.475 3.679 ;
      RECT 55.36 3.544 55.445 3.683 ;
      RECT 55.29 3.555 55.36 3.705 ;
      RECT 55.277 3.561 55.29 3.728 ;
      RECT 55.191 3.568 55.277 3.75 ;
      RECT 55.105 3.58 55.191 3.787 ;
      RECT 55.105 3.957 55.115 4.195 ;
      RECT 55.1 3.586 55.105 3.81 ;
      RECT 55.095 3.842 55.105 4.195 ;
      RECT 55.095 3.587 55.1 3.815 ;
      RECT 55.09 3.588 55.095 4.195 ;
      RECT 55.066 3.59 55.09 4.196 ;
      RECT 54.98 3.598 55.066 4.198 ;
      RECT 54.96 3.612 54.98 4.201 ;
      RECT 54.955 3.64 54.96 4.202 ;
      RECT 54.95 3.652 54.955 4.203 ;
      RECT 54.945 3.667 54.95 4.204 ;
      RECT 54.935 3.697 54.945 4.205 ;
      RECT 54.93 3.735 54.935 4.203 ;
      RECT 54.925 3.755 54.93 4.198 ;
      RECT 54.91 3.79 54.925 4.183 ;
      RECT 54.9 3.842 54.91 4.163 ;
      RECT 54.895 3.872 54.9 4.151 ;
      RECT 54.88 3.885 54.895 4.134 ;
      RECT 54.855 3.889 54.88 4.101 ;
      RECT 54.84 3.887 54.855 4.078 ;
      RECT 54.825 3.886 54.84 4.075 ;
      RECT 54.765 3.884 54.825 4.073 ;
      RECT 54.755 3.882 54.765 4.068 ;
      RECT 54.715 3.881 54.755 4.065 ;
      RECT 54.645 3.878 54.715 4.063 ;
      RECT 54.59 3.876 54.645 4.058 ;
      RECT 54.52 3.87 54.59 4.053 ;
      RECT 54.511 3.87 54.52 4.05 ;
      RECT 54.425 3.87 54.511 4.045 ;
      RECT 54.42 3.87 54.425 4.04 ;
      RECT 55.725 3.105 55.9 3.455 ;
      RECT 55.725 3.12 55.91 3.453 ;
      RECT 55.7 3.07 55.845 3.45 ;
      RECT 55.68 3.071 55.845 3.443 ;
      RECT 55.67 3.072 55.855 3.438 ;
      RECT 55.64 3.073 55.855 3.425 ;
      RECT 55.59 3.074 55.855 3.401 ;
      RECT 55.585 3.076 55.855 3.386 ;
      RECT 55.585 3.142 55.915 3.38 ;
      RECT 55.565 3.083 55.87 3.36 ;
      RECT 55.555 3.092 55.88 3.215 ;
      RECT 55.565 3.087 55.88 3.36 ;
      RECT 55.585 3.077 55.87 3.386 ;
      RECT 55.17 4.402 55.34 4.69 ;
      RECT 55.165 4.42 55.35 4.685 ;
      RECT 55.13 4.428 55.415 4.605 ;
      RECT 55.13 4.428 55.501 4.595 ;
      RECT 55.13 4.428 55.555 4.541 ;
      RECT 55.415 4.325 55.585 4.509 ;
      RECT 55.13 4.48 55.59 4.497 ;
      RECT 55.115 4.45 55.585 4.493 ;
      RECT 55.375 4.332 55.415 4.644 ;
      RECT 55.255 4.369 55.585 4.509 ;
      RECT 55.35 4.344 55.375 4.67 ;
      RECT 55.34 4.351 55.585 4.509 ;
      RECT 55.471 3.815 55.54 4.074 ;
      RECT 55.471 3.87 55.545 4.073 ;
      RECT 55.385 3.87 55.545 4.072 ;
      RECT 55.38 3.87 55.55 4.065 ;
      RECT 55.37 3.815 55.54 4.06 ;
      RECT 55.05 10.05 55.225 10.6 ;
      RECT 55.05 7.31 55.22 10.6 ;
      RECT 55.05 7.31 55.225 8.45 ;
      RECT 54.75 3.114 54.925 3.415 ;
      RECT 54.735 3.102 54.75 3.4 ;
      RECT 54.705 3.101 54.735 3.353 ;
      RECT 54.705 3.119 54.93 3.348 ;
      RECT 54.69 3.103 54.75 3.313 ;
      RECT 54.685 3.125 54.94 3.213 ;
      RECT 54.685 3.108 54.836 3.213 ;
      RECT 54.685 3.11 54.84 3.213 ;
      RECT 54.69 3.106 54.836 3.313 ;
      RECT 54.795 4.342 54.8 4.69 ;
      RECT 54.785 4.332 54.795 4.696 ;
      RECT 54.75 4.322 54.785 4.698 ;
      RECT 54.712 4.317 54.75 4.702 ;
      RECT 54.626 4.31 54.712 4.709 ;
      RECT 54.54 4.3 54.626 4.719 ;
      RECT 54.495 4.295 54.54 4.727 ;
      RECT 54.491 4.295 54.495 4.731 ;
      RECT 54.405 4.295 54.491 4.738 ;
      RECT 54.39 4.295 54.405 4.738 ;
      RECT 54.38 4.293 54.39 4.71 ;
      RECT 54.37 4.289 54.38 4.653 ;
      RECT 54.35 4.283 54.37 4.585 ;
      RECT 54.345 4.279 54.35 4.533 ;
      RECT 54.335 4.278 54.345 4.5 ;
      RECT 54.285 4.276 54.335 4.485 ;
      RECT 54.26 4.274 54.285 4.48 ;
      RECT 54.217 4.272 54.26 4.476 ;
      RECT 54.131 4.268 54.217 4.464 ;
      RECT 54.045 4.263 54.131 4.448 ;
      RECT 54.015 4.26 54.045 4.435 ;
      RECT 53.99 4.259 54.015 4.423 ;
      RECT 53.985 4.259 53.99 4.413 ;
      RECT 53.945 4.258 53.985 4.405 ;
      RECT 53.93 4.257 53.945 4.398 ;
      RECT 53.88 4.256 53.93 4.39 ;
      RECT 53.878 4.255 53.88 4.385 ;
      RECT 53.792 4.253 53.878 4.385 ;
      RECT 53.706 4.248 53.792 4.385 ;
      RECT 53.62 4.244 53.706 4.385 ;
      RECT 53.571 4.24 53.62 4.383 ;
      RECT 53.485 4.237 53.571 4.378 ;
      RECT 53.462 4.234 53.485 4.374 ;
      RECT 53.376 4.231 53.462 4.369 ;
      RECT 53.29 4.227 53.376 4.36 ;
      RECT 53.265 4.22 53.29 4.355 ;
      RECT 53.205 4.185 53.265 4.352 ;
      RECT 53.185 4.11 53.205 4.349 ;
      RECT 53.18 4.052 53.185 4.348 ;
      RECT 53.155 3.992 53.18 4.347 ;
      RECT 53.08 3.87 53.155 4.343 ;
      RECT 53.07 3.87 53.08 4.335 ;
      RECT 53.055 3.87 53.07 4.325 ;
      RECT 53.04 3.87 53.055 4.295 ;
      RECT 53.025 3.87 53.04 4.24 ;
      RECT 53.01 3.87 53.025 4.178 ;
      RECT 52.985 3.87 53.01 4.103 ;
      RECT 52.98 3.87 52.985 4.053 ;
      RECT 54.62 7.31 54.79 9.52 ;
      RECT 54.62 7.31 54.795 8.57 ;
      RECT 54.325 3.415 54.345 3.724 ;
      RECT 54.311 3.417 54.36 3.721 ;
      RECT 54.311 3.422 54.38 3.712 ;
      RECT 54.225 3.42 54.36 3.706 ;
      RECT 54.225 3.428 54.415 3.689 ;
      RECT 54.19 3.43 54.415 3.688 ;
      RECT 54.16 3.438 54.415 3.679 ;
      RECT 54.15 3.443 54.435 3.665 ;
      RECT 54.19 3.433 54.435 3.665 ;
      RECT 54.19 3.436 54.445 3.653 ;
      RECT 54.16 3.438 54.455 3.64 ;
      RECT 54.16 3.442 54.465 3.583 ;
      RECT 54.15 3.447 54.47 3.498 ;
      RECT 54.311 3.415 54.345 3.721 ;
      RECT 53.75 3.518 53.755 3.73 ;
      RECT 53.625 3.515 53.64 3.73 ;
      RECT 53.09 3.545 53.16 3.73 ;
      RECT 52.975 3.545 53.01 3.725 ;
      RECT 54.096 3.847 54.115 4.041 ;
      RECT 54.01 3.802 54.096 4.042 ;
      RECT 54 3.755 54.01 4.044 ;
      RECT 53.995 3.735 54 4.045 ;
      RECT 53.975 3.7 53.995 4.046 ;
      RECT 53.96 3.65 53.975 4.047 ;
      RECT 53.94 3.587 53.96 4.048 ;
      RECT 53.93 3.55 53.94 4.049 ;
      RECT 53.915 3.539 53.93 4.05 ;
      RECT 53.91 3.531 53.915 4.048 ;
      RECT 53.9 3.53 53.91 4.04 ;
      RECT 53.87 3.527 53.9 4.019 ;
      RECT 53.795 3.522 53.87 3.964 ;
      RECT 53.78 3.518 53.795 3.91 ;
      RECT 53.77 3.518 53.78 3.805 ;
      RECT 53.755 3.518 53.77 3.738 ;
      RECT 53.74 3.518 53.75 3.728 ;
      RECT 53.685 3.517 53.74 3.725 ;
      RECT 53.64 3.515 53.685 3.728 ;
      RECT 53.612 3.515 53.625 3.731 ;
      RECT 53.526 3.519 53.612 3.733 ;
      RECT 53.44 3.525 53.526 3.738 ;
      RECT 53.42 3.529 53.44 3.74 ;
      RECT 53.418 3.53 53.42 3.739 ;
      RECT 53.332 3.532 53.418 3.738 ;
      RECT 53.246 3.537 53.332 3.735 ;
      RECT 53.16 3.542 53.246 3.732 ;
      RECT 53.01 3.545 53.09 3.728 ;
      RECT 53.665 10.11 53.84 10.6 ;
      RECT 53.665 7.31 53.835 10.6 ;
      RECT 53.665 9.61 54.075 9.94 ;
      RECT 53.665 8.77 54.075 9.1 ;
      RECT 53.665 7.31 53.84 8.57 ;
      RECT 53.786 4.52 53.835 4.854 ;
      RECT 53.786 4.52 53.84 4.853 ;
      RECT 53.7 4.52 53.84 4.852 ;
      RECT 53.475 4.628 53.845 4.85 ;
      RECT 53.7 4.52 53.87 4.843 ;
      RECT 53.67 4.532 53.875 4.834 ;
      RECT 53.655 4.55 53.88 4.831 ;
      RECT 53.47 4.634 53.88 4.758 ;
      RECT 53.465 4.641 53.88 4.718 ;
      RECT 53.48 4.607 53.88 4.831 ;
      RECT 53.641 4.553 53.845 4.85 ;
      RECT 53.555 4.573 53.88 4.831 ;
      RECT 53.655 4.547 53.875 4.834 ;
      RECT 53.425 3.871 53.615 4.065 ;
      RECT 53.42 3.873 53.615 4.064 ;
      RECT 53.415 3.877 53.63 4.061 ;
      RECT 53.43 3.87 53.63 4.061 ;
      RECT 53.415 3.98 53.635 4.056 ;
      RECT 52.71 4.48 52.801 4.778 ;
      RECT 52.705 4.482 52.88 4.773 ;
      RECT 52.71 4.48 52.88 4.773 ;
      RECT 52.705 4.486 52.9 4.771 ;
      RECT 52.705 4.541 52.94 4.77 ;
      RECT 52.705 4.576 52.955 4.764 ;
      RECT 52.705 4.61 52.965 4.754 ;
      RECT 52.695 4.49 52.9 4.605 ;
      RECT 52.695 4.51 52.915 4.605 ;
      RECT 52.695 4.493 52.905 4.605 ;
      RECT 52.92 3.261 52.925 3.323 ;
      RECT 52.915 3.183 52.92 3.346 ;
      RECT 52.91 3.14 52.915 3.357 ;
      RECT 52.905 3.13 52.91 3.369 ;
      RECT 52.9 3.13 52.905 3.378 ;
      RECT 52.875 3.13 52.9 3.41 ;
      RECT 52.87 3.13 52.875 3.443 ;
      RECT 52.855 3.13 52.87 3.468 ;
      RECT 52.845 3.13 52.855 3.495 ;
      RECT 52.84 3.13 52.845 3.508 ;
      RECT 52.835 3.13 52.84 3.523 ;
      RECT 52.825 3.13 52.835 3.538 ;
      RECT 52.82 3.13 52.825 3.558 ;
      RECT 52.795 3.13 52.82 3.593 ;
      RECT 52.75 3.13 52.795 3.638 ;
      RECT 52.74 3.13 52.75 3.651 ;
      RECT 52.655 3.215 52.74 3.658 ;
      RECT 52.62 3.337 52.655 3.667 ;
      RECT 52.615 3.377 52.62 3.671 ;
      RECT 52.595 3.4 52.615 3.673 ;
      RECT 52.59 3.43 52.595 3.676 ;
      RECT 52.58 3.442 52.59 3.677 ;
      RECT 52.535 3.465 52.58 3.682 ;
      RECT 52.495 3.495 52.535 3.69 ;
      RECT 52.46 3.507 52.495 3.696 ;
      RECT 52.455 3.512 52.46 3.7 ;
      RECT 52.385 3.522 52.455 3.707 ;
      RECT 52.345 3.532 52.385 3.717 ;
      RECT 52.325 3.537 52.345 3.723 ;
      RECT 52.315 3.541 52.325 3.728 ;
      RECT 52.31 3.544 52.315 3.731 ;
      RECT 52.3 3.545 52.31 3.732 ;
      RECT 52.275 3.547 52.3 3.736 ;
      RECT 52.265 3.552 52.275 3.739 ;
      RECT 52.22 3.56 52.265 3.74 ;
      RECT 52.095 3.565 52.22 3.74 ;
      RECT 52.65 3.862 52.67 4.044 ;
      RECT 52.601 3.847 52.65 4.043 ;
      RECT 52.515 3.862 52.67 4.041 ;
      RECT 52.5 3.862 52.67 4.04 ;
      RECT 52.465 3.84 52.635 4.025 ;
      RECT 52.535 4.86 52.55 5.069 ;
      RECT 52.535 4.868 52.555 5.068 ;
      RECT 52.48 4.868 52.555 5.067 ;
      RECT 52.46 4.872 52.56 5.065 ;
      RECT 52.44 4.822 52.48 5.064 ;
      RECT 52.385 4.88 52.565 5.062 ;
      RECT 52.35 4.837 52.48 5.06 ;
      RECT 52.346 4.84 52.535 5.059 ;
      RECT 52.26 4.848 52.535 5.057 ;
      RECT 52.26 4.892 52.57 5.05 ;
      RECT 52.25 4.985 52.57 5.048 ;
      RECT 52.26 4.904 52.575 5.033 ;
      RECT 52.26 4.925 52.59 5.003 ;
      RECT 52.26 4.952 52.595 4.973 ;
      RECT 52.385 4.83 52.48 5.062 ;
      RECT 52.015 3.875 52.02 4.413 ;
      RECT 51.82 4.205 51.825 4.4 ;
      RECT 50.12 3.87 50.135 4.25 ;
      RECT 52.185 3.87 52.19 4.04 ;
      RECT 52.18 3.87 52.185 4.05 ;
      RECT 52.175 3.87 52.18 4.063 ;
      RECT 52.15 3.87 52.175 4.105 ;
      RECT 52.125 3.87 52.15 4.178 ;
      RECT 52.11 3.87 52.125 4.23 ;
      RECT 52.105 3.87 52.11 4.26 ;
      RECT 52.08 3.87 52.105 4.3 ;
      RECT 52.065 3.87 52.08 4.355 ;
      RECT 52.06 3.87 52.065 4.388 ;
      RECT 52.035 3.87 52.06 4.408 ;
      RECT 52.02 3.87 52.035 4.414 ;
      RECT 51.95 3.905 52.015 4.41 ;
      RECT 51.9 3.96 51.95 4.405 ;
      RECT 51.89 3.992 51.9 4.403 ;
      RECT 51.885 4.017 51.89 4.403 ;
      RECT 51.865 4.09 51.885 4.403 ;
      RECT 51.855 4.17 51.865 4.402 ;
      RECT 51.84 4.2 51.855 4.402 ;
      RECT 51.825 4.205 51.84 4.401 ;
      RECT 51.765 4.207 51.82 4.398 ;
      RECT 51.735 4.212 51.765 4.394 ;
      RECT 51.733 4.215 51.735 4.393 ;
      RECT 51.647 4.217 51.733 4.39 ;
      RECT 51.561 4.223 51.647 4.384 ;
      RECT 51.475 4.228 51.561 4.378 ;
      RECT 51.402 4.233 51.475 4.379 ;
      RECT 51.316 4.239 51.402 4.387 ;
      RECT 51.23 4.245 51.316 4.396 ;
      RECT 51.21 4.249 51.23 4.401 ;
      RECT 51.163 4.251 51.21 4.404 ;
      RECT 51.077 4.256 51.163 4.41 ;
      RECT 50.991 4.261 51.077 4.419 ;
      RECT 50.905 4.267 50.991 4.427 ;
      RECT 50.82 4.265 50.905 4.436 ;
      RECT 50.816 4.26 50.82 4.44 ;
      RECT 50.73 4.255 50.816 4.432 ;
      RECT 50.666 4.246 50.73 4.42 ;
      RECT 50.58 4.237 50.666 4.407 ;
      RECT 50.556 4.23 50.58 4.398 ;
      RECT 50.47 4.224 50.556 4.385 ;
      RECT 50.43 4.217 50.47 4.371 ;
      RECT 50.425 4.207 50.43 4.367 ;
      RECT 50.415 4.195 50.425 4.366 ;
      RECT 50.395 4.165 50.415 4.363 ;
      RECT 50.34 4.085 50.395 4.357 ;
      RECT 50.32 4.004 50.34 4.352 ;
      RECT 50.3 3.962 50.32 4.348 ;
      RECT 50.275 3.915 50.3 4.342 ;
      RECT 50.27 3.89 50.275 4.339 ;
      RECT 50.235 3.87 50.27 4.334 ;
      RECT 50.226 3.87 50.235 4.327 ;
      RECT 50.14 3.87 50.226 4.297 ;
      RECT 50.135 3.87 50.14 4.26 ;
      RECT 50.1 3.87 50.12 4.182 ;
      RECT 50.095 3.912 50.1 4.147 ;
      RECT 50.09 3.987 50.095 4.103 ;
      RECT 51.54 3.792 51.715 4.04 ;
      RECT 51.54 3.792 51.72 4.038 ;
      RECT 51.535 3.824 51.72 3.998 ;
      RECT 51.565 3.765 51.735 3.985 ;
      RECT 51.53 3.842 51.735 3.918 ;
      RECT 50.84 3.305 51.01 3.48 ;
      RECT 50.84 3.305 51.182 3.472 ;
      RECT 50.84 3.305 51.265 3.466 ;
      RECT 50.84 3.305 51.3 3.462 ;
      RECT 50.84 3.305 51.32 3.461 ;
      RECT 50.84 3.305 51.406 3.457 ;
      RECT 51.3 3.13 51.47 3.452 ;
      RECT 50.875 3.237 51.5 3.45 ;
      RECT 50.865 3.292 51.505 3.448 ;
      RECT 50.84 3.328 51.515 3.443 ;
      RECT 50.84 3.355 51.52 3.373 ;
      RECT 50.905 3.18 51.48 3.45 ;
      RECT 51.096 3.165 51.48 3.45 ;
      RECT 50.93 3.168 51.48 3.45 ;
      RECT 51.01 3.166 51.096 3.477 ;
      RECT 51.096 3.163 51.475 3.45 ;
      RECT 51.28 3.14 51.475 3.45 ;
      RECT 51.182 3.161 51.475 3.45 ;
      RECT 51.265 3.155 51.28 3.463 ;
      RECT 51.415 4.52 51.42 4.72 ;
      RECT 50.88 4.585 50.925 4.72 ;
      RECT 51.45 4.52 51.47 4.693 ;
      RECT 51.42 4.52 51.45 4.708 ;
      RECT 51.355 4.52 51.415 4.745 ;
      RECT 51.34 4.52 51.355 4.775 ;
      RECT 51.325 4.52 51.34 4.788 ;
      RECT 51.305 4.52 51.325 4.803 ;
      RECT 51.3 4.52 51.305 4.812 ;
      RECT 51.29 4.524 51.3 4.817 ;
      RECT 51.275 4.534 51.29 4.828 ;
      RECT 51.25 4.55 51.275 4.838 ;
      RECT 51.24 4.564 51.25 4.84 ;
      RECT 51.22 4.576 51.24 4.837 ;
      RECT 51.19 4.597 51.22 4.831 ;
      RECT 51.18 4.609 51.19 4.826 ;
      RECT 51.17 4.607 51.18 4.823 ;
      RECT 51.155 4.606 51.17 4.818 ;
      RECT 51.15 4.605 51.155 4.813 ;
      RECT 51.115 4.603 51.15 4.803 ;
      RECT 51.095 4.6 51.115 4.785 ;
      RECT 51.085 4.598 51.095 4.78 ;
      RECT 51.075 4.597 51.085 4.775 ;
      RECT 51.04 4.595 51.075 4.763 ;
      RECT 50.985 4.591 51.04 4.743 ;
      RECT 50.975 4.589 50.985 4.728 ;
      RECT 50.97 4.589 50.975 4.723 ;
      RECT 50.925 4.587 50.97 4.72 ;
      RECT 50.83 4.585 50.88 4.724 ;
      RECT 50.82 4.586 50.83 4.729 ;
      RECT 50.76 4.593 50.82 4.743 ;
      RECT 50.735 4.601 50.76 4.763 ;
      RECT 50.725 4.605 50.735 4.775 ;
      RECT 50.72 4.606 50.725 4.78 ;
      RECT 50.705 4.608 50.72 4.783 ;
      RECT 50.69 4.61 50.705 4.788 ;
      RECT 50.685 4.61 50.69 4.791 ;
      RECT 50.64 4.615 50.685 4.802 ;
      RECT 50.635 4.619 50.64 4.814 ;
      RECT 50.61 4.615 50.635 4.818 ;
      RECT 50.6 4.611 50.61 4.822 ;
      RECT 50.59 4.61 50.6 4.826 ;
      RECT 50.575 4.6 50.59 4.832 ;
      RECT 50.57 4.588 50.575 4.836 ;
      RECT 50.565 4.585 50.57 4.837 ;
      RECT 50.56 4.582 50.565 4.839 ;
      RECT 50.545 4.57 50.56 4.838 ;
      RECT 50.53 4.552 50.545 4.835 ;
      RECT 50.51 4.531 50.53 4.828 ;
      RECT 50.445 4.52 50.51 4.8 ;
      RECT 50.441 4.52 50.445 4.779 ;
      RECT 50.355 4.52 50.441 4.749 ;
      RECT 50.34 4.52 50.355 4.705 ;
      RECT 50.99 4.871 51.005 5.13 ;
      RECT 50.99 4.886 51.01 5.129 ;
      RECT 50.906 4.886 51.01 5.127 ;
      RECT 50.906 4.9 51.015 5.126 ;
      RECT 50.82 4.942 51.02 5.123 ;
      RECT 50.815 4.885 51.005 5.118 ;
      RECT 50.815 4.956 51.025 5.115 ;
      RECT 50.81 4.987 51.025 5.113 ;
      RECT 50.815 4.984 51.04 5.103 ;
      RECT 50.81 5.03 51.055 5.088 ;
      RECT 50.81 5.058 51.06 5.073 ;
      RECT 50.82 4.86 50.99 5.123 ;
      RECT 50.58 3.87 50.75 4.04 ;
      RECT 50.545 3.87 50.75 4.035 ;
      RECT 50.535 3.87 50.75 4.028 ;
      RECT 50.53 3.855 50.7 4.025 ;
      RECT 49.36 4.392 49.625 4.835 ;
      RECT 49.355 4.363 49.57 4.833 ;
      RECT 49.35 4.517 49.63 4.828 ;
      RECT 49.355 4.412 49.63 4.828 ;
      RECT 49.355 4.423 49.64 4.815 ;
      RECT 49.355 4.37 49.6 4.833 ;
      RECT 49.36 4.357 49.57 4.835 ;
      RECT 49.36 4.355 49.52 4.835 ;
      RECT 49.461 4.347 49.52 4.835 ;
      RECT 49.375 4.348 49.52 4.835 ;
      RECT 49.461 4.346 49.51 4.835 ;
      RECT 49.265 3.161 49.44 3.46 ;
      RECT 49.315 3.123 49.44 3.46 ;
      RECT 49.3 3.125 49.526 3.452 ;
      RECT 49.3 3.128 49.565 3.439 ;
      RECT 49.3 3.129 49.575 3.425 ;
      RECT 49.255 3.18 49.575 3.415 ;
      RECT 49.3 3.13 49.58 3.41 ;
      RECT 49.255 3.34 49.585 3.4 ;
      RECT 49.24 3.2 49.58 3.34 ;
      RECT 49.235 3.216 49.58 3.28 ;
      RECT 49.28 3.14 49.58 3.41 ;
      RECT 49.315 3.121 49.401 3.46 ;
      RECT 47.775 7.31 47.945 8.78 ;
      RECT 47.775 7.31 47.95 8.57 ;
      RECT 47.405 9.26 47.875 9.43 ;
      RECT 47.405 8.24 47.575 9.43 ;
      RECT 47.4 3.035 47.57 4.225 ;
      RECT 47.4 3.035 47.87 3.205 ;
      RECT 46.785 3.895 46.96 5.155 ;
      RECT 46.785 3.685 46.955 5.155 ;
      RECT 46.785 7.31 46.955 8.78 ;
      RECT 46.785 7.31 46.96 8.57 ;
      RECT 46.415 3.035 46.585 4.225 ;
      RECT 46.415 3.035 46.885 3.205 ;
      RECT 46.415 9.26 46.885 9.43 ;
      RECT 46.415 8.24 46.585 9.43 ;
      RECT 45.425 4.015 45.6 5.155 ;
      RECT 45.425 1.865 45.595 5.155 ;
      RECT 45.425 1.865 45.6 2.415 ;
      RECT 45.425 10.05 45.6 10.6 ;
      RECT 45.425 7.31 45.595 10.6 ;
      RECT 45.425 7.31 45.6 8.45 ;
      RECT 44.995 3.895 45.17 5.155 ;
      RECT 44.995 2.945 45.165 5.155 ;
      RECT 44.995 7.31 45.165 9.52 ;
      RECT 44.995 7.31 45.17 8.57 ;
      RECT 44.565 3.925 44.735 5.155 ;
      RECT 44.625 2.145 44.795 4.095 ;
      RECT 44.565 1.865 44.735 2.315 ;
      RECT 44.565 10.15 44.735 10.6 ;
      RECT 44.625 8.37 44.795 10.32 ;
      RECT 44.565 7.31 44.735 8.54 ;
      RECT 44.04 3.895 44.215 5.155 ;
      RECT 44.04 1.865 44.21 5.155 ;
      RECT 44.04 3.365 44.45 3.695 ;
      RECT 44.04 2.525 44.45 2.855 ;
      RECT 44.04 1.865 44.215 2.355 ;
      RECT 44.04 10.11 44.215 10.6 ;
      RECT 44.04 7.31 44.21 10.6 ;
      RECT 44.04 9.61 44.45 9.94 ;
      RECT 44.04 8.77 44.45 9.1 ;
      RECT 44.04 7.31 44.215 8.57 ;
      RECT 41.97 4.421 41.975 4.593 ;
      RECT 41.965 4.414 41.97 4.683 ;
      RECT 41.96 4.408 41.965 4.702 ;
      RECT 41.94 4.402 41.96 4.712 ;
      RECT 41.925 4.397 41.94 4.72 ;
      RECT 41.888 4.391 41.925 4.718 ;
      RECT 41.802 4.377 41.888 4.714 ;
      RECT 41.716 4.359 41.802 4.709 ;
      RECT 41.63 4.34 41.716 4.703 ;
      RECT 41.6 4.328 41.63 4.699 ;
      RECT 41.58 4.322 41.6 4.698 ;
      RECT 41.515 4.32 41.58 4.696 ;
      RECT 41.5 4.32 41.515 4.688 ;
      RECT 41.485 4.32 41.5 4.675 ;
      RECT 41.48 4.32 41.485 4.665 ;
      RECT 41.465 4.32 41.48 4.643 ;
      RECT 41.45 4.32 41.465 4.61 ;
      RECT 41.445 4.32 41.45 4.588 ;
      RECT 41.435 4.32 41.445 4.57 ;
      RECT 41.42 4.32 41.435 4.548 ;
      RECT 41.4 4.32 41.42 4.51 ;
      RECT 41.75 3.605 41.785 4.044 ;
      RECT 41.75 3.605 41.79 4.043 ;
      RECT 41.695 3.665 41.79 4.042 ;
      RECT 41.56 3.837 41.79 4.041 ;
      RECT 41.67 3.715 41.79 4.041 ;
      RECT 41.56 3.837 41.815 4.031 ;
      RECT 41.615 3.782 41.895 3.948 ;
      RECT 41.79 3.576 41.795 4.039 ;
      RECT 41.645 3.752 41.935 3.825 ;
      RECT 41.66 3.735 41.79 4.041 ;
      RECT 41.795 3.575 41.965 3.763 ;
      RECT 41.785 3.578 41.965 3.763 ;
      RECT 41.29 3.455 41.46 3.765 ;
      RECT 41.29 3.455 41.465 3.738 ;
      RECT 41.29 3.455 41.47 3.715 ;
      RECT 41.29 3.455 41.48 3.665 ;
      RECT 41.285 3.56 41.48 3.635 ;
      RECT 41.32 3.13 41.49 3.608 ;
      RECT 41.32 3.13 41.505 3.529 ;
      RECT 41.31 3.34 41.505 3.529 ;
      RECT 41.32 3.14 41.515 3.444 ;
      RECT 41.25 3.882 41.255 4.085 ;
      RECT 41.24 3.87 41.25 4.195 ;
      RECT 41.215 3.87 41.24 4.235 ;
      RECT 41.135 3.87 41.215 4.32 ;
      RECT 41.125 3.87 41.135 4.39 ;
      RECT 41.1 3.87 41.125 4.413 ;
      RECT 41.08 3.87 41.1 4.448 ;
      RECT 41.035 3.88 41.08 4.491 ;
      RECT 41.025 3.892 41.035 4.528 ;
      RECT 41.005 3.906 41.025 4.548 ;
      RECT 40.995 3.924 41.005 4.564 ;
      RECT 40.98 3.95 40.995 4.574 ;
      RECT 40.965 3.991 40.98 4.588 ;
      RECT 40.955 4.026 40.965 4.598 ;
      RECT 40.95 4.042 40.955 4.603 ;
      RECT 40.94 4.057 40.95 4.608 ;
      RECT 40.92 4.1 40.94 4.618 ;
      RECT 40.9 4.137 40.92 4.631 ;
      RECT 40.865 4.16 40.9 4.649 ;
      RECT 40.855 4.174 40.865 4.665 ;
      RECT 40.835 4.184 40.855 4.675 ;
      RECT 40.83 4.193 40.835 4.683 ;
      RECT 40.82 4.2 40.83 4.69 ;
      RECT 40.81 4.207 40.82 4.698 ;
      RECT 40.795 4.217 40.81 4.706 ;
      RECT 40.785 4.231 40.795 4.716 ;
      RECT 40.775 4.243 40.785 4.728 ;
      RECT 40.76 4.265 40.775 4.741 ;
      RECT 40.75 4.287 40.76 4.752 ;
      RECT 40.74 4.307 40.75 4.761 ;
      RECT 40.735 4.322 40.74 4.768 ;
      RECT 40.705 4.355 40.735 4.782 ;
      RECT 40.695 4.39 40.705 4.797 ;
      RECT 40.69 4.397 40.695 4.803 ;
      RECT 40.67 4.412 40.69 4.81 ;
      RECT 40.665 4.427 40.67 4.818 ;
      RECT 40.66 4.436 40.665 4.823 ;
      RECT 40.645 4.442 40.66 4.83 ;
      RECT 40.64 4.448 40.645 4.838 ;
      RECT 40.635 4.452 40.64 4.845 ;
      RECT 40.63 4.456 40.635 4.855 ;
      RECT 40.62 4.461 40.63 4.865 ;
      RECT 40.6 4.472 40.62 4.893 ;
      RECT 40.585 4.484 40.6 4.92 ;
      RECT 40.565 4.497 40.585 4.945 ;
      RECT 40.545 4.512 40.565 4.969 ;
      RECT 40.53 4.527 40.545 4.984 ;
      RECT 40.525 4.538 40.53 4.993 ;
      RECT 40.46 4.583 40.525 5.003 ;
      RECT 40.425 4.642 40.46 5.016 ;
      RECT 40.42 4.665 40.425 5.022 ;
      RECT 40.415 4.672 40.42 5.024 ;
      RECT 40.4 4.682 40.415 5.027 ;
      RECT 40.37 4.707 40.4 5.031 ;
      RECT 40.365 4.725 40.37 5.035 ;
      RECT 40.36 4.732 40.365 5.036 ;
      RECT 40.34 4.74 40.36 5.04 ;
      RECT 40.33 4.747 40.34 5.044 ;
      RECT 40.286 4.758 40.33 5.051 ;
      RECT 40.2 4.786 40.286 5.067 ;
      RECT 40.14 4.81 40.2 5.085 ;
      RECT 40.095 4.82 40.14 5.099 ;
      RECT 40.036 4.828 40.095 5.113 ;
      RECT 39.95 4.835 40.036 5.132 ;
      RECT 39.925 4.84 39.95 5.147 ;
      RECT 39.845 4.843 39.925 5.15 ;
      RECT 39.765 4.847 39.845 5.137 ;
      RECT 39.756 4.85 39.765 5.122 ;
      RECT 39.67 4.85 39.756 5.107 ;
      RECT 39.61 4.852 39.67 5.084 ;
      RECT 39.606 4.855 39.61 5.074 ;
      RECT 39.52 4.855 39.606 5.059 ;
      RECT 39.445 4.855 39.52 5.035 ;
      RECT 40.76 3.864 40.77 4.04 ;
      RECT 40.715 3.831 40.76 4.04 ;
      RECT 40.67 3.782 40.715 4.04 ;
      RECT 40.64 3.752 40.67 4.041 ;
      RECT 40.635 3.735 40.64 4.042 ;
      RECT 40.61 3.715 40.635 4.043 ;
      RECT 40.595 3.69 40.61 4.044 ;
      RECT 40.59 3.677 40.595 4.045 ;
      RECT 40.585 3.671 40.59 4.043 ;
      RECT 40.58 3.663 40.585 4.037 ;
      RECT 40.555 3.655 40.58 4.017 ;
      RECT 40.535 3.644 40.555 3.988 ;
      RECT 40.505 3.629 40.535 3.959 ;
      RECT 40.485 3.615 40.505 3.931 ;
      RECT 40.475 3.609 40.485 3.91 ;
      RECT 40.47 3.606 40.475 3.893 ;
      RECT 40.465 3.603 40.47 3.878 ;
      RECT 40.45 3.598 40.465 3.843 ;
      RECT 40.445 3.594 40.45 3.81 ;
      RECT 40.425 3.589 40.445 3.786 ;
      RECT 40.395 3.581 40.425 3.751 ;
      RECT 40.38 3.575 40.395 3.728 ;
      RECT 40.34 3.568 40.38 3.713 ;
      RECT 40.315 3.56 40.34 3.693 ;
      RECT 40.295 3.555 40.315 3.683 ;
      RECT 40.26 3.549 40.295 3.678 ;
      RECT 40.215 3.54 40.26 3.677 ;
      RECT 40.185 3.536 40.215 3.679 ;
      RECT 40.1 3.544 40.185 3.683 ;
      RECT 40.03 3.555 40.1 3.705 ;
      RECT 40.017 3.561 40.03 3.728 ;
      RECT 39.931 3.568 40.017 3.75 ;
      RECT 39.845 3.58 39.931 3.787 ;
      RECT 39.845 3.957 39.855 4.195 ;
      RECT 39.84 3.586 39.845 3.81 ;
      RECT 39.835 3.842 39.845 4.195 ;
      RECT 39.835 3.587 39.84 3.815 ;
      RECT 39.83 3.588 39.835 4.195 ;
      RECT 39.806 3.59 39.83 4.196 ;
      RECT 39.72 3.598 39.806 4.198 ;
      RECT 39.7 3.612 39.72 4.201 ;
      RECT 39.695 3.64 39.7 4.202 ;
      RECT 39.69 3.652 39.695 4.203 ;
      RECT 39.685 3.667 39.69 4.204 ;
      RECT 39.675 3.697 39.685 4.205 ;
      RECT 39.67 3.735 39.675 4.203 ;
      RECT 39.665 3.755 39.67 4.198 ;
      RECT 39.65 3.79 39.665 4.183 ;
      RECT 39.64 3.842 39.65 4.163 ;
      RECT 39.635 3.872 39.64 4.151 ;
      RECT 39.62 3.885 39.635 4.134 ;
      RECT 39.595 3.889 39.62 4.101 ;
      RECT 39.58 3.887 39.595 4.078 ;
      RECT 39.565 3.886 39.58 4.075 ;
      RECT 39.505 3.884 39.565 4.073 ;
      RECT 39.495 3.882 39.505 4.068 ;
      RECT 39.455 3.881 39.495 4.065 ;
      RECT 39.385 3.878 39.455 4.063 ;
      RECT 39.33 3.876 39.385 4.058 ;
      RECT 39.26 3.87 39.33 4.053 ;
      RECT 39.251 3.87 39.26 4.05 ;
      RECT 39.165 3.87 39.251 4.045 ;
      RECT 39.16 3.87 39.165 4.04 ;
      RECT 40.465 3.105 40.64 3.455 ;
      RECT 40.465 3.12 40.65 3.453 ;
      RECT 40.44 3.07 40.585 3.45 ;
      RECT 40.42 3.071 40.585 3.443 ;
      RECT 40.41 3.072 40.595 3.438 ;
      RECT 40.38 3.073 40.595 3.425 ;
      RECT 40.33 3.074 40.595 3.401 ;
      RECT 40.325 3.076 40.595 3.386 ;
      RECT 40.325 3.142 40.655 3.38 ;
      RECT 40.305 3.083 40.61 3.36 ;
      RECT 40.295 3.092 40.62 3.215 ;
      RECT 40.305 3.087 40.62 3.36 ;
      RECT 40.325 3.077 40.61 3.386 ;
      RECT 39.91 4.402 40.08 4.69 ;
      RECT 39.905 4.42 40.09 4.685 ;
      RECT 39.87 4.428 40.155 4.605 ;
      RECT 39.87 4.428 40.241 4.595 ;
      RECT 39.87 4.428 40.295 4.541 ;
      RECT 40.155 4.325 40.325 4.509 ;
      RECT 39.87 4.48 40.33 4.497 ;
      RECT 39.855 4.45 40.325 4.493 ;
      RECT 40.115 4.332 40.155 4.644 ;
      RECT 39.995 4.369 40.325 4.509 ;
      RECT 40.09 4.344 40.115 4.67 ;
      RECT 40.08 4.351 40.325 4.509 ;
      RECT 40.211 3.815 40.28 4.074 ;
      RECT 40.211 3.87 40.285 4.073 ;
      RECT 40.125 3.87 40.285 4.072 ;
      RECT 40.12 3.87 40.29 4.065 ;
      RECT 40.11 3.815 40.28 4.06 ;
      RECT 39.79 10.05 39.965 10.6 ;
      RECT 39.79 7.31 39.96 10.6 ;
      RECT 39.79 7.31 39.965 8.45 ;
      RECT 39.49 3.114 39.665 3.415 ;
      RECT 39.475 3.102 39.49 3.4 ;
      RECT 39.445 3.101 39.475 3.353 ;
      RECT 39.445 3.119 39.67 3.348 ;
      RECT 39.43 3.103 39.49 3.313 ;
      RECT 39.425 3.125 39.68 3.213 ;
      RECT 39.425 3.108 39.576 3.213 ;
      RECT 39.425 3.11 39.58 3.213 ;
      RECT 39.43 3.106 39.576 3.313 ;
      RECT 39.535 4.342 39.54 4.69 ;
      RECT 39.525 4.332 39.535 4.696 ;
      RECT 39.49 4.322 39.525 4.698 ;
      RECT 39.452 4.317 39.49 4.702 ;
      RECT 39.366 4.31 39.452 4.709 ;
      RECT 39.28 4.3 39.366 4.719 ;
      RECT 39.235 4.295 39.28 4.727 ;
      RECT 39.231 4.295 39.235 4.731 ;
      RECT 39.145 4.295 39.231 4.738 ;
      RECT 39.13 4.295 39.145 4.738 ;
      RECT 39.12 4.293 39.13 4.71 ;
      RECT 39.11 4.289 39.12 4.653 ;
      RECT 39.09 4.283 39.11 4.585 ;
      RECT 39.085 4.279 39.09 4.533 ;
      RECT 39.075 4.278 39.085 4.5 ;
      RECT 39.025 4.276 39.075 4.485 ;
      RECT 39 4.274 39.025 4.48 ;
      RECT 38.957 4.272 39 4.476 ;
      RECT 38.871 4.268 38.957 4.464 ;
      RECT 38.785 4.263 38.871 4.448 ;
      RECT 38.755 4.26 38.785 4.435 ;
      RECT 38.73 4.259 38.755 4.423 ;
      RECT 38.725 4.259 38.73 4.413 ;
      RECT 38.685 4.258 38.725 4.405 ;
      RECT 38.67 4.257 38.685 4.398 ;
      RECT 38.62 4.256 38.67 4.39 ;
      RECT 38.618 4.255 38.62 4.385 ;
      RECT 38.532 4.253 38.618 4.385 ;
      RECT 38.446 4.248 38.532 4.385 ;
      RECT 38.36 4.244 38.446 4.385 ;
      RECT 38.311 4.24 38.36 4.383 ;
      RECT 38.225 4.237 38.311 4.378 ;
      RECT 38.202 4.234 38.225 4.374 ;
      RECT 38.116 4.231 38.202 4.369 ;
      RECT 38.03 4.227 38.116 4.36 ;
      RECT 38.005 4.22 38.03 4.355 ;
      RECT 37.945 4.185 38.005 4.352 ;
      RECT 37.925 4.11 37.945 4.349 ;
      RECT 37.92 4.052 37.925 4.348 ;
      RECT 37.895 3.992 37.92 4.347 ;
      RECT 37.82 3.87 37.895 4.343 ;
      RECT 37.81 3.87 37.82 4.335 ;
      RECT 37.795 3.87 37.81 4.325 ;
      RECT 37.78 3.87 37.795 4.295 ;
      RECT 37.765 3.87 37.78 4.24 ;
      RECT 37.75 3.87 37.765 4.178 ;
      RECT 37.725 3.87 37.75 4.103 ;
      RECT 37.72 3.87 37.725 4.053 ;
      RECT 39.36 7.31 39.53 9.52 ;
      RECT 39.36 7.31 39.535 8.57 ;
      RECT 39.065 3.415 39.085 3.724 ;
      RECT 39.051 3.417 39.1 3.721 ;
      RECT 39.051 3.422 39.12 3.712 ;
      RECT 38.965 3.42 39.1 3.706 ;
      RECT 38.965 3.428 39.155 3.689 ;
      RECT 38.93 3.43 39.155 3.688 ;
      RECT 38.9 3.438 39.155 3.679 ;
      RECT 38.89 3.443 39.175 3.665 ;
      RECT 38.93 3.433 39.175 3.665 ;
      RECT 38.93 3.436 39.185 3.653 ;
      RECT 38.9 3.438 39.195 3.64 ;
      RECT 38.9 3.442 39.205 3.583 ;
      RECT 38.89 3.447 39.21 3.498 ;
      RECT 39.051 3.415 39.085 3.721 ;
      RECT 38.49 3.518 38.495 3.73 ;
      RECT 38.365 3.515 38.38 3.73 ;
      RECT 37.83 3.545 37.9 3.73 ;
      RECT 37.715 3.545 37.75 3.725 ;
      RECT 38.836 3.847 38.855 4.041 ;
      RECT 38.75 3.802 38.836 4.042 ;
      RECT 38.74 3.755 38.75 4.044 ;
      RECT 38.735 3.735 38.74 4.045 ;
      RECT 38.715 3.7 38.735 4.046 ;
      RECT 38.7 3.65 38.715 4.047 ;
      RECT 38.68 3.587 38.7 4.048 ;
      RECT 38.67 3.55 38.68 4.049 ;
      RECT 38.655 3.539 38.67 4.05 ;
      RECT 38.65 3.531 38.655 4.048 ;
      RECT 38.64 3.53 38.65 4.04 ;
      RECT 38.61 3.527 38.64 4.019 ;
      RECT 38.535 3.522 38.61 3.964 ;
      RECT 38.52 3.518 38.535 3.91 ;
      RECT 38.51 3.518 38.52 3.805 ;
      RECT 38.495 3.518 38.51 3.738 ;
      RECT 38.48 3.518 38.49 3.728 ;
      RECT 38.425 3.517 38.48 3.725 ;
      RECT 38.38 3.515 38.425 3.728 ;
      RECT 38.352 3.515 38.365 3.731 ;
      RECT 38.266 3.519 38.352 3.733 ;
      RECT 38.18 3.525 38.266 3.738 ;
      RECT 38.16 3.529 38.18 3.74 ;
      RECT 38.158 3.53 38.16 3.739 ;
      RECT 38.072 3.532 38.158 3.738 ;
      RECT 37.986 3.537 38.072 3.735 ;
      RECT 37.9 3.542 37.986 3.732 ;
      RECT 37.75 3.545 37.83 3.728 ;
      RECT 38.405 10.11 38.58 10.6 ;
      RECT 38.405 7.31 38.575 10.6 ;
      RECT 38.405 9.61 38.815 9.94 ;
      RECT 38.405 8.77 38.815 9.1 ;
      RECT 38.405 7.31 38.58 8.57 ;
      RECT 38.526 4.52 38.575 4.854 ;
      RECT 38.526 4.52 38.58 4.853 ;
      RECT 38.44 4.52 38.58 4.852 ;
      RECT 38.215 4.628 38.585 4.85 ;
      RECT 38.44 4.52 38.61 4.843 ;
      RECT 38.41 4.532 38.615 4.834 ;
      RECT 38.395 4.55 38.62 4.831 ;
      RECT 38.21 4.634 38.62 4.758 ;
      RECT 38.205 4.641 38.62 4.718 ;
      RECT 38.22 4.607 38.62 4.831 ;
      RECT 38.381 4.553 38.585 4.85 ;
      RECT 38.295 4.573 38.62 4.831 ;
      RECT 38.395 4.547 38.615 4.834 ;
      RECT 38.165 3.871 38.355 4.065 ;
      RECT 38.16 3.873 38.355 4.064 ;
      RECT 38.155 3.877 38.37 4.061 ;
      RECT 38.17 3.87 38.37 4.061 ;
      RECT 38.155 3.98 38.375 4.056 ;
      RECT 37.45 4.48 37.541 4.778 ;
      RECT 37.445 4.482 37.62 4.773 ;
      RECT 37.45 4.48 37.62 4.773 ;
      RECT 37.445 4.486 37.64 4.771 ;
      RECT 37.445 4.541 37.68 4.77 ;
      RECT 37.445 4.576 37.695 4.764 ;
      RECT 37.445 4.61 37.705 4.754 ;
      RECT 37.435 4.49 37.64 4.605 ;
      RECT 37.435 4.51 37.655 4.605 ;
      RECT 37.435 4.493 37.645 4.605 ;
      RECT 37.66 3.261 37.665 3.323 ;
      RECT 37.655 3.183 37.66 3.346 ;
      RECT 37.65 3.14 37.655 3.357 ;
      RECT 37.645 3.13 37.65 3.369 ;
      RECT 37.64 3.13 37.645 3.378 ;
      RECT 37.615 3.13 37.64 3.41 ;
      RECT 37.61 3.13 37.615 3.443 ;
      RECT 37.595 3.13 37.61 3.468 ;
      RECT 37.585 3.13 37.595 3.495 ;
      RECT 37.58 3.13 37.585 3.508 ;
      RECT 37.575 3.13 37.58 3.523 ;
      RECT 37.565 3.13 37.575 3.538 ;
      RECT 37.56 3.13 37.565 3.558 ;
      RECT 37.535 3.13 37.56 3.593 ;
      RECT 37.49 3.13 37.535 3.638 ;
      RECT 37.48 3.13 37.49 3.651 ;
      RECT 37.395 3.215 37.48 3.658 ;
      RECT 37.36 3.337 37.395 3.667 ;
      RECT 37.355 3.377 37.36 3.671 ;
      RECT 37.335 3.4 37.355 3.673 ;
      RECT 37.33 3.43 37.335 3.676 ;
      RECT 37.32 3.442 37.33 3.677 ;
      RECT 37.275 3.465 37.32 3.682 ;
      RECT 37.235 3.495 37.275 3.69 ;
      RECT 37.2 3.507 37.235 3.696 ;
      RECT 37.195 3.512 37.2 3.7 ;
      RECT 37.125 3.522 37.195 3.707 ;
      RECT 37.085 3.532 37.125 3.717 ;
      RECT 37.065 3.537 37.085 3.723 ;
      RECT 37.055 3.541 37.065 3.728 ;
      RECT 37.05 3.544 37.055 3.731 ;
      RECT 37.04 3.545 37.05 3.732 ;
      RECT 37.015 3.547 37.04 3.736 ;
      RECT 37.005 3.552 37.015 3.739 ;
      RECT 36.96 3.56 37.005 3.74 ;
      RECT 36.835 3.565 36.96 3.74 ;
      RECT 37.39 3.862 37.41 4.044 ;
      RECT 37.341 3.847 37.39 4.043 ;
      RECT 37.255 3.862 37.41 4.041 ;
      RECT 37.24 3.862 37.41 4.04 ;
      RECT 37.205 3.84 37.375 4.025 ;
      RECT 37.275 4.86 37.29 5.069 ;
      RECT 37.275 4.868 37.295 5.068 ;
      RECT 37.22 4.868 37.295 5.067 ;
      RECT 37.2 4.872 37.3 5.065 ;
      RECT 37.18 4.822 37.22 5.064 ;
      RECT 37.125 4.88 37.305 5.062 ;
      RECT 37.09 4.837 37.22 5.06 ;
      RECT 37.086 4.84 37.275 5.059 ;
      RECT 37 4.848 37.275 5.057 ;
      RECT 37 4.892 37.31 5.05 ;
      RECT 36.99 4.985 37.31 5.048 ;
      RECT 37 4.904 37.315 5.033 ;
      RECT 37 4.925 37.33 5.003 ;
      RECT 37 4.952 37.335 4.973 ;
      RECT 37.125 4.83 37.22 5.062 ;
      RECT 36.755 3.875 36.76 4.413 ;
      RECT 36.56 4.205 36.565 4.4 ;
      RECT 34.86 3.87 34.875 4.25 ;
      RECT 36.925 3.87 36.93 4.04 ;
      RECT 36.92 3.87 36.925 4.05 ;
      RECT 36.915 3.87 36.92 4.063 ;
      RECT 36.89 3.87 36.915 4.105 ;
      RECT 36.865 3.87 36.89 4.178 ;
      RECT 36.85 3.87 36.865 4.23 ;
      RECT 36.845 3.87 36.85 4.26 ;
      RECT 36.82 3.87 36.845 4.3 ;
      RECT 36.805 3.87 36.82 4.355 ;
      RECT 36.8 3.87 36.805 4.388 ;
      RECT 36.775 3.87 36.8 4.408 ;
      RECT 36.76 3.87 36.775 4.414 ;
      RECT 36.69 3.905 36.755 4.41 ;
      RECT 36.64 3.96 36.69 4.405 ;
      RECT 36.63 3.992 36.64 4.403 ;
      RECT 36.625 4.017 36.63 4.403 ;
      RECT 36.605 4.09 36.625 4.403 ;
      RECT 36.595 4.17 36.605 4.402 ;
      RECT 36.58 4.2 36.595 4.402 ;
      RECT 36.565 4.205 36.58 4.401 ;
      RECT 36.505 4.207 36.56 4.398 ;
      RECT 36.475 4.212 36.505 4.394 ;
      RECT 36.473 4.215 36.475 4.393 ;
      RECT 36.387 4.217 36.473 4.39 ;
      RECT 36.301 4.223 36.387 4.384 ;
      RECT 36.215 4.228 36.301 4.378 ;
      RECT 36.142 4.233 36.215 4.379 ;
      RECT 36.056 4.239 36.142 4.387 ;
      RECT 35.97 4.245 36.056 4.396 ;
      RECT 35.95 4.249 35.97 4.401 ;
      RECT 35.903 4.251 35.95 4.404 ;
      RECT 35.817 4.256 35.903 4.41 ;
      RECT 35.731 4.261 35.817 4.419 ;
      RECT 35.645 4.267 35.731 4.427 ;
      RECT 35.56 4.265 35.645 4.436 ;
      RECT 35.556 4.26 35.56 4.44 ;
      RECT 35.47 4.255 35.556 4.432 ;
      RECT 35.406 4.246 35.47 4.42 ;
      RECT 35.32 4.237 35.406 4.407 ;
      RECT 35.296 4.23 35.32 4.398 ;
      RECT 35.21 4.224 35.296 4.385 ;
      RECT 35.17 4.217 35.21 4.371 ;
      RECT 35.165 4.207 35.17 4.367 ;
      RECT 35.155 4.195 35.165 4.366 ;
      RECT 35.135 4.165 35.155 4.363 ;
      RECT 35.08 4.085 35.135 4.357 ;
      RECT 35.06 4.004 35.08 4.352 ;
      RECT 35.04 3.962 35.06 4.348 ;
      RECT 35.015 3.915 35.04 4.342 ;
      RECT 35.01 3.89 35.015 4.339 ;
      RECT 34.975 3.87 35.01 4.334 ;
      RECT 34.966 3.87 34.975 4.327 ;
      RECT 34.88 3.87 34.966 4.297 ;
      RECT 34.875 3.87 34.88 4.26 ;
      RECT 34.84 3.87 34.86 4.182 ;
      RECT 34.835 3.912 34.84 4.147 ;
      RECT 34.83 3.987 34.835 4.103 ;
      RECT 36.28 3.792 36.455 4.04 ;
      RECT 36.28 3.792 36.46 4.038 ;
      RECT 36.275 3.824 36.46 3.998 ;
      RECT 36.305 3.765 36.475 3.985 ;
      RECT 36.27 3.842 36.475 3.918 ;
      RECT 35.58 3.305 35.75 3.48 ;
      RECT 35.58 3.305 35.922 3.472 ;
      RECT 35.58 3.305 36.005 3.466 ;
      RECT 35.58 3.305 36.04 3.462 ;
      RECT 35.58 3.305 36.06 3.461 ;
      RECT 35.58 3.305 36.146 3.457 ;
      RECT 36.04 3.13 36.21 3.452 ;
      RECT 35.615 3.237 36.24 3.45 ;
      RECT 35.605 3.292 36.245 3.448 ;
      RECT 35.58 3.328 36.255 3.443 ;
      RECT 35.58 3.355 36.26 3.373 ;
      RECT 35.645 3.18 36.22 3.45 ;
      RECT 35.836 3.165 36.22 3.45 ;
      RECT 35.67 3.168 36.22 3.45 ;
      RECT 35.75 3.166 35.836 3.477 ;
      RECT 35.836 3.163 36.215 3.45 ;
      RECT 36.02 3.14 36.215 3.45 ;
      RECT 35.922 3.161 36.215 3.45 ;
      RECT 36.005 3.155 36.02 3.463 ;
      RECT 36.155 4.52 36.16 4.72 ;
      RECT 35.62 4.585 35.665 4.72 ;
      RECT 36.19 4.52 36.21 4.693 ;
      RECT 36.16 4.52 36.19 4.708 ;
      RECT 36.095 4.52 36.155 4.745 ;
      RECT 36.08 4.52 36.095 4.775 ;
      RECT 36.065 4.52 36.08 4.788 ;
      RECT 36.045 4.52 36.065 4.803 ;
      RECT 36.04 4.52 36.045 4.812 ;
      RECT 36.03 4.524 36.04 4.817 ;
      RECT 36.015 4.534 36.03 4.828 ;
      RECT 35.99 4.55 36.015 4.838 ;
      RECT 35.98 4.564 35.99 4.84 ;
      RECT 35.96 4.576 35.98 4.837 ;
      RECT 35.93 4.597 35.96 4.831 ;
      RECT 35.92 4.609 35.93 4.826 ;
      RECT 35.91 4.607 35.92 4.823 ;
      RECT 35.895 4.606 35.91 4.818 ;
      RECT 35.89 4.605 35.895 4.813 ;
      RECT 35.855 4.603 35.89 4.803 ;
      RECT 35.835 4.6 35.855 4.785 ;
      RECT 35.825 4.598 35.835 4.78 ;
      RECT 35.815 4.597 35.825 4.775 ;
      RECT 35.78 4.595 35.815 4.763 ;
      RECT 35.725 4.591 35.78 4.743 ;
      RECT 35.715 4.589 35.725 4.728 ;
      RECT 35.71 4.589 35.715 4.723 ;
      RECT 35.665 4.587 35.71 4.72 ;
      RECT 35.57 4.585 35.62 4.724 ;
      RECT 35.56 4.586 35.57 4.729 ;
      RECT 35.5 4.593 35.56 4.743 ;
      RECT 35.475 4.601 35.5 4.763 ;
      RECT 35.465 4.605 35.475 4.775 ;
      RECT 35.46 4.606 35.465 4.78 ;
      RECT 35.445 4.608 35.46 4.783 ;
      RECT 35.43 4.61 35.445 4.788 ;
      RECT 35.425 4.61 35.43 4.791 ;
      RECT 35.38 4.615 35.425 4.802 ;
      RECT 35.375 4.619 35.38 4.814 ;
      RECT 35.35 4.615 35.375 4.818 ;
      RECT 35.34 4.611 35.35 4.822 ;
      RECT 35.33 4.61 35.34 4.826 ;
      RECT 35.315 4.6 35.33 4.832 ;
      RECT 35.31 4.588 35.315 4.836 ;
      RECT 35.305 4.585 35.31 4.837 ;
      RECT 35.3 4.582 35.305 4.839 ;
      RECT 35.285 4.57 35.3 4.838 ;
      RECT 35.27 4.552 35.285 4.835 ;
      RECT 35.25 4.531 35.27 4.828 ;
      RECT 35.185 4.52 35.25 4.8 ;
      RECT 35.181 4.52 35.185 4.779 ;
      RECT 35.095 4.52 35.181 4.749 ;
      RECT 35.08 4.52 35.095 4.705 ;
      RECT 35.73 4.871 35.745 5.13 ;
      RECT 35.73 4.886 35.75 5.129 ;
      RECT 35.646 4.886 35.75 5.127 ;
      RECT 35.646 4.9 35.755 5.126 ;
      RECT 35.56 4.942 35.76 5.123 ;
      RECT 35.555 4.885 35.745 5.118 ;
      RECT 35.555 4.956 35.765 5.115 ;
      RECT 35.55 4.987 35.765 5.113 ;
      RECT 35.555 4.984 35.78 5.103 ;
      RECT 35.55 5.03 35.795 5.088 ;
      RECT 35.55 5.058 35.8 5.073 ;
      RECT 35.56 4.86 35.73 5.123 ;
      RECT 35.32 3.87 35.49 4.04 ;
      RECT 35.285 3.87 35.49 4.035 ;
      RECT 35.275 3.87 35.49 4.028 ;
      RECT 35.27 3.855 35.44 4.025 ;
      RECT 34.1 4.392 34.365 4.835 ;
      RECT 34.095 4.363 34.31 4.833 ;
      RECT 34.09 4.517 34.37 4.828 ;
      RECT 34.095 4.412 34.37 4.828 ;
      RECT 34.095 4.423 34.38 4.815 ;
      RECT 34.095 4.37 34.34 4.833 ;
      RECT 34.1 4.357 34.31 4.835 ;
      RECT 34.1 4.355 34.26 4.835 ;
      RECT 34.201 4.347 34.26 4.835 ;
      RECT 34.115 4.348 34.26 4.835 ;
      RECT 34.201 4.346 34.25 4.835 ;
      RECT 34.005 3.161 34.18 3.46 ;
      RECT 34.055 3.123 34.18 3.46 ;
      RECT 34.04 3.125 34.266 3.452 ;
      RECT 34.04 3.128 34.305 3.439 ;
      RECT 34.04 3.129 34.315 3.425 ;
      RECT 33.995 3.18 34.315 3.415 ;
      RECT 34.04 3.13 34.32 3.41 ;
      RECT 33.995 3.34 34.325 3.4 ;
      RECT 33.98 3.2 34.32 3.34 ;
      RECT 33.975 3.216 34.32 3.28 ;
      RECT 34.02 3.14 34.32 3.41 ;
      RECT 34.055 3.121 34.141 3.46 ;
      RECT 32.515 7.31 32.685 8.78 ;
      RECT 32.515 7.31 32.69 8.57 ;
      RECT 32.145 9.26 32.615 9.43 ;
      RECT 32.145 8.24 32.315 9.43 ;
      RECT 32.14 3.035 32.31 4.225 ;
      RECT 32.14 3.035 32.61 3.205 ;
      RECT 31.525 3.895 31.7 5.155 ;
      RECT 31.525 3.685 31.695 5.155 ;
      RECT 31.525 7.31 31.695 8.78 ;
      RECT 31.525 7.31 31.7 8.57 ;
      RECT 31.155 3.035 31.325 4.225 ;
      RECT 31.155 3.035 31.625 3.205 ;
      RECT 31.155 9.26 31.625 9.43 ;
      RECT 31.155 8.24 31.325 9.43 ;
      RECT 30.165 4.015 30.34 5.155 ;
      RECT 30.165 1.865 30.335 5.155 ;
      RECT 30.165 1.865 30.34 2.415 ;
      RECT 30.165 10.05 30.34 10.6 ;
      RECT 30.165 7.31 30.335 10.6 ;
      RECT 30.165 7.31 30.34 8.45 ;
      RECT 29.735 3.895 29.91 5.155 ;
      RECT 29.735 2.945 29.905 5.155 ;
      RECT 29.735 7.31 29.905 9.52 ;
      RECT 29.735 7.31 29.91 8.57 ;
      RECT 29.305 3.925 29.475 5.155 ;
      RECT 29.365 2.145 29.535 4.095 ;
      RECT 29.305 1.865 29.475 2.315 ;
      RECT 29.305 10.15 29.475 10.6 ;
      RECT 29.365 8.37 29.535 10.32 ;
      RECT 29.305 7.31 29.475 8.54 ;
      RECT 28.78 3.895 28.955 5.155 ;
      RECT 28.78 1.865 28.95 5.155 ;
      RECT 28.78 3.365 29.19 3.695 ;
      RECT 28.78 2.525 29.19 2.855 ;
      RECT 28.78 1.865 28.955 2.355 ;
      RECT 28.78 10.11 28.955 10.6 ;
      RECT 28.78 7.31 28.95 10.6 ;
      RECT 28.78 9.61 29.19 9.94 ;
      RECT 28.78 8.77 29.19 9.1 ;
      RECT 28.78 7.31 28.955 8.57 ;
      RECT 26.71 4.421 26.715 4.593 ;
      RECT 26.705 4.414 26.71 4.683 ;
      RECT 26.7 4.408 26.705 4.702 ;
      RECT 26.68 4.402 26.7 4.712 ;
      RECT 26.665 4.397 26.68 4.72 ;
      RECT 26.628 4.391 26.665 4.718 ;
      RECT 26.542 4.377 26.628 4.714 ;
      RECT 26.456 4.359 26.542 4.709 ;
      RECT 26.37 4.34 26.456 4.703 ;
      RECT 26.34 4.328 26.37 4.699 ;
      RECT 26.32 4.322 26.34 4.698 ;
      RECT 26.255 4.32 26.32 4.696 ;
      RECT 26.24 4.32 26.255 4.688 ;
      RECT 26.225 4.32 26.24 4.675 ;
      RECT 26.22 4.32 26.225 4.665 ;
      RECT 26.205 4.32 26.22 4.643 ;
      RECT 26.19 4.32 26.205 4.61 ;
      RECT 26.185 4.32 26.19 4.588 ;
      RECT 26.175 4.32 26.185 4.57 ;
      RECT 26.16 4.32 26.175 4.548 ;
      RECT 26.14 4.32 26.16 4.51 ;
      RECT 26.49 3.605 26.525 4.044 ;
      RECT 26.49 3.605 26.53 4.043 ;
      RECT 26.435 3.665 26.53 4.042 ;
      RECT 26.3 3.837 26.53 4.041 ;
      RECT 26.41 3.715 26.53 4.041 ;
      RECT 26.3 3.837 26.555 4.031 ;
      RECT 26.355 3.782 26.635 3.948 ;
      RECT 26.53 3.576 26.535 4.039 ;
      RECT 26.385 3.752 26.675 3.825 ;
      RECT 26.4 3.735 26.53 4.041 ;
      RECT 26.535 3.575 26.705 3.763 ;
      RECT 26.525 3.578 26.705 3.763 ;
      RECT 26.03 3.455 26.2 3.765 ;
      RECT 26.03 3.455 26.205 3.738 ;
      RECT 26.03 3.455 26.21 3.715 ;
      RECT 26.03 3.455 26.22 3.665 ;
      RECT 26.025 3.56 26.22 3.635 ;
      RECT 26.06 3.13 26.23 3.608 ;
      RECT 26.06 3.13 26.245 3.529 ;
      RECT 26.05 3.34 26.245 3.529 ;
      RECT 26.06 3.14 26.255 3.444 ;
      RECT 25.99 3.882 25.995 4.085 ;
      RECT 25.98 3.87 25.99 4.195 ;
      RECT 25.955 3.87 25.98 4.235 ;
      RECT 25.875 3.87 25.955 4.32 ;
      RECT 25.865 3.87 25.875 4.39 ;
      RECT 25.84 3.87 25.865 4.413 ;
      RECT 25.82 3.87 25.84 4.448 ;
      RECT 25.775 3.88 25.82 4.491 ;
      RECT 25.765 3.892 25.775 4.528 ;
      RECT 25.745 3.906 25.765 4.548 ;
      RECT 25.735 3.924 25.745 4.564 ;
      RECT 25.72 3.95 25.735 4.574 ;
      RECT 25.705 3.991 25.72 4.588 ;
      RECT 25.695 4.026 25.705 4.598 ;
      RECT 25.69 4.042 25.695 4.603 ;
      RECT 25.68 4.057 25.69 4.608 ;
      RECT 25.66 4.1 25.68 4.618 ;
      RECT 25.64 4.137 25.66 4.631 ;
      RECT 25.605 4.16 25.64 4.649 ;
      RECT 25.595 4.174 25.605 4.665 ;
      RECT 25.575 4.184 25.595 4.675 ;
      RECT 25.57 4.193 25.575 4.683 ;
      RECT 25.56 4.2 25.57 4.69 ;
      RECT 25.55 4.207 25.56 4.698 ;
      RECT 25.535 4.217 25.55 4.706 ;
      RECT 25.525 4.231 25.535 4.716 ;
      RECT 25.515 4.243 25.525 4.728 ;
      RECT 25.5 4.265 25.515 4.741 ;
      RECT 25.49 4.287 25.5 4.752 ;
      RECT 25.48 4.307 25.49 4.761 ;
      RECT 25.475 4.322 25.48 4.768 ;
      RECT 25.445 4.355 25.475 4.782 ;
      RECT 25.435 4.39 25.445 4.797 ;
      RECT 25.43 4.397 25.435 4.803 ;
      RECT 25.41 4.412 25.43 4.81 ;
      RECT 25.405 4.427 25.41 4.818 ;
      RECT 25.4 4.436 25.405 4.823 ;
      RECT 25.385 4.442 25.4 4.83 ;
      RECT 25.38 4.448 25.385 4.838 ;
      RECT 25.375 4.452 25.38 4.845 ;
      RECT 25.37 4.456 25.375 4.855 ;
      RECT 25.36 4.461 25.37 4.865 ;
      RECT 25.34 4.472 25.36 4.893 ;
      RECT 25.325 4.484 25.34 4.92 ;
      RECT 25.305 4.497 25.325 4.945 ;
      RECT 25.285 4.512 25.305 4.969 ;
      RECT 25.27 4.527 25.285 4.984 ;
      RECT 25.265 4.538 25.27 4.993 ;
      RECT 25.2 4.583 25.265 5.003 ;
      RECT 25.165 4.642 25.2 5.016 ;
      RECT 25.16 4.665 25.165 5.022 ;
      RECT 25.155 4.672 25.16 5.024 ;
      RECT 25.14 4.682 25.155 5.027 ;
      RECT 25.11 4.707 25.14 5.031 ;
      RECT 25.105 4.725 25.11 5.035 ;
      RECT 25.1 4.732 25.105 5.036 ;
      RECT 25.08 4.74 25.1 5.04 ;
      RECT 25.07 4.747 25.08 5.044 ;
      RECT 25.026 4.758 25.07 5.051 ;
      RECT 24.94 4.786 25.026 5.067 ;
      RECT 24.88 4.81 24.94 5.085 ;
      RECT 24.835 4.82 24.88 5.099 ;
      RECT 24.776 4.828 24.835 5.113 ;
      RECT 24.69 4.835 24.776 5.132 ;
      RECT 24.665 4.84 24.69 5.147 ;
      RECT 24.585 4.843 24.665 5.15 ;
      RECT 24.505 4.847 24.585 5.137 ;
      RECT 24.496 4.85 24.505 5.122 ;
      RECT 24.41 4.85 24.496 5.107 ;
      RECT 24.35 4.852 24.41 5.084 ;
      RECT 24.346 4.855 24.35 5.074 ;
      RECT 24.26 4.855 24.346 5.059 ;
      RECT 24.185 4.855 24.26 5.035 ;
      RECT 25.5 3.864 25.51 4.04 ;
      RECT 25.455 3.831 25.5 4.04 ;
      RECT 25.41 3.782 25.455 4.04 ;
      RECT 25.38 3.752 25.41 4.041 ;
      RECT 25.375 3.735 25.38 4.042 ;
      RECT 25.35 3.715 25.375 4.043 ;
      RECT 25.335 3.69 25.35 4.044 ;
      RECT 25.33 3.677 25.335 4.045 ;
      RECT 25.325 3.671 25.33 4.043 ;
      RECT 25.32 3.663 25.325 4.037 ;
      RECT 25.295 3.655 25.32 4.017 ;
      RECT 25.275 3.644 25.295 3.988 ;
      RECT 25.245 3.629 25.275 3.959 ;
      RECT 25.225 3.615 25.245 3.931 ;
      RECT 25.215 3.609 25.225 3.91 ;
      RECT 25.21 3.606 25.215 3.893 ;
      RECT 25.205 3.603 25.21 3.878 ;
      RECT 25.19 3.598 25.205 3.843 ;
      RECT 25.185 3.594 25.19 3.81 ;
      RECT 25.165 3.589 25.185 3.786 ;
      RECT 25.135 3.581 25.165 3.751 ;
      RECT 25.12 3.575 25.135 3.728 ;
      RECT 25.08 3.568 25.12 3.713 ;
      RECT 25.055 3.56 25.08 3.693 ;
      RECT 25.035 3.555 25.055 3.683 ;
      RECT 25 3.549 25.035 3.678 ;
      RECT 24.955 3.54 25 3.677 ;
      RECT 24.925 3.536 24.955 3.679 ;
      RECT 24.84 3.544 24.925 3.683 ;
      RECT 24.77 3.555 24.84 3.705 ;
      RECT 24.757 3.561 24.77 3.728 ;
      RECT 24.671 3.568 24.757 3.75 ;
      RECT 24.585 3.58 24.671 3.787 ;
      RECT 24.585 3.957 24.595 4.195 ;
      RECT 24.58 3.586 24.585 3.81 ;
      RECT 24.575 3.842 24.585 4.195 ;
      RECT 24.575 3.587 24.58 3.815 ;
      RECT 24.57 3.588 24.575 4.195 ;
      RECT 24.546 3.59 24.57 4.196 ;
      RECT 24.46 3.598 24.546 4.198 ;
      RECT 24.44 3.612 24.46 4.201 ;
      RECT 24.435 3.64 24.44 4.202 ;
      RECT 24.43 3.652 24.435 4.203 ;
      RECT 24.425 3.667 24.43 4.204 ;
      RECT 24.415 3.697 24.425 4.205 ;
      RECT 24.41 3.735 24.415 4.203 ;
      RECT 24.405 3.755 24.41 4.198 ;
      RECT 24.39 3.79 24.405 4.183 ;
      RECT 24.38 3.842 24.39 4.163 ;
      RECT 24.375 3.872 24.38 4.151 ;
      RECT 24.36 3.885 24.375 4.134 ;
      RECT 24.335 3.889 24.36 4.101 ;
      RECT 24.32 3.887 24.335 4.078 ;
      RECT 24.305 3.886 24.32 4.075 ;
      RECT 24.245 3.884 24.305 4.073 ;
      RECT 24.235 3.882 24.245 4.068 ;
      RECT 24.195 3.881 24.235 4.065 ;
      RECT 24.125 3.878 24.195 4.063 ;
      RECT 24.07 3.876 24.125 4.058 ;
      RECT 24 3.87 24.07 4.053 ;
      RECT 23.991 3.87 24 4.05 ;
      RECT 23.905 3.87 23.991 4.045 ;
      RECT 23.9 3.87 23.905 4.04 ;
      RECT 25.205 3.105 25.38 3.455 ;
      RECT 25.205 3.12 25.39 3.453 ;
      RECT 25.18 3.07 25.325 3.45 ;
      RECT 25.16 3.071 25.325 3.443 ;
      RECT 25.15 3.072 25.335 3.438 ;
      RECT 25.12 3.073 25.335 3.425 ;
      RECT 25.07 3.074 25.335 3.401 ;
      RECT 25.065 3.076 25.335 3.386 ;
      RECT 25.065 3.142 25.395 3.38 ;
      RECT 25.045 3.083 25.35 3.36 ;
      RECT 25.035 3.092 25.36 3.215 ;
      RECT 25.045 3.087 25.36 3.36 ;
      RECT 25.065 3.077 25.35 3.386 ;
      RECT 24.65 4.402 24.82 4.69 ;
      RECT 24.645 4.42 24.83 4.685 ;
      RECT 24.61 4.428 24.895 4.605 ;
      RECT 24.61 4.428 24.981 4.595 ;
      RECT 24.61 4.428 25.035 4.541 ;
      RECT 24.895 4.325 25.065 4.509 ;
      RECT 24.61 4.48 25.07 4.497 ;
      RECT 24.595 4.45 25.065 4.493 ;
      RECT 24.855 4.332 24.895 4.644 ;
      RECT 24.735 4.369 25.065 4.509 ;
      RECT 24.83 4.344 24.855 4.67 ;
      RECT 24.82 4.351 25.065 4.509 ;
      RECT 24.951 3.815 25.02 4.074 ;
      RECT 24.951 3.87 25.025 4.073 ;
      RECT 24.865 3.87 25.025 4.072 ;
      RECT 24.86 3.87 25.03 4.065 ;
      RECT 24.85 3.815 25.02 4.06 ;
      RECT 24.53 10.05 24.705 10.6 ;
      RECT 24.53 7.31 24.7 10.6 ;
      RECT 24.53 7.31 24.705 8.45 ;
      RECT 24.23 3.114 24.405 3.415 ;
      RECT 24.215 3.102 24.23 3.4 ;
      RECT 24.185 3.101 24.215 3.353 ;
      RECT 24.185 3.119 24.41 3.348 ;
      RECT 24.17 3.103 24.23 3.313 ;
      RECT 24.165 3.125 24.42 3.213 ;
      RECT 24.165 3.108 24.316 3.213 ;
      RECT 24.165 3.11 24.32 3.213 ;
      RECT 24.17 3.106 24.316 3.313 ;
      RECT 24.275 4.342 24.28 4.69 ;
      RECT 24.265 4.332 24.275 4.696 ;
      RECT 24.23 4.322 24.265 4.698 ;
      RECT 24.192 4.317 24.23 4.702 ;
      RECT 24.106 4.31 24.192 4.709 ;
      RECT 24.02 4.3 24.106 4.719 ;
      RECT 23.975 4.295 24.02 4.727 ;
      RECT 23.971 4.295 23.975 4.731 ;
      RECT 23.885 4.295 23.971 4.738 ;
      RECT 23.87 4.295 23.885 4.738 ;
      RECT 23.86 4.293 23.87 4.71 ;
      RECT 23.85 4.289 23.86 4.653 ;
      RECT 23.83 4.283 23.85 4.585 ;
      RECT 23.825 4.279 23.83 4.533 ;
      RECT 23.815 4.278 23.825 4.5 ;
      RECT 23.765 4.276 23.815 4.485 ;
      RECT 23.74 4.274 23.765 4.48 ;
      RECT 23.697 4.272 23.74 4.476 ;
      RECT 23.611 4.268 23.697 4.464 ;
      RECT 23.525 4.263 23.611 4.448 ;
      RECT 23.495 4.26 23.525 4.435 ;
      RECT 23.47 4.259 23.495 4.423 ;
      RECT 23.465 4.259 23.47 4.413 ;
      RECT 23.425 4.258 23.465 4.405 ;
      RECT 23.41 4.257 23.425 4.398 ;
      RECT 23.36 4.256 23.41 4.39 ;
      RECT 23.358 4.255 23.36 4.385 ;
      RECT 23.272 4.253 23.358 4.385 ;
      RECT 23.186 4.248 23.272 4.385 ;
      RECT 23.1 4.244 23.186 4.385 ;
      RECT 23.051 4.24 23.1 4.383 ;
      RECT 22.965 4.237 23.051 4.378 ;
      RECT 22.942 4.234 22.965 4.374 ;
      RECT 22.856 4.231 22.942 4.369 ;
      RECT 22.77 4.227 22.856 4.36 ;
      RECT 22.745 4.22 22.77 4.355 ;
      RECT 22.685 4.185 22.745 4.352 ;
      RECT 22.665 4.11 22.685 4.349 ;
      RECT 22.66 4.052 22.665 4.348 ;
      RECT 22.635 3.992 22.66 4.347 ;
      RECT 22.56 3.87 22.635 4.343 ;
      RECT 22.55 3.87 22.56 4.335 ;
      RECT 22.535 3.87 22.55 4.325 ;
      RECT 22.52 3.87 22.535 4.295 ;
      RECT 22.505 3.87 22.52 4.24 ;
      RECT 22.49 3.87 22.505 4.178 ;
      RECT 22.465 3.87 22.49 4.103 ;
      RECT 22.46 3.87 22.465 4.053 ;
      RECT 24.1 7.31 24.27 9.52 ;
      RECT 24.1 7.31 24.275 8.57 ;
      RECT 23.805 3.415 23.825 3.724 ;
      RECT 23.791 3.417 23.84 3.721 ;
      RECT 23.791 3.422 23.86 3.712 ;
      RECT 23.705 3.42 23.84 3.706 ;
      RECT 23.705 3.428 23.895 3.689 ;
      RECT 23.67 3.43 23.895 3.688 ;
      RECT 23.64 3.438 23.895 3.679 ;
      RECT 23.63 3.443 23.915 3.665 ;
      RECT 23.67 3.433 23.915 3.665 ;
      RECT 23.67 3.436 23.925 3.653 ;
      RECT 23.64 3.438 23.935 3.64 ;
      RECT 23.64 3.442 23.945 3.583 ;
      RECT 23.63 3.447 23.95 3.498 ;
      RECT 23.791 3.415 23.825 3.721 ;
      RECT 23.23 3.518 23.235 3.73 ;
      RECT 23.105 3.515 23.12 3.73 ;
      RECT 22.57 3.545 22.64 3.73 ;
      RECT 22.455 3.545 22.49 3.725 ;
      RECT 23.576 3.847 23.595 4.041 ;
      RECT 23.49 3.802 23.576 4.042 ;
      RECT 23.48 3.755 23.49 4.044 ;
      RECT 23.475 3.735 23.48 4.045 ;
      RECT 23.455 3.7 23.475 4.046 ;
      RECT 23.44 3.65 23.455 4.047 ;
      RECT 23.42 3.587 23.44 4.048 ;
      RECT 23.41 3.55 23.42 4.049 ;
      RECT 23.395 3.539 23.41 4.05 ;
      RECT 23.39 3.531 23.395 4.048 ;
      RECT 23.38 3.53 23.39 4.04 ;
      RECT 23.35 3.527 23.38 4.019 ;
      RECT 23.275 3.522 23.35 3.964 ;
      RECT 23.26 3.518 23.275 3.91 ;
      RECT 23.25 3.518 23.26 3.805 ;
      RECT 23.235 3.518 23.25 3.738 ;
      RECT 23.22 3.518 23.23 3.728 ;
      RECT 23.165 3.517 23.22 3.725 ;
      RECT 23.12 3.515 23.165 3.728 ;
      RECT 23.092 3.515 23.105 3.731 ;
      RECT 23.006 3.519 23.092 3.733 ;
      RECT 22.92 3.525 23.006 3.738 ;
      RECT 22.9 3.529 22.92 3.74 ;
      RECT 22.898 3.53 22.9 3.739 ;
      RECT 22.812 3.532 22.898 3.738 ;
      RECT 22.726 3.537 22.812 3.735 ;
      RECT 22.64 3.542 22.726 3.732 ;
      RECT 22.49 3.545 22.57 3.728 ;
      RECT 23.145 10.11 23.32 10.6 ;
      RECT 23.145 7.31 23.315 10.6 ;
      RECT 23.145 9.61 23.555 9.94 ;
      RECT 23.145 8.77 23.555 9.1 ;
      RECT 23.145 7.31 23.32 8.57 ;
      RECT 23.266 4.52 23.315 4.854 ;
      RECT 23.266 4.52 23.32 4.853 ;
      RECT 23.18 4.52 23.32 4.852 ;
      RECT 22.955 4.628 23.325 4.85 ;
      RECT 23.18 4.52 23.35 4.843 ;
      RECT 23.15 4.532 23.355 4.834 ;
      RECT 23.135 4.55 23.36 4.831 ;
      RECT 22.95 4.634 23.36 4.758 ;
      RECT 22.945 4.641 23.36 4.718 ;
      RECT 22.96 4.607 23.36 4.831 ;
      RECT 23.121 4.553 23.325 4.85 ;
      RECT 23.035 4.573 23.36 4.831 ;
      RECT 23.135 4.547 23.355 4.834 ;
      RECT 22.905 3.871 23.095 4.065 ;
      RECT 22.9 3.873 23.095 4.064 ;
      RECT 22.895 3.877 23.11 4.061 ;
      RECT 22.91 3.87 23.11 4.061 ;
      RECT 22.895 3.98 23.115 4.056 ;
      RECT 22.19 4.48 22.281 4.778 ;
      RECT 22.185 4.482 22.36 4.773 ;
      RECT 22.19 4.48 22.36 4.773 ;
      RECT 22.185 4.486 22.38 4.771 ;
      RECT 22.185 4.541 22.42 4.77 ;
      RECT 22.185 4.576 22.435 4.764 ;
      RECT 22.185 4.61 22.445 4.754 ;
      RECT 22.175 4.49 22.38 4.605 ;
      RECT 22.175 4.51 22.395 4.605 ;
      RECT 22.175 4.493 22.385 4.605 ;
      RECT 22.4 3.261 22.405 3.323 ;
      RECT 22.395 3.183 22.4 3.346 ;
      RECT 22.39 3.14 22.395 3.357 ;
      RECT 22.385 3.13 22.39 3.369 ;
      RECT 22.38 3.13 22.385 3.378 ;
      RECT 22.355 3.13 22.38 3.41 ;
      RECT 22.35 3.13 22.355 3.443 ;
      RECT 22.335 3.13 22.35 3.468 ;
      RECT 22.325 3.13 22.335 3.495 ;
      RECT 22.32 3.13 22.325 3.508 ;
      RECT 22.315 3.13 22.32 3.523 ;
      RECT 22.305 3.13 22.315 3.538 ;
      RECT 22.3 3.13 22.305 3.558 ;
      RECT 22.275 3.13 22.3 3.593 ;
      RECT 22.23 3.13 22.275 3.638 ;
      RECT 22.22 3.13 22.23 3.651 ;
      RECT 22.135 3.215 22.22 3.658 ;
      RECT 22.1 3.337 22.135 3.667 ;
      RECT 22.095 3.377 22.1 3.671 ;
      RECT 22.075 3.4 22.095 3.673 ;
      RECT 22.07 3.43 22.075 3.676 ;
      RECT 22.06 3.442 22.07 3.677 ;
      RECT 22.015 3.465 22.06 3.682 ;
      RECT 21.975 3.495 22.015 3.69 ;
      RECT 21.94 3.507 21.975 3.696 ;
      RECT 21.935 3.512 21.94 3.7 ;
      RECT 21.865 3.522 21.935 3.707 ;
      RECT 21.825 3.532 21.865 3.717 ;
      RECT 21.805 3.537 21.825 3.723 ;
      RECT 21.795 3.541 21.805 3.728 ;
      RECT 21.79 3.544 21.795 3.731 ;
      RECT 21.78 3.545 21.79 3.732 ;
      RECT 21.755 3.547 21.78 3.736 ;
      RECT 21.745 3.552 21.755 3.739 ;
      RECT 21.7 3.56 21.745 3.74 ;
      RECT 21.575 3.565 21.7 3.74 ;
      RECT 22.13 3.862 22.15 4.044 ;
      RECT 22.081 3.847 22.13 4.043 ;
      RECT 21.995 3.862 22.15 4.041 ;
      RECT 21.98 3.862 22.15 4.04 ;
      RECT 21.945 3.84 22.115 4.025 ;
      RECT 22.015 4.86 22.03 5.069 ;
      RECT 22.015 4.868 22.035 5.068 ;
      RECT 21.96 4.868 22.035 5.067 ;
      RECT 21.94 4.872 22.04 5.065 ;
      RECT 21.92 4.822 21.96 5.064 ;
      RECT 21.865 4.88 22.045 5.062 ;
      RECT 21.83 4.837 21.96 5.06 ;
      RECT 21.826 4.84 22.015 5.059 ;
      RECT 21.74 4.848 22.015 5.057 ;
      RECT 21.74 4.892 22.05 5.05 ;
      RECT 21.73 4.985 22.05 5.048 ;
      RECT 21.74 4.904 22.055 5.033 ;
      RECT 21.74 4.925 22.07 5.003 ;
      RECT 21.74 4.952 22.075 4.973 ;
      RECT 21.865 4.83 21.96 5.062 ;
      RECT 21.495 3.875 21.5 4.413 ;
      RECT 21.3 4.205 21.305 4.4 ;
      RECT 19.6 3.87 19.615 4.25 ;
      RECT 21.665 3.87 21.67 4.04 ;
      RECT 21.66 3.87 21.665 4.05 ;
      RECT 21.655 3.87 21.66 4.063 ;
      RECT 21.63 3.87 21.655 4.105 ;
      RECT 21.605 3.87 21.63 4.178 ;
      RECT 21.59 3.87 21.605 4.23 ;
      RECT 21.585 3.87 21.59 4.26 ;
      RECT 21.56 3.87 21.585 4.3 ;
      RECT 21.545 3.87 21.56 4.355 ;
      RECT 21.54 3.87 21.545 4.388 ;
      RECT 21.515 3.87 21.54 4.408 ;
      RECT 21.5 3.87 21.515 4.414 ;
      RECT 21.43 3.905 21.495 4.41 ;
      RECT 21.38 3.96 21.43 4.405 ;
      RECT 21.37 3.992 21.38 4.403 ;
      RECT 21.365 4.017 21.37 4.403 ;
      RECT 21.345 4.09 21.365 4.403 ;
      RECT 21.335 4.17 21.345 4.402 ;
      RECT 21.32 4.2 21.335 4.402 ;
      RECT 21.305 4.205 21.32 4.401 ;
      RECT 21.245 4.207 21.3 4.398 ;
      RECT 21.215 4.212 21.245 4.394 ;
      RECT 21.213 4.215 21.215 4.393 ;
      RECT 21.127 4.217 21.213 4.39 ;
      RECT 21.041 4.223 21.127 4.384 ;
      RECT 20.955 4.228 21.041 4.378 ;
      RECT 20.882 4.233 20.955 4.379 ;
      RECT 20.796 4.239 20.882 4.387 ;
      RECT 20.71 4.245 20.796 4.396 ;
      RECT 20.69 4.249 20.71 4.401 ;
      RECT 20.643 4.251 20.69 4.404 ;
      RECT 20.557 4.256 20.643 4.41 ;
      RECT 20.471 4.261 20.557 4.419 ;
      RECT 20.385 4.267 20.471 4.427 ;
      RECT 20.3 4.265 20.385 4.436 ;
      RECT 20.296 4.26 20.3 4.44 ;
      RECT 20.21 4.255 20.296 4.432 ;
      RECT 20.146 4.246 20.21 4.42 ;
      RECT 20.06 4.237 20.146 4.407 ;
      RECT 20.036 4.23 20.06 4.398 ;
      RECT 19.95 4.224 20.036 4.385 ;
      RECT 19.91 4.217 19.95 4.371 ;
      RECT 19.905 4.207 19.91 4.367 ;
      RECT 19.895 4.195 19.905 4.366 ;
      RECT 19.875 4.165 19.895 4.363 ;
      RECT 19.82 4.085 19.875 4.357 ;
      RECT 19.8 4.004 19.82 4.352 ;
      RECT 19.78 3.962 19.8 4.348 ;
      RECT 19.755 3.915 19.78 4.342 ;
      RECT 19.75 3.89 19.755 4.339 ;
      RECT 19.715 3.87 19.75 4.334 ;
      RECT 19.706 3.87 19.715 4.327 ;
      RECT 19.62 3.87 19.706 4.297 ;
      RECT 19.615 3.87 19.62 4.26 ;
      RECT 19.58 3.87 19.6 4.182 ;
      RECT 19.575 3.912 19.58 4.147 ;
      RECT 19.57 3.987 19.575 4.103 ;
      RECT 21.02 3.792 21.195 4.04 ;
      RECT 21.02 3.792 21.2 4.038 ;
      RECT 21.015 3.824 21.2 3.998 ;
      RECT 21.045 3.765 21.215 3.985 ;
      RECT 21.01 3.842 21.215 3.918 ;
      RECT 20.32 3.305 20.49 3.48 ;
      RECT 20.32 3.305 20.662 3.472 ;
      RECT 20.32 3.305 20.745 3.466 ;
      RECT 20.32 3.305 20.78 3.462 ;
      RECT 20.32 3.305 20.8 3.461 ;
      RECT 20.32 3.305 20.886 3.457 ;
      RECT 20.78 3.13 20.95 3.452 ;
      RECT 20.355 3.237 20.98 3.45 ;
      RECT 20.345 3.292 20.985 3.448 ;
      RECT 20.32 3.328 20.995 3.443 ;
      RECT 20.32 3.355 21 3.373 ;
      RECT 20.385 3.18 20.96 3.45 ;
      RECT 20.576 3.165 20.96 3.45 ;
      RECT 20.41 3.168 20.96 3.45 ;
      RECT 20.49 3.166 20.576 3.477 ;
      RECT 20.576 3.163 20.955 3.45 ;
      RECT 20.76 3.14 20.955 3.45 ;
      RECT 20.662 3.161 20.955 3.45 ;
      RECT 20.745 3.155 20.76 3.463 ;
      RECT 20.895 4.52 20.9 4.72 ;
      RECT 20.36 4.585 20.405 4.72 ;
      RECT 20.93 4.52 20.95 4.693 ;
      RECT 20.9 4.52 20.93 4.708 ;
      RECT 20.835 4.52 20.895 4.745 ;
      RECT 20.82 4.52 20.835 4.775 ;
      RECT 20.805 4.52 20.82 4.788 ;
      RECT 20.785 4.52 20.805 4.803 ;
      RECT 20.78 4.52 20.785 4.812 ;
      RECT 20.77 4.524 20.78 4.817 ;
      RECT 20.755 4.534 20.77 4.828 ;
      RECT 20.73 4.55 20.755 4.838 ;
      RECT 20.72 4.564 20.73 4.84 ;
      RECT 20.7 4.576 20.72 4.837 ;
      RECT 20.67 4.597 20.7 4.831 ;
      RECT 20.66 4.609 20.67 4.826 ;
      RECT 20.65 4.607 20.66 4.823 ;
      RECT 20.635 4.606 20.65 4.818 ;
      RECT 20.63 4.605 20.635 4.813 ;
      RECT 20.595 4.603 20.63 4.803 ;
      RECT 20.575 4.6 20.595 4.785 ;
      RECT 20.565 4.598 20.575 4.78 ;
      RECT 20.555 4.597 20.565 4.775 ;
      RECT 20.52 4.595 20.555 4.763 ;
      RECT 20.465 4.591 20.52 4.743 ;
      RECT 20.455 4.589 20.465 4.728 ;
      RECT 20.45 4.589 20.455 4.723 ;
      RECT 20.405 4.587 20.45 4.72 ;
      RECT 20.31 4.585 20.36 4.724 ;
      RECT 20.3 4.586 20.31 4.729 ;
      RECT 20.24 4.593 20.3 4.743 ;
      RECT 20.215 4.601 20.24 4.763 ;
      RECT 20.205 4.605 20.215 4.775 ;
      RECT 20.2 4.606 20.205 4.78 ;
      RECT 20.185 4.608 20.2 4.783 ;
      RECT 20.17 4.61 20.185 4.788 ;
      RECT 20.165 4.61 20.17 4.791 ;
      RECT 20.12 4.615 20.165 4.802 ;
      RECT 20.115 4.619 20.12 4.814 ;
      RECT 20.09 4.615 20.115 4.818 ;
      RECT 20.08 4.611 20.09 4.822 ;
      RECT 20.07 4.61 20.08 4.826 ;
      RECT 20.055 4.6 20.07 4.832 ;
      RECT 20.05 4.588 20.055 4.836 ;
      RECT 20.045 4.585 20.05 4.837 ;
      RECT 20.04 4.582 20.045 4.839 ;
      RECT 20.025 4.57 20.04 4.838 ;
      RECT 20.01 4.552 20.025 4.835 ;
      RECT 19.99 4.531 20.01 4.828 ;
      RECT 19.925 4.52 19.99 4.8 ;
      RECT 19.921 4.52 19.925 4.779 ;
      RECT 19.835 4.52 19.921 4.749 ;
      RECT 19.82 4.52 19.835 4.705 ;
      RECT 20.47 4.871 20.485 5.13 ;
      RECT 20.47 4.886 20.49 5.129 ;
      RECT 20.386 4.886 20.49 5.127 ;
      RECT 20.386 4.9 20.495 5.126 ;
      RECT 20.3 4.942 20.5 5.123 ;
      RECT 20.295 4.885 20.485 5.118 ;
      RECT 20.295 4.956 20.505 5.115 ;
      RECT 20.29 4.987 20.505 5.113 ;
      RECT 20.295 4.984 20.52 5.103 ;
      RECT 20.29 5.03 20.535 5.088 ;
      RECT 20.29 5.058 20.54 5.073 ;
      RECT 20.3 4.86 20.47 5.123 ;
      RECT 20.06 3.87 20.23 4.04 ;
      RECT 20.025 3.87 20.23 4.035 ;
      RECT 20.015 3.87 20.23 4.028 ;
      RECT 20.01 3.855 20.18 4.025 ;
      RECT 18.84 4.392 19.105 4.835 ;
      RECT 18.835 4.363 19.05 4.833 ;
      RECT 18.83 4.517 19.11 4.828 ;
      RECT 18.835 4.412 19.11 4.828 ;
      RECT 18.835 4.423 19.12 4.815 ;
      RECT 18.835 4.37 19.08 4.833 ;
      RECT 18.84 4.357 19.05 4.835 ;
      RECT 18.84 4.355 19 4.835 ;
      RECT 18.941 4.347 19 4.835 ;
      RECT 18.855 4.348 19 4.835 ;
      RECT 18.941 4.346 18.99 4.835 ;
      RECT 18.745 3.161 18.92 3.46 ;
      RECT 18.795 3.123 18.92 3.46 ;
      RECT 18.78 3.125 19.006 3.452 ;
      RECT 18.78 3.128 19.045 3.439 ;
      RECT 18.78 3.129 19.055 3.425 ;
      RECT 18.735 3.18 19.055 3.415 ;
      RECT 18.78 3.13 19.06 3.41 ;
      RECT 18.735 3.34 19.065 3.4 ;
      RECT 18.72 3.2 19.06 3.34 ;
      RECT 18.715 3.216 19.06 3.28 ;
      RECT 18.76 3.14 19.06 3.41 ;
      RECT 18.795 3.121 18.881 3.46 ;
      RECT 16.605 7.31 16.775 9.52 ;
      RECT 16.605 7.31 16.78 8.57 ;
      RECT 16.175 10.15 16.345 10.6 ;
      RECT 16.235 8.37 16.405 10.32 ;
      RECT 16.175 7.31 16.345 8.54 ;
      RECT 15.65 10.11 15.825 10.6 ;
      RECT 15.65 7.31 15.82 10.6 ;
      RECT 15.65 9.61 16.06 9.94 ;
      RECT 15.65 8.77 16.06 9.1 ;
      RECT 15.65 7.31 15.825 8.57 ;
      RECT 93.555 10.09 93.73 10.6 ;
      RECT 92.565 1.865 92.74 2.375 ;
      RECT 92.565 10.09 92.74 10.6 ;
      RECT 90.775 1.865 90.95 2.375 ;
      RECT 90.775 10.09 90.95 10.6 ;
      RECT 85.14 10.09 85.315 10.6 ;
      RECT 78.295 10.09 78.47 10.6 ;
      RECT 77.305 1.865 77.48 2.375 ;
      RECT 77.305 10.09 77.48 10.6 ;
      RECT 75.515 1.865 75.69 2.375 ;
      RECT 75.515 10.09 75.69 10.6 ;
      RECT 69.88 10.09 70.055 10.6 ;
      RECT 63.035 10.09 63.21 10.6 ;
      RECT 62.045 1.865 62.22 2.375 ;
      RECT 62.045 10.09 62.22 10.6 ;
      RECT 60.255 1.865 60.43 2.375 ;
      RECT 60.255 10.09 60.43 10.6 ;
      RECT 54.62 10.09 54.795 10.6 ;
      RECT 47.775 10.09 47.95 10.6 ;
      RECT 46.785 1.865 46.96 2.375 ;
      RECT 46.785 10.09 46.96 10.6 ;
      RECT 44.995 1.865 45.17 2.375 ;
      RECT 44.995 10.09 45.17 10.6 ;
      RECT 39.36 10.09 39.535 10.6 ;
      RECT 32.515 10.09 32.69 10.6 ;
      RECT 31.525 1.865 31.7 2.375 ;
      RECT 31.525 10.09 31.7 10.6 ;
      RECT 29.735 1.865 29.91 2.375 ;
      RECT 29.735 10.09 29.91 10.6 ;
      RECT 24.1 10.09 24.275 10.6 ;
      RECT 16.605 10.09 16.78 10.6 ;
  END
END sky130_osu_ring_oscillator_mpr2ya_8_b0r2

END LIBRARY
