magic
tech sky130A
magscale 1 2
timestamp 1712692843
<< nwell >>
rect 3010 1410 5944 1749
rect 8910 1636 8968 1694
rect 12622 1636 12680 1694
rect 16334 1636 16392 1694
rect 20046 1636 20104 1694
rect 3000 1090 22120 1410
rect 3001 1019 5944 1090
rect 7151 987 7209 1045
rect 10863 987 10921 1045
rect 14575 987 14633 1045
rect 18287 987 18345 1045
rect 21999 987 22057 1045
<< ndiff >>
rect 7162 442 7197 476
rect 10874 442 10909 476
rect 14586 442 14621 476
rect 18298 442 18333 476
rect 22010 442 22045 476
<< pdiff >>
rect 3046 1648 3080 1682
rect 5210 1647 5244 1681
rect 8910 1636 8968 1694
rect 12622 1636 12680 1694
rect 16334 1636 16392 1694
rect 20046 1636 20104 1694
<< locali >>
rect 1 2173 22120 2493
rect 3407 1410 3441 1473
rect 0 1090 22120 1410
rect 1 0 22120 320
<< viali >>
rect 3046 1648 3080 1682
rect 7162 442 7197 476
rect 10874 442 10909 476
rect 14586 442 14621 476
rect 18298 442 18333 476
rect 22010 442 22045 476
<< metal1 >>
rect 1 2173 22120 2493
rect 22043 1983 22046 2017
rect 22006 1977 22076 1983
rect 3303 1863 3309 1921
rect 3367 1863 3373 1921
rect 22006 1919 22012 1977
rect 22070 1919 22076 1977
rect 22006 1913 22076 1919
rect 7162 1853 7232 1859
rect 5599 1843 5669 1849
rect 5599 1785 5605 1843
rect 5663 1785 5669 1843
rect 7162 1795 7168 1853
rect 7226 1795 7232 1853
rect 10873 1854 10944 1861
rect 7162 1789 7232 1795
rect 9311 1844 9381 1850
rect 5599 1779 5669 1785
rect 9311 1786 9317 1844
rect 9375 1786 9381 1844
rect 10873 1796 10880 1854
rect 10938 1796 10944 1854
rect 14577 1853 14647 1859
rect 10873 1790 10944 1796
rect 13022 1845 13092 1851
rect 9311 1780 9381 1786
rect 13022 1787 13028 1845
rect 13086 1787 13092 1845
rect 14577 1795 14583 1853
rect 14641 1795 14647 1853
rect 18289 1853 18359 1859
rect 14577 1789 14647 1795
rect 16734 1844 16804 1850
rect 13022 1781 13092 1787
rect 16734 1786 16740 1844
rect 16798 1786 16804 1844
rect 18289 1795 18295 1853
rect 18353 1795 18359 1853
rect 18289 1789 18359 1795
rect 20446 1844 20516 1850
rect 16734 1780 16804 1786
rect 20446 1786 20452 1844
rect 20510 1786 20516 1844
rect 20446 1780 20516 1786
rect 3228 1715 3234 1773
rect 3292 1715 3298 1773
rect 3035 1682 3093 1687
rect 3035 1648 3046 1682
rect 3080 1648 3093 1682
rect 3035 1641 3093 1648
rect 0 1090 22120 1410
rect 1 0 22120 320
<< via1 >>
rect 3309 1863 3367 1921
rect 22012 1919 22070 1977
rect 5605 1785 5663 1843
rect 7168 1795 7226 1853
rect 9317 1786 9375 1844
rect 10880 1796 10938 1854
rect 13028 1787 13086 1845
rect 14583 1795 14641 1853
rect 16740 1786 16798 1844
rect 18295 1795 18353 1853
rect 20452 1786 20510 1844
rect 3234 1715 3292 1773
rect 5198 1636 5256 1694
rect 8910 1636 8968 1694
rect 12622 1636 12680 1694
rect 16334 1636 16392 1694
rect 20046 1636 20104 1694
rect 7151 987 7209 1045
rect 10863 987 10921 1045
rect 14575 987 14633 1045
rect 18287 987 18345 1045
rect 21999 987 22057 1045
<< metal2 >>
rect 3247 2138 22046 2172
rect 3247 1779 3281 2138
rect 22012 1983 22046 2138
rect 22006 1977 22076 1983
rect 3309 1921 3367 1927
rect 22006 1919 22012 1977
rect 22070 1919 22076 1977
rect 22006 1913 22076 1919
rect 3367 1868 3572 1902
rect 3309 1857 3367 1863
rect 3538 1829 3572 1868
rect 7162 1853 7232 1859
rect 5599 1843 5669 1849
rect 5599 1829 5605 1843
rect 3538 1795 5605 1829
rect 5599 1785 5605 1795
rect 5663 1785 5669 1843
rect 7162 1795 7168 1853
rect 7226 1835 7232 1853
rect 10874 1854 10944 1860
rect 9311 1844 9381 1850
rect 9311 1835 9317 1844
rect 7226 1795 9317 1835
rect 7162 1789 7232 1795
rect 5599 1779 5669 1785
rect 9311 1786 9317 1795
rect 9375 1786 9381 1844
rect 10874 1796 10880 1854
rect 10938 1836 10944 1854
rect 14577 1853 14647 1859
rect 13022 1845 13092 1851
rect 13022 1836 13028 1845
rect 10938 1796 13028 1836
rect 10874 1790 10944 1796
rect 9311 1780 9381 1786
rect 13022 1787 13028 1796
rect 13086 1787 13092 1845
rect 14577 1795 14583 1853
rect 14641 1835 14647 1853
rect 18289 1853 18359 1859
rect 16734 1844 16804 1850
rect 16734 1835 16740 1844
rect 14641 1795 16740 1835
rect 14577 1789 14647 1795
rect 13022 1781 13092 1787
rect 16734 1786 16740 1795
rect 16798 1786 16804 1844
rect 18289 1795 18295 1853
rect 18353 1835 18359 1853
rect 20446 1844 20516 1850
rect 20446 1835 20452 1844
rect 18353 1795 20452 1835
rect 18289 1789 18359 1795
rect 16734 1780 16804 1786
rect 20446 1786 20452 1795
rect 20510 1786 20516 1844
rect 20446 1780 20516 1786
rect 3234 1773 3292 1779
rect 3234 1709 3292 1715
<< via2 >>
rect 5198 1636 5256 1694
rect 8910 1636 8968 1694
rect 12622 1636 12680 1694
rect 16334 1636 16392 1694
rect 20046 1636 20104 1694
rect 7151 987 7209 1045
rect 10863 987 10921 1045
rect 14575 987 14633 1045
rect 18287 987 18345 1045
rect 21999 987 22057 1045
<< metal3 >>
rect 5194 1694 5259 2472
rect 8906 1694 8971 2472
rect 12618 1694 12683 2472
rect 16330 1694 16395 2472
rect 20042 1694 20107 2472
rect 7142 0 7218 987
rect 10854 0 10930 987
rect 14566 0 14642 987
rect 18278 0 18354 987
rect 21990 0 22066 987
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_0
timestamp 1710278372
transform 1 0 3010 0 -1 2234
box -10 0 552 902
use sky130_osu_single_mpr2et_8_b0r1  sky130_osu_single_mpr2et_8_b0r1_0
timestamp 1712692843
transform 1 0 18407 0 1 0
box 0 0 3716 2493
use sky130_osu_single_mpr2et_8_b0r1  sky130_osu_single_mpr2et_8_b0r1_1
timestamp 1712692843
transform 1 0 3559 0 1 0
box 0 0 3716 2493
use sky130_osu_single_mpr2et_8_b0r1  sky130_osu_single_mpr2et_8_b0r1_2
timestamp 1712692843
transform 1 0 7271 0 1 0
box 0 0 3716 2493
use sky130_osu_single_mpr2et_8_b0r1  sky130_osu_single_mpr2et_8_b0r1_3
timestamp 1712692843
transform 1 0 10983 0 1 0
box 0 0 3716 2493
use sky130_osu_single_mpr2et_8_b0r1  sky130_osu_single_mpr2et_8_b0r1_4
timestamp 1712692843
transform 1 0 14695 0 1 0
box 0 0 3716 2493
<< labels >>
flabel metal1 s 3035 1641 3093 1687 0 FreeSans 100 0 0 0 start
port 13 nsew signal input
flabel metal1 s 7162 442 7197 476 0 FreeSans 100 0 0 0 X1_Y1
port 6 s signal output
flabel metal1 s 10874 442 10909 476 0 FreeSans 100 0 0 0 X2_Y1
port 7 s signal output
flabel metal1 s 14586 442 14621 476 0 FreeSans 100 0 0 0 X3_Y1
port 8 s signal output
flabel metal1 s 18298 442 18333 476 0 FreeSans 100 0 0 0 X4_Y1
port 9 s signal output
flabel metal1 s 22010 442 22045 476 0 FreeSans 100 0 0 0 X5_Y1
port 10 s signal output
flabel metal1 s 1 2173 22120 2493 0 FreeSans 100 0 0 0 vssd1
port 14 nsew ground bidirectional
flabel metal1 s 0 1090 22120 1410 0 FreeSans 100 0 0 0 vccd1
port 15 nsew power bidirectional
flabel metal1 s 1 0 22120 320 0 FreeSans 100 0 0 0 vssd1
port 14 nsew ground bidirectional
flabel metal1 s 5209 1648 5243 1682 0 FreeSans 100 0 0 0 s1
port 1 n signal input
flabel metal1 s 8921 1648 8955 1682 0 FreeSans 100 0 0 0 s2
port 2 n signal input
flabel metal1 s 12633 1648 12667 1682 0 FreeSans 100 0 0 0 s3
port 3 n signal input
flabel metal1 s 16345 1648 16379 1682 0 FreeSans 100 0 0 0 s4
port 4 n signal input
flabel metal1 s 20057 1648 20091 1682 0 FreeSans 100 0 0 0 s5
port 5 n signal input
<< end >>
