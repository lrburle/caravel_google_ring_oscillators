VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1426.380 2924.800 1427.580 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3486.100 2.400 3487.300 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3224.980 2.400 3226.180 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2964.540 2.400 2965.740 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1692.260 2924.800 1693.460 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2703.420 2.400 2704.620 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2442.980 2.400 2444.180 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2182.540 2.400 2183.740 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1921.420 2.400 1922.620 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1660.980 2.400 1662.180 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 2.400 1401.060 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1139.420 2.400 1140.620 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 878.980 2.400 880.180 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 617.860 2.400 619.060 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1958.140 2924.800 1959.340 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2223.340 2924.800 2224.540 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2489.220 2924.800 2490.420 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2755.100 2924.800 2756.300 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3020.300 2924.800 3021.500 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3286.180 2924.800 3287.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 32.380 2924.800 33.580 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2289.980 2924.800 2291.180 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2555.860 2924.800 2557.060 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2821.060 2924.800 2822.260 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3086.940 2924.800 3088.140 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3352.820 2924.800 3354.020 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 230.940 2924.800 232.140 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3420.820 2.400 3422.020 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3159.700 2.400 3160.900 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2899.260 2.400 2900.460 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2638.820 2.400 2640.020 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2377.700 2.400 2378.900 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2117.260 2.400 2118.460 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 430.180 2924.800 431.380 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1856.140 2.400 1857.340 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1595.700 2.400 1596.900 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1335.260 2.400 1336.460 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1074.140 2.400 1075.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 813.700 2.400 814.900 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 552.580 2.400 553.780 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 357.420 2.400 358.620 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 161.580 2.400 162.780 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 629.420 2924.800 630.620 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 828.660 2924.800 829.860 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1027.900 2924.800 1029.100 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1227.140 2924.800 1228.340 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1493.020 2924.800 1494.220 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1758.900 2924.800 1760.100 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2024.100 2924.800 2025.300 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 164.980 2924.800 166.180 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2422.580 2924.800 2423.780 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2688.460 2924.800 2689.660 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2954.340 2924.800 2955.540 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3219.540 2924.800 3220.740 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3485.420 2924.800 3486.620 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 364.220 2924.800 365.420 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3290.260 2.400 3291.460 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3029.820 2.400 3031.020 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2768.700 2.400 2769.900 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2508.260 2.400 2509.460 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2247.140 2.400 2248.340 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1986.700 2.400 1987.900 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 563.460 2924.800 564.660 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1726.260 2.400 1727.460 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1465.140 2.400 1466.340 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1204.700 2.400 1205.900 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 943.580 2.400 944.780 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 683.140 2.400 684.340 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 422.700 2.400 423.900 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 226.860 2.400 228.060 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 31.700 2.400 32.900 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 762.700 2924.800 763.900 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 961.940 2924.800 963.140 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1161.180 2924.800 1162.380 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1360.420 2924.800 1361.620 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1625.620 2924.800 1626.820 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1891.500 2924.800 1892.700 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2157.380 2924.800 2158.580 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 98.340 2924.800 99.540 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2356.620 2924.800 2357.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2621.820 2924.800 2623.020 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2887.700 2924.800 2888.900 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3153.580 2924.800 3154.780 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3418.780 2924.800 3419.980 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 297.580 2924.800 298.780 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3355.540 2.400 3356.740 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3095.100 2.400 3096.300 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2833.980 2.400 2835.180 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2573.540 2.400 2574.740 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2312.420 2.400 2313.620 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2051.980 2.400 2053.180 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 496.820 2924.800 498.020 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1791.540 2.400 1792.740 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1530.420 2.400 1531.620 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1269.980 2.400 1271.180 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1008.860 2.400 1010.060 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 748.420 2.400 749.620 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 487.300 2.400 488.500 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 292.140 2.400 293.340 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 96.300 2.400 97.500 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 696.060 2924.800 697.260 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 895.300 2924.800 896.500 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1094.540 2924.800 1095.740 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1293.780 2924.800 1294.980 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1559.660 2924.800 1560.860 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1824.860 2924.800 1826.060 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2090.740 2924.800 2091.940 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.230 -4.800 629.790 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2402.530 -4.800 2403.090 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2420.010 -4.800 2420.570 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2437.950 -4.800 2438.510 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2455.430 -4.800 2455.990 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.370 -4.800 2473.930 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2490.850 -4.800 2491.410 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2508.790 -4.800 2509.350 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2526.730 -4.800 2527.290 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2544.210 -4.800 2544.770 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2562.150 -4.800 2562.710 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.330 -4.800 806.890 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2579.630 -4.800 2580.190 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2597.570 -4.800 2598.130 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2615.050 -4.800 2615.610 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2632.990 -4.800 2633.550 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2650.470 -4.800 2651.030 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2668.410 -4.800 2668.970 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2685.890 -4.800 2686.450 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2703.830 -4.800 2704.390 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2721.770 -4.800 2722.330 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2739.250 -4.800 2739.810 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.270 -4.800 824.830 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2757.190 -4.800 2757.750 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2774.670 -4.800 2775.230 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2792.610 -4.800 2793.170 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2810.090 -4.800 2810.650 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2828.030 -4.800 2828.590 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2845.510 -4.800 2846.070 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2863.450 -4.800 2864.010 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2881.390 -4.800 2881.950 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.750 -4.800 842.310 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.690 -4.800 860.250 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.170 -4.800 877.730 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.110 -4.800 895.670 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.530 -4.800 931.090 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.470 -4.800 949.030 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.710 -4.800 647.270 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.370 -4.800 1001.930 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.790 -4.800 1037.350 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.730 -4.800 1055.290 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.210 -4.800 1072.770 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.150 -4.800 1090.710 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.630 -4.800 1108.190 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.570 -4.800 1126.130 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.510 -4.800 1144.070 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.650 -4.800 665.210 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.990 -4.800 1161.550 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.930 -4.800 1179.490 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.410 -4.800 1196.970 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.350 -4.800 1214.910 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.830 -4.800 1232.390 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.770 -4.800 1250.330 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1267.250 -4.800 1267.810 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.190 -4.800 1285.750 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1303.130 -4.800 1303.690 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.610 -4.800 1321.170 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.130 -4.800 682.690 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.550 -4.800 1339.110 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.030 -4.800 1356.590 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.970 -4.800 1374.530 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.450 -4.800 1392.010 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.390 -4.800 1409.950 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.870 -4.800 1427.430 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.810 -4.800 1445.370 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.750 -4.800 1463.310 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1480.230 -4.800 1480.790 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1498.170 -4.800 1498.730 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.070 -4.800 700.630 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.650 -4.800 1516.210 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1533.590 -4.800 1534.150 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1551.070 -4.800 1551.630 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1569.010 -4.800 1569.570 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1586.490 -4.800 1587.050 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1604.430 -4.800 1604.990 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.910 -4.800 1622.470 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.850 -4.800 1640.410 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.790 -4.800 1658.350 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.270 -4.800 1675.830 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.550 -4.800 718.110 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.210 -4.800 1693.770 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.690 -4.800 1711.250 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.630 -4.800 1729.190 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1746.110 -4.800 1746.670 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.050 -4.800 1764.610 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1781.530 -4.800 1782.090 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.470 -4.800 1800.030 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1817.410 -4.800 1817.970 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1834.890 -4.800 1835.450 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1852.830 -4.800 1853.390 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.490 -4.800 736.050 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.310 -4.800 1870.870 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1888.250 -4.800 1888.810 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.670 -4.800 1924.230 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1976.570 -4.800 1977.130 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.510 -4.800 1995.070 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2029.930 -4.800 2030.490 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.970 -4.800 753.530 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2047.870 -4.800 2048.430 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2065.350 -4.800 2065.910 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2083.290 -4.800 2083.850 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2100.770 -4.800 2101.330 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.710 -4.800 2119.270 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2136.190 -4.800 2136.750 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2154.130 -4.800 2154.690 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2172.070 -4.800 2172.630 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2189.550 -4.800 2190.110 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2207.490 -4.800 2208.050 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.910 -4.800 771.470 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2224.970 -4.800 2225.530 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2242.910 -4.800 2243.470 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2260.390 -4.800 2260.950 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2278.330 -4.800 2278.890 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.810 -4.800 2296.370 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2313.750 -4.800 2314.310 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2331.230 -4.800 2331.790 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2349.170 -4.800 2349.730 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2367.110 -4.800 2367.670 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2384.590 -4.800 2385.150 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.850 -4.800 789.410 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.750 -4.800 635.310 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2408.510 -4.800 2409.070 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2425.990 -4.800 2426.550 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2443.930 -4.800 2444.490 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2461.410 -4.800 2461.970 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2479.350 -4.800 2479.910 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2496.830 -4.800 2497.390 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2514.770 -4.800 2515.330 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2532.250 -4.800 2532.810 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2550.190 -4.800 2550.750 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2567.670 -4.800 2568.230 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.310 -4.800 812.870 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2585.610 -4.800 2586.170 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2603.550 -4.800 2604.110 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2621.030 -4.800 2621.590 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2638.970 -4.800 2639.530 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2656.450 -4.800 2657.010 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2674.390 -4.800 2674.950 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2691.870 -4.800 2692.430 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2709.810 -4.800 2710.370 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2727.290 -4.800 2727.850 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2745.230 -4.800 2745.790 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.250 -4.800 830.810 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2763.170 -4.800 2763.730 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2780.650 -4.800 2781.210 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.590 -4.800 2799.150 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2816.070 -4.800 2816.630 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2834.010 -4.800 2834.570 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2851.490 -4.800 2852.050 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2869.430 -4.800 2869.990 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.730 -4.800 848.290 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.670 -4.800 866.230 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.150 -4.800 883.710 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.090 -4.800 901.650 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.510 -4.800 937.070 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.690 -4.800 653.250 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.410 -4.800 989.970 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.770 -4.800 1043.330 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.710 -4.800 1061.270 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.190 -4.800 1078.750 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.130 -4.800 1096.690 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.610 -4.800 1114.170 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.550 -4.800 1132.110 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.030 -4.800 1149.590 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.630 -4.800 671.190 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.970 -4.800 1167.530 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.910 -4.800 1185.470 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.390 -4.800 1202.950 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.330 -4.800 1220.890 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.810 -4.800 1238.370 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.750 -4.800 1256.310 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.230 -4.800 1273.790 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.170 -4.800 1291.730 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.650 -4.800 1309.210 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.590 -4.800 1327.150 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.110 -4.800 688.670 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.070 -4.800 1344.630 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.010 -4.800 1362.570 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.950 -4.800 1380.510 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.430 -4.800 1397.990 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.370 -4.800 1415.930 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.850 -4.800 1433.410 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1450.790 -4.800 1451.350 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.270 -4.800 1468.830 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.210 -4.800 1486.770 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.690 -4.800 1504.250 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.050 -4.800 706.610 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.630 -4.800 1522.190 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.570 -4.800 1540.130 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.050 -4.800 1557.610 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.990 -4.800 1575.550 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.470 -4.800 1593.030 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.410 -4.800 1610.970 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.890 -4.800 1628.450 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.830 -4.800 1646.390 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1663.310 -4.800 1663.870 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1681.250 -4.800 1681.810 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.530 -4.800 724.090 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1699.190 -4.800 1699.750 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.670 -4.800 1717.230 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1734.610 -4.800 1735.170 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1752.090 -4.800 1752.650 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.030 -4.800 1770.590 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.510 -4.800 1788.070 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1805.450 -4.800 1806.010 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.930 -4.800 1823.490 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1840.870 -4.800 1841.430 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.350 -4.800 1858.910 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.470 -4.800 742.030 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1876.290 -4.800 1876.850 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1894.230 -4.800 1894.790 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1929.650 -4.800 1930.210 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1982.550 -4.800 1983.110 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000.490 -4.800 2001.050 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2017.970 -4.800 2018.530 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.910 -4.800 2036.470 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.950 -4.800 759.510 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2053.850 -4.800 2054.410 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2071.330 -4.800 2071.890 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.270 -4.800 2089.830 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2106.750 -4.800 2107.310 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2124.690 -4.800 2125.250 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2142.170 -4.800 2142.730 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.110 -4.800 2160.670 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2177.590 -4.800 2178.150 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2195.530 -4.800 2196.090 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2213.010 -4.800 2213.570 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.890 -4.800 777.450 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.950 -4.800 2231.510 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2248.890 -4.800 2249.450 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2266.370 -4.800 2266.930 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2284.310 -4.800 2284.870 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.790 -4.800 2302.350 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2319.730 -4.800 2320.290 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2337.210 -4.800 2337.770 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2355.150 -4.800 2355.710 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2372.630 -4.800 2373.190 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2390.570 -4.800 2391.130 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.370 -4.800 794.930 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.730 -4.800 641.290 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2414.030 -4.800 2414.590 2.400 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2431.970 -4.800 2432.530 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2449.450 -4.800 2450.010 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2467.390 -4.800 2467.950 2.400 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2485.330 -4.800 2485.890 2.400 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2502.810 -4.800 2503.370 2.400 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2520.750 -4.800 2521.310 2.400 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2538.230 -4.800 2538.790 2.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2556.170 -4.800 2556.730 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2573.650 -4.800 2574.210 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.290 -4.800 818.850 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2591.590 -4.800 2592.150 2.400 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2609.070 -4.800 2609.630 2.400 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2627.010 -4.800 2627.570 2.400 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2644.950 -4.800 2645.510 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2662.430 -4.800 2662.990 2.400 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2680.370 -4.800 2680.930 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2697.850 -4.800 2698.410 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2715.790 -4.800 2716.350 2.400 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2733.270 -4.800 2733.830 2.400 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2751.210 -4.800 2751.770 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.770 -4.800 836.330 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2768.690 -4.800 2769.250 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2786.630 -4.800 2787.190 2.400 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2804.110 -4.800 2804.670 2.400 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2822.050 -4.800 2822.610 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2839.990 -4.800 2840.550 2.400 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2857.470 -4.800 2858.030 2.400 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2875.410 -4.800 2875.970 2.400 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.710 -4.800 854.270 2.400 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.190 -4.800 871.750 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.130 -4.800 889.690 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.070 -4.800 907.630 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.550 -4.800 925.110 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.490 -4.800 943.050 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.670 -4.800 659.230 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.390 -4.800 995.950 2.400 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.810 -4.800 1031.370 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.750 -4.800 1049.310 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.690 -4.800 1067.250 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.170 -4.800 1084.730 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.110 -4.800 1102.670 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.590 -4.800 1120.150 2.400 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.530 -4.800 1138.090 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.010 -4.800 1155.570 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.150 -4.800 676.710 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.950 -4.800 1173.510 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.430 -4.800 1190.990 2.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.370 -4.800 1208.930 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.850 -4.800 1226.410 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.790 -4.800 1244.350 2.400 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.730 -4.800 1262.290 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.210 -4.800 1279.770 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.150 -4.800 1297.710 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.630 -4.800 1315.190 2.400 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.570 -4.800 1333.130 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.090 -4.800 694.650 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1350.050 -4.800 1350.610 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.990 -4.800 1368.550 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.470 -4.800 1386.030 2.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.410 -4.800 1403.970 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.350 -4.800 1421.910 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.830 -4.800 1439.390 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.770 -4.800 1457.330 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.250 -4.800 1474.810 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.190 -4.800 1492.750 2.400 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1509.670 -4.800 1510.230 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.030 -4.800 712.590 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1527.610 -4.800 1528.170 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.090 -4.800 1545.650 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1563.030 -4.800 1563.590 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.970 -4.800 1581.530 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1598.450 -4.800 1599.010 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.390 -4.800 1616.950 2.400 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.870 -4.800 1634.430 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.810 -4.800 1652.370 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1669.290 -4.800 1669.850 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.230 -4.800 1687.790 2.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.510 -4.800 730.070 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.710 -4.800 1705.270 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.650 -4.800 1723.210 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1740.130 -4.800 1740.690 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.070 -4.800 1758.630 2.400 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.010 -4.800 1776.570 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.490 -4.800 1794.050 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1811.430 -4.800 1811.990 2.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.910 -4.800 1829.470 2.400 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1846.850 -4.800 1847.410 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.330 -4.800 1864.890 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.450 -4.800 748.010 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1882.270 -4.800 1882.830 2.400 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.630 -4.800 1936.190 2.400 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1988.530 -4.800 1989.090 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2023.950 -4.800 2024.510 2.400 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.890 -4.800 2042.450 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.930 -4.800 765.490 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2059.370 -4.800 2059.930 2.400 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2077.310 -4.800 2077.870 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2094.790 -4.800 2095.350 2.400 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.730 -4.800 2113.290 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.670 -4.800 2131.230 2.400 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2148.150 -4.800 2148.710 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2166.090 -4.800 2166.650 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.570 -4.800 2184.130 2.400 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2201.510 -4.800 2202.070 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.990 -4.800 2219.550 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.870 -4.800 783.430 2.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2236.930 -4.800 2237.490 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2254.410 -4.800 2254.970 2.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2272.350 -4.800 2272.910 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2290.290 -4.800 2290.850 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2307.770 -4.800 2308.330 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2325.710 -4.800 2326.270 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2343.190 -4.800 2343.750 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2361.130 -4.800 2361.690 2.400 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2378.610 -4.800 2379.170 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2396.550 -4.800 2397.110 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.350 -4.800 800.910 2.400 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -15.990 -10.630 -8.930 3530.310 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.030 -6.670 2935.610 -3.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -12.030 3523.250 2935.610 3526.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2928.550 -10.630 2935.610 3530.310 ;
    END
    PORT
      LAYER met4 ;
        RECT 5.720 -40.270 7.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 75.720 -40.270 77.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 145.720 -40.270 147.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 215.720 -40.270 217.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 285.720 -40.270 287.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 355.720 -40.270 357.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 425.720 -40.270 427.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 495.720 -40.270 497.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 565.720 -40.270 567.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.720 -40.270 637.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 705.720 -40.270 707.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 775.720 -40.270 777.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 845.720 -40.270 847.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 915.720 -40.270 917.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 985.720 -40.270 987.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1055.720 -40.270 1057.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1125.720 -40.270 1127.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1195.720 -40.270 1197.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1265.720 -40.270 1267.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1335.720 -40.270 1337.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1405.720 -40.270 1407.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1475.720 -40.270 1477.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1545.720 -40.270 1547.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1615.720 -40.270 1617.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1685.720 -40.270 1687.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1755.720 -40.270 1757.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1825.720 -40.270 1827.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1895.720 -40.270 1897.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1965.720 -40.270 1967.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2035.720 -40.270 2037.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2105.720 -40.270 2107.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2175.720 -40.270 2177.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2245.720 -40.270 2247.320 981.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 2245.720 1003.200 2247.320 1821.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 2245.720 1843.200 2247.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2315.720 -40.270 2317.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2385.720 -40.270 2387.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2455.720 -40.270 2457.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2525.720 -40.270 2527.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2595.720 -40.270 2597.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2665.720 -40.270 2667.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2735.720 -40.270 2737.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2805.720 -40.270 2807.320 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2875.720 -40.270 2877.320 3559.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 11.080 2996.930 12.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 81.080 2996.930 82.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 151.080 2996.930 152.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 221.080 2996.930 222.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 291.080 2996.930 292.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 361.080 2996.930 362.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 431.080 2996.930 432.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 501.080 2996.930 502.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 571.080 2996.930 572.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 641.080 2996.930 642.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 711.080 2996.930 712.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 781.080 2996.930 782.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 851.080 2996.930 852.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 921.080 2996.930 922.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 991.080 2996.930 992.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1061.080 2996.930 1062.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1131.080 2996.930 1132.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1201.080 2996.930 1202.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1271.080 2996.930 1272.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1341.080 2996.930 1342.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1411.080 2996.930 1412.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1481.080 2996.930 1482.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1551.080 2996.930 1552.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1621.080 2996.930 1622.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1691.080 2996.930 1692.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1761.080 2996.930 1762.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1831.080 2996.930 1832.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1901.080 2996.930 1902.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1971.080 2996.930 1972.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2041.080 2996.930 2042.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2111.080 2996.930 2112.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2181.080 2996.930 2182.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2251.080 2996.930 2252.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2321.080 2996.930 2322.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2391.080 2996.930 2392.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2461.080 2996.930 2462.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2531.080 2996.930 2532.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2601.080 2996.930 2602.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2671.080 2996.930 2672.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2741.080 2996.930 2742.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2811.080 2996.930 2812.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2881.080 2996.930 2882.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2951.080 2996.930 2952.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3021.080 2996.930 3022.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3091.080 2996.930 3092.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3161.080 2996.930 3162.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3231.080 2996.930 3232.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3301.080 2996.930 3302.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3371.080 2996.930 3372.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3441.080 2996.930 3442.680 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -33.510 -28.150 -26.450 3547.830 ;
    END
    PORT
      LAYER met5 ;
        RECT -21.630 -16.270 2941.250 -13.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -21.630 3532.850 2941.250 3535.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2946.070 -28.150 2953.130 3547.830 ;
    END
    PORT
      LAYER met4 ;
        RECT 23.040 -40.270 24.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 93.040 -40.270 94.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 163.040 -40.270 164.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.040 -40.270 234.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 303.040 -40.270 304.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 373.040 -40.270 374.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 443.040 -40.270 444.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 513.040 -40.270 514.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 583.040 -40.270 584.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 653.040 -40.270 654.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 723.040 -40.270 724.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 793.040 -40.270 794.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 863.040 -40.270 864.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 933.040 -40.270 934.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1003.040 -40.270 1004.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1073.040 -40.270 1074.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1143.040 -40.270 1144.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1213.040 -40.270 1214.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1283.040 -40.270 1284.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1353.040 -40.270 1354.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1423.040 -40.270 1424.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.040 -40.270 1494.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1563.040 -40.270 1564.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.040 -40.270 1634.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1703.040 -40.270 1704.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1773.040 -40.270 1774.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1843.040 -40.270 1844.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1913.040 -40.270 1914.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1983.040 -40.270 1984.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2053.040 -40.270 2054.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2123.040 -40.270 2124.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2193.040 -40.270 2194.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2263.040 -40.270 2264.640 981.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 2263.040 1003.200 2264.640 1821.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 2263.040 1843.200 2264.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2333.040 -40.270 2334.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2403.040 -40.270 2404.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2473.040 -40.270 2474.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2543.040 -40.270 2544.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2613.040 -40.270 2614.640 1200.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2613.040 1908.760 2614.640 2000.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2613.040 2108.760 2614.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2683.040 -40.270 2684.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2753.040 -40.270 2754.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2823.040 -40.270 2824.640 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2893.040 -40.270 2894.640 3559.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 21.750 2996.930 23.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 91.750 2996.930 93.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 161.750 2996.930 163.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 231.750 2996.930 233.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 301.750 2996.930 303.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 371.750 2996.930 373.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 441.750 2996.930 443.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 511.750 2996.930 513.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 581.750 2996.930 583.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 651.750 2996.930 653.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 721.750 2996.930 723.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 791.750 2996.930 793.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 861.750 2996.930 863.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 931.750 2996.930 933.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1001.750 2996.930 1003.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1071.750 2996.930 1073.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1141.750 2996.930 1143.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1211.750 2996.930 1213.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1281.750 2996.930 1283.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1351.750 2996.930 1353.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1421.750 2996.930 1423.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1491.750 2996.930 1493.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1561.750 2996.930 1563.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1631.750 2996.930 1633.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1701.750 2996.930 1703.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1771.750 2996.930 1773.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1841.750 2996.930 1843.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1911.750 2996.930 1913.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1981.750 2996.930 1983.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2051.750 2996.930 2053.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2121.750 2996.930 2123.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2191.750 2996.930 2193.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2261.750 2996.930 2263.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2331.750 2996.930 2333.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2401.750 2996.930 2403.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2471.750 2996.930 2473.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2541.750 2996.930 2543.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2611.750 2996.930 2613.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2681.750 2996.930 2683.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2751.750 2996.930 2753.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2821.750 2996.930 2823.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2891.750 2996.930 2893.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2961.750 2996.930 2963.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3031.750 2996.930 3033.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3101.750 2996.930 3103.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3171.750 2996.930 3173.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3241.750 2996.930 3243.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3311.750 2996.930 3313.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3381.750 2996.930 3383.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3451.750 2996.930 3453.350 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -51.030 -45.670 -43.970 3565.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -31.230 -25.870 2950.850 -22.770 ;
    END
    PORT
      LAYER met5 ;
        RECT -31.230 3542.450 2950.850 3545.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 2963.590 -45.670 2970.650 3565.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 40.360 -40.270 41.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 110.360 -40.270 111.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 180.360 -40.270 181.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 250.360 -40.270 251.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 320.360 -40.270 321.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 390.360 -40.270 391.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 460.360 -40.270 461.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 530.360 -40.270 531.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 600.360 -40.270 601.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 670.360 -40.270 671.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 740.360 -40.270 741.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 810.360 -40.270 811.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 880.360 -40.270 881.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 950.360 -40.270 951.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1020.360 -40.270 1021.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1090.360 -40.270 1091.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1160.360 -40.270 1161.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1230.360 -40.270 1231.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1300.360 -40.270 1301.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1370.360 -40.270 1371.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1440.360 -40.270 1441.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1510.360 -40.270 1511.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1580.360 -40.270 1581.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1650.360 -40.270 1651.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1720.360 -40.270 1721.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1790.360 -40.270 1791.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1860.360 -40.270 1861.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1930.360 -40.270 1931.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2000.360 -40.270 2001.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2070.360 -40.270 2071.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2140.360 -40.270 2141.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2210.360 -40.270 2211.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2280.360 -40.270 2281.960 981.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 2280.360 1003.200 2281.960 1821.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 2280.360 1843.200 2281.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2350.360 -40.270 2351.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2420.360 -40.270 2421.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2490.360 -40.270 2491.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2560.360 -40.270 2561.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2630.360 -40.270 2631.960 1200.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2630.360 1708.760 2631.960 1800.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2630.360 1908.760 2631.960 2000.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2630.360 2108.760 2631.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2700.360 -40.270 2701.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2770.360 -40.270 2771.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2840.360 -40.270 2841.960 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2910.360 -40.270 2911.960 3559.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 32.420 2996.930 34.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 102.420 2996.930 104.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 172.420 2996.930 174.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 242.420 2996.930 244.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 312.420 2996.930 314.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 382.420 2996.930 384.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 452.420 2996.930 454.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 522.420 2996.930 524.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 592.420 2996.930 594.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 662.420 2996.930 664.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 732.420 2996.930 734.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 802.420 2996.930 804.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 872.420 2996.930 874.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 942.420 2996.930 944.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1012.420 2996.930 1014.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1082.420 2996.930 1084.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1152.420 2996.930 1154.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1222.420 2996.930 1224.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1292.420 2996.930 1294.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1362.420 2996.930 1364.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1432.420 2996.930 1434.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1502.420 2996.930 1504.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1572.420 2996.930 1574.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1642.420 2996.930 1644.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1712.420 2996.930 1714.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1782.420 2996.930 1784.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1852.420 2996.930 1854.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1922.420 2996.930 1924.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1992.420 2996.930 1994.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2062.420 2996.930 2064.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2132.420 2996.930 2134.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2202.420 2996.930 2204.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2272.420 2996.930 2274.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2342.420 2996.930 2344.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2412.420 2996.930 2414.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2482.420 2996.930 2484.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2552.420 2996.930 2554.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2622.420 2996.930 2624.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2692.420 2996.930 2694.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2762.420 2996.930 2764.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2832.420 2996.930 2834.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2902.420 2996.930 2904.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2972.420 2996.930 2974.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3042.420 2996.930 3044.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3112.420 2996.930 3114.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3182.420 2996.930 3184.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3252.420 2996.930 3254.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3322.420 2996.930 3324.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3392.420 2996.930 3394.020 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3462.420 2996.930 3464.020 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -68.550 -63.190 -61.490 3582.870 ;
    END
    PORT
      LAYER met5 ;
        RECT -40.830 -35.470 2960.450 -32.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -40.830 3552.050 2960.450 3555.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2981.110 -63.190 2988.170 3582.870 ;
    END
    PORT
      LAYER met4 ;
        RECT 57.680 -40.270 59.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 127.680 -40.270 129.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 197.680 -40.270 199.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 267.680 -40.270 269.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 337.680 -40.270 339.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 407.680 -40.270 409.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 477.680 -40.270 479.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 547.680 -40.270 549.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 617.680 -40.270 619.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 687.680 -40.270 689.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 757.680 -40.270 759.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 827.680 -40.270 829.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 897.680 -40.270 899.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 967.680 -40.270 969.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1037.680 -40.270 1039.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1107.680 -40.270 1109.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1177.680 -40.270 1179.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1247.680 -40.270 1249.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1317.680 -40.270 1319.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1387.680 -40.270 1389.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1457.680 -40.270 1459.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1527.680 -40.270 1529.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1597.680 -40.270 1599.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1667.680 -40.270 1669.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1737.680 -40.270 1739.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1807.680 -40.270 1809.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1877.680 -40.270 1879.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1947.680 -40.270 1949.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.680 -40.270 2019.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2087.680 -40.270 2089.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2157.680 -40.270 2159.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2227.680 -40.270 2229.280 981.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 2227.680 1003.200 2229.280 1821.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 2227.680 1843.200 2229.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2297.680 -40.270 2299.280 981.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 2297.680 1003.200 2299.280 1821.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 2297.680 1843.200 2299.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2367.680 -40.270 2369.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2437.680 -40.270 2439.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2507.680 -40.270 2509.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2577.680 -40.270 2579.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2647.680 -40.270 2649.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2717.680 -40.270 2719.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2787.680 -40.270 2789.280 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2857.680 -40.270 2859.280 3559.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 43.090 2996.930 44.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 113.090 2996.930 114.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 183.090 2996.930 184.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 253.090 2996.930 254.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 323.090 2996.930 324.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 393.090 2996.930 394.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 463.090 2996.930 464.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 533.090 2996.930 534.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 603.090 2996.930 604.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 673.090 2996.930 674.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 743.090 2996.930 744.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 813.090 2996.930 814.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 883.090 2996.930 884.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 953.090 2996.930 954.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1023.090 2996.930 1024.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1093.090 2996.930 1094.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1163.090 2996.930 1164.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1233.090 2996.930 1234.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1303.090 2996.930 1304.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1373.090 2996.930 1374.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1443.090 2996.930 1444.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1513.090 2996.930 1514.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1583.090 2996.930 1584.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1653.090 2996.930 1654.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1723.090 2996.930 1724.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1793.090 2996.930 1794.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1863.090 2996.930 1864.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1933.090 2996.930 1934.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2003.090 2996.930 2004.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2073.090 2996.930 2074.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2143.090 2996.930 2144.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2213.090 2996.930 2214.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2283.090 2996.930 2284.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2353.090 2996.930 2354.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2423.090 2996.930 2424.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2493.090 2996.930 2494.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2563.090 2996.930 2564.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2633.090 2996.930 2634.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2703.090 2996.930 2704.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2773.090 2996.930 2774.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2843.090 2996.930 2844.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2913.090 2996.930 2914.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2983.090 2996.930 2984.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3053.090 2996.930 3054.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3123.090 2996.930 3124.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3193.090 2996.930 3194.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3263.090 2996.930 3264.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3333.090 2996.930 3334.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3403.090 2996.930 3404.690 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3473.090 2996.930 3474.690 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -59.790 -54.430 -52.730 3574.110 ;
    END
    PORT
      LAYER met5 ;
        RECT -36.030 -30.670 2955.650 -27.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -36.030 3547.250 2955.650 3550.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2972.350 -54.430 2979.410 3574.110 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.020 -40.270 50.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 119.020 -40.270 120.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 189.020 -40.270 190.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 259.020 -40.270 260.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 329.020 -40.270 330.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 399.020 -40.270 400.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 469.020 -40.270 470.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 539.020 -40.270 540.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 609.020 -40.270 610.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 679.020 -40.270 680.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 749.020 -40.270 750.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 819.020 -40.270 820.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 889.020 -40.270 890.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 959.020 -40.270 960.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1029.020 -40.270 1030.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1099.020 -40.270 1100.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1169.020 -40.270 1170.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1239.020 -40.270 1240.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1309.020 -40.270 1310.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1379.020 -40.270 1380.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1449.020 -40.270 1450.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1519.020 -40.270 1520.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1589.020 -40.270 1590.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1659.020 -40.270 1660.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1729.020 -40.270 1730.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1799.020 -40.270 1800.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1869.020 -40.270 1870.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1939.020 -40.270 1940.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2009.020 -40.270 2010.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2079.020 -40.270 2080.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2149.020 -40.270 2150.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2219.020 -40.270 2220.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2289.020 -40.270 2290.620 981.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 2289.020 1003.200 2290.620 1821.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 2289.020 1843.200 2290.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2359.020 -40.270 2360.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2429.020 -40.270 2430.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2499.020 -40.270 2500.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2569.020 -40.270 2570.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2639.020 -40.270 2640.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2709.020 -40.270 2710.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2779.020 -40.270 2780.620 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2849.020 -40.270 2850.620 3559.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 37.755 2996.930 39.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 107.755 2996.930 109.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 177.755 2996.930 179.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 247.755 2996.930 249.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 317.755 2996.930 319.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 387.755 2996.930 389.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 457.755 2996.930 459.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 527.755 2996.930 529.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 597.755 2996.930 599.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 667.755 2996.930 669.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 737.755 2996.930 739.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 807.755 2996.930 809.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 877.755 2996.930 879.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 947.755 2996.930 949.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1017.755 2996.930 1019.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1087.755 2996.930 1089.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1157.755 2996.930 1159.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1227.755 2996.930 1229.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1297.755 2996.930 1299.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1367.755 2996.930 1369.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1437.755 2996.930 1439.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1507.755 2996.930 1509.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1577.755 2996.930 1579.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1647.755 2996.930 1649.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1717.755 2996.930 1719.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1787.755 2996.930 1789.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1857.755 2996.930 1859.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1927.755 2996.930 1929.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1997.755 2996.930 1999.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2067.755 2996.930 2069.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2137.755 2996.930 2139.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2207.755 2996.930 2209.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2277.755 2996.930 2279.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2347.755 2996.930 2349.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2417.755 2996.930 2419.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2487.755 2996.930 2489.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2557.755 2996.930 2559.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2627.755 2996.930 2629.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2697.755 2996.930 2699.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2767.755 2996.930 2769.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2837.755 2996.930 2839.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2907.755 2996.930 2909.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2977.755 2996.930 2979.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3047.755 2996.930 3049.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3117.755 2996.930 3119.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3187.755 2996.930 3189.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3257.755 2996.930 3259.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3327.755 2996.930 3329.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3397.755 2996.930 3399.355 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3467.755 2996.930 3469.355 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -77.310 -71.950 -70.250 3591.630 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.630 -40.270 2965.250 -37.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.630 3556.850 2965.250 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2989.870 -71.950 2996.930 3591.630 ;
    END
    PORT
      LAYER met4 ;
        RECT 66.340 -40.270 67.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 136.340 -40.270 137.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 206.340 -40.270 207.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 276.340 -40.270 277.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.340 -40.270 347.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 416.340 -40.270 417.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 486.340 -40.270 487.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 556.340 -40.270 557.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 626.340 -40.270 627.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 696.340 -40.270 697.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 766.340 -40.270 767.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 836.340 -40.270 837.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 906.340 -40.270 907.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 976.340 -40.270 977.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1046.340 -40.270 1047.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1116.340 -40.270 1117.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1186.340 -40.270 1187.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1256.340 -40.270 1257.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.340 -40.270 1327.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1396.340 -40.270 1397.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1466.340 -40.270 1467.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1536.340 -40.270 1537.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1606.340 -40.270 1607.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1676.340 -40.270 1677.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1746.340 -40.270 1747.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1816.340 -40.270 1817.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1886.340 -40.270 1887.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1956.340 -40.270 1957.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2026.340 -40.270 2027.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2096.340 -40.270 2097.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2166.340 -40.270 2167.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2236.340 -40.270 2237.940 981.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 2236.340 1003.200 2237.940 1821.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 2236.340 1843.200 2237.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2306.340 -40.270 2307.940 981.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 2306.340 1003.200 2307.940 1821.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 2306.340 1843.200 2307.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2376.340 -40.270 2377.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2446.340 -40.270 2447.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2516.340 -40.270 2517.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2586.340 -40.270 2587.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2656.340 -40.270 2657.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2726.340 -40.270 2727.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2796.340 -40.270 2797.940 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2866.340 -40.270 2867.940 3559.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 48.425 2996.930 50.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 118.425 2996.930 120.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 188.425 2996.930 190.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 258.425 2996.930 260.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 328.425 2996.930 330.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 398.425 2996.930 400.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 468.425 2996.930 470.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 538.425 2996.930 540.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 608.425 2996.930 610.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 678.425 2996.930 680.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 748.425 2996.930 750.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 818.425 2996.930 820.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 888.425 2996.930 890.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 958.425 2996.930 960.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1028.425 2996.930 1030.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1098.425 2996.930 1100.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1168.425 2996.930 1170.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1238.425 2996.930 1240.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1308.425 2996.930 1310.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1378.425 2996.930 1380.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1448.425 2996.930 1450.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1518.425 2996.930 1520.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1588.425 2996.930 1590.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1658.425 2996.930 1660.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1728.425 2996.930 1730.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1798.425 2996.930 1800.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1868.425 2996.930 1870.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1938.425 2996.930 1940.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2008.425 2996.930 2010.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2078.425 2996.930 2080.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2148.425 2996.930 2150.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2218.425 2996.930 2220.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2288.425 2996.930 2290.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2358.425 2996.930 2360.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2428.425 2996.930 2430.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2498.425 2996.930 2500.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2568.425 2996.930 2570.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2638.425 2996.930 2640.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2708.425 2996.930 2710.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2778.425 2996.930 2780.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2848.425 2996.930 2850.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2918.425 2996.930 2920.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2988.425 2996.930 2990.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3058.425 2996.930 3060.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3128.425 2996.930 3130.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3198.425 2996.930 3200.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3268.425 2996.930 3270.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3338.425 2996.930 3340.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3408.425 2996.930 3410.025 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3478.425 2996.930 3480.025 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -24.750 -19.390 -17.690 3539.070 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.830 -11.470 2936.450 -8.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.830 3528.050 2936.450 3531.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2937.310 -19.390 2944.370 3539.070 ;
    END
    PORT
      LAYER met4 ;
        RECT 14.380 -40.270 15.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 84.380 -40.270 85.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 154.380 -40.270 155.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 224.380 -40.270 225.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 294.380 -40.270 295.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 364.380 -40.270 365.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 434.380 -40.270 435.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 504.380 -40.270 505.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 574.380 -40.270 575.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 644.380 -40.270 645.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 714.380 -40.270 715.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 784.380 -40.270 785.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 854.380 -40.270 855.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 924.380 -40.270 925.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 994.380 -40.270 995.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1064.380 -40.270 1065.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1134.380 -40.270 1135.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1204.380 -40.270 1205.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1274.380 -40.270 1275.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1344.380 -40.270 1345.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1414.380 -40.270 1415.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1484.380 -40.270 1485.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1554.380 -40.270 1555.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1624.380 -40.270 1625.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1694.380 -40.270 1695.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1764.380 -40.270 1765.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1834.380 -40.270 1835.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1904.380 -40.270 1905.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1974.380 -40.270 1975.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2044.380 -40.270 2045.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2114.380 -40.270 2115.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2184.380 -40.270 2185.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2254.380 -40.270 2255.980 981.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 2254.380 1003.200 2255.980 1821.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 2254.380 1843.200 2255.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2324.380 -40.270 2325.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2394.380 -40.270 2395.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2464.380 -40.270 2465.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2534.380 -40.270 2535.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2604.380 -40.270 2605.980 1200.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2604.380 2108.760 2605.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2674.380 -40.270 2675.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2744.380 -40.270 2745.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2814.380 -40.270 2815.980 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2884.380 -40.270 2885.980 3559.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 16.415 2996.930 18.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 86.415 2996.930 88.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 156.415 2996.930 158.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 226.415 2996.930 228.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 296.415 2996.930 298.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 366.415 2996.930 368.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 436.415 2996.930 438.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 506.415 2996.930 508.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 576.415 2996.930 578.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 646.415 2996.930 648.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 716.415 2996.930 718.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 786.415 2996.930 788.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 856.415 2996.930 858.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 926.415 2996.930 928.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 996.415 2996.930 998.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1066.415 2996.930 1068.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1136.415 2996.930 1138.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1206.415 2996.930 1208.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1276.415 2996.930 1278.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1346.415 2996.930 1348.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1416.415 2996.930 1418.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1486.415 2996.930 1488.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1556.415 2996.930 1558.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1626.415 2996.930 1628.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1696.415 2996.930 1698.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1766.415 2996.930 1768.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1836.415 2996.930 1838.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1906.415 2996.930 1908.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1976.415 2996.930 1978.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2046.415 2996.930 2048.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2116.415 2996.930 2118.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2186.415 2996.930 2188.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2256.415 2996.930 2258.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2326.415 2996.930 2328.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2396.415 2996.930 2398.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2466.415 2996.930 2468.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2536.415 2996.930 2538.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2606.415 2996.930 2608.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2676.415 2996.930 2678.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2746.415 2996.930 2748.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2816.415 2996.930 2818.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2886.415 2996.930 2888.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2956.415 2996.930 2958.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3026.415 2996.930 3028.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3096.415 2996.930 3098.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3166.415 2996.930 3168.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3236.415 2996.930 3238.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3306.415 2996.930 3308.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3376.415 2996.930 3378.015 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3446.415 2996.930 3448.015 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -42.270 -36.910 -35.210 3556.590 ;
    END
    PORT
      LAYER met5 ;
        RECT -26.430 -21.070 2946.050 -17.970 ;
    END
    PORT
      LAYER met5 ;
        RECT -26.430 3537.650 2946.050 3540.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2954.830 -36.910 2961.890 3556.590 ;
    END
    PORT
      LAYER met4 ;
        RECT 31.700 -40.270 33.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 101.700 -40.270 103.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 171.700 -40.270 173.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 241.700 -40.270 243.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 311.700 -40.270 313.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 381.700 -40.270 383.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 451.700 -40.270 453.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 521.700 -40.270 523.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 591.700 -40.270 593.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 661.700 -40.270 663.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 731.700 -40.270 733.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 801.700 -40.270 803.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 871.700 -40.270 873.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 941.700 -40.270 943.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1011.700 -40.270 1013.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1081.700 -40.270 1083.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1151.700 -40.270 1153.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1221.700 -40.270 1223.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1291.700 -40.270 1293.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1361.700 -40.270 1363.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1431.700 -40.270 1433.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1501.700 -40.270 1503.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1571.700 -40.270 1573.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1641.700 -40.270 1643.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1711.700 -40.270 1713.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1781.700 -40.270 1783.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1851.700 -40.270 1853.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1921.700 -40.270 1923.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1991.700 -40.270 1993.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2061.700 -40.270 2063.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2131.700 -40.270 2133.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2201.700 -40.270 2203.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2271.700 -40.270 2273.300 981.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 2271.700 1003.200 2273.300 1821.180 ;
    END
    PORT
      LAYER met4 ;
        RECT 2271.700 1843.200 2273.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2341.700 -40.270 2343.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2411.700 -40.270 2413.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2481.700 -40.270 2483.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2551.700 -40.270 2553.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2621.700 -40.270 2623.300 1200.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2621.700 1908.760 2623.300 2000.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 2621.700 2108.760 2623.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2691.700 -40.270 2693.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2761.700 -40.270 2763.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2831.700 -40.270 2833.300 3559.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2901.700 -40.270 2903.300 3559.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 27.085 2996.930 28.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 97.085 2996.930 98.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 167.085 2996.930 168.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 237.085 2996.930 238.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 307.085 2996.930 308.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 377.085 2996.930 378.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 447.085 2996.930 448.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 517.085 2996.930 518.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 587.085 2996.930 588.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 657.085 2996.930 658.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 727.085 2996.930 728.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 797.085 2996.930 798.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 867.085 2996.930 868.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 937.085 2996.930 938.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1007.085 2996.930 1008.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1077.085 2996.930 1078.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1147.085 2996.930 1148.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1217.085 2996.930 1218.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1287.085 2996.930 1288.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1357.085 2996.930 1358.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1427.085 2996.930 1428.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1497.085 2996.930 1498.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1567.085 2996.930 1568.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1637.085 2996.930 1638.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1707.085 2996.930 1708.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1777.085 2996.930 1778.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1847.085 2996.930 1848.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1917.085 2996.930 1918.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 1987.085 2996.930 1988.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2057.085 2996.930 2058.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2127.085 2996.930 2128.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2197.085 2996.930 2198.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2267.085 2996.930 2268.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2337.085 2996.930 2338.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2407.085 2996.930 2408.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2477.085 2996.930 2478.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2547.085 2996.930 2548.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2617.085 2996.930 2618.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2687.085 2996.930 2688.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2757.085 2996.930 2758.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2827.085 2996.930 2828.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2897.085 2996.930 2898.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 2967.085 2996.930 2968.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3037.085 2996.930 3038.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3107.085 2996.930 3108.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3177.085 2996.930 3178.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3247.085 2996.930 3248.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3317.085 2996.930 3318.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3387.085 2996.930 3388.685 ;
    END
    PORT
      LAYER met5 ;
        RECT -77.310 3457.085 2996.930 3458.685 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.150 -4.800 239.710 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.630 -4.800 257.190 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.570 -4.800 275.130 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.050 -4.800 292.610 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.990 -4.800 310.550 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.470 -4.800 328.030 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.410 -4.800 345.970 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.890 -4.800 363.450 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.830 -4.800 381.390 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.310 -4.800 398.870 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.590 -4.800 62.150 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.250 -4.800 416.810 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.190 -4.800 434.750 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.670 -4.800 452.230 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.610 -4.800 470.170 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.090 -4.800 487.650 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.030 -4.800 505.590 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.510 -4.800 523.070 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.450 -4.800 541.010 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.930 -4.800 558.490 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.870 -4.800 576.430 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.050 -4.800 85.610 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.810 -4.800 594.370 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.290 -4.800 611.850 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.970 -4.800 109.530 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.430 -4.800 132.990 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.370 -4.800 150.930 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.850 -4.800 168.410 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.790 -4.800 186.350 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.270 -4.800 203.830 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.210 -4.800 221.770 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.650 -4.800 44.210 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.670 -4.800 245.230 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.610 -4.800 263.170 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.090 -4.800 280.650 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.030 -4.800 298.590 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.970 -4.800 316.530 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.450 -4.800 334.010 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.390 -4.800 351.950 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.870 -4.800 369.430 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.810 -4.800 387.370 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.290 -4.800 404.850 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 -4.800 68.130 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.230 -4.800 422.790 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.710 -4.800 440.270 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.650 -4.800 458.210 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.590 -4.800 476.150 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.070 -4.800 493.630 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.010 -4.800 511.570 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.490 -4.800 529.050 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.430 -4.800 546.990 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.910 -4.800 564.470 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.850 -4.800 582.410 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.030 -4.800 91.590 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.330 -4.800 599.890 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.270 -4.800 617.830 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.950 -4.800 115.510 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.410 -4.800 138.970 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.350 -4.800 156.910 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.830 -4.800 174.390 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.770 -4.800 192.330 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.250 -4.800 209.810 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.190 -4.800 227.750 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.630 -4.800 50.190 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.650 -4.800 251.210 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.590 -4.800 269.150 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.070 -4.800 286.630 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.010 -4.800 304.570 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.490 -4.800 322.050 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.430 -4.800 339.990 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.370 -4.800 357.930 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.850 -4.800 375.410 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.790 -4.800 393.350 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.270 -4.800 410.830 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.550 -4.800 74.110 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.210 -4.800 428.770 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 -4.800 446.250 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.630 -4.800 464.190 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.110 -4.800 481.670 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.050 -4.800 499.610 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.530 -4.800 517.090 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.470 -4.800 535.030 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.410 -4.800 552.970 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.890 -4.800 570.450 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.830 -4.800 588.390 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.010 -4.800 97.570 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.310 -4.800 605.870 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.250 -4.800 623.810 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.930 -4.800 121.490 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.390 -4.800 144.950 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.870 -4.800 162.430 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.810 -4.800 180.370 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.750 -4.800 198.310 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.230 -4.800 215.790 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.170 -4.800 233.730 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.610 -4.800 56.170 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.530 -4.800 80.090 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.990 -4.800 103.550 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.450 -4.800 127.010 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 2207.000 884.000 2634.160 2458.315 ;
      LAYER met1 ;
        RECT 2207.000 884.000 2901.150 2463.260 ;
      LAYER met2 ;
        RECT 2220.050 32.795 2901.590 2464.845 ;
      LAYER met3 ;
        RECT 2220.025 2424.180 2917.600 2464.825 ;
        RECT 2220.025 2422.180 2917.200 2424.180 ;
        RECT 2220.025 2358.220 2917.600 2422.180 ;
        RECT 2220.025 2356.220 2917.200 2358.220 ;
        RECT 2220.025 2291.580 2917.600 2356.220 ;
        RECT 2220.025 2289.580 2917.200 2291.580 ;
        RECT 2220.025 2224.940 2917.600 2289.580 ;
        RECT 2220.025 2222.940 2917.200 2224.940 ;
        RECT 2220.025 2158.980 2917.600 2222.940 ;
        RECT 2220.025 2156.980 2917.200 2158.980 ;
        RECT 2220.025 2092.340 2917.600 2156.980 ;
        RECT 2220.025 2090.340 2917.200 2092.340 ;
        RECT 2220.025 2025.700 2917.600 2090.340 ;
        RECT 2220.025 2023.700 2917.200 2025.700 ;
        RECT 2220.025 1959.740 2917.600 2023.700 ;
        RECT 2220.025 1957.740 2917.200 1959.740 ;
        RECT 2220.025 1893.100 2917.600 1957.740 ;
        RECT 2220.025 1891.100 2917.200 1893.100 ;
        RECT 2220.025 1826.460 2917.600 1891.100 ;
        RECT 2220.025 1824.460 2917.200 1826.460 ;
        RECT 2220.025 1760.500 2917.600 1824.460 ;
        RECT 2220.025 1758.500 2917.200 1760.500 ;
        RECT 2220.025 1693.860 2917.600 1758.500 ;
        RECT 2220.025 1691.860 2917.200 1693.860 ;
        RECT 2220.025 1627.220 2917.600 1691.860 ;
        RECT 2220.025 1625.220 2917.200 1627.220 ;
        RECT 2220.025 1561.260 2917.600 1625.220 ;
        RECT 2220.025 1559.260 2917.200 1561.260 ;
        RECT 2220.025 1494.620 2917.600 1559.260 ;
        RECT 2220.025 1492.620 2917.200 1494.620 ;
        RECT 2220.025 1427.980 2917.600 1492.620 ;
        RECT 2220.025 1425.980 2917.200 1427.980 ;
        RECT 2220.025 1362.020 2917.600 1425.980 ;
        RECT 2220.025 1360.020 2917.200 1362.020 ;
        RECT 2220.025 1295.380 2917.600 1360.020 ;
        RECT 2220.025 1293.380 2917.200 1295.380 ;
        RECT 2220.025 1228.740 2917.600 1293.380 ;
        RECT 2220.025 1226.740 2917.200 1228.740 ;
        RECT 2220.025 1162.780 2917.600 1226.740 ;
        RECT 2220.025 1160.780 2917.200 1162.780 ;
        RECT 2220.025 1096.140 2917.600 1160.780 ;
        RECT 2220.025 1094.140 2917.200 1096.140 ;
        RECT 2220.025 1029.500 2917.600 1094.140 ;
        RECT 2220.025 1027.500 2917.200 1029.500 ;
        RECT 2220.025 963.540 2917.600 1027.500 ;
        RECT 2220.025 961.540 2917.200 963.540 ;
        RECT 2220.025 896.900 2917.600 961.540 ;
        RECT 2220.025 894.900 2917.200 896.900 ;
        RECT 2220.025 830.260 2917.600 894.900 ;
        RECT 2220.025 828.260 2917.200 830.260 ;
        RECT 2220.025 764.300 2917.600 828.260 ;
        RECT 2220.025 762.300 2917.200 764.300 ;
        RECT 2220.025 697.660 2917.600 762.300 ;
        RECT 2220.025 695.660 2917.200 697.660 ;
        RECT 2220.025 631.020 2917.600 695.660 ;
        RECT 2220.025 629.020 2917.200 631.020 ;
        RECT 2220.025 565.060 2917.600 629.020 ;
        RECT 2220.025 563.060 2917.200 565.060 ;
        RECT 2220.025 498.420 2917.600 563.060 ;
        RECT 2220.025 496.420 2917.200 498.420 ;
        RECT 2220.025 431.780 2917.600 496.420 ;
        RECT 2220.025 429.780 2917.200 431.780 ;
        RECT 2220.025 365.820 2917.600 429.780 ;
        RECT 2220.025 363.820 2917.200 365.820 ;
        RECT 2220.025 299.180 2917.600 363.820 ;
        RECT 2220.025 297.180 2917.200 299.180 ;
        RECT 2220.025 232.540 2917.600 297.180 ;
        RECT 2220.025 230.540 2917.200 232.540 ;
        RECT 2220.025 166.580 2917.600 230.540 ;
        RECT 2220.025 164.580 2917.200 166.580 ;
        RECT 2220.025 99.940 2917.600 164.580 ;
        RECT 2220.025 97.940 2917.200 99.940 ;
        RECT 2220.025 33.980 2917.600 97.940 ;
        RECT 2220.025 32.815 2917.200 33.980 ;
      LAYER met4 ;
        RECT 2238.340 1842.800 2245.320 2098.160 ;
        RECT 2247.720 1842.800 2253.980 2098.160 ;
        RECT 2256.380 1842.800 2262.640 2098.160 ;
        RECT 2265.040 1842.800 2271.300 2098.160 ;
        RECT 2273.700 1842.800 2279.960 2098.160 ;
        RECT 2282.360 1842.800 2288.620 2098.160 ;
        RECT 2291.020 1842.800 2297.280 2098.160 ;
        RECT 2299.680 1842.800 2305.940 2098.160 ;
        RECT 2308.340 1842.800 2315.320 2098.160 ;
        RECT 2237.645 1821.580 2315.320 1842.800 ;
        RECT 2238.340 1002.800 2245.320 1821.580 ;
        RECT 2247.720 1002.800 2253.980 1821.580 ;
        RECT 2256.380 1002.800 2262.640 1821.580 ;
        RECT 2265.040 1002.800 2271.300 1821.580 ;
        RECT 2273.700 1002.800 2279.960 1821.580 ;
        RECT 2282.360 1002.800 2288.620 1821.580 ;
        RECT 2291.020 1002.800 2297.280 1821.580 ;
        RECT 2299.680 1002.800 2305.940 1821.580 ;
        RECT 2308.340 1002.800 2315.320 1821.580 ;
        RECT 2237.645 991.780 2315.320 1002.800 ;
        RECT 2317.720 991.780 2323.980 2098.160 ;
        RECT 2326.380 991.780 2332.640 2098.160 ;
        RECT 2335.040 991.780 2341.300 2098.160 ;
        RECT 2343.700 991.780 2349.960 2098.160 ;
        RECT 2352.360 991.780 2358.620 2098.160 ;
        RECT 2361.020 991.780 2367.280 2098.160 ;
        RECT 2369.680 991.780 2375.940 2098.160 ;
        RECT 2378.340 991.780 2385.320 2098.160 ;
        RECT 2387.720 991.780 2393.980 2098.160 ;
        RECT 2396.380 991.780 2402.640 2098.160 ;
        RECT 2405.040 991.780 2411.300 2098.160 ;
        RECT 2413.700 991.780 2419.960 2098.160 ;
        RECT 2422.360 991.780 2428.620 2098.160 ;
        RECT 2431.020 991.780 2437.280 2098.160 ;
        RECT 2439.680 991.780 2445.940 2098.160 ;
        RECT 2448.340 991.780 2455.320 2098.160 ;
        RECT 2457.720 991.780 2463.980 2098.160 ;
        RECT 2466.380 991.780 2472.640 2098.160 ;
        RECT 2475.040 991.780 2481.300 2098.160 ;
        RECT 2483.700 991.780 2489.960 2098.160 ;
        RECT 2492.360 991.780 2498.620 2098.160 ;
        RECT 2501.020 991.780 2507.280 2098.160 ;
        RECT 2509.680 991.780 2515.940 2098.160 ;
        RECT 2518.340 991.780 2525.320 2098.160 ;
        RECT 2527.720 991.780 2533.980 2098.160 ;
        RECT 2536.380 991.780 2542.640 2098.160 ;
        RECT 2545.040 991.780 2551.300 2098.160 ;
        RECT 2553.700 991.780 2559.960 2098.160 ;
        RECT 2562.360 991.780 2568.620 2098.160 ;
        RECT 2571.020 991.780 2577.280 2098.160 ;
        RECT 2579.680 991.780 2585.940 2098.160 ;
        RECT 2588.340 991.780 2595.320 2098.160 ;
        RECT 2597.720 2000.440 2634.960 2098.160 ;
        RECT 2597.720 1908.360 2612.640 2000.440 ;
        RECT 2615.040 1908.360 2621.300 2000.440 ;
        RECT 2623.700 1908.360 2629.960 2000.440 ;
        RECT 2632.360 1908.360 2634.960 2000.440 ;
        RECT 2597.720 1800.440 2634.960 1908.360 ;
        RECT 2597.720 1708.360 2629.960 1800.440 ;
        RECT 2632.360 1708.360 2634.960 1800.440 ;
        RECT 2597.720 1200.440 2634.960 1708.360 ;
        RECT 2597.720 991.780 2603.980 1200.440 ;
        RECT 2606.380 991.780 2612.640 1200.440 ;
        RECT 2615.040 991.780 2621.300 1200.440 ;
        RECT 2623.700 991.780 2629.960 1200.440 ;
        RECT 2632.360 991.780 2634.960 1200.440 ;
  END
END user_project_wrapper
END LIBRARY

