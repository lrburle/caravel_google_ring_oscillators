magic
tech sky130A
magscale 1 2
timestamp 1712684334
<< nwell >>
rect 3003 1748 3202 1803
rect 3565 1748 3699 1749
rect 6979 1748 7136 1749
rect 10422 1748 10606 1749
rect 13867 1748 14021 1749
rect 17309 1748 17464 1749
rect 3003 1405 4282 1748
rect 3003 1283 4300 1405
rect 3003 1085 4325 1283
rect 3003 742 4282 1085
rect 5870 744 7693 1748
rect 9314 1406 11137 1748
rect 9255 1086 11187 1406
rect 9314 744 11137 1086
rect 12758 744 14581 1748
rect 16202 744 18025 1748
rect 19646 744 20785 1748
rect 6974 743 7017 744
rect 10420 743 10456 744
rect 13866 743 13896 744
rect 17299 743 17376 744
<< ndiff >>
rect 6899 441 6934 475
rect 10343 441 10378 475
rect 13787 441 13822 475
rect 17231 441 17266 475
rect 20675 441 20710 475
<< pdiff >>
rect 3050 1647 3084 1681
rect 3733 1646 3767 1680
rect 7177 1646 7211 1680
rect 10621 1646 10655 1680
rect 14065 1646 14099 1680
rect 17509 1646 17543 1680
<< locali >>
rect 0 2172 20785 2492
rect 3411 1405 3445 1475
rect 3 1283 4300 1405
rect 3 1085 4325 1283
rect 6973 1085 7011 1089
rect 9255 1086 11187 1406
rect 10417 1085 10456 1086
rect 13862 1085 13899 1087
rect 17306 1085 17344 1088
rect 3 0 20785 320
<< viali >>
rect 3050 1647 3084 1681
rect 6899 441 6934 475
rect 10343 441 10378 475
rect 13787 441 13822 475
rect 17231 441 17266 475
rect 20675 441 20710 475
<< metal1 >>
rect 0 2172 20785 2492
rect 20706 1982 20711 2014
rect 20670 1975 20735 1982
rect 20670 1923 20677 1975
rect 20729 1923 20735 1975
rect 3307 1862 3313 1918
rect 3369 1862 3375 1918
rect 20670 1917 20735 1923
rect 6901 1847 6966 1854
rect 6901 1795 6908 1847
rect 6960 1795 6966 1847
rect 6901 1789 6966 1795
rect 10345 1847 10410 1854
rect 10345 1795 10352 1847
rect 10404 1795 10410 1847
rect 10345 1789 10410 1795
rect 13789 1847 13854 1854
rect 13789 1795 13796 1847
rect 13848 1795 13854 1847
rect 13789 1789 13854 1795
rect 17233 1847 17298 1854
rect 17233 1795 17240 1847
rect 17292 1795 17298 1847
rect 17233 1789 17298 1795
rect 3232 1714 3238 1770
rect 3294 1714 3300 1770
rect 3039 1681 3097 1686
rect 3039 1647 3050 1681
rect 3084 1647 3097 1681
rect 3039 1640 3097 1647
rect 3 1283 4300 1405
rect 3 1085 4325 1283
rect 6973 1085 7011 1089
rect 9255 1086 11187 1406
rect 10417 1085 10456 1086
rect 13862 1085 13899 1087
rect 17306 1085 17344 1088
rect 3 0 20785 320
<< via1 >>
rect 20677 1923 20729 1975
rect 3313 1862 3369 1918
rect 6908 1795 6960 1847
rect 10352 1795 10404 1847
rect 13796 1795 13848 1847
rect 17240 1795 17292 1847
rect 3238 1714 3294 1770
rect 3719 1637 3775 1693
rect 7163 1637 7219 1693
rect 10607 1637 10663 1693
rect 14051 1637 14107 1693
rect 17495 1637 17551 1693
rect 6888 985 6946 1043
rect 10332 985 10390 1043
rect 13776 985 13834 1043
rect 17220 985 17278 1043
rect 20664 985 20722 1043
<< metal2 >>
rect 3249 2013 20711 2047
rect 3249 1776 3283 2013
rect 20677 1982 20711 2013
rect 20670 1975 20735 1982
rect 3313 1918 3369 1924
rect 20670 1923 20677 1975
rect 20729 1923 20735 1975
rect 20670 1917 20735 1923
rect 3369 1869 3555 1903
rect 3313 1856 3369 1862
rect 3521 1828 3555 1869
rect 6901 1847 6966 1854
rect 3521 1794 4090 1828
rect 6901 1795 6908 1847
rect 6960 1829 6966 1847
rect 10345 1847 10410 1854
rect 6960 1828 7083 1829
rect 6960 1795 7527 1828
rect 6901 1789 6966 1795
rect 7083 1794 7527 1795
rect 10345 1795 10352 1847
rect 10404 1829 10410 1847
rect 13789 1847 13854 1854
rect 10404 1828 10530 1829
rect 10404 1795 11029 1828
rect 10345 1789 10410 1795
rect 10735 1794 11029 1795
rect 13789 1795 13796 1847
rect 13848 1829 13854 1847
rect 17233 1847 17298 1854
rect 13848 1828 13978 1829
rect 13848 1795 14471 1828
rect 13789 1789 13854 1795
rect 13978 1794 14471 1795
rect 17233 1795 17240 1847
rect 17292 1829 17298 1847
rect 17292 1828 17431 1829
rect 17292 1795 17915 1828
rect 17233 1789 17298 1795
rect 17431 1794 17915 1795
rect 3238 1770 3294 1776
rect 3238 1708 3294 1714
<< via2 >>
rect 3719 1637 3775 1693
rect 7163 1637 7219 1693
rect 10607 1637 10663 1693
rect 14051 1637 14107 1693
rect 17495 1637 17551 1693
rect 6888 985 6946 1043
rect 10332 985 10390 1043
rect 13776 985 13834 1043
rect 17220 985 17278 1043
rect 20664 985 20722 1043
<< metal3 >>
rect 3714 1693 3780 2489
rect 7158 1693 7224 2489
rect 10602 1693 10668 2489
rect 14046 1693 14112 2489
rect 17490 1693 17556 2489
rect 6879 0 6955 985
rect 10323 0 10399 985
rect 13767 0 13843 985
rect 17211 0 17287 985
rect 20655 0 20731 985
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_0
timestamp 1710278372
transform 1 0 3014 0 -1 2233
box -10 0 552 902
use sky130_osu_single_mpr2ct_8_b0r1  sky130_osu_single_mpr2ct_8_b0r1_0
timestamp 1712684334
transform 1 0 19498 0 1 259
box -2159 -259 1287 2233
use sky130_osu_single_mpr2ct_8_b0r1  sky130_osu_single_mpr2ct_8_b0r1_1
timestamp 1712684334
transform 1 0 5722 0 1 259
box -2159 -259 1287 2233
use sky130_osu_single_mpr2ct_8_b0r1  sky130_osu_single_mpr2ct_8_b0r1_2
timestamp 1712684334
transform 1 0 9166 0 1 259
box -2159 -259 1287 2233
use sky130_osu_single_mpr2ct_8_b0r1  sky130_osu_single_mpr2ct_8_b0r1_3
timestamp 1712684334
transform 1 0 12610 0 1 259
box -2159 -259 1287 2233
use sky130_osu_single_mpr2ct_8_b0r1  sky130_osu_single_mpr2ct_8_b0r1_4
timestamp 1712684334
transform 1 0 16054 0 1 259
box -2159 -259 1287 2233
<< labels >>
flabel metal1 s 3039 1640 3097 1686 0 FreeSans 100 0 0 0 start
port 15 nsew signal input
flabel metal1 s 6899 441 6934 475 0 FreeSans 100 0 0 0 X1_Y1
port 10 s signal output
flabel metal1 s 10343 441 10378 475 0 FreeSans 100 0 0 0 X2_Y1
port 9 s signal output
flabel metal1 s 13787 441 13822 475 0 FreeSans 100 0 0 0 X3_Y1
port 8 s signal output
flabel metal1 s 17231 441 17266 475 0 FreeSans 100 0 0 0 X4_Y1
port 7 s signal output
flabel metal1 s 20675 441 20710 475 0 FreeSans 100 0 0 0 X5_Y1
port 6 s signal output
flabel metal1 s 5811 1086 7742 1406 0 FreeSans 100 0 0 0 vccd1
port 17 nsew power bidirectional
flabel metal1 s 9255 1086 11187 1406 0 FreeSans 100 0 0 0 vccd1
port 17 nsew power bidirectional
flabel metal1 s 12699 1086 14631 1406 0 FreeSans 100 0 0 0 vccd1
port 17 nsew power bidirectional
flabel metal1 s 16143 1086 18075 1406 0 FreeSans 100 0 0 0 vccd1
port 17 nsew power bidirectional
flabel metal1 s 19587 1086 20785 1406 0 FreeSans 100 0 0 0 vccd1
port 17 nsew power bidirectional
flabel metal1 s 0 2172 20785 2492 0 FreeSans 100 0 0 0 vssd1
port 16 nsew ground bidirectional
flabel metal1 s 3 1085 4300 1405 0 FreeSans 100 0 0 0 vccd1
port 17 nsew power bidirectional
flabel metal1 s 3 0 20785 320 0 FreeSans 100 0 0 0 vssd1
port 16 nsew ground bidirectional
flabel metal1 s 3732 1647 3766 1681 0 FreeSans 100 0 0 0 s1
port 1 n signal input
flabel metal1 s 7176 1647 7210 1681 0 FreeSans 100 0 0 0 s2
port 2 n signal input
flabel metal1 s 10620 1647 10654 1681 0 FreeSans 100 0 0 0 s3
port 3 n signal input
flabel metal1 s 14064 1647 14098 1681 0 FreeSans 100 0 0 0 s4
port 14 n signal input
flabel metal1 s 17508 1647 17542 1681 0 FreeSans 100 0 0 0 s5
port 13 n signal input
<< end >>
