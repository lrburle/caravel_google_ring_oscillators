magic
tech sky130A
magscale 1 2
timestamp 1714076846
<< nwell >>
rect -58 260 1418 826
<< pwell >>
rect -32 1066 106 1148
rect 488 1098 522 1104
rect 1132 1098 1166 1104
rect 488 1066 604 1098
rect 1132 1076 1258 1098
rect 1132 1066 1194 1076
rect -32 1028 1194 1066
rect 132 902 1194 1028
rect 132 884 322 902
rect 644 884 1194 902
rect -20 162 186 202
rect 452 162 642 202
rect -20 157 642 162
rect 918 157 1374 202
rect -20 60 1374 157
rect -32 26 1374 60
rect -32 -60 86 26
rect 456 21 1374 26
rect 672 -16 706 20
rect 1134 18 1168 20
rect 1132 16 1168 18
rect 1134 -16 1168 16
<< nmos >>
rect 58 92 88 176
<< scnmos >>
rect 214 910 244 1040
rect 322 928 352 1012
rect 406 928 436 1012
rect 742 910 772 1040
rect 814 910 844 1040
rect 1010 910 1040 1040
rect 1086 910 1116 1040
rect 266 52 296 136
rect 338 52 368 136
rect 418 52 448 136
rect 534 46 564 176
rect 722 46 752 130
rect 794 46 824 130
rect 866 46 896 130
rect 994 46 1024 176
rect 1182 46 1212 176
rect 1266 46 1296 176
<< scpmoshvt >>
rect 214 590 244 790
rect 730 590 760 790
rect 814 590 844 790
rect 1002 590 1032 790
rect 1086 590 1116 790
rect 260 310 290 394
rect 344 310 374 394
rect 440 296 470 380
rect 534 296 564 496
rect 722 300 752 384
rect 806 300 836 384
rect 900 300 930 384
rect 994 296 1024 496
rect 1182 296 1212 496
rect 1254 296 1284 496
<< pmoshvt >>
rect 322 590 352 674
rect 408 590 438 674
rect 58 412 88 496
<< ndiff >>
rect 158 1028 214 1040
rect 158 994 170 1028
rect 204 994 214 1028
rect 158 910 214 994
rect 244 1028 296 1040
rect 244 994 254 1028
rect 288 1012 296 1028
rect 670 1024 742 1040
rect 288 994 322 1012
rect 244 928 322 994
rect 352 928 406 1012
rect 436 998 492 1012
rect 436 964 446 998
rect 480 964 492 998
rect 436 928 492 964
rect 670 990 684 1024
rect 718 990 742 1024
rect 244 910 296 928
rect 670 910 742 990
rect 772 910 814 1040
rect 844 1020 896 1040
rect 844 986 854 1020
rect 888 986 896 1020
rect 844 910 896 986
rect 958 1020 1010 1040
rect 958 986 966 1020
rect 1000 986 1010 1020
rect 958 910 1010 986
rect 1040 910 1086 1040
rect 1116 1002 1168 1040
rect 1116 968 1126 1002
rect 1160 968 1168 1002
rect 1116 910 1168 968
rect 5 162 58 176
rect 5 128 13 162
rect 47 128 58 162
rect 5 92 58 128
rect 88 164 141 176
rect 88 130 99 164
rect 133 130 141 164
rect 478 136 534 176
rect 88 120 141 130
rect 88 92 139 120
rect 216 110 266 136
rect 214 98 266 110
rect 214 64 222 98
rect 256 64 266 98
rect 214 52 266 64
rect 296 52 338 136
rect 368 52 418 136
rect 448 108 534 136
rect 448 74 490 108
rect 524 74 534 108
rect 448 52 534 74
rect 482 46 534 52
rect 564 118 616 176
rect 944 130 994 176
rect 564 84 574 118
rect 608 84 616 118
rect 564 46 616 84
rect 670 92 722 130
rect 670 58 678 92
rect 712 58 722 92
rect 670 46 722 58
rect 752 46 794 130
rect 824 46 866 130
rect 896 108 994 130
rect 896 74 950 108
rect 984 74 994 108
rect 896 46 994 74
rect 1024 118 1076 176
rect 1024 84 1034 118
rect 1068 84 1076 118
rect 1024 46 1076 84
rect 1130 162 1182 176
rect 1130 128 1138 162
rect 1172 128 1182 162
rect 1130 94 1182 128
rect 1130 60 1138 94
rect 1172 60 1182 94
rect 1130 46 1182 60
rect 1212 162 1266 176
rect 1212 128 1222 162
rect 1256 128 1266 162
rect 1212 94 1266 128
rect 1212 60 1222 94
rect 1256 60 1266 94
rect 1212 46 1266 60
rect 1296 162 1348 176
rect 1296 128 1306 162
rect 1340 128 1348 162
rect 1296 94 1348 128
rect 1296 60 1306 94
rect 1340 60 1348 94
rect 1296 46 1348 60
<< pdiff >>
rect 120 704 214 790
rect 120 670 150 704
rect 184 670 214 704
rect 120 636 214 670
rect 120 602 150 636
rect 184 602 214 636
rect 120 590 214 602
rect 244 704 306 790
rect 244 670 254 704
rect 288 674 306 704
rect 670 700 730 790
rect 288 670 322 674
rect 244 636 322 670
rect 244 602 254 636
rect 288 602 322 636
rect 244 590 322 602
rect 352 644 408 674
rect 352 610 363 644
rect 397 610 408 644
rect 352 590 408 610
rect 438 636 495 674
rect 438 602 449 636
rect 483 602 495 636
rect 438 590 495 602
rect 670 666 686 700
rect 720 666 730 700
rect 670 632 730 666
rect 670 598 686 632
rect 720 598 730 632
rect 670 590 730 598
rect 760 704 814 790
rect 760 670 770 704
rect 804 670 814 704
rect 760 590 814 670
rect 844 636 896 790
rect 844 602 854 636
rect 888 602 896 636
rect 844 590 896 602
rect 950 636 1002 790
rect 950 602 958 636
rect 992 602 1002 636
rect 950 590 1002 602
rect 1032 712 1086 790
rect 1032 678 1042 712
rect 1076 678 1086 712
rect 1032 590 1086 678
rect 1116 772 1168 790
rect 1116 738 1126 772
rect 1160 738 1168 772
rect 1116 704 1168 738
rect 1116 670 1126 704
rect 1160 670 1168 704
rect 1116 636 1168 670
rect 1116 602 1126 636
rect 1160 602 1168 636
rect 1116 590 1168 602
rect 5 474 58 496
rect 5 440 13 474
rect 47 440 58 474
rect 5 412 58 440
rect 88 468 141 496
rect 88 434 99 468
rect 133 434 141 468
rect 88 422 141 434
rect 482 484 534 496
rect 482 450 490 484
rect 524 450 534 484
rect 482 438 534 450
rect 88 412 138 422
rect 210 380 260 394
rect 208 368 260 380
rect 208 334 216 368
rect 250 334 260 368
rect 208 310 260 334
rect 290 386 344 394
rect 290 352 300 386
rect 334 352 344 386
rect 290 310 344 352
rect 374 380 424 394
rect 485 380 534 438
rect 374 362 440 380
rect 374 328 394 362
rect 428 328 440 362
rect 374 310 440 328
rect 390 296 440 310
rect 470 296 534 380
rect 564 470 616 496
rect 564 436 574 470
rect 608 436 616 470
rect 564 402 616 436
rect 942 484 994 496
rect 942 450 950 484
rect 984 450 994 484
rect 942 438 994 450
rect 564 368 574 402
rect 608 368 616 402
rect 945 384 994 438
rect 564 296 616 368
rect 670 346 722 384
rect 670 312 678 346
rect 712 312 722 346
rect 670 300 722 312
rect 752 376 806 384
rect 752 342 762 376
rect 796 342 806 376
rect 752 300 806 342
rect 836 356 900 384
rect 836 322 856 356
rect 890 322 900 356
rect 836 300 900 322
rect 930 300 994 384
rect 945 296 994 300
rect 1024 470 1076 496
rect 1024 436 1034 470
rect 1068 436 1076 470
rect 1024 402 1076 436
rect 1024 368 1034 402
rect 1068 368 1076 402
rect 1024 296 1076 368
rect 1130 484 1182 496
rect 1130 450 1138 484
rect 1172 450 1182 484
rect 1130 416 1182 450
rect 1130 382 1138 416
rect 1172 382 1182 416
rect 1130 348 1182 382
rect 1130 314 1138 348
rect 1172 314 1182 348
rect 1130 296 1182 314
rect 1212 296 1254 496
rect 1284 484 1336 496
rect 1284 450 1294 484
rect 1328 450 1336 484
rect 1284 416 1336 450
rect 1284 382 1294 416
rect 1328 382 1336 416
rect 1284 348 1336 382
rect 1284 314 1294 348
rect 1328 314 1336 348
rect 1284 296 1336 314
<< ndiffc >>
rect 170 994 204 1028
rect 254 994 288 1028
rect 446 964 480 998
rect 684 990 718 1024
rect 854 986 888 1020
rect 966 986 1000 1020
rect 1126 968 1160 1002
rect 13 128 47 162
rect 99 130 133 164
rect 222 64 256 98
rect 490 74 524 108
rect 574 84 608 118
rect 678 58 712 92
rect 950 74 984 108
rect 1034 84 1068 118
rect 1138 128 1172 162
rect 1138 60 1172 94
rect 1222 128 1256 162
rect 1222 60 1256 94
rect 1306 128 1340 162
rect 1306 60 1340 94
<< pdiffc >>
rect 150 670 184 704
rect 150 602 184 636
rect 254 670 288 704
rect 254 602 288 636
rect 363 610 397 644
rect 449 602 483 636
rect 686 666 720 700
rect 686 598 720 632
rect 770 670 804 704
rect 854 602 888 636
rect 958 602 992 636
rect 1042 678 1076 712
rect 1126 738 1160 772
rect 1126 670 1160 704
rect 1126 602 1160 636
rect 13 440 47 474
rect 99 434 133 468
rect 490 450 524 484
rect 216 334 250 368
rect 300 352 334 386
rect 394 328 428 362
rect 574 436 608 470
rect 950 450 984 484
rect 574 368 608 402
rect 678 312 712 346
rect 762 342 796 376
rect 856 322 890 356
rect 1034 436 1068 470
rect 1034 368 1068 402
rect 1138 450 1172 484
rect 1138 382 1172 416
rect 1138 314 1172 348
rect 1294 450 1328 484
rect 1294 382 1328 416
rect 1294 314 1328 348
<< poly >>
rect 214 1040 244 1066
rect 742 1040 772 1066
rect 814 1040 844 1066
rect 1010 1040 1040 1066
rect 1086 1040 1116 1066
rect 322 1012 352 1038
rect 406 1012 436 1038
rect 214 888 244 910
rect 322 888 352 928
rect 178 872 244 888
rect 178 838 194 872
rect 228 838 244 872
rect 178 822 244 838
rect 286 872 352 888
rect 286 838 302 872
rect 336 838 352 872
rect 286 822 352 838
rect 406 888 436 928
rect 742 888 772 910
rect 406 872 494 888
rect 406 838 444 872
rect 478 838 494 872
rect 406 823 494 838
rect 407 822 494 823
rect 718 872 772 888
rect 718 838 728 872
rect 762 838 772 872
rect 718 822 772 838
rect 814 888 844 910
rect 1010 888 1040 910
rect 814 872 892 888
rect 814 838 844 872
rect 878 838 892 872
rect 814 822 892 838
rect 982 872 1040 888
rect 982 838 992 872
rect 1026 838 1040 872
rect 982 822 1040 838
rect 1086 888 1116 910
rect 1086 872 1140 888
rect 1086 838 1096 872
rect 1130 838 1140 872
rect 1086 822 1140 838
rect 214 790 244 822
rect 322 674 352 822
rect 408 674 438 822
rect 730 790 760 822
rect 814 790 844 822
rect 1002 790 1032 822
rect 1086 790 1116 822
rect 214 564 244 590
rect 322 564 352 590
rect 408 564 438 590
rect 730 564 760 590
rect 814 564 844 590
rect 1002 564 1032 590
rect 1086 564 1116 590
rect 58 496 88 522
rect 344 476 402 500
rect 534 496 564 522
rect 994 496 1024 522
rect 1182 496 1212 522
rect 1254 496 1284 522
rect 344 442 358 476
rect 392 442 402 476
rect 344 426 402 442
rect 58 338 88 412
rect 260 394 290 424
rect 344 394 374 426
rect 2 322 88 338
rect 2 288 14 322
rect 48 288 88 322
rect 440 380 470 406
rect 2 248 88 288
rect 260 264 290 310
rect 2 214 14 248
rect 48 214 88 248
rect 2 198 88 214
rect 212 248 296 264
rect 212 214 222 248
rect 256 214 296 248
rect 344 240 374 310
rect 806 476 860 492
rect 806 442 816 476
rect 850 442 860 476
rect 806 426 860 442
rect 722 384 752 424
rect 806 384 836 426
rect 900 384 930 410
rect 440 264 470 296
rect 534 264 564 296
rect 212 198 296 214
rect 58 176 88 198
rect 266 136 296 198
rect 338 202 374 240
rect 418 248 472 264
rect 418 214 428 248
rect 462 214 472 248
rect 338 136 368 202
rect 418 198 472 214
rect 514 248 568 264
rect 722 250 752 300
rect 806 282 836 300
rect 514 214 524 248
rect 558 214 568 248
rect 514 198 568 214
rect 668 202 752 250
rect 418 136 448 198
rect 534 176 564 198
rect 58 66 88 92
rect 266 26 296 52
rect 338 26 368 52
rect 418 26 448 52
rect 668 168 678 202
rect 712 168 752 202
rect 668 146 752 168
rect 722 130 752 146
rect 794 256 836 282
rect 900 258 930 300
rect 994 264 1024 296
rect 1182 264 1212 296
rect 794 130 824 256
rect 878 242 932 258
rect 878 226 888 242
rect 866 208 888 226
rect 922 208 932 242
rect 866 192 932 208
rect 974 248 1028 264
rect 974 214 984 248
rect 1018 214 1028 248
rect 974 198 1028 214
rect 1126 248 1212 264
rect 1126 214 1140 248
rect 1174 214 1212 248
rect 1254 264 1284 296
rect 1254 248 1358 264
rect 1254 234 1308 248
rect 1126 198 1212 214
rect 866 170 908 192
rect 994 176 1024 198
rect 1182 176 1212 198
rect 1266 214 1308 234
rect 1342 214 1358 248
rect 1266 198 1358 214
rect 1266 176 1296 198
rect 866 146 904 170
rect 866 130 896 146
rect 534 20 564 46
rect 722 20 752 46
rect 794 20 824 46
rect 866 20 896 46
rect 994 20 1024 46
rect 1182 20 1212 46
rect 1266 20 1296 46
<< polycont >>
rect 194 838 228 872
rect 302 838 336 872
rect 444 838 478 872
rect 728 838 762 872
rect 844 838 878 872
rect 992 838 1026 872
rect 1096 838 1130 872
rect 358 442 392 476
rect 14 288 48 322
rect 14 214 48 248
rect 222 214 256 248
rect 816 442 850 476
rect 428 214 462 248
rect 524 214 558 248
rect 678 168 712 202
rect 888 208 922 242
rect 984 214 1018 248
rect 1140 214 1174 248
rect 1308 214 1342 248
<< locali >>
rect -20 1070 8 1104
rect 42 1070 120 1104
rect 154 1070 212 1104
rect 246 1070 304 1104
rect 338 1070 396 1104
rect 430 1070 488 1104
rect 522 1070 580 1104
rect 614 1070 672 1104
rect 706 1070 764 1104
rect 798 1070 856 1104
rect 890 1070 948 1104
rect 982 1070 1040 1104
rect 1074 1070 1132 1104
rect 1166 1070 1224 1104
rect 1258 1070 1316 1104
rect 1350 1070 1380 1104
rect 108 1028 220 1036
rect 108 994 170 1028
rect 204 994 220 1028
rect 108 978 220 994
rect 254 1028 304 1070
rect 288 994 304 1028
rect 668 1024 734 1070
rect 254 978 304 994
rect 428 1010 480 1016
rect 428 998 494 1010
rect 108 704 158 978
rect 428 964 446 998
rect 480 964 494 998
rect 668 990 684 1024
rect 718 990 734 1024
rect 770 1020 1032 1036
rect 428 944 494 964
rect 770 986 854 1020
rect 888 986 966 1020
rect 1000 986 1032 1020
rect 1086 1002 1176 1070
rect 770 956 806 986
rect 1086 968 1126 1002
rect 1160 968 1176 1002
rect 216 906 494 944
rect 660 922 806 956
rect 216 888 250 906
rect 192 872 250 888
rect 192 838 194 872
rect 228 838 250 872
rect 192 822 250 838
rect 284 866 302 872
rect 284 832 288 866
rect 336 838 352 872
rect 322 832 352 838
rect 284 822 352 832
rect 396 838 444 872
rect 478 866 532 872
rect 478 838 492 866
rect 396 832 492 838
rect 526 832 532 866
rect 396 822 532 832
rect 216 772 250 822
rect 216 738 405 772
rect 478 750 532 822
rect 660 788 694 922
rect 728 872 794 888
rect 856 872 898 952
rect 762 866 794 872
rect 728 832 730 838
rect 764 832 794 866
rect 828 866 844 872
rect 828 832 832 866
rect 878 838 898 872
rect 866 832 898 838
rect 948 872 998 952
rect 1080 872 1170 934
rect 948 866 992 872
rect 948 832 968 866
rect 1026 838 1042 872
rect 1002 832 1042 838
rect 1080 838 1096 872
rect 1130 866 1170 872
rect 1080 832 1104 838
rect 1138 832 1170 866
rect 728 822 794 832
rect 828 788 1176 798
rect 660 772 1176 788
rect 660 762 1126 772
rect 660 754 872 762
rect 108 670 150 704
rect 184 670 200 704
rect 108 662 200 670
rect 108 636 152 662
rect 108 602 150 636
rect 186 628 200 662
rect 184 602 200 628
rect 108 594 200 602
rect 238 670 254 704
rect 288 670 304 704
rect 238 636 304 670
rect 238 602 254 636
rect 288 602 304 636
rect 238 560 304 602
rect 344 644 405 738
rect 1110 738 1126 762
rect 1160 738 1176 772
rect 900 720 1076 728
rect 670 700 724 716
rect 670 666 686 700
rect 720 666 724 700
rect 344 610 363 644
rect 397 610 405 644
rect 344 594 405 610
rect 441 636 497 652
rect 441 602 449 636
rect 483 602 497 636
rect 441 560 497 602
rect 670 632 724 666
rect 770 712 1076 720
rect 770 704 1042 712
rect 804 680 1042 704
rect 954 678 1042 680
rect 954 670 1076 678
rect 770 654 804 670
rect 1030 662 1076 670
rect 1110 704 1176 738
rect 1110 670 1126 704
rect 1160 670 1176 704
rect 1110 662 1176 670
rect 1110 636 1240 662
rect 670 598 686 632
rect 720 598 724 632
rect 670 560 724 598
rect 834 602 854 636
rect 888 602 908 636
rect 834 560 908 602
rect 942 602 958 636
rect 992 628 1008 636
rect 1110 628 1126 636
rect 992 602 1126 628
rect 1160 628 1240 636
rect 1160 602 1176 628
rect 942 594 1176 602
rect -20 526 8 560
rect 42 526 100 560
rect 134 526 212 560
rect 246 526 304 560
rect 338 526 396 560
rect 430 526 488 560
rect 522 526 580 560
rect 614 526 672 560
rect 706 526 764 560
rect 798 526 856 560
rect 890 526 948 560
rect 982 526 1040 560
rect 1074 526 1132 560
rect 1166 526 1224 560
rect 1258 526 1316 560
rect 1350 526 1380 560
rect -5 496 48 526
rect -5 474 47 496
rect -5 440 13 474
rect -5 424 47 440
rect 99 468 133 492
rect 99 424 133 434
rect 200 426 324 526
rect 98 412 133 424
rect -4 322 64 390
rect -4 288 14 322
rect 48 288 64 322
rect -4 254 64 288
rect -4 220 -2 254
rect 32 248 64 254
rect -4 214 14 220
rect 48 214 64 248
rect 98 248 132 412
rect 200 368 250 392
rect 200 334 216 368
rect 284 390 324 426
rect 358 476 452 492
rect 392 458 452 476
rect 358 424 390 442
rect 424 424 452 458
rect 486 484 530 526
rect 486 450 490 484
rect 524 450 530 484
rect 486 418 530 450
rect 572 470 626 492
rect 572 436 574 470
rect 608 436 626 470
rect 572 402 626 436
rect 284 386 350 390
rect 284 352 300 386
rect 334 352 350 386
rect 394 362 538 378
rect 200 318 250 334
rect 428 328 538 362
rect 572 368 574 402
rect 608 368 626 402
rect 660 396 782 526
rect 816 476 912 492
rect 850 458 912 476
rect 816 424 832 442
rect 866 424 912 458
rect 946 484 998 526
rect 946 450 950 484
rect 984 450 998 484
rect 946 418 998 450
rect 1032 470 1086 492
rect 1032 436 1034 470
rect 1068 436 1086 470
rect 1032 402 1086 436
rect 572 352 626 368
rect 746 390 784 396
rect 746 376 812 390
rect 394 318 538 328
rect 200 284 558 318
rect 98 214 222 248
rect 256 214 278 248
rect 98 198 278 214
rect 98 180 148 198
rect -4 162 47 180
rect -4 128 13 162
rect -4 70 47 128
rect 88 164 148 180
rect 88 130 99 164
rect 133 130 148 164
rect 88 96 148 130
rect 312 114 362 284
rect 512 248 558 284
rect 204 98 362 114
rect -4 18 48 70
rect 204 64 222 98
rect 256 64 362 98
rect 204 60 362 64
rect 396 214 428 248
rect 462 214 478 248
rect 396 186 478 214
rect 512 214 524 248
rect 512 198 558 214
rect 396 152 424 186
rect 458 152 478 186
rect 396 144 478 152
rect 592 186 626 352
rect 660 346 712 362
rect 660 312 678 346
rect 746 342 762 376
rect 796 342 812 376
rect 846 356 998 376
rect 846 326 856 356
rect 844 322 856 326
rect 890 322 998 356
rect 1032 368 1034 402
rect 1068 368 1086 402
rect 1032 352 1086 368
rect 844 320 998 322
rect 840 318 998 320
rect 840 314 1018 318
rect 836 312 1018 314
rect 660 272 712 312
rect 832 310 1018 312
rect 826 308 1018 310
rect 812 302 1018 308
rect 808 296 1018 302
rect 804 290 1018 296
rect 798 284 1018 290
rect 792 278 1018 284
rect 786 276 1018 278
rect 786 274 858 276
rect 786 272 856 274
rect 660 270 852 272
rect 660 268 850 270
rect 660 264 846 268
rect 660 262 844 264
rect 660 238 838 262
rect 972 248 1018 276
rect 592 146 626 152
rect 396 60 436 144
rect 574 118 626 146
rect 660 202 770 204
rect 660 168 678 202
rect 712 186 770 202
rect 660 152 696 168
rect 730 152 770 186
rect 660 126 770 152
rect 474 74 490 108
rect 524 74 540 108
rect 474 18 540 74
rect 608 84 626 118
rect 804 92 838 238
rect 574 52 626 84
rect 660 58 678 92
rect 712 58 838 92
rect 872 208 888 242
rect 922 208 938 242
rect 872 158 938 208
rect 972 214 984 248
rect 972 198 1018 214
rect 1052 254 1086 352
rect 1122 484 1188 490
rect 1122 450 1138 484
rect 1172 450 1188 484
rect 1122 416 1188 450
rect 1122 382 1138 416
rect 1172 382 1188 416
rect 1122 348 1188 382
rect 1122 314 1138 348
rect 1172 332 1188 348
rect 1294 484 1360 526
rect 1328 450 1360 484
rect 1294 416 1360 450
rect 1328 382 1360 416
rect 1294 348 1360 382
rect 1172 322 1258 332
rect 1172 314 1224 322
rect 1122 298 1224 314
rect 1328 314 1360 348
rect 1294 298 1360 314
rect 1120 254 1190 264
rect 1052 248 1190 254
rect 1052 220 1140 248
rect 872 120 916 158
rect 1052 146 1086 220
rect 1120 214 1140 220
rect 1174 214 1190 248
rect 1224 178 1258 288
rect 1292 254 1362 264
rect 1292 214 1308 254
rect 1342 214 1362 254
rect 872 86 878 120
rect 912 86 916 120
rect 872 60 916 86
rect 950 108 1000 124
rect 984 74 1000 108
rect 950 18 1000 74
rect 1034 122 1086 146
rect 1034 118 1036 122
rect 1070 88 1086 122
rect 1068 84 1086 88
rect 1034 52 1086 84
rect 1124 162 1172 178
rect 1124 128 1138 162
rect 1124 94 1172 128
rect 1124 60 1138 94
rect 1124 18 1172 60
rect 1206 162 1272 178
rect 1206 128 1222 162
rect 1256 128 1272 162
rect 1206 94 1272 128
rect 1206 60 1222 94
rect 1256 60 1272 94
rect 1206 52 1272 60
rect 1306 162 1360 178
rect 1340 128 1360 162
rect 1306 94 1360 128
rect 1340 60 1360 94
rect 1306 18 1360 60
rect -20 -16 8 18
rect 42 -16 100 18
rect 134 -16 212 18
rect 246 -16 304 18
rect 338 -16 396 18
rect 430 -16 488 18
rect 522 -16 580 18
rect 614 -16 672 18
rect 706 -16 764 18
rect 798 -16 856 18
rect 890 -16 948 18
rect 982 -16 1040 18
rect 1074 -16 1132 18
rect 1166 -16 1224 18
rect 1258 -16 1316 18
rect 1350 -16 1380 18
<< viali >>
rect 8 1070 42 1104
rect 120 1070 154 1104
rect 212 1070 246 1104
rect 304 1070 338 1104
rect 396 1070 430 1104
rect 488 1070 522 1104
rect 580 1070 614 1104
rect 672 1070 706 1104
rect 764 1070 798 1104
rect 856 1070 890 1104
rect 948 1070 982 1104
rect 1040 1070 1074 1104
rect 1132 1070 1166 1104
rect 1224 1070 1258 1104
rect 1316 1070 1350 1104
rect 288 838 302 866
rect 302 838 322 866
rect 288 832 322 838
rect 492 832 526 866
rect 730 838 762 866
rect 762 838 764 866
rect 730 832 764 838
rect 832 838 844 866
rect 844 838 866 866
rect 832 832 866 838
rect 968 838 992 866
rect 992 838 1002 866
rect 968 832 1002 838
rect 1104 838 1130 866
rect 1130 838 1138 866
rect 1104 832 1138 838
rect 152 636 186 662
rect 152 628 184 636
rect 184 628 186 636
rect 1240 628 1274 662
rect 8 526 42 560
rect 100 526 134 560
rect 212 526 246 560
rect 304 526 338 560
rect 396 526 430 560
rect 488 526 522 560
rect 580 526 614 560
rect 672 526 706 560
rect 764 526 798 560
rect 856 526 890 560
rect 948 526 982 560
rect 1040 526 1074 560
rect 1132 526 1166 560
rect 1224 526 1258 560
rect 1316 526 1350 560
rect -2 248 32 254
rect -2 220 14 248
rect 14 220 32 248
rect 390 442 392 458
rect 392 442 424 458
rect 390 424 424 442
rect 832 442 850 458
rect 850 442 866 458
rect 832 424 866 442
rect 424 152 458 186
rect 592 152 626 186
rect 696 168 712 186
rect 712 168 730 186
rect 696 152 730 168
rect 1224 288 1258 322
rect 1308 248 1342 254
rect 1308 220 1342 248
rect 878 86 912 120
rect 1036 118 1070 122
rect 1036 88 1068 118
rect 1068 88 1070 118
rect 8 -16 42 18
rect 100 -16 134 18
rect 212 -16 246 18
rect 304 -16 338 18
rect 396 -16 430 18
rect 488 -16 522 18
rect 580 -16 614 18
rect 672 -16 706 18
rect 764 -16 798 18
rect 856 -16 890 18
rect 948 -16 982 18
rect 1040 -16 1074 18
rect 1132 -16 1166 18
rect 1224 -16 1258 18
rect 1316 -16 1350 18
<< metal1 >>
rect -20 1104 1380 1136
rect -20 1070 8 1104
rect 42 1070 120 1104
rect 154 1070 212 1104
rect 246 1070 304 1104
rect 338 1070 396 1104
rect 430 1070 488 1104
rect 522 1070 580 1104
rect 614 1070 672 1104
rect 706 1070 764 1104
rect 798 1070 856 1104
rect 890 1070 948 1104
rect 982 1070 1040 1104
rect 1074 1070 1132 1104
rect 1166 1070 1224 1104
rect 1258 1070 1316 1104
rect 1350 1070 1380 1104
rect -20 1064 1380 1070
rect 478 1006 564 1008
rect 478 988 484 1006
rect 292 960 484 988
rect 292 872 320 960
rect 480 954 484 960
rect 536 988 564 1006
rect 536 960 762 988
rect 484 948 536 954
rect 276 866 334 872
rect 276 832 288 866
rect 322 832 334 866
rect 276 826 334 832
rect 480 866 538 872
rect 480 832 492 866
rect 526 864 538 866
rect 614 864 620 876
rect 526 836 620 864
rect 526 832 538 836
rect 480 826 538 832
rect 614 824 620 836
rect 672 824 678 876
rect 734 872 762 960
rect 718 866 776 872
rect 718 832 730 866
rect 764 832 776 866
rect 718 826 776 832
rect 818 824 824 876
rect 876 824 882 876
rect 956 866 1014 872
rect 956 832 968 866
rect 1002 832 1014 866
rect 956 826 1014 832
rect 632 796 660 824
rect 972 796 1000 826
rect 1090 824 1096 876
rect 1148 864 1154 876
rect 1148 836 1208 864
rect 1148 824 1154 836
rect 632 768 1000 796
rect 140 662 198 668
rect 140 628 152 662
rect 186 660 198 662
rect 682 660 688 672
rect 186 632 688 660
rect 186 628 198 632
rect 140 622 198 628
rect 682 620 688 632
rect 740 620 746 672
rect 1228 662 1300 672
rect 1228 628 1240 662
rect 1274 628 1300 662
rect 1228 620 1300 628
rect 1352 620 1358 672
rect 322 592 352 593
rect -20 560 1380 592
rect -20 526 8 560
rect 42 526 100 560
rect 134 526 212 560
rect 246 526 304 560
rect 338 526 396 560
rect 430 526 488 560
rect 522 526 580 560
rect 614 526 672 560
rect 706 526 764 560
rect 798 526 856 560
rect 890 526 948 560
rect 982 526 1040 560
rect 1074 526 1132 560
rect 1166 526 1224 560
rect 1258 526 1316 560
rect 1350 526 1380 560
rect -20 496 1380 526
rect 378 458 436 464
rect 378 424 390 458
rect 424 456 436 458
rect 820 458 878 464
rect 820 456 832 458
rect 424 428 832 456
rect 424 424 436 428
rect 378 418 436 424
rect 820 424 832 428
rect 866 456 878 458
rect 954 456 960 468
rect 866 428 960 456
rect 866 424 878 428
rect 820 418 878 424
rect 954 416 960 428
rect 1012 416 1018 468
rect 818 280 824 332
rect 876 320 882 332
rect 1212 322 1270 328
rect 1212 320 1224 322
rect 876 292 1224 320
rect 876 280 882 292
rect 1212 288 1224 292
rect 1258 288 1270 322
rect 1212 282 1270 288
rect -14 254 44 260
rect -14 220 -2 254
rect 32 252 44 254
rect 493 252 667 258
rect 954 252 960 264
rect 32 230 960 252
rect 32 224 521 230
rect 639 224 960 230
rect 32 220 44 224
rect -14 214 44 220
rect 954 212 960 224
rect 1012 212 1018 264
rect 1294 252 1300 264
rect 1238 224 1300 252
rect 1294 212 1300 224
rect 1352 212 1358 264
rect 412 186 470 192
rect 412 152 424 186
rect 458 152 470 186
rect 412 146 470 152
rect 428 106 456 146
rect 546 142 552 194
rect 604 192 610 194
rect 604 186 638 192
rect 626 184 638 186
rect 626 156 642 184
rect 626 152 638 156
rect 604 146 638 152
rect 604 142 610 146
rect 682 144 688 196
rect 740 184 746 196
rect 972 184 1000 212
rect 740 156 800 184
rect 972 156 1068 184
rect 740 144 746 156
rect 892 132 944 138
rect 886 128 892 132
rect 866 120 892 128
rect 866 106 878 120
rect 428 86 878 106
rect 428 80 892 86
rect 944 80 950 132
rect 1040 128 1068 156
rect 1024 122 1082 128
rect 1024 88 1036 122
rect 1070 88 1082 122
rect 1024 82 1082 88
rect 428 78 878 80
rect -20 18 1380 24
rect -20 -16 8 18
rect 42 -16 100 18
rect 134 -16 212 18
rect 246 -16 304 18
rect 338 -16 396 18
rect 430 -16 488 18
rect 522 -16 580 18
rect 614 -16 672 18
rect 706 -16 764 18
rect 798 -16 856 18
rect 890 -16 948 18
rect 982 -16 1040 18
rect 1074 -16 1132 18
rect 1166 -16 1224 18
rect 1258 -16 1316 18
rect 1350 -16 1380 18
rect -20 -48 1380 -16
<< via1 >>
rect 484 954 536 1006
rect 620 824 672 876
rect 824 866 876 876
rect 824 832 832 866
rect 832 832 866 866
rect 866 832 876 866
rect 824 824 876 832
rect 1096 866 1148 876
rect 1096 832 1104 866
rect 1104 832 1138 866
rect 1138 832 1148 866
rect 1096 824 1148 832
rect 688 620 740 672
rect 1300 620 1352 672
rect 960 416 1012 468
rect 824 280 876 332
rect 960 212 1012 264
rect 1300 254 1352 264
rect 1300 220 1308 254
rect 1308 220 1342 254
rect 1342 220 1352 254
rect 1300 212 1352 220
rect 552 186 604 194
rect 552 152 592 186
rect 592 152 604 186
rect 552 142 604 152
rect 688 186 740 196
rect 688 152 696 186
rect 696 152 730 186
rect 730 152 740 186
rect 688 144 740 152
rect 892 120 944 132
rect 892 86 912 120
rect 912 86 944 120
rect 892 80 944 86
<< metal2 >>
rect 480 1008 536 1018
rect 480 942 536 952
rect 614 882 670 887
rect 614 878 672 882
rect 670 876 672 878
rect 670 822 672 824
rect 614 818 672 822
rect 824 878 880 887
rect 1096 876 1148 882
rect 614 812 670 818
rect 824 812 880 822
rect 972 836 1096 864
rect 688 674 744 683
rect 688 608 744 618
rect 552 196 608 206
rect 700 202 728 608
rect 836 456 864 812
rect 972 479 1000 836
rect 1096 818 1148 824
rect 1300 672 1352 678
rect 1300 614 1352 620
rect 960 470 1016 479
rect 836 428 932 456
rect 820 334 876 343
rect 820 268 876 278
rect 552 130 608 140
rect 688 196 740 202
rect 688 138 740 144
rect 904 138 932 428
rect 960 404 1016 414
rect 960 266 1016 275
rect 1312 270 1340 614
rect 960 200 1016 210
rect 1300 264 1352 270
rect 1300 206 1352 212
rect 892 132 944 138
rect 892 70 944 80
<< via2 >>
rect 480 1006 536 1008
rect 480 954 484 1006
rect 484 954 536 1006
rect 480 952 536 954
rect 614 876 670 878
rect 614 824 620 876
rect 620 824 670 876
rect 614 822 670 824
rect 824 876 880 878
rect 824 824 876 876
rect 876 824 880 876
rect 824 822 880 824
rect 688 672 744 674
rect 688 620 740 672
rect 740 620 744 672
rect 688 618 744 620
rect 960 468 1016 470
rect 820 332 876 334
rect 820 280 824 332
rect 824 280 876 332
rect 820 278 876 280
rect 552 194 608 196
rect 552 142 604 194
rect 604 142 608 194
rect 552 140 608 142
rect 960 416 1012 468
rect 1012 416 1016 468
rect 960 414 1016 416
rect 960 264 1016 266
rect 960 212 1012 264
rect 1012 212 1016 264
rect 960 210 1016 212
<< metal3 >>
rect 468 1018 536 1038
rect 468 1016 540 1018
rect 380 1012 540 1016
rect 380 1008 541 1012
rect 380 956 480 1008
rect 472 952 480 956
rect 536 952 541 1008
rect 472 950 541 952
rect 474 944 541 950
rect 608 880 676 883
rect 516 878 676 880
rect 516 822 614 878
rect 670 822 676 878
rect 516 820 676 822
rect 608 814 676 820
rect 816 880 885 883
rect 816 878 978 880
rect 816 822 824 878
rect 880 822 978 878
rect 816 820 978 822
rect 816 816 885 820
rect 816 814 884 816
rect 680 676 749 679
rect 680 674 842 676
rect 680 618 688 674
rect 744 618 842 674
rect 680 616 842 618
rect 680 610 749 616
rect 954 474 1021 476
rect 952 472 1021 474
rect 952 470 1114 472
rect 952 414 960 470
rect 1016 414 1114 470
rect 952 412 1114 414
rect 952 406 1021 412
rect 956 398 1016 406
rect 814 336 882 340
rect 720 334 882 336
rect 720 278 820 334
rect 876 278 882 334
rect 720 276 882 278
rect 814 270 882 276
rect 954 270 1021 271
rect 952 268 1021 270
rect 952 266 1114 268
rect 952 210 960 266
rect 1016 210 1114 266
rect 952 208 1114 210
rect 952 204 1021 208
rect 952 202 1020 204
rect 544 200 613 202
rect 452 196 613 200
rect 452 140 552 196
rect 608 140 613 196
rect 524 138 613 140
rect 544 134 613 138
<< labels >>
rlabel metal3 s 954 204 1020 270 4 R3
port 17 nsew
rlabel metal3 s 814 272 880 338 4 R1
port 19 nsew
rlabel metal3 s 682 612 748 678 4 R0
port 20 nsew
rlabel metal3 s 954 408 1020 474 4 B1
port 16 nsew
rlabel metal3 s 474 952 540 1018 4 B0
port 21 nsew
rlabel metal3 s 818 816 884 882 4 A1
port 13 nsew
rlabel metal3 s 610 816 676 882 4 A0
port 22 nsew
rlabel metal1 s 546 136 612 202 4 R2
port 18 nsew
rlabel metal1 178 2 178 2 1 vgnd
port 23 n
rlabel viali 138 1086 138 1086 1 VNB
port 25 n
rlabel metal1 182 1086 182 1086 1 vgnd
port 23 n
rlabel viali 116 -2 116 -2 1 VNB
port 25 n
rlabel nwell 116 542 116 542 1 VPB
port 26 n
rlabel metal1 156 544 156 544 1 vpwr
port 24 n
<< properties >>
string FIXED_BBOX 0 0 1380 1088
string path 4.925 1.190 5.425 1.190 
<< end >>
