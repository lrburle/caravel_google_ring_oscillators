VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mux16x1_project
  CLASS BLOCK ;
  FOREIGN mux16x1_project ;
  ORIGIN 0.000 0.000 ;
  SIZE 50.000 BY 110.000 ;
  PIN data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 104.760 4.000 105.360 ;
    END
  END data_in[0]
  PIN data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 36.760 4.000 37.360 ;
    END
  END data_in[10]
  PIN data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 29.960 4.000 30.560 ;
    END
  END data_in[11]
  PIN data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.160 4.000 23.760 ;
    END
  END data_in[12]
  PIN data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END data_in[13]
  PIN data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 9.560 4.000 10.160 ;
    END
  END data_in[14]
  PIN data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.760 4.000 3.360 ;
    END
  END data_in[15]
  PIN data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END data_in[1]
  PIN data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END data_in[2]
  PIN data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 84.360 4.000 84.960 ;
    END
  END data_in[3]
  PIN data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END data_in[4]
  PIN data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END data_in[5]
  PIN data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 63.960 4.000 64.560 ;
    END
  END data_in[6]
  PIN data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.160 4.000 57.760 ;
    END
  END data_in[7]
  PIN data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END data_in[8]
  PIN data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END data_in[9]
  PIN select[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 6.070 106.000 6.350 110.000 ;
    END
  END select[0]
  PIN select[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 18.490 106.000 18.770 110.000 ;
    END
  END select[1]
  PIN select[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 30.910 106.000 31.190 110.000 ;
    END
  END select[2]
  PIN select[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 43.330 106.000 43.610 110.000 ;
    END
  END select[3]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.550 10.640 11.150 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 19.210 10.640 20.810 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 28.870 10.640 30.470 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 38.530 10.640 40.130 98.160 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 14.380 10.640 15.980 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 24.040 10.640 25.640 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 33.700 10.640 35.300 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 43.360 10.640 44.960 98.160 ;
    END
  END vssd1
  PIN y
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 46.000 54.440 50.000 55.040 ;
    END
  END y
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 44.160 98.005 ;
      LAYER met1 ;
        RECT 4.670 10.640 44.960 98.160 ;
      LAYER met2 ;
        RECT 4.690 105.720 5.790 106.490 ;
        RECT 6.630 105.720 18.210 106.490 ;
        RECT 19.050 105.720 30.630 106.490 ;
        RECT 31.470 105.720 43.050 106.490 ;
        RECT 43.890 105.720 44.930 106.490 ;
        RECT 4.690 3.555 44.930 105.720 ;
      LAYER met3 ;
        RECT 4.400 104.360 46.000 105.225 ;
        RECT 4.000 98.960 46.000 104.360 ;
        RECT 4.400 97.560 46.000 98.960 ;
        RECT 4.000 92.160 46.000 97.560 ;
        RECT 4.400 90.760 46.000 92.160 ;
        RECT 4.000 85.360 46.000 90.760 ;
        RECT 4.400 83.960 46.000 85.360 ;
        RECT 4.000 78.560 46.000 83.960 ;
        RECT 4.400 77.160 46.000 78.560 ;
        RECT 4.000 71.760 46.000 77.160 ;
        RECT 4.400 70.360 46.000 71.760 ;
        RECT 4.000 64.960 46.000 70.360 ;
        RECT 4.400 63.560 46.000 64.960 ;
        RECT 4.000 58.160 46.000 63.560 ;
        RECT 4.400 56.760 46.000 58.160 ;
        RECT 4.000 55.440 46.000 56.760 ;
        RECT 4.000 54.040 45.600 55.440 ;
        RECT 4.000 51.360 46.000 54.040 ;
        RECT 4.400 49.960 46.000 51.360 ;
        RECT 4.000 44.560 46.000 49.960 ;
        RECT 4.400 43.160 46.000 44.560 ;
        RECT 4.000 37.760 46.000 43.160 ;
        RECT 4.400 36.360 46.000 37.760 ;
        RECT 4.000 30.960 46.000 36.360 ;
        RECT 4.400 29.560 46.000 30.960 ;
        RECT 4.000 24.160 46.000 29.560 ;
        RECT 4.400 22.760 46.000 24.160 ;
        RECT 4.000 17.360 46.000 22.760 ;
        RECT 4.400 15.960 46.000 17.360 ;
        RECT 4.000 10.560 46.000 15.960 ;
        RECT 4.400 9.160 46.000 10.560 ;
        RECT 4.000 3.760 46.000 9.160 ;
        RECT 4.400 2.910 46.000 3.760 ;
  END
END mux16x1_project
END LIBRARY

