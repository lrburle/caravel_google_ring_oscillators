* NGSPICE file created from sky130_osu_ring_oscillator_mpr2ca_8_b0r1.ext - technology: sky130A

.subckt sky130_osu_sc_12T_hs__mux2_1 S0 Y A0 A1 vccd1 vssd1 
X0 Y S0 A0 vccd1 sky130_fd_pr__pfet_01v8 ad=0.1764 pd=1.54 as=0.3402 ps=3.06 w=1.26 l=0.15
X1 Y a_110_114# A0 vssd1  sky130_fd_pr__nfet_01v8_lvt ad=0.077 pd=0.83 as=0.1485 ps=1.64 w=0.55 l=0.15
X2 A1 a_110_114# Y vccd1 sky130_fd_pr__pfet_01v8 ad=0.3339 pd=3.05 as=0.1764 ps=1.54 w=1.26 l=0.15
X3 A1 S0 Y vssd1  sky130_fd_pr__nfet_01v8_lvt ad=0.14575 pd=1.63 as=0.077 ps=0.83 w=0.55 l=0.15
X4 a_110_114# S0 vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0.3339 pd=3.05 as=0.3402 ps=3.06 w=1.26 l=0.15
X5 a_110_114# S0 vssd1  vssd1  sky130_fd_pr__nfet_01v8_lvt ad=0.14575 pd=1.63 as=0.1485 ps=1.64 w=0.55 l=0.15
.ends

.subckt scs130hd_mpr2ca_8 A1 B1 R3 R2 R1 R0 B0 A0 vpwr VNB VPB VSUBS
X0 a_772_910# B0 VNB VSUBS sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.86 as=0.234 ps=2.02 w=0.65 l=0.15
X1 a_178_822# A0 a_352_928# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1176 pd=1.4 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 a_296_52# a_48_92# a_208_310# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1079 ps=1.36 w=0.42 l=0.15
X3 a_824_46# B1 a_752_46# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0441 ps=0.63 w=0.42 l=0.15
X4 VNB a_844_910# R1 VSUBS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 vpwr A1 a_670_46# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.140425 pd=1.335 as=0.0672 ps=0.74 w=0.42 l=0.15
X6 R3 a_670_46# vpwr VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.140425 ps=1.335 w=1 l=0.15
X7 a_352_928# B0 VNB VSUBS sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1118 ps=1.04 w=0.42 l=0.15
X8 vpwr A1 a_208_310# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.140425 pd=1.335 as=0.07525 ps=0.82 w=0.42 l=0.15
X9 a_368_52# B1 a_296_52# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0525 pd=0.67 as=0.0441 ps=0.63 w=0.42 l=0.15
X10 VNB A1 a_824_46# VSUBS sky130_fd_pr__nfet_01v8 ad=0.13165 pd=1.14 as=0.0441 ps=0.63 w=0.42 l=0.15
X11 vpwr a_178_822# R0 VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1718 pd=1.39 as=0.47 ps=2.94 w=1 l=0.15
X12 a_208_310# B1 vpwr VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07525 pd=0.82 as=0.0567 ps=0.69 w=0.42 l=0.15
X13 vpwr a_844_910# a_1212_296# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X14 vpwr a_48_92# a_208_310# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1085 ps=1.36 w=0.42 l=0.15
X15 a_178_822# B0 vpwr VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.1718 ps=1.39 w=0.42 l=0.15
X16 a_48_92# R3 vpwr VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11055 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X17 vpwr A1 a_760_590# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X18 a_670_46# B1 vpwr VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0672 pd=0.74 as=0.0567 ps=0.69 w=0.42 l=0.15
X19 a_1212_296# R3 R1 VPB sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X20 R2 a_208_310# VNB VSUBS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.1222 ps=1.08 w=0.65 l=0.15
X21 a_844_910# B1 a_760_590# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X22 vpwr R0 a_670_46# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X23 R3 a_670_46# VNB VSUBS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.13165 ps=1.14 w=0.65 l=0.15
X24 a_760_590# B0 vpwr VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.3 ps=2.6 w=1 l=0.15
X25 VNB A1 a_368_52# VSUBS sky130_fd_pr__nfet_01v8 ad=0.1222 pd=1.08 as=0.0525 ps=0.67 w=0.42 l=0.15
X26 VNB a_178_822# R0 VSUBS sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.182 ps=1.86 w=0.65 l=0.15
X27 a_1040_910# A0 a_844_910# VSUBS sky130_fd_pr__nfet_01v8 ad=0.07475 pd=0.88 as=0.169 ps=1.82 w=0.65 l=0.15
X28 vpwr A0 a_178_822# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1197 pd=1.41 as=0.0588 ps=0.7 w=0.42 l=0.15
X29 a_48_92# R3 VNB VSUBS sky130_fd_pr__nfet_01v8 ad=0.1099 pd=1.37 as=0.1113 ps=1.37 w=0.42 l=0.15
X30 R1 R3 VNB VSUBS sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X31 a_844_910# A1 a_772_910# VSUBS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.06825 ps=0.86 w=0.65 l=0.15
X32 R2 a_208_310# vpwr VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.140425 ps=1.335 w=1 l=0.15
X33 a_760_590# A0 a_844_910# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X34 a_752_46# R0 a_670_46# VSUBS sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X35 VNB B1 a_1040_910# VSUBS sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.07475 ps=0.88 w=0.65 l=0.15
.ends

.subckt sky130_osu_sc_12T_hs__inv_1 Y A vccd1 vssd1
X0 Y A vccd1 vccd1 sky130_fd_pr__pfet_01v8 ad=0.3339 pd=3.05 as=0.3402 ps=3.06 w=1.26 l=0.15
X1 Y A vssd1 vssd1 sky130_fd_pr__nfet_01v8_lvt ad=0.14575 pd=1.63 as=0.1485 ps=1.64 w=0.55 l=0.15
.ends

.subckt sky130_osu_single_mpr2ca_8_b0r1 vccd1 in Y0 Y1 sel scs130hd_mpr2ca_8_0/B1
+ vssd1
Xsky130_osu_sc_12T_hs__mux2_1_0 sel sky130_osu_sc_12T_hs__inv_1_1/A in scs130hd_mpr2ca_8_0/R1
+ vccd1 vssd1 sky130_osu_sc_12T_hs__mux2_1
Xscs130hd_mpr2ca_8_0 scs130hd_mpr2ca_8_0/B1 scs130hd_mpr2ca_8_0/B1 scs130hd_mpr2ca_8_0/R3
+ scs130hd_mpr2ca_8_0/R2 scs130hd_mpr2ca_8_0/R1 scs130hd_mpr2ca_8_0/R0 vssd1 scs130hd_mpr2ca_8_0/B1
+ vccd1 vssd1 vccd1 vssd1 scs130hd_mpr2ca_8
Xsky130_osu_sc_12T_hs__mux2_1_1 sel scs130hd_mpr2ca_8_0/B1 vssd1 in vccd1 vssd1 sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__inv_1_1 sky130_osu_sc_12T_hs__inv_1_2/A sky130_osu_sc_12T_hs__inv_1_1/A
+ vccd1 vssd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__inv_1_2 Y1 sky130_osu_sc_12T_hs__inv_1_2/A vccd1 vssd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__mux2_1_2 sel sky130_osu_sc_12T_hs__inv_1_4/A scs130hd_mpr2ca_8_0/R1
+ in vccd1 vssd1 sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_sc_12T_hs__inv_1_3 Y0 sky130_osu_sc_12T_hs__inv_1_4/Y vccd1 vssd1 sky130_osu_sc_12T_hs__inv_1
Xsky130_osu_sc_12T_hs__inv_1_4 sky130_osu_sc_12T_hs__inv_1_4/Y sky130_osu_sc_12T_hs__inv_1_4/A
+ vccd1 vssd1 sky130_osu_sc_12T_hs__inv_1
.ends

.subckt sky130_osu_ring_oscillator_mpr2ca_8_b0r1 s1 s2 s3 s4 s5 X5_Y1 X4_Y1 X3_Y1
+ X2_Y1 X1_Y1 start vccd1 vssd1
Xsky130_osu_single_mpr2ca_8_b0r1_0 vccd1 sky130_osu_single_mpr2ca_8_b0r1_4/Y0 sky130_osu_sc_12T_hs__mux2_1_0/A0
+ X5_Y1 s5 sky130_osu_single_mpr2ca_8_b0r1_0/scs130hd_mpr2ca_8_0/B1 vssd1 sky130_osu_single_mpr2ca_8_b0r1
Xsky130_osu_single_mpr2ca_8_b0r1_1 vccd1 sky130_osu_sc_12T_hs__mux2_1_0/Y sky130_osu_single_mpr2ca_8_b0r1_2/in
+ X1_Y1 s1 sky130_osu_single_mpr2ca_8_b0r1_1/scs130hd_mpr2ca_8_0/B1 vssd1 sky130_osu_single_mpr2ca_8_b0r1
Xsky130_osu_sc_12T_hs__mux2_1_0 start sky130_osu_sc_12T_hs__mux2_1_0/Y sky130_osu_sc_12T_hs__mux2_1_0/A0
+ vccd1 vccd1 vssd1 sky130_osu_sc_12T_hs__mux2_1
Xsky130_osu_single_mpr2ca_8_b0r1_2 vccd1 sky130_osu_single_mpr2ca_8_b0r1_2/in sky130_osu_single_mpr2ca_8_b0r1_3/in
+ X2_Y1 s2 sky130_osu_single_mpr2ca_8_b0r1_2/scs130hd_mpr2ca_8_0/B1 vssd1 sky130_osu_single_mpr2ca_8_b0r1
Xsky130_osu_single_mpr2ca_8_b0r1_3 vccd1 sky130_osu_single_mpr2ca_8_b0r1_3/in sky130_osu_single_mpr2ca_8_b0r1_4/in
+ X3_Y1 s3 sky130_osu_single_mpr2ca_8_b0r1_3/scs130hd_mpr2ca_8_0/B1 vssd1 sky130_osu_single_mpr2ca_8_b0r1
Xsky130_osu_single_mpr2ca_8_b0r1_4 vccd1 sky130_osu_single_mpr2ca_8_b0r1_4/in sky130_osu_single_mpr2ca_8_b0r1_4/Y0
+ X4_Y1 s4 sky130_osu_single_mpr2ca_8_b0r1_4/scs130hd_mpr2ca_8_0/B1 vssd1 sky130_osu_single_mpr2ca_8_b0r1
.ends

