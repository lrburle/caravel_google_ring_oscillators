magic
tech sky130A
magscale 1 2
timestamp 1699053139
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 580262 404968 580318 404977
rect 580262 404903 580318 404912
rect 486238 351928 486294 351937
rect 486238 351863 486294 351872
rect 484030 343768 484086 343777
rect 484030 343703 484086 343712
rect 484044 341986 484072 343703
rect 486252 342258 486280 351863
rect 580276 344321 580304 404903
rect 488998 344312 489054 344321
rect 488998 344247 489054 344256
rect 580262 344312 580318 344321
rect 580262 344247 580318 344256
rect 483736 341958 484072 341986
rect 486206 342230 486280 342258
rect 486206 341972 486234 342230
rect 489012 341986 489040 344247
rect 490562 343768 490618 343777
rect 490562 343703 490618 343712
rect 488704 341958 489040 341986
rect 480640 341414 481252 341442
rect 480640 245585 480668 341414
rect 490576 298761 490604 343703
rect 490562 298752 490618 298761
rect 490562 298687 490618 298696
rect 480626 245576 480682 245585
rect 480626 245511 480682 245520
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 580262 404912 580318 404968
rect 486238 351872 486294 351928
rect 484030 343712 484086 343768
rect 488998 344256 489054 344312
rect 580262 344256 580318 344312
rect 490562 343712 490618 343768
rect 490562 298696 490618 298752
rect 480626 245520 480682 245576
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 580257 404970 580323 404973
rect 583520 404970 584960 405060
rect 580257 404968 584960 404970
rect 580257 404912 580262 404968
rect 580318 404912 584960 404968
rect 580257 404910 584960 404912
rect 580257 404907 580323 404910
rect 583520 404820 584960 404910
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 486233 351930 486299 351933
rect 583520 351930 584960 352020
rect 486233 351928 584960 351930
rect 486233 351872 486238 351928
rect 486294 351872 584960 351928
rect 486233 351870 584960 351872
rect 486233 351867 486299 351870
rect 583520 351780 584960 351870
rect -960 345252 480 345492
rect 488993 344314 489059 344317
rect 580257 344314 580323 344317
rect 488993 344312 580323 344314
rect 488993 344256 488998 344312
rect 489054 344256 580262 344312
rect 580318 344256 580323 344312
rect 488993 344254 580323 344256
rect 488993 344251 489059 344254
rect 580257 344251 580323 344254
rect 484025 343770 484091 343773
rect 490557 343770 490623 343773
rect 484025 343768 490623 343770
rect 484025 343712 484030 343768
rect 484086 343712 490562 343768
rect 490618 343712 490623 343768
rect 484025 343710 490623 343712
rect 484025 343707 484091 343710
rect 490557 343707 490623 343710
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 491886 330986 491892 330988
rect 489900 330926 491892 330986
rect 491886 330924 491892 330926
rect 491956 330924 491962 330988
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 490557 298754 490623 298757
rect 583520 298754 584960 298844
rect 490557 298752 584960 298754
rect 490557 298696 490562 298752
rect 490618 298696 584960 298752
rect 490557 298694 584960 298696
rect 490557 298691 490623 298694
rect 583520 298604 584960 298694
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 480621 245578 480687 245581
rect 583520 245578 584960 245668
rect 480621 245576 584960 245578
rect 480621 245520 480626 245576
rect 480682 245520 584960 245576
rect 480621 245518 584960 245520
rect 480621 245515 480687 245518
rect 583520 245428 584960 245518
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 491886 19756 491892 19820
rect 491956 19818 491962 19820
rect 583520 19818 584960 19908
rect 491956 19758 584960 19818
rect 491956 19756 491962 19758
rect 583520 19668 584960 19758
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
<< via3 >>
rect 491892 330924 491956 330988
rect 491892 19756 491956 19820
<< metal4 >>
rect 1794 673054 2414 701760
rect 1794 672818 1826 673054
rect 2062 672818 2146 673054
rect 2382 672818 2414 673054
rect 1794 672734 2414 672818
rect 1794 672498 1826 672734
rect 2062 672498 2146 672734
rect 2382 672498 2414 672734
rect 1794 635854 2414 672498
rect 1794 635618 1826 635854
rect 2062 635618 2146 635854
rect 2382 635618 2414 635854
rect 1794 635534 2414 635618
rect 1794 635298 1826 635534
rect 2062 635298 2146 635534
rect 2382 635298 2414 635534
rect 1794 598654 2414 635298
rect 1794 598418 1826 598654
rect 2062 598418 2146 598654
rect 2382 598418 2414 598654
rect 1794 598334 2414 598418
rect 1794 598098 1826 598334
rect 2062 598098 2146 598334
rect 2382 598098 2414 598334
rect 1794 561454 2414 598098
rect 1794 561218 1826 561454
rect 2062 561218 2146 561454
rect 2382 561218 2414 561454
rect 1794 561134 2414 561218
rect 1794 560898 1826 561134
rect 2062 560898 2146 561134
rect 2382 560898 2414 561134
rect 1794 524254 2414 560898
rect 1794 524018 1826 524254
rect 2062 524018 2146 524254
rect 2382 524018 2414 524254
rect 1794 523934 2414 524018
rect 1794 523698 1826 523934
rect 2062 523698 2146 523934
rect 2382 523698 2414 523934
rect 1794 487054 2414 523698
rect 1794 486818 1826 487054
rect 2062 486818 2146 487054
rect 2382 486818 2414 487054
rect 1794 486734 2414 486818
rect 1794 486498 1826 486734
rect 2062 486498 2146 486734
rect 2382 486498 2414 486734
rect 1794 449854 2414 486498
rect 1794 449618 1826 449854
rect 2062 449618 2146 449854
rect 2382 449618 2414 449854
rect 1794 449534 2414 449618
rect 1794 449298 1826 449534
rect 2062 449298 2146 449534
rect 2382 449298 2414 449534
rect 1794 412654 2414 449298
rect 1794 412418 1826 412654
rect 2062 412418 2146 412654
rect 2382 412418 2414 412654
rect 1794 412334 2414 412418
rect 1794 412098 1826 412334
rect 2062 412098 2146 412334
rect 2382 412098 2414 412334
rect 1794 375454 2414 412098
rect 1794 375218 1826 375454
rect 2062 375218 2146 375454
rect 2382 375218 2414 375454
rect 1794 375134 2414 375218
rect 1794 374898 1826 375134
rect 2062 374898 2146 375134
rect 2382 374898 2414 375134
rect 1794 338254 2414 374898
rect 1794 338018 1826 338254
rect 2062 338018 2146 338254
rect 2382 338018 2414 338254
rect 1794 337934 2414 338018
rect 1794 337698 1826 337934
rect 2062 337698 2146 337934
rect 2382 337698 2414 337934
rect 1794 301054 2414 337698
rect 1794 300818 1826 301054
rect 2062 300818 2146 301054
rect 2382 300818 2414 301054
rect 1794 300734 2414 300818
rect 1794 300498 1826 300734
rect 2062 300498 2146 300734
rect 2382 300498 2414 300734
rect 1794 263854 2414 300498
rect 1794 263618 1826 263854
rect 2062 263618 2146 263854
rect 2382 263618 2414 263854
rect 1794 263534 2414 263618
rect 1794 263298 1826 263534
rect 2062 263298 2146 263534
rect 2382 263298 2414 263534
rect 1794 226654 2414 263298
rect 1794 226418 1826 226654
rect 2062 226418 2146 226654
rect 2382 226418 2414 226654
rect 1794 226334 2414 226418
rect 1794 226098 1826 226334
rect 2062 226098 2146 226334
rect 2382 226098 2414 226334
rect 1794 189454 2414 226098
rect 1794 189218 1826 189454
rect 2062 189218 2146 189454
rect 2382 189218 2414 189454
rect 1794 189134 2414 189218
rect 1794 188898 1826 189134
rect 2062 188898 2146 189134
rect 2382 188898 2414 189134
rect 1794 152254 2414 188898
rect 1794 152018 1826 152254
rect 2062 152018 2146 152254
rect 2382 152018 2414 152254
rect 1794 151934 2414 152018
rect 1794 151698 1826 151934
rect 2062 151698 2146 151934
rect 2382 151698 2414 151934
rect 1794 115054 2414 151698
rect 1794 114818 1826 115054
rect 2062 114818 2146 115054
rect 2382 114818 2414 115054
rect 1794 114734 2414 114818
rect 1794 114498 1826 114734
rect 2062 114498 2146 114734
rect 2382 114498 2414 114734
rect 1794 77854 2414 114498
rect 1794 77618 1826 77854
rect 2062 77618 2146 77854
rect 2382 77618 2414 77854
rect 1794 77534 2414 77618
rect 1794 77298 1826 77534
rect 2062 77298 2146 77534
rect 2382 77298 2414 77534
rect 1794 40654 2414 77298
rect 1794 40418 1826 40654
rect 2062 40418 2146 40654
rect 2382 40418 2414 40654
rect 1794 40334 2414 40418
rect 1794 40098 1826 40334
rect 2062 40098 2146 40334
rect 2382 40098 2414 40334
rect 1794 3454 2414 40098
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 2176 2414 2898
rect 5514 676774 6134 701760
rect 5514 676538 5546 676774
rect 5782 676538 5866 676774
rect 6102 676538 6134 676774
rect 5514 676454 6134 676538
rect 5514 676218 5546 676454
rect 5782 676218 5866 676454
rect 6102 676218 6134 676454
rect 5514 639574 6134 676218
rect 5514 639338 5546 639574
rect 5782 639338 5866 639574
rect 6102 639338 6134 639574
rect 5514 639254 6134 639338
rect 5514 639018 5546 639254
rect 5782 639018 5866 639254
rect 6102 639018 6134 639254
rect 5514 602374 6134 639018
rect 5514 602138 5546 602374
rect 5782 602138 5866 602374
rect 6102 602138 6134 602374
rect 5514 602054 6134 602138
rect 5514 601818 5546 602054
rect 5782 601818 5866 602054
rect 6102 601818 6134 602054
rect 5514 565174 6134 601818
rect 5514 564938 5546 565174
rect 5782 564938 5866 565174
rect 6102 564938 6134 565174
rect 5514 564854 6134 564938
rect 5514 564618 5546 564854
rect 5782 564618 5866 564854
rect 6102 564618 6134 564854
rect 5514 527974 6134 564618
rect 5514 527738 5546 527974
rect 5782 527738 5866 527974
rect 6102 527738 6134 527974
rect 5514 527654 6134 527738
rect 5514 527418 5546 527654
rect 5782 527418 5866 527654
rect 6102 527418 6134 527654
rect 5514 490774 6134 527418
rect 5514 490538 5546 490774
rect 5782 490538 5866 490774
rect 6102 490538 6134 490774
rect 5514 490454 6134 490538
rect 5514 490218 5546 490454
rect 5782 490218 5866 490454
rect 6102 490218 6134 490454
rect 5514 453574 6134 490218
rect 5514 453338 5546 453574
rect 5782 453338 5866 453574
rect 6102 453338 6134 453574
rect 5514 453254 6134 453338
rect 5514 453018 5546 453254
rect 5782 453018 5866 453254
rect 6102 453018 6134 453254
rect 5514 416374 6134 453018
rect 5514 416138 5546 416374
rect 5782 416138 5866 416374
rect 6102 416138 6134 416374
rect 5514 416054 6134 416138
rect 5514 415818 5546 416054
rect 5782 415818 5866 416054
rect 6102 415818 6134 416054
rect 5514 379174 6134 415818
rect 5514 378938 5546 379174
rect 5782 378938 5866 379174
rect 6102 378938 6134 379174
rect 5514 378854 6134 378938
rect 5514 378618 5546 378854
rect 5782 378618 5866 378854
rect 6102 378618 6134 378854
rect 5514 341974 6134 378618
rect 5514 341738 5546 341974
rect 5782 341738 5866 341974
rect 6102 341738 6134 341974
rect 5514 341654 6134 341738
rect 5514 341418 5546 341654
rect 5782 341418 5866 341654
rect 6102 341418 6134 341654
rect 5514 304774 6134 341418
rect 5514 304538 5546 304774
rect 5782 304538 5866 304774
rect 6102 304538 6134 304774
rect 5514 304454 6134 304538
rect 5514 304218 5546 304454
rect 5782 304218 5866 304454
rect 6102 304218 6134 304454
rect 5514 267574 6134 304218
rect 5514 267338 5546 267574
rect 5782 267338 5866 267574
rect 6102 267338 6134 267574
rect 5514 267254 6134 267338
rect 5514 267018 5546 267254
rect 5782 267018 5866 267254
rect 6102 267018 6134 267254
rect 5514 230374 6134 267018
rect 5514 230138 5546 230374
rect 5782 230138 5866 230374
rect 6102 230138 6134 230374
rect 5514 230054 6134 230138
rect 5514 229818 5546 230054
rect 5782 229818 5866 230054
rect 6102 229818 6134 230054
rect 5514 193174 6134 229818
rect 5514 192938 5546 193174
rect 5782 192938 5866 193174
rect 6102 192938 6134 193174
rect 5514 192854 6134 192938
rect 5514 192618 5546 192854
rect 5782 192618 5866 192854
rect 6102 192618 6134 192854
rect 5514 155974 6134 192618
rect 5514 155738 5546 155974
rect 5782 155738 5866 155974
rect 6102 155738 6134 155974
rect 5514 155654 6134 155738
rect 5514 155418 5546 155654
rect 5782 155418 5866 155654
rect 6102 155418 6134 155654
rect 5514 118774 6134 155418
rect 5514 118538 5546 118774
rect 5782 118538 5866 118774
rect 6102 118538 6134 118774
rect 5514 118454 6134 118538
rect 5514 118218 5546 118454
rect 5782 118218 5866 118454
rect 6102 118218 6134 118454
rect 5514 81574 6134 118218
rect 5514 81338 5546 81574
rect 5782 81338 5866 81574
rect 6102 81338 6134 81574
rect 5514 81254 6134 81338
rect 5514 81018 5546 81254
rect 5782 81018 5866 81254
rect 6102 81018 6134 81254
rect 5514 44374 6134 81018
rect 5514 44138 5546 44374
rect 5782 44138 5866 44374
rect 6102 44138 6134 44374
rect 5514 44054 6134 44138
rect 5514 43818 5546 44054
rect 5782 43818 5866 44054
rect 6102 43818 6134 44054
rect 5514 7174 6134 43818
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect 5514 2176 6134 6618
rect 9234 680494 9854 701760
rect 9234 680258 9266 680494
rect 9502 680258 9586 680494
rect 9822 680258 9854 680494
rect 9234 680174 9854 680258
rect 9234 679938 9266 680174
rect 9502 679938 9586 680174
rect 9822 679938 9854 680174
rect 9234 643294 9854 679938
rect 9234 643058 9266 643294
rect 9502 643058 9586 643294
rect 9822 643058 9854 643294
rect 9234 642974 9854 643058
rect 9234 642738 9266 642974
rect 9502 642738 9586 642974
rect 9822 642738 9854 642974
rect 9234 606094 9854 642738
rect 9234 605858 9266 606094
rect 9502 605858 9586 606094
rect 9822 605858 9854 606094
rect 9234 605774 9854 605858
rect 9234 605538 9266 605774
rect 9502 605538 9586 605774
rect 9822 605538 9854 605774
rect 9234 568894 9854 605538
rect 9234 568658 9266 568894
rect 9502 568658 9586 568894
rect 9822 568658 9854 568894
rect 9234 568574 9854 568658
rect 9234 568338 9266 568574
rect 9502 568338 9586 568574
rect 9822 568338 9854 568574
rect 9234 531694 9854 568338
rect 9234 531458 9266 531694
rect 9502 531458 9586 531694
rect 9822 531458 9854 531694
rect 9234 531374 9854 531458
rect 9234 531138 9266 531374
rect 9502 531138 9586 531374
rect 9822 531138 9854 531374
rect 9234 494494 9854 531138
rect 9234 494258 9266 494494
rect 9502 494258 9586 494494
rect 9822 494258 9854 494494
rect 9234 494174 9854 494258
rect 9234 493938 9266 494174
rect 9502 493938 9586 494174
rect 9822 493938 9854 494174
rect 9234 457294 9854 493938
rect 9234 457058 9266 457294
rect 9502 457058 9586 457294
rect 9822 457058 9854 457294
rect 9234 456974 9854 457058
rect 9234 456738 9266 456974
rect 9502 456738 9586 456974
rect 9822 456738 9854 456974
rect 9234 420094 9854 456738
rect 9234 419858 9266 420094
rect 9502 419858 9586 420094
rect 9822 419858 9854 420094
rect 9234 419774 9854 419858
rect 9234 419538 9266 419774
rect 9502 419538 9586 419774
rect 9822 419538 9854 419774
rect 9234 382894 9854 419538
rect 9234 382658 9266 382894
rect 9502 382658 9586 382894
rect 9822 382658 9854 382894
rect 9234 382574 9854 382658
rect 9234 382338 9266 382574
rect 9502 382338 9586 382574
rect 9822 382338 9854 382574
rect 9234 345694 9854 382338
rect 9234 345458 9266 345694
rect 9502 345458 9586 345694
rect 9822 345458 9854 345694
rect 9234 345374 9854 345458
rect 9234 345138 9266 345374
rect 9502 345138 9586 345374
rect 9822 345138 9854 345374
rect 9234 308494 9854 345138
rect 9234 308258 9266 308494
rect 9502 308258 9586 308494
rect 9822 308258 9854 308494
rect 9234 308174 9854 308258
rect 9234 307938 9266 308174
rect 9502 307938 9586 308174
rect 9822 307938 9854 308174
rect 9234 271294 9854 307938
rect 9234 271058 9266 271294
rect 9502 271058 9586 271294
rect 9822 271058 9854 271294
rect 9234 270974 9854 271058
rect 9234 270738 9266 270974
rect 9502 270738 9586 270974
rect 9822 270738 9854 270974
rect 9234 234094 9854 270738
rect 9234 233858 9266 234094
rect 9502 233858 9586 234094
rect 9822 233858 9854 234094
rect 9234 233774 9854 233858
rect 9234 233538 9266 233774
rect 9502 233538 9586 233774
rect 9822 233538 9854 233774
rect 9234 196894 9854 233538
rect 9234 196658 9266 196894
rect 9502 196658 9586 196894
rect 9822 196658 9854 196894
rect 9234 196574 9854 196658
rect 9234 196338 9266 196574
rect 9502 196338 9586 196574
rect 9822 196338 9854 196574
rect 9234 159694 9854 196338
rect 9234 159458 9266 159694
rect 9502 159458 9586 159694
rect 9822 159458 9854 159694
rect 9234 159374 9854 159458
rect 9234 159138 9266 159374
rect 9502 159138 9586 159374
rect 9822 159138 9854 159374
rect 9234 122494 9854 159138
rect 9234 122258 9266 122494
rect 9502 122258 9586 122494
rect 9822 122258 9854 122494
rect 9234 122174 9854 122258
rect 9234 121938 9266 122174
rect 9502 121938 9586 122174
rect 9822 121938 9854 122174
rect 9234 85294 9854 121938
rect 9234 85058 9266 85294
rect 9502 85058 9586 85294
rect 9822 85058 9854 85294
rect 9234 84974 9854 85058
rect 9234 84738 9266 84974
rect 9502 84738 9586 84974
rect 9822 84738 9854 84974
rect 9234 48094 9854 84738
rect 9234 47858 9266 48094
rect 9502 47858 9586 48094
rect 9822 47858 9854 48094
rect 9234 47774 9854 47858
rect 9234 47538 9266 47774
rect 9502 47538 9586 47774
rect 9822 47538 9854 47774
rect 9234 10894 9854 47538
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect 9234 2176 9854 10338
rect 12954 684214 13574 701760
rect 12954 683978 12986 684214
rect 13222 683978 13306 684214
rect 13542 683978 13574 684214
rect 12954 683894 13574 683978
rect 12954 683658 12986 683894
rect 13222 683658 13306 683894
rect 13542 683658 13574 683894
rect 12954 647014 13574 683658
rect 12954 646778 12986 647014
rect 13222 646778 13306 647014
rect 13542 646778 13574 647014
rect 12954 646694 13574 646778
rect 12954 646458 12986 646694
rect 13222 646458 13306 646694
rect 13542 646458 13574 646694
rect 12954 609814 13574 646458
rect 12954 609578 12986 609814
rect 13222 609578 13306 609814
rect 13542 609578 13574 609814
rect 12954 609494 13574 609578
rect 12954 609258 12986 609494
rect 13222 609258 13306 609494
rect 13542 609258 13574 609494
rect 12954 572614 13574 609258
rect 12954 572378 12986 572614
rect 13222 572378 13306 572614
rect 13542 572378 13574 572614
rect 12954 572294 13574 572378
rect 12954 572058 12986 572294
rect 13222 572058 13306 572294
rect 13542 572058 13574 572294
rect 12954 535414 13574 572058
rect 12954 535178 12986 535414
rect 13222 535178 13306 535414
rect 13542 535178 13574 535414
rect 12954 535094 13574 535178
rect 12954 534858 12986 535094
rect 13222 534858 13306 535094
rect 13542 534858 13574 535094
rect 12954 498214 13574 534858
rect 12954 497978 12986 498214
rect 13222 497978 13306 498214
rect 13542 497978 13574 498214
rect 12954 497894 13574 497978
rect 12954 497658 12986 497894
rect 13222 497658 13306 497894
rect 13542 497658 13574 497894
rect 12954 461014 13574 497658
rect 12954 460778 12986 461014
rect 13222 460778 13306 461014
rect 13542 460778 13574 461014
rect 12954 460694 13574 460778
rect 12954 460458 12986 460694
rect 13222 460458 13306 460694
rect 13542 460458 13574 460694
rect 12954 423814 13574 460458
rect 12954 423578 12986 423814
rect 13222 423578 13306 423814
rect 13542 423578 13574 423814
rect 12954 423494 13574 423578
rect 12954 423258 12986 423494
rect 13222 423258 13306 423494
rect 13542 423258 13574 423494
rect 12954 386614 13574 423258
rect 12954 386378 12986 386614
rect 13222 386378 13306 386614
rect 13542 386378 13574 386614
rect 12954 386294 13574 386378
rect 12954 386058 12986 386294
rect 13222 386058 13306 386294
rect 13542 386058 13574 386294
rect 12954 349414 13574 386058
rect 12954 349178 12986 349414
rect 13222 349178 13306 349414
rect 13542 349178 13574 349414
rect 12954 349094 13574 349178
rect 12954 348858 12986 349094
rect 13222 348858 13306 349094
rect 13542 348858 13574 349094
rect 12954 312214 13574 348858
rect 12954 311978 12986 312214
rect 13222 311978 13306 312214
rect 13542 311978 13574 312214
rect 12954 311894 13574 311978
rect 12954 311658 12986 311894
rect 13222 311658 13306 311894
rect 13542 311658 13574 311894
rect 12954 275014 13574 311658
rect 12954 274778 12986 275014
rect 13222 274778 13306 275014
rect 13542 274778 13574 275014
rect 12954 274694 13574 274778
rect 12954 274458 12986 274694
rect 13222 274458 13306 274694
rect 13542 274458 13574 274694
rect 12954 237814 13574 274458
rect 12954 237578 12986 237814
rect 13222 237578 13306 237814
rect 13542 237578 13574 237814
rect 12954 237494 13574 237578
rect 12954 237258 12986 237494
rect 13222 237258 13306 237494
rect 13542 237258 13574 237494
rect 12954 200614 13574 237258
rect 12954 200378 12986 200614
rect 13222 200378 13306 200614
rect 13542 200378 13574 200614
rect 12954 200294 13574 200378
rect 12954 200058 12986 200294
rect 13222 200058 13306 200294
rect 13542 200058 13574 200294
rect 12954 163414 13574 200058
rect 12954 163178 12986 163414
rect 13222 163178 13306 163414
rect 13542 163178 13574 163414
rect 12954 163094 13574 163178
rect 12954 162858 12986 163094
rect 13222 162858 13306 163094
rect 13542 162858 13574 163094
rect 12954 126214 13574 162858
rect 12954 125978 12986 126214
rect 13222 125978 13306 126214
rect 13542 125978 13574 126214
rect 12954 125894 13574 125978
rect 12954 125658 12986 125894
rect 13222 125658 13306 125894
rect 13542 125658 13574 125894
rect 12954 89014 13574 125658
rect 12954 88778 12986 89014
rect 13222 88778 13306 89014
rect 13542 88778 13574 89014
rect 12954 88694 13574 88778
rect 12954 88458 12986 88694
rect 13222 88458 13306 88694
rect 13542 88458 13574 88694
rect 12954 51814 13574 88458
rect 12954 51578 12986 51814
rect 13222 51578 13306 51814
rect 13542 51578 13574 51814
rect 12954 51494 13574 51578
rect 12954 51258 12986 51494
rect 13222 51258 13306 51494
rect 13542 51258 13574 51494
rect 12954 14614 13574 51258
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect 12954 2176 13574 14058
rect 16674 687934 17294 701760
rect 16674 687698 16706 687934
rect 16942 687698 17026 687934
rect 17262 687698 17294 687934
rect 16674 687614 17294 687698
rect 16674 687378 16706 687614
rect 16942 687378 17026 687614
rect 17262 687378 17294 687614
rect 16674 650734 17294 687378
rect 16674 650498 16706 650734
rect 16942 650498 17026 650734
rect 17262 650498 17294 650734
rect 16674 650414 17294 650498
rect 16674 650178 16706 650414
rect 16942 650178 17026 650414
rect 17262 650178 17294 650414
rect 16674 613534 17294 650178
rect 16674 613298 16706 613534
rect 16942 613298 17026 613534
rect 17262 613298 17294 613534
rect 16674 613214 17294 613298
rect 16674 612978 16706 613214
rect 16942 612978 17026 613214
rect 17262 612978 17294 613214
rect 16674 576334 17294 612978
rect 16674 576098 16706 576334
rect 16942 576098 17026 576334
rect 17262 576098 17294 576334
rect 16674 576014 17294 576098
rect 16674 575778 16706 576014
rect 16942 575778 17026 576014
rect 17262 575778 17294 576014
rect 16674 539134 17294 575778
rect 16674 538898 16706 539134
rect 16942 538898 17026 539134
rect 17262 538898 17294 539134
rect 16674 538814 17294 538898
rect 16674 538578 16706 538814
rect 16942 538578 17026 538814
rect 17262 538578 17294 538814
rect 16674 501934 17294 538578
rect 16674 501698 16706 501934
rect 16942 501698 17026 501934
rect 17262 501698 17294 501934
rect 16674 501614 17294 501698
rect 16674 501378 16706 501614
rect 16942 501378 17026 501614
rect 17262 501378 17294 501614
rect 16674 464734 17294 501378
rect 16674 464498 16706 464734
rect 16942 464498 17026 464734
rect 17262 464498 17294 464734
rect 16674 464414 17294 464498
rect 16674 464178 16706 464414
rect 16942 464178 17026 464414
rect 17262 464178 17294 464414
rect 16674 427534 17294 464178
rect 16674 427298 16706 427534
rect 16942 427298 17026 427534
rect 17262 427298 17294 427534
rect 16674 427214 17294 427298
rect 16674 426978 16706 427214
rect 16942 426978 17026 427214
rect 17262 426978 17294 427214
rect 16674 390334 17294 426978
rect 16674 390098 16706 390334
rect 16942 390098 17026 390334
rect 17262 390098 17294 390334
rect 16674 390014 17294 390098
rect 16674 389778 16706 390014
rect 16942 389778 17026 390014
rect 17262 389778 17294 390014
rect 16674 353134 17294 389778
rect 16674 352898 16706 353134
rect 16942 352898 17026 353134
rect 17262 352898 17294 353134
rect 16674 352814 17294 352898
rect 16674 352578 16706 352814
rect 16942 352578 17026 352814
rect 17262 352578 17294 352814
rect 16674 315934 17294 352578
rect 16674 315698 16706 315934
rect 16942 315698 17026 315934
rect 17262 315698 17294 315934
rect 16674 315614 17294 315698
rect 16674 315378 16706 315614
rect 16942 315378 17026 315614
rect 17262 315378 17294 315614
rect 16674 278734 17294 315378
rect 16674 278498 16706 278734
rect 16942 278498 17026 278734
rect 17262 278498 17294 278734
rect 16674 278414 17294 278498
rect 16674 278178 16706 278414
rect 16942 278178 17026 278414
rect 17262 278178 17294 278414
rect 16674 241534 17294 278178
rect 16674 241298 16706 241534
rect 16942 241298 17026 241534
rect 17262 241298 17294 241534
rect 16674 241214 17294 241298
rect 16674 240978 16706 241214
rect 16942 240978 17026 241214
rect 17262 240978 17294 241214
rect 16674 204334 17294 240978
rect 16674 204098 16706 204334
rect 16942 204098 17026 204334
rect 17262 204098 17294 204334
rect 16674 204014 17294 204098
rect 16674 203778 16706 204014
rect 16942 203778 17026 204014
rect 17262 203778 17294 204014
rect 16674 167134 17294 203778
rect 16674 166898 16706 167134
rect 16942 166898 17026 167134
rect 17262 166898 17294 167134
rect 16674 166814 17294 166898
rect 16674 166578 16706 166814
rect 16942 166578 17026 166814
rect 17262 166578 17294 166814
rect 16674 129934 17294 166578
rect 16674 129698 16706 129934
rect 16942 129698 17026 129934
rect 17262 129698 17294 129934
rect 16674 129614 17294 129698
rect 16674 129378 16706 129614
rect 16942 129378 17026 129614
rect 17262 129378 17294 129614
rect 16674 92734 17294 129378
rect 16674 92498 16706 92734
rect 16942 92498 17026 92734
rect 17262 92498 17294 92734
rect 16674 92414 17294 92498
rect 16674 92178 16706 92414
rect 16942 92178 17026 92414
rect 17262 92178 17294 92414
rect 16674 55534 17294 92178
rect 16674 55298 16706 55534
rect 16942 55298 17026 55534
rect 17262 55298 17294 55534
rect 16674 55214 17294 55298
rect 16674 54978 16706 55214
rect 16942 54978 17026 55214
rect 17262 54978 17294 55214
rect 16674 18334 17294 54978
rect 16674 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 17294 18334
rect 16674 18014 17294 18098
rect 16674 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 17294 18014
rect 16674 2176 17294 17778
rect 20394 691654 21014 701760
rect 20394 691418 20426 691654
rect 20662 691418 20746 691654
rect 20982 691418 21014 691654
rect 20394 691334 21014 691418
rect 20394 691098 20426 691334
rect 20662 691098 20746 691334
rect 20982 691098 21014 691334
rect 20394 654454 21014 691098
rect 20394 654218 20426 654454
rect 20662 654218 20746 654454
rect 20982 654218 21014 654454
rect 20394 654134 21014 654218
rect 20394 653898 20426 654134
rect 20662 653898 20746 654134
rect 20982 653898 21014 654134
rect 20394 617254 21014 653898
rect 20394 617018 20426 617254
rect 20662 617018 20746 617254
rect 20982 617018 21014 617254
rect 20394 616934 21014 617018
rect 20394 616698 20426 616934
rect 20662 616698 20746 616934
rect 20982 616698 21014 616934
rect 20394 580054 21014 616698
rect 20394 579818 20426 580054
rect 20662 579818 20746 580054
rect 20982 579818 21014 580054
rect 20394 579734 21014 579818
rect 20394 579498 20426 579734
rect 20662 579498 20746 579734
rect 20982 579498 21014 579734
rect 20394 542854 21014 579498
rect 20394 542618 20426 542854
rect 20662 542618 20746 542854
rect 20982 542618 21014 542854
rect 20394 542534 21014 542618
rect 20394 542298 20426 542534
rect 20662 542298 20746 542534
rect 20982 542298 21014 542534
rect 20394 505654 21014 542298
rect 20394 505418 20426 505654
rect 20662 505418 20746 505654
rect 20982 505418 21014 505654
rect 20394 505334 21014 505418
rect 20394 505098 20426 505334
rect 20662 505098 20746 505334
rect 20982 505098 21014 505334
rect 20394 468454 21014 505098
rect 20394 468218 20426 468454
rect 20662 468218 20746 468454
rect 20982 468218 21014 468454
rect 20394 468134 21014 468218
rect 20394 467898 20426 468134
rect 20662 467898 20746 468134
rect 20982 467898 21014 468134
rect 20394 431254 21014 467898
rect 20394 431018 20426 431254
rect 20662 431018 20746 431254
rect 20982 431018 21014 431254
rect 20394 430934 21014 431018
rect 20394 430698 20426 430934
rect 20662 430698 20746 430934
rect 20982 430698 21014 430934
rect 20394 394054 21014 430698
rect 20394 393818 20426 394054
rect 20662 393818 20746 394054
rect 20982 393818 21014 394054
rect 20394 393734 21014 393818
rect 20394 393498 20426 393734
rect 20662 393498 20746 393734
rect 20982 393498 21014 393734
rect 20394 356854 21014 393498
rect 20394 356618 20426 356854
rect 20662 356618 20746 356854
rect 20982 356618 21014 356854
rect 20394 356534 21014 356618
rect 20394 356298 20426 356534
rect 20662 356298 20746 356534
rect 20982 356298 21014 356534
rect 20394 319654 21014 356298
rect 20394 319418 20426 319654
rect 20662 319418 20746 319654
rect 20982 319418 21014 319654
rect 20394 319334 21014 319418
rect 20394 319098 20426 319334
rect 20662 319098 20746 319334
rect 20982 319098 21014 319334
rect 20394 282454 21014 319098
rect 20394 282218 20426 282454
rect 20662 282218 20746 282454
rect 20982 282218 21014 282454
rect 20394 282134 21014 282218
rect 20394 281898 20426 282134
rect 20662 281898 20746 282134
rect 20982 281898 21014 282134
rect 20394 245254 21014 281898
rect 20394 245018 20426 245254
rect 20662 245018 20746 245254
rect 20982 245018 21014 245254
rect 20394 244934 21014 245018
rect 20394 244698 20426 244934
rect 20662 244698 20746 244934
rect 20982 244698 21014 244934
rect 20394 208054 21014 244698
rect 20394 207818 20426 208054
rect 20662 207818 20746 208054
rect 20982 207818 21014 208054
rect 20394 207734 21014 207818
rect 20394 207498 20426 207734
rect 20662 207498 20746 207734
rect 20982 207498 21014 207734
rect 20394 170854 21014 207498
rect 20394 170618 20426 170854
rect 20662 170618 20746 170854
rect 20982 170618 21014 170854
rect 20394 170534 21014 170618
rect 20394 170298 20426 170534
rect 20662 170298 20746 170534
rect 20982 170298 21014 170534
rect 20394 133654 21014 170298
rect 20394 133418 20426 133654
rect 20662 133418 20746 133654
rect 20982 133418 21014 133654
rect 20394 133334 21014 133418
rect 20394 133098 20426 133334
rect 20662 133098 20746 133334
rect 20982 133098 21014 133334
rect 20394 96454 21014 133098
rect 20394 96218 20426 96454
rect 20662 96218 20746 96454
rect 20982 96218 21014 96454
rect 20394 96134 21014 96218
rect 20394 95898 20426 96134
rect 20662 95898 20746 96134
rect 20982 95898 21014 96134
rect 20394 59254 21014 95898
rect 20394 59018 20426 59254
rect 20662 59018 20746 59254
rect 20982 59018 21014 59254
rect 20394 58934 21014 59018
rect 20394 58698 20426 58934
rect 20662 58698 20746 58934
rect 20982 58698 21014 58934
rect 20394 22054 21014 58698
rect 20394 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 21014 22054
rect 20394 21734 21014 21818
rect 20394 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 21014 21734
rect 20394 2176 21014 21498
rect 24114 695374 24734 701760
rect 24114 695138 24146 695374
rect 24382 695138 24466 695374
rect 24702 695138 24734 695374
rect 24114 695054 24734 695138
rect 24114 694818 24146 695054
rect 24382 694818 24466 695054
rect 24702 694818 24734 695054
rect 24114 658174 24734 694818
rect 24114 657938 24146 658174
rect 24382 657938 24466 658174
rect 24702 657938 24734 658174
rect 24114 657854 24734 657938
rect 24114 657618 24146 657854
rect 24382 657618 24466 657854
rect 24702 657618 24734 657854
rect 24114 620974 24734 657618
rect 24114 620738 24146 620974
rect 24382 620738 24466 620974
rect 24702 620738 24734 620974
rect 24114 620654 24734 620738
rect 24114 620418 24146 620654
rect 24382 620418 24466 620654
rect 24702 620418 24734 620654
rect 24114 583774 24734 620418
rect 24114 583538 24146 583774
rect 24382 583538 24466 583774
rect 24702 583538 24734 583774
rect 24114 583454 24734 583538
rect 24114 583218 24146 583454
rect 24382 583218 24466 583454
rect 24702 583218 24734 583454
rect 24114 546574 24734 583218
rect 24114 546338 24146 546574
rect 24382 546338 24466 546574
rect 24702 546338 24734 546574
rect 24114 546254 24734 546338
rect 24114 546018 24146 546254
rect 24382 546018 24466 546254
rect 24702 546018 24734 546254
rect 24114 509374 24734 546018
rect 24114 509138 24146 509374
rect 24382 509138 24466 509374
rect 24702 509138 24734 509374
rect 24114 509054 24734 509138
rect 24114 508818 24146 509054
rect 24382 508818 24466 509054
rect 24702 508818 24734 509054
rect 24114 472174 24734 508818
rect 24114 471938 24146 472174
rect 24382 471938 24466 472174
rect 24702 471938 24734 472174
rect 24114 471854 24734 471938
rect 24114 471618 24146 471854
rect 24382 471618 24466 471854
rect 24702 471618 24734 471854
rect 24114 434974 24734 471618
rect 24114 434738 24146 434974
rect 24382 434738 24466 434974
rect 24702 434738 24734 434974
rect 24114 434654 24734 434738
rect 24114 434418 24146 434654
rect 24382 434418 24466 434654
rect 24702 434418 24734 434654
rect 24114 397774 24734 434418
rect 24114 397538 24146 397774
rect 24382 397538 24466 397774
rect 24702 397538 24734 397774
rect 24114 397454 24734 397538
rect 24114 397218 24146 397454
rect 24382 397218 24466 397454
rect 24702 397218 24734 397454
rect 24114 360574 24734 397218
rect 24114 360338 24146 360574
rect 24382 360338 24466 360574
rect 24702 360338 24734 360574
rect 24114 360254 24734 360338
rect 24114 360018 24146 360254
rect 24382 360018 24466 360254
rect 24702 360018 24734 360254
rect 24114 323374 24734 360018
rect 24114 323138 24146 323374
rect 24382 323138 24466 323374
rect 24702 323138 24734 323374
rect 24114 323054 24734 323138
rect 24114 322818 24146 323054
rect 24382 322818 24466 323054
rect 24702 322818 24734 323054
rect 24114 286174 24734 322818
rect 24114 285938 24146 286174
rect 24382 285938 24466 286174
rect 24702 285938 24734 286174
rect 24114 285854 24734 285938
rect 24114 285618 24146 285854
rect 24382 285618 24466 285854
rect 24702 285618 24734 285854
rect 24114 248974 24734 285618
rect 24114 248738 24146 248974
rect 24382 248738 24466 248974
rect 24702 248738 24734 248974
rect 24114 248654 24734 248738
rect 24114 248418 24146 248654
rect 24382 248418 24466 248654
rect 24702 248418 24734 248654
rect 24114 211774 24734 248418
rect 24114 211538 24146 211774
rect 24382 211538 24466 211774
rect 24702 211538 24734 211774
rect 24114 211454 24734 211538
rect 24114 211218 24146 211454
rect 24382 211218 24466 211454
rect 24702 211218 24734 211454
rect 24114 174574 24734 211218
rect 24114 174338 24146 174574
rect 24382 174338 24466 174574
rect 24702 174338 24734 174574
rect 24114 174254 24734 174338
rect 24114 174018 24146 174254
rect 24382 174018 24466 174254
rect 24702 174018 24734 174254
rect 24114 137374 24734 174018
rect 24114 137138 24146 137374
rect 24382 137138 24466 137374
rect 24702 137138 24734 137374
rect 24114 137054 24734 137138
rect 24114 136818 24146 137054
rect 24382 136818 24466 137054
rect 24702 136818 24734 137054
rect 24114 100174 24734 136818
rect 24114 99938 24146 100174
rect 24382 99938 24466 100174
rect 24702 99938 24734 100174
rect 24114 99854 24734 99938
rect 24114 99618 24146 99854
rect 24382 99618 24466 99854
rect 24702 99618 24734 99854
rect 24114 62974 24734 99618
rect 24114 62738 24146 62974
rect 24382 62738 24466 62974
rect 24702 62738 24734 62974
rect 24114 62654 24734 62738
rect 24114 62418 24146 62654
rect 24382 62418 24466 62654
rect 24702 62418 24734 62654
rect 24114 25774 24734 62418
rect 24114 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 24734 25774
rect 24114 25454 24734 25538
rect 24114 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 24734 25454
rect 24114 2176 24734 25218
rect 27834 699094 28454 701760
rect 27834 698858 27866 699094
rect 28102 698858 28186 699094
rect 28422 698858 28454 699094
rect 27834 698774 28454 698858
rect 27834 698538 27866 698774
rect 28102 698538 28186 698774
rect 28422 698538 28454 698774
rect 27834 661894 28454 698538
rect 27834 661658 27866 661894
rect 28102 661658 28186 661894
rect 28422 661658 28454 661894
rect 27834 661574 28454 661658
rect 27834 661338 27866 661574
rect 28102 661338 28186 661574
rect 28422 661338 28454 661574
rect 27834 624694 28454 661338
rect 27834 624458 27866 624694
rect 28102 624458 28186 624694
rect 28422 624458 28454 624694
rect 27834 624374 28454 624458
rect 27834 624138 27866 624374
rect 28102 624138 28186 624374
rect 28422 624138 28454 624374
rect 27834 587494 28454 624138
rect 27834 587258 27866 587494
rect 28102 587258 28186 587494
rect 28422 587258 28454 587494
rect 27834 587174 28454 587258
rect 27834 586938 27866 587174
rect 28102 586938 28186 587174
rect 28422 586938 28454 587174
rect 27834 550294 28454 586938
rect 27834 550058 27866 550294
rect 28102 550058 28186 550294
rect 28422 550058 28454 550294
rect 27834 549974 28454 550058
rect 27834 549738 27866 549974
rect 28102 549738 28186 549974
rect 28422 549738 28454 549974
rect 27834 513094 28454 549738
rect 27834 512858 27866 513094
rect 28102 512858 28186 513094
rect 28422 512858 28454 513094
rect 27834 512774 28454 512858
rect 27834 512538 27866 512774
rect 28102 512538 28186 512774
rect 28422 512538 28454 512774
rect 27834 475894 28454 512538
rect 27834 475658 27866 475894
rect 28102 475658 28186 475894
rect 28422 475658 28454 475894
rect 27834 475574 28454 475658
rect 27834 475338 27866 475574
rect 28102 475338 28186 475574
rect 28422 475338 28454 475574
rect 27834 438694 28454 475338
rect 27834 438458 27866 438694
rect 28102 438458 28186 438694
rect 28422 438458 28454 438694
rect 27834 438374 28454 438458
rect 27834 438138 27866 438374
rect 28102 438138 28186 438374
rect 28422 438138 28454 438374
rect 27834 401494 28454 438138
rect 27834 401258 27866 401494
rect 28102 401258 28186 401494
rect 28422 401258 28454 401494
rect 27834 401174 28454 401258
rect 27834 400938 27866 401174
rect 28102 400938 28186 401174
rect 28422 400938 28454 401174
rect 27834 364294 28454 400938
rect 27834 364058 27866 364294
rect 28102 364058 28186 364294
rect 28422 364058 28454 364294
rect 27834 363974 28454 364058
rect 27834 363738 27866 363974
rect 28102 363738 28186 363974
rect 28422 363738 28454 363974
rect 27834 327094 28454 363738
rect 27834 326858 27866 327094
rect 28102 326858 28186 327094
rect 28422 326858 28454 327094
rect 27834 326774 28454 326858
rect 27834 326538 27866 326774
rect 28102 326538 28186 326774
rect 28422 326538 28454 326774
rect 27834 289894 28454 326538
rect 27834 289658 27866 289894
rect 28102 289658 28186 289894
rect 28422 289658 28454 289894
rect 27834 289574 28454 289658
rect 27834 289338 27866 289574
rect 28102 289338 28186 289574
rect 28422 289338 28454 289574
rect 27834 252694 28454 289338
rect 27834 252458 27866 252694
rect 28102 252458 28186 252694
rect 28422 252458 28454 252694
rect 27834 252374 28454 252458
rect 27834 252138 27866 252374
rect 28102 252138 28186 252374
rect 28422 252138 28454 252374
rect 27834 215494 28454 252138
rect 27834 215258 27866 215494
rect 28102 215258 28186 215494
rect 28422 215258 28454 215494
rect 27834 215174 28454 215258
rect 27834 214938 27866 215174
rect 28102 214938 28186 215174
rect 28422 214938 28454 215174
rect 27834 178294 28454 214938
rect 27834 178058 27866 178294
rect 28102 178058 28186 178294
rect 28422 178058 28454 178294
rect 27834 177974 28454 178058
rect 27834 177738 27866 177974
rect 28102 177738 28186 177974
rect 28422 177738 28454 177974
rect 27834 141094 28454 177738
rect 27834 140858 27866 141094
rect 28102 140858 28186 141094
rect 28422 140858 28454 141094
rect 27834 140774 28454 140858
rect 27834 140538 27866 140774
rect 28102 140538 28186 140774
rect 28422 140538 28454 140774
rect 27834 103894 28454 140538
rect 27834 103658 27866 103894
rect 28102 103658 28186 103894
rect 28422 103658 28454 103894
rect 27834 103574 28454 103658
rect 27834 103338 27866 103574
rect 28102 103338 28186 103574
rect 28422 103338 28454 103574
rect 27834 66694 28454 103338
rect 27834 66458 27866 66694
rect 28102 66458 28186 66694
rect 28422 66458 28454 66694
rect 27834 66374 28454 66458
rect 27834 66138 27866 66374
rect 28102 66138 28186 66374
rect 28422 66138 28454 66374
rect 27834 29494 28454 66138
rect 27834 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 28454 29494
rect 27834 29174 28454 29258
rect 27834 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 28454 29174
rect 27834 2176 28454 28938
rect 38994 673054 39614 701760
rect 38994 672818 39026 673054
rect 39262 672818 39346 673054
rect 39582 672818 39614 673054
rect 38994 672734 39614 672818
rect 38994 672498 39026 672734
rect 39262 672498 39346 672734
rect 39582 672498 39614 672734
rect 38994 635854 39614 672498
rect 38994 635618 39026 635854
rect 39262 635618 39346 635854
rect 39582 635618 39614 635854
rect 38994 635534 39614 635618
rect 38994 635298 39026 635534
rect 39262 635298 39346 635534
rect 39582 635298 39614 635534
rect 38994 598654 39614 635298
rect 38994 598418 39026 598654
rect 39262 598418 39346 598654
rect 39582 598418 39614 598654
rect 38994 598334 39614 598418
rect 38994 598098 39026 598334
rect 39262 598098 39346 598334
rect 39582 598098 39614 598334
rect 38994 561454 39614 598098
rect 38994 561218 39026 561454
rect 39262 561218 39346 561454
rect 39582 561218 39614 561454
rect 38994 561134 39614 561218
rect 38994 560898 39026 561134
rect 39262 560898 39346 561134
rect 39582 560898 39614 561134
rect 38994 524254 39614 560898
rect 38994 524018 39026 524254
rect 39262 524018 39346 524254
rect 39582 524018 39614 524254
rect 38994 523934 39614 524018
rect 38994 523698 39026 523934
rect 39262 523698 39346 523934
rect 39582 523698 39614 523934
rect 38994 487054 39614 523698
rect 38994 486818 39026 487054
rect 39262 486818 39346 487054
rect 39582 486818 39614 487054
rect 38994 486734 39614 486818
rect 38994 486498 39026 486734
rect 39262 486498 39346 486734
rect 39582 486498 39614 486734
rect 38994 449854 39614 486498
rect 38994 449618 39026 449854
rect 39262 449618 39346 449854
rect 39582 449618 39614 449854
rect 38994 449534 39614 449618
rect 38994 449298 39026 449534
rect 39262 449298 39346 449534
rect 39582 449298 39614 449534
rect 38994 412654 39614 449298
rect 38994 412418 39026 412654
rect 39262 412418 39346 412654
rect 39582 412418 39614 412654
rect 38994 412334 39614 412418
rect 38994 412098 39026 412334
rect 39262 412098 39346 412334
rect 39582 412098 39614 412334
rect 38994 375454 39614 412098
rect 38994 375218 39026 375454
rect 39262 375218 39346 375454
rect 39582 375218 39614 375454
rect 38994 375134 39614 375218
rect 38994 374898 39026 375134
rect 39262 374898 39346 375134
rect 39582 374898 39614 375134
rect 38994 338254 39614 374898
rect 38994 338018 39026 338254
rect 39262 338018 39346 338254
rect 39582 338018 39614 338254
rect 38994 337934 39614 338018
rect 38994 337698 39026 337934
rect 39262 337698 39346 337934
rect 39582 337698 39614 337934
rect 38994 301054 39614 337698
rect 38994 300818 39026 301054
rect 39262 300818 39346 301054
rect 39582 300818 39614 301054
rect 38994 300734 39614 300818
rect 38994 300498 39026 300734
rect 39262 300498 39346 300734
rect 39582 300498 39614 300734
rect 38994 263854 39614 300498
rect 38994 263618 39026 263854
rect 39262 263618 39346 263854
rect 39582 263618 39614 263854
rect 38994 263534 39614 263618
rect 38994 263298 39026 263534
rect 39262 263298 39346 263534
rect 39582 263298 39614 263534
rect 38994 226654 39614 263298
rect 38994 226418 39026 226654
rect 39262 226418 39346 226654
rect 39582 226418 39614 226654
rect 38994 226334 39614 226418
rect 38994 226098 39026 226334
rect 39262 226098 39346 226334
rect 39582 226098 39614 226334
rect 38994 189454 39614 226098
rect 38994 189218 39026 189454
rect 39262 189218 39346 189454
rect 39582 189218 39614 189454
rect 38994 189134 39614 189218
rect 38994 188898 39026 189134
rect 39262 188898 39346 189134
rect 39582 188898 39614 189134
rect 38994 152254 39614 188898
rect 38994 152018 39026 152254
rect 39262 152018 39346 152254
rect 39582 152018 39614 152254
rect 38994 151934 39614 152018
rect 38994 151698 39026 151934
rect 39262 151698 39346 151934
rect 39582 151698 39614 151934
rect 38994 115054 39614 151698
rect 38994 114818 39026 115054
rect 39262 114818 39346 115054
rect 39582 114818 39614 115054
rect 38994 114734 39614 114818
rect 38994 114498 39026 114734
rect 39262 114498 39346 114734
rect 39582 114498 39614 114734
rect 38994 77854 39614 114498
rect 38994 77618 39026 77854
rect 39262 77618 39346 77854
rect 39582 77618 39614 77854
rect 38994 77534 39614 77618
rect 38994 77298 39026 77534
rect 39262 77298 39346 77534
rect 39582 77298 39614 77534
rect 38994 40654 39614 77298
rect 38994 40418 39026 40654
rect 39262 40418 39346 40654
rect 39582 40418 39614 40654
rect 38994 40334 39614 40418
rect 38994 40098 39026 40334
rect 39262 40098 39346 40334
rect 39582 40098 39614 40334
rect 38994 3454 39614 40098
rect 38994 3218 39026 3454
rect 39262 3218 39346 3454
rect 39582 3218 39614 3454
rect 38994 3134 39614 3218
rect 38994 2898 39026 3134
rect 39262 2898 39346 3134
rect 39582 2898 39614 3134
rect 38994 2176 39614 2898
rect 42714 676774 43334 701760
rect 42714 676538 42746 676774
rect 42982 676538 43066 676774
rect 43302 676538 43334 676774
rect 42714 676454 43334 676538
rect 42714 676218 42746 676454
rect 42982 676218 43066 676454
rect 43302 676218 43334 676454
rect 42714 639574 43334 676218
rect 42714 639338 42746 639574
rect 42982 639338 43066 639574
rect 43302 639338 43334 639574
rect 42714 639254 43334 639338
rect 42714 639018 42746 639254
rect 42982 639018 43066 639254
rect 43302 639018 43334 639254
rect 42714 602374 43334 639018
rect 42714 602138 42746 602374
rect 42982 602138 43066 602374
rect 43302 602138 43334 602374
rect 42714 602054 43334 602138
rect 42714 601818 42746 602054
rect 42982 601818 43066 602054
rect 43302 601818 43334 602054
rect 42714 565174 43334 601818
rect 42714 564938 42746 565174
rect 42982 564938 43066 565174
rect 43302 564938 43334 565174
rect 42714 564854 43334 564938
rect 42714 564618 42746 564854
rect 42982 564618 43066 564854
rect 43302 564618 43334 564854
rect 42714 527974 43334 564618
rect 42714 527738 42746 527974
rect 42982 527738 43066 527974
rect 43302 527738 43334 527974
rect 42714 527654 43334 527738
rect 42714 527418 42746 527654
rect 42982 527418 43066 527654
rect 43302 527418 43334 527654
rect 42714 490774 43334 527418
rect 42714 490538 42746 490774
rect 42982 490538 43066 490774
rect 43302 490538 43334 490774
rect 42714 490454 43334 490538
rect 42714 490218 42746 490454
rect 42982 490218 43066 490454
rect 43302 490218 43334 490454
rect 42714 453574 43334 490218
rect 42714 453338 42746 453574
rect 42982 453338 43066 453574
rect 43302 453338 43334 453574
rect 42714 453254 43334 453338
rect 42714 453018 42746 453254
rect 42982 453018 43066 453254
rect 43302 453018 43334 453254
rect 42714 416374 43334 453018
rect 42714 416138 42746 416374
rect 42982 416138 43066 416374
rect 43302 416138 43334 416374
rect 42714 416054 43334 416138
rect 42714 415818 42746 416054
rect 42982 415818 43066 416054
rect 43302 415818 43334 416054
rect 42714 379174 43334 415818
rect 42714 378938 42746 379174
rect 42982 378938 43066 379174
rect 43302 378938 43334 379174
rect 42714 378854 43334 378938
rect 42714 378618 42746 378854
rect 42982 378618 43066 378854
rect 43302 378618 43334 378854
rect 42714 341974 43334 378618
rect 42714 341738 42746 341974
rect 42982 341738 43066 341974
rect 43302 341738 43334 341974
rect 42714 341654 43334 341738
rect 42714 341418 42746 341654
rect 42982 341418 43066 341654
rect 43302 341418 43334 341654
rect 42714 304774 43334 341418
rect 42714 304538 42746 304774
rect 42982 304538 43066 304774
rect 43302 304538 43334 304774
rect 42714 304454 43334 304538
rect 42714 304218 42746 304454
rect 42982 304218 43066 304454
rect 43302 304218 43334 304454
rect 42714 267574 43334 304218
rect 42714 267338 42746 267574
rect 42982 267338 43066 267574
rect 43302 267338 43334 267574
rect 42714 267254 43334 267338
rect 42714 267018 42746 267254
rect 42982 267018 43066 267254
rect 43302 267018 43334 267254
rect 42714 230374 43334 267018
rect 42714 230138 42746 230374
rect 42982 230138 43066 230374
rect 43302 230138 43334 230374
rect 42714 230054 43334 230138
rect 42714 229818 42746 230054
rect 42982 229818 43066 230054
rect 43302 229818 43334 230054
rect 42714 193174 43334 229818
rect 42714 192938 42746 193174
rect 42982 192938 43066 193174
rect 43302 192938 43334 193174
rect 42714 192854 43334 192938
rect 42714 192618 42746 192854
rect 42982 192618 43066 192854
rect 43302 192618 43334 192854
rect 42714 155974 43334 192618
rect 42714 155738 42746 155974
rect 42982 155738 43066 155974
rect 43302 155738 43334 155974
rect 42714 155654 43334 155738
rect 42714 155418 42746 155654
rect 42982 155418 43066 155654
rect 43302 155418 43334 155654
rect 42714 118774 43334 155418
rect 42714 118538 42746 118774
rect 42982 118538 43066 118774
rect 43302 118538 43334 118774
rect 42714 118454 43334 118538
rect 42714 118218 42746 118454
rect 42982 118218 43066 118454
rect 43302 118218 43334 118454
rect 42714 81574 43334 118218
rect 42714 81338 42746 81574
rect 42982 81338 43066 81574
rect 43302 81338 43334 81574
rect 42714 81254 43334 81338
rect 42714 81018 42746 81254
rect 42982 81018 43066 81254
rect 43302 81018 43334 81254
rect 42714 44374 43334 81018
rect 42714 44138 42746 44374
rect 42982 44138 43066 44374
rect 43302 44138 43334 44374
rect 42714 44054 43334 44138
rect 42714 43818 42746 44054
rect 42982 43818 43066 44054
rect 43302 43818 43334 44054
rect 42714 7174 43334 43818
rect 42714 6938 42746 7174
rect 42982 6938 43066 7174
rect 43302 6938 43334 7174
rect 42714 6854 43334 6938
rect 42714 6618 42746 6854
rect 42982 6618 43066 6854
rect 43302 6618 43334 6854
rect 42714 2176 43334 6618
rect 46434 680494 47054 701760
rect 46434 680258 46466 680494
rect 46702 680258 46786 680494
rect 47022 680258 47054 680494
rect 46434 680174 47054 680258
rect 46434 679938 46466 680174
rect 46702 679938 46786 680174
rect 47022 679938 47054 680174
rect 46434 643294 47054 679938
rect 46434 643058 46466 643294
rect 46702 643058 46786 643294
rect 47022 643058 47054 643294
rect 46434 642974 47054 643058
rect 46434 642738 46466 642974
rect 46702 642738 46786 642974
rect 47022 642738 47054 642974
rect 46434 606094 47054 642738
rect 46434 605858 46466 606094
rect 46702 605858 46786 606094
rect 47022 605858 47054 606094
rect 46434 605774 47054 605858
rect 46434 605538 46466 605774
rect 46702 605538 46786 605774
rect 47022 605538 47054 605774
rect 46434 568894 47054 605538
rect 46434 568658 46466 568894
rect 46702 568658 46786 568894
rect 47022 568658 47054 568894
rect 46434 568574 47054 568658
rect 46434 568338 46466 568574
rect 46702 568338 46786 568574
rect 47022 568338 47054 568574
rect 46434 531694 47054 568338
rect 46434 531458 46466 531694
rect 46702 531458 46786 531694
rect 47022 531458 47054 531694
rect 46434 531374 47054 531458
rect 46434 531138 46466 531374
rect 46702 531138 46786 531374
rect 47022 531138 47054 531374
rect 46434 494494 47054 531138
rect 46434 494258 46466 494494
rect 46702 494258 46786 494494
rect 47022 494258 47054 494494
rect 46434 494174 47054 494258
rect 46434 493938 46466 494174
rect 46702 493938 46786 494174
rect 47022 493938 47054 494174
rect 46434 457294 47054 493938
rect 46434 457058 46466 457294
rect 46702 457058 46786 457294
rect 47022 457058 47054 457294
rect 46434 456974 47054 457058
rect 46434 456738 46466 456974
rect 46702 456738 46786 456974
rect 47022 456738 47054 456974
rect 46434 420094 47054 456738
rect 46434 419858 46466 420094
rect 46702 419858 46786 420094
rect 47022 419858 47054 420094
rect 46434 419774 47054 419858
rect 46434 419538 46466 419774
rect 46702 419538 46786 419774
rect 47022 419538 47054 419774
rect 46434 382894 47054 419538
rect 46434 382658 46466 382894
rect 46702 382658 46786 382894
rect 47022 382658 47054 382894
rect 46434 382574 47054 382658
rect 46434 382338 46466 382574
rect 46702 382338 46786 382574
rect 47022 382338 47054 382574
rect 46434 345694 47054 382338
rect 46434 345458 46466 345694
rect 46702 345458 46786 345694
rect 47022 345458 47054 345694
rect 46434 345374 47054 345458
rect 46434 345138 46466 345374
rect 46702 345138 46786 345374
rect 47022 345138 47054 345374
rect 46434 308494 47054 345138
rect 46434 308258 46466 308494
rect 46702 308258 46786 308494
rect 47022 308258 47054 308494
rect 46434 308174 47054 308258
rect 46434 307938 46466 308174
rect 46702 307938 46786 308174
rect 47022 307938 47054 308174
rect 46434 271294 47054 307938
rect 46434 271058 46466 271294
rect 46702 271058 46786 271294
rect 47022 271058 47054 271294
rect 46434 270974 47054 271058
rect 46434 270738 46466 270974
rect 46702 270738 46786 270974
rect 47022 270738 47054 270974
rect 46434 234094 47054 270738
rect 46434 233858 46466 234094
rect 46702 233858 46786 234094
rect 47022 233858 47054 234094
rect 46434 233774 47054 233858
rect 46434 233538 46466 233774
rect 46702 233538 46786 233774
rect 47022 233538 47054 233774
rect 46434 196894 47054 233538
rect 46434 196658 46466 196894
rect 46702 196658 46786 196894
rect 47022 196658 47054 196894
rect 46434 196574 47054 196658
rect 46434 196338 46466 196574
rect 46702 196338 46786 196574
rect 47022 196338 47054 196574
rect 46434 159694 47054 196338
rect 46434 159458 46466 159694
rect 46702 159458 46786 159694
rect 47022 159458 47054 159694
rect 46434 159374 47054 159458
rect 46434 159138 46466 159374
rect 46702 159138 46786 159374
rect 47022 159138 47054 159374
rect 46434 122494 47054 159138
rect 46434 122258 46466 122494
rect 46702 122258 46786 122494
rect 47022 122258 47054 122494
rect 46434 122174 47054 122258
rect 46434 121938 46466 122174
rect 46702 121938 46786 122174
rect 47022 121938 47054 122174
rect 46434 85294 47054 121938
rect 46434 85058 46466 85294
rect 46702 85058 46786 85294
rect 47022 85058 47054 85294
rect 46434 84974 47054 85058
rect 46434 84738 46466 84974
rect 46702 84738 46786 84974
rect 47022 84738 47054 84974
rect 46434 48094 47054 84738
rect 46434 47858 46466 48094
rect 46702 47858 46786 48094
rect 47022 47858 47054 48094
rect 46434 47774 47054 47858
rect 46434 47538 46466 47774
rect 46702 47538 46786 47774
rect 47022 47538 47054 47774
rect 46434 10894 47054 47538
rect 46434 10658 46466 10894
rect 46702 10658 46786 10894
rect 47022 10658 47054 10894
rect 46434 10574 47054 10658
rect 46434 10338 46466 10574
rect 46702 10338 46786 10574
rect 47022 10338 47054 10574
rect 46434 2176 47054 10338
rect 50154 684214 50774 701760
rect 50154 683978 50186 684214
rect 50422 683978 50506 684214
rect 50742 683978 50774 684214
rect 50154 683894 50774 683978
rect 50154 683658 50186 683894
rect 50422 683658 50506 683894
rect 50742 683658 50774 683894
rect 50154 647014 50774 683658
rect 50154 646778 50186 647014
rect 50422 646778 50506 647014
rect 50742 646778 50774 647014
rect 50154 646694 50774 646778
rect 50154 646458 50186 646694
rect 50422 646458 50506 646694
rect 50742 646458 50774 646694
rect 50154 609814 50774 646458
rect 50154 609578 50186 609814
rect 50422 609578 50506 609814
rect 50742 609578 50774 609814
rect 50154 609494 50774 609578
rect 50154 609258 50186 609494
rect 50422 609258 50506 609494
rect 50742 609258 50774 609494
rect 50154 572614 50774 609258
rect 50154 572378 50186 572614
rect 50422 572378 50506 572614
rect 50742 572378 50774 572614
rect 50154 572294 50774 572378
rect 50154 572058 50186 572294
rect 50422 572058 50506 572294
rect 50742 572058 50774 572294
rect 50154 535414 50774 572058
rect 50154 535178 50186 535414
rect 50422 535178 50506 535414
rect 50742 535178 50774 535414
rect 50154 535094 50774 535178
rect 50154 534858 50186 535094
rect 50422 534858 50506 535094
rect 50742 534858 50774 535094
rect 50154 498214 50774 534858
rect 50154 497978 50186 498214
rect 50422 497978 50506 498214
rect 50742 497978 50774 498214
rect 50154 497894 50774 497978
rect 50154 497658 50186 497894
rect 50422 497658 50506 497894
rect 50742 497658 50774 497894
rect 50154 461014 50774 497658
rect 50154 460778 50186 461014
rect 50422 460778 50506 461014
rect 50742 460778 50774 461014
rect 50154 460694 50774 460778
rect 50154 460458 50186 460694
rect 50422 460458 50506 460694
rect 50742 460458 50774 460694
rect 50154 423814 50774 460458
rect 50154 423578 50186 423814
rect 50422 423578 50506 423814
rect 50742 423578 50774 423814
rect 50154 423494 50774 423578
rect 50154 423258 50186 423494
rect 50422 423258 50506 423494
rect 50742 423258 50774 423494
rect 50154 386614 50774 423258
rect 50154 386378 50186 386614
rect 50422 386378 50506 386614
rect 50742 386378 50774 386614
rect 50154 386294 50774 386378
rect 50154 386058 50186 386294
rect 50422 386058 50506 386294
rect 50742 386058 50774 386294
rect 50154 349414 50774 386058
rect 50154 349178 50186 349414
rect 50422 349178 50506 349414
rect 50742 349178 50774 349414
rect 50154 349094 50774 349178
rect 50154 348858 50186 349094
rect 50422 348858 50506 349094
rect 50742 348858 50774 349094
rect 50154 312214 50774 348858
rect 50154 311978 50186 312214
rect 50422 311978 50506 312214
rect 50742 311978 50774 312214
rect 50154 311894 50774 311978
rect 50154 311658 50186 311894
rect 50422 311658 50506 311894
rect 50742 311658 50774 311894
rect 50154 275014 50774 311658
rect 50154 274778 50186 275014
rect 50422 274778 50506 275014
rect 50742 274778 50774 275014
rect 50154 274694 50774 274778
rect 50154 274458 50186 274694
rect 50422 274458 50506 274694
rect 50742 274458 50774 274694
rect 50154 237814 50774 274458
rect 50154 237578 50186 237814
rect 50422 237578 50506 237814
rect 50742 237578 50774 237814
rect 50154 237494 50774 237578
rect 50154 237258 50186 237494
rect 50422 237258 50506 237494
rect 50742 237258 50774 237494
rect 50154 200614 50774 237258
rect 50154 200378 50186 200614
rect 50422 200378 50506 200614
rect 50742 200378 50774 200614
rect 50154 200294 50774 200378
rect 50154 200058 50186 200294
rect 50422 200058 50506 200294
rect 50742 200058 50774 200294
rect 50154 163414 50774 200058
rect 50154 163178 50186 163414
rect 50422 163178 50506 163414
rect 50742 163178 50774 163414
rect 50154 163094 50774 163178
rect 50154 162858 50186 163094
rect 50422 162858 50506 163094
rect 50742 162858 50774 163094
rect 50154 126214 50774 162858
rect 50154 125978 50186 126214
rect 50422 125978 50506 126214
rect 50742 125978 50774 126214
rect 50154 125894 50774 125978
rect 50154 125658 50186 125894
rect 50422 125658 50506 125894
rect 50742 125658 50774 125894
rect 50154 89014 50774 125658
rect 50154 88778 50186 89014
rect 50422 88778 50506 89014
rect 50742 88778 50774 89014
rect 50154 88694 50774 88778
rect 50154 88458 50186 88694
rect 50422 88458 50506 88694
rect 50742 88458 50774 88694
rect 50154 51814 50774 88458
rect 50154 51578 50186 51814
rect 50422 51578 50506 51814
rect 50742 51578 50774 51814
rect 50154 51494 50774 51578
rect 50154 51258 50186 51494
rect 50422 51258 50506 51494
rect 50742 51258 50774 51494
rect 50154 14614 50774 51258
rect 50154 14378 50186 14614
rect 50422 14378 50506 14614
rect 50742 14378 50774 14614
rect 50154 14294 50774 14378
rect 50154 14058 50186 14294
rect 50422 14058 50506 14294
rect 50742 14058 50774 14294
rect 50154 2176 50774 14058
rect 53874 687934 54494 701760
rect 53874 687698 53906 687934
rect 54142 687698 54226 687934
rect 54462 687698 54494 687934
rect 53874 687614 54494 687698
rect 53874 687378 53906 687614
rect 54142 687378 54226 687614
rect 54462 687378 54494 687614
rect 53874 650734 54494 687378
rect 53874 650498 53906 650734
rect 54142 650498 54226 650734
rect 54462 650498 54494 650734
rect 53874 650414 54494 650498
rect 53874 650178 53906 650414
rect 54142 650178 54226 650414
rect 54462 650178 54494 650414
rect 53874 613534 54494 650178
rect 53874 613298 53906 613534
rect 54142 613298 54226 613534
rect 54462 613298 54494 613534
rect 53874 613214 54494 613298
rect 53874 612978 53906 613214
rect 54142 612978 54226 613214
rect 54462 612978 54494 613214
rect 53874 576334 54494 612978
rect 53874 576098 53906 576334
rect 54142 576098 54226 576334
rect 54462 576098 54494 576334
rect 53874 576014 54494 576098
rect 53874 575778 53906 576014
rect 54142 575778 54226 576014
rect 54462 575778 54494 576014
rect 53874 539134 54494 575778
rect 53874 538898 53906 539134
rect 54142 538898 54226 539134
rect 54462 538898 54494 539134
rect 53874 538814 54494 538898
rect 53874 538578 53906 538814
rect 54142 538578 54226 538814
rect 54462 538578 54494 538814
rect 53874 501934 54494 538578
rect 53874 501698 53906 501934
rect 54142 501698 54226 501934
rect 54462 501698 54494 501934
rect 53874 501614 54494 501698
rect 53874 501378 53906 501614
rect 54142 501378 54226 501614
rect 54462 501378 54494 501614
rect 53874 464734 54494 501378
rect 53874 464498 53906 464734
rect 54142 464498 54226 464734
rect 54462 464498 54494 464734
rect 53874 464414 54494 464498
rect 53874 464178 53906 464414
rect 54142 464178 54226 464414
rect 54462 464178 54494 464414
rect 53874 427534 54494 464178
rect 53874 427298 53906 427534
rect 54142 427298 54226 427534
rect 54462 427298 54494 427534
rect 53874 427214 54494 427298
rect 53874 426978 53906 427214
rect 54142 426978 54226 427214
rect 54462 426978 54494 427214
rect 53874 390334 54494 426978
rect 53874 390098 53906 390334
rect 54142 390098 54226 390334
rect 54462 390098 54494 390334
rect 53874 390014 54494 390098
rect 53874 389778 53906 390014
rect 54142 389778 54226 390014
rect 54462 389778 54494 390014
rect 53874 353134 54494 389778
rect 53874 352898 53906 353134
rect 54142 352898 54226 353134
rect 54462 352898 54494 353134
rect 53874 352814 54494 352898
rect 53874 352578 53906 352814
rect 54142 352578 54226 352814
rect 54462 352578 54494 352814
rect 53874 315934 54494 352578
rect 53874 315698 53906 315934
rect 54142 315698 54226 315934
rect 54462 315698 54494 315934
rect 53874 315614 54494 315698
rect 53874 315378 53906 315614
rect 54142 315378 54226 315614
rect 54462 315378 54494 315614
rect 53874 278734 54494 315378
rect 53874 278498 53906 278734
rect 54142 278498 54226 278734
rect 54462 278498 54494 278734
rect 53874 278414 54494 278498
rect 53874 278178 53906 278414
rect 54142 278178 54226 278414
rect 54462 278178 54494 278414
rect 53874 241534 54494 278178
rect 53874 241298 53906 241534
rect 54142 241298 54226 241534
rect 54462 241298 54494 241534
rect 53874 241214 54494 241298
rect 53874 240978 53906 241214
rect 54142 240978 54226 241214
rect 54462 240978 54494 241214
rect 53874 204334 54494 240978
rect 53874 204098 53906 204334
rect 54142 204098 54226 204334
rect 54462 204098 54494 204334
rect 53874 204014 54494 204098
rect 53874 203778 53906 204014
rect 54142 203778 54226 204014
rect 54462 203778 54494 204014
rect 53874 167134 54494 203778
rect 53874 166898 53906 167134
rect 54142 166898 54226 167134
rect 54462 166898 54494 167134
rect 53874 166814 54494 166898
rect 53874 166578 53906 166814
rect 54142 166578 54226 166814
rect 54462 166578 54494 166814
rect 53874 129934 54494 166578
rect 53874 129698 53906 129934
rect 54142 129698 54226 129934
rect 54462 129698 54494 129934
rect 53874 129614 54494 129698
rect 53874 129378 53906 129614
rect 54142 129378 54226 129614
rect 54462 129378 54494 129614
rect 53874 92734 54494 129378
rect 53874 92498 53906 92734
rect 54142 92498 54226 92734
rect 54462 92498 54494 92734
rect 53874 92414 54494 92498
rect 53874 92178 53906 92414
rect 54142 92178 54226 92414
rect 54462 92178 54494 92414
rect 53874 55534 54494 92178
rect 53874 55298 53906 55534
rect 54142 55298 54226 55534
rect 54462 55298 54494 55534
rect 53874 55214 54494 55298
rect 53874 54978 53906 55214
rect 54142 54978 54226 55214
rect 54462 54978 54494 55214
rect 53874 18334 54494 54978
rect 53874 18098 53906 18334
rect 54142 18098 54226 18334
rect 54462 18098 54494 18334
rect 53874 18014 54494 18098
rect 53874 17778 53906 18014
rect 54142 17778 54226 18014
rect 54462 17778 54494 18014
rect 53874 2176 54494 17778
rect 57594 691654 58214 701760
rect 57594 691418 57626 691654
rect 57862 691418 57946 691654
rect 58182 691418 58214 691654
rect 57594 691334 58214 691418
rect 57594 691098 57626 691334
rect 57862 691098 57946 691334
rect 58182 691098 58214 691334
rect 57594 654454 58214 691098
rect 57594 654218 57626 654454
rect 57862 654218 57946 654454
rect 58182 654218 58214 654454
rect 57594 654134 58214 654218
rect 57594 653898 57626 654134
rect 57862 653898 57946 654134
rect 58182 653898 58214 654134
rect 57594 617254 58214 653898
rect 57594 617018 57626 617254
rect 57862 617018 57946 617254
rect 58182 617018 58214 617254
rect 57594 616934 58214 617018
rect 57594 616698 57626 616934
rect 57862 616698 57946 616934
rect 58182 616698 58214 616934
rect 57594 580054 58214 616698
rect 57594 579818 57626 580054
rect 57862 579818 57946 580054
rect 58182 579818 58214 580054
rect 57594 579734 58214 579818
rect 57594 579498 57626 579734
rect 57862 579498 57946 579734
rect 58182 579498 58214 579734
rect 57594 542854 58214 579498
rect 57594 542618 57626 542854
rect 57862 542618 57946 542854
rect 58182 542618 58214 542854
rect 57594 542534 58214 542618
rect 57594 542298 57626 542534
rect 57862 542298 57946 542534
rect 58182 542298 58214 542534
rect 57594 505654 58214 542298
rect 57594 505418 57626 505654
rect 57862 505418 57946 505654
rect 58182 505418 58214 505654
rect 57594 505334 58214 505418
rect 57594 505098 57626 505334
rect 57862 505098 57946 505334
rect 58182 505098 58214 505334
rect 57594 468454 58214 505098
rect 57594 468218 57626 468454
rect 57862 468218 57946 468454
rect 58182 468218 58214 468454
rect 57594 468134 58214 468218
rect 57594 467898 57626 468134
rect 57862 467898 57946 468134
rect 58182 467898 58214 468134
rect 57594 431254 58214 467898
rect 57594 431018 57626 431254
rect 57862 431018 57946 431254
rect 58182 431018 58214 431254
rect 57594 430934 58214 431018
rect 57594 430698 57626 430934
rect 57862 430698 57946 430934
rect 58182 430698 58214 430934
rect 57594 394054 58214 430698
rect 57594 393818 57626 394054
rect 57862 393818 57946 394054
rect 58182 393818 58214 394054
rect 57594 393734 58214 393818
rect 57594 393498 57626 393734
rect 57862 393498 57946 393734
rect 58182 393498 58214 393734
rect 57594 356854 58214 393498
rect 57594 356618 57626 356854
rect 57862 356618 57946 356854
rect 58182 356618 58214 356854
rect 57594 356534 58214 356618
rect 57594 356298 57626 356534
rect 57862 356298 57946 356534
rect 58182 356298 58214 356534
rect 57594 319654 58214 356298
rect 57594 319418 57626 319654
rect 57862 319418 57946 319654
rect 58182 319418 58214 319654
rect 57594 319334 58214 319418
rect 57594 319098 57626 319334
rect 57862 319098 57946 319334
rect 58182 319098 58214 319334
rect 57594 282454 58214 319098
rect 57594 282218 57626 282454
rect 57862 282218 57946 282454
rect 58182 282218 58214 282454
rect 57594 282134 58214 282218
rect 57594 281898 57626 282134
rect 57862 281898 57946 282134
rect 58182 281898 58214 282134
rect 57594 245254 58214 281898
rect 57594 245018 57626 245254
rect 57862 245018 57946 245254
rect 58182 245018 58214 245254
rect 57594 244934 58214 245018
rect 57594 244698 57626 244934
rect 57862 244698 57946 244934
rect 58182 244698 58214 244934
rect 57594 208054 58214 244698
rect 57594 207818 57626 208054
rect 57862 207818 57946 208054
rect 58182 207818 58214 208054
rect 57594 207734 58214 207818
rect 57594 207498 57626 207734
rect 57862 207498 57946 207734
rect 58182 207498 58214 207734
rect 57594 170854 58214 207498
rect 57594 170618 57626 170854
rect 57862 170618 57946 170854
rect 58182 170618 58214 170854
rect 57594 170534 58214 170618
rect 57594 170298 57626 170534
rect 57862 170298 57946 170534
rect 58182 170298 58214 170534
rect 57594 133654 58214 170298
rect 57594 133418 57626 133654
rect 57862 133418 57946 133654
rect 58182 133418 58214 133654
rect 57594 133334 58214 133418
rect 57594 133098 57626 133334
rect 57862 133098 57946 133334
rect 58182 133098 58214 133334
rect 57594 96454 58214 133098
rect 57594 96218 57626 96454
rect 57862 96218 57946 96454
rect 58182 96218 58214 96454
rect 57594 96134 58214 96218
rect 57594 95898 57626 96134
rect 57862 95898 57946 96134
rect 58182 95898 58214 96134
rect 57594 59254 58214 95898
rect 57594 59018 57626 59254
rect 57862 59018 57946 59254
rect 58182 59018 58214 59254
rect 57594 58934 58214 59018
rect 57594 58698 57626 58934
rect 57862 58698 57946 58934
rect 58182 58698 58214 58934
rect 57594 22054 58214 58698
rect 57594 21818 57626 22054
rect 57862 21818 57946 22054
rect 58182 21818 58214 22054
rect 57594 21734 58214 21818
rect 57594 21498 57626 21734
rect 57862 21498 57946 21734
rect 58182 21498 58214 21734
rect 57594 2176 58214 21498
rect 61314 695374 61934 701760
rect 61314 695138 61346 695374
rect 61582 695138 61666 695374
rect 61902 695138 61934 695374
rect 61314 695054 61934 695138
rect 61314 694818 61346 695054
rect 61582 694818 61666 695054
rect 61902 694818 61934 695054
rect 61314 658174 61934 694818
rect 61314 657938 61346 658174
rect 61582 657938 61666 658174
rect 61902 657938 61934 658174
rect 61314 657854 61934 657938
rect 61314 657618 61346 657854
rect 61582 657618 61666 657854
rect 61902 657618 61934 657854
rect 61314 620974 61934 657618
rect 61314 620738 61346 620974
rect 61582 620738 61666 620974
rect 61902 620738 61934 620974
rect 61314 620654 61934 620738
rect 61314 620418 61346 620654
rect 61582 620418 61666 620654
rect 61902 620418 61934 620654
rect 61314 583774 61934 620418
rect 61314 583538 61346 583774
rect 61582 583538 61666 583774
rect 61902 583538 61934 583774
rect 61314 583454 61934 583538
rect 61314 583218 61346 583454
rect 61582 583218 61666 583454
rect 61902 583218 61934 583454
rect 61314 546574 61934 583218
rect 61314 546338 61346 546574
rect 61582 546338 61666 546574
rect 61902 546338 61934 546574
rect 61314 546254 61934 546338
rect 61314 546018 61346 546254
rect 61582 546018 61666 546254
rect 61902 546018 61934 546254
rect 61314 509374 61934 546018
rect 61314 509138 61346 509374
rect 61582 509138 61666 509374
rect 61902 509138 61934 509374
rect 61314 509054 61934 509138
rect 61314 508818 61346 509054
rect 61582 508818 61666 509054
rect 61902 508818 61934 509054
rect 61314 472174 61934 508818
rect 61314 471938 61346 472174
rect 61582 471938 61666 472174
rect 61902 471938 61934 472174
rect 61314 471854 61934 471938
rect 61314 471618 61346 471854
rect 61582 471618 61666 471854
rect 61902 471618 61934 471854
rect 61314 434974 61934 471618
rect 61314 434738 61346 434974
rect 61582 434738 61666 434974
rect 61902 434738 61934 434974
rect 61314 434654 61934 434738
rect 61314 434418 61346 434654
rect 61582 434418 61666 434654
rect 61902 434418 61934 434654
rect 61314 397774 61934 434418
rect 61314 397538 61346 397774
rect 61582 397538 61666 397774
rect 61902 397538 61934 397774
rect 61314 397454 61934 397538
rect 61314 397218 61346 397454
rect 61582 397218 61666 397454
rect 61902 397218 61934 397454
rect 61314 360574 61934 397218
rect 61314 360338 61346 360574
rect 61582 360338 61666 360574
rect 61902 360338 61934 360574
rect 61314 360254 61934 360338
rect 61314 360018 61346 360254
rect 61582 360018 61666 360254
rect 61902 360018 61934 360254
rect 61314 323374 61934 360018
rect 61314 323138 61346 323374
rect 61582 323138 61666 323374
rect 61902 323138 61934 323374
rect 61314 323054 61934 323138
rect 61314 322818 61346 323054
rect 61582 322818 61666 323054
rect 61902 322818 61934 323054
rect 61314 286174 61934 322818
rect 61314 285938 61346 286174
rect 61582 285938 61666 286174
rect 61902 285938 61934 286174
rect 61314 285854 61934 285938
rect 61314 285618 61346 285854
rect 61582 285618 61666 285854
rect 61902 285618 61934 285854
rect 61314 248974 61934 285618
rect 61314 248738 61346 248974
rect 61582 248738 61666 248974
rect 61902 248738 61934 248974
rect 61314 248654 61934 248738
rect 61314 248418 61346 248654
rect 61582 248418 61666 248654
rect 61902 248418 61934 248654
rect 61314 211774 61934 248418
rect 61314 211538 61346 211774
rect 61582 211538 61666 211774
rect 61902 211538 61934 211774
rect 61314 211454 61934 211538
rect 61314 211218 61346 211454
rect 61582 211218 61666 211454
rect 61902 211218 61934 211454
rect 61314 174574 61934 211218
rect 61314 174338 61346 174574
rect 61582 174338 61666 174574
rect 61902 174338 61934 174574
rect 61314 174254 61934 174338
rect 61314 174018 61346 174254
rect 61582 174018 61666 174254
rect 61902 174018 61934 174254
rect 61314 137374 61934 174018
rect 61314 137138 61346 137374
rect 61582 137138 61666 137374
rect 61902 137138 61934 137374
rect 61314 137054 61934 137138
rect 61314 136818 61346 137054
rect 61582 136818 61666 137054
rect 61902 136818 61934 137054
rect 61314 100174 61934 136818
rect 61314 99938 61346 100174
rect 61582 99938 61666 100174
rect 61902 99938 61934 100174
rect 61314 99854 61934 99938
rect 61314 99618 61346 99854
rect 61582 99618 61666 99854
rect 61902 99618 61934 99854
rect 61314 62974 61934 99618
rect 61314 62738 61346 62974
rect 61582 62738 61666 62974
rect 61902 62738 61934 62974
rect 61314 62654 61934 62738
rect 61314 62418 61346 62654
rect 61582 62418 61666 62654
rect 61902 62418 61934 62654
rect 61314 25774 61934 62418
rect 61314 25538 61346 25774
rect 61582 25538 61666 25774
rect 61902 25538 61934 25774
rect 61314 25454 61934 25538
rect 61314 25218 61346 25454
rect 61582 25218 61666 25454
rect 61902 25218 61934 25454
rect 61314 2176 61934 25218
rect 65034 699094 65654 701760
rect 65034 698858 65066 699094
rect 65302 698858 65386 699094
rect 65622 698858 65654 699094
rect 65034 698774 65654 698858
rect 65034 698538 65066 698774
rect 65302 698538 65386 698774
rect 65622 698538 65654 698774
rect 65034 661894 65654 698538
rect 65034 661658 65066 661894
rect 65302 661658 65386 661894
rect 65622 661658 65654 661894
rect 65034 661574 65654 661658
rect 65034 661338 65066 661574
rect 65302 661338 65386 661574
rect 65622 661338 65654 661574
rect 65034 624694 65654 661338
rect 65034 624458 65066 624694
rect 65302 624458 65386 624694
rect 65622 624458 65654 624694
rect 65034 624374 65654 624458
rect 65034 624138 65066 624374
rect 65302 624138 65386 624374
rect 65622 624138 65654 624374
rect 65034 587494 65654 624138
rect 65034 587258 65066 587494
rect 65302 587258 65386 587494
rect 65622 587258 65654 587494
rect 65034 587174 65654 587258
rect 65034 586938 65066 587174
rect 65302 586938 65386 587174
rect 65622 586938 65654 587174
rect 65034 550294 65654 586938
rect 65034 550058 65066 550294
rect 65302 550058 65386 550294
rect 65622 550058 65654 550294
rect 65034 549974 65654 550058
rect 65034 549738 65066 549974
rect 65302 549738 65386 549974
rect 65622 549738 65654 549974
rect 65034 513094 65654 549738
rect 65034 512858 65066 513094
rect 65302 512858 65386 513094
rect 65622 512858 65654 513094
rect 65034 512774 65654 512858
rect 65034 512538 65066 512774
rect 65302 512538 65386 512774
rect 65622 512538 65654 512774
rect 65034 475894 65654 512538
rect 65034 475658 65066 475894
rect 65302 475658 65386 475894
rect 65622 475658 65654 475894
rect 65034 475574 65654 475658
rect 65034 475338 65066 475574
rect 65302 475338 65386 475574
rect 65622 475338 65654 475574
rect 65034 438694 65654 475338
rect 65034 438458 65066 438694
rect 65302 438458 65386 438694
rect 65622 438458 65654 438694
rect 65034 438374 65654 438458
rect 65034 438138 65066 438374
rect 65302 438138 65386 438374
rect 65622 438138 65654 438374
rect 65034 401494 65654 438138
rect 65034 401258 65066 401494
rect 65302 401258 65386 401494
rect 65622 401258 65654 401494
rect 65034 401174 65654 401258
rect 65034 400938 65066 401174
rect 65302 400938 65386 401174
rect 65622 400938 65654 401174
rect 65034 364294 65654 400938
rect 65034 364058 65066 364294
rect 65302 364058 65386 364294
rect 65622 364058 65654 364294
rect 65034 363974 65654 364058
rect 65034 363738 65066 363974
rect 65302 363738 65386 363974
rect 65622 363738 65654 363974
rect 65034 327094 65654 363738
rect 65034 326858 65066 327094
rect 65302 326858 65386 327094
rect 65622 326858 65654 327094
rect 65034 326774 65654 326858
rect 65034 326538 65066 326774
rect 65302 326538 65386 326774
rect 65622 326538 65654 326774
rect 65034 289894 65654 326538
rect 65034 289658 65066 289894
rect 65302 289658 65386 289894
rect 65622 289658 65654 289894
rect 65034 289574 65654 289658
rect 65034 289338 65066 289574
rect 65302 289338 65386 289574
rect 65622 289338 65654 289574
rect 65034 252694 65654 289338
rect 65034 252458 65066 252694
rect 65302 252458 65386 252694
rect 65622 252458 65654 252694
rect 65034 252374 65654 252458
rect 65034 252138 65066 252374
rect 65302 252138 65386 252374
rect 65622 252138 65654 252374
rect 65034 215494 65654 252138
rect 65034 215258 65066 215494
rect 65302 215258 65386 215494
rect 65622 215258 65654 215494
rect 65034 215174 65654 215258
rect 65034 214938 65066 215174
rect 65302 214938 65386 215174
rect 65622 214938 65654 215174
rect 65034 178294 65654 214938
rect 65034 178058 65066 178294
rect 65302 178058 65386 178294
rect 65622 178058 65654 178294
rect 65034 177974 65654 178058
rect 65034 177738 65066 177974
rect 65302 177738 65386 177974
rect 65622 177738 65654 177974
rect 65034 141094 65654 177738
rect 65034 140858 65066 141094
rect 65302 140858 65386 141094
rect 65622 140858 65654 141094
rect 65034 140774 65654 140858
rect 65034 140538 65066 140774
rect 65302 140538 65386 140774
rect 65622 140538 65654 140774
rect 65034 103894 65654 140538
rect 65034 103658 65066 103894
rect 65302 103658 65386 103894
rect 65622 103658 65654 103894
rect 65034 103574 65654 103658
rect 65034 103338 65066 103574
rect 65302 103338 65386 103574
rect 65622 103338 65654 103574
rect 65034 66694 65654 103338
rect 65034 66458 65066 66694
rect 65302 66458 65386 66694
rect 65622 66458 65654 66694
rect 65034 66374 65654 66458
rect 65034 66138 65066 66374
rect 65302 66138 65386 66374
rect 65622 66138 65654 66374
rect 65034 29494 65654 66138
rect 65034 29258 65066 29494
rect 65302 29258 65386 29494
rect 65622 29258 65654 29494
rect 65034 29174 65654 29258
rect 65034 28938 65066 29174
rect 65302 28938 65386 29174
rect 65622 28938 65654 29174
rect 65034 2176 65654 28938
rect 76194 673054 76814 701760
rect 76194 672818 76226 673054
rect 76462 672818 76546 673054
rect 76782 672818 76814 673054
rect 76194 672734 76814 672818
rect 76194 672498 76226 672734
rect 76462 672498 76546 672734
rect 76782 672498 76814 672734
rect 76194 635854 76814 672498
rect 76194 635618 76226 635854
rect 76462 635618 76546 635854
rect 76782 635618 76814 635854
rect 76194 635534 76814 635618
rect 76194 635298 76226 635534
rect 76462 635298 76546 635534
rect 76782 635298 76814 635534
rect 76194 598654 76814 635298
rect 76194 598418 76226 598654
rect 76462 598418 76546 598654
rect 76782 598418 76814 598654
rect 76194 598334 76814 598418
rect 76194 598098 76226 598334
rect 76462 598098 76546 598334
rect 76782 598098 76814 598334
rect 76194 561454 76814 598098
rect 76194 561218 76226 561454
rect 76462 561218 76546 561454
rect 76782 561218 76814 561454
rect 76194 561134 76814 561218
rect 76194 560898 76226 561134
rect 76462 560898 76546 561134
rect 76782 560898 76814 561134
rect 76194 524254 76814 560898
rect 76194 524018 76226 524254
rect 76462 524018 76546 524254
rect 76782 524018 76814 524254
rect 76194 523934 76814 524018
rect 76194 523698 76226 523934
rect 76462 523698 76546 523934
rect 76782 523698 76814 523934
rect 76194 487054 76814 523698
rect 76194 486818 76226 487054
rect 76462 486818 76546 487054
rect 76782 486818 76814 487054
rect 76194 486734 76814 486818
rect 76194 486498 76226 486734
rect 76462 486498 76546 486734
rect 76782 486498 76814 486734
rect 76194 449854 76814 486498
rect 76194 449618 76226 449854
rect 76462 449618 76546 449854
rect 76782 449618 76814 449854
rect 76194 449534 76814 449618
rect 76194 449298 76226 449534
rect 76462 449298 76546 449534
rect 76782 449298 76814 449534
rect 76194 412654 76814 449298
rect 76194 412418 76226 412654
rect 76462 412418 76546 412654
rect 76782 412418 76814 412654
rect 76194 412334 76814 412418
rect 76194 412098 76226 412334
rect 76462 412098 76546 412334
rect 76782 412098 76814 412334
rect 76194 375454 76814 412098
rect 76194 375218 76226 375454
rect 76462 375218 76546 375454
rect 76782 375218 76814 375454
rect 76194 375134 76814 375218
rect 76194 374898 76226 375134
rect 76462 374898 76546 375134
rect 76782 374898 76814 375134
rect 76194 338254 76814 374898
rect 76194 338018 76226 338254
rect 76462 338018 76546 338254
rect 76782 338018 76814 338254
rect 76194 337934 76814 338018
rect 76194 337698 76226 337934
rect 76462 337698 76546 337934
rect 76782 337698 76814 337934
rect 76194 301054 76814 337698
rect 76194 300818 76226 301054
rect 76462 300818 76546 301054
rect 76782 300818 76814 301054
rect 76194 300734 76814 300818
rect 76194 300498 76226 300734
rect 76462 300498 76546 300734
rect 76782 300498 76814 300734
rect 76194 263854 76814 300498
rect 76194 263618 76226 263854
rect 76462 263618 76546 263854
rect 76782 263618 76814 263854
rect 76194 263534 76814 263618
rect 76194 263298 76226 263534
rect 76462 263298 76546 263534
rect 76782 263298 76814 263534
rect 76194 226654 76814 263298
rect 76194 226418 76226 226654
rect 76462 226418 76546 226654
rect 76782 226418 76814 226654
rect 76194 226334 76814 226418
rect 76194 226098 76226 226334
rect 76462 226098 76546 226334
rect 76782 226098 76814 226334
rect 76194 189454 76814 226098
rect 76194 189218 76226 189454
rect 76462 189218 76546 189454
rect 76782 189218 76814 189454
rect 76194 189134 76814 189218
rect 76194 188898 76226 189134
rect 76462 188898 76546 189134
rect 76782 188898 76814 189134
rect 76194 152254 76814 188898
rect 76194 152018 76226 152254
rect 76462 152018 76546 152254
rect 76782 152018 76814 152254
rect 76194 151934 76814 152018
rect 76194 151698 76226 151934
rect 76462 151698 76546 151934
rect 76782 151698 76814 151934
rect 76194 115054 76814 151698
rect 76194 114818 76226 115054
rect 76462 114818 76546 115054
rect 76782 114818 76814 115054
rect 76194 114734 76814 114818
rect 76194 114498 76226 114734
rect 76462 114498 76546 114734
rect 76782 114498 76814 114734
rect 76194 77854 76814 114498
rect 76194 77618 76226 77854
rect 76462 77618 76546 77854
rect 76782 77618 76814 77854
rect 76194 77534 76814 77618
rect 76194 77298 76226 77534
rect 76462 77298 76546 77534
rect 76782 77298 76814 77534
rect 76194 40654 76814 77298
rect 76194 40418 76226 40654
rect 76462 40418 76546 40654
rect 76782 40418 76814 40654
rect 76194 40334 76814 40418
rect 76194 40098 76226 40334
rect 76462 40098 76546 40334
rect 76782 40098 76814 40334
rect 76194 3454 76814 40098
rect 76194 3218 76226 3454
rect 76462 3218 76546 3454
rect 76782 3218 76814 3454
rect 76194 3134 76814 3218
rect 76194 2898 76226 3134
rect 76462 2898 76546 3134
rect 76782 2898 76814 3134
rect 76194 2176 76814 2898
rect 79914 676774 80534 701760
rect 79914 676538 79946 676774
rect 80182 676538 80266 676774
rect 80502 676538 80534 676774
rect 79914 676454 80534 676538
rect 79914 676218 79946 676454
rect 80182 676218 80266 676454
rect 80502 676218 80534 676454
rect 79914 639574 80534 676218
rect 79914 639338 79946 639574
rect 80182 639338 80266 639574
rect 80502 639338 80534 639574
rect 79914 639254 80534 639338
rect 79914 639018 79946 639254
rect 80182 639018 80266 639254
rect 80502 639018 80534 639254
rect 79914 602374 80534 639018
rect 79914 602138 79946 602374
rect 80182 602138 80266 602374
rect 80502 602138 80534 602374
rect 79914 602054 80534 602138
rect 79914 601818 79946 602054
rect 80182 601818 80266 602054
rect 80502 601818 80534 602054
rect 79914 565174 80534 601818
rect 79914 564938 79946 565174
rect 80182 564938 80266 565174
rect 80502 564938 80534 565174
rect 79914 564854 80534 564938
rect 79914 564618 79946 564854
rect 80182 564618 80266 564854
rect 80502 564618 80534 564854
rect 79914 527974 80534 564618
rect 79914 527738 79946 527974
rect 80182 527738 80266 527974
rect 80502 527738 80534 527974
rect 79914 527654 80534 527738
rect 79914 527418 79946 527654
rect 80182 527418 80266 527654
rect 80502 527418 80534 527654
rect 79914 490774 80534 527418
rect 79914 490538 79946 490774
rect 80182 490538 80266 490774
rect 80502 490538 80534 490774
rect 79914 490454 80534 490538
rect 79914 490218 79946 490454
rect 80182 490218 80266 490454
rect 80502 490218 80534 490454
rect 79914 453574 80534 490218
rect 79914 453338 79946 453574
rect 80182 453338 80266 453574
rect 80502 453338 80534 453574
rect 79914 453254 80534 453338
rect 79914 453018 79946 453254
rect 80182 453018 80266 453254
rect 80502 453018 80534 453254
rect 79914 416374 80534 453018
rect 79914 416138 79946 416374
rect 80182 416138 80266 416374
rect 80502 416138 80534 416374
rect 79914 416054 80534 416138
rect 79914 415818 79946 416054
rect 80182 415818 80266 416054
rect 80502 415818 80534 416054
rect 79914 379174 80534 415818
rect 79914 378938 79946 379174
rect 80182 378938 80266 379174
rect 80502 378938 80534 379174
rect 79914 378854 80534 378938
rect 79914 378618 79946 378854
rect 80182 378618 80266 378854
rect 80502 378618 80534 378854
rect 79914 341974 80534 378618
rect 79914 341738 79946 341974
rect 80182 341738 80266 341974
rect 80502 341738 80534 341974
rect 79914 341654 80534 341738
rect 79914 341418 79946 341654
rect 80182 341418 80266 341654
rect 80502 341418 80534 341654
rect 79914 304774 80534 341418
rect 79914 304538 79946 304774
rect 80182 304538 80266 304774
rect 80502 304538 80534 304774
rect 79914 304454 80534 304538
rect 79914 304218 79946 304454
rect 80182 304218 80266 304454
rect 80502 304218 80534 304454
rect 79914 267574 80534 304218
rect 79914 267338 79946 267574
rect 80182 267338 80266 267574
rect 80502 267338 80534 267574
rect 79914 267254 80534 267338
rect 79914 267018 79946 267254
rect 80182 267018 80266 267254
rect 80502 267018 80534 267254
rect 79914 230374 80534 267018
rect 79914 230138 79946 230374
rect 80182 230138 80266 230374
rect 80502 230138 80534 230374
rect 79914 230054 80534 230138
rect 79914 229818 79946 230054
rect 80182 229818 80266 230054
rect 80502 229818 80534 230054
rect 79914 193174 80534 229818
rect 79914 192938 79946 193174
rect 80182 192938 80266 193174
rect 80502 192938 80534 193174
rect 79914 192854 80534 192938
rect 79914 192618 79946 192854
rect 80182 192618 80266 192854
rect 80502 192618 80534 192854
rect 79914 155974 80534 192618
rect 79914 155738 79946 155974
rect 80182 155738 80266 155974
rect 80502 155738 80534 155974
rect 79914 155654 80534 155738
rect 79914 155418 79946 155654
rect 80182 155418 80266 155654
rect 80502 155418 80534 155654
rect 79914 118774 80534 155418
rect 79914 118538 79946 118774
rect 80182 118538 80266 118774
rect 80502 118538 80534 118774
rect 79914 118454 80534 118538
rect 79914 118218 79946 118454
rect 80182 118218 80266 118454
rect 80502 118218 80534 118454
rect 79914 81574 80534 118218
rect 79914 81338 79946 81574
rect 80182 81338 80266 81574
rect 80502 81338 80534 81574
rect 79914 81254 80534 81338
rect 79914 81018 79946 81254
rect 80182 81018 80266 81254
rect 80502 81018 80534 81254
rect 79914 44374 80534 81018
rect 79914 44138 79946 44374
rect 80182 44138 80266 44374
rect 80502 44138 80534 44374
rect 79914 44054 80534 44138
rect 79914 43818 79946 44054
rect 80182 43818 80266 44054
rect 80502 43818 80534 44054
rect 79914 7174 80534 43818
rect 79914 6938 79946 7174
rect 80182 6938 80266 7174
rect 80502 6938 80534 7174
rect 79914 6854 80534 6938
rect 79914 6618 79946 6854
rect 80182 6618 80266 6854
rect 80502 6618 80534 6854
rect 79914 2176 80534 6618
rect 83634 680494 84254 701760
rect 83634 680258 83666 680494
rect 83902 680258 83986 680494
rect 84222 680258 84254 680494
rect 83634 680174 84254 680258
rect 83634 679938 83666 680174
rect 83902 679938 83986 680174
rect 84222 679938 84254 680174
rect 83634 643294 84254 679938
rect 83634 643058 83666 643294
rect 83902 643058 83986 643294
rect 84222 643058 84254 643294
rect 83634 642974 84254 643058
rect 83634 642738 83666 642974
rect 83902 642738 83986 642974
rect 84222 642738 84254 642974
rect 83634 606094 84254 642738
rect 83634 605858 83666 606094
rect 83902 605858 83986 606094
rect 84222 605858 84254 606094
rect 83634 605774 84254 605858
rect 83634 605538 83666 605774
rect 83902 605538 83986 605774
rect 84222 605538 84254 605774
rect 83634 568894 84254 605538
rect 83634 568658 83666 568894
rect 83902 568658 83986 568894
rect 84222 568658 84254 568894
rect 83634 568574 84254 568658
rect 83634 568338 83666 568574
rect 83902 568338 83986 568574
rect 84222 568338 84254 568574
rect 83634 531694 84254 568338
rect 83634 531458 83666 531694
rect 83902 531458 83986 531694
rect 84222 531458 84254 531694
rect 83634 531374 84254 531458
rect 83634 531138 83666 531374
rect 83902 531138 83986 531374
rect 84222 531138 84254 531374
rect 83634 494494 84254 531138
rect 83634 494258 83666 494494
rect 83902 494258 83986 494494
rect 84222 494258 84254 494494
rect 83634 494174 84254 494258
rect 83634 493938 83666 494174
rect 83902 493938 83986 494174
rect 84222 493938 84254 494174
rect 83634 457294 84254 493938
rect 83634 457058 83666 457294
rect 83902 457058 83986 457294
rect 84222 457058 84254 457294
rect 83634 456974 84254 457058
rect 83634 456738 83666 456974
rect 83902 456738 83986 456974
rect 84222 456738 84254 456974
rect 83634 420094 84254 456738
rect 83634 419858 83666 420094
rect 83902 419858 83986 420094
rect 84222 419858 84254 420094
rect 83634 419774 84254 419858
rect 83634 419538 83666 419774
rect 83902 419538 83986 419774
rect 84222 419538 84254 419774
rect 83634 382894 84254 419538
rect 83634 382658 83666 382894
rect 83902 382658 83986 382894
rect 84222 382658 84254 382894
rect 83634 382574 84254 382658
rect 83634 382338 83666 382574
rect 83902 382338 83986 382574
rect 84222 382338 84254 382574
rect 83634 345694 84254 382338
rect 83634 345458 83666 345694
rect 83902 345458 83986 345694
rect 84222 345458 84254 345694
rect 83634 345374 84254 345458
rect 83634 345138 83666 345374
rect 83902 345138 83986 345374
rect 84222 345138 84254 345374
rect 83634 308494 84254 345138
rect 83634 308258 83666 308494
rect 83902 308258 83986 308494
rect 84222 308258 84254 308494
rect 83634 308174 84254 308258
rect 83634 307938 83666 308174
rect 83902 307938 83986 308174
rect 84222 307938 84254 308174
rect 83634 271294 84254 307938
rect 83634 271058 83666 271294
rect 83902 271058 83986 271294
rect 84222 271058 84254 271294
rect 83634 270974 84254 271058
rect 83634 270738 83666 270974
rect 83902 270738 83986 270974
rect 84222 270738 84254 270974
rect 83634 234094 84254 270738
rect 83634 233858 83666 234094
rect 83902 233858 83986 234094
rect 84222 233858 84254 234094
rect 83634 233774 84254 233858
rect 83634 233538 83666 233774
rect 83902 233538 83986 233774
rect 84222 233538 84254 233774
rect 83634 196894 84254 233538
rect 83634 196658 83666 196894
rect 83902 196658 83986 196894
rect 84222 196658 84254 196894
rect 83634 196574 84254 196658
rect 83634 196338 83666 196574
rect 83902 196338 83986 196574
rect 84222 196338 84254 196574
rect 83634 159694 84254 196338
rect 83634 159458 83666 159694
rect 83902 159458 83986 159694
rect 84222 159458 84254 159694
rect 83634 159374 84254 159458
rect 83634 159138 83666 159374
rect 83902 159138 83986 159374
rect 84222 159138 84254 159374
rect 83634 122494 84254 159138
rect 83634 122258 83666 122494
rect 83902 122258 83986 122494
rect 84222 122258 84254 122494
rect 83634 122174 84254 122258
rect 83634 121938 83666 122174
rect 83902 121938 83986 122174
rect 84222 121938 84254 122174
rect 83634 85294 84254 121938
rect 83634 85058 83666 85294
rect 83902 85058 83986 85294
rect 84222 85058 84254 85294
rect 83634 84974 84254 85058
rect 83634 84738 83666 84974
rect 83902 84738 83986 84974
rect 84222 84738 84254 84974
rect 83634 48094 84254 84738
rect 83634 47858 83666 48094
rect 83902 47858 83986 48094
rect 84222 47858 84254 48094
rect 83634 47774 84254 47858
rect 83634 47538 83666 47774
rect 83902 47538 83986 47774
rect 84222 47538 84254 47774
rect 83634 10894 84254 47538
rect 83634 10658 83666 10894
rect 83902 10658 83986 10894
rect 84222 10658 84254 10894
rect 83634 10574 84254 10658
rect 83634 10338 83666 10574
rect 83902 10338 83986 10574
rect 84222 10338 84254 10574
rect 83634 2176 84254 10338
rect 87354 684214 87974 701760
rect 87354 683978 87386 684214
rect 87622 683978 87706 684214
rect 87942 683978 87974 684214
rect 87354 683894 87974 683978
rect 87354 683658 87386 683894
rect 87622 683658 87706 683894
rect 87942 683658 87974 683894
rect 87354 647014 87974 683658
rect 87354 646778 87386 647014
rect 87622 646778 87706 647014
rect 87942 646778 87974 647014
rect 87354 646694 87974 646778
rect 87354 646458 87386 646694
rect 87622 646458 87706 646694
rect 87942 646458 87974 646694
rect 87354 609814 87974 646458
rect 87354 609578 87386 609814
rect 87622 609578 87706 609814
rect 87942 609578 87974 609814
rect 87354 609494 87974 609578
rect 87354 609258 87386 609494
rect 87622 609258 87706 609494
rect 87942 609258 87974 609494
rect 87354 572614 87974 609258
rect 87354 572378 87386 572614
rect 87622 572378 87706 572614
rect 87942 572378 87974 572614
rect 87354 572294 87974 572378
rect 87354 572058 87386 572294
rect 87622 572058 87706 572294
rect 87942 572058 87974 572294
rect 87354 535414 87974 572058
rect 87354 535178 87386 535414
rect 87622 535178 87706 535414
rect 87942 535178 87974 535414
rect 87354 535094 87974 535178
rect 87354 534858 87386 535094
rect 87622 534858 87706 535094
rect 87942 534858 87974 535094
rect 87354 498214 87974 534858
rect 87354 497978 87386 498214
rect 87622 497978 87706 498214
rect 87942 497978 87974 498214
rect 87354 497894 87974 497978
rect 87354 497658 87386 497894
rect 87622 497658 87706 497894
rect 87942 497658 87974 497894
rect 87354 461014 87974 497658
rect 87354 460778 87386 461014
rect 87622 460778 87706 461014
rect 87942 460778 87974 461014
rect 87354 460694 87974 460778
rect 87354 460458 87386 460694
rect 87622 460458 87706 460694
rect 87942 460458 87974 460694
rect 87354 423814 87974 460458
rect 87354 423578 87386 423814
rect 87622 423578 87706 423814
rect 87942 423578 87974 423814
rect 87354 423494 87974 423578
rect 87354 423258 87386 423494
rect 87622 423258 87706 423494
rect 87942 423258 87974 423494
rect 87354 386614 87974 423258
rect 87354 386378 87386 386614
rect 87622 386378 87706 386614
rect 87942 386378 87974 386614
rect 87354 386294 87974 386378
rect 87354 386058 87386 386294
rect 87622 386058 87706 386294
rect 87942 386058 87974 386294
rect 87354 349414 87974 386058
rect 87354 349178 87386 349414
rect 87622 349178 87706 349414
rect 87942 349178 87974 349414
rect 87354 349094 87974 349178
rect 87354 348858 87386 349094
rect 87622 348858 87706 349094
rect 87942 348858 87974 349094
rect 87354 312214 87974 348858
rect 87354 311978 87386 312214
rect 87622 311978 87706 312214
rect 87942 311978 87974 312214
rect 87354 311894 87974 311978
rect 87354 311658 87386 311894
rect 87622 311658 87706 311894
rect 87942 311658 87974 311894
rect 87354 275014 87974 311658
rect 87354 274778 87386 275014
rect 87622 274778 87706 275014
rect 87942 274778 87974 275014
rect 87354 274694 87974 274778
rect 87354 274458 87386 274694
rect 87622 274458 87706 274694
rect 87942 274458 87974 274694
rect 87354 237814 87974 274458
rect 87354 237578 87386 237814
rect 87622 237578 87706 237814
rect 87942 237578 87974 237814
rect 87354 237494 87974 237578
rect 87354 237258 87386 237494
rect 87622 237258 87706 237494
rect 87942 237258 87974 237494
rect 87354 200614 87974 237258
rect 87354 200378 87386 200614
rect 87622 200378 87706 200614
rect 87942 200378 87974 200614
rect 87354 200294 87974 200378
rect 87354 200058 87386 200294
rect 87622 200058 87706 200294
rect 87942 200058 87974 200294
rect 87354 163414 87974 200058
rect 87354 163178 87386 163414
rect 87622 163178 87706 163414
rect 87942 163178 87974 163414
rect 87354 163094 87974 163178
rect 87354 162858 87386 163094
rect 87622 162858 87706 163094
rect 87942 162858 87974 163094
rect 87354 126214 87974 162858
rect 87354 125978 87386 126214
rect 87622 125978 87706 126214
rect 87942 125978 87974 126214
rect 87354 125894 87974 125978
rect 87354 125658 87386 125894
rect 87622 125658 87706 125894
rect 87942 125658 87974 125894
rect 87354 89014 87974 125658
rect 87354 88778 87386 89014
rect 87622 88778 87706 89014
rect 87942 88778 87974 89014
rect 87354 88694 87974 88778
rect 87354 88458 87386 88694
rect 87622 88458 87706 88694
rect 87942 88458 87974 88694
rect 87354 51814 87974 88458
rect 87354 51578 87386 51814
rect 87622 51578 87706 51814
rect 87942 51578 87974 51814
rect 87354 51494 87974 51578
rect 87354 51258 87386 51494
rect 87622 51258 87706 51494
rect 87942 51258 87974 51494
rect 87354 14614 87974 51258
rect 87354 14378 87386 14614
rect 87622 14378 87706 14614
rect 87942 14378 87974 14614
rect 87354 14294 87974 14378
rect 87354 14058 87386 14294
rect 87622 14058 87706 14294
rect 87942 14058 87974 14294
rect 87354 2176 87974 14058
rect 91074 687934 91694 701760
rect 91074 687698 91106 687934
rect 91342 687698 91426 687934
rect 91662 687698 91694 687934
rect 91074 687614 91694 687698
rect 91074 687378 91106 687614
rect 91342 687378 91426 687614
rect 91662 687378 91694 687614
rect 91074 650734 91694 687378
rect 91074 650498 91106 650734
rect 91342 650498 91426 650734
rect 91662 650498 91694 650734
rect 91074 650414 91694 650498
rect 91074 650178 91106 650414
rect 91342 650178 91426 650414
rect 91662 650178 91694 650414
rect 91074 613534 91694 650178
rect 91074 613298 91106 613534
rect 91342 613298 91426 613534
rect 91662 613298 91694 613534
rect 91074 613214 91694 613298
rect 91074 612978 91106 613214
rect 91342 612978 91426 613214
rect 91662 612978 91694 613214
rect 91074 576334 91694 612978
rect 91074 576098 91106 576334
rect 91342 576098 91426 576334
rect 91662 576098 91694 576334
rect 91074 576014 91694 576098
rect 91074 575778 91106 576014
rect 91342 575778 91426 576014
rect 91662 575778 91694 576014
rect 91074 539134 91694 575778
rect 91074 538898 91106 539134
rect 91342 538898 91426 539134
rect 91662 538898 91694 539134
rect 91074 538814 91694 538898
rect 91074 538578 91106 538814
rect 91342 538578 91426 538814
rect 91662 538578 91694 538814
rect 91074 501934 91694 538578
rect 91074 501698 91106 501934
rect 91342 501698 91426 501934
rect 91662 501698 91694 501934
rect 91074 501614 91694 501698
rect 91074 501378 91106 501614
rect 91342 501378 91426 501614
rect 91662 501378 91694 501614
rect 91074 464734 91694 501378
rect 91074 464498 91106 464734
rect 91342 464498 91426 464734
rect 91662 464498 91694 464734
rect 91074 464414 91694 464498
rect 91074 464178 91106 464414
rect 91342 464178 91426 464414
rect 91662 464178 91694 464414
rect 91074 427534 91694 464178
rect 91074 427298 91106 427534
rect 91342 427298 91426 427534
rect 91662 427298 91694 427534
rect 91074 427214 91694 427298
rect 91074 426978 91106 427214
rect 91342 426978 91426 427214
rect 91662 426978 91694 427214
rect 91074 390334 91694 426978
rect 91074 390098 91106 390334
rect 91342 390098 91426 390334
rect 91662 390098 91694 390334
rect 91074 390014 91694 390098
rect 91074 389778 91106 390014
rect 91342 389778 91426 390014
rect 91662 389778 91694 390014
rect 91074 353134 91694 389778
rect 91074 352898 91106 353134
rect 91342 352898 91426 353134
rect 91662 352898 91694 353134
rect 91074 352814 91694 352898
rect 91074 352578 91106 352814
rect 91342 352578 91426 352814
rect 91662 352578 91694 352814
rect 91074 315934 91694 352578
rect 91074 315698 91106 315934
rect 91342 315698 91426 315934
rect 91662 315698 91694 315934
rect 91074 315614 91694 315698
rect 91074 315378 91106 315614
rect 91342 315378 91426 315614
rect 91662 315378 91694 315614
rect 91074 278734 91694 315378
rect 91074 278498 91106 278734
rect 91342 278498 91426 278734
rect 91662 278498 91694 278734
rect 91074 278414 91694 278498
rect 91074 278178 91106 278414
rect 91342 278178 91426 278414
rect 91662 278178 91694 278414
rect 91074 241534 91694 278178
rect 91074 241298 91106 241534
rect 91342 241298 91426 241534
rect 91662 241298 91694 241534
rect 91074 241214 91694 241298
rect 91074 240978 91106 241214
rect 91342 240978 91426 241214
rect 91662 240978 91694 241214
rect 91074 204334 91694 240978
rect 91074 204098 91106 204334
rect 91342 204098 91426 204334
rect 91662 204098 91694 204334
rect 91074 204014 91694 204098
rect 91074 203778 91106 204014
rect 91342 203778 91426 204014
rect 91662 203778 91694 204014
rect 91074 167134 91694 203778
rect 91074 166898 91106 167134
rect 91342 166898 91426 167134
rect 91662 166898 91694 167134
rect 91074 166814 91694 166898
rect 91074 166578 91106 166814
rect 91342 166578 91426 166814
rect 91662 166578 91694 166814
rect 91074 129934 91694 166578
rect 91074 129698 91106 129934
rect 91342 129698 91426 129934
rect 91662 129698 91694 129934
rect 91074 129614 91694 129698
rect 91074 129378 91106 129614
rect 91342 129378 91426 129614
rect 91662 129378 91694 129614
rect 91074 92734 91694 129378
rect 91074 92498 91106 92734
rect 91342 92498 91426 92734
rect 91662 92498 91694 92734
rect 91074 92414 91694 92498
rect 91074 92178 91106 92414
rect 91342 92178 91426 92414
rect 91662 92178 91694 92414
rect 91074 55534 91694 92178
rect 91074 55298 91106 55534
rect 91342 55298 91426 55534
rect 91662 55298 91694 55534
rect 91074 55214 91694 55298
rect 91074 54978 91106 55214
rect 91342 54978 91426 55214
rect 91662 54978 91694 55214
rect 91074 18334 91694 54978
rect 91074 18098 91106 18334
rect 91342 18098 91426 18334
rect 91662 18098 91694 18334
rect 91074 18014 91694 18098
rect 91074 17778 91106 18014
rect 91342 17778 91426 18014
rect 91662 17778 91694 18014
rect 91074 2176 91694 17778
rect 94794 691654 95414 701760
rect 94794 691418 94826 691654
rect 95062 691418 95146 691654
rect 95382 691418 95414 691654
rect 94794 691334 95414 691418
rect 94794 691098 94826 691334
rect 95062 691098 95146 691334
rect 95382 691098 95414 691334
rect 94794 654454 95414 691098
rect 94794 654218 94826 654454
rect 95062 654218 95146 654454
rect 95382 654218 95414 654454
rect 94794 654134 95414 654218
rect 94794 653898 94826 654134
rect 95062 653898 95146 654134
rect 95382 653898 95414 654134
rect 94794 617254 95414 653898
rect 94794 617018 94826 617254
rect 95062 617018 95146 617254
rect 95382 617018 95414 617254
rect 94794 616934 95414 617018
rect 94794 616698 94826 616934
rect 95062 616698 95146 616934
rect 95382 616698 95414 616934
rect 94794 580054 95414 616698
rect 94794 579818 94826 580054
rect 95062 579818 95146 580054
rect 95382 579818 95414 580054
rect 94794 579734 95414 579818
rect 94794 579498 94826 579734
rect 95062 579498 95146 579734
rect 95382 579498 95414 579734
rect 94794 542854 95414 579498
rect 94794 542618 94826 542854
rect 95062 542618 95146 542854
rect 95382 542618 95414 542854
rect 94794 542534 95414 542618
rect 94794 542298 94826 542534
rect 95062 542298 95146 542534
rect 95382 542298 95414 542534
rect 94794 505654 95414 542298
rect 94794 505418 94826 505654
rect 95062 505418 95146 505654
rect 95382 505418 95414 505654
rect 94794 505334 95414 505418
rect 94794 505098 94826 505334
rect 95062 505098 95146 505334
rect 95382 505098 95414 505334
rect 94794 468454 95414 505098
rect 94794 468218 94826 468454
rect 95062 468218 95146 468454
rect 95382 468218 95414 468454
rect 94794 468134 95414 468218
rect 94794 467898 94826 468134
rect 95062 467898 95146 468134
rect 95382 467898 95414 468134
rect 94794 431254 95414 467898
rect 94794 431018 94826 431254
rect 95062 431018 95146 431254
rect 95382 431018 95414 431254
rect 94794 430934 95414 431018
rect 94794 430698 94826 430934
rect 95062 430698 95146 430934
rect 95382 430698 95414 430934
rect 94794 394054 95414 430698
rect 94794 393818 94826 394054
rect 95062 393818 95146 394054
rect 95382 393818 95414 394054
rect 94794 393734 95414 393818
rect 94794 393498 94826 393734
rect 95062 393498 95146 393734
rect 95382 393498 95414 393734
rect 94794 356854 95414 393498
rect 94794 356618 94826 356854
rect 95062 356618 95146 356854
rect 95382 356618 95414 356854
rect 94794 356534 95414 356618
rect 94794 356298 94826 356534
rect 95062 356298 95146 356534
rect 95382 356298 95414 356534
rect 94794 319654 95414 356298
rect 94794 319418 94826 319654
rect 95062 319418 95146 319654
rect 95382 319418 95414 319654
rect 94794 319334 95414 319418
rect 94794 319098 94826 319334
rect 95062 319098 95146 319334
rect 95382 319098 95414 319334
rect 94794 282454 95414 319098
rect 94794 282218 94826 282454
rect 95062 282218 95146 282454
rect 95382 282218 95414 282454
rect 94794 282134 95414 282218
rect 94794 281898 94826 282134
rect 95062 281898 95146 282134
rect 95382 281898 95414 282134
rect 94794 245254 95414 281898
rect 94794 245018 94826 245254
rect 95062 245018 95146 245254
rect 95382 245018 95414 245254
rect 94794 244934 95414 245018
rect 94794 244698 94826 244934
rect 95062 244698 95146 244934
rect 95382 244698 95414 244934
rect 94794 208054 95414 244698
rect 94794 207818 94826 208054
rect 95062 207818 95146 208054
rect 95382 207818 95414 208054
rect 94794 207734 95414 207818
rect 94794 207498 94826 207734
rect 95062 207498 95146 207734
rect 95382 207498 95414 207734
rect 94794 170854 95414 207498
rect 94794 170618 94826 170854
rect 95062 170618 95146 170854
rect 95382 170618 95414 170854
rect 94794 170534 95414 170618
rect 94794 170298 94826 170534
rect 95062 170298 95146 170534
rect 95382 170298 95414 170534
rect 94794 133654 95414 170298
rect 94794 133418 94826 133654
rect 95062 133418 95146 133654
rect 95382 133418 95414 133654
rect 94794 133334 95414 133418
rect 94794 133098 94826 133334
rect 95062 133098 95146 133334
rect 95382 133098 95414 133334
rect 94794 96454 95414 133098
rect 94794 96218 94826 96454
rect 95062 96218 95146 96454
rect 95382 96218 95414 96454
rect 94794 96134 95414 96218
rect 94794 95898 94826 96134
rect 95062 95898 95146 96134
rect 95382 95898 95414 96134
rect 94794 59254 95414 95898
rect 94794 59018 94826 59254
rect 95062 59018 95146 59254
rect 95382 59018 95414 59254
rect 94794 58934 95414 59018
rect 94794 58698 94826 58934
rect 95062 58698 95146 58934
rect 95382 58698 95414 58934
rect 94794 22054 95414 58698
rect 94794 21818 94826 22054
rect 95062 21818 95146 22054
rect 95382 21818 95414 22054
rect 94794 21734 95414 21818
rect 94794 21498 94826 21734
rect 95062 21498 95146 21734
rect 95382 21498 95414 21734
rect 94794 2176 95414 21498
rect 98514 695374 99134 701760
rect 98514 695138 98546 695374
rect 98782 695138 98866 695374
rect 99102 695138 99134 695374
rect 98514 695054 99134 695138
rect 98514 694818 98546 695054
rect 98782 694818 98866 695054
rect 99102 694818 99134 695054
rect 98514 658174 99134 694818
rect 98514 657938 98546 658174
rect 98782 657938 98866 658174
rect 99102 657938 99134 658174
rect 98514 657854 99134 657938
rect 98514 657618 98546 657854
rect 98782 657618 98866 657854
rect 99102 657618 99134 657854
rect 98514 620974 99134 657618
rect 98514 620738 98546 620974
rect 98782 620738 98866 620974
rect 99102 620738 99134 620974
rect 98514 620654 99134 620738
rect 98514 620418 98546 620654
rect 98782 620418 98866 620654
rect 99102 620418 99134 620654
rect 98514 583774 99134 620418
rect 98514 583538 98546 583774
rect 98782 583538 98866 583774
rect 99102 583538 99134 583774
rect 98514 583454 99134 583538
rect 98514 583218 98546 583454
rect 98782 583218 98866 583454
rect 99102 583218 99134 583454
rect 98514 546574 99134 583218
rect 98514 546338 98546 546574
rect 98782 546338 98866 546574
rect 99102 546338 99134 546574
rect 98514 546254 99134 546338
rect 98514 546018 98546 546254
rect 98782 546018 98866 546254
rect 99102 546018 99134 546254
rect 98514 509374 99134 546018
rect 98514 509138 98546 509374
rect 98782 509138 98866 509374
rect 99102 509138 99134 509374
rect 98514 509054 99134 509138
rect 98514 508818 98546 509054
rect 98782 508818 98866 509054
rect 99102 508818 99134 509054
rect 98514 472174 99134 508818
rect 98514 471938 98546 472174
rect 98782 471938 98866 472174
rect 99102 471938 99134 472174
rect 98514 471854 99134 471938
rect 98514 471618 98546 471854
rect 98782 471618 98866 471854
rect 99102 471618 99134 471854
rect 98514 434974 99134 471618
rect 98514 434738 98546 434974
rect 98782 434738 98866 434974
rect 99102 434738 99134 434974
rect 98514 434654 99134 434738
rect 98514 434418 98546 434654
rect 98782 434418 98866 434654
rect 99102 434418 99134 434654
rect 98514 397774 99134 434418
rect 98514 397538 98546 397774
rect 98782 397538 98866 397774
rect 99102 397538 99134 397774
rect 98514 397454 99134 397538
rect 98514 397218 98546 397454
rect 98782 397218 98866 397454
rect 99102 397218 99134 397454
rect 98514 360574 99134 397218
rect 98514 360338 98546 360574
rect 98782 360338 98866 360574
rect 99102 360338 99134 360574
rect 98514 360254 99134 360338
rect 98514 360018 98546 360254
rect 98782 360018 98866 360254
rect 99102 360018 99134 360254
rect 98514 323374 99134 360018
rect 98514 323138 98546 323374
rect 98782 323138 98866 323374
rect 99102 323138 99134 323374
rect 98514 323054 99134 323138
rect 98514 322818 98546 323054
rect 98782 322818 98866 323054
rect 99102 322818 99134 323054
rect 98514 286174 99134 322818
rect 98514 285938 98546 286174
rect 98782 285938 98866 286174
rect 99102 285938 99134 286174
rect 98514 285854 99134 285938
rect 98514 285618 98546 285854
rect 98782 285618 98866 285854
rect 99102 285618 99134 285854
rect 98514 248974 99134 285618
rect 98514 248738 98546 248974
rect 98782 248738 98866 248974
rect 99102 248738 99134 248974
rect 98514 248654 99134 248738
rect 98514 248418 98546 248654
rect 98782 248418 98866 248654
rect 99102 248418 99134 248654
rect 98514 211774 99134 248418
rect 98514 211538 98546 211774
rect 98782 211538 98866 211774
rect 99102 211538 99134 211774
rect 98514 211454 99134 211538
rect 98514 211218 98546 211454
rect 98782 211218 98866 211454
rect 99102 211218 99134 211454
rect 98514 174574 99134 211218
rect 98514 174338 98546 174574
rect 98782 174338 98866 174574
rect 99102 174338 99134 174574
rect 98514 174254 99134 174338
rect 98514 174018 98546 174254
rect 98782 174018 98866 174254
rect 99102 174018 99134 174254
rect 98514 137374 99134 174018
rect 98514 137138 98546 137374
rect 98782 137138 98866 137374
rect 99102 137138 99134 137374
rect 98514 137054 99134 137138
rect 98514 136818 98546 137054
rect 98782 136818 98866 137054
rect 99102 136818 99134 137054
rect 98514 100174 99134 136818
rect 98514 99938 98546 100174
rect 98782 99938 98866 100174
rect 99102 99938 99134 100174
rect 98514 99854 99134 99938
rect 98514 99618 98546 99854
rect 98782 99618 98866 99854
rect 99102 99618 99134 99854
rect 98514 62974 99134 99618
rect 98514 62738 98546 62974
rect 98782 62738 98866 62974
rect 99102 62738 99134 62974
rect 98514 62654 99134 62738
rect 98514 62418 98546 62654
rect 98782 62418 98866 62654
rect 99102 62418 99134 62654
rect 98514 25774 99134 62418
rect 98514 25538 98546 25774
rect 98782 25538 98866 25774
rect 99102 25538 99134 25774
rect 98514 25454 99134 25538
rect 98514 25218 98546 25454
rect 98782 25218 98866 25454
rect 99102 25218 99134 25454
rect 98514 2176 99134 25218
rect 102234 699094 102854 701760
rect 102234 698858 102266 699094
rect 102502 698858 102586 699094
rect 102822 698858 102854 699094
rect 102234 698774 102854 698858
rect 102234 698538 102266 698774
rect 102502 698538 102586 698774
rect 102822 698538 102854 698774
rect 102234 661894 102854 698538
rect 102234 661658 102266 661894
rect 102502 661658 102586 661894
rect 102822 661658 102854 661894
rect 102234 661574 102854 661658
rect 102234 661338 102266 661574
rect 102502 661338 102586 661574
rect 102822 661338 102854 661574
rect 102234 624694 102854 661338
rect 102234 624458 102266 624694
rect 102502 624458 102586 624694
rect 102822 624458 102854 624694
rect 102234 624374 102854 624458
rect 102234 624138 102266 624374
rect 102502 624138 102586 624374
rect 102822 624138 102854 624374
rect 102234 587494 102854 624138
rect 102234 587258 102266 587494
rect 102502 587258 102586 587494
rect 102822 587258 102854 587494
rect 102234 587174 102854 587258
rect 102234 586938 102266 587174
rect 102502 586938 102586 587174
rect 102822 586938 102854 587174
rect 102234 550294 102854 586938
rect 102234 550058 102266 550294
rect 102502 550058 102586 550294
rect 102822 550058 102854 550294
rect 102234 549974 102854 550058
rect 102234 549738 102266 549974
rect 102502 549738 102586 549974
rect 102822 549738 102854 549974
rect 102234 513094 102854 549738
rect 102234 512858 102266 513094
rect 102502 512858 102586 513094
rect 102822 512858 102854 513094
rect 102234 512774 102854 512858
rect 102234 512538 102266 512774
rect 102502 512538 102586 512774
rect 102822 512538 102854 512774
rect 102234 475894 102854 512538
rect 102234 475658 102266 475894
rect 102502 475658 102586 475894
rect 102822 475658 102854 475894
rect 102234 475574 102854 475658
rect 102234 475338 102266 475574
rect 102502 475338 102586 475574
rect 102822 475338 102854 475574
rect 102234 438694 102854 475338
rect 102234 438458 102266 438694
rect 102502 438458 102586 438694
rect 102822 438458 102854 438694
rect 102234 438374 102854 438458
rect 102234 438138 102266 438374
rect 102502 438138 102586 438374
rect 102822 438138 102854 438374
rect 102234 401494 102854 438138
rect 102234 401258 102266 401494
rect 102502 401258 102586 401494
rect 102822 401258 102854 401494
rect 102234 401174 102854 401258
rect 102234 400938 102266 401174
rect 102502 400938 102586 401174
rect 102822 400938 102854 401174
rect 102234 364294 102854 400938
rect 102234 364058 102266 364294
rect 102502 364058 102586 364294
rect 102822 364058 102854 364294
rect 102234 363974 102854 364058
rect 102234 363738 102266 363974
rect 102502 363738 102586 363974
rect 102822 363738 102854 363974
rect 102234 327094 102854 363738
rect 102234 326858 102266 327094
rect 102502 326858 102586 327094
rect 102822 326858 102854 327094
rect 102234 326774 102854 326858
rect 102234 326538 102266 326774
rect 102502 326538 102586 326774
rect 102822 326538 102854 326774
rect 102234 289894 102854 326538
rect 102234 289658 102266 289894
rect 102502 289658 102586 289894
rect 102822 289658 102854 289894
rect 102234 289574 102854 289658
rect 102234 289338 102266 289574
rect 102502 289338 102586 289574
rect 102822 289338 102854 289574
rect 102234 252694 102854 289338
rect 102234 252458 102266 252694
rect 102502 252458 102586 252694
rect 102822 252458 102854 252694
rect 102234 252374 102854 252458
rect 102234 252138 102266 252374
rect 102502 252138 102586 252374
rect 102822 252138 102854 252374
rect 102234 215494 102854 252138
rect 102234 215258 102266 215494
rect 102502 215258 102586 215494
rect 102822 215258 102854 215494
rect 102234 215174 102854 215258
rect 102234 214938 102266 215174
rect 102502 214938 102586 215174
rect 102822 214938 102854 215174
rect 102234 178294 102854 214938
rect 102234 178058 102266 178294
rect 102502 178058 102586 178294
rect 102822 178058 102854 178294
rect 102234 177974 102854 178058
rect 102234 177738 102266 177974
rect 102502 177738 102586 177974
rect 102822 177738 102854 177974
rect 102234 141094 102854 177738
rect 102234 140858 102266 141094
rect 102502 140858 102586 141094
rect 102822 140858 102854 141094
rect 102234 140774 102854 140858
rect 102234 140538 102266 140774
rect 102502 140538 102586 140774
rect 102822 140538 102854 140774
rect 102234 103894 102854 140538
rect 102234 103658 102266 103894
rect 102502 103658 102586 103894
rect 102822 103658 102854 103894
rect 102234 103574 102854 103658
rect 102234 103338 102266 103574
rect 102502 103338 102586 103574
rect 102822 103338 102854 103574
rect 102234 66694 102854 103338
rect 102234 66458 102266 66694
rect 102502 66458 102586 66694
rect 102822 66458 102854 66694
rect 102234 66374 102854 66458
rect 102234 66138 102266 66374
rect 102502 66138 102586 66374
rect 102822 66138 102854 66374
rect 102234 29494 102854 66138
rect 102234 29258 102266 29494
rect 102502 29258 102586 29494
rect 102822 29258 102854 29494
rect 102234 29174 102854 29258
rect 102234 28938 102266 29174
rect 102502 28938 102586 29174
rect 102822 28938 102854 29174
rect 102234 2176 102854 28938
rect 113394 673054 114014 701760
rect 113394 672818 113426 673054
rect 113662 672818 113746 673054
rect 113982 672818 114014 673054
rect 113394 672734 114014 672818
rect 113394 672498 113426 672734
rect 113662 672498 113746 672734
rect 113982 672498 114014 672734
rect 113394 635854 114014 672498
rect 113394 635618 113426 635854
rect 113662 635618 113746 635854
rect 113982 635618 114014 635854
rect 113394 635534 114014 635618
rect 113394 635298 113426 635534
rect 113662 635298 113746 635534
rect 113982 635298 114014 635534
rect 113394 598654 114014 635298
rect 113394 598418 113426 598654
rect 113662 598418 113746 598654
rect 113982 598418 114014 598654
rect 113394 598334 114014 598418
rect 113394 598098 113426 598334
rect 113662 598098 113746 598334
rect 113982 598098 114014 598334
rect 113394 561454 114014 598098
rect 113394 561218 113426 561454
rect 113662 561218 113746 561454
rect 113982 561218 114014 561454
rect 113394 561134 114014 561218
rect 113394 560898 113426 561134
rect 113662 560898 113746 561134
rect 113982 560898 114014 561134
rect 113394 524254 114014 560898
rect 113394 524018 113426 524254
rect 113662 524018 113746 524254
rect 113982 524018 114014 524254
rect 113394 523934 114014 524018
rect 113394 523698 113426 523934
rect 113662 523698 113746 523934
rect 113982 523698 114014 523934
rect 113394 487054 114014 523698
rect 113394 486818 113426 487054
rect 113662 486818 113746 487054
rect 113982 486818 114014 487054
rect 113394 486734 114014 486818
rect 113394 486498 113426 486734
rect 113662 486498 113746 486734
rect 113982 486498 114014 486734
rect 113394 449854 114014 486498
rect 113394 449618 113426 449854
rect 113662 449618 113746 449854
rect 113982 449618 114014 449854
rect 113394 449534 114014 449618
rect 113394 449298 113426 449534
rect 113662 449298 113746 449534
rect 113982 449298 114014 449534
rect 113394 412654 114014 449298
rect 113394 412418 113426 412654
rect 113662 412418 113746 412654
rect 113982 412418 114014 412654
rect 113394 412334 114014 412418
rect 113394 412098 113426 412334
rect 113662 412098 113746 412334
rect 113982 412098 114014 412334
rect 113394 375454 114014 412098
rect 113394 375218 113426 375454
rect 113662 375218 113746 375454
rect 113982 375218 114014 375454
rect 113394 375134 114014 375218
rect 113394 374898 113426 375134
rect 113662 374898 113746 375134
rect 113982 374898 114014 375134
rect 113394 338254 114014 374898
rect 113394 338018 113426 338254
rect 113662 338018 113746 338254
rect 113982 338018 114014 338254
rect 113394 337934 114014 338018
rect 113394 337698 113426 337934
rect 113662 337698 113746 337934
rect 113982 337698 114014 337934
rect 113394 301054 114014 337698
rect 113394 300818 113426 301054
rect 113662 300818 113746 301054
rect 113982 300818 114014 301054
rect 113394 300734 114014 300818
rect 113394 300498 113426 300734
rect 113662 300498 113746 300734
rect 113982 300498 114014 300734
rect 113394 263854 114014 300498
rect 113394 263618 113426 263854
rect 113662 263618 113746 263854
rect 113982 263618 114014 263854
rect 113394 263534 114014 263618
rect 113394 263298 113426 263534
rect 113662 263298 113746 263534
rect 113982 263298 114014 263534
rect 113394 226654 114014 263298
rect 113394 226418 113426 226654
rect 113662 226418 113746 226654
rect 113982 226418 114014 226654
rect 113394 226334 114014 226418
rect 113394 226098 113426 226334
rect 113662 226098 113746 226334
rect 113982 226098 114014 226334
rect 113394 189454 114014 226098
rect 113394 189218 113426 189454
rect 113662 189218 113746 189454
rect 113982 189218 114014 189454
rect 113394 189134 114014 189218
rect 113394 188898 113426 189134
rect 113662 188898 113746 189134
rect 113982 188898 114014 189134
rect 113394 152254 114014 188898
rect 113394 152018 113426 152254
rect 113662 152018 113746 152254
rect 113982 152018 114014 152254
rect 113394 151934 114014 152018
rect 113394 151698 113426 151934
rect 113662 151698 113746 151934
rect 113982 151698 114014 151934
rect 113394 115054 114014 151698
rect 113394 114818 113426 115054
rect 113662 114818 113746 115054
rect 113982 114818 114014 115054
rect 113394 114734 114014 114818
rect 113394 114498 113426 114734
rect 113662 114498 113746 114734
rect 113982 114498 114014 114734
rect 113394 77854 114014 114498
rect 113394 77618 113426 77854
rect 113662 77618 113746 77854
rect 113982 77618 114014 77854
rect 113394 77534 114014 77618
rect 113394 77298 113426 77534
rect 113662 77298 113746 77534
rect 113982 77298 114014 77534
rect 113394 40654 114014 77298
rect 113394 40418 113426 40654
rect 113662 40418 113746 40654
rect 113982 40418 114014 40654
rect 113394 40334 114014 40418
rect 113394 40098 113426 40334
rect 113662 40098 113746 40334
rect 113982 40098 114014 40334
rect 113394 3454 114014 40098
rect 113394 3218 113426 3454
rect 113662 3218 113746 3454
rect 113982 3218 114014 3454
rect 113394 3134 114014 3218
rect 113394 2898 113426 3134
rect 113662 2898 113746 3134
rect 113982 2898 114014 3134
rect 113394 2176 114014 2898
rect 117114 676774 117734 701760
rect 117114 676538 117146 676774
rect 117382 676538 117466 676774
rect 117702 676538 117734 676774
rect 117114 676454 117734 676538
rect 117114 676218 117146 676454
rect 117382 676218 117466 676454
rect 117702 676218 117734 676454
rect 117114 639574 117734 676218
rect 117114 639338 117146 639574
rect 117382 639338 117466 639574
rect 117702 639338 117734 639574
rect 117114 639254 117734 639338
rect 117114 639018 117146 639254
rect 117382 639018 117466 639254
rect 117702 639018 117734 639254
rect 117114 602374 117734 639018
rect 117114 602138 117146 602374
rect 117382 602138 117466 602374
rect 117702 602138 117734 602374
rect 117114 602054 117734 602138
rect 117114 601818 117146 602054
rect 117382 601818 117466 602054
rect 117702 601818 117734 602054
rect 117114 565174 117734 601818
rect 117114 564938 117146 565174
rect 117382 564938 117466 565174
rect 117702 564938 117734 565174
rect 117114 564854 117734 564938
rect 117114 564618 117146 564854
rect 117382 564618 117466 564854
rect 117702 564618 117734 564854
rect 117114 527974 117734 564618
rect 117114 527738 117146 527974
rect 117382 527738 117466 527974
rect 117702 527738 117734 527974
rect 117114 527654 117734 527738
rect 117114 527418 117146 527654
rect 117382 527418 117466 527654
rect 117702 527418 117734 527654
rect 117114 490774 117734 527418
rect 117114 490538 117146 490774
rect 117382 490538 117466 490774
rect 117702 490538 117734 490774
rect 117114 490454 117734 490538
rect 117114 490218 117146 490454
rect 117382 490218 117466 490454
rect 117702 490218 117734 490454
rect 117114 453574 117734 490218
rect 117114 453338 117146 453574
rect 117382 453338 117466 453574
rect 117702 453338 117734 453574
rect 117114 453254 117734 453338
rect 117114 453018 117146 453254
rect 117382 453018 117466 453254
rect 117702 453018 117734 453254
rect 117114 416374 117734 453018
rect 117114 416138 117146 416374
rect 117382 416138 117466 416374
rect 117702 416138 117734 416374
rect 117114 416054 117734 416138
rect 117114 415818 117146 416054
rect 117382 415818 117466 416054
rect 117702 415818 117734 416054
rect 117114 379174 117734 415818
rect 117114 378938 117146 379174
rect 117382 378938 117466 379174
rect 117702 378938 117734 379174
rect 117114 378854 117734 378938
rect 117114 378618 117146 378854
rect 117382 378618 117466 378854
rect 117702 378618 117734 378854
rect 117114 341974 117734 378618
rect 117114 341738 117146 341974
rect 117382 341738 117466 341974
rect 117702 341738 117734 341974
rect 117114 341654 117734 341738
rect 117114 341418 117146 341654
rect 117382 341418 117466 341654
rect 117702 341418 117734 341654
rect 117114 304774 117734 341418
rect 117114 304538 117146 304774
rect 117382 304538 117466 304774
rect 117702 304538 117734 304774
rect 117114 304454 117734 304538
rect 117114 304218 117146 304454
rect 117382 304218 117466 304454
rect 117702 304218 117734 304454
rect 117114 267574 117734 304218
rect 117114 267338 117146 267574
rect 117382 267338 117466 267574
rect 117702 267338 117734 267574
rect 117114 267254 117734 267338
rect 117114 267018 117146 267254
rect 117382 267018 117466 267254
rect 117702 267018 117734 267254
rect 117114 230374 117734 267018
rect 117114 230138 117146 230374
rect 117382 230138 117466 230374
rect 117702 230138 117734 230374
rect 117114 230054 117734 230138
rect 117114 229818 117146 230054
rect 117382 229818 117466 230054
rect 117702 229818 117734 230054
rect 117114 193174 117734 229818
rect 117114 192938 117146 193174
rect 117382 192938 117466 193174
rect 117702 192938 117734 193174
rect 117114 192854 117734 192938
rect 117114 192618 117146 192854
rect 117382 192618 117466 192854
rect 117702 192618 117734 192854
rect 117114 155974 117734 192618
rect 117114 155738 117146 155974
rect 117382 155738 117466 155974
rect 117702 155738 117734 155974
rect 117114 155654 117734 155738
rect 117114 155418 117146 155654
rect 117382 155418 117466 155654
rect 117702 155418 117734 155654
rect 117114 118774 117734 155418
rect 117114 118538 117146 118774
rect 117382 118538 117466 118774
rect 117702 118538 117734 118774
rect 117114 118454 117734 118538
rect 117114 118218 117146 118454
rect 117382 118218 117466 118454
rect 117702 118218 117734 118454
rect 117114 81574 117734 118218
rect 117114 81338 117146 81574
rect 117382 81338 117466 81574
rect 117702 81338 117734 81574
rect 117114 81254 117734 81338
rect 117114 81018 117146 81254
rect 117382 81018 117466 81254
rect 117702 81018 117734 81254
rect 117114 44374 117734 81018
rect 117114 44138 117146 44374
rect 117382 44138 117466 44374
rect 117702 44138 117734 44374
rect 117114 44054 117734 44138
rect 117114 43818 117146 44054
rect 117382 43818 117466 44054
rect 117702 43818 117734 44054
rect 117114 7174 117734 43818
rect 117114 6938 117146 7174
rect 117382 6938 117466 7174
rect 117702 6938 117734 7174
rect 117114 6854 117734 6938
rect 117114 6618 117146 6854
rect 117382 6618 117466 6854
rect 117702 6618 117734 6854
rect 117114 2176 117734 6618
rect 120834 680494 121454 701760
rect 120834 680258 120866 680494
rect 121102 680258 121186 680494
rect 121422 680258 121454 680494
rect 120834 680174 121454 680258
rect 120834 679938 120866 680174
rect 121102 679938 121186 680174
rect 121422 679938 121454 680174
rect 120834 643294 121454 679938
rect 120834 643058 120866 643294
rect 121102 643058 121186 643294
rect 121422 643058 121454 643294
rect 120834 642974 121454 643058
rect 120834 642738 120866 642974
rect 121102 642738 121186 642974
rect 121422 642738 121454 642974
rect 120834 606094 121454 642738
rect 120834 605858 120866 606094
rect 121102 605858 121186 606094
rect 121422 605858 121454 606094
rect 120834 605774 121454 605858
rect 120834 605538 120866 605774
rect 121102 605538 121186 605774
rect 121422 605538 121454 605774
rect 120834 568894 121454 605538
rect 120834 568658 120866 568894
rect 121102 568658 121186 568894
rect 121422 568658 121454 568894
rect 120834 568574 121454 568658
rect 120834 568338 120866 568574
rect 121102 568338 121186 568574
rect 121422 568338 121454 568574
rect 120834 531694 121454 568338
rect 120834 531458 120866 531694
rect 121102 531458 121186 531694
rect 121422 531458 121454 531694
rect 120834 531374 121454 531458
rect 120834 531138 120866 531374
rect 121102 531138 121186 531374
rect 121422 531138 121454 531374
rect 120834 494494 121454 531138
rect 120834 494258 120866 494494
rect 121102 494258 121186 494494
rect 121422 494258 121454 494494
rect 120834 494174 121454 494258
rect 120834 493938 120866 494174
rect 121102 493938 121186 494174
rect 121422 493938 121454 494174
rect 120834 457294 121454 493938
rect 120834 457058 120866 457294
rect 121102 457058 121186 457294
rect 121422 457058 121454 457294
rect 120834 456974 121454 457058
rect 120834 456738 120866 456974
rect 121102 456738 121186 456974
rect 121422 456738 121454 456974
rect 120834 420094 121454 456738
rect 120834 419858 120866 420094
rect 121102 419858 121186 420094
rect 121422 419858 121454 420094
rect 120834 419774 121454 419858
rect 120834 419538 120866 419774
rect 121102 419538 121186 419774
rect 121422 419538 121454 419774
rect 120834 382894 121454 419538
rect 120834 382658 120866 382894
rect 121102 382658 121186 382894
rect 121422 382658 121454 382894
rect 120834 382574 121454 382658
rect 120834 382338 120866 382574
rect 121102 382338 121186 382574
rect 121422 382338 121454 382574
rect 120834 345694 121454 382338
rect 120834 345458 120866 345694
rect 121102 345458 121186 345694
rect 121422 345458 121454 345694
rect 120834 345374 121454 345458
rect 120834 345138 120866 345374
rect 121102 345138 121186 345374
rect 121422 345138 121454 345374
rect 120834 308494 121454 345138
rect 120834 308258 120866 308494
rect 121102 308258 121186 308494
rect 121422 308258 121454 308494
rect 120834 308174 121454 308258
rect 120834 307938 120866 308174
rect 121102 307938 121186 308174
rect 121422 307938 121454 308174
rect 120834 271294 121454 307938
rect 120834 271058 120866 271294
rect 121102 271058 121186 271294
rect 121422 271058 121454 271294
rect 120834 270974 121454 271058
rect 120834 270738 120866 270974
rect 121102 270738 121186 270974
rect 121422 270738 121454 270974
rect 120834 234094 121454 270738
rect 120834 233858 120866 234094
rect 121102 233858 121186 234094
rect 121422 233858 121454 234094
rect 120834 233774 121454 233858
rect 120834 233538 120866 233774
rect 121102 233538 121186 233774
rect 121422 233538 121454 233774
rect 120834 196894 121454 233538
rect 120834 196658 120866 196894
rect 121102 196658 121186 196894
rect 121422 196658 121454 196894
rect 120834 196574 121454 196658
rect 120834 196338 120866 196574
rect 121102 196338 121186 196574
rect 121422 196338 121454 196574
rect 120834 159694 121454 196338
rect 120834 159458 120866 159694
rect 121102 159458 121186 159694
rect 121422 159458 121454 159694
rect 120834 159374 121454 159458
rect 120834 159138 120866 159374
rect 121102 159138 121186 159374
rect 121422 159138 121454 159374
rect 120834 122494 121454 159138
rect 120834 122258 120866 122494
rect 121102 122258 121186 122494
rect 121422 122258 121454 122494
rect 120834 122174 121454 122258
rect 120834 121938 120866 122174
rect 121102 121938 121186 122174
rect 121422 121938 121454 122174
rect 120834 85294 121454 121938
rect 120834 85058 120866 85294
rect 121102 85058 121186 85294
rect 121422 85058 121454 85294
rect 120834 84974 121454 85058
rect 120834 84738 120866 84974
rect 121102 84738 121186 84974
rect 121422 84738 121454 84974
rect 120834 48094 121454 84738
rect 120834 47858 120866 48094
rect 121102 47858 121186 48094
rect 121422 47858 121454 48094
rect 120834 47774 121454 47858
rect 120834 47538 120866 47774
rect 121102 47538 121186 47774
rect 121422 47538 121454 47774
rect 120834 10894 121454 47538
rect 120834 10658 120866 10894
rect 121102 10658 121186 10894
rect 121422 10658 121454 10894
rect 120834 10574 121454 10658
rect 120834 10338 120866 10574
rect 121102 10338 121186 10574
rect 121422 10338 121454 10574
rect 120834 2176 121454 10338
rect 124554 684214 125174 701760
rect 124554 683978 124586 684214
rect 124822 683978 124906 684214
rect 125142 683978 125174 684214
rect 124554 683894 125174 683978
rect 124554 683658 124586 683894
rect 124822 683658 124906 683894
rect 125142 683658 125174 683894
rect 124554 647014 125174 683658
rect 124554 646778 124586 647014
rect 124822 646778 124906 647014
rect 125142 646778 125174 647014
rect 124554 646694 125174 646778
rect 124554 646458 124586 646694
rect 124822 646458 124906 646694
rect 125142 646458 125174 646694
rect 124554 609814 125174 646458
rect 124554 609578 124586 609814
rect 124822 609578 124906 609814
rect 125142 609578 125174 609814
rect 124554 609494 125174 609578
rect 124554 609258 124586 609494
rect 124822 609258 124906 609494
rect 125142 609258 125174 609494
rect 124554 572614 125174 609258
rect 124554 572378 124586 572614
rect 124822 572378 124906 572614
rect 125142 572378 125174 572614
rect 124554 572294 125174 572378
rect 124554 572058 124586 572294
rect 124822 572058 124906 572294
rect 125142 572058 125174 572294
rect 124554 535414 125174 572058
rect 124554 535178 124586 535414
rect 124822 535178 124906 535414
rect 125142 535178 125174 535414
rect 124554 535094 125174 535178
rect 124554 534858 124586 535094
rect 124822 534858 124906 535094
rect 125142 534858 125174 535094
rect 124554 498214 125174 534858
rect 124554 497978 124586 498214
rect 124822 497978 124906 498214
rect 125142 497978 125174 498214
rect 124554 497894 125174 497978
rect 124554 497658 124586 497894
rect 124822 497658 124906 497894
rect 125142 497658 125174 497894
rect 124554 461014 125174 497658
rect 124554 460778 124586 461014
rect 124822 460778 124906 461014
rect 125142 460778 125174 461014
rect 124554 460694 125174 460778
rect 124554 460458 124586 460694
rect 124822 460458 124906 460694
rect 125142 460458 125174 460694
rect 124554 423814 125174 460458
rect 124554 423578 124586 423814
rect 124822 423578 124906 423814
rect 125142 423578 125174 423814
rect 124554 423494 125174 423578
rect 124554 423258 124586 423494
rect 124822 423258 124906 423494
rect 125142 423258 125174 423494
rect 124554 386614 125174 423258
rect 124554 386378 124586 386614
rect 124822 386378 124906 386614
rect 125142 386378 125174 386614
rect 124554 386294 125174 386378
rect 124554 386058 124586 386294
rect 124822 386058 124906 386294
rect 125142 386058 125174 386294
rect 124554 349414 125174 386058
rect 124554 349178 124586 349414
rect 124822 349178 124906 349414
rect 125142 349178 125174 349414
rect 124554 349094 125174 349178
rect 124554 348858 124586 349094
rect 124822 348858 124906 349094
rect 125142 348858 125174 349094
rect 124554 312214 125174 348858
rect 124554 311978 124586 312214
rect 124822 311978 124906 312214
rect 125142 311978 125174 312214
rect 124554 311894 125174 311978
rect 124554 311658 124586 311894
rect 124822 311658 124906 311894
rect 125142 311658 125174 311894
rect 124554 275014 125174 311658
rect 124554 274778 124586 275014
rect 124822 274778 124906 275014
rect 125142 274778 125174 275014
rect 124554 274694 125174 274778
rect 124554 274458 124586 274694
rect 124822 274458 124906 274694
rect 125142 274458 125174 274694
rect 124554 237814 125174 274458
rect 124554 237578 124586 237814
rect 124822 237578 124906 237814
rect 125142 237578 125174 237814
rect 124554 237494 125174 237578
rect 124554 237258 124586 237494
rect 124822 237258 124906 237494
rect 125142 237258 125174 237494
rect 124554 200614 125174 237258
rect 124554 200378 124586 200614
rect 124822 200378 124906 200614
rect 125142 200378 125174 200614
rect 124554 200294 125174 200378
rect 124554 200058 124586 200294
rect 124822 200058 124906 200294
rect 125142 200058 125174 200294
rect 124554 163414 125174 200058
rect 124554 163178 124586 163414
rect 124822 163178 124906 163414
rect 125142 163178 125174 163414
rect 124554 163094 125174 163178
rect 124554 162858 124586 163094
rect 124822 162858 124906 163094
rect 125142 162858 125174 163094
rect 124554 126214 125174 162858
rect 124554 125978 124586 126214
rect 124822 125978 124906 126214
rect 125142 125978 125174 126214
rect 124554 125894 125174 125978
rect 124554 125658 124586 125894
rect 124822 125658 124906 125894
rect 125142 125658 125174 125894
rect 124554 89014 125174 125658
rect 124554 88778 124586 89014
rect 124822 88778 124906 89014
rect 125142 88778 125174 89014
rect 124554 88694 125174 88778
rect 124554 88458 124586 88694
rect 124822 88458 124906 88694
rect 125142 88458 125174 88694
rect 124554 51814 125174 88458
rect 124554 51578 124586 51814
rect 124822 51578 124906 51814
rect 125142 51578 125174 51814
rect 124554 51494 125174 51578
rect 124554 51258 124586 51494
rect 124822 51258 124906 51494
rect 125142 51258 125174 51494
rect 124554 14614 125174 51258
rect 124554 14378 124586 14614
rect 124822 14378 124906 14614
rect 125142 14378 125174 14614
rect 124554 14294 125174 14378
rect 124554 14058 124586 14294
rect 124822 14058 124906 14294
rect 125142 14058 125174 14294
rect 124554 2176 125174 14058
rect 128274 687934 128894 701760
rect 128274 687698 128306 687934
rect 128542 687698 128626 687934
rect 128862 687698 128894 687934
rect 128274 687614 128894 687698
rect 128274 687378 128306 687614
rect 128542 687378 128626 687614
rect 128862 687378 128894 687614
rect 128274 650734 128894 687378
rect 128274 650498 128306 650734
rect 128542 650498 128626 650734
rect 128862 650498 128894 650734
rect 128274 650414 128894 650498
rect 128274 650178 128306 650414
rect 128542 650178 128626 650414
rect 128862 650178 128894 650414
rect 128274 613534 128894 650178
rect 128274 613298 128306 613534
rect 128542 613298 128626 613534
rect 128862 613298 128894 613534
rect 128274 613214 128894 613298
rect 128274 612978 128306 613214
rect 128542 612978 128626 613214
rect 128862 612978 128894 613214
rect 128274 576334 128894 612978
rect 128274 576098 128306 576334
rect 128542 576098 128626 576334
rect 128862 576098 128894 576334
rect 128274 576014 128894 576098
rect 128274 575778 128306 576014
rect 128542 575778 128626 576014
rect 128862 575778 128894 576014
rect 128274 539134 128894 575778
rect 128274 538898 128306 539134
rect 128542 538898 128626 539134
rect 128862 538898 128894 539134
rect 128274 538814 128894 538898
rect 128274 538578 128306 538814
rect 128542 538578 128626 538814
rect 128862 538578 128894 538814
rect 128274 501934 128894 538578
rect 128274 501698 128306 501934
rect 128542 501698 128626 501934
rect 128862 501698 128894 501934
rect 128274 501614 128894 501698
rect 128274 501378 128306 501614
rect 128542 501378 128626 501614
rect 128862 501378 128894 501614
rect 128274 464734 128894 501378
rect 128274 464498 128306 464734
rect 128542 464498 128626 464734
rect 128862 464498 128894 464734
rect 128274 464414 128894 464498
rect 128274 464178 128306 464414
rect 128542 464178 128626 464414
rect 128862 464178 128894 464414
rect 128274 427534 128894 464178
rect 128274 427298 128306 427534
rect 128542 427298 128626 427534
rect 128862 427298 128894 427534
rect 128274 427214 128894 427298
rect 128274 426978 128306 427214
rect 128542 426978 128626 427214
rect 128862 426978 128894 427214
rect 128274 390334 128894 426978
rect 128274 390098 128306 390334
rect 128542 390098 128626 390334
rect 128862 390098 128894 390334
rect 128274 390014 128894 390098
rect 128274 389778 128306 390014
rect 128542 389778 128626 390014
rect 128862 389778 128894 390014
rect 128274 353134 128894 389778
rect 128274 352898 128306 353134
rect 128542 352898 128626 353134
rect 128862 352898 128894 353134
rect 128274 352814 128894 352898
rect 128274 352578 128306 352814
rect 128542 352578 128626 352814
rect 128862 352578 128894 352814
rect 128274 315934 128894 352578
rect 128274 315698 128306 315934
rect 128542 315698 128626 315934
rect 128862 315698 128894 315934
rect 128274 315614 128894 315698
rect 128274 315378 128306 315614
rect 128542 315378 128626 315614
rect 128862 315378 128894 315614
rect 128274 278734 128894 315378
rect 128274 278498 128306 278734
rect 128542 278498 128626 278734
rect 128862 278498 128894 278734
rect 128274 278414 128894 278498
rect 128274 278178 128306 278414
rect 128542 278178 128626 278414
rect 128862 278178 128894 278414
rect 128274 241534 128894 278178
rect 128274 241298 128306 241534
rect 128542 241298 128626 241534
rect 128862 241298 128894 241534
rect 128274 241214 128894 241298
rect 128274 240978 128306 241214
rect 128542 240978 128626 241214
rect 128862 240978 128894 241214
rect 128274 204334 128894 240978
rect 128274 204098 128306 204334
rect 128542 204098 128626 204334
rect 128862 204098 128894 204334
rect 128274 204014 128894 204098
rect 128274 203778 128306 204014
rect 128542 203778 128626 204014
rect 128862 203778 128894 204014
rect 128274 167134 128894 203778
rect 128274 166898 128306 167134
rect 128542 166898 128626 167134
rect 128862 166898 128894 167134
rect 128274 166814 128894 166898
rect 128274 166578 128306 166814
rect 128542 166578 128626 166814
rect 128862 166578 128894 166814
rect 128274 129934 128894 166578
rect 128274 129698 128306 129934
rect 128542 129698 128626 129934
rect 128862 129698 128894 129934
rect 128274 129614 128894 129698
rect 128274 129378 128306 129614
rect 128542 129378 128626 129614
rect 128862 129378 128894 129614
rect 128274 92734 128894 129378
rect 128274 92498 128306 92734
rect 128542 92498 128626 92734
rect 128862 92498 128894 92734
rect 128274 92414 128894 92498
rect 128274 92178 128306 92414
rect 128542 92178 128626 92414
rect 128862 92178 128894 92414
rect 128274 55534 128894 92178
rect 128274 55298 128306 55534
rect 128542 55298 128626 55534
rect 128862 55298 128894 55534
rect 128274 55214 128894 55298
rect 128274 54978 128306 55214
rect 128542 54978 128626 55214
rect 128862 54978 128894 55214
rect 128274 18334 128894 54978
rect 128274 18098 128306 18334
rect 128542 18098 128626 18334
rect 128862 18098 128894 18334
rect 128274 18014 128894 18098
rect 128274 17778 128306 18014
rect 128542 17778 128626 18014
rect 128862 17778 128894 18014
rect 128274 2176 128894 17778
rect 131994 691654 132614 701760
rect 131994 691418 132026 691654
rect 132262 691418 132346 691654
rect 132582 691418 132614 691654
rect 131994 691334 132614 691418
rect 131994 691098 132026 691334
rect 132262 691098 132346 691334
rect 132582 691098 132614 691334
rect 131994 654454 132614 691098
rect 131994 654218 132026 654454
rect 132262 654218 132346 654454
rect 132582 654218 132614 654454
rect 131994 654134 132614 654218
rect 131994 653898 132026 654134
rect 132262 653898 132346 654134
rect 132582 653898 132614 654134
rect 131994 617254 132614 653898
rect 131994 617018 132026 617254
rect 132262 617018 132346 617254
rect 132582 617018 132614 617254
rect 131994 616934 132614 617018
rect 131994 616698 132026 616934
rect 132262 616698 132346 616934
rect 132582 616698 132614 616934
rect 131994 580054 132614 616698
rect 131994 579818 132026 580054
rect 132262 579818 132346 580054
rect 132582 579818 132614 580054
rect 131994 579734 132614 579818
rect 131994 579498 132026 579734
rect 132262 579498 132346 579734
rect 132582 579498 132614 579734
rect 131994 542854 132614 579498
rect 131994 542618 132026 542854
rect 132262 542618 132346 542854
rect 132582 542618 132614 542854
rect 131994 542534 132614 542618
rect 131994 542298 132026 542534
rect 132262 542298 132346 542534
rect 132582 542298 132614 542534
rect 131994 505654 132614 542298
rect 131994 505418 132026 505654
rect 132262 505418 132346 505654
rect 132582 505418 132614 505654
rect 131994 505334 132614 505418
rect 131994 505098 132026 505334
rect 132262 505098 132346 505334
rect 132582 505098 132614 505334
rect 131994 468454 132614 505098
rect 131994 468218 132026 468454
rect 132262 468218 132346 468454
rect 132582 468218 132614 468454
rect 131994 468134 132614 468218
rect 131994 467898 132026 468134
rect 132262 467898 132346 468134
rect 132582 467898 132614 468134
rect 131994 431254 132614 467898
rect 131994 431018 132026 431254
rect 132262 431018 132346 431254
rect 132582 431018 132614 431254
rect 131994 430934 132614 431018
rect 131994 430698 132026 430934
rect 132262 430698 132346 430934
rect 132582 430698 132614 430934
rect 131994 394054 132614 430698
rect 131994 393818 132026 394054
rect 132262 393818 132346 394054
rect 132582 393818 132614 394054
rect 131994 393734 132614 393818
rect 131994 393498 132026 393734
rect 132262 393498 132346 393734
rect 132582 393498 132614 393734
rect 131994 356854 132614 393498
rect 131994 356618 132026 356854
rect 132262 356618 132346 356854
rect 132582 356618 132614 356854
rect 131994 356534 132614 356618
rect 131994 356298 132026 356534
rect 132262 356298 132346 356534
rect 132582 356298 132614 356534
rect 131994 319654 132614 356298
rect 131994 319418 132026 319654
rect 132262 319418 132346 319654
rect 132582 319418 132614 319654
rect 131994 319334 132614 319418
rect 131994 319098 132026 319334
rect 132262 319098 132346 319334
rect 132582 319098 132614 319334
rect 131994 282454 132614 319098
rect 131994 282218 132026 282454
rect 132262 282218 132346 282454
rect 132582 282218 132614 282454
rect 131994 282134 132614 282218
rect 131994 281898 132026 282134
rect 132262 281898 132346 282134
rect 132582 281898 132614 282134
rect 131994 245254 132614 281898
rect 131994 245018 132026 245254
rect 132262 245018 132346 245254
rect 132582 245018 132614 245254
rect 131994 244934 132614 245018
rect 131994 244698 132026 244934
rect 132262 244698 132346 244934
rect 132582 244698 132614 244934
rect 131994 208054 132614 244698
rect 131994 207818 132026 208054
rect 132262 207818 132346 208054
rect 132582 207818 132614 208054
rect 131994 207734 132614 207818
rect 131994 207498 132026 207734
rect 132262 207498 132346 207734
rect 132582 207498 132614 207734
rect 131994 170854 132614 207498
rect 131994 170618 132026 170854
rect 132262 170618 132346 170854
rect 132582 170618 132614 170854
rect 131994 170534 132614 170618
rect 131994 170298 132026 170534
rect 132262 170298 132346 170534
rect 132582 170298 132614 170534
rect 131994 133654 132614 170298
rect 131994 133418 132026 133654
rect 132262 133418 132346 133654
rect 132582 133418 132614 133654
rect 131994 133334 132614 133418
rect 131994 133098 132026 133334
rect 132262 133098 132346 133334
rect 132582 133098 132614 133334
rect 131994 96454 132614 133098
rect 131994 96218 132026 96454
rect 132262 96218 132346 96454
rect 132582 96218 132614 96454
rect 131994 96134 132614 96218
rect 131994 95898 132026 96134
rect 132262 95898 132346 96134
rect 132582 95898 132614 96134
rect 131994 59254 132614 95898
rect 131994 59018 132026 59254
rect 132262 59018 132346 59254
rect 132582 59018 132614 59254
rect 131994 58934 132614 59018
rect 131994 58698 132026 58934
rect 132262 58698 132346 58934
rect 132582 58698 132614 58934
rect 131994 22054 132614 58698
rect 131994 21818 132026 22054
rect 132262 21818 132346 22054
rect 132582 21818 132614 22054
rect 131994 21734 132614 21818
rect 131994 21498 132026 21734
rect 132262 21498 132346 21734
rect 132582 21498 132614 21734
rect 131994 2176 132614 21498
rect 135714 695374 136334 701760
rect 135714 695138 135746 695374
rect 135982 695138 136066 695374
rect 136302 695138 136334 695374
rect 135714 695054 136334 695138
rect 135714 694818 135746 695054
rect 135982 694818 136066 695054
rect 136302 694818 136334 695054
rect 135714 658174 136334 694818
rect 135714 657938 135746 658174
rect 135982 657938 136066 658174
rect 136302 657938 136334 658174
rect 135714 657854 136334 657938
rect 135714 657618 135746 657854
rect 135982 657618 136066 657854
rect 136302 657618 136334 657854
rect 135714 620974 136334 657618
rect 135714 620738 135746 620974
rect 135982 620738 136066 620974
rect 136302 620738 136334 620974
rect 135714 620654 136334 620738
rect 135714 620418 135746 620654
rect 135982 620418 136066 620654
rect 136302 620418 136334 620654
rect 135714 583774 136334 620418
rect 135714 583538 135746 583774
rect 135982 583538 136066 583774
rect 136302 583538 136334 583774
rect 135714 583454 136334 583538
rect 135714 583218 135746 583454
rect 135982 583218 136066 583454
rect 136302 583218 136334 583454
rect 135714 546574 136334 583218
rect 135714 546338 135746 546574
rect 135982 546338 136066 546574
rect 136302 546338 136334 546574
rect 135714 546254 136334 546338
rect 135714 546018 135746 546254
rect 135982 546018 136066 546254
rect 136302 546018 136334 546254
rect 135714 509374 136334 546018
rect 135714 509138 135746 509374
rect 135982 509138 136066 509374
rect 136302 509138 136334 509374
rect 135714 509054 136334 509138
rect 135714 508818 135746 509054
rect 135982 508818 136066 509054
rect 136302 508818 136334 509054
rect 135714 472174 136334 508818
rect 135714 471938 135746 472174
rect 135982 471938 136066 472174
rect 136302 471938 136334 472174
rect 135714 471854 136334 471938
rect 135714 471618 135746 471854
rect 135982 471618 136066 471854
rect 136302 471618 136334 471854
rect 135714 434974 136334 471618
rect 135714 434738 135746 434974
rect 135982 434738 136066 434974
rect 136302 434738 136334 434974
rect 135714 434654 136334 434738
rect 135714 434418 135746 434654
rect 135982 434418 136066 434654
rect 136302 434418 136334 434654
rect 135714 397774 136334 434418
rect 135714 397538 135746 397774
rect 135982 397538 136066 397774
rect 136302 397538 136334 397774
rect 135714 397454 136334 397538
rect 135714 397218 135746 397454
rect 135982 397218 136066 397454
rect 136302 397218 136334 397454
rect 135714 360574 136334 397218
rect 135714 360338 135746 360574
rect 135982 360338 136066 360574
rect 136302 360338 136334 360574
rect 135714 360254 136334 360338
rect 135714 360018 135746 360254
rect 135982 360018 136066 360254
rect 136302 360018 136334 360254
rect 135714 323374 136334 360018
rect 135714 323138 135746 323374
rect 135982 323138 136066 323374
rect 136302 323138 136334 323374
rect 135714 323054 136334 323138
rect 135714 322818 135746 323054
rect 135982 322818 136066 323054
rect 136302 322818 136334 323054
rect 135714 286174 136334 322818
rect 135714 285938 135746 286174
rect 135982 285938 136066 286174
rect 136302 285938 136334 286174
rect 135714 285854 136334 285938
rect 135714 285618 135746 285854
rect 135982 285618 136066 285854
rect 136302 285618 136334 285854
rect 135714 248974 136334 285618
rect 135714 248738 135746 248974
rect 135982 248738 136066 248974
rect 136302 248738 136334 248974
rect 135714 248654 136334 248738
rect 135714 248418 135746 248654
rect 135982 248418 136066 248654
rect 136302 248418 136334 248654
rect 135714 211774 136334 248418
rect 135714 211538 135746 211774
rect 135982 211538 136066 211774
rect 136302 211538 136334 211774
rect 135714 211454 136334 211538
rect 135714 211218 135746 211454
rect 135982 211218 136066 211454
rect 136302 211218 136334 211454
rect 135714 174574 136334 211218
rect 135714 174338 135746 174574
rect 135982 174338 136066 174574
rect 136302 174338 136334 174574
rect 135714 174254 136334 174338
rect 135714 174018 135746 174254
rect 135982 174018 136066 174254
rect 136302 174018 136334 174254
rect 135714 137374 136334 174018
rect 135714 137138 135746 137374
rect 135982 137138 136066 137374
rect 136302 137138 136334 137374
rect 135714 137054 136334 137138
rect 135714 136818 135746 137054
rect 135982 136818 136066 137054
rect 136302 136818 136334 137054
rect 135714 100174 136334 136818
rect 135714 99938 135746 100174
rect 135982 99938 136066 100174
rect 136302 99938 136334 100174
rect 135714 99854 136334 99938
rect 135714 99618 135746 99854
rect 135982 99618 136066 99854
rect 136302 99618 136334 99854
rect 135714 62974 136334 99618
rect 135714 62738 135746 62974
rect 135982 62738 136066 62974
rect 136302 62738 136334 62974
rect 135714 62654 136334 62738
rect 135714 62418 135746 62654
rect 135982 62418 136066 62654
rect 136302 62418 136334 62654
rect 135714 25774 136334 62418
rect 135714 25538 135746 25774
rect 135982 25538 136066 25774
rect 136302 25538 136334 25774
rect 135714 25454 136334 25538
rect 135714 25218 135746 25454
rect 135982 25218 136066 25454
rect 136302 25218 136334 25454
rect 135714 2176 136334 25218
rect 139434 699094 140054 701760
rect 139434 698858 139466 699094
rect 139702 698858 139786 699094
rect 140022 698858 140054 699094
rect 139434 698774 140054 698858
rect 139434 698538 139466 698774
rect 139702 698538 139786 698774
rect 140022 698538 140054 698774
rect 139434 661894 140054 698538
rect 139434 661658 139466 661894
rect 139702 661658 139786 661894
rect 140022 661658 140054 661894
rect 139434 661574 140054 661658
rect 139434 661338 139466 661574
rect 139702 661338 139786 661574
rect 140022 661338 140054 661574
rect 139434 624694 140054 661338
rect 139434 624458 139466 624694
rect 139702 624458 139786 624694
rect 140022 624458 140054 624694
rect 139434 624374 140054 624458
rect 139434 624138 139466 624374
rect 139702 624138 139786 624374
rect 140022 624138 140054 624374
rect 139434 587494 140054 624138
rect 139434 587258 139466 587494
rect 139702 587258 139786 587494
rect 140022 587258 140054 587494
rect 139434 587174 140054 587258
rect 139434 586938 139466 587174
rect 139702 586938 139786 587174
rect 140022 586938 140054 587174
rect 139434 550294 140054 586938
rect 139434 550058 139466 550294
rect 139702 550058 139786 550294
rect 140022 550058 140054 550294
rect 139434 549974 140054 550058
rect 139434 549738 139466 549974
rect 139702 549738 139786 549974
rect 140022 549738 140054 549974
rect 139434 513094 140054 549738
rect 139434 512858 139466 513094
rect 139702 512858 139786 513094
rect 140022 512858 140054 513094
rect 139434 512774 140054 512858
rect 139434 512538 139466 512774
rect 139702 512538 139786 512774
rect 140022 512538 140054 512774
rect 139434 475894 140054 512538
rect 139434 475658 139466 475894
rect 139702 475658 139786 475894
rect 140022 475658 140054 475894
rect 139434 475574 140054 475658
rect 139434 475338 139466 475574
rect 139702 475338 139786 475574
rect 140022 475338 140054 475574
rect 139434 438694 140054 475338
rect 139434 438458 139466 438694
rect 139702 438458 139786 438694
rect 140022 438458 140054 438694
rect 139434 438374 140054 438458
rect 139434 438138 139466 438374
rect 139702 438138 139786 438374
rect 140022 438138 140054 438374
rect 139434 401494 140054 438138
rect 139434 401258 139466 401494
rect 139702 401258 139786 401494
rect 140022 401258 140054 401494
rect 139434 401174 140054 401258
rect 139434 400938 139466 401174
rect 139702 400938 139786 401174
rect 140022 400938 140054 401174
rect 139434 364294 140054 400938
rect 139434 364058 139466 364294
rect 139702 364058 139786 364294
rect 140022 364058 140054 364294
rect 139434 363974 140054 364058
rect 139434 363738 139466 363974
rect 139702 363738 139786 363974
rect 140022 363738 140054 363974
rect 139434 327094 140054 363738
rect 139434 326858 139466 327094
rect 139702 326858 139786 327094
rect 140022 326858 140054 327094
rect 139434 326774 140054 326858
rect 139434 326538 139466 326774
rect 139702 326538 139786 326774
rect 140022 326538 140054 326774
rect 139434 289894 140054 326538
rect 139434 289658 139466 289894
rect 139702 289658 139786 289894
rect 140022 289658 140054 289894
rect 139434 289574 140054 289658
rect 139434 289338 139466 289574
rect 139702 289338 139786 289574
rect 140022 289338 140054 289574
rect 139434 252694 140054 289338
rect 139434 252458 139466 252694
rect 139702 252458 139786 252694
rect 140022 252458 140054 252694
rect 139434 252374 140054 252458
rect 139434 252138 139466 252374
rect 139702 252138 139786 252374
rect 140022 252138 140054 252374
rect 139434 215494 140054 252138
rect 139434 215258 139466 215494
rect 139702 215258 139786 215494
rect 140022 215258 140054 215494
rect 139434 215174 140054 215258
rect 139434 214938 139466 215174
rect 139702 214938 139786 215174
rect 140022 214938 140054 215174
rect 139434 178294 140054 214938
rect 139434 178058 139466 178294
rect 139702 178058 139786 178294
rect 140022 178058 140054 178294
rect 139434 177974 140054 178058
rect 139434 177738 139466 177974
rect 139702 177738 139786 177974
rect 140022 177738 140054 177974
rect 139434 141094 140054 177738
rect 139434 140858 139466 141094
rect 139702 140858 139786 141094
rect 140022 140858 140054 141094
rect 139434 140774 140054 140858
rect 139434 140538 139466 140774
rect 139702 140538 139786 140774
rect 140022 140538 140054 140774
rect 139434 103894 140054 140538
rect 139434 103658 139466 103894
rect 139702 103658 139786 103894
rect 140022 103658 140054 103894
rect 139434 103574 140054 103658
rect 139434 103338 139466 103574
rect 139702 103338 139786 103574
rect 140022 103338 140054 103574
rect 139434 66694 140054 103338
rect 139434 66458 139466 66694
rect 139702 66458 139786 66694
rect 140022 66458 140054 66694
rect 139434 66374 140054 66458
rect 139434 66138 139466 66374
rect 139702 66138 139786 66374
rect 140022 66138 140054 66374
rect 139434 29494 140054 66138
rect 139434 29258 139466 29494
rect 139702 29258 139786 29494
rect 140022 29258 140054 29494
rect 139434 29174 140054 29258
rect 139434 28938 139466 29174
rect 139702 28938 139786 29174
rect 140022 28938 140054 29174
rect 139434 2176 140054 28938
rect 150594 673054 151214 701760
rect 150594 672818 150626 673054
rect 150862 672818 150946 673054
rect 151182 672818 151214 673054
rect 150594 672734 151214 672818
rect 150594 672498 150626 672734
rect 150862 672498 150946 672734
rect 151182 672498 151214 672734
rect 150594 635854 151214 672498
rect 150594 635618 150626 635854
rect 150862 635618 150946 635854
rect 151182 635618 151214 635854
rect 150594 635534 151214 635618
rect 150594 635298 150626 635534
rect 150862 635298 150946 635534
rect 151182 635298 151214 635534
rect 150594 598654 151214 635298
rect 150594 598418 150626 598654
rect 150862 598418 150946 598654
rect 151182 598418 151214 598654
rect 150594 598334 151214 598418
rect 150594 598098 150626 598334
rect 150862 598098 150946 598334
rect 151182 598098 151214 598334
rect 150594 561454 151214 598098
rect 150594 561218 150626 561454
rect 150862 561218 150946 561454
rect 151182 561218 151214 561454
rect 150594 561134 151214 561218
rect 150594 560898 150626 561134
rect 150862 560898 150946 561134
rect 151182 560898 151214 561134
rect 150594 524254 151214 560898
rect 150594 524018 150626 524254
rect 150862 524018 150946 524254
rect 151182 524018 151214 524254
rect 150594 523934 151214 524018
rect 150594 523698 150626 523934
rect 150862 523698 150946 523934
rect 151182 523698 151214 523934
rect 150594 487054 151214 523698
rect 150594 486818 150626 487054
rect 150862 486818 150946 487054
rect 151182 486818 151214 487054
rect 150594 486734 151214 486818
rect 150594 486498 150626 486734
rect 150862 486498 150946 486734
rect 151182 486498 151214 486734
rect 150594 449854 151214 486498
rect 150594 449618 150626 449854
rect 150862 449618 150946 449854
rect 151182 449618 151214 449854
rect 150594 449534 151214 449618
rect 150594 449298 150626 449534
rect 150862 449298 150946 449534
rect 151182 449298 151214 449534
rect 150594 412654 151214 449298
rect 150594 412418 150626 412654
rect 150862 412418 150946 412654
rect 151182 412418 151214 412654
rect 150594 412334 151214 412418
rect 150594 412098 150626 412334
rect 150862 412098 150946 412334
rect 151182 412098 151214 412334
rect 150594 375454 151214 412098
rect 150594 375218 150626 375454
rect 150862 375218 150946 375454
rect 151182 375218 151214 375454
rect 150594 375134 151214 375218
rect 150594 374898 150626 375134
rect 150862 374898 150946 375134
rect 151182 374898 151214 375134
rect 150594 338254 151214 374898
rect 150594 338018 150626 338254
rect 150862 338018 150946 338254
rect 151182 338018 151214 338254
rect 150594 337934 151214 338018
rect 150594 337698 150626 337934
rect 150862 337698 150946 337934
rect 151182 337698 151214 337934
rect 150594 301054 151214 337698
rect 150594 300818 150626 301054
rect 150862 300818 150946 301054
rect 151182 300818 151214 301054
rect 150594 300734 151214 300818
rect 150594 300498 150626 300734
rect 150862 300498 150946 300734
rect 151182 300498 151214 300734
rect 150594 263854 151214 300498
rect 150594 263618 150626 263854
rect 150862 263618 150946 263854
rect 151182 263618 151214 263854
rect 150594 263534 151214 263618
rect 150594 263298 150626 263534
rect 150862 263298 150946 263534
rect 151182 263298 151214 263534
rect 150594 226654 151214 263298
rect 150594 226418 150626 226654
rect 150862 226418 150946 226654
rect 151182 226418 151214 226654
rect 150594 226334 151214 226418
rect 150594 226098 150626 226334
rect 150862 226098 150946 226334
rect 151182 226098 151214 226334
rect 150594 189454 151214 226098
rect 150594 189218 150626 189454
rect 150862 189218 150946 189454
rect 151182 189218 151214 189454
rect 150594 189134 151214 189218
rect 150594 188898 150626 189134
rect 150862 188898 150946 189134
rect 151182 188898 151214 189134
rect 150594 152254 151214 188898
rect 150594 152018 150626 152254
rect 150862 152018 150946 152254
rect 151182 152018 151214 152254
rect 150594 151934 151214 152018
rect 150594 151698 150626 151934
rect 150862 151698 150946 151934
rect 151182 151698 151214 151934
rect 150594 115054 151214 151698
rect 150594 114818 150626 115054
rect 150862 114818 150946 115054
rect 151182 114818 151214 115054
rect 150594 114734 151214 114818
rect 150594 114498 150626 114734
rect 150862 114498 150946 114734
rect 151182 114498 151214 114734
rect 150594 77854 151214 114498
rect 150594 77618 150626 77854
rect 150862 77618 150946 77854
rect 151182 77618 151214 77854
rect 150594 77534 151214 77618
rect 150594 77298 150626 77534
rect 150862 77298 150946 77534
rect 151182 77298 151214 77534
rect 150594 40654 151214 77298
rect 150594 40418 150626 40654
rect 150862 40418 150946 40654
rect 151182 40418 151214 40654
rect 150594 40334 151214 40418
rect 150594 40098 150626 40334
rect 150862 40098 150946 40334
rect 151182 40098 151214 40334
rect 150594 3454 151214 40098
rect 150594 3218 150626 3454
rect 150862 3218 150946 3454
rect 151182 3218 151214 3454
rect 150594 3134 151214 3218
rect 150594 2898 150626 3134
rect 150862 2898 150946 3134
rect 151182 2898 151214 3134
rect 150594 2176 151214 2898
rect 154314 676774 154934 701760
rect 154314 676538 154346 676774
rect 154582 676538 154666 676774
rect 154902 676538 154934 676774
rect 154314 676454 154934 676538
rect 154314 676218 154346 676454
rect 154582 676218 154666 676454
rect 154902 676218 154934 676454
rect 154314 639574 154934 676218
rect 154314 639338 154346 639574
rect 154582 639338 154666 639574
rect 154902 639338 154934 639574
rect 154314 639254 154934 639338
rect 154314 639018 154346 639254
rect 154582 639018 154666 639254
rect 154902 639018 154934 639254
rect 154314 602374 154934 639018
rect 154314 602138 154346 602374
rect 154582 602138 154666 602374
rect 154902 602138 154934 602374
rect 154314 602054 154934 602138
rect 154314 601818 154346 602054
rect 154582 601818 154666 602054
rect 154902 601818 154934 602054
rect 154314 565174 154934 601818
rect 154314 564938 154346 565174
rect 154582 564938 154666 565174
rect 154902 564938 154934 565174
rect 154314 564854 154934 564938
rect 154314 564618 154346 564854
rect 154582 564618 154666 564854
rect 154902 564618 154934 564854
rect 154314 527974 154934 564618
rect 154314 527738 154346 527974
rect 154582 527738 154666 527974
rect 154902 527738 154934 527974
rect 154314 527654 154934 527738
rect 154314 527418 154346 527654
rect 154582 527418 154666 527654
rect 154902 527418 154934 527654
rect 154314 490774 154934 527418
rect 154314 490538 154346 490774
rect 154582 490538 154666 490774
rect 154902 490538 154934 490774
rect 154314 490454 154934 490538
rect 154314 490218 154346 490454
rect 154582 490218 154666 490454
rect 154902 490218 154934 490454
rect 154314 453574 154934 490218
rect 154314 453338 154346 453574
rect 154582 453338 154666 453574
rect 154902 453338 154934 453574
rect 154314 453254 154934 453338
rect 154314 453018 154346 453254
rect 154582 453018 154666 453254
rect 154902 453018 154934 453254
rect 154314 416374 154934 453018
rect 154314 416138 154346 416374
rect 154582 416138 154666 416374
rect 154902 416138 154934 416374
rect 154314 416054 154934 416138
rect 154314 415818 154346 416054
rect 154582 415818 154666 416054
rect 154902 415818 154934 416054
rect 154314 379174 154934 415818
rect 154314 378938 154346 379174
rect 154582 378938 154666 379174
rect 154902 378938 154934 379174
rect 154314 378854 154934 378938
rect 154314 378618 154346 378854
rect 154582 378618 154666 378854
rect 154902 378618 154934 378854
rect 154314 341974 154934 378618
rect 154314 341738 154346 341974
rect 154582 341738 154666 341974
rect 154902 341738 154934 341974
rect 154314 341654 154934 341738
rect 154314 341418 154346 341654
rect 154582 341418 154666 341654
rect 154902 341418 154934 341654
rect 154314 304774 154934 341418
rect 154314 304538 154346 304774
rect 154582 304538 154666 304774
rect 154902 304538 154934 304774
rect 154314 304454 154934 304538
rect 154314 304218 154346 304454
rect 154582 304218 154666 304454
rect 154902 304218 154934 304454
rect 154314 267574 154934 304218
rect 154314 267338 154346 267574
rect 154582 267338 154666 267574
rect 154902 267338 154934 267574
rect 154314 267254 154934 267338
rect 154314 267018 154346 267254
rect 154582 267018 154666 267254
rect 154902 267018 154934 267254
rect 154314 230374 154934 267018
rect 154314 230138 154346 230374
rect 154582 230138 154666 230374
rect 154902 230138 154934 230374
rect 154314 230054 154934 230138
rect 154314 229818 154346 230054
rect 154582 229818 154666 230054
rect 154902 229818 154934 230054
rect 154314 193174 154934 229818
rect 154314 192938 154346 193174
rect 154582 192938 154666 193174
rect 154902 192938 154934 193174
rect 154314 192854 154934 192938
rect 154314 192618 154346 192854
rect 154582 192618 154666 192854
rect 154902 192618 154934 192854
rect 154314 155974 154934 192618
rect 154314 155738 154346 155974
rect 154582 155738 154666 155974
rect 154902 155738 154934 155974
rect 154314 155654 154934 155738
rect 154314 155418 154346 155654
rect 154582 155418 154666 155654
rect 154902 155418 154934 155654
rect 154314 118774 154934 155418
rect 154314 118538 154346 118774
rect 154582 118538 154666 118774
rect 154902 118538 154934 118774
rect 154314 118454 154934 118538
rect 154314 118218 154346 118454
rect 154582 118218 154666 118454
rect 154902 118218 154934 118454
rect 154314 81574 154934 118218
rect 154314 81338 154346 81574
rect 154582 81338 154666 81574
rect 154902 81338 154934 81574
rect 154314 81254 154934 81338
rect 154314 81018 154346 81254
rect 154582 81018 154666 81254
rect 154902 81018 154934 81254
rect 154314 44374 154934 81018
rect 154314 44138 154346 44374
rect 154582 44138 154666 44374
rect 154902 44138 154934 44374
rect 154314 44054 154934 44138
rect 154314 43818 154346 44054
rect 154582 43818 154666 44054
rect 154902 43818 154934 44054
rect 154314 7174 154934 43818
rect 154314 6938 154346 7174
rect 154582 6938 154666 7174
rect 154902 6938 154934 7174
rect 154314 6854 154934 6938
rect 154314 6618 154346 6854
rect 154582 6618 154666 6854
rect 154902 6618 154934 6854
rect 154314 2176 154934 6618
rect 158034 680494 158654 701760
rect 158034 680258 158066 680494
rect 158302 680258 158386 680494
rect 158622 680258 158654 680494
rect 158034 680174 158654 680258
rect 158034 679938 158066 680174
rect 158302 679938 158386 680174
rect 158622 679938 158654 680174
rect 158034 643294 158654 679938
rect 158034 643058 158066 643294
rect 158302 643058 158386 643294
rect 158622 643058 158654 643294
rect 158034 642974 158654 643058
rect 158034 642738 158066 642974
rect 158302 642738 158386 642974
rect 158622 642738 158654 642974
rect 158034 606094 158654 642738
rect 158034 605858 158066 606094
rect 158302 605858 158386 606094
rect 158622 605858 158654 606094
rect 158034 605774 158654 605858
rect 158034 605538 158066 605774
rect 158302 605538 158386 605774
rect 158622 605538 158654 605774
rect 158034 568894 158654 605538
rect 158034 568658 158066 568894
rect 158302 568658 158386 568894
rect 158622 568658 158654 568894
rect 158034 568574 158654 568658
rect 158034 568338 158066 568574
rect 158302 568338 158386 568574
rect 158622 568338 158654 568574
rect 158034 531694 158654 568338
rect 158034 531458 158066 531694
rect 158302 531458 158386 531694
rect 158622 531458 158654 531694
rect 158034 531374 158654 531458
rect 158034 531138 158066 531374
rect 158302 531138 158386 531374
rect 158622 531138 158654 531374
rect 158034 494494 158654 531138
rect 158034 494258 158066 494494
rect 158302 494258 158386 494494
rect 158622 494258 158654 494494
rect 158034 494174 158654 494258
rect 158034 493938 158066 494174
rect 158302 493938 158386 494174
rect 158622 493938 158654 494174
rect 158034 457294 158654 493938
rect 158034 457058 158066 457294
rect 158302 457058 158386 457294
rect 158622 457058 158654 457294
rect 158034 456974 158654 457058
rect 158034 456738 158066 456974
rect 158302 456738 158386 456974
rect 158622 456738 158654 456974
rect 158034 420094 158654 456738
rect 158034 419858 158066 420094
rect 158302 419858 158386 420094
rect 158622 419858 158654 420094
rect 158034 419774 158654 419858
rect 158034 419538 158066 419774
rect 158302 419538 158386 419774
rect 158622 419538 158654 419774
rect 158034 382894 158654 419538
rect 158034 382658 158066 382894
rect 158302 382658 158386 382894
rect 158622 382658 158654 382894
rect 158034 382574 158654 382658
rect 158034 382338 158066 382574
rect 158302 382338 158386 382574
rect 158622 382338 158654 382574
rect 158034 345694 158654 382338
rect 158034 345458 158066 345694
rect 158302 345458 158386 345694
rect 158622 345458 158654 345694
rect 158034 345374 158654 345458
rect 158034 345138 158066 345374
rect 158302 345138 158386 345374
rect 158622 345138 158654 345374
rect 158034 308494 158654 345138
rect 158034 308258 158066 308494
rect 158302 308258 158386 308494
rect 158622 308258 158654 308494
rect 158034 308174 158654 308258
rect 158034 307938 158066 308174
rect 158302 307938 158386 308174
rect 158622 307938 158654 308174
rect 158034 271294 158654 307938
rect 158034 271058 158066 271294
rect 158302 271058 158386 271294
rect 158622 271058 158654 271294
rect 158034 270974 158654 271058
rect 158034 270738 158066 270974
rect 158302 270738 158386 270974
rect 158622 270738 158654 270974
rect 158034 234094 158654 270738
rect 158034 233858 158066 234094
rect 158302 233858 158386 234094
rect 158622 233858 158654 234094
rect 158034 233774 158654 233858
rect 158034 233538 158066 233774
rect 158302 233538 158386 233774
rect 158622 233538 158654 233774
rect 158034 196894 158654 233538
rect 158034 196658 158066 196894
rect 158302 196658 158386 196894
rect 158622 196658 158654 196894
rect 158034 196574 158654 196658
rect 158034 196338 158066 196574
rect 158302 196338 158386 196574
rect 158622 196338 158654 196574
rect 158034 159694 158654 196338
rect 158034 159458 158066 159694
rect 158302 159458 158386 159694
rect 158622 159458 158654 159694
rect 158034 159374 158654 159458
rect 158034 159138 158066 159374
rect 158302 159138 158386 159374
rect 158622 159138 158654 159374
rect 158034 122494 158654 159138
rect 158034 122258 158066 122494
rect 158302 122258 158386 122494
rect 158622 122258 158654 122494
rect 158034 122174 158654 122258
rect 158034 121938 158066 122174
rect 158302 121938 158386 122174
rect 158622 121938 158654 122174
rect 158034 85294 158654 121938
rect 158034 85058 158066 85294
rect 158302 85058 158386 85294
rect 158622 85058 158654 85294
rect 158034 84974 158654 85058
rect 158034 84738 158066 84974
rect 158302 84738 158386 84974
rect 158622 84738 158654 84974
rect 158034 48094 158654 84738
rect 158034 47858 158066 48094
rect 158302 47858 158386 48094
rect 158622 47858 158654 48094
rect 158034 47774 158654 47858
rect 158034 47538 158066 47774
rect 158302 47538 158386 47774
rect 158622 47538 158654 47774
rect 158034 10894 158654 47538
rect 158034 10658 158066 10894
rect 158302 10658 158386 10894
rect 158622 10658 158654 10894
rect 158034 10574 158654 10658
rect 158034 10338 158066 10574
rect 158302 10338 158386 10574
rect 158622 10338 158654 10574
rect 158034 2176 158654 10338
rect 161754 684214 162374 701760
rect 161754 683978 161786 684214
rect 162022 683978 162106 684214
rect 162342 683978 162374 684214
rect 161754 683894 162374 683978
rect 161754 683658 161786 683894
rect 162022 683658 162106 683894
rect 162342 683658 162374 683894
rect 161754 647014 162374 683658
rect 161754 646778 161786 647014
rect 162022 646778 162106 647014
rect 162342 646778 162374 647014
rect 161754 646694 162374 646778
rect 161754 646458 161786 646694
rect 162022 646458 162106 646694
rect 162342 646458 162374 646694
rect 161754 609814 162374 646458
rect 161754 609578 161786 609814
rect 162022 609578 162106 609814
rect 162342 609578 162374 609814
rect 161754 609494 162374 609578
rect 161754 609258 161786 609494
rect 162022 609258 162106 609494
rect 162342 609258 162374 609494
rect 161754 572614 162374 609258
rect 161754 572378 161786 572614
rect 162022 572378 162106 572614
rect 162342 572378 162374 572614
rect 161754 572294 162374 572378
rect 161754 572058 161786 572294
rect 162022 572058 162106 572294
rect 162342 572058 162374 572294
rect 161754 535414 162374 572058
rect 161754 535178 161786 535414
rect 162022 535178 162106 535414
rect 162342 535178 162374 535414
rect 161754 535094 162374 535178
rect 161754 534858 161786 535094
rect 162022 534858 162106 535094
rect 162342 534858 162374 535094
rect 161754 498214 162374 534858
rect 161754 497978 161786 498214
rect 162022 497978 162106 498214
rect 162342 497978 162374 498214
rect 161754 497894 162374 497978
rect 161754 497658 161786 497894
rect 162022 497658 162106 497894
rect 162342 497658 162374 497894
rect 161754 461014 162374 497658
rect 161754 460778 161786 461014
rect 162022 460778 162106 461014
rect 162342 460778 162374 461014
rect 161754 460694 162374 460778
rect 161754 460458 161786 460694
rect 162022 460458 162106 460694
rect 162342 460458 162374 460694
rect 161754 423814 162374 460458
rect 161754 423578 161786 423814
rect 162022 423578 162106 423814
rect 162342 423578 162374 423814
rect 161754 423494 162374 423578
rect 161754 423258 161786 423494
rect 162022 423258 162106 423494
rect 162342 423258 162374 423494
rect 161754 386614 162374 423258
rect 161754 386378 161786 386614
rect 162022 386378 162106 386614
rect 162342 386378 162374 386614
rect 161754 386294 162374 386378
rect 161754 386058 161786 386294
rect 162022 386058 162106 386294
rect 162342 386058 162374 386294
rect 161754 349414 162374 386058
rect 161754 349178 161786 349414
rect 162022 349178 162106 349414
rect 162342 349178 162374 349414
rect 161754 349094 162374 349178
rect 161754 348858 161786 349094
rect 162022 348858 162106 349094
rect 162342 348858 162374 349094
rect 161754 312214 162374 348858
rect 161754 311978 161786 312214
rect 162022 311978 162106 312214
rect 162342 311978 162374 312214
rect 161754 311894 162374 311978
rect 161754 311658 161786 311894
rect 162022 311658 162106 311894
rect 162342 311658 162374 311894
rect 161754 275014 162374 311658
rect 161754 274778 161786 275014
rect 162022 274778 162106 275014
rect 162342 274778 162374 275014
rect 161754 274694 162374 274778
rect 161754 274458 161786 274694
rect 162022 274458 162106 274694
rect 162342 274458 162374 274694
rect 161754 237814 162374 274458
rect 161754 237578 161786 237814
rect 162022 237578 162106 237814
rect 162342 237578 162374 237814
rect 161754 237494 162374 237578
rect 161754 237258 161786 237494
rect 162022 237258 162106 237494
rect 162342 237258 162374 237494
rect 161754 200614 162374 237258
rect 161754 200378 161786 200614
rect 162022 200378 162106 200614
rect 162342 200378 162374 200614
rect 161754 200294 162374 200378
rect 161754 200058 161786 200294
rect 162022 200058 162106 200294
rect 162342 200058 162374 200294
rect 161754 163414 162374 200058
rect 161754 163178 161786 163414
rect 162022 163178 162106 163414
rect 162342 163178 162374 163414
rect 161754 163094 162374 163178
rect 161754 162858 161786 163094
rect 162022 162858 162106 163094
rect 162342 162858 162374 163094
rect 161754 126214 162374 162858
rect 161754 125978 161786 126214
rect 162022 125978 162106 126214
rect 162342 125978 162374 126214
rect 161754 125894 162374 125978
rect 161754 125658 161786 125894
rect 162022 125658 162106 125894
rect 162342 125658 162374 125894
rect 161754 89014 162374 125658
rect 161754 88778 161786 89014
rect 162022 88778 162106 89014
rect 162342 88778 162374 89014
rect 161754 88694 162374 88778
rect 161754 88458 161786 88694
rect 162022 88458 162106 88694
rect 162342 88458 162374 88694
rect 161754 51814 162374 88458
rect 161754 51578 161786 51814
rect 162022 51578 162106 51814
rect 162342 51578 162374 51814
rect 161754 51494 162374 51578
rect 161754 51258 161786 51494
rect 162022 51258 162106 51494
rect 162342 51258 162374 51494
rect 161754 14614 162374 51258
rect 161754 14378 161786 14614
rect 162022 14378 162106 14614
rect 162342 14378 162374 14614
rect 161754 14294 162374 14378
rect 161754 14058 161786 14294
rect 162022 14058 162106 14294
rect 162342 14058 162374 14294
rect 161754 2176 162374 14058
rect 165474 687934 166094 701760
rect 165474 687698 165506 687934
rect 165742 687698 165826 687934
rect 166062 687698 166094 687934
rect 165474 687614 166094 687698
rect 165474 687378 165506 687614
rect 165742 687378 165826 687614
rect 166062 687378 166094 687614
rect 165474 650734 166094 687378
rect 165474 650498 165506 650734
rect 165742 650498 165826 650734
rect 166062 650498 166094 650734
rect 165474 650414 166094 650498
rect 165474 650178 165506 650414
rect 165742 650178 165826 650414
rect 166062 650178 166094 650414
rect 165474 613534 166094 650178
rect 165474 613298 165506 613534
rect 165742 613298 165826 613534
rect 166062 613298 166094 613534
rect 165474 613214 166094 613298
rect 165474 612978 165506 613214
rect 165742 612978 165826 613214
rect 166062 612978 166094 613214
rect 165474 576334 166094 612978
rect 165474 576098 165506 576334
rect 165742 576098 165826 576334
rect 166062 576098 166094 576334
rect 165474 576014 166094 576098
rect 165474 575778 165506 576014
rect 165742 575778 165826 576014
rect 166062 575778 166094 576014
rect 165474 539134 166094 575778
rect 165474 538898 165506 539134
rect 165742 538898 165826 539134
rect 166062 538898 166094 539134
rect 165474 538814 166094 538898
rect 165474 538578 165506 538814
rect 165742 538578 165826 538814
rect 166062 538578 166094 538814
rect 165474 501934 166094 538578
rect 165474 501698 165506 501934
rect 165742 501698 165826 501934
rect 166062 501698 166094 501934
rect 165474 501614 166094 501698
rect 165474 501378 165506 501614
rect 165742 501378 165826 501614
rect 166062 501378 166094 501614
rect 165474 464734 166094 501378
rect 165474 464498 165506 464734
rect 165742 464498 165826 464734
rect 166062 464498 166094 464734
rect 165474 464414 166094 464498
rect 165474 464178 165506 464414
rect 165742 464178 165826 464414
rect 166062 464178 166094 464414
rect 165474 427534 166094 464178
rect 165474 427298 165506 427534
rect 165742 427298 165826 427534
rect 166062 427298 166094 427534
rect 165474 427214 166094 427298
rect 165474 426978 165506 427214
rect 165742 426978 165826 427214
rect 166062 426978 166094 427214
rect 165474 390334 166094 426978
rect 165474 390098 165506 390334
rect 165742 390098 165826 390334
rect 166062 390098 166094 390334
rect 165474 390014 166094 390098
rect 165474 389778 165506 390014
rect 165742 389778 165826 390014
rect 166062 389778 166094 390014
rect 165474 353134 166094 389778
rect 165474 352898 165506 353134
rect 165742 352898 165826 353134
rect 166062 352898 166094 353134
rect 165474 352814 166094 352898
rect 165474 352578 165506 352814
rect 165742 352578 165826 352814
rect 166062 352578 166094 352814
rect 165474 315934 166094 352578
rect 165474 315698 165506 315934
rect 165742 315698 165826 315934
rect 166062 315698 166094 315934
rect 165474 315614 166094 315698
rect 165474 315378 165506 315614
rect 165742 315378 165826 315614
rect 166062 315378 166094 315614
rect 165474 278734 166094 315378
rect 165474 278498 165506 278734
rect 165742 278498 165826 278734
rect 166062 278498 166094 278734
rect 165474 278414 166094 278498
rect 165474 278178 165506 278414
rect 165742 278178 165826 278414
rect 166062 278178 166094 278414
rect 165474 241534 166094 278178
rect 165474 241298 165506 241534
rect 165742 241298 165826 241534
rect 166062 241298 166094 241534
rect 165474 241214 166094 241298
rect 165474 240978 165506 241214
rect 165742 240978 165826 241214
rect 166062 240978 166094 241214
rect 165474 204334 166094 240978
rect 165474 204098 165506 204334
rect 165742 204098 165826 204334
rect 166062 204098 166094 204334
rect 165474 204014 166094 204098
rect 165474 203778 165506 204014
rect 165742 203778 165826 204014
rect 166062 203778 166094 204014
rect 165474 167134 166094 203778
rect 165474 166898 165506 167134
rect 165742 166898 165826 167134
rect 166062 166898 166094 167134
rect 165474 166814 166094 166898
rect 165474 166578 165506 166814
rect 165742 166578 165826 166814
rect 166062 166578 166094 166814
rect 165474 129934 166094 166578
rect 165474 129698 165506 129934
rect 165742 129698 165826 129934
rect 166062 129698 166094 129934
rect 165474 129614 166094 129698
rect 165474 129378 165506 129614
rect 165742 129378 165826 129614
rect 166062 129378 166094 129614
rect 165474 92734 166094 129378
rect 165474 92498 165506 92734
rect 165742 92498 165826 92734
rect 166062 92498 166094 92734
rect 165474 92414 166094 92498
rect 165474 92178 165506 92414
rect 165742 92178 165826 92414
rect 166062 92178 166094 92414
rect 165474 55534 166094 92178
rect 165474 55298 165506 55534
rect 165742 55298 165826 55534
rect 166062 55298 166094 55534
rect 165474 55214 166094 55298
rect 165474 54978 165506 55214
rect 165742 54978 165826 55214
rect 166062 54978 166094 55214
rect 165474 18334 166094 54978
rect 165474 18098 165506 18334
rect 165742 18098 165826 18334
rect 166062 18098 166094 18334
rect 165474 18014 166094 18098
rect 165474 17778 165506 18014
rect 165742 17778 165826 18014
rect 166062 17778 166094 18014
rect 165474 2176 166094 17778
rect 169194 691654 169814 701760
rect 169194 691418 169226 691654
rect 169462 691418 169546 691654
rect 169782 691418 169814 691654
rect 169194 691334 169814 691418
rect 169194 691098 169226 691334
rect 169462 691098 169546 691334
rect 169782 691098 169814 691334
rect 169194 654454 169814 691098
rect 169194 654218 169226 654454
rect 169462 654218 169546 654454
rect 169782 654218 169814 654454
rect 169194 654134 169814 654218
rect 169194 653898 169226 654134
rect 169462 653898 169546 654134
rect 169782 653898 169814 654134
rect 169194 617254 169814 653898
rect 169194 617018 169226 617254
rect 169462 617018 169546 617254
rect 169782 617018 169814 617254
rect 169194 616934 169814 617018
rect 169194 616698 169226 616934
rect 169462 616698 169546 616934
rect 169782 616698 169814 616934
rect 169194 580054 169814 616698
rect 169194 579818 169226 580054
rect 169462 579818 169546 580054
rect 169782 579818 169814 580054
rect 169194 579734 169814 579818
rect 169194 579498 169226 579734
rect 169462 579498 169546 579734
rect 169782 579498 169814 579734
rect 169194 542854 169814 579498
rect 169194 542618 169226 542854
rect 169462 542618 169546 542854
rect 169782 542618 169814 542854
rect 169194 542534 169814 542618
rect 169194 542298 169226 542534
rect 169462 542298 169546 542534
rect 169782 542298 169814 542534
rect 169194 505654 169814 542298
rect 169194 505418 169226 505654
rect 169462 505418 169546 505654
rect 169782 505418 169814 505654
rect 169194 505334 169814 505418
rect 169194 505098 169226 505334
rect 169462 505098 169546 505334
rect 169782 505098 169814 505334
rect 169194 468454 169814 505098
rect 169194 468218 169226 468454
rect 169462 468218 169546 468454
rect 169782 468218 169814 468454
rect 169194 468134 169814 468218
rect 169194 467898 169226 468134
rect 169462 467898 169546 468134
rect 169782 467898 169814 468134
rect 169194 431254 169814 467898
rect 169194 431018 169226 431254
rect 169462 431018 169546 431254
rect 169782 431018 169814 431254
rect 169194 430934 169814 431018
rect 169194 430698 169226 430934
rect 169462 430698 169546 430934
rect 169782 430698 169814 430934
rect 169194 394054 169814 430698
rect 169194 393818 169226 394054
rect 169462 393818 169546 394054
rect 169782 393818 169814 394054
rect 169194 393734 169814 393818
rect 169194 393498 169226 393734
rect 169462 393498 169546 393734
rect 169782 393498 169814 393734
rect 169194 356854 169814 393498
rect 169194 356618 169226 356854
rect 169462 356618 169546 356854
rect 169782 356618 169814 356854
rect 169194 356534 169814 356618
rect 169194 356298 169226 356534
rect 169462 356298 169546 356534
rect 169782 356298 169814 356534
rect 169194 319654 169814 356298
rect 169194 319418 169226 319654
rect 169462 319418 169546 319654
rect 169782 319418 169814 319654
rect 169194 319334 169814 319418
rect 169194 319098 169226 319334
rect 169462 319098 169546 319334
rect 169782 319098 169814 319334
rect 169194 282454 169814 319098
rect 169194 282218 169226 282454
rect 169462 282218 169546 282454
rect 169782 282218 169814 282454
rect 169194 282134 169814 282218
rect 169194 281898 169226 282134
rect 169462 281898 169546 282134
rect 169782 281898 169814 282134
rect 169194 245254 169814 281898
rect 169194 245018 169226 245254
rect 169462 245018 169546 245254
rect 169782 245018 169814 245254
rect 169194 244934 169814 245018
rect 169194 244698 169226 244934
rect 169462 244698 169546 244934
rect 169782 244698 169814 244934
rect 169194 208054 169814 244698
rect 169194 207818 169226 208054
rect 169462 207818 169546 208054
rect 169782 207818 169814 208054
rect 169194 207734 169814 207818
rect 169194 207498 169226 207734
rect 169462 207498 169546 207734
rect 169782 207498 169814 207734
rect 169194 170854 169814 207498
rect 169194 170618 169226 170854
rect 169462 170618 169546 170854
rect 169782 170618 169814 170854
rect 169194 170534 169814 170618
rect 169194 170298 169226 170534
rect 169462 170298 169546 170534
rect 169782 170298 169814 170534
rect 169194 133654 169814 170298
rect 169194 133418 169226 133654
rect 169462 133418 169546 133654
rect 169782 133418 169814 133654
rect 169194 133334 169814 133418
rect 169194 133098 169226 133334
rect 169462 133098 169546 133334
rect 169782 133098 169814 133334
rect 169194 96454 169814 133098
rect 169194 96218 169226 96454
rect 169462 96218 169546 96454
rect 169782 96218 169814 96454
rect 169194 96134 169814 96218
rect 169194 95898 169226 96134
rect 169462 95898 169546 96134
rect 169782 95898 169814 96134
rect 169194 59254 169814 95898
rect 169194 59018 169226 59254
rect 169462 59018 169546 59254
rect 169782 59018 169814 59254
rect 169194 58934 169814 59018
rect 169194 58698 169226 58934
rect 169462 58698 169546 58934
rect 169782 58698 169814 58934
rect 169194 22054 169814 58698
rect 169194 21818 169226 22054
rect 169462 21818 169546 22054
rect 169782 21818 169814 22054
rect 169194 21734 169814 21818
rect 169194 21498 169226 21734
rect 169462 21498 169546 21734
rect 169782 21498 169814 21734
rect 169194 2176 169814 21498
rect 172914 695374 173534 701760
rect 172914 695138 172946 695374
rect 173182 695138 173266 695374
rect 173502 695138 173534 695374
rect 172914 695054 173534 695138
rect 172914 694818 172946 695054
rect 173182 694818 173266 695054
rect 173502 694818 173534 695054
rect 172914 658174 173534 694818
rect 172914 657938 172946 658174
rect 173182 657938 173266 658174
rect 173502 657938 173534 658174
rect 172914 657854 173534 657938
rect 172914 657618 172946 657854
rect 173182 657618 173266 657854
rect 173502 657618 173534 657854
rect 172914 620974 173534 657618
rect 172914 620738 172946 620974
rect 173182 620738 173266 620974
rect 173502 620738 173534 620974
rect 172914 620654 173534 620738
rect 172914 620418 172946 620654
rect 173182 620418 173266 620654
rect 173502 620418 173534 620654
rect 172914 583774 173534 620418
rect 172914 583538 172946 583774
rect 173182 583538 173266 583774
rect 173502 583538 173534 583774
rect 172914 583454 173534 583538
rect 172914 583218 172946 583454
rect 173182 583218 173266 583454
rect 173502 583218 173534 583454
rect 172914 546574 173534 583218
rect 172914 546338 172946 546574
rect 173182 546338 173266 546574
rect 173502 546338 173534 546574
rect 172914 546254 173534 546338
rect 172914 546018 172946 546254
rect 173182 546018 173266 546254
rect 173502 546018 173534 546254
rect 172914 509374 173534 546018
rect 172914 509138 172946 509374
rect 173182 509138 173266 509374
rect 173502 509138 173534 509374
rect 172914 509054 173534 509138
rect 172914 508818 172946 509054
rect 173182 508818 173266 509054
rect 173502 508818 173534 509054
rect 172914 472174 173534 508818
rect 172914 471938 172946 472174
rect 173182 471938 173266 472174
rect 173502 471938 173534 472174
rect 172914 471854 173534 471938
rect 172914 471618 172946 471854
rect 173182 471618 173266 471854
rect 173502 471618 173534 471854
rect 172914 434974 173534 471618
rect 172914 434738 172946 434974
rect 173182 434738 173266 434974
rect 173502 434738 173534 434974
rect 172914 434654 173534 434738
rect 172914 434418 172946 434654
rect 173182 434418 173266 434654
rect 173502 434418 173534 434654
rect 172914 397774 173534 434418
rect 172914 397538 172946 397774
rect 173182 397538 173266 397774
rect 173502 397538 173534 397774
rect 172914 397454 173534 397538
rect 172914 397218 172946 397454
rect 173182 397218 173266 397454
rect 173502 397218 173534 397454
rect 172914 360574 173534 397218
rect 172914 360338 172946 360574
rect 173182 360338 173266 360574
rect 173502 360338 173534 360574
rect 172914 360254 173534 360338
rect 172914 360018 172946 360254
rect 173182 360018 173266 360254
rect 173502 360018 173534 360254
rect 172914 323374 173534 360018
rect 172914 323138 172946 323374
rect 173182 323138 173266 323374
rect 173502 323138 173534 323374
rect 172914 323054 173534 323138
rect 172914 322818 172946 323054
rect 173182 322818 173266 323054
rect 173502 322818 173534 323054
rect 172914 286174 173534 322818
rect 172914 285938 172946 286174
rect 173182 285938 173266 286174
rect 173502 285938 173534 286174
rect 172914 285854 173534 285938
rect 172914 285618 172946 285854
rect 173182 285618 173266 285854
rect 173502 285618 173534 285854
rect 172914 248974 173534 285618
rect 172914 248738 172946 248974
rect 173182 248738 173266 248974
rect 173502 248738 173534 248974
rect 172914 248654 173534 248738
rect 172914 248418 172946 248654
rect 173182 248418 173266 248654
rect 173502 248418 173534 248654
rect 172914 211774 173534 248418
rect 172914 211538 172946 211774
rect 173182 211538 173266 211774
rect 173502 211538 173534 211774
rect 172914 211454 173534 211538
rect 172914 211218 172946 211454
rect 173182 211218 173266 211454
rect 173502 211218 173534 211454
rect 172914 174574 173534 211218
rect 172914 174338 172946 174574
rect 173182 174338 173266 174574
rect 173502 174338 173534 174574
rect 172914 174254 173534 174338
rect 172914 174018 172946 174254
rect 173182 174018 173266 174254
rect 173502 174018 173534 174254
rect 172914 137374 173534 174018
rect 172914 137138 172946 137374
rect 173182 137138 173266 137374
rect 173502 137138 173534 137374
rect 172914 137054 173534 137138
rect 172914 136818 172946 137054
rect 173182 136818 173266 137054
rect 173502 136818 173534 137054
rect 172914 100174 173534 136818
rect 172914 99938 172946 100174
rect 173182 99938 173266 100174
rect 173502 99938 173534 100174
rect 172914 99854 173534 99938
rect 172914 99618 172946 99854
rect 173182 99618 173266 99854
rect 173502 99618 173534 99854
rect 172914 62974 173534 99618
rect 172914 62738 172946 62974
rect 173182 62738 173266 62974
rect 173502 62738 173534 62974
rect 172914 62654 173534 62738
rect 172914 62418 172946 62654
rect 173182 62418 173266 62654
rect 173502 62418 173534 62654
rect 172914 25774 173534 62418
rect 172914 25538 172946 25774
rect 173182 25538 173266 25774
rect 173502 25538 173534 25774
rect 172914 25454 173534 25538
rect 172914 25218 172946 25454
rect 173182 25218 173266 25454
rect 173502 25218 173534 25454
rect 172914 2176 173534 25218
rect 176634 699094 177254 701760
rect 176634 698858 176666 699094
rect 176902 698858 176986 699094
rect 177222 698858 177254 699094
rect 176634 698774 177254 698858
rect 176634 698538 176666 698774
rect 176902 698538 176986 698774
rect 177222 698538 177254 698774
rect 176634 661894 177254 698538
rect 176634 661658 176666 661894
rect 176902 661658 176986 661894
rect 177222 661658 177254 661894
rect 176634 661574 177254 661658
rect 176634 661338 176666 661574
rect 176902 661338 176986 661574
rect 177222 661338 177254 661574
rect 176634 624694 177254 661338
rect 176634 624458 176666 624694
rect 176902 624458 176986 624694
rect 177222 624458 177254 624694
rect 176634 624374 177254 624458
rect 176634 624138 176666 624374
rect 176902 624138 176986 624374
rect 177222 624138 177254 624374
rect 176634 587494 177254 624138
rect 176634 587258 176666 587494
rect 176902 587258 176986 587494
rect 177222 587258 177254 587494
rect 176634 587174 177254 587258
rect 176634 586938 176666 587174
rect 176902 586938 176986 587174
rect 177222 586938 177254 587174
rect 176634 550294 177254 586938
rect 176634 550058 176666 550294
rect 176902 550058 176986 550294
rect 177222 550058 177254 550294
rect 176634 549974 177254 550058
rect 176634 549738 176666 549974
rect 176902 549738 176986 549974
rect 177222 549738 177254 549974
rect 176634 513094 177254 549738
rect 176634 512858 176666 513094
rect 176902 512858 176986 513094
rect 177222 512858 177254 513094
rect 176634 512774 177254 512858
rect 176634 512538 176666 512774
rect 176902 512538 176986 512774
rect 177222 512538 177254 512774
rect 176634 475894 177254 512538
rect 176634 475658 176666 475894
rect 176902 475658 176986 475894
rect 177222 475658 177254 475894
rect 176634 475574 177254 475658
rect 176634 475338 176666 475574
rect 176902 475338 176986 475574
rect 177222 475338 177254 475574
rect 176634 438694 177254 475338
rect 176634 438458 176666 438694
rect 176902 438458 176986 438694
rect 177222 438458 177254 438694
rect 176634 438374 177254 438458
rect 176634 438138 176666 438374
rect 176902 438138 176986 438374
rect 177222 438138 177254 438374
rect 176634 401494 177254 438138
rect 176634 401258 176666 401494
rect 176902 401258 176986 401494
rect 177222 401258 177254 401494
rect 176634 401174 177254 401258
rect 176634 400938 176666 401174
rect 176902 400938 176986 401174
rect 177222 400938 177254 401174
rect 176634 364294 177254 400938
rect 176634 364058 176666 364294
rect 176902 364058 176986 364294
rect 177222 364058 177254 364294
rect 176634 363974 177254 364058
rect 176634 363738 176666 363974
rect 176902 363738 176986 363974
rect 177222 363738 177254 363974
rect 176634 327094 177254 363738
rect 176634 326858 176666 327094
rect 176902 326858 176986 327094
rect 177222 326858 177254 327094
rect 176634 326774 177254 326858
rect 176634 326538 176666 326774
rect 176902 326538 176986 326774
rect 177222 326538 177254 326774
rect 176634 289894 177254 326538
rect 176634 289658 176666 289894
rect 176902 289658 176986 289894
rect 177222 289658 177254 289894
rect 176634 289574 177254 289658
rect 176634 289338 176666 289574
rect 176902 289338 176986 289574
rect 177222 289338 177254 289574
rect 176634 252694 177254 289338
rect 176634 252458 176666 252694
rect 176902 252458 176986 252694
rect 177222 252458 177254 252694
rect 176634 252374 177254 252458
rect 176634 252138 176666 252374
rect 176902 252138 176986 252374
rect 177222 252138 177254 252374
rect 176634 215494 177254 252138
rect 176634 215258 176666 215494
rect 176902 215258 176986 215494
rect 177222 215258 177254 215494
rect 176634 215174 177254 215258
rect 176634 214938 176666 215174
rect 176902 214938 176986 215174
rect 177222 214938 177254 215174
rect 176634 178294 177254 214938
rect 176634 178058 176666 178294
rect 176902 178058 176986 178294
rect 177222 178058 177254 178294
rect 176634 177974 177254 178058
rect 176634 177738 176666 177974
rect 176902 177738 176986 177974
rect 177222 177738 177254 177974
rect 176634 141094 177254 177738
rect 176634 140858 176666 141094
rect 176902 140858 176986 141094
rect 177222 140858 177254 141094
rect 176634 140774 177254 140858
rect 176634 140538 176666 140774
rect 176902 140538 176986 140774
rect 177222 140538 177254 140774
rect 176634 103894 177254 140538
rect 176634 103658 176666 103894
rect 176902 103658 176986 103894
rect 177222 103658 177254 103894
rect 176634 103574 177254 103658
rect 176634 103338 176666 103574
rect 176902 103338 176986 103574
rect 177222 103338 177254 103574
rect 176634 66694 177254 103338
rect 176634 66458 176666 66694
rect 176902 66458 176986 66694
rect 177222 66458 177254 66694
rect 176634 66374 177254 66458
rect 176634 66138 176666 66374
rect 176902 66138 176986 66374
rect 177222 66138 177254 66374
rect 176634 29494 177254 66138
rect 176634 29258 176666 29494
rect 176902 29258 176986 29494
rect 177222 29258 177254 29494
rect 176634 29174 177254 29258
rect 176634 28938 176666 29174
rect 176902 28938 176986 29174
rect 177222 28938 177254 29174
rect 176634 2176 177254 28938
rect 187794 673054 188414 701760
rect 187794 672818 187826 673054
rect 188062 672818 188146 673054
rect 188382 672818 188414 673054
rect 187794 672734 188414 672818
rect 187794 672498 187826 672734
rect 188062 672498 188146 672734
rect 188382 672498 188414 672734
rect 187794 635854 188414 672498
rect 187794 635618 187826 635854
rect 188062 635618 188146 635854
rect 188382 635618 188414 635854
rect 187794 635534 188414 635618
rect 187794 635298 187826 635534
rect 188062 635298 188146 635534
rect 188382 635298 188414 635534
rect 187794 598654 188414 635298
rect 187794 598418 187826 598654
rect 188062 598418 188146 598654
rect 188382 598418 188414 598654
rect 187794 598334 188414 598418
rect 187794 598098 187826 598334
rect 188062 598098 188146 598334
rect 188382 598098 188414 598334
rect 187794 561454 188414 598098
rect 187794 561218 187826 561454
rect 188062 561218 188146 561454
rect 188382 561218 188414 561454
rect 187794 561134 188414 561218
rect 187794 560898 187826 561134
rect 188062 560898 188146 561134
rect 188382 560898 188414 561134
rect 187794 524254 188414 560898
rect 187794 524018 187826 524254
rect 188062 524018 188146 524254
rect 188382 524018 188414 524254
rect 187794 523934 188414 524018
rect 187794 523698 187826 523934
rect 188062 523698 188146 523934
rect 188382 523698 188414 523934
rect 187794 487054 188414 523698
rect 187794 486818 187826 487054
rect 188062 486818 188146 487054
rect 188382 486818 188414 487054
rect 187794 486734 188414 486818
rect 187794 486498 187826 486734
rect 188062 486498 188146 486734
rect 188382 486498 188414 486734
rect 187794 449854 188414 486498
rect 187794 449618 187826 449854
rect 188062 449618 188146 449854
rect 188382 449618 188414 449854
rect 187794 449534 188414 449618
rect 187794 449298 187826 449534
rect 188062 449298 188146 449534
rect 188382 449298 188414 449534
rect 187794 412654 188414 449298
rect 187794 412418 187826 412654
rect 188062 412418 188146 412654
rect 188382 412418 188414 412654
rect 187794 412334 188414 412418
rect 187794 412098 187826 412334
rect 188062 412098 188146 412334
rect 188382 412098 188414 412334
rect 187794 375454 188414 412098
rect 187794 375218 187826 375454
rect 188062 375218 188146 375454
rect 188382 375218 188414 375454
rect 187794 375134 188414 375218
rect 187794 374898 187826 375134
rect 188062 374898 188146 375134
rect 188382 374898 188414 375134
rect 187794 338254 188414 374898
rect 187794 338018 187826 338254
rect 188062 338018 188146 338254
rect 188382 338018 188414 338254
rect 187794 337934 188414 338018
rect 187794 337698 187826 337934
rect 188062 337698 188146 337934
rect 188382 337698 188414 337934
rect 187794 301054 188414 337698
rect 187794 300818 187826 301054
rect 188062 300818 188146 301054
rect 188382 300818 188414 301054
rect 187794 300734 188414 300818
rect 187794 300498 187826 300734
rect 188062 300498 188146 300734
rect 188382 300498 188414 300734
rect 187794 263854 188414 300498
rect 187794 263618 187826 263854
rect 188062 263618 188146 263854
rect 188382 263618 188414 263854
rect 187794 263534 188414 263618
rect 187794 263298 187826 263534
rect 188062 263298 188146 263534
rect 188382 263298 188414 263534
rect 187794 226654 188414 263298
rect 187794 226418 187826 226654
rect 188062 226418 188146 226654
rect 188382 226418 188414 226654
rect 187794 226334 188414 226418
rect 187794 226098 187826 226334
rect 188062 226098 188146 226334
rect 188382 226098 188414 226334
rect 187794 189454 188414 226098
rect 187794 189218 187826 189454
rect 188062 189218 188146 189454
rect 188382 189218 188414 189454
rect 187794 189134 188414 189218
rect 187794 188898 187826 189134
rect 188062 188898 188146 189134
rect 188382 188898 188414 189134
rect 187794 152254 188414 188898
rect 187794 152018 187826 152254
rect 188062 152018 188146 152254
rect 188382 152018 188414 152254
rect 187794 151934 188414 152018
rect 187794 151698 187826 151934
rect 188062 151698 188146 151934
rect 188382 151698 188414 151934
rect 187794 115054 188414 151698
rect 187794 114818 187826 115054
rect 188062 114818 188146 115054
rect 188382 114818 188414 115054
rect 187794 114734 188414 114818
rect 187794 114498 187826 114734
rect 188062 114498 188146 114734
rect 188382 114498 188414 114734
rect 187794 77854 188414 114498
rect 187794 77618 187826 77854
rect 188062 77618 188146 77854
rect 188382 77618 188414 77854
rect 187794 77534 188414 77618
rect 187794 77298 187826 77534
rect 188062 77298 188146 77534
rect 188382 77298 188414 77534
rect 187794 40654 188414 77298
rect 187794 40418 187826 40654
rect 188062 40418 188146 40654
rect 188382 40418 188414 40654
rect 187794 40334 188414 40418
rect 187794 40098 187826 40334
rect 188062 40098 188146 40334
rect 188382 40098 188414 40334
rect 187794 3454 188414 40098
rect 187794 3218 187826 3454
rect 188062 3218 188146 3454
rect 188382 3218 188414 3454
rect 187794 3134 188414 3218
rect 187794 2898 187826 3134
rect 188062 2898 188146 3134
rect 188382 2898 188414 3134
rect 187794 2176 188414 2898
rect 191514 676774 192134 701760
rect 191514 676538 191546 676774
rect 191782 676538 191866 676774
rect 192102 676538 192134 676774
rect 191514 676454 192134 676538
rect 191514 676218 191546 676454
rect 191782 676218 191866 676454
rect 192102 676218 192134 676454
rect 191514 639574 192134 676218
rect 191514 639338 191546 639574
rect 191782 639338 191866 639574
rect 192102 639338 192134 639574
rect 191514 639254 192134 639338
rect 191514 639018 191546 639254
rect 191782 639018 191866 639254
rect 192102 639018 192134 639254
rect 191514 602374 192134 639018
rect 191514 602138 191546 602374
rect 191782 602138 191866 602374
rect 192102 602138 192134 602374
rect 191514 602054 192134 602138
rect 191514 601818 191546 602054
rect 191782 601818 191866 602054
rect 192102 601818 192134 602054
rect 191514 565174 192134 601818
rect 191514 564938 191546 565174
rect 191782 564938 191866 565174
rect 192102 564938 192134 565174
rect 191514 564854 192134 564938
rect 191514 564618 191546 564854
rect 191782 564618 191866 564854
rect 192102 564618 192134 564854
rect 191514 527974 192134 564618
rect 191514 527738 191546 527974
rect 191782 527738 191866 527974
rect 192102 527738 192134 527974
rect 191514 527654 192134 527738
rect 191514 527418 191546 527654
rect 191782 527418 191866 527654
rect 192102 527418 192134 527654
rect 191514 490774 192134 527418
rect 191514 490538 191546 490774
rect 191782 490538 191866 490774
rect 192102 490538 192134 490774
rect 191514 490454 192134 490538
rect 191514 490218 191546 490454
rect 191782 490218 191866 490454
rect 192102 490218 192134 490454
rect 191514 453574 192134 490218
rect 191514 453338 191546 453574
rect 191782 453338 191866 453574
rect 192102 453338 192134 453574
rect 191514 453254 192134 453338
rect 191514 453018 191546 453254
rect 191782 453018 191866 453254
rect 192102 453018 192134 453254
rect 191514 416374 192134 453018
rect 191514 416138 191546 416374
rect 191782 416138 191866 416374
rect 192102 416138 192134 416374
rect 191514 416054 192134 416138
rect 191514 415818 191546 416054
rect 191782 415818 191866 416054
rect 192102 415818 192134 416054
rect 191514 379174 192134 415818
rect 191514 378938 191546 379174
rect 191782 378938 191866 379174
rect 192102 378938 192134 379174
rect 191514 378854 192134 378938
rect 191514 378618 191546 378854
rect 191782 378618 191866 378854
rect 192102 378618 192134 378854
rect 191514 341974 192134 378618
rect 191514 341738 191546 341974
rect 191782 341738 191866 341974
rect 192102 341738 192134 341974
rect 191514 341654 192134 341738
rect 191514 341418 191546 341654
rect 191782 341418 191866 341654
rect 192102 341418 192134 341654
rect 191514 304774 192134 341418
rect 191514 304538 191546 304774
rect 191782 304538 191866 304774
rect 192102 304538 192134 304774
rect 191514 304454 192134 304538
rect 191514 304218 191546 304454
rect 191782 304218 191866 304454
rect 192102 304218 192134 304454
rect 191514 267574 192134 304218
rect 191514 267338 191546 267574
rect 191782 267338 191866 267574
rect 192102 267338 192134 267574
rect 191514 267254 192134 267338
rect 191514 267018 191546 267254
rect 191782 267018 191866 267254
rect 192102 267018 192134 267254
rect 191514 230374 192134 267018
rect 191514 230138 191546 230374
rect 191782 230138 191866 230374
rect 192102 230138 192134 230374
rect 191514 230054 192134 230138
rect 191514 229818 191546 230054
rect 191782 229818 191866 230054
rect 192102 229818 192134 230054
rect 191514 193174 192134 229818
rect 191514 192938 191546 193174
rect 191782 192938 191866 193174
rect 192102 192938 192134 193174
rect 191514 192854 192134 192938
rect 191514 192618 191546 192854
rect 191782 192618 191866 192854
rect 192102 192618 192134 192854
rect 191514 155974 192134 192618
rect 191514 155738 191546 155974
rect 191782 155738 191866 155974
rect 192102 155738 192134 155974
rect 191514 155654 192134 155738
rect 191514 155418 191546 155654
rect 191782 155418 191866 155654
rect 192102 155418 192134 155654
rect 191514 118774 192134 155418
rect 191514 118538 191546 118774
rect 191782 118538 191866 118774
rect 192102 118538 192134 118774
rect 191514 118454 192134 118538
rect 191514 118218 191546 118454
rect 191782 118218 191866 118454
rect 192102 118218 192134 118454
rect 191514 81574 192134 118218
rect 191514 81338 191546 81574
rect 191782 81338 191866 81574
rect 192102 81338 192134 81574
rect 191514 81254 192134 81338
rect 191514 81018 191546 81254
rect 191782 81018 191866 81254
rect 192102 81018 192134 81254
rect 191514 44374 192134 81018
rect 191514 44138 191546 44374
rect 191782 44138 191866 44374
rect 192102 44138 192134 44374
rect 191514 44054 192134 44138
rect 191514 43818 191546 44054
rect 191782 43818 191866 44054
rect 192102 43818 192134 44054
rect 191514 7174 192134 43818
rect 191514 6938 191546 7174
rect 191782 6938 191866 7174
rect 192102 6938 192134 7174
rect 191514 6854 192134 6938
rect 191514 6618 191546 6854
rect 191782 6618 191866 6854
rect 192102 6618 192134 6854
rect 191514 2176 192134 6618
rect 195234 680494 195854 701760
rect 195234 680258 195266 680494
rect 195502 680258 195586 680494
rect 195822 680258 195854 680494
rect 195234 680174 195854 680258
rect 195234 679938 195266 680174
rect 195502 679938 195586 680174
rect 195822 679938 195854 680174
rect 195234 643294 195854 679938
rect 195234 643058 195266 643294
rect 195502 643058 195586 643294
rect 195822 643058 195854 643294
rect 195234 642974 195854 643058
rect 195234 642738 195266 642974
rect 195502 642738 195586 642974
rect 195822 642738 195854 642974
rect 195234 606094 195854 642738
rect 195234 605858 195266 606094
rect 195502 605858 195586 606094
rect 195822 605858 195854 606094
rect 195234 605774 195854 605858
rect 195234 605538 195266 605774
rect 195502 605538 195586 605774
rect 195822 605538 195854 605774
rect 195234 568894 195854 605538
rect 195234 568658 195266 568894
rect 195502 568658 195586 568894
rect 195822 568658 195854 568894
rect 195234 568574 195854 568658
rect 195234 568338 195266 568574
rect 195502 568338 195586 568574
rect 195822 568338 195854 568574
rect 195234 531694 195854 568338
rect 195234 531458 195266 531694
rect 195502 531458 195586 531694
rect 195822 531458 195854 531694
rect 195234 531374 195854 531458
rect 195234 531138 195266 531374
rect 195502 531138 195586 531374
rect 195822 531138 195854 531374
rect 195234 494494 195854 531138
rect 195234 494258 195266 494494
rect 195502 494258 195586 494494
rect 195822 494258 195854 494494
rect 195234 494174 195854 494258
rect 195234 493938 195266 494174
rect 195502 493938 195586 494174
rect 195822 493938 195854 494174
rect 195234 457294 195854 493938
rect 195234 457058 195266 457294
rect 195502 457058 195586 457294
rect 195822 457058 195854 457294
rect 195234 456974 195854 457058
rect 195234 456738 195266 456974
rect 195502 456738 195586 456974
rect 195822 456738 195854 456974
rect 195234 420094 195854 456738
rect 195234 419858 195266 420094
rect 195502 419858 195586 420094
rect 195822 419858 195854 420094
rect 195234 419774 195854 419858
rect 195234 419538 195266 419774
rect 195502 419538 195586 419774
rect 195822 419538 195854 419774
rect 195234 382894 195854 419538
rect 195234 382658 195266 382894
rect 195502 382658 195586 382894
rect 195822 382658 195854 382894
rect 195234 382574 195854 382658
rect 195234 382338 195266 382574
rect 195502 382338 195586 382574
rect 195822 382338 195854 382574
rect 195234 345694 195854 382338
rect 195234 345458 195266 345694
rect 195502 345458 195586 345694
rect 195822 345458 195854 345694
rect 195234 345374 195854 345458
rect 195234 345138 195266 345374
rect 195502 345138 195586 345374
rect 195822 345138 195854 345374
rect 195234 308494 195854 345138
rect 195234 308258 195266 308494
rect 195502 308258 195586 308494
rect 195822 308258 195854 308494
rect 195234 308174 195854 308258
rect 195234 307938 195266 308174
rect 195502 307938 195586 308174
rect 195822 307938 195854 308174
rect 195234 271294 195854 307938
rect 195234 271058 195266 271294
rect 195502 271058 195586 271294
rect 195822 271058 195854 271294
rect 195234 270974 195854 271058
rect 195234 270738 195266 270974
rect 195502 270738 195586 270974
rect 195822 270738 195854 270974
rect 195234 234094 195854 270738
rect 195234 233858 195266 234094
rect 195502 233858 195586 234094
rect 195822 233858 195854 234094
rect 195234 233774 195854 233858
rect 195234 233538 195266 233774
rect 195502 233538 195586 233774
rect 195822 233538 195854 233774
rect 195234 196894 195854 233538
rect 195234 196658 195266 196894
rect 195502 196658 195586 196894
rect 195822 196658 195854 196894
rect 195234 196574 195854 196658
rect 195234 196338 195266 196574
rect 195502 196338 195586 196574
rect 195822 196338 195854 196574
rect 195234 159694 195854 196338
rect 195234 159458 195266 159694
rect 195502 159458 195586 159694
rect 195822 159458 195854 159694
rect 195234 159374 195854 159458
rect 195234 159138 195266 159374
rect 195502 159138 195586 159374
rect 195822 159138 195854 159374
rect 195234 122494 195854 159138
rect 195234 122258 195266 122494
rect 195502 122258 195586 122494
rect 195822 122258 195854 122494
rect 195234 122174 195854 122258
rect 195234 121938 195266 122174
rect 195502 121938 195586 122174
rect 195822 121938 195854 122174
rect 195234 85294 195854 121938
rect 195234 85058 195266 85294
rect 195502 85058 195586 85294
rect 195822 85058 195854 85294
rect 195234 84974 195854 85058
rect 195234 84738 195266 84974
rect 195502 84738 195586 84974
rect 195822 84738 195854 84974
rect 195234 48094 195854 84738
rect 195234 47858 195266 48094
rect 195502 47858 195586 48094
rect 195822 47858 195854 48094
rect 195234 47774 195854 47858
rect 195234 47538 195266 47774
rect 195502 47538 195586 47774
rect 195822 47538 195854 47774
rect 195234 10894 195854 47538
rect 195234 10658 195266 10894
rect 195502 10658 195586 10894
rect 195822 10658 195854 10894
rect 195234 10574 195854 10658
rect 195234 10338 195266 10574
rect 195502 10338 195586 10574
rect 195822 10338 195854 10574
rect 195234 2176 195854 10338
rect 198954 684214 199574 701760
rect 198954 683978 198986 684214
rect 199222 683978 199306 684214
rect 199542 683978 199574 684214
rect 198954 683894 199574 683978
rect 198954 683658 198986 683894
rect 199222 683658 199306 683894
rect 199542 683658 199574 683894
rect 198954 647014 199574 683658
rect 198954 646778 198986 647014
rect 199222 646778 199306 647014
rect 199542 646778 199574 647014
rect 198954 646694 199574 646778
rect 198954 646458 198986 646694
rect 199222 646458 199306 646694
rect 199542 646458 199574 646694
rect 198954 609814 199574 646458
rect 198954 609578 198986 609814
rect 199222 609578 199306 609814
rect 199542 609578 199574 609814
rect 198954 609494 199574 609578
rect 198954 609258 198986 609494
rect 199222 609258 199306 609494
rect 199542 609258 199574 609494
rect 198954 572614 199574 609258
rect 198954 572378 198986 572614
rect 199222 572378 199306 572614
rect 199542 572378 199574 572614
rect 198954 572294 199574 572378
rect 198954 572058 198986 572294
rect 199222 572058 199306 572294
rect 199542 572058 199574 572294
rect 198954 535414 199574 572058
rect 198954 535178 198986 535414
rect 199222 535178 199306 535414
rect 199542 535178 199574 535414
rect 198954 535094 199574 535178
rect 198954 534858 198986 535094
rect 199222 534858 199306 535094
rect 199542 534858 199574 535094
rect 198954 498214 199574 534858
rect 198954 497978 198986 498214
rect 199222 497978 199306 498214
rect 199542 497978 199574 498214
rect 198954 497894 199574 497978
rect 198954 497658 198986 497894
rect 199222 497658 199306 497894
rect 199542 497658 199574 497894
rect 198954 461014 199574 497658
rect 198954 460778 198986 461014
rect 199222 460778 199306 461014
rect 199542 460778 199574 461014
rect 198954 460694 199574 460778
rect 198954 460458 198986 460694
rect 199222 460458 199306 460694
rect 199542 460458 199574 460694
rect 198954 423814 199574 460458
rect 198954 423578 198986 423814
rect 199222 423578 199306 423814
rect 199542 423578 199574 423814
rect 198954 423494 199574 423578
rect 198954 423258 198986 423494
rect 199222 423258 199306 423494
rect 199542 423258 199574 423494
rect 198954 386614 199574 423258
rect 198954 386378 198986 386614
rect 199222 386378 199306 386614
rect 199542 386378 199574 386614
rect 198954 386294 199574 386378
rect 198954 386058 198986 386294
rect 199222 386058 199306 386294
rect 199542 386058 199574 386294
rect 198954 349414 199574 386058
rect 198954 349178 198986 349414
rect 199222 349178 199306 349414
rect 199542 349178 199574 349414
rect 198954 349094 199574 349178
rect 198954 348858 198986 349094
rect 199222 348858 199306 349094
rect 199542 348858 199574 349094
rect 198954 312214 199574 348858
rect 198954 311978 198986 312214
rect 199222 311978 199306 312214
rect 199542 311978 199574 312214
rect 198954 311894 199574 311978
rect 198954 311658 198986 311894
rect 199222 311658 199306 311894
rect 199542 311658 199574 311894
rect 198954 275014 199574 311658
rect 198954 274778 198986 275014
rect 199222 274778 199306 275014
rect 199542 274778 199574 275014
rect 198954 274694 199574 274778
rect 198954 274458 198986 274694
rect 199222 274458 199306 274694
rect 199542 274458 199574 274694
rect 198954 237814 199574 274458
rect 198954 237578 198986 237814
rect 199222 237578 199306 237814
rect 199542 237578 199574 237814
rect 198954 237494 199574 237578
rect 198954 237258 198986 237494
rect 199222 237258 199306 237494
rect 199542 237258 199574 237494
rect 198954 200614 199574 237258
rect 198954 200378 198986 200614
rect 199222 200378 199306 200614
rect 199542 200378 199574 200614
rect 198954 200294 199574 200378
rect 198954 200058 198986 200294
rect 199222 200058 199306 200294
rect 199542 200058 199574 200294
rect 198954 163414 199574 200058
rect 198954 163178 198986 163414
rect 199222 163178 199306 163414
rect 199542 163178 199574 163414
rect 198954 163094 199574 163178
rect 198954 162858 198986 163094
rect 199222 162858 199306 163094
rect 199542 162858 199574 163094
rect 198954 126214 199574 162858
rect 198954 125978 198986 126214
rect 199222 125978 199306 126214
rect 199542 125978 199574 126214
rect 198954 125894 199574 125978
rect 198954 125658 198986 125894
rect 199222 125658 199306 125894
rect 199542 125658 199574 125894
rect 198954 89014 199574 125658
rect 198954 88778 198986 89014
rect 199222 88778 199306 89014
rect 199542 88778 199574 89014
rect 198954 88694 199574 88778
rect 198954 88458 198986 88694
rect 199222 88458 199306 88694
rect 199542 88458 199574 88694
rect 198954 51814 199574 88458
rect 198954 51578 198986 51814
rect 199222 51578 199306 51814
rect 199542 51578 199574 51814
rect 198954 51494 199574 51578
rect 198954 51258 198986 51494
rect 199222 51258 199306 51494
rect 199542 51258 199574 51494
rect 198954 14614 199574 51258
rect 198954 14378 198986 14614
rect 199222 14378 199306 14614
rect 199542 14378 199574 14614
rect 198954 14294 199574 14378
rect 198954 14058 198986 14294
rect 199222 14058 199306 14294
rect 199542 14058 199574 14294
rect 198954 2176 199574 14058
rect 202674 687934 203294 701760
rect 202674 687698 202706 687934
rect 202942 687698 203026 687934
rect 203262 687698 203294 687934
rect 202674 687614 203294 687698
rect 202674 687378 202706 687614
rect 202942 687378 203026 687614
rect 203262 687378 203294 687614
rect 202674 650734 203294 687378
rect 202674 650498 202706 650734
rect 202942 650498 203026 650734
rect 203262 650498 203294 650734
rect 202674 650414 203294 650498
rect 202674 650178 202706 650414
rect 202942 650178 203026 650414
rect 203262 650178 203294 650414
rect 202674 613534 203294 650178
rect 202674 613298 202706 613534
rect 202942 613298 203026 613534
rect 203262 613298 203294 613534
rect 202674 613214 203294 613298
rect 202674 612978 202706 613214
rect 202942 612978 203026 613214
rect 203262 612978 203294 613214
rect 202674 576334 203294 612978
rect 202674 576098 202706 576334
rect 202942 576098 203026 576334
rect 203262 576098 203294 576334
rect 202674 576014 203294 576098
rect 202674 575778 202706 576014
rect 202942 575778 203026 576014
rect 203262 575778 203294 576014
rect 202674 539134 203294 575778
rect 202674 538898 202706 539134
rect 202942 538898 203026 539134
rect 203262 538898 203294 539134
rect 202674 538814 203294 538898
rect 202674 538578 202706 538814
rect 202942 538578 203026 538814
rect 203262 538578 203294 538814
rect 202674 501934 203294 538578
rect 202674 501698 202706 501934
rect 202942 501698 203026 501934
rect 203262 501698 203294 501934
rect 202674 501614 203294 501698
rect 202674 501378 202706 501614
rect 202942 501378 203026 501614
rect 203262 501378 203294 501614
rect 202674 464734 203294 501378
rect 202674 464498 202706 464734
rect 202942 464498 203026 464734
rect 203262 464498 203294 464734
rect 202674 464414 203294 464498
rect 202674 464178 202706 464414
rect 202942 464178 203026 464414
rect 203262 464178 203294 464414
rect 202674 427534 203294 464178
rect 202674 427298 202706 427534
rect 202942 427298 203026 427534
rect 203262 427298 203294 427534
rect 202674 427214 203294 427298
rect 202674 426978 202706 427214
rect 202942 426978 203026 427214
rect 203262 426978 203294 427214
rect 202674 390334 203294 426978
rect 202674 390098 202706 390334
rect 202942 390098 203026 390334
rect 203262 390098 203294 390334
rect 202674 390014 203294 390098
rect 202674 389778 202706 390014
rect 202942 389778 203026 390014
rect 203262 389778 203294 390014
rect 202674 353134 203294 389778
rect 202674 352898 202706 353134
rect 202942 352898 203026 353134
rect 203262 352898 203294 353134
rect 202674 352814 203294 352898
rect 202674 352578 202706 352814
rect 202942 352578 203026 352814
rect 203262 352578 203294 352814
rect 202674 315934 203294 352578
rect 202674 315698 202706 315934
rect 202942 315698 203026 315934
rect 203262 315698 203294 315934
rect 202674 315614 203294 315698
rect 202674 315378 202706 315614
rect 202942 315378 203026 315614
rect 203262 315378 203294 315614
rect 202674 278734 203294 315378
rect 202674 278498 202706 278734
rect 202942 278498 203026 278734
rect 203262 278498 203294 278734
rect 202674 278414 203294 278498
rect 202674 278178 202706 278414
rect 202942 278178 203026 278414
rect 203262 278178 203294 278414
rect 202674 241534 203294 278178
rect 202674 241298 202706 241534
rect 202942 241298 203026 241534
rect 203262 241298 203294 241534
rect 202674 241214 203294 241298
rect 202674 240978 202706 241214
rect 202942 240978 203026 241214
rect 203262 240978 203294 241214
rect 202674 204334 203294 240978
rect 202674 204098 202706 204334
rect 202942 204098 203026 204334
rect 203262 204098 203294 204334
rect 202674 204014 203294 204098
rect 202674 203778 202706 204014
rect 202942 203778 203026 204014
rect 203262 203778 203294 204014
rect 202674 167134 203294 203778
rect 202674 166898 202706 167134
rect 202942 166898 203026 167134
rect 203262 166898 203294 167134
rect 202674 166814 203294 166898
rect 202674 166578 202706 166814
rect 202942 166578 203026 166814
rect 203262 166578 203294 166814
rect 202674 129934 203294 166578
rect 202674 129698 202706 129934
rect 202942 129698 203026 129934
rect 203262 129698 203294 129934
rect 202674 129614 203294 129698
rect 202674 129378 202706 129614
rect 202942 129378 203026 129614
rect 203262 129378 203294 129614
rect 202674 92734 203294 129378
rect 202674 92498 202706 92734
rect 202942 92498 203026 92734
rect 203262 92498 203294 92734
rect 202674 92414 203294 92498
rect 202674 92178 202706 92414
rect 202942 92178 203026 92414
rect 203262 92178 203294 92414
rect 202674 55534 203294 92178
rect 202674 55298 202706 55534
rect 202942 55298 203026 55534
rect 203262 55298 203294 55534
rect 202674 55214 203294 55298
rect 202674 54978 202706 55214
rect 202942 54978 203026 55214
rect 203262 54978 203294 55214
rect 202674 18334 203294 54978
rect 202674 18098 202706 18334
rect 202942 18098 203026 18334
rect 203262 18098 203294 18334
rect 202674 18014 203294 18098
rect 202674 17778 202706 18014
rect 202942 17778 203026 18014
rect 203262 17778 203294 18014
rect 202674 2176 203294 17778
rect 206394 691654 207014 701760
rect 206394 691418 206426 691654
rect 206662 691418 206746 691654
rect 206982 691418 207014 691654
rect 206394 691334 207014 691418
rect 206394 691098 206426 691334
rect 206662 691098 206746 691334
rect 206982 691098 207014 691334
rect 206394 654454 207014 691098
rect 206394 654218 206426 654454
rect 206662 654218 206746 654454
rect 206982 654218 207014 654454
rect 206394 654134 207014 654218
rect 206394 653898 206426 654134
rect 206662 653898 206746 654134
rect 206982 653898 207014 654134
rect 206394 617254 207014 653898
rect 206394 617018 206426 617254
rect 206662 617018 206746 617254
rect 206982 617018 207014 617254
rect 206394 616934 207014 617018
rect 206394 616698 206426 616934
rect 206662 616698 206746 616934
rect 206982 616698 207014 616934
rect 206394 580054 207014 616698
rect 206394 579818 206426 580054
rect 206662 579818 206746 580054
rect 206982 579818 207014 580054
rect 206394 579734 207014 579818
rect 206394 579498 206426 579734
rect 206662 579498 206746 579734
rect 206982 579498 207014 579734
rect 206394 542854 207014 579498
rect 206394 542618 206426 542854
rect 206662 542618 206746 542854
rect 206982 542618 207014 542854
rect 206394 542534 207014 542618
rect 206394 542298 206426 542534
rect 206662 542298 206746 542534
rect 206982 542298 207014 542534
rect 206394 505654 207014 542298
rect 206394 505418 206426 505654
rect 206662 505418 206746 505654
rect 206982 505418 207014 505654
rect 206394 505334 207014 505418
rect 206394 505098 206426 505334
rect 206662 505098 206746 505334
rect 206982 505098 207014 505334
rect 206394 468454 207014 505098
rect 206394 468218 206426 468454
rect 206662 468218 206746 468454
rect 206982 468218 207014 468454
rect 206394 468134 207014 468218
rect 206394 467898 206426 468134
rect 206662 467898 206746 468134
rect 206982 467898 207014 468134
rect 206394 431254 207014 467898
rect 206394 431018 206426 431254
rect 206662 431018 206746 431254
rect 206982 431018 207014 431254
rect 206394 430934 207014 431018
rect 206394 430698 206426 430934
rect 206662 430698 206746 430934
rect 206982 430698 207014 430934
rect 206394 394054 207014 430698
rect 206394 393818 206426 394054
rect 206662 393818 206746 394054
rect 206982 393818 207014 394054
rect 206394 393734 207014 393818
rect 206394 393498 206426 393734
rect 206662 393498 206746 393734
rect 206982 393498 207014 393734
rect 206394 356854 207014 393498
rect 206394 356618 206426 356854
rect 206662 356618 206746 356854
rect 206982 356618 207014 356854
rect 206394 356534 207014 356618
rect 206394 356298 206426 356534
rect 206662 356298 206746 356534
rect 206982 356298 207014 356534
rect 206394 319654 207014 356298
rect 206394 319418 206426 319654
rect 206662 319418 206746 319654
rect 206982 319418 207014 319654
rect 206394 319334 207014 319418
rect 206394 319098 206426 319334
rect 206662 319098 206746 319334
rect 206982 319098 207014 319334
rect 206394 282454 207014 319098
rect 206394 282218 206426 282454
rect 206662 282218 206746 282454
rect 206982 282218 207014 282454
rect 206394 282134 207014 282218
rect 206394 281898 206426 282134
rect 206662 281898 206746 282134
rect 206982 281898 207014 282134
rect 206394 245254 207014 281898
rect 206394 245018 206426 245254
rect 206662 245018 206746 245254
rect 206982 245018 207014 245254
rect 206394 244934 207014 245018
rect 206394 244698 206426 244934
rect 206662 244698 206746 244934
rect 206982 244698 207014 244934
rect 206394 208054 207014 244698
rect 206394 207818 206426 208054
rect 206662 207818 206746 208054
rect 206982 207818 207014 208054
rect 206394 207734 207014 207818
rect 206394 207498 206426 207734
rect 206662 207498 206746 207734
rect 206982 207498 207014 207734
rect 206394 170854 207014 207498
rect 206394 170618 206426 170854
rect 206662 170618 206746 170854
rect 206982 170618 207014 170854
rect 206394 170534 207014 170618
rect 206394 170298 206426 170534
rect 206662 170298 206746 170534
rect 206982 170298 207014 170534
rect 206394 133654 207014 170298
rect 206394 133418 206426 133654
rect 206662 133418 206746 133654
rect 206982 133418 207014 133654
rect 206394 133334 207014 133418
rect 206394 133098 206426 133334
rect 206662 133098 206746 133334
rect 206982 133098 207014 133334
rect 206394 96454 207014 133098
rect 206394 96218 206426 96454
rect 206662 96218 206746 96454
rect 206982 96218 207014 96454
rect 206394 96134 207014 96218
rect 206394 95898 206426 96134
rect 206662 95898 206746 96134
rect 206982 95898 207014 96134
rect 206394 59254 207014 95898
rect 206394 59018 206426 59254
rect 206662 59018 206746 59254
rect 206982 59018 207014 59254
rect 206394 58934 207014 59018
rect 206394 58698 206426 58934
rect 206662 58698 206746 58934
rect 206982 58698 207014 58934
rect 206394 22054 207014 58698
rect 206394 21818 206426 22054
rect 206662 21818 206746 22054
rect 206982 21818 207014 22054
rect 206394 21734 207014 21818
rect 206394 21498 206426 21734
rect 206662 21498 206746 21734
rect 206982 21498 207014 21734
rect 206394 2176 207014 21498
rect 210114 695374 210734 701760
rect 210114 695138 210146 695374
rect 210382 695138 210466 695374
rect 210702 695138 210734 695374
rect 210114 695054 210734 695138
rect 210114 694818 210146 695054
rect 210382 694818 210466 695054
rect 210702 694818 210734 695054
rect 210114 658174 210734 694818
rect 210114 657938 210146 658174
rect 210382 657938 210466 658174
rect 210702 657938 210734 658174
rect 210114 657854 210734 657938
rect 210114 657618 210146 657854
rect 210382 657618 210466 657854
rect 210702 657618 210734 657854
rect 210114 620974 210734 657618
rect 210114 620738 210146 620974
rect 210382 620738 210466 620974
rect 210702 620738 210734 620974
rect 210114 620654 210734 620738
rect 210114 620418 210146 620654
rect 210382 620418 210466 620654
rect 210702 620418 210734 620654
rect 210114 583774 210734 620418
rect 210114 583538 210146 583774
rect 210382 583538 210466 583774
rect 210702 583538 210734 583774
rect 210114 583454 210734 583538
rect 210114 583218 210146 583454
rect 210382 583218 210466 583454
rect 210702 583218 210734 583454
rect 210114 546574 210734 583218
rect 210114 546338 210146 546574
rect 210382 546338 210466 546574
rect 210702 546338 210734 546574
rect 210114 546254 210734 546338
rect 210114 546018 210146 546254
rect 210382 546018 210466 546254
rect 210702 546018 210734 546254
rect 210114 509374 210734 546018
rect 210114 509138 210146 509374
rect 210382 509138 210466 509374
rect 210702 509138 210734 509374
rect 210114 509054 210734 509138
rect 210114 508818 210146 509054
rect 210382 508818 210466 509054
rect 210702 508818 210734 509054
rect 210114 472174 210734 508818
rect 210114 471938 210146 472174
rect 210382 471938 210466 472174
rect 210702 471938 210734 472174
rect 210114 471854 210734 471938
rect 210114 471618 210146 471854
rect 210382 471618 210466 471854
rect 210702 471618 210734 471854
rect 210114 434974 210734 471618
rect 210114 434738 210146 434974
rect 210382 434738 210466 434974
rect 210702 434738 210734 434974
rect 210114 434654 210734 434738
rect 210114 434418 210146 434654
rect 210382 434418 210466 434654
rect 210702 434418 210734 434654
rect 210114 397774 210734 434418
rect 210114 397538 210146 397774
rect 210382 397538 210466 397774
rect 210702 397538 210734 397774
rect 210114 397454 210734 397538
rect 210114 397218 210146 397454
rect 210382 397218 210466 397454
rect 210702 397218 210734 397454
rect 210114 360574 210734 397218
rect 210114 360338 210146 360574
rect 210382 360338 210466 360574
rect 210702 360338 210734 360574
rect 210114 360254 210734 360338
rect 210114 360018 210146 360254
rect 210382 360018 210466 360254
rect 210702 360018 210734 360254
rect 210114 323374 210734 360018
rect 210114 323138 210146 323374
rect 210382 323138 210466 323374
rect 210702 323138 210734 323374
rect 210114 323054 210734 323138
rect 210114 322818 210146 323054
rect 210382 322818 210466 323054
rect 210702 322818 210734 323054
rect 210114 286174 210734 322818
rect 210114 285938 210146 286174
rect 210382 285938 210466 286174
rect 210702 285938 210734 286174
rect 210114 285854 210734 285938
rect 210114 285618 210146 285854
rect 210382 285618 210466 285854
rect 210702 285618 210734 285854
rect 210114 248974 210734 285618
rect 210114 248738 210146 248974
rect 210382 248738 210466 248974
rect 210702 248738 210734 248974
rect 210114 248654 210734 248738
rect 210114 248418 210146 248654
rect 210382 248418 210466 248654
rect 210702 248418 210734 248654
rect 210114 211774 210734 248418
rect 210114 211538 210146 211774
rect 210382 211538 210466 211774
rect 210702 211538 210734 211774
rect 210114 211454 210734 211538
rect 210114 211218 210146 211454
rect 210382 211218 210466 211454
rect 210702 211218 210734 211454
rect 210114 174574 210734 211218
rect 210114 174338 210146 174574
rect 210382 174338 210466 174574
rect 210702 174338 210734 174574
rect 210114 174254 210734 174338
rect 210114 174018 210146 174254
rect 210382 174018 210466 174254
rect 210702 174018 210734 174254
rect 210114 137374 210734 174018
rect 210114 137138 210146 137374
rect 210382 137138 210466 137374
rect 210702 137138 210734 137374
rect 210114 137054 210734 137138
rect 210114 136818 210146 137054
rect 210382 136818 210466 137054
rect 210702 136818 210734 137054
rect 210114 100174 210734 136818
rect 210114 99938 210146 100174
rect 210382 99938 210466 100174
rect 210702 99938 210734 100174
rect 210114 99854 210734 99938
rect 210114 99618 210146 99854
rect 210382 99618 210466 99854
rect 210702 99618 210734 99854
rect 210114 62974 210734 99618
rect 210114 62738 210146 62974
rect 210382 62738 210466 62974
rect 210702 62738 210734 62974
rect 210114 62654 210734 62738
rect 210114 62418 210146 62654
rect 210382 62418 210466 62654
rect 210702 62418 210734 62654
rect 210114 25774 210734 62418
rect 210114 25538 210146 25774
rect 210382 25538 210466 25774
rect 210702 25538 210734 25774
rect 210114 25454 210734 25538
rect 210114 25218 210146 25454
rect 210382 25218 210466 25454
rect 210702 25218 210734 25454
rect 210114 2176 210734 25218
rect 213834 699094 214454 701760
rect 213834 698858 213866 699094
rect 214102 698858 214186 699094
rect 214422 698858 214454 699094
rect 213834 698774 214454 698858
rect 213834 698538 213866 698774
rect 214102 698538 214186 698774
rect 214422 698538 214454 698774
rect 213834 661894 214454 698538
rect 213834 661658 213866 661894
rect 214102 661658 214186 661894
rect 214422 661658 214454 661894
rect 213834 661574 214454 661658
rect 213834 661338 213866 661574
rect 214102 661338 214186 661574
rect 214422 661338 214454 661574
rect 213834 624694 214454 661338
rect 213834 624458 213866 624694
rect 214102 624458 214186 624694
rect 214422 624458 214454 624694
rect 213834 624374 214454 624458
rect 213834 624138 213866 624374
rect 214102 624138 214186 624374
rect 214422 624138 214454 624374
rect 213834 587494 214454 624138
rect 213834 587258 213866 587494
rect 214102 587258 214186 587494
rect 214422 587258 214454 587494
rect 213834 587174 214454 587258
rect 213834 586938 213866 587174
rect 214102 586938 214186 587174
rect 214422 586938 214454 587174
rect 213834 550294 214454 586938
rect 213834 550058 213866 550294
rect 214102 550058 214186 550294
rect 214422 550058 214454 550294
rect 213834 549974 214454 550058
rect 213834 549738 213866 549974
rect 214102 549738 214186 549974
rect 214422 549738 214454 549974
rect 213834 513094 214454 549738
rect 213834 512858 213866 513094
rect 214102 512858 214186 513094
rect 214422 512858 214454 513094
rect 213834 512774 214454 512858
rect 213834 512538 213866 512774
rect 214102 512538 214186 512774
rect 214422 512538 214454 512774
rect 213834 475894 214454 512538
rect 213834 475658 213866 475894
rect 214102 475658 214186 475894
rect 214422 475658 214454 475894
rect 213834 475574 214454 475658
rect 213834 475338 213866 475574
rect 214102 475338 214186 475574
rect 214422 475338 214454 475574
rect 213834 438694 214454 475338
rect 213834 438458 213866 438694
rect 214102 438458 214186 438694
rect 214422 438458 214454 438694
rect 213834 438374 214454 438458
rect 213834 438138 213866 438374
rect 214102 438138 214186 438374
rect 214422 438138 214454 438374
rect 213834 401494 214454 438138
rect 213834 401258 213866 401494
rect 214102 401258 214186 401494
rect 214422 401258 214454 401494
rect 213834 401174 214454 401258
rect 213834 400938 213866 401174
rect 214102 400938 214186 401174
rect 214422 400938 214454 401174
rect 213834 364294 214454 400938
rect 213834 364058 213866 364294
rect 214102 364058 214186 364294
rect 214422 364058 214454 364294
rect 213834 363974 214454 364058
rect 213834 363738 213866 363974
rect 214102 363738 214186 363974
rect 214422 363738 214454 363974
rect 213834 327094 214454 363738
rect 213834 326858 213866 327094
rect 214102 326858 214186 327094
rect 214422 326858 214454 327094
rect 213834 326774 214454 326858
rect 213834 326538 213866 326774
rect 214102 326538 214186 326774
rect 214422 326538 214454 326774
rect 213834 289894 214454 326538
rect 213834 289658 213866 289894
rect 214102 289658 214186 289894
rect 214422 289658 214454 289894
rect 213834 289574 214454 289658
rect 213834 289338 213866 289574
rect 214102 289338 214186 289574
rect 214422 289338 214454 289574
rect 213834 252694 214454 289338
rect 213834 252458 213866 252694
rect 214102 252458 214186 252694
rect 214422 252458 214454 252694
rect 213834 252374 214454 252458
rect 213834 252138 213866 252374
rect 214102 252138 214186 252374
rect 214422 252138 214454 252374
rect 213834 215494 214454 252138
rect 213834 215258 213866 215494
rect 214102 215258 214186 215494
rect 214422 215258 214454 215494
rect 213834 215174 214454 215258
rect 213834 214938 213866 215174
rect 214102 214938 214186 215174
rect 214422 214938 214454 215174
rect 213834 178294 214454 214938
rect 213834 178058 213866 178294
rect 214102 178058 214186 178294
rect 214422 178058 214454 178294
rect 213834 177974 214454 178058
rect 213834 177738 213866 177974
rect 214102 177738 214186 177974
rect 214422 177738 214454 177974
rect 213834 141094 214454 177738
rect 213834 140858 213866 141094
rect 214102 140858 214186 141094
rect 214422 140858 214454 141094
rect 213834 140774 214454 140858
rect 213834 140538 213866 140774
rect 214102 140538 214186 140774
rect 214422 140538 214454 140774
rect 213834 103894 214454 140538
rect 213834 103658 213866 103894
rect 214102 103658 214186 103894
rect 214422 103658 214454 103894
rect 213834 103574 214454 103658
rect 213834 103338 213866 103574
rect 214102 103338 214186 103574
rect 214422 103338 214454 103574
rect 213834 66694 214454 103338
rect 213834 66458 213866 66694
rect 214102 66458 214186 66694
rect 214422 66458 214454 66694
rect 213834 66374 214454 66458
rect 213834 66138 213866 66374
rect 214102 66138 214186 66374
rect 214422 66138 214454 66374
rect 213834 29494 214454 66138
rect 213834 29258 213866 29494
rect 214102 29258 214186 29494
rect 214422 29258 214454 29494
rect 213834 29174 214454 29258
rect 213834 28938 213866 29174
rect 214102 28938 214186 29174
rect 214422 28938 214454 29174
rect 213834 2176 214454 28938
rect 224994 673054 225614 701760
rect 224994 672818 225026 673054
rect 225262 672818 225346 673054
rect 225582 672818 225614 673054
rect 224994 672734 225614 672818
rect 224994 672498 225026 672734
rect 225262 672498 225346 672734
rect 225582 672498 225614 672734
rect 224994 635854 225614 672498
rect 224994 635618 225026 635854
rect 225262 635618 225346 635854
rect 225582 635618 225614 635854
rect 224994 635534 225614 635618
rect 224994 635298 225026 635534
rect 225262 635298 225346 635534
rect 225582 635298 225614 635534
rect 224994 598654 225614 635298
rect 224994 598418 225026 598654
rect 225262 598418 225346 598654
rect 225582 598418 225614 598654
rect 224994 598334 225614 598418
rect 224994 598098 225026 598334
rect 225262 598098 225346 598334
rect 225582 598098 225614 598334
rect 224994 561454 225614 598098
rect 224994 561218 225026 561454
rect 225262 561218 225346 561454
rect 225582 561218 225614 561454
rect 224994 561134 225614 561218
rect 224994 560898 225026 561134
rect 225262 560898 225346 561134
rect 225582 560898 225614 561134
rect 224994 524254 225614 560898
rect 224994 524018 225026 524254
rect 225262 524018 225346 524254
rect 225582 524018 225614 524254
rect 224994 523934 225614 524018
rect 224994 523698 225026 523934
rect 225262 523698 225346 523934
rect 225582 523698 225614 523934
rect 224994 487054 225614 523698
rect 224994 486818 225026 487054
rect 225262 486818 225346 487054
rect 225582 486818 225614 487054
rect 224994 486734 225614 486818
rect 224994 486498 225026 486734
rect 225262 486498 225346 486734
rect 225582 486498 225614 486734
rect 224994 449854 225614 486498
rect 224994 449618 225026 449854
rect 225262 449618 225346 449854
rect 225582 449618 225614 449854
rect 224994 449534 225614 449618
rect 224994 449298 225026 449534
rect 225262 449298 225346 449534
rect 225582 449298 225614 449534
rect 224994 412654 225614 449298
rect 224994 412418 225026 412654
rect 225262 412418 225346 412654
rect 225582 412418 225614 412654
rect 224994 412334 225614 412418
rect 224994 412098 225026 412334
rect 225262 412098 225346 412334
rect 225582 412098 225614 412334
rect 224994 375454 225614 412098
rect 224994 375218 225026 375454
rect 225262 375218 225346 375454
rect 225582 375218 225614 375454
rect 224994 375134 225614 375218
rect 224994 374898 225026 375134
rect 225262 374898 225346 375134
rect 225582 374898 225614 375134
rect 224994 338254 225614 374898
rect 224994 338018 225026 338254
rect 225262 338018 225346 338254
rect 225582 338018 225614 338254
rect 224994 337934 225614 338018
rect 224994 337698 225026 337934
rect 225262 337698 225346 337934
rect 225582 337698 225614 337934
rect 224994 301054 225614 337698
rect 224994 300818 225026 301054
rect 225262 300818 225346 301054
rect 225582 300818 225614 301054
rect 224994 300734 225614 300818
rect 224994 300498 225026 300734
rect 225262 300498 225346 300734
rect 225582 300498 225614 300734
rect 224994 263854 225614 300498
rect 224994 263618 225026 263854
rect 225262 263618 225346 263854
rect 225582 263618 225614 263854
rect 224994 263534 225614 263618
rect 224994 263298 225026 263534
rect 225262 263298 225346 263534
rect 225582 263298 225614 263534
rect 224994 226654 225614 263298
rect 224994 226418 225026 226654
rect 225262 226418 225346 226654
rect 225582 226418 225614 226654
rect 224994 226334 225614 226418
rect 224994 226098 225026 226334
rect 225262 226098 225346 226334
rect 225582 226098 225614 226334
rect 224994 189454 225614 226098
rect 224994 189218 225026 189454
rect 225262 189218 225346 189454
rect 225582 189218 225614 189454
rect 224994 189134 225614 189218
rect 224994 188898 225026 189134
rect 225262 188898 225346 189134
rect 225582 188898 225614 189134
rect 224994 152254 225614 188898
rect 224994 152018 225026 152254
rect 225262 152018 225346 152254
rect 225582 152018 225614 152254
rect 224994 151934 225614 152018
rect 224994 151698 225026 151934
rect 225262 151698 225346 151934
rect 225582 151698 225614 151934
rect 224994 115054 225614 151698
rect 224994 114818 225026 115054
rect 225262 114818 225346 115054
rect 225582 114818 225614 115054
rect 224994 114734 225614 114818
rect 224994 114498 225026 114734
rect 225262 114498 225346 114734
rect 225582 114498 225614 114734
rect 224994 77854 225614 114498
rect 224994 77618 225026 77854
rect 225262 77618 225346 77854
rect 225582 77618 225614 77854
rect 224994 77534 225614 77618
rect 224994 77298 225026 77534
rect 225262 77298 225346 77534
rect 225582 77298 225614 77534
rect 224994 40654 225614 77298
rect 224994 40418 225026 40654
rect 225262 40418 225346 40654
rect 225582 40418 225614 40654
rect 224994 40334 225614 40418
rect 224994 40098 225026 40334
rect 225262 40098 225346 40334
rect 225582 40098 225614 40334
rect 224994 3454 225614 40098
rect 224994 3218 225026 3454
rect 225262 3218 225346 3454
rect 225582 3218 225614 3454
rect 224994 3134 225614 3218
rect 224994 2898 225026 3134
rect 225262 2898 225346 3134
rect 225582 2898 225614 3134
rect 224994 2176 225614 2898
rect 228714 676774 229334 701760
rect 228714 676538 228746 676774
rect 228982 676538 229066 676774
rect 229302 676538 229334 676774
rect 228714 676454 229334 676538
rect 228714 676218 228746 676454
rect 228982 676218 229066 676454
rect 229302 676218 229334 676454
rect 228714 639574 229334 676218
rect 228714 639338 228746 639574
rect 228982 639338 229066 639574
rect 229302 639338 229334 639574
rect 228714 639254 229334 639338
rect 228714 639018 228746 639254
rect 228982 639018 229066 639254
rect 229302 639018 229334 639254
rect 228714 602374 229334 639018
rect 228714 602138 228746 602374
rect 228982 602138 229066 602374
rect 229302 602138 229334 602374
rect 228714 602054 229334 602138
rect 228714 601818 228746 602054
rect 228982 601818 229066 602054
rect 229302 601818 229334 602054
rect 228714 565174 229334 601818
rect 228714 564938 228746 565174
rect 228982 564938 229066 565174
rect 229302 564938 229334 565174
rect 228714 564854 229334 564938
rect 228714 564618 228746 564854
rect 228982 564618 229066 564854
rect 229302 564618 229334 564854
rect 228714 527974 229334 564618
rect 228714 527738 228746 527974
rect 228982 527738 229066 527974
rect 229302 527738 229334 527974
rect 228714 527654 229334 527738
rect 228714 527418 228746 527654
rect 228982 527418 229066 527654
rect 229302 527418 229334 527654
rect 228714 490774 229334 527418
rect 228714 490538 228746 490774
rect 228982 490538 229066 490774
rect 229302 490538 229334 490774
rect 228714 490454 229334 490538
rect 228714 490218 228746 490454
rect 228982 490218 229066 490454
rect 229302 490218 229334 490454
rect 228714 453574 229334 490218
rect 228714 453338 228746 453574
rect 228982 453338 229066 453574
rect 229302 453338 229334 453574
rect 228714 453254 229334 453338
rect 228714 453018 228746 453254
rect 228982 453018 229066 453254
rect 229302 453018 229334 453254
rect 228714 416374 229334 453018
rect 228714 416138 228746 416374
rect 228982 416138 229066 416374
rect 229302 416138 229334 416374
rect 228714 416054 229334 416138
rect 228714 415818 228746 416054
rect 228982 415818 229066 416054
rect 229302 415818 229334 416054
rect 228714 379174 229334 415818
rect 228714 378938 228746 379174
rect 228982 378938 229066 379174
rect 229302 378938 229334 379174
rect 228714 378854 229334 378938
rect 228714 378618 228746 378854
rect 228982 378618 229066 378854
rect 229302 378618 229334 378854
rect 228714 341974 229334 378618
rect 228714 341738 228746 341974
rect 228982 341738 229066 341974
rect 229302 341738 229334 341974
rect 228714 341654 229334 341738
rect 228714 341418 228746 341654
rect 228982 341418 229066 341654
rect 229302 341418 229334 341654
rect 228714 304774 229334 341418
rect 228714 304538 228746 304774
rect 228982 304538 229066 304774
rect 229302 304538 229334 304774
rect 228714 304454 229334 304538
rect 228714 304218 228746 304454
rect 228982 304218 229066 304454
rect 229302 304218 229334 304454
rect 228714 267574 229334 304218
rect 228714 267338 228746 267574
rect 228982 267338 229066 267574
rect 229302 267338 229334 267574
rect 228714 267254 229334 267338
rect 228714 267018 228746 267254
rect 228982 267018 229066 267254
rect 229302 267018 229334 267254
rect 228714 230374 229334 267018
rect 228714 230138 228746 230374
rect 228982 230138 229066 230374
rect 229302 230138 229334 230374
rect 228714 230054 229334 230138
rect 228714 229818 228746 230054
rect 228982 229818 229066 230054
rect 229302 229818 229334 230054
rect 228714 193174 229334 229818
rect 228714 192938 228746 193174
rect 228982 192938 229066 193174
rect 229302 192938 229334 193174
rect 228714 192854 229334 192938
rect 228714 192618 228746 192854
rect 228982 192618 229066 192854
rect 229302 192618 229334 192854
rect 228714 155974 229334 192618
rect 228714 155738 228746 155974
rect 228982 155738 229066 155974
rect 229302 155738 229334 155974
rect 228714 155654 229334 155738
rect 228714 155418 228746 155654
rect 228982 155418 229066 155654
rect 229302 155418 229334 155654
rect 228714 118774 229334 155418
rect 228714 118538 228746 118774
rect 228982 118538 229066 118774
rect 229302 118538 229334 118774
rect 228714 118454 229334 118538
rect 228714 118218 228746 118454
rect 228982 118218 229066 118454
rect 229302 118218 229334 118454
rect 228714 81574 229334 118218
rect 228714 81338 228746 81574
rect 228982 81338 229066 81574
rect 229302 81338 229334 81574
rect 228714 81254 229334 81338
rect 228714 81018 228746 81254
rect 228982 81018 229066 81254
rect 229302 81018 229334 81254
rect 228714 44374 229334 81018
rect 228714 44138 228746 44374
rect 228982 44138 229066 44374
rect 229302 44138 229334 44374
rect 228714 44054 229334 44138
rect 228714 43818 228746 44054
rect 228982 43818 229066 44054
rect 229302 43818 229334 44054
rect 228714 7174 229334 43818
rect 228714 6938 228746 7174
rect 228982 6938 229066 7174
rect 229302 6938 229334 7174
rect 228714 6854 229334 6938
rect 228714 6618 228746 6854
rect 228982 6618 229066 6854
rect 229302 6618 229334 6854
rect 228714 2176 229334 6618
rect 232434 680494 233054 701760
rect 232434 680258 232466 680494
rect 232702 680258 232786 680494
rect 233022 680258 233054 680494
rect 232434 680174 233054 680258
rect 232434 679938 232466 680174
rect 232702 679938 232786 680174
rect 233022 679938 233054 680174
rect 232434 643294 233054 679938
rect 232434 643058 232466 643294
rect 232702 643058 232786 643294
rect 233022 643058 233054 643294
rect 232434 642974 233054 643058
rect 232434 642738 232466 642974
rect 232702 642738 232786 642974
rect 233022 642738 233054 642974
rect 232434 606094 233054 642738
rect 232434 605858 232466 606094
rect 232702 605858 232786 606094
rect 233022 605858 233054 606094
rect 232434 605774 233054 605858
rect 232434 605538 232466 605774
rect 232702 605538 232786 605774
rect 233022 605538 233054 605774
rect 232434 568894 233054 605538
rect 232434 568658 232466 568894
rect 232702 568658 232786 568894
rect 233022 568658 233054 568894
rect 232434 568574 233054 568658
rect 232434 568338 232466 568574
rect 232702 568338 232786 568574
rect 233022 568338 233054 568574
rect 232434 531694 233054 568338
rect 232434 531458 232466 531694
rect 232702 531458 232786 531694
rect 233022 531458 233054 531694
rect 232434 531374 233054 531458
rect 232434 531138 232466 531374
rect 232702 531138 232786 531374
rect 233022 531138 233054 531374
rect 232434 494494 233054 531138
rect 232434 494258 232466 494494
rect 232702 494258 232786 494494
rect 233022 494258 233054 494494
rect 232434 494174 233054 494258
rect 232434 493938 232466 494174
rect 232702 493938 232786 494174
rect 233022 493938 233054 494174
rect 232434 457294 233054 493938
rect 232434 457058 232466 457294
rect 232702 457058 232786 457294
rect 233022 457058 233054 457294
rect 232434 456974 233054 457058
rect 232434 456738 232466 456974
rect 232702 456738 232786 456974
rect 233022 456738 233054 456974
rect 232434 420094 233054 456738
rect 232434 419858 232466 420094
rect 232702 419858 232786 420094
rect 233022 419858 233054 420094
rect 232434 419774 233054 419858
rect 232434 419538 232466 419774
rect 232702 419538 232786 419774
rect 233022 419538 233054 419774
rect 232434 382894 233054 419538
rect 232434 382658 232466 382894
rect 232702 382658 232786 382894
rect 233022 382658 233054 382894
rect 232434 382574 233054 382658
rect 232434 382338 232466 382574
rect 232702 382338 232786 382574
rect 233022 382338 233054 382574
rect 232434 345694 233054 382338
rect 232434 345458 232466 345694
rect 232702 345458 232786 345694
rect 233022 345458 233054 345694
rect 232434 345374 233054 345458
rect 232434 345138 232466 345374
rect 232702 345138 232786 345374
rect 233022 345138 233054 345374
rect 232434 308494 233054 345138
rect 232434 308258 232466 308494
rect 232702 308258 232786 308494
rect 233022 308258 233054 308494
rect 232434 308174 233054 308258
rect 232434 307938 232466 308174
rect 232702 307938 232786 308174
rect 233022 307938 233054 308174
rect 232434 271294 233054 307938
rect 232434 271058 232466 271294
rect 232702 271058 232786 271294
rect 233022 271058 233054 271294
rect 232434 270974 233054 271058
rect 232434 270738 232466 270974
rect 232702 270738 232786 270974
rect 233022 270738 233054 270974
rect 232434 234094 233054 270738
rect 232434 233858 232466 234094
rect 232702 233858 232786 234094
rect 233022 233858 233054 234094
rect 232434 233774 233054 233858
rect 232434 233538 232466 233774
rect 232702 233538 232786 233774
rect 233022 233538 233054 233774
rect 232434 196894 233054 233538
rect 232434 196658 232466 196894
rect 232702 196658 232786 196894
rect 233022 196658 233054 196894
rect 232434 196574 233054 196658
rect 232434 196338 232466 196574
rect 232702 196338 232786 196574
rect 233022 196338 233054 196574
rect 232434 159694 233054 196338
rect 232434 159458 232466 159694
rect 232702 159458 232786 159694
rect 233022 159458 233054 159694
rect 232434 159374 233054 159458
rect 232434 159138 232466 159374
rect 232702 159138 232786 159374
rect 233022 159138 233054 159374
rect 232434 122494 233054 159138
rect 232434 122258 232466 122494
rect 232702 122258 232786 122494
rect 233022 122258 233054 122494
rect 232434 122174 233054 122258
rect 232434 121938 232466 122174
rect 232702 121938 232786 122174
rect 233022 121938 233054 122174
rect 232434 85294 233054 121938
rect 232434 85058 232466 85294
rect 232702 85058 232786 85294
rect 233022 85058 233054 85294
rect 232434 84974 233054 85058
rect 232434 84738 232466 84974
rect 232702 84738 232786 84974
rect 233022 84738 233054 84974
rect 232434 48094 233054 84738
rect 232434 47858 232466 48094
rect 232702 47858 232786 48094
rect 233022 47858 233054 48094
rect 232434 47774 233054 47858
rect 232434 47538 232466 47774
rect 232702 47538 232786 47774
rect 233022 47538 233054 47774
rect 232434 10894 233054 47538
rect 232434 10658 232466 10894
rect 232702 10658 232786 10894
rect 233022 10658 233054 10894
rect 232434 10574 233054 10658
rect 232434 10338 232466 10574
rect 232702 10338 232786 10574
rect 233022 10338 233054 10574
rect 232434 2176 233054 10338
rect 236154 684214 236774 701760
rect 236154 683978 236186 684214
rect 236422 683978 236506 684214
rect 236742 683978 236774 684214
rect 236154 683894 236774 683978
rect 236154 683658 236186 683894
rect 236422 683658 236506 683894
rect 236742 683658 236774 683894
rect 236154 647014 236774 683658
rect 236154 646778 236186 647014
rect 236422 646778 236506 647014
rect 236742 646778 236774 647014
rect 236154 646694 236774 646778
rect 236154 646458 236186 646694
rect 236422 646458 236506 646694
rect 236742 646458 236774 646694
rect 236154 609814 236774 646458
rect 236154 609578 236186 609814
rect 236422 609578 236506 609814
rect 236742 609578 236774 609814
rect 236154 609494 236774 609578
rect 236154 609258 236186 609494
rect 236422 609258 236506 609494
rect 236742 609258 236774 609494
rect 236154 572614 236774 609258
rect 236154 572378 236186 572614
rect 236422 572378 236506 572614
rect 236742 572378 236774 572614
rect 236154 572294 236774 572378
rect 236154 572058 236186 572294
rect 236422 572058 236506 572294
rect 236742 572058 236774 572294
rect 236154 535414 236774 572058
rect 236154 535178 236186 535414
rect 236422 535178 236506 535414
rect 236742 535178 236774 535414
rect 236154 535094 236774 535178
rect 236154 534858 236186 535094
rect 236422 534858 236506 535094
rect 236742 534858 236774 535094
rect 236154 498214 236774 534858
rect 236154 497978 236186 498214
rect 236422 497978 236506 498214
rect 236742 497978 236774 498214
rect 236154 497894 236774 497978
rect 236154 497658 236186 497894
rect 236422 497658 236506 497894
rect 236742 497658 236774 497894
rect 236154 461014 236774 497658
rect 236154 460778 236186 461014
rect 236422 460778 236506 461014
rect 236742 460778 236774 461014
rect 236154 460694 236774 460778
rect 236154 460458 236186 460694
rect 236422 460458 236506 460694
rect 236742 460458 236774 460694
rect 236154 423814 236774 460458
rect 236154 423578 236186 423814
rect 236422 423578 236506 423814
rect 236742 423578 236774 423814
rect 236154 423494 236774 423578
rect 236154 423258 236186 423494
rect 236422 423258 236506 423494
rect 236742 423258 236774 423494
rect 236154 386614 236774 423258
rect 236154 386378 236186 386614
rect 236422 386378 236506 386614
rect 236742 386378 236774 386614
rect 236154 386294 236774 386378
rect 236154 386058 236186 386294
rect 236422 386058 236506 386294
rect 236742 386058 236774 386294
rect 236154 349414 236774 386058
rect 236154 349178 236186 349414
rect 236422 349178 236506 349414
rect 236742 349178 236774 349414
rect 236154 349094 236774 349178
rect 236154 348858 236186 349094
rect 236422 348858 236506 349094
rect 236742 348858 236774 349094
rect 236154 312214 236774 348858
rect 236154 311978 236186 312214
rect 236422 311978 236506 312214
rect 236742 311978 236774 312214
rect 236154 311894 236774 311978
rect 236154 311658 236186 311894
rect 236422 311658 236506 311894
rect 236742 311658 236774 311894
rect 236154 275014 236774 311658
rect 236154 274778 236186 275014
rect 236422 274778 236506 275014
rect 236742 274778 236774 275014
rect 236154 274694 236774 274778
rect 236154 274458 236186 274694
rect 236422 274458 236506 274694
rect 236742 274458 236774 274694
rect 236154 237814 236774 274458
rect 236154 237578 236186 237814
rect 236422 237578 236506 237814
rect 236742 237578 236774 237814
rect 236154 237494 236774 237578
rect 236154 237258 236186 237494
rect 236422 237258 236506 237494
rect 236742 237258 236774 237494
rect 236154 200614 236774 237258
rect 236154 200378 236186 200614
rect 236422 200378 236506 200614
rect 236742 200378 236774 200614
rect 236154 200294 236774 200378
rect 236154 200058 236186 200294
rect 236422 200058 236506 200294
rect 236742 200058 236774 200294
rect 236154 163414 236774 200058
rect 236154 163178 236186 163414
rect 236422 163178 236506 163414
rect 236742 163178 236774 163414
rect 236154 163094 236774 163178
rect 236154 162858 236186 163094
rect 236422 162858 236506 163094
rect 236742 162858 236774 163094
rect 236154 126214 236774 162858
rect 236154 125978 236186 126214
rect 236422 125978 236506 126214
rect 236742 125978 236774 126214
rect 236154 125894 236774 125978
rect 236154 125658 236186 125894
rect 236422 125658 236506 125894
rect 236742 125658 236774 125894
rect 236154 89014 236774 125658
rect 236154 88778 236186 89014
rect 236422 88778 236506 89014
rect 236742 88778 236774 89014
rect 236154 88694 236774 88778
rect 236154 88458 236186 88694
rect 236422 88458 236506 88694
rect 236742 88458 236774 88694
rect 236154 51814 236774 88458
rect 236154 51578 236186 51814
rect 236422 51578 236506 51814
rect 236742 51578 236774 51814
rect 236154 51494 236774 51578
rect 236154 51258 236186 51494
rect 236422 51258 236506 51494
rect 236742 51258 236774 51494
rect 236154 14614 236774 51258
rect 236154 14378 236186 14614
rect 236422 14378 236506 14614
rect 236742 14378 236774 14614
rect 236154 14294 236774 14378
rect 236154 14058 236186 14294
rect 236422 14058 236506 14294
rect 236742 14058 236774 14294
rect 236154 2176 236774 14058
rect 239874 687934 240494 701760
rect 239874 687698 239906 687934
rect 240142 687698 240226 687934
rect 240462 687698 240494 687934
rect 239874 687614 240494 687698
rect 239874 687378 239906 687614
rect 240142 687378 240226 687614
rect 240462 687378 240494 687614
rect 239874 650734 240494 687378
rect 239874 650498 239906 650734
rect 240142 650498 240226 650734
rect 240462 650498 240494 650734
rect 239874 650414 240494 650498
rect 239874 650178 239906 650414
rect 240142 650178 240226 650414
rect 240462 650178 240494 650414
rect 239874 613534 240494 650178
rect 239874 613298 239906 613534
rect 240142 613298 240226 613534
rect 240462 613298 240494 613534
rect 239874 613214 240494 613298
rect 239874 612978 239906 613214
rect 240142 612978 240226 613214
rect 240462 612978 240494 613214
rect 239874 576334 240494 612978
rect 239874 576098 239906 576334
rect 240142 576098 240226 576334
rect 240462 576098 240494 576334
rect 239874 576014 240494 576098
rect 239874 575778 239906 576014
rect 240142 575778 240226 576014
rect 240462 575778 240494 576014
rect 239874 539134 240494 575778
rect 239874 538898 239906 539134
rect 240142 538898 240226 539134
rect 240462 538898 240494 539134
rect 239874 538814 240494 538898
rect 239874 538578 239906 538814
rect 240142 538578 240226 538814
rect 240462 538578 240494 538814
rect 239874 501934 240494 538578
rect 239874 501698 239906 501934
rect 240142 501698 240226 501934
rect 240462 501698 240494 501934
rect 239874 501614 240494 501698
rect 239874 501378 239906 501614
rect 240142 501378 240226 501614
rect 240462 501378 240494 501614
rect 239874 464734 240494 501378
rect 239874 464498 239906 464734
rect 240142 464498 240226 464734
rect 240462 464498 240494 464734
rect 239874 464414 240494 464498
rect 239874 464178 239906 464414
rect 240142 464178 240226 464414
rect 240462 464178 240494 464414
rect 239874 427534 240494 464178
rect 239874 427298 239906 427534
rect 240142 427298 240226 427534
rect 240462 427298 240494 427534
rect 239874 427214 240494 427298
rect 239874 426978 239906 427214
rect 240142 426978 240226 427214
rect 240462 426978 240494 427214
rect 239874 390334 240494 426978
rect 239874 390098 239906 390334
rect 240142 390098 240226 390334
rect 240462 390098 240494 390334
rect 239874 390014 240494 390098
rect 239874 389778 239906 390014
rect 240142 389778 240226 390014
rect 240462 389778 240494 390014
rect 239874 353134 240494 389778
rect 239874 352898 239906 353134
rect 240142 352898 240226 353134
rect 240462 352898 240494 353134
rect 239874 352814 240494 352898
rect 239874 352578 239906 352814
rect 240142 352578 240226 352814
rect 240462 352578 240494 352814
rect 239874 315934 240494 352578
rect 239874 315698 239906 315934
rect 240142 315698 240226 315934
rect 240462 315698 240494 315934
rect 239874 315614 240494 315698
rect 239874 315378 239906 315614
rect 240142 315378 240226 315614
rect 240462 315378 240494 315614
rect 239874 278734 240494 315378
rect 239874 278498 239906 278734
rect 240142 278498 240226 278734
rect 240462 278498 240494 278734
rect 239874 278414 240494 278498
rect 239874 278178 239906 278414
rect 240142 278178 240226 278414
rect 240462 278178 240494 278414
rect 239874 241534 240494 278178
rect 239874 241298 239906 241534
rect 240142 241298 240226 241534
rect 240462 241298 240494 241534
rect 239874 241214 240494 241298
rect 239874 240978 239906 241214
rect 240142 240978 240226 241214
rect 240462 240978 240494 241214
rect 239874 204334 240494 240978
rect 239874 204098 239906 204334
rect 240142 204098 240226 204334
rect 240462 204098 240494 204334
rect 239874 204014 240494 204098
rect 239874 203778 239906 204014
rect 240142 203778 240226 204014
rect 240462 203778 240494 204014
rect 239874 167134 240494 203778
rect 239874 166898 239906 167134
rect 240142 166898 240226 167134
rect 240462 166898 240494 167134
rect 239874 166814 240494 166898
rect 239874 166578 239906 166814
rect 240142 166578 240226 166814
rect 240462 166578 240494 166814
rect 239874 129934 240494 166578
rect 239874 129698 239906 129934
rect 240142 129698 240226 129934
rect 240462 129698 240494 129934
rect 239874 129614 240494 129698
rect 239874 129378 239906 129614
rect 240142 129378 240226 129614
rect 240462 129378 240494 129614
rect 239874 92734 240494 129378
rect 239874 92498 239906 92734
rect 240142 92498 240226 92734
rect 240462 92498 240494 92734
rect 239874 92414 240494 92498
rect 239874 92178 239906 92414
rect 240142 92178 240226 92414
rect 240462 92178 240494 92414
rect 239874 55534 240494 92178
rect 239874 55298 239906 55534
rect 240142 55298 240226 55534
rect 240462 55298 240494 55534
rect 239874 55214 240494 55298
rect 239874 54978 239906 55214
rect 240142 54978 240226 55214
rect 240462 54978 240494 55214
rect 239874 18334 240494 54978
rect 239874 18098 239906 18334
rect 240142 18098 240226 18334
rect 240462 18098 240494 18334
rect 239874 18014 240494 18098
rect 239874 17778 239906 18014
rect 240142 17778 240226 18014
rect 240462 17778 240494 18014
rect 239874 2176 240494 17778
rect 243594 691654 244214 701760
rect 243594 691418 243626 691654
rect 243862 691418 243946 691654
rect 244182 691418 244214 691654
rect 243594 691334 244214 691418
rect 243594 691098 243626 691334
rect 243862 691098 243946 691334
rect 244182 691098 244214 691334
rect 243594 654454 244214 691098
rect 243594 654218 243626 654454
rect 243862 654218 243946 654454
rect 244182 654218 244214 654454
rect 243594 654134 244214 654218
rect 243594 653898 243626 654134
rect 243862 653898 243946 654134
rect 244182 653898 244214 654134
rect 243594 617254 244214 653898
rect 243594 617018 243626 617254
rect 243862 617018 243946 617254
rect 244182 617018 244214 617254
rect 243594 616934 244214 617018
rect 243594 616698 243626 616934
rect 243862 616698 243946 616934
rect 244182 616698 244214 616934
rect 243594 580054 244214 616698
rect 243594 579818 243626 580054
rect 243862 579818 243946 580054
rect 244182 579818 244214 580054
rect 243594 579734 244214 579818
rect 243594 579498 243626 579734
rect 243862 579498 243946 579734
rect 244182 579498 244214 579734
rect 243594 542854 244214 579498
rect 243594 542618 243626 542854
rect 243862 542618 243946 542854
rect 244182 542618 244214 542854
rect 243594 542534 244214 542618
rect 243594 542298 243626 542534
rect 243862 542298 243946 542534
rect 244182 542298 244214 542534
rect 243594 505654 244214 542298
rect 243594 505418 243626 505654
rect 243862 505418 243946 505654
rect 244182 505418 244214 505654
rect 243594 505334 244214 505418
rect 243594 505098 243626 505334
rect 243862 505098 243946 505334
rect 244182 505098 244214 505334
rect 243594 468454 244214 505098
rect 243594 468218 243626 468454
rect 243862 468218 243946 468454
rect 244182 468218 244214 468454
rect 243594 468134 244214 468218
rect 243594 467898 243626 468134
rect 243862 467898 243946 468134
rect 244182 467898 244214 468134
rect 243594 431254 244214 467898
rect 243594 431018 243626 431254
rect 243862 431018 243946 431254
rect 244182 431018 244214 431254
rect 243594 430934 244214 431018
rect 243594 430698 243626 430934
rect 243862 430698 243946 430934
rect 244182 430698 244214 430934
rect 243594 394054 244214 430698
rect 243594 393818 243626 394054
rect 243862 393818 243946 394054
rect 244182 393818 244214 394054
rect 243594 393734 244214 393818
rect 243594 393498 243626 393734
rect 243862 393498 243946 393734
rect 244182 393498 244214 393734
rect 243594 356854 244214 393498
rect 243594 356618 243626 356854
rect 243862 356618 243946 356854
rect 244182 356618 244214 356854
rect 243594 356534 244214 356618
rect 243594 356298 243626 356534
rect 243862 356298 243946 356534
rect 244182 356298 244214 356534
rect 243594 319654 244214 356298
rect 243594 319418 243626 319654
rect 243862 319418 243946 319654
rect 244182 319418 244214 319654
rect 243594 319334 244214 319418
rect 243594 319098 243626 319334
rect 243862 319098 243946 319334
rect 244182 319098 244214 319334
rect 243594 282454 244214 319098
rect 243594 282218 243626 282454
rect 243862 282218 243946 282454
rect 244182 282218 244214 282454
rect 243594 282134 244214 282218
rect 243594 281898 243626 282134
rect 243862 281898 243946 282134
rect 244182 281898 244214 282134
rect 243594 245254 244214 281898
rect 243594 245018 243626 245254
rect 243862 245018 243946 245254
rect 244182 245018 244214 245254
rect 243594 244934 244214 245018
rect 243594 244698 243626 244934
rect 243862 244698 243946 244934
rect 244182 244698 244214 244934
rect 243594 208054 244214 244698
rect 243594 207818 243626 208054
rect 243862 207818 243946 208054
rect 244182 207818 244214 208054
rect 243594 207734 244214 207818
rect 243594 207498 243626 207734
rect 243862 207498 243946 207734
rect 244182 207498 244214 207734
rect 243594 170854 244214 207498
rect 243594 170618 243626 170854
rect 243862 170618 243946 170854
rect 244182 170618 244214 170854
rect 243594 170534 244214 170618
rect 243594 170298 243626 170534
rect 243862 170298 243946 170534
rect 244182 170298 244214 170534
rect 243594 133654 244214 170298
rect 243594 133418 243626 133654
rect 243862 133418 243946 133654
rect 244182 133418 244214 133654
rect 243594 133334 244214 133418
rect 243594 133098 243626 133334
rect 243862 133098 243946 133334
rect 244182 133098 244214 133334
rect 243594 96454 244214 133098
rect 243594 96218 243626 96454
rect 243862 96218 243946 96454
rect 244182 96218 244214 96454
rect 243594 96134 244214 96218
rect 243594 95898 243626 96134
rect 243862 95898 243946 96134
rect 244182 95898 244214 96134
rect 243594 59254 244214 95898
rect 243594 59018 243626 59254
rect 243862 59018 243946 59254
rect 244182 59018 244214 59254
rect 243594 58934 244214 59018
rect 243594 58698 243626 58934
rect 243862 58698 243946 58934
rect 244182 58698 244214 58934
rect 243594 22054 244214 58698
rect 243594 21818 243626 22054
rect 243862 21818 243946 22054
rect 244182 21818 244214 22054
rect 243594 21734 244214 21818
rect 243594 21498 243626 21734
rect 243862 21498 243946 21734
rect 244182 21498 244214 21734
rect 243594 2176 244214 21498
rect 247314 695374 247934 701760
rect 247314 695138 247346 695374
rect 247582 695138 247666 695374
rect 247902 695138 247934 695374
rect 247314 695054 247934 695138
rect 247314 694818 247346 695054
rect 247582 694818 247666 695054
rect 247902 694818 247934 695054
rect 247314 658174 247934 694818
rect 247314 657938 247346 658174
rect 247582 657938 247666 658174
rect 247902 657938 247934 658174
rect 247314 657854 247934 657938
rect 247314 657618 247346 657854
rect 247582 657618 247666 657854
rect 247902 657618 247934 657854
rect 247314 620974 247934 657618
rect 247314 620738 247346 620974
rect 247582 620738 247666 620974
rect 247902 620738 247934 620974
rect 247314 620654 247934 620738
rect 247314 620418 247346 620654
rect 247582 620418 247666 620654
rect 247902 620418 247934 620654
rect 247314 583774 247934 620418
rect 247314 583538 247346 583774
rect 247582 583538 247666 583774
rect 247902 583538 247934 583774
rect 247314 583454 247934 583538
rect 247314 583218 247346 583454
rect 247582 583218 247666 583454
rect 247902 583218 247934 583454
rect 247314 546574 247934 583218
rect 247314 546338 247346 546574
rect 247582 546338 247666 546574
rect 247902 546338 247934 546574
rect 247314 546254 247934 546338
rect 247314 546018 247346 546254
rect 247582 546018 247666 546254
rect 247902 546018 247934 546254
rect 247314 509374 247934 546018
rect 247314 509138 247346 509374
rect 247582 509138 247666 509374
rect 247902 509138 247934 509374
rect 247314 509054 247934 509138
rect 247314 508818 247346 509054
rect 247582 508818 247666 509054
rect 247902 508818 247934 509054
rect 247314 472174 247934 508818
rect 247314 471938 247346 472174
rect 247582 471938 247666 472174
rect 247902 471938 247934 472174
rect 247314 471854 247934 471938
rect 247314 471618 247346 471854
rect 247582 471618 247666 471854
rect 247902 471618 247934 471854
rect 247314 434974 247934 471618
rect 247314 434738 247346 434974
rect 247582 434738 247666 434974
rect 247902 434738 247934 434974
rect 247314 434654 247934 434738
rect 247314 434418 247346 434654
rect 247582 434418 247666 434654
rect 247902 434418 247934 434654
rect 247314 397774 247934 434418
rect 247314 397538 247346 397774
rect 247582 397538 247666 397774
rect 247902 397538 247934 397774
rect 247314 397454 247934 397538
rect 247314 397218 247346 397454
rect 247582 397218 247666 397454
rect 247902 397218 247934 397454
rect 247314 360574 247934 397218
rect 247314 360338 247346 360574
rect 247582 360338 247666 360574
rect 247902 360338 247934 360574
rect 247314 360254 247934 360338
rect 247314 360018 247346 360254
rect 247582 360018 247666 360254
rect 247902 360018 247934 360254
rect 247314 323374 247934 360018
rect 247314 323138 247346 323374
rect 247582 323138 247666 323374
rect 247902 323138 247934 323374
rect 247314 323054 247934 323138
rect 247314 322818 247346 323054
rect 247582 322818 247666 323054
rect 247902 322818 247934 323054
rect 247314 286174 247934 322818
rect 247314 285938 247346 286174
rect 247582 285938 247666 286174
rect 247902 285938 247934 286174
rect 247314 285854 247934 285938
rect 247314 285618 247346 285854
rect 247582 285618 247666 285854
rect 247902 285618 247934 285854
rect 247314 248974 247934 285618
rect 247314 248738 247346 248974
rect 247582 248738 247666 248974
rect 247902 248738 247934 248974
rect 247314 248654 247934 248738
rect 247314 248418 247346 248654
rect 247582 248418 247666 248654
rect 247902 248418 247934 248654
rect 247314 211774 247934 248418
rect 247314 211538 247346 211774
rect 247582 211538 247666 211774
rect 247902 211538 247934 211774
rect 247314 211454 247934 211538
rect 247314 211218 247346 211454
rect 247582 211218 247666 211454
rect 247902 211218 247934 211454
rect 247314 174574 247934 211218
rect 247314 174338 247346 174574
rect 247582 174338 247666 174574
rect 247902 174338 247934 174574
rect 247314 174254 247934 174338
rect 247314 174018 247346 174254
rect 247582 174018 247666 174254
rect 247902 174018 247934 174254
rect 247314 137374 247934 174018
rect 247314 137138 247346 137374
rect 247582 137138 247666 137374
rect 247902 137138 247934 137374
rect 247314 137054 247934 137138
rect 247314 136818 247346 137054
rect 247582 136818 247666 137054
rect 247902 136818 247934 137054
rect 247314 100174 247934 136818
rect 247314 99938 247346 100174
rect 247582 99938 247666 100174
rect 247902 99938 247934 100174
rect 247314 99854 247934 99938
rect 247314 99618 247346 99854
rect 247582 99618 247666 99854
rect 247902 99618 247934 99854
rect 247314 62974 247934 99618
rect 247314 62738 247346 62974
rect 247582 62738 247666 62974
rect 247902 62738 247934 62974
rect 247314 62654 247934 62738
rect 247314 62418 247346 62654
rect 247582 62418 247666 62654
rect 247902 62418 247934 62654
rect 247314 25774 247934 62418
rect 247314 25538 247346 25774
rect 247582 25538 247666 25774
rect 247902 25538 247934 25774
rect 247314 25454 247934 25538
rect 247314 25218 247346 25454
rect 247582 25218 247666 25454
rect 247902 25218 247934 25454
rect 247314 2176 247934 25218
rect 251034 699094 251654 701760
rect 251034 698858 251066 699094
rect 251302 698858 251386 699094
rect 251622 698858 251654 699094
rect 251034 698774 251654 698858
rect 251034 698538 251066 698774
rect 251302 698538 251386 698774
rect 251622 698538 251654 698774
rect 251034 661894 251654 698538
rect 251034 661658 251066 661894
rect 251302 661658 251386 661894
rect 251622 661658 251654 661894
rect 251034 661574 251654 661658
rect 251034 661338 251066 661574
rect 251302 661338 251386 661574
rect 251622 661338 251654 661574
rect 251034 624694 251654 661338
rect 251034 624458 251066 624694
rect 251302 624458 251386 624694
rect 251622 624458 251654 624694
rect 251034 624374 251654 624458
rect 251034 624138 251066 624374
rect 251302 624138 251386 624374
rect 251622 624138 251654 624374
rect 251034 587494 251654 624138
rect 251034 587258 251066 587494
rect 251302 587258 251386 587494
rect 251622 587258 251654 587494
rect 251034 587174 251654 587258
rect 251034 586938 251066 587174
rect 251302 586938 251386 587174
rect 251622 586938 251654 587174
rect 251034 550294 251654 586938
rect 251034 550058 251066 550294
rect 251302 550058 251386 550294
rect 251622 550058 251654 550294
rect 251034 549974 251654 550058
rect 251034 549738 251066 549974
rect 251302 549738 251386 549974
rect 251622 549738 251654 549974
rect 251034 513094 251654 549738
rect 251034 512858 251066 513094
rect 251302 512858 251386 513094
rect 251622 512858 251654 513094
rect 251034 512774 251654 512858
rect 251034 512538 251066 512774
rect 251302 512538 251386 512774
rect 251622 512538 251654 512774
rect 251034 475894 251654 512538
rect 251034 475658 251066 475894
rect 251302 475658 251386 475894
rect 251622 475658 251654 475894
rect 251034 475574 251654 475658
rect 251034 475338 251066 475574
rect 251302 475338 251386 475574
rect 251622 475338 251654 475574
rect 251034 438694 251654 475338
rect 251034 438458 251066 438694
rect 251302 438458 251386 438694
rect 251622 438458 251654 438694
rect 251034 438374 251654 438458
rect 251034 438138 251066 438374
rect 251302 438138 251386 438374
rect 251622 438138 251654 438374
rect 251034 401494 251654 438138
rect 251034 401258 251066 401494
rect 251302 401258 251386 401494
rect 251622 401258 251654 401494
rect 251034 401174 251654 401258
rect 251034 400938 251066 401174
rect 251302 400938 251386 401174
rect 251622 400938 251654 401174
rect 251034 364294 251654 400938
rect 251034 364058 251066 364294
rect 251302 364058 251386 364294
rect 251622 364058 251654 364294
rect 251034 363974 251654 364058
rect 251034 363738 251066 363974
rect 251302 363738 251386 363974
rect 251622 363738 251654 363974
rect 251034 327094 251654 363738
rect 251034 326858 251066 327094
rect 251302 326858 251386 327094
rect 251622 326858 251654 327094
rect 251034 326774 251654 326858
rect 251034 326538 251066 326774
rect 251302 326538 251386 326774
rect 251622 326538 251654 326774
rect 251034 289894 251654 326538
rect 251034 289658 251066 289894
rect 251302 289658 251386 289894
rect 251622 289658 251654 289894
rect 251034 289574 251654 289658
rect 251034 289338 251066 289574
rect 251302 289338 251386 289574
rect 251622 289338 251654 289574
rect 251034 252694 251654 289338
rect 251034 252458 251066 252694
rect 251302 252458 251386 252694
rect 251622 252458 251654 252694
rect 251034 252374 251654 252458
rect 251034 252138 251066 252374
rect 251302 252138 251386 252374
rect 251622 252138 251654 252374
rect 251034 215494 251654 252138
rect 251034 215258 251066 215494
rect 251302 215258 251386 215494
rect 251622 215258 251654 215494
rect 251034 215174 251654 215258
rect 251034 214938 251066 215174
rect 251302 214938 251386 215174
rect 251622 214938 251654 215174
rect 251034 178294 251654 214938
rect 251034 178058 251066 178294
rect 251302 178058 251386 178294
rect 251622 178058 251654 178294
rect 251034 177974 251654 178058
rect 251034 177738 251066 177974
rect 251302 177738 251386 177974
rect 251622 177738 251654 177974
rect 251034 141094 251654 177738
rect 251034 140858 251066 141094
rect 251302 140858 251386 141094
rect 251622 140858 251654 141094
rect 251034 140774 251654 140858
rect 251034 140538 251066 140774
rect 251302 140538 251386 140774
rect 251622 140538 251654 140774
rect 251034 103894 251654 140538
rect 251034 103658 251066 103894
rect 251302 103658 251386 103894
rect 251622 103658 251654 103894
rect 251034 103574 251654 103658
rect 251034 103338 251066 103574
rect 251302 103338 251386 103574
rect 251622 103338 251654 103574
rect 251034 66694 251654 103338
rect 251034 66458 251066 66694
rect 251302 66458 251386 66694
rect 251622 66458 251654 66694
rect 251034 66374 251654 66458
rect 251034 66138 251066 66374
rect 251302 66138 251386 66374
rect 251622 66138 251654 66374
rect 251034 29494 251654 66138
rect 251034 29258 251066 29494
rect 251302 29258 251386 29494
rect 251622 29258 251654 29494
rect 251034 29174 251654 29258
rect 251034 28938 251066 29174
rect 251302 28938 251386 29174
rect 251622 28938 251654 29174
rect 251034 2176 251654 28938
rect 262194 673054 262814 701760
rect 262194 672818 262226 673054
rect 262462 672818 262546 673054
rect 262782 672818 262814 673054
rect 262194 672734 262814 672818
rect 262194 672498 262226 672734
rect 262462 672498 262546 672734
rect 262782 672498 262814 672734
rect 262194 635854 262814 672498
rect 262194 635618 262226 635854
rect 262462 635618 262546 635854
rect 262782 635618 262814 635854
rect 262194 635534 262814 635618
rect 262194 635298 262226 635534
rect 262462 635298 262546 635534
rect 262782 635298 262814 635534
rect 262194 598654 262814 635298
rect 262194 598418 262226 598654
rect 262462 598418 262546 598654
rect 262782 598418 262814 598654
rect 262194 598334 262814 598418
rect 262194 598098 262226 598334
rect 262462 598098 262546 598334
rect 262782 598098 262814 598334
rect 262194 561454 262814 598098
rect 262194 561218 262226 561454
rect 262462 561218 262546 561454
rect 262782 561218 262814 561454
rect 262194 561134 262814 561218
rect 262194 560898 262226 561134
rect 262462 560898 262546 561134
rect 262782 560898 262814 561134
rect 262194 524254 262814 560898
rect 262194 524018 262226 524254
rect 262462 524018 262546 524254
rect 262782 524018 262814 524254
rect 262194 523934 262814 524018
rect 262194 523698 262226 523934
rect 262462 523698 262546 523934
rect 262782 523698 262814 523934
rect 262194 487054 262814 523698
rect 262194 486818 262226 487054
rect 262462 486818 262546 487054
rect 262782 486818 262814 487054
rect 262194 486734 262814 486818
rect 262194 486498 262226 486734
rect 262462 486498 262546 486734
rect 262782 486498 262814 486734
rect 262194 449854 262814 486498
rect 262194 449618 262226 449854
rect 262462 449618 262546 449854
rect 262782 449618 262814 449854
rect 262194 449534 262814 449618
rect 262194 449298 262226 449534
rect 262462 449298 262546 449534
rect 262782 449298 262814 449534
rect 262194 412654 262814 449298
rect 262194 412418 262226 412654
rect 262462 412418 262546 412654
rect 262782 412418 262814 412654
rect 262194 412334 262814 412418
rect 262194 412098 262226 412334
rect 262462 412098 262546 412334
rect 262782 412098 262814 412334
rect 262194 375454 262814 412098
rect 262194 375218 262226 375454
rect 262462 375218 262546 375454
rect 262782 375218 262814 375454
rect 262194 375134 262814 375218
rect 262194 374898 262226 375134
rect 262462 374898 262546 375134
rect 262782 374898 262814 375134
rect 262194 338254 262814 374898
rect 262194 338018 262226 338254
rect 262462 338018 262546 338254
rect 262782 338018 262814 338254
rect 262194 337934 262814 338018
rect 262194 337698 262226 337934
rect 262462 337698 262546 337934
rect 262782 337698 262814 337934
rect 262194 301054 262814 337698
rect 262194 300818 262226 301054
rect 262462 300818 262546 301054
rect 262782 300818 262814 301054
rect 262194 300734 262814 300818
rect 262194 300498 262226 300734
rect 262462 300498 262546 300734
rect 262782 300498 262814 300734
rect 262194 263854 262814 300498
rect 262194 263618 262226 263854
rect 262462 263618 262546 263854
rect 262782 263618 262814 263854
rect 262194 263534 262814 263618
rect 262194 263298 262226 263534
rect 262462 263298 262546 263534
rect 262782 263298 262814 263534
rect 262194 226654 262814 263298
rect 262194 226418 262226 226654
rect 262462 226418 262546 226654
rect 262782 226418 262814 226654
rect 262194 226334 262814 226418
rect 262194 226098 262226 226334
rect 262462 226098 262546 226334
rect 262782 226098 262814 226334
rect 262194 189454 262814 226098
rect 262194 189218 262226 189454
rect 262462 189218 262546 189454
rect 262782 189218 262814 189454
rect 262194 189134 262814 189218
rect 262194 188898 262226 189134
rect 262462 188898 262546 189134
rect 262782 188898 262814 189134
rect 262194 152254 262814 188898
rect 262194 152018 262226 152254
rect 262462 152018 262546 152254
rect 262782 152018 262814 152254
rect 262194 151934 262814 152018
rect 262194 151698 262226 151934
rect 262462 151698 262546 151934
rect 262782 151698 262814 151934
rect 262194 115054 262814 151698
rect 262194 114818 262226 115054
rect 262462 114818 262546 115054
rect 262782 114818 262814 115054
rect 262194 114734 262814 114818
rect 262194 114498 262226 114734
rect 262462 114498 262546 114734
rect 262782 114498 262814 114734
rect 262194 77854 262814 114498
rect 262194 77618 262226 77854
rect 262462 77618 262546 77854
rect 262782 77618 262814 77854
rect 262194 77534 262814 77618
rect 262194 77298 262226 77534
rect 262462 77298 262546 77534
rect 262782 77298 262814 77534
rect 262194 40654 262814 77298
rect 262194 40418 262226 40654
rect 262462 40418 262546 40654
rect 262782 40418 262814 40654
rect 262194 40334 262814 40418
rect 262194 40098 262226 40334
rect 262462 40098 262546 40334
rect 262782 40098 262814 40334
rect 262194 3454 262814 40098
rect 262194 3218 262226 3454
rect 262462 3218 262546 3454
rect 262782 3218 262814 3454
rect 262194 3134 262814 3218
rect 262194 2898 262226 3134
rect 262462 2898 262546 3134
rect 262782 2898 262814 3134
rect 262194 2176 262814 2898
rect 265914 676774 266534 701760
rect 265914 676538 265946 676774
rect 266182 676538 266266 676774
rect 266502 676538 266534 676774
rect 265914 676454 266534 676538
rect 265914 676218 265946 676454
rect 266182 676218 266266 676454
rect 266502 676218 266534 676454
rect 265914 639574 266534 676218
rect 265914 639338 265946 639574
rect 266182 639338 266266 639574
rect 266502 639338 266534 639574
rect 265914 639254 266534 639338
rect 265914 639018 265946 639254
rect 266182 639018 266266 639254
rect 266502 639018 266534 639254
rect 265914 602374 266534 639018
rect 265914 602138 265946 602374
rect 266182 602138 266266 602374
rect 266502 602138 266534 602374
rect 265914 602054 266534 602138
rect 265914 601818 265946 602054
rect 266182 601818 266266 602054
rect 266502 601818 266534 602054
rect 265914 565174 266534 601818
rect 265914 564938 265946 565174
rect 266182 564938 266266 565174
rect 266502 564938 266534 565174
rect 265914 564854 266534 564938
rect 265914 564618 265946 564854
rect 266182 564618 266266 564854
rect 266502 564618 266534 564854
rect 265914 527974 266534 564618
rect 265914 527738 265946 527974
rect 266182 527738 266266 527974
rect 266502 527738 266534 527974
rect 265914 527654 266534 527738
rect 265914 527418 265946 527654
rect 266182 527418 266266 527654
rect 266502 527418 266534 527654
rect 265914 490774 266534 527418
rect 265914 490538 265946 490774
rect 266182 490538 266266 490774
rect 266502 490538 266534 490774
rect 265914 490454 266534 490538
rect 265914 490218 265946 490454
rect 266182 490218 266266 490454
rect 266502 490218 266534 490454
rect 265914 453574 266534 490218
rect 265914 453338 265946 453574
rect 266182 453338 266266 453574
rect 266502 453338 266534 453574
rect 265914 453254 266534 453338
rect 265914 453018 265946 453254
rect 266182 453018 266266 453254
rect 266502 453018 266534 453254
rect 265914 416374 266534 453018
rect 265914 416138 265946 416374
rect 266182 416138 266266 416374
rect 266502 416138 266534 416374
rect 265914 416054 266534 416138
rect 265914 415818 265946 416054
rect 266182 415818 266266 416054
rect 266502 415818 266534 416054
rect 265914 379174 266534 415818
rect 265914 378938 265946 379174
rect 266182 378938 266266 379174
rect 266502 378938 266534 379174
rect 265914 378854 266534 378938
rect 265914 378618 265946 378854
rect 266182 378618 266266 378854
rect 266502 378618 266534 378854
rect 265914 341974 266534 378618
rect 265914 341738 265946 341974
rect 266182 341738 266266 341974
rect 266502 341738 266534 341974
rect 265914 341654 266534 341738
rect 265914 341418 265946 341654
rect 266182 341418 266266 341654
rect 266502 341418 266534 341654
rect 265914 304774 266534 341418
rect 265914 304538 265946 304774
rect 266182 304538 266266 304774
rect 266502 304538 266534 304774
rect 265914 304454 266534 304538
rect 265914 304218 265946 304454
rect 266182 304218 266266 304454
rect 266502 304218 266534 304454
rect 265914 267574 266534 304218
rect 265914 267338 265946 267574
rect 266182 267338 266266 267574
rect 266502 267338 266534 267574
rect 265914 267254 266534 267338
rect 265914 267018 265946 267254
rect 266182 267018 266266 267254
rect 266502 267018 266534 267254
rect 265914 230374 266534 267018
rect 265914 230138 265946 230374
rect 266182 230138 266266 230374
rect 266502 230138 266534 230374
rect 265914 230054 266534 230138
rect 265914 229818 265946 230054
rect 266182 229818 266266 230054
rect 266502 229818 266534 230054
rect 265914 193174 266534 229818
rect 265914 192938 265946 193174
rect 266182 192938 266266 193174
rect 266502 192938 266534 193174
rect 265914 192854 266534 192938
rect 265914 192618 265946 192854
rect 266182 192618 266266 192854
rect 266502 192618 266534 192854
rect 265914 155974 266534 192618
rect 265914 155738 265946 155974
rect 266182 155738 266266 155974
rect 266502 155738 266534 155974
rect 265914 155654 266534 155738
rect 265914 155418 265946 155654
rect 266182 155418 266266 155654
rect 266502 155418 266534 155654
rect 265914 118774 266534 155418
rect 265914 118538 265946 118774
rect 266182 118538 266266 118774
rect 266502 118538 266534 118774
rect 265914 118454 266534 118538
rect 265914 118218 265946 118454
rect 266182 118218 266266 118454
rect 266502 118218 266534 118454
rect 265914 81574 266534 118218
rect 265914 81338 265946 81574
rect 266182 81338 266266 81574
rect 266502 81338 266534 81574
rect 265914 81254 266534 81338
rect 265914 81018 265946 81254
rect 266182 81018 266266 81254
rect 266502 81018 266534 81254
rect 265914 44374 266534 81018
rect 265914 44138 265946 44374
rect 266182 44138 266266 44374
rect 266502 44138 266534 44374
rect 265914 44054 266534 44138
rect 265914 43818 265946 44054
rect 266182 43818 266266 44054
rect 266502 43818 266534 44054
rect 265914 7174 266534 43818
rect 265914 6938 265946 7174
rect 266182 6938 266266 7174
rect 266502 6938 266534 7174
rect 265914 6854 266534 6938
rect 265914 6618 265946 6854
rect 266182 6618 266266 6854
rect 266502 6618 266534 6854
rect 265914 2176 266534 6618
rect 269634 680494 270254 701760
rect 269634 680258 269666 680494
rect 269902 680258 269986 680494
rect 270222 680258 270254 680494
rect 269634 680174 270254 680258
rect 269634 679938 269666 680174
rect 269902 679938 269986 680174
rect 270222 679938 270254 680174
rect 269634 643294 270254 679938
rect 269634 643058 269666 643294
rect 269902 643058 269986 643294
rect 270222 643058 270254 643294
rect 269634 642974 270254 643058
rect 269634 642738 269666 642974
rect 269902 642738 269986 642974
rect 270222 642738 270254 642974
rect 269634 606094 270254 642738
rect 269634 605858 269666 606094
rect 269902 605858 269986 606094
rect 270222 605858 270254 606094
rect 269634 605774 270254 605858
rect 269634 605538 269666 605774
rect 269902 605538 269986 605774
rect 270222 605538 270254 605774
rect 269634 568894 270254 605538
rect 269634 568658 269666 568894
rect 269902 568658 269986 568894
rect 270222 568658 270254 568894
rect 269634 568574 270254 568658
rect 269634 568338 269666 568574
rect 269902 568338 269986 568574
rect 270222 568338 270254 568574
rect 269634 531694 270254 568338
rect 269634 531458 269666 531694
rect 269902 531458 269986 531694
rect 270222 531458 270254 531694
rect 269634 531374 270254 531458
rect 269634 531138 269666 531374
rect 269902 531138 269986 531374
rect 270222 531138 270254 531374
rect 269634 494494 270254 531138
rect 269634 494258 269666 494494
rect 269902 494258 269986 494494
rect 270222 494258 270254 494494
rect 269634 494174 270254 494258
rect 269634 493938 269666 494174
rect 269902 493938 269986 494174
rect 270222 493938 270254 494174
rect 269634 457294 270254 493938
rect 269634 457058 269666 457294
rect 269902 457058 269986 457294
rect 270222 457058 270254 457294
rect 269634 456974 270254 457058
rect 269634 456738 269666 456974
rect 269902 456738 269986 456974
rect 270222 456738 270254 456974
rect 269634 420094 270254 456738
rect 269634 419858 269666 420094
rect 269902 419858 269986 420094
rect 270222 419858 270254 420094
rect 269634 419774 270254 419858
rect 269634 419538 269666 419774
rect 269902 419538 269986 419774
rect 270222 419538 270254 419774
rect 269634 382894 270254 419538
rect 269634 382658 269666 382894
rect 269902 382658 269986 382894
rect 270222 382658 270254 382894
rect 269634 382574 270254 382658
rect 269634 382338 269666 382574
rect 269902 382338 269986 382574
rect 270222 382338 270254 382574
rect 269634 345694 270254 382338
rect 269634 345458 269666 345694
rect 269902 345458 269986 345694
rect 270222 345458 270254 345694
rect 269634 345374 270254 345458
rect 269634 345138 269666 345374
rect 269902 345138 269986 345374
rect 270222 345138 270254 345374
rect 269634 308494 270254 345138
rect 269634 308258 269666 308494
rect 269902 308258 269986 308494
rect 270222 308258 270254 308494
rect 269634 308174 270254 308258
rect 269634 307938 269666 308174
rect 269902 307938 269986 308174
rect 270222 307938 270254 308174
rect 269634 271294 270254 307938
rect 269634 271058 269666 271294
rect 269902 271058 269986 271294
rect 270222 271058 270254 271294
rect 269634 270974 270254 271058
rect 269634 270738 269666 270974
rect 269902 270738 269986 270974
rect 270222 270738 270254 270974
rect 269634 234094 270254 270738
rect 269634 233858 269666 234094
rect 269902 233858 269986 234094
rect 270222 233858 270254 234094
rect 269634 233774 270254 233858
rect 269634 233538 269666 233774
rect 269902 233538 269986 233774
rect 270222 233538 270254 233774
rect 269634 196894 270254 233538
rect 269634 196658 269666 196894
rect 269902 196658 269986 196894
rect 270222 196658 270254 196894
rect 269634 196574 270254 196658
rect 269634 196338 269666 196574
rect 269902 196338 269986 196574
rect 270222 196338 270254 196574
rect 269634 159694 270254 196338
rect 269634 159458 269666 159694
rect 269902 159458 269986 159694
rect 270222 159458 270254 159694
rect 269634 159374 270254 159458
rect 269634 159138 269666 159374
rect 269902 159138 269986 159374
rect 270222 159138 270254 159374
rect 269634 122494 270254 159138
rect 269634 122258 269666 122494
rect 269902 122258 269986 122494
rect 270222 122258 270254 122494
rect 269634 122174 270254 122258
rect 269634 121938 269666 122174
rect 269902 121938 269986 122174
rect 270222 121938 270254 122174
rect 269634 85294 270254 121938
rect 269634 85058 269666 85294
rect 269902 85058 269986 85294
rect 270222 85058 270254 85294
rect 269634 84974 270254 85058
rect 269634 84738 269666 84974
rect 269902 84738 269986 84974
rect 270222 84738 270254 84974
rect 269634 48094 270254 84738
rect 269634 47858 269666 48094
rect 269902 47858 269986 48094
rect 270222 47858 270254 48094
rect 269634 47774 270254 47858
rect 269634 47538 269666 47774
rect 269902 47538 269986 47774
rect 270222 47538 270254 47774
rect 269634 10894 270254 47538
rect 269634 10658 269666 10894
rect 269902 10658 269986 10894
rect 270222 10658 270254 10894
rect 269634 10574 270254 10658
rect 269634 10338 269666 10574
rect 269902 10338 269986 10574
rect 270222 10338 270254 10574
rect 269634 2176 270254 10338
rect 273354 684214 273974 701760
rect 273354 683978 273386 684214
rect 273622 683978 273706 684214
rect 273942 683978 273974 684214
rect 273354 683894 273974 683978
rect 273354 683658 273386 683894
rect 273622 683658 273706 683894
rect 273942 683658 273974 683894
rect 273354 647014 273974 683658
rect 273354 646778 273386 647014
rect 273622 646778 273706 647014
rect 273942 646778 273974 647014
rect 273354 646694 273974 646778
rect 273354 646458 273386 646694
rect 273622 646458 273706 646694
rect 273942 646458 273974 646694
rect 273354 609814 273974 646458
rect 273354 609578 273386 609814
rect 273622 609578 273706 609814
rect 273942 609578 273974 609814
rect 273354 609494 273974 609578
rect 273354 609258 273386 609494
rect 273622 609258 273706 609494
rect 273942 609258 273974 609494
rect 273354 572614 273974 609258
rect 273354 572378 273386 572614
rect 273622 572378 273706 572614
rect 273942 572378 273974 572614
rect 273354 572294 273974 572378
rect 273354 572058 273386 572294
rect 273622 572058 273706 572294
rect 273942 572058 273974 572294
rect 273354 535414 273974 572058
rect 273354 535178 273386 535414
rect 273622 535178 273706 535414
rect 273942 535178 273974 535414
rect 273354 535094 273974 535178
rect 273354 534858 273386 535094
rect 273622 534858 273706 535094
rect 273942 534858 273974 535094
rect 273354 498214 273974 534858
rect 273354 497978 273386 498214
rect 273622 497978 273706 498214
rect 273942 497978 273974 498214
rect 273354 497894 273974 497978
rect 273354 497658 273386 497894
rect 273622 497658 273706 497894
rect 273942 497658 273974 497894
rect 273354 461014 273974 497658
rect 273354 460778 273386 461014
rect 273622 460778 273706 461014
rect 273942 460778 273974 461014
rect 273354 460694 273974 460778
rect 273354 460458 273386 460694
rect 273622 460458 273706 460694
rect 273942 460458 273974 460694
rect 273354 423814 273974 460458
rect 273354 423578 273386 423814
rect 273622 423578 273706 423814
rect 273942 423578 273974 423814
rect 273354 423494 273974 423578
rect 273354 423258 273386 423494
rect 273622 423258 273706 423494
rect 273942 423258 273974 423494
rect 273354 386614 273974 423258
rect 273354 386378 273386 386614
rect 273622 386378 273706 386614
rect 273942 386378 273974 386614
rect 273354 386294 273974 386378
rect 273354 386058 273386 386294
rect 273622 386058 273706 386294
rect 273942 386058 273974 386294
rect 273354 349414 273974 386058
rect 273354 349178 273386 349414
rect 273622 349178 273706 349414
rect 273942 349178 273974 349414
rect 273354 349094 273974 349178
rect 273354 348858 273386 349094
rect 273622 348858 273706 349094
rect 273942 348858 273974 349094
rect 273354 312214 273974 348858
rect 273354 311978 273386 312214
rect 273622 311978 273706 312214
rect 273942 311978 273974 312214
rect 273354 311894 273974 311978
rect 273354 311658 273386 311894
rect 273622 311658 273706 311894
rect 273942 311658 273974 311894
rect 273354 275014 273974 311658
rect 273354 274778 273386 275014
rect 273622 274778 273706 275014
rect 273942 274778 273974 275014
rect 273354 274694 273974 274778
rect 273354 274458 273386 274694
rect 273622 274458 273706 274694
rect 273942 274458 273974 274694
rect 273354 237814 273974 274458
rect 273354 237578 273386 237814
rect 273622 237578 273706 237814
rect 273942 237578 273974 237814
rect 273354 237494 273974 237578
rect 273354 237258 273386 237494
rect 273622 237258 273706 237494
rect 273942 237258 273974 237494
rect 273354 200614 273974 237258
rect 273354 200378 273386 200614
rect 273622 200378 273706 200614
rect 273942 200378 273974 200614
rect 273354 200294 273974 200378
rect 273354 200058 273386 200294
rect 273622 200058 273706 200294
rect 273942 200058 273974 200294
rect 273354 163414 273974 200058
rect 273354 163178 273386 163414
rect 273622 163178 273706 163414
rect 273942 163178 273974 163414
rect 273354 163094 273974 163178
rect 273354 162858 273386 163094
rect 273622 162858 273706 163094
rect 273942 162858 273974 163094
rect 273354 126214 273974 162858
rect 273354 125978 273386 126214
rect 273622 125978 273706 126214
rect 273942 125978 273974 126214
rect 273354 125894 273974 125978
rect 273354 125658 273386 125894
rect 273622 125658 273706 125894
rect 273942 125658 273974 125894
rect 273354 89014 273974 125658
rect 273354 88778 273386 89014
rect 273622 88778 273706 89014
rect 273942 88778 273974 89014
rect 273354 88694 273974 88778
rect 273354 88458 273386 88694
rect 273622 88458 273706 88694
rect 273942 88458 273974 88694
rect 273354 51814 273974 88458
rect 273354 51578 273386 51814
rect 273622 51578 273706 51814
rect 273942 51578 273974 51814
rect 273354 51494 273974 51578
rect 273354 51258 273386 51494
rect 273622 51258 273706 51494
rect 273942 51258 273974 51494
rect 273354 14614 273974 51258
rect 273354 14378 273386 14614
rect 273622 14378 273706 14614
rect 273942 14378 273974 14614
rect 273354 14294 273974 14378
rect 273354 14058 273386 14294
rect 273622 14058 273706 14294
rect 273942 14058 273974 14294
rect 273354 2176 273974 14058
rect 277074 687934 277694 701760
rect 277074 687698 277106 687934
rect 277342 687698 277426 687934
rect 277662 687698 277694 687934
rect 277074 687614 277694 687698
rect 277074 687378 277106 687614
rect 277342 687378 277426 687614
rect 277662 687378 277694 687614
rect 277074 650734 277694 687378
rect 277074 650498 277106 650734
rect 277342 650498 277426 650734
rect 277662 650498 277694 650734
rect 277074 650414 277694 650498
rect 277074 650178 277106 650414
rect 277342 650178 277426 650414
rect 277662 650178 277694 650414
rect 277074 613534 277694 650178
rect 277074 613298 277106 613534
rect 277342 613298 277426 613534
rect 277662 613298 277694 613534
rect 277074 613214 277694 613298
rect 277074 612978 277106 613214
rect 277342 612978 277426 613214
rect 277662 612978 277694 613214
rect 277074 576334 277694 612978
rect 277074 576098 277106 576334
rect 277342 576098 277426 576334
rect 277662 576098 277694 576334
rect 277074 576014 277694 576098
rect 277074 575778 277106 576014
rect 277342 575778 277426 576014
rect 277662 575778 277694 576014
rect 277074 539134 277694 575778
rect 277074 538898 277106 539134
rect 277342 538898 277426 539134
rect 277662 538898 277694 539134
rect 277074 538814 277694 538898
rect 277074 538578 277106 538814
rect 277342 538578 277426 538814
rect 277662 538578 277694 538814
rect 277074 501934 277694 538578
rect 277074 501698 277106 501934
rect 277342 501698 277426 501934
rect 277662 501698 277694 501934
rect 277074 501614 277694 501698
rect 277074 501378 277106 501614
rect 277342 501378 277426 501614
rect 277662 501378 277694 501614
rect 277074 464734 277694 501378
rect 277074 464498 277106 464734
rect 277342 464498 277426 464734
rect 277662 464498 277694 464734
rect 277074 464414 277694 464498
rect 277074 464178 277106 464414
rect 277342 464178 277426 464414
rect 277662 464178 277694 464414
rect 277074 427534 277694 464178
rect 277074 427298 277106 427534
rect 277342 427298 277426 427534
rect 277662 427298 277694 427534
rect 277074 427214 277694 427298
rect 277074 426978 277106 427214
rect 277342 426978 277426 427214
rect 277662 426978 277694 427214
rect 277074 390334 277694 426978
rect 277074 390098 277106 390334
rect 277342 390098 277426 390334
rect 277662 390098 277694 390334
rect 277074 390014 277694 390098
rect 277074 389778 277106 390014
rect 277342 389778 277426 390014
rect 277662 389778 277694 390014
rect 277074 353134 277694 389778
rect 277074 352898 277106 353134
rect 277342 352898 277426 353134
rect 277662 352898 277694 353134
rect 277074 352814 277694 352898
rect 277074 352578 277106 352814
rect 277342 352578 277426 352814
rect 277662 352578 277694 352814
rect 277074 315934 277694 352578
rect 277074 315698 277106 315934
rect 277342 315698 277426 315934
rect 277662 315698 277694 315934
rect 277074 315614 277694 315698
rect 277074 315378 277106 315614
rect 277342 315378 277426 315614
rect 277662 315378 277694 315614
rect 277074 278734 277694 315378
rect 277074 278498 277106 278734
rect 277342 278498 277426 278734
rect 277662 278498 277694 278734
rect 277074 278414 277694 278498
rect 277074 278178 277106 278414
rect 277342 278178 277426 278414
rect 277662 278178 277694 278414
rect 277074 241534 277694 278178
rect 277074 241298 277106 241534
rect 277342 241298 277426 241534
rect 277662 241298 277694 241534
rect 277074 241214 277694 241298
rect 277074 240978 277106 241214
rect 277342 240978 277426 241214
rect 277662 240978 277694 241214
rect 277074 204334 277694 240978
rect 277074 204098 277106 204334
rect 277342 204098 277426 204334
rect 277662 204098 277694 204334
rect 277074 204014 277694 204098
rect 277074 203778 277106 204014
rect 277342 203778 277426 204014
rect 277662 203778 277694 204014
rect 277074 167134 277694 203778
rect 277074 166898 277106 167134
rect 277342 166898 277426 167134
rect 277662 166898 277694 167134
rect 277074 166814 277694 166898
rect 277074 166578 277106 166814
rect 277342 166578 277426 166814
rect 277662 166578 277694 166814
rect 277074 129934 277694 166578
rect 277074 129698 277106 129934
rect 277342 129698 277426 129934
rect 277662 129698 277694 129934
rect 277074 129614 277694 129698
rect 277074 129378 277106 129614
rect 277342 129378 277426 129614
rect 277662 129378 277694 129614
rect 277074 92734 277694 129378
rect 277074 92498 277106 92734
rect 277342 92498 277426 92734
rect 277662 92498 277694 92734
rect 277074 92414 277694 92498
rect 277074 92178 277106 92414
rect 277342 92178 277426 92414
rect 277662 92178 277694 92414
rect 277074 55534 277694 92178
rect 277074 55298 277106 55534
rect 277342 55298 277426 55534
rect 277662 55298 277694 55534
rect 277074 55214 277694 55298
rect 277074 54978 277106 55214
rect 277342 54978 277426 55214
rect 277662 54978 277694 55214
rect 277074 18334 277694 54978
rect 277074 18098 277106 18334
rect 277342 18098 277426 18334
rect 277662 18098 277694 18334
rect 277074 18014 277694 18098
rect 277074 17778 277106 18014
rect 277342 17778 277426 18014
rect 277662 17778 277694 18014
rect 277074 2176 277694 17778
rect 280794 691654 281414 701760
rect 280794 691418 280826 691654
rect 281062 691418 281146 691654
rect 281382 691418 281414 691654
rect 280794 691334 281414 691418
rect 280794 691098 280826 691334
rect 281062 691098 281146 691334
rect 281382 691098 281414 691334
rect 280794 654454 281414 691098
rect 280794 654218 280826 654454
rect 281062 654218 281146 654454
rect 281382 654218 281414 654454
rect 280794 654134 281414 654218
rect 280794 653898 280826 654134
rect 281062 653898 281146 654134
rect 281382 653898 281414 654134
rect 280794 617254 281414 653898
rect 280794 617018 280826 617254
rect 281062 617018 281146 617254
rect 281382 617018 281414 617254
rect 280794 616934 281414 617018
rect 280794 616698 280826 616934
rect 281062 616698 281146 616934
rect 281382 616698 281414 616934
rect 280794 580054 281414 616698
rect 280794 579818 280826 580054
rect 281062 579818 281146 580054
rect 281382 579818 281414 580054
rect 280794 579734 281414 579818
rect 280794 579498 280826 579734
rect 281062 579498 281146 579734
rect 281382 579498 281414 579734
rect 280794 542854 281414 579498
rect 280794 542618 280826 542854
rect 281062 542618 281146 542854
rect 281382 542618 281414 542854
rect 280794 542534 281414 542618
rect 280794 542298 280826 542534
rect 281062 542298 281146 542534
rect 281382 542298 281414 542534
rect 280794 505654 281414 542298
rect 280794 505418 280826 505654
rect 281062 505418 281146 505654
rect 281382 505418 281414 505654
rect 280794 505334 281414 505418
rect 280794 505098 280826 505334
rect 281062 505098 281146 505334
rect 281382 505098 281414 505334
rect 280794 468454 281414 505098
rect 280794 468218 280826 468454
rect 281062 468218 281146 468454
rect 281382 468218 281414 468454
rect 280794 468134 281414 468218
rect 280794 467898 280826 468134
rect 281062 467898 281146 468134
rect 281382 467898 281414 468134
rect 280794 431254 281414 467898
rect 280794 431018 280826 431254
rect 281062 431018 281146 431254
rect 281382 431018 281414 431254
rect 280794 430934 281414 431018
rect 280794 430698 280826 430934
rect 281062 430698 281146 430934
rect 281382 430698 281414 430934
rect 280794 394054 281414 430698
rect 280794 393818 280826 394054
rect 281062 393818 281146 394054
rect 281382 393818 281414 394054
rect 280794 393734 281414 393818
rect 280794 393498 280826 393734
rect 281062 393498 281146 393734
rect 281382 393498 281414 393734
rect 280794 356854 281414 393498
rect 280794 356618 280826 356854
rect 281062 356618 281146 356854
rect 281382 356618 281414 356854
rect 280794 356534 281414 356618
rect 280794 356298 280826 356534
rect 281062 356298 281146 356534
rect 281382 356298 281414 356534
rect 280794 319654 281414 356298
rect 280794 319418 280826 319654
rect 281062 319418 281146 319654
rect 281382 319418 281414 319654
rect 280794 319334 281414 319418
rect 280794 319098 280826 319334
rect 281062 319098 281146 319334
rect 281382 319098 281414 319334
rect 280794 282454 281414 319098
rect 280794 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 281414 282454
rect 280794 282134 281414 282218
rect 280794 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 281414 282134
rect 280794 245254 281414 281898
rect 280794 245018 280826 245254
rect 281062 245018 281146 245254
rect 281382 245018 281414 245254
rect 280794 244934 281414 245018
rect 280794 244698 280826 244934
rect 281062 244698 281146 244934
rect 281382 244698 281414 244934
rect 280794 208054 281414 244698
rect 280794 207818 280826 208054
rect 281062 207818 281146 208054
rect 281382 207818 281414 208054
rect 280794 207734 281414 207818
rect 280794 207498 280826 207734
rect 281062 207498 281146 207734
rect 281382 207498 281414 207734
rect 280794 170854 281414 207498
rect 280794 170618 280826 170854
rect 281062 170618 281146 170854
rect 281382 170618 281414 170854
rect 280794 170534 281414 170618
rect 280794 170298 280826 170534
rect 281062 170298 281146 170534
rect 281382 170298 281414 170534
rect 280794 133654 281414 170298
rect 280794 133418 280826 133654
rect 281062 133418 281146 133654
rect 281382 133418 281414 133654
rect 280794 133334 281414 133418
rect 280794 133098 280826 133334
rect 281062 133098 281146 133334
rect 281382 133098 281414 133334
rect 280794 96454 281414 133098
rect 280794 96218 280826 96454
rect 281062 96218 281146 96454
rect 281382 96218 281414 96454
rect 280794 96134 281414 96218
rect 280794 95898 280826 96134
rect 281062 95898 281146 96134
rect 281382 95898 281414 96134
rect 280794 59254 281414 95898
rect 280794 59018 280826 59254
rect 281062 59018 281146 59254
rect 281382 59018 281414 59254
rect 280794 58934 281414 59018
rect 280794 58698 280826 58934
rect 281062 58698 281146 58934
rect 281382 58698 281414 58934
rect 280794 22054 281414 58698
rect 280794 21818 280826 22054
rect 281062 21818 281146 22054
rect 281382 21818 281414 22054
rect 280794 21734 281414 21818
rect 280794 21498 280826 21734
rect 281062 21498 281146 21734
rect 281382 21498 281414 21734
rect 280794 2176 281414 21498
rect 284514 695374 285134 701760
rect 284514 695138 284546 695374
rect 284782 695138 284866 695374
rect 285102 695138 285134 695374
rect 284514 695054 285134 695138
rect 284514 694818 284546 695054
rect 284782 694818 284866 695054
rect 285102 694818 285134 695054
rect 284514 658174 285134 694818
rect 284514 657938 284546 658174
rect 284782 657938 284866 658174
rect 285102 657938 285134 658174
rect 284514 657854 285134 657938
rect 284514 657618 284546 657854
rect 284782 657618 284866 657854
rect 285102 657618 285134 657854
rect 284514 620974 285134 657618
rect 284514 620738 284546 620974
rect 284782 620738 284866 620974
rect 285102 620738 285134 620974
rect 284514 620654 285134 620738
rect 284514 620418 284546 620654
rect 284782 620418 284866 620654
rect 285102 620418 285134 620654
rect 284514 583774 285134 620418
rect 284514 583538 284546 583774
rect 284782 583538 284866 583774
rect 285102 583538 285134 583774
rect 284514 583454 285134 583538
rect 284514 583218 284546 583454
rect 284782 583218 284866 583454
rect 285102 583218 285134 583454
rect 284514 546574 285134 583218
rect 284514 546338 284546 546574
rect 284782 546338 284866 546574
rect 285102 546338 285134 546574
rect 284514 546254 285134 546338
rect 284514 546018 284546 546254
rect 284782 546018 284866 546254
rect 285102 546018 285134 546254
rect 284514 509374 285134 546018
rect 284514 509138 284546 509374
rect 284782 509138 284866 509374
rect 285102 509138 285134 509374
rect 284514 509054 285134 509138
rect 284514 508818 284546 509054
rect 284782 508818 284866 509054
rect 285102 508818 285134 509054
rect 284514 472174 285134 508818
rect 284514 471938 284546 472174
rect 284782 471938 284866 472174
rect 285102 471938 285134 472174
rect 284514 471854 285134 471938
rect 284514 471618 284546 471854
rect 284782 471618 284866 471854
rect 285102 471618 285134 471854
rect 284514 434974 285134 471618
rect 284514 434738 284546 434974
rect 284782 434738 284866 434974
rect 285102 434738 285134 434974
rect 284514 434654 285134 434738
rect 284514 434418 284546 434654
rect 284782 434418 284866 434654
rect 285102 434418 285134 434654
rect 284514 397774 285134 434418
rect 284514 397538 284546 397774
rect 284782 397538 284866 397774
rect 285102 397538 285134 397774
rect 284514 397454 285134 397538
rect 284514 397218 284546 397454
rect 284782 397218 284866 397454
rect 285102 397218 285134 397454
rect 284514 360574 285134 397218
rect 284514 360338 284546 360574
rect 284782 360338 284866 360574
rect 285102 360338 285134 360574
rect 284514 360254 285134 360338
rect 284514 360018 284546 360254
rect 284782 360018 284866 360254
rect 285102 360018 285134 360254
rect 284514 323374 285134 360018
rect 284514 323138 284546 323374
rect 284782 323138 284866 323374
rect 285102 323138 285134 323374
rect 284514 323054 285134 323138
rect 284514 322818 284546 323054
rect 284782 322818 284866 323054
rect 285102 322818 285134 323054
rect 284514 286174 285134 322818
rect 284514 285938 284546 286174
rect 284782 285938 284866 286174
rect 285102 285938 285134 286174
rect 284514 285854 285134 285938
rect 284514 285618 284546 285854
rect 284782 285618 284866 285854
rect 285102 285618 285134 285854
rect 284514 248974 285134 285618
rect 284514 248738 284546 248974
rect 284782 248738 284866 248974
rect 285102 248738 285134 248974
rect 284514 248654 285134 248738
rect 284514 248418 284546 248654
rect 284782 248418 284866 248654
rect 285102 248418 285134 248654
rect 284514 211774 285134 248418
rect 284514 211538 284546 211774
rect 284782 211538 284866 211774
rect 285102 211538 285134 211774
rect 284514 211454 285134 211538
rect 284514 211218 284546 211454
rect 284782 211218 284866 211454
rect 285102 211218 285134 211454
rect 284514 174574 285134 211218
rect 284514 174338 284546 174574
rect 284782 174338 284866 174574
rect 285102 174338 285134 174574
rect 284514 174254 285134 174338
rect 284514 174018 284546 174254
rect 284782 174018 284866 174254
rect 285102 174018 285134 174254
rect 284514 137374 285134 174018
rect 284514 137138 284546 137374
rect 284782 137138 284866 137374
rect 285102 137138 285134 137374
rect 284514 137054 285134 137138
rect 284514 136818 284546 137054
rect 284782 136818 284866 137054
rect 285102 136818 285134 137054
rect 284514 100174 285134 136818
rect 284514 99938 284546 100174
rect 284782 99938 284866 100174
rect 285102 99938 285134 100174
rect 284514 99854 285134 99938
rect 284514 99618 284546 99854
rect 284782 99618 284866 99854
rect 285102 99618 285134 99854
rect 284514 62974 285134 99618
rect 284514 62738 284546 62974
rect 284782 62738 284866 62974
rect 285102 62738 285134 62974
rect 284514 62654 285134 62738
rect 284514 62418 284546 62654
rect 284782 62418 284866 62654
rect 285102 62418 285134 62654
rect 284514 25774 285134 62418
rect 284514 25538 284546 25774
rect 284782 25538 284866 25774
rect 285102 25538 285134 25774
rect 284514 25454 285134 25538
rect 284514 25218 284546 25454
rect 284782 25218 284866 25454
rect 285102 25218 285134 25454
rect 284514 2176 285134 25218
rect 288234 699094 288854 701760
rect 288234 698858 288266 699094
rect 288502 698858 288586 699094
rect 288822 698858 288854 699094
rect 288234 698774 288854 698858
rect 288234 698538 288266 698774
rect 288502 698538 288586 698774
rect 288822 698538 288854 698774
rect 288234 661894 288854 698538
rect 288234 661658 288266 661894
rect 288502 661658 288586 661894
rect 288822 661658 288854 661894
rect 288234 661574 288854 661658
rect 288234 661338 288266 661574
rect 288502 661338 288586 661574
rect 288822 661338 288854 661574
rect 288234 624694 288854 661338
rect 288234 624458 288266 624694
rect 288502 624458 288586 624694
rect 288822 624458 288854 624694
rect 288234 624374 288854 624458
rect 288234 624138 288266 624374
rect 288502 624138 288586 624374
rect 288822 624138 288854 624374
rect 288234 587494 288854 624138
rect 288234 587258 288266 587494
rect 288502 587258 288586 587494
rect 288822 587258 288854 587494
rect 288234 587174 288854 587258
rect 288234 586938 288266 587174
rect 288502 586938 288586 587174
rect 288822 586938 288854 587174
rect 288234 550294 288854 586938
rect 288234 550058 288266 550294
rect 288502 550058 288586 550294
rect 288822 550058 288854 550294
rect 288234 549974 288854 550058
rect 288234 549738 288266 549974
rect 288502 549738 288586 549974
rect 288822 549738 288854 549974
rect 288234 513094 288854 549738
rect 288234 512858 288266 513094
rect 288502 512858 288586 513094
rect 288822 512858 288854 513094
rect 288234 512774 288854 512858
rect 288234 512538 288266 512774
rect 288502 512538 288586 512774
rect 288822 512538 288854 512774
rect 288234 475894 288854 512538
rect 288234 475658 288266 475894
rect 288502 475658 288586 475894
rect 288822 475658 288854 475894
rect 288234 475574 288854 475658
rect 288234 475338 288266 475574
rect 288502 475338 288586 475574
rect 288822 475338 288854 475574
rect 288234 438694 288854 475338
rect 288234 438458 288266 438694
rect 288502 438458 288586 438694
rect 288822 438458 288854 438694
rect 288234 438374 288854 438458
rect 288234 438138 288266 438374
rect 288502 438138 288586 438374
rect 288822 438138 288854 438374
rect 288234 401494 288854 438138
rect 288234 401258 288266 401494
rect 288502 401258 288586 401494
rect 288822 401258 288854 401494
rect 288234 401174 288854 401258
rect 288234 400938 288266 401174
rect 288502 400938 288586 401174
rect 288822 400938 288854 401174
rect 288234 364294 288854 400938
rect 288234 364058 288266 364294
rect 288502 364058 288586 364294
rect 288822 364058 288854 364294
rect 288234 363974 288854 364058
rect 288234 363738 288266 363974
rect 288502 363738 288586 363974
rect 288822 363738 288854 363974
rect 288234 327094 288854 363738
rect 288234 326858 288266 327094
rect 288502 326858 288586 327094
rect 288822 326858 288854 327094
rect 288234 326774 288854 326858
rect 288234 326538 288266 326774
rect 288502 326538 288586 326774
rect 288822 326538 288854 326774
rect 288234 289894 288854 326538
rect 288234 289658 288266 289894
rect 288502 289658 288586 289894
rect 288822 289658 288854 289894
rect 288234 289574 288854 289658
rect 288234 289338 288266 289574
rect 288502 289338 288586 289574
rect 288822 289338 288854 289574
rect 288234 252694 288854 289338
rect 288234 252458 288266 252694
rect 288502 252458 288586 252694
rect 288822 252458 288854 252694
rect 288234 252374 288854 252458
rect 288234 252138 288266 252374
rect 288502 252138 288586 252374
rect 288822 252138 288854 252374
rect 288234 215494 288854 252138
rect 288234 215258 288266 215494
rect 288502 215258 288586 215494
rect 288822 215258 288854 215494
rect 288234 215174 288854 215258
rect 288234 214938 288266 215174
rect 288502 214938 288586 215174
rect 288822 214938 288854 215174
rect 288234 178294 288854 214938
rect 288234 178058 288266 178294
rect 288502 178058 288586 178294
rect 288822 178058 288854 178294
rect 288234 177974 288854 178058
rect 288234 177738 288266 177974
rect 288502 177738 288586 177974
rect 288822 177738 288854 177974
rect 288234 141094 288854 177738
rect 288234 140858 288266 141094
rect 288502 140858 288586 141094
rect 288822 140858 288854 141094
rect 288234 140774 288854 140858
rect 288234 140538 288266 140774
rect 288502 140538 288586 140774
rect 288822 140538 288854 140774
rect 288234 103894 288854 140538
rect 288234 103658 288266 103894
rect 288502 103658 288586 103894
rect 288822 103658 288854 103894
rect 288234 103574 288854 103658
rect 288234 103338 288266 103574
rect 288502 103338 288586 103574
rect 288822 103338 288854 103574
rect 288234 66694 288854 103338
rect 288234 66458 288266 66694
rect 288502 66458 288586 66694
rect 288822 66458 288854 66694
rect 288234 66374 288854 66458
rect 288234 66138 288266 66374
rect 288502 66138 288586 66374
rect 288822 66138 288854 66374
rect 288234 29494 288854 66138
rect 288234 29258 288266 29494
rect 288502 29258 288586 29494
rect 288822 29258 288854 29494
rect 288234 29174 288854 29258
rect 288234 28938 288266 29174
rect 288502 28938 288586 29174
rect 288822 28938 288854 29174
rect 288234 2176 288854 28938
rect 299394 673054 300014 701760
rect 299394 672818 299426 673054
rect 299662 672818 299746 673054
rect 299982 672818 300014 673054
rect 299394 672734 300014 672818
rect 299394 672498 299426 672734
rect 299662 672498 299746 672734
rect 299982 672498 300014 672734
rect 299394 635854 300014 672498
rect 299394 635618 299426 635854
rect 299662 635618 299746 635854
rect 299982 635618 300014 635854
rect 299394 635534 300014 635618
rect 299394 635298 299426 635534
rect 299662 635298 299746 635534
rect 299982 635298 300014 635534
rect 299394 598654 300014 635298
rect 299394 598418 299426 598654
rect 299662 598418 299746 598654
rect 299982 598418 300014 598654
rect 299394 598334 300014 598418
rect 299394 598098 299426 598334
rect 299662 598098 299746 598334
rect 299982 598098 300014 598334
rect 299394 561454 300014 598098
rect 299394 561218 299426 561454
rect 299662 561218 299746 561454
rect 299982 561218 300014 561454
rect 299394 561134 300014 561218
rect 299394 560898 299426 561134
rect 299662 560898 299746 561134
rect 299982 560898 300014 561134
rect 299394 524254 300014 560898
rect 299394 524018 299426 524254
rect 299662 524018 299746 524254
rect 299982 524018 300014 524254
rect 299394 523934 300014 524018
rect 299394 523698 299426 523934
rect 299662 523698 299746 523934
rect 299982 523698 300014 523934
rect 299394 487054 300014 523698
rect 299394 486818 299426 487054
rect 299662 486818 299746 487054
rect 299982 486818 300014 487054
rect 299394 486734 300014 486818
rect 299394 486498 299426 486734
rect 299662 486498 299746 486734
rect 299982 486498 300014 486734
rect 299394 449854 300014 486498
rect 299394 449618 299426 449854
rect 299662 449618 299746 449854
rect 299982 449618 300014 449854
rect 299394 449534 300014 449618
rect 299394 449298 299426 449534
rect 299662 449298 299746 449534
rect 299982 449298 300014 449534
rect 299394 412654 300014 449298
rect 299394 412418 299426 412654
rect 299662 412418 299746 412654
rect 299982 412418 300014 412654
rect 299394 412334 300014 412418
rect 299394 412098 299426 412334
rect 299662 412098 299746 412334
rect 299982 412098 300014 412334
rect 299394 375454 300014 412098
rect 299394 375218 299426 375454
rect 299662 375218 299746 375454
rect 299982 375218 300014 375454
rect 299394 375134 300014 375218
rect 299394 374898 299426 375134
rect 299662 374898 299746 375134
rect 299982 374898 300014 375134
rect 299394 338254 300014 374898
rect 299394 338018 299426 338254
rect 299662 338018 299746 338254
rect 299982 338018 300014 338254
rect 299394 337934 300014 338018
rect 299394 337698 299426 337934
rect 299662 337698 299746 337934
rect 299982 337698 300014 337934
rect 299394 301054 300014 337698
rect 299394 300818 299426 301054
rect 299662 300818 299746 301054
rect 299982 300818 300014 301054
rect 299394 300734 300014 300818
rect 299394 300498 299426 300734
rect 299662 300498 299746 300734
rect 299982 300498 300014 300734
rect 299394 263854 300014 300498
rect 299394 263618 299426 263854
rect 299662 263618 299746 263854
rect 299982 263618 300014 263854
rect 299394 263534 300014 263618
rect 299394 263298 299426 263534
rect 299662 263298 299746 263534
rect 299982 263298 300014 263534
rect 299394 226654 300014 263298
rect 299394 226418 299426 226654
rect 299662 226418 299746 226654
rect 299982 226418 300014 226654
rect 299394 226334 300014 226418
rect 299394 226098 299426 226334
rect 299662 226098 299746 226334
rect 299982 226098 300014 226334
rect 299394 189454 300014 226098
rect 299394 189218 299426 189454
rect 299662 189218 299746 189454
rect 299982 189218 300014 189454
rect 299394 189134 300014 189218
rect 299394 188898 299426 189134
rect 299662 188898 299746 189134
rect 299982 188898 300014 189134
rect 299394 152254 300014 188898
rect 299394 152018 299426 152254
rect 299662 152018 299746 152254
rect 299982 152018 300014 152254
rect 299394 151934 300014 152018
rect 299394 151698 299426 151934
rect 299662 151698 299746 151934
rect 299982 151698 300014 151934
rect 299394 115054 300014 151698
rect 299394 114818 299426 115054
rect 299662 114818 299746 115054
rect 299982 114818 300014 115054
rect 299394 114734 300014 114818
rect 299394 114498 299426 114734
rect 299662 114498 299746 114734
rect 299982 114498 300014 114734
rect 299394 77854 300014 114498
rect 299394 77618 299426 77854
rect 299662 77618 299746 77854
rect 299982 77618 300014 77854
rect 299394 77534 300014 77618
rect 299394 77298 299426 77534
rect 299662 77298 299746 77534
rect 299982 77298 300014 77534
rect 299394 40654 300014 77298
rect 299394 40418 299426 40654
rect 299662 40418 299746 40654
rect 299982 40418 300014 40654
rect 299394 40334 300014 40418
rect 299394 40098 299426 40334
rect 299662 40098 299746 40334
rect 299982 40098 300014 40334
rect 299394 3454 300014 40098
rect 299394 3218 299426 3454
rect 299662 3218 299746 3454
rect 299982 3218 300014 3454
rect 299394 3134 300014 3218
rect 299394 2898 299426 3134
rect 299662 2898 299746 3134
rect 299982 2898 300014 3134
rect 299394 2176 300014 2898
rect 303114 676774 303734 701760
rect 303114 676538 303146 676774
rect 303382 676538 303466 676774
rect 303702 676538 303734 676774
rect 303114 676454 303734 676538
rect 303114 676218 303146 676454
rect 303382 676218 303466 676454
rect 303702 676218 303734 676454
rect 303114 639574 303734 676218
rect 303114 639338 303146 639574
rect 303382 639338 303466 639574
rect 303702 639338 303734 639574
rect 303114 639254 303734 639338
rect 303114 639018 303146 639254
rect 303382 639018 303466 639254
rect 303702 639018 303734 639254
rect 303114 602374 303734 639018
rect 303114 602138 303146 602374
rect 303382 602138 303466 602374
rect 303702 602138 303734 602374
rect 303114 602054 303734 602138
rect 303114 601818 303146 602054
rect 303382 601818 303466 602054
rect 303702 601818 303734 602054
rect 303114 565174 303734 601818
rect 303114 564938 303146 565174
rect 303382 564938 303466 565174
rect 303702 564938 303734 565174
rect 303114 564854 303734 564938
rect 303114 564618 303146 564854
rect 303382 564618 303466 564854
rect 303702 564618 303734 564854
rect 303114 527974 303734 564618
rect 303114 527738 303146 527974
rect 303382 527738 303466 527974
rect 303702 527738 303734 527974
rect 303114 527654 303734 527738
rect 303114 527418 303146 527654
rect 303382 527418 303466 527654
rect 303702 527418 303734 527654
rect 303114 490774 303734 527418
rect 303114 490538 303146 490774
rect 303382 490538 303466 490774
rect 303702 490538 303734 490774
rect 303114 490454 303734 490538
rect 303114 490218 303146 490454
rect 303382 490218 303466 490454
rect 303702 490218 303734 490454
rect 303114 453574 303734 490218
rect 303114 453338 303146 453574
rect 303382 453338 303466 453574
rect 303702 453338 303734 453574
rect 303114 453254 303734 453338
rect 303114 453018 303146 453254
rect 303382 453018 303466 453254
rect 303702 453018 303734 453254
rect 303114 416374 303734 453018
rect 303114 416138 303146 416374
rect 303382 416138 303466 416374
rect 303702 416138 303734 416374
rect 303114 416054 303734 416138
rect 303114 415818 303146 416054
rect 303382 415818 303466 416054
rect 303702 415818 303734 416054
rect 303114 379174 303734 415818
rect 303114 378938 303146 379174
rect 303382 378938 303466 379174
rect 303702 378938 303734 379174
rect 303114 378854 303734 378938
rect 303114 378618 303146 378854
rect 303382 378618 303466 378854
rect 303702 378618 303734 378854
rect 303114 341974 303734 378618
rect 303114 341738 303146 341974
rect 303382 341738 303466 341974
rect 303702 341738 303734 341974
rect 303114 341654 303734 341738
rect 303114 341418 303146 341654
rect 303382 341418 303466 341654
rect 303702 341418 303734 341654
rect 303114 304774 303734 341418
rect 303114 304538 303146 304774
rect 303382 304538 303466 304774
rect 303702 304538 303734 304774
rect 303114 304454 303734 304538
rect 303114 304218 303146 304454
rect 303382 304218 303466 304454
rect 303702 304218 303734 304454
rect 303114 267574 303734 304218
rect 303114 267338 303146 267574
rect 303382 267338 303466 267574
rect 303702 267338 303734 267574
rect 303114 267254 303734 267338
rect 303114 267018 303146 267254
rect 303382 267018 303466 267254
rect 303702 267018 303734 267254
rect 303114 230374 303734 267018
rect 303114 230138 303146 230374
rect 303382 230138 303466 230374
rect 303702 230138 303734 230374
rect 303114 230054 303734 230138
rect 303114 229818 303146 230054
rect 303382 229818 303466 230054
rect 303702 229818 303734 230054
rect 303114 193174 303734 229818
rect 303114 192938 303146 193174
rect 303382 192938 303466 193174
rect 303702 192938 303734 193174
rect 303114 192854 303734 192938
rect 303114 192618 303146 192854
rect 303382 192618 303466 192854
rect 303702 192618 303734 192854
rect 303114 155974 303734 192618
rect 303114 155738 303146 155974
rect 303382 155738 303466 155974
rect 303702 155738 303734 155974
rect 303114 155654 303734 155738
rect 303114 155418 303146 155654
rect 303382 155418 303466 155654
rect 303702 155418 303734 155654
rect 303114 118774 303734 155418
rect 303114 118538 303146 118774
rect 303382 118538 303466 118774
rect 303702 118538 303734 118774
rect 303114 118454 303734 118538
rect 303114 118218 303146 118454
rect 303382 118218 303466 118454
rect 303702 118218 303734 118454
rect 303114 81574 303734 118218
rect 303114 81338 303146 81574
rect 303382 81338 303466 81574
rect 303702 81338 303734 81574
rect 303114 81254 303734 81338
rect 303114 81018 303146 81254
rect 303382 81018 303466 81254
rect 303702 81018 303734 81254
rect 303114 44374 303734 81018
rect 303114 44138 303146 44374
rect 303382 44138 303466 44374
rect 303702 44138 303734 44374
rect 303114 44054 303734 44138
rect 303114 43818 303146 44054
rect 303382 43818 303466 44054
rect 303702 43818 303734 44054
rect 303114 7174 303734 43818
rect 303114 6938 303146 7174
rect 303382 6938 303466 7174
rect 303702 6938 303734 7174
rect 303114 6854 303734 6938
rect 303114 6618 303146 6854
rect 303382 6618 303466 6854
rect 303702 6618 303734 6854
rect 303114 2176 303734 6618
rect 306834 680494 307454 701760
rect 306834 680258 306866 680494
rect 307102 680258 307186 680494
rect 307422 680258 307454 680494
rect 306834 680174 307454 680258
rect 306834 679938 306866 680174
rect 307102 679938 307186 680174
rect 307422 679938 307454 680174
rect 306834 643294 307454 679938
rect 306834 643058 306866 643294
rect 307102 643058 307186 643294
rect 307422 643058 307454 643294
rect 306834 642974 307454 643058
rect 306834 642738 306866 642974
rect 307102 642738 307186 642974
rect 307422 642738 307454 642974
rect 306834 606094 307454 642738
rect 306834 605858 306866 606094
rect 307102 605858 307186 606094
rect 307422 605858 307454 606094
rect 306834 605774 307454 605858
rect 306834 605538 306866 605774
rect 307102 605538 307186 605774
rect 307422 605538 307454 605774
rect 306834 568894 307454 605538
rect 306834 568658 306866 568894
rect 307102 568658 307186 568894
rect 307422 568658 307454 568894
rect 306834 568574 307454 568658
rect 306834 568338 306866 568574
rect 307102 568338 307186 568574
rect 307422 568338 307454 568574
rect 306834 531694 307454 568338
rect 306834 531458 306866 531694
rect 307102 531458 307186 531694
rect 307422 531458 307454 531694
rect 306834 531374 307454 531458
rect 306834 531138 306866 531374
rect 307102 531138 307186 531374
rect 307422 531138 307454 531374
rect 306834 494494 307454 531138
rect 306834 494258 306866 494494
rect 307102 494258 307186 494494
rect 307422 494258 307454 494494
rect 306834 494174 307454 494258
rect 306834 493938 306866 494174
rect 307102 493938 307186 494174
rect 307422 493938 307454 494174
rect 306834 457294 307454 493938
rect 306834 457058 306866 457294
rect 307102 457058 307186 457294
rect 307422 457058 307454 457294
rect 306834 456974 307454 457058
rect 306834 456738 306866 456974
rect 307102 456738 307186 456974
rect 307422 456738 307454 456974
rect 306834 420094 307454 456738
rect 306834 419858 306866 420094
rect 307102 419858 307186 420094
rect 307422 419858 307454 420094
rect 306834 419774 307454 419858
rect 306834 419538 306866 419774
rect 307102 419538 307186 419774
rect 307422 419538 307454 419774
rect 306834 382894 307454 419538
rect 306834 382658 306866 382894
rect 307102 382658 307186 382894
rect 307422 382658 307454 382894
rect 306834 382574 307454 382658
rect 306834 382338 306866 382574
rect 307102 382338 307186 382574
rect 307422 382338 307454 382574
rect 306834 345694 307454 382338
rect 306834 345458 306866 345694
rect 307102 345458 307186 345694
rect 307422 345458 307454 345694
rect 306834 345374 307454 345458
rect 306834 345138 306866 345374
rect 307102 345138 307186 345374
rect 307422 345138 307454 345374
rect 306834 308494 307454 345138
rect 306834 308258 306866 308494
rect 307102 308258 307186 308494
rect 307422 308258 307454 308494
rect 306834 308174 307454 308258
rect 306834 307938 306866 308174
rect 307102 307938 307186 308174
rect 307422 307938 307454 308174
rect 306834 271294 307454 307938
rect 306834 271058 306866 271294
rect 307102 271058 307186 271294
rect 307422 271058 307454 271294
rect 306834 270974 307454 271058
rect 306834 270738 306866 270974
rect 307102 270738 307186 270974
rect 307422 270738 307454 270974
rect 306834 234094 307454 270738
rect 306834 233858 306866 234094
rect 307102 233858 307186 234094
rect 307422 233858 307454 234094
rect 306834 233774 307454 233858
rect 306834 233538 306866 233774
rect 307102 233538 307186 233774
rect 307422 233538 307454 233774
rect 306834 196894 307454 233538
rect 306834 196658 306866 196894
rect 307102 196658 307186 196894
rect 307422 196658 307454 196894
rect 306834 196574 307454 196658
rect 306834 196338 306866 196574
rect 307102 196338 307186 196574
rect 307422 196338 307454 196574
rect 306834 159694 307454 196338
rect 306834 159458 306866 159694
rect 307102 159458 307186 159694
rect 307422 159458 307454 159694
rect 306834 159374 307454 159458
rect 306834 159138 306866 159374
rect 307102 159138 307186 159374
rect 307422 159138 307454 159374
rect 306834 122494 307454 159138
rect 306834 122258 306866 122494
rect 307102 122258 307186 122494
rect 307422 122258 307454 122494
rect 306834 122174 307454 122258
rect 306834 121938 306866 122174
rect 307102 121938 307186 122174
rect 307422 121938 307454 122174
rect 306834 85294 307454 121938
rect 306834 85058 306866 85294
rect 307102 85058 307186 85294
rect 307422 85058 307454 85294
rect 306834 84974 307454 85058
rect 306834 84738 306866 84974
rect 307102 84738 307186 84974
rect 307422 84738 307454 84974
rect 306834 48094 307454 84738
rect 306834 47858 306866 48094
rect 307102 47858 307186 48094
rect 307422 47858 307454 48094
rect 306834 47774 307454 47858
rect 306834 47538 306866 47774
rect 307102 47538 307186 47774
rect 307422 47538 307454 47774
rect 306834 10894 307454 47538
rect 306834 10658 306866 10894
rect 307102 10658 307186 10894
rect 307422 10658 307454 10894
rect 306834 10574 307454 10658
rect 306834 10338 306866 10574
rect 307102 10338 307186 10574
rect 307422 10338 307454 10574
rect 306834 2176 307454 10338
rect 310554 684214 311174 701760
rect 310554 683978 310586 684214
rect 310822 683978 310906 684214
rect 311142 683978 311174 684214
rect 310554 683894 311174 683978
rect 310554 683658 310586 683894
rect 310822 683658 310906 683894
rect 311142 683658 311174 683894
rect 310554 647014 311174 683658
rect 310554 646778 310586 647014
rect 310822 646778 310906 647014
rect 311142 646778 311174 647014
rect 310554 646694 311174 646778
rect 310554 646458 310586 646694
rect 310822 646458 310906 646694
rect 311142 646458 311174 646694
rect 310554 609814 311174 646458
rect 310554 609578 310586 609814
rect 310822 609578 310906 609814
rect 311142 609578 311174 609814
rect 310554 609494 311174 609578
rect 310554 609258 310586 609494
rect 310822 609258 310906 609494
rect 311142 609258 311174 609494
rect 310554 572614 311174 609258
rect 310554 572378 310586 572614
rect 310822 572378 310906 572614
rect 311142 572378 311174 572614
rect 310554 572294 311174 572378
rect 310554 572058 310586 572294
rect 310822 572058 310906 572294
rect 311142 572058 311174 572294
rect 310554 535414 311174 572058
rect 310554 535178 310586 535414
rect 310822 535178 310906 535414
rect 311142 535178 311174 535414
rect 310554 535094 311174 535178
rect 310554 534858 310586 535094
rect 310822 534858 310906 535094
rect 311142 534858 311174 535094
rect 310554 498214 311174 534858
rect 310554 497978 310586 498214
rect 310822 497978 310906 498214
rect 311142 497978 311174 498214
rect 310554 497894 311174 497978
rect 310554 497658 310586 497894
rect 310822 497658 310906 497894
rect 311142 497658 311174 497894
rect 310554 461014 311174 497658
rect 310554 460778 310586 461014
rect 310822 460778 310906 461014
rect 311142 460778 311174 461014
rect 310554 460694 311174 460778
rect 310554 460458 310586 460694
rect 310822 460458 310906 460694
rect 311142 460458 311174 460694
rect 310554 423814 311174 460458
rect 310554 423578 310586 423814
rect 310822 423578 310906 423814
rect 311142 423578 311174 423814
rect 310554 423494 311174 423578
rect 310554 423258 310586 423494
rect 310822 423258 310906 423494
rect 311142 423258 311174 423494
rect 310554 386614 311174 423258
rect 310554 386378 310586 386614
rect 310822 386378 310906 386614
rect 311142 386378 311174 386614
rect 310554 386294 311174 386378
rect 310554 386058 310586 386294
rect 310822 386058 310906 386294
rect 311142 386058 311174 386294
rect 310554 349414 311174 386058
rect 310554 349178 310586 349414
rect 310822 349178 310906 349414
rect 311142 349178 311174 349414
rect 310554 349094 311174 349178
rect 310554 348858 310586 349094
rect 310822 348858 310906 349094
rect 311142 348858 311174 349094
rect 310554 312214 311174 348858
rect 310554 311978 310586 312214
rect 310822 311978 310906 312214
rect 311142 311978 311174 312214
rect 310554 311894 311174 311978
rect 310554 311658 310586 311894
rect 310822 311658 310906 311894
rect 311142 311658 311174 311894
rect 310554 275014 311174 311658
rect 310554 274778 310586 275014
rect 310822 274778 310906 275014
rect 311142 274778 311174 275014
rect 310554 274694 311174 274778
rect 310554 274458 310586 274694
rect 310822 274458 310906 274694
rect 311142 274458 311174 274694
rect 310554 237814 311174 274458
rect 310554 237578 310586 237814
rect 310822 237578 310906 237814
rect 311142 237578 311174 237814
rect 310554 237494 311174 237578
rect 310554 237258 310586 237494
rect 310822 237258 310906 237494
rect 311142 237258 311174 237494
rect 310554 200614 311174 237258
rect 310554 200378 310586 200614
rect 310822 200378 310906 200614
rect 311142 200378 311174 200614
rect 310554 200294 311174 200378
rect 310554 200058 310586 200294
rect 310822 200058 310906 200294
rect 311142 200058 311174 200294
rect 310554 163414 311174 200058
rect 310554 163178 310586 163414
rect 310822 163178 310906 163414
rect 311142 163178 311174 163414
rect 310554 163094 311174 163178
rect 310554 162858 310586 163094
rect 310822 162858 310906 163094
rect 311142 162858 311174 163094
rect 310554 126214 311174 162858
rect 310554 125978 310586 126214
rect 310822 125978 310906 126214
rect 311142 125978 311174 126214
rect 310554 125894 311174 125978
rect 310554 125658 310586 125894
rect 310822 125658 310906 125894
rect 311142 125658 311174 125894
rect 310554 89014 311174 125658
rect 310554 88778 310586 89014
rect 310822 88778 310906 89014
rect 311142 88778 311174 89014
rect 310554 88694 311174 88778
rect 310554 88458 310586 88694
rect 310822 88458 310906 88694
rect 311142 88458 311174 88694
rect 310554 51814 311174 88458
rect 310554 51578 310586 51814
rect 310822 51578 310906 51814
rect 311142 51578 311174 51814
rect 310554 51494 311174 51578
rect 310554 51258 310586 51494
rect 310822 51258 310906 51494
rect 311142 51258 311174 51494
rect 310554 14614 311174 51258
rect 310554 14378 310586 14614
rect 310822 14378 310906 14614
rect 311142 14378 311174 14614
rect 310554 14294 311174 14378
rect 310554 14058 310586 14294
rect 310822 14058 310906 14294
rect 311142 14058 311174 14294
rect 310554 2176 311174 14058
rect 314274 687934 314894 701760
rect 314274 687698 314306 687934
rect 314542 687698 314626 687934
rect 314862 687698 314894 687934
rect 314274 687614 314894 687698
rect 314274 687378 314306 687614
rect 314542 687378 314626 687614
rect 314862 687378 314894 687614
rect 314274 650734 314894 687378
rect 314274 650498 314306 650734
rect 314542 650498 314626 650734
rect 314862 650498 314894 650734
rect 314274 650414 314894 650498
rect 314274 650178 314306 650414
rect 314542 650178 314626 650414
rect 314862 650178 314894 650414
rect 314274 613534 314894 650178
rect 314274 613298 314306 613534
rect 314542 613298 314626 613534
rect 314862 613298 314894 613534
rect 314274 613214 314894 613298
rect 314274 612978 314306 613214
rect 314542 612978 314626 613214
rect 314862 612978 314894 613214
rect 314274 576334 314894 612978
rect 314274 576098 314306 576334
rect 314542 576098 314626 576334
rect 314862 576098 314894 576334
rect 314274 576014 314894 576098
rect 314274 575778 314306 576014
rect 314542 575778 314626 576014
rect 314862 575778 314894 576014
rect 314274 539134 314894 575778
rect 314274 538898 314306 539134
rect 314542 538898 314626 539134
rect 314862 538898 314894 539134
rect 314274 538814 314894 538898
rect 314274 538578 314306 538814
rect 314542 538578 314626 538814
rect 314862 538578 314894 538814
rect 314274 501934 314894 538578
rect 314274 501698 314306 501934
rect 314542 501698 314626 501934
rect 314862 501698 314894 501934
rect 314274 501614 314894 501698
rect 314274 501378 314306 501614
rect 314542 501378 314626 501614
rect 314862 501378 314894 501614
rect 314274 464734 314894 501378
rect 314274 464498 314306 464734
rect 314542 464498 314626 464734
rect 314862 464498 314894 464734
rect 314274 464414 314894 464498
rect 314274 464178 314306 464414
rect 314542 464178 314626 464414
rect 314862 464178 314894 464414
rect 314274 427534 314894 464178
rect 314274 427298 314306 427534
rect 314542 427298 314626 427534
rect 314862 427298 314894 427534
rect 314274 427214 314894 427298
rect 314274 426978 314306 427214
rect 314542 426978 314626 427214
rect 314862 426978 314894 427214
rect 314274 390334 314894 426978
rect 314274 390098 314306 390334
rect 314542 390098 314626 390334
rect 314862 390098 314894 390334
rect 314274 390014 314894 390098
rect 314274 389778 314306 390014
rect 314542 389778 314626 390014
rect 314862 389778 314894 390014
rect 314274 353134 314894 389778
rect 314274 352898 314306 353134
rect 314542 352898 314626 353134
rect 314862 352898 314894 353134
rect 314274 352814 314894 352898
rect 314274 352578 314306 352814
rect 314542 352578 314626 352814
rect 314862 352578 314894 352814
rect 314274 315934 314894 352578
rect 314274 315698 314306 315934
rect 314542 315698 314626 315934
rect 314862 315698 314894 315934
rect 314274 315614 314894 315698
rect 314274 315378 314306 315614
rect 314542 315378 314626 315614
rect 314862 315378 314894 315614
rect 314274 278734 314894 315378
rect 314274 278498 314306 278734
rect 314542 278498 314626 278734
rect 314862 278498 314894 278734
rect 314274 278414 314894 278498
rect 314274 278178 314306 278414
rect 314542 278178 314626 278414
rect 314862 278178 314894 278414
rect 314274 241534 314894 278178
rect 314274 241298 314306 241534
rect 314542 241298 314626 241534
rect 314862 241298 314894 241534
rect 314274 241214 314894 241298
rect 314274 240978 314306 241214
rect 314542 240978 314626 241214
rect 314862 240978 314894 241214
rect 314274 204334 314894 240978
rect 314274 204098 314306 204334
rect 314542 204098 314626 204334
rect 314862 204098 314894 204334
rect 314274 204014 314894 204098
rect 314274 203778 314306 204014
rect 314542 203778 314626 204014
rect 314862 203778 314894 204014
rect 314274 167134 314894 203778
rect 314274 166898 314306 167134
rect 314542 166898 314626 167134
rect 314862 166898 314894 167134
rect 314274 166814 314894 166898
rect 314274 166578 314306 166814
rect 314542 166578 314626 166814
rect 314862 166578 314894 166814
rect 314274 129934 314894 166578
rect 314274 129698 314306 129934
rect 314542 129698 314626 129934
rect 314862 129698 314894 129934
rect 314274 129614 314894 129698
rect 314274 129378 314306 129614
rect 314542 129378 314626 129614
rect 314862 129378 314894 129614
rect 314274 92734 314894 129378
rect 314274 92498 314306 92734
rect 314542 92498 314626 92734
rect 314862 92498 314894 92734
rect 314274 92414 314894 92498
rect 314274 92178 314306 92414
rect 314542 92178 314626 92414
rect 314862 92178 314894 92414
rect 314274 55534 314894 92178
rect 314274 55298 314306 55534
rect 314542 55298 314626 55534
rect 314862 55298 314894 55534
rect 314274 55214 314894 55298
rect 314274 54978 314306 55214
rect 314542 54978 314626 55214
rect 314862 54978 314894 55214
rect 314274 18334 314894 54978
rect 314274 18098 314306 18334
rect 314542 18098 314626 18334
rect 314862 18098 314894 18334
rect 314274 18014 314894 18098
rect 314274 17778 314306 18014
rect 314542 17778 314626 18014
rect 314862 17778 314894 18014
rect 314274 2176 314894 17778
rect 317994 691654 318614 701760
rect 317994 691418 318026 691654
rect 318262 691418 318346 691654
rect 318582 691418 318614 691654
rect 317994 691334 318614 691418
rect 317994 691098 318026 691334
rect 318262 691098 318346 691334
rect 318582 691098 318614 691334
rect 317994 654454 318614 691098
rect 317994 654218 318026 654454
rect 318262 654218 318346 654454
rect 318582 654218 318614 654454
rect 317994 654134 318614 654218
rect 317994 653898 318026 654134
rect 318262 653898 318346 654134
rect 318582 653898 318614 654134
rect 317994 617254 318614 653898
rect 317994 617018 318026 617254
rect 318262 617018 318346 617254
rect 318582 617018 318614 617254
rect 317994 616934 318614 617018
rect 317994 616698 318026 616934
rect 318262 616698 318346 616934
rect 318582 616698 318614 616934
rect 317994 580054 318614 616698
rect 317994 579818 318026 580054
rect 318262 579818 318346 580054
rect 318582 579818 318614 580054
rect 317994 579734 318614 579818
rect 317994 579498 318026 579734
rect 318262 579498 318346 579734
rect 318582 579498 318614 579734
rect 317994 542854 318614 579498
rect 317994 542618 318026 542854
rect 318262 542618 318346 542854
rect 318582 542618 318614 542854
rect 317994 542534 318614 542618
rect 317994 542298 318026 542534
rect 318262 542298 318346 542534
rect 318582 542298 318614 542534
rect 317994 505654 318614 542298
rect 317994 505418 318026 505654
rect 318262 505418 318346 505654
rect 318582 505418 318614 505654
rect 317994 505334 318614 505418
rect 317994 505098 318026 505334
rect 318262 505098 318346 505334
rect 318582 505098 318614 505334
rect 317994 468454 318614 505098
rect 317994 468218 318026 468454
rect 318262 468218 318346 468454
rect 318582 468218 318614 468454
rect 317994 468134 318614 468218
rect 317994 467898 318026 468134
rect 318262 467898 318346 468134
rect 318582 467898 318614 468134
rect 317994 431254 318614 467898
rect 317994 431018 318026 431254
rect 318262 431018 318346 431254
rect 318582 431018 318614 431254
rect 317994 430934 318614 431018
rect 317994 430698 318026 430934
rect 318262 430698 318346 430934
rect 318582 430698 318614 430934
rect 317994 394054 318614 430698
rect 317994 393818 318026 394054
rect 318262 393818 318346 394054
rect 318582 393818 318614 394054
rect 317994 393734 318614 393818
rect 317994 393498 318026 393734
rect 318262 393498 318346 393734
rect 318582 393498 318614 393734
rect 317994 356854 318614 393498
rect 317994 356618 318026 356854
rect 318262 356618 318346 356854
rect 318582 356618 318614 356854
rect 317994 356534 318614 356618
rect 317994 356298 318026 356534
rect 318262 356298 318346 356534
rect 318582 356298 318614 356534
rect 317994 319654 318614 356298
rect 317994 319418 318026 319654
rect 318262 319418 318346 319654
rect 318582 319418 318614 319654
rect 317994 319334 318614 319418
rect 317994 319098 318026 319334
rect 318262 319098 318346 319334
rect 318582 319098 318614 319334
rect 317994 282454 318614 319098
rect 317994 282218 318026 282454
rect 318262 282218 318346 282454
rect 318582 282218 318614 282454
rect 317994 282134 318614 282218
rect 317994 281898 318026 282134
rect 318262 281898 318346 282134
rect 318582 281898 318614 282134
rect 317994 245254 318614 281898
rect 317994 245018 318026 245254
rect 318262 245018 318346 245254
rect 318582 245018 318614 245254
rect 317994 244934 318614 245018
rect 317994 244698 318026 244934
rect 318262 244698 318346 244934
rect 318582 244698 318614 244934
rect 317994 208054 318614 244698
rect 317994 207818 318026 208054
rect 318262 207818 318346 208054
rect 318582 207818 318614 208054
rect 317994 207734 318614 207818
rect 317994 207498 318026 207734
rect 318262 207498 318346 207734
rect 318582 207498 318614 207734
rect 317994 170854 318614 207498
rect 317994 170618 318026 170854
rect 318262 170618 318346 170854
rect 318582 170618 318614 170854
rect 317994 170534 318614 170618
rect 317994 170298 318026 170534
rect 318262 170298 318346 170534
rect 318582 170298 318614 170534
rect 317994 133654 318614 170298
rect 317994 133418 318026 133654
rect 318262 133418 318346 133654
rect 318582 133418 318614 133654
rect 317994 133334 318614 133418
rect 317994 133098 318026 133334
rect 318262 133098 318346 133334
rect 318582 133098 318614 133334
rect 317994 96454 318614 133098
rect 317994 96218 318026 96454
rect 318262 96218 318346 96454
rect 318582 96218 318614 96454
rect 317994 96134 318614 96218
rect 317994 95898 318026 96134
rect 318262 95898 318346 96134
rect 318582 95898 318614 96134
rect 317994 59254 318614 95898
rect 317994 59018 318026 59254
rect 318262 59018 318346 59254
rect 318582 59018 318614 59254
rect 317994 58934 318614 59018
rect 317994 58698 318026 58934
rect 318262 58698 318346 58934
rect 318582 58698 318614 58934
rect 317994 22054 318614 58698
rect 317994 21818 318026 22054
rect 318262 21818 318346 22054
rect 318582 21818 318614 22054
rect 317994 21734 318614 21818
rect 317994 21498 318026 21734
rect 318262 21498 318346 21734
rect 318582 21498 318614 21734
rect 317994 2176 318614 21498
rect 321714 695374 322334 701760
rect 321714 695138 321746 695374
rect 321982 695138 322066 695374
rect 322302 695138 322334 695374
rect 321714 695054 322334 695138
rect 321714 694818 321746 695054
rect 321982 694818 322066 695054
rect 322302 694818 322334 695054
rect 321714 658174 322334 694818
rect 321714 657938 321746 658174
rect 321982 657938 322066 658174
rect 322302 657938 322334 658174
rect 321714 657854 322334 657938
rect 321714 657618 321746 657854
rect 321982 657618 322066 657854
rect 322302 657618 322334 657854
rect 321714 620974 322334 657618
rect 321714 620738 321746 620974
rect 321982 620738 322066 620974
rect 322302 620738 322334 620974
rect 321714 620654 322334 620738
rect 321714 620418 321746 620654
rect 321982 620418 322066 620654
rect 322302 620418 322334 620654
rect 321714 583774 322334 620418
rect 321714 583538 321746 583774
rect 321982 583538 322066 583774
rect 322302 583538 322334 583774
rect 321714 583454 322334 583538
rect 321714 583218 321746 583454
rect 321982 583218 322066 583454
rect 322302 583218 322334 583454
rect 321714 546574 322334 583218
rect 321714 546338 321746 546574
rect 321982 546338 322066 546574
rect 322302 546338 322334 546574
rect 321714 546254 322334 546338
rect 321714 546018 321746 546254
rect 321982 546018 322066 546254
rect 322302 546018 322334 546254
rect 321714 509374 322334 546018
rect 321714 509138 321746 509374
rect 321982 509138 322066 509374
rect 322302 509138 322334 509374
rect 321714 509054 322334 509138
rect 321714 508818 321746 509054
rect 321982 508818 322066 509054
rect 322302 508818 322334 509054
rect 321714 472174 322334 508818
rect 321714 471938 321746 472174
rect 321982 471938 322066 472174
rect 322302 471938 322334 472174
rect 321714 471854 322334 471938
rect 321714 471618 321746 471854
rect 321982 471618 322066 471854
rect 322302 471618 322334 471854
rect 321714 434974 322334 471618
rect 321714 434738 321746 434974
rect 321982 434738 322066 434974
rect 322302 434738 322334 434974
rect 321714 434654 322334 434738
rect 321714 434418 321746 434654
rect 321982 434418 322066 434654
rect 322302 434418 322334 434654
rect 321714 397774 322334 434418
rect 321714 397538 321746 397774
rect 321982 397538 322066 397774
rect 322302 397538 322334 397774
rect 321714 397454 322334 397538
rect 321714 397218 321746 397454
rect 321982 397218 322066 397454
rect 322302 397218 322334 397454
rect 321714 360574 322334 397218
rect 321714 360338 321746 360574
rect 321982 360338 322066 360574
rect 322302 360338 322334 360574
rect 321714 360254 322334 360338
rect 321714 360018 321746 360254
rect 321982 360018 322066 360254
rect 322302 360018 322334 360254
rect 321714 323374 322334 360018
rect 321714 323138 321746 323374
rect 321982 323138 322066 323374
rect 322302 323138 322334 323374
rect 321714 323054 322334 323138
rect 321714 322818 321746 323054
rect 321982 322818 322066 323054
rect 322302 322818 322334 323054
rect 321714 286174 322334 322818
rect 321714 285938 321746 286174
rect 321982 285938 322066 286174
rect 322302 285938 322334 286174
rect 321714 285854 322334 285938
rect 321714 285618 321746 285854
rect 321982 285618 322066 285854
rect 322302 285618 322334 285854
rect 321714 248974 322334 285618
rect 321714 248738 321746 248974
rect 321982 248738 322066 248974
rect 322302 248738 322334 248974
rect 321714 248654 322334 248738
rect 321714 248418 321746 248654
rect 321982 248418 322066 248654
rect 322302 248418 322334 248654
rect 321714 211774 322334 248418
rect 321714 211538 321746 211774
rect 321982 211538 322066 211774
rect 322302 211538 322334 211774
rect 321714 211454 322334 211538
rect 321714 211218 321746 211454
rect 321982 211218 322066 211454
rect 322302 211218 322334 211454
rect 321714 174574 322334 211218
rect 321714 174338 321746 174574
rect 321982 174338 322066 174574
rect 322302 174338 322334 174574
rect 321714 174254 322334 174338
rect 321714 174018 321746 174254
rect 321982 174018 322066 174254
rect 322302 174018 322334 174254
rect 321714 137374 322334 174018
rect 321714 137138 321746 137374
rect 321982 137138 322066 137374
rect 322302 137138 322334 137374
rect 321714 137054 322334 137138
rect 321714 136818 321746 137054
rect 321982 136818 322066 137054
rect 322302 136818 322334 137054
rect 321714 100174 322334 136818
rect 321714 99938 321746 100174
rect 321982 99938 322066 100174
rect 322302 99938 322334 100174
rect 321714 99854 322334 99938
rect 321714 99618 321746 99854
rect 321982 99618 322066 99854
rect 322302 99618 322334 99854
rect 321714 62974 322334 99618
rect 321714 62738 321746 62974
rect 321982 62738 322066 62974
rect 322302 62738 322334 62974
rect 321714 62654 322334 62738
rect 321714 62418 321746 62654
rect 321982 62418 322066 62654
rect 322302 62418 322334 62654
rect 321714 25774 322334 62418
rect 321714 25538 321746 25774
rect 321982 25538 322066 25774
rect 322302 25538 322334 25774
rect 321714 25454 322334 25538
rect 321714 25218 321746 25454
rect 321982 25218 322066 25454
rect 322302 25218 322334 25454
rect 321714 2176 322334 25218
rect 325434 699094 326054 701760
rect 325434 698858 325466 699094
rect 325702 698858 325786 699094
rect 326022 698858 326054 699094
rect 325434 698774 326054 698858
rect 325434 698538 325466 698774
rect 325702 698538 325786 698774
rect 326022 698538 326054 698774
rect 325434 661894 326054 698538
rect 325434 661658 325466 661894
rect 325702 661658 325786 661894
rect 326022 661658 326054 661894
rect 325434 661574 326054 661658
rect 325434 661338 325466 661574
rect 325702 661338 325786 661574
rect 326022 661338 326054 661574
rect 325434 624694 326054 661338
rect 325434 624458 325466 624694
rect 325702 624458 325786 624694
rect 326022 624458 326054 624694
rect 325434 624374 326054 624458
rect 325434 624138 325466 624374
rect 325702 624138 325786 624374
rect 326022 624138 326054 624374
rect 325434 587494 326054 624138
rect 325434 587258 325466 587494
rect 325702 587258 325786 587494
rect 326022 587258 326054 587494
rect 325434 587174 326054 587258
rect 325434 586938 325466 587174
rect 325702 586938 325786 587174
rect 326022 586938 326054 587174
rect 325434 550294 326054 586938
rect 325434 550058 325466 550294
rect 325702 550058 325786 550294
rect 326022 550058 326054 550294
rect 325434 549974 326054 550058
rect 325434 549738 325466 549974
rect 325702 549738 325786 549974
rect 326022 549738 326054 549974
rect 325434 513094 326054 549738
rect 325434 512858 325466 513094
rect 325702 512858 325786 513094
rect 326022 512858 326054 513094
rect 325434 512774 326054 512858
rect 325434 512538 325466 512774
rect 325702 512538 325786 512774
rect 326022 512538 326054 512774
rect 325434 475894 326054 512538
rect 325434 475658 325466 475894
rect 325702 475658 325786 475894
rect 326022 475658 326054 475894
rect 325434 475574 326054 475658
rect 325434 475338 325466 475574
rect 325702 475338 325786 475574
rect 326022 475338 326054 475574
rect 325434 438694 326054 475338
rect 325434 438458 325466 438694
rect 325702 438458 325786 438694
rect 326022 438458 326054 438694
rect 325434 438374 326054 438458
rect 325434 438138 325466 438374
rect 325702 438138 325786 438374
rect 326022 438138 326054 438374
rect 325434 401494 326054 438138
rect 325434 401258 325466 401494
rect 325702 401258 325786 401494
rect 326022 401258 326054 401494
rect 325434 401174 326054 401258
rect 325434 400938 325466 401174
rect 325702 400938 325786 401174
rect 326022 400938 326054 401174
rect 325434 364294 326054 400938
rect 325434 364058 325466 364294
rect 325702 364058 325786 364294
rect 326022 364058 326054 364294
rect 325434 363974 326054 364058
rect 325434 363738 325466 363974
rect 325702 363738 325786 363974
rect 326022 363738 326054 363974
rect 325434 327094 326054 363738
rect 325434 326858 325466 327094
rect 325702 326858 325786 327094
rect 326022 326858 326054 327094
rect 325434 326774 326054 326858
rect 325434 326538 325466 326774
rect 325702 326538 325786 326774
rect 326022 326538 326054 326774
rect 325434 289894 326054 326538
rect 325434 289658 325466 289894
rect 325702 289658 325786 289894
rect 326022 289658 326054 289894
rect 325434 289574 326054 289658
rect 325434 289338 325466 289574
rect 325702 289338 325786 289574
rect 326022 289338 326054 289574
rect 325434 252694 326054 289338
rect 325434 252458 325466 252694
rect 325702 252458 325786 252694
rect 326022 252458 326054 252694
rect 325434 252374 326054 252458
rect 325434 252138 325466 252374
rect 325702 252138 325786 252374
rect 326022 252138 326054 252374
rect 325434 215494 326054 252138
rect 325434 215258 325466 215494
rect 325702 215258 325786 215494
rect 326022 215258 326054 215494
rect 325434 215174 326054 215258
rect 325434 214938 325466 215174
rect 325702 214938 325786 215174
rect 326022 214938 326054 215174
rect 325434 178294 326054 214938
rect 325434 178058 325466 178294
rect 325702 178058 325786 178294
rect 326022 178058 326054 178294
rect 325434 177974 326054 178058
rect 325434 177738 325466 177974
rect 325702 177738 325786 177974
rect 326022 177738 326054 177974
rect 325434 141094 326054 177738
rect 325434 140858 325466 141094
rect 325702 140858 325786 141094
rect 326022 140858 326054 141094
rect 325434 140774 326054 140858
rect 325434 140538 325466 140774
rect 325702 140538 325786 140774
rect 326022 140538 326054 140774
rect 325434 103894 326054 140538
rect 325434 103658 325466 103894
rect 325702 103658 325786 103894
rect 326022 103658 326054 103894
rect 325434 103574 326054 103658
rect 325434 103338 325466 103574
rect 325702 103338 325786 103574
rect 326022 103338 326054 103574
rect 325434 66694 326054 103338
rect 325434 66458 325466 66694
rect 325702 66458 325786 66694
rect 326022 66458 326054 66694
rect 325434 66374 326054 66458
rect 325434 66138 325466 66374
rect 325702 66138 325786 66374
rect 326022 66138 326054 66374
rect 325434 29494 326054 66138
rect 325434 29258 325466 29494
rect 325702 29258 325786 29494
rect 326022 29258 326054 29494
rect 325434 29174 326054 29258
rect 325434 28938 325466 29174
rect 325702 28938 325786 29174
rect 326022 28938 326054 29174
rect 325434 2176 326054 28938
rect 336594 673054 337214 701760
rect 336594 672818 336626 673054
rect 336862 672818 336946 673054
rect 337182 672818 337214 673054
rect 336594 672734 337214 672818
rect 336594 672498 336626 672734
rect 336862 672498 336946 672734
rect 337182 672498 337214 672734
rect 336594 635854 337214 672498
rect 336594 635618 336626 635854
rect 336862 635618 336946 635854
rect 337182 635618 337214 635854
rect 336594 635534 337214 635618
rect 336594 635298 336626 635534
rect 336862 635298 336946 635534
rect 337182 635298 337214 635534
rect 336594 598654 337214 635298
rect 336594 598418 336626 598654
rect 336862 598418 336946 598654
rect 337182 598418 337214 598654
rect 336594 598334 337214 598418
rect 336594 598098 336626 598334
rect 336862 598098 336946 598334
rect 337182 598098 337214 598334
rect 336594 561454 337214 598098
rect 336594 561218 336626 561454
rect 336862 561218 336946 561454
rect 337182 561218 337214 561454
rect 336594 561134 337214 561218
rect 336594 560898 336626 561134
rect 336862 560898 336946 561134
rect 337182 560898 337214 561134
rect 336594 524254 337214 560898
rect 336594 524018 336626 524254
rect 336862 524018 336946 524254
rect 337182 524018 337214 524254
rect 336594 523934 337214 524018
rect 336594 523698 336626 523934
rect 336862 523698 336946 523934
rect 337182 523698 337214 523934
rect 336594 487054 337214 523698
rect 336594 486818 336626 487054
rect 336862 486818 336946 487054
rect 337182 486818 337214 487054
rect 336594 486734 337214 486818
rect 336594 486498 336626 486734
rect 336862 486498 336946 486734
rect 337182 486498 337214 486734
rect 336594 449854 337214 486498
rect 336594 449618 336626 449854
rect 336862 449618 336946 449854
rect 337182 449618 337214 449854
rect 336594 449534 337214 449618
rect 336594 449298 336626 449534
rect 336862 449298 336946 449534
rect 337182 449298 337214 449534
rect 336594 412654 337214 449298
rect 336594 412418 336626 412654
rect 336862 412418 336946 412654
rect 337182 412418 337214 412654
rect 336594 412334 337214 412418
rect 336594 412098 336626 412334
rect 336862 412098 336946 412334
rect 337182 412098 337214 412334
rect 336594 375454 337214 412098
rect 336594 375218 336626 375454
rect 336862 375218 336946 375454
rect 337182 375218 337214 375454
rect 336594 375134 337214 375218
rect 336594 374898 336626 375134
rect 336862 374898 336946 375134
rect 337182 374898 337214 375134
rect 336594 338254 337214 374898
rect 336594 338018 336626 338254
rect 336862 338018 336946 338254
rect 337182 338018 337214 338254
rect 336594 337934 337214 338018
rect 336594 337698 336626 337934
rect 336862 337698 336946 337934
rect 337182 337698 337214 337934
rect 336594 301054 337214 337698
rect 336594 300818 336626 301054
rect 336862 300818 336946 301054
rect 337182 300818 337214 301054
rect 336594 300734 337214 300818
rect 336594 300498 336626 300734
rect 336862 300498 336946 300734
rect 337182 300498 337214 300734
rect 336594 263854 337214 300498
rect 336594 263618 336626 263854
rect 336862 263618 336946 263854
rect 337182 263618 337214 263854
rect 336594 263534 337214 263618
rect 336594 263298 336626 263534
rect 336862 263298 336946 263534
rect 337182 263298 337214 263534
rect 336594 226654 337214 263298
rect 336594 226418 336626 226654
rect 336862 226418 336946 226654
rect 337182 226418 337214 226654
rect 336594 226334 337214 226418
rect 336594 226098 336626 226334
rect 336862 226098 336946 226334
rect 337182 226098 337214 226334
rect 336594 189454 337214 226098
rect 336594 189218 336626 189454
rect 336862 189218 336946 189454
rect 337182 189218 337214 189454
rect 336594 189134 337214 189218
rect 336594 188898 336626 189134
rect 336862 188898 336946 189134
rect 337182 188898 337214 189134
rect 336594 152254 337214 188898
rect 336594 152018 336626 152254
rect 336862 152018 336946 152254
rect 337182 152018 337214 152254
rect 336594 151934 337214 152018
rect 336594 151698 336626 151934
rect 336862 151698 336946 151934
rect 337182 151698 337214 151934
rect 336594 115054 337214 151698
rect 336594 114818 336626 115054
rect 336862 114818 336946 115054
rect 337182 114818 337214 115054
rect 336594 114734 337214 114818
rect 336594 114498 336626 114734
rect 336862 114498 336946 114734
rect 337182 114498 337214 114734
rect 336594 77854 337214 114498
rect 336594 77618 336626 77854
rect 336862 77618 336946 77854
rect 337182 77618 337214 77854
rect 336594 77534 337214 77618
rect 336594 77298 336626 77534
rect 336862 77298 336946 77534
rect 337182 77298 337214 77534
rect 336594 40654 337214 77298
rect 336594 40418 336626 40654
rect 336862 40418 336946 40654
rect 337182 40418 337214 40654
rect 336594 40334 337214 40418
rect 336594 40098 336626 40334
rect 336862 40098 336946 40334
rect 337182 40098 337214 40334
rect 336594 3454 337214 40098
rect 336594 3218 336626 3454
rect 336862 3218 336946 3454
rect 337182 3218 337214 3454
rect 336594 3134 337214 3218
rect 336594 2898 336626 3134
rect 336862 2898 336946 3134
rect 337182 2898 337214 3134
rect 336594 2176 337214 2898
rect 340314 676774 340934 701760
rect 340314 676538 340346 676774
rect 340582 676538 340666 676774
rect 340902 676538 340934 676774
rect 340314 676454 340934 676538
rect 340314 676218 340346 676454
rect 340582 676218 340666 676454
rect 340902 676218 340934 676454
rect 340314 639574 340934 676218
rect 340314 639338 340346 639574
rect 340582 639338 340666 639574
rect 340902 639338 340934 639574
rect 340314 639254 340934 639338
rect 340314 639018 340346 639254
rect 340582 639018 340666 639254
rect 340902 639018 340934 639254
rect 340314 602374 340934 639018
rect 340314 602138 340346 602374
rect 340582 602138 340666 602374
rect 340902 602138 340934 602374
rect 340314 602054 340934 602138
rect 340314 601818 340346 602054
rect 340582 601818 340666 602054
rect 340902 601818 340934 602054
rect 340314 565174 340934 601818
rect 340314 564938 340346 565174
rect 340582 564938 340666 565174
rect 340902 564938 340934 565174
rect 340314 564854 340934 564938
rect 340314 564618 340346 564854
rect 340582 564618 340666 564854
rect 340902 564618 340934 564854
rect 340314 527974 340934 564618
rect 340314 527738 340346 527974
rect 340582 527738 340666 527974
rect 340902 527738 340934 527974
rect 340314 527654 340934 527738
rect 340314 527418 340346 527654
rect 340582 527418 340666 527654
rect 340902 527418 340934 527654
rect 340314 490774 340934 527418
rect 340314 490538 340346 490774
rect 340582 490538 340666 490774
rect 340902 490538 340934 490774
rect 340314 490454 340934 490538
rect 340314 490218 340346 490454
rect 340582 490218 340666 490454
rect 340902 490218 340934 490454
rect 340314 453574 340934 490218
rect 340314 453338 340346 453574
rect 340582 453338 340666 453574
rect 340902 453338 340934 453574
rect 340314 453254 340934 453338
rect 340314 453018 340346 453254
rect 340582 453018 340666 453254
rect 340902 453018 340934 453254
rect 340314 416374 340934 453018
rect 340314 416138 340346 416374
rect 340582 416138 340666 416374
rect 340902 416138 340934 416374
rect 340314 416054 340934 416138
rect 340314 415818 340346 416054
rect 340582 415818 340666 416054
rect 340902 415818 340934 416054
rect 340314 379174 340934 415818
rect 340314 378938 340346 379174
rect 340582 378938 340666 379174
rect 340902 378938 340934 379174
rect 340314 378854 340934 378938
rect 340314 378618 340346 378854
rect 340582 378618 340666 378854
rect 340902 378618 340934 378854
rect 340314 341974 340934 378618
rect 340314 341738 340346 341974
rect 340582 341738 340666 341974
rect 340902 341738 340934 341974
rect 340314 341654 340934 341738
rect 340314 341418 340346 341654
rect 340582 341418 340666 341654
rect 340902 341418 340934 341654
rect 340314 304774 340934 341418
rect 340314 304538 340346 304774
rect 340582 304538 340666 304774
rect 340902 304538 340934 304774
rect 340314 304454 340934 304538
rect 340314 304218 340346 304454
rect 340582 304218 340666 304454
rect 340902 304218 340934 304454
rect 340314 267574 340934 304218
rect 340314 267338 340346 267574
rect 340582 267338 340666 267574
rect 340902 267338 340934 267574
rect 340314 267254 340934 267338
rect 340314 267018 340346 267254
rect 340582 267018 340666 267254
rect 340902 267018 340934 267254
rect 340314 230374 340934 267018
rect 340314 230138 340346 230374
rect 340582 230138 340666 230374
rect 340902 230138 340934 230374
rect 340314 230054 340934 230138
rect 340314 229818 340346 230054
rect 340582 229818 340666 230054
rect 340902 229818 340934 230054
rect 340314 193174 340934 229818
rect 340314 192938 340346 193174
rect 340582 192938 340666 193174
rect 340902 192938 340934 193174
rect 340314 192854 340934 192938
rect 340314 192618 340346 192854
rect 340582 192618 340666 192854
rect 340902 192618 340934 192854
rect 340314 155974 340934 192618
rect 340314 155738 340346 155974
rect 340582 155738 340666 155974
rect 340902 155738 340934 155974
rect 340314 155654 340934 155738
rect 340314 155418 340346 155654
rect 340582 155418 340666 155654
rect 340902 155418 340934 155654
rect 340314 118774 340934 155418
rect 340314 118538 340346 118774
rect 340582 118538 340666 118774
rect 340902 118538 340934 118774
rect 340314 118454 340934 118538
rect 340314 118218 340346 118454
rect 340582 118218 340666 118454
rect 340902 118218 340934 118454
rect 340314 81574 340934 118218
rect 340314 81338 340346 81574
rect 340582 81338 340666 81574
rect 340902 81338 340934 81574
rect 340314 81254 340934 81338
rect 340314 81018 340346 81254
rect 340582 81018 340666 81254
rect 340902 81018 340934 81254
rect 340314 44374 340934 81018
rect 340314 44138 340346 44374
rect 340582 44138 340666 44374
rect 340902 44138 340934 44374
rect 340314 44054 340934 44138
rect 340314 43818 340346 44054
rect 340582 43818 340666 44054
rect 340902 43818 340934 44054
rect 340314 7174 340934 43818
rect 340314 6938 340346 7174
rect 340582 6938 340666 7174
rect 340902 6938 340934 7174
rect 340314 6854 340934 6938
rect 340314 6618 340346 6854
rect 340582 6618 340666 6854
rect 340902 6618 340934 6854
rect 340314 2176 340934 6618
rect 344034 680494 344654 701760
rect 344034 680258 344066 680494
rect 344302 680258 344386 680494
rect 344622 680258 344654 680494
rect 344034 680174 344654 680258
rect 344034 679938 344066 680174
rect 344302 679938 344386 680174
rect 344622 679938 344654 680174
rect 344034 643294 344654 679938
rect 344034 643058 344066 643294
rect 344302 643058 344386 643294
rect 344622 643058 344654 643294
rect 344034 642974 344654 643058
rect 344034 642738 344066 642974
rect 344302 642738 344386 642974
rect 344622 642738 344654 642974
rect 344034 606094 344654 642738
rect 344034 605858 344066 606094
rect 344302 605858 344386 606094
rect 344622 605858 344654 606094
rect 344034 605774 344654 605858
rect 344034 605538 344066 605774
rect 344302 605538 344386 605774
rect 344622 605538 344654 605774
rect 344034 568894 344654 605538
rect 344034 568658 344066 568894
rect 344302 568658 344386 568894
rect 344622 568658 344654 568894
rect 344034 568574 344654 568658
rect 344034 568338 344066 568574
rect 344302 568338 344386 568574
rect 344622 568338 344654 568574
rect 344034 531694 344654 568338
rect 344034 531458 344066 531694
rect 344302 531458 344386 531694
rect 344622 531458 344654 531694
rect 344034 531374 344654 531458
rect 344034 531138 344066 531374
rect 344302 531138 344386 531374
rect 344622 531138 344654 531374
rect 344034 494494 344654 531138
rect 344034 494258 344066 494494
rect 344302 494258 344386 494494
rect 344622 494258 344654 494494
rect 344034 494174 344654 494258
rect 344034 493938 344066 494174
rect 344302 493938 344386 494174
rect 344622 493938 344654 494174
rect 344034 457294 344654 493938
rect 344034 457058 344066 457294
rect 344302 457058 344386 457294
rect 344622 457058 344654 457294
rect 344034 456974 344654 457058
rect 344034 456738 344066 456974
rect 344302 456738 344386 456974
rect 344622 456738 344654 456974
rect 344034 420094 344654 456738
rect 344034 419858 344066 420094
rect 344302 419858 344386 420094
rect 344622 419858 344654 420094
rect 344034 419774 344654 419858
rect 344034 419538 344066 419774
rect 344302 419538 344386 419774
rect 344622 419538 344654 419774
rect 344034 382894 344654 419538
rect 344034 382658 344066 382894
rect 344302 382658 344386 382894
rect 344622 382658 344654 382894
rect 344034 382574 344654 382658
rect 344034 382338 344066 382574
rect 344302 382338 344386 382574
rect 344622 382338 344654 382574
rect 344034 345694 344654 382338
rect 344034 345458 344066 345694
rect 344302 345458 344386 345694
rect 344622 345458 344654 345694
rect 344034 345374 344654 345458
rect 344034 345138 344066 345374
rect 344302 345138 344386 345374
rect 344622 345138 344654 345374
rect 344034 308494 344654 345138
rect 344034 308258 344066 308494
rect 344302 308258 344386 308494
rect 344622 308258 344654 308494
rect 344034 308174 344654 308258
rect 344034 307938 344066 308174
rect 344302 307938 344386 308174
rect 344622 307938 344654 308174
rect 344034 271294 344654 307938
rect 344034 271058 344066 271294
rect 344302 271058 344386 271294
rect 344622 271058 344654 271294
rect 344034 270974 344654 271058
rect 344034 270738 344066 270974
rect 344302 270738 344386 270974
rect 344622 270738 344654 270974
rect 344034 234094 344654 270738
rect 344034 233858 344066 234094
rect 344302 233858 344386 234094
rect 344622 233858 344654 234094
rect 344034 233774 344654 233858
rect 344034 233538 344066 233774
rect 344302 233538 344386 233774
rect 344622 233538 344654 233774
rect 344034 196894 344654 233538
rect 344034 196658 344066 196894
rect 344302 196658 344386 196894
rect 344622 196658 344654 196894
rect 344034 196574 344654 196658
rect 344034 196338 344066 196574
rect 344302 196338 344386 196574
rect 344622 196338 344654 196574
rect 344034 159694 344654 196338
rect 344034 159458 344066 159694
rect 344302 159458 344386 159694
rect 344622 159458 344654 159694
rect 344034 159374 344654 159458
rect 344034 159138 344066 159374
rect 344302 159138 344386 159374
rect 344622 159138 344654 159374
rect 344034 122494 344654 159138
rect 344034 122258 344066 122494
rect 344302 122258 344386 122494
rect 344622 122258 344654 122494
rect 344034 122174 344654 122258
rect 344034 121938 344066 122174
rect 344302 121938 344386 122174
rect 344622 121938 344654 122174
rect 344034 85294 344654 121938
rect 344034 85058 344066 85294
rect 344302 85058 344386 85294
rect 344622 85058 344654 85294
rect 344034 84974 344654 85058
rect 344034 84738 344066 84974
rect 344302 84738 344386 84974
rect 344622 84738 344654 84974
rect 344034 48094 344654 84738
rect 344034 47858 344066 48094
rect 344302 47858 344386 48094
rect 344622 47858 344654 48094
rect 344034 47774 344654 47858
rect 344034 47538 344066 47774
rect 344302 47538 344386 47774
rect 344622 47538 344654 47774
rect 344034 10894 344654 47538
rect 344034 10658 344066 10894
rect 344302 10658 344386 10894
rect 344622 10658 344654 10894
rect 344034 10574 344654 10658
rect 344034 10338 344066 10574
rect 344302 10338 344386 10574
rect 344622 10338 344654 10574
rect 344034 2176 344654 10338
rect 347754 684214 348374 701760
rect 347754 683978 347786 684214
rect 348022 683978 348106 684214
rect 348342 683978 348374 684214
rect 347754 683894 348374 683978
rect 347754 683658 347786 683894
rect 348022 683658 348106 683894
rect 348342 683658 348374 683894
rect 347754 647014 348374 683658
rect 347754 646778 347786 647014
rect 348022 646778 348106 647014
rect 348342 646778 348374 647014
rect 347754 646694 348374 646778
rect 347754 646458 347786 646694
rect 348022 646458 348106 646694
rect 348342 646458 348374 646694
rect 347754 609814 348374 646458
rect 347754 609578 347786 609814
rect 348022 609578 348106 609814
rect 348342 609578 348374 609814
rect 347754 609494 348374 609578
rect 347754 609258 347786 609494
rect 348022 609258 348106 609494
rect 348342 609258 348374 609494
rect 347754 572614 348374 609258
rect 347754 572378 347786 572614
rect 348022 572378 348106 572614
rect 348342 572378 348374 572614
rect 347754 572294 348374 572378
rect 347754 572058 347786 572294
rect 348022 572058 348106 572294
rect 348342 572058 348374 572294
rect 347754 535414 348374 572058
rect 347754 535178 347786 535414
rect 348022 535178 348106 535414
rect 348342 535178 348374 535414
rect 347754 535094 348374 535178
rect 347754 534858 347786 535094
rect 348022 534858 348106 535094
rect 348342 534858 348374 535094
rect 347754 498214 348374 534858
rect 347754 497978 347786 498214
rect 348022 497978 348106 498214
rect 348342 497978 348374 498214
rect 347754 497894 348374 497978
rect 347754 497658 347786 497894
rect 348022 497658 348106 497894
rect 348342 497658 348374 497894
rect 347754 461014 348374 497658
rect 347754 460778 347786 461014
rect 348022 460778 348106 461014
rect 348342 460778 348374 461014
rect 347754 460694 348374 460778
rect 347754 460458 347786 460694
rect 348022 460458 348106 460694
rect 348342 460458 348374 460694
rect 347754 423814 348374 460458
rect 347754 423578 347786 423814
rect 348022 423578 348106 423814
rect 348342 423578 348374 423814
rect 347754 423494 348374 423578
rect 347754 423258 347786 423494
rect 348022 423258 348106 423494
rect 348342 423258 348374 423494
rect 347754 386614 348374 423258
rect 347754 386378 347786 386614
rect 348022 386378 348106 386614
rect 348342 386378 348374 386614
rect 347754 386294 348374 386378
rect 347754 386058 347786 386294
rect 348022 386058 348106 386294
rect 348342 386058 348374 386294
rect 347754 349414 348374 386058
rect 347754 349178 347786 349414
rect 348022 349178 348106 349414
rect 348342 349178 348374 349414
rect 347754 349094 348374 349178
rect 347754 348858 347786 349094
rect 348022 348858 348106 349094
rect 348342 348858 348374 349094
rect 347754 312214 348374 348858
rect 347754 311978 347786 312214
rect 348022 311978 348106 312214
rect 348342 311978 348374 312214
rect 347754 311894 348374 311978
rect 347754 311658 347786 311894
rect 348022 311658 348106 311894
rect 348342 311658 348374 311894
rect 347754 275014 348374 311658
rect 347754 274778 347786 275014
rect 348022 274778 348106 275014
rect 348342 274778 348374 275014
rect 347754 274694 348374 274778
rect 347754 274458 347786 274694
rect 348022 274458 348106 274694
rect 348342 274458 348374 274694
rect 347754 237814 348374 274458
rect 347754 237578 347786 237814
rect 348022 237578 348106 237814
rect 348342 237578 348374 237814
rect 347754 237494 348374 237578
rect 347754 237258 347786 237494
rect 348022 237258 348106 237494
rect 348342 237258 348374 237494
rect 347754 200614 348374 237258
rect 347754 200378 347786 200614
rect 348022 200378 348106 200614
rect 348342 200378 348374 200614
rect 347754 200294 348374 200378
rect 347754 200058 347786 200294
rect 348022 200058 348106 200294
rect 348342 200058 348374 200294
rect 347754 163414 348374 200058
rect 347754 163178 347786 163414
rect 348022 163178 348106 163414
rect 348342 163178 348374 163414
rect 347754 163094 348374 163178
rect 347754 162858 347786 163094
rect 348022 162858 348106 163094
rect 348342 162858 348374 163094
rect 347754 126214 348374 162858
rect 347754 125978 347786 126214
rect 348022 125978 348106 126214
rect 348342 125978 348374 126214
rect 347754 125894 348374 125978
rect 347754 125658 347786 125894
rect 348022 125658 348106 125894
rect 348342 125658 348374 125894
rect 347754 89014 348374 125658
rect 347754 88778 347786 89014
rect 348022 88778 348106 89014
rect 348342 88778 348374 89014
rect 347754 88694 348374 88778
rect 347754 88458 347786 88694
rect 348022 88458 348106 88694
rect 348342 88458 348374 88694
rect 347754 51814 348374 88458
rect 347754 51578 347786 51814
rect 348022 51578 348106 51814
rect 348342 51578 348374 51814
rect 347754 51494 348374 51578
rect 347754 51258 347786 51494
rect 348022 51258 348106 51494
rect 348342 51258 348374 51494
rect 347754 14614 348374 51258
rect 347754 14378 347786 14614
rect 348022 14378 348106 14614
rect 348342 14378 348374 14614
rect 347754 14294 348374 14378
rect 347754 14058 347786 14294
rect 348022 14058 348106 14294
rect 348342 14058 348374 14294
rect 347754 2176 348374 14058
rect 351474 687934 352094 701760
rect 351474 687698 351506 687934
rect 351742 687698 351826 687934
rect 352062 687698 352094 687934
rect 351474 687614 352094 687698
rect 351474 687378 351506 687614
rect 351742 687378 351826 687614
rect 352062 687378 352094 687614
rect 351474 650734 352094 687378
rect 351474 650498 351506 650734
rect 351742 650498 351826 650734
rect 352062 650498 352094 650734
rect 351474 650414 352094 650498
rect 351474 650178 351506 650414
rect 351742 650178 351826 650414
rect 352062 650178 352094 650414
rect 351474 613534 352094 650178
rect 351474 613298 351506 613534
rect 351742 613298 351826 613534
rect 352062 613298 352094 613534
rect 351474 613214 352094 613298
rect 351474 612978 351506 613214
rect 351742 612978 351826 613214
rect 352062 612978 352094 613214
rect 351474 576334 352094 612978
rect 351474 576098 351506 576334
rect 351742 576098 351826 576334
rect 352062 576098 352094 576334
rect 351474 576014 352094 576098
rect 351474 575778 351506 576014
rect 351742 575778 351826 576014
rect 352062 575778 352094 576014
rect 351474 539134 352094 575778
rect 351474 538898 351506 539134
rect 351742 538898 351826 539134
rect 352062 538898 352094 539134
rect 351474 538814 352094 538898
rect 351474 538578 351506 538814
rect 351742 538578 351826 538814
rect 352062 538578 352094 538814
rect 351474 501934 352094 538578
rect 351474 501698 351506 501934
rect 351742 501698 351826 501934
rect 352062 501698 352094 501934
rect 351474 501614 352094 501698
rect 351474 501378 351506 501614
rect 351742 501378 351826 501614
rect 352062 501378 352094 501614
rect 351474 464734 352094 501378
rect 351474 464498 351506 464734
rect 351742 464498 351826 464734
rect 352062 464498 352094 464734
rect 351474 464414 352094 464498
rect 351474 464178 351506 464414
rect 351742 464178 351826 464414
rect 352062 464178 352094 464414
rect 351474 427534 352094 464178
rect 351474 427298 351506 427534
rect 351742 427298 351826 427534
rect 352062 427298 352094 427534
rect 351474 427214 352094 427298
rect 351474 426978 351506 427214
rect 351742 426978 351826 427214
rect 352062 426978 352094 427214
rect 351474 390334 352094 426978
rect 351474 390098 351506 390334
rect 351742 390098 351826 390334
rect 352062 390098 352094 390334
rect 351474 390014 352094 390098
rect 351474 389778 351506 390014
rect 351742 389778 351826 390014
rect 352062 389778 352094 390014
rect 351474 353134 352094 389778
rect 351474 352898 351506 353134
rect 351742 352898 351826 353134
rect 352062 352898 352094 353134
rect 351474 352814 352094 352898
rect 351474 352578 351506 352814
rect 351742 352578 351826 352814
rect 352062 352578 352094 352814
rect 351474 315934 352094 352578
rect 351474 315698 351506 315934
rect 351742 315698 351826 315934
rect 352062 315698 352094 315934
rect 351474 315614 352094 315698
rect 351474 315378 351506 315614
rect 351742 315378 351826 315614
rect 352062 315378 352094 315614
rect 351474 278734 352094 315378
rect 351474 278498 351506 278734
rect 351742 278498 351826 278734
rect 352062 278498 352094 278734
rect 351474 278414 352094 278498
rect 351474 278178 351506 278414
rect 351742 278178 351826 278414
rect 352062 278178 352094 278414
rect 351474 241534 352094 278178
rect 351474 241298 351506 241534
rect 351742 241298 351826 241534
rect 352062 241298 352094 241534
rect 351474 241214 352094 241298
rect 351474 240978 351506 241214
rect 351742 240978 351826 241214
rect 352062 240978 352094 241214
rect 351474 204334 352094 240978
rect 351474 204098 351506 204334
rect 351742 204098 351826 204334
rect 352062 204098 352094 204334
rect 351474 204014 352094 204098
rect 351474 203778 351506 204014
rect 351742 203778 351826 204014
rect 352062 203778 352094 204014
rect 351474 167134 352094 203778
rect 351474 166898 351506 167134
rect 351742 166898 351826 167134
rect 352062 166898 352094 167134
rect 351474 166814 352094 166898
rect 351474 166578 351506 166814
rect 351742 166578 351826 166814
rect 352062 166578 352094 166814
rect 351474 129934 352094 166578
rect 351474 129698 351506 129934
rect 351742 129698 351826 129934
rect 352062 129698 352094 129934
rect 351474 129614 352094 129698
rect 351474 129378 351506 129614
rect 351742 129378 351826 129614
rect 352062 129378 352094 129614
rect 351474 92734 352094 129378
rect 351474 92498 351506 92734
rect 351742 92498 351826 92734
rect 352062 92498 352094 92734
rect 351474 92414 352094 92498
rect 351474 92178 351506 92414
rect 351742 92178 351826 92414
rect 352062 92178 352094 92414
rect 351474 55534 352094 92178
rect 351474 55298 351506 55534
rect 351742 55298 351826 55534
rect 352062 55298 352094 55534
rect 351474 55214 352094 55298
rect 351474 54978 351506 55214
rect 351742 54978 351826 55214
rect 352062 54978 352094 55214
rect 351474 18334 352094 54978
rect 351474 18098 351506 18334
rect 351742 18098 351826 18334
rect 352062 18098 352094 18334
rect 351474 18014 352094 18098
rect 351474 17778 351506 18014
rect 351742 17778 351826 18014
rect 352062 17778 352094 18014
rect 351474 2176 352094 17778
rect 355194 691654 355814 701760
rect 355194 691418 355226 691654
rect 355462 691418 355546 691654
rect 355782 691418 355814 691654
rect 355194 691334 355814 691418
rect 355194 691098 355226 691334
rect 355462 691098 355546 691334
rect 355782 691098 355814 691334
rect 355194 654454 355814 691098
rect 355194 654218 355226 654454
rect 355462 654218 355546 654454
rect 355782 654218 355814 654454
rect 355194 654134 355814 654218
rect 355194 653898 355226 654134
rect 355462 653898 355546 654134
rect 355782 653898 355814 654134
rect 355194 617254 355814 653898
rect 355194 617018 355226 617254
rect 355462 617018 355546 617254
rect 355782 617018 355814 617254
rect 355194 616934 355814 617018
rect 355194 616698 355226 616934
rect 355462 616698 355546 616934
rect 355782 616698 355814 616934
rect 355194 580054 355814 616698
rect 355194 579818 355226 580054
rect 355462 579818 355546 580054
rect 355782 579818 355814 580054
rect 355194 579734 355814 579818
rect 355194 579498 355226 579734
rect 355462 579498 355546 579734
rect 355782 579498 355814 579734
rect 355194 542854 355814 579498
rect 355194 542618 355226 542854
rect 355462 542618 355546 542854
rect 355782 542618 355814 542854
rect 355194 542534 355814 542618
rect 355194 542298 355226 542534
rect 355462 542298 355546 542534
rect 355782 542298 355814 542534
rect 355194 505654 355814 542298
rect 355194 505418 355226 505654
rect 355462 505418 355546 505654
rect 355782 505418 355814 505654
rect 355194 505334 355814 505418
rect 355194 505098 355226 505334
rect 355462 505098 355546 505334
rect 355782 505098 355814 505334
rect 355194 468454 355814 505098
rect 355194 468218 355226 468454
rect 355462 468218 355546 468454
rect 355782 468218 355814 468454
rect 355194 468134 355814 468218
rect 355194 467898 355226 468134
rect 355462 467898 355546 468134
rect 355782 467898 355814 468134
rect 355194 431254 355814 467898
rect 355194 431018 355226 431254
rect 355462 431018 355546 431254
rect 355782 431018 355814 431254
rect 355194 430934 355814 431018
rect 355194 430698 355226 430934
rect 355462 430698 355546 430934
rect 355782 430698 355814 430934
rect 355194 394054 355814 430698
rect 355194 393818 355226 394054
rect 355462 393818 355546 394054
rect 355782 393818 355814 394054
rect 355194 393734 355814 393818
rect 355194 393498 355226 393734
rect 355462 393498 355546 393734
rect 355782 393498 355814 393734
rect 355194 356854 355814 393498
rect 355194 356618 355226 356854
rect 355462 356618 355546 356854
rect 355782 356618 355814 356854
rect 355194 356534 355814 356618
rect 355194 356298 355226 356534
rect 355462 356298 355546 356534
rect 355782 356298 355814 356534
rect 355194 319654 355814 356298
rect 355194 319418 355226 319654
rect 355462 319418 355546 319654
rect 355782 319418 355814 319654
rect 355194 319334 355814 319418
rect 355194 319098 355226 319334
rect 355462 319098 355546 319334
rect 355782 319098 355814 319334
rect 355194 282454 355814 319098
rect 355194 282218 355226 282454
rect 355462 282218 355546 282454
rect 355782 282218 355814 282454
rect 355194 282134 355814 282218
rect 355194 281898 355226 282134
rect 355462 281898 355546 282134
rect 355782 281898 355814 282134
rect 355194 245254 355814 281898
rect 355194 245018 355226 245254
rect 355462 245018 355546 245254
rect 355782 245018 355814 245254
rect 355194 244934 355814 245018
rect 355194 244698 355226 244934
rect 355462 244698 355546 244934
rect 355782 244698 355814 244934
rect 355194 208054 355814 244698
rect 355194 207818 355226 208054
rect 355462 207818 355546 208054
rect 355782 207818 355814 208054
rect 355194 207734 355814 207818
rect 355194 207498 355226 207734
rect 355462 207498 355546 207734
rect 355782 207498 355814 207734
rect 355194 170854 355814 207498
rect 355194 170618 355226 170854
rect 355462 170618 355546 170854
rect 355782 170618 355814 170854
rect 355194 170534 355814 170618
rect 355194 170298 355226 170534
rect 355462 170298 355546 170534
rect 355782 170298 355814 170534
rect 355194 133654 355814 170298
rect 355194 133418 355226 133654
rect 355462 133418 355546 133654
rect 355782 133418 355814 133654
rect 355194 133334 355814 133418
rect 355194 133098 355226 133334
rect 355462 133098 355546 133334
rect 355782 133098 355814 133334
rect 355194 96454 355814 133098
rect 355194 96218 355226 96454
rect 355462 96218 355546 96454
rect 355782 96218 355814 96454
rect 355194 96134 355814 96218
rect 355194 95898 355226 96134
rect 355462 95898 355546 96134
rect 355782 95898 355814 96134
rect 355194 59254 355814 95898
rect 355194 59018 355226 59254
rect 355462 59018 355546 59254
rect 355782 59018 355814 59254
rect 355194 58934 355814 59018
rect 355194 58698 355226 58934
rect 355462 58698 355546 58934
rect 355782 58698 355814 58934
rect 355194 22054 355814 58698
rect 355194 21818 355226 22054
rect 355462 21818 355546 22054
rect 355782 21818 355814 22054
rect 355194 21734 355814 21818
rect 355194 21498 355226 21734
rect 355462 21498 355546 21734
rect 355782 21498 355814 21734
rect 355194 2176 355814 21498
rect 358914 695374 359534 701760
rect 358914 695138 358946 695374
rect 359182 695138 359266 695374
rect 359502 695138 359534 695374
rect 358914 695054 359534 695138
rect 358914 694818 358946 695054
rect 359182 694818 359266 695054
rect 359502 694818 359534 695054
rect 358914 658174 359534 694818
rect 358914 657938 358946 658174
rect 359182 657938 359266 658174
rect 359502 657938 359534 658174
rect 358914 657854 359534 657938
rect 358914 657618 358946 657854
rect 359182 657618 359266 657854
rect 359502 657618 359534 657854
rect 358914 620974 359534 657618
rect 358914 620738 358946 620974
rect 359182 620738 359266 620974
rect 359502 620738 359534 620974
rect 358914 620654 359534 620738
rect 358914 620418 358946 620654
rect 359182 620418 359266 620654
rect 359502 620418 359534 620654
rect 358914 583774 359534 620418
rect 358914 583538 358946 583774
rect 359182 583538 359266 583774
rect 359502 583538 359534 583774
rect 358914 583454 359534 583538
rect 358914 583218 358946 583454
rect 359182 583218 359266 583454
rect 359502 583218 359534 583454
rect 358914 546574 359534 583218
rect 358914 546338 358946 546574
rect 359182 546338 359266 546574
rect 359502 546338 359534 546574
rect 358914 546254 359534 546338
rect 358914 546018 358946 546254
rect 359182 546018 359266 546254
rect 359502 546018 359534 546254
rect 358914 509374 359534 546018
rect 358914 509138 358946 509374
rect 359182 509138 359266 509374
rect 359502 509138 359534 509374
rect 358914 509054 359534 509138
rect 358914 508818 358946 509054
rect 359182 508818 359266 509054
rect 359502 508818 359534 509054
rect 358914 472174 359534 508818
rect 358914 471938 358946 472174
rect 359182 471938 359266 472174
rect 359502 471938 359534 472174
rect 358914 471854 359534 471938
rect 358914 471618 358946 471854
rect 359182 471618 359266 471854
rect 359502 471618 359534 471854
rect 358914 434974 359534 471618
rect 358914 434738 358946 434974
rect 359182 434738 359266 434974
rect 359502 434738 359534 434974
rect 358914 434654 359534 434738
rect 358914 434418 358946 434654
rect 359182 434418 359266 434654
rect 359502 434418 359534 434654
rect 358914 397774 359534 434418
rect 358914 397538 358946 397774
rect 359182 397538 359266 397774
rect 359502 397538 359534 397774
rect 358914 397454 359534 397538
rect 358914 397218 358946 397454
rect 359182 397218 359266 397454
rect 359502 397218 359534 397454
rect 358914 360574 359534 397218
rect 358914 360338 358946 360574
rect 359182 360338 359266 360574
rect 359502 360338 359534 360574
rect 358914 360254 359534 360338
rect 358914 360018 358946 360254
rect 359182 360018 359266 360254
rect 359502 360018 359534 360254
rect 358914 323374 359534 360018
rect 358914 323138 358946 323374
rect 359182 323138 359266 323374
rect 359502 323138 359534 323374
rect 358914 323054 359534 323138
rect 358914 322818 358946 323054
rect 359182 322818 359266 323054
rect 359502 322818 359534 323054
rect 358914 286174 359534 322818
rect 358914 285938 358946 286174
rect 359182 285938 359266 286174
rect 359502 285938 359534 286174
rect 358914 285854 359534 285938
rect 358914 285618 358946 285854
rect 359182 285618 359266 285854
rect 359502 285618 359534 285854
rect 358914 248974 359534 285618
rect 358914 248738 358946 248974
rect 359182 248738 359266 248974
rect 359502 248738 359534 248974
rect 358914 248654 359534 248738
rect 358914 248418 358946 248654
rect 359182 248418 359266 248654
rect 359502 248418 359534 248654
rect 358914 211774 359534 248418
rect 358914 211538 358946 211774
rect 359182 211538 359266 211774
rect 359502 211538 359534 211774
rect 358914 211454 359534 211538
rect 358914 211218 358946 211454
rect 359182 211218 359266 211454
rect 359502 211218 359534 211454
rect 358914 174574 359534 211218
rect 358914 174338 358946 174574
rect 359182 174338 359266 174574
rect 359502 174338 359534 174574
rect 358914 174254 359534 174338
rect 358914 174018 358946 174254
rect 359182 174018 359266 174254
rect 359502 174018 359534 174254
rect 358914 137374 359534 174018
rect 358914 137138 358946 137374
rect 359182 137138 359266 137374
rect 359502 137138 359534 137374
rect 358914 137054 359534 137138
rect 358914 136818 358946 137054
rect 359182 136818 359266 137054
rect 359502 136818 359534 137054
rect 358914 100174 359534 136818
rect 358914 99938 358946 100174
rect 359182 99938 359266 100174
rect 359502 99938 359534 100174
rect 358914 99854 359534 99938
rect 358914 99618 358946 99854
rect 359182 99618 359266 99854
rect 359502 99618 359534 99854
rect 358914 62974 359534 99618
rect 358914 62738 358946 62974
rect 359182 62738 359266 62974
rect 359502 62738 359534 62974
rect 358914 62654 359534 62738
rect 358914 62418 358946 62654
rect 359182 62418 359266 62654
rect 359502 62418 359534 62654
rect 358914 25774 359534 62418
rect 358914 25538 358946 25774
rect 359182 25538 359266 25774
rect 359502 25538 359534 25774
rect 358914 25454 359534 25538
rect 358914 25218 358946 25454
rect 359182 25218 359266 25454
rect 359502 25218 359534 25454
rect 358914 2176 359534 25218
rect 362634 699094 363254 701760
rect 362634 698858 362666 699094
rect 362902 698858 362986 699094
rect 363222 698858 363254 699094
rect 362634 698774 363254 698858
rect 362634 698538 362666 698774
rect 362902 698538 362986 698774
rect 363222 698538 363254 698774
rect 362634 661894 363254 698538
rect 362634 661658 362666 661894
rect 362902 661658 362986 661894
rect 363222 661658 363254 661894
rect 362634 661574 363254 661658
rect 362634 661338 362666 661574
rect 362902 661338 362986 661574
rect 363222 661338 363254 661574
rect 362634 624694 363254 661338
rect 362634 624458 362666 624694
rect 362902 624458 362986 624694
rect 363222 624458 363254 624694
rect 362634 624374 363254 624458
rect 362634 624138 362666 624374
rect 362902 624138 362986 624374
rect 363222 624138 363254 624374
rect 362634 587494 363254 624138
rect 362634 587258 362666 587494
rect 362902 587258 362986 587494
rect 363222 587258 363254 587494
rect 362634 587174 363254 587258
rect 362634 586938 362666 587174
rect 362902 586938 362986 587174
rect 363222 586938 363254 587174
rect 362634 550294 363254 586938
rect 362634 550058 362666 550294
rect 362902 550058 362986 550294
rect 363222 550058 363254 550294
rect 362634 549974 363254 550058
rect 362634 549738 362666 549974
rect 362902 549738 362986 549974
rect 363222 549738 363254 549974
rect 362634 513094 363254 549738
rect 362634 512858 362666 513094
rect 362902 512858 362986 513094
rect 363222 512858 363254 513094
rect 362634 512774 363254 512858
rect 362634 512538 362666 512774
rect 362902 512538 362986 512774
rect 363222 512538 363254 512774
rect 362634 475894 363254 512538
rect 362634 475658 362666 475894
rect 362902 475658 362986 475894
rect 363222 475658 363254 475894
rect 362634 475574 363254 475658
rect 362634 475338 362666 475574
rect 362902 475338 362986 475574
rect 363222 475338 363254 475574
rect 362634 438694 363254 475338
rect 362634 438458 362666 438694
rect 362902 438458 362986 438694
rect 363222 438458 363254 438694
rect 362634 438374 363254 438458
rect 362634 438138 362666 438374
rect 362902 438138 362986 438374
rect 363222 438138 363254 438374
rect 362634 401494 363254 438138
rect 362634 401258 362666 401494
rect 362902 401258 362986 401494
rect 363222 401258 363254 401494
rect 362634 401174 363254 401258
rect 362634 400938 362666 401174
rect 362902 400938 362986 401174
rect 363222 400938 363254 401174
rect 362634 364294 363254 400938
rect 362634 364058 362666 364294
rect 362902 364058 362986 364294
rect 363222 364058 363254 364294
rect 362634 363974 363254 364058
rect 362634 363738 362666 363974
rect 362902 363738 362986 363974
rect 363222 363738 363254 363974
rect 362634 327094 363254 363738
rect 362634 326858 362666 327094
rect 362902 326858 362986 327094
rect 363222 326858 363254 327094
rect 362634 326774 363254 326858
rect 362634 326538 362666 326774
rect 362902 326538 362986 326774
rect 363222 326538 363254 326774
rect 362634 289894 363254 326538
rect 362634 289658 362666 289894
rect 362902 289658 362986 289894
rect 363222 289658 363254 289894
rect 362634 289574 363254 289658
rect 362634 289338 362666 289574
rect 362902 289338 362986 289574
rect 363222 289338 363254 289574
rect 362634 252694 363254 289338
rect 362634 252458 362666 252694
rect 362902 252458 362986 252694
rect 363222 252458 363254 252694
rect 362634 252374 363254 252458
rect 362634 252138 362666 252374
rect 362902 252138 362986 252374
rect 363222 252138 363254 252374
rect 362634 215494 363254 252138
rect 362634 215258 362666 215494
rect 362902 215258 362986 215494
rect 363222 215258 363254 215494
rect 362634 215174 363254 215258
rect 362634 214938 362666 215174
rect 362902 214938 362986 215174
rect 363222 214938 363254 215174
rect 362634 178294 363254 214938
rect 362634 178058 362666 178294
rect 362902 178058 362986 178294
rect 363222 178058 363254 178294
rect 362634 177974 363254 178058
rect 362634 177738 362666 177974
rect 362902 177738 362986 177974
rect 363222 177738 363254 177974
rect 362634 141094 363254 177738
rect 362634 140858 362666 141094
rect 362902 140858 362986 141094
rect 363222 140858 363254 141094
rect 362634 140774 363254 140858
rect 362634 140538 362666 140774
rect 362902 140538 362986 140774
rect 363222 140538 363254 140774
rect 362634 103894 363254 140538
rect 362634 103658 362666 103894
rect 362902 103658 362986 103894
rect 363222 103658 363254 103894
rect 362634 103574 363254 103658
rect 362634 103338 362666 103574
rect 362902 103338 362986 103574
rect 363222 103338 363254 103574
rect 362634 66694 363254 103338
rect 362634 66458 362666 66694
rect 362902 66458 362986 66694
rect 363222 66458 363254 66694
rect 362634 66374 363254 66458
rect 362634 66138 362666 66374
rect 362902 66138 362986 66374
rect 363222 66138 363254 66374
rect 362634 29494 363254 66138
rect 362634 29258 362666 29494
rect 362902 29258 362986 29494
rect 363222 29258 363254 29494
rect 362634 29174 363254 29258
rect 362634 28938 362666 29174
rect 362902 28938 362986 29174
rect 363222 28938 363254 29174
rect 362634 2176 363254 28938
rect 373794 673054 374414 701760
rect 373794 672818 373826 673054
rect 374062 672818 374146 673054
rect 374382 672818 374414 673054
rect 373794 672734 374414 672818
rect 373794 672498 373826 672734
rect 374062 672498 374146 672734
rect 374382 672498 374414 672734
rect 373794 635854 374414 672498
rect 373794 635618 373826 635854
rect 374062 635618 374146 635854
rect 374382 635618 374414 635854
rect 373794 635534 374414 635618
rect 373794 635298 373826 635534
rect 374062 635298 374146 635534
rect 374382 635298 374414 635534
rect 373794 598654 374414 635298
rect 373794 598418 373826 598654
rect 374062 598418 374146 598654
rect 374382 598418 374414 598654
rect 373794 598334 374414 598418
rect 373794 598098 373826 598334
rect 374062 598098 374146 598334
rect 374382 598098 374414 598334
rect 373794 561454 374414 598098
rect 373794 561218 373826 561454
rect 374062 561218 374146 561454
rect 374382 561218 374414 561454
rect 373794 561134 374414 561218
rect 373794 560898 373826 561134
rect 374062 560898 374146 561134
rect 374382 560898 374414 561134
rect 373794 524254 374414 560898
rect 373794 524018 373826 524254
rect 374062 524018 374146 524254
rect 374382 524018 374414 524254
rect 373794 523934 374414 524018
rect 373794 523698 373826 523934
rect 374062 523698 374146 523934
rect 374382 523698 374414 523934
rect 373794 487054 374414 523698
rect 373794 486818 373826 487054
rect 374062 486818 374146 487054
rect 374382 486818 374414 487054
rect 373794 486734 374414 486818
rect 373794 486498 373826 486734
rect 374062 486498 374146 486734
rect 374382 486498 374414 486734
rect 373794 449854 374414 486498
rect 373794 449618 373826 449854
rect 374062 449618 374146 449854
rect 374382 449618 374414 449854
rect 373794 449534 374414 449618
rect 373794 449298 373826 449534
rect 374062 449298 374146 449534
rect 374382 449298 374414 449534
rect 373794 412654 374414 449298
rect 373794 412418 373826 412654
rect 374062 412418 374146 412654
rect 374382 412418 374414 412654
rect 373794 412334 374414 412418
rect 373794 412098 373826 412334
rect 374062 412098 374146 412334
rect 374382 412098 374414 412334
rect 373794 375454 374414 412098
rect 373794 375218 373826 375454
rect 374062 375218 374146 375454
rect 374382 375218 374414 375454
rect 373794 375134 374414 375218
rect 373794 374898 373826 375134
rect 374062 374898 374146 375134
rect 374382 374898 374414 375134
rect 373794 338254 374414 374898
rect 373794 338018 373826 338254
rect 374062 338018 374146 338254
rect 374382 338018 374414 338254
rect 373794 337934 374414 338018
rect 373794 337698 373826 337934
rect 374062 337698 374146 337934
rect 374382 337698 374414 337934
rect 373794 301054 374414 337698
rect 373794 300818 373826 301054
rect 374062 300818 374146 301054
rect 374382 300818 374414 301054
rect 373794 300734 374414 300818
rect 373794 300498 373826 300734
rect 374062 300498 374146 300734
rect 374382 300498 374414 300734
rect 373794 263854 374414 300498
rect 373794 263618 373826 263854
rect 374062 263618 374146 263854
rect 374382 263618 374414 263854
rect 373794 263534 374414 263618
rect 373794 263298 373826 263534
rect 374062 263298 374146 263534
rect 374382 263298 374414 263534
rect 373794 226654 374414 263298
rect 373794 226418 373826 226654
rect 374062 226418 374146 226654
rect 374382 226418 374414 226654
rect 373794 226334 374414 226418
rect 373794 226098 373826 226334
rect 374062 226098 374146 226334
rect 374382 226098 374414 226334
rect 373794 189454 374414 226098
rect 373794 189218 373826 189454
rect 374062 189218 374146 189454
rect 374382 189218 374414 189454
rect 373794 189134 374414 189218
rect 373794 188898 373826 189134
rect 374062 188898 374146 189134
rect 374382 188898 374414 189134
rect 373794 152254 374414 188898
rect 373794 152018 373826 152254
rect 374062 152018 374146 152254
rect 374382 152018 374414 152254
rect 373794 151934 374414 152018
rect 373794 151698 373826 151934
rect 374062 151698 374146 151934
rect 374382 151698 374414 151934
rect 373794 115054 374414 151698
rect 373794 114818 373826 115054
rect 374062 114818 374146 115054
rect 374382 114818 374414 115054
rect 373794 114734 374414 114818
rect 373794 114498 373826 114734
rect 374062 114498 374146 114734
rect 374382 114498 374414 114734
rect 373794 77854 374414 114498
rect 373794 77618 373826 77854
rect 374062 77618 374146 77854
rect 374382 77618 374414 77854
rect 373794 77534 374414 77618
rect 373794 77298 373826 77534
rect 374062 77298 374146 77534
rect 374382 77298 374414 77534
rect 373794 40654 374414 77298
rect 373794 40418 373826 40654
rect 374062 40418 374146 40654
rect 374382 40418 374414 40654
rect 373794 40334 374414 40418
rect 373794 40098 373826 40334
rect 374062 40098 374146 40334
rect 374382 40098 374414 40334
rect 373794 3454 374414 40098
rect 373794 3218 373826 3454
rect 374062 3218 374146 3454
rect 374382 3218 374414 3454
rect 373794 3134 374414 3218
rect 373794 2898 373826 3134
rect 374062 2898 374146 3134
rect 374382 2898 374414 3134
rect 373794 2176 374414 2898
rect 377514 676774 378134 701760
rect 377514 676538 377546 676774
rect 377782 676538 377866 676774
rect 378102 676538 378134 676774
rect 377514 676454 378134 676538
rect 377514 676218 377546 676454
rect 377782 676218 377866 676454
rect 378102 676218 378134 676454
rect 377514 639574 378134 676218
rect 377514 639338 377546 639574
rect 377782 639338 377866 639574
rect 378102 639338 378134 639574
rect 377514 639254 378134 639338
rect 377514 639018 377546 639254
rect 377782 639018 377866 639254
rect 378102 639018 378134 639254
rect 377514 602374 378134 639018
rect 377514 602138 377546 602374
rect 377782 602138 377866 602374
rect 378102 602138 378134 602374
rect 377514 602054 378134 602138
rect 377514 601818 377546 602054
rect 377782 601818 377866 602054
rect 378102 601818 378134 602054
rect 377514 565174 378134 601818
rect 377514 564938 377546 565174
rect 377782 564938 377866 565174
rect 378102 564938 378134 565174
rect 377514 564854 378134 564938
rect 377514 564618 377546 564854
rect 377782 564618 377866 564854
rect 378102 564618 378134 564854
rect 377514 527974 378134 564618
rect 377514 527738 377546 527974
rect 377782 527738 377866 527974
rect 378102 527738 378134 527974
rect 377514 527654 378134 527738
rect 377514 527418 377546 527654
rect 377782 527418 377866 527654
rect 378102 527418 378134 527654
rect 377514 490774 378134 527418
rect 377514 490538 377546 490774
rect 377782 490538 377866 490774
rect 378102 490538 378134 490774
rect 377514 490454 378134 490538
rect 377514 490218 377546 490454
rect 377782 490218 377866 490454
rect 378102 490218 378134 490454
rect 377514 453574 378134 490218
rect 377514 453338 377546 453574
rect 377782 453338 377866 453574
rect 378102 453338 378134 453574
rect 377514 453254 378134 453338
rect 377514 453018 377546 453254
rect 377782 453018 377866 453254
rect 378102 453018 378134 453254
rect 377514 416374 378134 453018
rect 377514 416138 377546 416374
rect 377782 416138 377866 416374
rect 378102 416138 378134 416374
rect 377514 416054 378134 416138
rect 377514 415818 377546 416054
rect 377782 415818 377866 416054
rect 378102 415818 378134 416054
rect 377514 379174 378134 415818
rect 377514 378938 377546 379174
rect 377782 378938 377866 379174
rect 378102 378938 378134 379174
rect 377514 378854 378134 378938
rect 377514 378618 377546 378854
rect 377782 378618 377866 378854
rect 378102 378618 378134 378854
rect 377514 341974 378134 378618
rect 377514 341738 377546 341974
rect 377782 341738 377866 341974
rect 378102 341738 378134 341974
rect 377514 341654 378134 341738
rect 377514 341418 377546 341654
rect 377782 341418 377866 341654
rect 378102 341418 378134 341654
rect 377514 304774 378134 341418
rect 377514 304538 377546 304774
rect 377782 304538 377866 304774
rect 378102 304538 378134 304774
rect 377514 304454 378134 304538
rect 377514 304218 377546 304454
rect 377782 304218 377866 304454
rect 378102 304218 378134 304454
rect 377514 267574 378134 304218
rect 377514 267338 377546 267574
rect 377782 267338 377866 267574
rect 378102 267338 378134 267574
rect 377514 267254 378134 267338
rect 377514 267018 377546 267254
rect 377782 267018 377866 267254
rect 378102 267018 378134 267254
rect 377514 230374 378134 267018
rect 377514 230138 377546 230374
rect 377782 230138 377866 230374
rect 378102 230138 378134 230374
rect 377514 230054 378134 230138
rect 377514 229818 377546 230054
rect 377782 229818 377866 230054
rect 378102 229818 378134 230054
rect 377514 193174 378134 229818
rect 377514 192938 377546 193174
rect 377782 192938 377866 193174
rect 378102 192938 378134 193174
rect 377514 192854 378134 192938
rect 377514 192618 377546 192854
rect 377782 192618 377866 192854
rect 378102 192618 378134 192854
rect 377514 155974 378134 192618
rect 377514 155738 377546 155974
rect 377782 155738 377866 155974
rect 378102 155738 378134 155974
rect 377514 155654 378134 155738
rect 377514 155418 377546 155654
rect 377782 155418 377866 155654
rect 378102 155418 378134 155654
rect 377514 118774 378134 155418
rect 377514 118538 377546 118774
rect 377782 118538 377866 118774
rect 378102 118538 378134 118774
rect 377514 118454 378134 118538
rect 377514 118218 377546 118454
rect 377782 118218 377866 118454
rect 378102 118218 378134 118454
rect 377514 81574 378134 118218
rect 377514 81338 377546 81574
rect 377782 81338 377866 81574
rect 378102 81338 378134 81574
rect 377514 81254 378134 81338
rect 377514 81018 377546 81254
rect 377782 81018 377866 81254
rect 378102 81018 378134 81254
rect 377514 44374 378134 81018
rect 377514 44138 377546 44374
rect 377782 44138 377866 44374
rect 378102 44138 378134 44374
rect 377514 44054 378134 44138
rect 377514 43818 377546 44054
rect 377782 43818 377866 44054
rect 378102 43818 378134 44054
rect 377514 7174 378134 43818
rect 377514 6938 377546 7174
rect 377782 6938 377866 7174
rect 378102 6938 378134 7174
rect 377514 6854 378134 6938
rect 377514 6618 377546 6854
rect 377782 6618 377866 6854
rect 378102 6618 378134 6854
rect 377514 2176 378134 6618
rect 381234 680494 381854 701760
rect 381234 680258 381266 680494
rect 381502 680258 381586 680494
rect 381822 680258 381854 680494
rect 381234 680174 381854 680258
rect 381234 679938 381266 680174
rect 381502 679938 381586 680174
rect 381822 679938 381854 680174
rect 381234 643294 381854 679938
rect 381234 643058 381266 643294
rect 381502 643058 381586 643294
rect 381822 643058 381854 643294
rect 381234 642974 381854 643058
rect 381234 642738 381266 642974
rect 381502 642738 381586 642974
rect 381822 642738 381854 642974
rect 381234 606094 381854 642738
rect 381234 605858 381266 606094
rect 381502 605858 381586 606094
rect 381822 605858 381854 606094
rect 381234 605774 381854 605858
rect 381234 605538 381266 605774
rect 381502 605538 381586 605774
rect 381822 605538 381854 605774
rect 381234 568894 381854 605538
rect 381234 568658 381266 568894
rect 381502 568658 381586 568894
rect 381822 568658 381854 568894
rect 381234 568574 381854 568658
rect 381234 568338 381266 568574
rect 381502 568338 381586 568574
rect 381822 568338 381854 568574
rect 381234 531694 381854 568338
rect 381234 531458 381266 531694
rect 381502 531458 381586 531694
rect 381822 531458 381854 531694
rect 381234 531374 381854 531458
rect 381234 531138 381266 531374
rect 381502 531138 381586 531374
rect 381822 531138 381854 531374
rect 381234 494494 381854 531138
rect 381234 494258 381266 494494
rect 381502 494258 381586 494494
rect 381822 494258 381854 494494
rect 381234 494174 381854 494258
rect 381234 493938 381266 494174
rect 381502 493938 381586 494174
rect 381822 493938 381854 494174
rect 381234 457294 381854 493938
rect 381234 457058 381266 457294
rect 381502 457058 381586 457294
rect 381822 457058 381854 457294
rect 381234 456974 381854 457058
rect 381234 456738 381266 456974
rect 381502 456738 381586 456974
rect 381822 456738 381854 456974
rect 381234 420094 381854 456738
rect 381234 419858 381266 420094
rect 381502 419858 381586 420094
rect 381822 419858 381854 420094
rect 381234 419774 381854 419858
rect 381234 419538 381266 419774
rect 381502 419538 381586 419774
rect 381822 419538 381854 419774
rect 381234 382894 381854 419538
rect 381234 382658 381266 382894
rect 381502 382658 381586 382894
rect 381822 382658 381854 382894
rect 381234 382574 381854 382658
rect 381234 382338 381266 382574
rect 381502 382338 381586 382574
rect 381822 382338 381854 382574
rect 381234 345694 381854 382338
rect 381234 345458 381266 345694
rect 381502 345458 381586 345694
rect 381822 345458 381854 345694
rect 381234 345374 381854 345458
rect 381234 345138 381266 345374
rect 381502 345138 381586 345374
rect 381822 345138 381854 345374
rect 381234 308494 381854 345138
rect 381234 308258 381266 308494
rect 381502 308258 381586 308494
rect 381822 308258 381854 308494
rect 381234 308174 381854 308258
rect 381234 307938 381266 308174
rect 381502 307938 381586 308174
rect 381822 307938 381854 308174
rect 381234 271294 381854 307938
rect 381234 271058 381266 271294
rect 381502 271058 381586 271294
rect 381822 271058 381854 271294
rect 381234 270974 381854 271058
rect 381234 270738 381266 270974
rect 381502 270738 381586 270974
rect 381822 270738 381854 270974
rect 381234 234094 381854 270738
rect 381234 233858 381266 234094
rect 381502 233858 381586 234094
rect 381822 233858 381854 234094
rect 381234 233774 381854 233858
rect 381234 233538 381266 233774
rect 381502 233538 381586 233774
rect 381822 233538 381854 233774
rect 381234 196894 381854 233538
rect 381234 196658 381266 196894
rect 381502 196658 381586 196894
rect 381822 196658 381854 196894
rect 381234 196574 381854 196658
rect 381234 196338 381266 196574
rect 381502 196338 381586 196574
rect 381822 196338 381854 196574
rect 381234 159694 381854 196338
rect 381234 159458 381266 159694
rect 381502 159458 381586 159694
rect 381822 159458 381854 159694
rect 381234 159374 381854 159458
rect 381234 159138 381266 159374
rect 381502 159138 381586 159374
rect 381822 159138 381854 159374
rect 381234 122494 381854 159138
rect 381234 122258 381266 122494
rect 381502 122258 381586 122494
rect 381822 122258 381854 122494
rect 381234 122174 381854 122258
rect 381234 121938 381266 122174
rect 381502 121938 381586 122174
rect 381822 121938 381854 122174
rect 381234 85294 381854 121938
rect 381234 85058 381266 85294
rect 381502 85058 381586 85294
rect 381822 85058 381854 85294
rect 381234 84974 381854 85058
rect 381234 84738 381266 84974
rect 381502 84738 381586 84974
rect 381822 84738 381854 84974
rect 381234 48094 381854 84738
rect 381234 47858 381266 48094
rect 381502 47858 381586 48094
rect 381822 47858 381854 48094
rect 381234 47774 381854 47858
rect 381234 47538 381266 47774
rect 381502 47538 381586 47774
rect 381822 47538 381854 47774
rect 381234 10894 381854 47538
rect 381234 10658 381266 10894
rect 381502 10658 381586 10894
rect 381822 10658 381854 10894
rect 381234 10574 381854 10658
rect 381234 10338 381266 10574
rect 381502 10338 381586 10574
rect 381822 10338 381854 10574
rect 381234 2176 381854 10338
rect 384954 684214 385574 701760
rect 384954 683978 384986 684214
rect 385222 683978 385306 684214
rect 385542 683978 385574 684214
rect 384954 683894 385574 683978
rect 384954 683658 384986 683894
rect 385222 683658 385306 683894
rect 385542 683658 385574 683894
rect 384954 647014 385574 683658
rect 384954 646778 384986 647014
rect 385222 646778 385306 647014
rect 385542 646778 385574 647014
rect 384954 646694 385574 646778
rect 384954 646458 384986 646694
rect 385222 646458 385306 646694
rect 385542 646458 385574 646694
rect 384954 609814 385574 646458
rect 384954 609578 384986 609814
rect 385222 609578 385306 609814
rect 385542 609578 385574 609814
rect 384954 609494 385574 609578
rect 384954 609258 384986 609494
rect 385222 609258 385306 609494
rect 385542 609258 385574 609494
rect 384954 572614 385574 609258
rect 384954 572378 384986 572614
rect 385222 572378 385306 572614
rect 385542 572378 385574 572614
rect 384954 572294 385574 572378
rect 384954 572058 384986 572294
rect 385222 572058 385306 572294
rect 385542 572058 385574 572294
rect 384954 535414 385574 572058
rect 384954 535178 384986 535414
rect 385222 535178 385306 535414
rect 385542 535178 385574 535414
rect 384954 535094 385574 535178
rect 384954 534858 384986 535094
rect 385222 534858 385306 535094
rect 385542 534858 385574 535094
rect 384954 498214 385574 534858
rect 384954 497978 384986 498214
rect 385222 497978 385306 498214
rect 385542 497978 385574 498214
rect 384954 497894 385574 497978
rect 384954 497658 384986 497894
rect 385222 497658 385306 497894
rect 385542 497658 385574 497894
rect 384954 461014 385574 497658
rect 384954 460778 384986 461014
rect 385222 460778 385306 461014
rect 385542 460778 385574 461014
rect 384954 460694 385574 460778
rect 384954 460458 384986 460694
rect 385222 460458 385306 460694
rect 385542 460458 385574 460694
rect 384954 423814 385574 460458
rect 384954 423578 384986 423814
rect 385222 423578 385306 423814
rect 385542 423578 385574 423814
rect 384954 423494 385574 423578
rect 384954 423258 384986 423494
rect 385222 423258 385306 423494
rect 385542 423258 385574 423494
rect 384954 386614 385574 423258
rect 384954 386378 384986 386614
rect 385222 386378 385306 386614
rect 385542 386378 385574 386614
rect 384954 386294 385574 386378
rect 384954 386058 384986 386294
rect 385222 386058 385306 386294
rect 385542 386058 385574 386294
rect 384954 349414 385574 386058
rect 384954 349178 384986 349414
rect 385222 349178 385306 349414
rect 385542 349178 385574 349414
rect 384954 349094 385574 349178
rect 384954 348858 384986 349094
rect 385222 348858 385306 349094
rect 385542 348858 385574 349094
rect 384954 312214 385574 348858
rect 384954 311978 384986 312214
rect 385222 311978 385306 312214
rect 385542 311978 385574 312214
rect 384954 311894 385574 311978
rect 384954 311658 384986 311894
rect 385222 311658 385306 311894
rect 385542 311658 385574 311894
rect 384954 275014 385574 311658
rect 384954 274778 384986 275014
rect 385222 274778 385306 275014
rect 385542 274778 385574 275014
rect 384954 274694 385574 274778
rect 384954 274458 384986 274694
rect 385222 274458 385306 274694
rect 385542 274458 385574 274694
rect 384954 237814 385574 274458
rect 384954 237578 384986 237814
rect 385222 237578 385306 237814
rect 385542 237578 385574 237814
rect 384954 237494 385574 237578
rect 384954 237258 384986 237494
rect 385222 237258 385306 237494
rect 385542 237258 385574 237494
rect 384954 200614 385574 237258
rect 384954 200378 384986 200614
rect 385222 200378 385306 200614
rect 385542 200378 385574 200614
rect 384954 200294 385574 200378
rect 384954 200058 384986 200294
rect 385222 200058 385306 200294
rect 385542 200058 385574 200294
rect 384954 163414 385574 200058
rect 384954 163178 384986 163414
rect 385222 163178 385306 163414
rect 385542 163178 385574 163414
rect 384954 163094 385574 163178
rect 384954 162858 384986 163094
rect 385222 162858 385306 163094
rect 385542 162858 385574 163094
rect 384954 126214 385574 162858
rect 384954 125978 384986 126214
rect 385222 125978 385306 126214
rect 385542 125978 385574 126214
rect 384954 125894 385574 125978
rect 384954 125658 384986 125894
rect 385222 125658 385306 125894
rect 385542 125658 385574 125894
rect 384954 89014 385574 125658
rect 384954 88778 384986 89014
rect 385222 88778 385306 89014
rect 385542 88778 385574 89014
rect 384954 88694 385574 88778
rect 384954 88458 384986 88694
rect 385222 88458 385306 88694
rect 385542 88458 385574 88694
rect 384954 51814 385574 88458
rect 384954 51578 384986 51814
rect 385222 51578 385306 51814
rect 385542 51578 385574 51814
rect 384954 51494 385574 51578
rect 384954 51258 384986 51494
rect 385222 51258 385306 51494
rect 385542 51258 385574 51494
rect 384954 14614 385574 51258
rect 384954 14378 384986 14614
rect 385222 14378 385306 14614
rect 385542 14378 385574 14614
rect 384954 14294 385574 14378
rect 384954 14058 384986 14294
rect 385222 14058 385306 14294
rect 385542 14058 385574 14294
rect 384954 2176 385574 14058
rect 388674 687934 389294 701760
rect 388674 687698 388706 687934
rect 388942 687698 389026 687934
rect 389262 687698 389294 687934
rect 388674 687614 389294 687698
rect 388674 687378 388706 687614
rect 388942 687378 389026 687614
rect 389262 687378 389294 687614
rect 388674 650734 389294 687378
rect 388674 650498 388706 650734
rect 388942 650498 389026 650734
rect 389262 650498 389294 650734
rect 388674 650414 389294 650498
rect 388674 650178 388706 650414
rect 388942 650178 389026 650414
rect 389262 650178 389294 650414
rect 388674 613534 389294 650178
rect 388674 613298 388706 613534
rect 388942 613298 389026 613534
rect 389262 613298 389294 613534
rect 388674 613214 389294 613298
rect 388674 612978 388706 613214
rect 388942 612978 389026 613214
rect 389262 612978 389294 613214
rect 388674 576334 389294 612978
rect 388674 576098 388706 576334
rect 388942 576098 389026 576334
rect 389262 576098 389294 576334
rect 388674 576014 389294 576098
rect 388674 575778 388706 576014
rect 388942 575778 389026 576014
rect 389262 575778 389294 576014
rect 388674 539134 389294 575778
rect 388674 538898 388706 539134
rect 388942 538898 389026 539134
rect 389262 538898 389294 539134
rect 388674 538814 389294 538898
rect 388674 538578 388706 538814
rect 388942 538578 389026 538814
rect 389262 538578 389294 538814
rect 388674 501934 389294 538578
rect 388674 501698 388706 501934
rect 388942 501698 389026 501934
rect 389262 501698 389294 501934
rect 388674 501614 389294 501698
rect 388674 501378 388706 501614
rect 388942 501378 389026 501614
rect 389262 501378 389294 501614
rect 388674 464734 389294 501378
rect 388674 464498 388706 464734
rect 388942 464498 389026 464734
rect 389262 464498 389294 464734
rect 388674 464414 389294 464498
rect 388674 464178 388706 464414
rect 388942 464178 389026 464414
rect 389262 464178 389294 464414
rect 388674 427534 389294 464178
rect 388674 427298 388706 427534
rect 388942 427298 389026 427534
rect 389262 427298 389294 427534
rect 388674 427214 389294 427298
rect 388674 426978 388706 427214
rect 388942 426978 389026 427214
rect 389262 426978 389294 427214
rect 388674 390334 389294 426978
rect 388674 390098 388706 390334
rect 388942 390098 389026 390334
rect 389262 390098 389294 390334
rect 388674 390014 389294 390098
rect 388674 389778 388706 390014
rect 388942 389778 389026 390014
rect 389262 389778 389294 390014
rect 388674 353134 389294 389778
rect 388674 352898 388706 353134
rect 388942 352898 389026 353134
rect 389262 352898 389294 353134
rect 388674 352814 389294 352898
rect 388674 352578 388706 352814
rect 388942 352578 389026 352814
rect 389262 352578 389294 352814
rect 388674 315934 389294 352578
rect 388674 315698 388706 315934
rect 388942 315698 389026 315934
rect 389262 315698 389294 315934
rect 388674 315614 389294 315698
rect 388674 315378 388706 315614
rect 388942 315378 389026 315614
rect 389262 315378 389294 315614
rect 388674 278734 389294 315378
rect 388674 278498 388706 278734
rect 388942 278498 389026 278734
rect 389262 278498 389294 278734
rect 388674 278414 389294 278498
rect 388674 278178 388706 278414
rect 388942 278178 389026 278414
rect 389262 278178 389294 278414
rect 388674 241534 389294 278178
rect 388674 241298 388706 241534
rect 388942 241298 389026 241534
rect 389262 241298 389294 241534
rect 388674 241214 389294 241298
rect 388674 240978 388706 241214
rect 388942 240978 389026 241214
rect 389262 240978 389294 241214
rect 388674 204334 389294 240978
rect 388674 204098 388706 204334
rect 388942 204098 389026 204334
rect 389262 204098 389294 204334
rect 388674 204014 389294 204098
rect 388674 203778 388706 204014
rect 388942 203778 389026 204014
rect 389262 203778 389294 204014
rect 388674 167134 389294 203778
rect 388674 166898 388706 167134
rect 388942 166898 389026 167134
rect 389262 166898 389294 167134
rect 388674 166814 389294 166898
rect 388674 166578 388706 166814
rect 388942 166578 389026 166814
rect 389262 166578 389294 166814
rect 388674 129934 389294 166578
rect 388674 129698 388706 129934
rect 388942 129698 389026 129934
rect 389262 129698 389294 129934
rect 388674 129614 389294 129698
rect 388674 129378 388706 129614
rect 388942 129378 389026 129614
rect 389262 129378 389294 129614
rect 388674 92734 389294 129378
rect 388674 92498 388706 92734
rect 388942 92498 389026 92734
rect 389262 92498 389294 92734
rect 388674 92414 389294 92498
rect 388674 92178 388706 92414
rect 388942 92178 389026 92414
rect 389262 92178 389294 92414
rect 388674 55534 389294 92178
rect 388674 55298 388706 55534
rect 388942 55298 389026 55534
rect 389262 55298 389294 55534
rect 388674 55214 389294 55298
rect 388674 54978 388706 55214
rect 388942 54978 389026 55214
rect 389262 54978 389294 55214
rect 388674 18334 389294 54978
rect 388674 18098 388706 18334
rect 388942 18098 389026 18334
rect 389262 18098 389294 18334
rect 388674 18014 389294 18098
rect 388674 17778 388706 18014
rect 388942 17778 389026 18014
rect 389262 17778 389294 18014
rect 388674 2176 389294 17778
rect 392394 691654 393014 701760
rect 392394 691418 392426 691654
rect 392662 691418 392746 691654
rect 392982 691418 393014 691654
rect 392394 691334 393014 691418
rect 392394 691098 392426 691334
rect 392662 691098 392746 691334
rect 392982 691098 393014 691334
rect 392394 654454 393014 691098
rect 392394 654218 392426 654454
rect 392662 654218 392746 654454
rect 392982 654218 393014 654454
rect 392394 654134 393014 654218
rect 392394 653898 392426 654134
rect 392662 653898 392746 654134
rect 392982 653898 393014 654134
rect 392394 617254 393014 653898
rect 392394 617018 392426 617254
rect 392662 617018 392746 617254
rect 392982 617018 393014 617254
rect 392394 616934 393014 617018
rect 392394 616698 392426 616934
rect 392662 616698 392746 616934
rect 392982 616698 393014 616934
rect 392394 580054 393014 616698
rect 392394 579818 392426 580054
rect 392662 579818 392746 580054
rect 392982 579818 393014 580054
rect 392394 579734 393014 579818
rect 392394 579498 392426 579734
rect 392662 579498 392746 579734
rect 392982 579498 393014 579734
rect 392394 542854 393014 579498
rect 392394 542618 392426 542854
rect 392662 542618 392746 542854
rect 392982 542618 393014 542854
rect 392394 542534 393014 542618
rect 392394 542298 392426 542534
rect 392662 542298 392746 542534
rect 392982 542298 393014 542534
rect 392394 505654 393014 542298
rect 392394 505418 392426 505654
rect 392662 505418 392746 505654
rect 392982 505418 393014 505654
rect 392394 505334 393014 505418
rect 392394 505098 392426 505334
rect 392662 505098 392746 505334
rect 392982 505098 393014 505334
rect 392394 468454 393014 505098
rect 392394 468218 392426 468454
rect 392662 468218 392746 468454
rect 392982 468218 393014 468454
rect 392394 468134 393014 468218
rect 392394 467898 392426 468134
rect 392662 467898 392746 468134
rect 392982 467898 393014 468134
rect 392394 431254 393014 467898
rect 392394 431018 392426 431254
rect 392662 431018 392746 431254
rect 392982 431018 393014 431254
rect 392394 430934 393014 431018
rect 392394 430698 392426 430934
rect 392662 430698 392746 430934
rect 392982 430698 393014 430934
rect 392394 394054 393014 430698
rect 392394 393818 392426 394054
rect 392662 393818 392746 394054
rect 392982 393818 393014 394054
rect 392394 393734 393014 393818
rect 392394 393498 392426 393734
rect 392662 393498 392746 393734
rect 392982 393498 393014 393734
rect 392394 356854 393014 393498
rect 392394 356618 392426 356854
rect 392662 356618 392746 356854
rect 392982 356618 393014 356854
rect 392394 356534 393014 356618
rect 392394 356298 392426 356534
rect 392662 356298 392746 356534
rect 392982 356298 393014 356534
rect 392394 319654 393014 356298
rect 392394 319418 392426 319654
rect 392662 319418 392746 319654
rect 392982 319418 393014 319654
rect 392394 319334 393014 319418
rect 392394 319098 392426 319334
rect 392662 319098 392746 319334
rect 392982 319098 393014 319334
rect 392394 282454 393014 319098
rect 392394 282218 392426 282454
rect 392662 282218 392746 282454
rect 392982 282218 393014 282454
rect 392394 282134 393014 282218
rect 392394 281898 392426 282134
rect 392662 281898 392746 282134
rect 392982 281898 393014 282134
rect 392394 245254 393014 281898
rect 392394 245018 392426 245254
rect 392662 245018 392746 245254
rect 392982 245018 393014 245254
rect 392394 244934 393014 245018
rect 392394 244698 392426 244934
rect 392662 244698 392746 244934
rect 392982 244698 393014 244934
rect 392394 208054 393014 244698
rect 392394 207818 392426 208054
rect 392662 207818 392746 208054
rect 392982 207818 393014 208054
rect 392394 207734 393014 207818
rect 392394 207498 392426 207734
rect 392662 207498 392746 207734
rect 392982 207498 393014 207734
rect 392394 170854 393014 207498
rect 392394 170618 392426 170854
rect 392662 170618 392746 170854
rect 392982 170618 393014 170854
rect 392394 170534 393014 170618
rect 392394 170298 392426 170534
rect 392662 170298 392746 170534
rect 392982 170298 393014 170534
rect 392394 133654 393014 170298
rect 392394 133418 392426 133654
rect 392662 133418 392746 133654
rect 392982 133418 393014 133654
rect 392394 133334 393014 133418
rect 392394 133098 392426 133334
rect 392662 133098 392746 133334
rect 392982 133098 393014 133334
rect 392394 96454 393014 133098
rect 392394 96218 392426 96454
rect 392662 96218 392746 96454
rect 392982 96218 393014 96454
rect 392394 96134 393014 96218
rect 392394 95898 392426 96134
rect 392662 95898 392746 96134
rect 392982 95898 393014 96134
rect 392394 59254 393014 95898
rect 392394 59018 392426 59254
rect 392662 59018 392746 59254
rect 392982 59018 393014 59254
rect 392394 58934 393014 59018
rect 392394 58698 392426 58934
rect 392662 58698 392746 58934
rect 392982 58698 393014 58934
rect 392394 22054 393014 58698
rect 392394 21818 392426 22054
rect 392662 21818 392746 22054
rect 392982 21818 393014 22054
rect 392394 21734 393014 21818
rect 392394 21498 392426 21734
rect 392662 21498 392746 21734
rect 392982 21498 393014 21734
rect 392394 2176 393014 21498
rect 396114 695374 396734 701760
rect 396114 695138 396146 695374
rect 396382 695138 396466 695374
rect 396702 695138 396734 695374
rect 396114 695054 396734 695138
rect 396114 694818 396146 695054
rect 396382 694818 396466 695054
rect 396702 694818 396734 695054
rect 396114 658174 396734 694818
rect 396114 657938 396146 658174
rect 396382 657938 396466 658174
rect 396702 657938 396734 658174
rect 396114 657854 396734 657938
rect 396114 657618 396146 657854
rect 396382 657618 396466 657854
rect 396702 657618 396734 657854
rect 396114 620974 396734 657618
rect 396114 620738 396146 620974
rect 396382 620738 396466 620974
rect 396702 620738 396734 620974
rect 396114 620654 396734 620738
rect 396114 620418 396146 620654
rect 396382 620418 396466 620654
rect 396702 620418 396734 620654
rect 396114 583774 396734 620418
rect 396114 583538 396146 583774
rect 396382 583538 396466 583774
rect 396702 583538 396734 583774
rect 396114 583454 396734 583538
rect 396114 583218 396146 583454
rect 396382 583218 396466 583454
rect 396702 583218 396734 583454
rect 396114 546574 396734 583218
rect 396114 546338 396146 546574
rect 396382 546338 396466 546574
rect 396702 546338 396734 546574
rect 396114 546254 396734 546338
rect 396114 546018 396146 546254
rect 396382 546018 396466 546254
rect 396702 546018 396734 546254
rect 396114 509374 396734 546018
rect 396114 509138 396146 509374
rect 396382 509138 396466 509374
rect 396702 509138 396734 509374
rect 396114 509054 396734 509138
rect 396114 508818 396146 509054
rect 396382 508818 396466 509054
rect 396702 508818 396734 509054
rect 396114 472174 396734 508818
rect 396114 471938 396146 472174
rect 396382 471938 396466 472174
rect 396702 471938 396734 472174
rect 396114 471854 396734 471938
rect 396114 471618 396146 471854
rect 396382 471618 396466 471854
rect 396702 471618 396734 471854
rect 396114 434974 396734 471618
rect 396114 434738 396146 434974
rect 396382 434738 396466 434974
rect 396702 434738 396734 434974
rect 396114 434654 396734 434738
rect 396114 434418 396146 434654
rect 396382 434418 396466 434654
rect 396702 434418 396734 434654
rect 396114 397774 396734 434418
rect 396114 397538 396146 397774
rect 396382 397538 396466 397774
rect 396702 397538 396734 397774
rect 396114 397454 396734 397538
rect 396114 397218 396146 397454
rect 396382 397218 396466 397454
rect 396702 397218 396734 397454
rect 396114 360574 396734 397218
rect 396114 360338 396146 360574
rect 396382 360338 396466 360574
rect 396702 360338 396734 360574
rect 396114 360254 396734 360338
rect 396114 360018 396146 360254
rect 396382 360018 396466 360254
rect 396702 360018 396734 360254
rect 396114 323374 396734 360018
rect 396114 323138 396146 323374
rect 396382 323138 396466 323374
rect 396702 323138 396734 323374
rect 396114 323054 396734 323138
rect 396114 322818 396146 323054
rect 396382 322818 396466 323054
rect 396702 322818 396734 323054
rect 396114 286174 396734 322818
rect 396114 285938 396146 286174
rect 396382 285938 396466 286174
rect 396702 285938 396734 286174
rect 396114 285854 396734 285938
rect 396114 285618 396146 285854
rect 396382 285618 396466 285854
rect 396702 285618 396734 285854
rect 396114 248974 396734 285618
rect 396114 248738 396146 248974
rect 396382 248738 396466 248974
rect 396702 248738 396734 248974
rect 396114 248654 396734 248738
rect 396114 248418 396146 248654
rect 396382 248418 396466 248654
rect 396702 248418 396734 248654
rect 396114 211774 396734 248418
rect 396114 211538 396146 211774
rect 396382 211538 396466 211774
rect 396702 211538 396734 211774
rect 396114 211454 396734 211538
rect 396114 211218 396146 211454
rect 396382 211218 396466 211454
rect 396702 211218 396734 211454
rect 396114 174574 396734 211218
rect 396114 174338 396146 174574
rect 396382 174338 396466 174574
rect 396702 174338 396734 174574
rect 396114 174254 396734 174338
rect 396114 174018 396146 174254
rect 396382 174018 396466 174254
rect 396702 174018 396734 174254
rect 396114 137374 396734 174018
rect 396114 137138 396146 137374
rect 396382 137138 396466 137374
rect 396702 137138 396734 137374
rect 396114 137054 396734 137138
rect 396114 136818 396146 137054
rect 396382 136818 396466 137054
rect 396702 136818 396734 137054
rect 396114 100174 396734 136818
rect 396114 99938 396146 100174
rect 396382 99938 396466 100174
rect 396702 99938 396734 100174
rect 396114 99854 396734 99938
rect 396114 99618 396146 99854
rect 396382 99618 396466 99854
rect 396702 99618 396734 99854
rect 396114 62974 396734 99618
rect 396114 62738 396146 62974
rect 396382 62738 396466 62974
rect 396702 62738 396734 62974
rect 396114 62654 396734 62738
rect 396114 62418 396146 62654
rect 396382 62418 396466 62654
rect 396702 62418 396734 62654
rect 396114 25774 396734 62418
rect 396114 25538 396146 25774
rect 396382 25538 396466 25774
rect 396702 25538 396734 25774
rect 396114 25454 396734 25538
rect 396114 25218 396146 25454
rect 396382 25218 396466 25454
rect 396702 25218 396734 25454
rect 396114 2176 396734 25218
rect 399834 699094 400454 701760
rect 399834 698858 399866 699094
rect 400102 698858 400186 699094
rect 400422 698858 400454 699094
rect 399834 698774 400454 698858
rect 399834 698538 399866 698774
rect 400102 698538 400186 698774
rect 400422 698538 400454 698774
rect 399834 661894 400454 698538
rect 399834 661658 399866 661894
rect 400102 661658 400186 661894
rect 400422 661658 400454 661894
rect 399834 661574 400454 661658
rect 399834 661338 399866 661574
rect 400102 661338 400186 661574
rect 400422 661338 400454 661574
rect 399834 624694 400454 661338
rect 399834 624458 399866 624694
rect 400102 624458 400186 624694
rect 400422 624458 400454 624694
rect 399834 624374 400454 624458
rect 399834 624138 399866 624374
rect 400102 624138 400186 624374
rect 400422 624138 400454 624374
rect 399834 587494 400454 624138
rect 399834 587258 399866 587494
rect 400102 587258 400186 587494
rect 400422 587258 400454 587494
rect 399834 587174 400454 587258
rect 399834 586938 399866 587174
rect 400102 586938 400186 587174
rect 400422 586938 400454 587174
rect 399834 550294 400454 586938
rect 399834 550058 399866 550294
rect 400102 550058 400186 550294
rect 400422 550058 400454 550294
rect 399834 549974 400454 550058
rect 399834 549738 399866 549974
rect 400102 549738 400186 549974
rect 400422 549738 400454 549974
rect 399834 513094 400454 549738
rect 399834 512858 399866 513094
rect 400102 512858 400186 513094
rect 400422 512858 400454 513094
rect 399834 512774 400454 512858
rect 399834 512538 399866 512774
rect 400102 512538 400186 512774
rect 400422 512538 400454 512774
rect 399834 475894 400454 512538
rect 399834 475658 399866 475894
rect 400102 475658 400186 475894
rect 400422 475658 400454 475894
rect 399834 475574 400454 475658
rect 399834 475338 399866 475574
rect 400102 475338 400186 475574
rect 400422 475338 400454 475574
rect 399834 438694 400454 475338
rect 399834 438458 399866 438694
rect 400102 438458 400186 438694
rect 400422 438458 400454 438694
rect 399834 438374 400454 438458
rect 399834 438138 399866 438374
rect 400102 438138 400186 438374
rect 400422 438138 400454 438374
rect 399834 401494 400454 438138
rect 399834 401258 399866 401494
rect 400102 401258 400186 401494
rect 400422 401258 400454 401494
rect 399834 401174 400454 401258
rect 399834 400938 399866 401174
rect 400102 400938 400186 401174
rect 400422 400938 400454 401174
rect 399834 364294 400454 400938
rect 399834 364058 399866 364294
rect 400102 364058 400186 364294
rect 400422 364058 400454 364294
rect 399834 363974 400454 364058
rect 399834 363738 399866 363974
rect 400102 363738 400186 363974
rect 400422 363738 400454 363974
rect 399834 327094 400454 363738
rect 399834 326858 399866 327094
rect 400102 326858 400186 327094
rect 400422 326858 400454 327094
rect 399834 326774 400454 326858
rect 399834 326538 399866 326774
rect 400102 326538 400186 326774
rect 400422 326538 400454 326774
rect 399834 289894 400454 326538
rect 399834 289658 399866 289894
rect 400102 289658 400186 289894
rect 400422 289658 400454 289894
rect 399834 289574 400454 289658
rect 399834 289338 399866 289574
rect 400102 289338 400186 289574
rect 400422 289338 400454 289574
rect 399834 252694 400454 289338
rect 399834 252458 399866 252694
rect 400102 252458 400186 252694
rect 400422 252458 400454 252694
rect 399834 252374 400454 252458
rect 399834 252138 399866 252374
rect 400102 252138 400186 252374
rect 400422 252138 400454 252374
rect 399834 215494 400454 252138
rect 399834 215258 399866 215494
rect 400102 215258 400186 215494
rect 400422 215258 400454 215494
rect 399834 215174 400454 215258
rect 399834 214938 399866 215174
rect 400102 214938 400186 215174
rect 400422 214938 400454 215174
rect 399834 178294 400454 214938
rect 399834 178058 399866 178294
rect 400102 178058 400186 178294
rect 400422 178058 400454 178294
rect 399834 177974 400454 178058
rect 399834 177738 399866 177974
rect 400102 177738 400186 177974
rect 400422 177738 400454 177974
rect 399834 141094 400454 177738
rect 399834 140858 399866 141094
rect 400102 140858 400186 141094
rect 400422 140858 400454 141094
rect 399834 140774 400454 140858
rect 399834 140538 399866 140774
rect 400102 140538 400186 140774
rect 400422 140538 400454 140774
rect 399834 103894 400454 140538
rect 399834 103658 399866 103894
rect 400102 103658 400186 103894
rect 400422 103658 400454 103894
rect 399834 103574 400454 103658
rect 399834 103338 399866 103574
rect 400102 103338 400186 103574
rect 400422 103338 400454 103574
rect 399834 66694 400454 103338
rect 399834 66458 399866 66694
rect 400102 66458 400186 66694
rect 400422 66458 400454 66694
rect 399834 66374 400454 66458
rect 399834 66138 399866 66374
rect 400102 66138 400186 66374
rect 400422 66138 400454 66374
rect 399834 29494 400454 66138
rect 399834 29258 399866 29494
rect 400102 29258 400186 29494
rect 400422 29258 400454 29494
rect 399834 29174 400454 29258
rect 399834 28938 399866 29174
rect 400102 28938 400186 29174
rect 400422 28938 400454 29174
rect 399834 2176 400454 28938
rect 410994 673054 411614 701760
rect 410994 672818 411026 673054
rect 411262 672818 411346 673054
rect 411582 672818 411614 673054
rect 410994 672734 411614 672818
rect 410994 672498 411026 672734
rect 411262 672498 411346 672734
rect 411582 672498 411614 672734
rect 410994 635854 411614 672498
rect 410994 635618 411026 635854
rect 411262 635618 411346 635854
rect 411582 635618 411614 635854
rect 410994 635534 411614 635618
rect 410994 635298 411026 635534
rect 411262 635298 411346 635534
rect 411582 635298 411614 635534
rect 410994 598654 411614 635298
rect 410994 598418 411026 598654
rect 411262 598418 411346 598654
rect 411582 598418 411614 598654
rect 410994 598334 411614 598418
rect 410994 598098 411026 598334
rect 411262 598098 411346 598334
rect 411582 598098 411614 598334
rect 410994 561454 411614 598098
rect 410994 561218 411026 561454
rect 411262 561218 411346 561454
rect 411582 561218 411614 561454
rect 410994 561134 411614 561218
rect 410994 560898 411026 561134
rect 411262 560898 411346 561134
rect 411582 560898 411614 561134
rect 410994 524254 411614 560898
rect 410994 524018 411026 524254
rect 411262 524018 411346 524254
rect 411582 524018 411614 524254
rect 410994 523934 411614 524018
rect 410994 523698 411026 523934
rect 411262 523698 411346 523934
rect 411582 523698 411614 523934
rect 410994 487054 411614 523698
rect 410994 486818 411026 487054
rect 411262 486818 411346 487054
rect 411582 486818 411614 487054
rect 410994 486734 411614 486818
rect 410994 486498 411026 486734
rect 411262 486498 411346 486734
rect 411582 486498 411614 486734
rect 410994 449854 411614 486498
rect 410994 449618 411026 449854
rect 411262 449618 411346 449854
rect 411582 449618 411614 449854
rect 410994 449534 411614 449618
rect 410994 449298 411026 449534
rect 411262 449298 411346 449534
rect 411582 449298 411614 449534
rect 410994 412654 411614 449298
rect 410994 412418 411026 412654
rect 411262 412418 411346 412654
rect 411582 412418 411614 412654
rect 410994 412334 411614 412418
rect 410994 412098 411026 412334
rect 411262 412098 411346 412334
rect 411582 412098 411614 412334
rect 410994 375454 411614 412098
rect 410994 375218 411026 375454
rect 411262 375218 411346 375454
rect 411582 375218 411614 375454
rect 410994 375134 411614 375218
rect 410994 374898 411026 375134
rect 411262 374898 411346 375134
rect 411582 374898 411614 375134
rect 410994 338254 411614 374898
rect 410994 338018 411026 338254
rect 411262 338018 411346 338254
rect 411582 338018 411614 338254
rect 410994 337934 411614 338018
rect 410994 337698 411026 337934
rect 411262 337698 411346 337934
rect 411582 337698 411614 337934
rect 410994 301054 411614 337698
rect 410994 300818 411026 301054
rect 411262 300818 411346 301054
rect 411582 300818 411614 301054
rect 410994 300734 411614 300818
rect 410994 300498 411026 300734
rect 411262 300498 411346 300734
rect 411582 300498 411614 300734
rect 410994 263854 411614 300498
rect 410994 263618 411026 263854
rect 411262 263618 411346 263854
rect 411582 263618 411614 263854
rect 410994 263534 411614 263618
rect 410994 263298 411026 263534
rect 411262 263298 411346 263534
rect 411582 263298 411614 263534
rect 410994 226654 411614 263298
rect 410994 226418 411026 226654
rect 411262 226418 411346 226654
rect 411582 226418 411614 226654
rect 410994 226334 411614 226418
rect 410994 226098 411026 226334
rect 411262 226098 411346 226334
rect 411582 226098 411614 226334
rect 410994 189454 411614 226098
rect 410994 189218 411026 189454
rect 411262 189218 411346 189454
rect 411582 189218 411614 189454
rect 410994 189134 411614 189218
rect 410994 188898 411026 189134
rect 411262 188898 411346 189134
rect 411582 188898 411614 189134
rect 410994 152254 411614 188898
rect 410994 152018 411026 152254
rect 411262 152018 411346 152254
rect 411582 152018 411614 152254
rect 410994 151934 411614 152018
rect 410994 151698 411026 151934
rect 411262 151698 411346 151934
rect 411582 151698 411614 151934
rect 410994 115054 411614 151698
rect 410994 114818 411026 115054
rect 411262 114818 411346 115054
rect 411582 114818 411614 115054
rect 410994 114734 411614 114818
rect 410994 114498 411026 114734
rect 411262 114498 411346 114734
rect 411582 114498 411614 114734
rect 410994 77854 411614 114498
rect 410994 77618 411026 77854
rect 411262 77618 411346 77854
rect 411582 77618 411614 77854
rect 410994 77534 411614 77618
rect 410994 77298 411026 77534
rect 411262 77298 411346 77534
rect 411582 77298 411614 77534
rect 410994 40654 411614 77298
rect 410994 40418 411026 40654
rect 411262 40418 411346 40654
rect 411582 40418 411614 40654
rect 410994 40334 411614 40418
rect 410994 40098 411026 40334
rect 411262 40098 411346 40334
rect 411582 40098 411614 40334
rect 410994 3454 411614 40098
rect 410994 3218 411026 3454
rect 411262 3218 411346 3454
rect 411582 3218 411614 3454
rect 410994 3134 411614 3218
rect 410994 2898 411026 3134
rect 411262 2898 411346 3134
rect 411582 2898 411614 3134
rect 410994 2176 411614 2898
rect 414714 676774 415334 701760
rect 414714 676538 414746 676774
rect 414982 676538 415066 676774
rect 415302 676538 415334 676774
rect 414714 676454 415334 676538
rect 414714 676218 414746 676454
rect 414982 676218 415066 676454
rect 415302 676218 415334 676454
rect 414714 639574 415334 676218
rect 414714 639338 414746 639574
rect 414982 639338 415066 639574
rect 415302 639338 415334 639574
rect 414714 639254 415334 639338
rect 414714 639018 414746 639254
rect 414982 639018 415066 639254
rect 415302 639018 415334 639254
rect 414714 602374 415334 639018
rect 414714 602138 414746 602374
rect 414982 602138 415066 602374
rect 415302 602138 415334 602374
rect 414714 602054 415334 602138
rect 414714 601818 414746 602054
rect 414982 601818 415066 602054
rect 415302 601818 415334 602054
rect 414714 565174 415334 601818
rect 414714 564938 414746 565174
rect 414982 564938 415066 565174
rect 415302 564938 415334 565174
rect 414714 564854 415334 564938
rect 414714 564618 414746 564854
rect 414982 564618 415066 564854
rect 415302 564618 415334 564854
rect 414714 527974 415334 564618
rect 414714 527738 414746 527974
rect 414982 527738 415066 527974
rect 415302 527738 415334 527974
rect 414714 527654 415334 527738
rect 414714 527418 414746 527654
rect 414982 527418 415066 527654
rect 415302 527418 415334 527654
rect 414714 490774 415334 527418
rect 414714 490538 414746 490774
rect 414982 490538 415066 490774
rect 415302 490538 415334 490774
rect 414714 490454 415334 490538
rect 414714 490218 414746 490454
rect 414982 490218 415066 490454
rect 415302 490218 415334 490454
rect 414714 453574 415334 490218
rect 414714 453338 414746 453574
rect 414982 453338 415066 453574
rect 415302 453338 415334 453574
rect 414714 453254 415334 453338
rect 414714 453018 414746 453254
rect 414982 453018 415066 453254
rect 415302 453018 415334 453254
rect 414714 416374 415334 453018
rect 414714 416138 414746 416374
rect 414982 416138 415066 416374
rect 415302 416138 415334 416374
rect 414714 416054 415334 416138
rect 414714 415818 414746 416054
rect 414982 415818 415066 416054
rect 415302 415818 415334 416054
rect 414714 379174 415334 415818
rect 414714 378938 414746 379174
rect 414982 378938 415066 379174
rect 415302 378938 415334 379174
rect 414714 378854 415334 378938
rect 414714 378618 414746 378854
rect 414982 378618 415066 378854
rect 415302 378618 415334 378854
rect 414714 341974 415334 378618
rect 414714 341738 414746 341974
rect 414982 341738 415066 341974
rect 415302 341738 415334 341974
rect 414714 341654 415334 341738
rect 414714 341418 414746 341654
rect 414982 341418 415066 341654
rect 415302 341418 415334 341654
rect 414714 304774 415334 341418
rect 414714 304538 414746 304774
rect 414982 304538 415066 304774
rect 415302 304538 415334 304774
rect 414714 304454 415334 304538
rect 414714 304218 414746 304454
rect 414982 304218 415066 304454
rect 415302 304218 415334 304454
rect 414714 267574 415334 304218
rect 414714 267338 414746 267574
rect 414982 267338 415066 267574
rect 415302 267338 415334 267574
rect 414714 267254 415334 267338
rect 414714 267018 414746 267254
rect 414982 267018 415066 267254
rect 415302 267018 415334 267254
rect 414714 230374 415334 267018
rect 414714 230138 414746 230374
rect 414982 230138 415066 230374
rect 415302 230138 415334 230374
rect 414714 230054 415334 230138
rect 414714 229818 414746 230054
rect 414982 229818 415066 230054
rect 415302 229818 415334 230054
rect 414714 193174 415334 229818
rect 414714 192938 414746 193174
rect 414982 192938 415066 193174
rect 415302 192938 415334 193174
rect 414714 192854 415334 192938
rect 414714 192618 414746 192854
rect 414982 192618 415066 192854
rect 415302 192618 415334 192854
rect 414714 155974 415334 192618
rect 414714 155738 414746 155974
rect 414982 155738 415066 155974
rect 415302 155738 415334 155974
rect 414714 155654 415334 155738
rect 414714 155418 414746 155654
rect 414982 155418 415066 155654
rect 415302 155418 415334 155654
rect 414714 118774 415334 155418
rect 414714 118538 414746 118774
rect 414982 118538 415066 118774
rect 415302 118538 415334 118774
rect 414714 118454 415334 118538
rect 414714 118218 414746 118454
rect 414982 118218 415066 118454
rect 415302 118218 415334 118454
rect 414714 81574 415334 118218
rect 414714 81338 414746 81574
rect 414982 81338 415066 81574
rect 415302 81338 415334 81574
rect 414714 81254 415334 81338
rect 414714 81018 414746 81254
rect 414982 81018 415066 81254
rect 415302 81018 415334 81254
rect 414714 44374 415334 81018
rect 414714 44138 414746 44374
rect 414982 44138 415066 44374
rect 415302 44138 415334 44374
rect 414714 44054 415334 44138
rect 414714 43818 414746 44054
rect 414982 43818 415066 44054
rect 415302 43818 415334 44054
rect 414714 7174 415334 43818
rect 414714 6938 414746 7174
rect 414982 6938 415066 7174
rect 415302 6938 415334 7174
rect 414714 6854 415334 6938
rect 414714 6618 414746 6854
rect 414982 6618 415066 6854
rect 415302 6618 415334 6854
rect 414714 2176 415334 6618
rect 418434 680494 419054 701760
rect 418434 680258 418466 680494
rect 418702 680258 418786 680494
rect 419022 680258 419054 680494
rect 418434 680174 419054 680258
rect 418434 679938 418466 680174
rect 418702 679938 418786 680174
rect 419022 679938 419054 680174
rect 418434 643294 419054 679938
rect 418434 643058 418466 643294
rect 418702 643058 418786 643294
rect 419022 643058 419054 643294
rect 418434 642974 419054 643058
rect 418434 642738 418466 642974
rect 418702 642738 418786 642974
rect 419022 642738 419054 642974
rect 418434 606094 419054 642738
rect 418434 605858 418466 606094
rect 418702 605858 418786 606094
rect 419022 605858 419054 606094
rect 418434 605774 419054 605858
rect 418434 605538 418466 605774
rect 418702 605538 418786 605774
rect 419022 605538 419054 605774
rect 418434 568894 419054 605538
rect 418434 568658 418466 568894
rect 418702 568658 418786 568894
rect 419022 568658 419054 568894
rect 418434 568574 419054 568658
rect 418434 568338 418466 568574
rect 418702 568338 418786 568574
rect 419022 568338 419054 568574
rect 418434 531694 419054 568338
rect 418434 531458 418466 531694
rect 418702 531458 418786 531694
rect 419022 531458 419054 531694
rect 418434 531374 419054 531458
rect 418434 531138 418466 531374
rect 418702 531138 418786 531374
rect 419022 531138 419054 531374
rect 418434 494494 419054 531138
rect 418434 494258 418466 494494
rect 418702 494258 418786 494494
rect 419022 494258 419054 494494
rect 418434 494174 419054 494258
rect 418434 493938 418466 494174
rect 418702 493938 418786 494174
rect 419022 493938 419054 494174
rect 418434 457294 419054 493938
rect 418434 457058 418466 457294
rect 418702 457058 418786 457294
rect 419022 457058 419054 457294
rect 418434 456974 419054 457058
rect 418434 456738 418466 456974
rect 418702 456738 418786 456974
rect 419022 456738 419054 456974
rect 418434 420094 419054 456738
rect 418434 419858 418466 420094
rect 418702 419858 418786 420094
rect 419022 419858 419054 420094
rect 418434 419774 419054 419858
rect 418434 419538 418466 419774
rect 418702 419538 418786 419774
rect 419022 419538 419054 419774
rect 418434 382894 419054 419538
rect 418434 382658 418466 382894
rect 418702 382658 418786 382894
rect 419022 382658 419054 382894
rect 418434 382574 419054 382658
rect 418434 382338 418466 382574
rect 418702 382338 418786 382574
rect 419022 382338 419054 382574
rect 418434 345694 419054 382338
rect 418434 345458 418466 345694
rect 418702 345458 418786 345694
rect 419022 345458 419054 345694
rect 418434 345374 419054 345458
rect 418434 345138 418466 345374
rect 418702 345138 418786 345374
rect 419022 345138 419054 345374
rect 418434 308494 419054 345138
rect 418434 308258 418466 308494
rect 418702 308258 418786 308494
rect 419022 308258 419054 308494
rect 418434 308174 419054 308258
rect 418434 307938 418466 308174
rect 418702 307938 418786 308174
rect 419022 307938 419054 308174
rect 418434 271294 419054 307938
rect 418434 271058 418466 271294
rect 418702 271058 418786 271294
rect 419022 271058 419054 271294
rect 418434 270974 419054 271058
rect 418434 270738 418466 270974
rect 418702 270738 418786 270974
rect 419022 270738 419054 270974
rect 418434 234094 419054 270738
rect 418434 233858 418466 234094
rect 418702 233858 418786 234094
rect 419022 233858 419054 234094
rect 418434 233774 419054 233858
rect 418434 233538 418466 233774
rect 418702 233538 418786 233774
rect 419022 233538 419054 233774
rect 418434 196894 419054 233538
rect 418434 196658 418466 196894
rect 418702 196658 418786 196894
rect 419022 196658 419054 196894
rect 418434 196574 419054 196658
rect 418434 196338 418466 196574
rect 418702 196338 418786 196574
rect 419022 196338 419054 196574
rect 418434 159694 419054 196338
rect 418434 159458 418466 159694
rect 418702 159458 418786 159694
rect 419022 159458 419054 159694
rect 418434 159374 419054 159458
rect 418434 159138 418466 159374
rect 418702 159138 418786 159374
rect 419022 159138 419054 159374
rect 418434 122494 419054 159138
rect 418434 122258 418466 122494
rect 418702 122258 418786 122494
rect 419022 122258 419054 122494
rect 418434 122174 419054 122258
rect 418434 121938 418466 122174
rect 418702 121938 418786 122174
rect 419022 121938 419054 122174
rect 418434 85294 419054 121938
rect 418434 85058 418466 85294
rect 418702 85058 418786 85294
rect 419022 85058 419054 85294
rect 418434 84974 419054 85058
rect 418434 84738 418466 84974
rect 418702 84738 418786 84974
rect 419022 84738 419054 84974
rect 418434 48094 419054 84738
rect 418434 47858 418466 48094
rect 418702 47858 418786 48094
rect 419022 47858 419054 48094
rect 418434 47774 419054 47858
rect 418434 47538 418466 47774
rect 418702 47538 418786 47774
rect 419022 47538 419054 47774
rect 418434 10894 419054 47538
rect 418434 10658 418466 10894
rect 418702 10658 418786 10894
rect 419022 10658 419054 10894
rect 418434 10574 419054 10658
rect 418434 10338 418466 10574
rect 418702 10338 418786 10574
rect 419022 10338 419054 10574
rect 418434 2176 419054 10338
rect 422154 684214 422774 701760
rect 422154 683978 422186 684214
rect 422422 683978 422506 684214
rect 422742 683978 422774 684214
rect 422154 683894 422774 683978
rect 422154 683658 422186 683894
rect 422422 683658 422506 683894
rect 422742 683658 422774 683894
rect 422154 647014 422774 683658
rect 422154 646778 422186 647014
rect 422422 646778 422506 647014
rect 422742 646778 422774 647014
rect 422154 646694 422774 646778
rect 422154 646458 422186 646694
rect 422422 646458 422506 646694
rect 422742 646458 422774 646694
rect 422154 609814 422774 646458
rect 422154 609578 422186 609814
rect 422422 609578 422506 609814
rect 422742 609578 422774 609814
rect 422154 609494 422774 609578
rect 422154 609258 422186 609494
rect 422422 609258 422506 609494
rect 422742 609258 422774 609494
rect 422154 572614 422774 609258
rect 422154 572378 422186 572614
rect 422422 572378 422506 572614
rect 422742 572378 422774 572614
rect 422154 572294 422774 572378
rect 422154 572058 422186 572294
rect 422422 572058 422506 572294
rect 422742 572058 422774 572294
rect 422154 535414 422774 572058
rect 422154 535178 422186 535414
rect 422422 535178 422506 535414
rect 422742 535178 422774 535414
rect 422154 535094 422774 535178
rect 422154 534858 422186 535094
rect 422422 534858 422506 535094
rect 422742 534858 422774 535094
rect 422154 498214 422774 534858
rect 422154 497978 422186 498214
rect 422422 497978 422506 498214
rect 422742 497978 422774 498214
rect 422154 497894 422774 497978
rect 422154 497658 422186 497894
rect 422422 497658 422506 497894
rect 422742 497658 422774 497894
rect 422154 461014 422774 497658
rect 422154 460778 422186 461014
rect 422422 460778 422506 461014
rect 422742 460778 422774 461014
rect 422154 460694 422774 460778
rect 422154 460458 422186 460694
rect 422422 460458 422506 460694
rect 422742 460458 422774 460694
rect 422154 423814 422774 460458
rect 422154 423578 422186 423814
rect 422422 423578 422506 423814
rect 422742 423578 422774 423814
rect 422154 423494 422774 423578
rect 422154 423258 422186 423494
rect 422422 423258 422506 423494
rect 422742 423258 422774 423494
rect 422154 386614 422774 423258
rect 422154 386378 422186 386614
rect 422422 386378 422506 386614
rect 422742 386378 422774 386614
rect 422154 386294 422774 386378
rect 422154 386058 422186 386294
rect 422422 386058 422506 386294
rect 422742 386058 422774 386294
rect 422154 349414 422774 386058
rect 422154 349178 422186 349414
rect 422422 349178 422506 349414
rect 422742 349178 422774 349414
rect 422154 349094 422774 349178
rect 422154 348858 422186 349094
rect 422422 348858 422506 349094
rect 422742 348858 422774 349094
rect 422154 312214 422774 348858
rect 422154 311978 422186 312214
rect 422422 311978 422506 312214
rect 422742 311978 422774 312214
rect 422154 311894 422774 311978
rect 422154 311658 422186 311894
rect 422422 311658 422506 311894
rect 422742 311658 422774 311894
rect 422154 275014 422774 311658
rect 422154 274778 422186 275014
rect 422422 274778 422506 275014
rect 422742 274778 422774 275014
rect 422154 274694 422774 274778
rect 422154 274458 422186 274694
rect 422422 274458 422506 274694
rect 422742 274458 422774 274694
rect 422154 237814 422774 274458
rect 422154 237578 422186 237814
rect 422422 237578 422506 237814
rect 422742 237578 422774 237814
rect 422154 237494 422774 237578
rect 422154 237258 422186 237494
rect 422422 237258 422506 237494
rect 422742 237258 422774 237494
rect 422154 200614 422774 237258
rect 422154 200378 422186 200614
rect 422422 200378 422506 200614
rect 422742 200378 422774 200614
rect 422154 200294 422774 200378
rect 422154 200058 422186 200294
rect 422422 200058 422506 200294
rect 422742 200058 422774 200294
rect 422154 163414 422774 200058
rect 422154 163178 422186 163414
rect 422422 163178 422506 163414
rect 422742 163178 422774 163414
rect 422154 163094 422774 163178
rect 422154 162858 422186 163094
rect 422422 162858 422506 163094
rect 422742 162858 422774 163094
rect 422154 126214 422774 162858
rect 422154 125978 422186 126214
rect 422422 125978 422506 126214
rect 422742 125978 422774 126214
rect 422154 125894 422774 125978
rect 422154 125658 422186 125894
rect 422422 125658 422506 125894
rect 422742 125658 422774 125894
rect 422154 89014 422774 125658
rect 422154 88778 422186 89014
rect 422422 88778 422506 89014
rect 422742 88778 422774 89014
rect 422154 88694 422774 88778
rect 422154 88458 422186 88694
rect 422422 88458 422506 88694
rect 422742 88458 422774 88694
rect 422154 51814 422774 88458
rect 422154 51578 422186 51814
rect 422422 51578 422506 51814
rect 422742 51578 422774 51814
rect 422154 51494 422774 51578
rect 422154 51258 422186 51494
rect 422422 51258 422506 51494
rect 422742 51258 422774 51494
rect 422154 14614 422774 51258
rect 422154 14378 422186 14614
rect 422422 14378 422506 14614
rect 422742 14378 422774 14614
rect 422154 14294 422774 14378
rect 422154 14058 422186 14294
rect 422422 14058 422506 14294
rect 422742 14058 422774 14294
rect 422154 2176 422774 14058
rect 425874 687934 426494 701760
rect 425874 687698 425906 687934
rect 426142 687698 426226 687934
rect 426462 687698 426494 687934
rect 425874 687614 426494 687698
rect 425874 687378 425906 687614
rect 426142 687378 426226 687614
rect 426462 687378 426494 687614
rect 425874 650734 426494 687378
rect 425874 650498 425906 650734
rect 426142 650498 426226 650734
rect 426462 650498 426494 650734
rect 425874 650414 426494 650498
rect 425874 650178 425906 650414
rect 426142 650178 426226 650414
rect 426462 650178 426494 650414
rect 425874 613534 426494 650178
rect 425874 613298 425906 613534
rect 426142 613298 426226 613534
rect 426462 613298 426494 613534
rect 425874 613214 426494 613298
rect 425874 612978 425906 613214
rect 426142 612978 426226 613214
rect 426462 612978 426494 613214
rect 425874 576334 426494 612978
rect 425874 576098 425906 576334
rect 426142 576098 426226 576334
rect 426462 576098 426494 576334
rect 425874 576014 426494 576098
rect 425874 575778 425906 576014
rect 426142 575778 426226 576014
rect 426462 575778 426494 576014
rect 425874 539134 426494 575778
rect 425874 538898 425906 539134
rect 426142 538898 426226 539134
rect 426462 538898 426494 539134
rect 425874 538814 426494 538898
rect 425874 538578 425906 538814
rect 426142 538578 426226 538814
rect 426462 538578 426494 538814
rect 425874 501934 426494 538578
rect 425874 501698 425906 501934
rect 426142 501698 426226 501934
rect 426462 501698 426494 501934
rect 425874 501614 426494 501698
rect 425874 501378 425906 501614
rect 426142 501378 426226 501614
rect 426462 501378 426494 501614
rect 425874 464734 426494 501378
rect 425874 464498 425906 464734
rect 426142 464498 426226 464734
rect 426462 464498 426494 464734
rect 425874 464414 426494 464498
rect 425874 464178 425906 464414
rect 426142 464178 426226 464414
rect 426462 464178 426494 464414
rect 425874 427534 426494 464178
rect 425874 427298 425906 427534
rect 426142 427298 426226 427534
rect 426462 427298 426494 427534
rect 425874 427214 426494 427298
rect 425874 426978 425906 427214
rect 426142 426978 426226 427214
rect 426462 426978 426494 427214
rect 425874 390334 426494 426978
rect 425874 390098 425906 390334
rect 426142 390098 426226 390334
rect 426462 390098 426494 390334
rect 425874 390014 426494 390098
rect 425874 389778 425906 390014
rect 426142 389778 426226 390014
rect 426462 389778 426494 390014
rect 425874 353134 426494 389778
rect 425874 352898 425906 353134
rect 426142 352898 426226 353134
rect 426462 352898 426494 353134
rect 425874 352814 426494 352898
rect 425874 352578 425906 352814
rect 426142 352578 426226 352814
rect 426462 352578 426494 352814
rect 425874 315934 426494 352578
rect 425874 315698 425906 315934
rect 426142 315698 426226 315934
rect 426462 315698 426494 315934
rect 425874 315614 426494 315698
rect 425874 315378 425906 315614
rect 426142 315378 426226 315614
rect 426462 315378 426494 315614
rect 425874 278734 426494 315378
rect 425874 278498 425906 278734
rect 426142 278498 426226 278734
rect 426462 278498 426494 278734
rect 425874 278414 426494 278498
rect 425874 278178 425906 278414
rect 426142 278178 426226 278414
rect 426462 278178 426494 278414
rect 425874 241534 426494 278178
rect 425874 241298 425906 241534
rect 426142 241298 426226 241534
rect 426462 241298 426494 241534
rect 425874 241214 426494 241298
rect 425874 240978 425906 241214
rect 426142 240978 426226 241214
rect 426462 240978 426494 241214
rect 425874 204334 426494 240978
rect 425874 204098 425906 204334
rect 426142 204098 426226 204334
rect 426462 204098 426494 204334
rect 425874 204014 426494 204098
rect 425874 203778 425906 204014
rect 426142 203778 426226 204014
rect 426462 203778 426494 204014
rect 425874 167134 426494 203778
rect 425874 166898 425906 167134
rect 426142 166898 426226 167134
rect 426462 166898 426494 167134
rect 425874 166814 426494 166898
rect 425874 166578 425906 166814
rect 426142 166578 426226 166814
rect 426462 166578 426494 166814
rect 425874 129934 426494 166578
rect 425874 129698 425906 129934
rect 426142 129698 426226 129934
rect 426462 129698 426494 129934
rect 425874 129614 426494 129698
rect 425874 129378 425906 129614
rect 426142 129378 426226 129614
rect 426462 129378 426494 129614
rect 425874 92734 426494 129378
rect 425874 92498 425906 92734
rect 426142 92498 426226 92734
rect 426462 92498 426494 92734
rect 425874 92414 426494 92498
rect 425874 92178 425906 92414
rect 426142 92178 426226 92414
rect 426462 92178 426494 92414
rect 425874 55534 426494 92178
rect 425874 55298 425906 55534
rect 426142 55298 426226 55534
rect 426462 55298 426494 55534
rect 425874 55214 426494 55298
rect 425874 54978 425906 55214
rect 426142 54978 426226 55214
rect 426462 54978 426494 55214
rect 425874 18334 426494 54978
rect 425874 18098 425906 18334
rect 426142 18098 426226 18334
rect 426462 18098 426494 18334
rect 425874 18014 426494 18098
rect 425874 17778 425906 18014
rect 426142 17778 426226 18014
rect 426462 17778 426494 18014
rect 425874 2176 426494 17778
rect 429594 691654 430214 701760
rect 429594 691418 429626 691654
rect 429862 691418 429946 691654
rect 430182 691418 430214 691654
rect 429594 691334 430214 691418
rect 429594 691098 429626 691334
rect 429862 691098 429946 691334
rect 430182 691098 430214 691334
rect 429594 654454 430214 691098
rect 429594 654218 429626 654454
rect 429862 654218 429946 654454
rect 430182 654218 430214 654454
rect 429594 654134 430214 654218
rect 429594 653898 429626 654134
rect 429862 653898 429946 654134
rect 430182 653898 430214 654134
rect 429594 617254 430214 653898
rect 429594 617018 429626 617254
rect 429862 617018 429946 617254
rect 430182 617018 430214 617254
rect 429594 616934 430214 617018
rect 429594 616698 429626 616934
rect 429862 616698 429946 616934
rect 430182 616698 430214 616934
rect 429594 580054 430214 616698
rect 429594 579818 429626 580054
rect 429862 579818 429946 580054
rect 430182 579818 430214 580054
rect 429594 579734 430214 579818
rect 429594 579498 429626 579734
rect 429862 579498 429946 579734
rect 430182 579498 430214 579734
rect 429594 542854 430214 579498
rect 429594 542618 429626 542854
rect 429862 542618 429946 542854
rect 430182 542618 430214 542854
rect 429594 542534 430214 542618
rect 429594 542298 429626 542534
rect 429862 542298 429946 542534
rect 430182 542298 430214 542534
rect 429594 505654 430214 542298
rect 429594 505418 429626 505654
rect 429862 505418 429946 505654
rect 430182 505418 430214 505654
rect 429594 505334 430214 505418
rect 429594 505098 429626 505334
rect 429862 505098 429946 505334
rect 430182 505098 430214 505334
rect 429594 468454 430214 505098
rect 429594 468218 429626 468454
rect 429862 468218 429946 468454
rect 430182 468218 430214 468454
rect 429594 468134 430214 468218
rect 429594 467898 429626 468134
rect 429862 467898 429946 468134
rect 430182 467898 430214 468134
rect 429594 431254 430214 467898
rect 429594 431018 429626 431254
rect 429862 431018 429946 431254
rect 430182 431018 430214 431254
rect 429594 430934 430214 431018
rect 429594 430698 429626 430934
rect 429862 430698 429946 430934
rect 430182 430698 430214 430934
rect 429594 394054 430214 430698
rect 429594 393818 429626 394054
rect 429862 393818 429946 394054
rect 430182 393818 430214 394054
rect 429594 393734 430214 393818
rect 429594 393498 429626 393734
rect 429862 393498 429946 393734
rect 430182 393498 430214 393734
rect 429594 356854 430214 393498
rect 429594 356618 429626 356854
rect 429862 356618 429946 356854
rect 430182 356618 430214 356854
rect 429594 356534 430214 356618
rect 429594 356298 429626 356534
rect 429862 356298 429946 356534
rect 430182 356298 430214 356534
rect 429594 319654 430214 356298
rect 429594 319418 429626 319654
rect 429862 319418 429946 319654
rect 430182 319418 430214 319654
rect 429594 319334 430214 319418
rect 429594 319098 429626 319334
rect 429862 319098 429946 319334
rect 430182 319098 430214 319334
rect 429594 282454 430214 319098
rect 429594 282218 429626 282454
rect 429862 282218 429946 282454
rect 430182 282218 430214 282454
rect 429594 282134 430214 282218
rect 429594 281898 429626 282134
rect 429862 281898 429946 282134
rect 430182 281898 430214 282134
rect 429594 245254 430214 281898
rect 429594 245018 429626 245254
rect 429862 245018 429946 245254
rect 430182 245018 430214 245254
rect 429594 244934 430214 245018
rect 429594 244698 429626 244934
rect 429862 244698 429946 244934
rect 430182 244698 430214 244934
rect 429594 208054 430214 244698
rect 429594 207818 429626 208054
rect 429862 207818 429946 208054
rect 430182 207818 430214 208054
rect 429594 207734 430214 207818
rect 429594 207498 429626 207734
rect 429862 207498 429946 207734
rect 430182 207498 430214 207734
rect 429594 170854 430214 207498
rect 429594 170618 429626 170854
rect 429862 170618 429946 170854
rect 430182 170618 430214 170854
rect 429594 170534 430214 170618
rect 429594 170298 429626 170534
rect 429862 170298 429946 170534
rect 430182 170298 430214 170534
rect 429594 133654 430214 170298
rect 429594 133418 429626 133654
rect 429862 133418 429946 133654
rect 430182 133418 430214 133654
rect 429594 133334 430214 133418
rect 429594 133098 429626 133334
rect 429862 133098 429946 133334
rect 430182 133098 430214 133334
rect 429594 96454 430214 133098
rect 429594 96218 429626 96454
rect 429862 96218 429946 96454
rect 430182 96218 430214 96454
rect 429594 96134 430214 96218
rect 429594 95898 429626 96134
rect 429862 95898 429946 96134
rect 430182 95898 430214 96134
rect 429594 59254 430214 95898
rect 429594 59018 429626 59254
rect 429862 59018 429946 59254
rect 430182 59018 430214 59254
rect 429594 58934 430214 59018
rect 429594 58698 429626 58934
rect 429862 58698 429946 58934
rect 430182 58698 430214 58934
rect 429594 22054 430214 58698
rect 429594 21818 429626 22054
rect 429862 21818 429946 22054
rect 430182 21818 430214 22054
rect 429594 21734 430214 21818
rect 429594 21498 429626 21734
rect 429862 21498 429946 21734
rect 430182 21498 430214 21734
rect 429594 2176 430214 21498
rect 433314 695374 433934 701760
rect 433314 695138 433346 695374
rect 433582 695138 433666 695374
rect 433902 695138 433934 695374
rect 433314 695054 433934 695138
rect 433314 694818 433346 695054
rect 433582 694818 433666 695054
rect 433902 694818 433934 695054
rect 433314 658174 433934 694818
rect 433314 657938 433346 658174
rect 433582 657938 433666 658174
rect 433902 657938 433934 658174
rect 433314 657854 433934 657938
rect 433314 657618 433346 657854
rect 433582 657618 433666 657854
rect 433902 657618 433934 657854
rect 433314 620974 433934 657618
rect 433314 620738 433346 620974
rect 433582 620738 433666 620974
rect 433902 620738 433934 620974
rect 433314 620654 433934 620738
rect 433314 620418 433346 620654
rect 433582 620418 433666 620654
rect 433902 620418 433934 620654
rect 433314 583774 433934 620418
rect 433314 583538 433346 583774
rect 433582 583538 433666 583774
rect 433902 583538 433934 583774
rect 433314 583454 433934 583538
rect 433314 583218 433346 583454
rect 433582 583218 433666 583454
rect 433902 583218 433934 583454
rect 433314 546574 433934 583218
rect 433314 546338 433346 546574
rect 433582 546338 433666 546574
rect 433902 546338 433934 546574
rect 433314 546254 433934 546338
rect 433314 546018 433346 546254
rect 433582 546018 433666 546254
rect 433902 546018 433934 546254
rect 433314 509374 433934 546018
rect 433314 509138 433346 509374
rect 433582 509138 433666 509374
rect 433902 509138 433934 509374
rect 433314 509054 433934 509138
rect 433314 508818 433346 509054
rect 433582 508818 433666 509054
rect 433902 508818 433934 509054
rect 433314 472174 433934 508818
rect 433314 471938 433346 472174
rect 433582 471938 433666 472174
rect 433902 471938 433934 472174
rect 433314 471854 433934 471938
rect 433314 471618 433346 471854
rect 433582 471618 433666 471854
rect 433902 471618 433934 471854
rect 433314 434974 433934 471618
rect 433314 434738 433346 434974
rect 433582 434738 433666 434974
rect 433902 434738 433934 434974
rect 433314 434654 433934 434738
rect 433314 434418 433346 434654
rect 433582 434418 433666 434654
rect 433902 434418 433934 434654
rect 433314 397774 433934 434418
rect 433314 397538 433346 397774
rect 433582 397538 433666 397774
rect 433902 397538 433934 397774
rect 433314 397454 433934 397538
rect 433314 397218 433346 397454
rect 433582 397218 433666 397454
rect 433902 397218 433934 397454
rect 433314 360574 433934 397218
rect 433314 360338 433346 360574
rect 433582 360338 433666 360574
rect 433902 360338 433934 360574
rect 433314 360254 433934 360338
rect 433314 360018 433346 360254
rect 433582 360018 433666 360254
rect 433902 360018 433934 360254
rect 433314 323374 433934 360018
rect 433314 323138 433346 323374
rect 433582 323138 433666 323374
rect 433902 323138 433934 323374
rect 433314 323054 433934 323138
rect 433314 322818 433346 323054
rect 433582 322818 433666 323054
rect 433902 322818 433934 323054
rect 433314 286174 433934 322818
rect 433314 285938 433346 286174
rect 433582 285938 433666 286174
rect 433902 285938 433934 286174
rect 433314 285854 433934 285938
rect 433314 285618 433346 285854
rect 433582 285618 433666 285854
rect 433902 285618 433934 285854
rect 433314 248974 433934 285618
rect 433314 248738 433346 248974
rect 433582 248738 433666 248974
rect 433902 248738 433934 248974
rect 433314 248654 433934 248738
rect 433314 248418 433346 248654
rect 433582 248418 433666 248654
rect 433902 248418 433934 248654
rect 433314 211774 433934 248418
rect 433314 211538 433346 211774
rect 433582 211538 433666 211774
rect 433902 211538 433934 211774
rect 433314 211454 433934 211538
rect 433314 211218 433346 211454
rect 433582 211218 433666 211454
rect 433902 211218 433934 211454
rect 433314 174574 433934 211218
rect 433314 174338 433346 174574
rect 433582 174338 433666 174574
rect 433902 174338 433934 174574
rect 433314 174254 433934 174338
rect 433314 174018 433346 174254
rect 433582 174018 433666 174254
rect 433902 174018 433934 174254
rect 433314 137374 433934 174018
rect 433314 137138 433346 137374
rect 433582 137138 433666 137374
rect 433902 137138 433934 137374
rect 433314 137054 433934 137138
rect 433314 136818 433346 137054
rect 433582 136818 433666 137054
rect 433902 136818 433934 137054
rect 433314 100174 433934 136818
rect 433314 99938 433346 100174
rect 433582 99938 433666 100174
rect 433902 99938 433934 100174
rect 433314 99854 433934 99938
rect 433314 99618 433346 99854
rect 433582 99618 433666 99854
rect 433902 99618 433934 99854
rect 433314 62974 433934 99618
rect 433314 62738 433346 62974
rect 433582 62738 433666 62974
rect 433902 62738 433934 62974
rect 433314 62654 433934 62738
rect 433314 62418 433346 62654
rect 433582 62418 433666 62654
rect 433902 62418 433934 62654
rect 433314 25774 433934 62418
rect 433314 25538 433346 25774
rect 433582 25538 433666 25774
rect 433902 25538 433934 25774
rect 433314 25454 433934 25538
rect 433314 25218 433346 25454
rect 433582 25218 433666 25454
rect 433902 25218 433934 25454
rect 433314 2176 433934 25218
rect 437034 699094 437654 701760
rect 437034 698858 437066 699094
rect 437302 698858 437386 699094
rect 437622 698858 437654 699094
rect 437034 698774 437654 698858
rect 437034 698538 437066 698774
rect 437302 698538 437386 698774
rect 437622 698538 437654 698774
rect 437034 661894 437654 698538
rect 437034 661658 437066 661894
rect 437302 661658 437386 661894
rect 437622 661658 437654 661894
rect 437034 661574 437654 661658
rect 437034 661338 437066 661574
rect 437302 661338 437386 661574
rect 437622 661338 437654 661574
rect 437034 624694 437654 661338
rect 437034 624458 437066 624694
rect 437302 624458 437386 624694
rect 437622 624458 437654 624694
rect 437034 624374 437654 624458
rect 437034 624138 437066 624374
rect 437302 624138 437386 624374
rect 437622 624138 437654 624374
rect 437034 587494 437654 624138
rect 437034 587258 437066 587494
rect 437302 587258 437386 587494
rect 437622 587258 437654 587494
rect 437034 587174 437654 587258
rect 437034 586938 437066 587174
rect 437302 586938 437386 587174
rect 437622 586938 437654 587174
rect 437034 550294 437654 586938
rect 437034 550058 437066 550294
rect 437302 550058 437386 550294
rect 437622 550058 437654 550294
rect 437034 549974 437654 550058
rect 437034 549738 437066 549974
rect 437302 549738 437386 549974
rect 437622 549738 437654 549974
rect 437034 513094 437654 549738
rect 437034 512858 437066 513094
rect 437302 512858 437386 513094
rect 437622 512858 437654 513094
rect 437034 512774 437654 512858
rect 437034 512538 437066 512774
rect 437302 512538 437386 512774
rect 437622 512538 437654 512774
rect 437034 475894 437654 512538
rect 437034 475658 437066 475894
rect 437302 475658 437386 475894
rect 437622 475658 437654 475894
rect 437034 475574 437654 475658
rect 437034 475338 437066 475574
rect 437302 475338 437386 475574
rect 437622 475338 437654 475574
rect 437034 438694 437654 475338
rect 437034 438458 437066 438694
rect 437302 438458 437386 438694
rect 437622 438458 437654 438694
rect 437034 438374 437654 438458
rect 437034 438138 437066 438374
rect 437302 438138 437386 438374
rect 437622 438138 437654 438374
rect 437034 401494 437654 438138
rect 437034 401258 437066 401494
rect 437302 401258 437386 401494
rect 437622 401258 437654 401494
rect 437034 401174 437654 401258
rect 437034 400938 437066 401174
rect 437302 400938 437386 401174
rect 437622 400938 437654 401174
rect 437034 364294 437654 400938
rect 437034 364058 437066 364294
rect 437302 364058 437386 364294
rect 437622 364058 437654 364294
rect 437034 363974 437654 364058
rect 437034 363738 437066 363974
rect 437302 363738 437386 363974
rect 437622 363738 437654 363974
rect 437034 327094 437654 363738
rect 437034 326858 437066 327094
rect 437302 326858 437386 327094
rect 437622 326858 437654 327094
rect 437034 326774 437654 326858
rect 437034 326538 437066 326774
rect 437302 326538 437386 326774
rect 437622 326538 437654 326774
rect 437034 289894 437654 326538
rect 437034 289658 437066 289894
rect 437302 289658 437386 289894
rect 437622 289658 437654 289894
rect 437034 289574 437654 289658
rect 437034 289338 437066 289574
rect 437302 289338 437386 289574
rect 437622 289338 437654 289574
rect 437034 252694 437654 289338
rect 437034 252458 437066 252694
rect 437302 252458 437386 252694
rect 437622 252458 437654 252694
rect 437034 252374 437654 252458
rect 437034 252138 437066 252374
rect 437302 252138 437386 252374
rect 437622 252138 437654 252374
rect 437034 215494 437654 252138
rect 437034 215258 437066 215494
rect 437302 215258 437386 215494
rect 437622 215258 437654 215494
rect 437034 215174 437654 215258
rect 437034 214938 437066 215174
rect 437302 214938 437386 215174
rect 437622 214938 437654 215174
rect 437034 178294 437654 214938
rect 437034 178058 437066 178294
rect 437302 178058 437386 178294
rect 437622 178058 437654 178294
rect 437034 177974 437654 178058
rect 437034 177738 437066 177974
rect 437302 177738 437386 177974
rect 437622 177738 437654 177974
rect 437034 141094 437654 177738
rect 437034 140858 437066 141094
rect 437302 140858 437386 141094
rect 437622 140858 437654 141094
rect 437034 140774 437654 140858
rect 437034 140538 437066 140774
rect 437302 140538 437386 140774
rect 437622 140538 437654 140774
rect 437034 103894 437654 140538
rect 437034 103658 437066 103894
rect 437302 103658 437386 103894
rect 437622 103658 437654 103894
rect 437034 103574 437654 103658
rect 437034 103338 437066 103574
rect 437302 103338 437386 103574
rect 437622 103338 437654 103574
rect 437034 66694 437654 103338
rect 437034 66458 437066 66694
rect 437302 66458 437386 66694
rect 437622 66458 437654 66694
rect 437034 66374 437654 66458
rect 437034 66138 437066 66374
rect 437302 66138 437386 66374
rect 437622 66138 437654 66374
rect 437034 29494 437654 66138
rect 437034 29258 437066 29494
rect 437302 29258 437386 29494
rect 437622 29258 437654 29494
rect 437034 29174 437654 29258
rect 437034 28938 437066 29174
rect 437302 28938 437386 29174
rect 437622 28938 437654 29174
rect 437034 2176 437654 28938
rect 448194 673054 448814 701760
rect 448194 672818 448226 673054
rect 448462 672818 448546 673054
rect 448782 672818 448814 673054
rect 448194 672734 448814 672818
rect 448194 672498 448226 672734
rect 448462 672498 448546 672734
rect 448782 672498 448814 672734
rect 448194 635854 448814 672498
rect 448194 635618 448226 635854
rect 448462 635618 448546 635854
rect 448782 635618 448814 635854
rect 448194 635534 448814 635618
rect 448194 635298 448226 635534
rect 448462 635298 448546 635534
rect 448782 635298 448814 635534
rect 448194 598654 448814 635298
rect 448194 598418 448226 598654
rect 448462 598418 448546 598654
rect 448782 598418 448814 598654
rect 448194 598334 448814 598418
rect 448194 598098 448226 598334
rect 448462 598098 448546 598334
rect 448782 598098 448814 598334
rect 448194 561454 448814 598098
rect 448194 561218 448226 561454
rect 448462 561218 448546 561454
rect 448782 561218 448814 561454
rect 448194 561134 448814 561218
rect 448194 560898 448226 561134
rect 448462 560898 448546 561134
rect 448782 560898 448814 561134
rect 448194 524254 448814 560898
rect 448194 524018 448226 524254
rect 448462 524018 448546 524254
rect 448782 524018 448814 524254
rect 448194 523934 448814 524018
rect 448194 523698 448226 523934
rect 448462 523698 448546 523934
rect 448782 523698 448814 523934
rect 448194 487054 448814 523698
rect 448194 486818 448226 487054
rect 448462 486818 448546 487054
rect 448782 486818 448814 487054
rect 448194 486734 448814 486818
rect 448194 486498 448226 486734
rect 448462 486498 448546 486734
rect 448782 486498 448814 486734
rect 448194 449854 448814 486498
rect 448194 449618 448226 449854
rect 448462 449618 448546 449854
rect 448782 449618 448814 449854
rect 448194 449534 448814 449618
rect 448194 449298 448226 449534
rect 448462 449298 448546 449534
rect 448782 449298 448814 449534
rect 448194 412654 448814 449298
rect 448194 412418 448226 412654
rect 448462 412418 448546 412654
rect 448782 412418 448814 412654
rect 448194 412334 448814 412418
rect 448194 412098 448226 412334
rect 448462 412098 448546 412334
rect 448782 412098 448814 412334
rect 448194 375454 448814 412098
rect 448194 375218 448226 375454
rect 448462 375218 448546 375454
rect 448782 375218 448814 375454
rect 448194 375134 448814 375218
rect 448194 374898 448226 375134
rect 448462 374898 448546 375134
rect 448782 374898 448814 375134
rect 448194 338254 448814 374898
rect 448194 338018 448226 338254
rect 448462 338018 448546 338254
rect 448782 338018 448814 338254
rect 448194 337934 448814 338018
rect 448194 337698 448226 337934
rect 448462 337698 448546 337934
rect 448782 337698 448814 337934
rect 448194 301054 448814 337698
rect 448194 300818 448226 301054
rect 448462 300818 448546 301054
rect 448782 300818 448814 301054
rect 448194 300734 448814 300818
rect 448194 300498 448226 300734
rect 448462 300498 448546 300734
rect 448782 300498 448814 300734
rect 448194 263854 448814 300498
rect 448194 263618 448226 263854
rect 448462 263618 448546 263854
rect 448782 263618 448814 263854
rect 448194 263534 448814 263618
rect 448194 263298 448226 263534
rect 448462 263298 448546 263534
rect 448782 263298 448814 263534
rect 448194 226654 448814 263298
rect 448194 226418 448226 226654
rect 448462 226418 448546 226654
rect 448782 226418 448814 226654
rect 448194 226334 448814 226418
rect 448194 226098 448226 226334
rect 448462 226098 448546 226334
rect 448782 226098 448814 226334
rect 448194 189454 448814 226098
rect 448194 189218 448226 189454
rect 448462 189218 448546 189454
rect 448782 189218 448814 189454
rect 448194 189134 448814 189218
rect 448194 188898 448226 189134
rect 448462 188898 448546 189134
rect 448782 188898 448814 189134
rect 448194 152254 448814 188898
rect 448194 152018 448226 152254
rect 448462 152018 448546 152254
rect 448782 152018 448814 152254
rect 448194 151934 448814 152018
rect 448194 151698 448226 151934
rect 448462 151698 448546 151934
rect 448782 151698 448814 151934
rect 448194 115054 448814 151698
rect 448194 114818 448226 115054
rect 448462 114818 448546 115054
rect 448782 114818 448814 115054
rect 448194 114734 448814 114818
rect 448194 114498 448226 114734
rect 448462 114498 448546 114734
rect 448782 114498 448814 114734
rect 448194 77854 448814 114498
rect 448194 77618 448226 77854
rect 448462 77618 448546 77854
rect 448782 77618 448814 77854
rect 448194 77534 448814 77618
rect 448194 77298 448226 77534
rect 448462 77298 448546 77534
rect 448782 77298 448814 77534
rect 448194 40654 448814 77298
rect 448194 40418 448226 40654
rect 448462 40418 448546 40654
rect 448782 40418 448814 40654
rect 448194 40334 448814 40418
rect 448194 40098 448226 40334
rect 448462 40098 448546 40334
rect 448782 40098 448814 40334
rect 448194 3454 448814 40098
rect 448194 3218 448226 3454
rect 448462 3218 448546 3454
rect 448782 3218 448814 3454
rect 448194 3134 448814 3218
rect 448194 2898 448226 3134
rect 448462 2898 448546 3134
rect 448782 2898 448814 3134
rect 448194 2176 448814 2898
rect 451914 676774 452534 701760
rect 451914 676538 451946 676774
rect 452182 676538 452266 676774
rect 452502 676538 452534 676774
rect 451914 676454 452534 676538
rect 451914 676218 451946 676454
rect 452182 676218 452266 676454
rect 452502 676218 452534 676454
rect 451914 639574 452534 676218
rect 451914 639338 451946 639574
rect 452182 639338 452266 639574
rect 452502 639338 452534 639574
rect 451914 639254 452534 639338
rect 451914 639018 451946 639254
rect 452182 639018 452266 639254
rect 452502 639018 452534 639254
rect 451914 602374 452534 639018
rect 451914 602138 451946 602374
rect 452182 602138 452266 602374
rect 452502 602138 452534 602374
rect 451914 602054 452534 602138
rect 451914 601818 451946 602054
rect 452182 601818 452266 602054
rect 452502 601818 452534 602054
rect 451914 565174 452534 601818
rect 451914 564938 451946 565174
rect 452182 564938 452266 565174
rect 452502 564938 452534 565174
rect 451914 564854 452534 564938
rect 451914 564618 451946 564854
rect 452182 564618 452266 564854
rect 452502 564618 452534 564854
rect 451914 527974 452534 564618
rect 451914 527738 451946 527974
rect 452182 527738 452266 527974
rect 452502 527738 452534 527974
rect 451914 527654 452534 527738
rect 451914 527418 451946 527654
rect 452182 527418 452266 527654
rect 452502 527418 452534 527654
rect 451914 490774 452534 527418
rect 451914 490538 451946 490774
rect 452182 490538 452266 490774
rect 452502 490538 452534 490774
rect 451914 490454 452534 490538
rect 451914 490218 451946 490454
rect 452182 490218 452266 490454
rect 452502 490218 452534 490454
rect 451914 453574 452534 490218
rect 451914 453338 451946 453574
rect 452182 453338 452266 453574
rect 452502 453338 452534 453574
rect 451914 453254 452534 453338
rect 451914 453018 451946 453254
rect 452182 453018 452266 453254
rect 452502 453018 452534 453254
rect 451914 416374 452534 453018
rect 451914 416138 451946 416374
rect 452182 416138 452266 416374
rect 452502 416138 452534 416374
rect 451914 416054 452534 416138
rect 451914 415818 451946 416054
rect 452182 415818 452266 416054
rect 452502 415818 452534 416054
rect 451914 379174 452534 415818
rect 451914 378938 451946 379174
rect 452182 378938 452266 379174
rect 452502 378938 452534 379174
rect 451914 378854 452534 378938
rect 451914 378618 451946 378854
rect 452182 378618 452266 378854
rect 452502 378618 452534 378854
rect 451914 341974 452534 378618
rect 451914 341738 451946 341974
rect 452182 341738 452266 341974
rect 452502 341738 452534 341974
rect 451914 341654 452534 341738
rect 451914 341418 451946 341654
rect 452182 341418 452266 341654
rect 452502 341418 452534 341654
rect 451914 304774 452534 341418
rect 451914 304538 451946 304774
rect 452182 304538 452266 304774
rect 452502 304538 452534 304774
rect 451914 304454 452534 304538
rect 451914 304218 451946 304454
rect 452182 304218 452266 304454
rect 452502 304218 452534 304454
rect 451914 267574 452534 304218
rect 451914 267338 451946 267574
rect 452182 267338 452266 267574
rect 452502 267338 452534 267574
rect 451914 267254 452534 267338
rect 451914 267018 451946 267254
rect 452182 267018 452266 267254
rect 452502 267018 452534 267254
rect 451914 230374 452534 267018
rect 451914 230138 451946 230374
rect 452182 230138 452266 230374
rect 452502 230138 452534 230374
rect 451914 230054 452534 230138
rect 451914 229818 451946 230054
rect 452182 229818 452266 230054
rect 452502 229818 452534 230054
rect 451914 193174 452534 229818
rect 451914 192938 451946 193174
rect 452182 192938 452266 193174
rect 452502 192938 452534 193174
rect 451914 192854 452534 192938
rect 451914 192618 451946 192854
rect 452182 192618 452266 192854
rect 452502 192618 452534 192854
rect 451914 155974 452534 192618
rect 451914 155738 451946 155974
rect 452182 155738 452266 155974
rect 452502 155738 452534 155974
rect 451914 155654 452534 155738
rect 451914 155418 451946 155654
rect 452182 155418 452266 155654
rect 452502 155418 452534 155654
rect 451914 118774 452534 155418
rect 451914 118538 451946 118774
rect 452182 118538 452266 118774
rect 452502 118538 452534 118774
rect 451914 118454 452534 118538
rect 451914 118218 451946 118454
rect 452182 118218 452266 118454
rect 452502 118218 452534 118454
rect 451914 81574 452534 118218
rect 451914 81338 451946 81574
rect 452182 81338 452266 81574
rect 452502 81338 452534 81574
rect 451914 81254 452534 81338
rect 451914 81018 451946 81254
rect 452182 81018 452266 81254
rect 452502 81018 452534 81254
rect 451914 44374 452534 81018
rect 451914 44138 451946 44374
rect 452182 44138 452266 44374
rect 452502 44138 452534 44374
rect 451914 44054 452534 44138
rect 451914 43818 451946 44054
rect 452182 43818 452266 44054
rect 452502 43818 452534 44054
rect 451914 7174 452534 43818
rect 451914 6938 451946 7174
rect 452182 6938 452266 7174
rect 452502 6938 452534 7174
rect 451914 6854 452534 6938
rect 451914 6618 451946 6854
rect 452182 6618 452266 6854
rect 452502 6618 452534 6854
rect 451914 2176 452534 6618
rect 455634 680494 456254 701760
rect 455634 680258 455666 680494
rect 455902 680258 455986 680494
rect 456222 680258 456254 680494
rect 455634 680174 456254 680258
rect 455634 679938 455666 680174
rect 455902 679938 455986 680174
rect 456222 679938 456254 680174
rect 455634 643294 456254 679938
rect 455634 643058 455666 643294
rect 455902 643058 455986 643294
rect 456222 643058 456254 643294
rect 455634 642974 456254 643058
rect 455634 642738 455666 642974
rect 455902 642738 455986 642974
rect 456222 642738 456254 642974
rect 455634 606094 456254 642738
rect 455634 605858 455666 606094
rect 455902 605858 455986 606094
rect 456222 605858 456254 606094
rect 455634 605774 456254 605858
rect 455634 605538 455666 605774
rect 455902 605538 455986 605774
rect 456222 605538 456254 605774
rect 455634 568894 456254 605538
rect 455634 568658 455666 568894
rect 455902 568658 455986 568894
rect 456222 568658 456254 568894
rect 455634 568574 456254 568658
rect 455634 568338 455666 568574
rect 455902 568338 455986 568574
rect 456222 568338 456254 568574
rect 455634 531694 456254 568338
rect 455634 531458 455666 531694
rect 455902 531458 455986 531694
rect 456222 531458 456254 531694
rect 455634 531374 456254 531458
rect 455634 531138 455666 531374
rect 455902 531138 455986 531374
rect 456222 531138 456254 531374
rect 455634 494494 456254 531138
rect 455634 494258 455666 494494
rect 455902 494258 455986 494494
rect 456222 494258 456254 494494
rect 455634 494174 456254 494258
rect 455634 493938 455666 494174
rect 455902 493938 455986 494174
rect 456222 493938 456254 494174
rect 455634 457294 456254 493938
rect 455634 457058 455666 457294
rect 455902 457058 455986 457294
rect 456222 457058 456254 457294
rect 455634 456974 456254 457058
rect 455634 456738 455666 456974
rect 455902 456738 455986 456974
rect 456222 456738 456254 456974
rect 455634 420094 456254 456738
rect 455634 419858 455666 420094
rect 455902 419858 455986 420094
rect 456222 419858 456254 420094
rect 455634 419774 456254 419858
rect 455634 419538 455666 419774
rect 455902 419538 455986 419774
rect 456222 419538 456254 419774
rect 455634 382894 456254 419538
rect 455634 382658 455666 382894
rect 455902 382658 455986 382894
rect 456222 382658 456254 382894
rect 455634 382574 456254 382658
rect 455634 382338 455666 382574
rect 455902 382338 455986 382574
rect 456222 382338 456254 382574
rect 455634 345694 456254 382338
rect 455634 345458 455666 345694
rect 455902 345458 455986 345694
rect 456222 345458 456254 345694
rect 455634 345374 456254 345458
rect 455634 345138 455666 345374
rect 455902 345138 455986 345374
rect 456222 345138 456254 345374
rect 455634 308494 456254 345138
rect 455634 308258 455666 308494
rect 455902 308258 455986 308494
rect 456222 308258 456254 308494
rect 455634 308174 456254 308258
rect 455634 307938 455666 308174
rect 455902 307938 455986 308174
rect 456222 307938 456254 308174
rect 455634 271294 456254 307938
rect 455634 271058 455666 271294
rect 455902 271058 455986 271294
rect 456222 271058 456254 271294
rect 455634 270974 456254 271058
rect 455634 270738 455666 270974
rect 455902 270738 455986 270974
rect 456222 270738 456254 270974
rect 455634 234094 456254 270738
rect 455634 233858 455666 234094
rect 455902 233858 455986 234094
rect 456222 233858 456254 234094
rect 455634 233774 456254 233858
rect 455634 233538 455666 233774
rect 455902 233538 455986 233774
rect 456222 233538 456254 233774
rect 455634 196894 456254 233538
rect 455634 196658 455666 196894
rect 455902 196658 455986 196894
rect 456222 196658 456254 196894
rect 455634 196574 456254 196658
rect 455634 196338 455666 196574
rect 455902 196338 455986 196574
rect 456222 196338 456254 196574
rect 455634 159694 456254 196338
rect 455634 159458 455666 159694
rect 455902 159458 455986 159694
rect 456222 159458 456254 159694
rect 455634 159374 456254 159458
rect 455634 159138 455666 159374
rect 455902 159138 455986 159374
rect 456222 159138 456254 159374
rect 455634 122494 456254 159138
rect 455634 122258 455666 122494
rect 455902 122258 455986 122494
rect 456222 122258 456254 122494
rect 455634 122174 456254 122258
rect 455634 121938 455666 122174
rect 455902 121938 455986 122174
rect 456222 121938 456254 122174
rect 455634 85294 456254 121938
rect 455634 85058 455666 85294
rect 455902 85058 455986 85294
rect 456222 85058 456254 85294
rect 455634 84974 456254 85058
rect 455634 84738 455666 84974
rect 455902 84738 455986 84974
rect 456222 84738 456254 84974
rect 455634 48094 456254 84738
rect 455634 47858 455666 48094
rect 455902 47858 455986 48094
rect 456222 47858 456254 48094
rect 455634 47774 456254 47858
rect 455634 47538 455666 47774
rect 455902 47538 455986 47774
rect 456222 47538 456254 47774
rect 455634 10894 456254 47538
rect 455634 10658 455666 10894
rect 455902 10658 455986 10894
rect 456222 10658 456254 10894
rect 455634 10574 456254 10658
rect 455634 10338 455666 10574
rect 455902 10338 455986 10574
rect 456222 10338 456254 10574
rect 455634 2176 456254 10338
rect 459354 684214 459974 701760
rect 459354 683978 459386 684214
rect 459622 683978 459706 684214
rect 459942 683978 459974 684214
rect 459354 683894 459974 683978
rect 459354 683658 459386 683894
rect 459622 683658 459706 683894
rect 459942 683658 459974 683894
rect 459354 647014 459974 683658
rect 459354 646778 459386 647014
rect 459622 646778 459706 647014
rect 459942 646778 459974 647014
rect 459354 646694 459974 646778
rect 459354 646458 459386 646694
rect 459622 646458 459706 646694
rect 459942 646458 459974 646694
rect 459354 609814 459974 646458
rect 459354 609578 459386 609814
rect 459622 609578 459706 609814
rect 459942 609578 459974 609814
rect 459354 609494 459974 609578
rect 459354 609258 459386 609494
rect 459622 609258 459706 609494
rect 459942 609258 459974 609494
rect 459354 572614 459974 609258
rect 459354 572378 459386 572614
rect 459622 572378 459706 572614
rect 459942 572378 459974 572614
rect 459354 572294 459974 572378
rect 459354 572058 459386 572294
rect 459622 572058 459706 572294
rect 459942 572058 459974 572294
rect 459354 535414 459974 572058
rect 459354 535178 459386 535414
rect 459622 535178 459706 535414
rect 459942 535178 459974 535414
rect 459354 535094 459974 535178
rect 459354 534858 459386 535094
rect 459622 534858 459706 535094
rect 459942 534858 459974 535094
rect 459354 498214 459974 534858
rect 459354 497978 459386 498214
rect 459622 497978 459706 498214
rect 459942 497978 459974 498214
rect 459354 497894 459974 497978
rect 459354 497658 459386 497894
rect 459622 497658 459706 497894
rect 459942 497658 459974 497894
rect 459354 461014 459974 497658
rect 459354 460778 459386 461014
rect 459622 460778 459706 461014
rect 459942 460778 459974 461014
rect 459354 460694 459974 460778
rect 459354 460458 459386 460694
rect 459622 460458 459706 460694
rect 459942 460458 459974 460694
rect 459354 423814 459974 460458
rect 459354 423578 459386 423814
rect 459622 423578 459706 423814
rect 459942 423578 459974 423814
rect 459354 423494 459974 423578
rect 459354 423258 459386 423494
rect 459622 423258 459706 423494
rect 459942 423258 459974 423494
rect 459354 386614 459974 423258
rect 459354 386378 459386 386614
rect 459622 386378 459706 386614
rect 459942 386378 459974 386614
rect 459354 386294 459974 386378
rect 459354 386058 459386 386294
rect 459622 386058 459706 386294
rect 459942 386058 459974 386294
rect 459354 349414 459974 386058
rect 459354 349178 459386 349414
rect 459622 349178 459706 349414
rect 459942 349178 459974 349414
rect 459354 349094 459974 349178
rect 459354 348858 459386 349094
rect 459622 348858 459706 349094
rect 459942 348858 459974 349094
rect 459354 312214 459974 348858
rect 459354 311978 459386 312214
rect 459622 311978 459706 312214
rect 459942 311978 459974 312214
rect 459354 311894 459974 311978
rect 459354 311658 459386 311894
rect 459622 311658 459706 311894
rect 459942 311658 459974 311894
rect 459354 275014 459974 311658
rect 459354 274778 459386 275014
rect 459622 274778 459706 275014
rect 459942 274778 459974 275014
rect 459354 274694 459974 274778
rect 459354 274458 459386 274694
rect 459622 274458 459706 274694
rect 459942 274458 459974 274694
rect 459354 237814 459974 274458
rect 459354 237578 459386 237814
rect 459622 237578 459706 237814
rect 459942 237578 459974 237814
rect 459354 237494 459974 237578
rect 459354 237258 459386 237494
rect 459622 237258 459706 237494
rect 459942 237258 459974 237494
rect 459354 200614 459974 237258
rect 459354 200378 459386 200614
rect 459622 200378 459706 200614
rect 459942 200378 459974 200614
rect 459354 200294 459974 200378
rect 459354 200058 459386 200294
rect 459622 200058 459706 200294
rect 459942 200058 459974 200294
rect 459354 163414 459974 200058
rect 459354 163178 459386 163414
rect 459622 163178 459706 163414
rect 459942 163178 459974 163414
rect 459354 163094 459974 163178
rect 459354 162858 459386 163094
rect 459622 162858 459706 163094
rect 459942 162858 459974 163094
rect 459354 126214 459974 162858
rect 459354 125978 459386 126214
rect 459622 125978 459706 126214
rect 459942 125978 459974 126214
rect 459354 125894 459974 125978
rect 459354 125658 459386 125894
rect 459622 125658 459706 125894
rect 459942 125658 459974 125894
rect 459354 89014 459974 125658
rect 459354 88778 459386 89014
rect 459622 88778 459706 89014
rect 459942 88778 459974 89014
rect 459354 88694 459974 88778
rect 459354 88458 459386 88694
rect 459622 88458 459706 88694
rect 459942 88458 459974 88694
rect 459354 51814 459974 88458
rect 459354 51578 459386 51814
rect 459622 51578 459706 51814
rect 459942 51578 459974 51814
rect 459354 51494 459974 51578
rect 459354 51258 459386 51494
rect 459622 51258 459706 51494
rect 459942 51258 459974 51494
rect 459354 14614 459974 51258
rect 459354 14378 459386 14614
rect 459622 14378 459706 14614
rect 459942 14378 459974 14614
rect 459354 14294 459974 14378
rect 459354 14058 459386 14294
rect 459622 14058 459706 14294
rect 459942 14058 459974 14294
rect 459354 2176 459974 14058
rect 463074 687934 463694 701760
rect 463074 687698 463106 687934
rect 463342 687698 463426 687934
rect 463662 687698 463694 687934
rect 463074 687614 463694 687698
rect 463074 687378 463106 687614
rect 463342 687378 463426 687614
rect 463662 687378 463694 687614
rect 463074 650734 463694 687378
rect 463074 650498 463106 650734
rect 463342 650498 463426 650734
rect 463662 650498 463694 650734
rect 463074 650414 463694 650498
rect 463074 650178 463106 650414
rect 463342 650178 463426 650414
rect 463662 650178 463694 650414
rect 463074 613534 463694 650178
rect 463074 613298 463106 613534
rect 463342 613298 463426 613534
rect 463662 613298 463694 613534
rect 463074 613214 463694 613298
rect 463074 612978 463106 613214
rect 463342 612978 463426 613214
rect 463662 612978 463694 613214
rect 463074 576334 463694 612978
rect 463074 576098 463106 576334
rect 463342 576098 463426 576334
rect 463662 576098 463694 576334
rect 463074 576014 463694 576098
rect 463074 575778 463106 576014
rect 463342 575778 463426 576014
rect 463662 575778 463694 576014
rect 463074 539134 463694 575778
rect 463074 538898 463106 539134
rect 463342 538898 463426 539134
rect 463662 538898 463694 539134
rect 463074 538814 463694 538898
rect 463074 538578 463106 538814
rect 463342 538578 463426 538814
rect 463662 538578 463694 538814
rect 463074 501934 463694 538578
rect 463074 501698 463106 501934
rect 463342 501698 463426 501934
rect 463662 501698 463694 501934
rect 463074 501614 463694 501698
rect 463074 501378 463106 501614
rect 463342 501378 463426 501614
rect 463662 501378 463694 501614
rect 463074 464734 463694 501378
rect 463074 464498 463106 464734
rect 463342 464498 463426 464734
rect 463662 464498 463694 464734
rect 463074 464414 463694 464498
rect 463074 464178 463106 464414
rect 463342 464178 463426 464414
rect 463662 464178 463694 464414
rect 463074 427534 463694 464178
rect 463074 427298 463106 427534
rect 463342 427298 463426 427534
rect 463662 427298 463694 427534
rect 463074 427214 463694 427298
rect 463074 426978 463106 427214
rect 463342 426978 463426 427214
rect 463662 426978 463694 427214
rect 463074 390334 463694 426978
rect 463074 390098 463106 390334
rect 463342 390098 463426 390334
rect 463662 390098 463694 390334
rect 463074 390014 463694 390098
rect 463074 389778 463106 390014
rect 463342 389778 463426 390014
rect 463662 389778 463694 390014
rect 463074 353134 463694 389778
rect 463074 352898 463106 353134
rect 463342 352898 463426 353134
rect 463662 352898 463694 353134
rect 463074 352814 463694 352898
rect 463074 352578 463106 352814
rect 463342 352578 463426 352814
rect 463662 352578 463694 352814
rect 463074 315934 463694 352578
rect 463074 315698 463106 315934
rect 463342 315698 463426 315934
rect 463662 315698 463694 315934
rect 463074 315614 463694 315698
rect 463074 315378 463106 315614
rect 463342 315378 463426 315614
rect 463662 315378 463694 315614
rect 463074 278734 463694 315378
rect 463074 278498 463106 278734
rect 463342 278498 463426 278734
rect 463662 278498 463694 278734
rect 463074 278414 463694 278498
rect 463074 278178 463106 278414
rect 463342 278178 463426 278414
rect 463662 278178 463694 278414
rect 463074 241534 463694 278178
rect 463074 241298 463106 241534
rect 463342 241298 463426 241534
rect 463662 241298 463694 241534
rect 463074 241214 463694 241298
rect 463074 240978 463106 241214
rect 463342 240978 463426 241214
rect 463662 240978 463694 241214
rect 463074 204334 463694 240978
rect 463074 204098 463106 204334
rect 463342 204098 463426 204334
rect 463662 204098 463694 204334
rect 463074 204014 463694 204098
rect 463074 203778 463106 204014
rect 463342 203778 463426 204014
rect 463662 203778 463694 204014
rect 463074 167134 463694 203778
rect 463074 166898 463106 167134
rect 463342 166898 463426 167134
rect 463662 166898 463694 167134
rect 463074 166814 463694 166898
rect 463074 166578 463106 166814
rect 463342 166578 463426 166814
rect 463662 166578 463694 166814
rect 463074 129934 463694 166578
rect 463074 129698 463106 129934
rect 463342 129698 463426 129934
rect 463662 129698 463694 129934
rect 463074 129614 463694 129698
rect 463074 129378 463106 129614
rect 463342 129378 463426 129614
rect 463662 129378 463694 129614
rect 463074 92734 463694 129378
rect 463074 92498 463106 92734
rect 463342 92498 463426 92734
rect 463662 92498 463694 92734
rect 463074 92414 463694 92498
rect 463074 92178 463106 92414
rect 463342 92178 463426 92414
rect 463662 92178 463694 92414
rect 463074 55534 463694 92178
rect 463074 55298 463106 55534
rect 463342 55298 463426 55534
rect 463662 55298 463694 55534
rect 463074 55214 463694 55298
rect 463074 54978 463106 55214
rect 463342 54978 463426 55214
rect 463662 54978 463694 55214
rect 463074 18334 463694 54978
rect 463074 18098 463106 18334
rect 463342 18098 463426 18334
rect 463662 18098 463694 18334
rect 463074 18014 463694 18098
rect 463074 17778 463106 18014
rect 463342 17778 463426 18014
rect 463662 17778 463694 18014
rect 463074 2176 463694 17778
rect 466794 691654 467414 701760
rect 466794 691418 466826 691654
rect 467062 691418 467146 691654
rect 467382 691418 467414 691654
rect 466794 691334 467414 691418
rect 466794 691098 466826 691334
rect 467062 691098 467146 691334
rect 467382 691098 467414 691334
rect 466794 654454 467414 691098
rect 466794 654218 466826 654454
rect 467062 654218 467146 654454
rect 467382 654218 467414 654454
rect 466794 654134 467414 654218
rect 466794 653898 466826 654134
rect 467062 653898 467146 654134
rect 467382 653898 467414 654134
rect 466794 617254 467414 653898
rect 466794 617018 466826 617254
rect 467062 617018 467146 617254
rect 467382 617018 467414 617254
rect 466794 616934 467414 617018
rect 466794 616698 466826 616934
rect 467062 616698 467146 616934
rect 467382 616698 467414 616934
rect 466794 580054 467414 616698
rect 466794 579818 466826 580054
rect 467062 579818 467146 580054
rect 467382 579818 467414 580054
rect 466794 579734 467414 579818
rect 466794 579498 466826 579734
rect 467062 579498 467146 579734
rect 467382 579498 467414 579734
rect 466794 542854 467414 579498
rect 466794 542618 466826 542854
rect 467062 542618 467146 542854
rect 467382 542618 467414 542854
rect 466794 542534 467414 542618
rect 466794 542298 466826 542534
rect 467062 542298 467146 542534
rect 467382 542298 467414 542534
rect 466794 505654 467414 542298
rect 466794 505418 466826 505654
rect 467062 505418 467146 505654
rect 467382 505418 467414 505654
rect 466794 505334 467414 505418
rect 466794 505098 466826 505334
rect 467062 505098 467146 505334
rect 467382 505098 467414 505334
rect 466794 468454 467414 505098
rect 466794 468218 466826 468454
rect 467062 468218 467146 468454
rect 467382 468218 467414 468454
rect 466794 468134 467414 468218
rect 466794 467898 466826 468134
rect 467062 467898 467146 468134
rect 467382 467898 467414 468134
rect 466794 431254 467414 467898
rect 466794 431018 466826 431254
rect 467062 431018 467146 431254
rect 467382 431018 467414 431254
rect 466794 430934 467414 431018
rect 466794 430698 466826 430934
rect 467062 430698 467146 430934
rect 467382 430698 467414 430934
rect 466794 394054 467414 430698
rect 466794 393818 466826 394054
rect 467062 393818 467146 394054
rect 467382 393818 467414 394054
rect 466794 393734 467414 393818
rect 466794 393498 466826 393734
rect 467062 393498 467146 393734
rect 467382 393498 467414 393734
rect 466794 356854 467414 393498
rect 466794 356618 466826 356854
rect 467062 356618 467146 356854
rect 467382 356618 467414 356854
rect 466794 356534 467414 356618
rect 466794 356298 466826 356534
rect 467062 356298 467146 356534
rect 467382 356298 467414 356534
rect 466794 319654 467414 356298
rect 466794 319418 466826 319654
rect 467062 319418 467146 319654
rect 467382 319418 467414 319654
rect 466794 319334 467414 319418
rect 466794 319098 466826 319334
rect 467062 319098 467146 319334
rect 467382 319098 467414 319334
rect 466794 282454 467414 319098
rect 466794 282218 466826 282454
rect 467062 282218 467146 282454
rect 467382 282218 467414 282454
rect 466794 282134 467414 282218
rect 466794 281898 466826 282134
rect 467062 281898 467146 282134
rect 467382 281898 467414 282134
rect 466794 245254 467414 281898
rect 466794 245018 466826 245254
rect 467062 245018 467146 245254
rect 467382 245018 467414 245254
rect 466794 244934 467414 245018
rect 466794 244698 466826 244934
rect 467062 244698 467146 244934
rect 467382 244698 467414 244934
rect 466794 208054 467414 244698
rect 466794 207818 466826 208054
rect 467062 207818 467146 208054
rect 467382 207818 467414 208054
rect 466794 207734 467414 207818
rect 466794 207498 466826 207734
rect 467062 207498 467146 207734
rect 467382 207498 467414 207734
rect 466794 170854 467414 207498
rect 466794 170618 466826 170854
rect 467062 170618 467146 170854
rect 467382 170618 467414 170854
rect 466794 170534 467414 170618
rect 466794 170298 466826 170534
rect 467062 170298 467146 170534
rect 467382 170298 467414 170534
rect 466794 133654 467414 170298
rect 466794 133418 466826 133654
rect 467062 133418 467146 133654
rect 467382 133418 467414 133654
rect 466794 133334 467414 133418
rect 466794 133098 466826 133334
rect 467062 133098 467146 133334
rect 467382 133098 467414 133334
rect 466794 96454 467414 133098
rect 466794 96218 466826 96454
rect 467062 96218 467146 96454
rect 467382 96218 467414 96454
rect 466794 96134 467414 96218
rect 466794 95898 466826 96134
rect 467062 95898 467146 96134
rect 467382 95898 467414 96134
rect 466794 59254 467414 95898
rect 466794 59018 466826 59254
rect 467062 59018 467146 59254
rect 467382 59018 467414 59254
rect 466794 58934 467414 59018
rect 466794 58698 466826 58934
rect 467062 58698 467146 58934
rect 467382 58698 467414 58934
rect 466794 22054 467414 58698
rect 466794 21818 466826 22054
rect 467062 21818 467146 22054
rect 467382 21818 467414 22054
rect 466794 21734 467414 21818
rect 466794 21498 466826 21734
rect 467062 21498 467146 21734
rect 467382 21498 467414 21734
rect 466794 2176 467414 21498
rect 470514 695374 471134 701760
rect 470514 695138 470546 695374
rect 470782 695138 470866 695374
rect 471102 695138 471134 695374
rect 470514 695054 471134 695138
rect 470514 694818 470546 695054
rect 470782 694818 470866 695054
rect 471102 694818 471134 695054
rect 470514 658174 471134 694818
rect 470514 657938 470546 658174
rect 470782 657938 470866 658174
rect 471102 657938 471134 658174
rect 470514 657854 471134 657938
rect 470514 657618 470546 657854
rect 470782 657618 470866 657854
rect 471102 657618 471134 657854
rect 470514 620974 471134 657618
rect 470514 620738 470546 620974
rect 470782 620738 470866 620974
rect 471102 620738 471134 620974
rect 470514 620654 471134 620738
rect 470514 620418 470546 620654
rect 470782 620418 470866 620654
rect 471102 620418 471134 620654
rect 470514 583774 471134 620418
rect 470514 583538 470546 583774
rect 470782 583538 470866 583774
rect 471102 583538 471134 583774
rect 470514 583454 471134 583538
rect 470514 583218 470546 583454
rect 470782 583218 470866 583454
rect 471102 583218 471134 583454
rect 470514 546574 471134 583218
rect 470514 546338 470546 546574
rect 470782 546338 470866 546574
rect 471102 546338 471134 546574
rect 470514 546254 471134 546338
rect 470514 546018 470546 546254
rect 470782 546018 470866 546254
rect 471102 546018 471134 546254
rect 470514 509374 471134 546018
rect 470514 509138 470546 509374
rect 470782 509138 470866 509374
rect 471102 509138 471134 509374
rect 470514 509054 471134 509138
rect 470514 508818 470546 509054
rect 470782 508818 470866 509054
rect 471102 508818 471134 509054
rect 470514 472174 471134 508818
rect 470514 471938 470546 472174
rect 470782 471938 470866 472174
rect 471102 471938 471134 472174
rect 470514 471854 471134 471938
rect 470514 471618 470546 471854
rect 470782 471618 470866 471854
rect 471102 471618 471134 471854
rect 470514 434974 471134 471618
rect 470514 434738 470546 434974
rect 470782 434738 470866 434974
rect 471102 434738 471134 434974
rect 470514 434654 471134 434738
rect 470514 434418 470546 434654
rect 470782 434418 470866 434654
rect 471102 434418 471134 434654
rect 470514 397774 471134 434418
rect 470514 397538 470546 397774
rect 470782 397538 470866 397774
rect 471102 397538 471134 397774
rect 470514 397454 471134 397538
rect 470514 397218 470546 397454
rect 470782 397218 470866 397454
rect 471102 397218 471134 397454
rect 470514 360574 471134 397218
rect 470514 360338 470546 360574
rect 470782 360338 470866 360574
rect 471102 360338 471134 360574
rect 470514 360254 471134 360338
rect 470514 360018 470546 360254
rect 470782 360018 470866 360254
rect 471102 360018 471134 360254
rect 470514 323374 471134 360018
rect 470514 323138 470546 323374
rect 470782 323138 470866 323374
rect 471102 323138 471134 323374
rect 470514 323054 471134 323138
rect 470514 322818 470546 323054
rect 470782 322818 470866 323054
rect 471102 322818 471134 323054
rect 470514 286174 471134 322818
rect 470514 285938 470546 286174
rect 470782 285938 470866 286174
rect 471102 285938 471134 286174
rect 470514 285854 471134 285938
rect 470514 285618 470546 285854
rect 470782 285618 470866 285854
rect 471102 285618 471134 285854
rect 470514 248974 471134 285618
rect 470514 248738 470546 248974
rect 470782 248738 470866 248974
rect 471102 248738 471134 248974
rect 470514 248654 471134 248738
rect 470514 248418 470546 248654
rect 470782 248418 470866 248654
rect 471102 248418 471134 248654
rect 470514 211774 471134 248418
rect 470514 211538 470546 211774
rect 470782 211538 470866 211774
rect 471102 211538 471134 211774
rect 470514 211454 471134 211538
rect 470514 211218 470546 211454
rect 470782 211218 470866 211454
rect 471102 211218 471134 211454
rect 470514 174574 471134 211218
rect 470514 174338 470546 174574
rect 470782 174338 470866 174574
rect 471102 174338 471134 174574
rect 470514 174254 471134 174338
rect 470514 174018 470546 174254
rect 470782 174018 470866 174254
rect 471102 174018 471134 174254
rect 470514 137374 471134 174018
rect 470514 137138 470546 137374
rect 470782 137138 470866 137374
rect 471102 137138 471134 137374
rect 470514 137054 471134 137138
rect 470514 136818 470546 137054
rect 470782 136818 470866 137054
rect 471102 136818 471134 137054
rect 470514 100174 471134 136818
rect 470514 99938 470546 100174
rect 470782 99938 470866 100174
rect 471102 99938 471134 100174
rect 470514 99854 471134 99938
rect 470514 99618 470546 99854
rect 470782 99618 470866 99854
rect 471102 99618 471134 99854
rect 470514 62974 471134 99618
rect 470514 62738 470546 62974
rect 470782 62738 470866 62974
rect 471102 62738 471134 62974
rect 470514 62654 471134 62738
rect 470514 62418 470546 62654
rect 470782 62418 470866 62654
rect 471102 62418 471134 62654
rect 470514 25774 471134 62418
rect 470514 25538 470546 25774
rect 470782 25538 470866 25774
rect 471102 25538 471134 25774
rect 470514 25454 471134 25538
rect 470514 25218 470546 25454
rect 470782 25218 470866 25454
rect 471102 25218 471134 25454
rect 470514 2176 471134 25218
rect 474234 699094 474854 701760
rect 474234 698858 474266 699094
rect 474502 698858 474586 699094
rect 474822 698858 474854 699094
rect 474234 698774 474854 698858
rect 474234 698538 474266 698774
rect 474502 698538 474586 698774
rect 474822 698538 474854 698774
rect 474234 661894 474854 698538
rect 474234 661658 474266 661894
rect 474502 661658 474586 661894
rect 474822 661658 474854 661894
rect 474234 661574 474854 661658
rect 474234 661338 474266 661574
rect 474502 661338 474586 661574
rect 474822 661338 474854 661574
rect 474234 624694 474854 661338
rect 474234 624458 474266 624694
rect 474502 624458 474586 624694
rect 474822 624458 474854 624694
rect 474234 624374 474854 624458
rect 474234 624138 474266 624374
rect 474502 624138 474586 624374
rect 474822 624138 474854 624374
rect 474234 587494 474854 624138
rect 474234 587258 474266 587494
rect 474502 587258 474586 587494
rect 474822 587258 474854 587494
rect 474234 587174 474854 587258
rect 474234 586938 474266 587174
rect 474502 586938 474586 587174
rect 474822 586938 474854 587174
rect 474234 550294 474854 586938
rect 474234 550058 474266 550294
rect 474502 550058 474586 550294
rect 474822 550058 474854 550294
rect 474234 549974 474854 550058
rect 474234 549738 474266 549974
rect 474502 549738 474586 549974
rect 474822 549738 474854 549974
rect 474234 513094 474854 549738
rect 474234 512858 474266 513094
rect 474502 512858 474586 513094
rect 474822 512858 474854 513094
rect 474234 512774 474854 512858
rect 474234 512538 474266 512774
rect 474502 512538 474586 512774
rect 474822 512538 474854 512774
rect 474234 475894 474854 512538
rect 474234 475658 474266 475894
rect 474502 475658 474586 475894
rect 474822 475658 474854 475894
rect 474234 475574 474854 475658
rect 474234 475338 474266 475574
rect 474502 475338 474586 475574
rect 474822 475338 474854 475574
rect 474234 438694 474854 475338
rect 474234 438458 474266 438694
rect 474502 438458 474586 438694
rect 474822 438458 474854 438694
rect 474234 438374 474854 438458
rect 474234 438138 474266 438374
rect 474502 438138 474586 438374
rect 474822 438138 474854 438374
rect 474234 401494 474854 438138
rect 474234 401258 474266 401494
rect 474502 401258 474586 401494
rect 474822 401258 474854 401494
rect 474234 401174 474854 401258
rect 474234 400938 474266 401174
rect 474502 400938 474586 401174
rect 474822 400938 474854 401174
rect 474234 364294 474854 400938
rect 474234 364058 474266 364294
rect 474502 364058 474586 364294
rect 474822 364058 474854 364294
rect 474234 363974 474854 364058
rect 474234 363738 474266 363974
rect 474502 363738 474586 363974
rect 474822 363738 474854 363974
rect 474234 327094 474854 363738
rect 485394 673054 486014 701760
rect 485394 672818 485426 673054
rect 485662 672818 485746 673054
rect 485982 672818 486014 673054
rect 485394 672734 486014 672818
rect 485394 672498 485426 672734
rect 485662 672498 485746 672734
rect 485982 672498 486014 672734
rect 485394 635854 486014 672498
rect 485394 635618 485426 635854
rect 485662 635618 485746 635854
rect 485982 635618 486014 635854
rect 485394 635534 486014 635618
rect 485394 635298 485426 635534
rect 485662 635298 485746 635534
rect 485982 635298 486014 635534
rect 485394 598654 486014 635298
rect 485394 598418 485426 598654
rect 485662 598418 485746 598654
rect 485982 598418 486014 598654
rect 485394 598334 486014 598418
rect 485394 598098 485426 598334
rect 485662 598098 485746 598334
rect 485982 598098 486014 598334
rect 485394 561454 486014 598098
rect 485394 561218 485426 561454
rect 485662 561218 485746 561454
rect 485982 561218 486014 561454
rect 485394 561134 486014 561218
rect 485394 560898 485426 561134
rect 485662 560898 485746 561134
rect 485982 560898 486014 561134
rect 485394 524254 486014 560898
rect 485394 524018 485426 524254
rect 485662 524018 485746 524254
rect 485982 524018 486014 524254
rect 485394 523934 486014 524018
rect 485394 523698 485426 523934
rect 485662 523698 485746 523934
rect 485982 523698 486014 523934
rect 485394 487054 486014 523698
rect 485394 486818 485426 487054
rect 485662 486818 485746 487054
rect 485982 486818 486014 487054
rect 485394 486734 486014 486818
rect 485394 486498 485426 486734
rect 485662 486498 485746 486734
rect 485982 486498 486014 486734
rect 485394 449854 486014 486498
rect 485394 449618 485426 449854
rect 485662 449618 485746 449854
rect 485982 449618 486014 449854
rect 485394 449534 486014 449618
rect 485394 449298 485426 449534
rect 485662 449298 485746 449534
rect 485982 449298 486014 449534
rect 485394 412654 486014 449298
rect 485394 412418 485426 412654
rect 485662 412418 485746 412654
rect 485982 412418 486014 412654
rect 485394 412334 486014 412418
rect 485394 412098 485426 412334
rect 485662 412098 485746 412334
rect 485982 412098 486014 412334
rect 485394 375454 486014 412098
rect 485394 375218 485426 375454
rect 485662 375218 485746 375454
rect 485982 375218 486014 375454
rect 485394 375134 486014 375218
rect 485394 374898 485426 375134
rect 485662 374898 485746 375134
rect 485982 374898 486014 375134
rect 485394 341772 486014 374898
rect 489114 676774 489734 701760
rect 489114 676538 489146 676774
rect 489382 676538 489466 676774
rect 489702 676538 489734 676774
rect 489114 676454 489734 676538
rect 489114 676218 489146 676454
rect 489382 676218 489466 676454
rect 489702 676218 489734 676454
rect 489114 639574 489734 676218
rect 489114 639338 489146 639574
rect 489382 639338 489466 639574
rect 489702 639338 489734 639574
rect 489114 639254 489734 639338
rect 489114 639018 489146 639254
rect 489382 639018 489466 639254
rect 489702 639018 489734 639254
rect 489114 602374 489734 639018
rect 489114 602138 489146 602374
rect 489382 602138 489466 602374
rect 489702 602138 489734 602374
rect 489114 602054 489734 602138
rect 489114 601818 489146 602054
rect 489382 601818 489466 602054
rect 489702 601818 489734 602054
rect 489114 565174 489734 601818
rect 489114 564938 489146 565174
rect 489382 564938 489466 565174
rect 489702 564938 489734 565174
rect 489114 564854 489734 564938
rect 489114 564618 489146 564854
rect 489382 564618 489466 564854
rect 489702 564618 489734 564854
rect 489114 527974 489734 564618
rect 489114 527738 489146 527974
rect 489382 527738 489466 527974
rect 489702 527738 489734 527974
rect 489114 527654 489734 527738
rect 489114 527418 489146 527654
rect 489382 527418 489466 527654
rect 489702 527418 489734 527654
rect 489114 490774 489734 527418
rect 489114 490538 489146 490774
rect 489382 490538 489466 490774
rect 489702 490538 489734 490774
rect 489114 490454 489734 490538
rect 489114 490218 489146 490454
rect 489382 490218 489466 490454
rect 489702 490218 489734 490454
rect 489114 453574 489734 490218
rect 489114 453338 489146 453574
rect 489382 453338 489466 453574
rect 489702 453338 489734 453574
rect 489114 453254 489734 453338
rect 489114 453018 489146 453254
rect 489382 453018 489466 453254
rect 489702 453018 489734 453254
rect 489114 416374 489734 453018
rect 489114 416138 489146 416374
rect 489382 416138 489466 416374
rect 489702 416138 489734 416374
rect 489114 416054 489734 416138
rect 489114 415818 489146 416054
rect 489382 415818 489466 416054
rect 489702 415818 489734 416054
rect 489114 379174 489734 415818
rect 489114 378938 489146 379174
rect 489382 378938 489466 379174
rect 489702 378938 489734 379174
rect 489114 378854 489734 378938
rect 489114 378618 489146 378854
rect 489382 378618 489466 378854
rect 489702 378618 489734 378854
rect 489114 341974 489734 378618
rect 489114 341738 489146 341974
rect 489382 341738 489466 341974
rect 489702 341738 489734 341974
rect 489114 341654 489734 341738
rect 489114 341418 489146 341654
rect 489382 341418 489466 341654
rect 489702 341418 489734 341654
rect 489114 341386 489734 341418
rect 492834 680494 493454 701760
rect 492834 680258 492866 680494
rect 493102 680258 493186 680494
rect 493422 680258 493454 680494
rect 492834 680174 493454 680258
rect 492834 679938 492866 680174
rect 493102 679938 493186 680174
rect 493422 679938 493454 680174
rect 492834 643294 493454 679938
rect 492834 643058 492866 643294
rect 493102 643058 493186 643294
rect 493422 643058 493454 643294
rect 492834 642974 493454 643058
rect 492834 642738 492866 642974
rect 493102 642738 493186 642974
rect 493422 642738 493454 642974
rect 492834 606094 493454 642738
rect 492834 605858 492866 606094
rect 493102 605858 493186 606094
rect 493422 605858 493454 606094
rect 492834 605774 493454 605858
rect 492834 605538 492866 605774
rect 493102 605538 493186 605774
rect 493422 605538 493454 605774
rect 492834 568894 493454 605538
rect 492834 568658 492866 568894
rect 493102 568658 493186 568894
rect 493422 568658 493454 568894
rect 492834 568574 493454 568658
rect 492834 568338 492866 568574
rect 493102 568338 493186 568574
rect 493422 568338 493454 568574
rect 492834 531694 493454 568338
rect 492834 531458 492866 531694
rect 493102 531458 493186 531694
rect 493422 531458 493454 531694
rect 492834 531374 493454 531458
rect 492834 531138 492866 531374
rect 493102 531138 493186 531374
rect 493422 531138 493454 531374
rect 492834 494494 493454 531138
rect 492834 494258 492866 494494
rect 493102 494258 493186 494494
rect 493422 494258 493454 494494
rect 492834 494174 493454 494258
rect 492834 493938 492866 494174
rect 493102 493938 493186 494174
rect 493422 493938 493454 494174
rect 492834 457294 493454 493938
rect 492834 457058 492866 457294
rect 493102 457058 493186 457294
rect 493422 457058 493454 457294
rect 492834 456974 493454 457058
rect 492834 456738 492866 456974
rect 493102 456738 493186 456974
rect 493422 456738 493454 456974
rect 492834 420094 493454 456738
rect 492834 419858 492866 420094
rect 493102 419858 493186 420094
rect 493422 419858 493454 420094
rect 492834 419774 493454 419858
rect 492834 419538 492866 419774
rect 493102 419538 493186 419774
rect 493422 419538 493454 419774
rect 492834 382894 493454 419538
rect 492834 382658 492866 382894
rect 493102 382658 493186 382894
rect 493422 382658 493454 382894
rect 492834 382574 493454 382658
rect 492834 382338 492866 382574
rect 493102 382338 493186 382574
rect 493422 382338 493454 382574
rect 492834 345694 493454 382338
rect 492834 345458 492866 345694
rect 493102 345458 493186 345694
rect 493422 345458 493454 345694
rect 492834 345374 493454 345458
rect 492834 345138 492866 345374
rect 493102 345138 493186 345374
rect 493422 345138 493454 345374
rect 481910 338254 482230 338286
rect 481910 338018 481952 338254
rect 482188 338018 482230 338254
rect 481910 337934 482230 338018
rect 481910 337698 481952 337934
rect 482188 337698 482230 337934
rect 481910 337666 482230 337698
rect 483842 338254 484162 338286
rect 483842 338018 483884 338254
rect 484120 338018 484162 338254
rect 483842 337934 484162 338018
rect 483842 337698 483884 337934
rect 484120 337698 484162 337934
rect 483842 337666 484162 337698
rect 485774 338254 486094 338286
rect 485774 338018 485816 338254
rect 486052 338018 486094 338254
rect 485774 337934 486094 338018
rect 485774 337698 485816 337934
rect 486052 337698 486094 337934
rect 485774 337666 486094 337698
rect 487706 338254 488026 338286
rect 487706 338018 487748 338254
rect 487984 338018 488026 338254
rect 487706 337934 488026 338018
rect 487706 337698 487748 337934
rect 487984 337698 488026 337934
rect 487706 337666 488026 337698
rect 491891 330988 491957 330989
rect 491891 330924 491892 330988
rect 491956 330924 491957 330988
rect 491891 330923 491957 330924
rect 474234 326858 474266 327094
rect 474502 326858 474586 327094
rect 474822 326858 474854 327094
rect 474234 326774 474854 326858
rect 474234 326538 474266 326774
rect 474502 326538 474586 326774
rect 474822 326538 474854 326774
rect 474234 289894 474854 326538
rect 474234 289658 474266 289894
rect 474502 289658 474586 289894
rect 474822 289658 474854 289894
rect 474234 289574 474854 289658
rect 474234 289338 474266 289574
rect 474502 289338 474586 289574
rect 474822 289338 474854 289574
rect 474234 252694 474854 289338
rect 474234 252458 474266 252694
rect 474502 252458 474586 252694
rect 474822 252458 474854 252694
rect 474234 252374 474854 252458
rect 474234 252138 474266 252374
rect 474502 252138 474586 252374
rect 474822 252138 474854 252374
rect 474234 215494 474854 252138
rect 474234 215258 474266 215494
rect 474502 215258 474586 215494
rect 474822 215258 474854 215494
rect 474234 215174 474854 215258
rect 474234 214938 474266 215174
rect 474502 214938 474586 215174
rect 474822 214938 474854 215174
rect 474234 178294 474854 214938
rect 474234 178058 474266 178294
rect 474502 178058 474586 178294
rect 474822 178058 474854 178294
rect 474234 177974 474854 178058
rect 474234 177738 474266 177974
rect 474502 177738 474586 177974
rect 474822 177738 474854 177974
rect 474234 141094 474854 177738
rect 474234 140858 474266 141094
rect 474502 140858 474586 141094
rect 474822 140858 474854 141094
rect 474234 140774 474854 140858
rect 474234 140538 474266 140774
rect 474502 140538 474586 140774
rect 474822 140538 474854 140774
rect 474234 103894 474854 140538
rect 474234 103658 474266 103894
rect 474502 103658 474586 103894
rect 474822 103658 474854 103894
rect 474234 103574 474854 103658
rect 474234 103338 474266 103574
rect 474502 103338 474586 103574
rect 474822 103338 474854 103574
rect 474234 66694 474854 103338
rect 474234 66458 474266 66694
rect 474502 66458 474586 66694
rect 474822 66458 474854 66694
rect 474234 66374 474854 66458
rect 474234 66138 474266 66374
rect 474502 66138 474586 66374
rect 474822 66138 474854 66374
rect 474234 29494 474854 66138
rect 474234 29258 474266 29494
rect 474502 29258 474586 29494
rect 474822 29258 474854 29494
rect 474234 29174 474854 29258
rect 474234 28938 474266 29174
rect 474502 28938 474586 29174
rect 474822 28938 474854 29174
rect 474234 2176 474854 28938
rect 485394 301054 486014 319988
rect 485394 300818 485426 301054
rect 485662 300818 485746 301054
rect 485982 300818 486014 301054
rect 485394 300734 486014 300818
rect 485394 300498 485426 300734
rect 485662 300498 485746 300734
rect 485982 300498 486014 300734
rect 485394 263854 486014 300498
rect 485394 263618 485426 263854
rect 485662 263618 485746 263854
rect 485982 263618 486014 263854
rect 485394 263534 486014 263618
rect 485394 263298 485426 263534
rect 485662 263298 485746 263534
rect 485982 263298 486014 263534
rect 485394 226654 486014 263298
rect 485394 226418 485426 226654
rect 485662 226418 485746 226654
rect 485982 226418 486014 226654
rect 485394 226334 486014 226418
rect 485394 226098 485426 226334
rect 485662 226098 485746 226334
rect 485982 226098 486014 226334
rect 485394 189454 486014 226098
rect 485394 189218 485426 189454
rect 485662 189218 485746 189454
rect 485982 189218 486014 189454
rect 485394 189134 486014 189218
rect 485394 188898 485426 189134
rect 485662 188898 485746 189134
rect 485982 188898 486014 189134
rect 485394 152254 486014 188898
rect 485394 152018 485426 152254
rect 485662 152018 485746 152254
rect 485982 152018 486014 152254
rect 485394 151934 486014 152018
rect 485394 151698 485426 151934
rect 485662 151698 485746 151934
rect 485982 151698 486014 151934
rect 485394 115054 486014 151698
rect 485394 114818 485426 115054
rect 485662 114818 485746 115054
rect 485982 114818 486014 115054
rect 485394 114734 486014 114818
rect 485394 114498 485426 114734
rect 485662 114498 485746 114734
rect 485982 114498 486014 114734
rect 485394 77854 486014 114498
rect 485394 77618 485426 77854
rect 485662 77618 485746 77854
rect 485982 77618 486014 77854
rect 485394 77534 486014 77618
rect 485394 77298 485426 77534
rect 485662 77298 485746 77534
rect 485982 77298 486014 77534
rect 485394 40654 486014 77298
rect 485394 40418 485426 40654
rect 485662 40418 485746 40654
rect 485982 40418 486014 40654
rect 485394 40334 486014 40418
rect 485394 40098 485426 40334
rect 485662 40098 485746 40334
rect 485982 40098 486014 40334
rect 485394 3454 486014 40098
rect 485394 3218 485426 3454
rect 485662 3218 485746 3454
rect 485982 3218 486014 3454
rect 485394 3134 486014 3218
rect 485394 2898 485426 3134
rect 485662 2898 485746 3134
rect 485982 2898 486014 3134
rect 485394 2176 486014 2898
rect 489114 304774 489734 319988
rect 489114 304538 489146 304774
rect 489382 304538 489466 304774
rect 489702 304538 489734 304774
rect 489114 304454 489734 304538
rect 489114 304218 489146 304454
rect 489382 304218 489466 304454
rect 489702 304218 489734 304454
rect 489114 267574 489734 304218
rect 489114 267338 489146 267574
rect 489382 267338 489466 267574
rect 489702 267338 489734 267574
rect 489114 267254 489734 267338
rect 489114 267018 489146 267254
rect 489382 267018 489466 267254
rect 489702 267018 489734 267254
rect 489114 230374 489734 267018
rect 489114 230138 489146 230374
rect 489382 230138 489466 230374
rect 489702 230138 489734 230374
rect 489114 230054 489734 230138
rect 489114 229818 489146 230054
rect 489382 229818 489466 230054
rect 489702 229818 489734 230054
rect 489114 193174 489734 229818
rect 489114 192938 489146 193174
rect 489382 192938 489466 193174
rect 489702 192938 489734 193174
rect 489114 192854 489734 192938
rect 489114 192618 489146 192854
rect 489382 192618 489466 192854
rect 489702 192618 489734 192854
rect 489114 155974 489734 192618
rect 489114 155738 489146 155974
rect 489382 155738 489466 155974
rect 489702 155738 489734 155974
rect 489114 155654 489734 155738
rect 489114 155418 489146 155654
rect 489382 155418 489466 155654
rect 489702 155418 489734 155654
rect 489114 118774 489734 155418
rect 489114 118538 489146 118774
rect 489382 118538 489466 118774
rect 489702 118538 489734 118774
rect 489114 118454 489734 118538
rect 489114 118218 489146 118454
rect 489382 118218 489466 118454
rect 489702 118218 489734 118454
rect 489114 81574 489734 118218
rect 489114 81338 489146 81574
rect 489382 81338 489466 81574
rect 489702 81338 489734 81574
rect 489114 81254 489734 81338
rect 489114 81018 489146 81254
rect 489382 81018 489466 81254
rect 489702 81018 489734 81254
rect 489114 44374 489734 81018
rect 489114 44138 489146 44374
rect 489382 44138 489466 44374
rect 489702 44138 489734 44374
rect 489114 44054 489734 44138
rect 489114 43818 489146 44054
rect 489382 43818 489466 44054
rect 489702 43818 489734 44054
rect 489114 7174 489734 43818
rect 491894 19821 491954 330923
rect 492834 308494 493454 345138
rect 492834 308258 492866 308494
rect 493102 308258 493186 308494
rect 493422 308258 493454 308494
rect 492834 308174 493454 308258
rect 492834 307938 492866 308174
rect 493102 307938 493186 308174
rect 493422 307938 493454 308174
rect 492834 271294 493454 307938
rect 492834 271058 492866 271294
rect 493102 271058 493186 271294
rect 493422 271058 493454 271294
rect 492834 270974 493454 271058
rect 492834 270738 492866 270974
rect 493102 270738 493186 270974
rect 493422 270738 493454 270974
rect 492834 234094 493454 270738
rect 492834 233858 492866 234094
rect 493102 233858 493186 234094
rect 493422 233858 493454 234094
rect 492834 233774 493454 233858
rect 492834 233538 492866 233774
rect 493102 233538 493186 233774
rect 493422 233538 493454 233774
rect 492834 196894 493454 233538
rect 492834 196658 492866 196894
rect 493102 196658 493186 196894
rect 493422 196658 493454 196894
rect 492834 196574 493454 196658
rect 492834 196338 492866 196574
rect 493102 196338 493186 196574
rect 493422 196338 493454 196574
rect 492834 159694 493454 196338
rect 492834 159458 492866 159694
rect 493102 159458 493186 159694
rect 493422 159458 493454 159694
rect 492834 159374 493454 159458
rect 492834 159138 492866 159374
rect 493102 159138 493186 159374
rect 493422 159138 493454 159374
rect 492834 122494 493454 159138
rect 492834 122258 492866 122494
rect 493102 122258 493186 122494
rect 493422 122258 493454 122494
rect 492834 122174 493454 122258
rect 492834 121938 492866 122174
rect 493102 121938 493186 122174
rect 493422 121938 493454 122174
rect 492834 85294 493454 121938
rect 492834 85058 492866 85294
rect 493102 85058 493186 85294
rect 493422 85058 493454 85294
rect 492834 84974 493454 85058
rect 492834 84738 492866 84974
rect 493102 84738 493186 84974
rect 493422 84738 493454 84974
rect 492834 48094 493454 84738
rect 492834 47858 492866 48094
rect 493102 47858 493186 48094
rect 493422 47858 493454 48094
rect 492834 47774 493454 47858
rect 492834 47538 492866 47774
rect 493102 47538 493186 47774
rect 493422 47538 493454 47774
rect 491891 19820 491957 19821
rect 491891 19756 491892 19820
rect 491956 19756 491957 19820
rect 491891 19755 491957 19756
rect 489114 6938 489146 7174
rect 489382 6938 489466 7174
rect 489702 6938 489734 7174
rect 489114 6854 489734 6938
rect 489114 6618 489146 6854
rect 489382 6618 489466 6854
rect 489702 6618 489734 6854
rect 489114 2176 489734 6618
rect 492834 10894 493454 47538
rect 492834 10658 492866 10894
rect 493102 10658 493186 10894
rect 493422 10658 493454 10894
rect 492834 10574 493454 10658
rect 492834 10338 492866 10574
rect 493102 10338 493186 10574
rect 493422 10338 493454 10574
rect 492834 2176 493454 10338
rect 496554 684214 497174 701760
rect 496554 683978 496586 684214
rect 496822 683978 496906 684214
rect 497142 683978 497174 684214
rect 496554 683894 497174 683978
rect 496554 683658 496586 683894
rect 496822 683658 496906 683894
rect 497142 683658 497174 683894
rect 496554 647014 497174 683658
rect 496554 646778 496586 647014
rect 496822 646778 496906 647014
rect 497142 646778 497174 647014
rect 496554 646694 497174 646778
rect 496554 646458 496586 646694
rect 496822 646458 496906 646694
rect 497142 646458 497174 646694
rect 496554 609814 497174 646458
rect 496554 609578 496586 609814
rect 496822 609578 496906 609814
rect 497142 609578 497174 609814
rect 496554 609494 497174 609578
rect 496554 609258 496586 609494
rect 496822 609258 496906 609494
rect 497142 609258 497174 609494
rect 496554 572614 497174 609258
rect 496554 572378 496586 572614
rect 496822 572378 496906 572614
rect 497142 572378 497174 572614
rect 496554 572294 497174 572378
rect 496554 572058 496586 572294
rect 496822 572058 496906 572294
rect 497142 572058 497174 572294
rect 496554 535414 497174 572058
rect 496554 535178 496586 535414
rect 496822 535178 496906 535414
rect 497142 535178 497174 535414
rect 496554 535094 497174 535178
rect 496554 534858 496586 535094
rect 496822 534858 496906 535094
rect 497142 534858 497174 535094
rect 496554 498214 497174 534858
rect 496554 497978 496586 498214
rect 496822 497978 496906 498214
rect 497142 497978 497174 498214
rect 496554 497894 497174 497978
rect 496554 497658 496586 497894
rect 496822 497658 496906 497894
rect 497142 497658 497174 497894
rect 496554 461014 497174 497658
rect 496554 460778 496586 461014
rect 496822 460778 496906 461014
rect 497142 460778 497174 461014
rect 496554 460694 497174 460778
rect 496554 460458 496586 460694
rect 496822 460458 496906 460694
rect 497142 460458 497174 460694
rect 496554 423814 497174 460458
rect 496554 423578 496586 423814
rect 496822 423578 496906 423814
rect 497142 423578 497174 423814
rect 496554 423494 497174 423578
rect 496554 423258 496586 423494
rect 496822 423258 496906 423494
rect 497142 423258 497174 423494
rect 496554 386614 497174 423258
rect 496554 386378 496586 386614
rect 496822 386378 496906 386614
rect 497142 386378 497174 386614
rect 496554 386294 497174 386378
rect 496554 386058 496586 386294
rect 496822 386058 496906 386294
rect 497142 386058 497174 386294
rect 496554 349414 497174 386058
rect 496554 349178 496586 349414
rect 496822 349178 496906 349414
rect 497142 349178 497174 349414
rect 496554 349094 497174 349178
rect 496554 348858 496586 349094
rect 496822 348858 496906 349094
rect 497142 348858 497174 349094
rect 496554 312214 497174 348858
rect 496554 311978 496586 312214
rect 496822 311978 496906 312214
rect 497142 311978 497174 312214
rect 496554 311894 497174 311978
rect 496554 311658 496586 311894
rect 496822 311658 496906 311894
rect 497142 311658 497174 311894
rect 496554 275014 497174 311658
rect 496554 274778 496586 275014
rect 496822 274778 496906 275014
rect 497142 274778 497174 275014
rect 496554 274694 497174 274778
rect 496554 274458 496586 274694
rect 496822 274458 496906 274694
rect 497142 274458 497174 274694
rect 496554 237814 497174 274458
rect 496554 237578 496586 237814
rect 496822 237578 496906 237814
rect 497142 237578 497174 237814
rect 496554 237494 497174 237578
rect 496554 237258 496586 237494
rect 496822 237258 496906 237494
rect 497142 237258 497174 237494
rect 496554 200614 497174 237258
rect 496554 200378 496586 200614
rect 496822 200378 496906 200614
rect 497142 200378 497174 200614
rect 496554 200294 497174 200378
rect 496554 200058 496586 200294
rect 496822 200058 496906 200294
rect 497142 200058 497174 200294
rect 496554 163414 497174 200058
rect 496554 163178 496586 163414
rect 496822 163178 496906 163414
rect 497142 163178 497174 163414
rect 496554 163094 497174 163178
rect 496554 162858 496586 163094
rect 496822 162858 496906 163094
rect 497142 162858 497174 163094
rect 496554 126214 497174 162858
rect 496554 125978 496586 126214
rect 496822 125978 496906 126214
rect 497142 125978 497174 126214
rect 496554 125894 497174 125978
rect 496554 125658 496586 125894
rect 496822 125658 496906 125894
rect 497142 125658 497174 125894
rect 496554 89014 497174 125658
rect 496554 88778 496586 89014
rect 496822 88778 496906 89014
rect 497142 88778 497174 89014
rect 496554 88694 497174 88778
rect 496554 88458 496586 88694
rect 496822 88458 496906 88694
rect 497142 88458 497174 88694
rect 496554 51814 497174 88458
rect 496554 51578 496586 51814
rect 496822 51578 496906 51814
rect 497142 51578 497174 51814
rect 496554 51494 497174 51578
rect 496554 51258 496586 51494
rect 496822 51258 496906 51494
rect 497142 51258 497174 51494
rect 496554 14614 497174 51258
rect 496554 14378 496586 14614
rect 496822 14378 496906 14614
rect 497142 14378 497174 14614
rect 496554 14294 497174 14378
rect 496554 14058 496586 14294
rect 496822 14058 496906 14294
rect 497142 14058 497174 14294
rect 496554 2176 497174 14058
rect 500274 687934 500894 701760
rect 500274 687698 500306 687934
rect 500542 687698 500626 687934
rect 500862 687698 500894 687934
rect 500274 687614 500894 687698
rect 500274 687378 500306 687614
rect 500542 687378 500626 687614
rect 500862 687378 500894 687614
rect 500274 650734 500894 687378
rect 500274 650498 500306 650734
rect 500542 650498 500626 650734
rect 500862 650498 500894 650734
rect 500274 650414 500894 650498
rect 500274 650178 500306 650414
rect 500542 650178 500626 650414
rect 500862 650178 500894 650414
rect 500274 613534 500894 650178
rect 500274 613298 500306 613534
rect 500542 613298 500626 613534
rect 500862 613298 500894 613534
rect 500274 613214 500894 613298
rect 500274 612978 500306 613214
rect 500542 612978 500626 613214
rect 500862 612978 500894 613214
rect 500274 576334 500894 612978
rect 500274 576098 500306 576334
rect 500542 576098 500626 576334
rect 500862 576098 500894 576334
rect 500274 576014 500894 576098
rect 500274 575778 500306 576014
rect 500542 575778 500626 576014
rect 500862 575778 500894 576014
rect 500274 539134 500894 575778
rect 500274 538898 500306 539134
rect 500542 538898 500626 539134
rect 500862 538898 500894 539134
rect 500274 538814 500894 538898
rect 500274 538578 500306 538814
rect 500542 538578 500626 538814
rect 500862 538578 500894 538814
rect 500274 501934 500894 538578
rect 500274 501698 500306 501934
rect 500542 501698 500626 501934
rect 500862 501698 500894 501934
rect 500274 501614 500894 501698
rect 500274 501378 500306 501614
rect 500542 501378 500626 501614
rect 500862 501378 500894 501614
rect 500274 464734 500894 501378
rect 500274 464498 500306 464734
rect 500542 464498 500626 464734
rect 500862 464498 500894 464734
rect 500274 464414 500894 464498
rect 500274 464178 500306 464414
rect 500542 464178 500626 464414
rect 500862 464178 500894 464414
rect 500274 427534 500894 464178
rect 500274 427298 500306 427534
rect 500542 427298 500626 427534
rect 500862 427298 500894 427534
rect 500274 427214 500894 427298
rect 500274 426978 500306 427214
rect 500542 426978 500626 427214
rect 500862 426978 500894 427214
rect 500274 390334 500894 426978
rect 500274 390098 500306 390334
rect 500542 390098 500626 390334
rect 500862 390098 500894 390334
rect 500274 390014 500894 390098
rect 500274 389778 500306 390014
rect 500542 389778 500626 390014
rect 500862 389778 500894 390014
rect 500274 353134 500894 389778
rect 500274 352898 500306 353134
rect 500542 352898 500626 353134
rect 500862 352898 500894 353134
rect 500274 352814 500894 352898
rect 500274 352578 500306 352814
rect 500542 352578 500626 352814
rect 500862 352578 500894 352814
rect 500274 315934 500894 352578
rect 500274 315698 500306 315934
rect 500542 315698 500626 315934
rect 500862 315698 500894 315934
rect 500274 315614 500894 315698
rect 500274 315378 500306 315614
rect 500542 315378 500626 315614
rect 500862 315378 500894 315614
rect 500274 278734 500894 315378
rect 500274 278498 500306 278734
rect 500542 278498 500626 278734
rect 500862 278498 500894 278734
rect 500274 278414 500894 278498
rect 500274 278178 500306 278414
rect 500542 278178 500626 278414
rect 500862 278178 500894 278414
rect 500274 241534 500894 278178
rect 500274 241298 500306 241534
rect 500542 241298 500626 241534
rect 500862 241298 500894 241534
rect 500274 241214 500894 241298
rect 500274 240978 500306 241214
rect 500542 240978 500626 241214
rect 500862 240978 500894 241214
rect 500274 204334 500894 240978
rect 500274 204098 500306 204334
rect 500542 204098 500626 204334
rect 500862 204098 500894 204334
rect 500274 204014 500894 204098
rect 500274 203778 500306 204014
rect 500542 203778 500626 204014
rect 500862 203778 500894 204014
rect 500274 167134 500894 203778
rect 500274 166898 500306 167134
rect 500542 166898 500626 167134
rect 500862 166898 500894 167134
rect 500274 166814 500894 166898
rect 500274 166578 500306 166814
rect 500542 166578 500626 166814
rect 500862 166578 500894 166814
rect 500274 129934 500894 166578
rect 500274 129698 500306 129934
rect 500542 129698 500626 129934
rect 500862 129698 500894 129934
rect 500274 129614 500894 129698
rect 500274 129378 500306 129614
rect 500542 129378 500626 129614
rect 500862 129378 500894 129614
rect 500274 92734 500894 129378
rect 500274 92498 500306 92734
rect 500542 92498 500626 92734
rect 500862 92498 500894 92734
rect 500274 92414 500894 92498
rect 500274 92178 500306 92414
rect 500542 92178 500626 92414
rect 500862 92178 500894 92414
rect 500274 55534 500894 92178
rect 500274 55298 500306 55534
rect 500542 55298 500626 55534
rect 500862 55298 500894 55534
rect 500274 55214 500894 55298
rect 500274 54978 500306 55214
rect 500542 54978 500626 55214
rect 500862 54978 500894 55214
rect 500274 18334 500894 54978
rect 500274 18098 500306 18334
rect 500542 18098 500626 18334
rect 500862 18098 500894 18334
rect 500274 18014 500894 18098
rect 500274 17778 500306 18014
rect 500542 17778 500626 18014
rect 500862 17778 500894 18014
rect 500274 2176 500894 17778
rect 503994 691654 504614 701760
rect 503994 691418 504026 691654
rect 504262 691418 504346 691654
rect 504582 691418 504614 691654
rect 503994 691334 504614 691418
rect 503994 691098 504026 691334
rect 504262 691098 504346 691334
rect 504582 691098 504614 691334
rect 503994 654454 504614 691098
rect 503994 654218 504026 654454
rect 504262 654218 504346 654454
rect 504582 654218 504614 654454
rect 503994 654134 504614 654218
rect 503994 653898 504026 654134
rect 504262 653898 504346 654134
rect 504582 653898 504614 654134
rect 503994 617254 504614 653898
rect 503994 617018 504026 617254
rect 504262 617018 504346 617254
rect 504582 617018 504614 617254
rect 503994 616934 504614 617018
rect 503994 616698 504026 616934
rect 504262 616698 504346 616934
rect 504582 616698 504614 616934
rect 503994 580054 504614 616698
rect 503994 579818 504026 580054
rect 504262 579818 504346 580054
rect 504582 579818 504614 580054
rect 503994 579734 504614 579818
rect 503994 579498 504026 579734
rect 504262 579498 504346 579734
rect 504582 579498 504614 579734
rect 503994 542854 504614 579498
rect 503994 542618 504026 542854
rect 504262 542618 504346 542854
rect 504582 542618 504614 542854
rect 503994 542534 504614 542618
rect 503994 542298 504026 542534
rect 504262 542298 504346 542534
rect 504582 542298 504614 542534
rect 503994 505654 504614 542298
rect 503994 505418 504026 505654
rect 504262 505418 504346 505654
rect 504582 505418 504614 505654
rect 503994 505334 504614 505418
rect 503994 505098 504026 505334
rect 504262 505098 504346 505334
rect 504582 505098 504614 505334
rect 503994 468454 504614 505098
rect 503994 468218 504026 468454
rect 504262 468218 504346 468454
rect 504582 468218 504614 468454
rect 503994 468134 504614 468218
rect 503994 467898 504026 468134
rect 504262 467898 504346 468134
rect 504582 467898 504614 468134
rect 503994 431254 504614 467898
rect 503994 431018 504026 431254
rect 504262 431018 504346 431254
rect 504582 431018 504614 431254
rect 503994 430934 504614 431018
rect 503994 430698 504026 430934
rect 504262 430698 504346 430934
rect 504582 430698 504614 430934
rect 503994 394054 504614 430698
rect 503994 393818 504026 394054
rect 504262 393818 504346 394054
rect 504582 393818 504614 394054
rect 503994 393734 504614 393818
rect 503994 393498 504026 393734
rect 504262 393498 504346 393734
rect 504582 393498 504614 393734
rect 503994 356854 504614 393498
rect 503994 356618 504026 356854
rect 504262 356618 504346 356854
rect 504582 356618 504614 356854
rect 503994 356534 504614 356618
rect 503994 356298 504026 356534
rect 504262 356298 504346 356534
rect 504582 356298 504614 356534
rect 503994 319654 504614 356298
rect 503994 319418 504026 319654
rect 504262 319418 504346 319654
rect 504582 319418 504614 319654
rect 503994 319334 504614 319418
rect 503994 319098 504026 319334
rect 504262 319098 504346 319334
rect 504582 319098 504614 319334
rect 503994 282454 504614 319098
rect 503994 282218 504026 282454
rect 504262 282218 504346 282454
rect 504582 282218 504614 282454
rect 503994 282134 504614 282218
rect 503994 281898 504026 282134
rect 504262 281898 504346 282134
rect 504582 281898 504614 282134
rect 503994 245254 504614 281898
rect 503994 245018 504026 245254
rect 504262 245018 504346 245254
rect 504582 245018 504614 245254
rect 503994 244934 504614 245018
rect 503994 244698 504026 244934
rect 504262 244698 504346 244934
rect 504582 244698 504614 244934
rect 503994 208054 504614 244698
rect 503994 207818 504026 208054
rect 504262 207818 504346 208054
rect 504582 207818 504614 208054
rect 503994 207734 504614 207818
rect 503994 207498 504026 207734
rect 504262 207498 504346 207734
rect 504582 207498 504614 207734
rect 503994 170854 504614 207498
rect 503994 170618 504026 170854
rect 504262 170618 504346 170854
rect 504582 170618 504614 170854
rect 503994 170534 504614 170618
rect 503994 170298 504026 170534
rect 504262 170298 504346 170534
rect 504582 170298 504614 170534
rect 503994 133654 504614 170298
rect 503994 133418 504026 133654
rect 504262 133418 504346 133654
rect 504582 133418 504614 133654
rect 503994 133334 504614 133418
rect 503994 133098 504026 133334
rect 504262 133098 504346 133334
rect 504582 133098 504614 133334
rect 503994 96454 504614 133098
rect 503994 96218 504026 96454
rect 504262 96218 504346 96454
rect 504582 96218 504614 96454
rect 503994 96134 504614 96218
rect 503994 95898 504026 96134
rect 504262 95898 504346 96134
rect 504582 95898 504614 96134
rect 503994 59254 504614 95898
rect 503994 59018 504026 59254
rect 504262 59018 504346 59254
rect 504582 59018 504614 59254
rect 503994 58934 504614 59018
rect 503994 58698 504026 58934
rect 504262 58698 504346 58934
rect 504582 58698 504614 58934
rect 503994 22054 504614 58698
rect 503994 21818 504026 22054
rect 504262 21818 504346 22054
rect 504582 21818 504614 22054
rect 503994 21734 504614 21818
rect 503994 21498 504026 21734
rect 504262 21498 504346 21734
rect 504582 21498 504614 21734
rect 503994 2176 504614 21498
rect 507714 695374 508334 701760
rect 507714 695138 507746 695374
rect 507982 695138 508066 695374
rect 508302 695138 508334 695374
rect 507714 695054 508334 695138
rect 507714 694818 507746 695054
rect 507982 694818 508066 695054
rect 508302 694818 508334 695054
rect 507714 658174 508334 694818
rect 507714 657938 507746 658174
rect 507982 657938 508066 658174
rect 508302 657938 508334 658174
rect 507714 657854 508334 657938
rect 507714 657618 507746 657854
rect 507982 657618 508066 657854
rect 508302 657618 508334 657854
rect 507714 620974 508334 657618
rect 507714 620738 507746 620974
rect 507982 620738 508066 620974
rect 508302 620738 508334 620974
rect 507714 620654 508334 620738
rect 507714 620418 507746 620654
rect 507982 620418 508066 620654
rect 508302 620418 508334 620654
rect 507714 583774 508334 620418
rect 507714 583538 507746 583774
rect 507982 583538 508066 583774
rect 508302 583538 508334 583774
rect 507714 583454 508334 583538
rect 507714 583218 507746 583454
rect 507982 583218 508066 583454
rect 508302 583218 508334 583454
rect 507714 546574 508334 583218
rect 507714 546338 507746 546574
rect 507982 546338 508066 546574
rect 508302 546338 508334 546574
rect 507714 546254 508334 546338
rect 507714 546018 507746 546254
rect 507982 546018 508066 546254
rect 508302 546018 508334 546254
rect 507714 509374 508334 546018
rect 507714 509138 507746 509374
rect 507982 509138 508066 509374
rect 508302 509138 508334 509374
rect 507714 509054 508334 509138
rect 507714 508818 507746 509054
rect 507982 508818 508066 509054
rect 508302 508818 508334 509054
rect 507714 472174 508334 508818
rect 507714 471938 507746 472174
rect 507982 471938 508066 472174
rect 508302 471938 508334 472174
rect 507714 471854 508334 471938
rect 507714 471618 507746 471854
rect 507982 471618 508066 471854
rect 508302 471618 508334 471854
rect 507714 434974 508334 471618
rect 507714 434738 507746 434974
rect 507982 434738 508066 434974
rect 508302 434738 508334 434974
rect 507714 434654 508334 434738
rect 507714 434418 507746 434654
rect 507982 434418 508066 434654
rect 508302 434418 508334 434654
rect 507714 397774 508334 434418
rect 507714 397538 507746 397774
rect 507982 397538 508066 397774
rect 508302 397538 508334 397774
rect 507714 397454 508334 397538
rect 507714 397218 507746 397454
rect 507982 397218 508066 397454
rect 508302 397218 508334 397454
rect 507714 360574 508334 397218
rect 507714 360338 507746 360574
rect 507982 360338 508066 360574
rect 508302 360338 508334 360574
rect 507714 360254 508334 360338
rect 507714 360018 507746 360254
rect 507982 360018 508066 360254
rect 508302 360018 508334 360254
rect 507714 323374 508334 360018
rect 507714 323138 507746 323374
rect 507982 323138 508066 323374
rect 508302 323138 508334 323374
rect 507714 323054 508334 323138
rect 507714 322818 507746 323054
rect 507982 322818 508066 323054
rect 508302 322818 508334 323054
rect 507714 286174 508334 322818
rect 507714 285938 507746 286174
rect 507982 285938 508066 286174
rect 508302 285938 508334 286174
rect 507714 285854 508334 285938
rect 507714 285618 507746 285854
rect 507982 285618 508066 285854
rect 508302 285618 508334 285854
rect 507714 248974 508334 285618
rect 507714 248738 507746 248974
rect 507982 248738 508066 248974
rect 508302 248738 508334 248974
rect 507714 248654 508334 248738
rect 507714 248418 507746 248654
rect 507982 248418 508066 248654
rect 508302 248418 508334 248654
rect 507714 211774 508334 248418
rect 507714 211538 507746 211774
rect 507982 211538 508066 211774
rect 508302 211538 508334 211774
rect 507714 211454 508334 211538
rect 507714 211218 507746 211454
rect 507982 211218 508066 211454
rect 508302 211218 508334 211454
rect 507714 174574 508334 211218
rect 507714 174338 507746 174574
rect 507982 174338 508066 174574
rect 508302 174338 508334 174574
rect 507714 174254 508334 174338
rect 507714 174018 507746 174254
rect 507982 174018 508066 174254
rect 508302 174018 508334 174254
rect 507714 137374 508334 174018
rect 507714 137138 507746 137374
rect 507982 137138 508066 137374
rect 508302 137138 508334 137374
rect 507714 137054 508334 137138
rect 507714 136818 507746 137054
rect 507982 136818 508066 137054
rect 508302 136818 508334 137054
rect 507714 100174 508334 136818
rect 507714 99938 507746 100174
rect 507982 99938 508066 100174
rect 508302 99938 508334 100174
rect 507714 99854 508334 99938
rect 507714 99618 507746 99854
rect 507982 99618 508066 99854
rect 508302 99618 508334 99854
rect 507714 62974 508334 99618
rect 507714 62738 507746 62974
rect 507982 62738 508066 62974
rect 508302 62738 508334 62974
rect 507714 62654 508334 62738
rect 507714 62418 507746 62654
rect 507982 62418 508066 62654
rect 508302 62418 508334 62654
rect 507714 25774 508334 62418
rect 507714 25538 507746 25774
rect 507982 25538 508066 25774
rect 508302 25538 508334 25774
rect 507714 25454 508334 25538
rect 507714 25218 507746 25454
rect 507982 25218 508066 25454
rect 508302 25218 508334 25454
rect 507714 2176 508334 25218
rect 511434 699094 512054 701760
rect 511434 698858 511466 699094
rect 511702 698858 511786 699094
rect 512022 698858 512054 699094
rect 511434 698774 512054 698858
rect 511434 698538 511466 698774
rect 511702 698538 511786 698774
rect 512022 698538 512054 698774
rect 511434 661894 512054 698538
rect 511434 661658 511466 661894
rect 511702 661658 511786 661894
rect 512022 661658 512054 661894
rect 511434 661574 512054 661658
rect 511434 661338 511466 661574
rect 511702 661338 511786 661574
rect 512022 661338 512054 661574
rect 511434 624694 512054 661338
rect 511434 624458 511466 624694
rect 511702 624458 511786 624694
rect 512022 624458 512054 624694
rect 511434 624374 512054 624458
rect 511434 624138 511466 624374
rect 511702 624138 511786 624374
rect 512022 624138 512054 624374
rect 511434 587494 512054 624138
rect 511434 587258 511466 587494
rect 511702 587258 511786 587494
rect 512022 587258 512054 587494
rect 511434 587174 512054 587258
rect 511434 586938 511466 587174
rect 511702 586938 511786 587174
rect 512022 586938 512054 587174
rect 511434 550294 512054 586938
rect 511434 550058 511466 550294
rect 511702 550058 511786 550294
rect 512022 550058 512054 550294
rect 511434 549974 512054 550058
rect 511434 549738 511466 549974
rect 511702 549738 511786 549974
rect 512022 549738 512054 549974
rect 511434 513094 512054 549738
rect 511434 512858 511466 513094
rect 511702 512858 511786 513094
rect 512022 512858 512054 513094
rect 511434 512774 512054 512858
rect 511434 512538 511466 512774
rect 511702 512538 511786 512774
rect 512022 512538 512054 512774
rect 511434 475894 512054 512538
rect 511434 475658 511466 475894
rect 511702 475658 511786 475894
rect 512022 475658 512054 475894
rect 511434 475574 512054 475658
rect 511434 475338 511466 475574
rect 511702 475338 511786 475574
rect 512022 475338 512054 475574
rect 511434 438694 512054 475338
rect 511434 438458 511466 438694
rect 511702 438458 511786 438694
rect 512022 438458 512054 438694
rect 511434 438374 512054 438458
rect 511434 438138 511466 438374
rect 511702 438138 511786 438374
rect 512022 438138 512054 438374
rect 511434 401494 512054 438138
rect 511434 401258 511466 401494
rect 511702 401258 511786 401494
rect 512022 401258 512054 401494
rect 511434 401174 512054 401258
rect 511434 400938 511466 401174
rect 511702 400938 511786 401174
rect 512022 400938 512054 401174
rect 511434 364294 512054 400938
rect 511434 364058 511466 364294
rect 511702 364058 511786 364294
rect 512022 364058 512054 364294
rect 511434 363974 512054 364058
rect 511434 363738 511466 363974
rect 511702 363738 511786 363974
rect 512022 363738 512054 363974
rect 511434 327094 512054 363738
rect 511434 326858 511466 327094
rect 511702 326858 511786 327094
rect 512022 326858 512054 327094
rect 511434 326774 512054 326858
rect 511434 326538 511466 326774
rect 511702 326538 511786 326774
rect 512022 326538 512054 326774
rect 511434 289894 512054 326538
rect 511434 289658 511466 289894
rect 511702 289658 511786 289894
rect 512022 289658 512054 289894
rect 511434 289574 512054 289658
rect 511434 289338 511466 289574
rect 511702 289338 511786 289574
rect 512022 289338 512054 289574
rect 511434 252694 512054 289338
rect 511434 252458 511466 252694
rect 511702 252458 511786 252694
rect 512022 252458 512054 252694
rect 511434 252374 512054 252458
rect 511434 252138 511466 252374
rect 511702 252138 511786 252374
rect 512022 252138 512054 252374
rect 511434 215494 512054 252138
rect 511434 215258 511466 215494
rect 511702 215258 511786 215494
rect 512022 215258 512054 215494
rect 511434 215174 512054 215258
rect 511434 214938 511466 215174
rect 511702 214938 511786 215174
rect 512022 214938 512054 215174
rect 511434 178294 512054 214938
rect 511434 178058 511466 178294
rect 511702 178058 511786 178294
rect 512022 178058 512054 178294
rect 511434 177974 512054 178058
rect 511434 177738 511466 177974
rect 511702 177738 511786 177974
rect 512022 177738 512054 177974
rect 511434 141094 512054 177738
rect 511434 140858 511466 141094
rect 511702 140858 511786 141094
rect 512022 140858 512054 141094
rect 511434 140774 512054 140858
rect 511434 140538 511466 140774
rect 511702 140538 511786 140774
rect 512022 140538 512054 140774
rect 511434 103894 512054 140538
rect 511434 103658 511466 103894
rect 511702 103658 511786 103894
rect 512022 103658 512054 103894
rect 511434 103574 512054 103658
rect 511434 103338 511466 103574
rect 511702 103338 511786 103574
rect 512022 103338 512054 103574
rect 511434 66694 512054 103338
rect 511434 66458 511466 66694
rect 511702 66458 511786 66694
rect 512022 66458 512054 66694
rect 511434 66374 512054 66458
rect 511434 66138 511466 66374
rect 511702 66138 511786 66374
rect 512022 66138 512054 66374
rect 511434 29494 512054 66138
rect 511434 29258 511466 29494
rect 511702 29258 511786 29494
rect 512022 29258 512054 29494
rect 511434 29174 512054 29258
rect 511434 28938 511466 29174
rect 511702 28938 511786 29174
rect 512022 28938 512054 29174
rect 511434 2176 512054 28938
rect 522594 673054 523214 701760
rect 522594 672818 522626 673054
rect 522862 672818 522946 673054
rect 523182 672818 523214 673054
rect 522594 672734 523214 672818
rect 522594 672498 522626 672734
rect 522862 672498 522946 672734
rect 523182 672498 523214 672734
rect 522594 635854 523214 672498
rect 522594 635618 522626 635854
rect 522862 635618 522946 635854
rect 523182 635618 523214 635854
rect 522594 635534 523214 635618
rect 522594 635298 522626 635534
rect 522862 635298 522946 635534
rect 523182 635298 523214 635534
rect 522594 598654 523214 635298
rect 522594 598418 522626 598654
rect 522862 598418 522946 598654
rect 523182 598418 523214 598654
rect 522594 598334 523214 598418
rect 522594 598098 522626 598334
rect 522862 598098 522946 598334
rect 523182 598098 523214 598334
rect 522594 561454 523214 598098
rect 522594 561218 522626 561454
rect 522862 561218 522946 561454
rect 523182 561218 523214 561454
rect 522594 561134 523214 561218
rect 522594 560898 522626 561134
rect 522862 560898 522946 561134
rect 523182 560898 523214 561134
rect 522594 524254 523214 560898
rect 522594 524018 522626 524254
rect 522862 524018 522946 524254
rect 523182 524018 523214 524254
rect 522594 523934 523214 524018
rect 522594 523698 522626 523934
rect 522862 523698 522946 523934
rect 523182 523698 523214 523934
rect 522594 487054 523214 523698
rect 522594 486818 522626 487054
rect 522862 486818 522946 487054
rect 523182 486818 523214 487054
rect 522594 486734 523214 486818
rect 522594 486498 522626 486734
rect 522862 486498 522946 486734
rect 523182 486498 523214 486734
rect 522594 449854 523214 486498
rect 522594 449618 522626 449854
rect 522862 449618 522946 449854
rect 523182 449618 523214 449854
rect 522594 449534 523214 449618
rect 522594 449298 522626 449534
rect 522862 449298 522946 449534
rect 523182 449298 523214 449534
rect 522594 412654 523214 449298
rect 522594 412418 522626 412654
rect 522862 412418 522946 412654
rect 523182 412418 523214 412654
rect 522594 412334 523214 412418
rect 522594 412098 522626 412334
rect 522862 412098 522946 412334
rect 523182 412098 523214 412334
rect 522594 375454 523214 412098
rect 522594 375218 522626 375454
rect 522862 375218 522946 375454
rect 523182 375218 523214 375454
rect 522594 375134 523214 375218
rect 522594 374898 522626 375134
rect 522862 374898 522946 375134
rect 523182 374898 523214 375134
rect 522594 338254 523214 374898
rect 522594 338018 522626 338254
rect 522862 338018 522946 338254
rect 523182 338018 523214 338254
rect 522594 337934 523214 338018
rect 522594 337698 522626 337934
rect 522862 337698 522946 337934
rect 523182 337698 523214 337934
rect 522594 301054 523214 337698
rect 522594 300818 522626 301054
rect 522862 300818 522946 301054
rect 523182 300818 523214 301054
rect 522594 300734 523214 300818
rect 522594 300498 522626 300734
rect 522862 300498 522946 300734
rect 523182 300498 523214 300734
rect 522594 263854 523214 300498
rect 522594 263618 522626 263854
rect 522862 263618 522946 263854
rect 523182 263618 523214 263854
rect 522594 263534 523214 263618
rect 522594 263298 522626 263534
rect 522862 263298 522946 263534
rect 523182 263298 523214 263534
rect 522594 226654 523214 263298
rect 522594 226418 522626 226654
rect 522862 226418 522946 226654
rect 523182 226418 523214 226654
rect 522594 226334 523214 226418
rect 522594 226098 522626 226334
rect 522862 226098 522946 226334
rect 523182 226098 523214 226334
rect 522594 189454 523214 226098
rect 522594 189218 522626 189454
rect 522862 189218 522946 189454
rect 523182 189218 523214 189454
rect 522594 189134 523214 189218
rect 522594 188898 522626 189134
rect 522862 188898 522946 189134
rect 523182 188898 523214 189134
rect 522594 152254 523214 188898
rect 522594 152018 522626 152254
rect 522862 152018 522946 152254
rect 523182 152018 523214 152254
rect 522594 151934 523214 152018
rect 522594 151698 522626 151934
rect 522862 151698 522946 151934
rect 523182 151698 523214 151934
rect 522594 115054 523214 151698
rect 522594 114818 522626 115054
rect 522862 114818 522946 115054
rect 523182 114818 523214 115054
rect 522594 114734 523214 114818
rect 522594 114498 522626 114734
rect 522862 114498 522946 114734
rect 523182 114498 523214 114734
rect 522594 77854 523214 114498
rect 522594 77618 522626 77854
rect 522862 77618 522946 77854
rect 523182 77618 523214 77854
rect 522594 77534 523214 77618
rect 522594 77298 522626 77534
rect 522862 77298 522946 77534
rect 523182 77298 523214 77534
rect 522594 40654 523214 77298
rect 522594 40418 522626 40654
rect 522862 40418 522946 40654
rect 523182 40418 523214 40654
rect 522594 40334 523214 40418
rect 522594 40098 522626 40334
rect 522862 40098 522946 40334
rect 523182 40098 523214 40334
rect 522594 3454 523214 40098
rect 522594 3218 522626 3454
rect 522862 3218 522946 3454
rect 523182 3218 523214 3454
rect 522594 3134 523214 3218
rect 522594 2898 522626 3134
rect 522862 2898 522946 3134
rect 523182 2898 523214 3134
rect 522594 2176 523214 2898
rect 526314 676774 526934 701760
rect 526314 676538 526346 676774
rect 526582 676538 526666 676774
rect 526902 676538 526934 676774
rect 526314 676454 526934 676538
rect 526314 676218 526346 676454
rect 526582 676218 526666 676454
rect 526902 676218 526934 676454
rect 526314 639574 526934 676218
rect 526314 639338 526346 639574
rect 526582 639338 526666 639574
rect 526902 639338 526934 639574
rect 526314 639254 526934 639338
rect 526314 639018 526346 639254
rect 526582 639018 526666 639254
rect 526902 639018 526934 639254
rect 526314 602374 526934 639018
rect 526314 602138 526346 602374
rect 526582 602138 526666 602374
rect 526902 602138 526934 602374
rect 526314 602054 526934 602138
rect 526314 601818 526346 602054
rect 526582 601818 526666 602054
rect 526902 601818 526934 602054
rect 526314 565174 526934 601818
rect 526314 564938 526346 565174
rect 526582 564938 526666 565174
rect 526902 564938 526934 565174
rect 526314 564854 526934 564938
rect 526314 564618 526346 564854
rect 526582 564618 526666 564854
rect 526902 564618 526934 564854
rect 526314 527974 526934 564618
rect 526314 527738 526346 527974
rect 526582 527738 526666 527974
rect 526902 527738 526934 527974
rect 526314 527654 526934 527738
rect 526314 527418 526346 527654
rect 526582 527418 526666 527654
rect 526902 527418 526934 527654
rect 526314 490774 526934 527418
rect 526314 490538 526346 490774
rect 526582 490538 526666 490774
rect 526902 490538 526934 490774
rect 526314 490454 526934 490538
rect 526314 490218 526346 490454
rect 526582 490218 526666 490454
rect 526902 490218 526934 490454
rect 526314 453574 526934 490218
rect 526314 453338 526346 453574
rect 526582 453338 526666 453574
rect 526902 453338 526934 453574
rect 526314 453254 526934 453338
rect 526314 453018 526346 453254
rect 526582 453018 526666 453254
rect 526902 453018 526934 453254
rect 526314 416374 526934 453018
rect 526314 416138 526346 416374
rect 526582 416138 526666 416374
rect 526902 416138 526934 416374
rect 526314 416054 526934 416138
rect 526314 415818 526346 416054
rect 526582 415818 526666 416054
rect 526902 415818 526934 416054
rect 526314 379174 526934 415818
rect 526314 378938 526346 379174
rect 526582 378938 526666 379174
rect 526902 378938 526934 379174
rect 526314 378854 526934 378938
rect 526314 378618 526346 378854
rect 526582 378618 526666 378854
rect 526902 378618 526934 378854
rect 526314 341974 526934 378618
rect 526314 341738 526346 341974
rect 526582 341738 526666 341974
rect 526902 341738 526934 341974
rect 526314 341654 526934 341738
rect 526314 341418 526346 341654
rect 526582 341418 526666 341654
rect 526902 341418 526934 341654
rect 526314 304774 526934 341418
rect 526314 304538 526346 304774
rect 526582 304538 526666 304774
rect 526902 304538 526934 304774
rect 526314 304454 526934 304538
rect 526314 304218 526346 304454
rect 526582 304218 526666 304454
rect 526902 304218 526934 304454
rect 526314 267574 526934 304218
rect 526314 267338 526346 267574
rect 526582 267338 526666 267574
rect 526902 267338 526934 267574
rect 526314 267254 526934 267338
rect 526314 267018 526346 267254
rect 526582 267018 526666 267254
rect 526902 267018 526934 267254
rect 526314 230374 526934 267018
rect 526314 230138 526346 230374
rect 526582 230138 526666 230374
rect 526902 230138 526934 230374
rect 526314 230054 526934 230138
rect 526314 229818 526346 230054
rect 526582 229818 526666 230054
rect 526902 229818 526934 230054
rect 526314 193174 526934 229818
rect 526314 192938 526346 193174
rect 526582 192938 526666 193174
rect 526902 192938 526934 193174
rect 526314 192854 526934 192938
rect 526314 192618 526346 192854
rect 526582 192618 526666 192854
rect 526902 192618 526934 192854
rect 526314 155974 526934 192618
rect 526314 155738 526346 155974
rect 526582 155738 526666 155974
rect 526902 155738 526934 155974
rect 526314 155654 526934 155738
rect 526314 155418 526346 155654
rect 526582 155418 526666 155654
rect 526902 155418 526934 155654
rect 526314 118774 526934 155418
rect 526314 118538 526346 118774
rect 526582 118538 526666 118774
rect 526902 118538 526934 118774
rect 526314 118454 526934 118538
rect 526314 118218 526346 118454
rect 526582 118218 526666 118454
rect 526902 118218 526934 118454
rect 526314 81574 526934 118218
rect 526314 81338 526346 81574
rect 526582 81338 526666 81574
rect 526902 81338 526934 81574
rect 526314 81254 526934 81338
rect 526314 81018 526346 81254
rect 526582 81018 526666 81254
rect 526902 81018 526934 81254
rect 526314 44374 526934 81018
rect 526314 44138 526346 44374
rect 526582 44138 526666 44374
rect 526902 44138 526934 44374
rect 526314 44054 526934 44138
rect 526314 43818 526346 44054
rect 526582 43818 526666 44054
rect 526902 43818 526934 44054
rect 526314 7174 526934 43818
rect 526314 6938 526346 7174
rect 526582 6938 526666 7174
rect 526902 6938 526934 7174
rect 526314 6854 526934 6938
rect 526314 6618 526346 6854
rect 526582 6618 526666 6854
rect 526902 6618 526934 6854
rect 526314 2176 526934 6618
rect 530034 680494 530654 701760
rect 530034 680258 530066 680494
rect 530302 680258 530386 680494
rect 530622 680258 530654 680494
rect 530034 680174 530654 680258
rect 530034 679938 530066 680174
rect 530302 679938 530386 680174
rect 530622 679938 530654 680174
rect 530034 643294 530654 679938
rect 530034 643058 530066 643294
rect 530302 643058 530386 643294
rect 530622 643058 530654 643294
rect 530034 642974 530654 643058
rect 530034 642738 530066 642974
rect 530302 642738 530386 642974
rect 530622 642738 530654 642974
rect 530034 606094 530654 642738
rect 530034 605858 530066 606094
rect 530302 605858 530386 606094
rect 530622 605858 530654 606094
rect 530034 605774 530654 605858
rect 530034 605538 530066 605774
rect 530302 605538 530386 605774
rect 530622 605538 530654 605774
rect 530034 568894 530654 605538
rect 530034 568658 530066 568894
rect 530302 568658 530386 568894
rect 530622 568658 530654 568894
rect 530034 568574 530654 568658
rect 530034 568338 530066 568574
rect 530302 568338 530386 568574
rect 530622 568338 530654 568574
rect 530034 531694 530654 568338
rect 530034 531458 530066 531694
rect 530302 531458 530386 531694
rect 530622 531458 530654 531694
rect 530034 531374 530654 531458
rect 530034 531138 530066 531374
rect 530302 531138 530386 531374
rect 530622 531138 530654 531374
rect 530034 494494 530654 531138
rect 530034 494258 530066 494494
rect 530302 494258 530386 494494
rect 530622 494258 530654 494494
rect 530034 494174 530654 494258
rect 530034 493938 530066 494174
rect 530302 493938 530386 494174
rect 530622 493938 530654 494174
rect 530034 457294 530654 493938
rect 530034 457058 530066 457294
rect 530302 457058 530386 457294
rect 530622 457058 530654 457294
rect 530034 456974 530654 457058
rect 530034 456738 530066 456974
rect 530302 456738 530386 456974
rect 530622 456738 530654 456974
rect 530034 420094 530654 456738
rect 530034 419858 530066 420094
rect 530302 419858 530386 420094
rect 530622 419858 530654 420094
rect 530034 419774 530654 419858
rect 530034 419538 530066 419774
rect 530302 419538 530386 419774
rect 530622 419538 530654 419774
rect 530034 382894 530654 419538
rect 530034 382658 530066 382894
rect 530302 382658 530386 382894
rect 530622 382658 530654 382894
rect 530034 382574 530654 382658
rect 530034 382338 530066 382574
rect 530302 382338 530386 382574
rect 530622 382338 530654 382574
rect 530034 345694 530654 382338
rect 530034 345458 530066 345694
rect 530302 345458 530386 345694
rect 530622 345458 530654 345694
rect 530034 345374 530654 345458
rect 530034 345138 530066 345374
rect 530302 345138 530386 345374
rect 530622 345138 530654 345374
rect 530034 308494 530654 345138
rect 530034 308258 530066 308494
rect 530302 308258 530386 308494
rect 530622 308258 530654 308494
rect 530034 308174 530654 308258
rect 530034 307938 530066 308174
rect 530302 307938 530386 308174
rect 530622 307938 530654 308174
rect 530034 271294 530654 307938
rect 530034 271058 530066 271294
rect 530302 271058 530386 271294
rect 530622 271058 530654 271294
rect 530034 270974 530654 271058
rect 530034 270738 530066 270974
rect 530302 270738 530386 270974
rect 530622 270738 530654 270974
rect 530034 234094 530654 270738
rect 530034 233858 530066 234094
rect 530302 233858 530386 234094
rect 530622 233858 530654 234094
rect 530034 233774 530654 233858
rect 530034 233538 530066 233774
rect 530302 233538 530386 233774
rect 530622 233538 530654 233774
rect 530034 196894 530654 233538
rect 530034 196658 530066 196894
rect 530302 196658 530386 196894
rect 530622 196658 530654 196894
rect 530034 196574 530654 196658
rect 530034 196338 530066 196574
rect 530302 196338 530386 196574
rect 530622 196338 530654 196574
rect 530034 159694 530654 196338
rect 530034 159458 530066 159694
rect 530302 159458 530386 159694
rect 530622 159458 530654 159694
rect 530034 159374 530654 159458
rect 530034 159138 530066 159374
rect 530302 159138 530386 159374
rect 530622 159138 530654 159374
rect 530034 122494 530654 159138
rect 530034 122258 530066 122494
rect 530302 122258 530386 122494
rect 530622 122258 530654 122494
rect 530034 122174 530654 122258
rect 530034 121938 530066 122174
rect 530302 121938 530386 122174
rect 530622 121938 530654 122174
rect 530034 85294 530654 121938
rect 530034 85058 530066 85294
rect 530302 85058 530386 85294
rect 530622 85058 530654 85294
rect 530034 84974 530654 85058
rect 530034 84738 530066 84974
rect 530302 84738 530386 84974
rect 530622 84738 530654 84974
rect 530034 48094 530654 84738
rect 530034 47858 530066 48094
rect 530302 47858 530386 48094
rect 530622 47858 530654 48094
rect 530034 47774 530654 47858
rect 530034 47538 530066 47774
rect 530302 47538 530386 47774
rect 530622 47538 530654 47774
rect 530034 10894 530654 47538
rect 530034 10658 530066 10894
rect 530302 10658 530386 10894
rect 530622 10658 530654 10894
rect 530034 10574 530654 10658
rect 530034 10338 530066 10574
rect 530302 10338 530386 10574
rect 530622 10338 530654 10574
rect 530034 2176 530654 10338
rect 533754 684214 534374 701760
rect 533754 683978 533786 684214
rect 534022 683978 534106 684214
rect 534342 683978 534374 684214
rect 533754 683894 534374 683978
rect 533754 683658 533786 683894
rect 534022 683658 534106 683894
rect 534342 683658 534374 683894
rect 533754 647014 534374 683658
rect 533754 646778 533786 647014
rect 534022 646778 534106 647014
rect 534342 646778 534374 647014
rect 533754 646694 534374 646778
rect 533754 646458 533786 646694
rect 534022 646458 534106 646694
rect 534342 646458 534374 646694
rect 533754 609814 534374 646458
rect 533754 609578 533786 609814
rect 534022 609578 534106 609814
rect 534342 609578 534374 609814
rect 533754 609494 534374 609578
rect 533754 609258 533786 609494
rect 534022 609258 534106 609494
rect 534342 609258 534374 609494
rect 533754 572614 534374 609258
rect 533754 572378 533786 572614
rect 534022 572378 534106 572614
rect 534342 572378 534374 572614
rect 533754 572294 534374 572378
rect 533754 572058 533786 572294
rect 534022 572058 534106 572294
rect 534342 572058 534374 572294
rect 533754 535414 534374 572058
rect 533754 535178 533786 535414
rect 534022 535178 534106 535414
rect 534342 535178 534374 535414
rect 533754 535094 534374 535178
rect 533754 534858 533786 535094
rect 534022 534858 534106 535094
rect 534342 534858 534374 535094
rect 533754 498214 534374 534858
rect 533754 497978 533786 498214
rect 534022 497978 534106 498214
rect 534342 497978 534374 498214
rect 533754 497894 534374 497978
rect 533754 497658 533786 497894
rect 534022 497658 534106 497894
rect 534342 497658 534374 497894
rect 533754 461014 534374 497658
rect 533754 460778 533786 461014
rect 534022 460778 534106 461014
rect 534342 460778 534374 461014
rect 533754 460694 534374 460778
rect 533754 460458 533786 460694
rect 534022 460458 534106 460694
rect 534342 460458 534374 460694
rect 533754 423814 534374 460458
rect 533754 423578 533786 423814
rect 534022 423578 534106 423814
rect 534342 423578 534374 423814
rect 533754 423494 534374 423578
rect 533754 423258 533786 423494
rect 534022 423258 534106 423494
rect 534342 423258 534374 423494
rect 533754 386614 534374 423258
rect 533754 386378 533786 386614
rect 534022 386378 534106 386614
rect 534342 386378 534374 386614
rect 533754 386294 534374 386378
rect 533754 386058 533786 386294
rect 534022 386058 534106 386294
rect 534342 386058 534374 386294
rect 533754 349414 534374 386058
rect 533754 349178 533786 349414
rect 534022 349178 534106 349414
rect 534342 349178 534374 349414
rect 533754 349094 534374 349178
rect 533754 348858 533786 349094
rect 534022 348858 534106 349094
rect 534342 348858 534374 349094
rect 533754 312214 534374 348858
rect 533754 311978 533786 312214
rect 534022 311978 534106 312214
rect 534342 311978 534374 312214
rect 533754 311894 534374 311978
rect 533754 311658 533786 311894
rect 534022 311658 534106 311894
rect 534342 311658 534374 311894
rect 533754 275014 534374 311658
rect 533754 274778 533786 275014
rect 534022 274778 534106 275014
rect 534342 274778 534374 275014
rect 533754 274694 534374 274778
rect 533754 274458 533786 274694
rect 534022 274458 534106 274694
rect 534342 274458 534374 274694
rect 533754 237814 534374 274458
rect 533754 237578 533786 237814
rect 534022 237578 534106 237814
rect 534342 237578 534374 237814
rect 533754 237494 534374 237578
rect 533754 237258 533786 237494
rect 534022 237258 534106 237494
rect 534342 237258 534374 237494
rect 533754 200614 534374 237258
rect 533754 200378 533786 200614
rect 534022 200378 534106 200614
rect 534342 200378 534374 200614
rect 533754 200294 534374 200378
rect 533754 200058 533786 200294
rect 534022 200058 534106 200294
rect 534342 200058 534374 200294
rect 533754 163414 534374 200058
rect 533754 163178 533786 163414
rect 534022 163178 534106 163414
rect 534342 163178 534374 163414
rect 533754 163094 534374 163178
rect 533754 162858 533786 163094
rect 534022 162858 534106 163094
rect 534342 162858 534374 163094
rect 533754 126214 534374 162858
rect 533754 125978 533786 126214
rect 534022 125978 534106 126214
rect 534342 125978 534374 126214
rect 533754 125894 534374 125978
rect 533754 125658 533786 125894
rect 534022 125658 534106 125894
rect 534342 125658 534374 125894
rect 533754 89014 534374 125658
rect 533754 88778 533786 89014
rect 534022 88778 534106 89014
rect 534342 88778 534374 89014
rect 533754 88694 534374 88778
rect 533754 88458 533786 88694
rect 534022 88458 534106 88694
rect 534342 88458 534374 88694
rect 533754 51814 534374 88458
rect 533754 51578 533786 51814
rect 534022 51578 534106 51814
rect 534342 51578 534374 51814
rect 533754 51494 534374 51578
rect 533754 51258 533786 51494
rect 534022 51258 534106 51494
rect 534342 51258 534374 51494
rect 533754 14614 534374 51258
rect 533754 14378 533786 14614
rect 534022 14378 534106 14614
rect 534342 14378 534374 14614
rect 533754 14294 534374 14378
rect 533754 14058 533786 14294
rect 534022 14058 534106 14294
rect 534342 14058 534374 14294
rect 533754 2176 534374 14058
rect 537474 687934 538094 701760
rect 537474 687698 537506 687934
rect 537742 687698 537826 687934
rect 538062 687698 538094 687934
rect 537474 687614 538094 687698
rect 537474 687378 537506 687614
rect 537742 687378 537826 687614
rect 538062 687378 538094 687614
rect 537474 650734 538094 687378
rect 537474 650498 537506 650734
rect 537742 650498 537826 650734
rect 538062 650498 538094 650734
rect 537474 650414 538094 650498
rect 537474 650178 537506 650414
rect 537742 650178 537826 650414
rect 538062 650178 538094 650414
rect 537474 613534 538094 650178
rect 537474 613298 537506 613534
rect 537742 613298 537826 613534
rect 538062 613298 538094 613534
rect 537474 613214 538094 613298
rect 537474 612978 537506 613214
rect 537742 612978 537826 613214
rect 538062 612978 538094 613214
rect 537474 576334 538094 612978
rect 537474 576098 537506 576334
rect 537742 576098 537826 576334
rect 538062 576098 538094 576334
rect 537474 576014 538094 576098
rect 537474 575778 537506 576014
rect 537742 575778 537826 576014
rect 538062 575778 538094 576014
rect 537474 539134 538094 575778
rect 537474 538898 537506 539134
rect 537742 538898 537826 539134
rect 538062 538898 538094 539134
rect 537474 538814 538094 538898
rect 537474 538578 537506 538814
rect 537742 538578 537826 538814
rect 538062 538578 538094 538814
rect 537474 501934 538094 538578
rect 537474 501698 537506 501934
rect 537742 501698 537826 501934
rect 538062 501698 538094 501934
rect 537474 501614 538094 501698
rect 537474 501378 537506 501614
rect 537742 501378 537826 501614
rect 538062 501378 538094 501614
rect 537474 464734 538094 501378
rect 537474 464498 537506 464734
rect 537742 464498 537826 464734
rect 538062 464498 538094 464734
rect 537474 464414 538094 464498
rect 537474 464178 537506 464414
rect 537742 464178 537826 464414
rect 538062 464178 538094 464414
rect 537474 427534 538094 464178
rect 537474 427298 537506 427534
rect 537742 427298 537826 427534
rect 538062 427298 538094 427534
rect 537474 427214 538094 427298
rect 537474 426978 537506 427214
rect 537742 426978 537826 427214
rect 538062 426978 538094 427214
rect 537474 390334 538094 426978
rect 537474 390098 537506 390334
rect 537742 390098 537826 390334
rect 538062 390098 538094 390334
rect 537474 390014 538094 390098
rect 537474 389778 537506 390014
rect 537742 389778 537826 390014
rect 538062 389778 538094 390014
rect 537474 353134 538094 389778
rect 537474 352898 537506 353134
rect 537742 352898 537826 353134
rect 538062 352898 538094 353134
rect 537474 352814 538094 352898
rect 537474 352578 537506 352814
rect 537742 352578 537826 352814
rect 538062 352578 538094 352814
rect 537474 315934 538094 352578
rect 537474 315698 537506 315934
rect 537742 315698 537826 315934
rect 538062 315698 538094 315934
rect 537474 315614 538094 315698
rect 537474 315378 537506 315614
rect 537742 315378 537826 315614
rect 538062 315378 538094 315614
rect 537474 278734 538094 315378
rect 537474 278498 537506 278734
rect 537742 278498 537826 278734
rect 538062 278498 538094 278734
rect 537474 278414 538094 278498
rect 537474 278178 537506 278414
rect 537742 278178 537826 278414
rect 538062 278178 538094 278414
rect 537474 241534 538094 278178
rect 537474 241298 537506 241534
rect 537742 241298 537826 241534
rect 538062 241298 538094 241534
rect 537474 241214 538094 241298
rect 537474 240978 537506 241214
rect 537742 240978 537826 241214
rect 538062 240978 538094 241214
rect 537474 204334 538094 240978
rect 537474 204098 537506 204334
rect 537742 204098 537826 204334
rect 538062 204098 538094 204334
rect 537474 204014 538094 204098
rect 537474 203778 537506 204014
rect 537742 203778 537826 204014
rect 538062 203778 538094 204014
rect 537474 167134 538094 203778
rect 537474 166898 537506 167134
rect 537742 166898 537826 167134
rect 538062 166898 538094 167134
rect 537474 166814 538094 166898
rect 537474 166578 537506 166814
rect 537742 166578 537826 166814
rect 538062 166578 538094 166814
rect 537474 129934 538094 166578
rect 537474 129698 537506 129934
rect 537742 129698 537826 129934
rect 538062 129698 538094 129934
rect 537474 129614 538094 129698
rect 537474 129378 537506 129614
rect 537742 129378 537826 129614
rect 538062 129378 538094 129614
rect 537474 92734 538094 129378
rect 537474 92498 537506 92734
rect 537742 92498 537826 92734
rect 538062 92498 538094 92734
rect 537474 92414 538094 92498
rect 537474 92178 537506 92414
rect 537742 92178 537826 92414
rect 538062 92178 538094 92414
rect 537474 55534 538094 92178
rect 537474 55298 537506 55534
rect 537742 55298 537826 55534
rect 538062 55298 538094 55534
rect 537474 55214 538094 55298
rect 537474 54978 537506 55214
rect 537742 54978 537826 55214
rect 538062 54978 538094 55214
rect 537474 18334 538094 54978
rect 537474 18098 537506 18334
rect 537742 18098 537826 18334
rect 538062 18098 538094 18334
rect 537474 18014 538094 18098
rect 537474 17778 537506 18014
rect 537742 17778 537826 18014
rect 538062 17778 538094 18014
rect 537474 2176 538094 17778
rect 541194 691654 541814 701760
rect 541194 691418 541226 691654
rect 541462 691418 541546 691654
rect 541782 691418 541814 691654
rect 541194 691334 541814 691418
rect 541194 691098 541226 691334
rect 541462 691098 541546 691334
rect 541782 691098 541814 691334
rect 541194 654454 541814 691098
rect 541194 654218 541226 654454
rect 541462 654218 541546 654454
rect 541782 654218 541814 654454
rect 541194 654134 541814 654218
rect 541194 653898 541226 654134
rect 541462 653898 541546 654134
rect 541782 653898 541814 654134
rect 541194 617254 541814 653898
rect 541194 617018 541226 617254
rect 541462 617018 541546 617254
rect 541782 617018 541814 617254
rect 541194 616934 541814 617018
rect 541194 616698 541226 616934
rect 541462 616698 541546 616934
rect 541782 616698 541814 616934
rect 541194 580054 541814 616698
rect 541194 579818 541226 580054
rect 541462 579818 541546 580054
rect 541782 579818 541814 580054
rect 541194 579734 541814 579818
rect 541194 579498 541226 579734
rect 541462 579498 541546 579734
rect 541782 579498 541814 579734
rect 541194 542854 541814 579498
rect 541194 542618 541226 542854
rect 541462 542618 541546 542854
rect 541782 542618 541814 542854
rect 541194 542534 541814 542618
rect 541194 542298 541226 542534
rect 541462 542298 541546 542534
rect 541782 542298 541814 542534
rect 541194 505654 541814 542298
rect 541194 505418 541226 505654
rect 541462 505418 541546 505654
rect 541782 505418 541814 505654
rect 541194 505334 541814 505418
rect 541194 505098 541226 505334
rect 541462 505098 541546 505334
rect 541782 505098 541814 505334
rect 541194 468454 541814 505098
rect 541194 468218 541226 468454
rect 541462 468218 541546 468454
rect 541782 468218 541814 468454
rect 541194 468134 541814 468218
rect 541194 467898 541226 468134
rect 541462 467898 541546 468134
rect 541782 467898 541814 468134
rect 541194 431254 541814 467898
rect 541194 431018 541226 431254
rect 541462 431018 541546 431254
rect 541782 431018 541814 431254
rect 541194 430934 541814 431018
rect 541194 430698 541226 430934
rect 541462 430698 541546 430934
rect 541782 430698 541814 430934
rect 541194 394054 541814 430698
rect 541194 393818 541226 394054
rect 541462 393818 541546 394054
rect 541782 393818 541814 394054
rect 541194 393734 541814 393818
rect 541194 393498 541226 393734
rect 541462 393498 541546 393734
rect 541782 393498 541814 393734
rect 541194 356854 541814 393498
rect 541194 356618 541226 356854
rect 541462 356618 541546 356854
rect 541782 356618 541814 356854
rect 541194 356534 541814 356618
rect 541194 356298 541226 356534
rect 541462 356298 541546 356534
rect 541782 356298 541814 356534
rect 541194 319654 541814 356298
rect 541194 319418 541226 319654
rect 541462 319418 541546 319654
rect 541782 319418 541814 319654
rect 541194 319334 541814 319418
rect 541194 319098 541226 319334
rect 541462 319098 541546 319334
rect 541782 319098 541814 319334
rect 541194 282454 541814 319098
rect 541194 282218 541226 282454
rect 541462 282218 541546 282454
rect 541782 282218 541814 282454
rect 541194 282134 541814 282218
rect 541194 281898 541226 282134
rect 541462 281898 541546 282134
rect 541782 281898 541814 282134
rect 541194 245254 541814 281898
rect 541194 245018 541226 245254
rect 541462 245018 541546 245254
rect 541782 245018 541814 245254
rect 541194 244934 541814 245018
rect 541194 244698 541226 244934
rect 541462 244698 541546 244934
rect 541782 244698 541814 244934
rect 541194 208054 541814 244698
rect 541194 207818 541226 208054
rect 541462 207818 541546 208054
rect 541782 207818 541814 208054
rect 541194 207734 541814 207818
rect 541194 207498 541226 207734
rect 541462 207498 541546 207734
rect 541782 207498 541814 207734
rect 541194 170854 541814 207498
rect 541194 170618 541226 170854
rect 541462 170618 541546 170854
rect 541782 170618 541814 170854
rect 541194 170534 541814 170618
rect 541194 170298 541226 170534
rect 541462 170298 541546 170534
rect 541782 170298 541814 170534
rect 541194 133654 541814 170298
rect 541194 133418 541226 133654
rect 541462 133418 541546 133654
rect 541782 133418 541814 133654
rect 541194 133334 541814 133418
rect 541194 133098 541226 133334
rect 541462 133098 541546 133334
rect 541782 133098 541814 133334
rect 541194 96454 541814 133098
rect 541194 96218 541226 96454
rect 541462 96218 541546 96454
rect 541782 96218 541814 96454
rect 541194 96134 541814 96218
rect 541194 95898 541226 96134
rect 541462 95898 541546 96134
rect 541782 95898 541814 96134
rect 541194 59254 541814 95898
rect 541194 59018 541226 59254
rect 541462 59018 541546 59254
rect 541782 59018 541814 59254
rect 541194 58934 541814 59018
rect 541194 58698 541226 58934
rect 541462 58698 541546 58934
rect 541782 58698 541814 58934
rect 541194 22054 541814 58698
rect 541194 21818 541226 22054
rect 541462 21818 541546 22054
rect 541782 21818 541814 22054
rect 541194 21734 541814 21818
rect 541194 21498 541226 21734
rect 541462 21498 541546 21734
rect 541782 21498 541814 21734
rect 541194 2176 541814 21498
rect 544914 695374 545534 701760
rect 544914 695138 544946 695374
rect 545182 695138 545266 695374
rect 545502 695138 545534 695374
rect 544914 695054 545534 695138
rect 544914 694818 544946 695054
rect 545182 694818 545266 695054
rect 545502 694818 545534 695054
rect 544914 658174 545534 694818
rect 544914 657938 544946 658174
rect 545182 657938 545266 658174
rect 545502 657938 545534 658174
rect 544914 657854 545534 657938
rect 544914 657618 544946 657854
rect 545182 657618 545266 657854
rect 545502 657618 545534 657854
rect 544914 620974 545534 657618
rect 544914 620738 544946 620974
rect 545182 620738 545266 620974
rect 545502 620738 545534 620974
rect 544914 620654 545534 620738
rect 544914 620418 544946 620654
rect 545182 620418 545266 620654
rect 545502 620418 545534 620654
rect 544914 583774 545534 620418
rect 544914 583538 544946 583774
rect 545182 583538 545266 583774
rect 545502 583538 545534 583774
rect 544914 583454 545534 583538
rect 544914 583218 544946 583454
rect 545182 583218 545266 583454
rect 545502 583218 545534 583454
rect 544914 546574 545534 583218
rect 544914 546338 544946 546574
rect 545182 546338 545266 546574
rect 545502 546338 545534 546574
rect 544914 546254 545534 546338
rect 544914 546018 544946 546254
rect 545182 546018 545266 546254
rect 545502 546018 545534 546254
rect 544914 509374 545534 546018
rect 544914 509138 544946 509374
rect 545182 509138 545266 509374
rect 545502 509138 545534 509374
rect 544914 509054 545534 509138
rect 544914 508818 544946 509054
rect 545182 508818 545266 509054
rect 545502 508818 545534 509054
rect 544914 472174 545534 508818
rect 544914 471938 544946 472174
rect 545182 471938 545266 472174
rect 545502 471938 545534 472174
rect 544914 471854 545534 471938
rect 544914 471618 544946 471854
rect 545182 471618 545266 471854
rect 545502 471618 545534 471854
rect 544914 434974 545534 471618
rect 544914 434738 544946 434974
rect 545182 434738 545266 434974
rect 545502 434738 545534 434974
rect 544914 434654 545534 434738
rect 544914 434418 544946 434654
rect 545182 434418 545266 434654
rect 545502 434418 545534 434654
rect 544914 397774 545534 434418
rect 544914 397538 544946 397774
rect 545182 397538 545266 397774
rect 545502 397538 545534 397774
rect 544914 397454 545534 397538
rect 544914 397218 544946 397454
rect 545182 397218 545266 397454
rect 545502 397218 545534 397454
rect 544914 360574 545534 397218
rect 544914 360338 544946 360574
rect 545182 360338 545266 360574
rect 545502 360338 545534 360574
rect 544914 360254 545534 360338
rect 544914 360018 544946 360254
rect 545182 360018 545266 360254
rect 545502 360018 545534 360254
rect 544914 323374 545534 360018
rect 544914 323138 544946 323374
rect 545182 323138 545266 323374
rect 545502 323138 545534 323374
rect 544914 323054 545534 323138
rect 544914 322818 544946 323054
rect 545182 322818 545266 323054
rect 545502 322818 545534 323054
rect 544914 286174 545534 322818
rect 544914 285938 544946 286174
rect 545182 285938 545266 286174
rect 545502 285938 545534 286174
rect 544914 285854 545534 285938
rect 544914 285618 544946 285854
rect 545182 285618 545266 285854
rect 545502 285618 545534 285854
rect 544914 248974 545534 285618
rect 544914 248738 544946 248974
rect 545182 248738 545266 248974
rect 545502 248738 545534 248974
rect 544914 248654 545534 248738
rect 544914 248418 544946 248654
rect 545182 248418 545266 248654
rect 545502 248418 545534 248654
rect 544914 211774 545534 248418
rect 544914 211538 544946 211774
rect 545182 211538 545266 211774
rect 545502 211538 545534 211774
rect 544914 211454 545534 211538
rect 544914 211218 544946 211454
rect 545182 211218 545266 211454
rect 545502 211218 545534 211454
rect 544914 174574 545534 211218
rect 544914 174338 544946 174574
rect 545182 174338 545266 174574
rect 545502 174338 545534 174574
rect 544914 174254 545534 174338
rect 544914 174018 544946 174254
rect 545182 174018 545266 174254
rect 545502 174018 545534 174254
rect 544914 137374 545534 174018
rect 544914 137138 544946 137374
rect 545182 137138 545266 137374
rect 545502 137138 545534 137374
rect 544914 137054 545534 137138
rect 544914 136818 544946 137054
rect 545182 136818 545266 137054
rect 545502 136818 545534 137054
rect 544914 100174 545534 136818
rect 544914 99938 544946 100174
rect 545182 99938 545266 100174
rect 545502 99938 545534 100174
rect 544914 99854 545534 99938
rect 544914 99618 544946 99854
rect 545182 99618 545266 99854
rect 545502 99618 545534 99854
rect 544914 62974 545534 99618
rect 544914 62738 544946 62974
rect 545182 62738 545266 62974
rect 545502 62738 545534 62974
rect 544914 62654 545534 62738
rect 544914 62418 544946 62654
rect 545182 62418 545266 62654
rect 545502 62418 545534 62654
rect 544914 25774 545534 62418
rect 544914 25538 544946 25774
rect 545182 25538 545266 25774
rect 545502 25538 545534 25774
rect 544914 25454 545534 25538
rect 544914 25218 544946 25454
rect 545182 25218 545266 25454
rect 545502 25218 545534 25454
rect 544914 2176 545534 25218
rect 548634 699094 549254 701760
rect 548634 698858 548666 699094
rect 548902 698858 548986 699094
rect 549222 698858 549254 699094
rect 548634 698774 549254 698858
rect 548634 698538 548666 698774
rect 548902 698538 548986 698774
rect 549222 698538 549254 698774
rect 548634 661894 549254 698538
rect 548634 661658 548666 661894
rect 548902 661658 548986 661894
rect 549222 661658 549254 661894
rect 548634 661574 549254 661658
rect 548634 661338 548666 661574
rect 548902 661338 548986 661574
rect 549222 661338 549254 661574
rect 548634 624694 549254 661338
rect 548634 624458 548666 624694
rect 548902 624458 548986 624694
rect 549222 624458 549254 624694
rect 548634 624374 549254 624458
rect 548634 624138 548666 624374
rect 548902 624138 548986 624374
rect 549222 624138 549254 624374
rect 548634 587494 549254 624138
rect 548634 587258 548666 587494
rect 548902 587258 548986 587494
rect 549222 587258 549254 587494
rect 548634 587174 549254 587258
rect 548634 586938 548666 587174
rect 548902 586938 548986 587174
rect 549222 586938 549254 587174
rect 548634 550294 549254 586938
rect 548634 550058 548666 550294
rect 548902 550058 548986 550294
rect 549222 550058 549254 550294
rect 548634 549974 549254 550058
rect 548634 549738 548666 549974
rect 548902 549738 548986 549974
rect 549222 549738 549254 549974
rect 548634 513094 549254 549738
rect 548634 512858 548666 513094
rect 548902 512858 548986 513094
rect 549222 512858 549254 513094
rect 548634 512774 549254 512858
rect 548634 512538 548666 512774
rect 548902 512538 548986 512774
rect 549222 512538 549254 512774
rect 548634 475894 549254 512538
rect 548634 475658 548666 475894
rect 548902 475658 548986 475894
rect 549222 475658 549254 475894
rect 548634 475574 549254 475658
rect 548634 475338 548666 475574
rect 548902 475338 548986 475574
rect 549222 475338 549254 475574
rect 548634 438694 549254 475338
rect 548634 438458 548666 438694
rect 548902 438458 548986 438694
rect 549222 438458 549254 438694
rect 548634 438374 549254 438458
rect 548634 438138 548666 438374
rect 548902 438138 548986 438374
rect 549222 438138 549254 438374
rect 548634 401494 549254 438138
rect 548634 401258 548666 401494
rect 548902 401258 548986 401494
rect 549222 401258 549254 401494
rect 548634 401174 549254 401258
rect 548634 400938 548666 401174
rect 548902 400938 548986 401174
rect 549222 400938 549254 401174
rect 548634 364294 549254 400938
rect 548634 364058 548666 364294
rect 548902 364058 548986 364294
rect 549222 364058 549254 364294
rect 548634 363974 549254 364058
rect 548634 363738 548666 363974
rect 548902 363738 548986 363974
rect 549222 363738 549254 363974
rect 548634 327094 549254 363738
rect 548634 326858 548666 327094
rect 548902 326858 548986 327094
rect 549222 326858 549254 327094
rect 548634 326774 549254 326858
rect 548634 326538 548666 326774
rect 548902 326538 548986 326774
rect 549222 326538 549254 326774
rect 548634 289894 549254 326538
rect 548634 289658 548666 289894
rect 548902 289658 548986 289894
rect 549222 289658 549254 289894
rect 548634 289574 549254 289658
rect 548634 289338 548666 289574
rect 548902 289338 548986 289574
rect 549222 289338 549254 289574
rect 548634 252694 549254 289338
rect 548634 252458 548666 252694
rect 548902 252458 548986 252694
rect 549222 252458 549254 252694
rect 548634 252374 549254 252458
rect 548634 252138 548666 252374
rect 548902 252138 548986 252374
rect 549222 252138 549254 252374
rect 548634 215494 549254 252138
rect 548634 215258 548666 215494
rect 548902 215258 548986 215494
rect 549222 215258 549254 215494
rect 548634 215174 549254 215258
rect 548634 214938 548666 215174
rect 548902 214938 548986 215174
rect 549222 214938 549254 215174
rect 548634 178294 549254 214938
rect 548634 178058 548666 178294
rect 548902 178058 548986 178294
rect 549222 178058 549254 178294
rect 548634 177974 549254 178058
rect 548634 177738 548666 177974
rect 548902 177738 548986 177974
rect 549222 177738 549254 177974
rect 548634 141094 549254 177738
rect 548634 140858 548666 141094
rect 548902 140858 548986 141094
rect 549222 140858 549254 141094
rect 548634 140774 549254 140858
rect 548634 140538 548666 140774
rect 548902 140538 548986 140774
rect 549222 140538 549254 140774
rect 548634 103894 549254 140538
rect 548634 103658 548666 103894
rect 548902 103658 548986 103894
rect 549222 103658 549254 103894
rect 548634 103574 549254 103658
rect 548634 103338 548666 103574
rect 548902 103338 548986 103574
rect 549222 103338 549254 103574
rect 548634 66694 549254 103338
rect 548634 66458 548666 66694
rect 548902 66458 548986 66694
rect 549222 66458 549254 66694
rect 548634 66374 549254 66458
rect 548634 66138 548666 66374
rect 548902 66138 548986 66374
rect 549222 66138 549254 66374
rect 548634 29494 549254 66138
rect 548634 29258 548666 29494
rect 548902 29258 548986 29494
rect 549222 29258 549254 29494
rect 548634 29174 549254 29258
rect 548634 28938 548666 29174
rect 548902 28938 548986 29174
rect 549222 28938 549254 29174
rect 548634 2176 549254 28938
rect 559794 673054 560414 701760
rect 559794 672818 559826 673054
rect 560062 672818 560146 673054
rect 560382 672818 560414 673054
rect 559794 672734 560414 672818
rect 559794 672498 559826 672734
rect 560062 672498 560146 672734
rect 560382 672498 560414 672734
rect 559794 635854 560414 672498
rect 559794 635618 559826 635854
rect 560062 635618 560146 635854
rect 560382 635618 560414 635854
rect 559794 635534 560414 635618
rect 559794 635298 559826 635534
rect 560062 635298 560146 635534
rect 560382 635298 560414 635534
rect 559794 598654 560414 635298
rect 559794 598418 559826 598654
rect 560062 598418 560146 598654
rect 560382 598418 560414 598654
rect 559794 598334 560414 598418
rect 559794 598098 559826 598334
rect 560062 598098 560146 598334
rect 560382 598098 560414 598334
rect 559794 561454 560414 598098
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 524254 560414 560898
rect 559794 524018 559826 524254
rect 560062 524018 560146 524254
rect 560382 524018 560414 524254
rect 559794 523934 560414 524018
rect 559794 523698 559826 523934
rect 560062 523698 560146 523934
rect 560382 523698 560414 523934
rect 559794 487054 560414 523698
rect 559794 486818 559826 487054
rect 560062 486818 560146 487054
rect 560382 486818 560414 487054
rect 559794 486734 560414 486818
rect 559794 486498 559826 486734
rect 560062 486498 560146 486734
rect 560382 486498 560414 486734
rect 559794 449854 560414 486498
rect 559794 449618 559826 449854
rect 560062 449618 560146 449854
rect 560382 449618 560414 449854
rect 559794 449534 560414 449618
rect 559794 449298 559826 449534
rect 560062 449298 560146 449534
rect 560382 449298 560414 449534
rect 559794 412654 560414 449298
rect 559794 412418 559826 412654
rect 560062 412418 560146 412654
rect 560382 412418 560414 412654
rect 559794 412334 560414 412418
rect 559794 412098 559826 412334
rect 560062 412098 560146 412334
rect 560382 412098 560414 412334
rect 559794 375454 560414 412098
rect 559794 375218 559826 375454
rect 560062 375218 560146 375454
rect 560382 375218 560414 375454
rect 559794 375134 560414 375218
rect 559794 374898 559826 375134
rect 560062 374898 560146 375134
rect 560382 374898 560414 375134
rect 559794 338254 560414 374898
rect 559794 338018 559826 338254
rect 560062 338018 560146 338254
rect 560382 338018 560414 338254
rect 559794 337934 560414 338018
rect 559794 337698 559826 337934
rect 560062 337698 560146 337934
rect 560382 337698 560414 337934
rect 559794 301054 560414 337698
rect 559794 300818 559826 301054
rect 560062 300818 560146 301054
rect 560382 300818 560414 301054
rect 559794 300734 560414 300818
rect 559794 300498 559826 300734
rect 560062 300498 560146 300734
rect 560382 300498 560414 300734
rect 559794 263854 560414 300498
rect 559794 263618 559826 263854
rect 560062 263618 560146 263854
rect 560382 263618 560414 263854
rect 559794 263534 560414 263618
rect 559794 263298 559826 263534
rect 560062 263298 560146 263534
rect 560382 263298 560414 263534
rect 559794 226654 560414 263298
rect 559794 226418 559826 226654
rect 560062 226418 560146 226654
rect 560382 226418 560414 226654
rect 559794 226334 560414 226418
rect 559794 226098 559826 226334
rect 560062 226098 560146 226334
rect 560382 226098 560414 226334
rect 559794 189454 560414 226098
rect 559794 189218 559826 189454
rect 560062 189218 560146 189454
rect 560382 189218 560414 189454
rect 559794 189134 560414 189218
rect 559794 188898 559826 189134
rect 560062 188898 560146 189134
rect 560382 188898 560414 189134
rect 559794 152254 560414 188898
rect 559794 152018 559826 152254
rect 560062 152018 560146 152254
rect 560382 152018 560414 152254
rect 559794 151934 560414 152018
rect 559794 151698 559826 151934
rect 560062 151698 560146 151934
rect 560382 151698 560414 151934
rect 559794 115054 560414 151698
rect 559794 114818 559826 115054
rect 560062 114818 560146 115054
rect 560382 114818 560414 115054
rect 559794 114734 560414 114818
rect 559794 114498 559826 114734
rect 560062 114498 560146 114734
rect 560382 114498 560414 114734
rect 559794 77854 560414 114498
rect 559794 77618 559826 77854
rect 560062 77618 560146 77854
rect 560382 77618 560414 77854
rect 559794 77534 560414 77618
rect 559794 77298 559826 77534
rect 560062 77298 560146 77534
rect 560382 77298 560414 77534
rect 559794 40654 560414 77298
rect 559794 40418 559826 40654
rect 560062 40418 560146 40654
rect 560382 40418 560414 40654
rect 559794 40334 560414 40418
rect 559794 40098 559826 40334
rect 560062 40098 560146 40334
rect 560382 40098 560414 40334
rect 559794 3454 560414 40098
rect 559794 3218 559826 3454
rect 560062 3218 560146 3454
rect 560382 3218 560414 3454
rect 559794 3134 560414 3218
rect 559794 2898 559826 3134
rect 560062 2898 560146 3134
rect 560382 2898 560414 3134
rect 559794 2176 560414 2898
rect 563514 676774 564134 701760
rect 563514 676538 563546 676774
rect 563782 676538 563866 676774
rect 564102 676538 564134 676774
rect 563514 676454 564134 676538
rect 563514 676218 563546 676454
rect 563782 676218 563866 676454
rect 564102 676218 564134 676454
rect 563514 639574 564134 676218
rect 563514 639338 563546 639574
rect 563782 639338 563866 639574
rect 564102 639338 564134 639574
rect 563514 639254 564134 639338
rect 563514 639018 563546 639254
rect 563782 639018 563866 639254
rect 564102 639018 564134 639254
rect 563514 602374 564134 639018
rect 563514 602138 563546 602374
rect 563782 602138 563866 602374
rect 564102 602138 564134 602374
rect 563514 602054 564134 602138
rect 563514 601818 563546 602054
rect 563782 601818 563866 602054
rect 564102 601818 564134 602054
rect 563514 565174 564134 601818
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 527974 564134 564618
rect 563514 527738 563546 527974
rect 563782 527738 563866 527974
rect 564102 527738 564134 527974
rect 563514 527654 564134 527738
rect 563514 527418 563546 527654
rect 563782 527418 563866 527654
rect 564102 527418 564134 527654
rect 563514 490774 564134 527418
rect 563514 490538 563546 490774
rect 563782 490538 563866 490774
rect 564102 490538 564134 490774
rect 563514 490454 564134 490538
rect 563514 490218 563546 490454
rect 563782 490218 563866 490454
rect 564102 490218 564134 490454
rect 563514 453574 564134 490218
rect 563514 453338 563546 453574
rect 563782 453338 563866 453574
rect 564102 453338 564134 453574
rect 563514 453254 564134 453338
rect 563514 453018 563546 453254
rect 563782 453018 563866 453254
rect 564102 453018 564134 453254
rect 563514 416374 564134 453018
rect 563514 416138 563546 416374
rect 563782 416138 563866 416374
rect 564102 416138 564134 416374
rect 563514 416054 564134 416138
rect 563514 415818 563546 416054
rect 563782 415818 563866 416054
rect 564102 415818 564134 416054
rect 563514 379174 564134 415818
rect 563514 378938 563546 379174
rect 563782 378938 563866 379174
rect 564102 378938 564134 379174
rect 563514 378854 564134 378938
rect 563514 378618 563546 378854
rect 563782 378618 563866 378854
rect 564102 378618 564134 378854
rect 563514 341974 564134 378618
rect 563514 341738 563546 341974
rect 563782 341738 563866 341974
rect 564102 341738 564134 341974
rect 563514 341654 564134 341738
rect 563514 341418 563546 341654
rect 563782 341418 563866 341654
rect 564102 341418 564134 341654
rect 563514 304774 564134 341418
rect 563514 304538 563546 304774
rect 563782 304538 563866 304774
rect 564102 304538 564134 304774
rect 563514 304454 564134 304538
rect 563514 304218 563546 304454
rect 563782 304218 563866 304454
rect 564102 304218 564134 304454
rect 563514 267574 564134 304218
rect 563514 267338 563546 267574
rect 563782 267338 563866 267574
rect 564102 267338 564134 267574
rect 563514 267254 564134 267338
rect 563514 267018 563546 267254
rect 563782 267018 563866 267254
rect 564102 267018 564134 267254
rect 563514 230374 564134 267018
rect 563514 230138 563546 230374
rect 563782 230138 563866 230374
rect 564102 230138 564134 230374
rect 563514 230054 564134 230138
rect 563514 229818 563546 230054
rect 563782 229818 563866 230054
rect 564102 229818 564134 230054
rect 563514 193174 564134 229818
rect 563514 192938 563546 193174
rect 563782 192938 563866 193174
rect 564102 192938 564134 193174
rect 563514 192854 564134 192938
rect 563514 192618 563546 192854
rect 563782 192618 563866 192854
rect 564102 192618 564134 192854
rect 563514 155974 564134 192618
rect 563514 155738 563546 155974
rect 563782 155738 563866 155974
rect 564102 155738 564134 155974
rect 563514 155654 564134 155738
rect 563514 155418 563546 155654
rect 563782 155418 563866 155654
rect 564102 155418 564134 155654
rect 563514 118774 564134 155418
rect 563514 118538 563546 118774
rect 563782 118538 563866 118774
rect 564102 118538 564134 118774
rect 563514 118454 564134 118538
rect 563514 118218 563546 118454
rect 563782 118218 563866 118454
rect 564102 118218 564134 118454
rect 563514 81574 564134 118218
rect 563514 81338 563546 81574
rect 563782 81338 563866 81574
rect 564102 81338 564134 81574
rect 563514 81254 564134 81338
rect 563514 81018 563546 81254
rect 563782 81018 563866 81254
rect 564102 81018 564134 81254
rect 563514 44374 564134 81018
rect 563514 44138 563546 44374
rect 563782 44138 563866 44374
rect 564102 44138 564134 44374
rect 563514 44054 564134 44138
rect 563514 43818 563546 44054
rect 563782 43818 563866 44054
rect 564102 43818 564134 44054
rect 563514 7174 564134 43818
rect 563514 6938 563546 7174
rect 563782 6938 563866 7174
rect 564102 6938 564134 7174
rect 563514 6854 564134 6938
rect 563514 6618 563546 6854
rect 563782 6618 563866 6854
rect 564102 6618 564134 6854
rect 563514 2176 564134 6618
rect 567234 680494 567854 701760
rect 567234 680258 567266 680494
rect 567502 680258 567586 680494
rect 567822 680258 567854 680494
rect 567234 680174 567854 680258
rect 567234 679938 567266 680174
rect 567502 679938 567586 680174
rect 567822 679938 567854 680174
rect 567234 643294 567854 679938
rect 567234 643058 567266 643294
rect 567502 643058 567586 643294
rect 567822 643058 567854 643294
rect 567234 642974 567854 643058
rect 567234 642738 567266 642974
rect 567502 642738 567586 642974
rect 567822 642738 567854 642974
rect 567234 606094 567854 642738
rect 567234 605858 567266 606094
rect 567502 605858 567586 606094
rect 567822 605858 567854 606094
rect 567234 605774 567854 605858
rect 567234 605538 567266 605774
rect 567502 605538 567586 605774
rect 567822 605538 567854 605774
rect 567234 568894 567854 605538
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 531694 567854 568338
rect 567234 531458 567266 531694
rect 567502 531458 567586 531694
rect 567822 531458 567854 531694
rect 567234 531374 567854 531458
rect 567234 531138 567266 531374
rect 567502 531138 567586 531374
rect 567822 531138 567854 531374
rect 567234 494494 567854 531138
rect 567234 494258 567266 494494
rect 567502 494258 567586 494494
rect 567822 494258 567854 494494
rect 567234 494174 567854 494258
rect 567234 493938 567266 494174
rect 567502 493938 567586 494174
rect 567822 493938 567854 494174
rect 567234 457294 567854 493938
rect 567234 457058 567266 457294
rect 567502 457058 567586 457294
rect 567822 457058 567854 457294
rect 567234 456974 567854 457058
rect 567234 456738 567266 456974
rect 567502 456738 567586 456974
rect 567822 456738 567854 456974
rect 567234 420094 567854 456738
rect 567234 419858 567266 420094
rect 567502 419858 567586 420094
rect 567822 419858 567854 420094
rect 567234 419774 567854 419858
rect 567234 419538 567266 419774
rect 567502 419538 567586 419774
rect 567822 419538 567854 419774
rect 567234 382894 567854 419538
rect 567234 382658 567266 382894
rect 567502 382658 567586 382894
rect 567822 382658 567854 382894
rect 567234 382574 567854 382658
rect 567234 382338 567266 382574
rect 567502 382338 567586 382574
rect 567822 382338 567854 382574
rect 567234 345694 567854 382338
rect 567234 345458 567266 345694
rect 567502 345458 567586 345694
rect 567822 345458 567854 345694
rect 567234 345374 567854 345458
rect 567234 345138 567266 345374
rect 567502 345138 567586 345374
rect 567822 345138 567854 345374
rect 567234 308494 567854 345138
rect 567234 308258 567266 308494
rect 567502 308258 567586 308494
rect 567822 308258 567854 308494
rect 567234 308174 567854 308258
rect 567234 307938 567266 308174
rect 567502 307938 567586 308174
rect 567822 307938 567854 308174
rect 567234 271294 567854 307938
rect 567234 271058 567266 271294
rect 567502 271058 567586 271294
rect 567822 271058 567854 271294
rect 567234 270974 567854 271058
rect 567234 270738 567266 270974
rect 567502 270738 567586 270974
rect 567822 270738 567854 270974
rect 567234 234094 567854 270738
rect 567234 233858 567266 234094
rect 567502 233858 567586 234094
rect 567822 233858 567854 234094
rect 567234 233774 567854 233858
rect 567234 233538 567266 233774
rect 567502 233538 567586 233774
rect 567822 233538 567854 233774
rect 567234 196894 567854 233538
rect 567234 196658 567266 196894
rect 567502 196658 567586 196894
rect 567822 196658 567854 196894
rect 567234 196574 567854 196658
rect 567234 196338 567266 196574
rect 567502 196338 567586 196574
rect 567822 196338 567854 196574
rect 567234 159694 567854 196338
rect 567234 159458 567266 159694
rect 567502 159458 567586 159694
rect 567822 159458 567854 159694
rect 567234 159374 567854 159458
rect 567234 159138 567266 159374
rect 567502 159138 567586 159374
rect 567822 159138 567854 159374
rect 567234 122494 567854 159138
rect 567234 122258 567266 122494
rect 567502 122258 567586 122494
rect 567822 122258 567854 122494
rect 567234 122174 567854 122258
rect 567234 121938 567266 122174
rect 567502 121938 567586 122174
rect 567822 121938 567854 122174
rect 567234 85294 567854 121938
rect 567234 85058 567266 85294
rect 567502 85058 567586 85294
rect 567822 85058 567854 85294
rect 567234 84974 567854 85058
rect 567234 84738 567266 84974
rect 567502 84738 567586 84974
rect 567822 84738 567854 84974
rect 567234 48094 567854 84738
rect 567234 47858 567266 48094
rect 567502 47858 567586 48094
rect 567822 47858 567854 48094
rect 567234 47774 567854 47858
rect 567234 47538 567266 47774
rect 567502 47538 567586 47774
rect 567822 47538 567854 47774
rect 567234 10894 567854 47538
rect 567234 10658 567266 10894
rect 567502 10658 567586 10894
rect 567822 10658 567854 10894
rect 567234 10574 567854 10658
rect 567234 10338 567266 10574
rect 567502 10338 567586 10574
rect 567822 10338 567854 10574
rect 567234 2176 567854 10338
rect 570954 684214 571574 701760
rect 570954 683978 570986 684214
rect 571222 683978 571306 684214
rect 571542 683978 571574 684214
rect 570954 683894 571574 683978
rect 570954 683658 570986 683894
rect 571222 683658 571306 683894
rect 571542 683658 571574 683894
rect 570954 647014 571574 683658
rect 570954 646778 570986 647014
rect 571222 646778 571306 647014
rect 571542 646778 571574 647014
rect 570954 646694 571574 646778
rect 570954 646458 570986 646694
rect 571222 646458 571306 646694
rect 571542 646458 571574 646694
rect 570954 609814 571574 646458
rect 570954 609578 570986 609814
rect 571222 609578 571306 609814
rect 571542 609578 571574 609814
rect 570954 609494 571574 609578
rect 570954 609258 570986 609494
rect 571222 609258 571306 609494
rect 571542 609258 571574 609494
rect 570954 572614 571574 609258
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 535414 571574 572058
rect 570954 535178 570986 535414
rect 571222 535178 571306 535414
rect 571542 535178 571574 535414
rect 570954 535094 571574 535178
rect 570954 534858 570986 535094
rect 571222 534858 571306 535094
rect 571542 534858 571574 535094
rect 570954 498214 571574 534858
rect 570954 497978 570986 498214
rect 571222 497978 571306 498214
rect 571542 497978 571574 498214
rect 570954 497894 571574 497978
rect 570954 497658 570986 497894
rect 571222 497658 571306 497894
rect 571542 497658 571574 497894
rect 570954 461014 571574 497658
rect 570954 460778 570986 461014
rect 571222 460778 571306 461014
rect 571542 460778 571574 461014
rect 570954 460694 571574 460778
rect 570954 460458 570986 460694
rect 571222 460458 571306 460694
rect 571542 460458 571574 460694
rect 570954 423814 571574 460458
rect 570954 423578 570986 423814
rect 571222 423578 571306 423814
rect 571542 423578 571574 423814
rect 570954 423494 571574 423578
rect 570954 423258 570986 423494
rect 571222 423258 571306 423494
rect 571542 423258 571574 423494
rect 570954 386614 571574 423258
rect 570954 386378 570986 386614
rect 571222 386378 571306 386614
rect 571542 386378 571574 386614
rect 570954 386294 571574 386378
rect 570954 386058 570986 386294
rect 571222 386058 571306 386294
rect 571542 386058 571574 386294
rect 570954 349414 571574 386058
rect 570954 349178 570986 349414
rect 571222 349178 571306 349414
rect 571542 349178 571574 349414
rect 570954 349094 571574 349178
rect 570954 348858 570986 349094
rect 571222 348858 571306 349094
rect 571542 348858 571574 349094
rect 570954 312214 571574 348858
rect 570954 311978 570986 312214
rect 571222 311978 571306 312214
rect 571542 311978 571574 312214
rect 570954 311894 571574 311978
rect 570954 311658 570986 311894
rect 571222 311658 571306 311894
rect 571542 311658 571574 311894
rect 570954 275014 571574 311658
rect 570954 274778 570986 275014
rect 571222 274778 571306 275014
rect 571542 274778 571574 275014
rect 570954 274694 571574 274778
rect 570954 274458 570986 274694
rect 571222 274458 571306 274694
rect 571542 274458 571574 274694
rect 570954 237814 571574 274458
rect 570954 237578 570986 237814
rect 571222 237578 571306 237814
rect 571542 237578 571574 237814
rect 570954 237494 571574 237578
rect 570954 237258 570986 237494
rect 571222 237258 571306 237494
rect 571542 237258 571574 237494
rect 570954 200614 571574 237258
rect 570954 200378 570986 200614
rect 571222 200378 571306 200614
rect 571542 200378 571574 200614
rect 570954 200294 571574 200378
rect 570954 200058 570986 200294
rect 571222 200058 571306 200294
rect 571542 200058 571574 200294
rect 570954 163414 571574 200058
rect 570954 163178 570986 163414
rect 571222 163178 571306 163414
rect 571542 163178 571574 163414
rect 570954 163094 571574 163178
rect 570954 162858 570986 163094
rect 571222 162858 571306 163094
rect 571542 162858 571574 163094
rect 570954 126214 571574 162858
rect 570954 125978 570986 126214
rect 571222 125978 571306 126214
rect 571542 125978 571574 126214
rect 570954 125894 571574 125978
rect 570954 125658 570986 125894
rect 571222 125658 571306 125894
rect 571542 125658 571574 125894
rect 570954 89014 571574 125658
rect 570954 88778 570986 89014
rect 571222 88778 571306 89014
rect 571542 88778 571574 89014
rect 570954 88694 571574 88778
rect 570954 88458 570986 88694
rect 571222 88458 571306 88694
rect 571542 88458 571574 88694
rect 570954 51814 571574 88458
rect 570954 51578 570986 51814
rect 571222 51578 571306 51814
rect 571542 51578 571574 51814
rect 570954 51494 571574 51578
rect 570954 51258 570986 51494
rect 571222 51258 571306 51494
rect 571542 51258 571574 51494
rect 570954 14614 571574 51258
rect 570954 14378 570986 14614
rect 571222 14378 571306 14614
rect 571542 14378 571574 14614
rect 570954 14294 571574 14378
rect 570954 14058 570986 14294
rect 571222 14058 571306 14294
rect 571542 14058 571574 14294
rect 570954 2176 571574 14058
rect 574674 687934 575294 701760
rect 574674 687698 574706 687934
rect 574942 687698 575026 687934
rect 575262 687698 575294 687934
rect 574674 687614 575294 687698
rect 574674 687378 574706 687614
rect 574942 687378 575026 687614
rect 575262 687378 575294 687614
rect 574674 650734 575294 687378
rect 574674 650498 574706 650734
rect 574942 650498 575026 650734
rect 575262 650498 575294 650734
rect 574674 650414 575294 650498
rect 574674 650178 574706 650414
rect 574942 650178 575026 650414
rect 575262 650178 575294 650414
rect 574674 613534 575294 650178
rect 574674 613298 574706 613534
rect 574942 613298 575026 613534
rect 575262 613298 575294 613534
rect 574674 613214 575294 613298
rect 574674 612978 574706 613214
rect 574942 612978 575026 613214
rect 575262 612978 575294 613214
rect 574674 576334 575294 612978
rect 574674 576098 574706 576334
rect 574942 576098 575026 576334
rect 575262 576098 575294 576334
rect 574674 576014 575294 576098
rect 574674 575778 574706 576014
rect 574942 575778 575026 576014
rect 575262 575778 575294 576014
rect 574674 539134 575294 575778
rect 574674 538898 574706 539134
rect 574942 538898 575026 539134
rect 575262 538898 575294 539134
rect 574674 538814 575294 538898
rect 574674 538578 574706 538814
rect 574942 538578 575026 538814
rect 575262 538578 575294 538814
rect 574674 501934 575294 538578
rect 574674 501698 574706 501934
rect 574942 501698 575026 501934
rect 575262 501698 575294 501934
rect 574674 501614 575294 501698
rect 574674 501378 574706 501614
rect 574942 501378 575026 501614
rect 575262 501378 575294 501614
rect 574674 464734 575294 501378
rect 574674 464498 574706 464734
rect 574942 464498 575026 464734
rect 575262 464498 575294 464734
rect 574674 464414 575294 464498
rect 574674 464178 574706 464414
rect 574942 464178 575026 464414
rect 575262 464178 575294 464414
rect 574674 427534 575294 464178
rect 574674 427298 574706 427534
rect 574942 427298 575026 427534
rect 575262 427298 575294 427534
rect 574674 427214 575294 427298
rect 574674 426978 574706 427214
rect 574942 426978 575026 427214
rect 575262 426978 575294 427214
rect 574674 390334 575294 426978
rect 574674 390098 574706 390334
rect 574942 390098 575026 390334
rect 575262 390098 575294 390334
rect 574674 390014 575294 390098
rect 574674 389778 574706 390014
rect 574942 389778 575026 390014
rect 575262 389778 575294 390014
rect 574674 353134 575294 389778
rect 574674 352898 574706 353134
rect 574942 352898 575026 353134
rect 575262 352898 575294 353134
rect 574674 352814 575294 352898
rect 574674 352578 574706 352814
rect 574942 352578 575026 352814
rect 575262 352578 575294 352814
rect 574674 315934 575294 352578
rect 574674 315698 574706 315934
rect 574942 315698 575026 315934
rect 575262 315698 575294 315934
rect 574674 315614 575294 315698
rect 574674 315378 574706 315614
rect 574942 315378 575026 315614
rect 575262 315378 575294 315614
rect 574674 278734 575294 315378
rect 574674 278498 574706 278734
rect 574942 278498 575026 278734
rect 575262 278498 575294 278734
rect 574674 278414 575294 278498
rect 574674 278178 574706 278414
rect 574942 278178 575026 278414
rect 575262 278178 575294 278414
rect 574674 241534 575294 278178
rect 574674 241298 574706 241534
rect 574942 241298 575026 241534
rect 575262 241298 575294 241534
rect 574674 241214 575294 241298
rect 574674 240978 574706 241214
rect 574942 240978 575026 241214
rect 575262 240978 575294 241214
rect 574674 204334 575294 240978
rect 574674 204098 574706 204334
rect 574942 204098 575026 204334
rect 575262 204098 575294 204334
rect 574674 204014 575294 204098
rect 574674 203778 574706 204014
rect 574942 203778 575026 204014
rect 575262 203778 575294 204014
rect 574674 167134 575294 203778
rect 574674 166898 574706 167134
rect 574942 166898 575026 167134
rect 575262 166898 575294 167134
rect 574674 166814 575294 166898
rect 574674 166578 574706 166814
rect 574942 166578 575026 166814
rect 575262 166578 575294 166814
rect 574674 129934 575294 166578
rect 574674 129698 574706 129934
rect 574942 129698 575026 129934
rect 575262 129698 575294 129934
rect 574674 129614 575294 129698
rect 574674 129378 574706 129614
rect 574942 129378 575026 129614
rect 575262 129378 575294 129614
rect 574674 92734 575294 129378
rect 574674 92498 574706 92734
rect 574942 92498 575026 92734
rect 575262 92498 575294 92734
rect 574674 92414 575294 92498
rect 574674 92178 574706 92414
rect 574942 92178 575026 92414
rect 575262 92178 575294 92414
rect 574674 55534 575294 92178
rect 574674 55298 574706 55534
rect 574942 55298 575026 55534
rect 575262 55298 575294 55534
rect 574674 55214 575294 55298
rect 574674 54978 574706 55214
rect 574942 54978 575026 55214
rect 575262 54978 575294 55214
rect 574674 18334 575294 54978
rect 574674 18098 574706 18334
rect 574942 18098 575026 18334
rect 575262 18098 575294 18334
rect 574674 18014 575294 18098
rect 574674 17778 574706 18014
rect 574942 17778 575026 18014
rect 575262 17778 575294 18014
rect 574674 2176 575294 17778
rect 578394 691654 579014 701760
rect 578394 691418 578426 691654
rect 578662 691418 578746 691654
rect 578982 691418 579014 691654
rect 578394 691334 579014 691418
rect 578394 691098 578426 691334
rect 578662 691098 578746 691334
rect 578982 691098 579014 691334
rect 578394 654454 579014 691098
rect 578394 654218 578426 654454
rect 578662 654218 578746 654454
rect 578982 654218 579014 654454
rect 578394 654134 579014 654218
rect 578394 653898 578426 654134
rect 578662 653898 578746 654134
rect 578982 653898 579014 654134
rect 578394 617254 579014 653898
rect 578394 617018 578426 617254
rect 578662 617018 578746 617254
rect 578982 617018 579014 617254
rect 578394 616934 579014 617018
rect 578394 616698 578426 616934
rect 578662 616698 578746 616934
rect 578982 616698 579014 616934
rect 578394 580054 579014 616698
rect 578394 579818 578426 580054
rect 578662 579818 578746 580054
rect 578982 579818 579014 580054
rect 578394 579734 579014 579818
rect 578394 579498 578426 579734
rect 578662 579498 578746 579734
rect 578982 579498 579014 579734
rect 578394 542854 579014 579498
rect 578394 542618 578426 542854
rect 578662 542618 578746 542854
rect 578982 542618 579014 542854
rect 578394 542534 579014 542618
rect 578394 542298 578426 542534
rect 578662 542298 578746 542534
rect 578982 542298 579014 542534
rect 578394 505654 579014 542298
rect 578394 505418 578426 505654
rect 578662 505418 578746 505654
rect 578982 505418 579014 505654
rect 578394 505334 579014 505418
rect 578394 505098 578426 505334
rect 578662 505098 578746 505334
rect 578982 505098 579014 505334
rect 578394 468454 579014 505098
rect 578394 468218 578426 468454
rect 578662 468218 578746 468454
rect 578982 468218 579014 468454
rect 578394 468134 579014 468218
rect 578394 467898 578426 468134
rect 578662 467898 578746 468134
rect 578982 467898 579014 468134
rect 578394 431254 579014 467898
rect 578394 431018 578426 431254
rect 578662 431018 578746 431254
rect 578982 431018 579014 431254
rect 578394 430934 579014 431018
rect 578394 430698 578426 430934
rect 578662 430698 578746 430934
rect 578982 430698 579014 430934
rect 578394 394054 579014 430698
rect 578394 393818 578426 394054
rect 578662 393818 578746 394054
rect 578982 393818 579014 394054
rect 578394 393734 579014 393818
rect 578394 393498 578426 393734
rect 578662 393498 578746 393734
rect 578982 393498 579014 393734
rect 578394 356854 579014 393498
rect 578394 356618 578426 356854
rect 578662 356618 578746 356854
rect 578982 356618 579014 356854
rect 578394 356534 579014 356618
rect 578394 356298 578426 356534
rect 578662 356298 578746 356534
rect 578982 356298 579014 356534
rect 578394 319654 579014 356298
rect 578394 319418 578426 319654
rect 578662 319418 578746 319654
rect 578982 319418 579014 319654
rect 578394 319334 579014 319418
rect 578394 319098 578426 319334
rect 578662 319098 578746 319334
rect 578982 319098 579014 319334
rect 578394 282454 579014 319098
rect 578394 282218 578426 282454
rect 578662 282218 578746 282454
rect 578982 282218 579014 282454
rect 578394 282134 579014 282218
rect 578394 281898 578426 282134
rect 578662 281898 578746 282134
rect 578982 281898 579014 282134
rect 578394 245254 579014 281898
rect 578394 245018 578426 245254
rect 578662 245018 578746 245254
rect 578982 245018 579014 245254
rect 578394 244934 579014 245018
rect 578394 244698 578426 244934
rect 578662 244698 578746 244934
rect 578982 244698 579014 244934
rect 578394 208054 579014 244698
rect 578394 207818 578426 208054
rect 578662 207818 578746 208054
rect 578982 207818 579014 208054
rect 578394 207734 579014 207818
rect 578394 207498 578426 207734
rect 578662 207498 578746 207734
rect 578982 207498 579014 207734
rect 578394 170854 579014 207498
rect 578394 170618 578426 170854
rect 578662 170618 578746 170854
rect 578982 170618 579014 170854
rect 578394 170534 579014 170618
rect 578394 170298 578426 170534
rect 578662 170298 578746 170534
rect 578982 170298 579014 170534
rect 578394 133654 579014 170298
rect 578394 133418 578426 133654
rect 578662 133418 578746 133654
rect 578982 133418 579014 133654
rect 578394 133334 579014 133418
rect 578394 133098 578426 133334
rect 578662 133098 578746 133334
rect 578982 133098 579014 133334
rect 578394 96454 579014 133098
rect 578394 96218 578426 96454
rect 578662 96218 578746 96454
rect 578982 96218 579014 96454
rect 578394 96134 579014 96218
rect 578394 95898 578426 96134
rect 578662 95898 578746 96134
rect 578982 95898 579014 96134
rect 578394 59254 579014 95898
rect 578394 59018 578426 59254
rect 578662 59018 578746 59254
rect 578982 59018 579014 59254
rect 578394 58934 579014 59018
rect 578394 58698 578426 58934
rect 578662 58698 578746 58934
rect 578982 58698 579014 58934
rect 578394 22054 579014 58698
rect 578394 21818 578426 22054
rect 578662 21818 578746 22054
rect 578982 21818 579014 22054
rect 578394 21734 579014 21818
rect 578394 21498 578426 21734
rect 578662 21498 578746 21734
rect 578982 21498 579014 21734
rect 578394 2176 579014 21498
rect 582114 695374 582734 701760
rect 582114 695138 582146 695374
rect 582382 695138 582466 695374
rect 582702 695138 582734 695374
rect 582114 695054 582734 695138
rect 582114 694818 582146 695054
rect 582382 694818 582466 695054
rect 582702 694818 582734 695054
rect 582114 658174 582734 694818
rect 582114 657938 582146 658174
rect 582382 657938 582466 658174
rect 582702 657938 582734 658174
rect 582114 657854 582734 657938
rect 582114 657618 582146 657854
rect 582382 657618 582466 657854
rect 582702 657618 582734 657854
rect 582114 620974 582734 657618
rect 582114 620738 582146 620974
rect 582382 620738 582466 620974
rect 582702 620738 582734 620974
rect 582114 620654 582734 620738
rect 582114 620418 582146 620654
rect 582382 620418 582466 620654
rect 582702 620418 582734 620654
rect 582114 583774 582734 620418
rect 582114 583538 582146 583774
rect 582382 583538 582466 583774
rect 582702 583538 582734 583774
rect 582114 583454 582734 583538
rect 582114 583218 582146 583454
rect 582382 583218 582466 583454
rect 582702 583218 582734 583454
rect 582114 546574 582734 583218
rect 582114 546338 582146 546574
rect 582382 546338 582466 546574
rect 582702 546338 582734 546574
rect 582114 546254 582734 546338
rect 582114 546018 582146 546254
rect 582382 546018 582466 546254
rect 582702 546018 582734 546254
rect 582114 509374 582734 546018
rect 582114 509138 582146 509374
rect 582382 509138 582466 509374
rect 582702 509138 582734 509374
rect 582114 509054 582734 509138
rect 582114 508818 582146 509054
rect 582382 508818 582466 509054
rect 582702 508818 582734 509054
rect 582114 472174 582734 508818
rect 582114 471938 582146 472174
rect 582382 471938 582466 472174
rect 582702 471938 582734 472174
rect 582114 471854 582734 471938
rect 582114 471618 582146 471854
rect 582382 471618 582466 471854
rect 582702 471618 582734 471854
rect 582114 434974 582734 471618
rect 582114 434738 582146 434974
rect 582382 434738 582466 434974
rect 582702 434738 582734 434974
rect 582114 434654 582734 434738
rect 582114 434418 582146 434654
rect 582382 434418 582466 434654
rect 582702 434418 582734 434654
rect 582114 397774 582734 434418
rect 582114 397538 582146 397774
rect 582382 397538 582466 397774
rect 582702 397538 582734 397774
rect 582114 397454 582734 397538
rect 582114 397218 582146 397454
rect 582382 397218 582466 397454
rect 582702 397218 582734 397454
rect 582114 360574 582734 397218
rect 582114 360338 582146 360574
rect 582382 360338 582466 360574
rect 582702 360338 582734 360574
rect 582114 360254 582734 360338
rect 582114 360018 582146 360254
rect 582382 360018 582466 360254
rect 582702 360018 582734 360254
rect 582114 323374 582734 360018
rect 582114 323138 582146 323374
rect 582382 323138 582466 323374
rect 582702 323138 582734 323374
rect 582114 323054 582734 323138
rect 582114 322818 582146 323054
rect 582382 322818 582466 323054
rect 582702 322818 582734 323054
rect 582114 286174 582734 322818
rect 582114 285938 582146 286174
rect 582382 285938 582466 286174
rect 582702 285938 582734 286174
rect 582114 285854 582734 285938
rect 582114 285618 582146 285854
rect 582382 285618 582466 285854
rect 582702 285618 582734 285854
rect 582114 248974 582734 285618
rect 582114 248738 582146 248974
rect 582382 248738 582466 248974
rect 582702 248738 582734 248974
rect 582114 248654 582734 248738
rect 582114 248418 582146 248654
rect 582382 248418 582466 248654
rect 582702 248418 582734 248654
rect 582114 211774 582734 248418
rect 582114 211538 582146 211774
rect 582382 211538 582466 211774
rect 582702 211538 582734 211774
rect 582114 211454 582734 211538
rect 582114 211218 582146 211454
rect 582382 211218 582466 211454
rect 582702 211218 582734 211454
rect 582114 174574 582734 211218
rect 582114 174338 582146 174574
rect 582382 174338 582466 174574
rect 582702 174338 582734 174574
rect 582114 174254 582734 174338
rect 582114 174018 582146 174254
rect 582382 174018 582466 174254
rect 582702 174018 582734 174254
rect 582114 137374 582734 174018
rect 582114 137138 582146 137374
rect 582382 137138 582466 137374
rect 582702 137138 582734 137374
rect 582114 137054 582734 137138
rect 582114 136818 582146 137054
rect 582382 136818 582466 137054
rect 582702 136818 582734 137054
rect 582114 100174 582734 136818
rect 582114 99938 582146 100174
rect 582382 99938 582466 100174
rect 582702 99938 582734 100174
rect 582114 99854 582734 99938
rect 582114 99618 582146 99854
rect 582382 99618 582466 99854
rect 582702 99618 582734 99854
rect 582114 62974 582734 99618
rect 582114 62738 582146 62974
rect 582382 62738 582466 62974
rect 582702 62738 582734 62974
rect 582114 62654 582734 62738
rect 582114 62418 582146 62654
rect 582382 62418 582466 62654
rect 582702 62418 582734 62654
rect 582114 25774 582734 62418
rect 582114 25538 582146 25774
rect 582382 25538 582466 25774
rect 582702 25538 582734 25774
rect 582114 25454 582734 25538
rect 582114 25218 582146 25454
rect 582382 25218 582466 25454
rect 582702 25218 582734 25454
rect 582114 2176 582734 25218
<< via4 >>
rect 1826 672818 2062 673054
rect 2146 672818 2382 673054
rect 1826 672498 2062 672734
rect 2146 672498 2382 672734
rect 1826 635618 2062 635854
rect 2146 635618 2382 635854
rect 1826 635298 2062 635534
rect 2146 635298 2382 635534
rect 1826 598418 2062 598654
rect 2146 598418 2382 598654
rect 1826 598098 2062 598334
rect 2146 598098 2382 598334
rect 1826 561218 2062 561454
rect 2146 561218 2382 561454
rect 1826 560898 2062 561134
rect 2146 560898 2382 561134
rect 1826 524018 2062 524254
rect 2146 524018 2382 524254
rect 1826 523698 2062 523934
rect 2146 523698 2382 523934
rect 1826 486818 2062 487054
rect 2146 486818 2382 487054
rect 1826 486498 2062 486734
rect 2146 486498 2382 486734
rect 1826 449618 2062 449854
rect 2146 449618 2382 449854
rect 1826 449298 2062 449534
rect 2146 449298 2382 449534
rect 1826 412418 2062 412654
rect 2146 412418 2382 412654
rect 1826 412098 2062 412334
rect 2146 412098 2382 412334
rect 1826 375218 2062 375454
rect 2146 375218 2382 375454
rect 1826 374898 2062 375134
rect 2146 374898 2382 375134
rect 1826 338018 2062 338254
rect 2146 338018 2382 338254
rect 1826 337698 2062 337934
rect 2146 337698 2382 337934
rect 1826 300818 2062 301054
rect 2146 300818 2382 301054
rect 1826 300498 2062 300734
rect 2146 300498 2382 300734
rect 1826 263618 2062 263854
rect 2146 263618 2382 263854
rect 1826 263298 2062 263534
rect 2146 263298 2382 263534
rect 1826 226418 2062 226654
rect 2146 226418 2382 226654
rect 1826 226098 2062 226334
rect 2146 226098 2382 226334
rect 1826 189218 2062 189454
rect 2146 189218 2382 189454
rect 1826 188898 2062 189134
rect 2146 188898 2382 189134
rect 1826 152018 2062 152254
rect 2146 152018 2382 152254
rect 1826 151698 2062 151934
rect 2146 151698 2382 151934
rect 1826 114818 2062 115054
rect 2146 114818 2382 115054
rect 1826 114498 2062 114734
rect 2146 114498 2382 114734
rect 1826 77618 2062 77854
rect 2146 77618 2382 77854
rect 1826 77298 2062 77534
rect 2146 77298 2382 77534
rect 1826 40418 2062 40654
rect 2146 40418 2382 40654
rect 1826 40098 2062 40334
rect 2146 40098 2382 40334
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 5546 676538 5782 676774
rect 5866 676538 6102 676774
rect 5546 676218 5782 676454
rect 5866 676218 6102 676454
rect 5546 639338 5782 639574
rect 5866 639338 6102 639574
rect 5546 639018 5782 639254
rect 5866 639018 6102 639254
rect 5546 602138 5782 602374
rect 5866 602138 6102 602374
rect 5546 601818 5782 602054
rect 5866 601818 6102 602054
rect 5546 564938 5782 565174
rect 5866 564938 6102 565174
rect 5546 564618 5782 564854
rect 5866 564618 6102 564854
rect 5546 527738 5782 527974
rect 5866 527738 6102 527974
rect 5546 527418 5782 527654
rect 5866 527418 6102 527654
rect 5546 490538 5782 490774
rect 5866 490538 6102 490774
rect 5546 490218 5782 490454
rect 5866 490218 6102 490454
rect 5546 453338 5782 453574
rect 5866 453338 6102 453574
rect 5546 453018 5782 453254
rect 5866 453018 6102 453254
rect 5546 416138 5782 416374
rect 5866 416138 6102 416374
rect 5546 415818 5782 416054
rect 5866 415818 6102 416054
rect 5546 378938 5782 379174
rect 5866 378938 6102 379174
rect 5546 378618 5782 378854
rect 5866 378618 6102 378854
rect 5546 341738 5782 341974
rect 5866 341738 6102 341974
rect 5546 341418 5782 341654
rect 5866 341418 6102 341654
rect 5546 304538 5782 304774
rect 5866 304538 6102 304774
rect 5546 304218 5782 304454
rect 5866 304218 6102 304454
rect 5546 267338 5782 267574
rect 5866 267338 6102 267574
rect 5546 267018 5782 267254
rect 5866 267018 6102 267254
rect 5546 230138 5782 230374
rect 5866 230138 6102 230374
rect 5546 229818 5782 230054
rect 5866 229818 6102 230054
rect 5546 192938 5782 193174
rect 5866 192938 6102 193174
rect 5546 192618 5782 192854
rect 5866 192618 6102 192854
rect 5546 155738 5782 155974
rect 5866 155738 6102 155974
rect 5546 155418 5782 155654
rect 5866 155418 6102 155654
rect 5546 118538 5782 118774
rect 5866 118538 6102 118774
rect 5546 118218 5782 118454
rect 5866 118218 6102 118454
rect 5546 81338 5782 81574
rect 5866 81338 6102 81574
rect 5546 81018 5782 81254
rect 5866 81018 6102 81254
rect 5546 44138 5782 44374
rect 5866 44138 6102 44374
rect 5546 43818 5782 44054
rect 5866 43818 6102 44054
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect 9266 680258 9502 680494
rect 9586 680258 9822 680494
rect 9266 679938 9502 680174
rect 9586 679938 9822 680174
rect 9266 643058 9502 643294
rect 9586 643058 9822 643294
rect 9266 642738 9502 642974
rect 9586 642738 9822 642974
rect 9266 605858 9502 606094
rect 9586 605858 9822 606094
rect 9266 605538 9502 605774
rect 9586 605538 9822 605774
rect 9266 568658 9502 568894
rect 9586 568658 9822 568894
rect 9266 568338 9502 568574
rect 9586 568338 9822 568574
rect 9266 531458 9502 531694
rect 9586 531458 9822 531694
rect 9266 531138 9502 531374
rect 9586 531138 9822 531374
rect 9266 494258 9502 494494
rect 9586 494258 9822 494494
rect 9266 493938 9502 494174
rect 9586 493938 9822 494174
rect 9266 457058 9502 457294
rect 9586 457058 9822 457294
rect 9266 456738 9502 456974
rect 9586 456738 9822 456974
rect 9266 419858 9502 420094
rect 9586 419858 9822 420094
rect 9266 419538 9502 419774
rect 9586 419538 9822 419774
rect 9266 382658 9502 382894
rect 9586 382658 9822 382894
rect 9266 382338 9502 382574
rect 9586 382338 9822 382574
rect 9266 345458 9502 345694
rect 9586 345458 9822 345694
rect 9266 345138 9502 345374
rect 9586 345138 9822 345374
rect 9266 308258 9502 308494
rect 9586 308258 9822 308494
rect 9266 307938 9502 308174
rect 9586 307938 9822 308174
rect 9266 271058 9502 271294
rect 9586 271058 9822 271294
rect 9266 270738 9502 270974
rect 9586 270738 9822 270974
rect 9266 233858 9502 234094
rect 9586 233858 9822 234094
rect 9266 233538 9502 233774
rect 9586 233538 9822 233774
rect 9266 196658 9502 196894
rect 9586 196658 9822 196894
rect 9266 196338 9502 196574
rect 9586 196338 9822 196574
rect 9266 159458 9502 159694
rect 9586 159458 9822 159694
rect 9266 159138 9502 159374
rect 9586 159138 9822 159374
rect 9266 122258 9502 122494
rect 9586 122258 9822 122494
rect 9266 121938 9502 122174
rect 9586 121938 9822 122174
rect 9266 85058 9502 85294
rect 9586 85058 9822 85294
rect 9266 84738 9502 84974
rect 9586 84738 9822 84974
rect 9266 47858 9502 48094
rect 9586 47858 9822 48094
rect 9266 47538 9502 47774
rect 9586 47538 9822 47774
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect 12986 683978 13222 684214
rect 13306 683978 13542 684214
rect 12986 683658 13222 683894
rect 13306 683658 13542 683894
rect 12986 646778 13222 647014
rect 13306 646778 13542 647014
rect 12986 646458 13222 646694
rect 13306 646458 13542 646694
rect 12986 609578 13222 609814
rect 13306 609578 13542 609814
rect 12986 609258 13222 609494
rect 13306 609258 13542 609494
rect 12986 572378 13222 572614
rect 13306 572378 13542 572614
rect 12986 572058 13222 572294
rect 13306 572058 13542 572294
rect 12986 535178 13222 535414
rect 13306 535178 13542 535414
rect 12986 534858 13222 535094
rect 13306 534858 13542 535094
rect 12986 497978 13222 498214
rect 13306 497978 13542 498214
rect 12986 497658 13222 497894
rect 13306 497658 13542 497894
rect 12986 460778 13222 461014
rect 13306 460778 13542 461014
rect 12986 460458 13222 460694
rect 13306 460458 13542 460694
rect 12986 423578 13222 423814
rect 13306 423578 13542 423814
rect 12986 423258 13222 423494
rect 13306 423258 13542 423494
rect 12986 386378 13222 386614
rect 13306 386378 13542 386614
rect 12986 386058 13222 386294
rect 13306 386058 13542 386294
rect 12986 349178 13222 349414
rect 13306 349178 13542 349414
rect 12986 348858 13222 349094
rect 13306 348858 13542 349094
rect 12986 311978 13222 312214
rect 13306 311978 13542 312214
rect 12986 311658 13222 311894
rect 13306 311658 13542 311894
rect 12986 274778 13222 275014
rect 13306 274778 13542 275014
rect 12986 274458 13222 274694
rect 13306 274458 13542 274694
rect 12986 237578 13222 237814
rect 13306 237578 13542 237814
rect 12986 237258 13222 237494
rect 13306 237258 13542 237494
rect 12986 200378 13222 200614
rect 13306 200378 13542 200614
rect 12986 200058 13222 200294
rect 13306 200058 13542 200294
rect 12986 163178 13222 163414
rect 13306 163178 13542 163414
rect 12986 162858 13222 163094
rect 13306 162858 13542 163094
rect 12986 125978 13222 126214
rect 13306 125978 13542 126214
rect 12986 125658 13222 125894
rect 13306 125658 13542 125894
rect 12986 88778 13222 89014
rect 13306 88778 13542 89014
rect 12986 88458 13222 88694
rect 13306 88458 13542 88694
rect 12986 51578 13222 51814
rect 13306 51578 13542 51814
rect 12986 51258 13222 51494
rect 13306 51258 13542 51494
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect 16706 687698 16942 687934
rect 17026 687698 17262 687934
rect 16706 687378 16942 687614
rect 17026 687378 17262 687614
rect 16706 650498 16942 650734
rect 17026 650498 17262 650734
rect 16706 650178 16942 650414
rect 17026 650178 17262 650414
rect 16706 613298 16942 613534
rect 17026 613298 17262 613534
rect 16706 612978 16942 613214
rect 17026 612978 17262 613214
rect 16706 576098 16942 576334
rect 17026 576098 17262 576334
rect 16706 575778 16942 576014
rect 17026 575778 17262 576014
rect 16706 538898 16942 539134
rect 17026 538898 17262 539134
rect 16706 538578 16942 538814
rect 17026 538578 17262 538814
rect 16706 501698 16942 501934
rect 17026 501698 17262 501934
rect 16706 501378 16942 501614
rect 17026 501378 17262 501614
rect 16706 464498 16942 464734
rect 17026 464498 17262 464734
rect 16706 464178 16942 464414
rect 17026 464178 17262 464414
rect 16706 427298 16942 427534
rect 17026 427298 17262 427534
rect 16706 426978 16942 427214
rect 17026 426978 17262 427214
rect 16706 390098 16942 390334
rect 17026 390098 17262 390334
rect 16706 389778 16942 390014
rect 17026 389778 17262 390014
rect 16706 352898 16942 353134
rect 17026 352898 17262 353134
rect 16706 352578 16942 352814
rect 17026 352578 17262 352814
rect 16706 315698 16942 315934
rect 17026 315698 17262 315934
rect 16706 315378 16942 315614
rect 17026 315378 17262 315614
rect 16706 278498 16942 278734
rect 17026 278498 17262 278734
rect 16706 278178 16942 278414
rect 17026 278178 17262 278414
rect 16706 241298 16942 241534
rect 17026 241298 17262 241534
rect 16706 240978 16942 241214
rect 17026 240978 17262 241214
rect 16706 204098 16942 204334
rect 17026 204098 17262 204334
rect 16706 203778 16942 204014
rect 17026 203778 17262 204014
rect 16706 166898 16942 167134
rect 17026 166898 17262 167134
rect 16706 166578 16942 166814
rect 17026 166578 17262 166814
rect 16706 129698 16942 129934
rect 17026 129698 17262 129934
rect 16706 129378 16942 129614
rect 17026 129378 17262 129614
rect 16706 92498 16942 92734
rect 17026 92498 17262 92734
rect 16706 92178 16942 92414
rect 17026 92178 17262 92414
rect 16706 55298 16942 55534
rect 17026 55298 17262 55534
rect 16706 54978 16942 55214
rect 17026 54978 17262 55214
rect 16706 18098 16942 18334
rect 17026 18098 17262 18334
rect 16706 17778 16942 18014
rect 17026 17778 17262 18014
rect 20426 691418 20662 691654
rect 20746 691418 20982 691654
rect 20426 691098 20662 691334
rect 20746 691098 20982 691334
rect 20426 654218 20662 654454
rect 20746 654218 20982 654454
rect 20426 653898 20662 654134
rect 20746 653898 20982 654134
rect 20426 617018 20662 617254
rect 20746 617018 20982 617254
rect 20426 616698 20662 616934
rect 20746 616698 20982 616934
rect 20426 579818 20662 580054
rect 20746 579818 20982 580054
rect 20426 579498 20662 579734
rect 20746 579498 20982 579734
rect 20426 542618 20662 542854
rect 20746 542618 20982 542854
rect 20426 542298 20662 542534
rect 20746 542298 20982 542534
rect 20426 505418 20662 505654
rect 20746 505418 20982 505654
rect 20426 505098 20662 505334
rect 20746 505098 20982 505334
rect 20426 468218 20662 468454
rect 20746 468218 20982 468454
rect 20426 467898 20662 468134
rect 20746 467898 20982 468134
rect 20426 431018 20662 431254
rect 20746 431018 20982 431254
rect 20426 430698 20662 430934
rect 20746 430698 20982 430934
rect 20426 393818 20662 394054
rect 20746 393818 20982 394054
rect 20426 393498 20662 393734
rect 20746 393498 20982 393734
rect 20426 356618 20662 356854
rect 20746 356618 20982 356854
rect 20426 356298 20662 356534
rect 20746 356298 20982 356534
rect 20426 319418 20662 319654
rect 20746 319418 20982 319654
rect 20426 319098 20662 319334
rect 20746 319098 20982 319334
rect 20426 282218 20662 282454
rect 20746 282218 20982 282454
rect 20426 281898 20662 282134
rect 20746 281898 20982 282134
rect 20426 245018 20662 245254
rect 20746 245018 20982 245254
rect 20426 244698 20662 244934
rect 20746 244698 20982 244934
rect 20426 207818 20662 208054
rect 20746 207818 20982 208054
rect 20426 207498 20662 207734
rect 20746 207498 20982 207734
rect 20426 170618 20662 170854
rect 20746 170618 20982 170854
rect 20426 170298 20662 170534
rect 20746 170298 20982 170534
rect 20426 133418 20662 133654
rect 20746 133418 20982 133654
rect 20426 133098 20662 133334
rect 20746 133098 20982 133334
rect 20426 96218 20662 96454
rect 20746 96218 20982 96454
rect 20426 95898 20662 96134
rect 20746 95898 20982 96134
rect 20426 59018 20662 59254
rect 20746 59018 20982 59254
rect 20426 58698 20662 58934
rect 20746 58698 20982 58934
rect 20426 21818 20662 22054
rect 20746 21818 20982 22054
rect 20426 21498 20662 21734
rect 20746 21498 20982 21734
rect 24146 695138 24382 695374
rect 24466 695138 24702 695374
rect 24146 694818 24382 695054
rect 24466 694818 24702 695054
rect 24146 657938 24382 658174
rect 24466 657938 24702 658174
rect 24146 657618 24382 657854
rect 24466 657618 24702 657854
rect 24146 620738 24382 620974
rect 24466 620738 24702 620974
rect 24146 620418 24382 620654
rect 24466 620418 24702 620654
rect 24146 583538 24382 583774
rect 24466 583538 24702 583774
rect 24146 583218 24382 583454
rect 24466 583218 24702 583454
rect 24146 546338 24382 546574
rect 24466 546338 24702 546574
rect 24146 546018 24382 546254
rect 24466 546018 24702 546254
rect 24146 509138 24382 509374
rect 24466 509138 24702 509374
rect 24146 508818 24382 509054
rect 24466 508818 24702 509054
rect 24146 471938 24382 472174
rect 24466 471938 24702 472174
rect 24146 471618 24382 471854
rect 24466 471618 24702 471854
rect 24146 434738 24382 434974
rect 24466 434738 24702 434974
rect 24146 434418 24382 434654
rect 24466 434418 24702 434654
rect 24146 397538 24382 397774
rect 24466 397538 24702 397774
rect 24146 397218 24382 397454
rect 24466 397218 24702 397454
rect 24146 360338 24382 360574
rect 24466 360338 24702 360574
rect 24146 360018 24382 360254
rect 24466 360018 24702 360254
rect 24146 323138 24382 323374
rect 24466 323138 24702 323374
rect 24146 322818 24382 323054
rect 24466 322818 24702 323054
rect 24146 285938 24382 286174
rect 24466 285938 24702 286174
rect 24146 285618 24382 285854
rect 24466 285618 24702 285854
rect 24146 248738 24382 248974
rect 24466 248738 24702 248974
rect 24146 248418 24382 248654
rect 24466 248418 24702 248654
rect 24146 211538 24382 211774
rect 24466 211538 24702 211774
rect 24146 211218 24382 211454
rect 24466 211218 24702 211454
rect 24146 174338 24382 174574
rect 24466 174338 24702 174574
rect 24146 174018 24382 174254
rect 24466 174018 24702 174254
rect 24146 137138 24382 137374
rect 24466 137138 24702 137374
rect 24146 136818 24382 137054
rect 24466 136818 24702 137054
rect 24146 99938 24382 100174
rect 24466 99938 24702 100174
rect 24146 99618 24382 99854
rect 24466 99618 24702 99854
rect 24146 62738 24382 62974
rect 24466 62738 24702 62974
rect 24146 62418 24382 62654
rect 24466 62418 24702 62654
rect 24146 25538 24382 25774
rect 24466 25538 24702 25774
rect 24146 25218 24382 25454
rect 24466 25218 24702 25454
rect 27866 698858 28102 699094
rect 28186 698858 28422 699094
rect 27866 698538 28102 698774
rect 28186 698538 28422 698774
rect 27866 661658 28102 661894
rect 28186 661658 28422 661894
rect 27866 661338 28102 661574
rect 28186 661338 28422 661574
rect 27866 624458 28102 624694
rect 28186 624458 28422 624694
rect 27866 624138 28102 624374
rect 28186 624138 28422 624374
rect 27866 587258 28102 587494
rect 28186 587258 28422 587494
rect 27866 586938 28102 587174
rect 28186 586938 28422 587174
rect 27866 550058 28102 550294
rect 28186 550058 28422 550294
rect 27866 549738 28102 549974
rect 28186 549738 28422 549974
rect 27866 512858 28102 513094
rect 28186 512858 28422 513094
rect 27866 512538 28102 512774
rect 28186 512538 28422 512774
rect 27866 475658 28102 475894
rect 28186 475658 28422 475894
rect 27866 475338 28102 475574
rect 28186 475338 28422 475574
rect 27866 438458 28102 438694
rect 28186 438458 28422 438694
rect 27866 438138 28102 438374
rect 28186 438138 28422 438374
rect 27866 401258 28102 401494
rect 28186 401258 28422 401494
rect 27866 400938 28102 401174
rect 28186 400938 28422 401174
rect 27866 364058 28102 364294
rect 28186 364058 28422 364294
rect 27866 363738 28102 363974
rect 28186 363738 28422 363974
rect 27866 326858 28102 327094
rect 28186 326858 28422 327094
rect 27866 326538 28102 326774
rect 28186 326538 28422 326774
rect 27866 289658 28102 289894
rect 28186 289658 28422 289894
rect 27866 289338 28102 289574
rect 28186 289338 28422 289574
rect 27866 252458 28102 252694
rect 28186 252458 28422 252694
rect 27866 252138 28102 252374
rect 28186 252138 28422 252374
rect 27866 215258 28102 215494
rect 28186 215258 28422 215494
rect 27866 214938 28102 215174
rect 28186 214938 28422 215174
rect 27866 178058 28102 178294
rect 28186 178058 28422 178294
rect 27866 177738 28102 177974
rect 28186 177738 28422 177974
rect 27866 140858 28102 141094
rect 28186 140858 28422 141094
rect 27866 140538 28102 140774
rect 28186 140538 28422 140774
rect 27866 103658 28102 103894
rect 28186 103658 28422 103894
rect 27866 103338 28102 103574
rect 28186 103338 28422 103574
rect 27866 66458 28102 66694
rect 28186 66458 28422 66694
rect 27866 66138 28102 66374
rect 28186 66138 28422 66374
rect 27866 29258 28102 29494
rect 28186 29258 28422 29494
rect 27866 28938 28102 29174
rect 28186 28938 28422 29174
rect 39026 672818 39262 673054
rect 39346 672818 39582 673054
rect 39026 672498 39262 672734
rect 39346 672498 39582 672734
rect 39026 635618 39262 635854
rect 39346 635618 39582 635854
rect 39026 635298 39262 635534
rect 39346 635298 39582 635534
rect 39026 598418 39262 598654
rect 39346 598418 39582 598654
rect 39026 598098 39262 598334
rect 39346 598098 39582 598334
rect 39026 561218 39262 561454
rect 39346 561218 39582 561454
rect 39026 560898 39262 561134
rect 39346 560898 39582 561134
rect 39026 524018 39262 524254
rect 39346 524018 39582 524254
rect 39026 523698 39262 523934
rect 39346 523698 39582 523934
rect 39026 486818 39262 487054
rect 39346 486818 39582 487054
rect 39026 486498 39262 486734
rect 39346 486498 39582 486734
rect 39026 449618 39262 449854
rect 39346 449618 39582 449854
rect 39026 449298 39262 449534
rect 39346 449298 39582 449534
rect 39026 412418 39262 412654
rect 39346 412418 39582 412654
rect 39026 412098 39262 412334
rect 39346 412098 39582 412334
rect 39026 375218 39262 375454
rect 39346 375218 39582 375454
rect 39026 374898 39262 375134
rect 39346 374898 39582 375134
rect 39026 338018 39262 338254
rect 39346 338018 39582 338254
rect 39026 337698 39262 337934
rect 39346 337698 39582 337934
rect 39026 300818 39262 301054
rect 39346 300818 39582 301054
rect 39026 300498 39262 300734
rect 39346 300498 39582 300734
rect 39026 263618 39262 263854
rect 39346 263618 39582 263854
rect 39026 263298 39262 263534
rect 39346 263298 39582 263534
rect 39026 226418 39262 226654
rect 39346 226418 39582 226654
rect 39026 226098 39262 226334
rect 39346 226098 39582 226334
rect 39026 189218 39262 189454
rect 39346 189218 39582 189454
rect 39026 188898 39262 189134
rect 39346 188898 39582 189134
rect 39026 152018 39262 152254
rect 39346 152018 39582 152254
rect 39026 151698 39262 151934
rect 39346 151698 39582 151934
rect 39026 114818 39262 115054
rect 39346 114818 39582 115054
rect 39026 114498 39262 114734
rect 39346 114498 39582 114734
rect 39026 77618 39262 77854
rect 39346 77618 39582 77854
rect 39026 77298 39262 77534
rect 39346 77298 39582 77534
rect 39026 40418 39262 40654
rect 39346 40418 39582 40654
rect 39026 40098 39262 40334
rect 39346 40098 39582 40334
rect 39026 3218 39262 3454
rect 39346 3218 39582 3454
rect 39026 2898 39262 3134
rect 39346 2898 39582 3134
rect 42746 676538 42982 676774
rect 43066 676538 43302 676774
rect 42746 676218 42982 676454
rect 43066 676218 43302 676454
rect 42746 639338 42982 639574
rect 43066 639338 43302 639574
rect 42746 639018 42982 639254
rect 43066 639018 43302 639254
rect 42746 602138 42982 602374
rect 43066 602138 43302 602374
rect 42746 601818 42982 602054
rect 43066 601818 43302 602054
rect 42746 564938 42982 565174
rect 43066 564938 43302 565174
rect 42746 564618 42982 564854
rect 43066 564618 43302 564854
rect 42746 527738 42982 527974
rect 43066 527738 43302 527974
rect 42746 527418 42982 527654
rect 43066 527418 43302 527654
rect 42746 490538 42982 490774
rect 43066 490538 43302 490774
rect 42746 490218 42982 490454
rect 43066 490218 43302 490454
rect 42746 453338 42982 453574
rect 43066 453338 43302 453574
rect 42746 453018 42982 453254
rect 43066 453018 43302 453254
rect 42746 416138 42982 416374
rect 43066 416138 43302 416374
rect 42746 415818 42982 416054
rect 43066 415818 43302 416054
rect 42746 378938 42982 379174
rect 43066 378938 43302 379174
rect 42746 378618 42982 378854
rect 43066 378618 43302 378854
rect 42746 341738 42982 341974
rect 43066 341738 43302 341974
rect 42746 341418 42982 341654
rect 43066 341418 43302 341654
rect 42746 304538 42982 304774
rect 43066 304538 43302 304774
rect 42746 304218 42982 304454
rect 43066 304218 43302 304454
rect 42746 267338 42982 267574
rect 43066 267338 43302 267574
rect 42746 267018 42982 267254
rect 43066 267018 43302 267254
rect 42746 230138 42982 230374
rect 43066 230138 43302 230374
rect 42746 229818 42982 230054
rect 43066 229818 43302 230054
rect 42746 192938 42982 193174
rect 43066 192938 43302 193174
rect 42746 192618 42982 192854
rect 43066 192618 43302 192854
rect 42746 155738 42982 155974
rect 43066 155738 43302 155974
rect 42746 155418 42982 155654
rect 43066 155418 43302 155654
rect 42746 118538 42982 118774
rect 43066 118538 43302 118774
rect 42746 118218 42982 118454
rect 43066 118218 43302 118454
rect 42746 81338 42982 81574
rect 43066 81338 43302 81574
rect 42746 81018 42982 81254
rect 43066 81018 43302 81254
rect 42746 44138 42982 44374
rect 43066 44138 43302 44374
rect 42746 43818 42982 44054
rect 43066 43818 43302 44054
rect 42746 6938 42982 7174
rect 43066 6938 43302 7174
rect 42746 6618 42982 6854
rect 43066 6618 43302 6854
rect 46466 680258 46702 680494
rect 46786 680258 47022 680494
rect 46466 679938 46702 680174
rect 46786 679938 47022 680174
rect 46466 643058 46702 643294
rect 46786 643058 47022 643294
rect 46466 642738 46702 642974
rect 46786 642738 47022 642974
rect 46466 605858 46702 606094
rect 46786 605858 47022 606094
rect 46466 605538 46702 605774
rect 46786 605538 47022 605774
rect 46466 568658 46702 568894
rect 46786 568658 47022 568894
rect 46466 568338 46702 568574
rect 46786 568338 47022 568574
rect 46466 531458 46702 531694
rect 46786 531458 47022 531694
rect 46466 531138 46702 531374
rect 46786 531138 47022 531374
rect 46466 494258 46702 494494
rect 46786 494258 47022 494494
rect 46466 493938 46702 494174
rect 46786 493938 47022 494174
rect 46466 457058 46702 457294
rect 46786 457058 47022 457294
rect 46466 456738 46702 456974
rect 46786 456738 47022 456974
rect 46466 419858 46702 420094
rect 46786 419858 47022 420094
rect 46466 419538 46702 419774
rect 46786 419538 47022 419774
rect 46466 382658 46702 382894
rect 46786 382658 47022 382894
rect 46466 382338 46702 382574
rect 46786 382338 47022 382574
rect 46466 345458 46702 345694
rect 46786 345458 47022 345694
rect 46466 345138 46702 345374
rect 46786 345138 47022 345374
rect 46466 308258 46702 308494
rect 46786 308258 47022 308494
rect 46466 307938 46702 308174
rect 46786 307938 47022 308174
rect 46466 271058 46702 271294
rect 46786 271058 47022 271294
rect 46466 270738 46702 270974
rect 46786 270738 47022 270974
rect 46466 233858 46702 234094
rect 46786 233858 47022 234094
rect 46466 233538 46702 233774
rect 46786 233538 47022 233774
rect 46466 196658 46702 196894
rect 46786 196658 47022 196894
rect 46466 196338 46702 196574
rect 46786 196338 47022 196574
rect 46466 159458 46702 159694
rect 46786 159458 47022 159694
rect 46466 159138 46702 159374
rect 46786 159138 47022 159374
rect 46466 122258 46702 122494
rect 46786 122258 47022 122494
rect 46466 121938 46702 122174
rect 46786 121938 47022 122174
rect 46466 85058 46702 85294
rect 46786 85058 47022 85294
rect 46466 84738 46702 84974
rect 46786 84738 47022 84974
rect 46466 47858 46702 48094
rect 46786 47858 47022 48094
rect 46466 47538 46702 47774
rect 46786 47538 47022 47774
rect 46466 10658 46702 10894
rect 46786 10658 47022 10894
rect 46466 10338 46702 10574
rect 46786 10338 47022 10574
rect 50186 683978 50422 684214
rect 50506 683978 50742 684214
rect 50186 683658 50422 683894
rect 50506 683658 50742 683894
rect 50186 646778 50422 647014
rect 50506 646778 50742 647014
rect 50186 646458 50422 646694
rect 50506 646458 50742 646694
rect 50186 609578 50422 609814
rect 50506 609578 50742 609814
rect 50186 609258 50422 609494
rect 50506 609258 50742 609494
rect 50186 572378 50422 572614
rect 50506 572378 50742 572614
rect 50186 572058 50422 572294
rect 50506 572058 50742 572294
rect 50186 535178 50422 535414
rect 50506 535178 50742 535414
rect 50186 534858 50422 535094
rect 50506 534858 50742 535094
rect 50186 497978 50422 498214
rect 50506 497978 50742 498214
rect 50186 497658 50422 497894
rect 50506 497658 50742 497894
rect 50186 460778 50422 461014
rect 50506 460778 50742 461014
rect 50186 460458 50422 460694
rect 50506 460458 50742 460694
rect 50186 423578 50422 423814
rect 50506 423578 50742 423814
rect 50186 423258 50422 423494
rect 50506 423258 50742 423494
rect 50186 386378 50422 386614
rect 50506 386378 50742 386614
rect 50186 386058 50422 386294
rect 50506 386058 50742 386294
rect 50186 349178 50422 349414
rect 50506 349178 50742 349414
rect 50186 348858 50422 349094
rect 50506 348858 50742 349094
rect 50186 311978 50422 312214
rect 50506 311978 50742 312214
rect 50186 311658 50422 311894
rect 50506 311658 50742 311894
rect 50186 274778 50422 275014
rect 50506 274778 50742 275014
rect 50186 274458 50422 274694
rect 50506 274458 50742 274694
rect 50186 237578 50422 237814
rect 50506 237578 50742 237814
rect 50186 237258 50422 237494
rect 50506 237258 50742 237494
rect 50186 200378 50422 200614
rect 50506 200378 50742 200614
rect 50186 200058 50422 200294
rect 50506 200058 50742 200294
rect 50186 163178 50422 163414
rect 50506 163178 50742 163414
rect 50186 162858 50422 163094
rect 50506 162858 50742 163094
rect 50186 125978 50422 126214
rect 50506 125978 50742 126214
rect 50186 125658 50422 125894
rect 50506 125658 50742 125894
rect 50186 88778 50422 89014
rect 50506 88778 50742 89014
rect 50186 88458 50422 88694
rect 50506 88458 50742 88694
rect 50186 51578 50422 51814
rect 50506 51578 50742 51814
rect 50186 51258 50422 51494
rect 50506 51258 50742 51494
rect 50186 14378 50422 14614
rect 50506 14378 50742 14614
rect 50186 14058 50422 14294
rect 50506 14058 50742 14294
rect 53906 687698 54142 687934
rect 54226 687698 54462 687934
rect 53906 687378 54142 687614
rect 54226 687378 54462 687614
rect 53906 650498 54142 650734
rect 54226 650498 54462 650734
rect 53906 650178 54142 650414
rect 54226 650178 54462 650414
rect 53906 613298 54142 613534
rect 54226 613298 54462 613534
rect 53906 612978 54142 613214
rect 54226 612978 54462 613214
rect 53906 576098 54142 576334
rect 54226 576098 54462 576334
rect 53906 575778 54142 576014
rect 54226 575778 54462 576014
rect 53906 538898 54142 539134
rect 54226 538898 54462 539134
rect 53906 538578 54142 538814
rect 54226 538578 54462 538814
rect 53906 501698 54142 501934
rect 54226 501698 54462 501934
rect 53906 501378 54142 501614
rect 54226 501378 54462 501614
rect 53906 464498 54142 464734
rect 54226 464498 54462 464734
rect 53906 464178 54142 464414
rect 54226 464178 54462 464414
rect 53906 427298 54142 427534
rect 54226 427298 54462 427534
rect 53906 426978 54142 427214
rect 54226 426978 54462 427214
rect 53906 390098 54142 390334
rect 54226 390098 54462 390334
rect 53906 389778 54142 390014
rect 54226 389778 54462 390014
rect 53906 352898 54142 353134
rect 54226 352898 54462 353134
rect 53906 352578 54142 352814
rect 54226 352578 54462 352814
rect 53906 315698 54142 315934
rect 54226 315698 54462 315934
rect 53906 315378 54142 315614
rect 54226 315378 54462 315614
rect 53906 278498 54142 278734
rect 54226 278498 54462 278734
rect 53906 278178 54142 278414
rect 54226 278178 54462 278414
rect 53906 241298 54142 241534
rect 54226 241298 54462 241534
rect 53906 240978 54142 241214
rect 54226 240978 54462 241214
rect 53906 204098 54142 204334
rect 54226 204098 54462 204334
rect 53906 203778 54142 204014
rect 54226 203778 54462 204014
rect 53906 166898 54142 167134
rect 54226 166898 54462 167134
rect 53906 166578 54142 166814
rect 54226 166578 54462 166814
rect 53906 129698 54142 129934
rect 54226 129698 54462 129934
rect 53906 129378 54142 129614
rect 54226 129378 54462 129614
rect 53906 92498 54142 92734
rect 54226 92498 54462 92734
rect 53906 92178 54142 92414
rect 54226 92178 54462 92414
rect 53906 55298 54142 55534
rect 54226 55298 54462 55534
rect 53906 54978 54142 55214
rect 54226 54978 54462 55214
rect 53906 18098 54142 18334
rect 54226 18098 54462 18334
rect 53906 17778 54142 18014
rect 54226 17778 54462 18014
rect 57626 691418 57862 691654
rect 57946 691418 58182 691654
rect 57626 691098 57862 691334
rect 57946 691098 58182 691334
rect 57626 654218 57862 654454
rect 57946 654218 58182 654454
rect 57626 653898 57862 654134
rect 57946 653898 58182 654134
rect 57626 617018 57862 617254
rect 57946 617018 58182 617254
rect 57626 616698 57862 616934
rect 57946 616698 58182 616934
rect 57626 579818 57862 580054
rect 57946 579818 58182 580054
rect 57626 579498 57862 579734
rect 57946 579498 58182 579734
rect 57626 542618 57862 542854
rect 57946 542618 58182 542854
rect 57626 542298 57862 542534
rect 57946 542298 58182 542534
rect 57626 505418 57862 505654
rect 57946 505418 58182 505654
rect 57626 505098 57862 505334
rect 57946 505098 58182 505334
rect 57626 468218 57862 468454
rect 57946 468218 58182 468454
rect 57626 467898 57862 468134
rect 57946 467898 58182 468134
rect 57626 431018 57862 431254
rect 57946 431018 58182 431254
rect 57626 430698 57862 430934
rect 57946 430698 58182 430934
rect 57626 393818 57862 394054
rect 57946 393818 58182 394054
rect 57626 393498 57862 393734
rect 57946 393498 58182 393734
rect 57626 356618 57862 356854
rect 57946 356618 58182 356854
rect 57626 356298 57862 356534
rect 57946 356298 58182 356534
rect 57626 319418 57862 319654
rect 57946 319418 58182 319654
rect 57626 319098 57862 319334
rect 57946 319098 58182 319334
rect 57626 282218 57862 282454
rect 57946 282218 58182 282454
rect 57626 281898 57862 282134
rect 57946 281898 58182 282134
rect 57626 245018 57862 245254
rect 57946 245018 58182 245254
rect 57626 244698 57862 244934
rect 57946 244698 58182 244934
rect 57626 207818 57862 208054
rect 57946 207818 58182 208054
rect 57626 207498 57862 207734
rect 57946 207498 58182 207734
rect 57626 170618 57862 170854
rect 57946 170618 58182 170854
rect 57626 170298 57862 170534
rect 57946 170298 58182 170534
rect 57626 133418 57862 133654
rect 57946 133418 58182 133654
rect 57626 133098 57862 133334
rect 57946 133098 58182 133334
rect 57626 96218 57862 96454
rect 57946 96218 58182 96454
rect 57626 95898 57862 96134
rect 57946 95898 58182 96134
rect 57626 59018 57862 59254
rect 57946 59018 58182 59254
rect 57626 58698 57862 58934
rect 57946 58698 58182 58934
rect 57626 21818 57862 22054
rect 57946 21818 58182 22054
rect 57626 21498 57862 21734
rect 57946 21498 58182 21734
rect 61346 695138 61582 695374
rect 61666 695138 61902 695374
rect 61346 694818 61582 695054
rect 61666 694818 61902 695054
rect 61346 657938 61582 658174
rect 61666 657938 61902 658174
rect 61346 657618 61582 657854
rect 61666 657618 61902 657854
rect 61346 620738 61582 620974
rect 61666 620738 61902 620974
rect 61346 620418 61582 620654
rect 61666 620418 61902 620654
rect 61346 583538 61582 583774
rect 61666 583538 61902 583774
rect 61346 583218 61582 583454
rect 61666 583218 61902 583454
rect 61346 546338 61582 546574
rect 61666 546338 61902 546574
rect 61346 546018 61582 546254
rect 61666 546018 61902 546254
rect 61346 509138 61582 509374
rect 61666 509138 61902 509374
rect 61346 508818 61582 509054
rect 61666 508818 61902 509054
rect 61346 471938 61582 472174
rect 61666 471938 61902 472174
rect 61346 471618 61582 471854
rect 61666 471618 61902 471854
rect 61346 434738 61582 434974
rect 61666 434738 61902 434974
rect 61346 434418 61582 434654
rect 61666 434418 61902 434654
rect 61346 397538 61582 397774
rect 61666 397538 61902 397774
rect 61346 397218 61582 397454
rect 61666 397218 61902 397454
rect 61346 360338 61582 360574
rect 61666 360338 61902 360574
rect 61346 360018 61582 360254
rect 61666 360018 61902 360254
rect 61346 323138 61582 323374
rect 61666 323138 61902 323374
rect 61346 322818 61582 323054
rect 61666 322818 61902 323054
rect 61346 285938 61582 286174
rect 61666 285938 61902 286174
rect 61346 285618 61582 285854
rect 61666 285618 61902 285854
rect 61346 248738 61582 248974
rect 61666 248738 61902 248974
rect 61346 248418 61582 248654
rect 61666 248418 61902 248654
rect 61346 211538 61582 211774
rect 61666 211538 61902 211774
rect 61346 211218 61582 211454
rect 61666 211218 61902 211454
rect 61346 174338 61582 174574
rect 61666 174338 61902 174574
rect 61346 174018 61582 174254
rect 61666 174018 61902 174254
rect 61346 137138 61582 137374
rect 61666 137138 61902 137374
rect 61346 136818 61582 137054
rect 61666 136818 61902 137054
rect 61346 99938 61582 100174
rect 61666 99938 61902 100174
rect 61346 99618 61582 99854
rect 61666 99618 61902 99854
rect 61346 62738 61582 62974
rect 61666 62738 61902 62974
rect 61346 62418 61582 62654
rect 61666 62418 61902 62654
rect 61346 25538 61582 25774
rect 61666 25538 61902 25774
rect 61346 25218 61582 25454
rect 61666 25218 61902 25454
rect 65066 698858 65302 699094
rect 65386 698858 65622 699094
rect 65066 698538 65302 698774
rect 65386 698538 65622 698774
rect 65066 661658 65302 661894
rect 65386 661658 65622 661894
rect 65066 661338 65302 661574
rect 65386 661338 65622 661574
rect 65066 624458 65302 624694
rect 65386 624458 65622 624694
rect 65066 624138 65302 624374
rect 65386 624138 65622 624374
rect 65066 587258 65302 587494
rect 65386 587258 65622 587494
rect 65066 586938 65302 587174
rect 65386 586938 65622 587174
rect 65066 550058 65302 550294
rect 65386 550058 65622 550294
rect 65066 549738 65302 549974
rect 65386 549738 65622 549974
rect 65066 512858 65302 513094
rect 65386 512858 65622 513094
rect 65066 512538 65302 512774
rect 65386 512538 65622 512774
rect 65066 475658 65302 475894
rect 65386 475658 65622 475894
rect 65066 475338 65302 475574
rect 65386 475338 65622 475574
rect 65066 438458 65302 438694
rect 65386 438458 65622 438694
rect 65066 438138 65302 438374
rect 65386 438138 65622 438374
rect 65066 401258 65302 401494
rect 65386 401258 65622 401494
rect 65066 400938 65302 401174
rect 65386 400938 65622 401174
rect 65066 364058 65302 364294
rect 65386 364058 65622 364294
rect 65066 363738 65302 363974
rect 65386 363738 65622 363974
rect 65066 326858 65302 327094
rect 65386 326858 65622 327094
rect 65066 326538 65302 326774
rect 65386 326538 65622 326774
rect 65066 289658 65302 289894
rect 65386 289658 65622 289894
rect 65066 289338 65302 289574
rect 65386 289338 65622 289574
rect 65066 252458 65302 252694
rect 65386 252458 65622 252694
rect 65066 252138 65302 252374
rect 65386 252138 65622 252374
rect 65066 215258 65302 215494
rect 65386 215258 65622 215494
rect 65066 214938 65302 215174
rect 65386 214938 65622 215174
rect 65066 178058 65302 178294
rect 65386 178058 65622 178294
rect 65066 177738 65302 177974
rect 65386 177738 65622 177974
rect 65066 140858 65302 141094
rect 65386 140858 65622 141094
rect 65066 140538 65302 140774
rect 65386 140538 65622 140774
rect 65066 103658 65302 103894
rect 65386 103658 65622 103894
rect 65066 103338 65302 103574
rect 65386 103338 65622 103574
rect 65066 66458 65302 66694
rect 65386 66458 65622 66694
rect 65066 66138 65302 66374
rect 65386 66138 65622 66374
rect 65066 29258 65302 29494
rect 65386 29258 65622 29494
rect 65066 28938 65302 29174
rect 65386 28938 65622 29174
rect 76226 672818 76462 673054
rect 76546 672818 76782 673054
rect 76226 672498 76462 672734
rect 76546 672498 76782 672734
rect 76226 635618 76462 635854
rect 76546 635618 76782 635854
rect 76226 635298 76462 635534
rect 76546 635298 76782 635534
rect 76226 598418 76462 598654
rect 76546 598418 76782 598654
rect 76226 598098 76462 598334
rect 76546 598098 76782 598334
rect 76226 561218 76462 561454
rect 76546 561218 76782 561454
rect 76226 560898 76462 561134
rect 76546 560898 76782 561134
rect 76226 524018 76462 524254
rect 76546 524018 76782 524254
rect 76226 523698 76462 523934
rect 76546 523698 76782 523934
rect 76226 486818 76462 487054
rect 76546 486818 76782 487054
rect 76226 486498 76462 486734
rect 76546 486498 76782 486734
rect 76226 449618 76462 449854
rect 76546 449618 76782 449854
rect 76226 449298 76462 449534
rect 76546 449298 76782 449534
rect 76226 412418 76462 412654
rect 76546 412418 76782 412654
rect 76226 412098 76462 412334
rect 76546 412098 76782 412334
rect 76226 375218 76462 375454
rect 76546 375218 76782 375454
rect 76226 374898 76462 375134
rect 76546 374898 76782 375134
rect 76226 338018 76462 338254
rect 76546 338018 76782 338254
rect 76226 337698 76462 337934
rect 76546 337698 76782 337934
rect 76226 300818 76462 301054
rect 76546 300818 76782 301054
rect 76226 300498 76462 300734
rect 76546 300498 76782 300734
rect 76226 263618 76462 263854
rect 76546 263618 76782 263854
rect 76226 263298 76462 263534
rect 76546 263298 76782 263534
rect 76226 226418 76462 226654
rect 76546 226418 76782 226654
rect 76226 226098 76462 226334
rect 76546 226098 76782 226334
rect 76226 189218 76462 189454
rect 76546 189218 76782 189454
rect 76226 188898 76462 189134
rect 76546 188898 76782 189134
rect 76226 152018 76462 152254
rect 76546 152018 76782 152254
rect 76226 151698 76462 151934
rect 76546 151698 76782 151934
rect 76226 114818 76462 115054
rect 76546 114818 76782 115054
rect 76226 114498 76462 114734
rect 76546 114498 76782 114734
rect 76226 77618 76462 77854
rect 76546 77618 76782 77854
rect 76226 77298 76462 77534
rect 76546 77298 76782 77534
rect 76226 40418 76462 40654
rect 76546 40418 76782 40654
rect 76226 40098 76462 40334
rect 76546 40098 76782 40334
rect 76226 3218 76462 3454
rect 76546 3218 76782 3454
rect 76226 2898 76462 3134
rect 76546 2898 76782 3134
rect 79946 676538 80182 676774
rect 80266 676538 80502 676774
rect 79946 676218 80182 676454
rect 80266 676218 80502 676454
rect 79946 639338 80182 639574
rect 80266 639338 80502 639574
rect 79946 639018 80182 639254
rect 80266 639018 80502 639254
rect 79946 602138 80182 602374
rect 80266 602138 80502 602374
rect 79946 601818 80182 602054
rect 80266 601818 80502 602054
rect 79946 564938 80182 565174
rect 80266 564938 80502 565174
rect 79946 564618 80182 564854
rect 80266 564618 80502 564854
rect 79946 527738 80182 527974
rect 80266 527738 80502 527974
rect 79946 527418 80182 527654
rect 80266 527418 80502 527654
rect 79946 490538 80182 490774
rect 80266 490538 80502 490774
rect 79946 490218 80182 490454
rect 80266 490218 80502 490454
rect 79946 453338 80182 453574
rect 80266 453338 80502 453574
rect 79946 453018 80182 453254
rect 80266 453018 80502 453254
rect 79946 416138 80182 416374
rect 80266 416138 80502 416374
rect 79946 415818 80182 416054
rect 80266 415818 80502 416054
rect 79946 378938 80182 379174
rect 80266 378938 80502 379174
rect 79946 378618 80182 378854
rect 80266 378618 80502 378854
rect 79946 341738 80182 341974
rect 80266 341738 80502 341974
rect 79946 341418 80182 341654
rect 80266 341418 80502 341654
rect 79946 304538 80182 304774
rect 80266 304538 80502 304774
rect 79946 304218 80182 304454
rect 80266 304218 80502 304454
rect 79946 267338 80182 267574
rect 80266 267338 80502 267574
rect 79946 267018 80182 267254
rect 80266 267018 80502 267254
rect 79946 230138 80182 230374
rect 80266 230138 80502 230374
rect 79946 229818 80182 230054
rect 80266 229818 80502 230054
rect 79946 192938 80182 193174
rect 80266 192938 80502 193174
rect 79946 192618 80182 192854
rect 80266 192618 80502 192854
rect 79946 155738 80182 155974
rect 80266 155738 80502 155974
rect 79946 155418 80182 155654
rect 80266 155418 80502 155654
rect 79946 118538 80182 118774
rect 80266 118538 80502 118774
rect 79946 118218 80182 118454
rect 80266 118218 80502 118454
rect 79946 81338 80182 81574
rect 80266 81338 80502 81574
rect 79946 81018 80182 81254
rect 80266 81018 80502 81254
rect 79946 44138 80182 44374
rect 80266 44138 80502 44374
rect 79946 43818 80182 44054
rect 80266 43818 80502 44054
rect 79946 6938 80182 7174
rect 80266 6938 80502 7174
rect 79946 6618 80182 6854
rect 80266 6618 80502 6854
rect 83666 680258 83902 680494
rect 83986 680258 84222 680494
rect 83666 679938 83902 680174
rect 83986 679938 84222 680174
rect 83666 643058 83902 643294
rect 83986 643058 84222 643294
rect 83666 642738 83902 642974
rect 83986 642738 84222 642974
rect 83666 605858 83902 606094
rect 83986 605858 84222 606094
rect 83666 605538 83902 605774
rect 83986 605538 84222 605774
rect 83666 568658 83902 568894
rect 83986 568658 84222 568894
rect 83666 568338 83902 568574
rect 83986 568338 84222 568574
rect 83666 531458 83902 531694
rect 83986 531458 84222 531694
rect 83666 531138 83902 531374
rect 83986 531138 84222 531374
rect 83666 494258 83902 494494
rect 83986 494258 84222 494494
rect 83666 493938 83902 494174
rect 83986 493938 84222 494174
rect 83666 457058 83902 457294
rect 83986 457058 84222 457294
rect 83666 456738 83902 456974
rect 83986 456738 84222 456974
rect 83666 419858 83902 420094
rect 83986 419858 84222 420094
rect 83666 419538 83902 419774
rect 83986 419538 84222 419774
rect 83666 382658 83902 382894
rect 83986 382658 84222 382894
rect 83666 382338 83902 382574
rect 83986 382338 84222 382574
rect 83666 345458 83902 345694
rect 83986 345458 84222 345694
rect 83666 345138 83902 345374
rect 83986 345138 84222 345374
rect 83666 308258 83902 308494
rect 83986 308258 84222 308494
rect 83666 307938 83902 308174
rect 83986 307938 84222 308174
rect 83666 271058 83902 271294
rect 83986 271058 84222 271294
rect 83666 270738 83902 270974
rect 83986 270738 84222 270974
rect 83666 233858 83902 234094
rect 83986 233858 84222 234094
rect 83666 233538 83902 233774
rect 83986 233538 84222 233774
rect 83666 196658 83902 196894
rect 83986 196658 84222 196894
rect 83666 196338 83902 196574
rect 83986 196338 84222 196574
rect 83666 159458 83902 159694
rect 83986 159458 84222 159694
rect 83666 159138 83902 159374
rect 83986 159138 84222 159374
rect 83666 122258 83902 122494
rect 83986 122258 84222 122494
rect 83666 121938 83902 122174
rect 83986 121938 84222 122174
rect 83666 85058 83902 85294
rect 83986 85058 84222 85294
rect 83666 84738 83902 84974
rect 83986 84738 84222 84974
rect 83666 47858 83902 48094
rect 83986 47858 84222 48094
rect 83666 47538 83902 47774
rect 83986 47538 84222 47774
rect 83666 10658 83902 10894
rect 83986 10658 84222 10894
rect 83666 10338 83902 10574
rect 83986 10338 84222 10574
rect 87386 683978 87622 684214
rect 87706 683978 87942 684214
rect 87386 683658 87622 683894
rect 87706 683658 87942 683894
rect 87386 646778 87622 647014
rect 87706 646778 87942 647014
rect 87386 646458 87622 646694
rect 87706 646458 87942 646694
rect 87386 609578 87622 609814
rect 87706 609578 87942 609814
rect 87386 609258 87622 609494
rect 87706 609258 87942 609494
rect 87386 572378 87622 572614
rect 87706 572378 87942 572614
rect 87386 572058 87622 572294
rect 87706 572058 87942 572294
rect 87386 535178 87622 535414
rect 87706 535178 87942 535414
rect 87386 534858 87622 535094
rect 87706 534858 87942 535094
rect 87386 497978 87622 498214
rect 87706 497978 87942 498214
rect 87386 497658 87622 497894
rect 87706 497658 87942 497894
rect 87386 460778 87622 461014
rect 87706 460778 87942 461014
rect 87386 460458 87622 460694
rect 87706 460458 87942 460694
rect 87386 423578 87622 423814
rect 87706 423578 87942 423814
rect 87386 423258 87622 423494
rect 87706 423258 87942 423494
rect 87386 386378 87622 386614
rect 87706 386378 87942 386614
rect 87386 386058 87622 386294
rect 87706 386058 87942 386294
rect 87386 349178 87622 349414
rect 87706 349178 87942 349414
rect 87386 348858 87622 349094
rect 87706 348858 87942 349094
rect 87386 311978 87622 312214
rect 87706 311978 87942 312214
rect 87386 311658 87622 311894
rect 87706 311658 87942 311894
rect 87386 274778 87622 275014
rect 87706 274778 87942 275014
rect 87386 274458 87622 274694
rect 87706 274458 87942 274694
rect 87386 237578 87622 237814
rect 87706 237578 87942 237814
rect 87386 237258 87622 237494
rect 87706 237258 87942 237494
rect 87386 200378 87622 200614
rect 87706 200378 87942 200614
rect 87386 200058 87622 200294
rect 87706 200058 87942 200294
rect 87386 163178 87622 163414
rect 87706 163178 87942 163414
rect 87386 162858 87622 163094
rect 87706 162858 87942 163094
rect 87386 125978 87622 126214
rect 87706 125978 87942 126214
rect 87386 125658 87622 125894
rect 87706 125658 87942 125894
rect 87386 88778 87622 89014
rect 87706 88778 87942 89014
rect 87386 88458 87622 88694
rect 87706 88458 87942 88694
rect 87386 51578 87622 51814
rect 87706 51578 87942 51814
rect 87386 51258 87622 51494
rect 87706 51258 87942 51494
rect 87386 14378 87622 14614
rect 87706 14378 87942 14614
rect 87386 14058 87622 14294
rect 87706 14058 87942 14294
rect 91106 687698 91342 687934
rect 91426 687698 91662 687934
rect 91106 687378 91342 687614
rect 91426 687378 91662 687614
rect 91106 650498 91342 650734
rect 91426 650498 91662 650734
rect 91106 650178 91342 650414
rect 91426 650178 91662 650414
rect 91106 613298 91342 613534
rect 91426 613298 91662 613534
rect 91106 612978 91342 613214
rect 91426 612978 91662 613214
rect 91106 576098 91342 576334
rect 91426 576098 91662 576334
rect 91106 575778 91342 576014
rect 91426 575778 91662 576014
rect 91106 538898 91342 539134
rect 91426 538898 91662 539134
rect 91106 538578 91342 538814
rect 91426 538578 91662 538814
rect 91106 501698 91342 501934
rect 91426 501698 91662 501934
rect 91106 501378 91342 501614
rect 91426 501378 91662 501614
rect 91106 464498 91342 464734
rect 91426 464498 91662 464734
rect 91106 464178 91342 464414
rect 91426 464178 91662 464414
rect 91106 427298 91342 427534
rect 91426 427298 91662 427534
rect 91106 426978 91342 427214
rect 91426 426978 91662 427214
rect 91106 390098 91342 390334
rect 91426 390098 91662 390334
rect 91106 389778 91342 390014
rect 91426 389778 91662 390014
rect 91106 352898 91342 353134
rect 91426 352898 91662 353134
rect 91106 352578 91342 352814
rect 91426 352578 91662 352814
rect 91106 315698 91342 315934
rect 91426 315698 91662 315934
rect 91106 315378 91342 315614
rect 91426 315378 91662 315614
rect 91106 278498 91342 278734
rect 91426 278498 91662 278734
rect 91106 278178 91342 278414
rect 91426 278178 91662 278414
rect 91106 241298 91342 241534
rect 91426 241298 91662 241534
rect 91106 240978 91342 241214
rect 91426 240978 91662 241214
rect 91106 204098 91342 204334
rect 91426 204098 91662 204334
rect 91106 203778 91342 204014
rect 91426 203778 91662 204014
rect 91106 166898 91342 167134
rect 91426 166898 91662 167134
rect 91106 166578 91342 166814
rect 91426 166578 91662 166814
rect 91106 129698 91342 129934
rect 91426 129698 91662 129934
rect 91106 129378 91342 129614
rect 91426 129378 91662 129614
rect 91106 92498 91342 92734
rect 91426 92498 91662 92734
rect 91106 92178 91342 92414
rect 91426 92178 91662 92414
rect 91106 55298 91342 55534
rect 91426 55298 91662 55534
rect 91106 54978 91342 55214
rect 91426 54978 91662 55214
rect 91106 18098 91342 18334
rect 91426 18098 91662 18334
rect 91106 17778 91342 18014
rect 91426 17778 91662 18014
rect 94826 691418 95062 691654
rect 95146 691418 95382 691654
rect 94826 691098 95062 691334
rect 95146 691098 95382 691334
rect 94826 654218 95062 654454
rect 95146 654218 95382 654454
rect 94826 653898 95062 654134
rect 95146 653898 95382 654134
rect 94826 617018 95062 617254
rect 95146 617018 95382 617254
rect 94826 616698 95062 616934
rect 95146 616698 95382 616934
rect 94826 579818 95062 580054
rect 95146 579818 95382 580054
rect 94826 579498 95062 579734
rect 95146 579498 95382 579734
rect 94826 542618 95062 542854
rect 95146 542618 95382 542854
rect 94826 542298 95062 542534
rect 95146 542298 95382 542534
rect 94826 505418 95062 505654
rect 95146 505418 95382 505654
rect 94826 505098 95062 505334
rect 95146 505098 95382 505334
rect 94826 468218 95062 468454
rect 95146 468218 95382 468454
rect 94826 467898 95062 468134
rect 95146 467898 95382 468134
rect 94826 431018 95062 431254
rect 95146 431018 95382 431254
rect 94826 430698 95062 430934
rect 95146 430698 95382 430934
rect 94826 393818 95062 394054
rect 95146 393818 95382 394054
rect 94826 393498 95062 393734
rect 95146 393498 95382 393734
rect 94826 356618 95062 356854
rect 95146 356618 95382 356854
rect 94826 356298 95062 356534
rect 95146 356298 95382 356534
rect 94826 319418 95062 319654
rect 95146 319418 95382 319654
rect 94826 319098 95062 319334
rect 95146 319098 95382 319334
rect 94826 282218 95062 282454
rect 95146 282218 95382 282454
rect 94826 281898 95062 282134
rect 95146 281898 95382 282134
rect 94826 245018 95062 245254
rect 95146 245018 95382 245254
rect 94826 244698 95062 244934
rect 95146 244698 95382 244934
rect 94826 207818 95062 208054
rect 95146 207818 95382 208054
rect 94826 207498 95062 207734
rect 95146 207498 95382 207734
rect 94826 170618 95062 170854
rect 95146 170618 95382 170854
rect 94826 170298 95062 170534
rect 95146 170298 95382 170534
rect 94826 133418 95062 133654
rect 95146 133418 95382 133654
rect 94826 133098 95062 133334
rect 95146 133098 95382 133334
rect 94826 96218 95062 96454
rect 95146 96218 95382 96454
rect 94826 95898 95062 96134
rect 95146 95898 95382 96134
rect 94826 59018 95062 59254
rect 95146 59018 95382 59254
rect 94826 58698 95062 58934
rect 95146 58698 95382 58934
rect 94826 21818 95062 22054
rect 95146 21818 95382 22054
rect 94826 21498 95062 21734
rect 95146 21498 95382 21734
rect 98546 695138 98782 695374
rect 98866 695138 99102 695374
rect 98546 694818 98782 695054
rect 98866 694818 99102 695054
rect 98546 657938 98782 658174
rect 98866 657938 99102 658174
rect 98546 657618 98782 657854
rect 98866 657618 99102 657854
rect 98546 620738 98782 620974
rect 98866 620738 99102 620974
rect 98546 620418 98782 620654
rect 98866 620418 99102 620654
rect 98546 583538 98782 583774
rect 98866 583538 99102 583774
rect 98546 583218 98782 583454
rect 98866 583218 99102 583454
rect 98546 546338 98782 546574
rect 98866 546338 99102 546574
rect 98546 546018 98782 546254
rect 98866 546018 99102 546254
rect 98546 509138 98782 509374
rect 98866 509138 99102 509374
rect 98546 508818 98782 509054
rect 98866 508818 99102 509054
rect 98546 471938 98782 472174
rect 98866 471938 99102 472174
rect 98546 471618 98782 471854
rect 98866 471618 99102 471854
rect 98546 434738 98782 434974
rect 98866 434738 99102 434974
rect 98546 434418 98782 434654
rect 98866 434418 99102 434654
rect 98546 397538 98782 397774
rect 98866 397538 99102 397774
rect 98546 397218 98782 397454
rect 98866 397218 99102 397454
rect 98546 360338 98782 360574
rect 98866 360338 99102 360574
rect 98546 360018 98782 360254
rect 98866 360018 99102 360254
rect 98546 323138 98782 323374
rect 98866 323138 99102 323374
rect 98546 322818 98782 323054
rect 98866 322818 99102 323054
rect 98546 285938 98782 286174
rect 98866 285938 99102 286174
rect 98546 285618 98782 285854
rect 98866 285618 99102 285854
rect 98546 248738 98782 248974
rect 98866 248738 99102 248974
rect 98546 248418 98782 248654
rect 98866 248418 99102 248654
rect 98546 211538 98782 211774
rect 98866 211538 99102 211774
rect 98546 211218 98782 211454
rect 98866 211218 99102 211454
rect 98546 174338 98782 174574
rect 98866 174338 99102 174574
rect 98546 174018 98782 174254
rect 98866 174018 99102 174254
rect 98546 137138 98782 137374
rect 98866 137138 99102 137374
rect 98546 136818 98782 137054
rect 98866 136818 99102 137054
rect 98546 99938 98782 100174
rect 98866 99938 99102 100174
rect 98546 99618 98782 99854
rect 98866 99618 99102 99854
rect 98546 62738 98782 62974
rect 98866 62738 99102 62974
rect 98546 62418 98782 62654
rect 98866 62418 99102 62654
rect 98546 25538 98782 25774
rect 98866 25538 99102 25774
rect 98546 25218 98782 25454
rect 98866 25218 99102 25454
rect 102266 698858 102502 699094
rect 102586 698858 102822 699094
rect 102266 698538 102502 698774
rect 102586 698538 102822 698774
rect 102266 661658 102502 661894
rect 102586 661658 102822 661894
rect 102266 661338 102502 661574
rect 102586 661338 102822 661574
rect 102266 624458 102502 624694
rect 102586 624458 102822 624694
rect 102266 624138 102502 624374
rect 102586 624138 102822 624374
rect 102266 587258 102502 587494
rect 102586 587258 102822 587494
rect 102266 586938 102502 587174
rect 102586 586938 102822 587174
rect 102266 550058 102502 550294
rect 102586 550058 102822 550294
rect 102266 549738 102502 549974
rect 102586 549738 102822 549974
rect 102266 512858 102502 513094
rect 102586 512858 102822 513094
rect 102266 512538 102502 512774
rect 102586 512538 102822 512774
rect 102266 475658 102502 475894
rect 102586 475658 102822 475894
rect 102266 475338 102502 475574
rect 102586 475338 102822 475574
rect 102266 438458 102502 438694
rect 102586 438458 102822 438694
rect 102266 438138 102502 438374
rect 102586 438138 102822 438374
rect 102266 401258 102502 401494
rect 102586 401258 102822 401494
rect 102266 400938 102502 401174
rect 102586 400938 102822 401174
rect 102266 364058 102502 364294
rect 102586 364058 102822 364294
rect 102266 363738 102502 363974
rect 102586 363738 102822 363974
rect 102266 326858 102502 327094
rect 102586 326858 102822 327094
rect 102266 326538 102502 326774
rect 102586 326538 102822 326774
rect 102266 289658 102502 289894
rect 102586 289658 102822 289894
rect 102266 289338 102502 289574
rect 102586 289338 102822 289574
rect 102266 252458 102502 252694
rect 102586 252458 102822 252694
rect 102266 252138 102502 252374
rect 102586 252138 102822 252374
rect 102266 215258 102502 215494
rect 102586 215258 102822 215494
rect 102266 214938 102502 215174
rect 102586 214938 102822 215174
rect 102266 178058 102502 178294
rect 102586 178058 102822 178294
rect 102266 177738 102502 177974
rect 102586 177738 102822 177974
rect 102266 140858 102502 141094
rect 102586 140858 102822 141094
rect 102266 140538 102502 140774
rect 102586 140538 102822 140774
rect 102266 103658 102502 103894
rect 102586 103658 102822 103894
rect 102266 103338 102502 103574
rect 102586 103338 102822 103574
rect 102266 66458 102502 66694
rect 102586 66458 102822 66694
rect 102266 66138 102502 66374
rect 102586 66138 102822 66374
rect 102266 29258 102502 29494
rect 102586 29258 102822 29494
rect 102266 28938 102502 29174
rect 102586 28938 102822 29174
rect 113426 672818 113662 673054
rect 113746 672818 113982 673054
rect 113426 672498 113662 672734
rect 113746 672498 113982 672734
rect 113426 635618 113662 635854
rect 113746 635618 113982 635854
rect 113426 635298 113662 635534
rect 113746 635298 113982 635534
rect 113426 598418 113662 598654
rect 113746 598418 113982 598654
rect 113426 598098 113662 598334
rect 113746 598098 113982 598334
rect 113426 561218 113662 561454
rect 113746 561218 113982 561454
rect 113426 560898 113662 561134
rect 113746 560898 113982 561134
rect 113426 524018 113662 524254
rect 113746 524018 113982 524254
rect 113426 523698 113662 523934
rect 113746 523698 113982 523934
rect 113426 486818 113662 487054
rect 113746 486818 113982 487054
rect 113426 486498 113662 486734
rect 113746 486498 113982 486734
rect 113426 449618 113662 449854
rect 113746 449618 113982 449854
rect 113426 449298 113662 449534
rect 113746 449298 113982 449534
rect 113426 412418 113662 412654
rect 113746 412418 113982 412654
rect 113426 412098 113662 412334
rect 113746 412098 113982 412334
rect 113426 375218 113662 375454
rect 113746 375218 113982 375454
rect 113426 374898 113662 375134
rect 113746 374898 113982 375134
rect 113426 338018 113662 338254
rect 113746 338018 113982 338254
rect 113426 337698 113662 337934
rect 113746 337698 113982 337934
rect 113426 300818 113662 301054
rect 113746 300818 113982 301054
rect 113426 300498 113662 300734
rect 113746 300498 113982 300734
rect 113426 263618 113662 263854
rect 113746 263618 113982 263854
rect 113426 263298 113662 263534
rect 113746 263298 113982 263534
rect 113426 226418 113662 226654
rect 113746 226418 113982 226654
rect 113426 226098 113662 226334
rect 113746 226098 113982 226334
rect 113426 189218 113662 189454
rect 113746 189218 113982 189454
rect 113426 188898 113662 189134
rect 113746 188898 113982 189134
rect 113426 152018 113662 152254
rect 113746 152018 113982 152254
rect 113426 151698 113662 151934
rect 113746 151698 113982 151934
rect 113426 114818 113662 115054
rect 113746 114818 113982 115054
rect 113426 114498 113662 114734
rect 113746 114498 113982 114734
rect 113426 77618 113662 77854
rect 113746 77618 113982 77854
rect 113426 77298 113662 77534
rect 113746 77298 113982 77534
rect 113426 40418 113662 40654
rect 113746 40418 113982 40654
rect 113426 40098 113662 40334
rect 113746 40098 113982 40334
rect 113426 3218 113662 3454
rect 113746 3218 113982 3454
rect 113426 2898 113662 3134
rect 113746 2898 113982 3134
rect 117146 676538 117382 676774
rect 117466 676538 117702 676774
rect 117146 676218 117382 676454
rect 117466 676218 117702 676454
rect 117146 639338 117382 639574
rect 117466 639338 117702 639574
rect 117146 639018 117382 639254
rect 117466 639018 117702 639254
rect 117146 602138 117382 602374
rect 117466 602138 117702 602374
rect 117146 601818 117382 602054
rect 117466 601818 117702 602054
rect 117146 564938 117382 565174
rect 117466 564938 117702 565174
rect 117146 564618 117382 564854
rect 117466 564618 117702 564854
rect 117146 527738 117382 527974
rect 117466 527738 117702 527974
rect 117146 527418 117382 527654
rect 117466 527418 117702 527654
rect 117146 490538 117382 490774
rect 117466 490538 117702 490774
rect 117146 490218 117382 490454
rect 117466 490218 117702 490454
rect 117146 453338 117382 453574
rect 117466 453338 117702 453574
rect 117146 453018 117382 453254
rect 117466 453018 117702 453254
rect 117146 416138 117382 416374
rect 117466 416138 117702 416374
rect 117146 415818 117382 416054
rect 117466 415818 117702 416054
rect 117146 378938 117382 379174
rect 117466 378938 117702 379174
rect 117146 378618 117382 378854
rect 117466 378618 117702 378854
rect 117146 341738 117382 341974
rect 117466 341738 117702 341974
rect 117146 341418 117382 341654
rect 117466 341418 117702 341654
rect 117146 304538 117382 304774
rect 117466 304538 117702 304774
rect 117146 304218 117382 304454
rect 117466 304218 117702 304454
rect 117146 267338 117382 267574
rect 117466 267338 117702 267574
rect 117146 267018 117382 267254
rect 117466 267018 117702 267254
rect 117146 230138 117382 230374
rect 117466 230138 117702 230374
rect 117146 229818 117382 230054
rect 117466 229818 117702 230054
rect 117146 192938 117382 193174
rect 117466 192938 117702 193174
rect 117146 192618 117382 192854
rect 117466 192618 117702 192854
rect 117146 155738 117382 155974
rect 117466 155738 117702 155974
rect 117146 155418 117382 155654
rect 117466 155418 117702 155654
rect 117146 118538 117382 118774
rect 117466 118538 117702 118774
rect 117146 118218 117382 118454
rect 117466 118218 117702 118454
rect 117146 81338 117382 81574
rect 117466 81338 117702 81574
rect 117146 81018 117382 81254
rect 117466 81018 117702 81254
rect 117146 44138 117382 44374
rect 117466 44138 117702 44374
rect 117146 43818 117382 44054
rect 117466 43818 117702 44054
rect 117146 6938 117382 7174
rect 117466 6938 117702 7174
rect 117146 6618 117382 6854
rect 117466 6618 117702 6854
rect 120866 680258 121102 680494
rect 121186 680258 121422 680494
rect 120866 679938 121102 680174
rect 121186 679938 121422 680174
rect 120866 643058 121102 643294
rect 121186 643058 121422 643294
rect 120866 642738 121102 642974
rect 121186 642738 121422 642974
rect 120866 605858 121102 606094
rect 121186 605858 121422 606094
rect 120866 605538 121102 605774
rect 121186 605538 121422 605774
rect 120866 568658 121102 568894
rect 121186 568658 121422 568894
rect 120866 568338 121102 568574
rect 121186 568338 121422 568574
rect 120866 531458 121102 531694
rect 121186 531458 121422 531694
rect 120866 531138 121102 531374
rect 121186 531138 121422 531374
rect 120866 494258 121102 494494
rect 121186 494258 121422 494494
rect 120866 493938 121102 494174
rect 121186 493938 121422 494174
rect 120866 457058 121102 457294
rect 121186 457058 121422 457294
rect 120866 456738 121102 456974
rect 121186 456738 121422 456974
rect 120866 419858 121102 420094
rect 121186 419858 121422 420094
rect 120866 419538 121102 419774
rect 121186 419538 121422 419774
rect 120866 382658 121102 382894
rect 121186 382658 121422 382894
rect 120866 382338 121102 382574
rect 121186 382338 121422 382574
rect 120866 345458 121102 345694
rect 121186 345458 121422 345694
rect 120866 345138 121102 345374
rect 121186 345138 121422 345374
rect 120866 308258 121102 308494
rect 121186 308258 121422 308494
rect 120866 307938 121102 308174
rect 121186 307938 121422 308174
rect 120866 271058 121102 271294
rect 121186 271058 121422 271294
rect 120866 270738 121102 270974
rect 121186 270738 121422 270974
rect 120866 233858 121102 234094
rect 121186 233858 121422 234094
rect 120866 233538 121102 233774
rect 121186 233538 121422 233774
rect 120866 196658 121102 196894
rect 121186 196658 121422 196894
rect 120866 196338 121102 196574
rect 121186 196338 121422 196574
rect 120866 159458 121102 159694
rect 121186 159458 121422 159694
rect 120866 159138 121102 159374
rect 121186 159138 121422 159374
rect 120866 122258 121102 122494
rect 121186 122258 121422 122494
rect 120866 121938 121102 122174
rect 121186 121938 121422 122174
rect 120866 85058 121102 85294
rect 121186 85058 121422 85294
rect 120866 84738 121102 84974
rect 121186 84738 121422 84974
rect 120866 47858 121102 48094
rect 121186 47858 121422 48094
rect 120866 47538 121102 47774
rect 121186 47538 121422 47774
rect 120866 10658 121102 10894
rect 121186 10658 121422 10894
rect 120866 10338 121102 10574
rect 121186 10338 121422 10574
rect 124586 683978 124822 684214
rect 124906 683978 125142 684214
rect 124586 683658 124822 683894
rect 124906 683658 125142 683894
rect 124586 646778 124822 647014
rect 124906 646778 125142 647014
rect 124586 646458 124822 646694
rect 124906 646458 125142 646694
rect 124586 609578 124822 609814
rect 124906 609578 125142 609814
rect 124586 609258 124822 609494
rect 124906 609258 125142 609494
rect 124586 572378 124822 572614
rect 124906 572378 125142 572614
rect 124586 572058 124822 572294
rect 124906 572058 125142 572294
rect 124586 535178 124822 535414
rect 124906 535178 125142 535414
rect 124586 534858 124822 535094
rect 124906 534858 125142 535094
rect 124586 497978 124822 498214
rect 124906 497978 125142 498214
rect 124586 497658 124822 497894
rect 124906 497658 125142 497894
rect 124586 460778 124822 461014
rect 124906 460778 125142 461014
rect 124586 460458 124822 460694
rect 124906 460458 125142 460694
rect 124586 423578 124822 423814
rect 124906 423578 125142 423814
rect 124586 423258 124822 423494
rect 124906 423258 125142 423494
rect 124586 386378 124822 386614
rect 124906 386378 125142 386614
rect 124586 386058 124822 386294
rect 124906 386058 125142 386294
rect 124586 349178 124822 349414
rect 124906 349178 125142 349414
rect 124586 348858 124822 349094
rect 124906 348858 125142 349094
rect 124586 311978 124822 312214
rect 124906 311978 125142 312214
rect 124586 311658 124822 311894
rect 124906 311658 125142 311894
rect 124586 274778 124822 275014
rect 124906 274778 125142 275014
rect 124586 274458 124822 274694
rect 124906 274458 125142 274694
rect 124586 237578 124822 237814
rect 124906 237578 125142 237814
rect 124586 237258 124822 237494
rect 124906 237258 125142 237494
rect 124586 200378 124822 200614
rect 124906 200378 125142 200614
rect 124586 200058 124822 200294
rect 124906 200058 125142 200294
rect 124586 163178 124822 163414
rect 124906 163178 125142 163414
rect 124586 162858 124822 163094
rect 124906 162858 125142 163094
rect 124586 125978 124822 126214
rect 124906 125978 125142 126214
rect 124586 125658 124822 125894
rect 124906 125658 125142 125894
rect 124586 88778 124822 89014
rect 124906 88778 125142 89014
rect 124586 88458 124822 88694
rect 124906 88458 125142 88694
rect 124586 51578 124822 51814
rect 124906 51578 125142 51814
rect 124586 51258 124822 51494
rect 124906 51258 125142 51494
rect 124586 14378 124822 14614
rect 124906 14378 125142 14614
rect 124586 14058 124822 14294
rect 124906 14058 125142 14294
rect 128306 687698 128542 687934
rect 128626 687698 128862 687934
rect 128306 687378 128542 687614
rect 128626 687378 128862 687614
rect 128306 650498 128542 650734
rect 128626 650498 128862 650734
rect 128306 650178 128542 650414
rect 128626 650178 128862 650414
rect 128306 613298 128542 613534
rect 128626 613298 128862 613534
rect 128306 612978 128542 613214
rect 128626 612978 128862 613214
rect 128306 576098 128542 576334
rect 128626 576098 128862 576334
rect 128306 575778 128542 576014
rect 128626 575778 128862 576014
rect 128306 538898 128542 539134
rect 128626 538898 128862 539134
rect 128306 538578 128542 538814
rect 128626 538578 128862 538814
rect 128306 501698 128542 501934
rect 128626 501698 128862 501934
rect 128306 501378 128542 501614
rect 128626 501378 128862 501614
rect 128306 464498 128542 464734
rect 128626 464498 128862 464734
rect 128306 464178 128542 464414
rect 128626 464178 128862 464414
rect 128306 427298 128542 427534
rect 128626 427298 128862 427534
rect 128306 426978 128542 427214
rect 128626 426978 128862 427214
rect 128306 390098 128542 390334
rect 128626 390098 128862 390334
rect 128306 389778 128542 390014
rect 128626 389778 128862 390014
rect 128306 352898 128542 353134
rect 128626 352898 128862 353134
rect 128306 352578 128542 352814
rect 128626 352578 128862 352814
rect 128306 315698 128542 315934
rect 128626 315698 128862 315934
rect 128306 315378 128542 315614
rect 128626 315378 128862 315614
rect 128306 278498 128542 278734
rect 128626 278498 128862 278734
rect 128306 278178 128542 278414
rect 128626 278178 128862 278414
rect 128306 241298 128542 241534
rect 128626 241298 128862 241534
rect 128306 240978 128542 241214
rect 128626 240978 128862 241214
rect 128306 204098 128542 204334
rect 128626 204098 128862 204334
rect 128306 203778 128542 204014
rect 128626 203778 128862 204014
rect 128306 166898 128542 167134
rect 128626 166898 128862 167134
rect 128306 166578 128542 166814
rect 128626 166578 128862 166814
rect 128306 129698 128542 129934
rect 128626 129698 128862 129934
rect 128306 129378 128542 129614
rect 128626 129378 128862 129614
rect 128306 92498 128542 92734
rect 128626 92498 128862 92734
rect 128306 92178 128542 92414
rect 128626 92178 128862 92414
rect 128306 55298 128542 55534
rect 128626 55298 128862 55534
rect 128306 54978 128542 55214
rect 128626 54978 128862 55214
rect 128306 18098 128542 18334
rect 128626 18098 128862 18334
rect 128306 17778 128542 18014
rect 128626 17778 128862 18014
rect 132026 691418 132262 691654
rect 132346 691418 132582 691654
rect 132026 691098 132262 691334
rect 132346 691098 132582 691334
rect 132026 654218 132262 654454
rect 132346 654218 132582 654454
rect 132026 653898 132262 654134
rect 132346 653898 132582 654134
rect 132026 617018 132262 617254
rect 132346 617018 132582 617254
rect 132026 616698 132262 616934
rect 132346 616698 132582 616934
rect 132026 579818 132262 580054
rect 132346 579818 132582 580054
rect 132026 579498 132262 579734
rect 132346 579498 132582 579734
rect 132026 542618 132262 542854
rect 132346 542618 132582 542854
rect 132026 542298 132262 542534
rect 132346 542298 132582 542534
rect 132026 505418 132262 505654
rect 132346 505418 132582 505654
rect 132026 505098 132262 505334
rect 132346 505098 132582 505334
rect 132026 468218 132262 468454
rect 132346 468218 132582 468454
rect 132026 467898 132262 468134
rect 132346 467898 132582 468134
rect 132026 431018 132262 431254
rect 132346 431018 132582 431254
rect 132026 430698 132262 430934
rect 132346 430698 132582 430934
rect 132026 393818 132262 394054
rect 132346 393818 132582 394054
rect 132026 393498 132262 393734
rect 132346 393498 132582 393734
rect 132026 356618 132262 356854
rect 132346 356618 132582 356854
rect 132026 356298 132262 356534
rect 132346 356298 132582 356534
rect 132026 319418 132262 319654
rect 132346 319418 132582 319654
rect 132026 319098 132262 319334
rect 132346 319098 132582 319334
rect 132026 282218 132262 282454
rect 132346 282218 132582 282454
rect 132026 281898 132262 282134
rect 132346 281898 132582 282134
rect 132026 245018 132262 245254
rect 132346 245018 132582 245254
rect 132026 244698 132262 244934
rect 132346 244698 132582 244934
rect 132026 207818 132262 208054
rect 132346 207818 132582 208054
rect 132026 207498 132262 207734
rect 132346 207498 132582 207734
rect 132026 170618 132262 170854
rect 132346 170618 132582 170854
rect 132026 170298 132262 170534
rect 132346 170298 132582 170534
rect 132026 133418 132262 133654
rect 132346 133418 132582 133654
rect 132026 133098 132262 133334
rect 132346 133098 132582 133334
rect 132026 96218 132262 96454
rect 132346 96218 132582 96454
rect 132026 95898 132262 96134
rect 132346 95898 132582 96134
rect 132026 59018 132262 59254
rect 132346 59018 132582 59254
rect 132026 58698 132262 58934
rect 132346 58698 132582 58934
rect 132026 21818 132262 22054
rect 132346 21818 132582 22054
rect 132026 21498 132262 21734
rect 132346 21498 132582 21734
rect 135746 695138 135982 695374
rect 136066 695138 136302 695374
rect 135746 694818 135982 695054
rect 136066 694818 136302 695054
rect 135746 657938 135982 658174
rect 136066 657938 136302 658174
rect 135746 657618 135982 657854
rect 136066 657618 136302 657854
rect 135746 620738 135982 620974
rect 136066 620738 136302 620974
rect 135746 620418 135982 620654
rect 136066 620418 136302 620654
rect 135746 583538 135982 583774
rect 136066 583538 136302 583774
rect 135746 583218 135982 583454
rect 136066 583218 136302 583454
rect 135746 546338 135982 546574
rect 136066 546338 136302 546574
rect 135746 546018 135982 546254
rect 136066 546018 136302 546254
rect 135746 509138 135982 509374
rect 136066 509138 136302 509374
rect 135746 508818 135982 509054
rect 136066 508818 136302 509054
rect 135746 471938 135982 472174
rect 136066 471938 136302 472174
rect 135746 471618 135982 471854
rect 136066 471618 136302 471854
rect 135746 434738 135982 434974
rect 136066 434738 136302 434974
rect 135746 434418 135982 434654
rect 136066 434418 136302 434654
rect 135746 397538 135982 397774
rect 136066 397538 136302 397774
rect 135746 397218 135982 397454
rect 136066 397218 136302 397454
rect 135746 360338 135982 360574
rect 136066 360338 136302 360574
rect 135746 360018 135982 360254
rect 136066 360018 136302 360254
rect 135746 323138 135982 323374
rect 136066 323138 136302 323374
rect 135746 322818 135982 323054
rect 136066 322818 136302 323054
rect 135746 285938 135982 286174
rect 136066 285938 136302 286174
rect 135746 285618 135982 285854
rect 136066 285618 136302 285854
rect 135746 248738 135982 248974
rect 136066 248738 136302 248974
rect 135746 248418 135982 248654
rect 136066 248418 136302 248654
rect 135746 211538 135982 211774
rect 136066 211538 136302 211774
rect 135746 211218 135982 211454
rect 136066 211218 136302 211454
rect 135746 174338 135982 174574
rect 136066 174338 136302 174574
rect 135746 174018 135982 174254
rect 136066 174018 136302 174254
rect 135746 137138 135982 137374
rect 136066 137138 136302 137374
rect 135746 136818 135982 137054
rect 136066 136818 136302 137054
rect 135746 99938 135982 100174
rect 136066 99938 136302 100174
rect 135746 99618 135982 99854
rect 136066 99618 136302 99854
rect 135746 62738 135982 62974
rect 136066 62738 136302 62974
rect 135746 62418 135982 62654
rect 136066 62418 136302 62654
rect 135746 25538 135982 25774
rect 136066 25538 136302 25774
rect 135746 25218 135982 25454
rect 136066 25218 136302 25454
rect 139466 698858 139702 699094
rect 139786 698858 140022 699094
rect 139466 698538 139702 698774
rect 139786 698538 140022 698774
rect 139466 661658 139702 661894
rect 139786 661658 140022 661894
rect 139466 661338 139702 661574
rect 139786 661338 140022 661574
rect 139466 624458 139702 624694
rect 139786 624458 140022 624694
rect 139466 624138 139702 624374
rect 139786 624138 140022 624374
rect 139466 587258 139702 587494
rect 139786 587258 140022 587494
rect 139466 586938 139702 587174
rect 139786 586938 140022 587174
rect 139466 550058 139702 550294
rect 139786 550058 140022 550294
rect 139466 549738 139702 549974
rect 139786 549738 140022 549974
rect 139466 512858 139702 513094
rect 139786 512858 140022 513094
rect 139466 512538 139702 512774
rect 139786 512538 140022 512774
rect 139466 475658 139702 475894
rect 139786 475658 140022 475894
rect 139466 475338 139702 475574
rect 139786 475338 140022 475574
rect 139466 438458 139702 438694
rect 139786 438458 140022 438694
rect 139466 438138 139702 438374
rect 139786 438138 140022 438374
rect 139466 401258 139702 401494
rect 139786 401258 140022 401494
rect 139466 400938 139702 401174
rect 139786 400938 140022 401174
rect 139466 364058 139702 364294
rect 139786 364058 140022 364294
rect 139466 363738 139702 363974
rect 139786 363738 140022 363974
rect 139466 326858 139702 327094
rect 139786 326858 140022 327094
rect 139466 326538 139702 326774
rect 139786 326538 140022 326774
rect 139466 289658 139702 289894
rect 139786 289658 140022 289894
rect 139466 289338 139702 289574
rect 139786 289338 140022 289574
rect 139466 252458 139702 252694
rect 139786 252458 140022 252694
rect 139466 252138 139702 252374
rect 139786 252138 140022 252374
rect 139466 215258 139702 215494
rect 139786 215258 140022 215494
rect 139466 214938 139702 215174
rect 139786 214938 140022 215174
rect 139466 178058 139702 178294
rect 139786 178058 140022 178294
rect 139466 177738 139702 177974
rect 139786 177738 140022 177974
rect 139466 140858 139702 141094
rect 139786 140858 140022 141094
rect 139466 140538 139702 140774
rect 139786 140538 140022 140774
rect 139466 103658 139702 103894
rect 139786 103658 140022 103894
rect 139466 103338 139702 103574
rect 139786 103338 140022 103574
rect 139466 66458 139702 66694
rect 139786 66458 140022 66694
rect 139466 66138 139702 66374
rect 139786 66138 140022 66374
rect 139466 29258 139702 29494
rect 139786 29258 140022 29494
rect 139466 28938 139702 29174
rect 139786 28938 140022 29174
rect 150626 672818 150862 673054
rect 150946 672818 151182 673054
rect 150626 672498 150862 672734
rect 150946 672498 151182 672734
rect 150626 635618 150862 635854
rect 150946 635618 151182 635854
rect 150626 635298 150862 635534
rect 150946 635298 151182 635534
rect 150626 598418 150862 598654
rect 150946 598418 151182 598654
rect 150626 598098 150862 598334
rect 150946 598098 151182 598334
rect 150626 561218 150862 561454
rect 150946 561218 151182 561454
rect 150626 560898 150862 561134
rect 150946 560898 151182 561134
rect 150626 524018 150862 524254
rect 150946 524018 151182 524254
rect 150626 523698 150862 523934
rect 150946 523698 151182 523934
rect 150626 486818 150862 487054
rect 150946 486818 151182 487054
rect 150626 486498 150862 486734
rect 150946 486498 151182 486734
rect 150626 449618 150862 449854
rect 150946 449618 151182 449854
rect 150626 449298 150862 449534
rect 150946 449298 151182 449534
rect 150626 412418 150862 412654
rect 150946 412418 151182 412654
rect 150626 412098 150862 412334
rect 150946 412098 151182 412334
rect 150626 375218 150862 375454
rect 150946 375218 151182 375454
rect 150626 374898 150862 375134
rect 150946 374898 151182 375134
rect 150626 338018 150862 338254
rect 150946 338018 151182 338254
rect 150626 337698 150862 337934
rect 150946 337698 151182 337934
rect 150626 300818 150862 301054
rect 150946 300818 151182 301054
rect 150626 300498 150862 300734
rect 150946 300498 151182 300734
rect 150626 263618 150862 263854
rect 150946 263618 151182 263854
rect 150626 263298 150862 263534
rect 150946 263298 151182 263534
rect 150626 226418 150862 226654
rect 150946 226418 151182 226654
rect 150626 226098 150862 226334
rect 150946 226098 151182 226334
rect 150626 189218 150862 189454
rect 150946 189218 151182 189454
rect 150626 188898 150862 189134
rect 150946 188898 151182 189134
rect 150626 152018 150862 152254
rect 150946 152018 151182 152254
rect 150626 151698 150862 151934
rect 150946 151698 151182 151934
rect 150626 114818 150862 115054
rect 150946 114818 151182 115054
rect 150626 114498 150862 114734
rect 150946 114498 151182 114734
rect 150626 77618 150862 77854
rect 150946 77618 151182 77854
rect 150626 77298 150862 77534
rect 150946 77298 151182 77534
rect 150626 40418 150862 40654
rect 150946 40418 151182 40654
rect 150626 40098 150862 40334
rect 150946 40098 151182 40334
rect 150626 3218 150862 3454
rect 150946 3218 151182 3454
rect 150626 2898 150862 3134
rect 150946 2898 151182 3134
rect 154346 676538 154582 676774
rect 154666 676538 154902 676774
rect 154346 676218 154582 676454
rect 154666 676218 154902 676454
rect 154346 639338 154582 639574
rect 154666 639338 154902 639574
rect 154346 639018 154582 639254
rect 154666 639018 154902 639254
rect 154346 602138 154582 602374
rect 154666 602138 154902 602374
rect 154346 601818 154582 602054
rect 154666 601818 154902 602054
rect 154346 564938 154582 565174
rect 154666 564938 154902 565174
rect 154346 564618 154582 564854
rect 154666 564618 154902 564854
rect 154346 527738 154582 527974
rect 154666 527738 154902 527974
rect 154346 527418 154582 527654
rect 154666 527418 154902 527654
rect 154346 490538 154582 490774
rect 154666 490538 154902 490774
rect 154346 490218 154582 490454
rect 154666 490218 154902 490454
rect 154346 453338 154582 453574
rect 154666 453338 154902 453574
rect 154346 453018 154582 453254
rect 154666 453018 154902 453254
rect 154346 416138 154582 416374
rect 154666 416138 154902 416374
rect 154346 415818 154582 416054
rect 154666 415818 154902 416054
rect 154346 378938 154582 379174
rect 154666 378938 154902 379174
rect 154346 378618 154582 378854
rect 154666 378618 154902 378854
rect 154346 341738 154582 341974
rect 154666 341738 154902 341974
rect 154346 341418 154582 341654
rect 154666 341418 154902 341654
rect 154346 304538 154582 304774
rect 154666 304538 154902 304774
rect 154346 304218 154582 304454
rect 154666 304218 154902 304454
rect 154346 267338 154582 267574
rect 154666 267338 154902 267574
rect 154346 267018 154582 267254
rect 154666 267018 154902 267254
rect 154346 230138 154582 230374
rect 154666 230138 154902 230374
rect 154346 229818 154582 230054
rect 154666 229818 154902 230054
rect 154346 192938 154582 193174
rect 154666 192938 154902 193174
rect 154346 192618 154582 192854
rect 154666 192618 154902 192854
rect 154346 155738 154582 155974
rect 154666 155738 154902 155974
rect 154346 155418 154582 155654
rect 154666 155418 154902 155654
rect 154346 118538 154582 118774
rect 154666 118538 154902 118774
rect 154346 118218 154582 118454
rect 154666 118218 154902 118454
rect 154346 81338 154582 81574
rect 154666 81338 154902 81574
rect 154346 81018 154582 81254
rect 154666 81018 154902 81254
rect 154346 44138 154582 44374
rect 154666 44138 154902 44374
rect 154346 43818 154582 44054
rect 154666 43818 154902 44054
rect 154346 6938 154582 7174
rect 154666 6938 154902 7174
rect 154346 6618 154582 6854
rect 154666 6618 154902 6854
rect 158066 680258 158302 680494
rect 158386 680258 158622 680494
rect 158066 679938 158302 680174
rect 158386 679938 158622 680174
rect 158066 643058 158302 643294
rect 158386 643058 158622 643294
rect 158066 642738 158302 642974
rect 158386 642738 158622 642974
rect 158066 605858 158302 606094
rect 158386 605858 158622 606094
rect 158066 605538 158302 605774
rect 158386 605538 158622 605774
rect 158066 568658 158302 568894
rect 158386 568658 158622 568894
rect 158066 568338 158302 568574
rect 158386 568338 158622 568574
rect 158066 531458 158302 531694
rect 158386 531458 158622 531694
rect 158066 531138 158302 531374
rect 158386 531138 158622 531374
rect 158066 494258 158302 494494
rect 158386 494258 158622 494494
rect 158066 493938 158302 494174
rect 158386 493938 158622 494174
rect 158066 457058 158302 457294
rect 158386 457058 158622 457294
rect 158066 456738 158302 456974
rect 158386 456738 158622 456974
rect 158066 419858 158302 420094
rect 158386 419858 158622 420094
rect 158066 419538 158302 419774
rect 158386 419538 158622 419774
rect 158066 382658 158302 382894
rect 158386 382658 158622 382894
rect 158066 382338 158302 382574
rect 158386 382338 158622 382574
rect 158066 345458 158302 345694
rect 158386 345458 158622 345694
rect 158066 345138 158302 345374
rect 158386 345138 158622 345374
rect 158066 308258 158302 308494
rect 158386 308258 158622 308494
rect 158066 307938 158302 308174
rect 158386 307938 158622 308174
rect 158066 271058 158302 271294
rect 158386 271058 158622 271294
rect 158066 270738 158302 270974
rect 158386 270738 158622 270974
rect 158066 233858 158302 234094
rect 158386 233858 158622 234094
rect 158066 233538 158302 233774
rect 158386 233538 158622 233774
rect 158066 196658 158302 196894
rect 158386 196658 158622 196894
rect 158066 196338 158302 196574
rect 158386 196338 158622 196574
rect 158066 159458 158302 159694
rect 158386 159458 158622 159694
rect 158066 159138 158302 159374
rect 158386 159138 158622 159374
rect 158066 122258 158302 122494
rect 158386 122258 158622 122494
rect 158066 121938 158302 122174
rect 158386 121938 158622 122174
rect 158066 85058 158302 85294
rect 158386 85058 158622 85294
rect 158066 84738 158302 84974
rect 158386 84738 158622 84974
rect 158066 47858 158302 48094
rect 158386 47858 158622 48094
rect 158066 47538 158302 47774
rect 158386 47538 158622 47774
rect 158066 10658 158302 10894
rect 158386 10658 158622 10894
rect 158066 10338 158302 10574
rect 158386 10338 158622 10574
rect 161786 683978 162022 684214
rect 162106 683978 162342 684214
rect 161786 683658 162022 683894
rect 162106 683658 162342 683894
rect 161786 646778 162022 647014
rect 162106 646778 162342 647014
rect 161786 646458 162022 646694
rect 162106 646458 162342 646694
rect 161786 609578 162022 609814
rect 162106 609578 162342 609814
rect 161786 609258 162022 609494
rect 162106 609258 162342 609494
rect 161786 572378 162022 572614
rect 162106 572378 162342 572614
rect 161786 572058 162022 572294
rect 162106 572058 162342 572294
rect 161786 535178 162022 535414
rect 162106 535178 162342 535414
rect 161786 534858 162022 535094
rect 162106 534858 162342 535094
rect 161786 497978 162022 498214
rect 162106 497978 162342 498214
rect 161786 497658 162022 497894
rect 162106 497658 162342 497894
rect 161786 460778 162022 461014
rect 162106 460778 162342 461014
rect 161786 460458 162022 460694
rect 162106 460458 162342 460694
rect 161786 423578 162022 423814
rect 162106 423578 162342 423814
rect 161786 423258 162022 423494
rect 162106 423258 162342 423494
rect 161786 386378 162022 386614
rect 162106 386378 162342 386614
rect 161786 386058 162022 386294
rect 162106 386058 162342 386294
rect 161786 349178 162022 349414
rect 162106 349178 162342 349414
rect 161786 348858 162022 349094
rect 162106 348858 162342 349094
rect 161786 311978 162022 312214
rect 162106 311978 162342 312214
rect 161786 311658 162022 311894
rect 162106 311658 162342 311894
rect 161786 274778 162022 275014
rect 162106 274778 162342 275014
rect 161786 274458 162022 274694
rect 162106 274458 162342 274694
rect 161786 237578 162022 237814
rect 162106 237578 162342 237814
rect 161786 237258 162022 237494
rect 162106 237258 162342 237494
rect 161786 200378 162022 200614
rect 162106 200378 162342 200614
rect 161786 200058 162022 200294
rect 162106 200058 162342 200294
rect 161786 163178 162022 163414
rect 162106 163178 162342 163414
rect 161786 162858 162022 163094
rect 162106 162858 162342 163094
rect 161786 125978 162022 126214
rect 162106 125978 162342 126214
rect 161786 125658 162022 125894
rect 162106 125658 162342 125894
rect 161786 88778 162022 89014
rect 162106 88778 162342 89014
rect 161786 88458 162022 88694
rect 162106 88458 162342 88694
rect 161786 51578 162022 51814
rect 162106 51578 162342 51814
rect 161786 51258 162022 51494
rect 162106 51258 162342 51494
rect 161786 14378 162022 14614
rect 162106 14378 162342 14614
rect 161786 14058 162022 14294
rect 162106 14058 162342 14294
rect 165506 687698 165742 687934
rect 165826 687698 166062 687934
rect 165506 687378 165742 687614
rect 165826 687378 166062 687614
rect 165506 650498 165742 650734
rect 165826 650498 166062 650734
rect 165506 650178 165742 650414
rect 165826 650178 166062 650414
rect 165506 613298 165742 613534
rect 165826 613298 166062 613534
rect 165506 612978 165742 613214
rect 165826 612978 166062 613214
rect 165506 576098 165742 576334
rect 165826 576098 166062 576334
rect 165506 575778 165742 576014
rect 165826 575778 166062 576014
rect 165506 538898 165742 539134
rect 165826 538898 166062 539134
rect 165506 538578 165742 538814
rect 165826 538578 166062 538814
rect 165506 501698 165742 501934
rect 165826 501698 166062 501934
rect 165506 501378 165742 501614
rect 165826 501378 166062 501614
rect 165506 464498 165742 464734
rect 165826 464498 166062 464734
rect 165506 464178 165742 464414
rect 165826 464178 166062 464414
rect 165506 427298 165742 427534
rect 165826 427298 166062 427534
rect 165506 426978 165742 427214
rect 165826 426978 166062 427214
rect 165506 390098 165742 390334
rect 165826 390098 166062 390334
rect 165506 389778 165742 390014
rect 165826 389778 166062 390014
rect 165506 352898 165742 353134
rect 165826 352898 166062 353134
rect 165506 352578 165742 352814
rect 165826 352578 166062 352814
rect 165506 315698 165742 315934
rect 165826 315698 166062 315934
rect 165506 315378 165742 315614
rect 165826 315378 166062 315614
rect 165506 278498 165742 278734
rect 165826 278498 166062 278734
rect 165506 278178 165742 278414
rect 165826 278178 166062 278414
rect 165506 241298 165742 241534
rect 165826 241298 166062 241534
rect 165506 240978 165742 241214
rect 165826 240978 166062 241214
rect 165506 204098 165742 204334
rect 165826 204098 166062 204334
rect 165506 203778 165742 204014
rect 165826 203778 166062 204014
rect 165506 166898 165742 167134
rect 165826 166898 166062 167134
rect 165506 166578 165742 166814
rect 165826 166578 166062 166814
rect 165506 129698 165742 129934
rect 165826 129698 166062 129934
rect 165506 129378 165742 129614
rect 165826 129378 166062 129614
rect 165506 92498 165742 92734
rect 165826 92498 166062 92734
rect 165506 92178 165742 92414
rect 165826 92178 166062 92414
rect 165506 55298 165742 55534
rect 165826 55298 166062 55534
rect 165506 54978 165742 55214
rect 165826 54978 166062 55214
rect 165506 18098 165742 18334
rect 165826 18098 166062 18334
rect 165506 17778 165742 18014
rect 165826 17778 166062 18014
rect 169226 691418 169462 691654
rect 169546 691418 169782 691654
rect 169226 691098 169462 691334
rect 169546 691098 169782 691334
rect 169226 654218 169462 654454
rect 169546 654218 169782 654454
rect 169226 653898 169462 654134
rect 169546 653898 169782 654134
rect 169226 617018 169462 617254
rect 169546 617018 169782 617254
rect 169226 616698 169462 616934
rect 169546 616698 169782 616934
rect 169226 579818 169462 580054
rect 169546 579818 169782 580054
rect 169226 579498 169462 579734
rect 169546 579498 169782 579734
rect 169226 542618 169462 542854
rect 169546 542618 169782 542854
rect 169226 542298 169462 542534
rect 169546 542298 169782 542534
rect 169226 505418 169462 505654
rect 169546 505418 169782 505654
rect 169226 505098 169462 505334
rect 169546 505098 169782 505334
rect 169226 468218 169462 468454
rect 169546 468218 169782 468454
rect 169226 467898 169462 468134
rect 169546 467898 169782 468134
rect 169226 431018 169462 431254
rect 169546 431018 169782 431254
rect 169226 430698 169462 430934
rect 169546 430698 169782 430934
rect 169226 393818 169462 394054
rect 169546 393818 169782 394054
rect 169226 393498 169462 393734
rect 169546 393498 169782 393734
rect 169226 356618 169462 356854
rect 169546 356618 169782 356854
rect 169226 356298 169462 356534
rect 169546 356298 169782 356534
rect 169226 319418 169462 319654
rect 169546 319418 169782 319654
rect 169226 319098 169462 319334
rect 169546 319098 169782 319334
rect 169226 282218 169462 282454
rect 169546 282218 169782 282454
rect 169226 281898 169462 282134
rect 169546 281898 169782 282134
rect 169226 245018 169462 245254
rect 169546 245018 169782 245254
rect 169226 244698 169462 244934
rect 169546 244698 169782 244934
rect 169226 207818 169462 208054
rect 169546 207818 169782 208054
rect 169226 207498 169462 207734
rect 169546 207498 169782 207734
rect 169226 170618 169462 170854
rect 169546 170618 169782 170854
rect 169226 170298 169462 170534
rect 169546 170298 169782 170534
rect 169226 133418 169462 133654
rect 169546 133418 169782 133654
rect 169226 133098 169462 133334
rect 169546 133098 169782 133334
rect 169226 96218 169462 96454
rect 169546 96218 169782 96454
rect 169226 95898 169462 96134
rect 169546 95898 169782 96134
rect 169226 59018 169462 59254
rect 169546 59018 169782 59254
rect 169226 58698 169462 58934
rect 169546 58698 169782 58934
rect 169226 21818 169462 22054
rect 169546 21818 169782 22054
rect 169226 21498 169462 21734
rect 169546 21498 169782 21734
rect 172946 695138 173182 695374
rect 173266 695138 173502 695374
rect 172946 694818 173182 695054
rect 173266 694818 173502 695054
rect 172946 657938 173182 658174
rect 173266 657938 173502 658174
rect 172946 657618 173182 657854
rect 173266 657618 173502 657854
rect 172946 620738 173182 620974
rect 173266 620738 173502 620974
rect 172946 620418 173182 620654
rect 173266 620418 173502 620654
rect 172946 583538 173182 583774
rect 173266 583538 173502 583774
rect 172946 583218 173182 583454
rect 173266 583218 173502 583454
rect 172946 546338 173182 546574
rect 173266 546338 173502 546574
rect 172946 546018 173182 546254
rect 173266 546018 173502 546254
rect 172946 509138 173182 509374
rect 173266 509138 173502 509374
rect 172946 508818 173182 509054
rect 173266 508818 173502 509054
rect 172946 471938 173182 472174
rect 173266 471938 173502 472174
rect 172946 471618 173182 471854
rect 173266 471618 173502 471854
rect 172946 434738 173182 434974
rect 173266 434738 173502 434974
rect 172946 434418 173182 434654
rect 173266 434418 173502 434654
rect 172946 397538 173182 397774
rect 173266 397538 173502 397774
rect 172946 397218 173182 397454
rect 173266 397218 173502 397454
rect 172946 360338 173182 360574
rect 173266 360338 173502 360574
rect 172946 360018 173182 360254
rect 173266 360018 173502 360254
rect 172946 323138 173182 323374
rect 173266 323138 173502 323374
rect 172946 322818 173182 323054
rect 173266 322818 173502 323054
rect 172946 285938 173182 286174
rect 173266 285938 173502 286174
rect 172946 285618 173182 285854
rect 173266 285618 173502 285854
rect 172946 248738 173182 248974
rect 173266 248738 173502 248974
rect 172946 248418 173182 248654
rect 173266 248418 173502 248654
rect 172946 211538 173182 211774
rect 173266 211538 173502 211774
rect 172946 211218 173182 211454
rect 173266 211218 173502 211454
rect 172946 174338 173182 174574
rect 173266 174338 173502 174574
rect 172946 174018 173182 174254
rect 173266 174018 173502 174254
rect 172946 137138 173182 137374
rect 173266 137138 173502 137374
rect 172946 136818 173182 137054
rect 173266 136818 173502 137054
rect 172946 99938 173182 100174
rect 173266 99938 173502 100174
rect 172946 99618 173182 99854
rect 173266 99618 173502 99854
rect 172946 62738 173182 62974
rect 173266 62738 173502 62974
rect 172946 62418 173182 62654
rect 173266 62418 173502 62654
rect 172946 25538 173182 25774
rect 173266 25538 173502 25774
rect 172946 25218 173182 25454
rect 173266 25218 173502 25454
rect 176666 698858 176902 699094
rect 176986 698858 177222 699094
rect 176666 698538 176902 698774
rect 176986 698538 177222 698774
rect 176666 661658 176902 661894
rect 176986 661658 177222 661894
rect 176666 661338 176902 661574
rect 176986 661338 177222 661574
rect 176666 624458 176902 624694
rect 176986 624458 177222 624694
rect 176666 624138 176902 624374
rect 176986 624138 177222 624374
rect 176666 587258 176902 587494
rect 176986 587258 177222 587494
rect 176666 586938 176902 587174
rect 176986 586938 177222 587174
rect 176666 550058 176902 550294
rect 176986 550058 177222 550294
rect 176666 549738 176902 549974
rect 176986 549738 177222 549974
rect 176666 512858 176902 513094
rect 176986 512858 177222 513094
rect 176666 512538 176902 512774
rect 176986 512538 177222 512774
rect 176666 475658 176902 475894
rect 176986 475658 177222 475894
rect 176666 475338 176902 475574
rect 176986 475338 177222 475574
rect 176666 438458 176902 438694
rect 176986 438458 177222 438694
rect 176666 438138 176902 438374
rect 176986 438138 177222 438374
rect 176666 401258 176902 401494
rect 176986 401258 177222 401494
rect 176666 400938 176902 401174
rect 176986 400938 177222 401174
rect 176666 364058 176902 364294
rect 176986 364058 177222 364294
rect 176666 363738 176902 363974
rect 176986 363738 177222 363974
rect 176666 326858 176902 327094
rect 176986 326858 177222 327094
rect 176666 326538 176902 326774
rect 176986 326538 177222 326774
rect 176666 289658 176902 289894
rect 176986 289658 177222 289894
rect 176666 289338 176902 289574
rect 176986 289338 177222 289574
rect 176666 252458 176902 252694
rect 176986 252458 177222 252694
rect 176666 252138 176902 252374
rect 176986 252138 177222 252374
rect 176666 215258 176902 215494
rect 176986 215258 177222 215494
rect 176666 214938 176902 215174
rect 176986 214938 177222 215174
rect 176666 178058 176902 178294
rect 176986 178058 177222 178294
rect 176666 177738 176902 177974
rect 176986 177738 177222 177974
rect 176666 140858 176902 141094
rect 176986 140858 177222 141094
rect 176666 140538 176902 140774
rect 176986 140538 177222 140774
rect 176666 103658 176902 103894
rect 176986 103658 177222 103894
rect 176666 103338 176902 103574
rect 176986 103338 177222 103574
rect 176666 66458 176902 66694
rect 176986 66458 177222 66694
rect 176666 66138 176902 66374
rect 176986 66138 177222 66374
rect 176666 29258 176902 29494
rect 176986 29258 177222 29494
rect 176666 28938 176902 29174
rect 176986 28938 177222 29174
rect 187826 672818 188062 673054
rect 188146 672818 188382 673054
rect 187826 672498 188062 672734
rect 188146 672498 188382 672734
rect 187826 635618 188062 635854
rect 188146 635618 188382 635854
rect 187826 635298 188062 635534
rect 188146 635298 188382 635534
rect 187826 598418 188062 598654
rect 188146 598418 188382 598654
rect 187826 598098 188062 598334
rect 188146 598098 188382 598334
rect 187826 561218 188062 561454
rect 188146 561218 188382 561454
rect 187826 560898 188062 561134
rect 188146 560898 188382 561134
rect 187826 524018 188062 524254
rect 188146 524018 188382 524254
rect 187826 523698 188062 523934
rect 188146 523698 188382 523934
rect 187826 486818 188062 487054
rect 188146 486818 188382 487054
rect 187826 486498 188062 486734
rect 188146 486498 188382 486734
rect 187826 449618 188062 449854
rect 188146 449618 188382 449854
rect 187826 449298 188062 449534
rect 188146 449298 188382 449534
rect 187826 412418 188062 412654
rect 188146 412418 188382 412654
rect 187826 412098 188062 412334
rect 188146 412098 188382 412334
rect 187826 375218 188062 375454
rect 188146 375218 188382 375454
rect 187826 374898 188062 375134
rect 188146 374898 188382 375134
rect 187826 338018 188062 338254
rect 188146 338018 188382 338254
rect 187826 337698 188062 337934
rect 188146 337698 188382 337934
rect 187826 300818 188062 301054
rect 188146 300818 188382 301054
rect 187826 300498 188062 300734
rect 188146 300498 188382 300734
rect 187826 263618 188062 263854
rect 188146 263618 188382 263854
rect 187826 263298 188062 263534
rect 188146 263298 188382 263534
rect 187826 226418 188062 226654
rect 188146 226418 188382 226654
rect 187826 226098 188062 226334
rect 188146 226098 188382 226334
rect 187826 189218 188062 189454
rect 188146 189218 188382 189454
rect 187826 188898 188062 189134
rect 188146 188898 188382 189134
rect 187826 152018 188062 152254
rect 188146 152018 188382 152254
rect 187826 151698 188062 151934
rect 188146 151698 188382 151934
rect 187826 114818 188062 115054
rect 188146 114818 188382 115054
rect 187826 114498 188062 114734
rect 188146 114498 188382 114734
rect 187826 77618 188062 77854
rect 188146 77618 188382 77854
rect 187826 77298 188062 77534
rect 188146 77298 188382 77534
rect 187826 40418 188062 40654
rect 188146 40418 188382 40654
rect 187826 40098 188062 40334
rect 188146 40098 188382 40334
rect 187826 3218 188062 3454
rect 188146 3218 188382 3454
rect 187826 2898 188062 3134
rect 188146 2898 188382 3134
rect 191546 676538 191782 676774
rect 191866 676538 192102 676774
rect 191546 676218 191782 676454
rect 191866 676218 192102 676454
rect 191546 639338 191782 639574
rect 191866 639338 192102 639574
rect 191546 639018 191782 639254
rect 191866 639018 192102 639254
rect 191546 602138 191782 602374
rect 191866 602138 192102 602374
rect 191546 601818 191782 602054
rect 191866 601818 192102 602054
rect 191546 564938 191782 565174
rect 191866 564938 192102 565174
rect 191546 564618 191782 564854
rect 191866 564618 192102 564854
rect 191546 527738 191782 527974
rect 191866 527738 192102 527974
rect 191546 527418 191782 527654
rect 191866 527418 192102 527654
rect 191546 490538 191782 490774
rect 191866 490538 192102 490774
rect 191546 490218 191782 490454
rect 191866 490218 192102 490454
rect 191546 453338 191782 453574
rect 191866 453338 192102 453574
rect 191546 453018 191782 453254
rect 191866 453018 192102 453254
rect 191546 416138 191782 416374
rect 191866 416138 192102 416374
rect 191546 415818 191782 416054
rect 191866 415818 192102 416054
rect 191546 378938 191782 379174
rect 191866 378938 192102 379174
rect 191546 378618 191782 378854
rect 191866 378618 192102 378854
rect 191546 341738 191782 341974
rect 191866 341738 192102 341974
rect 191546 341418 191782 341654
rect 191866 341418 192102 341654
rect 191546 304538 191782 304774
rect 191866 304538 192102 304774
rect 191546 304218 191782 304454
rect 191866 304218 192102 304454
rect 191546 267338 191782 267574
rect 191866 267338 192102 267574
rect 191546 267018 191782 267254
rect 191866 267018 192102 267254
rect 191546 230138 191782 230374
rect 191866 230138 192102 230374
rect 191546 229818 191782 230054
rect 191866 229818 192102 230054
rect 191546 192938 191782 193174
rect 191866 192938 192102 193174
rect 191546 192618 191782 192854
rect 191866 192618 192102 192854
rect 191546 155738 191782 155974
rect 191866 155738 192102 155974
rect 191546 155418 191782 155654
rect 191866 155418 192102 155654
rect 191546 118538 191782 118774
rect 191866 118538 192102 118774
rect 191546 118218 191782 118454
rect 191866 118218 192102 118454
rect 191546 81338 191782 81574
rect 191866 81338 192102 81574
rect 191546 81018 191782 81254
rect 191866 81018 192102 81254
rect 191546 44138 191782 44374
rect 191866 44138 192102 44374
rect 191546 43818 191782 44054
rect 191866 43818 192102 44054
rect 191546 6938 191782 7174
rect 191866 6938 192102 7174
rect 191546 6618 191782 6854
rect 191866 6618 192102 6854
rect 195266 680258 195502 680494
rect 195586 680258 195822 680494
rect 195266 679938 195502 680174
rect 195586 679938 195822 680174
rect 195266 643058 195502 643294
rect 195586 643058 195822 643294
rect 195266 642738 195502 642974
rect 195586 642738 195822 642974
rect 195266 605858 195502 606094
rect 195586 605858 195822 606094
rect 195266 605538 195502 605774
rect 195586 605538 195822 605774
rect 195266 568658 195502 568894
rect 195586 568658 195822 568894
rect 195266 568338 195502 568574
rect 195586 568338 195822 568574
rect 195266 531458 195502 531694
rect 195586 531458 195822 531694
rect 195266 531138 195502 531374
rect 195586 531138 195822 531374
rect 195266 494258 195502 494494
rect 195586 494258 195822 494494
rect 195266 493938 195502 494174
rect 195586 493938 195822 494174
rect 195266 457058 195502 457294
rect 195586 457058 195822 457294
rect 195266 456738 195502 456974
rect 195586 456738 195822 456974
rect 195266 419858 195502 420094
rect 195586 419858 195822 420094
rect 195266 419538 195502 419774
rect 195586 419538 195822 419774
rect 195266 382658 195502 382894
rect 195586 382658 195822 382894
rect 195266 382338 195502 382574
rect 195586 382338 195822 382574
rect 195266 345458 195502 345694
rect 195586 345458 195822 345694
rect 195266 345138 195502 345374
rect 195586 345138 195822 345374
rect 195266 308258 195502 308494
rect 195586 308258 195822 308494
rect 195266 307938 195502 308174
rect 195586 307938 195822 308174
rect 195266 271058 195502 271294
rect 195586 271058 195822 271294
rect 195266 270738 195502 270974
rect 195586 270738 195822 270974
rect 195266 233858 195502 234094
rect 195586 233858 195822 234094
rect 195266 233538 195502 233774
rect 195586 233538 195822 233774
rect 195266 196658 195502 196894
rect 195586 196658 195822 196894
rect 195266 196338 195502 196574
rect 195586 196338 195822 196574
rect 195266 159458 195502 159694
rect 195586 159458 195822 159694
rect 195266 159138 195502 159374
rect 195586 159138 195822 159374
rect 195266 122258 195502 122494
rect 195586 122258 195822 122494
rect 195266 121938 195502 122174
rect 195586 121938 195822 122174
rect 195266 85058 195502 85294
rect 195586 85058 195822 85294
rect 195266 84738 195502 84974
rect 195586 84738 195822 84974
rect 195266 47858 195502 48094
rect 195586 47858 195822 48094
rect 195266 47538 195502 47774
rect 195586 47538 195822 47774
rect 195266 10658 195502 10894
rect 195586 10658 195822 10894
rect 195266 10338 195502 10574
rect 195586 10338 195822 10574
rect 198986 683978 199222 684214
rect 199306 683978 199542 684214
rect 198986 683658 199222 683894
rect 199306 683658 199542 683894
rect 198986 646778 199222 647014
rect 199306 646778 199542 647014
rect 198986 646458 199222 646694
rect 199306 646458 199542 646694
rect 198986 609578 199222 609814
rect 199306 609578 199542 609814
rect 198986 609258 199222 609494
rect 199306 609258 199542 609494
rect 198986 572378 199222 572614
rect 199306 572378 199542 572614
rect 198986 572058 199222 572294
rect 199306 572058 199542 572294
rect 198986 535178 199222 535414
rect 199306 535178 199542 535414
rect 198986 534858 199222 535094
rect 199306 534858 199542 535094
rect 198986 497978 199222 498214
rect 199306 497978 199542 498214
rect 198986 497658 199222 497894
rect 199306 497658 199542 497894
rect 198986 460778 199222 461014
rect 199306 460778 199542 461014
rect 198986 460458 199222 460694
rect 199306 460458 199542 460694
rect 198986 423578 199222 423814
rect 199306 423578 199542 423814
rect 198986 423258 199222 423494
rect 199306 423258 199542 423494
rect 198986 386378 199222 386614
rect 199306 386378 199542 386614
rect 198986 386058 199222 386294
rect 199306 386058 199542 386294
rect 198986 349178 199222 349414
rect 199306 349178 199542 349414
rect 198986 348858 199222 349094
rect 199306 348858 199542 349094
rect 198986 311978 199222 312214
rect 199306 311978 199542 312214
rect 198986 311658 199222 311894
rect 199306 311658 199542 311894
rect 198986 274778 199222 275014
rect 199306 274778 199542 275014
rect 198986 274458 199222 274694
rect 199306 274458 199542 274694
rect 198986 237578 199222 237814
rect 199306 237578 199542 237814
rect 198986 237258 199222 237494
rect 199306 237258 199542 237494
rect 198986 200378 199222 200614
rect 199306 200378 199542 200614
rect 198986 200058 199222 200294
rect 199306 200058 199542 200294
rect 198986 163178 199222 163414
rect 199306 163178 199542 163414
rect 198986 162858 199222 163094
rect 199306 162858 199542 163094
rect 198986 125978 199222 126214
rect 199306 125978 199542 126214
rect 198986 125658 199222 125894
rect 199306 125658 199542 125894
rect 198986 88778 199222 89014
rect 199306 88778 199542 89014
rect 198986 88458 199222 88694
rect 199306 88458 199542 88694
rect 198986 51578 199222 51814
rect 199306 51578 199542 51814
rect 198986 51258 199222 51494
rect 199306 51258 199542 51494
rect 198986 14378 199222 14614
rect 199306 14378 199542 14614
rect 198986 14058 199222 14294
rect 199306 14058 199542 14294
rect 202706 687698 202942 687934
rect 203026 687698 203262 687934
rect 202706 687378 202942 687614
rect 203026 687378 203262 687614
rect 202706 650498 202942 650734
rect 203026 650498 203262 650734
rect 202706 650178 202942 650414
rect 203026 650178 203262 650414
rect 202706 613298 202942 613534
rect 203026 613298 203262 613534
rect 202706 612978 202942 613214
rect 203026 612978 203262 613214
rect 202706 576098 202942 576334
rect 203026 576098 203262 576334
rect 202706 575778 202942 576014
rect 203026 575778 203262 576014
rect 202706 538898 202942 539134
rect 203026 538898 203262 539134
rect 202706 538578 202942 538814
rect 203026 538578 203262 538814
rect 202706 501698 202942 501934
rect 203026 501698 203262 501934
rect 202706 501378 202942 501614
rect 203026 501378 203262 501614
rect 202706 464498 202942 464734
rect 203026 464498 203262 464734
rect 202706 464178 202942 464414
rect 203026 464178 203262 464414
rect 202706 427298 202942 427534
rect 203026 427298 203262 427534
rect 202706 426978 202942 427214
rect 203026 426978 203262 427214
rect 202706 390098 202942 390334
rect 203026 390098 203262 390334
rect 202706 389778 202942 390014
rect 203026 389778 203262 390014
rect 202706 352898 202942 353134
rect 203026 352898 203262 353134
rect 202706 352578 202942 352814
rect 203026 352578 203262 352814
rect 202706 315698 202942 315934
rect 203026 315698 203262 315934
rect 202706 315378 202942 315614
rect 203026 315378 203262 315614
rect 202706 278498 202942 278734
rect 203026 278498 203262 278734
rect 202706 278178 202942 278414
rect 203026 278178 203262 278414
rect 202706 241298 202942 241534
rect 203026 241298 203262 241534
rect 202706 240978 202942 241214
rect 203026 240978 203262 241214
rect 202706 204098 202942 204334
rect 203026 204098 203262 204334
rect 202706 203778 202942 204014
rect 203026 203778 203262 204014
rect 202706 166898 202942 167134
rect 203026 166898 203262 167134
rect 202706 166578 202942 166814
rect 203026 166578 203262 166814
rect 202706 129698 202942 129934
rect 203026 129698 203262 129934
rect 202706 129378 202942 129614
rect 203026 129378 203262 129614
rect 202706 92498 202942 92734
rect 203026 92498 203262 92734
rect 202706 92178 202942 92414
rect 203026 92178 203262 92414
rect 202706 55298 202942 55534
rect 203026 55298 203262 55534
rect 202706 54978 202942 55214
rect 203026 54978 203262 55214
rect 202706 18098 202942 18334
rect 203026 18098 203262 18334
rect 202706 17778 202942 18014
rect 203026 17778 203262 18014
rect 206426 691418 206662 691654
rect 206746 691418 206982 691654
rect 206426 691098 206662 691334
rect 206746 691098 206982 691334
rect 206426 654218 206662 654454
rect 206746 654218 206982 654454
rect 206426 653898 206662 654134
rect 206746 653898 206982 654134
rect 206426 617018 206662 617254
rect 206746 617018 206982 617254
rect 206426 616698 206662 616934
rect 206746 616698 206982 616934
rect 206426 579818 206662 580054
rect 206746 579818 206982 580054
rect 206426 579498 206662 579734
rect 206746 579498 206982 579734
rect 206426 542618 206662 542854
rect 206746 542618 206982 542854
rect 206426 542298 206662 542534
rect 206746 542298 206982 542534
rect 206426 505418 206662 505654
rect 206746 505418 206982 505654
rect 206426 505098 206662 505334
rect 206746 505098 206982 505334
rect 206426 468218 206662 468454
rect 206746 468218 206982 468454
rect 206426 467898 206662 468134
rect 206746 467898 206982 468134
rect 206426 431018 206662 431254
rect 206746 431018 206982 431254
rect 206426 430698 206662 430934
rect 206746 430698 206982 430934
rect 206426 393818 206662 394054
rect 206746 393818 206982 394054
rect 206426 393498 206662 393734
rect 206746 393498 206982 393734
rect 206426 356618 206662 356854
rect 206746 356618 206982 356854
rect 206426 356298 206662 356534
rect 206746 356298 206982 356534
rect 206426 319418 206662 319654
rect 206746 319418 206982 319654
rect 206426 319098 206662 319334
rect 206746 319098 206982 319334
rect 206426 282218 206662 282454
rect 206746 282218 206982 282454
rect 206426 281898 206662 282134
rect 206746 281898 206982 282134
rect 206426 245018 206662 245254
rect 206746 245018 206982 245254
rect 206426 244698 206662 244934
rect 206746 244698 206982 244934
rect 206426 207818 206662 208054
rect 206746 207818 206982 208054
rect 206426 207498 206662 207734
rect 206746 207498 206982 207734
rect 206426 170618 206662 170854
rect 206746 170618 206982 170854
rect 206426 170298 206662 170534
rect 206746 170298 206982 170534
rect 206426 133418 206662 133654
rect 206746 133418 206982 133654
rect 206426 133098 206662 133334
rect 206746 133098 206982 133334
rect 206426 96218 206662 96454
rect 206746 96218 206982 96454
rect 206426 95898 206662 96134
rect 206746 95898 206982 96134
rect 206426 59018 206662 59254
rect 206746 59018 206982 59254
rect 206426 58698 206662 58934
rect 206746 58698 206982 58934
rect 206426 21818 206662 22054
rect 206746 21818 206982 22054
rect 206426 21498 206662 21734
rect 206746 21498 206982 21734
rect 210146 695138 210382 695374
rect 210466 695138 210702 695374
rect 210146 694818 210382 695054
rect 210466 694818 210702 695054
rect 210146 657938 210382 658174
rect 210466 657938 210702 658174
rect 210146 657618 210382 657854
rect 210466 657618 210702 657854
rect 210146 620738 210382 620974
rect 210466 620738 210702 620974
rect 210146 620418 210382 620654
rect 210466 620418 210702 620654
rect 210146 583538 210382 583774
rect 210466 583538 210702 583774
rect 210146 583218 210382 583454
rect 210466 583218 210702 583454
rect 210146 546338 210382 546574
rect 210466 546338 210702 546574
rect 210146 546018 210382 546254
rect 210466 546018 210702 546254
rect 210146 509138 210382 509374
rect 210466 509138 210702 509374
rect 210146 508818 210382 509054
rect 210466 508818 210702 509054
rect 210146 471938 210382 472174
rect 210466 471938 210702 472174
rect 210146 471618 210382 471854
rect 210466 471618 210702 471854
rect 210146 434738 210382 434974
rect 210466 434738 210702 434974
rect 210146 434418 210382 434654
rect 210466 434418 210702 434654
rect 210146 397538 210382 397774
rect 210466 397538 210702 397774
rect 210146 397218 210382 397454
rect 210466 397218 210702 397454
rect 210146 360338 210382 360574
rect 210466 360338 210702 360574
rect 210146 360018 210382 360254
rect 210466 360018 210702 360254
rect 210146 323138 210382 323374
rect 210466 323138 210702 323374
rect 210146 322818 210382 323054
rect 210466 322818 210702 323054
rect 210146 285938 210382 286174
rect 210466 285938 210702 286174
rect 210146 285618 210382 285854
rect 210466 285618 210702 285854
rect 210146 248738 210382 248974
rect 210466 248738 210702 248974
rect 210146 248418 210382 248654
rect 210466 248418 210702 248654
rect 210146 211538 210382 211774
rect 210466 211538 210702 211774
rect 210146 211218 210382 211454
rect 210466 211218 210702 211454
rect 210146 174338 210382 174574
rect 210466 174338 210702 174574
rect 210146 174018 210382 174254
rect 210466 174018 210702 174254
rect 210146 137138 210382 137374
rect 210466 137138 210702 137374
rect 210146 136818 210382 137054
rect 210466 136818 210702 137054
rect 210146 99938 210382 100174
rect 210466 99938 210702 100174
rect 210146 99618 210382 99854
rect 210466 99618 210702 99854
rect 210146 62738 210382 62974
rect 210466 62738 210702 62974
rect 210146 62418 210382 62654
rect 210466 62418 210702 62654
rect 210146 25538 210382 25774
rect 210466 25538 210702 25774
rect 210146 25218 210382 25454
rect 210466 25218 210702 25454
rect 213866 698858 214102 699094
rect 214186 698858 214422 699094
rect 213866 698538 214102 698774
rect 214186 698538 214422 698774
rect 213866 661658 214102 661894
rect 214186 661658 214422 661894
rect 213866 661338 214102 661574
rect 214186 661338 214422 661574
rect 213866 624458 214102 624694
rect 214186 624458 214422 624694
rect 213866 624138 214102 624374
rect 214186 624138 214422 624374
rect 213866 587258 214102 587494
rect 214186 587258 214422 587494
rect 213866 586938 214102 587174
rect 214186 586938 214422 587174
rect 213866 550058 214102 550294
rect 214186 550058 214422 550294
rect 213866 549738 214102 549974
rect 214186 549738 214422 549974
rect 213866 512858 214102 513094
rect 214186 512858 214422 513094
rect 213866 512538 214102 512774
rect 214186 512538 214422 512774
rect 213866 475658 214102 475894
rect 214186 475658 214422 475894
rect 213866 475338 214102 475574
rect 214186 475338 214422 475574
rect 213866 438458 214102 438694
rect 214186 438458 214422 438694
rect 213866 438138 214102 438374
rect 214186 438138 214422 438374
rect 213866 401258 214102 401494
rect 214186 401258 214422 401494
rect 213866 400938 214102 401174
rect 214186 400938 214422 401174
rect 213866 364058 214102 364294
rect 214186 364058 214422 364294
rect 213866 363738 214102 363974
rect 214186 363738 214422 363974
rect 213866 326858 214102 327094
rect 214186 326858 214422 327094
rect 213866 326538 214102 326774
rect 214186 326538 214422 326774
rect 213866 289658 214102 289894
rect 214186 289658 214422 289894
rect 213866 289338 214102 289574
rect 214186 289338 214422 289574
rect 213866 252458 214102 252694
rect 214186 252458 214422 252694
rect 213866 252138 214102 252374
rect 214186 252138 214422 252374
rect 213866 215258 214102 215494
rect 214186 215258 214422 215494
rect 213866 214938 214102 215174
rect 214186 214938 214422 215174
rect 213866 178058 214102 178294
rect 214186 178058 214422 178294
rect 213866 177738 214102 177974
rect 214186 177738 214422 177974
rect 213866 140858 214102 141094
rect 214186 140858 214422 141094
rect 213866 140538 214102 140774
rect 214186 140538 214422 140774
rect 213866 103658 214102 103894
rect 214186 103658 214422 103894
rect 213866 103338 214102 103574
rect 214186 103338 214422 103574
rect 213866 66458 214102 66694
rect 214186 66458 214422 66694
rect 213866 66138 214102 66374
rect 214186 66138 214422 66374
rect 213866 29258 214102 29494
rect 214186 29258 214422 29494
rect 213866 28938 214102 29174
rect 214186 28938 214422 29174
rect 225026 672818 225262 673054
rect 225346 672818 225582 673054
rect 225026 672498 225262 672734
rect 225346 672498 225582 672734
rect 225026 635618 225262 635854
rect 225346 635618 225582 635854
rect 225026 635298 225262 635534
rect 225346 635298 225582 635534
rect 225026 598418 225262 598654
rect 225346 598418 225582 598654
rect 225026 598098 225262 598334
rect 225346 598098 225582 598334
rect 225026 561218 225262 561454
rect 225346 561218 225582 561454
rect 225026 560898 225262 561134
rect 225346 560898 225582 561134
rect 225026 524018 225262 524254
rect 225346 524018 225582 524254
rect 225026 523698 225262 523934
rect 225346 523698 225582 523934
rect 225026 486818 225262 487054
rect 225346 486818 225582 487054
rect 225026 486498 225262 486734
rect 225346 486498 225582 486734
rect 225026 449618 225262 449854
rect 225346 449618 225582 449854
rect 225026 449298 225262 449534
rect 225346 449298 225582 449534
rect 225026 412418 225262 412654
rect 225346 412418 225582 412654
rect 225026 412098 225262 412334
rect 225346 412098 225582 412334
rect 225026 375218 225262 375454
rect 225346 375218 225582 375454
rect 225026 374898 225262 375134
rect 225346 374898 225582 375134
rect 225026 338018 225262 338254
rect 225346 338018 225582 338254
rect 225026 337698 225262 337934
rect 225346 337698 225582 337934
rect 225026 300818 225262 301054
rect 225346 300818 225582 301054
rect 225026 300498 225262 300734
rect 225346 300498 225582 300734
rect 225026 263618 225262 263854
rect 225346 263618 225582 263854
rect 225026 263298 225262 263534
rect 225346 263298 225582 263534
rect 225026 226418 225262 226654
rect 225346 226418 225582 226654
rect 225026 226098 225262 226334
rect 225346 226098 225582 226334
rect 225026 189218 225262 189454
rect 225346 189218 225582 189454
rect 225026 188898 225262 189134
rect 225346 188898 225582 189134
rect 225026 152018 225262 152254
rect 225346 152018 225582 152254
rect 225026 151698 225262 151934
rect 225346 151698 225582 151934
rect 225026 114818 225262 115054
rect 225346 114818 225582 115054
rect 225026 114498 225262 114734
rect 225346 114498 225582 114734
rect 225026 77618 225262 77854
rect 225346 77618 225582 77854
rect 225026 77298 225262 77534
rect 225346 77298 225582 77534
rect 225026 40418 225262 40654
rect 225346 40418 225582 40654
rect 225026 40098 225262 40334
rect 225346 40098 225582 40334
rect 225026 3218 225262 3454
rect 225346 3218 225582 3454
rect 225026 2898 225262 3134
rect 225346 2898 225582 3134
rect 228746 676538 228982 676774
rect 229066 676538 229302 676774
rect 228746 676218 228982 676454
rect 229066 676218 229302 676454
rect 228746 639338 228982 639574
rect 229066 639338 229302 639574
rect 228746 639018 228982 639254
rect 229066 639018 229302 639254
rect 228746 602138 228982 602374
rect 229066 602138 229302 602374
rect 228746 601818 228982 602054
rect 229066 601818 229302 602054
rect 228746 564938 228982 565174
rect 229066 564938 229302 565174
rect 228746 564618 228982 564854
rect 229066 564618 229302 564854
rect 228746 527738 228982 527974
rect 229066 527738 229302 527974
rect 228746 527418 228982 527654
rect 229066 527418 229302 527654
rect 228746 490538 228982 490774
rect 229066 490538 229302 490774
rect 228746 490218 228982 490454
rect 229066 490218 229302 490454
rect 228746 453338 228982 453574
rect 229066 453338 229302 453574
rect 228746 453018 228982 453254
rect 229066 453018 229302 453254
rect 228746 416138 228982 416374
rect 229066 416138 229302 416374
rect 228746 415818 228982 416054
rect 229066 415818 229302 416054
rect 228746 378938 228982 379174
rect 229066 378938 229302 379174
rect 228746 378618 228982 378854
rect 229066 378618 229302 378854
rect 228746 341738 228982 341974
rect 229066 341738 229302 341974
rect 228746 341418 228982 341654
rect 229066 341418 229302 341654
rect 228746 304538 228982 304774
rect 229066 304538 229302 304774
rect 228746 304218 228982 304454
rect 229066 304218 229302 304454
rect 228746 267338 228982 267574
rect 229066 267338 229302 267574
rect 228746 267018 228982 267254
rect 229066 267018 229302 267254
rect 228746 230138 228982 230374
rect 229066 230138 229302 230374
rect 228746 229818 228982 230054
rect 229066 229818 229302 230054
rect 228746 192938 228982 193174
rect 229066 192938 229302 193174
rect 228746 192618 228982 192854
rect 229066 192618 229302 192854
rect 228746 155738 228982 155974
rect 229066 155738 229302 155974
rect 228746 155418 228982 155654
rect 229066 155418 229302 155654
rect 228746 118538 228982 118774
rect 229066 118538 229302 118774
rect 228746 118218 228982 118454
rect 229066 118218 229302 118454
rect 228746 81338 228982 81574
rect 229066 81338 229302 81574
rect 228746 81018 228982 81254
rect 229066 81018 229302 81254
rect 228746 44138 228982 44374
rect 229066 44138 229302 44374
rect 228746 43818 228982 44054
rect 229066 43818 229302 44054
rect 228746 6938 228982 7174
rect 229066 6938 229302 7174
rect 228746 6618 228982 6854
rect 229066 6618 229302 6854
rect 232466 680258 232702 680494
rect 232786 680258 233022 680494
rect 232466 679938 232702 680174
rect 232786 679938 233022 680174
rect 232466 643058 232702 643294
rect 232786 643058 233022 643294
rect 232466 642738 232702 642974
rect 232786 642738 233022 642974
rect 232466 605858 232702 606094
rect 232786 605858 233022 606094
rect 232466 605538 232702 605774
rect 232786 605538 233022 605774
rect 232466 568658 232702 568894
rect 232786 568658 233022 568894
rect 232466 568338 232702 568574
rect 232786 568338 233022 568574
rect 232466 531458 232702 531694
rect 232786 531458 233022 531694
rect 232466 531138 232702 531374
rect 232786 531138 233022 531374
rect 232466 494258 232702 494494
rect 232786 494258 233022 494494
rect 232466 493938 232702 494174
rect 232786 493938 233022 494174
rect 232466 457058 232702 457294
rect 232786 457058 233022 457294
rect 232466 456738 232702 456974
rect 232786 456738 233022 456974
rect 232466 419858 232702 420094
rect 232786 419858 233022 420094
rect 232466 419538 232702 419774
rect 232786 419538 233022 419774
rect 232466 382658 232702 382894
rect 232786 382658 233022 382894
rect 232466 382338 232702 382574
rect 232786 382338 233022 382574
rect 232466 345458 232702 345694
rect 232786 345458 233022 345694
rect 232466 345138 232702 345374
rect 232786 345138 233022 345374
rect 232466 308258 232702 308494
rect 232786 308258 233022 308494
rect 232466 307938 232702 308174
rect 232786 307938 233022 308174
rect 232466 271058 232702 271294
rect 232786 271058 233022 271294
rect 232466 270738 232702 270974
rect 232786 270738 233022 270974
rect 232466 233858 232702 234094
rect 232786 233858 233022 234094
rect 232466 233538 232702 233774
rect 232786 233538 233022 233774
rect 232466 196658 232702 196894
rect 232786 196658 233022 196894
rect 232466 196338 232702 196574
rect 232786 196338 233022 196574
rect 232466 159458 232702 159694
rect 232786 159458 233022 159694
rect 232466 159138 232702 159374
rect 232786 159138 233022 159374
rect 232466 122258 232702 122494
rect 232786 122258 233022 122494
rect 232466 121938 232702 122174
rect 232786 121938 233022 122174
rect 232466 85058 232702 85294
rect 232786 85058 233022 85294
rect 232466 84738 232702 84974
rect 232786 84738 233022 84974
rect 232466 47858 232702 48094
rect 232786 47858 233022 48094
rect 232466 47538 232702 47774
rect 232786 47538 233022 47774
rect 232466 10658 232702 10894
rect 232786 10658 233022 10894
rect 232466 10338 232702 10574
rect 232786 10338 233022 10574
rect 236186 683978 236422 684214
rect 236506 683978 236742 684214
rect 236186 683658 236422 683894
rect 236506 683658 236742 683894
rect 236186 646778 236422 647014
rect 236506 646778 236742 647014
rect 236186 646458 236422 646694
rect 236506 646458 236742 646694
rect 236186 609578 236422 609814
rect 236506 609578 236742 609814
rect 236186 609258 236422 609494
rect 236506 609258 236742 609494
rect 236186 572378 236422 572614
rect 236506 572378 236742 572614
rect 236186 572058 236422 572294
rect 236506 572058 236742 572294
rect 236186 535178 236422 535414
rect 236506 535178 236742 535414
rect 236186 534858 236422 535094
rect 236506 534858 236742 535094
rect 236186 497978 236422 498214
rect 236506 497978 236742 498214
rect 236186 497658 236422 497894
rect 236506 497658 236742 497894
rect 236186 460778 236422 461014
rect 236506 460778 236742 461014
rect 236186 460458 236422 460694
rect 236506 460458 236742 460694
rect 236186 423578 236422 423814
rect 236506 423578 236742 423814
rect 236186 423258 236422 423494
rect 236506 423258 236742 423494
rect 236186 386378 236422 386614
rect 236506 386378 236742 386614
rect 236186 386058 236422 386294
rect 236506 386058 236742 386294
rect 236186 349178 236422 349414
rect 236506 349178 236742 349414
rect 236186 348858 236422 349094
rect 236506 348858 236742 349094
rect 236186 311978 236422 312214
rect 236506 311978 236742 312214
rect 236186 311658 236422 311894
rect 236506 311658 236742 311894
rect 236186 274778 236422 275014
rect 236506 274778 236742 275014
rect 236186 274458 236422 274694
rect 236506 274458 236742 274694
rect 236186 237578 236422 237814
rect 236506 237578 236742 237814
rect 236186 237258 236422 237494
rect 236506 237258 236742 237494
rect 236186 200378 236422 200614
rect 236506 200378 236742 200614
rect 236186 200058 236422 200294
rect 236506 200058 236742 200294
rect 236186 163178 236422 163414
rect 236506 163178 236742 163414
rect 236186 162858 236422 163094
rect 236506 162858 236742 163094
rect 236186 125978 236422 126214
rect 236506 125978 236742 126214
rect 236186 125658 236422 125894
rect 236506 125658 236742 125894
rect 236186 88778 236422 89014
rect 236506 88778 236742 89014
rect 236186 88458 236422 88694
rect 236506 88458 236742 88694
rect 236186 51578 236422 51814
rect 236506 51578 236742 51814
rect 236186 51258 236422 51494
rect 236506 51258 236742 51494
rect 236186 14378 236422 14614
rect 236506 14378 236742 14614
rect 236186 14058 236422 14294
rect 236506 14058 236742 14294
rect 239906 687698 240142 687934
rect 240226 687698 240462 687934
rect 239906 687378 240142 687614
rect 240226 687378 240462 687614
rect 239906 650498 240142 650734
rect 240226 650498 240462 650734
rect 239906 650178 240142 650414
rect 240226 650178 240462 650414
rect 239906 613298 240142 613534
rect 240226 613298 240462 613534
rect 239906 612978 240142 613214
rect 240226 612978 240462 613214
rect 239906 576098 240142 576334
rect 240226 576098 240462 576334
rect 239906 575778 240142 576014
rect 240226 575778 240462 576014
rect 239906 538898 240142 539134
rect 240226 538898 240462 539134
rect 239906 538578 240142 538814
rect 240226 538578 240462 538814
rect 239906 501698 240142 501934
rect 240226 501698 240462 501934
rect 239906 501378 240142 501614
rect 240226 501378 240462 501614
rect 239906 464498 240142 464734
rect 240226 464498 240462 464734
rect 239906 464178 240142 464414
rect 240226 464178 240462 464414
rect 239906 427298 240142 427534
rect 240226 427298 240462 427534
rect 239906 426978 240142 427214
rect 240226 426978 240462 427214
rect 239906 390098 240142 390334
rect 240226 390098 240462 390334
rect 239906 389778 240142 390014
rect 240226 389778 240462 390014
rect 239906 352898 240142 353134
rect 240226 352898 240462 353134
rect 239906 352578 240142 352814
rect 240226 352578 240462 352814
rect 239906 315698 240142 315934
rect 240226 315698 240462 315934
rect 239906 315378 240142 315614
rect 240226 315378 240462 315614
rect 239906 278498 240142 278734
rect 240226 278498 240462 278734
rect 239906 278178 240142 278414
rect 240226 278178 240462 278414
rect 239906 241298 240142 241534
rect 240226 241298 240462 241534
rect 239906 240978 240142 241214
rect 240226 240978 240462 241214
rect 239906 204098 240142 204334
rect 240226 204098 240462 204334
rect 239906 203778 240142 204014
rect 240226 203778 240462 204014
rect 239906 166898 240142 167134
rect 240226 166898 240462 167134
rect 239906 166578 240142 166814
rect 240226 166578 240462 166814
rect 239906 129698 240142 129934
rect 240226 129698 240462 129934
rect 239906 129378 240142 129614
rect 240226 129378 240462 129614
rect 239906 92498 240142 92734
rect 240226 92498 240462 92734
rect 239906 92178 240142 92414
rect 240226 92178 240462 92414
rect 239906 55298 240142 55534
rect 240226 55298 240462 55534
rect 239906 54978 240142 55214
rect 240226 54978 240462 55214
rect 239906 18098 240142 18334
rect 240226 18098 240462 18334
rect 239906 17778 240142 18014
rect 240226 17778 240462 18014
rect 243626 691418 243862 691654
rect 243946 691418 244182 691654
rect 243626 691098 243862 691334
rect 243946 691098 244182 691334
rect 243626 654218 243862 654454
rect 243946 654218 244182 654454
rect 243626 653898 243862 654134
rect 243946 653898 244182 654134
rect 243626 617018 243862 617254
rect 243946 617018 244182 617254
rect 243626 616698 243862 616934
rect 243946 616698 244182 616934
rect 243626 579818 243862 580054
rect 243946 579818 244182 580054
rect 243626 579498 243862 579734
rect 243946 579498 244182 579734
rect 243626 542618 243862 542854
rect 243946 542618 244182 542854
rect 243626 542298 243862 542534
rect 243946 542298 244182 542534
rect 243626 505418 243862 505654
rect 243946 505418 244182 505654
rect 243626 505098 243862 505334
rect 243946 505098 244182 505334
rect 243626 468218 243862 468454
rect 243946 468218 244182 468454
rect 243626 467898 243862 468134
rect 243946 467898 244182 468134
rect 243626 431018 243862 431254
rect 243946 431018 244182 431254
rect 243626 430698 243862 430934
rect 243946 430698 244182 430934
rect 243626 393818 243862 394054
rect 243946 393818 244182 394054
rect 243626 393498 243862 393734
rect 243946 393498 244182 393734
rect 243626 356618 243862 356854
rect 243946 356618 244182 356854
rect 243626 356298 243862 356534
rect 243946 356298 244182 356534
rect 243626 319418 243862 319654
rect 243946 319418 244182 319654
rect 243626 319098 243862 319334
rect 243946 319098 244182 319334
rect 243626 282218 243862 282454
rect 243946 282218 244182 282454
rect 243626 281898 243862 282134
rect 243946 281898 244182 282134
rect 243626 245018 243862 245254
rect 243946 245018 244182 245254
rect 243626 244698 243862 244934
rect 243946 244698 244182 244934
rect 243626 207818 243862 208054
rect 243946 207818 244182 208054
rect 243626 207498 243862 207734
rect 243946 207498 244182 207734
rect 243626 170618 243862 170854
rect 243946 170618 244182 170854
rect 243626 170298 243862 170534
rect 243946 170298 244182 170534
rect 243626 133418 243862 133654
rect 243946 133418 244182 133654
rect 243626 133098 243862 133334
rect 243946 133098 244182 133334
rect 243626 96218 243862 96454
rect 243946 96218 244182 96454
rect 243626 95898 243862 96134
rect 243946 95898 244182 96134
rect 243626 59018 243862 59254
rect 243946 59018 244182 59254
rect 243626 58698 243862 58934
rect 243946 58698 244182 58934
rect 243626 21818 243862 22054
rect 243946 21818 244182 22054
rect 243626 21498 243862 21734
rect 243946 21498 244182 21734
rect 247346 695138 247582 695374
rect 247666 695138 247902 695374
rect 247346 694818 247582 695054
rect 247666 694818 247902 695054
rect 247346 657938 247582 658174
rect 247666 657938 247902 658174
rect 247346 657618 247582 657854
rect 247666 657618 247902 657854
rect 247346 620738 247582 620974
rect 247666 620738 247902 620974
rect 247346 620418 247582 620654
rect 247666 620418 247902 620654
rect 247346 583538 247582 583774
rect 247666 583538 247902 583774
rect 247346 583218 247582 583454
rect 247666 583218 247902 583454
rect 247346 546338 247582 546574
rect 247666 546338 247902 546574
rect 247346 546018 247582 546254
rect 247666 546018 247902 546254
rect 247346 509138 247582 509374
rect 247666 509138 247902 509374
rect 247346 508818 247582 509054
rect 247666 508818 247902 509054
rect 247346 471938 247582 472174
rect 247666 471938 247902 472174
rect 247346 471618 247582 471854
rect 247666 471618 247902 471854
rect 247346 434738 247582 434974
rect 247666 434738 247902 434974
rect 247346 434418 247582 434654
rect 247666 434418 247902 434654
rect 247346 397538 247582 397774
rect 247666 397538 247902 397774
rect 247346 397218 247582 397454
rect 247666 397218 247902 397454
rect 247346 360338 247582 360574
rect 247666 360338 247902 360574
rect 247346 360018 247582 360254
rect 247666 360018 247902 360254
rect 247346 323138 247582 323374
rect 247666 323138 247902 323374
rect 247346 322818 247582 323054
rect 247666 322818 247902 323054
rect 247346 285938 247582 286174
rect 247666 285938 247902 286174
rect 247346 285618 247582 285854
rect 247666 285618 247902 285854
rect 247346 248738 247582 248974
rect 247666 248738 247902 248974
rect 247346 248418 247582 248654
rect 247666 248418 247902 248654
rect 247346 211538 247582 211774
rect 247666 211538 247902 211774
rect 247346 211218 247582 211454
rect 247666 211218 247902 211454
rect 247346 174338 247582 174574
rect 247666 174338 247902 174574
rect 247346 174018 247582 174254
rect 247666 174018 247902 174254
rect 247346 137138 247582 137374
rect 247666 137138 247902 137374
rect 247346 136818 247582 137054
rect 247666 136818 247902 137054
rect 247346 99938 247582 100174
rect 247666 99938 247902 100174
rect 247346 99618 247582 99854
rect 247666 99618 247902 99854
rect 247346 62738 247582 62974
rect 247666 62738 247902 62974
rect 247346 62418 247582 62654
rect 247666 62418 247902 62654
rect 247346 25538 247582 25774
rect 247666 25538 247902 25774
rect 247346 25218 247582 25454
rect 247666 25218 247902 25454
rect 251066 698858 251302 699094
rect 251386 698858 251622 699094
rect 251066 698538 251302 698774
rect 251386 698538 251622 698774
rect 251066 661658 251302 661894
rect 251386 661658 251622 661894
rect 251066 661338 251302 661574
rect 251386 661338 251622 661574
rect 251066 624458 251302 624694
rect 251386 624458 251622 624694
rect 251066 624138 251302 624374
rect 251386 624138 251622 624374
rect 251066 587258 251302 587494
rect 251386 587258 251622 587494
rect 251066 586938 251302 587174
rect 251386 586938 251622 587174
rect 251066 550058 251302 550294
rect 251386 550058 251622 550294
rect 251066 549738 251302 549974
rect 251386 549738 251622 549974
rect 251066 512858 251302 513094
rect 251386 512858 251622 513094
rect 251066 512538 251302 512774
rect 251386 512538 251622 512774
rect 251066 475658 251302 475894
rect 251386 475658 251622 475894
rect 251066 475338 251302 475574
rect 251386 475338 251622 475574
rect 251066 438458 251302 438694
rect 251386 438458 251622 438694
rect 251066 438138 251302 438374
rect 251386 438138 251622 438374
rect 251066 401258 251302 401494
rect 251386 401258 251622 401494
rect 251066 400938 251302 401174
rect 251386 400938 251622 401174
rect 251066 364058 251302 364294
rect 251386 364058 251622 364294
rect 251066 363738 251302 363974
rect 251386 363738 251622 363974
rect 251066 326858 251302 327094
rect 251386 326858 251622 327094
rect 251066 326538 251302 326774
rect 251386 326538 251622 326774
rect 251066 289658 251302 289894
rect 251386 289658 251622 289894
rect 251066 289338 251302 289574
rect 251386 289338 251622 289574
rect 251066 252458 251302 252694
rect 251386 252458 251622 252694
rect 251066 252138 251302 252374
rect 251386 252138 251622 252374
rect 251066 215258 251302 215494
rect 251386 215258 251622 215494
rect 251066 214938 251302 215174
rect 251386 214938 251622 215174
rect 251066 178058 251302 178294
rect 251386 178058 251622 178294
rect 251066 177738 251302 177974
rect 251386 177738 251622 177974
rect 251066 140858 251302 141094
rect 251386 140858 251622 141094
rect 251066 140538 251302 140774
rect 251386 140538 251622 140774
rect 251066 103658 251302 103894
rect 251386 103658 251622 103894
rect 251066 103338 251302 103574
rect 251386 103338 251622 103574
rect 251066 66458 251302 66694
rect 251386 66458 251622 66694
rect 251066 66138 251302 66374
rect 251386 66138 251622 66374
rect 251066 29258 251302 29494
rect 251386 29258 251622 29494
rect 251066 28938 251302 29174
rect 251386 28938 251622 29174
rect 262226 672818 262462 673054
rect 262546 672818 262782 673054
rect 262226 672498 262462 672734
rect 262546 672498 262782 672734
rect 262226 635618 262462 635854
rect 262546 635618 262782 635854
rect 262226 635298 262462 635534
rect 262546 635298 262782 635534
rect 262226 598418 262462 598654
rect 262546 598418 262782 598654
rect 262226 598098 262462 598334
rect 262546 598098 262782 598334
rect 262226 561218 262462 561454
rect 262546 561218 262782 561454
rect 262226 560898 262462 561134
rect 262546 560898 262782 561134
rect 262226 524018 262462 524254
rect 262546 524018 262782 524254
rect 262226 523698 262462 523934
rect 262546 523698 262782 523934
rect 262226 486818 262462 487054
rect 262546 486818 262782 487054
rect 262226 486498 262462 486734
rect 262546 486498 262782 486734
rect 262226 449618 262462 449854
rect 262546 449618 262782 449854
rect 262226 449298 262462 449534
rect 262546 449298 262782 449534
rect 262226 412418 262462 412654
rect 262546 412418 262782 412654
rect 262226 412098 262462 412334
rect 262546 412098 262782 412334
rect 262226 375218 262462 375454
rect 262546 375218 262782 375454
rect 262226 374898 262462 375134
rect 262546 374898 262782 375134
rect 262226 338018 262462 338254
rect 262546 338018 262782 338254
rect 262226 337698 262462 337934
rect 262546 337698 262782 337934
rect 262226 300818 262462 301054
rect 262546 300818 262782 301054
rect 262226 300498 262462 300734
rect 262546 300498 262782 300734
rect 262226 263618 262462 263854
rect 262546 263618 262782 263854
rect 262226 263298 262462 263534
rect 262546 263298 262782 263534
rect 262226 226418 262462 226654
rect 262546 226418 262782 226654
rect 262226 226098 262462 226334
rect 262546 226098 262782 226334
rect 262226 189218 262462 189454
rect 262546 189218 262782 189454
rect 262226 188898 262462 189134
rect 262546 188898 262782 189134
rect 262226 152018 262462 152254
rect 262546 152018 262782 152254
rect 262226 151698 262462 151934
rect 262546 151698 262782 151934
rect 262226 114818 262462 115054
rect 262546 114818 262782 115054
rect 262226 114498 262462 114734
rect 262546 114498 262782 114734
rect 262226 77618 262462 77854
rect 262546 77618 262782 77854
rect 262226 77298 262462 77534
rect 262546 77298 262782 77534
rect 262226 40418 262462 40654
rect 262546 40418 262782 40654
rect 262226 40098 262462 40334
rect 262546 40098 262782 40334
rect 262226 3218 262462 3454
rect 262546 3218 262782 3454
rect 262226 2898 262462 3134
rect 262546 2898 262782 3134
rect 265946 676538 266182 676774
rect 266266 676538 266502 676774
rect 265946 676218 266182 676454
rect 266266 676218 266502 676454
rect 265946 639338 266182 639574
rect 266266 639338 266502 639574
rect 265946 639018 266182 639254
rect 266266 639018 266502 639254
rect 265946 602138 266182 602374
rect 266266 602138 266502 602374
rect 265946 601818 266182 602054
rect 266266 601818 266502 602054
rect 265946 564938 266182 565174
rect 266266 564938 266502 565174
rect 265946 564618 266182 564854
rect 266266 564618 266502 564854
rect 265946 527738 266182 527974
rect 266266 527738 266502 527974
rect 265946 527418 266182 527654
rect 266266 527418 266502 527654
rect 265946 490538 266182 490774
rect 266266 490538 266502 490774
rect 265946 490218 266182 490454
rect 266266 490218 266502 490454
rect 265946 453338 266182 453574
rect 266266 453338 266502 453574
rect 265946 453018 266182 453254
rect 266266 453018 266502 453254
rect 265946 416138 266182 416374
rect 266266 416138 266502 416374
rect 265946 415818 266182 416054
rect 266266 415818 266502 416054
rect 265946 378938 266182 379174
rect 266266 378938 266502 379174
rect 265946 378618 266182 378854
rect 266266 378618 266502 378854
rect 265946 341738 266182 341974
rect 266266 341738 266502 341974
rect 265946 341418 266182 341654
rect 266266 341418 266502 341654
rect 265946 304538 266182 304774
rect 266266 304538 266502 304774
rect 265946 304218 266182 304454
rect 266266 304218 266502 304454
rect 265946 267338 266182 267574
rect 266266 267338 266502 267574
rect 265946 267018 266182 267254
rect 266266 267018 266502 267254
rect 265946 230138 266182 230374
rect 266266 230138 266502 230374
rect 265946 229818 266182 230054
rect 266266 229818 266502 230054
rect 265946 192938 266182 193174
rect 266266 192938 266502 193174
rect 265946 192618 266182 192854
rect 266266 192618 266502 192854
rect 265946 155738 266182 155974
rect 266266 155738 266502 155974
rect 265946 155418 266182 155654
rect 266266 155418 266502 155654
rect 265946 118538 266182 118774
rect 266266 118538 266502 118774
rect 265946 118218 266182 118454
rect 266266 118218 266502 118454
rect 265946 81338 266182 81574
rect 266266 81338 266502 81574
rect 265946 81018 266182 81254
rect 266266 81018 266502 81254
rect 265946 44138 266182 44374
rect 266266 44138 266502 44374
rect 265946 43818 266182 44054
rect 266266 43818 266502 44054
rect 265946 6938 266182 7174
rect 266266 6938 266502 7174
rect 265946 6618 266182 6854
rect 266266 6618 266502 6854
rect 269666 680258 269902 680494
rect 269986 680258 270222 680494
rect 269666 679938 269902 680174
rect 269986 679938 270222 680174
rect 269666 643058 269902 643294
rect 269986 643058 270222 643294
rect 269666 642738 269902 642974
rect 269986 642738 270222 642974
rect 269666 605858 269902 606094
rect 269986 605858 270222 606094
rect 269666 605538 269902 605774
rect 269986 605538 270222 605774
rect 269666 568658 269902 568894
rect 269986 568658 270222 568894
rect 269666 568338 269902 568574
rect 269986 568338 270222 568574
rect 269666 531458 269902 531694
rect 269986 531458 270222 531694
rect 269666 531138 269902 531374
rect 269986 531138 270222 531374
rect 269666 494258 269902 494494
rect 269986 494258 270222 494494
rect 269666 493938 269902 494174
rect 269986 493938 270222 494174
rect 269666 457058 269902 457294
rect 269986 457058 270222 457294
rect 269666 456738 269902 456974
rect 269986 456738 270222 456974
rect 269666 419858 269902 420094
rect 269986 419858 270222 420094
rect 269666 419538 269902 419774
rect 269986 419538 270222 419774
rect 269666 382658 269902 382894
rect 269986 382658 270222 382894
rect 269666 382338 269902 382574
rect 269986 382338 270222 382574
rect 269666 345458 269902 345694
rect 269986 345458 270222 345694
rect 269666 345138 269902 345374
rect 269986 345138 270222 345374
rect 269666 308258 269902 308494
rect 269986 308258 270222 308494
rect 269666 307938 269902 308174
rect 269986 307938 270222 308174
rect 269666 271058 269902 271294
rect 269986 271058 270222 271294
rect 269666 270738 269902 270974
rect 269986 270738 270222 270974
rect 269666 233858 269902 234094
rect 269986 233858 270222 234094
rect 269666 233538 269902 233774
rect 269986 233538 270222 233774
rect 269666 196658 269902 196894
rect 269986 196658 270222 196894
rect 269666 196338 269902 196574
rect 269986 196338 270222 196574
rect 269666 159458 269902 159694
rect 269986 159458 270222 159694
rect 269666 159138 269902 159374
rect 269986 159138 270222 159374
rect 269666 122258 269902 122494
rect 269986 122258 270222 122494
rect 269666 121938 269902 122174
rect 269986 121938 270222 122174
rect 269666 85058 269902 85294
rect 269986 85058 270222 85294
rect 269666 84738 269902 84974
rect 269986 84738 270222 84974
rect 269666 47858 269902 48094
rect 269986 47858 270222 48094
rect 269666 47538 269902 47774
rect 269986 47538 270222 47774
rect 269666 10658 269902 10894
rect 269986 10658 270222 10894
rect 269666 10338 269902 10574
rect 269986 10338 270222 10574
rect 273386 683978 273622 684214
rect 273706 683978 273942 684214
rect 273386 683658 273622 683894
rect 273706 683658 273942 683894
rect 273386 646778 273622 647014
rect 273706 646778 273942 647014
rect 273386 646458 273622 646694
rect 273706 646458 273942 646694
rect 273386 609578 273622 609814
rect 273706 609578 273942 609814
rect 273386 609258 273622 609494
rect 273706 609258 273942 609494
rect 273386 572378 273622 572614
rect 273706 572378 273942 572614
rect 273386 572058 273622 572294
rect 273706 572058 273942 572294
rect 273386 535178 273622 535414
rect 273706 535178 273942 535414
rect 273386 534858 273622 535094
rect 273706 534858 273942 535094
rect 273386 497978 273622 498214
rect 273706 497978 273942 498214
rect 273386 497658 273622 497894
rect 273706 497658 273942 497894
rect 273386 460778 273622 461014
rect 273706 460778 273942 461014
rect 273386 460458 273622 460694
rect 273706 460458 273942 460694
rect 273386 423578 273622 423814
rect 273706 423578 273942 423814
rect 273386 423258 273622 423494
rect 273706 423258 273942 423494
rect 273386 386378 273622 386614
rect 273706 386378 273942 386614
rect 273386 386058 273622 386294
rect 273706 386058 273942 386294
rect 273386 349178 273622 349414
rect 273706 349178 273942 349414
rect 273386 348858 273622 349094
rect 273706 348858 273942 349094
rect 273386 311978 273622 312214
rect 273706 311978 273942 312214
rect 273386 311658 273622 311894
rect 273706 311658 273942 311894
rect 273386 274778 273622 275014
rect 273706 274778 273942 275014
rect 273386 274458 273622 274694
rect 273706 274458 273942 274694
rect 273386 237578 273622 237814
rect 273706 237578 273942 237814
rect 273386 237258 273622 237494
rect 273706 237258 273942 237494
rect 273386 200378 273622 200614
rect 273706 200378 273942 200614
rect 273386 200058 273622 200294
rect 273706 200058 273942 200294
rect 273386 163178 273622 163414
rect 273706 163178 273942 163414
rect 273386 162858 273622 163094
rect 273706 162858 273942 163094
rect 273386 125978 273622 126214
rect 273706 125978 273942 126214
rect 273386 125658 273622 125894
rect 273706 125658 273942 125894
rect 273386 88778 273622 89014
rect 273706 88778 273942 89014
rect 273386 88458 273622 88694
rect 273706 88458 273942 88694
rect 273386 51578 273622 51814
rect 273706 51578 273942 51814
rect 273386 51258 273622 51494
rect 273706 51258 273942 51494
rect 273386 14378 273622 14614
rect 273706 14378 273942 14614
rect 273386 14058 273622 14294
rect 273706 14058 273942 14294
rect 277106 687698 277342 687934
rect 277426 687698 277662 687934
rect 277106 687378 277342 687614
rect 277426 687378 277662 687614
rect 277106 650498 277342 650734
rect 277426 650498 277662 650734
rect 277106 650178 277342 650414
rect 277426 650178 277662 650414
rect 277106 613298 277342 613534
rect 277426 613298 277662 613534
rect 277106 612978 277342 613214
rect 277426 612978 277662 613214
rect 277106 576098 277342 576334
rect 277426 576098 277662 576334
rect 277106 575778 277342 576014
rect 277426 575778 277662 576014
rect 277106 538898 277342 539134
rect 277426 538898 277662 539134
rect 277106 538578 277342 538814
rect 277426 538578 277662 538814
rect 277106 501698 277342 501934
rect 277426 501698 277662 501934
rect 277106 501378 277342 501614
rect 277426 501378 277662 501614
rect 277106 464498 277342 464734
rect 277426 464498 277662 464734
rect 277106 464178 277342 464414
rect 277426 464178 277662 464414
rect 277106 427298 277342 427534
rect 277426 427298 277662 427534
rect 277106 426978 277342 427214
rect 277426 426978 277662 427214
rect 277106 390098 277342 390334
rect 277426 390098 277662 390334
rect 277106 389778 277342 390014
rect 277426 389778 277662 390014
rect 277106 352898 277342 353134
rect 277426 352898 277662 353134
rect 277106 352578 277342 352814
rect 277426 352578 277662 352814
rect 277106 315698 277342 315934
rect 277426 315698 277662 315934
rect 277106 315378 277342 315614
rect 277426 315378 277662 315614
rect 277106 278498 277342 278734
rect 277426 278498 277662 278734
rect 277106 278178 277342 278414
rect 277426 278178 277662 278414
rect 277106 241298 277342 241534
rect 277426 241298 277662 241534
rect 277106 240978 277342 241214
rect 277426 240978 277662 241214
rect 277106 204098 277342 204334
rect 277426 204098 277662 204334
rect 277106 203778 277342 204014
rect 277426 203778 277662 204014
rect 277106 166898 277342 167134
rect 277426 166898 277662 167134
rect 277106 166578 277342 166814
rect 277426 166578 277662 166814
rect 277106 129698 277342 129934
rect 277426 129698 277662 129934
rect 277106 129378 277342 129614
rect 277426 129378 277662 129614
rect 277106 92498 277342 92734
rect 277426 92498 277662 92734
rect 277106 92178 277342 92414
rect 277426 92178 277662 92414
rect 277106 55298 277342 55534
rect 277426 55298 277662 55534
rect 277106 54978 277342 55214
rect 277426 54978 277662 55214
rect 277106 18098 277342 18334
rect 277426 18098 277662 18334
rect 277106 17778 277342 18014
rect 277426 17778 277662 18014
rect 280826 691418 281062 691654
rect 281146 691418 281382 691654
rect 280826 691098 281062 691334
rect 281146 691098 281382 691334
rect 280826 654218 281062 654454
rect 281146 654218 281382 654454
rect 280826 653898 281062 654134
rect 281146 653898 281382 654134
rect 280826 617018 281062 617254
rect 281146 617018 281382 617254
rect 280826 616698 281062 616934
rect 281146 616698 281382 616934
rect 280826 579818 281062 580054
rect 281146 579818 281382 580054
rect 280826 579498 281062 579734
rect 281146 579498 281382 579734
rect 280826 542618 281062 542854
rect 281146 542618 281382 542854
rect 280826 542298 281062 542534
rect 281146 542298 281382 542534
rect 280826 505418 281062 505654
rect 281146 505418 281382 505654
rect 280826 505098 281062 505334
rect 281146 505098 281382 505334
rect 280826 468218 281062 468454
rect 281146 468218 281382 468454
rect 280826 467898 281062 468134
rect 281146 467898 281382 468134
rect 280826 431018 281062 431254
rect 281146 431018 281382 431254
rect 280826 430698 281062 430934
rect 281146 430698 281382 430934
rect 280826 393818 281062 394054
rect 281146 393818 281382 394054
rect 280826 393498 281062 393734
rect 281146 393498 281382 393734
rect 280826 356618 281062 356854
rect 281146 356618 281382 356854
rect 280826 356298 281062 356534
rect 281146 356298 281382 356534
rect 280826 319418 281062 319654
rect 281146 319418 281382 319654
rect 280826 319098 281062 319334
rect 281146 319098 281382 319334
rect 280826 282218 281062 282454
rect 281146 282218 281382 282454
rect 280826 281898 281062 282134
rect 281146 281898 281382 282134
rect 280826 245018 281062 245254
rect 281146 245018 281382 245254
rect 280826 244698 281062 244934
rect 281146 244698 281382 244934
rect 280826 207818 281062 208054
rect 281146 207818 281382 208054
rect 280826 207498 281062 207734
rect 281146 207498 281382 207734
rect 280826 170618 281062 170854
rect 281146 170618 281382 170854
rect 280826 170298 281062 170534
rect 281146 170298 281382 170534
rect 280826 133418 281062 133654
rect 281146 133418 281382 133654
rect 280826 133098 281062 133334
rect 281146 133098 281382 133334
rect 280826 96218 281062 96454
rect 281146 96218 281382 96454
rect 280826 95898 281062 96134
rect 281146 95898 281382 96134
rect 280826 59018 281062 59254
rect 281146 59018 281382 59254
rect 280826 58698 281062 58934
rect 281146 58698 281382 58934
rect 280826 21818 281062 22054
rect 281146 21818 281382 22054
rect 280826 21498 281062 21734
rect 281146 21498 281382 21734
rect 284546 695138 284782 695374
rect 284866 695138 285102 695374
rect 284546 694818 284782 695054
rect 284866 694818 285102 695054
rect 284546 657938 284782 658174
rect 284866 657938 285102 658174
rect 284546 657618 284782 657854
rect 284866 657618 285102 657854
rect 284546 620738 284782 620974
rect 284866 620738 285102 620974
rect 284546 620418 284782 620654
rect 284866 620418 285102 620654
rect 284546 583538 284782 583774
rect 284866 583538 285102 583774
rect 284546 583218 284782 583454
rect 284866 583218 285102 583454
rect 284546 546338 284782 546574
rect 284866 546338 285102 546574
rect 284546 546018 284782 546254
rect 284866 546018 285102 546254
rect 284546 509138 284782 509374
rect 284866 509138 285102 509374
rect 284546 508818 284782 509054
rect 284866 508818 285102 509054
rect 284546 471938 284782 472174
rect 284866 471938 285102 472174
rect 284546 471618 284782 471854
rect 284866 471618 285102 471854
rect 284546 434738 284782 434974
rect 284866 434738 285102 434974
rect 284546 434418 284782 434654
rect 284866 434418 285102 434654
rect 284546 397538 284782 397774
rect 284866 397538 285102 397774
rect 284546 397218 284782 397454
rect 284866 397218 285102 397454
rect 284546 360338 284782 360574
rect 284866 360338 285102 360574
rect 284546 360018 284782 360254
rect 284866 360018 285102 360254
rect 284546 323138 284782 323374
rect 284866 323138 285102 323374
rect 284546 322818 284782 323054
rect 284866 322818 285102 323054
rect 284546 285938 284782 286174
rect 284866 285938 285102 286174
rect 284546 285618 284782 285854
rect 284866 285618 285102 285854
rect 284546 248738 284782 248974
rect 284866 248738 285102 248974
rect 284546 248418 284782 248654
rect 284866 248418 285102 248654
rect 284546 211538 284782 211774
rect 284866 211538 285102 211774
rect 284546 211218 284782 211454
rect 284866 211218 285102 211454
rect 284546 174338 284782 174574
rect 284866 174338 285102 174574
rect 284546 174018 284782 174254
rect 284866 174018 285102 174254
rect 284546 137138 284782 137374
rect 284866 137138 285102 137374
rect 284546 136818 284782 137054
rect 284866 136818 285102 137054
rect 284546 99938 284782 100174
rect 284866 99938 285102 100174
rect 284546 99618 284782 99854
rect 284866 99618 285102 99854
rect 284546 62738 284782 62974
rect 284866 62738 285102 62974
rect 284546 62418 284782 62654
rect 284866 62418 285102 62654
rect 284546 25538 284782 25774
rect 284866 25538 285102 25774
rect 284546 25218 284782 25454
rect 284866 25218 285102 25454
rect 288266 698858 288502 699094
rect 288586 698858 288822 699094
rect 288266 698538 288502 698774
rect 288586 698538 288822 698774
rect 288266 661658 288502 661894
rect 288586 661658 288822 661894
rect 288266 661338 288502 661574
rect 288586 661338 288822 661574
rect 288266 624458 288502 624694
rect 288586 624458 288822 624694
rect 288266 624138 288502 624374
rect 288586 624138 288822 624374
rect 288266 587258 288502 587494
rect 288586 587258 288822 587494
rect 288266 586938 288502 587174
rect 288586 586938 288822 587174
rect 288266 550058 288502 550294
rect 288586 550058 288822 550294
rect 288266 549738 288502 549974
rect 288586 549738 288822 549974
rect 288266 512858 288502 513094
rect 288586 512858 288822 513094
rect 288266 512538 288502 512774
rect 288586 512538 288822 512774
rect 288266 475658 288502 475894
rect 288586 475658 288822 475894
rect 288266 475338 288502 475574
rect 288586 475338 288822 475574
rect 288266 438458 288502 438694
rect 288586 438458 288822 438694
rect 288266 438138 288502 438374
rect 288586 438138 288822 438374
rect 288266 401258 288502 401494
rect 288586 401258 288822 401494
rect 288266 400938 288502 401174
rect 288586 400938 288822 401174
rect 288266 364058 288502 364294
rect 288586 364058 288822 364294
rect 288266 363738 288502 363974
rect 288586 363738 288822 363974
rect 288266 326858 288502 327094
rect 288586 326858 288822 327094
rect 288266 326538 288502 326774
rect 288586 326538 288822 326774
rect 288266 289658 288502 289894
rect 288586 289658 288822 289894
rect 288266 289338 288502 289574
rect 288586 289338 288822 289574
rect 288266 252458 288502 252694
rect 288586 252458 288822 252694
rect 288266 252138 288502 252374
rect 288586 252138 288822 252374
rect 288266 215258 288502 215494
rect 288586 215258 288822 215494
rect 288266 214938 288502 215174
rect 288586 214938 288822 215174
rect 288266 178058 288502 178294
rect 288586 178058 288822 178294
rect 288266 177738 288502 177974
rect 288586 177738 288822 177974
rect 288266 140858 288502 141094
rect 288586 140858 288822 141094
rect 288266 140538 288502 140774
rect 288586 140538 288822 140774
rect 288266 103658 288502 103894
rect 288586 103658 288822 103894
rect 288266 103338 288502 103574
rect 288586 103338 288822 103574
rect 288266 66458 288502 66694
rect 288586 66458 288822 66694
rect 288266 66138 288502 66374
rect 288586 66138 288822 66374
rect 288266 29258 288502 29494
rect 288586 29258 288822 29494
rect 288266 28938 288502 29174
rect 288586 28938 288822 29174
rect 299426 672818 299662 673054
rect 299746 672818 299982 673054
rect 299426 672498 299662 672734
rect 299746 672498 299982 672734
rect 299426 635618 299662 635854
rect 299746 635618 299982 635854
rect 299426 635298 299662 635534
rect 299746 635298 299982 635534
rect 299426 598418 299662 598654
rect 299746 598418 299982 598654
rect 299426 598098 299662 598334
rect 299746 598098 299982 598334
rect 299426 561218 299662 561454
rect 299746 561218 299982 561454
rect 299426 560898 299662 561134
rect 299746 560898 299982 561134
rect 299426 524018 299662 524254
rect 299746 524018 299982 524254
rect 299426 523698 299662 523934
rect 299746 523698 299982 523934
rect 299426 486818 299662 487054
rect 299746 486818 299982 487054
rect 299426 486498 299662 486734
rect 299746 486498 299982 486734
rect 299426 449618 299662 449854
rect 299746 449618 299982 449854
rect 299426 449298 299662 449534
rect 299746 449298 299982 449534
rect 299426 412418 299662 412654
rect 299746 412418 299982 412654
rect 299426 412098 299662 412334
rect 299746 412098 299982 412334
rect 299426 375218 299662 375454
rect 299746 375218 299982 375454
rect 299426 374898 299662 375134
rect 299746 374898 299982 375134
rect 299426 338018 299662 338254
rect 299746 338018 299982 338254
rect 299426 337698 299662 337934
rect 299746 337698 299982 337934
rect 299426 300818 299662 301054
rect 299746 300818 299982 301054
rect 299426 300498 299662 300734
rect 299746 300498 299982 300734
rect 299426 263618 299662 263854
rect 299746 263618 299982 263854
rect 299426 263298 299662 263534
rect 299746 263298 299982 263534
rect 299426 226418 299662 226654
rect 299746 226418 299982 226654
rect 299426 226098 299662 226334
rect 299746 226098 299982 226334
rect 299426 189218 299662 189454
rect 299746 189218 299982 189454
rect 299426 188898 299662 189134
rect 299746 188898 299982 189134
rect 299426 152018 299662 152254
rect 299746 152018 299982 152254
rect 299426 151698 299662 151934
rect 299746 151698 299982 151934
rect 299426 114818 299662 115054
rect 299746 114818 299982 115054
rect 299426 114498 299662 114734
rect 299746 114498 299982 114734
rect 299426 77618 299662 77854
rect 299746 77618 299982 77854
rect 299426 77298 299662 77534
rect 299746 77298 299982 77534
rect 299426 40418 299662 40654
rect 299746 40418 299982 40654
rect 299426 40098 299662 40334
rect 299746 40098 299982 40334
rect 299426 3218 299662 3454
rect 299746 3218 299982 3454
rect 299426 2898 299662 3134
rect 299746 2898 299982 3134
rect 303146 676538 303382 676774
rect 303466 676538 303702 676774
rect 303146 676218 303382 676454
rect 303466 676218 303702 676454
rect 303146 639338 303382 639574
rect 303466 639338 303702 639574
rect 303146 639018 303382 639254
rect 303466 639018 303702 639254
rect 303146 602138 303382 602374
rect 303466 602138 303702 602374
rect 303146 601818 303382 602054
rect 303466 601818 303702 602054
rect 303146 564938 303382 565174
rect 303466 564938 303702 565174
rect 303146 564618 303382 564854
rect 303466 564618 303702 564854
rect 303146 527738 303382 527974
rect 303466 527738 303702 527974
rect 303146 527418 303382 527654
rect 303466 527418 303702 527654
rect 303146 490538 303382 490774
rect 303466 490538 303702 490774
rect 303146 490218 303382 490454
rect 303466 490218 303702 490454
rect 303146 453338 303382 453574
rect 303466 453338 303702 453574
rect 303146 453018 303382 453254
rect 303466 453018 303702 453254
rect 303146 416138 303382 416374
rect 303466 416138 303702 416374
rect 303146 415818 303382 416054
rect 303466 415818 303702 416054
rect 303146 378938 303382 379174
rect 303466 378938 303702 379174
rect 303146 378618 303382 378854
rect 303466 378618 303702 378854
rect 303146 341738 303382 341974
rect 303466 341738 303702 341974
rect 303146 341418 303382 341654
rect 303466 341418 303702 341654
rect 303146 304538 303382 304774
rect 303466 304538 303702 304774
rect 303146 304218 303382 304454
rect 303466 304218 303702 304454
rect 303146 267338 303382 267574
rect 303466 267338 303702 267574
rect 303146 267018 303382 267254
rect 303466 267018 303702 267254
rect 303146 230138 303382 230374
rect 303466 230138 303702 230374
rect 303146 229818 303382 230054
rect 303466 229818 303702 230054
rect 303146 192938 303382 193174
rect 303466 192938 303702 193174
rect 303146 192618 303382 192854
rect 303466 192618 303702 192854
rect 303146 155738 303382 155974
rect 303466 155738 303702 155974
rect 303146 155418 303382 155654
rect 303466 155418 303702 155654
rect 303146 118538 303382 118774
rect 303466 118538 303702 118774
rect 303146 118218 303382 118454
rect 303466 118218 303702 118454
rect 303146 81338 303382 81574
rect 303466 81338 303702 81574
rect 303146 81018 303382 81254
rect 303466 81018 303702 81254
rect 303146 44138 303382 44374
rect 303466 44138 303702 44374
rect 303146 43818 303382 44054
rect 303466 43818 303702 44054
rect 303146 6938 303382 7174
rect 303466 6938 303702 7174
rect 303146 6618 303382 6854
rect 303466 6618 303702 6854
rect 306866 680258 307102 680494
rect 307186 680258 307422 680494
rect 306866 679938 307102 680174
rect 307186 679938 307422 680174
rect 306866 643058 307102 643294
rect 307186 643058 307422 643294
rect 306866 642738 307102 642974
rect 307186 642738 307422 642974
rect 306866 605858 307102 606094
rect 307186 605858 307422 606094
rect 306866 605538 307102 605774
rect 307186 605538 307422 605774
rect 306866 568658 307102 568894
rect 307186 568658 307422 568894
rect 306866 568338 307102 568574
rect 307186 568338 307422 568574
rect 306866 531458 307102 531694
rect 307186 531458 307422 531694
rect 306866 531138 307102 531374
rect 307186 531138 307422 531374
rect 306866 494258 307102 494494
rect 307186 494258 307422 494494
rect 306866 493938 307102 494174
rect 307186 493938 307422 494174
rect 306866 457058 307102 457294
rect 307186 457058 307422 457294
rect 306866 456738 307102 456974
rect 307186 456738 307422 456974
rect 306866 419858 307102 420094
rect 307186 419858 307422 420094
rect 306866 419538 307102 419774
rect 307186 419538 307422 419774
rect 306866 382658 307102 382894
rect 307186 382658 307422 382894
rect 306866 382338 307102 382574
rect 307186 382338 307422 382574
rect 306866 345458 307102 345694
rect 307186 345458 307422 345694
rect 306866 345138 307102 345374
rect 307186 345138 307422 345374
rect 306866 308258 307102 308494
rect 307186 308258 307422 308494
rect 306866 307938 307102 308174
rect 307186 307938 307422 308174
rect 306866 271058 307102 271294
rect 307186 271058 307422 271294
rect 306866 270738 307102 270974
rect 307186 270738 307422 270974
rect 306866 233858 307102 234094
rect 307186 233858 307422 234094
rect 306866 233538 307102 233774
rect 307186 233538 307422 233774
rect 306866 196658 307102 196894
rect 307186 196658 307422 196894
rect 306866 196338 307102 196574
rect 307186 196338 307422 196574
rect 306866 159458 307102 159694
rect 307186 159458 307422 159694
rect 306866 159138 307102 159374
rect 307186 159138 307422 159374
rect 306866 122258 307102 122494
rect 307186 122258 307422 122494
rect 306866 121938 307102 122174
rect 307186 121938 307422 122174
rect 306866 85058 307102 85294
rect 307186 85058 307422 85294
rect 306866 84738 307102 84974
rect 307186 84738 307422 84974
rect 306866 47858 307102 48094
rect 307186 47858 307422 48094
rect 306866 47538 307102 47774
rect 307186 47538 307422 47774
rect 306866 10658 307102 10894
rect 307186 10658 307422 10894
rect 306866 10338 307102 10574
rect 307186 10338 307422 10574
rect 310586 683978 310822 684214
rect 310906 683978 311142 684214
rect 310586 683658 310822 683894
rect 310906 683658 311142 683894
rect 310586 646778 310822 647014
rect 310906 646778 311142 647014
rect 310586 646458 310822 646694
rect 310906 646458 311142 646694
rect 310586 609578 310822 609814
rect 310906 609578 311142 609814
rect 310586 609258 310822 609494
rect 310906 609258 311142 609494
rect 310586 572378 310822 572614
rect 310906 572378 311142 572614
rect 310586 572058 310822 572294
rect 310906 572058 311142 572294
rect 310586 535178 310822 535414
rect 310906 535178 311142 535414
rect 310586 534858 310822 535094
rect 310906 534858 311142 535094
rect 310586 497978 310822 498214
rect 310906 497978 311142 498214
rect 310586 497658 310822 497894
rect 310906 497658 311142 497894
rect 310586 460778 310822 461014
rect 310906 460778 311142 461014
rect 310586 460458 310822 460694
rect 310906 460458 311142 460694
rect 310586 423578 310822 423814
rect 310906 423578 311142 423814
rect 310586 423258 310822 423494
rect 310906 423258 311142 423494
rect 310586 386378 310822 386614
rect 310906 386378 311142 386614
rect 310586 386058 310822 386294
rect 310906 386058 311142 386294
rect 310586 349178 310822 349414
rect 310906 349178 311142 349414
rect 310586 348858 310822 349094
rect 310906 348858 311142 349094
rect 310586 311978 310822 312214
rect 310906 311978 311142 312214
rect 310586 311658 310822 311894
rect 310906 311658 311142 311894
rect 310586 274778 310822 275014
rect 310906 274778 311142 275014
rect 310586 274458 310822 274694
rect 310906 274458 311142 274694
rect 310586 237578 310822 237814
rect 310906 237578 311142 237814
rect 310586 237258 310822 237494
rect 310906 237258 311142 237494
rect 310586 200378 310822 200614
rect 310906 200378 311142 200614
rect 310586 200058 310822 200294
rect 310906 200058 311142 200294
rect 310586 163178 310822 163414
rect 310906 163178 311142 163414
rect 310586 162858 310822 163094
rect 310906 162858 311142 163094
rect 310586 125978 310822 126214
rect 310906 125978 311142 126214
rect 310586 125658 310822 125894
rect 310906 125658 311142 125894
rect 310586 88778 310822 89014
rect 310906 88778 311142 89014
rect 310586 88458 310822 88694
rect 310906 88458 311142 88694
rect 310586 51578 310822 51814
rect 310906 51578 311142 51814
rect 310586 51258 310822 51494
rect 310906 51258 311142 51494
rect 310586 14378 310822 14614
rect 310906 14378 311142 14614
rect 310586 14058 310822 14294
rect 310906 14058 311142 14294
rect 314306 687698 314542 687934
rect 314626 687698 314862 687934
rect 314306 687378 314542 687614
rect 314626 687378 314862 687614
rect 314306 650498 314542 650734
rect 314626 650498 314862 650734
rect 314306 650178 314542 650414
rect 314626 650178 314862 650414
rect 314306 613298 314542 613534
rect 314626 613298 314862 613534
rect 314306 612978 314542 613214
rect 314626 612978 314862 613214
rect 314306 576098 314542 576334
rect 314626 576098 314862 576334
rect 314306 575778 314542 576014
rect 314626 575778 314862 576014
rect 314306 538898 314542 539134
rect 314626 538898 314862 539134
rect 314306 538578 314542 538814
rect 314626 538578 314862 538814
rect 314306 501698 314542 501934
rect 314626 501698 314862 501934
rect 314306 501378 314542 501614
rect 314626 501378 314862 501614
rect 314306 464498 314542 464734
rect 314626 464498 314862 464734
rect 314306 464178 314542 464414
rect 314626 464178 314862 464414
rect 314306 427298 314542 427534
rect 314626 427298 314862 427534
rect 314306 426978 314542 427214
rect 314626 426978 314862 427214
rect 314306 390098 314542 390334
rect 314626 390098 314862 390334
rect 314306 389778 314542 390014
rect 314626 389778 314862 390014
rect 314306 352898 314542 353134
rect 314626 352898 314862 353134
rect 314306 352578 314542 352814
rect 314626 352578 314862 352814
rect 314306 315698 314542 315934
rect 314626 315698 314862 315934
rect 314306 315378 314542 315614
rect 314626 315378 314862 315614
rect 314306 278498 314542 278734
rect 314626 278498 314862 278734
rect 314306 278178 314542 278414
rect 314626 278178 314862 278414
rect 314306 241298 314542 241534
rect 314626 241298 314862 241534
rect 314306 240978 314542 241214
rect 314626 240978 314862 241214
rect 314306 204098 314542 204334
rect 314626 204098 314862 204334
rect 314306 203778 314542 204014
rect 314626 203778 314862 204014
rect 314306 166898 314542 167134
rect 314626 166898 314862 167134
rect 314306 166578 314542 166814
rect 314626 166578 314862 166814
rect 314306 129698 314542 129934
rect 314626 129698 314862 129934
rect 314306 129378 314542 129614
rect 314626 129378 314862 129614
rect 314306 92498 314542 92734
rect 314626 92498 314862 92734
rect 314306 92178 314542 92414
rect 314626 92178 314862 92414
rect 314306 55298 314542 55534
rect 314626 55298 314862 55534
rect 314306 54978 314542 55214
rect 314626 54978 314862 55214
rect 314306 18098 314542 18334
rect 314626 18098 314862 18334
rect 314306 17778 314542 18014
rect 314626 17778 314862 18014
rect 318026 691418 318262 691654
rect 318346 691418 318582 691654
rect 318026 691098 318262 691334
rect 318346 691098 318582 691334
rect 318026 654218 318262 654454
rect 318346 654218 318582 654454
rect 318026 653898 318262 654134
rect 318346 653898 318582 654134
rect 318026 617018 318262 617254
rect 318346 617018 318582 617254
rect 318026 616698 318262 616934
rect 318346 616698 318582 616934
rect 318026 579818 318262 580054
rect 318346 579818 318582 580054
rect 318026 579498 318262 579734
rect 318346 579498 318582 579734
rect 318026 542618 318262 542854
rect 318346 542618 318582 542854
rect 318026 542298 318262 542534
rect 318346 542298 318582 542534
rect 318026 505418 318262 505654
rect 318346 505418 318582 505654
rect 318026 505098 318262 505334
rect 318346 505098 318582 505334
rect 318026 468218 318262 468454
rect 318346 468218 318582 468454
rect 318026 467898 318262 468134
rect 318346 467898 318582 468134
rect 318026 431018 318262 431254
rect 318346 431018 318582 431254
rect 318026 430698 318262 430934
rect 318346 430698 318582 430934
rect 318026 393818 318262 394054
rect 318346 393818 318582 394054
rect 318026 393498 318262 393734
rect 318346 393498 318582 393734
rect 318026 356618 318262 356854
rect 318346 356618 318582 356854
rect 318026 356298 318262 356534
rect 318346 356298 318582 356534
rect 318026 319418 318262 319654
rect 318346 319418 318582 319654
rect 318026 319098 318262 319334
rect 318346 319098 318582 319334
rect 318026 282218 318262 282454
rect 318346 282218 318582 282454
rect 318026 281898 318262 282134
rect 318346 281898 318582 282134
rect 318026 245018 318262 245254
rect 318346 245018 318582 245254
rect 318026 244698 318262 244934
rect 318346 244698 318582 244934
rect 318026 207818 318262 208054
rect 318346 207818 318582 208054
rect 318026 207498 318262 207734
rect 318346 207498 318582 207734
rect 318026 170618 318262 170854
rect 318346 170618 318582 170854
rect 318026 170298 318262 170534
rect 318346 170298 318582 170534
rect 318026 133418 318262 133654
rect 318346 133418 318582 133654
rect 318026 133098 318262 133334
rect 318346 133098 318582 133334
rect 318026 96218 318262 96454
rect 318346 96218 318582 96454
rect 318026 95898 318262 96134
rect 318346 95898 318582 96134
rect 318026 59018 318262 59254
rect 318346 59018 318582 59254
rect 318026 58698 318262 58934
rect 318346 58698 318582 58934
rect 318026 21818 318262 22054
rect 318346 21818 318582 22054
rect 318026 21498 318262 21734
rect 318346 21498 318582 21734
rect 321746 695138 321982 695374
rect 322066 695138 322302 695374
rect 321746 694818 321982 695054
rect 322066 694818 322302 695054
rect 321746 657938 321982 658174
rect 322066 657938 322302 658174
rect 321746 657618 321982 657854
rect 322066 657618 322302 657854
rect 321746 620738 321982 620974
rect 322066 620738 322302 620974
rect 321746 620418 321982 620654
rect 322066 620418 322302 620654
rect 321746 583538 321982 583774
rect 322066 583538 322302 583774
rect 321746 583218 321982 583454
rect 322066 583218 322302 583454
rect 321746 546338 321982 546574
rect 322066 546338 322302 546574
rect 321746 546018 321982 546254
rect 322066 546018 322302 546254
rect 321746 509138 321982 509374
rect 322066 509138 322302 509374
rect 321746 508818 321982 509054
rect 322066 508818 322302 509054
rect 321746 471938 321982 472174
rect 322066 471938 322302 472174
rect 321746 471618 321982 471854
rect 322066 471618 322302 471854
rect 321746 434738 321982 434974
rect 322066 434738 322302 434974
rect 321746 434418 321982 434654
rect 322066 434418 322302 434654
rect 321746 397538 321982 397774
rect 322066 397538 322302 397774
rect 321746 397218 321982 397454
rect 322066 397218 322302 397454
rect 321746 360338 321982 360574
rect 322066 360338 322302 360574
rect 321746 360018 321982 360254
rect 322066 360018 322302 360254
rect 321746 323138 321982 323374
rect 322066 323138 322302 323374
rect 321746 322818 321982 323054
rect 322066 322818 322302 323054
rect 321746 285938 321982 286174
rect 322066 285938 322302 286174
rect 321746 285618 321982 285854
rect 322066 285618 322302 285854
rect 321746 248738 321982 248974
rect 322066 248738 322302 248974
rect 321746 248418 321982 248654
rect 322066 248418 322302 248654
rect 321746 211538 321982 211774
rect 322066 211538 322302 211774
rect 321746 211218 321982 211454
rect 322066 211218 322302 211454
rect 321746 174338 321982 174574
rect 322066 174338 322302 174574
rect 321746 174018 321982 174254
rect 322066 174018 322302 174254
rect 321746 137138 321982 137374
rect 322066 137138 322302 137374
rect 321746 136818 321982 137054
rect 322066 136818 322302 137054
rect 321746 99938 321982 100174
rect 322066 99938 322302 100174
rect 321746 99618 321982 99854
rect 322066 99618 322302 99854
rect 321746 62738 321982 62974
rect 322066 62738 322302 62974
rect 321746 62418 321982 62654
rect 322066 62418 322302 62654
rect 321746 25538 321982 25774
rect 322066 25538 322302 25774
rect 321746 25218 321982 25454
rect 322066 25218 322302 25454
rect 325466 698858 325702 699094
rect 325786 698858 326022 699094
rect 325466 698538 325702 698774
rect 325786 698538 326022 698774
rect 325466 661658 325702 661894
rect 325786 661658 326022 661894
rect 325466 661338 325702 661574
rect 325786 661338 326022 661574
rect 325466 624458 325702 624694
rect 325786 624458 326022 624694
rect 325466 624138 325702 624374
rect 325786 624138 326022 624374
rect 325466 587258 325702 587494
rect 325786 587258 326022 587494
rect 325466 586938 325702 587174
rect 325786 586938 326022 587174
rect 325466 550058 325702 550294
rect 325786 550058 326022 550294
rect 325466 549738 325702 549974
rect 325786 549738 326022 549974
rect 325466 512858 325702 513094
rect 325786 512858 326022 513094
rect 325466 512538 325702 512774
rect 325786 512538 326022 512774
rect 325466 475658 325702 475894
rect 325786 475658 326022 475894
rect 325466 475338 325702 475574
rect 325786 475338 326022 475574
rect 325466 438458 325702 438694
rect 325786 438458 326022 438694
rect 325466 438138 325702 438374
rect 325786 438138 326022 438374
rect 325466 401258 325702 401494
rect 325786 401258 326022 401494
rect 325466 400938 325702 401174
rect 325786 400938 326022 401174
rect 325466 364058 325702 364294
rect 325786 364058 326022 364294
rect 325466 363738 325702 363974
rect 325786 363738 326022 363974
rect 325466 326858 325702 327094
rect 325786 326858 326022 327094
rect 325466 326538 325702 326774
rect 325786 326538 326022 326774
rect 325466 289658 325702 289894
rect 325786 289658 326022 289894
rect 325466 289338 325702 289574
rect 325786 289338 326022 289574
rect 325466 252458 325702 252694
rect 325786 252458 326022 252694
rect 325466 252138 325702 252374
rect 325786 252138 326022 252374
rect 325466 215258 325702 215494
rect 325786 215258 326022 215494
rect 325466 214938 325702 215174
rect 325786 214938 326022 215174
rect 325466 178058 325702 178294
rect 325786 178058 326022 178294
rect 325466 177738 325702 177974
rect 325786 177738 326022 177974
rect 325466 140858 325702 141094
rect 325786 140858 326022 141094
rect 325466 140538 325702 140774
rect 325786 140538 326022 140774
rect 325466 103658 325702 103894
rect 325786 103658 326022 103894
rect 325466 103338 325702 103574
rect 325786 103338 326022 103574
rect 325466 66458 325702 66694
rect 325786 66458 326022 66694
rect 325466 66138 325702 66374
rect 325786 66138 326022 66374
rect 325466 29258 325702 29494
rect 325786 29258 326022 29494
rect 325466 28938 325702 29174
rect 325786 28938 326022 29174
rect 336626 672818 336862 673054
rect 336946 672818 337182 673054
rect 336626 672498 336862 672734
rect 336946 672498 337182 672734
rect 336626 635618 336862 635854
rect 336946 635618 337182 635854
rect 336626 635298 336862 635534
rect 336946 635298 337182 635534
rect 336626 598418 336862 598654
rect 336946 598418 337182 598654
rect 336626 598098 336862 598334
rect 336946 598098 337182 598334
rect 336626 561218 336862 561454
rect 336946 561218 337182 561454
rect 336626 560898 336862 561134
rect 336946 560898 337182 561134
rect 336626 524018 336862 524254
rect 336946 524018 337182 524254
rect 336626 523698 336862 523934
rect 336946 523698 337182 523934
rect 336626 486818 336862 487054
rect 336946 486818 337182 487054
rect 336626 486498 336862 486734
rect 336946 486498 337182 486734
rect 336626 449618 336862 449854
rect 336946 449618 337182 449854
rect 336626 449298 336862 449534
rect 336946 449298 337182 449534
rect 336626 412418 336862 412654
rect 336946 412418 337182 412654
rect 336626 412098 336862 412334
rect 336946 412098 337182 412334
rect 336626 375218 336862 375454
rect 336946 375218 337182 375454
rect 336626 374898 336862 375134
rect 336946 374898 337182 375134
rect 336626 338018 336862 338254
rect 336946 338018 337182 338254
rect 336626 337698 336862 337934
rect 336946 337698 337182 337934
rect 336626 300818 336862 301054
rect 336946 300818 337182 301054
rect 336626 300498 336862 300734
rect 336946 300498 337182 300734
rect 336626 263618 336862 263854
rect 336946 263618 337182 263854
rect 336626 263298 336862 263534
rect 336946 263298 337182 263534
rect 336626 226418 336862 226654
rect 336946 226418 337182 226654
rect 336626 226098 336862 226334
rect 336946 226098 337182 226334
rect 336626 189218 336862 189454
rect 336946 189218 337182 189454
rect 336626 188898 336862 189134
rect 336946 188898 337182 189134
rect 336626 152018 336862 152254
rect 336946 152018 337182 152254
rect 336626 151698 336862 151934
rect 336946 151698 337182 151934
rect 336626 114818 336862 115054
rect 336946 114818 337182 115054
rect 336626 114498 336862 114734
rect 336946 114498 337182 114734
rect 336626 77618 336862 77854
rect 336946 77618 337182 77854
rect 336626 77298 336862 77534
rect 336946 77298 337182 77534
rect 336626 40418 336862 40654
rect 336946 40418 337182 40654
rect 336626 40098 336862 40334
rect 336946 40098 337182 40334
rect 336626 3218 336862 3454
rect 336946 3218 337182 3454
rect 336626 2898 336862 3134
rect 336946 2898 337182 3134
rect 340346 676538 340582 676774
rect 340666 676538 340902 676774
rect 340346 676218 340582 676454
rect 340666 676218 340902 676454
rect 340346 639338 340582 639574
rect 340666 639338 340902 639574
rect 340346 639018 340582 639254
rect 340666 639018 340902 639254
rect 340346 602138 340582 602374
rect 340666 602138 340902 602374
rect 340346 601818 340582 602054
rect 340666 601818 340902 602054
rect 340346 564938 340582 565174
rect 340666 564938 340902 565174
rect 340346 564618 340582 564854
rect 340666 564618 340902 564854
rect 340346 527738 340582 527974
rect 340666 527738 340902 527974
rect 340346 527418 340582 527654
rect 340666 527418 340902 527654
rect 340346 490538 340582 490774
rect 340666 490538 340902 490774
rect 340346 490218 340582 490454
rect 340666 490218 340902 490454
rect 340346 453338 340582 453574
rect 340666 453338 340902 453574
rect 340346 453018 340582 453254
rect 340666 453018 340902 453254
rect 340346 416138 340582 416374
rect 340666 416138 340902 416374
rect 340346 415818 340582 416054
rect 340666 415818 340902 416054
rect 340346 378938 340582 379174
rect 340666 378938 340902 379174
rect 340346 378618 340582 378854
rect 340666 378618 340902 378854
rect 340346 341738 340582 341974
rect 340666 341738 340902 341974
rect 340346 341418 340582 341654
rect 340666 341418 340902 341654
rect 340346 304538 340582 304774
rect 340666 304538 340902 304774
rect 340346 304218 340582 304454
rect 340666 304218 340902 304454
rect 340346 267338 340582 267574
rect 340666 267338 340902 267574
rect 340346 267018 340582 267254
rect 340666 267018 340902 267254
rect 340346 230138 340582 230374
rect 340666 230138 340902 230374
rect 340346 229818 340582 230054
rect 340666 229818 340902 230054
rect 340346 192938 340582 193174
rect 340666 192938 340902 193174
rect 340346 192618 340582 192854
rect 340666 192618 340902 192854
rect 340346 155738 340582 155974
rect 340666 155738 340902 155974
rect 340346 155418 340582 155654
rect 340666 155418 340902 155654
rect 340346 118538 340582 118774
rect 340666 118538 340902 118774
rect 340346 118218 340582 118454
rect 340666 118218 340902 118454
rect 340346 81338 340582 81574
rect 340666 81338 340902 81574
rect 340346 81018 340582 81254
rect 340666 81018 340902 81254
rect 340346 44138 340582 44374
rect 340666 44138 340902 44374
rect 340346 43818 340582 44054
rect 340666 43818 340902 44054
rect 340346 6938 340582 7174
rect 340666 6938 340902 7174
rect 340346 6618 340582 6854
rect 340666 6618 340902 6854
rect 344066 680258 344302 680494
rect 344386 680258 344622 680494
rect 344066 679938 344302 680174
rect 344386 679938 344622 680174
rect 344066 643058 344302 643294
rect 344386 643058 344622 643294
rect 344066 642738 344302 642974
rect 344386 642738 344622 642974
rect 344066 605858 344302 606094
rect 344386 605858 344622 606094
rect 344066 605538 344302 605774
rect 344386 605538 344622 605774
rect 344066 568658 344302 568894
rect 344386 568658 344622 568894
rect 344066 568338 344302 568574
rect 344386 568338 344622 568574
rect 344066 531458 344302 531694
rect 344386 531458 344622 531694
rect 344066 531138 344302 531374
rect 344386 531138 344622 531374
rect 344066 494258 344302 494494
rect 344386 494258 344622 494494
rect 344066 493938 344302 494174
rect 344386 493938 344622 494174
rect 344066 457058 344302 457294
rect 344386 457058 344622 457294
rect 344066 456738 344302 456974
rect 344386 456738 344622 456974
rect 344066 419858 344302 420094
rect 344386 419858 344622 420094
rect 344066 419538 344302 419774
rect 344386 419538 344622 419774
rect 344066 382658 344302 382894
rect 344386 382658 344622 382894
rect 344066 382338 344302 382574
rect 344386 382338 344622 382574
rect 344066 345458 344302 345694
rect 344386 345458 344622 345694
rect 344066 345138 344302 345374
rect 344386 345138 344622 345374
rect 344066 308258 344302 308494
rect 344386 308258 344622 308494
rect 344066 307938 344302 308174
rect 344386 307938 344622 308174
rect 344066 271058 344302 271294
rect 344386 271058 344622 271294
rect 344066 270738 344302 270974
rect 344386 270738 344622 270974
rect 344066 233858 344302 234094
rect 344386 233858 344622 234094
rect 344066 233538 344302 233774
rect 344386 233538 344622 233774
rect 344066 196658 344302 196894
rect 344386 196658 344622 196894
rect 344066 196338 344302 196574
rect 344386 196338 344622 196574
rect 344066 159458 344302 159694
rect 344386 159458 344622 159694
rect 344066 159138 344302 159374
rect 344386 159138 344622 159374
rect 344066 122258 344302 122494
rect 344386 122258 344622 122494
rect 344066 121938 344302 122174
rect 344386 121938 344622 122174
rect 344066 85058 344302 85294
rect 344386 85058 344622 85294
rect 344066 84738 344302 84974
rect 344386 84738 344622 84974
rect 344066 47858 344302 48094
rect 344386 47858 344622 48094
rect 344066 47538 344302 47774
rect 344386 47538 344622 47774
rect 344066 10658 344302 10894
rect 344386 10658 344622 10894
rect 344066 10338 344302 10574
rect 344386 10338 344622 10574
rect 347786 683978 348022 684214
rect 348106 683978 348342 684214
rect 347786 683658 348022 683894
rect 348106 683658 348342 683894
rect 347786 646778 348022 647014
rect 348106 646778 348342 647014
rect 347786 646458 348022 646694
rect 348106 646458 348342 646694
rect 347786 609578 348022 609814
rect 348106 609578 348342 609814
rect 347786 609258 348022 609494
rect 348106 609258 348342 609494
rect 347786 572378 348022 572614
rect 348106 572378 348342 572614
rect 347786 572058 348022 572294
rect 348106 572058 348342 572294
rect 347786 535178 348022 535414
rect 348106 535178 348342 535414
rect 347786 534858 348022 535094
rect 348106 534858 348342 535094
rect 347786 497978 348022 498214
rect 348106 497978 348342 498214
rect 347786 497658 348022 497894
rect 348106 497658 348342 497894
rect 347786 460778 348022 461014
rect 348106 460778 348342 461014
rect 347786 460458 348022 460694
rect 348106 460458 348342 460694
rect 347786 423578 348022 423814
rect 348106 423578 348342 423814
rect 347786 423258 348022 423494
rect 348106 423258 348342 423494
rect 347786 386378 348022 386614
rect 348106 386378 348342 386614
rect 347786 386058 348022 386294
rect 348106 386058 348342 386294
rect 347786 349178 348022 349414
rect 348106 349178 348342 349414
rect 347786 348858 348022 349094
rect 348106 348858 348342 349094
rect 347786 311978 348022 312214
rect 348106 311978 348342 312214
rect 347786 311658 348022 311894
rect 348106 311658 348342 311894
rect 347786 274778 348022 275014
rect 348106 274778 348342 275014
rect 347786 274458 348022 274694
rect 348106 274458 348342 274694
rect 347786 237578 348022 237814
rect 348106 237578 348342 237814
rect 347786 237258 348022 237494
rect 348106 237258 348342 237494
rect 347786 200378 348022 200614
rect 348106 200378 348342 200614
rect 347786 200058 348022 200294
rect 348106 200058 348342 200294
rect 347786 163178 348022 163414
rect 348106 163178 348342 163414
rect 347786 162858 348022 163094
rect 348106 162858 348342 163094
rect 347786 125978 348022 126214
rect 348106 125978 348342 126214
rect 347786 125658 348022 125894
rect 348106 125658 348342 125894
rect 347786 88778 348022 89014
rect 348106 88778 348342 89014
rect 347786 88458 348022 88694
rect 348106 88458 348342 88694
rect 347786 51578 348022 51814
rect 348106 51578 348342 51814
rect 347786 51258 348022 51494
rect 348106 51258 348342 51494
rect 347786 14378 348022 14614
rect 348106 14378 348342 14614
rect 347786 14058 348022 14294
rect 348106 14058 348342 14294
rect 351506 687698 351742 687934
rect 351826 687698 352062 687934
rect 351506 687378 351742 687614
rect 351826 687378 352062 687614
rect 351506 650498 351742 650734
rect 351826 650498 352062 650734
rect 351506 650178 351742 650414
rect 351826 650178 352062 650414
rect 351506 613298 351742 613534
rect 351826 613298 352062 613534
rect 351506 612978 351742 613214
rect 351826 612978 352062 613214
rect 351506 576098 351742 576334
rect 351826 576098 352062 576334
rect 351506 575778 351742 576014
rect 351826 575778 352062 576014
rect 351506 538898 351742 539134
rect 351826 538898 352062 539134
rect 351506 538578 351742 538814
rect 351826 538578 352062 538814
rect 351506 501698 351742 501934
rect 351826 501698 352062 501934
rect 351506 501378 351742 501614
rect 351826 501378 352062 501614
rect 351506 464498 351742 464734
rect 351826 464498 352062 464734
rect 351506 464178 351742 464414
rect 351826 464178 352062 464414
rect 351506 427298 351742 427534
rect 351826 427298 352062 427534
rect 351506 426978 351742 427214
rect 351826 426978 352062 427214
rect 351506 390098 351742 390334
rect 351826 390098 352062 390334
rect 351506 389778 351742 390014
rect 351826 389778 352062 390014
rect 351506 352898 351742 353134
rect 351826 352898 352062 353134
rect 351506 352578 351742 352814
rect 351826 352578 352062 352814
rect 351506 315698 351742 315934
rect 351826 315698 352062 315934
rect 351506 315378 351742 315614
rect 351826 315378 352062 315614
rect 351506 278498 351742 278734
rect 351826 278498 352062 278734
rect 351506 278178 351742 278414
rect 351826 278178 352062 278414
rect 351506 241298 351742 241534
rect 351826 241298 352062 241534
rect 351506 240978 351742 241214
rect 351826 240978 352062 241214
rect 351506 204098 351742 204334
rect 351826 204098 352062 204334
rect 351506 203778 351742 204014
rect 351826 203778 352062 204014
rect 351506 166898 351742 167134
rect 351826 166898 352062 167134
rect 351506 166578 351742 166814
rect 351826 166578 352062 166814
rect 351506 129698 351742 129934
rect 351826 129698 352062 129934
rect 351506 129378 351742 129614
rect 351826 129378 352062 129614
rect 351506 92498 351742 92734
rect 351826 92498 352062 92734
rect 351506 92178 351742 92414
rect 351826 92178 352062 92414
rect 351506 55298 351742 55534
rect 351826 55298 352062 55534
rect 351506 54978 351742 55214
rect 351826 54978 352062 55214
rect 351506 18098 351742 18334
rect 351826 18098 352062 18334
rect 351506 17778 351742 18014
rect 351826 17778 352062 18014
rect 355226 691418 355462 691654
rect 355546 691418 355782 691654
rect 355226 691098 355462 691334
rect 355546 691098 355782 691334
rect 355226 654218 355462 654454
rect 355546 654218 355782 654454
rect 355226 653898 355462 654134
rect 355546 653898 355782 654134
rect 355226 617018 355462 617254
rect 355546 617018 355782 617254
rect 355226 616698 355462 616934
rect 355546 616698 355782 616934
rect 355226 579818 355462 580054
rect 355546 579818 355782 580054
rect 355226 579498 355462 579734
rect 355546 579498 355782 579734
rect 355226 542618 355462 542854
rect 355546 542618 355782 542854
rect 355226 542298 355462 542534
rect 355546 542298 355782 542534
rect 355226 505418 355462 505654
rect 355546 505418 355782 505654
rect 355226 505098 355462 505334
rect 355546 505098 355782 505334
rect 355226 468218 355462 468454
rect 355546 468218 355782 468454
rect 355226 467898 355462 468134
rect 355546 467898 355782 468134
rect 355226 431018 355462 431254
rect 355546 431018 355782 431254
rect 355226 430698 355462 430934
rect 355546 430698 355782 430934
rect 355226 393818 355462 394054
rect 355546 393818 355782 394054
rect 355226 393498 355462 393734
rect 355546 393498 355782 393734
rect 355226 356618 355462 356854
rect 355546 356618 355782 356854
rect 355226 356298 355462 356534
rect 355546 356298 355782 356534
rect 355226 319418 355462 319654
rect 355546 319418 355782 319654
rect 355226 319098 355462 319334
rect 355546 319098 355782 319334
rect 355226 282218 355462 282454
rect 355546 282218 355782 282454
rect 355226 281898 355462 282134
rect 355546 281898 355782 282134
rect 355226 245018 355462 245254
rect 355546 245018 355782 245254
rect 355226 244698 355462 244934
rect 355546 244698 355782 244934
rect 355226 207818 355462 208054
rect 355546 207818 355782 208054
rect 355226 207498 355462 207734
rect 355546 207498 355782 207734
rect 355226 170618 355462 170854
rect 355546 170618 355782 170854
rect 355226 170298 355462 170534
rect 355546 170298 355782 170534
rect 355226 133418 355462 133654
rect 355546 133418 355782 133654
rect 355226 133098 355462 133334
rect 355546 133098 355782 133334
rect 355226 96218 355462 96454
rect 355546 96218 355782 96454
rect 355226 95898 355462 96134
rect 355546 95898 355782 96134
rect 355226 59018 355462 59254
rect 355546 59018 355782 59254
rect 355226 58698 355462 58934
rect 355546 58698 355782 58934
rect 355226 21818 355462 22054
rect 355546 21818 355782 22054
rect 355226 21498 355462 21734
rect 355546 21498 355782 21734
rect 358946 695138 359182 695374
rect 359266 695138 359502 695374
rect 358946 694818 359182 695054
rect 359266 694818 359502 695054
rect 358946 657938 359182 658174
rect 359266 657938 359502 658174
rect 358946 657618 359182 657854
rect 359266 657618 359502 657854
rect 358946 620738 359182 620974
rect 359266 620738 359502 620974
rect 358946 620418 359182 620654
rect 359266 620418 359502 620654
rect 358946 583538 359182 583774
rect 359266 583538 359502 583774
rect 358946 583218 359182 583454
rect 359266 583218 359502 583454
rect 358946 546338 359182 546574
rect 359266 546338 359502 546574
rect 358946 546018 359182 546254
rect 359266 546018 359502 546254
rect 358946 509138 359182 509374
rect 359266 509138 359502 509374
rect 358946 508818 359182 509054
rect 359266 508818 359502 509054
rect 358946 471938 359182 472174
rect 359266 471938 359502 472174
rect 358946 471618 359182 471854
rect 359266 471618 359502 471854
rect 358946 434738 359182 434974
rect 359266 434738 359502 434974
rect 358946 434418 359182 434654
rect 359266 434418 359502 434654
rect 358946 397538 359182 397774
rect 359266 397538 359502 397774
rect 358946 397218 359182 397454
rect 359266 397218 359502 397454
rect 358946 360338 359182 360574
rect 359266 360338 359502 360574
rect 358946 360018 359182 360254
rect 359266 360018 359502 360254
rect 358946 323138 359182 323374
rect 359266 323138 359502 323374
rect 358946 322818 359182 323054
rect 359266 322818 359502 323054
rect 358946 285938 359182 286174
rect 359266 285938 359502 286174
rect 358946 285618 359182 285854
rect 359266 285618 359502 285854
rect 358946 248738 359182 248974
rect 359266 248738 359502 248974
rect 358946 248418 359182 248654
rect 359266 248418 359502 248654
rect 358946 211538 359182 211774
rect 359266 211538 359502 211774
rect 358946 211218 359182 211454
rect 359266 211218 359502 211454
rect 358946 174338 359182 174574
rect 359266 174338 359502 174574
rect 358946 174018 359182 174254
rect 359266 174018 359502 174254
rect 358946 137138 359182 137374
rect 359266 137138 359502 137374
rect 358946 136818 359182 137054
rect 359266 136818 359502 137054
rect 358946 99938 359182 100174
rect 359266 99938 359502 100174
rect 358946 99618 359182 99854
rect 359266 99618 359502 99854
rect 358946 62738 359182 62974
rect 359266 62738 359502 62974
rect 358946 62418 359182 62654
rect 359266 62418 359502 62654
rect 358946 25538 359182 25774
rect 359266 25538 359502 25774
rect 358946 25218 359182 25454
rect 359266 25218 359502 25454
rect 362666 698858 362902 699094
rect 362986 698858 363222 699094
rect 362666 698538 362902 698774
rect 362986 698538 363222 698774
rect 362666 661658 362902 661894
rect 362986 661658 363222 661894
rect 362666 661338 362902 661574
rect 362986 661338 363222 661574
rect 362666 624458 362902 624694
rect 362986 624458 363222 624694
rect 362666 624138 362902 624374
rect 362986 624138 363222 624374
rect 362666 587258 362902 587494
rect 362986 587258 363222 587494
rect 362666 586938 362902 587174
rect 362986 586938 363222 587174
rect 362666 550058 362902 550294
rect 362986 550058 363222 550294
rect 362666 549738 362902 549974
rect 362986 549738 363222 549974
rect 362666 512858 362902 513094
rect 362986 512858 363222 513094
rect 362666 512538 362902 512774
rect 362986 512538 363222 512774
rect 362666 475658 362902 475894
rect 362986 475658 363222 475894
rect 362666 475338 362902 475574
rect 362986 475338 363222 475574
rect 362666 438458 362902 438694
rect 362986 438458 363222 438694
rect 362666 438138 362902 438374
rect 362986 438138 363222 438374
rect 362666 401258 362902 401494
rect 362986 401258 363222 401494
rect 362666 400938 362902 401174
rect 362986 400938 363222 401174
rect 362666 364058 362902 364294
rect 362986 364058 363222 364294
rect 362666 363738 362902 363974
rect 362986 363738 363222 363974
rect 362666 326858 362902 327094
rect 362986 326858 363222 327094
rect 362666 326538 362902 326774
rect 362986 326538 363222 326774
rect 362666 289658 362902 289894
rect 362986 289658 363222 289894
rect 362666 289338 362902 289574
rect 362986 289338 363222 289574
rect 362666 252458 362902 252694
rect 362986 252458 363222 252694
rect 362666 252138 362902 252374
rect 362986 252138 363222 252374
rect 362666 215258 362902 215494
rect 362986 215258 363222 215494
rect 362666 214938 362902 215174
rect 362986 214938 363222 215174
rect 362666 178058 362902 178294
rect 362986 178058 363222 178294
rect 362666 177738 362902 177974
rect 362986 177738 363222 177974
rect 362666 140858 362902 141094
rect 362986 140858 363222 141094
rect 362666 140538 362902 140774
rect 362986 140538 363222 140774
rect 362666 103658 362902 103894
rect 362986 103658 363222 103894
rect 362666 103338 362902 103574
rect 362986 103338 363222 103574
rect 362666 66458 362902 66694
rect 362986 66458 363222 66694
rect 362666 66138 362902 66374
rect 362986 66138 363222 66374
rect 362666 29258 362902 29494
rect 362986 29258 363222 29494
rect 362666 28938 362902 29174
rect 362986 28938 363222 29174
rect 373826 672818 374062 673054
rect 374146 672818 374382 673054
rect 373826 672498 374062 672734
rect 374146 672498 374382 672734
rect 373826 635618 374062 635854
rect 374146 635618 374382 635854
rect 373826 635298 374062 635534
rect 374146 635298 374382 635534
rect 373826 598418 374062 598654
rect 374146 598418 374382 598654
rect 373826 598098 374062 598334
rect 374146 598098 374382 598334
rect 373826 561218 374062 561454
rect 374146 561218 374382 561454
rect 373826 560898 374062 561134
rect 374146 560898 374382 561134
rect 373826 524018 374062 524254
rect 374146 524018 374382 524254
rect 373826 523698 374062 523934
rect 374146 523698 374382 523934
rect 373826 486818 374062 487054
rect 374146 486818 374382 487054
rect 373826 486498 374062 486734
rect 374146 486498 374382 486734
rect 373826 449618 374062 449854
rect 374146 449618 374382 449854
rect 373826 449298 374062 449534
rect 374146 449298 374382 449534
rect 373826 412418 374062 412654
rect 374146 412418 374382 412654
rect 373826 412098 374062 412334
rect 374146 412098 374382 412334
rect 373826 375218 374062 375454
rect 374146 375218 374382 375454
rect 373826 374898 374062 375134
rect 374146 374898 374382 375134
rect 373826 338018 374062 338254
rect 374146 338018 374382 338254
rect 373826 337698 374062 337934
rect 374146 337698 374382 337934
rect 373826 300818 374062 301054
rect 374146 300818 374382 301054
rect 373826 300498 374062 300734
rect 374146 300498 374382 300734
rect 373826 263618 374062 263854
rect 374146 263618 374382 263854
rect 373826 263298 374062 263534
rect 374146 263298 374382 263534
rect 373826 226418 374062 226654
rect 374146 226418 374382 226654
rect 373826 226098 374062 226334
rect 374146 226098 374382 226334
rect 373826 189218 374062 189454
rect 374146 189218 374382 189454
rect 373826 188898 374062 189134
rect 374146 188898 374382 189134
rect 373826 152018 374062 152254
rect 374146 152018 374382 152254
rect 373826 151698 374062 151934
rect 374146 151698 374382 151934
rect 373826 114818 374062 115054
rect 374146 114818 374382 115054
rect 373826 114498 374062 114734
rect 374146 114498 374382 114734
rect 373826 77618 374062 77854
rect 374146 77618 374382 77854
rect 373826 77298 374062 77534
rect 374146 77298 374382 77534
rect 373826 40418 374062 40654
rect 374146 40418 374382 40654
rect 373826 40098 374062 40334
rect 374146 40098 374382 40334
rect 373826 3218 374062 3454
rect 374146 3218 374382 3454
rect 373826 2898 374062 3134
rect 374146 2898 374382 3134
rect 377546 676538 377782 676774
rect 377866 676538 378102 676774
rect 377546 676218 377782 676454
rect 377866 676218 378102 676454
rect 377546 639338 377782 639574
rect 377866 639338 378102 639574
rect 377546 639018 377782 639254
rect 377866 639018 378102 639254
rect 377546 602138 377782 602374
rect 377866 602138 378102 602374
rect 377546 601818 377782 602054
rect 377866 601818 378102 602054
rect 377546 564938 377782 565174
rect 377866 564938 378102 565174
rect 377546 564618 377782 564854
rect 377866 564618 378102 564854
rect 377546 527738 377782 527974
rect 377866 527738 378102 527974
rect 377546 527418 377782 527654
rect 377866 527418 378102 527654
rect 377546 490538 377782 490774
rect 377866 490538 378102 490774
rect 377546 490218 377782 490454
rect 377866 490218 378102 490454
rect 377546 453338 377782 453574
rect 377866 453338 378102 453574
rect 377546 453018 377782 453254
rect 377866 453018 378102 453254
rect 377546 416138 377782 416374
rect 377866 416138 378102 416374
rect 377546 415818 377782 416054
rect 377866 415818 378102 416054
rect 377546 378938 377782 379174
rect 377866 378938 378102 379174
rect 377546 378618 377782 378854
rect 377866 378618 378102 378854
rect 377546 341738 377782 341974
rect 377866 341738 378102 341974
rect 377546 341418 377782 341654
rect 377866 341418 378102 341654
rect 377546 304538 377782 304774
rect 377866 304538 378102 304774
rect 377546 304218 377782 304454
rect 377866 304218 378102 304454
rect 377546 267338 377782 267574
rect 377866 267338 378102 267574
rect 377546 267018 377782 267254
rect 377866 267018 378102 267254
rect 377546 230138 377782 230374
rect 377866 230138 378102 230374
rect 377546 229818 377782 230054
rect 377866 229818 378102 230054
rect 377546 192938 377782 193174
rect 377866 192938 378102 193174
rect 377546 192618 377782 192854
rect 377866 192618 378102 192854
rect 377546 155738 377782 155974
rect 377866 155738 378102 155974
rect 377546 155418 377782 155654
rect 377866 155418 378102 155654
rect 377546 118538 377782 118774
rect 377866 118538 378102 118774
rect 377546 118218 377782 118454
rect 377866 118218 378102 118454
rect 377546 81338 377782 81574
rect 377866 81338 378102 81574
rect 377546 81018 377782 81254
rect 377866 81018 378102 81254
rect 377546 44138 377782 44374
rect 377866 44138 378102 44374
rect 377546 43818 377782 44054
rect 377866 43818 378102 44054
rect 377546 6938 377782 7174
rect 377866 6938 378102 7174
rect 377546 6618 377782 6854
rect 377866 6618 378102 6854
rect 381266 680258 381502 680494
rect 381586 680258 381822 680494
rect 381266 679938 381502 680174
rect 381586 679938 381822 680174
rect 381266 643058 381502 643294
rect 381586 643058 381822 643294
rect 381266 642738 381502 642974
rect 381586 642738 381822 642974
rect 381266 605858 381502 606094
rect 381586 605858 381822 606094
rect 381266 605538 381502 605774
rect 381586 605538 381822 605774
rect 381266 568658 381502 568894
rect 381586 568658 381822 568894
rect 381266 568338 381502 568574
rect 381586 568338 381822 568574
rect 381266 531458 381502 531694
rect 381586 531458 381822 531694
rect 381266 531138 381502 531374
rect 381586 531138 381822 531374
rect 381266 494258 381502 494494
rect 381586 494258 381822 494494
rect 381266 493938 381502 494174
rect 381586 493938 381822 494174
rect 381266 457058 381502 457294
rect 381586 457058 381822 457294
rect 381266 456738 381502 456974
rect 381586 456738 381822 456974
rect 381266 419858 381502 420094
rect 381586 419858 381822 420094
rect 381266 419538 381502 419774
rect 381586 419538 381822 419774
rect 381266 382658 381502 382894
rect 381586 382658 381822 382894
rect 381266 382338 381502 382574
rect 381586 382338 381822 382574
rect 381266 345458 381502 345694
rect 381586 345458 381822 345694
rect 381266 345138 381502 345374
rect 381586 345138 381822 345374
rect 381266 308258 381502 308494
rect 381586 308258 381822 308494
rect 381266 307938 381502 308174
rect 381586 307938 381822 308174
rect 381266 271058 381502 271294
rect 381586 271058 381822 271294
rect 381266 270738 381502 270974
rect 381586 270738 381822 270974
rect 381266 233858 381502 234094
rect 381586 233858 381822 234094
rect 381266 233538 381502 233774
rect 381586 233538 381822 233774
rect 381266 196658 381502 196894
rect 381586 196658 381822 196894
rect 381266 196338 381502 196574
rect 381586 196338 381822 196574
rect 381266 159458 381502 159694
rect 381586 159458 381822 159694
rect 381266 159138 381502 159374
rect 381586 159138 381822 159374
rect 381266 122258 381502 122494
rect 381586 122258 381822 122494
rect 381266 121938 381502 122174
rect 381586 121938 381822 122174
rect 381266 85058 381502 85294
rect 381586 85058 381822 85294
rect 381266 84738 381502 84974
rect 381586 84738 381822 84974
rect 381266 47858 381502 48094
rect 381586 47858 381822 48094
rect 381266 47538 381502 47774
rect 381586 47538 381822 47774
rect 381266 10658 381502 10894
rect 381586 10658 381822 10894
rect 381266 10338 381502 10574
rect 381586 10338 381822 10574
rect 384986 683978 385222 684214
rect 385306 683978 385542 684214
rect 384986 683658 385222 683894
rect 385306 683658 385542 683894
rect 384986 646778 385222 647014
rect 385306 646778 385542 647014
rect 384986 646458 385222 646694
rect 385306 646458 385542 646694
rect 384986 609578 385222 609814
rect 385306 609578 385542 609814
rect 384986 609258 385222 609494
rect 385306 609258 385542 609494
rect 384986 572378 385222 572614
rect 385306 572378 385542 572614
rect 384986 572058 385222 572294
rect 385306 572058 385542 572294
rect 384986 535178 385222 535414
rect 385306 535178 385542 535414
rect 384986 534858 385222 535094
rect 385306 534858 385542 535094
rect 384986 497978 385222 498214
rect 385306 497978 385542 498214
rect 384986 497658 385222 497894
rect 385306 497658 385542 497894
rect 384986 460778 385222 461014
rect 385306 460778 385542 461014
rect 384986 460458 385222 460694
rect 385306 460458 385542 460694
rect 384986 423578 385222 423814
rect 385306 423578 385542 423814
rect 384986 423258 385222 423494
rect 385306 423258 385542 423494
rect 384986 386378 385222 386614
rect 385306 386378 385542 386614
rect 384986 386058 385222 386294
rect 385306 386058 385542 386294
rect 384986 349178 385222 349414
rect 385306 349178 385542 349414
rect 384986 348858 385222 349094
rect 385306 348858 385542 349094
rect 384986 311978 385222 312214
rect 385306 311978 385542 312214
rect 384986 311658 385222 311894
rect 385306 311658 385542 311894
rect 384986 274778 385222 275014
rect 385306 274778 385542 275014
rect 384986 274458 385222 274694
rect 385306 274458 385542 274694
rect 384986 237578 385222 237814
rect 385306 237578 385542 237814
rect 384986 237258 385222 237494
rect 385306 237258 385542 237494
rect 384986 200378 385222 200614
rect 385306 200378 385542 200614
rect 384986 200058 385222 200294
rect 385306 200058 385542 200294
rect 384986 163178 385222 163414
rect 385306 163178 385542 163414
rect 384986 162858 385222 163094
rect 385306 162858 385542 163094
rect 384986 125978 385222 126214
rect 385306 125978 385542 126214
rect 384986 125658 385222 125894
rect 385306 125658 385542 125894
rect 384986 88778 385222 89014
rect 385306 88778 385542 89014
rect 384986 88458 385222 88694
rect 385306 88458 385542 88694
rect 384986 51578 385222 51814
rect 385306 51578 385542 51814
rect 384986 51258 385222 51494
rect 385306 51258 385542 51494
rect 384986 14378 385222 14614
rect 385306 14378 385542 14614
rect 384986 14058 385222 14294
rect 385306 14058 385542 14294
rect 388706 687698 388942 687934
rect 389026 687698 389262 687934
rect 388706 687378 388942 687614
rect 389026 687378 389262 687614
rect 388706 650498 388942 650734
rect 389026 650498 389262 650734
rect 388706 650178 388942 650414
rect 389026 650178 389262 650414
rect 388706 613298 388942 613534
rect 389026 613298 389262 613534
rect 388706 612978 388942 613214
rect 389026 612978 389262 613214
rect 388706 576098 388942 576334
rect 389026 576098 389262 576334
rect 388706 575778 388942 576014
rect 389026 575778 389262 576014
rect 388706 538898 388942 539134
rect 389026 538898 389262 539134
rect 388706 538578 388942 538814
rect 389026 538578 389262 538814
rect 388706 501698 388942 501934
rect 389026 501698 389262 501934
rect 388706 501378 388942 501614
rect 389026 501378 389262 501614
rect 388706 464498 388942 464734
rect 389026 464498 389262 464734
rect 388706 464178 388942 464414
rect 389026 464178 389262 464414
rect 388706 427298 388942 427534
rect 389026 427298 389262 427534
rect 388706 426978 388942 427214
rect 389026 426978 389262 427214
rect 388706 390098 388942 390334
rect 389026 390098 389262 390334
rect 388706 389778 388942 390014
rect 389026 389778 389262 390014
rect 388706 352898 388942 353134
rect 389026 352898 389262 353134
rect 388706 352578 388942 352814
rect 389026 352578 389262 352814
rect 388706 315698 388942 315934
rect 389026 315698 389262 315934
rect 388706 315378 388942 315614
rect 389026 315378 389262 315614
rect 388706 278498 388942 278734
rect 389026 278498 389262 278734
rect 388706 278178 388942 278414
rect 389026 278178 389262 278414
rect 388706 241298 388942 241534
rect 389026 241298 389262 241534
rect 388706 240978 388942 241214
rect 389026 240978 389262 241214
rect 388706 204098 388942 204334
rect 389026 204098 389262 204334
rect 388706 203778 388942 204014
rect 389026 203778 389262 204014
rect 388706 166898 388942 167134
rect 389026 166898 389262 167134
rect 388706 166578 388942 166814
rect 389026 166578 389262 166814
rect 388706 129698 388942 129934
rect 389026 129698 389262 129934
rect 388706 129378 388942 129614
rect 389026 129378 389262 129614
rect 388706 92498 388942 92734
rect 389026 92498 389262 92734
rect 388706 92178 388942 92414
rect 389026 92178 389262 92414
rect 388706 55298 388942 55534
rect 389026 55298 389262 55534
rect 388706 54978 388942 55214
rect 389026 54978 389262 55214
rect 388706 18098 388942 18334
rect 389026 18098 389262 18334
rect 388706 17778 388942 18014
rect 389026 17778 389262 18014
rect 392426 691418 392662 691654
rect 392746 691418 392982 691654
rect 392426 691098 392662 691334
rect 392746 691098 392982 691334
rect 392426 654218 392662 654454
rect 392746 654218 392982 654454
rect 392426 653898 392662 654134
rect 392746 653898 392982 654134
rect 392426 617018 392662 617254
rect 392746 617018 392982 617254
rect 392426 616698 392662 616934
rect 392746 616698 392982 616934
rect 392426 579818 392662 580054
rect 392746 579818 392982 580054
rect 392426 579498 392662 579734
rect 392746 579498 392982 579734
rect 392426 542618 392662 542854
rect 392746 542618 392982 542854
rect 392426 542298 392662 542534
rect 392746 542298 392982 542534
rect 392426 505418 392662 505654
rect 392746 505418 392982 505654
rect 392426 505098 392662 505334
rect 392746 505098 392982 505334
rect 392426 468218 392662 468454
rect 392746 468218 392982 468454
rect 392426 467898 392662 468134
rect 392746 467898 392982 468134
rect 392426 431018 392662 431254
rect 392746 431018 392982 431254
rect 392426 430698 392662 430934
rect 392746 430698 392982 430934
rect 392426 393818 392662 394054
rect 392746 393818 392982 394054
rect 392426 393498 392662 393734
rect 392746 393498 392982 393734
rect 392426 356618 392662 356854
rect 392746 356618 392982 356854
rect 392426 356298 392662 356534
rect 392746 356298 392982 356534
rect 392426 319418 392662 319654
rect 392746 319418 392982 319654
rect 392426 319098 392662 319334
rect 392746 319098 392982 319334
rect 392426 282218 392662 282454
rect 392746 282218 392982 282454
rect 392426 281898 392662 282134
rect 392746 281898 392982 282134
rect 392426 245018 392662 245254
rect 392746 245018 392982 245254
rect 392426 244698 392662 244934
rect 392746 244698 392982 244934
rect 392426 207818 392662 208054
rect 392746 207818 392982 208054
rect 392426 207498 392662 207734
rect 392746 207498 392982 207734
rect 392426 170618 392662 170854
rect 392746 170618 392982 170854
rect 392426 170298 392662 170534
rect 392746 170298 392982 170534
rect 392426 133418 392662 133654
rect 392746 133418 392982 133654
rect 392426 133098 392662 133334
rect 392746 133098 392982 133334
rect 392426 96218 392662 96454
rect 392746 96218 392982 96454
rect 392426 95898 392662 96134
rect 392746 95898 392982 96134
rect 392426 59018 392662 59254
rect 392746 59018 392982 59254
rect 392426 58698 392662 58934
rect 392746 58698 392982 58934
rect 392426 21818 392662 22054
rect 392746 21818 392982 22054
rect 392426 21498 392662 21734
rect 392746 21498 392982 21734
rect 396146 695138 396382 695374
rect 396466 695138 396702 695374
rect 396146 694818 396382 695054
rect 396466 694818 396702 695054
rect 396146 657938 396382 658174
rect 396466 657938 396702 658174
rect 396146 657618 396382 657854
rect 396466 657618 396702 657854
rect 396146 620738 396382 620974
rect 396466 620738 396702 620974
rect 396146 620418 396382 620654
rect 396466 620418 396702 620654
rect 396146 583538 396382 583774
rect 396466 583538 396702 583774
rect 396146 583218 396382 583454
rect 396466 583218 396702 583454
rect 396146 546338 396382 546574
rect 396466 546338 396702 546574
rect 396146 546018 396382 546254
rect 396466 546018 396702 546254
rect 396146 509138 396382 509374
rect 396466 509138 396702 509374
rect 396146 508818 396382 509054
rect 396466 508818 396702 509054
rect 396146 471938 396382 472174
rect 396466 471938 396702 472174
rect 396146 471618 396382 471854
rect 396466 471618 396702 471854
rect 396146 434738 396382 434974
rect 396466 434738 396702 434974
rect 396146 434418 396382 434654
rect 396466 434418 396702 434654
rect 396146 397538 396382 397774
rect 396466 397538 396702 397774
rect 396146 397218 396382 397454
rect 396466 397218 396702 397454
rect 396146 360338 396382 360574
rect 396466 360338 396702 360574
rect 396146 360018 396382 360254
rect 396466 360018 396702 360254
rect 396146 323138 396382 323374
rect 396466 323138 396702 323374
rect 396146 322818 396382 323054
rect 396466 322818 396702 323054
rect 396146 285938 396382 286174
rect 396466 285938 396702 286174
rect 396146 285618 396382 285854
rect 396466 285618 396702 285854
rect 396146 248738 396382 248974
rect 396466 248738 396702 248974
rect 396146 248418 396382 248654
rect 396466 248418 396702 248654
rect 396146 211538 396382 211774
rect 396466 211538 396702 211774
rect 396146 211218 396382 211454
rect 396466 211218 396702 211454
rect 396146 174338 396382 174574
rect 396466 174338 396702 174574
rect 396146 174018 396382 174254
rect 396466 174018 396702 174254
rect 396146 137138 396382 137374
rect 396466 137138 396702 137374
rect 396146 136818 396382 137054
rect 396466 136818 396702 137054
rect 396146 99938 396382 100174
rect 396466 99938 396702 100174
rect 396146 99618 396382 99854
rect 396466 99618 396702 99854
rect 396146 62738 396382 62974
rect 396466 62738 396702 62974
rect 396146 62418 396382 62654
rect 396466 62418 396702 62654
rect 396146 25538 396382 25774
rect 396466 25538 396702 25774
rect 396146 25218 396382 25454
rect 396466 25218 396702 25454
rect 399866 698858 400102 699094
rect 400186 698858 400422 699094
rect 399866 698538 400102 698774
rect 400186 698538 400422 698774
rect 399866 661658 400102 661894
rect 400186 661658 400422 661894
rect 399866 661338 400102 661574
rect 400186 661338 400422 661574
rect 399866 624458 400102 624694
rect 400186 624458 400422 624694
rect 399866 624138 400102 624374
rect 400186 624138 400422 624374
rect 399866 587258 400102 587494
rect 400186 587258 400422 587494
rect 399866 586938 400102 587174
rect 400186 586938 400422 587174
rect 399866 550058 400102 550294
rect 400186 550058 400422 550294
rect 399866 549738 400102 549974
rect 400186 549738 400422 549974
rect 399866 512858 400102 513094
rect 400186 512858 400422 513094
rect 399866 512538 400102 512774
rect 400186 512538 400422 512774
rect 399866 475658 400102 475894
rect 400186 475658 400422 475894
rect 399866 475338 400102 475574
rect 400186 475338 400422 475574
rect 399866 438458 400102 438694
rect 400186 438458 400422 438694
rect 399866 438138 400102 438374
rect 400186 438138 400422 438374
rect 399866 401258 400102 401494
rect 400186 401258 400422 401494
rect 399866 400938 400102 401174
rect 400186 400938 400422 401174
rect 399866 364058 400102 364294
rect 400186 364058 400422 364294
rect 399866 363738 400102 363974
rect 400186 363738 400422 363974
rect 399866 326858 400102 327094
rect 400186 326858 400422 327094
rect 399866 326538 400102 326774
rect 400186 326538 400422 326774
rect 399866 289658 400102 289894
rect 400186 289658 400422 289894
rect 399866 289338 400102 289574
rect 400186 289338 400422 289574
rect 399866 252458 400102 252694
rect 400186 252458 400422 252694
rect 399866 252138 400102 252374
rect 400186 252138 400422 252374
rect 399866 215258 400102 215494
rect 400186 215258 400422 215494
rect 399866 214938 400102 215174
rect 400186 214938 400422 215174
rect 399866 178058 400102 178294
rect 400186 178058 400422 178294
rect 399866 177738 400102 177974
rect 400186 177738 400422 177974
rect 399866 140858 400102 141094
rect 400186 140858 400422 141094
rect 399866 140538 400102 140774
rect 400186 140538 400422 140774
rect 399866 103658 400102 103894
rect 400186 103658 400422 103894
rect 399866 103338 400102 103574
rect 400186 103338 400422 103574
rect 399866 66458 400102 66694
rect 400186 66458 400422 66694
rect 399866 66138 400102 66374
rect 400186 66138 400422 66374
rect 399866 29258 400102 29494
rect 400186 29258 400422 29494
rect 399866 28938 400102 29174
rect 400186 28938 400422 29174
rect 411026 672818 411262 673054
rect 411346 672818 411582 673054
rect 411026 672498 411262 672734
rect 411346 672498 411582 672734
rect 411026 635618 411262 635854
rect 411346 635618 411582 635854
rect 411026 635298 411262 635534
rect 411346 635298 411582 635534
rect 411026 598418 411262 598654
rect 411346 598418 411582 598654
rect 411026 598098 411262 598334
rect 411346 598098 411582 598334
rect 411026 561218 411262 561454
rect 411346 561218 411582 561454
rect 411026 560898 411262 561134
rect 411346 560898 411582 561134
rect 411026 524018 411262 524254
rect 411346 524018 411582 524254
rect 411026 523698 411262 523934
rect 411346 523698 411582 523934
rect 411026 486818 411262 487054
rect 411346 486818 411582 487054
rect 411026 486498 411262 486734
rect 411346 486498 411582 486734
rect 411026 449618 411262 449854
rect 411346 449618 411582 449854
rect 411026 449298 411262 449534
rect 411346 449298 411582 449534
rect 411026 412418 411262 412654
rect 411346 412418 411582 412654
rect 411026 412098 411262 412334
rect 411346 412098 411582 412334
rect 411026 375218 411262 375454
rect 411346 375218 411582 375454
rect 411026 374898 411262 375134
rect 411346 374898 411582 375134
rect 411026 338018 411262 338254
rect 411346 338018 411582 338254
rect 411026 337698 411262 337934
rect 411346 337698 411582 337934
rect 411026 300818 411262 301054
rect 411346 300818 411582 301054
rect 411026 300498 411262 300734
rect 411346 300498 411582 300734
rect 411026 263618 411262 263854
rect 411346 263618 411582 263854
rect 411026 263298 411262 263534
rect 411346 263298 411582 263534
rect 411026 226418 411262 226654
rect 411346 226418 411582 226654
rect 411026 226098 411262 226334
rect 411346 226098 411582 226334
rect 411026 189218 411262 189454
rect 411346 189218 411582 189454
rect 411026 188898 411262 189134
rect 411346 188898 411582 189134
rect 411026 152018 411262 152254
rect 411346 152018 411582 152254
rect 411026 151698 411262 151934
rect 411346 151698 411582 151934
rect 411026 114818 411262 115054
rect 411346 114818 411582 115054
rect 411026 114498 411262 114734
rect 411346 114498 411582 114734
rect 411026 77618 411262 77854
rect 411346 77618 411582 77854
rect 411026 77298 411262 77534
rect 411346 77298 411582 77534
rect 411026 40418 411262 40654
rect 411346 40418 411582 40654
rect 411026 40098 411262 40334
rect 411346 40098 411582 40334
rect 411026 3218 411262 3454
rect 411346 3218 411582 3454
rect 411026 2898 411262 3134
rect 411346 2898 411582 3134
rect 414746 676538 414982 676774
rect 415066 676538 415302 676774
rect 414746 676218 414982 676454
rect 415066 676218 415302 676454
rect 414746 639338 414982 639574
rect 415066 639338 415302 639574
rect 414746 639018 414982 639254
rect 415066 639018 415302 639254
rect 414746 602138 414982 602374
rect 415066 602138 415302 602374
rect 414746 601818 414982 602054
rect 415066 601818 415302 602054
rect 414746 564938 414982 565174
rect 415066 564938 415302 565174
rect 414746 564618 414982 564854
rect 415066 564618 415302 564854
rect 414746 527738 414982 527974
rect 415066 527738 415302 527974
rect 414746 527418 414982 527654
rect 415066 527418 415302 527654
rect 414746 490538 414982 490774
rect 415066 490538 415302 490774
rect 414746 490218 414982 490454
rect 415066 490218 415302 490454
rect 414746 453338 414982 453574
rect 415066 453338 415302 453574
rect 414746 453018 414982 453254
rect 415066 453018 415302 453254
rect 414746 416138 414982 416374
rect 415066 416138 415302 416374
rect 414746 415818 414982 416054
rect 415066 415818 415302 416054
rect 414746 378938 414982 379174
rect 415066 378938 415302 379174
rect 414746 378618 414982 378854
rect 415066 378618 415302 378854
rect 414746 341738 414982 341974
rect 415066 341738 415302 341974
rect 414746 341418 414982 341654
rect 415066 341418 415302 341654
rect 414746 304538 414982 304774
rect 415066 304538 415302 304774
rect 414746 304218 414982 304454
rect 415066 304218 415302 304454
rect 414746 267338 414982 267574
rect 415066 267338 415302 267574
rect 414746 267018 414982 267254
rect 415066 267018 415302 267254
rect 414746 230138 414982 230374
rect 415066 230138 415302 230374
rect 414746 229818 414982 230054
rect 415066 229818 415302 230054
rect 414746 192938 414982 193174
rect 415066 192938 415302 193174
rect 414746 192618 414982 192854
rect 415066 192618 415302 192854
rect 414746 155738 414982 155974
rect 415066 155738 415302 155974
rect 414746 155418 414982 155654
rect 415066 155418 415302 155654
rect 414746 118538 414982 118774
rect 415066 118538 415302 118774
rect 414746 118218 414982 118454
rect 415066 118218 415302 118454
rect 414746 81338 414982 81574
rect 415066 81338 415302 81574
rect 414746 81018 414982 81254
rect 415066 81018 415302 81254
rect 414746 44138 414982 44374
rect 415066 44138 415302 44374
rect 414746 43818 414982 44054
rect 415066 43818 415302 44054
rect 414746 6938 414982 7174
rect 415066 6938 415302 7174
rect 414746 6618 414982 6854
rect 415066 6618 415302 6854
rect 418466 680258 418702 680494
rect 418786 680258 419022 680494
rect 418466 679938 418702 680174
rect 418786 679938 419022 680174
rect 418466 643058 418702 643294
rect 418786 643058 419022 643294
rect 418466 642738 418702 642974
rect 418786 642738 419022 642974
rect 418466 605858 418702 606094
rect 418786 605858 419022 606094
rect 418466 605538 418702 605774
rect 418786 605538 419022 605774
rect 418466 568658 418702 568894
rect 418786 568658 419022 568894
rect 418466 568338 418702 568574
rect 418786 568338 419022 568574
rect 418466 531458 418702 531694
rect 418786 531458 419022 531694
rect 418466 531138 418702 531374
rect 418786 531138 419022 531374
rect 418466 494258 418702 494494
rect 418786 494258 419022 494494
rect 418466 493938 418702 494174
rect 418786 493938 419022 494174
rect 418466 457058 418702 457294
rect 418786 457058 419022 457294
rect 418466 456738 418702 456974
rect 418786 456738 419022 456974
rect 418466 419858 418702 420094
rect 418786 419858 419022 420094
rect 418466 419538 418702 419774
rect 418786 419538 419022 419774
rect 418466 382658 418702 382894
rect 418786 382658 419022 382894
rect 418466 382338 418702 382574
rect 418786 382338 419022 382574
rect 418466 345458 418702 345694
rect 418786 345458 419022 345694
rect 418466 345138 418702 345374
rect 418786 345138 419022 345374
rect 418466 308258 418702 308494
rect 418786 308258 419022 308494
rect 418466 307938 418702 308174
rect 418786 307938 419022 308174
rect 418466 271058 418702 271294
rect 418786 271058 419022 271294
rect 418466 270738 418702 270974
rect 418786 270738 419022 270974
rect 418466 233858 418702 234094
rect 418786 233858 419022 234094
rect 418466 233538 418702 233774
rect 418786 233538 419022 233774
rect 418466 196658 418702 196894
rect 418786 196658 419022 196894
rect 418466 196338 418702 196574
rect 418786 196338 419022 196574
rect 418466 159458 418702 159694
rect 418786 159458 419022 159694
rect 418466 159138 418702 159374
rect 418786 159138 419022 159374
rect 418466 122258 418702 122494
rect 418786 122258 419022 122494
rect 418466 121938 418702 122174
rect 418786 121938 419022 122174
rect 418466 85058 418702 85294
rect 418786 85058 419022 85294
rect 418466 84738 418702 84974
rect 418786 84738 419022 84974
rect 418466 47858 418702 48094
rect 418786 47858 419022 48094
rect 418466 47538 418702 47774
rect 418786 47538 419022 47774
rect 418466 10658 418702 10894
rect 418786 10658 419022 10894
rect 418466 10338 418702 10574
rect 418786 10338 419022 10574
rect 422186 683978 422422 684214
rect 422506 683978 422742 684214
rect 422186 683658 422422 683894
rect 422506 683658 422742 683894
rect 422186 646778 422422 647014
rect 422506 646778 422742 647014
rect 422186 646458 422422 646694
rect 422506 646458 422742 646694
rect 422186 609578 422422 609814
rect 422506 609578 422742 609814
rect 422186 609258 422422 609494
rect 422506 609258 422742 609494
rect 422186 572378 422422 572614
rect 422506 572378 422742 572614
rect 422186 572058 422422 572294
rect 422506 572058 422742 572294
rect 422186 535178 422422 535414
rect 422506 535178 422742 535414
rect 422186 534858 422422 535094
rect 422506 534858 422742 535094
rect 422186 497978 422422 498214
rect 422506 497978 422742 498214
rect 422186 497658 422422 497894
rect 422506 497658 422742 497894
rect 422186 460778 422422 461014
rect 422506 460778 422742 461014
rect 422186 460458 422422 460694
rect 422506 460458 422742 460694
rect 422186 423578 422422 423814
rect 422506 423578 422742 423814
rect 422186 423258 422422 423494
rect 422506 423258 422742 423494
rect 422186 386378 422422 386614
rect 422506 386378 422742 386614
rect 422186 386058 422422 386294
rect 422506 386058 422742 386294
rect 422186 349178 422422 349414
rect 422506 349178 422742 349414
rect 422186 348858 422422 349094
rect 422506 348858 422742 349094
rect 422186 311978 422422 312214
rect 422506 311978 422742 312214
rect 422186 311658 422422 311894
rect 422506 311658 422742 311894
rect 422186 274778 422422 275014
rect 422506 274778 422742 275014
rect 422186 274458 422422 274694
rect 422506 274458 422742 274694
rect 422186 237578 422422 237814
rect 422506 237578 422742 237814
rect 422186 237258 422422 237494
rect 422506 237258 422742 237494
rect 422186 200378 422422 200614
rect 422506 200378 422742 200614
rect 422186 200058 422422 200294
rect 422506 200058 422742 200294
rect 422186 163178 422422 163414
rect 422506 163178 422742 163414
rect 422186 162858 422422 163094
rect 422506 162858 422742 163094
rect 422186 125978 422422 126214
rect 422506 125978 422742 126214
rect 422186 125658 422422 125894
rect 422506 125658 422742 125894
rect 422186 88778 422422 89014
rect 422506 88778 422742 89014
rect 422186 88458 422422 88694
rect 422506 88458 422742 88694
rect 422186 51578 422422 51814
rect 422506 51578 422742 51814
rect 422186 51258 422422 51494
rect 422506 51258 422742 51494
rect 422186 14378 422422 14614
rect 422506 14378 422742 14614
rect 422186 14058 422422 14294
rect 422506 14058 422742 14294
rect 425906 687698 426142 687934
rect 426226 687698 426462 687934
rect 425906 687378 426142 687614
rect 426226 687378 426462 687614
rect 425906 650498 426142 650734
rect 426226 650498 426462 650734
rect 425906 650178 426142 650414
rect 426226 650178 426462 650414
rect 425906 613298 426142 613534
rect 426226 613298 426462 613534
rect 425906 612978 426142 613214
rect 426226 612978 426462 613214
rect 425906 576098 426142 576334
rect 426226 576098 426462 576334
rect 425906 575778 426142 576014
rect 426226 575778 426462 576014
rect 425906 538898 426142 539134
rect 426226 538898 426462 539134
rect 425906 538578 426142 538814
rect 426226 538578 426462 538814
rect 425906 501698 426142 501934
rect 426226 501698 426462 501934
rect 425906 501378 426142 501614
rect 426226 501378 426462 501614
rect 425906 464498 426142 464734
rect 426226 464498 426462 464734
rect 425906 464178 426142 464414
rect 426226 464178 426462 464414
rect 425906 427298 426142 427534
rect 426226 427298 426462 427534
rect 425906 426978 426142 427214
rect 426226 426978 426462 427214
rect 425906 390098 426142 390334
rect 426226 390098 426462 390334
rect 425906 389778 426142 390014
rect 426226 389778 426462 390014
rect 425906 352898 426142 353134
rect 426226 352898 426462 353134
rect 425906 352578 426142 352814
rect 426226 352578 426462 352814
rect 425906 315698 426142 315934
rect 426226 315698 426462 315934
rect 425906 315378 426142 315614
rect 426226 315378 426462 315614
rect 425906 278498 426142 278734
rect 426226 278498 426462 278734
rect 425906 278178 426142 278414
rect 426226 278178 426462 278414
rect 425906 241298 426142 241534
rect 426226 241298 426462 241534
rect 425906 240978 426142 241214
rect 426226 240978 426462 241214
rect 425906 204098 426142 204334
rect 426226 204098 426462 204334
rect 425906 203778 426142 204014
rect 426226 203778 426462 204014
rect 425906 166898 426142 167134
rect 426226 166898 426462 167134
rect 425906 166578 426142 166814
rect 426226 166578 426462 166814
rect 425906 129698 426142 129934
rect 426226 129698 426462 129934
rect 425906 129378 426142 129614
rect 426226 129378 426462 129614
rect 425906 92498 426142 92734
rect 426226 92498 426462 92734
rect 425906 92178 426142 92414
rect 426226 92178 426462 92414
rect 425906 55298 426142 55534
rect 426226 55298 426462 55534
rect 425906 54978 426142 55214
rect 426226 54978 426462 55214
rect 425906 18098 426142 18334
rect 426226 18098 426462 18334
rect 425906 17778 426142 18014
rect 426226 17778 426462 18014
rect 429626 691418 429862 691654
rect 429946 691418 430182 691654
rect 429626 691098 429862 691334
rect 429946 691098 430182 691334
rect 429626 654218 429862 654454
rect 429946 654218 430182 654454
rect 429626 653898 429862 654134
rect 429946 653898 430182 654134
rect 429626 617018 429862 617254
rect 429946 617018 430182 617254
rect 429626 616698 429862 616934
rect 429946 616698 430182 616934
rect 429626 579818 429862 580054
rect 429946 579818 430182 580054
rect 429626 579498 429862 579734
rect 429946 579498 430182 579734
rect 429626 542618 429862 542854
rect 429946 542618 430182 542854
rect 429626 542298 429862 542534
rect 429946 542298 430182 542534
rect 429626 505418 429862 505654
rect 429946 505418 430182 505654
rect 429626 505098 429862 505334
rect 429946 505098 430182 505334
rect 429626 468218 429862 468454
rect 429946 468218 430182 468454
rect 429626 467898 429862 468134
rect 429946 467898 430182 468134
rect 429626 431018 429862 431254
rect 429946 431018 430182 431254
rect 429626 430698 429862 430934
rect 429946 430698 430182 430934
rect 429626 393818 429862 394054
rect 429946 393818 430182 394054
rect 429626 393498 429862 393734
rect 429946 393498 430182 393734
rect 429626 356618 429862 356854
rect 429946 356618 430182 356854
rect 429626 356298 429862 356534
rect 429946 356298 430182 356534
rect 429626 319418 429862 319654
rect 429946 319418 430182 319654
rect 429626 319098 429862 319334
rect 429946 319098 430182 319334
rect 429626 282218 429862 282454
rect 429946 282218 430182 282454
rect 429626 281898 429862 282134
rect 429946 281898 430182 282134
rect 429626 245018 429862 245254
rect 429946 245018 430182 245254
rect 429626 244698 429862 244934
rect 429946 244698 430182 244934
rect 429626 207818 429862 208054
rect 429946 207818 430182 208054
rect 429626 207498 429862 207734
rect 429946 207498 430182 207734
rect 429626 170618 429862 170854
rect 429946 170618 430182 170854
rect 429626 170298 429862 170534
rect 429946 170298 430182 170534
rect 429626 133418 429862 133654
rect 429946 133418 430182 133654
rect 429626 133098 429862 133334
rect 429946 133098 430182 133334
rect 429626 96218 429862 96454
rect 429946 96218 430182 96454
rect 429626 95898 429862 96134
rect 429946 95898 430182 96134
rect 429626 59018 429862 59254
rect 429946 59018 430182 59254
rect 429626 58698 429862 58934
rect 429946 58698 430182 58934
rect 429626 21818 429862 22054
rect 429946 21818 430182 22054
rect 429626 21498 429862 21734
rect 429946 21498 430182 21734
rect 433346 695138 433582 695374
rect 433666 695138 433902 695374
rect 433346 694818 433582 695054
rect 433666 694818 433902 695054
rect 433346 657938 433582 658174
rect 433666 657938 433902 658174
rect 433346 657618 433582 657854
rect 433666 657618 433902 657854
rect 433346 620738 433582 620974
rect 433666 620738 433902 620974
rect 433346 620418 433582 620654
rect 433666 620418 433902 620654
rect 433346 583538 433582 583774
rect 433666 583538 433902 583774
rect 433346 583218 433582 583454
rect 433666 583218 433902 583454
rect 433346 546338 433582 546574
rect 433666 546338 433902 546574
rect 433346 546018 433582 546254
rect 433666 546018 433902 546254
rect 433346 509138 433582 509374
rect 433666 509138 433902 509374
rect 433346 508818 433582 509054
rect 433666 508818 433902 509054
rect 433346 471938 433582 472174
rect 433666 471938 433902 472174
rect 433346 471618 433582 471854
rect 433666 471618 433902 471854
rect 433346 434738 433582 434974
rect 433666 434738 433902 434974
rect 433346 434418 433582 434654
rect 433666 434418 433902 434654
rect 433346 397538 433582 397774
rect 433666 397538 433902 397774
rect 433346 397218 433582 397454
rect 433666 397218 433902 397454
rect 433346 360338 433582 360574
rect 433666 360338 433902 360574
rect 433346 360018 433582 360254
rect 433666 360018 433902 360254
rect 433346 323138 433582 323374
rect 433666 323138 433902 323374
rect 433346 322818 433582 323054
rect 433666 322818 433902 323054
rect 433346 285938 433582 286174
rect 433666 285938 433902 286174
rect 433346 285618 433582 285854
rect 433666 285618 433902 285854
rect 433346 248738 433582 248974
rect 433666 248738 433902 248974
rect 433346 248418 433582 248654
rect 433666 248418 433902 248654
rect 433346 211538 433582 211774
rect 433666 211538 433902 211774
rect 433346 211218 433582 211454
rect 433666 211218 433902 211454
rect 433346 174338 433582 174574
rect 433666 174338 433902 174574
rect 433346 174018 433582 174254
rect 433666 174018 433902 174254
rect 433346 137138 433582 137374
rect 433666 137138 433902 137374
rect 433346 136818 433582 137054
rect 433666 136818 433902 137054
rect 433346 99938 433582 100174
rect 433666 99938 433902 100174
rect 433346 99618 433582 99854
rect 433666 99618 433902 99854
rect 433346 62738 433582 62974
rect 433666 62738 433902 62974
rect 433346 62418 433582 62654
rect 433666 62418 433902 62654
rect 433346 25538 433582 25774
rect 433666 25538 433902 25774
rect 433346 25218 433582 25454
rect 433666 25218 433902 25454
rect 437066 698858 437302 699094
rect 437386 698858 437622 699094
rect 437066 698538 437302 698774
rect 437386 698538 437622 698774
rect 437066 661658 437302 661894
rect 437386 661658 437622 661894
rect 437066 661338 437302 661574
rect 437386 661338 437622 661574
rect 437066 624458 437302 624694
rect 437386 624458 437622 624694
rect 437066 624138 437302 624374
rect 437386 624138 437622 624374
rect 437066 587258 437302 587494
rect 437386 587258 437622 587494
rect 437066 586938 437302 587174
rect 437386 586938 437622 587174
rect 437066 550058 437302 550294
rect 437386 550058 437622 550294
rect 437066 549738 437302 549974
rect 437386 549738 437622 549974
rect 437066 512858 437302 513094
rect 437386 512858 437622 513094
rect 437066 512538 437302 512774
rect 437386 512538 437622 512774
rect 437066 475658 437302 475894
rect 437386 475658 437622 475894
rect 437066 475338 437302 475574
rect 437386 475338 437622 475574
rect 437066 438458 437302 438694
rect 437386 438458 437622 438694
rect 437066 438138 437302 438374
rect 437386 438138 437622 438374
rect 437066 401258 437302 401494
rect 437386 401258 437622 401494
rect 437066 400938 437302 401174
rect 437386 400938 437622 401174
rect 437066 364058 437302 364294
rect 437386 364058 437622 364294
rect 437066 363738 437302 363974
rect 437386 363738 437622 363974
rect 437066 326858 437302 327094
rect 437386 326858 437622 327094
rect 437066 326538 437302 326774
rect 437386 326538 437622 326774
rect 437066 289658 437302 289894
rect 437386 289658 437622 289894
rect 437066 289338 437302 289574
rect 437386 289338 437622 289574
rect 437066 252458 437302 252694
rect 437386 252458 437622 252694
rect 437066 252138 437302 252374
rect 437386 252138 437622 252374
rect 437066 215258 437302 215494
rect 437386 215258 437622 215494
rect 437066 214938 437302 215174
rect 437386 214938 437622 215174
rect 437066 178058 437302 178294
rect 437386 178058 437622 178294
rect 437066 177738 437302 177974
rect 437386 177738 437622 177974
rect 437066 140858 437302 141094
rect 437386 140858 437622 141094
rect 437066 140538 437302 140774
rect 437386 140538 437622 140774
rect 437066 103658 437302 103894
rect 437386 103658 437622 103894
rect 437066 103338 437302 103574
rect 437386 103338 437622 103574
rect 437066 66458 437302 66694
rect 437386 66458 437622 66694
rect 437066 66138 437302 66374
rect 437386 66138 437622 66374
rect 437066 29258 437302 29494
rect 437386 29258 437622 29494
rect 437066 28938 437302 29174
rect 437386 28938 437622 29174
rect 448226 672818 448462 673054
rect 448546 672818 448782 673054
rect 448226 672498 448462 672734
rect 448546 672498 448782 672734
rect 448226 635618 448462 635854
rect 448546 635618 448782 635854
rect 448226 635298 448462 635534
rect 448546 635298 448782 635534
rect 448226 598418 448462 598654
rect 448546 598418 448782 598654
rect 448226 598098 448462 598334
rect 448546 598098 448782 598334
rect 448226 561218 448462 561454
rect 448546 561218 448782 561454
rect 448226 560898 448462 561134
rect 448546 560898 448782 561134
rect 448226 524018 448462 524254
rect 448546 524018 448782 524254
rect 448226 523698 448462 523934
rect 448546 523698 448782 523934
rect 448226 486818 448462 487054
rect 448546 486818 448782 487054
rect 448226 486498 448462 486734
rect 448546 486498 448782 486734
rect 448226 449618 448462 449854
rect 448546 449618 448782 449854
rect 448226 449298 448462 449534
rect 448546 449298 448782 449534
rect 448226 412418 448462 412654
rect 448546 412418 448782 412654
rect 448226 412098 448462 412334
rect 448546 412098 448782 412334
rect 448226 375218 448462 375454
rect 448546 375218 448782 375454
rect 448226 374898 448462 375134
rect 448546 374898 448782 375134
rect 448226 338018 448462 338254
rect 448546 338018 448782 338254
rect 448226 337698 448462 337934
rect 448546 337698 448782 337934
rect 448226 300818 448462 301054
rect 448546 300818 448782 301054
rect 448226 300498 448462 300734
rect 448546 300498 448782 300734
rect 448226 263618 448462 263854
rect 448546 263618 448782 263854
rect 448226 263298 448462 263534
rect 448546 263298 448782 263534
rect 448226 226418 448462 226654
rect 448546 226418 448782 226654
rect 448226 226098 448462 226334
rect 448546 226098 448782 226334
rect 448226 189218 448462 189454
rect 448546 189218 448782 189454
rect 448226 188898 448462 189134
rect 448546 188898 448782 189134
rect 448226 152018 448462 152254
rect 448546 152018 448782 152254
rect 448226 151698 448462 151934
rect 448546 151698 448782 151934
rect 448226 114818 448462 115054
rect 448546 114818 448782 115054
rect 448226 114498 448462 114734
rect 448546 114498 448782 114734
rect 448226 77618 448462 77854
rect 448546 77618 448782 77854
rect 448226 77298 448462 77534
rect 448546 77298 448782 77534
rect 448226 40418 448462 40654
rect 448546 40418 448782 40654
rect 448226 40098 448462 40334
rect 448546 40098 448782 40334
rect 448226 3218 448462 3454
rect 448546 3218 448782 3454
rect 448226 2898 448462 3134
rect 448546 2898 448782 3134
rect 451946 676538 452182 676774
rect 452266 676538 452502 676774
rect 451946 676218 452182 676454
rect 452266 676218 452502 676454
rect 451946 639338 452182 639574
rect 452266 639338 452502 639574
rect 451946 639018 452182 639254
rect 452266 639018 452502 639254
rect 451946 602138 452182 602374
rect 452266 602138 452502 602374
rect 451946 601818 452182 602054
rect 452266 601818 452502 602054
rect 451946 564938 452182 565174
rect 452266 564938 452502 565174
rect 451946 564618 452182 564854
rect 452266 564618 452502 564854
rect 451946 527738 452182 527974
rect 452266 527738 452502 527974
rect 451946 527418 452182 527654
rect 452266 527418 452502 527654
rect 451946 490538 452182 490774
rect 452266 490538 452502 490774
rect 451946 490218 452182 490454
rect 452266 490218 452502 490454
rect 451946 453338 452182 453574
rect 452266 453338 452502 453574
rect 451946 453018 452182 453254
rect 452266 453018 452502 453254
rect 451946 416138 452182 416374
rect 452266 416138 452502 416374
rect 451946 415818 452182 416054
rect 452266 415818 452502 416054
rect 451946 378938 452182 379174
rect 452266 378938 452502 379174
rect 451946 378618 452182 378854
rect 452266 378618 452502 378854
rect 451946 341738 452182 341974
rect 452266 341738 452502 341974
rect 451946 341418 452182 341654
rect 452266 341418 452502 341654
rect 451946 304538 452182 304774
rect 452266 304538 452502 304774
rect 451946 304218 452182 304454
rect 452266 304218 452502 304454
rect 451946 267338 452182 267574
rect 452266 267338 452502 267574
rect 451946 267018 452182 267254
rect 452266 267018 452502 267254
rect 451946 230138 452182 230374
rect 452266 230138 452502 230374
rect 451946 229818 452182 230054
rect 452266 229818 452502 230054
rect 451946 192938 452182 193174
rect 452266 192938 452502 193174
rect 451946 192618 452182 192854
rect 452266 192618 452502 192854
rect 451946 155738 452182 155974
rect 452266 155738 452502 155974
rect 451946 155418 452182 155654
rect 452266 155418 452502 155654
rect 451946 118538 452182 118774
rect 452266 118538 452502 118774
rect 451946 118218 452182 118454
rect 452266 118218 452502 118454
rect 451946 81338 452182 81574
rect 452266 81338 452502 81574
rect 451946 81018 452182 81254
rect 452266 81018 452502 81254
rect 451946 44138 452182 44374
rect 452266 44138 452502 44374
rect 451946 43818 452182 44054
rect 452266 43818 452502 44054
rect 451946 6938 452182 7174
rect 452266 6938 452502 7174
rect 451946 6618 452182 6854
rect 452266 6618 452502 6854
rect 455666 680258 455902 680494
rect 455986 680258 456222 680494
rect 455666 679938 455902 680174
rect 455986 679938 456222 680174
rect 455666 643058 455902 643294
rect 455986 643058 456222 643294
rect 455666 642738 455902 642974
rect 455986 642738 456222 642974
rect 455666 605858 455902 606094
rect 455986 605858 456222 606094
rect 455666 605538 455902 605774
rect 455986 605538 456222 605774
rect 455666 568658 455902 568894
rect 455986 568658 456222 568894
rect 455666 568338 455902 568574
rect 455986 568338 456222 568574
rect 455666 531458 455902 531694
rect 455986 531458 456222 531694
rect 455666 531138 455902 531374
rect 455986 531138 456222 531374
rect 455666 494258 455902 494494
rect 455986 494258 456222 494494
rect 455666 493938 455902 494174
rect 455986 493938 456222 494174
rect 455666 457058 455902 457294
rect 455986 457058 456222 457294
rect 455666 456738 455902 456974
rect 455986 456738 456222 456974
rect 455666 419858 455902 420094
rect 455986 419858 456222 420094
rect 455666 419538 455902 419774
rect 455986 419538 456222 419774
rect 455666 382658 455902 382894
rect 455986 382658 456222 382894
rect 455666 382338 455902 382574
rect 455986 382338 456222 382574
rect 455666 345458 455902 345694
rect 455986 345458 456222 345694
rect 455666 345138 455902 345374
rect 455986 345138 456222 345374
rect 455666 308258 455902 308494
rect 455986 308258 456222 308494
rect 455666 307938 455902 308174
rect 455986 307938 456222 308174
rect 455666 271058 455902 271294
rect 455986 271058 456222 271294
rect 455666 270738 455902 270974
rect 455986 270738 456222 270974
rect 455666 233858 455902 234094
rect 455986 233858 456222 234094
rect 455666 233538 455902 233774
rect 455986 233538 456222 233774
rect 455666 196658 455902 196894
rect 455986 196658 456222 196894
rect 455666 196338 455902 196574
rect 455986 196338 456222 196574
rect 455666 159458 455902 159694
rect 455986 159458 456222 159694
rect 455666 159138 455902 159374
rect 455986 159138 456222 159374
rect 455666 122258 455902 122494
rect 455986 122258 456222 122494
rect 455666 121938 455902 122174
rect 455986 121938 456222 122174
rect 455666 85058 455902 85294
rect 455986 85058 456222 85294
rect 455666 84738 455902 84974
rect 455986 84738 456222 84974
rect 455666 47858 455902 48094
rect 455986 47858 456222 48094
rect 455666 47538 455902 47774
rect 455986 47538 456222 47774
rect 455666 10658 455902 10894
rect 455986 10658 456222 10894
rect 455666 10338 455902 10574
rect 455986 10338 456222 10574
rect 459386 683978 459622 684214
rect 459706 683978 459942 684214
rect 459386 683658 459622 683894
rect 459706 683658 459942 683894
rect 459386 646778 459622 647014
rect 459706 646778 459942 647014
rect 459386 646458 459622 646694
rect 459706 646458 459942 646694
rect 459386 609578 459622 609814
rect 459706 609578 459942 609814
rect 459386 609258 459622 609494
rect 459706 609258 459942 609494
rect 459386 572378 459622 572614
rect 459706 572378 459942 572614
rect 459386 572058 459622 572294
rect 459706 572058 459942 572294
rect 459386 535178 459622 535414
rect 459706 535178 459942 535414
rect 459386 534858 459622 535094
rect 459706 534858 459942 535094
rect 459386 497978 459622 498214
rect 459706 497978 459942 498214
rect 459386 497658 459622 497894
rect 459706 497658 459942 497894
rect 459386 460778 459622 461014
rect 459706 460778 459942 461014
rect 459386 460458 459622 460694
rect 459706 460458 459942 460694
rect 459386 423578 459622 423814
rect 459706 423578 459942 423814
rect 459386 423258 459622 423494
rect 459706 423258 459942 423494
rect 459386 386378 459622 386614
rect 459706 386378 459942 386614
rect 459386 386058 459622 386294
rect 459706 386058 459942 386294
rect 459386 349178 459622 349414
rect 459706 349178 459942 349414
rect 459386 348858 459622 349094
rect 459706 348858 459942 349094
rect 459386 311978 459622 312214
rect 459706 311978 459942 312214
rect 459386 311658 459622 311894
rect 459706 311658 459942 311894
rect 459386 274778 459622 275014
rect 459706 274778 459942 275014
rect 459386 274458 459622 274694
rect 459706 274458 459942 274694
rect 459386 237578 459622 237814
rect 459706 237578 459942 237814
rect 459386 237258 459622 237494
rect 459706 237258 459942 237494
rect 459386 200378 459622 200614
rect 459706 200378 459942 200614
rect 459386 200058 459622 200294
rect 459706 200058 459942 200294
rect 459386 163178 459622 163414
rect 459706 163178 459942 163414
rect 459386 162858 459622 163094
rect 459706 162858 459942 163094
rect 459386 125978 459622 126214
rect 459706 125978 459942 126214
rect 459386 125658 459622 125894
rect 459706 125658 459942 125894
rect 459386 88778 459622 89014
rect 459706 88778 459942 89014
rect 459386 88458 459622 88694
rect 459706 88458 459942 88694
rect 459386 51578 459622 51814
rect 459706 51578 459942 51814
rect 459386 51258 459622 51494
rect 459706 51258 459942 51494
rect 459386 14378 459622 14614
rect 459706 14378 459942 14614
rect 459386 14058 459622 14294
rect 459706 14058 459942 14294
rect 463106 687698 463342 687934
rect 463426 687698 463662 687934
rect 463106 687378 463342 687614
rect 463426 687378 463662 687614
rect 463106 650498 463342 650734
rect 463426 650498 463662 650734
rect 463106 650178 463342 650414
rect 463426 650178 463662 650414
rect 463106 613298 463342 613534
rect 463426 613298 463662 613534
rect 463106 612978 463342 613214
rect 463426 612978 463662 613214
rect 463106 576098 463342 576334
rect 463426 576098 463662 576334
rect 463106 575778 463342 576014
rect 463426 575778 463662 576014
rect 463106 538898 463342 539134
rect 463426 538898 463662 539134
rect 463106 538578 463342 538814
rect 463426 538578 463662 538814
rect 463106 501698 463342 501934
rect 463426 501698 463662 501934
rect 463106 501378 463342 501614
rect 463426 501378 463662 501614
rect 463106 464498 463342 464734
rect 463426 464498 463662 464734
rect 463106 464178 463342 464414
rect 463426 464178 463662 464414
rect 463106 427298 463342 427534
rect 463426 427298 463662 427534
rect 463106 426978 463342 427214
rect 463426 426978 463662 427214
rect 463106 390098 463342 390334
rect 463426 390098 463662 390334
rect 463106 389778 463342 390014
rect 463426 389778 463662 390014
rect 463106 352898 463342 353134
rect 463426 352898 463662 353134
rect 463106 352578 463342 352814
rect 463426 352578 463662 352814
rect 463106 315698 463342 315934
rect 463426 315698 463662 315934
rect 463106 315378 463342 315614
rect 463426 315378 463662 315614
rect 463106 278498 463342 278734
rect 463426 278498 463662 278734
rect 463106 278178 463342 278414
rect 463426 278178 463662 278414
rect 463106 241298 463342 241534
rect 463426 241298 463662 241534
rect 463106 240978 463342 241214
rect 463426 240978 463662 241214
rect 463106 204098 463342 204334
rect 463426 204098 463662 204334
rect 463106 203778 463342 204014
rect 463426 203778 463662 204014
rect 463106 166898 463342 167134
rect 463426 166898 463662 167134
rect 463106 166578 463342 166814
rect 463426 166578 463662 166814
rect 463106 129698 463342 129934
rect 463426 129698 463662 129934
rect 463106 129378 463342 129614
rect 463426 129378 463662 129614
rect 463106 92498 463342 92734
rect 463426 92498 463662 92734
rect 463106 92178 463342 92414
rect 463426 92178 463662 92414
rect 463106 55298 463342 55534
rect 463426 55298 463662 55534
rect 463106 54978 463342 55214
rect 463426 54978 463662 55214
rect 463106 18098 463342 18334
rect 463426 18098 463662 18334
rect 463106 17778 463342 18014
rect 463426 17778 463662 18014
rect 466826 691418 467062 691654
rect 467146 691418 467382 691654
rect 466826 691098 467062 691334
rect 467146 691098 467382 691334
rect 466826 654218 467062 654454
rect 467146 654218 467382 654454
rect 466826 653898 467062 654134
rect 467146 653898 467382 654134
rect 466826 617018 467062 617254
rect 467146 617018 467382 617254
rect 466826 616698 467062 616934
rect 467146 616698 467382 616934
rect 466826 579818 467062 580054
rect 467146 579818 467382 580054
rect 466826 579498 467062 579734
rect 467146 579498 467382 579734
rect 466826 542618 467062 542854
rect 467146 542618 467382 542854
rect 466826 542298 467062 542534
rect 467146 542298 467382 542534
rect 466826 505418 467062 505654
rect 467146 505418 467382 505654
rect 466826 505098 467062 505334
rect 467146 505098 467382 505334
rect 466826 468218 467062 468454
rect 467146 468218 467382 468454
rect 466826 467898 467062 468134
rect 467146 467898 467382 468134
rect 466826 431018 467062 431254
rect 467146 431018 467382 431254
rect 466826 430698 467062 430934
rect 467146 430698 467382 430934
rect 466826 393818 467062 394054
rect 467146 393818 467382 394054
rect 466826 393498 467062 393734
rect 467146 393498 467382 393734
rect 466826 356618 467062 356854
rect 467146 356618 467382 356854
rect 466826 356298 467062 356534
rect 467146 356298 467382 356534
rect 466826 319418 467062 319654
rect 467146 319418 467382 319654
rect 466826 319098 467062 319334
rect 467146 319098 467382 319334
rect 466826 282218 467062 282454
rect 467146 282218 467382 282454
rect 466826 281898 467062 282134
rect 467146 281898 467382 282134
rect 466826 245018 467062 245254
rect 467146 245018 467382 245254
rect 466826 244698 467062 244934
rect 467146 244698 467382 244934
rect 466826 207818 467062 208054
rect 467146 207818 467382 208054
rect 466826 207498 467062 207734
rect 467146 207498 467382 207734
rect 466826 170618 467062 170854
rect 467146 170618 467382 170854
rect 466826 170298 467062 170534
rect 467146 170298 467382 170534
rect 466826 133418 467062 133654
rect 467146 133418 467382 133654
rect 466826 133098 467062 133334
rect 467146 133098 467382 133334
rect 466826 96218 467062 96454
rect 467146 96218 467382 96454
rect 466826 95898 467062 96134
rect 467146 95898 467382 96134
rect 466826 59018 467062 59254
rect 467146 59018 467382 59254
rect 466826 58698 467062 58934
rect 467146 58698 467382 58934
rect 466826 21818 467062 22054
rect 467146 21818 467382 22054
rect 466826 21498 467062 21734
rect 467146 21498 467382 21734
rect 470546 695138 470782 695374
rect 470866 695138 471102 695374
rect 470546 694818 470782 695054
rect 470866 694818 471102 695054
rect 470546 657938 470782 658174
rect 470866 657938 471102 658174
rect 470546 657618 470782 657854
rect 470866 657618 471102 657854
rect 470546 620738 470782 620974
rect 470866 620738 471102 620974
rect 470546 620418 470782 620654
rect 470866 620418 471102 620654
rect 470546 583538 470782 583774
rect 470866 583538 471102 583774
rect 470546 583218 470782 583454
rect 470866 583218 471102 583454
rect 470546 546338 470782 546574
rect 470866 546338 471102 546574
rect 470546 546018 470782 546254
rect 470866 546018 471102 546254
rect 470546 509138 470782 509374
rect 470866 509138 471102 509374
rect 470546 508818 470782 509054
rect 470866 508818 471102 509054
rect 470546 471938 470782 472174
rect 470866 471938 471102 472174
rect 470546 471618 470782 471854
rect 470866 471618 471102 471854
rect 470546 434738 470782 434974
rect 470866 434738 471102 434974
rect 470546 434418 470782 434654
rect 470866 434418 471102 434654
rect 470546 397538 470782 397774
rect 470866 397538 471102 397774
rect 470546 397218 470782 397454
rect 470866 397218 471102 397454
rect 470546 360338 470782 360574
rect 470866 360338 471102 360574
rect 470546 360018 470782 360254
rect 470866 360018 471102 360254
rect 470546 323138 470782 323374
rect 470866 323138 471102 323374
rect 470546 322818 470782 323054
rect 470866 322818 471102 323054
rect 470546 285938 470782 286174
rect 470866 285938 471102 286174
rect 470546 285618 470782 285854
rect 470866 285618 471102 285854
rect 470546 248738 470782 248974
rect 470866 248738 471102 248974
rect 470546 248418 470782 248654
rect 470866 248418 471102 248654
rect 470546 211538 470782 211774
rect 470866 211538 471102 211774
rect 470546 211218 470782 211454
rect 470866 211218 471102 211454
rect 470546 174338 470782 174574
rect 470866 174338 471102 174574
rect 470546 174018 470782 174254
rect 470866 174018 471102 174254
rect 470546 137138 470782 137374
rect 470866 137138 471102 137374
rect 470546 136818 470782 137054
rect 470866 136818 471102 137054
rect 470546 99938 470782 100174
rect 470866 99938 471102 100174
rect 470546 99618 470782 99854
rect 470866 99618 471102 99854
rect 470546 62738 470782 62974
rect 470866 62738 471102 62974
rect 470546 62418 470782 62654
rect 470866 62418 471102 62654
rect 470546 25538 470782 25774
rect 470866 25538 471102 25774
rect 470546 25218 470782 25454
rect 470866 25218 471102 25454
rect 474266 698858 474502 699094
rect 474586 698858 474822 699094
rect 474266 698538 474502 698774
rect 474586 698538 474822 698774
rect 474266 661658 474502 661894
rect 474586 661658 474822 661894
rect 474266 661338 474502 661574
rect 474586 661338 474822 661574
rect 474266 624458 474502 624694
rect 474586 624458 474822 624694
rect 474266 624138 474502 624374
rect 474586 624138 474822 624374
rect 474266 587258 474502 587494
rect 474586 587258 474822 587494
rect 474266 586938 474502 587174
rect 474586 586938 474822 587174
rect 474266 550058 474502 550294
rect 474586 550058 474822 550294
rect 474266 549738 474502 549974
rect 474586 549738 474822 549974
rect 474266 512858 474502 513094
rect 474586 512858 474822 513094
rect 474266 512538 474502 512774
rect 474586 512538 474822 512774
rect 474266 475658 474502 475894
rect 474586 475658 474822 475894
rect 474266 475338 474502 475574
rect 474586 475338 474822 475574
rect 474266 438458 474502 438694
rect 474586 438458 474822 438694
rect 474266 438138 474502 438374
rect 474586 438138 474822 438374
rect 474266 401258 474502 401494
rect 474586 401258 474822 401494
rect 474266 400938 474502 401174
rect 474586 400938 474822 401174
rect 474266 364058 474502 364294
rect 474586 364058 474822 364294
rect 474266 363738 474502 363974
rect 474586 363738 474822 363974
rect 485426 672818 485662 673054
rect 485746 672818 485982 673054
rect 485426 672498 485662 672734
rect 485746 672498 485982 672734
rect 485426 635618 485662 635854
rect 485746 635618 485982 635854
rect 485426 635298 485662 635534
rect 485746 635298 485982 635534
rect 485426 598418 485662 598654
rect 485746 598418 485982 598654
rect 485426 598098 485662 598334
rect 485746 598098 485982 598334
rect 485426 561218 485662 561454
rect 485746 561218 485982 561454
rect 485426 560898 485662 561134
rect 485746 560898 485982 561134
rect 485426 524018 485662 524254
rect 485746 524018 485982 524254
rect 485426 523698 485662 523934
rect 485746 523698 485982 523934
rect 485426 486818 485662 487054
rect 485746 486818 485982 487054
rect 485426 486498 485662 486734
rect 485746 486498 485982 486734
rect 485426 449618 485662 449854
rect 485746 449618 485982 449854
rect 485426 449298 485662 449534
rect 485746 449298 485982 449534
rect 485426 412418 485662 412654
rect 485746 412418 485982 412654
rect 485426 412098 485662 412334
rect 485746 412098 485982 412334
rect 485426 375218 485662 375454
rect 485746 375218 485982 375454
rect 485426 374898 485662 375134
rect 485746 374898 485982 375134
rect 489146 676538 489382 676774
rect 489466 676538 489702 676774
rect 489146 676218 489382 676454
rect 489466 676218 489702 676454
rect 489146 639338 489382 639574
rect 489466 639338 489702 639574
rect 489146 639018 489382 639254
rect 489466 639018 489702 639254
rect 489146 602138 489382 602374
rect 489466 602138 489702 602374
rect 489146 601818 489382 602054
rect 489466 601818 489702 602054
rect 489146 564938 489382 565174
rect 489466 564938 489702 565174
rect 489146 564618 489382 564854
rect 489466 564618 489702 564854
rect 489146 527738 489382 527974
rect 489466 527738 489702 527974
rect 489146 527418 489382 527654
rect 489466 527418 489702 527654
rect 489146 490538 489382 490774
rect 489466 490538 489702 490774
rect 489146 490218 489382 490454
rect 489466 490218 489702 490454
rect 489146 453338 489382 453574
rect 489466 453338 489702 453574
rect 489146 453018 489382 453254
rect 489466 453018 489702 453254
rect 489146 416138 489382 416374
rect 489466 416138 489702 416374
rect 489146 415818 489382 416054
rect 489466 415818 489702 416054
rect 489146 378938 489382 379174
rect 489466 378938 489702 379174
rect 489146 378618 489382 378854
rect 489466 378618 489702 378854
rect 489146 341738 489382 341974
rect 489466 341738 489702 341974
rect 489146 341418 489382 341654
rect 489466 341418 489702 341654
rect 492866 680258 493102 680494
rect 493186 680258 493422 680494
rect 492866 679938 493102 680174
rect 493186 679938 493422 680174
rect 492866 643058 493102 643294
rect 493186 643058 493422 643294
rect 492866 642738 493102 642974
rect 493186 642738 493422 642974
rect 492866 605858 493102 606094
rect 493186 605858 493422 606094
rect 492866 605538 493102 605774
rect 493186 605538 493422 605774
rect 492866 568658 493102 568894
rect 493186 568658 493422 568894
rect 492866 568338 493102 568574
rect 493186 568338 493422 568574
rect 492866 531458 493102 531694
rect 493186 531458 493422 531694
rect 492866 531138 493102 531374
rect 493186 531138 493422 531374
rect 492866 494258 493102 494494
rect 493186 494258 493422 494494
rect 492866 493938 493102 494174
rect 493186 493938 493422 494174
rect 492866 457058 493102 457294
rect 493186 457058 493422 457294
rect 492866 456738 493102 456974
rect 493186 456738 493422 456974
rect 492866 419858 493102 420094
rect 493186 419858 493422 420094
rect 492866 419538 493102 419774
rect 493186 419538 493422 419774
rect 492866 382658 493102 382894
rect 493186 382658 493422 382894
rect 492866 382338 493102 382574
rect 493186 382338 493422 382574
rect 492866 345458 493102 345694
rect 493186 345458 493422 345694
rect 492866 345138 493102 345374
rect 493186 345138 493422 345374
rect 481952 338018 482188 338254
rect 481952 337698 482188 337934
rect 483884 338018 484120 338254
rect 483884 337698 484120 337934
rect 485816 338018 486052 338254
rect 485816 337698 486052 337934
rect 487748 338018 487984 338254
rect 487748 337698 487984 337934
rect 474266 326858 474502 327094
rect 474586 326858 474822 327094
rect 474266 326538 474502 326774
rect 474586 326538 474822 326774
rect 474266 289658 474502 289894
rect 474586 289658 474822 289894
rect 474266 289338 474502 289574
rect 474586 289338 474822 289574
rect 474266 252458 474502 252694
rect 474586 252458 474822 252694
rect 474266 252138 474502 252374
rect 474586 252138 474822 252374
rect 474266 215258 474502 215494
rect 474586 215258 474822 215494
rect 474266 214938 474502 215174
rect 474586 214938 474822 215174
rect 474266 178058 474502 178294
rect 474586 178058 474822 178294
rect 474266 177738 474502 177974
rect 474586 177738 474822 177974
rect 474266 140858 474502 141094
rect 474586 140858 474822 141094
rect 474266 140538 474502 140774
rect 474586 140538 474822 140774
rect 474266 103658 474502 103894
rect 474586 103658 474822 103894
rect 474266 103338 474502 103574
rect 474586 103338 474822 103574
rect 474266 66458 474502 66694
rect 474586 66458 474822 66694
rect 474266 66138 474502 66374
rect 474586 66138 474822 66374
rect 474266 29258 474502 29494
rect 474586 29258 474822 29494
rect 474266 28938 474502 29174
rect 474586 28938 474822 29174
rect 485426 300818 485662 301054
rect 485746 300818 485982 301054
rect 485426 300498 485662 300734
rect 485746 300498 485982 300734
rect 485426 263618 485662 263854
rect 485746 263618 485982 263854
rect 485426 263298 485662 263534
rect 485746 263298 485982 263534
rect 485426 226418 485662 226654
rect 485746 226418 485982 226654
rect 485426 226098 485662 226334
rect 485746 226098 485982 226334
rect 485426 189218 485662 189454
rect 485746 189218 485982 189454
rect 485426 188898 485662 189134
rect 485746 188898 485982 189134
rect 485426 152018 485662 152254
rect 485746 152018 485982 152254
rect 485426 151698 485662 151934
rect 485746 151698 485982 151934
rect 485426 114818 485662 115054
rect 485746 114818 485982 115054
rect 485426 114498 485662 114734
rect 485746 114498 485982 114734
rect 485426 77618 485662 77854
rect 485746 77618 485982 77854
rect 485426 77298 485662 77534
rect 485746 77298 485982 77534
rect 485426 40418 485662 40654
rect 485746 40418 485982 40654
rect 485426 40098 485662 40334
rect 485746 40098 485982 40334
rect 485426 3218 485662 3454
rect 485746 3218 485982 3454
rect 485426 2898 485662 3134
rect 485746 2898 485982 3134
rect 489146 304538 489382 304774
rect 489466 304538 489702 304774
rect 489146 304218 489382 304454
rect 489466 304218 489702 304454
rect 489146 267338 489382 267574
rect 489466 267338 489702 267574
rect 489146 267018 489382 267254
rect 489466 267018 489702 267254
rect 489146 230138 489382 230374
rect 489466 230138 489702 230374
rect 489146 229818 489382 230054
rect 489466 229818 489702 230054
rect 489146 192938 489382 193174
rect 489466 192938 489702 193174
rect 489146 192618 489382 192854
rect 489466 192618 489702 192854
rect 489146 155738 489382 155974
rect 489466 155738 489702 155974
rect 489146 155418 489382 155654
rect 489466 155418 489702 155654
rect 489146 118538 489382 118774
rect 489466 118538 489702 118774
rect 489146 118218 489382 118454
rect 489466 118218 489702 118454
rect 489146 81338 489382 81574
rect 489466 81338 489702 81574
rect 489146 81018 489382 81254
rect 489466 81018 489702 81254
rect 489146 44138 489382 44374
rect 489466 44138 489702 44374
rect 489146 43818 489382 44054
rect 489466 43818 489702 44054
rect 492866 308258 493102 308494
rect 493186 308258 493422 308494
rect 492866 307938 493102 308174
rect 493186 307938 493422 308174
rect 492866 271058 493102 271294
rect 493186 271058 493422 271294
rect 492866 270738 493102 270974
rect 493186 270738 493422 270974
rect 492866 233858 493102 234094
rect 493186 233858 493422 234094
rect 492866 233538 493102 233774
rect 493186 233538 493422 233774
rect 492866 196658 493102 196894
rect 493186 196658 493422 196894
rect 492866 196338 493102 196574
rect 493186 196338 493422 196574
rect 492866 159458 493102 159694
rect 493186 159458 493422 159694
rect 492866 159138 493102 159374
rect 493186 159138 493422 159374
rect 492866 122258 493102 122494
rect 493186 122258 493422 122494
rect 492866 121938 493102 122174
rect 493186 121938 493422 122174
rect 492866 85058 493102 85294
rect 493186 85058 493422 85294
rect 492866 84738 493102 84974
rect 493186 84738 493422 84974
rect 492866 47858 493102 48094
rect 493186 47858 493422 48094
rect 492866 47538 493102 47774
rect 493186 47538 493422 47774
rect 489146 6938 489382 7174
rect 489466 6938 489702 7174
rect 489146 6618 489382 6854
rect 489466 6618 489702 6854
rect 492866 10658 493102 10894
rect 493186 10658 493422 10894
rect 492866 10338 493102 10574
rect 493186 10338 493422 10574
rect 496586 683978 496822 684214
rect 496906 683978 497142 684214
rect 496586 683658 496822 683894
rect 496906 683658 497142 683894
rect 496586 646778 496822 647014
rect 496906 646778 497142 647014
rect 496586 646458 496822 646694
rect 496906 646458 497142 646694
rect 496586 609578 496822 609814
rect 496906 609578 497142 609814
rect 496586 609258 496822 609494
rect 496906 609258 497142 609494
rect 496586 572378 496822 572614
rect 496906 572378 497142 572614
rect 496586 572058 496822 572294
rect 496906 572058 497142 572294
rect 496586 535178 496822 535414
rect 496906 535178 497142 535414
rect 496586 534858 496822 535094
rect 496906 534858 497142 535094
rect 496586 497978 496822 498214
rect 496906 497978 497142 498214
rect 496586 497658 496822 497894
rect 496906 497658 497142 497894
rect 496586 460778 496822 461014
rect 496906 460778 497142 461014
rect 496586 460458 496822 460694
rect 496906 460458 497142 460694
rect 496586 423578 496822 423814
rect 496906 423578 497142 423814
rect 496586 423258 496822 423494
rect 496906 423258 497142 423494
rect 496586 386378 496822 386614
rect 496906 386378 497142 386614
rect 496586 386058 496822 386294
rect 496906 386058 497142 386294
rect 496586 349178 496822 349414
rect 496906 349178 497142 349414
rect 496586 348858 496822 349094
rect 496906 348858 497142 349094
rect 496586 311978 496822 312214
rect 496906 311978 497142 312214
rect 496586 311658 496822 311894
rect 496906 311658 497142 311894
rect 496586 274778 496822 275014
rect 496906 274778 497142 275014
rect 496586 274458 496822 274694
rect 496906 274458 497142 274694
rect 496586 237578 496822 237814
rect 496906 237578 497142 237814
rect 496586 237258 496822 237494
rect 496906 237258 497142 237494
rect 496586 200378 496822 200614
rect 496906 200378 497142 200614
rect 496586 200058 496822 200294
rect 496906 200058 497142 200294
rect 496586 163178 496822 163414
rect 496906 163178 497142 163414
rect 496586 162858 496822 163094
rect 496906 162858 497142 163094
rect 496586 125978 496822 126214
rect 496906 125978 497142 126214
rect 496586 125658 496822 125894
rect 496906 125658 497142 125894
rect 496586 88778 496822 89014
rect 496906 88778 497142 89014
rect 496586 88458 496822 88694
rect 496906 88458 497142 88694
rect 496586 51578 496822 51814
rect 496906 51578 497142 51814
rect 496586 51258 496822 51494
rect 496906 51258 497142 51494
rect 496586 14378 496822 14614
rect 496906 14378 497142 14614
rect 496586 14058 496822 14294
rect 496906 14058 497142 14294
rect 500306 687698 500542 687934
rect 500626 687698 500862 687934
rect 500306 687378 500542 687614
rect 500626 687378 500862 687614
rect 500306 650498 500542 650734
rect 500626 650498 500862 650734
rect 500306 650178 500542 650414
rect 500626 650178 500862 650414
rect 500306 613298 500542 613534
rect 500626 613298 500862 613534
rect 500306 612978 500542 613214
rect 500626 612978 500862 613214
rect 500306 576098 500542 576334
rect 500626 576098 500862 576334
rect 500306 575778 500542 576014
rect 500626 575778 500862 576014
rect 500306 538898 500542 539134
rect 500626 538898 500862 539134
rect 500306 538578 500542 538814
rect 500626 538578 500862 538814
rect 500306 501698 500542 501934
rect 500626 501698 500862 501934
rect 500306 501378 500542 501614
rect 500626 501378 500862 501614
rect 500306 464498 500542 464734
rect 500626 464498 500862 464734
rect 500306 464178 500542 464414
rect 500626 464178 500862 464414
rect 500306 427298 500542 427534
rect 500626 427298 500862 427534
rect 500306 426978 500542 427214
rect 500626 426978 500862 427214
rect 500306 390098 500542 390334
rect 500626 390098 500862 390334
rect 500306 389778 500542 390014
rect 500626 389778 500862 390014
rect 500306 352898 500542 353134
rect 500626 352898 500862 353134
rect 500306 352578 500542 352814
rect 500626 352578 500862 352814
rect 500306 315698 500542 315934
rect 500626 315698 500862 315934
rect 500306 315378 500542 315614
rect 500626 315378 500862 315614
rect 500306 278498 500542 278734
rect 500626 278498 500862 278734
rect 500306 278178 500542 278414
rect 500626 278178 500862 278414
rect 500306 241298 500542 241534
rect 500626 241298 500862 241534
rect 500306 240978 500542 241214
rect 500626 240978 500862 241214
rect 500306 204098 500542 204334
rect 500626 204098 500862 204334
rect 500306 203778 500542 204014
rect 500626 203778 500862 204014
rect 500306 166898 500542 167134
rect 500626 166898 500862 167134
rect 500306 166578 500542 166814
rect 500626 166578 500862 166814
rect 500306 129698 500542 129934
rect 500626 129698 500862 129934
rect 500306 129378 500542 129614
rect 500626 129378 500862 129614
rect 500306 92498 500542 92734
rect 500626 92498 500862 92734
rect 500306 92178 500542 92414
rect 500626 92178 500862 92414
rect 500306 55298 500542 55534
rect 500626 55298 500862 55534
rect 500306 54978 500542 55214
rect 500626 54978 500862 55214
rect 500306 18098 500542 18334
rect 500626 18098 500862 18334
rect 500306 17778 500542 18014
rect 500626 17778 500862 18014
rect 504026 691418 504262 691654
rect 504346 691418 504582 691654
rect 504026 691098 504262 691334
rect 504346 691098 504582 691334
rect 504026 654218 504262 654454
rect 504346 654218 504582 654454
rect 504026 653898 504262 654134
rect 504346 653898 504582 654134
rect 504026 617018 504262 617254
rect 504346 617018 504582 617254
rect 504026 616698 504262 616934
rect 504346 616698 504582 616934
rect 504026 579818 504262 580054
rect 504346 579818 504582 580054
rect 504026 579498 504262 579734
rect 504346 579498 504582 579734
rect 504026 542618 504262 542854
rect 504346 542618 504582 542854
rect 504026 542298 504262 542534
rect 504346 542298 504582 542534
rect 504026 505418 504262 505654
rect 504346 505418 504582 505654
rect 504026 505098 504262 505334
rect 504346 505098 504582 505334
rect 504026 468218 504262 468454
rect 504346 468218 504582 468454
rect 504026 467898 504262 468134
rect 504346 467898 504582 468134
rect 504026 431018 504262 431254
rect 504346 431018 504582 431254
rect 504026 430698 504262 430934
rect 504346 430698 504582 430934
rect 504026 393818 504262 394054
rect 504346 393818 504582 394054
rect 504026 393498 504262 393734
rect 504346 393498 504582 393734
rect 504026 356618 504262 356854
rect 504346 356618 504582 356854
rect 504026 356298 504262 356534
rect 504346 356298 504582 356534
rect 504026 319418 504262 319654
rect 504346 319418 504582 319654
rect 504026 319098 504262 319334
rect 504346 319098 504582 319334
rect 504026 282218 504262 282454
rect 504346 282218 504582 282454
rect 504026 281898 504262 282134
rect 504346 281898 504582 282134
rect 504026 245018 504262 245254
rect 504346 245018 504582 245254
rect 504026 244698 504262 244934
rect 504346 244698 504582 244934
rect 504026 207818 504262 208054
rect 504346 207818 504582 208054
rect 504026 207498 504262 207734
rect 504346 207498 504582 207734
rect 504026 170618 504262 170854
rect 504346 170618 504582 170854
rect 504026 170298 504262 170534
rect 504346 170298 504582 170534
rect 504026 133418 504262 133654
rect 504346 133418 504582 133654
rect 504026 133098 504262 133334
rect 504346 133098 504582 133334
rect 504026 96218 504262 96454
rect 504346 96218 504582 96454
rect 504026 95898 504262 96134
rect 504346 95898 504582 96134
rect 504026 59018 504262 59254
rect 504346 59018 504582 59254
rect 504026 58698 504262 58934
rect 504346 58698 504582 58934
rect 504026 21818 504262 22054
rect 504346 21818 504582 22054
rect 504026 21498 504262 21734
rect 504346 21498 504582 21734
rect 507746 695138 507982 695374
rect 508066 695138 508302 695374
rect 507746 694818 507982 695054
rect 508066 694818 508302 695054
rect 507746 657938 507982 658174
rect 508066 657938 508302 658174
rect 507746 657618 507982 657854
rect 508066 657618 508302 657854
rect 507746 620738 507982 620974
rect 508066 620738 508302 620974
rect 507746 620418 507982 620654
rect 508066 620418 508302 620654
rect 507746 583538 507982 583774
rect 508066 583538 508302 583774
rect 507746 583218 507982 583454
rect 508066 583218 508302 583454
rect 507746 546338 507982 546574
rect 508066 546338 508302 546574
rect 507746 546018 507982 546254
rect 508066 546018 508302 546254
rect 507746 509138 507982 509374
rect 508066 509138 508302 509374
rect 507746 508818 507982 509054
rect 508066 508818 508302 509054
rect 507746 471938 507982 472174
rect 508066 471938 508302 472174
rect 507746 471618 507982 471854
rect 508066 471618 508302 471854
rect 507746 434738 507982 434974
rect 508066 434738 508302 434974
rect 507746 434418 507982 434654
rect 508066 434418 508302 434654
rect 507746 397538 507982 397774
rect 508066 397538 508302 397774
rect 507746 397218 507982 397454
rect 508066 397218 508302 397454
rect 507746 360338 507982 360574
rect 508066 360338 508302 360574
rect 507746 360018 507982 360254
rect 508066 360018 508302 360254
rect 507746 323138 507982 323374
rect 508066 323138 508302 323374
rect 507746 322818 507982 323054
rect 508066 322818 508302 323054
rect 507746 285938 507982 286174
rect 508066 285938 508302 286174
rect 507746 285618 507982 285854
rect 508066 285618 508302 285854
rect 507746 248738 507982 248974
rect 508066 248738 508302 248974
rect 507746 248418 507982 248654
rect 508066 248418 508302 248654
rect 507746 211538 507982 211774
rect 508066 211538 508302 211774
rect 507746 211218 507982 211454
rect 508066 211218 508302 211454
rect 507746 174338 507982 174574
rect 508066 174338 508302 174574
rect 507746 174018 507982 174254
rect 508066 174018 508302 174254
rect 507746 137138 507982 137374
rect 508066 137138 508302 137374
rect 507746 136818 507982 137054
rect 508066 136818 508302 137054
rect 507746 99938 507982 100174
rect 508066 99938 508302 100174
rect 507746 99618 507982 99854
rect 508066 99618 508302 99854
rect 507746 62738 507982 62974
rect 508066 62738 508302 62974
rect 507746 62418 507982 62654
rect 508066 62418 508302 62654
rect 507746 25538 507982 25774
rect 508066 25538 508302 25774
rect 507746 25218 507982 25454
rect 508066 25218 508302 25454
rect 511466 698858 511702 699094
rect 511786 698858 512022 699094
rect 511466 698538 511702 698774
rect 511786 698538 512022 698774
rect 511466 661658 511702 661894
rect 511786 661658 512022 661894
rect 511466 661338 511702 661574
rect 511786 661338 512022 661574
rect 511466 624458 511702 624694
rect 511786 624458 512022 624694
rect 511466 624138 511702 624374
rect 511786 624138 512022 624374
rect 511466 587258 511702 587494
rect 511786 587258 512022 587494
rect 511466 586938 511702 587174
rect 511786 586938 512022 587174
rect 511466 550058 511702 550294
rect 511786 550058 512022 550294
rect 511466 549738 511702 549974
rect 511786 549738 512022 549974
rect 511466 512858 511702 513094
rect 511786 512858 512022 513094
rect 511466 512538 511702 512774
rect 511786 512538 512022 512774
rect 511466 475658 511702 475894
rect 511786 475658 512022 475894
rect 511466 475338 511702 475574
rect 511786 475338 512022 475574
rect 511466 438458 511702 438694
rect 511786 438458 512022 438694
rect 511466 438138 511702 438374
rect 511786 438138 512022 438374
rect 511466 401258 511702 401494
rect 511786 401258 512022 401494
rect 511466 400938 511702 401174
rect 511786 400938 512022 401174
rect 511466 364058 511702 364294
rect 511786 364058 512022 364294
rect 511466 363738 511702 363974
rect 511786 363738 512022 363974
rect 511466 326858 511702 327094
rect 511786 326858 512022 327094
rect 511466 326538 511702 326774
rect 511786 326538 512022 326774
rect 511466 289658 511702 289894
rect 511786 289658 512022 289894
rect 511466 289338 511702 289574
rect 511786 289338 512022 289574
rect 511466 252458 511702 252694
rect 511786 252458 512022 252694
rect 511466 252138 511702 252374
rect 511786 252138 512022 252374
rect 511466 215258 511702 215494
rect 511786 215258 512022 215494
rect 511466 214938 511702 215174
rect 511786 214938 512022 215174
rect 511466 178058 511702 178294
rect 511786 178058 512022 178294
rect 511466 177738 511702 177974
rect 511786 177738 512022 177974
rect 511466 140858 511702 141094
rect 511786 140858 512022 141094
rect 511466 140538 511702 140774
rect 511786 140538 512022 140774
rect 511466 103658 511702 103894
rect 511786 103658 512022 103894
rect 511466 103338 511702 103574
rect 511786 103338 512022 103574
rect 511466 66458 511702 66694
rect 511786 66458 512022 66694
rect 511466 66138 511702 66374
rect 511786 66138 512022 66374
rect 511466 29258 511702 29494
rect 511786 29258 512022 29494
rect 511466 28938 511702 29174
rect 511786 28938 512022 29174
rect 522626 672818 522862 673054
rect 522946 672818 523182 673054
rect 522626 672498 522862 672734
rect 522946 672498 523182 672734
rect 522626 635618 522862 635854
rect 522946 635618 523182 635854
rect 522626 635298 522862 635534
rect 522946 635298 523182 635534
rect 522626 598418 522862 598654
rect 522946 598418 523182 598654
rect 522626 598098 522862 598334
rect 522946 598098 523182 598334
rect 522626 561218 522862 561454
rect 522946 561218 523182 561454
rect 522626 560898 522862 561134
rect 522946 560898 523182 561134
rect 522626 524018 522862 524254
rect 522946 524018 523182 524254
rect 522626 523698 522862 523934
rect 522946 523698 523182 523934
rect 522626 486818 522862 487054
rect 522946 486818 523182 487054
rect 522626 486498 522862 486734
rect 522946 486498 523182 486734
rect 522626 449618 522862 449854
rect 522946 449618 523182 449854
rect 522626 449298 522862 449534
rect 522946 449298 523182 449534
rect 522626 412418 522862 412654
rect 522946 412418 523182 412654
rect 522626 412098 522862 412334
rect 522946 412098 523182 412334
rect 522626 375218 522862 375454
rect 522946 375218 523182 375454
rect 522626 374898 522862 375134
rect 522946 374898 523182 375134
rect 522626 338018 522862 338254
rect 522946 338018 523182 338254
rect 522626 337698 522862 337934
rect 522946 337698 523182 337934
rect 522626 300818 522862 301054
rect 522946 300818 523182 301054
rect 522626 300498 522862 300734
rect 522946 300498 523182 300734
rect 522626 263618 522862 263854
rect 522946 263618 523182 263854
rect 522626 263298 522862 263534
rect 522946 263298 523182 263534
rect 522626 226418 522862 226654
rect 522946 226418 523182 226654
rect 522626 226098 522862 226334
rect 522946 226098 523182 226334
rect 522626 189218 522862 189454
rect 522946 189218 523182 189454
rect 522626 188898 522862 189134
rect 522946 188898 523182 189134
rect 522626 152018 522862 152254
rect 522946 152018 523182 152254
rect 522626 151698 522862 151934
rect 522946 151698 523182 151934
rect 522626 114818 522862 115054
rect 522946 114818 523182 115054
rect 522626 114498 522862 114734
rect 522946 114498 523182 114734
rect 522626 77618 522862 77854
rect 522946 77618 523182 77854
rect 522626 77298 522862 77534
rect 522946 77298 523182 77534
rect 522626 40418 522862 40654
rect 522946 40418 523182 40654
rect 522626 40098 522862 40334
rect 522946 40098 523182 40334
rect 522626 3218 522862 3454
rect 522946 3218 523182 3454
rect 522626 2898 522862 3134
rect 522946 2898 523182 3134
rect 526346 676538 526582 676774
rect 526666 676538 526902 676774
rect 526346 676218 526582 676454
rect 526666 676218 526902 676454
rect 526346 639338 526582 639574
rect 526666 639338 526902 639574
rect 526346 639018 526582 639254
rect 526666 639018 526902 639254
rect 526346 602138 526582 602374
rect 526666 602138 526902 602374
rect 526346 601818 526582 602054
rect 526666 601818 526902 602054
rect 526346 564938 526582 565174
rect 526666 564938 526902 565174
rect 526346 564618 526582 564854
rect 526666 564618 526902 564854
rect 526346 527738 526582 527974
rect 526666 527738 526902 527974
rect 526346 527418 526582 527654
rect 526666 527418 526902 527654
rect 526346 490538 526582 490774
rect 526666 490538 526902 490774
rect 526346 490218 526582 490454
rect 526666 490218 526902 490454
rect 526346 453338 526582 453574
rect 526666 453338 526902 453574
rect 526346 453018 526582 453254
rect 526666 453018 526902 453254
rect 526346 416138 526582 416374
rect 526666 416138 526902 416374
rect 526346 415818 526582 416054
rect 526666 415818 526902 416054
rect 526346 378938 526582 379174
rect 526666 378938 526902 379174
rect 526346 378618 526582 378854
rect 526666 378618 526902 378854
rect 526346 341738 526582 341974
rect 526666 341738 526902 341974
rect 526346 341418 526582 341654
rect 526666 341418 526902 341654
rect 526346 304538 526582 304774
rect 526666 304538 526902 304774
rect 526346 304218 526582 304454
rect 526666 304218 526902 304454
rect 526346 267338 526582 267574
rect 526666 267338 526902 267574
rect 526346 267018 526582 267254
rect 526666 267018 526902 267254
rect 526346 230138 526582 230374
rect 526666 230138 526902 230374
rect 526346 229818 526582 230054
rect 526666 229818 526902 230054
rect 526346 192938 526582 193174
rect 526666 192938 526902 193174
rect 526346 192618 526582 192854
rect 526666 192618 526902 192854
rect 526346 155738 526582 155974
rect 526666 155738 526902 155974
rect 526346 155418 526582 155654
rect 526666 155418 526902 155654
rect 526346 118538 526582 118774
rect 526666 118538 526902 118774
rect 526346 118218 526582 118454
rect 526666 118218 526902 118454
rect 526346 81338 526582 81574
rect 526666 81338 526902 81574
rect 526346 81018 526582 81254
rect 526666 81018 526902 81254
rect 526346 44138 526582 44374
rect 526666 44138 526902 44374
rect 526346 43818 526582 44054
rect 526666 43818 526902 44054
rect 526346 6938 526582 7174
rect 526666 6938 526902 7174
rect 526346 6618 526582 6854
rect 526666 6618 526902 6854
rect 530066 680258 530302 680494
rect 530386 680258 530622 680494
rect 530066 679938 530302 680174
rect 530386 679938 530622 680174
rect 530066 643058 530302 643294
rect 530386 643058 530622 643294
rect 530066 642738 530302 642974
rect 530386 642738 530622 642974
rect 530066 605858 530302 606094
rect 530386 605858 530622 606094
rect 530066 605538 530302 605774
rect 530386 605538 530622 605774
rect 530066 568658 530302 568894
rect 530386 568658 530622 568894
rect 530066 568338 530302 568574
rect 530386 568338 530622 568574
rect 530066 531458 530302 531694
rect 530386 531458 530622 531694
rect 530066 531138 530302 531374
rect 530386 531138 530622 531374
rect 530066 494258 530302 494494
rect 530386 494258 530622 494494
rect 530066 493938 530302 494174
rect 530386 493938 530622 494174
rect 530066 457058 530302 457294
rect 530386 457058 530622 457294
rect 530066 456738 530302 456974
rect 530386 456738 530622 456974
rect 530066 419858 530302 420094
rect 530386 419858 530622 420094
rect 530066 419538 530302 419774
rect 530386 419538 530622 419774
rect 530066 382658 530302 382894
rect 530386 382658 530622 382894
rect 530066 382338 530302 382574
rect 530386 382338 530622 382574
rect 530066 345458 530302 345694
rect 530386 345458 530622 345694
rect 530066 345138 530302 345374
rect 530386 345138 530622 345374
rect 530066 308258 530302 308494
rect 530386 308258 530622 308494
rect 530066 307938 530302 308174
rect 530386 307938 530622 308174
rect 530066 271058 530302 271294
rect 530386 271058 530622 271294
rect 530066 270738 530302 270974
rect 530386 270738 530622 270974
rect 530066 233858 530302 234094
rect 530386 233858 530622 234094
rect 530066 233538 530302 233774
rect 530386 233538 530622 233774
rect 530066 196658 530302 196894
rect 530386 196658 530622 196894
rect 530066 196338 530302 196574
rect 530386 196338 530622 196574
rect 530066 159458 530302 159694
rect 530386 159458 530622 159694
rect 530066 159138 530302 159374
rect 530386 159138 530622 159374
rect 530066 122258 530302 122494
rect 530386 122258 530622 122494
rect 530066 121938 530302 122174
rect 530386 121938 530622 122174
rect 530066 85058 530302 85294
rect 530386 85058 530622 85294
rect 530066 84738 530302 84974
rect 530386 84738 530622 84974
rect 530066 47858 530302 48094
rect 530386 47858 530622 48094
rect 530066 47538 530302 47774
rect 530386 47538 530622 47774
rect 530066 10658 530302 10894
rect 530386 10658 530622 10894
rect 530066 10338 530302 10574
rect 530386 10338 530622 10574
rect 533786 683978 534022 684214
rect 534106 683978 534342 684214
rect 533786 683658 534022 683894
rect 534106 683658 534342 683894
rect 533786 646778 534022 647014
rect 534106 646778 534342 647014
rect 533786 646458 534022 646694
rect 534106 646458 534342 646694
rect 533786 609578 534022 609814
rect 534106 609578 534342 609814
rect 533786 609258 534022 609494
rect 534106 609258 534342 609494
rect 533786 572378 534022 572614
rect 534106 572378 534342 572614
rect 533786 572058 534022 572294
rect 534106 572058 534342 572294
rect 533786 535178 534022 535414
rect 534106 535178 534342 535414
rect 533786 534858 534022 535094
rect 534106 534858 534342 535094
rect 533786 497978 534022 498214
rect 534106 497978 534342 498214
rect 533786 497658 534022 497894
rect 534106 497658 534342 497894
rect 533786 460778 534022 461014
rect 534106 460778 534342 461014
rect 533786 460458 534022 460694
rect 534106 460458 534342 460694
rect 533786 423578 534022 423814
rect 534106 423578 534342 423814
rect 533786 423258 534022 423494
rect 534106 423258 534342 423494
rect 533786 386378 534022 386614
rect 534106 386378 534342 386614
rect 533786 386058 534022 386294
rect 534106 386058 534342 386294
rect 533786 349178 534022 349414
rect 534106 349178 534342 349414
rect 533786 348858 534022 349094
rect 534106 348858 534342 349094
rect 533786 311978 534022 312214
rect 534106 311978 534342 312214
rect 533786 311658 534022 311894
rect 534106 311658 534342 311894
rect 533786 274778 534022 275014
rect 534106 274778 534342 275014
rect 533786 274458 534022 274694
rect 534106 274458 534342 274694
rect 533786 237578 534022 237814
rect 534106 237578 534342 237814
rect 533786 237258 534022 237494
rect 534106 237258 534342 237494
rect 533786 200378 534022 200614
rect 534106 200378 534342 200614
rect 533786 200058 534022 200294
rect 534106 200058 534342 200294
rect 533786 163178 534022 163414
rect 534106 163178 534342 163414
rect 533786 162858 534022 163094
rect 534106 162858 534342 163094
rect 533786 125978 534022 126214
rect 534106 125978 534342 126214
rect 533786 125658 534022 125894
rect 534106 125658 534342 125894
rect 533786 88778 534022 89014
rect 534106 88778 534342 89014
rect 533786 88458 534022 88694
rect 534106 88458 534342 88694
rect 533786 51578 534022 51814
rect 534106 51578 534342 51814
rect 533786 51258 534022 51494
rect 534106 51258 534342 51494
rect 533786 14378 534022 14614
rect 534106 14378 534342 14614
rect 533786 14058 534022 14294
rect 534106 14058 534342 14294
rect 537506 687698 537742 687934
rect 537826 687698 538062 687934
rect 537506 687378 537742 687614
rect 537826 687378 538062 687614
rect 537506 650498 537742 650734
rect 537826 650498 538062 650734
rect 537506 650178 537742 650414
rect 537826 650178 538062 650414
rect 537506 613298 537742 613534
rect 537826 613298 538062 613534
rect 537506 612978 537742 613214
rect 537826 612978 538062 613214
rect 537506 576098 537742 576334
rect 537826 576098 538062 576334
rect 537506 575778 537742 576014
rect 537826 575778 538062 576014
rect 537506 538898 537742 539134
rect 537826 538898 538062 539134
rect 537506 538578 537742 538814
rect 537826 538578 538062 538814
rect 537506 501698 537742 501934
rect 537826 501698 538062 501934
rect 537506 501378 537742 501614
rect 537826 501378 538062 501614
rect 537506 464498 537742 464734
rect 537826 464498 538062 464734
rect 537506 464178 537742 464414
rect 537826 464178 538062 464414
rect 537506 427298 537742 427534
rect 537826 427298 538062 427534
rect 537506 426978 537742 427214
rect 537826 426978 538062 427214
rect 537506 390098 537742 390334
rect 537826 390098 538062 390334
rect 537506 389778 537742 390014
rect 537826 389778 538062 390014
rect 537506 352898 537742 353134
rect 537826 352898 538062 353134
rect 537506 352578 537742 352814
rect 537826 352578 538062 352814
rect 537506 315698 537742 315934
rect 537826 315698 538062 315934
rect 537506 315378 537742 315614
rect 537826 315378 538062 315614
rect 537506 278498 537742 278734
rect 537826 278498 538062 278734
rect 537506 278178 537742 278414
rect 537826 278178 538062 278414
rect 537506 241298 537742 241534
rect 537826 241298 538062 241534
rect 537506 240978 537742 241214
rect 537826 240978 538062 241214
rect 537506 204098 537742 204334
rect 537826 204098 538062 204334
rect 537506 203778 537742 204014
rect 537826 203778 538062 204014
rect 537506 166898 537742 167134
rect 537826 166898 538062 167134
rect 537506 166578 537742 166814
rect 537826 166578 538062 166814
rect 537506 129698 537742 129934
rect 537826 129698 538062 129934
rect 537506 129378 537742 129614
rect 537826 129378 538062 129614
rect 537506 92498 537742 92734
rect 537826 92498 538062 92734
rect 537506 92178 537742 92414
rect 537826 92178 538062 92414
rect 537506 55298 537742 55534
rect 537826 55298 538062 55534
rect 537506 54978 537742 55214
rect 537826 54978 538062 55214
rect 537506 18098 537742 18334
rect 537826 18098 538062 18334
rect 537506 17778 537742 18014
rect 537826 17778 538062 18014
rect 541226 691418 541462 691654
rect 541546 691418 541782 691654
rect 541226 691098 541462 691334
rect 541546 691098 541782 691334
rect 541226 654218 541462 654454
rect 541546 654218 541782 654454
rect 541226 653898 541462 654134
rect 541546 653898 541782 654134
rect 541226 617018 541462 617254
rect 541546 617018 541782 617254
rect 541226 616698 541462 616934
rect 541546 616698 541782 616934
rect 541226 579818 541462 580054
rect 541546 579818 541782 580054
rect 541226 579498 541462 579734
rect 541546 579498 541782 579734
rect 541226 542618 541462 542854
rect 541546 542618 541782 542854
rect 541226 542298 541462 542534
rect 541546 542298 541782 542534
rect 541226 505418 541462 505654
rect 541546 505418 541782 505654
rect 541226 505098 541462 505334
rect 541546 505098 541782 505334
rect 541226 468218 541462 468454
rect 541546 468218 541782 468454
rect 541226 467898 541462 468134
rect 541546 467898 541782 468134
rect 541226 431018 541462 431254
rect 541546 431018 541782 431254
rect 541226 430698 541462 430934
rect 541546 430698 541782 430934
rect 541226 393818 541462 394054
rect 541546 393818 541782 394054
rect 541226 393498 541462 393734
rect 541546 393498 541782 393734
rect 541226 356618 541462 356854
rect 541546 356618 541782 356854
rect 541226 356298 541462 356534
rect 541546 356298 541782 356534
rect 541226 319418 541462 319654
rect 541546 319418 541782 319654
rect 541226 319098 541462 319334
rect 541546 319098 541782 319334
rect 541226 282218 541462 282454
rect 541546 282218 541782 282454
rect 541226 281898 541462 282134
rect 541546 281898 541782 282134
rect 541226 245018 541462 245254
rect 541546 245018 541782 245254
rect 541226 244698 541462 244934
rect 541546 244698 541782 244934
rect 541226 207818 541462 208054
rect 541546 207818 541782 208054
rect 541226 207498 541462 207734
rect 541546 207498 541782 207734
rect 541226 170618 541462 170854
rect 541546 170618 541782 170854
rect 541226 170298 541462 170534
rect 541546 170298 541782 170534
rect 541226 133418 541462 133654
rect 541546 133418 541782 133654
rect 541226 133098 541462 133334
rect 541546 133098 541782 133334
rect 541226 96218 541462 96454
rect 541546 96218 541782 96454
rect 541226 95898 541462 96134
rect 541546 95898 541782 96134
rect 541226 59018 541462 59254
rect 541546 59018 541782 59254
rect 541226 58698 541462 58934
rect 541546 58698 541782 58934
rect 541226 21818 541462 22054
rect 541546 21818 541782 22054
rect 541226 21498 541462 21734
rect 541546 21498 541782 21734
rect 544946 695138 545182 695374
rect 545266 695138 545502 695374
rect 544946 694818 545182 695054
rect 545266 694818 545502 695054
rect 544946 657938 545182 658174
rect 545266 657938 545502 658174
rect 544946 657618 545182 657854
rect 545266 657618 545502 657854
rect 544946 620738 545182 620974
rect 545266 620738 545502 620974
rect 544946 620418 545182 620654
rect 545266 620418 545502 620654
rect 544946 583538 545182 583774
rect 545266 583538 545502 583774
rect 544946 583218 545182 583454
rect 545266 583218 545502 583454
rect 544946 546338 545182 546574
rect 545266 546338 545502 546574
rect 544946 546018 545182 546254
rect 545266 546018 545502 546254
rect 544946 509138 545182 509374
rect 545266 509138 545502 509374
rect 544946 508818 545182 509054
rect 545266 508818 545502 509054
rect 544946 471938 545182 472174
rect 545266 471938 545502 472174
rect 544946 471618 545182 471854
rect 545266 471618 545502 471854
rect 544946 434738 545182 434974
rect 545266 434738 545502 434974
rect 544946 434418 545182 434654
rect 545266 434418 545502 434654
rect 544946 397538 545182 397774
rect 545266 397538 545502 397774
rect 544946 397218 545182 397454
rect 545266 397218 545502 397454
rect 544946 360338 545182 360574
rect 545266 360338 545502 360574
rect 544946 360018 545182 360254
rect 545266 360018 545502 360254
rect 544946 323138 545182 323374
rect 545266 323138 545502 323374
rect 544946 322818 545182 323054
rect 545266 322818 545502 323054
rect 544946 285938 545182 286174
rect 545266 285938 545502 286174
rect 544946 285618 545182 285854
rect 545266 285618 545502 285854
rect 544946 248738 545182 248974
rect 545266 248738 545502 248974
rect 544946 248418 545182 248654
rect 545266 248418 545502 248654
rect 544946 211538 545182 211774
rect 545266 211538 545502 211774
rect 544946 211218 545182 211454
rect 545266 211218 545502 211454
rect 544946 174338 545182 174574
rect 545266 174338 545502 174574
rect 544946 174018 545182 174254
rect 545266 174018 545502 174254
rect 544946 137138 545182 137374
rect 545266 137138 545502 137374
rect 544946 136818 545182 137054
rect 545266 136818 545502 137054
rect 544946 99938 545182 100174
rect 545266 99938 545502 100174
rect 544946 99618 545182 99854
rect 545266 99618 545502 99854
rect 544946 62738 545182 62974
rect 545266 62738 545502 62974
rect 544946 62418 545182 62654
rect 545266 62418 545502 62654
rect 544946 25538 545182 25774
rect 545266 25538 545502 25774
rect 544946 25218 545182 25454
rect 545266 25218 545502 25454
rect 548666 698858 548902 699094
rect 548986 698858 549222 699094
rect 548666 698538 548902 698774
rect 548986 698538 549222 698774
rect 548666 661658 548902 661894
rect 548986 661658 549222 661894
rect 548666 661338 548902 661574
rect 548986 661338 549222 661574
rect 548666 624458 548902 624694
rect 548986 624458 549222 624694
rect 548666 624138 548902 624374
rect 548986 624138 549222 624374
rect 548666 587258 548902 587494
rect 548986 587258 549222 587494
rect 548666 586938 548902 587174
rect 548986 586938 549222 587174
rect 548666 550058 548902 550294
rect 548986 550058 549222 550294
rect 548666 549738 548902 549974
rect 548986 549738 549222 549974
rect 548666 512858 548902 513094
rect 548986 512858 549222 513094
rect 548666 512538 548902 512774
rect 548986 512538 549222 512774
rect 548666 475658 548902 475894
rect 548986 475658 549222 475894
rect 548666 475338 548902 475574
rect 548986 475338 549222 475574
rect 548666 438458 548902 438694
rect 548986 438458 549222 438694
rect 548666 438138 548902 438374
rect 548986 438138 549222 438374
rect 548666 401258 548902 401494
rect 548986 401258 549222 401494
rect 548666 400938 548902 401174
rect 548986 400938 549222 401174
rect 548666 364058 548902 364294
rect 548986 364058 549222 364294
rect 548666 363738 548902 363974
rect 548986 363738 549222 363974
rect 548666 326858 548902 327094
rect 548986 326858 549222 327094
rect 548666 326538 548902 326774
rect 548986 326538 549222 326774
rect 548666 289658 548902 289894
rect 548986 289658 549222 289894
rect 548666 289338 548902 289574
rect 548986 289338 549222 289574
rect 548666 252458 548902 252694
rect 548986 252458 549222 252694
rect 548666 252138 548902 252374
rect 548986 252138 549222 252374
rect 548666 215258 548902 215494
rect 548986 215258 549222 215494
rect 548666 214938 548902 215174
rect 548986 214938 549222 215174
rect 548666 178058 548902 178294
rect 548986 178058 549222 178294
rect 548666 177738 548902 177974
rect 548986 177738 549222 177974
rect 548666 140858 548902 141094
rect 548986 140858 549222 141094
rect 548666 140538 548902 140774
rect 548986 140538 549222 140774
rect 548666 103658 548902 103894
rect 548986 103658 549222 103894
rect 548666 103338 548902 103574
rect 548986 103338 549222 103574
rect 548666 66458 548902 66694
rect 548986 66458 549222 66694
rect 548666 66138 548902 66374
rect 548986 66138 549222 66374
rect 548666 29258 548902 29494
rect 548986 29258 549222 29494
rect 548666 28938 548902 29174
rect 548986 28938 549222 29174
rect 559826 672818 560062 673054
rect 560146 672818 560382 673054
rect 559826 672498 560062 672734
rect 560146 672498 560382 672734
rect 559826 635618 560062 635854
rect 560146 635618 560382 635854
rect 559826 635298 560062 635534
rect 560146 635298 560382 635534
rect 559826 598418 560062 598654
rect 560146 598418 560382 598654
rect 559826 598098 560062 598334
rect 560146 598098 560382 598334
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 524018 560062 524254
rect 560146 524018 560382 524254
rect 559826 523698 560062 523934
rect 560146 523698 560382 523934
rect 559826 486818 560062 487054
rect 560146 486818 560382 487054
rect 559826 486498 560062 486734
rect 560146 486498 560382 486734
rect 559826 449618 560062 449854
rect 560146 449618 560382 449854
rect 559826 449298 560062 449534
rect 560146 449298 560382 449534
rect 559826 412418 560062 412654
rect 560146 412418 560382 412654
rect 559826 412098 560062 412334
rect 560146 412098 560382 412334
rect 559826 375218 560062 375454
rect 560146 375218 560382 375454
rect 559826 374898 560062 375134
rect 560146 374898 560382 375134
rect 559826 338018 560062 338254
rect 560146 338018 560382 338254
rect 559826 337698 560062 337934
rect 560146 337698 560382 337934
rect 559826 300818 560062 301054
rect 560146 300818 560382 301054
rect 559826 300498 560062 300734
rect 560146 300498 560382 300734
rect 559826 263618 560062 263854
rect 560146 263618 560382 263854
rect 559826 263298 560062 263534
rect 560146 263298 560382 263534
rect 559826 226418 560062 226654
rect 560146 226418 560382 226654
rect 559826 226098 560062 226334
rect 560146 226098 560382 226334
rect 559826 189218 560062 189454
rect 560146 189218 560382 189454
rect 559826 188898 560062 189134
rect 560146 188898 560382 189134
rect 559826 152018 560062 152254
rect 560146 152018 560382 152254
rect 559826 151698 560062 151934
rect 560146 151698 560382 151934
rect 559826 114818 560062 115054
rect 560146 114818 560382 115054
rect 559826 114498 560062 114734
rect 560146 114498 560382 114734
rect 559826 77618 560062 77854
rect 560146 77618 560382 77854
rect 559826 77298 560062 77534
rect 560146 77298 560382 77534
rect 559826 40418 560062 40654
rect 560146 40418 560382 40654
rect 559826 40098 560062 40334
rect 560146 40098 560382 40334
rect 559826 3218 560062 3454
rect 560146 3218 560382 3454
rect 559826 2898 560062 3134
rect 560146 2898 560382 3134
rect 563546 676538 563782 676774
rect 563866 676538 564102 676774
rect 563546 676218 563782 676454
rect 563866 676218 564102 676454
rect 563546 639338 563782 639574
rect 563866 639338 564102 639574
rect 563546 639018 563782 639254
rect 563866 639018 564102 639254
rect 563546 602138 563782 602374
rect 563866 602138 564102 602374
rect 563546 601818 563782 602054
rect 563866 601818 564102 602054
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 527738 563782 527974
rect 563866 527738 564102 527974
rect 563546 527418 563782 527654
rect 563866 527418 564102 527654
rect 563546 490538 563782 490774
rect 563866 490538 564102 490774
rect 563546 490218 563782 490454
rect 563866 490218 564102 490454
rect 563546 453338 563782 453574
rect 563866 453338 564102 453574
rect 563546 453018 563782 453254
rect 563866 453018 564102 453254
rect 563546 416138 563782 416374
rect 563866 416138 564102 416374
rect 563546 415818 563782 416054
rect 563866 415818 564102 416054
rect 563546 378938 563782 379174
rect 563866 378938 564102 379174
rect 563546 378618 563782 378854
rect 563866 378618 564102 378854
rect 563546 341738 563782 341974
rect 563866 341738 564102 341974
rect 563546 341418 563782 341654
rect 563866 341418 564102 341654
rect 563546 304538 563782 304774
rect 563866 304538 564102 304774
rect 563546 304218 563782 304454
rect 563866 304218 564102 304454
rect 563546 267338 563782 267574
rect 563866 267338 564102 267574
rect 563546 267018 563782 267254
rect 563866 267018 564102 267254
rect 563546 230138 563782 230374
rect 563866 230138 564102 230374
rect 563546 229818 563782 230054
rect 563866 229818 564102 230054
rect 563546 192938 563782 193174
rect 563866 192938 564102 193174
rect 563546 192618 563782 192854
rect 563866 192618 564102 192854
rect 563546 155738 563782 155974
rect 563866 155738 564102 155974
rect 563546 155418 563782 155654
rect 563866 155418 564102 155654
rect 563546 118538 563782 118774
rect 563866 118538 564102 118774
rect 563546 118218 563782 118454
rect 563866 118218 564102 118454
rect 563546 81338 563782 81574
rect 563866 81338 564102 81574
rect 563546 81018 563782 81254
rect 563866 81018 564102 81254
rect 563546 44138 563782 44374
rect 563866 44138 564102 44374
rect 563546 43818 563782 44054
rect 563866 43818 564102 44054
rect 563546 6938 563782 7174
rect 563866 6938 564102 7174
rect 563546 6618 563782 6854
rect 563866 6618 564102 6854
rect 567266 680258 567502 680494
rect 567586 680258 567822 680494
rect 567266 679938 567502 680174
rect 567586 679938 567822 680174
rect 567266 643058 567502 643294
rect 567586 643058 567822 643294
rect 567266 642738 567502 642974
rect 567586 642738 567822 642974
rect 567266 605858 567502 606094
rect 567586 605858 567822 606094
rect 567266 605538 567502 605774
rect 567586 605538 567822 605774
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 531458 567502 531694
rect 567586 531458 567822 531694
rect 567266 531138 567502 531374
rect 567586 531138 567822 531374
rect 567266 494258 567502 494494
rect 567586 494258 567822 494494
rect 567266 493938 567502 494174
rect 567586 493938 567822 494174
rect 567266 457058 567502 457294
rect 567586 457058 567822 457294
rect 567266 456738 567502 456974
rect 567586 456738 567822 456974
rect 567266 419858 567502 420094
rect 567586 419858 567822 420094
rect 567266 419538 567502 419774
rect 567586 419538 567822 419774
rect 567266 382658 567502 382894
rect 567586 382658 567822 382894
rect 567266 382338 567502 382574
rect 567586 382338 567822 382574
rect 567266 345458 567502 345694
rect 567586 345458 567822 345694
rect 567266 345138 567502 345374
rect 567586 345138 567822 345374
rect 567266 308258 567502 308494
rect 567586 308258 567822 308494
rect 567266 307938 567502 308174
rect 567586 307938 567822 308174
rect 567266 271058 567502 271294
rect 567586 271058 567822 271294
rect 567266 270738 567502 270974
rect 567586 270738 567822 270974
rect 567266 233858 567502 234094
rect 567586 233858 567822 234094
rect 567266 233538 567502 233774
rect 567586 233538 567822 233774
rect 567266 196658 567502 196894
rect 567586 196658 567822 196894
rect 567266 196338 567502 196574
rect 567586 196338 567822 196574
rect 567266 159458 567502 159694
rect 567586 159458 567822 159694
rect 567266 159138 567502 159374
rect 567586 159138 567822 159374
rect 567266 122258 567502 122494
rect 567586 122258 567822 122494
rect 567266 121938 567502 122174
rect 567586 121938 567822 122174
rect 567266 85058 567502 85294
rect 567586 85058 567822 85294
rect 567266 84738 567502 84974
rect 567586 84738 567822 84974
rect 567266 47858 567502 48094
rect 567586 47858 567822 48094
rect 567266 47538 567502 47774
rect 567586 47538 567822 47774
rect 567266 10658 567502 10894
rect 567586 10658 567822 10894
rect 567266 10338 567502 10574
rect 567586 10338 567822 10574
rect 570986 683978 571222 684214
rect 571306 683978 571542 684214
rect 570986 683658 571222 683894
rect 571306 683658 571542 683894
rect 570986 646778 571222 647014
rect 571306 646778 571542 647014
rect 570986 646458 571222 646694
rect 571306 646458 571542 646694
rect 570986 609578 571222 609814
rect 571306 609578 571542 609814
rect 570986 609258 571222 609494
rect 571306 609258 571542 609494
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 535178 571222 535414
rect 571306 535178 571542 535414
rect 570986 534858 571222 535094
rect 571306 534858 571542 535094
rect 570986 497978 571222 498214
rect 571306 497978 571542 498214
rect 570986 497658 571222 497894
rect 571306 497658 571542 497894
rect 570986 460778 571222 461014
rect 571306 460778 571542 461014
rect 570986 460458 571222 460694
rect 571306 460458 571542 460694
rect 570986 423578 571222 423814
rect 571306 423578 571542 423814
rect 570986 423258 571222 423494
rect 571306 423258 571542 423494
rect 570986 386378 571222 386614
rect 571306 386378 571542 386614
rect 570986 386058 571222 386294
rect 571306 386058 571542 386294
rect 570986 349178 571222 349414
rect 571306 349178 571542 349414
rect 570986 348858 571222 349094
rect 571306 348858 571542 349094
rect 570986 311978 571222 312214
rect 571306 311978 571542 312214
rect 570986 311658 571222 311894
rect 571306 311658 571542 311894
rect 570986 274778 571222 275014
rect 571306 274778 571542 275014
rect 570986 274458 571222 274694
rect 571306 274458 571542 274694
rect 570986 237578 571222 237814
rect 571306 237578 571542 237814
rect 570986 237258 571222 237494
rect 571306 237258 571542 237494
rect 570986 200378 571222 200614
rect 571306 200378 571542 200614
rect 570986 200058 571222 200294
rect 571306 200058 571542 200294
rect 570986 163178 571222 163414
rect 571306 163178 571542 163414
rect 570986 162858 571222 163094
rect 571306 162858 571542 163094
rect 570986 125978 571222 126214
rect 571306 125978 571542 126214
rect 570986 125658 571222 125894
rect 571306 125658 571542 125894
rect 570986 88778 571222 89014
rect 571306 88778 571542 89014
rect 570986 88458 571222 88694
rect 571306 88458 571542 88694
rect 570986 51578 571222 51814
rect 571306 51578 571542 51814
rect 570986 51258 571222 51494
rect 571306 51258 571542 51494
rect 570986 14378 571222 14614
rect 571306 14378 571542 14614
rect 570986 14058 571222 14294
rect 571306 14058 571542 14294
rect 574706 687698 574942 687934
rect 575026 687698 575262 687934
rect 574706 687378 574942 687614
rect 575026 687378 575262 687614
rect 574706 650498 574942 650734
rect 575026 650498 575262 650734
rect 574706 650178 574942 650414
rect 575026 650178 575262 650414
rect 574706 613298 574942 613534
rect 575026 613298 575262 613534
rect 574706 612978 574942 613214
rect 575026 612978 575262 613214
rect 574706 576098 574942 576334
rect 575026 576098 575262 576334
rect 574706 575778 574942 576014
rect 575026 575778 575262 576014
rect 574706 538898 574942 539134
rect 575026 538898 575262 539134
rect 574706 538578 574942 538814
rect 575026 538578 575262 538814
rect 574706 501698 574942 501934
rect 575026 501698 575262 501934
rect 574706 501378 574942 501614
rect 575026 501378 575262 501614
rect 574706 464498 574942 464734
rect 575026 464498 575262 464734
rect 574706 464178 574942 464414
rect 575026 464178 575262 464414
rect 574706 427298 574942 427534
rect 575026 427298 575262 427534
rect 574706 426978 574942 427214
rect 575026 426978 575262 427214
rect 574706 390098 574942 390334
rect 575026 390098 575262 390334
rect 574706 389778 574942 390014
rect 575026 389778 575262 390014
rect 574706 352898 574942 353134
rect 575026 352898 575262 353134
rect 574706 352578 574942 352814
rect 575026 352578 575262 352814
rect 574706 315698 574942 315934
rect 575026 315698 575262 315934
rect 574706 315378 574942 315614
rect 575026 315378 575262 315614
rect 574706 278498 574942 278734
rect 575026 278498 575262 278734
rect 574706 278178 574942 278414
rect 575026 278178 575262 278414
rect 574706 241298 574942 241534
rect 575026 241298 575262 241534
rect 574706 240978 574942 241214
rect 575026 240978 575262 241214
rect 574706 204098 574942 204334
rect 575026 204098 575262 204334
rect 574706 203778 574942 204014
rect 575026 203778 575262 204014
rect 574706 166898 574942 167134
rect 575026 166898 575262 167134
rect 574706 166578 574942 166814
rect 575026 166578 575262 166814
rect 574706 129698 574942 129934
rect 575026 129698 575262 129934
rect 574706 129378 574942 129614
rect 575026 129378 575262 129614
rect 574706 92498 574942 92734
rect 575026 92498 575262 92734
rect 574706 92178 574942 92414
rect 575026 92178 575262 92414
rect 574706 55298 574942 55534
rect 575026 55298 575262 55534
rect 574706 54978 574942 55214
rect 575026 54978 575262 55214
rect 574706 18098 574942 18334
rect 575026 18098 575262 18334
rect 574706 17778 574942 18014
rect 575026 17778 575262 18014
rect 578426 691418 578662 691654
rect 578746 691418 578982 691654
rect 578426 691098 578662 691334
rect 578746 691098 578982 691334
rect 578426 654218 578662 654454
rect 578746 654218 578982 654454
rect 578426 653898 578662 654134
rect 578746 653898 578982 654134
rect 578426 617018 578662 617254
rect 578746 617018 578982 617254
rect 578426 616698 578662 616934
rect 578746 616698 578982 616934
rect 578426 579818 578662 580054
rect 578746 579818 578982 580054
rect 578426 579498 578662 579734
rect 578746 579498 578982 579734
rect 578426 542618 578662 542854
rect 578746 542618 578982 542854
rect 578426 542298 578662 542534
rect 578746 542298 578982 542534
rect 578426 505418 578662 505654
rect 578746 505418 578982 505654
rect 578426 505098 578662 505334
rect 578746 505098 578982 505334
rect 578426 468218 578662 468454
rect 578746 468218 578982 468454
rect 578426 467898 578662 468134
rect 578746 467898 578982 468134
rect 578426 431018 578662 431254
rect 578746 431018 578982 431254
rect 578426 430698 578662 430934
rect 578746 430698 578982 430934
rect 578426 393818 578662 394054
rect 578746 393818 578982 394054
rect 578426 393498 578662 393734
rect 578746 393498 578982 393734
rect 578426 356618 578662 356854
rect 578746 356618 578982 356854
rect 578426 356298 578662 356534
rect 578746 356298 578982 356534
rect 578426 319418 578662 319654
rect 578746 319418 578982 319654
rect 578426 319098 578662 319334
rect 578746 319098 578982 319334
rect 578426 282218 578662 282454
rect 578746 282218 578982 282454
rect 578426 281898 578662 282134
rect 578746 281898 578982 282134
rect 578426 245018 578662 245254
rect 578746 245018 578982 245254
rect 578426 244698 578662 244934
rect 578746 244698 578982 244934
rect 578426 207818 578662 208054
rect 578746 207818 578982 208054
rect 578426 207498 578662 207734
rect 578746 207498 578982 207734
rect 578426 170618 578662 170854
rect 578746 170618 578982 170854
rect 578426 170298 578662 170534
rect 578746 170298 578982 170534
rect 578426 133418 578662 133654
rect 578746 133418 578982 133654
rect 578426 133098 578662 133334
rect 578746 133098 578982 133334
rect 578426 96218 578662 96454
rect 578746 96218 578982 96454
rect 578426 95898 578662 96134
rect 578746 95898 578982 96134
rect 578426 59018 578662 59254
rect 578746 59018 578982 59254
rect 578426 58698 578662 58934
rect 578746 58698 578982 58934
rect 578426 21818 578662 22054
rect 578746 21818 578982 22054
rect 578426 21498 578662 21734
rect 578746 21498 578982 21734
rect 582146 695138 582382 695374
rect 582466 695138 582702 695374
rect 582146 694818 582382 695054
rect 582466 694818 582702 695054
rect 582146 657938 582382 658174
rect 582466 657938 582702 658174
rect 582146 657618 582382 657854
rect 582466 657618 582702 657854
rect 582146 620738 582382 620974
rect 582466 620738 582702 620974
rect 582146 620418 582382 620654
rect 582466 620418 582702 620654
rect 582146 583538 582382 583774
rect 582466 583538 582702 583774
rect 582146 583218 582382 583454
rect 582466 583218 582702 583454
rect 582146 546338 582382 546574
rect 582466 546338 582702 546574
rect 582146 546018 582382 546254
rect 582466 546018 582702 546254
rect 582146 509138 582382 509374
rect 582466 509138 582702 509374
rect 582146 508818 582382 509054
rect 582466 508818 582702 509054
rect 582146 471938 582382 472174
rect 582466 471938 582702 472174
rect 582146 471618 582382 471854
rect 582466 471618 582702 471854
rect 582146 434738 582382 434974
rect 582466 434738 582702 434974
rect 582146 434418 582382 434654
rect 582466 434418 582702 434654
rect 582146 397538 582382 397774
rect 582466 397538 582702 397774
rect 582146 397218 582382 397454
rect 582466 397218 582702 397454
rect 582146 360338 582382 360574
rect 582466 360338 582702 360574
rect 582146 360018 582382 360254
rect 582466 360018 582702 360254
rect 582146 323138 582382 323374
rect 582466 323138 582702 323374
rect 582146 322818 582382 323054
rect 582466 322818 582702 323054
rect 582146 285938 582382 286174
rect 582466 285938 582702 286174
rect 582146 285618 582382 285854
rect 582466 285618 582702 285854
rect 582146 248738 582382 248974
rect 582466 248738 582702 248974
rect 582146 248418 582382 248654
rect 582466 248418 582702 248654
rect 582146 211538 582382 211774
rect 582466 211538 582702 211774
rect 582146 211218 582382 211454
rect 582466 211218 582702 211454
rect 582146 174338 582382 174574
rect 582466 174338 582702 174574
rect 582146 174018 582382 174254
rect 582466 174018 582702 174254
rect 582146 137138 582382 137374
rect 582466 137138 582702 137374
rect 582146 136818 582382 137054
rect 582466 136818 582702 137054
rect 582146 99938 582382 100174
rect 582466 99938 582702 100174
rect 582146 99618 582382 99854
rect 582466 99618 582702 99854
rect 582146 62738 582382 62974
rect 582466 62738 582702 62974
rect 582146 62418 582382 62654
rect 582466 62418 582702 62654
rect 582146 25538 582382 25774
rect 582466 25538 582702 25774
rect 582146 25218 582382 25454
rect 582466 25218 582702 25454
<< metal5 >>
rect 1104 699094 582820 699126
rect 1104 698858 27866 699094
rect 28102 698858 28186 699094
rect 28422 698858 65066 699094
rect 65302 698858 65386 699094
rect 65622 698858 102266 699094
rect 102502 698858 102586 699094
rect 102822 698858 139466 699094
rect 139702 698858 139786 699094
rect 140022 698858 176666 699094
rect 176902 698858 176986 699094
rect 177222 698858 213866 699094
rect 214102 698858 214186 699094
rect 214422 698858 251066 699094
rect 251302 698858 251386 699094
rect 251622 698858 288266 699094
rect 288502 698858 288586 699094
rect 288822 698858 325466 699094
rect 325702 698858 325786 699094
rect 326022 698858 362666 699094
rect 362902 698858 362986 699094
rect 363222 698858 399866 699094
rect 400102 698858 400186 699094
rect 400422 698858 437066 699094
rect 437302 698858 437386 699094
rect 437622 698858 474266 699094
rect 474502 698858 474586 699094
rect 474822 698858 511466 699094
rect 511702 698858 511786 699094
rect 512022 698858 548666 699094
rect 548902 698858 548986 699094
rect 549222 698858 582820 699094
rect 1104 698774 582820 698858
rect 1104 698538 27866 698774
rect 28102 698538 28186 698774
rect 28422 698538 65066 698774
rect 65302 698538 65386 698774
rect 65622 698538 102266 698774
rect 102502 698538 102586 698774
rect 102822 698538 139466 698774
rect 139702 698538 139786 698774
rect 140022 698538 176666 698774
rect 176902 698538 176986 698774
rect 177222 698538 213866 698774
rect 214102 698538 214186 698774
rect 214422 698538 251066 698774
rect 251302 698538 251386 698774
rect 251622 698538 288266 698774
rect 288502 698538 288586 698774
rect 288822 698538 325466 698774
rect 325702 698538 325786 698774
rect 326022 698538 362666 698774
rect 362902 698538 362986 698774
rect 363222 698538 399866 698774
rect 400102 698538 400186 698774
rect 400422 698538 437066 698774
rect 437302 698538 437386 698774
rect 437622 698538 474266 698774
rect 474502 698538 474586 698774
rect 474822 698538 511466 698774
rect 511702 698538 511786 698774
rect 512022 698538 548666 698774
rect 548902 698538 548986 698774
rect 549222 698538 582820 698774
rect 1104 698506 582820 698538
rect 1104 695374 582820 695406
rect 1104 695138 24146 695374
rect 24382 695138 24466 695374
rect 24702 695138 61346 695374
rect 61582 695138 61666 695374
rect 61902 695138 98546 695374
rect 98782 695138 98866 695374
rect 99102 695138 135746 695374
rect 135982 695138 136066 695374
rect 136302 695138 172946 695374
rect 173182 695138 173266 695374
rect 173502 695138 210146 695374
rect 210382 695138 210466 695374
rect 210702 695138 247346 695374
rect 247582 695138 247666 695374
rect 247902 695138 284546 695374
rect 284782 695138 284866 695374
rect 285102 695138 321746 695374
rect 321982 695138 322066 695374
rect 322302 695138 358946 695374
rect 359182 695138 359266 695374
rect 359502 695138 396146 695374
rect 396382 695138 396466 695374
rect 396702 695138 433346 695374
rect 433582 695138 433666 695374
rect 433902 695138 470546 695374
rect 470782 695138 470866 695374
rect 471102 695138 507746 695374
rect 507982 695138 508066 695374
rect 508302 695138 544946 695374
rect 545182 695138 545266 695374
rect 545502 695138 582146 695374
rect 582382 695138 582466 695374
rect 582702 695138 582820 695374
rect 1104 695054 582820 695138
rect 1104 694818 24146 695054
rect 24382 694818 24466 695054
rect 24702 694818 61346 695054
rect 61582 694818 61666 695054
rect 61902 694818 98546 695054
rect 98782 694818 98866 695054
rect 99102 694818 135746 695054
rect 135982 694818 136066 695054
rect 136302 694818 172946 695054
rect 173182 694818 173266 695054
rect 173502 694818 210146 695054
rect 210382 694818 210466 695054
rect 210702 694818 247346 695054
rect 247582 694818 247666 695054
rect 247902 694818 284546 695054
rect 284782 694818 284866 695054
rect 285102 694818 321746 695054
rect 321982 694818 322066 695054
rect 322302 694818 358946 695054
rect 359182 694818 359266 695054
rect 359502 694818 396146 695054
rect 396382 694818 396466 695054
rect 396702 694818 433346 695054
rect 433582 694818 433666 695054
rect 433902 694818 470546 695054
rect 470782 694818 470866 695054
rect 471102 694818 507746 695054
rect 507982 694818 508066 695054
rect 508302 694818 544946 695054
rect 545182 694818 545266 695054
rect 545502 694818 582146 695054
rect 582382 694818 582466 695054
rect 582702 694818 582820 695054
rect 1104 694786 582820 694818
rect 1104 691654 582820 691686
rect 1104 691418 20426 691654
rect 20662 691418 20746 691654
rect 20982 691418 57626 691654
rect 57862 691418 57946 691654
rect 58182 691418 94826 691654
rect 95062 691418 95146 691654
rect 95382 691418 132026 691654
rect 132262 691418 132346 691654
rect 132582 691418 169226 691654
rect 169462 691418 169546 691654
rect 169782 691418 206426 691654
rect 206662 691418 206746 691654
rect 206982 691418 243626 691654
rect 243862 691418 243946 691654
rect 244182 691418 280826 691654
rect 281062 691418 281146 691654
rect 281382 691418 318026 691654
rect 318262 691418 318346 691654
rect 318582 691418 355226 691654
rect 355462 691418 355546 691654
rect 355782 691418 392426 691654
rect 392662 691418 392746 691654
rect 392982 691418 429626 691654
rect 429862 691418 429946 691654
rect 430182 691418 466826 691654
rect 467062 691418 467146 691654
rect 467382 691418 504026 691654
rect 504262 691418 504346 691654
rect 504582 691418 541226 691654
rect 541462 691418 541546 691654
rect 541782 691418 578426 691654
rect 578662 691418 578746 691654
rect 578982 691418 582820 691654
rect 1104 691334 582820 691418
rect 1104 691098 20426 691334
rect 20662 691098 20746 691334
rect 20982 691098 57626 691334
rect 57862 691098 57946 691334
rect 58182 691098 94826 691334
rect 95062 691098 95146 691334
rect 95382 691098 132026 691334
rect 132262 691098 132346 691334
rect 132582 691098 169226 691334
rect 169462 691098 169546 691334
rect 169782 691098 206426 691334
rect 206662 691098 206746 691334
rect 206982 691098 243626 691334
rect 243862 691098 243946 691334
rect 244182 691098 280826 691334
rect 281062 691098 281146 691334
rect 281382 691098 318026 691334
rect 318262 691098 318346 691334
rect 318582 691098 355226 691334
rect 355462 691098 355546 691334
rect 355782 691098 392426 691334
rect 392662 691098 392746 691334
rect 392982 691098 429626 691334
rect 429862 691098 429946 691334
rect 430182 691098 466826 691334
rect 467062 691098 467146 691334
rect 467382 691098 504026 691334
rect 504262 691098 504346 691334
rect 504582 691098 541226 691334
rect 541462 691098 541546 691334
rect 541782 691098 578426 691334
rect 578662 691098 578746 691334
rect 578982 691098 582820 691334
rect 1104 691066 582820 691098
rect 1104 687934 582820 687966
rect 1104 687698 16706 687934
rect 16942 687698 17026 687934
rect 17262 687698 53906 687934
rect 54142 687698 54226 687934
rect 54462 687698 91106 687934
rect 91342 687698 91426 687934
rect 91662 687698 128306 687934
rect 128542 687698 128626 687934
rect 128862 687698 165506 687934
rect 165742 687698 165826 687934
rect 166062 687698 202706 687934
rect 202942 687698 203026 687934
rect 203262 687698 239906 687934
rect 240142 687698 240226 687934
rect 240462 687698 277106 687934
rect 277342 687698 277426 687934
rect 277662 687698 314306 687934
rect 314542 687698 314626 687934
rect 314862 687698 351506 687934
rect 351742 687698 351826 687934
rect 352062 687698 388706 687934
rect 388942 687698 389026 687934
rect 389262 687698 425906 687934
rect 426142 687698 426226 687934
rect 426462 687698 463106 687934
rect 463342 687698 463426 687934
rect 463662 687698 500306 687934
rect 500542 687698 500626 687934
rect 500862 687698 537506 687934
rect 537742 687698 537826 687934
rect 538062 687698 574706 687934
rect 574942 687698 575026 687934
rect 575262 687698 582820 687934
rect 1104 687614 582820 687698
rect 1104 687378 16706 687614
rect 16942 687378 17026 687614
rect 17262 687378 53906 687614
rect 54142 687378 54226 687614
rect 54462 687378 91106 687614
rect 91342 687378 91426 687614
rect 91662 687378 128306 687614
rect 128542 687378 128626 687614
rect 128862 687378 165506 687614
rect 165742 687378 165826 687614
rect 166062 687378 202706 687614
rect 202942 687378 203026 687614
rect 203262 687378 239906 687614
rect 240142 687378 240226 687614
rect 240462 687378 277106 687614
rect 277342 687378 277426 687614
rect 277662 687378 314306 687614
rect 314542 687378 314626 687614
rect 314862 687378 351506 687614
rect 351742 687378 351826 687614
rect 352062 687378 388706 687614
rect 388942 687378 389026 687614
rect 389262 687378 425906 687614
rect 426142 687378 426226 687614
rect 426462 687378 463106 687614
rect 463342 687378 463426 687614
rect 463662 687378 500306 687614
rect 500542 687378 500626 687614
rect 500862 687378 537506 687614
rect 537742 687378 537826 687614
rect 538062 687378 574706 687614
rect 574942 687378 575026 687614
rect 575262 687378 582820 687614
rect 1104 687346 582820 687378
rect 1104 684214 582820 684246
rect 1104 683978 12986 684214
rect 13222 683978 13306 684214
rect 13542 683978 50186 684214
rect 50422 683978 50506 684214
rect 50742 683978 87386 684214
rect 87622 683978 87706 684214
rect 87942 683978 124586 684214
rect 124822 683978 124906 684214
rect 125142 683978 161786 684214
rect 162022 683978 162106 684214
rect 162342 683978 198986 684214
rect 199222 683978 199306 684214
rect 199542 683978 236186 684214
rect 236422 683978 236506 684214
rect 236742 683978 273386 684214
rect 273622 683978 273706 684214
rect 273942 683978 310586 684214
rect 310822 683978 310906 684214
rect 311142 683978 347786 684214
rect 348022 683978 348106 684214
rect 348342 683978 384986 684214
rect 385222 683978 385306 684214
rect 385542 683978 422186 684214
rect 422422 683978 422506 684214
rect 422742 683978 459386 684214
rect 459622 683978 459706 684214
rect 459942 683978 496586 684214
rect 496822 683978 496906 684214
rect 497142 683978 533786 684214
rect 534022 683978 534106 684214
rect 534342 683978 570986 684214
rect 571222 683978 571306 684214
rect 571542 683978 582820 684214
rect 1104 683894 582820 683978
rect 1104 683658 12986 683894
rect 13222 683658 13306 683894
rect 13542 683658 50186 683894
rect 50422 683658 50506 683894
rect 50742 683658 87386 683894
rect 87622 683658 87706 683894
rect 87942 683658 124586 683894
rect 124822 683658 124906 683894
rect 125142 683658 161786 683894
rect 162022 683658 162106 683894
rect 162342 683658 198986 683894
rect 199222 683658 199306 683894
rect 199542 683658 236186 683894
rect 236422 683658 236506 683894
rect 236742 683658 273386 683894
rect 273622 683658 273706 683894
rect 273942 683658 310586 683894
rect 310822 683658 310906 683894
rect 311142 683658 347786 683894
rect 348022 683658 348106 683894
rect 348342 683658 384986 683894
rect 385222 683658 385306 683894
rect 385542 683658 422186 683894
rect 422422 683658 422506 683894
rect 422742 683658 459386 683894
rect 459622 683658 459706 683894
rect 459942 683658 496586 683894
rect 496822 683658 496906 683894
rect 497142 683658 533786 683894
rect 534022 683658 534106 683894
rect 534342 683658 570986 683894
rect 571222 683658 571306 683894
rect 571542 683658 582820 683894
rect 1104 683626 582820 683658
rect 1104 680494 582820 680526
rect 1104 680258 9266 680494
rect 9502 680258 9586 680494
rect 9822 680258 46466 680494
rect 46702 680258 46786 680494
rect 47022 680258 83666 680494
rect 83902 680258 83986 680494
rect 84222 680258 120866 680494
rect 121102 680258 121186 680494
rect 121422 680258 158066 680494
rect 158302 680258 158386 680494
rect 158622 680258 195266 680494
rect 195502 680258 195586 680494
rect 195822 680258 232466 680494
rect 232702 680258 232786 680494
rect 233022 680258 269666 680494
rect 269902 680258 269986 680494
rect 270222 680258 306866 680494
rect 307102 680258 307186 680494
rect 307422 680258 344066 680494
rect 344302 680258 344386 680494
rect 344622 680258 381266 680494
rect 381502 680258 381586 680494
rect 381822 680258 418466 680494
rect 418702 680258 418786 680494
rect 419022 680258 455666 680494
rect 455902 680258 455986 680494
rect 456222 680258 492866 680494
rect 493102 680258 493186 680494
rect 493422 680258 530066 680494
rect 530302 680258 530386 680494
rect 530622 680258 567266 680494
rect 567502 680258 567586 680494
rect 567822 680258 582820 680494
rect 1104 680174 582820 680258
rect 1104 679938 9266 680174
rect 9502 679938 9586 680174
rect 9822 679938 46466 680174
rect 46702 679938 46786 680174
rect 47022 679938 83666 680174
rect 83902 679938 83986 680174
rect 84222 679938 120866 680174
rect 121102 679938 121186 680174
rect 121422 679938 158066 680174
rect 158302 679938 158386 680174
rect 158622 679938 195266 680174
rect 195502 679938 195586 680174
rect 195822 679938 232466 680174
rect 232702 679938 232786 680174
rect 233022 679938 269666 680174
rect 269902 679938 269986 680174
rect 270222 679938 306866 680174
rect 307102 679938 307186 680174
rect 307422 679938 344066 680174
rect 344302 679938 344386 680174
rect 344622 679938 381266 680174
rect 381502 679938 381586 680174
rect 381822 679938 418466 680174
rect 418702 679938 418786 680174
rect 419022 679938 455666 680174
rect 455902 679938 455986 680174
rect 456222 679938 492866 680174
rect 493102 679938 493186 680174
rect 493422 679938 530066 680174
rect 530302 679938 530386 680174
rect 530622 679938 567266 680174
rect 567502 679938 567586 680174
rect 567822 679938 582820 680174
rect 1104 679906 582820 679938
rect 1104 676774 582820 676806
rect 1104 676538 5546 676774
rect 5782 676538 5866 676774
rect 6102 676538 42746 676774
rect 42982 676538 43066 676774
rect 43302 676538 79946 676774
rect 80182 676538 80266 676774
rect 80502 676538 117146 676774
rect 117382 676538 117466 676774
rect 117702 676538 154346 676774
rect 154582 676538 154666 676774
rect 154902 676538 191546 676774
rect 191782 676538 191866 676774
rect 192102 676538 228746 676774
rect 228982 676538 229066 676774
rect 229302 676538 265946 676774
rect 266182 676538 266266 676774
rect 266502 676538 303146 676774
rect 303382 676538 303466 676774
rect 303702 676538 340346 676774
rect 340582 676538 340666 676774
rect 340902 676538 377546 676774
rect 377782 676538 377866 676774
rect 378102 676538 414746 676774
rect 414982 676538 415066 676774
rect 415302 676538 451946 676774
rect 452182 676538 452266 676774
rect 452502 676538 489146 676774
rect 489382 676538 489466 676774
rect 489702 676538 526346 676774
rect 526582 676538 526666 676774
rect 526902 676538 563546 676774
rect 563782 676538 563866 676774
rect 564102 676538 582820 676774
rect 1104 676454 582820 676538
rect 1104 676218 5546 676454
rect 5782 676218 5866 676454
rect 6102 676218 42746 676454
rect 42982 676218 43066 676454
rect 43302 676218 79946 676454
rect 80182 676218 80266 676454
rect 80502 676218 117146 676454
rect 117382 676218 117466 676454
rect 117702 676218 154346 676454
rect 154582 676218 154666 676454
rect 154902 676218 191546 676454
rect 191782 676218 191866 676454
rect 192102 676218 228746 676454
rect 228982 676218 229066 676454
rect 229302 676218 265946 676454
rect 266182 676218 266266 676454
rect 266502 676218 303146 676454
rect 303382 676218 303466 676454
rect 303702 676218 340346 676454
rect 340582 676218 340666 676454
rect 340902 676218 377546 676454
rect 377782 676218 377866 676454
rect 378102 676218 414746 676454
rect 414982 676218 415066 676454
rect 415302 676218 451946 676454
rect 452182 676218 452266 676454
rect 452502 676218 489146 676454
rect 489382 676218 489466 676454
rect 489702 676218 526346 676454
rect 526582 676218 526666 676454
rect 526902 676218 563546 676454
rect 563782 676218 563866 676454
rect 564102 676218 582820 676454
rect 1104 676186 582820 676218
rect 1104 673054 582820 673086
rect 1104 672818 1826 673054
rect 2062 672818 2146 673054
rect 2382 672818 39026 673054
rect 39262 672818 39346 673054
rect 39582 672818 76226 673054
rect 76462 672818 76546 673054
rect 76782 672818 113426 673054
rect 113662 672818 113746 673054
rect 113982 672818 150626 673054
rect 150862 672818 150946 673054
rect 151182 672818 187826 673054
rect 188062 672818 188146 673054
rect 188382 672818 225026 673054
rect 225262 672818 225346 673054
rect 225582 672818 262226 673054
rect 262462 672818 262546 673054
rect 262782 672818 299426 673054
rect 299662 672818 299746 673054
rect 299982 672818 336626 673054
rect 336862 672818 336946 673054
rect 337182 672818 373826 673054
rect 374062 672818 374146 673054
rect 374382 672818 411026 673054
rect 411262 672818 411346 673054
rect 411582 672818 448226 673054
rect 448462 672818 448546 673054
rect 448782 672818 485426 673054
rect 485662 672818 485746 673054
rect 485982 672818 522626 673054
rect 522862 672818 522946 673054
rect 523182 672818 559826 673054
rect 560062 672818 560146 673054
rect 560382 672818 582820 673054
rect 1104 672734 582820 672818
rect 1104 672498 1826 672734
rect 2062 672498 2146 672734
rect 2382 672498 39026 672734
rect 39262 672498 39346 672734
rect 39582 672498 76226 672734
rect 76462 672498 76546 672734
rect 76782 672498 113426 672734
rect 113662 672498 113746 672734
rect 113982 672498 150626 672734
rect 150862 672498 150946 672734
rect 151182 672498 187826 672734
rect 188062 672498 188146 672734
rect 188382 672498 225026 672734
rect 225262 672498 225346 672734
rect 225582 672498 262226 672734
rect 262462 672498 262546 672734
rect 262782 672498 299426 672734
rect 299662 672498 299746 672734
rect 299982 672498 336626 672734
rect 336862 672498 336946 672734
rect 337182 672498 373826 672734
rect 374062 672498 374146 672734
rect 374382 672498 411026 672734
rect 411262 672498 411346 672734
rect 411582 672498 448226 672734
rect 448462 672498 448546 672734
rect 448782 672498 485426 672734
rect 485662 672498 485746 672734
rect 485982 672498 522626 672734
rect 522862 672498 522946 672734
rect 523182 672498 559826 672734
rect 560062 672498 560146 672734
rect 560382 672498 582820 672734
rect 1104 672466 582820 672498
rect 1104 661894 582820 661926
rect 1104 661658 27866 661894
rect 28102 661658 28186 661894
rect 28422 661658 65066 661894
rect 65302 661658 65386 661894
rect 65622 661658 102266 661894
rect 102502 661658 102586 661894
rect 102822 661658 139466 661894
rect 139702 661658 139786 661894
rect 140022 661658 176666 661894
rect 176902 661658 176986 661894
rect 177222 661658 213866 661894
rect 214102 661658 214186 661894
rect 214422 661658 251066 661894
rect 251302 661658 251386 661894
rect 251622 661658 288266 661894
rect 288502 661658 288586 661894
rect 288822 661658 325466 661894
rect 325702 661658 325786 661894
rect 326022 661658 362666 661894
rect 362902 661658 362986 661894
rect 363222 661658 399866 661894
rect 400102 661658 400186 661894
rect 400422 661658 437066 661894
rect 437302 661658 437386 661894
rect 437622 661658 474266 661894
rect 474502 661658 474586 661894
rect 474822 661658 511466 661894
rect 511702 661658 511786 661894
rect 512022 661658 548666 661894
rect 548902 661658 548986 661894
rect 549222 661658 582820 661894
rect 1104 661574 582820 661658
rect 1104 661338 27866 661574
rect 28102 661338 28186 661574
rect 28422 661338 65066 661574
rect 65302 661338 65386 661574
rect 65622 661338 102266 661574
rect 102502 661338 102586 661574
rect 102822 661338 139466 661574
rect 139702 661338 139786 661574
rect 140022 661338 176666 661574
rect 176902 661338 176986 661574
rect 177222 661338 213866 661574
rect 214102 661338 214186 661574
rect 214422 661338 251066 661574
rect 251302 661338 251386 661574
rect 251622 661338 288266 661574
rect 288502 661338 288586 661574
rect 288822 661338 325466 661574
rect 325702 661338 325786 661574
rect 326022 661338 362666 661574
rect 362902 661338 362986 661574
rect 363222 661338 399866 661574
rect 400102 661338 400186 661574
rect 400422 661338 437066 661574
rect 437302 661338 437386 661574
rect 437622 661338 474266 661574
rect 474502 661338 474586 661574
rect 474822 661338 511466 661574
rect 511702 661338 511786 661574
rect 512022 661338 548666 661574
rect 548902 661338 548986 661574
rect 549222 661338 582820 661574
rect 1104 661306 582820 661338
rect 1104 658174 582820 658206
rect 1104 657938 24146 658174
rect 24382 657938 24466 658174
rect 24702 657938 61346 658174
rect 61582 657938 61666 658174
rect 61902 657938 98546 658174
rect 98782 657938 98866 658174
rect 99102 657938 135746 658174
rect 135982 657938 136066 658174
rect 136302 657938 172946 658174
rect 173182 657938 173266 658174
rect 173502 657938 210146 658174
rect 210382 657938 210466 658174
rect 210702 657938 247346 658174
rect 247582 657938 247666 658174
rect 247902 657938 284546 658174
rect 284782 657938 284866 658174
rect 285102 657938 321746 658174
rect 321982 657938 322066 658174
rect 322302 657938 358946 658174
rect 359182 657938 359266 658174
rect 359502 657938 396146 658174
rect 396382 657938 396466 658174
rect 396702 657938 433346 658174
rect 433582 657938 433666 658174
rect 433902 657938 470546 658174
rect 470782 657938 470866 658174
rect 471102 657938 507746 658174
rect 507982 657938 508066 658174
rect 508302 657938 544946 658174
rect 545182 657938 545266 658174
rect 545502 657938 582146 658174
rect 582382 657938 582466 658174
rect 582702 657938 582820 658174
rect 1104 657854 582820 657938
rect 1104 657618 24146 657854
rect 24382 657618 24466 657854
rect 24702 657618 61346 657854
rect 61582 657618 61666 657854
rect 61902 657618 98546 657854
rect 98782 657618 98866 657854
rect 99102 657618 135746 657854
rect 135982 657618 136066 657854
rect 136302 657618 172946 657854
rect 173182 657618 173266 657854
rect 173502 657618 210146 657854
rect 210382 657618 210466 657854
rect 210702 657618 247346 657854
rect 247582 657618 247666 657854
rect 247902 657618 284546 657854
rect 284782 657618 284866 657854
rect 285102 657618 321746 657854
rect 321982 657618 322066 657854
rect 322302 657618 358946 657854
rect 359182 657618 359266 657854
rect 359502 657618 396146 657854
rect 396382 657618 396466 657854
rect 396702 657618 433346 657854
rect 433582 657618 433666 657854
rect 433902 657618 470546 657854
rect 470782 657618 470866 657854
rect 471102 657618 507746 657854
rect 507982 657618 508066 657854
rect 508302 657618 544946 657854
rect 545182 657618 545266 657854
rect 545502 657618 582146 657854
rect 582382 657618 582466 657854
rect 582702 657618 582820 657854
rect 1104 657586 582820 657618
rect 1104 654454 582820 654486
rect 1104 654218 20426 654454
rect 20662 654218 20746 654454
rect 20982 654218 57626 654454
rect 57862 654218 57946 654454
rect 58182 654218 94826 654454
rect 95062 654218 95146 654454
rect 95382 654218 132026 654454
rect 132262 654218 132346 654454
rect 132582 654218 169226 654454
rect 169462 654218 169546 654454
rect 169782 654218 206426 654454
rect 206662 654218 206746 654454
rect 206982 654218 243626 654454
rect 243862 654218 243946 654454
rect 244182 654218 280826 654454
rect 281062 654218 281146 654454
rect 281382 654218 318026 654454
rect 318262 654218 318346 654454
rect 318582 654218 355226 654454
rect 355462 654218 355546 654454
rect 355782 654218 392426 654454
rect 392662 654218 392746 654454
rect 392982 654218 429626 654454
rect 429862 654218 429946 654454
rect 430182 654218 466826 654454
rect 467062 654218 467146 654454
rect 467382 654218 504026 654454
rect 504262 654218 504346 654454
rect 504582 654218 541226 654454
rect 541462 654218 541546 654454
rect 541782 654218 578426 654454
rect 578662 654218 578746 654454
rect 578982 654218 582820 654454
rect 1104 654134 582820 654218
rect 1104 653898 20426 654134
rect 20662 653898 20746 654134
rect 20982 653898 57626 654134
rect 57862 653898 57946 654134
rect 58182 653898 94826 654134
rect 95062 653898 95146 654134
rect 95382 653898 132026 654134
rect 132262 653898 132346 654134
rect 132582 653898 169226 654134
rect 169462 653898 169546 654134
rect 169782 653898 206426 654134
rect 206662 653898 206746 654134
rect 206982 653898 243626 654134
rect 243862 653898 243946 654134
rect 244182 653898 280826 654134
rect 281062 653898 281146 654134
rect 281382 653898 318026 654134
rect 318262 653898 318346 654134
rect 318582 653898 355226 654134
rect 355462 653898 355546 654134
rect 355782 653898 392426 654134
rect 392662 653898 392746 654134
rect 392982 653898 429626 654134
rect 429862 653898 429946 654134
rect 430182 653898 466826 654134
rect 467062 653898 467146 654134
rect 467382 653898 504026 654134
rect 504262 653898 504346 654134
rect 504582 653898 541226 654134
rect 541462 653898 541546 654134
rect 541782 653898 578426 654134
rect 578662 653898 578746 654134
rect 578982 653898 582820 654134
rect 1104 653866 582820 653898
rect 1104 650734 582820 650766
rect 1104 650498 16706 650734
rect 16942 650498 17026 650734
rect 17262 650498 53906 650734
rect 54142 650498 54226 650734
rect 54462 650498 91106 650734
rect 91342 650498 91426 650734
rect 91662 650498 128306 650734
rect 128542 650498 128626 650734
rect 128862 650498 165506 650734
rect 165742 650498 165826 650734
rect 166062 650498 202706 650734
rect 202942 650498 203026 650734
rect 203262 650498 239906 650734
rect 240142 650498 240226 650734
rect 240462 650498 277106 650734
rect 277342 650498 277426 650734
rect 277662 650498 314306 650734
rect 314542 650498 314626 650734
rect 314862 650498 351506 650734
rect 351742 650498 351826 650734
rect 352062 650498 388706 650734
rect 388942 650498 389026 650734
rect 389262 650498 425906 650734
rect 426142 650498 426226 650734
rect 426462 650498 463106 650734
rect 463342 650498 463426 650734
rect 463662 650498 500306 650734
rect 500542 650498 500626 650734
rect 500862 650498 537506 650734
rect 537742 650498 537826 650734
rect 538062 650498 574706 650734
rect 574942 650498 575026 650734
rect 575262 650498 582820 650734
rect 1104 650414 582820 650498
rect 1104 650178 16706 650414
rect 16942 650178 17026 650414
rect 17262 650178 53906 650414
rect 54142 650178 54226 650414
rect 54462 650178 91106 650414
rect 91342 650178 91426 650414
rect 91662 650178 128306 650414
rect 128542 650178 128626 650414
rect 128862 650178 165506 650414
rect 165742 650178 165826 650414
rect 166062 650178 202706 650414
rect 202942 650178 203026 650414
rect 203262 650178 239906 650414
rect 240142 650178 240226 650414
rect 240462 650178 277106 650414
rect 277342 650178 277426 650414
rect 277662 650178 314306 650414
rect 314542 650178 314626 650414
rect 314862 650178 351506 650414
rect 351742 650178 351826 650414
rect 352062 650178 388706 650414
rect 388942 650178 389026 650414
rect 389262 650178 425906 650414
rect 426142 650178 426226 650414
rect 426462 650178 463106 650414
rect 463342 650178 463426 650414
rect 463662 650178 500306 650414
rect 500542 650178 500626 650414
rect 500862 650178 537506 650414
rect 537742 650178 537826 650414
rect 538062 650178 574706 650414
rect 574942 650178 575026 650414
rect 575262 650178 582820 650414
rect 1104 650146 582820 650178
rect 1104 647014 582820 647046
rect 1104 646778 12986 647014
rect 13222 646778 13306 647014
rect 13542 646778 50186 647014
rect 50422 646778 50506 647014
rect 50742 646778 87386 647014
rect 87622 646778 87706 647014
rect 87942 646778 124586 647014
rect 124822 646778 124906 647014
rect 125142 646778 161786 647014
rect 162022 646778 162106 647014
rect 162342 646778 198986 647014
rect 199222 646778 199306 647014
rect 199542 646778 236186 647014
rect 236422 646778 236506 647014
rect 236742 646778 273386 647014
rect 273622 646778 273706 647014
rect 273942 646778 310586 647014
rect 310822 646778 310906 647014
rect 311142 646778 347786 647014
rect 348022 646778 348106 647014
rect 348342 646778 384986 647014
rect 385222 646778 385306 647014
rect 385542 646778 422186 647014
rect 422422 646778 422506 647014
rect 422742 646778 459386 647014
rect 459622 646778 459706 647014
rect 459942 646778 496586 647014
rect 496822 646778 496906 647014
rect 497142 646778 533786 647014
rect 534022 646778 534106 647014
rect 534342 646778 570986 647014
rect 571222 646778 571306 647014
rect 571542 646778 582820 647014
rect 1104 646694 582820 646778
rect 1104 646458 12986 646694
rect 13222 646458 13306 646694
rect 13542 646458 50186 646694
rect 50422 646458 50506 646694
rect 50742 646458 87386 646694
rect 87622 646458 87706 646694
rect 87942 646458 124586 646694
rect 124822 646458 124906 646694
rect 125142 646458 161786 646694
rect 162022 646458 162106 646694
rect 162342 646458 198986 646694
rect 199222 646458 199306 646694
rect 199542 646458 236186 646694
rect 236422 646458 236506 646694
rect 236742 646458 273386 646694
rect 273622 646458 273706 646694
rect 273942 646458 310586 646694
rect 310822 646458 310906 646694
rect 311142 646458 347786 646694
rect 348022 646458 348106 646694
rect 348342 646458 384986 646694
rect 385222 646458 385306 646694
rect 385542 646458 422186 646694
rect 422422 646458 422506 646694
rect 422742 646458 459386 646694
rect 459622 646458 459706 646694
rect 459942 646458 496586 646694
rect 496822 646458 496906 646694
rect 497142 646458 533786 646694
rect 534022 646458 534106 646694
rect 534342 646458 570986 646694
rect 571222 646458 571306 646694
rect 571542 646458 582820 646694
rect 1104 646426 582820 646458
rect 1104 643294 582820 643326
rect 1104 643058 9266 643294
rect 9502 643058 9586 643294
rect 9822 643058 46466 643294
rect 46702 643058 46786 643294
rect 47022 643058 83666 643294
rect 83902 643058 83986 643294
rect 84222 643058 120866 643294
rect 121102 643058 121186 643294
rect 121422 643058 158066 643294
rect 158302 643058 158386 643294
rect 158622 643058 195266 643294
rect 195502 643058 195586 643294
rect 195822 643058 232466 643294
rect 232702 643058 232786 643294
rect 233022 643058 269666 643294
rect 269902 643058 269986 643294
rect 270222 643058 306866 643294
rect 307102 643058 307186 643294
rect 307422 643058 344066 643294
rect 344302 643058 344386 643294
rect 344622 643058 381266 643294
rect 381502 643058 381586 643294
rect 381822 643058 418466 643294
rect 418702 643058 418786 643294
rect 419022 643058 455666 643294
rect 455902 643058 455986 643294
rect 456222 643058 492866 643294
rect 493102 643058 493186 643294
rect 493422 643058 530066 643294
rect 530302 643058 530386 643294
rect 530622 643058 567266 643294
rect 567502 643058 567586 643294
rect 567822 643058 582820 643294
rect 1104 642974 582820 643058
rect 1104 642738 9266 642974
rect 9502 642738 9586 642974
rect 9822 642738 46466 642974
rect 46702 642738 46786 642974
rect 47022 642738 83666 642974
rect 83902 642738 83986 642974
rect 84222 642738 120866 642974
rect 121102 642738 121186 642974
rect 121422 642738 158066 642974
rect 158302 642738 158386 642974
rect 158622 642738 195266 642974
rect 195502 642738 195586 642974
rect 195822 642738 232466 642974
rect 232702 642738 232786 642974
rect 233022 642738 269666 642974
rect 269902 642738 269986 642974
rect 270222 642738 306866 642974
rect 307102 642738 307186 642974
rect 307422 642738 344066 642974
rect 344302 642738 344386 642974
rect 344622 642738 381266 642974
rect 381502 642738 381586 642974
rect 381822 642738 418466 642974
rect 418702 642738 418786 642974
rect 419022 642738 455666 642974
rect 455902 642738 455986 642974
rect 456222 642738 492866 642974
rect 493102 642738 493186 642974
rect 493422 642738 530066 642974
rect 530302 642738 530386 642974
rect 530622 642738 567266 642974
rect 567502 642738 567586 642974
rect 567822 642738 582820 642974
rect 1104 642706 582820 642738
rect 1104 639574 582820 639606
rect 1104 639338 5546 639574
rect 5782 639338 5866 639574
rect 6102 639338 42746 639574
rect 42982 639338 43066 639574
rect 43302 639338 79946 639574
rect 80182 639338 80266 639574
rect 80502 639338 117146 639574
rect 117382 639338 117466 639574
rect 117702 639338 154346 639574
rect 154582 639338 154666 639574
rect 154902 639338 191546 639574
rect 191782 639338 191866 639574
rect 192102 639338 228746 639574
rect 228982 639338 229066 639574
rect 229302 639338 265946 639574
rect 266182 639338 266266 639574
rect 266502 639338 303146 639574
rect 303382 639338 303466 639574
rect 303702 639338 340346 639574
rect 340582 639338 340666 639574
rect 340902 639338 377546 639574
rect 377782 639338 377866 639574
rect 378102 639338 414746 639574
rect 414982 639338 415066 639574
rect 415302 639338 451946 639574
rect 452182 639338 452266 639574
rect 452502 639338 489146 639574
rect 489382 639338 489466 639574
rect 489702 639338 526346 639574
rect 526582 639338 526666 639574
rect 526902 639338 563546 639574
rect 563782 639338 563866 639574
rect 564102 639338 582820 639574
rect 1104 639254 582820 639338
rect 1104 639018 5546 639254
rect 5782 639018 5866 639254
rect 6102 639018 42746 639254
rect 42982 639018 43066 639254
rect 43302 639018 79946 639254
rect 80182 639018 80266 639254
rect 80502 639018 117146 639254
rect 117382 639018 117466 639254
rect 117702 639018 154346 639254
rect 154582 639018 154666 639254
rect 154902 639018 191546 639254
rect 191782 639018 191866 639254
rect 192102 639018 228746 639254
rect 228982 639018 229066 639254
rect 229302 639018 265946 639254
rect 266182 639018 266266 639254
rect 266502 639018 303146 639254
rect 303382 639018 303466 639254
rect 303702 639018 340346 639254
rect 340582 639018 340666 639254
rect 340902 639018 377546 639254
rect 377782 639018 377866 639254
rect 378102 639018 414746 639254
rect 414982 639018 415066 639254
rect 415302 639018 451946 639254
rect 452182 639018 452266 639254
rect 452502 639018 489146 639254
rect 489382 639018 489466 639254
rect 489702 639018 526346 639254
rect 526582 639018 526666 639254
rect 526902 639018 563546 639254
rect 563782 639018 563866 639254
rect 564102 639018 582820 639254
rect 1104 638986 582820 639018
rect 1104 635854 582820 635886
rect 1104 635618 1826 635854
rect 2062 635618 2146 635854
rect 2382 635618 39026 635854
rect 39262 635618 39346 635854
rect 39582 635618 76226 635854
rect 76462 635618 76546 635854
rect 76782 635618 113426 635854
rect 113662 635618 113746 635854
rect 113982 635618 150626 635854
rect 150862 635618 150946 635854
rect 151182 635618 187826 635854
rect 188062 635618 188146 635854
rect 188382 635618 225026 635854
rect 225262 635618 225346 635854
rect 225582 635618 262226 635854
rect 262462 635618 262546 635854
rect 262782 635618 299426 635854
rect 299662 635618 299746 635854
rect 299982 635618 336626 635854
rect 336862 635618 336946 635854
rect 337182 635618 373826 635854
rect 374062 635618 374146 635854
rect 374382 635618 411026 635854
rect 411262 635618 411346 635854
rect 411582 635618 448226 635854
rect 448462 635618 448546 635854
rect 448782 635618 485426 635854
rect 485662 635618 485746 635854
rect 485982 635618 522626 635854
rect 522862 635618 522946 635854
rect 523182 635618 559826 635854
rect 560062 635618 560146 635854
rect 560382 635618 582820 635854
rect 1104 635534 582820 635618
rect 1104 635298 1826 635534
rect 2062 635298 2146 635534
rect 2382 635298 39026 635534
rect 39262 635298 39346 635534
rect 39582 635298 76226 635534
rect 76462 635298 76546 635534
rect 76782 635298 113426 635534
rect 113662 635298 113746 635534
rect 113982 635298 150626 635534
rect 150862 635298 150946 635534
rect 151182 635298 187826 635534
rect 188062 635298 188146 635534
rect 188382 635298 225026 635534
rect 225262 635298 225346 635534
rect 225582 635298 262226 635534
rect 262462 635298 262546 635534
rect 262782 635298 299426 635534
rect 299662 635298 299746 635534
rect 299982 635298 336626 635534
rect 336862 635298 336946 635534
rect 337182 635298 373826 635534
rect 374062 635298 374146 635534
rect 374382 635298 411026 635534
rect 411262 635298 411346 635534
rect 411582 635298 448226 635534
rect 448462 635298 448546 635534
rect 448782 635298 485426 635534
rect 485662 635298 485746 635534
rect 485982 635298 522626 635534
rect 522862 635298 522946 635534
rect 523182 635298 559826 635534
rect 560062 635298 560146 635534
rect 560382 635298 582820 635534
rect 1104 635266 582820 635298
rect 1104 624694 582820 624726
rect 1104 624458 27866 624694
rect 28102 624458 28186 624694
rect 28422 624458 65066 624694
rect 65302 624458 65386 624694
rect 65622 624458 102266 624694
rect 102502 624458 102586 624694
rect 102822 624458 139466 624694
rect 139702 624458 139786 624694
rect 140022 624458 176666 624694
rect 176902 624458 176986 624694
rect 177222 624458 213866 624694
rect 214102 624458 214186 624694
rect 214422 624458 251066 624694
rect 251302 624458 251386 624694
rect 251622 624458 288266 624694
rect 288502 624458 288586 624694
rect 288822 624458 325466 624694
rect 325702 624458 325786 624694
rect 326022 624458 362666 624694
rect 362902 624458 362986 624694
rect 363222 624458 399866 624694
rect 400102 624458 400186 624694
rect 400422 624458 437066 624694
rect 437302 624458 437386 624694
rect 437622 624458 474266 624694
rect 474502 624458 474586 624694
rect 474822 624458 511466 624694
rect 511702 624458 511786 624694
rect 512022 624458 548666 624694
rect 548902 624458 548986 624694
rect 549222 624458 582820 624694
rect 1104 624374 582820 624458
rect 1104 624138 27866 624374
rect 28102 624138 28186 624374
rect 28422 624138 65066 624374
rect 65302 624138 65386 624374
rect 65622 624138 102266 624374
rect 102502 624138 102586 624374
rect 102822 624138 139466 624374
rect 139702 624138 139786 624374
rect 140022 624138 176666 624374
rect 176902 624138 176986 624374
rect 177222 624138 213866 624374
rect 214102 624138 214186 624374
rect 214422 624138 251066 624374
rect 251302 624138 251386 624374
rect 251622 624138 288266 624374
rect 288502 624138 288586 624374
rect 288822 624138 325466 624374
rect 325702 624138 325786 624374
rect 326022 624138 362666 624374
rect 362902 624138 362986 624374
rect 363222 624138 399866 624374
rect 400102 624138 400186 624374
rect 400422 624138 437066 624374
rect 437302 624138 437386 624374
rect 437622 624138 474266 624374
rect 474502 624138 474586 624374
rect 474822 624138 511466 624374
rect 511702 624138 511786 624374
rect 512022 624138 548666 624374
rect 548902 624138 548986 624374
rect 549222 624138 582820 624374
rect 1104 624106 582820 624138
rect 1104 620974 582820 621006
rect 1104 620738 24146 620974
rect 24382 620738 24466 620974
rect 24702 620738 61346 620974
rect 61582 620738 61666 620974
rect 61902 620738 98546 620974
rect 98782 620738 98866 620974
rect 99102 620738 135746 620974
rect 135982 620738 136066 620974
rect 136302 620738 172946 620974
rect 173182 620738 173266 620974
rect 173502 620738 210146 620974
rect 210382 620738 210466 620974
rect 210702 620738 247346 620974
rect 247582 620738 247666 620974
rect 247902 620738 284546 620974
rect 284782 620738 284866 620974
rect 285102 620738 321746 620974
rect 321982 620738 322066 620974
rect 322302 620738 358946 620974
rect 359182 620738 359266 620974
rect 359502 620738 396146 620974
rect 396382 620738 396466 620974
rect 396702 620738 433346 620974
rect 433582 620738 433666 620974
rect 433902 620738 470546 620974
rect 470782 620738 470866 620974
rect 471102 620738 507746 620974
rect 507982 620738 508066 620974
rect 508302 620738 544946 620974
rect 545182 620738 545266 620974
rect 545502 620738 582146 620974
rect 582382 620738 582466 620974
rect 582702 620738 582820 620974
rect 1104 620654 582820 620738
rect 1104 620418 24146 620654
rect 24382 620418 24466 620654
rect 24702 620418 61346 620654
rect 61582 620418 61666 620654
rect 61902 620418 98546 620654
rect 98782 620418 98866 620654
rect 99102 620418 135746 620654
rect 135982 620418 136066 620654
rect 136302 620418 172946 620654
rect 173182 620418 173266 620654
rect 173502 620418 210146 620654
rect 210382 620418 210466 620654
rect 210702 620418 247346 620654
rect 247582 620418 247666 620654
rect 247902 620418 284546 620654
rect 284782 620418 284866 620654
rect 285102 620418 321746 620654
rect 321982 620418 322066 620654
rect 322302 620418 358946 620654
rect 359182 620418 359266 620654
rect 359502 620418 396146 620654
rect 396382 620418 396466 620654
rect 396702 620418 433346 620654
rect 433582 620418 433666 620654
rect 433902 620418 470546 620654
rect 470782 620418 470866 620654
rect 471102 620418 507746 620654
rect 507982 620418 508066 620654
rect 508302 620418 544946 620654
rect 545182 620418 545266 620654
rect 545502 620418 582146 620654
rect 582382 620418 582466 620654
rect 582702 620418 582820 620654
rect 1104 620386 582820 620418
rect 1104 617254 582820 617286
rect 1104 617018 20426 617254
rect 20662 617018 20746 617254
rect 20982 617018 57626 617254
rect 57862 617018 57946 617254
rect 58182 617018 94826 617254
rect 95062 617018 95146 617254
rect 95382 617018 132026 617254
rect 132262 617018 132346 617254
rect 132582 617018 169226 617254
rect 169462 617018 169546 617254
rect 169782 617018 206426 617254
rect 206662 617018 206746 617254
rect 206982 617018 243626 617254
rect 243862 617018 243946 617254
rect 244182 617018 280826 617254
rect 281062 617018 281146 617254
rect 281382 617018 318026 617254
rect 318262 617018 318346 617254
rect 318582 617018 355226 617254
rect 355462 617018 355546 617254
rect 355782 617018 392426 617254
rect 392662 617018 392746 617254
rect 392982 617018 429626 617254
rect 429862 617018 429946 617254
rect 430182 617018 466826 617254
rect 467062 617018 467146 617254
rect 467382 617018 504026 617254
rect 504262 617018 504346 617254
rect 504582 617018 541226 617254
rect 541462 617018 541546 617254
rect 541782 617018 578426 617254
rect 578662 617018 578746 617254
rect 578982 617018 582820 617254
rect 1104 616934 582820 617018
rect 1104 616698 20426 616934
rect 20662 616698 20746 616934
rect 20982 616698 57626 616934
rect 57862 616698 57946 616934
rect 58182 616698 94826 616934
rect 95062 616698 95146 616934
rect 95382 616698 132026 616934
rect 132262 616698 132346 616934
rect 132582 616698 169226 616934
rect 169462 616698 169546 616934
rect 169782 616698 206426 616934
rect 206662 616698 206746 616934
rect 206982 616698 243626 616934
rect 243862 616698 243946 616934
rect 244182 616698 280826 616934
rect 281062 616698 281146 616934
rect 281382 616698 318026 616934
rect 318262 616698 318346 616934
rect 318582 616698 355226 616934
rect 355462 616698 355546 616934
rect 355782 616698 392426 616934
rect 392662 616698 392746 616934
rect 392982 616698 429626 616934
rect 429862 616698 429946 616934
rect 430182 616698 466826 616934
rect 467062 616698 467146 616934
rect 467382 616698 504026 616934
rect 504262 616698 504346 616934
rect 504582 616698 541226 616934
rect 541462 616698 541546 616934
rect 541782 616698 578426 616934
rect 578662 616698 578746 616934
rect 578982 616698 582820 616934
rect 1104 616666 582820 616698
rect 1104 613534 582820 613566
rect 1104 613298 16706 613534
rect 16942 613298 17026 613534
rect 17262 613298 53906 613534
rect 54142 613298 54226 613534
rect 54462 613298 91106 613534
rect 91342 613298 91426 613534
rect 91662 613298 128306 613534
rect 128542 613298 128626 613534
rect 128862 613298 165506 613534
rect 165742 613298 165826 613534
rect 166062 613298 202706 613534
rect 202942 613298 203026 613534
rect 203262 613298 239906 613534
rect 240142 613298 240226 613534
rect 240462 613298 277106 613534
rect 277342 613298 277426 613534
rect 277662 613298 314306 613534
rect 314542 613298 314626 613534
rect 314862 613298 351506 613534
rect 351742 613298 351826 613534
rect 352062 613298 388706 613534
rect 388942 613298 389026 613534
rect 389262 613298 425906 613534
rect 426142 613298 426226 613534
rect 426462 613298 463106 613534
rect 463342 613298 463426 613534
rect 463662 613298 500306 613534
rect 500542 613298 500626 613534
rect 500862 613298 537506 613534
rect 537742 613298 537826 613534
rect 538062 613298 574706 613534
rect 574942 613298 575026 613534
rect 575262 613298 582820 613534
rect 1104 613214 582820 613298
rect 1104 612978 16706 613214
rect 16942 612978 17026 613214
rect 17262 612978 53906 613214
rect 54142 612978 54226 613214
rect 54462 612978 91106 613214
rect 91342 612978 91426 613214
rect 91662 612978 128306 613214
rect 128542 612978 128626 613214
rect 128862 612978 165506 613214
rect 165742 612978 165826 613214
rect 166062 612978 202706 613214
rect 202942 612978 203026 613214
rect 203262 612978 239906 613214
rect 240142 612978 240226 613214
rect 240462 612978 277106 613214
rect 277342 612978 277426 613214
rect 277662 612978 314306 613214
rect 314542 612978 314626 613214
rect 314862 612978 351506 613214
rect 351742 612978 351826 613214
rect 352062 612978 388706 613214
rect 388942 612978 389026 613214
rect 389262 612978 425906 613214
rect 426142 612978 426226 613214
rect 426462 612978 463106 613214
rect 463342 612978 463426 613214
rect 463662 612978 500306 613214
rect 500542 612978 500626 613214
rect 500862 612978 537506 613214
rect 537742 612978 537826 613214
rect 538062 612978 574706 613214
rect 574942 612978 575026 613214
rect 575262 612978 582820 613214
rect 1104 612946 582820 612978
rect 1104 609814 582820 609846
rect 1104 609578 12986 609814
rect 13222 609578 13306 609814
rect 13542 609578 50186 609814
rect 50422 609578 50506 609814
rect 50742 609578 87386 609814
rect 87622 609578 87706 609814
rect 87942 609578 124586 609814
rect 124822 609578 124906 609814
rect 125142 609578 161786 609814
rect 162022 609578 162106 609814
rect 162342 609578 198986 609814
rect 199222 609578 199306 609814
rect 199542 609578 236186 609814
rect 236422 609578 236506 609814
rect 236742 609578 273386 609814
rect 273622 609578 273706 609814
rect 273942 609578 310586 609814
rect 310822 609578 310906 609814
rect 311142 609578 347786 609814
rect 348022 609578 348106 609814
rect 348342 609578 384986 609814
rect 385222 609578 385306 609814
rect 385542 609578 422186 609814
rect 422422 609578 422506 609814
rect 422742 609578 459386 609814
rect 459622 609578 459706 609814
rect 459942 609578 496586 609814
rect 496822 609578 496906 609814
rect 497142 609578 533786 609814
rect 534022 609578 534106 609814
rect 534342 609578 570986 609814
rect 571222 609578 571306 609814
rect 571542 609578 582820 609814
rect 1104 609494 582820 609578
rect 1104 609258 12986 609494
rect 13222 609258 13306 609494
rect 13542 609258 50186 609494
rect 50422 609258 50506 609494
rect 50742 609258 87386 609494
rect 87622 609258 87706 609494
rect 87942 609258 124586 609494
rect 124822 609258 124906 609494
rect 125142 609258 161786 609494
rect 162022 609258 162106 609494
rect 162342 609258 198986 609494
rect 199222 609258 199306 609494
rect 199542 609258 236186 609494
rect 236422 609258 236506 609494
rect 236742 609258 273386 609494
rect 273622 609258 273706 609494
rect 273942 609258 310586 609494
rect 310822 609258 310906 609494
rect 311142 609258 347786 609494
rect 348022 609258 348106 609494
rect 348342 609258 384986 609494
rect 385222 609258 385306 609494
rect 385542 609258 422186 609494
rect 422422 609258 422506 609494
rect 422742 609258 459386 609494
rect 459622 609258 459706 609494
rect 459942 609258 496586 609494
rect 496822 609258 496906 609494
rect 497142 609258 533786 609494
rect 534022 609258 534106 609494
rect 534342 609258 570986 609494
rect 571222 609258 571306 609494
rect 571542 609258 582820 609494
rect 1104 609226 582820 609258
rect 1104 606094 582820 606126
rect 1104 605858 9266 606094
rect 9502 605858 9586 606094
rect 9822 605858 46466 606094
rect 46702 605858 46786 606094
rect 47022 605858 83666 606094
rect 83902 605858 83986 606094
rect 84222 605858 120866 606094
rect 121102 605858 121186 606094
rect 121422 605858 158066 606094
rect 158302 605858 158386 606094
rect 158622 605858 195266 606094
rect 195502 605858 195586 606094
rect 195822 605858 232466 606094
rect 232702 605858 232786 606094
rect 233022 605858 269666 606094
rect 269902 605858 269986 606094
rect 270222 605858 306866 606094
rect 307102 605858 307186 606094
rect 307422 605858 344066 606094
rect 344302 605858 344386 606094
rect 344622 605858 381266 606094
rect 381502 605858 381586 606094
rect 381822 605858 418466 606094
rect 418702 605858 418786 606094
rect 419022 605858 455666 606094
rect 455902 605858 455986 606094
rect 456222 605858 492866 606094
rect 493102 605858 493186 606094
rect 493422 605858 530066 606094
rect 530302 605858 530386 606094
rect 530622 605858 567266 606094
rect 567502 605858 567586 606094
rect 567822 605858 582820 606094
rect 1104 605774 582820 605858
rect 1104 605538 9266 605774
rect 9502 605538 9586 605774
rect 9822 605538 46466 605774
rect 46702 605538 46786 605774
rect 47022 605538 83666 605774
rect 83902 605538 83986 605774
rect 84222 605538 120866 605774
rect 121102 605538 121186 605774
rect 121422 605538 158066 605774
rect 158302 605538 158386 605774
rect 158622 605538 195266 605774
rect 195502 605538 195586 605774
rect 195822 605538 232466 605774
rect 232702 605538 232786 605774
rect 233022 605538 269666 605774
rect 269902 605538 269986 605774
rect 270222 605538 306866 605774
rect 307102 605538 307186 605774
rect 307422 605538 344066 605774
rect 344302 605538 344386 605774
rect 344622 605538 381266 605774
rect 381502 605538 381586 605774
rect 381822 605538 418466 605774
rect 418702 605538 418786 605774
rect 419022 605538 455666 605774
rect 455902 605538 455986 605774
rect 456222 605538 492866 605774
rect 493102 605538 493186 605774
rect 493422 605538 530066 605774
rect 530302 605538 530386 605774
rect 530622 605538 567266 605774
rect 567502 605538 567586 605774
rect 567822 605538 582820 605774
rect 1104 605506 582820 605538
rect 1104 602374 582820 602406
rect 1104 602138 5546 602374
rect 5782 602138 5866 602374
rect 6102 602138 42746 602374
rect 42982 602138 43066 602374
rect 43302 602138 79946 602374
rect 80182 602138 80266 602374
rect 80502 602138 117146 602374
rect 117382 602138 117466 602374
rect 117702 602138 154346 602374
rect 154582 602138 154666 602374
rect 154902 602138 191546 602374
rect 191782 602138 191866 602374
rect 192102 602138 228746 602374
rect 228982 602138 229066 602374
rect 229302 602138 265946 602374
rect 266182 602138 266266 602374
rect 266502 602138 303146 602374
rect 303382 602138 303466 602374
rect 303702 602138 340346 602374
rect 340582 602138 340666 602374
rect 340902 602138 377546 602374
rect 377782 602138 377866 602374
rect 378102 602138 414746 602374
rect 414982 602138 415066 602374
rect 415302 602138 451946 602374
rect 452182 602138 452266 602374
rect 452502 602138 489146 602374
rect 489382 602138 489466 602374
rect 489702 602138 526346 602374
rect 526582 602138 526666 602374
rect 526902 602138 563546 602374
rect 563782 602138 563866 602374
rect 564102 602138 582820 602374
rect 1104 602054 582820 602138
rect 1104 601818 5546 602054
rect 5782 601818 5866 602054
rect 6102 601818 42746 602054
rect 42982 601818 43066 602054
rect 43302 601818 79946 602054
rect 80182 601818 80266 602054
rect 80502 601818 117146 602054
rect 117382 601818 117466 602054
rect 117702 601818 154346 602054
rect 154582 601818 154666 602054
rect 154902 601818 191546 602054
rect 191782 601818 191866 602054
rect 192102 601818 228746 602054
rect 228982 601818 229066 602054
rect 229302 601818 265946 602054
rect 266182 601818 266266 602054
rect 266502 601818 303146 602054
rect 303382 601818 303466 602054
rect 303702 601818 340346 602054
rect 340582 601818 340666 602054
rect 340902 601818 377546 602054
rect 377782 601818 377866 602054
rect 378102 601818 414746 602054
rect 414982 601818 415066 602054
rect 415302 601818 451946 602054
rect 452182 601818 452266 602054
rect 452502 601818 489146 602054
rect 489382 601818 489466 602054
rect 489702 601818 526346 602054
rect 526582 601818 526666 602054
rect 526902 601818 563546 602054
rect 563782 601818 563866 602054
rect 564102 601818 582820 602054
rect 1104 601786 582820 601818
rect 1104 598654 582820 598686
rect 1104 598418 1826 598654
rect 2062 598418 2146 598654
rect 2382 598418 39026 598654
rect 39262 598418 39346 598654
rect 39582 598418 76226 598654
rect 76462 598418 76546 598654
rect 76782 598418 113426 598654
rect 113662 598418 113746 598654
rect 113982 598418 150626 598654
rect 150862 598418 150946 598654
rect 151182 598418 187826 598654
rect 188062 598418 188146 598654
rect 188382 598418 225026 598654
rect 225262 598418 225346 598654
rect 225582 598418 262226 598654
rect 262462 598418 262546 598654
rect 262782 598418 299426 598654
rect 299662 598418 299746 598654
rect 299982 598418 336626 598654
rect 336862 598418 336946 598654
rect 337182 598418 373826 598654
rect 374062 598418 374146 598654
rect 374382 598418 411026 598654
rect 411262 598418 411346 598654
rect 411582 598418 448226 598654
rect 448462 598418 448546 598654
rect 448782 598418 485426 598654
rect 485662 598418 485746 598654
rect 485982 598418 522626 598654
rect 522862 598418 522946 598654
rect 523182 598418 559826 598654
rect 560062 598418 560146 598654
rect 560382 598418 582820 598654
rect 1104 598334 582820 598418
rect 1104 598098 1826 598334
rect 2062 598098 2146 598334
rect 2382 598098 39026 598334
rect 39262 598098 39346 598334
rect 39582 598098 76226 598334
rect 76462 598098 76546 598334
rect 76782 598098 113426 598334
rect 113662 598098 113746 598334
rect 113982 598098 150626 598334
rect 150862 598098 150946 598334
rect 151182 598098 187826 598334
rect 188062 598098 188146 598334
rect 188382 598098 225026 598334
rect 225262 598098 225346 598334
rect 225582 598098 262226 598334
rect 262462 598098 262546 598334
rect 262782 598098 299426 598334
rect 299662 598098 299746 598334
rect 299982 598098 336626 598334
rect 336862 598098 336946 598334
rect 337182 598098 373826 598334
rect 374062 598098 374146 598334
rect 374382 598098 411026 598334
rect 411262 598098 411346 598334
rect 411582 598098 448226 598334
rect 448462 598098 448546 598334
rect 448782 598098 485426 598334
rect 485662 598098 485746 598334
rect 485982 598098 522626 598334
rect 522862 598098 522946 598334
rect 523182 598098 559826 598334
rect 560062 598098 560146 598334
rect 560382 598098 582820 598334
rect 1104 598066 582820 598098
rect 1104 587494 582820 587526
rect 1104 587258 27866 587494
rect 28102 587258 28186 587494
rect 28422 587258 65066 587494
rect 65302 587258 65386 587494
rect 65622 587258 102266 587494
rect 102502 587258 102586 587494
rect 102822 587258 139466 587494
rect 139702 587258 139786 587494
rect 140022 587258 176666 587494
rect 176902 587258 176986 587494
rect 177222 587258 213866 587494
rect 214102 587258 214186 587494
rect 214422 587258 251066 587494
rect 251302 587258 251386 587494
rect 251622 587258 288266 587494
rect 288502 587258 288586 587494
rect 288822 587258 325466 587494
rect 325702 587258 325786 587494
rect 326022 587258 362666 587494
rect 362902 587258 362986 587494
rect 363222 587258 399866 587494
rect 400102 587258 400186 587494
rect 400422 587258 437066 587494
rect 437302 587258 437386 587494
rect 437622 587258 474266 587494
rect 474502 587258 474586 587494
rect 474822 587258 511466 587494
rect 511702 587258 511786 587494
rect 512022 587258 548666 587494
rect 548902 587258 548986 587494
rect 549222 587258 582820 587494
rect 1104 587174 582820 587258
rect 1104 586938 27866 587174
rect 28102 586938 28186 587174
rect 28422 586938 65066 587174
rect 65302 586938 65386 587174
rect 65622 586938 102266 587174
rect 102502 586938 102586 587174
rect 102822 586938 139466 587174
rect 139702 586938 139786 587174
rect 140022 586938 176666 587174
rect 176902 586938 176986 587174
rect 177222 586938 213866 587174
rect 214102 586938 214186 587174
rect 214422 586938 251066 587174
rect 251302 586938 251386 587174
rect 251622 586938 288266 587174
rect 288502 586938 288586 587174
rect 288822 586938 325466 587174
rect 325702 586938 325786 587174
rect 326022 586938 362666 587174
rect 362902 586938 362986 587174
rect 363222 586938 399866 587174
rect 400102 586938 400186 587174
rect 400422 586938 437066 587174
rect 437302 586938 437386 587174
rect 437622 586938 474266 587174
rect 474502 586938 474586 587174
rect 474822 586938 511466 587174
rect 511702 586938 511786 587174
rect 512022 586938 548666 587174
rect 548902 586938 548986 587174
rect 549222 586938 582820 587174
rect 1104 586906 582820 586938
rect 1104 583774 582820 583806
rect 1104 583538 24146 583774
rect 24382 583538 24466 583774
rect 24702 583538 61346 583774
rect 61582 583538 61666 583774
rect 61902 583538 98546 583774
rect 98782 583538 98866 583774
rect 99102 583538 135746 583774
rect 135982 583538 136066 583774
rect 136302 583538 172946 583774
rect 173182 583538 173266 583774
rect 173502 583538 210146 583774
rect 210382 583538 210466 583774
rect 210702 583538 247346 583774
rect 247582 583538 247666 583774
rect 247902 583538 284546 583774
rect 284782 583538 284866 583774
rect 285102 583538 321746 583774
rect 321982 583538 322066 583774
rect 322302 583538 358946 583774
rect 359182 583538 359266 583774
rect 359502 583538 396146 583774
rect 396382 583538 396466 583774
rect 396702 583538 433346 583774
rect 433582 583538 433666 583774
rect 433902 583538 470546 583774
rect 470782 583538 470866 583774
rect 471102 583538 507746 583774
rect 507982 583538 508066 583774
rect 508302 583538 544946 583774
rect 545182 583538 545266 583774
rect 545502 583538 582146 583774
rect 582382 583538 582466 583774
rect 582702 583538 582820 583774
rect 1104 583454 582820 583538
rect 1104 583218 24146 583454
rect 24382 583218 24466 583454
rect 24702 583218 61346 583454
rect 61582 583218 61666 583454
rect 61902 583218 98546 583454
rect 98782 583218 98866 583454
rect 99102 583218 135746 583454
rect 135982 583218 136066 583454
rect 136302 583218 172946 583454
rect 173182 583218 173266 583454
rect 173502 583218 210146 583454
rect 210382 583218 210466 583454
rect 210702 583218 247346 583454
rect 247582 583218 247666 583454
rect 247902 583218 284546 583454
rect 284782 583218 284866 583454
rect 285102 583218 321746 583454
rect 321982 583218 322066 583454
rect 322302 583218 358946 583454
rect 359182 583218 359266 583454
rect 359502 583218 396146 583454
rect 396382 583218 396466 583454
rect 396702 583218 433346 583454
rect 433582 583218 433666 583454
rect 433902 583218 470546 583454
rect 470782 583218 470866 583454
rect 471102 583218 507746 583454
rect 507982 583218 508066 583454
rect 508302 583218 544946 583454
rect 545182 583218 545266 583454
rect 545502 583218 582146 583454
rect 582382 583218 582466 583454
rect 582702 583218 582820 583454
rect 1104 583186 582820 583218
rect 1104 580054 582820 580086
rect 1104 579818 20426 580054
rect 20662 579818 20746 580054
rect 20982 579818 57626 580054
rect 57862 579818 57946 580054
rect 58182 579818 94826 580054
rect 95062 579818 95146 580054
rect 95382 579818 132026 580054
rect 132262 579818 132346 580054
rect 132582 579818 169226 580054
rect 169462 579818 169546 580054
rect 169782 579818 206426 580054
rect 206662 579818 206746 580054
rect 206982 579818 243626 580054
rect 243862 579818 243946 580054
rect 244182 579818 280826 580054
rect 281062 579818 281146 580054
rect 281382 579818 318026 580054
rect 318262 579818 318346 580054
rect 318582 579818 355226 580054
rect 355462 579818 355546 580054
rect 355782 579818 392426 580054
rect 392662 579818 392746 580054
rect 392982 579818 429626 580054
rect 429862 579818 429946 580054
rect 430182 579818 466826 580054
rect 467062 579818 467146 580054
rect 467382 579818 504026 580054
rect 504262 579818 504346 580054
rect 504582 579818 541226 580054
rect 541462 579818 541546 580054
rect 541782 579818 578426 580054
rect 578662 579818 578746 580054
rect 578982 579818 582820 580054
rect 1104 579734 582820 579818
rect 1104 579498 20426 579734
rect 20662 579498 20746 579734
rect 20982 579498 57626 579734
rect 57862 579498 57946 579734
rect 58182 579498 94826 579734
rect 95062 579498 95146 579734
rect 95382 579498 132026 579734
rect 132262 579498 132346 579734
rect 132582 579498 169226 579734
rect 169462 579498 169546 579734
rect 169782 579498 206426 579734
rect 206662 579498 206746 579734
rect 206982 579498 243626 579734
rect 243862 579498 243946 579734
rect 244182 579498 280826 579734
rect 281062 579498 281146 579734
rect 281382 579498 318026 579734
rect 318262 579498 318346 579734
rect 318582 579498 355226 579734
rect 355462 579498 355546 579734
rect 355782 579498 392426 579734
rect 392662 579498 392746 579734
rect 392982 579498 429626 579734
rect 429862 579498 429946 579734
rect 430182 579498 466826 579734
rect 467062 579498 467146 579734
rect 467382 579498 504026 579734
rect 504262 579498 504346 579734
rect 504582 579498 541226 579734
rect 541462 579498 541546 579734
rect 541782 579498 578426 579734
rect 578662 579498 578746 579734
rect 578982 579498 582820 579734
rect 1104 579466 582820 579498
rect 1104 576334 582820 576366
rect 1104 576098 16706 576334
rect 16942 576098 17026 576334
rect 17262 576098 53906 576334
rect 54142 576098 54226 576334
rect 54462 576098 91106 576334
rect 91342 576098 91426 576334
rect 91662 576098 128306 576334
rect 128542 576098 128626 576334
rect 128862 576098 165506 576334
rect 165742 576098 165826 576334
rect 166062 576098 202706 576334
rect 202942 576098 203026 576334
rect 203262 576098 239906 576334
rect 240142 576098 240226 576334
rect 240462 576098 277106 576334
rect 277342 576098 277426 576334
rect 277662 576098 314306 576334
rect 314542 576098 314626 576334
rect 314862 576098 351506 576334
rect 351742 576098 351826 576334
rect 352062 576098 388706 576334
rect 388942 576098 389026 576334
rect 389262 576098 425906 576334
rect 426142 576098 426226 576334
rect 426462 576098 463106 576334
rect 463342 576098 463426 576334
rect 463662 576098 500306 576334
rect 500542 576098 500626 576334
rect 500862 576098 537506 576334
rect 537742 576098 537826 576334
rect 538062 576098 574706 576334
rect 574942 576098 575026 576334
rect 575262 576098 582820 576334
rect 1104 576014 582820 576098
rect 1104 575778 16706 576014
rect 16942 575778 17026 576014
rect 17262 575778 53906 576014
rect 54142 575778 54226 576014
rect 54462 575778 91106 576014
rect 91342 575778 91426 576014
rect 91662 575778 128306 576014
rect 128542 575778 128626 576014
rect 128862 575778 165506 576014
rect 165742 575778 165826 576014
rect 166062 575778 202706 576014
rect 202942 575778 203026 576014
rect 203262 575778 239906 576014
rect 240142 575778 240226 576014
rect 240462 575778 277106 576014
rect 277342 575778 277426 576014
rect 277662 575778 314306 576014
rect 314542 575778 314626 576014
rect 314862 575778 351506 576014
rect 351742 575778 351826 576014
rect 352062 575778 388706 576014
rect 388942 575778 389026 576014
rect 389262 575778 425906 576014
rect 426142 575778 426226 576014
rect 426462 575778 463106 576014
rect 463342 575778 463426 576014
rect 463662 575778 500306 576014
rect 500542 575778 500626 576014
rect 500862 575778 537506 576014
rect 537742 575778 537826 576014
rect 538062 575778 574706 576014
rect 574942 575778 575026 576014
rect 575262 575778 582820 576014
rect 1104 575746 582820 575778
rect 1104 572614 582820 572646
rect 1104 572378 12986 572614
rect 13222 572378 13306 572614
rect 13542 572378 50186 572614
rect 50422 572378 50506 572614
rect 50742 572378 87386 572614
rect 87622 572378 87706 572614
rect 87942 572378 124586 572614
rect 124822 572378 124906 572614
rect 125142 572378 161786 572614
rect 162022 572378 162106 572614
rect 162342 572378 198986 572614
rect 199222 572378 199306 572614
rect 199542 572378 236186 572614
rect 236422 572378 236506 572614
rect 236742 572378 273386 572614
rect 273622 572378 273706 572614
rect 273942 572378 310586 572614
rect 310822 572378 310906 572614
rect 311142 572378 347786 572614
rect 348022 572378 348106 572614
rect 348342 572378 384986 572614
rect 385222 572378 385306 572614
rect 385542 572378 422186 572614
rect 422422 572378 422506 572614
rect 422742 572378 459386 572614
rect 459622 572378 459706 572614
rect 459942 572378 496586 572614
rect 496822 572378 496906 572614
rect 497142 572378 533786 572614
rect 534022 572378 534106 572614
rect 534342 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 582820 572614
rect 1104 572294 582820 572378
rect 1104 572058 12986 572294
rect 13222 572058 13306 572294
rect 13542 572058 50186 572294
rect 50422 572058 50506 572294
rect 50742 572058 87386 572294
rect 87622 572058 87706 572294
rect 87942 572058 124586 572294
rect 124822 572058 124906 572294
rect 125142 572058 161786 572294
rect 162022 572058 162106 572294
rect 162342 572058 198986 572294
rect 199222 572058 199306 572294
rect 199542 572058 236186 572294
rect 236422 572058 236506 572294
rect 236742 572058 273386 572294
rect 273622 572058 273706 572294
rect 273942 572058 310586 572294
rect 310822 572058 310906 572294
rect 311142 572058 347786 572294
rect 348022 572058 348106 572294
rect 348342 572058 384986 572294
rect 385222 572058 385306 572294
rect 385542 572058 422186 572294
rect 422422 572058 422506 572294
rect 422742 572058 459386 572294
rect 459622 572058 459706 572294
rect 459942 572058 496586 572294
rect 496822 572058 496906 572294
rect 497142 572058 533786 572294
rect 534022 572058 534106 572294
rect 534342 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 582820 572294
rect 1104 572026 582820 572058
rect 1104 568894 582820 568926
rect 1104 568658 9266 568894
rect 9502 568658 9586 568894
rect 9822 568658 46466 568894
rect 46702 568658 46786 568894
rect 47022 568658 83666 568894
rect 83902 568658 83986 568894
rect 84222 568658 120866 568894
rect 121102 568658 121186 568894
rect 121422 568658 158066 568894
rect 158302 568658 158386 568894
rect 158622 568658 195266 568894
rect 195502 568658 195586 568894
rect 195822 568658 232466 568894
rect 232702 568658 232786 568894
rect 233022 568658 269666 568894
rect 269902 568658 269986 568894
rect 270222 568658 306866 568894
rect 307102 568658 307186 568894
rect 307422 568658 344066 568894
rect 344302 568658 344386 568894
rect 344622 568658 381266 568894
rect 381502 568658 381586 568894
rect 381822 568658 418466 568894
rect 418702 568658 418786 568894
rect 419022 568658 455666 568894
rect 455902 568658 455986 568894
rect 456222 568658 492866 568894
rect 493102 568658 493186 568894
rect 493422 568658 530066 568894
rect 530302 568658 530386 568894
rect 530622 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 582820 568894
rect 1104 568574 582820 568658
rect 1104 568338 9266 568574
rect 9502 568338 9586 568574
rect 9822 568338 46466 568574
rect 46702 568338 46786 568574
rect 47022 568338 83666 568574
rect 83902 568338 83986 568574
rect 84222 568338 120866 568574
rect 121102 568338 121186 568574
rect 121422 568338 158066 568574
rect 158302 568338 158386 568574
rect 158622 568338 195266 568574
rect 195502 568338 195586 568574
rect 195822 568338 232466 568574
rect 232702 568338 232786 568574
rect 233022 568338 269666 568574
rect 269902 568338 269986 568574
rect 270222 568338 306866 568574
rect 307102 568338 307186 568574
rect 307422 568338 344066 568574
rect 344302 568338 344386 568574
rect 344622 568338 381266 568574
rect 381502 568338 381586 568574
rect 381822 568338 418466 568574
rect 418702 568338 418786 568574
rect 419022 568338 455666 568574
rect 455902 568338 455986 568574
rect 456222 568338 492866 568574
rect 493102 568338 493186 568574
rect 493422 568338 530066 568574
rect 530302 568338 530386 568574
rect 530622 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 582820 568574
rect 1104 568306 582820 568338
rect 1104 565174 582820 565206
rect 1104 564938 5546 565174
rect 5782 564938 5866 565174
rect 6102 564938 42746 565174
rect 42982 564938 43066 565174
rect 43302 564938 79946 565174
rect 80182 564938 80266 565174
rect 80502 564938 117146 565174
rect 117382 564938 117466 565174
rect 117702 564938 154346 565174
rect 154582 564938 154666 565174
rect 154902 564938 191546 565174
rect 191782 564938 191866 565174
rect 192102 564938 228746 565174
rect 228982 564938 229066 565174
rect 229302 564938 265946 565174
rect 266182 564938 266266 565174
rect 266502 564938 303146 565174
rect 303382 564938 303466 565174
rect 303702 564938 340346 565174
rect 340582 564938 340666 565174
rect 340902 564938 377546 565174
rect 377782 564938 377866 565174
rect 378102 564938 414746 565174
rect 414982 564938 415066 565174
rect 415302 564938 451946 565174
rect 452182 564938 452266 565174
rect 452502 564938 489146 565174
rect 489382 564938 489466 565174
rect 489702 564938 526346 565174
rect 526582 564938 526666 565174
rect 526902 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 582820 565174
rect 1104 564854 582820 564938
rect 1104 564618 5546 564854
rect 5782 564618 5866 564854
rect 6102 564618 42746 564854
rect 42982 564618 43066 564854
rect 43302 564618 79946 564854
rect 80182 564618 80266 564854
rect 80502 564618 117146 564854
rect 117382 564618 117466 564854
rect 117702 564618 154346 564854
rect 154582 564618 154666 564854
rect 154902 564618 191546 564854
rect 191782 564618 191866 564854
rect 192102 564618 228746 564854
rect 228982 564618 229066 564854
rect 229302 564618 265946 564854
rect 266182 564618 266266 564854
rect 266502 564618 303146 564854
rect 303382 564618 303466 564854
rect 303702 564618 340346 564854
rect 340582 564618 340666 564854
rect 340902 564618 377546 564854
rect 377782 564618 377866 564854
rect 378102 564618 414746 564854
rect 414982 564618 415066 564854
rect 415302 564618 451946 564854
rect 452182 564618 452266 564854
rect 452502 564618 489146 564854
rect 489382 564618 489466 564854
rect 489702 564618 526346 564854
rect 526582 564618 526666 564854
rect 526902 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 582820 564854
rect 1104 564586 582820 564618
rect 1104 561454 582820 561486
rect 1104 561218 1826 561454
rect 2062 561218 2146 561454
rect 2382 561218 39026 561454
rect 39262 561218 39346 561454
rect 39582 561218 76226 561454
rect 76462 561218 76546 561454
rect 76782 561218 113426 561454
rect 113662 561218 113746 561454
rect 113982 561218 150626 561454
rect 150862 561218 150946 561454
rect 151182 561218 187826 561454
rect 188062 561218 188146 561454
rect 188382 561218 225026 561454
rect 225262 561218 225346 561454
rect 225582 561218 262226 561454
rect 262462 561218 262546 561454
rect 262782 561218 299426 561454
rect 299662 561218 299746 561454
rect 299982 561218 336626 561454
rect 336862 561218 336946 561454
rect 337182 561218 373826 561454
rect 374062 561218 374146 561454
rect 374382 561218 411026 561454
rect 411262 561218 411346 561454
rect 411582 561218 448226 561454
rect 448462 561218 448546 561454
rect 448782 561218 485426 561454
rect 485662 561218 485746 561454
rect 485982 561218 522626 561454
rect 522862 561218 522946 561454
rect 523182 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 582820 561454
rect 1104 561134 582820 561218
rect 1104 560898 1826 561134
rect 2062 560898 2146 561134
rect 2382 560898 39026 561134
rect 39262 560898 39346 561134
rect 39582 560898 76226 561134
rect 76462 560898 76546 561134
rect 76782 560898 113426 561134
rect 113662 560898 113746 561134
rect 113982 560898 150626 561134
rect 150862 560898 150946 561134
rect 151182 560898 187826 561134
rect 188062 560898 188146 561134
rect 188382 560898 225026 561134
rect 225262 560898 225346 561134
rect 225582 560898 262226 561134
rect 262462 560898 262546 561134
rect 262782 560898 299426 561134
rect 299662 560898 299746 561134
rect 299982 560898 336626 561134
rect 336862 560898 336946 561134
rect 337182 560898 373826 561134
rect 374062 560898 374146 561134
rect 374382 560898 411026 561134
rect 411262 560898 411346 561134
rect 411582 560898 448226 561134
rect 448462 560898 448546 561134
rect 448782 560898 485426 561134
rect 485662 560898 485746 561134
rect 485982 560898 522626 561134
rect 522862 560898 522946 561134
rect 523182 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 582820 561134
rect 1104 560866 582820 560898
rect 1104 550294 582820 550326
rect 1104 550058 27866 550294
rect 28102 550058 28186 550294
rect 28422 550058 65066 550294
rect 65302 550058 65386 550294
rect 65622 550058 102266 550294
rect 102502 550058 102586 550294
rect 102822 550058 139466 550294
rect 139702 550058 139786 550294
rect 140022 550058 176666 550294
rect 176902 550058 176986 550294
rect 177222 550058 213866 550294
rect 214102 550058 214186 550294
rect 214422 550058 251066 550294
rect 251302 550058 251386 550294
rect 251622 550058 288266 550294
rect 288502 550058 288586 550294
rect 288822 550058 325466 550294
rect 325702 550058 325786 550294
rect 326022 550058 362666 550294
rect 362902 550058 362986 550294
rect 363222 550058 399866 550294
rect 400102 550058 400186 550294
rect 400422 550058 437066 550294
rect 437302 550058 437386 550294
rect 437622 550058 474266 550294
rect 474502 550058 474586 550294
rect 474822 550058 511466 550294
rect 511702 550058 511786 550294
rect 512022 550058 548666 550294
rect 548902 550058 548986 550294
rect 549222 550058 582820 550294
rect 1104 549974 582820 550058
rect 1104 549738 27866 549974
rect 28102 549738 28186 549974
rect 28422 549738 65066 549974
rect 65302 549738 65386 549974
rect 65622 549738 102266 549974
rect 102502 549738 102586 549974
rect 102822 549738 139466 549974
rect 139702 549738 139786 549974
rect 140022 549738 176666 549974
rect 176902 549738 176986 549974
rect 177222 549738 213866 549974
rect 214102 549738 214186 549974
rect 214422 549738 251066 549974
rect 251302 549738 251386 549974
rect 251622 549738 288266 549974
rect 288502 549738 288586 549974
rect 288822 549738 325466 549974
rect 325702 549738 325786 549974
rect 326022 549738 362666 549974
rect 362902 549738 362986 549974
rect 363222 549738 399866 549974
rect 400102 549738 400186 549974
rect 400422 549738 437066 549974
rect 437302 549738 437386 549974
rect 437622 549738 474266 549974
rect 474502 549738 474586 549974
rect 474822 549738 511466 549974
rect 511702 549738 511786 549974
rect 512022 549738 548666 549974
rect 548902 549738 548986 549974
rect 549222 549738 582820 549974
rect 1104 549706 582820 549738
rect 1104 546574 582820 546606
rect 1104 546338 24146 546574
rect 24382 546338 24466 546574
rect 24702 546338 61346 546574
rect 61582 546338 61666 546574
rect 61902 546338 98546 546574
rect 98782 546338 98866 546574
rect 99102 546338 135746 546574
rect 135982 546338 136066 546574
rect 136302 546338 172946 546574
rect 173182 546338 173266 546574
rect 173502 546338 210146 546574
rect 210382 546338 210466 546574
rect 210702 546338 247346 546574
rect 247582 546338 247666 546574
rect 247902 546338 284546 546574
rect 284782 546338 284866 546574
rect 285102 546338 321746 546574
rect 321982 546338 322066 546574
rect 322302 546338 358946 546574
rect 359182 546338 359266 546574
rect 359502 546338 396146 546574
rect 396382 546338 396466 546574
rect 396702 546338 433346 546574
rect 433582 546338 433666 546574
rect 433902 546338 470546 546574
rect 470782 546338 470866 546574
rect 471102 546338 507746 546574
rect 507982 546338 508066 546574
rect 508302 546338 544946 546574
rect 545182 546338 545266 546574
rect 545502 546338 582146 546574
rect 582382 546338 582466 546574
rect 582702 546338 582820 546574
rect 1104 546254 582820 546338
rect 1104 546018 24146 546254
rect 24382 546018 24466 546254
rect 24702 546018 61346 546254
rect 61582 546018 61666 546254
rect 61902 546018 98546 546254
rect 98782 546018 98866 546254
rect 99102 546018 135746 546254
rect 135982 546018 136066 546254
rect 136302 546018 172946 546254
rect 173182 546018 173266 546254
rect 173502 546018 210146 546254
rect 210382 546018 210466 546254
rect 210702 546018 247346 546254
rect 247582 546018 247666 546254
rect 247902 546018 284546 546254
rect 284782 546018 284866 546254
rect 285102 546018 321746 546254
rect 321982 546018 322066 546254
rect 322302 546018 358946 546254
rect 359182 546018 359266 546254
rect 359502 546018 396146 546254
rect 396382 546018 396466 546254
rect 396702 546018 433346 546254
rect 433582 546018 433666 546254
rect 433902 546018 470546 546254
rect 470782 546018 470866 546254
rect 471102 546018 507746 546254
rect 507982 546018 508066 546254
rect 508302 546018 544946 546254
rect 545182 546018 545266 546254
rect 545502 546018 582146 546254
rect 582382 546018 582466 546254
rect 582702 546018 582820 546254
rect 1104 545986 582820 546018
rect 1104 542854 582820 542886
rect 1104 542618 20426 542854
rect 20662 542618 20746 542854
rect 20982 542618 57626 542854
rect 57862 542618 57946 542854
rect 58182 542618 94826 542854
rect 95062 542618 95146 542854
rect 95382 542618 132026 542854
rect 132262 542618 132346 542854
rect 132582 542618 169226 542854
rect 169462 542618 169546 542854
rect 169782 542618 206426 542854
rect 206662 542618 206746 542854
rect 206982 542618 243626 542854
rect 243862 542618 243946 542854
rect 244182 542618 280826 542854
rect 281062 542618 281146 542854
rect 281382 542618 318026 542854
rect 318262 542618 318346 542854
rect 318582 542618 355226 542854
rect 355462 542618 355546 542854
rect 355782 542618 392426 542854
rect 392662 542618 392746 542854
rect 392982 542618 429626 542854
rect 429862 542618 429946 542854
rect 430182 542618 466826 542854
rect 467062 542618 467146 542854
rect 467382 542618 504026 542854
rect 504262 542618 504346 542854
rect 504582 542618 541226 542854
rect 541462 542618 541546 542854
rect 541782 542618 578426 542854
rect 578662 542618 578746 542854
rect 578982 542618 582820 542854
rect 1104 542534 582820 542618
rect 1104 542298 20426 542534
rect 20662 542298 20746 542534
rect 20982 542298 57626 542534
rect 57862 542298 57946 542534
rect 58182 542298 94826 542534
rect 95062 542298 95146 542534
rect 95382 542298 132026 542534
rect 132262 542298 132346 542534
rect 132582 542298 169226 542534
rect 169462 542298 169546 542534
rect 169782 542298 206426 542534
rect 206662 542298 206746 542534
rect 206982 542298 243626 542534
rect 243862 542298 243946 542534
rect 244182 542298 280826 542534
rect 281062 542298 281146 542534
rect 281382 542298 318026 542534
rect 318262 542298 318346 542534
rect 318582 542298 355226 542534
rect 355462 542298 355546 542534
rect 355782 542298 392426 542534
rect 392662 542298 392746 542534
rect 392982 542298 429626 542534
rect 429862 542298 429946 542534
rect 430182 542298 466826 542534
rect 467062 542298 467146 542534
rect 467382 542298 504026 542534
rect 504262 542298 504346 542534
rect 504582 542298 541226 542534
rect 541462 542298 541546 542534
rect 541782 542298 578426 542534
rect 578662 542298 578746 542534
rect 578982 542298 582820 542534
rect 1104 542266 582820 542298
rect 1104 539134 582820 539166
rect 1104 538898 16706 539134
rect 16942 538898 17026 539134
rect 17262 538898 53906 539134
rect 54142 538898 54226 539134
rect 54462 538898 91106 539134
rect 91342 538898 91426 539134
rect 91662 538898 128306 539134
rect 128542 538898 128626 539134
rect 128862 538898 165506 539134
rect 165742 538898 165826 539134
rect 166062 538898 202706 539134
rect 202942 538898 203026 539134
rect 203262 538898 239906 539134
rect 240142 538898 240226 539134
rect 240462 538898 277106 539134
rect 277342 538898 277426 539134
rect 277662 538898 314306 539134
rect 314542 538898 314626 539134
rect 314862 538898 351506 539134
rect 351742 538898 351826 539134
rect 352062 538898 388706 539134
rect 388942 538898 389026 539134
rect 389262 538898 425906 539134
rect 426142 538898 426226 539134
rect 426462 538898 463106 539134
rect 463342 538898 463426 539134
rect 463662 538898 500306 539134
rect 500542 538898 500626 539134
rect 500862 538898 537506 539134
rect 537742 538898 537826 539134
rect 538062 538898 574706 539134
rect 574942 538898 575026 539134
rect 575262 538898 582820 539134
rect 1104 538814 582820 538898
rect 1104 538578 16706 538814
rect 16942 538578 17026 538814
rect 17262 538578 53906 538814
rect 54142 538578 54226 538814
rect 54462 538578 91106 538814
rect 91342 538578 91426 538814
rect 91662 538578 128306 538814
rect 128542 538578 128626 538814
rect 128862 538578 165506 538814
rect 165742 538578 165826 538814
rect 166062 538578 202706 538814
rect 202942 538578 203026 538814
rect 203262 538578 239906 538814
rect 240142 538578 240226 538814
rect 240462 538578 277106 538814
rect 277342 538578 277426 538814
rect 277662 538578 314306 538814
rect 314542 538578 314626 538814
rect 314862 538578 351506 538814
rect 351742 538578 351826 538814
rect 352062 538578 388706 538814
rect 388942 538578 389026 538814
rect 389262 538578 425906 538814
rect 426142 538578 426226 538814
rect 426462 538578 463106 538814
rect 463342 538578 463426 538814
rect 463662 538578 500306 538814
rect 500542 538578 500626 538814
rect 500862 538578 537506 538814
rect 537742 538578 537826 538814
rect 538062 538578 574706 538814
rect 574942 538578 575026 538814
rect 575262 538578 582820 538814
rect 1104 538546 582820 538578
rect 1104 535414 582820 535446
rect 1104 535178 12986 535414
rect 13222 535178 13306 535414
rect 13542 535178 50186 535414
rect 50422 535178 50506 535414
rect 50742 535178 87386 535414
rect 87622 535178 87706 535414
rect 87942 535178 124586 535414
rect 124822 535178 124906 535414
rect 125142 535178 161786 535414
rect 162022 535178 162106 535414
rect 162342 535178 198986 535414
rect 199222 535178 199306 535414
rect 199542 535178 236186 535414
rect 236422 535178 236506 535414
rect 236742 535178 273386 535414
rect 273622 535178 273706 535414
rect 273942 535178 310586 535414
rect 310822 535178 310906 535414
rect 311142 535178 347786 535414
rect 348022 535178 348106 535414
rect 348342 535178 384986 535414
rect 385222 535178 385306 535414
rect 385542 535178 422186 535414
rect 422422 535178 422506 535414
rect 422742 535178 459386 535414
rect 459622 535178 459706 535414
rect 459942 535178 496586 535414
rect 496822 535178 496906 535414
rect 497142 535178 533786 535414
rect 534022 535178 534106 535414
rect 534342 535178 570986 535414
rect 571222 535178 571306 535414
rect 571542 535178 582820 535414
rect 1104 535094 582820 535178
rect 1104 534858 12986 535094
rect 13222 534858 13306 535094
rect 13542 534858 50186 535094
rect 50422 534858 50506 535094
rect 50742 534858 87386 535094
rect 87622 534858 87706 535094
rect 87942 534858 124586 535094
rect 124822 534858 124906 535094
rect 125142 534858 161786 535094
rect 162022 534858 162106 535094
rect 162342 534858 198986 535094
rect 199222 534858 199306 535094
rect 199542 534858 236186 535094
rect 236422 534858 236506 535094
rect 236742 534858 273386 535094
rect 273622 534858 273706 535094
rect 273942 534858 310586 535094
rect 310822 534858 310906 535094
rect 311142 534858 347786 535094
rect 348022 534858 348106 535094
rect 348342 534858 384986 535094
rect 385222 534858 385306 535094
rect 385542 534858 422186 535094
rect 422422 534858 422506 535094
rect 422742 534858 459386 535094
rect 459622 534858 459706 535094
rect 459942 534858 496586 535094
rect 496822 534858 496906 535094
rect 497142 534858 533786 535094
rect 534022 534858 534106 535094
rect 534342 534858 570986 535094
rect 571222 534858 571306 535094
rect 571542 534858 582820 535094
rect 1104 534826 582820 534858
rect 1104 531694 582820 531726
rect 1104 531458 9266 531694
rect 9502 531458 9586 531694
rect 9822 531458 46466 531694
rect 46702 531458 46786 531694
rect 47022 531458 83666 531694
rect 83902 531458 83986 531694
rect 84222 531458 120866 531694
rect 121102 531458 121186 531694
rect 121422 531458 158066 531694
rect 158302 531458 158386 531694
rect 158622 531458 195266 531694
rect 195502 531458 195586 531694
rect 195822 531458 232466 531694
rect 232702 531458 232786 531694
rect 233022 531458 269666 531694
rect 269902 531458 269986 531694
rect 270222 531458 306866 531694
rect 307102 531458 307186 531694
rect 307422 531458 344066 531694
rect 344302 531458 344386 531694
rect 344622 531458 381266 531694
rect 381502 531458 381586 531694
rect 381822 531458 418466 531694
rect 418702 531458 418786 531694
rect 419022 531458 455666 531694
rect 455902 531458 455986 531694
rect 456222 531458 492866 531694
rect 493102 531458 493186 531694
rect 493422 531458 530066 531694
rect 530302 531458 530386 531694
rect 530622 531458 567266 531694
rect 567502 531458 567586 531694
rect 567822 531458 582820 531694
rect 1104 531374 582820 531458
rect 1104 531138 9266 531374
rect 9502 531138 9586 531374
rect 9822 531138 46466 531374
rect 46702 531138 46786 531374
rect 47022 531138 83666 531374
rect 83902 531138 83986 531374
rect 84222 531138 120866 531374
rect 121102 531138 121186 531374
rect 121422 531138 158066 531374
rect 158302 531138 158386 531374
rect 158622 531138 195266 531374
rect 195502 531138 195586 531374
rect 195822 531138 232466 531374
rect 232702 531138 232786 531374
rect 233022 531138 269666 531374
rect 269902 531138 269986 531374
rect 270222 531138 306866 531374
rect 307102 531138 307186 531374
rect 307422 531138 344066 531374
rect 344302 531138 344386 531374
rect 344622 531138 381266 531374
rect 381502 531138 381586 531374
rect 381822 531138 418466 531374
rect 418702 531138 418786 531374
rect 419022 531138 455666 531374
rect 455902 531138 455986 531374
rect 456222 531138 492866 531374
rect 493102 531138 493186 531374
rect 493422 531138 530066 531374
rect 530302 531138 530386 531374
rect 530622 531138 567266 531374
rect 567502 531138 567586 531374
rect 567822 531138 582820 531374
rect 1104 531106 582820 531138
rect 1104 527974 582820 528006
rect 1104 527738 5546 527974
rect 5782 527738 5866 527974
rect 6102 527738 42746 527974
rect 42982 527738 43066 527974
rect 43302 527738 79946 527974
rect 80182 527738 80266 527974
rect 80502 527738 117146 527974
rect 117382 527738 117466 527974
rect 117702 527738 154346 527974
rect 154582 527738 154666 527974
rect 154902 527738 191546 527974
rect 191782 527738 191866 527974
rect 192102 527738 228746 527974
rect 228982 527738 229066 527974
rect 229302 527738 265946 527974
rect 266182 527738 266266 527974
rect 266502 527738 303146 527974
rect 303382 527738 303466 527974
rect 303702 527738 340346 527974
rect 340582 527738 340666 527974
rect 340902 527738 377546 527974
rect 377782 527738 377866 527974
rect 378102 527738 414746 527974
rect 414982 527738 415066 527974
rect 415302 527738 451946 527974
rect 452182 527738 452266 527974
rect 452502 527738 489146 527974
rect 489382 527738 489466 527974
rect 489702 527738 526346 527974
rect 526582 527738 526666 527974
rect 526902 527738 563546 527974
rect 563782 527738 563866 527974
rect 564102 527738 582820 527974
rect 1104 527654 582820 527738
rect 1104 527418 5546 527654
rect 5782 527418 5866 527654
rect 6102 527418 42746 527654
rect 42982 527418 43066 527654
rect 43302 527418 79946 527654
rect 80182 527418 80266 527654
rect 80502 527418 117146 527654
rect 117382 527418 117466 527654
rect 117702 527418 154346 527654
rect 154582 527418 154666 527654
rect 154902 527418 191546 527654
rect 191782 527418 191866 527654
rect 192102 527418 228746 527654
rect 228982 527418 229066 527654
rect 229302 527418 265946 527654
rect 266182 527418 266266 527654
rect 266502 527418 303146 527654
rect 303382 527418 303466 527654
rect 303702 527418 340346 527654
rect 340582 527418 340666 527654
rect 340902 527418 377546 527654
rect 377782 527418 377866 527654
rect 378102 527418 414746 527654
rect 414982 527418 415066 527654
rect 415302 527418 451946 527654
rect 452182 527418 452266 527654
rect 452502 527418 489146 527654
rect 489382 527418 489466 527654
rect 489702 527418 526346 527654
rect 526582 527418 526666 527654
rect 526902 527418 563546 527654
rect 563782 527418 563866 527654
rect 564102 527418 582820 527654
rect 1104 527386 582820 527418
rect 1104 524254 582820 524286
rect 1104 524018 1826 524254
rect 2062 524018 2146 524254
rect 2382 524018 39026 524254
rect 39262 524018 39346 524254
rect 39582 524018 76226 524254
rect 76462 524018 76546 524254
rect 76782 524018 113426 524254
rect 113662 524018 113746 524254
rect 113982 524018 150626 524254
rect 150862 524018 150946 524254
rect 151182 524018 187826 524254
rect 188062 524018 188146 524254
rect 188382 524018 225026 524254
rect 225262 524018 225346 524254
rect 225582 524018 262226 524254
rect 262462 524018 262546 524254
rect 262782 524018 299426 524254
rect 299662 524018 299746 524254
rect 299982 524018 336626 524254
rect 336862 524018 336946 524254
rect 337182 524018 373826 524254
rect 374062 524018 374146 524254
rect 374382 524018 411026 524254
rect 411262 524018 411346 524254
rect 411582 524018 448226 524254
rect 448462 524018 448546 524254
rect 448782 524018 485426 524254
rect 485662 524018 485746 524254
rect 485982 524018 522626 524254
rect 522862 524018 522946 524254
rect 523182 524018 559826 524254
rect 560062 524018 560146 524254
rect 560382 524018 582820 524254
rect 1104 523934 582820 524018
rect 1104 523698 1826 523934
rect 2062 523698 2146 523934
rect 2382 523698 39026 523934
rect 39262 523698 39346 523934
rect 39582 523698 76226 523934
rect 76462 523698 76546 523934
rect 76782 523698 113426 523934
rect 113662 523698 113746 523934
rect 113982 523698 150626 523934
rect 150862 523698 150946 523934
rect 151182 523698 187826 523934
rect 188062 523698 188146 523934
rect 188382 523698 225026 523934
rect 225262 523698 225346 523934
rect 225582 523698 262226 523934
rect 262462 523698 262546 523934
rect 262782 523698 299426 523934
rect 299662 523698 299746 523934
rect 299982 523698 336626 523934
rect 336862 523698 336946 523934
rect 337182 523698 373826 523934
rect 374062 523698 374146 523934
rect 374382 523698 411026 523934
rect 411262 523698 411346 523934
rect 411582 523698 448226 523934
rect 448462 523698 448546 523934
rect 448782 523698 485426 523934
rect 485662 523698 485746 523934
rect 485982 523698 522626 523934
rect 522862 523698 522946 523934
rect 523182 523698 559826 523934
rect 560062 523698 560146 523934
rect 560382 523698 582820 523934
rect 1104 523666 582820 523698
rect 1104 513094 582820 513126
rect 1104 512858 27866 513094
rect 28102 512858 28186 513094
rect 28422 512858 65066 513094
rect 65302 512858 65386 513094
rect 65622 512858 102266 513094
rect 102502 512858 102586 513094
rect 102822 512858 139466 513094
rect 139702 512858 139786 513094
rect 140022 512858 176666 513094
rect 176902 512858 176986 513094
rect 177222 512858 213866 513094
rect 214102 512858 214186 513094
rect 214422 512858 251066 513094
rect 251302 512858 251386 513094
rect 251622 512858 288266 513094
rect 288502 512858 288586 513094
rect 288822 512858 325466 513094
rect 325702 512858 325786 513094
rect 326022 512858 362666 513094
rect 362902 512858 362986 513094
rect 363222 512858 399866 513094
rect 400102 512858 400186 513094
rect 400422 512858 437066 513094
rect 437302 512858 437386 513094
rect 437622 512858 474266 513094
rect 474502 512858 474586 513094
rect 474822 512858 511466 513094
rect 511702 512858 511786 513094
rect 512022 512858 548666 513094
rect 548902 512858 548986 513094
rect 549222 512858 582820 513094
rect 1104 512774 582820 512858
rect 1104 512538 27866 512774
rect 28102 512538 28186 512774
rect 28422 512538 65066 512774
rect 65302 512538 65386 512774
rect 65622 512538 102266 512774
rect 102502 512538 102586 512774
rect 102822 512538 139466 512774
rect 139702 512538 139786 512774
rect 140022 512538 176666 512774
rect 176902 512538 176986 512774
rect 177222 512538 213866 512774
rect 214102 512538 214186 512774
rect 214422 512538 251066 512774
rect 251302 512538 251386 512774
rect 251622 512538 288266 512774
rect 288502 512538 288586 512774
rect 288822 512538 325466 512774
rect 325702 512538 325786 512774
rect 326022 512538 362666 512774
rect 362902 512538 362986 512774
rect 363222 512538 399866 512774
rect 400102 512538 400186 512774
rect 400422 512538 437066 512774
rect 437302 512538 437386 512774
rect 437622 512538 474266 512774
rect 474502 512538 474586 512774
rect 474822 512538 511466 512774
rect 511702 512538 511786 512774
rect 512022 512538 548666 512774
rect 548902 512538 548986 512774
rect 549222 512538 582820 512774
rect 1104 512506 582820 512538
rect 1104 509374 582820 509406
rect 1104 509138 24146 509374
rect 24382 509138 24466 509374
rect 24702 509138 61346 509374
rect 61582 509138 61666 509374
rect 61902 509138 98546 509374
rect 98782 509138 98866 509374
rect 99102 509138 135746 509374
rect 135982 509138 136066 509374
rect 136302 509138 172946 509374
rect 173182 509138 173266 509374
rect 173502 509138 210146 509374
rect 210382 509138 210466 509374
rect 210702 509138 247346 509374
rect 247582 509138 247666 509374
rect 247902 509138 284546 509374
rect 284782 509138 284866 509374
rect 285102 509138 321746 509374
rect 321982 509138 322066 509374
rect 322302 509138 358946 509374
rect 359182 509138 359266 509374
rect 359502 509138 396146 509374
rect 396382 509138 396466 509374
rect 396702 509138 433346 509374
rect 433582 509138 433666 509374
rect 433902 509138 470546 509374
rect 470782 509138 470866 509374
rect 471102 509138 507746 509374
rect 507982 509138 508066 509374
rect 508302 509138 544946 509374
rect 545182 509138 545266 509374
rect 545502 509138 582146 509374
rect 582382 509138 582466 509374
rect 582702 509138 582820 509374
rect 1104 509054 582820 509138
rect 1104 508818 24146 509054
rect 24382 508818 24466 509054
rect 24702 508818 61346 509054
rect 61582 508818 61666 509054
rect 61902 508818 98546 509054
rect 98782 508818 98866 509054
rect 99102 508818 135746 509054
rect 135982 508818 136066 509054
rect 136302 508818 172946 509054
rect 173182 508818 173266 509054
rect 173502 508818 210146 509054
rect 210382 508818 210466 509054
rect 210702 508818 247346 509054
rect 247582 508818 247666 509054
rect 247902 508818 284546 509054
rect 284782 508818 284866 509054
rect 285102 508818 321746 509054
rect 321982 508818 322066 509054
rect 322302 508818 358946 509054
rect 359182 508818 359266 509054
rect 359502 508818 396146 509054
rect 396382 508818 396466 509054
rect 396702 508818 433346 509054
rect 433582 508818 433666 509054
rect 433902 508818 470546 509054
rect 470782 508818 470866 509054
rect 471102 508818 507746 509054
rect 507982 508818 508066 509054
rect 508302 508818 544946 509054
rect 545182 508818 545266 509054
rect 545502 508818 582146 509054
rect 582382 508818 582466 509054
rect 582702 508818 582820 509054
rect 1104 508786 582820 508818
rect 1104 505654 582820 505686
rect 1104 505418 20426 505654
rect 20662 505418 20746 505654
rect 20982 505418 57626 505654
rect 57862 505418 57946 505654
rect 58182 505418 94826 505654
rect 95062 505418 95146 505654
rect 95382 505418 132026 505654
rect 132262 505418 132346 505654
rect 132582 505418 169226 505654
rect 169462 505418 169546 505654
rect 169782 505418 206426 505654
rect 206662 505418 206746 505654
rect 206982 505418 243626 505654
rect 243862 505418 243946 505654
rect 244182 505418 280826 505654
rect 281062 505418 281146 505654
rect 281382 505418 318026 505654
rect 318262 505418 318346 505654
rect 318582 505418 355226 505654
rect 355462 505418 355546 505654
rect 355782 505418 392426 505654
rect 392662 505418 392746 505654
rect 392982 505418 429626 505654
rect 429862 505418 429946 505654
rect 430182 505418 466826 505654
rect 467062 505418 467146 505654
rect 467382 505418 504026 505654
rect 504262 505418 504346 505654
rect 504582 505418 541226 505654
rect 541462 505418 541546 505654
rect 541782 505418 578426 505654
rect 578662 505418 578746 505654
rect 578982 505418 582820 505654
rect 1104 505334 582820 505418
rect 1104 505098 20426 505334
rect 20662 505098 20746 505334
rect 20982 505098 57626 505334
rect 57862 505098 57946 505334
rect 58182 505098 94826 505334
rect 95062 505098 95146 505334
rect 95382 505098 132026 505334
rect 132262 505098 132346 505334
rect 132582 505098 169226 505334
rect 169462 505098 169546 505334
rect 169782 505098 206426 505334
rect 206662 505098 206746 505334
rect 206982 505098 243626 505334
rect 243862 505098 243946 505334
rect 244182 505098 280826 505334
rect 281062 505098 281146 505334
rect 281382 505098 318026 505334
rect 318262 505098 318346 505334
rect 318582 505098 355226 505334
rect 355462 505098 355546 505334
rect 355782 505098 392426 505334
rect 392662 505098 392746 505334
rect 392982 505098 429626 505334
rect 429862 505098 429946 505334
rect 430182 505098 466826 505334
rect 467062 505098 467146 505334
rect 467382 505098 504026 505334
rect 504262 505098 504346 505334
rect 504582 505098 541226 505334
rect 541462 505098 541546 505334
rect 541782 505098 578426 505334
rect 578662 505098 578746 505334
rect 578982 505098 582820 505334
rect 1104 505066 582820 505098
rect 1104 501934 582820 501966
rect 1104 501698 16706 501934
rect 16942 501698 17026 501934
rect 17262 501698 53906 501934
rect 54142 501698 54226 501934
rect 54462 501698 91106 501934
rect 91342 501698 91426 501934
rect 91662 501698 128306 501934
rect 128542 501698 128626 501934
rect 128862 501698 165506 501934
rect 165742 501698 165826 501934
rect 166062 501698 202706 501934
rect 202942 501698 203026 501934
rect 203262 501698 239906 501934
rect 240142 501698 240226 501934
rect 240462 501698 277106 501934
rect 277342 501698 277426 501934
rect 277662 501698 314306 501934
rect 314542 501698 314626 501934
rect 314862 501698 351506 501934
rect 351742 501698 351826 501934
rect 352062 501698 388706 501934
rect 388942 501698 389026 501934
rect 389262 501698 425906 501934
rect 426142 501698 426226 501934
rect 426462 501698 463106 501934
rect 463342 501698 463426 501934
rect 463662 501698 500306 501934
rect 500542 501698 500626 501934
rect 500862 501698 537506 501934
rect 537742 501698 537826 501934
rect 538062 501698 574706 501934
rect 574942 501698 575026 501934
rect 575262 501698 582820 501934
rect 1104 501614 582820 501698
rect 1104 501378 16706 501614
rect 16942 501378 17026 501614
rect 17262 501378 53906 501614
rect 54142 501378 54226 501614
rect 54462 501378 91106 501614
rect 91342 501378 91426 501614
rect 91662 501378 128306 501614
rect 128542 501378 128626 501614
rect 128862 501378 165506 501614
rect 165742 501378 165826 501614
rect 166062 501378 202706 501614
rect 202942 501378 203026 501614
rect 203262 501378 239906 501614
rect 240142 501378 240226 501614
rect 240462 501378 277106 501614
rect 277342 501378 277426 501614
rect 277662 501378 314306 501614
rect 314542 501378 314626 501614
rect 314862 501378 351506 501614
rect 351742 501378 351826 501614
rect 352062 501378 388706 501614
rect 388942 501378 389026 501614
rect 389262 501378 425906 501614
rect 426142 501378 426226 501614
rect 426462 501378 463106 501614
rect 463342 501378 463426 501614
rect 463662 501378 500306 501614
rect 500542 501378 500626 501614
rect 500862 501378 537506 501614
rect 537742 501378 537826 501614
rect 538062 501378 574706 501614
rect 574942 501378 575026 501614
rect 575262 501378 582820 501614
rect 1104 501346 582820 501378
rect 1104 498214 582820 498246
rect 1104 497978 12986 498214
rect 13222 497978 13306 498214
rect 13542 497978 50186 498214
rect 50422 497978 50506 498214
rect 50742 497978 87386 498214
rect 87622 497978 87706 498214
rect 87942 497978 124586 498214
rect 124822 497978 124906 498214
rect 125142 497978 161786 498214
rect 162022 497978 162106 498214
rect 162342 497978 198986 498214
rect 199222 497978 199306 498214
rect 199542 497978 236186 498214
rect 236422 497978 236506 498214
rect 236742 497978 273386 498214
rect 273622 497978 273706 498214
rect 273942 497978 310586 498214
rect 310822 497978 310906 498214
rect 311142 497978 347786 498214
rect 348022 497978 348106 498214
rect 348342 497978 384986 498214
rect 385222 497978 385306 498214
rect 385542 497978 422186 498214
rect 422422 497978 422506 498214
rect 422742 497978 459386 498214
rect 459622 497978 459706 498214
rect 459942 497978 496586 498214
rect 496822 497978 496906 498214
rect 497142 497978 533786 498214
rect 534022 497978 534106 498214
rect 534342 497978 570986 498214
rect 571222 497978 571306 498214
rect 571542 497978 582820 498214
rect 1104 497894 582820 497978
rect 1104 497658 12986 497894
rect 13222 497658 13306 497894
rect 13542 497658 50186 497894
rect 50422 497658 50506 497894
rect 50742 497658 87386 497894
rect 87622 497658 87706 497894
rect 87942 497658 124586 497894
rect 124822 497658 124906 497894
rect 125142 497658 161786 497894
rect 162022 497658 162106 497894
rect 162342 497658 198986 497894
rect 199222 497658 199306 497894
rect 199542 497658 236186 497894
rect 236422 497658 236506 497894
rect 236742 497658 273386 497894
rect 273622 497658 273706 497894
rect 273942 497658 310586 497894
rect 310822 497658 310906 497894
rect 311142 497658 347786 497894
rect 348022 497658 348106 497894
rect 348342 497658 384986 497894
rect 385222 497658 385306 497894
rect 385542 497658 422186 497894
rect 422422 497658 422506 497894
rect 422742 497658 459386 497894
rect 459622 497658 459706 497894
rect 459942 497658 496586 497894
rect 496822 497658 496906 497894
rect 497142 497658 533786 497894
rect 534022 497658 534106 497894
rect 534342 497658 570986 497894
rect 571222 497658 571306 497894
rect 571542 497658 582820 497894
rect 1104 497626 582820 497658
rect 1104 494494 582820 494526
rect 1104 494258 9266 494494
rect 9502 494258 9586 494494
rect 9822 494258 46466 494494
rect 46702 494258 46786 494494
rect 47022 494258 83666 494494
rect 83902 494258 83986 494494
rect 84222 494258 120866 494494
rect 121102 494258 121186 494494
rect 121422 494258 158066 494494
rect 158302 494258 158386 494494
rect 158622 494258 195266 494494
rect 195502 494258 195586 494494
rect 195822 494258 232466 494494
rect 232702 494258 232786 494494
rect 233022 494258 269666 494494
rect 269902 494258 269986 494494
rect 270222 494258 306866 494494
rect 307102 494258 307186 494494
rect 307422 494258 344066 494494
rect 344302 494258 344386 494494
rect 344622 494258 381266 494494
rect 381502 494258 381586 494494
rect 381822 494258 418466 494494
rect 418702 494258 418786 494494
rect 419022 494258 455666 494494
rect 455902 494258 455986 494494
rect 456222 494258 492866 494494
rect 493102 494258 493186 494494
rect 493422 494258 530066 494494
rect 530302 494258 530386 494494
rect 530622 494258 567266 494494
rect 567502 494258 567586 494494
rect 567822 494258 582820 494494
rect 1104 494174 582820 494258
rect 1104 493938 9266 494174
rect 9502 493938 9586 494174
rect 9822 493938 46466 494174
rect 46702 493938 46786 494174
rect 47022 493938 83666 494174
rect 83902 493938 83986 494174
rect 84222 493938 120866 494174
rect 121102 493938 121186 494174
rect 121422 493938 158066 494174
rect 158302 493938 158386 494174
rect 158622 493938 195266 494174
rect 195502 493938 195586 494174
rect 195822 493938 232466 494174
rect 232702 493938 232786 494174
rect 233022 493938 269666 494174
rect 269902 493938 269986 494174
rect 270222 493938 306866 494174
rect 307102 493938 307186 494174
rect 307422 493938 344066 494174
rect 344302 493938 344386 494174
rect 344622 493938 381266 494174
rect 381502 493938 381586 494174
rect 381822 493938 418466 494174
rect 418702 493938 418786 494174
rect 419022 493938 455666 494174
rect 455902 493938 455986 494174
rect 456222 493938 492866 494174
rect 493102 493938 493186 494174
rect 493422 493938 530066 494174
rect 530302 493938 530386 494174
rect 530622 493938 567266 494174
rect 567502 493938 567586 494174
rect 567822 493938 582820 494174
rect 1104 493906 582820 493938
rect 1104 490774 582820 490806
rect 1104 490538 5546 490774
rect 5782 490538 5866 490774
rect 6102 490538 42746 490774
rect 42982 490538 43066 490774
rect 43302 490538 79946 490774
rect 80182 490538 80266 490774
rect 80502 490538 117146 490774
rect 117382 490538 117466 490774
rect 117702 490538 154346 490774
rect 154582 490538 154666 490774
rect 154902 490538 191546 490774
rect 191782 490538 191866 490774
rect 192102 490538 228746 490774
rect 228982 490538 229066 490774
rect 229302 490538 265946 490774
rect 266182 490538 266266 490774
rect 266502 490538 303146 490774
rect 303382 490538 303466 490774
rect 303702 490538 340346 490774
rect 340582 490538 340666 490774
rect 340902 490538 377546 490774
rect 377782 490538 377866 490774
rect 378102 490538 414746 490774
rect 414982 490538 415066 490774
rect 415302 490538 451946 490774
rect 452182 490538 452266 490774
rect 452502 490538 489146 490774
rect 489382 490538 489466 490774
rect 489702 490538 526346 490774
rect 526582 490538 526666 490774
rect 526902 490538 563546 490774
rect 563782 490538 563866 490774
rect 564102 490538 582820 490774
rect 1104 490454 582820 490538
rect 1104 490218 5546 490454
rect 5782 490218 5866 490454
rect 6102 490218 42746 490454
rect 42982 490218 43066 490454
rect 43302 490218 79946 490454
rect 80182 490218 80266 490454
rect 80502 490218 117146 490454
rect 117382 490218 117466 490454
rect 117702 490218 154346 490454
rect 154582 490218 154666 490454
rect 154902 490218 191546 490454
rect 191782 490218 191866 490454
rect 192102 490218 228746 490454
rect 228982 490218 229066 490454
rect 229302 490218 265946 490454
rect 266182 490218 266266 490454
rect 266502 490218 303146 490454
rect 303382 490218 303466 490454
rect 303702 490218 340346 490454
rect 340582 490218 340666 490454
rect 340902 490218 377546 490454
rect 377782 490218 377866 490454
rect 378102 490218 414746 490454
rect 414982 490218 415066 490454
rect 415302 490218 451946 490454
rect 452182 490218 452266 490454
rect 452502 490218 489146 490454
rect 489382 490218 489466 490454
rect 489702 490218 526346 490454
rect 526582 490218 526666 490454
rect 526902 490218 563546 490454
rect 563782 490218 563866 490454
rect 564102 490218 582820 490454
rect 1104 490186 582820 490218
rect 1104 487054 582820 487086
rect 1104 486818 1826 487054
rect 2062 486818 2146 487054
rect 2382 486818 39026 487054
rect 39262 486818 39346 487054
rect 39582 486818 76226 487054
rect 76462 486818 76546 487054
rect 76782 486818 113426 487054
rect 113662 486818 113746 487054
rect 113982 486818 150626 487054
rect 150862 486818 150946 487054
rect 151182 486818 187826 487054
rect 188062 486818 188146 487054
rect 188382 486818 225026 487054
rect 225262 486818 225346 487054
rect 225582 486818 262226 487054
rect 262462 486818 262546 487054
rect 262782 486818 299426 487054
rect 299662 486818 299746 487054
rect 299982 486818 336626 487054
rect 336862 486818 336946 487054
rect 337182 486818 373826 487054
rect 374062 486818 374146 487054
rect 374382 486818 411026 487054
rect 411262 486818 411346 487054
rect 411582 486818 448226 487054
rect 448462 486818 448546 487054
rect 448782 486818 485426 487054
rect 485662 486818 485746 487054
rect 485982 486818 522626 487054
rect 522862 486818 522946 487054
rect 523182 486818 559826 487054
rect 560062 486818 560146 487054
rect 560382 486818 582820 487054
rect 1104 486734 582820 486818
rect 1104 486498 1826 486734
rect 2062 486498 2146 486734
rect 2382 486498 39026 486734
rect 39262 486498 39346 486734
rect 39582 486498 76226 486734
rect 76462 486498 76546 486734
rect 76782 486498 113426 486734
rect 113662 486498 113746 486734
rect 113982 486498 150626 486734
rect 150862 486498 150946 486734
rect 151182 486498 187826 486734
rect 188062 486498 188146 486734
rect 188382 486498 225026 486734
rect 225262 486498 225346 486734
rect 225582 486498 262226 486734
rect 262462 486498 262546 486734
rect 262782 486498 299426 486734
rect 299662 486498 299746 486734
rect 299982 486498 336626 486734
rect 336862 486498 336946 486734
rect 337182 486498 373826 486734
rect 374062 486498 374146 486734
rect 374382 486498 411026 486734
rect 411262 486498 411346 486734
rect 411582 486498 448226 486734
rect 448462 486498 448546 486734
rect 448782 486498 485426 486734
rect 485662 486498 485746 486734
rect 485982 486498 522626 486734
rect 522862 486498 522946 486734
rect 523182 486498 559826 486734
rect 560062 486498 560146 486734
rect 560382 486498 582820 486734
rect 1104 486466 582820 486498
rect 1104 475894 582820 475926
rect 1104 475658 27866 475894
rect 28102 475658 28186 475894
rect 28422 475658 65066 475894
rect 65302 475658 65386 475894
rect 65622 475658 102266 475894
rect 102502 475658 102586 475894
rect 102822 475658 139466 475894
rect 139702 475658 139786 475894
rect 140022 475658 176666 475894
rect 176902 475658 176986 475894
rect 177222 475658 213866 475894
rect 214102 475658 214186 475894
rect 214422 475658 251066 475894
rect 251302 475658 251386 475894
rect 251622 475658 288266 475894
rect 288502 475658 288586 475894
rect 288822 475658 325466 475894
rect 325702 475658 325786 475894
rect 326022 475658 362666 475894
rect 362902 475658 362986 475894
rect 363222 475658 399866 475894
rect 400102 475658 400186 475894
rect 400422 475658 437066 475894
rect 437302 475658 437386 475894
rect 437622 475658 474266 475894
rect 474502 475658 474586 475894
rect 474822 475658 511466 475894
rect 511702 475658 511786 475894
rect 512022 475658 548666 475894
rect 548902 475658 548986 475894
rect 549222 475658 582820 475894
rect 1104 475574 582820 475658
rect 1104 475338 27866 475574
rect 28102 475338 28186 475574
rect 28422 475338 65066 475574
rect 65302 475338 65386 475574
rect 65622 475338 102266 475574
rect 102502 475338 102586 475574
rect 102822 475338 139466 475574
rect 139702 475338 139786 475574
rect 140022 475338 176666 475574
rect 176902 475338 176986 475574
rect 177222 475338 213866 475574
rect 214102 475338 214186 475574
rect 214422 475338 251066 475574
rect 251302 475338 251386 475574
rect 251622 475338 288266 475574
rect 288502 475338 288586 475574
rect 288822 475338 325466 475574
rect 325702 475338 325786 475574
rect 326022 475338 362666 475574
rect 362902 475338 362986 475574
rect 363222 475338 399866 475574
rect 400102 475338 400186 475574
rect 400422 475338 437066 475574
rect 437302 475338 437386 475574
rect 437622 475338 474266 475574
rect 474502 475338 474586 475574
rect 474822 475338 511466 475574
rect 511702 475338 511786 475574
rect 512022 475338 548666 475574
rect 548902 475338 548986 475574
rect 549222 475338 582820 475574
rect 1104 475306 582820 475338
rect 1104 472174 582820 472206
rect 1104 471938 24146 472174
rect 24382 471938 24466 472174
rect 24702 471938 61346 472174
rect 61582 471938 61666 472174
rect 61902 471938 98546 472174
rect 98782 471938 98866 472174
rect 99102 471938 135746 472174
rect 135982 471938 136066 472174
rect 136302 471938 172946 472174
rect 173182 471938 173266 472174
rect 173502 471938 210146 472174
rect 210382 471938 210466 472174
rect 210702 471938 247346 472174
rect 247582 471938 247666 472174
rect 247902 471938 284546 472174
rect 284782 471938 284866 472174
rect 285102 471938 321746 472174
rect 321982 471938 322066 472174
rect 322302 471938 358946 472174
rect 359182 471938 359266 472174
rect 359502 471938 396146 472174
rect 396382 471938 396466 472174
rect 396702 471938 433346 472174
rect 433582 471938 433666 472174
rect 433902 471938 470546 472174
rect 470782 471938 470866 472174
rect 471102 471938 507746 472174
rect 507982 471938 508066 472174
rect 508302 471938 544946 472174
rect 545182 471938 545266 472174
rect 545502 471938 582146 472174
rect 582382 471938 582466 472174
rect 582702 471938 582820 472174
rect 1104 471854 582820 471938
rect 1104 471618 24146 471854
rect 24382 471618 24466 471854
rect 24702 471618 61346 471854
rect 61582 471618 61666 471854
rect 61902 471618 98546 471854
rect 98782 471618 98866 471854
rect 99102 471618 135746 471854
rect 135982 471618 136066 471854
rect 136302 471618 172946 471854
rect 173182 471618 173266 471854
rect 173502 471618 210146 471854
rect 210382 471618 210466 471854
rect 210702 471618 247346 471854
rect 247582 471618 247666 471854
rect 247902 471618 284546 471854
rect 284782 471618 284866 471854
rect 285102 471618 321746 471854
rect 321982 471618 322066 471854
rect 322302 471618 358946 471854
rect 359182 471618 359266 471854
rect 359502 471618 396146 471854
rect 396382 471618 396466 471854
rect 396702 471618 433346 471854
rect 433582 471618 433666 471854
rect 433902 471618 470546 471854
rect 470782 471618 470866 471854
rect 471102 471618 507746 471854
rect 507982 471618 508066 471854
rect 508302 471618 544946 471854
rect 545182 471618 545266 471854
rect 545502 471618 582146 471854
rect 582382 471618 582466 471854
rect 582702 471618 582820 471854
rect 1104 471586 582820 471618
rect 1104 468454 582820 468486
rect 1104 468218 20426 468454
rect 20662 468218 20746 468454
rect 20982 468218 57626 468454
rect 57862 468218 57946 468454
rect 58182 468218 94826 468454
rect 95062 468218 95146 468454
rect 95382 468218 132026 468454
rect 132262 468218 132346 468454
rect 132582 468218 169226 468454
rect 169462 468218 169546 468454
rect 169782 468218 206426 468454
rect 206662 468218 206746 468454
rect 206982 468218 243626 468454
rect 243862 468218 243946 468454
rect 244182 468218 280826 468454
rect 281062 468218 281146 468454
rect 281382 468218 318026 468454
rect 318262 468218 318346 468454
rect 318582 468218 355226 468454
rect 355462 468218 355546 468454
rect 355782 468218 392426 468454
rect 392662 468218 392746 468454
rect 392982 468218 429626 468454
rect 429862 468218 429946 468454
rect 430182 468218 466826 468454
rect 467062 468218 467146 468454
rect 467382 468218 504026 468454
rect 504262 468218 504346 468454
rect 504582 468218 541226 468454
rect 541462 468218 541546 468454
rect 541782 468218 578426 468454
rect 578662 468218 578746 468454
rect 578982 468218 582820 468454
rect 1104 468134 582820 468218
rect 1104 467898 20426 468134
rect 20662 467898 20746 468134
rect 20982 467898 57626 468134
rect 57862 467898 57946 468134
rect 58182 467898 94826 468134
rect 95062 467898 95146 468134
rect 95382 467898 132026 468134
rect 132262 467898 132346 468134
rect 132582 467898 169226 468134
rect 169462 467898 169546 468134
rect 169782 467898 206426 468134
rect 206662 467898 206746 468134
rect 206982 467898 243626 468134
rect 243862 467898 243946 468134
rect 244182 467898 280826 468134
rect 281062 467898 281146 468134
rect 281382 467898 318026 468134
rect 318262 467898 318346 468134
rect 318582 467898 355226 468134
rect 355462 467898 355546 468134
rect 355782 467898 392426 468134
rect 392662 467898 392746 468134
rect 392982 467898 429626 468134
rect 429862 467898 429946 468134
rect 430182 467898 466826 468134
rect 467062 467898 467146 468134
rect 467382 467898 504026 468134
rect 504262 467898 504346 468134
rect 504582 467898 541226 468134
rect 541462 467898 541546 468134
rect 541782 467898 578426 468134
rect 578662 467898 578746 468134
rect 578982 467898 582820 468134
rect 1104 467866 582820 467898
rect 1104 464734 582820 464766
rect 1104 464498 16706 464734
rect 16942 464498 17026 464734
rect 17262 464498 53906 464734
rect 54142 464498 54226 464734
rect 54462 464498 91106 464734
rect 91342 464498 91426 464734
rect 91662 464498 128306 464734
rect 128542 464498 128626 464734
rect 128862 464498 165506 464734
rect 165742 464498 165826 464734
rect 166062 464498 202706 464734
rect 202942 464498 203026 464734
rect 203262 464498 239906 464734
rect 240142 464498 240226 464734
rect 240462 464498 277106 464734
rect 277342 464498 277426 464734
rect 277662 464498 314306 464734
rect 314542 464498 314626 464734
rect 314862 464498 351506 464734
rect 351742 464498 351826 464734
rect 352062 464498 388706 464734
rect 388942 464498 389026 464734
rect 389262 464498 425906 464734
rect 426142 464498 426226 464734
rect 426462 464498 463106 464734
rect 463342 464498 463426 464734
rect 463662 464498 500306 464734
rect 500542 464498 500626 464734
rect 500862 464498 537506 464734
rect 537742 464498 537826 464734
rect 538062 464498 574706 464734
rect 574942 464498 575026 464734
rect 575262 464498 582820 464734
rect 1104 464414 582820 464498
rect 1104 464178 16706 464414
rect 16942 464178 17026 464414
rect 17262 464178 53906 464414
rect 54142 464178 54226 464414
rect 54462 464178 91106 464414
rect 91342 464178 91426 464414
rect 91662 464178 128306 464414
rect 128542 464178 128626 464414
rect 128862 464178 165506 464414
rect 165742 464178 165826 464414
rect 166062 464178 202706 464414
rect 202942 464178 203026 464414
rect 203262 464178 239906 464414
rect 240142 464178 240226 464414
rect 240462 464178 277106 464414
rect 277342 464178 277426 464414
rect 277662 464178 314306 464414
rect 314542 464178 314626 464414
rect 314862 464178 351506 464414
rect 351742 464178 351826 464414
rect 352062 464178 388706 464414
rect 388942 464178 389026 464414
rect 389262 464178 425906 464414
rect 426142 464178 426226 464414
rect 426462 464178 463106 464414
rect 463342 464178 463426 464414
rect 463662 464178 500306 464414
rect 500542 464178 500626 464414
rect 500862 464178 537506 464414
rect 537742 464178 537826 464414
rect 538062 464178 574706 464414
rect 574942 464178 575026 464414
rect 575262 464178 582820 464414
rect 1104 464146 582820 464178
rect 1104 461014 582820 461046
rect 1104 460778 12986 461014
rect 13222 460778 13306 461014
rect 13542 460778 50186 461014
rect 50422 460778 50506 461014
rect 50742 460778 87386 461014
rect 87622 460778 87706 461014
rect 87942 460778 124586 461014
rect 124822 460778 124906 461014
rect 125142 460778 161786 461014
rect 162022 460778 162106 461014
rect 162342 460778 198986 461014
rect 199222 460778 199306 461014
rect 199542 460778 236186 461014
rect 236422 460778 236506 461014
rect 236742 460778 273386 461014
rect 273622 460778 273706 461014
rect 273942 460778 310586 461014
rect 310822 460778 310906 461014
rect 311142 460778 347786 461014
rect 348022 460778 348106 461014
rect 348342 460778 384986 461014
rect 385222 460778 385306 461014
rect 385542 460778 422186 461014
rect 422422 460778 422506 461014
rect 422742 460778 459386 461014
rect 459622 460778 459706 461014
rect 459942 460778 496586 461014
rect 496822 460778 496906 461014
rect 497142 460778 533786 461014
rect 534022 460778 534106 461014
rect 534342 460778 570986 461014
rect 571222 460778 571306 461014
rect 571542 460778 582820 461014
rect 1104 460694 582820 460778
rect 1104 460458 12986 460694
rect 13222 460458 13306 460694
rect 13542 460458 50186 460694
rect 50422 460458 50506 460694
rect 50742 460458 87386 460694
rect 87622 460458 87706 460694
rect 87942 460458 124586 460694
rect 124822 460458 124906 460694
rect 125142 460458 161786 460694
rect 162022 460458 162106 460694
rect 162342 460458 198986 460694
rect 199222 460458 199306 460694
rect 199542 460458 236186 460694
rect 236422 460458 236506 460694
rect 236742 460458 273386 460694
rect 273622 460458 273706 460694
rect 273942 460458 310586 460694
rect 310822 460458 310906 460694
rect 311142 460458 347786 460694
rect 348022 460458 348106 460694
rect 348342 460458 384986 460694
rect 385222 460458 385306 460694
rect 385542 460458 422186 460694
rect 422422 460458 422506 460694
rect 422742 460458 459386 460694
rect 459622 460458 459706 460694
rect 459942 460458 496586 460694
rect 496822 460458 496906 460694
rect 497142 460458 533786 460694
rect 534022 460458 534106 460694
rect 534342 460458 570986 460694
rect 571222 460458 571306 460694
rect 571542 460458 582820 460694
rect 1104 460426 582820 460458
rect 1104 457294 582820 457326
rect 1104 457058 9266 457294
rect 9502 457058 9586 457294
rect 9822 457058 46466 457294
rect 46702 457058 46786 457294
rect 47022 457058 83666 457294
rect 83902 457058 83986 457294
rect 84222 457058 120866 457294
rect 121102 457058 121186 457294
rect 121422 457058 158066 457294
rect 158302 457058 158386 457294
rect 158622 457058 195266 457294
rect 195502 457058 195586 457294
rect 195822 457058 232466 457294
rect 232702 457058 232786 457294
rect 233022 457058 269666 457294
rect 269902 457058 269986 457294
rect 270222 457058 306866 457294
rect 307102 457058 307186 457294
rect 307422 457058 344066 457294
rect 344302 457058 344386 457294
rect 344622 457058 381266 457294
rect 381502 457058 381586 457294
rect 381822 457058 418466 457294
rect 418702 457058 418786 457294
rect 419022 457058 455666 457294
rect 455902 457058 455986 457294
rect 456222 457058 492866 457294
rect 493102 457058 493186 457294
rect 493422 457058 530066 457294
rect 530302 457058 530386 457294
rect 530622 457058 567266 457294
rect 567502 457058 567586 457294
rect 567822 457058 582820 457294
rect 1104 456974 582820 457058
rect 1104 456738 9266 456974
rect 9502 456738 9586 456974
rect 9822 456738 46466 456974
rect 46702 456738 46786 456974
rect 47022 456738 83666 456974
rect 83902 456738 83986 456974
rect 84222 456738 120866 456974
rect 121102 456738 121186 456974
rect 121422 456738 158066 456974
rect 158302 456738 158386 456974
rect 158622 456738 195266 456974
rect 195502 456738 195586 456974
rect 195822 456738 232466 456974
rect 232702 456738 232786 456974
rect 233022 456738 269666 456974
rect 269902 456738 269986 456974
rect 270222 456738 306866 456974
rect 307102 456738 307186 456974
rect 307422 456738 344066 456974
rect 344302 456738 344386 456974
rect 344622 456738 381266 456974
rect 381502 456738 381586 456974
rect 381822 456738 418466 456974
rect 418702 456738 418786 456974
rect 419022 456738 455666 456974
rect 455902 456738 455986 456974
rect 456222 456738 492866 456974
rect 493102 456738 493186 456974
rect 493422 456738 530066 456974
rect 530302 456738 530386 456974
rect 530622 456738 567266 456974
rect 567502 456738 567586 456974
rect 567822 456738 582820 456974
rect 1104 456706 582820 456738
rect 1104 453574 582820 453606
rect 1104 453338 5546 453574
rect 5782 453338 5866 453574
rect 6102 453338 42746 453574
rect 42982 453338 43066 453574
rect 43302 453338 79946 453574
rect 80182 453338 80266 453574
rect 80502 453338 117146 453574
rect 117382 453338 117466 453574
rect 117702 453338 154346 453574
rect 154582 453338 154666 453574
rect 154902 453338 191546 453574
rect 191782 453338 191866 453574
rect 192102 453338 228746 453574
rect 228982 453338 229066 453574
rect 229302 453338 265946 453574
rect 266182 453338 266266 453574
rect 266502 453338 303146 453574
rect 303382 453338 303466 453574
rect 303702 453338 340346 453574
rect 340582 453338 340666 453574
rect 340902 453338 377546 453574
rect 377782 453338 377866 453574
rect 378102 453338 414746 453574
rect 414982 453338 415066 453574
rect 415302 453338 451946 453574
rect 452182 453338 452266 453574
rect 452502 453338 489146 453574
rect 489382 453338 489466 453574
rect 489702 453338 526346 453574
rect 526582 453338 526666 453574
rect 526902 453338 563546 453574
rect 563782 453338 563866 453574
rect 564102 453338 582820 453574
rect 1104 453254 582820 453338
rect 1104 453018 5546 453254
rect 5782 453018 5866 453254
rect 6102 453018 42746 453254
rect 42982 453018 43066 453254
rect 43302 453018 79946 453254
rect 80182 453018 80266 453254
rect 80502 453018 117146 453254
rect 117382 453018 117466 453254
rect 117702 453018 154346 453254
rect 154582 453018 154666 453254
rect 154902 453018 191546 453254
rect 191782 453018 191866 453254
rect 192102 453018 228746 453254
rect 228982 453018 229066 453254
rect 229302 453018 265946 453254
rect 266182 453018 266266 453254
rect 266502 453018 303146 453254
rect 303382 453018 303466 453254
rect 303702 453018 340346 453254
rect 340582 453018 340666 453254
rect 340902 453018 377546 453254
rect 377782 453018 377866 453254
rect 378102 453018 414746 453254
rect 414982 453018 415066 453254
rect 415302 453018 451946 453254
rect 452182 453018 452266 453254
rect 452502 453018 489146 453254
rect 489382 453018 489466 453254
rect 489702 453018 526346 453254
rect 526582 453018 526666 453254
rect 526902 453018 563546 453254
rect 563782 453018 563866 453254
rect 564102 453018 582820 453254
rect 1104 452986 582820 453018
rect 1104 449854 582820 449886
rect 1104 449618 1826 449854
rect 2062 449618 2146 449854
rect 2382 449618 39026 449854
rect 39262 449618 39346 449854
rect 39582 449618 76226 449854
rect 76462 449618 76546 449854
rect 76782 449618 113426 449854
rect 113662 449618 113746 449854
rect 113982 449618 150626 449854
rect 150862 449618 150946 449854
rect 151182 449618 187826 449854
rect 188062 449618 188146 449854
rect 188382 449618 225026 449854
rect 225262 449618 225346 449854
rect 225582 449618 262226 449854
rect 262462 449618 262546 449854
rect 262782 449618 299426 449854
rect 299662 449618 299746 449854
rect 299982 449618 336626 449854
rect 336862 449618 336946 449854
rect 337182 449618 373826 449854
rect 374062 449618 374146 449854
rect 374382 449618 411026 449854
rect 411262 449618 411346 449854
rect 411582 449618 448226 449854
rect 448462 449618 448546 449854
rect 448782 449618 485426 449854
rect 485662 449618 485746 449854
rect 485982 449618 522626 449854
rect 522862 449618 522946 449854
rect 523182 449618 559826 449854
rect 560062 449618 560146 449854
rect 560382 449618 582820 449854
rect 1104 449534 582820 449618
rect 1104 449298 1826 449534
rect 2062 449298 2146 449534
rect 2382 449298 39026 449534
rect 39262 449298 39346 449534
rect 39582 449298 76226 449534
rect 76462 449298 76546 449534
rect 76782 449298 113426 449534
rect 113662 449298 113746 449534
rect 113982 449298 150626 449534
rect 150862 449298 150946 449534
rect 151182 449298 187826 449534
rect 188062 449298 188146 449534
rect 188382 449298 225026 449534
rect 225262 449298 225346 449534
rect 225582 449298 262226 449534
rect 262462 449298 262546 449534
rect 262782 449298 299426 449534
rect 299662 449298 299746 449534
rect 299982 449298 336626 449534
rect 336862 449298 336946 449534
rect 337182 449298 373826 449534
rect 374062 449298 374146 449534
rect 374382 449298 411026 449534
rect 411262 449298 411346 449534
rect 411582 449298 448226 449534
rect 448462 449298 448546 449534
rect 448782 449298 485426 449534
rect 485662 449298 485746 449534
rect 485982 449298 522626 449534
rect 522862 449298 522946 449534
rect 523182 449298 559826 449534
rect 560062 449298 560146 449534
rect 560382 449298 582820 449534
rect 1104 449266 582820 449298
rect 1104 438694 582820 438726
rect 1104 438458 27866 438694
rect 28102 438458 28186 438694
rect 28422 438458 65066 438694
rect 65302 438458 65386 438694
rect 65622 438458 102266 438694
rect 102502 438458 102586 438694
rect 102822 438458 139466 438694
rect 139702 438458 139786 438694
rect 140022 438458 176666 438694
rect 176902 438458 176986 438694
rect 177222 438458 213866 438694
rect 214102 438458 214186 438694
rect 214422 438458 251066 438694
rect 251302 438458 251386 438694
rect 251622 438458 288266 438694
rect 288502 438458 288586 438694
rect 288822 438458 325466 438694
rect 325702 438458 325786 438694
rect 326022 438458 362666 438694
rect 362902 438458 362986 438694
rect 363222 438458 399866 438694
rect 400102 438458 400186 438694
rect 400422 438458 437066 438694
rect 437302 438458 437386 438694
rect 437622 438458 474266 438694
rect 474502 438458 474586 438694
rect 474822 438458 511466 438694
rect 511702 438458 511786 438694
rect 512022 438458 548666 438694
rect 548902 438458 548986 438694
rect 549222 438458 582820 438694
rect 1104 438374 582820 438458
rect 1104 438138 27866 438374
rect 28102 438138 28186 438374
rect 28422 438138 65066 438374
rect 65302 438138 65386 438374
rect 65622 438138 102266 438374
rect 102502 438138 102586 438374
rect 102822 438138 139466 438374
rect 139702 438138 139786 438374
rect 140022 438138 176666 438374
rect 176902 438138 176986 438374
rect 177222 438138 213866 438374
rect 214102 438138 214186 438374
rect 214422 438138 251066 438374
rect 251302 438138 251386 438374
rect 251622 438138 288266 438374
rect 288502 438138 288586 438374
rect 288822 438138 325466 438374
rect 325702 438138 325786 438374
rect 326022 438138 362666 438374
rect 362902 438138 362986 438374
rect 363222 438138 399866 438374
rect 400102 438138 400186 438374
rect 400422 438138 437066 438374
rect 437302 438138 437386 438374
rect 437622 438138 474266 438374
rect 474502 438138 474586 438374
rect 474822 438138 511466 438374
rect 511702 438138 511786 438374
rect 512022 438138 548666 438374
rect 548902 438138 548986 438374
rect 549222 438138 582820 438374
rect 1104 438106 582820 438138
rect 1104 434974 582820 435006
rect 1104 434738 24146 434974
rect 24382 434738 24466 434974
rect 24702 434738 61346 434974
rect 61582 434738 61666 434974
rect 61902 434738 98546 434974
rect 98782 434738 98866 434974
rect 99102 434738 135746 434974
rect 135982 434738 136066 434974
rect 136302 434738 172946 434974
rect 173182 434738 173266 434974
rect 173502 434738 210146 434974
rect 210382 434738 210466 434974
rect 210702 434738 247346 434974
rect 247582 434738 247666 434974
rect 247902 434738 284546 434974
rect 284782 434738 284866 434974
rect 285102 434738 321746 434974
rect 321982 434738 322066 434974
rect 322302 434738 358946 434974
rect 359182 434738 359266 434974
rect 359502 434738 396146 434974
rect 396382 434738 396466 434974
rect 396702 434738 433346 434974
rect 433582 434738 433666 434974
rect 433902 434738 470546 434974
rect 470782 434738 470866 434974
rect 471102 434738 507746 434974
rect 507982 434738 508066 434974
rect 508302 434738 544946 434974
rect 545182 434738 545266 434974
rect 545502 434738 582146 434974
rect 582382 434738 582466 434974
rect 582702 434738 582820 434974
rect 1104 434654 582820 434738
rect 1104 434418 24146 434654
rect 24382 434418 24466 434654
rect 24702 434418 61346 434654
rect 61582 434418 61666 434654
rect 61902 434418 98546 434654
rect 98782 434418 98866 434654
rect 99102 434418 135746 434654
rect 135982 434418 136066 434654
rect 136302 434418 172946 434654
rect 173182 434418 173266 434654
rect 173502 434418 210146 434654
rect 210382 434418 210466 434654
rect 210702 434418 247346 434654
rect 247582 434418 247666 434654
rect 247902 434418 284546 434654
rect 284782 434418 284866 434654
rect 285102 434418 321746 434654
rect 321982 434418 322066 434654
rect 322302 434418 358946 434654
rect 359182 434418 359266 434654
rect 359502 434418 396146 434654
rect 396382 434418 396466 434654
rect 396702 434418 433346 434654
rect 433582 434418 433666 434654
rect 433902 434418 470546 434654
rect 470782 434418 470866 434654
rect 471102 434418 507746 434654
rect 507982 434418 508066 434654
rect 508302 434418 544946 434654
rect 545182 434418 545266 434654
rect 545502 434418 582146 434654
rect 582382 434418 582466 434654
rect 582702 434418 582820 434654
rect 1104 434386 582820 434418
rect 1104 431254 582820 431286
rect 1104 431018 20426 431254
rect 20662 431018 20746 431254
rect 20982 431018 57626 431254
rect 57862 431018 57946 431254
rect 58182 431018 94826 431254
rect 95062 431018 95146 431254
rect 95382 431018 132026 431254
rect 132262 431018 132346 431254
rect 132582 431018 169226 431254
rect 169462 431018 169546 431254
rect 169782 431018 206426 431254
rect 206662 431018 206746 431254
rect 206982 431018 243626 431254
rect 243862 431018 243946 431254
rect 244182 431018 280826 431254
rect 281062 431018 281146 431254
rect 281382 431018 318026 431254
rect 318262 431018 318346 431254
rect 318582 431018 355226 431254
rect 355462 431018 355546 431254
rect 355782 431018 392426 431254
rect 392662 431018 392746 431254
rect 392982 431018 429626 431254
rect 429862 431018 429946 431254
rect 430182 431018 466826 431254
rect 467062 431018 467146 431254
rect 467382 431018 504026 431254
rect 504262 431018 504346 431254
rect 504582 431018 541226 431254
rect 541462 431018 541546 431254
rect 541782 431018 578426 431254
rect 578662 431018 578746 431254
rect 578982 431018 582820 431254
rect 1104 430934 582820 431018
rect 1104 430698 20426 430934
rect 20662 430698 20746 430934
rect 20982 430698 57626 430934
rect 57862 430698 57946 430934
rect 58182 430698 94826 430934
rect 95062 430698 95146 430934
rect 95382 430698 132026 430934
rect 132262 430698 132346 430934
rect 132582 430698 169226 430934
rect 169462 430698 169546 430934
rect 169782 430698 206426 430934
rect 206662 430698 206746 430934
rect 206982 430698 243626 430934
rect 243862 430698 243946 430934
rect 244182 430698 280826 430934
rect 281062 430698 281146 430934
rect 281382 430698 318026 430934
rect 318262 430698 318346 430934
rect 318582 430698 355226 430934
rect 355462 430698 355546 430934
rect 355782 430698 392426 430934
rect 392662 430698 392746 430934
rect 392982 430698 429626 430934
rect 429862 430698 429946 430934
rect 430182 430698 466826 430934
rect 467062 430698 467146 430934
rect 467382 430698 504026 430934
rect 504262 430698 504346 430934
rect 504582 430698 541226 430934
rect 541462 430698 541546 430934
rect 541782 430698 578426 430934
rect 578662 430698 578746 430934
rect 578982 430698 582820 430934
rect 1104 430666 582820 430698
rect 1104 427534 582820 427566
rect 1104 427298 16706 427534
rect 16942 427298 17026 427534
rect 17262 427298 53906 427534
rect 54142 427298 54226 427534
rect 54462 427298 91106 427534
rect 91342 427298 91426 427534
rect 91662 427298 128306 427534
rect 128542 427298 128626 427534
rect 128862 427298 165506 427534
rect 165742 427298 165826 427534
rect 166062 427298 202706 427534
rect 202942 427298 203026 427534
rect 203262 427298 239906 427534
rect 240142 427298 240226 427534
rect 240462 427298 277106 427534
rect 277342 427298 277426 427534
rect 277662 427298 314306 427534
rect 314542 427298 314626 427534
rect 314862 427298 351506 427534
rect 351742 427298 351826 427534
rect 352062 427298 388706 427534
rect 388942 427298 389026 427534
rect 389262 427298 425906 427534
rect 426142 427298 426226 427534
rect 426462 427298 463106 427534
rect 463342 427298 463426 427534
rect 463662 427298 500306 427534
rect 500542 427298 500626 427534
rect 500862 427298 537506 427534
rect 537742 427298 537826 427534
rect 538062 427298 574706 427534
rect 574942 427298 575026 427534
rect 575262 427298 582820 427534
rect 1104 427214 582820 427298
rect 1104 426978 16706 427214
rect 16942 426978 17026 427214
rect 17262 426978 53906 427214
rect 54142 426978 54226 427214
rect 54462 426978 91106 427214
rect 91342 426978 91426 427214
rect 91662 426978 128306 427214
rect 128542 426978 128626 427214
rect 128862 426978 165506 427214
rect 165742 426978 165826 427214
rect 166062 426978 202706 427214
rect 202942 426978 203026 427214
rect 203262 426978 239906 427214
rect 240142 426978 240226 427214
rect 240462 426978 277106 427214
rect 277342 426978 277426 427214
rect 277662 426978 314306 427214
rect 314542 426978 314626 427214
rect 314862 426978 351506 427214
rect 351742 426978 351826 427214
rect 352062 426978 388706 427214
rect 388942 426978 389026 427214
rect 389262 426978 425906 427214
rect 426142 426978 426226 427214
rect 426462 426978 463106 427214
rect 463342 426978 463426 427214
rect 463662 426978 500306 427214
rect 500542 426978 500626 427214
rect 500862 426978 537506 427214
rect 537742 426978 537826 427214
rect 538062 426978 574706 427214
rect 574942 426978 575026 427214
rect 575262 426978 582820 427214
rect 1104 426946 582820 426978
rect 1104 423814 582820 423846
rect 1104 423578 12986 423814
rect 13222 423578 13306 423814
rect 13542 423578 50186 423814
rect 50422 423578 50506 423814
rect 50742 423578 87386 423814
rect 87622 423578 87706 423814
rect 87942 423578 124586 423814
rect 124822 423578 124906 423814
rect 125142 423578 161786 423814
rect 162022 423578 162106 423814
rect 162342 423578 198986 423814
rect 199222 423578 199306 423814
rect 199542 423578 236186 423814
rect 236422 423578 236506 423814
rect 236742 423578 273386 423814
rect 273622 423578 273706 423814
rect 273942 423578 310586 423814
rect 310822 423578 310906 423814
rect 311142 423578 347786 423814
rect 348022 423578 348106 423814
rect 348342 423578 384986 423814
rect 385222 423578 385306 423814
rect 385542 423578 422186 423814
rect 422422 423578 422506 423814
rect 422742 423578 459386 423814
rect 459622 423578 459706 423814
rect 459942 423578 496586 423814
rect 496822 423578 496906 423814
rect 497142 423578 533786 423814
rect 534022 423578 534106 423814
rect 534342 423578 570986 423814
rect 571222 423578 571306 423814
rect 571542 423578 582820 423814
rect 1104 423494 582820 423578
rect 1104 423258 12986 423494
rect 13222 423258 13306 423494
rect 13542 423258 50186 423494
rect 50422 423258 50506 423494
rect 50742 423258 87386 423494
rect 87622 423258 87706 423494
rect 87942 423258 124586 423494
rect 124822 423258 124906 423494
rect 125142 423258 161786 423494
rect 162022 423258 162106 423494
rect 162342 423258 198986 423494
rect 199222 423258 199306 423494
rect 199542 423258 236186 423494
rect 236422 423258 236506 423494
rect 236742 423258 273386 423494
rect 273622 423258 273706 423494
rect 273942 423258 310586 423494
rect 310822 423258 310906 423494
rect 311142 423258 347786 423494
rect 348022 423258 348106 423494
rect 348342 423258 384986 423494
rect 385222 423258 385306 423494
rect 385542 423258 422186 423494
rect 422422 423258 422506 423494
rect 422742 423258 459386 423494
rect 459622 423258 459706 423494
rect 459942 423258 496586 423494
rect 496822 423258 496906 423494
rect 497142 423258 533786 423494
rect 534022 423258 534106 423494
rect 534342 423258 570986 423494
rect 571222 423258 571306 423494
rect 571542 423258 582820 423494
rect 1104 423226 582820 423258
rect 1104 420094 582820 420126
rect 1104 419858 9266 420094
rect 9502 419858 9586 420094
rect 9822 419858 46466 420094
rect 46702 419858 46786 420094
rect 47022 419858 83666 420094
rect 83902 419858 83986 420094
rect 84222 419858 120866 420094
rect 121102 419858 121186 420094
rect 121422 419858 158066 420094
rect 158302 419858 158386 420094
rect 158622 419858 195266 420094
rect 195502 419858 195586 420094
rect 195822 419858 232466 420094
rect 232702 419858 232786 420094
rect 233022 419858 269666 420094
rect 269902 419858 269986 420094
rect 270222 419858 306866 420094
rect 307102 419858 307186 420094
rect 307422 419858 344066 420094
rect 344302 419858 344386 420094
rect 344622 419858 381266 420094
rect 381502 419858 381586 420094
rect 381822 419858 418466 420094
rect 418702 419858 418786 420094
rect 419022 419858 455666 420094
rect 455902 419858 455986 420094
rect 456222 419858 492866 420094
rect 493102 419858 493186 420094
rect 493422 419858 530066 420094
rect 530302 419858 530386 420094
rect 530622 419858 567266 420094
rect 567502 419858 567586 420094
rect 567822 419858 582820 420094
rect 1104 419774 582820 419858
rect 1104 419538 9266 419774
rect 9502 419538 9586 419774
rect 9822 419538 46466 419774
rect 46702 419538 46786 419774
rect 47022 419538 83666 419774
rect 83902 419538 83986 419774
rect 84222 419538 120866 419774
rect 121102 419538 121186 419774
rect 121422 419538 158066 419774
rect 158302 419538 158386 419774
rect 158622 419538 195266 419774
rect 195502 419538 195586 419774
rect 195822 419538 232466 419774
rect 232702 419538 232786 419774
rect 233022 419538 269666 419774
rect 269902 419538 269986 419774
rect 270222 419538 306866 419774
rect 307102 419538 307186 419774
rect 307422 419538 344066 419774
rect 344302 419538 344386 419774
rect 344622 419538 381266 419774
rect 381502 419538 381586 419774
rect 381822 419538 418466 419774
rect 418702 419538 418786 419774
rect 419022 419538 455666 419774
rect 455902 419538 455986 419774
rect 456222 419538 492866 419774
rect 493102 419538 493186 419774
rect 493422 419538 530066 419774
rect 530302 419538 530386 419774
rect 530622 419538 567266 419774
rect 567502 419538 567586 419774
rect 567822 419538 582820 419774
rect 1104 419506 582820 419538
rect 1104 416374 582820 416406
rect 1104 416138 5546 416374
rect 5782 416138 5866 416374
rect 6102 416138 42746 416374
rect 42982 416138 43066 416374
rect 43302 416138 79946 416374
rect 80182 416138 80266 416374
rect 80502 416138 117146 416374
rect 117382 416138 117466 416374
rect 117702 416138 154346 416374
rect 154582 416138 154666 416374
rect 154902 416138 191546 416374
rect 191782 416138 191866 416374
rect 192102 416138 228746 416374
rect 228982 416138 229066 416374
rect 229302 416138 265946 416374
rect 266182 416138 266266 416374
rect 266502 416138 303146 416374
rect 303382 416138 303466 416374
rect 303702 416138 340346 416374
rect 340582 416138 340666 416374
rect 340902 416138 377546 416374
rect 377782 416138 377866 416374
rect 378102 416138 414746 416374
rect 414982 416138 415066 416374
rect 415302 416138 451946 416374
rect 452182 416138 452266 416374
rect 452502 416138 489146 416374
rect 489382 416138 489466 416374
rect 489702 416138 526346 416374
rect 526582 416138 526666 416374
rect 526902 416138 563546 416374
rect 563782 416138 563866 416374
rect 564102 416138 582820 416374
rect 1104 416054 582820 416138
rect 1104 415818 5546 416054
rect 5782 415818 5866 416054
rect 6102 415818 42746 416054
rect 42982 415818 43066 416054
rect 43302 415818 79946 416054
rect 80182 415818 80266 416054
rect 80502 415818 117146 416054
rect 117382 415818 117466 416054
rect 117702 415818 154346 416054
rect 154582 415818 154666 416054
rect 154902 415818 191546 416054
rect 191782 415818 191866 416054
rect 192102 415818 228746 416054
rect 228982 415818 229066 416054
rect 229302 415818 265946 416054
rect 266182 415818 266266 416054
rect 266502 415818 303146 416054
rect 303382 415818 303466 416054
rect 303702 415818 340346 416054
rect 340582 415818 340666 416054
rect 340902 415818 377546 416054
rect 377782 415818 377866 416054
rect 378102 415818 414746 416054
rect 414982 415818 415066 416054
rect 415302 415818 451946 416054
rect 452182 415818 452266 416054
rect 452502 415818 489146 416054
rect 489382 415818 489466 416054
rect 489702 415818 526346 416054
rect 526582 415818 526666 416054
rect 526902 415818 563546 416054
rect 563782 415818 563866 416054
rect 564102 415818 582820 416054
rect 1104 415786 582820 415818
rect 1104 412654 582820 412686
rect 1104 412418 1826 412654
rect 2062 412418 2146 412654
rect 2382 412418 39026 412654
rect 39262 412418 39346 412654
rect 39582 412418 76226 412654
rect 76462 412418 76546 412654
rect 76782 412418 113426 412654
rect 113662 412418 113746 412654
rect 113982 412418 150626 412654
rect 150862 412418 150946 412654
rect 151182 412418 187826 412654
rect 188062 412418 188146 412654
rect 188382 412418 225026 412654
rect 225262 412418 225346 412654
rect 225582 412418 262226 412654
rect 262462 412418 262546 412654
rect 262782 412418 299426 412654
rect 299662 412418 299746 412654
rect 299982 412418 336626 412654
rect 336862 412418 336946 412654
rect 337182 412418 373826 412654
rect 374062 412418 374146 412654
rect 374382 412418 411026 412654
rect 411262 412418 411346 412654
rect 411582 412418 448226 412654
rect 448462 412418 448546 412654
rect 448782 412418 485426 412654
rect 485662 412418 485746 412654
rect 485982 412418 522626 412654
rect 522862 412418 522946 412654
rect 523182 412418 559826 412654
rect 560062 412418 560146 412654
rect 560382 412418 582820 412654
rect 1104 412334 582820 412418
rect 1104 412098 1826 412334
rect 2062 412098 2146 412334
rect 2382 412098 39026 412334
rect 39262 412098 39346 412334
rect 39582 412098 76226 412334
rect 76462 412098 76546 412334
rect 76782 412098 113426 412334
rect 113662 412098 113746 412334
rect 113982 412098 150626 412334
rect 150862 412098 150946 412334
rect 151182 412098 187826 412334
rect 188062 412098 188146 412334
rect 188382 412098 225026 412334
rect 225262 412098 225346 412334
rect 225582 412098 262226 412334
rect 262462 412098 262546 412334
rect 262782 412098 299426 412334
rect 299662 412098 299746 412334
rect 299982 412098 336626 412334
rect 336862 412098 336946 412334
rect 337182 412098 373826 412334
rect 374062 412098 374146 412334
rect 374382 412098 411026 412334
rect 411262 412098 411346 412334
rect 411582 412098 448226 412334
rect 448462 412098 448546 412334
rect 448782 412098 485426 412334
rect 485662 412098 485746 412334
rect 485982 412098 522626 412334
rect 522862 412098 522946 412334
rect 523182 412098 559826 412334
rect 560062 412098 560146 412334
rect 560382 412098 582820 412334
rect 1104 412066 582820 412098
rect 1104 401494 582820 401526
rect 1104 401258 27866 401494
rect 28102 401258 28186 401494
rect 28422 401258 65066 401494
rect 65302 401258 65386 401494
rect 65622 401258 102266 401494
rect 102502 401258 102586 401494
rect 102822 401258 139466 401494
rect 139702 401258 139786 401494
rect 140022 401258 176666 401494
rect 176902 401258 176986 401494
rect 177222 401258 213866 401494
rect 214102 401258 214186 401494
rect 214422 401258 251066 401494
rect 251302 401258 251386 401494
rect 251622 401258 288266 401494
rect 288502 401258 288586 401494
rect 288822 401258 325466 401494
rect 325702 401258 325786 401494
rect 326022 401258 362666 401494
rect 362902 401258 362986 401494
rect 363222 401258 399866 401494
rect 400102 401258 400186 401494
rect 400422 401258 437066 401494
rect 437302 401258 437386 401494
rect 437622 401258 474266 401494
rect 474502 401258 474586 401494
rect 474822 401258 511466 401494
rect 511702 401258 511786 401494
rect 512022 401258 548666 401494
rect 548902 401258 548986 401494
rect 549222 401258 582820 401494
rect 1104 401174 582820 401258
rect 1104 400938 27866 401174
rect 28102 400938 28186 401174
rect 28422 400938 65066 401174
rect 65302 400938 65386 401174
rect 65622 400938 102266 401174
rect 102502 400938 102586 401174
rect 102822 400938 139466 401174
rect 139702 400938 139786 401174
rect 140022 400938 176666 401174
rect 176902 400938 176986 401174
rect 177222 400938 213866 401174
rect 214102 400938 214186 401174
rect 214422 400938 251066 401174
rect 251302 400938 251386 401174
rect 251622 400938 288266 401174
rect 288502 400938 288586 401174
rect 288822 400938 325466 401174
rect 325702 400938 325786 401174
rect 326022 400938 362666 401174
rect 362902 400938 362986 401174
rect 363222 400938 399866 401174
rect 400102 400938 400186 401174
rect 400422 400938 437066 401174
rect 437302 400938 437386 401174
rect 437622 400938 474266 401174
rect 474502 400938 474586 401174
rect 474822 400938 511466 401174
rect 511702 400938 511786 401174
rect 512022 400938 548666 401174
rect 548902 400938 548986 401174
rect 549222 400938 582820 401174
rect 1104 400906 582820 400938
rect 1104 397774 582820 397806
rect 1104 397538 24146 397774
rect 24382 397538 24466 397774
rect 24702 397538 61346 397774
rect 61582 397538 61666 397774
rect 61902 397538 98546 397774
rect 98782 397538 98866 397774
rect 99102 397538 135746 397774
rect 135982 397538 136066 397774
rect 136302 397538 172946 397774
rect 173182 397538 173266 397774
rect 173502 397538 210146 397774
rect 210382 397538 210466 397774
rect 210702 397538 247346 397774
rect 247582 397538 247666 397774
rect 247902 397538 284546 397774
rect 284782 397538 284866 397774
rect 285102 397538 321746 397774
rect 321982 397538 322066 397774
rect 322302 397538 358946 397774
rect 359182 397538 359266 397774
rect 359502 397538 396146 397774
rect 396382 397538 396466 397774
rect 396702 397538 433346 397774
rect 433582 397538 433666 397774
rect 433902 397538 470546 397774
rect 470782 397538 470866 397774
rect 471102 397538 507746 397774
rect 507982 397538 508066 397774
rect 508302 397538 544946 397774
rect 545182 397538 545266 397774
rect 545502 397538 582146 397774
rect 582382 397538 582466 397774
rect 582702 397538 582820 397774
rect 1104 397454 582820 397538
rect 1104 397218 24146 397454
rect 24382 397218 24466 397454
rect 24702 397218 61346 397454
rect 61582 397218 61666 397454
rect 61902 397218 98546 397454
rect 98782 397218 98866 397454
rect 99102 397218 135746 397454
rect 135982 397218 136066 397454
rect 136302 397218 172946 397454
rect 173182 397218 173266 397454
rect 173502 397218 210146 397454
rect 210382 397218 210466 397454
rect 210702 397218 247346 397454
rect 247582 397218 247666 397454
rect 247902 397218 284546 397454
rect 284782 397218 284866 397454
rect 285102 397218 321746 397454
rect 321982 397218 322066 397454
rect 322302 397218 358946 397454
rect 359182 397218 359266 397454
rect 359502 397218 396146 397454
rect 396382 397218 396466 397454
rect 396702 397218 433346 397454
rect 433582 397218 433666 397454
rect 433902 397218 470546 397454
rect 470782 397218 470866 397454
rect 471102 397218 507746 397454
rect 507982 397218 508066 397454
rect 508302 397218 544946 397454
rect 545182 397218 545266 397454
rect 545502 397218 582146 397454
rect 582382 397218 582466 397454
rect 582702 397218 582820 397454
rect 1104 397186 582820 397218
rect 1104 394054 582820 394086
rect 1104 393818 20426 394054
rect 20662 393818 20746 394054
rect 20982 393818 57626 394054
rect 57862 393818 57946 394054
rect 58182 393818 94826 394054
rect 95062 393818 95146 394054
rect 95382 393818 132026 394054
rect 132262 393818 132346 394054
rect 132582 393818 169226 394054
rect 169462 393818 169546 394054
rect 169782 393818 206426 394054
rect 206662 393818 206746 394054
rect 206982 393818 243626 394054
rect 243862 393818 243946 394054
rect 244182 393818 280826 394054
rect 281062 393818 281146 394054
rect 281382 393818 318026 394054
rect 318262 393818 318346 394054
rect 318582 393818 355226 394054
rect 355462 393818 355546 394054
rect 355782 393818 392426 394054
rect 392662 393818 392746 394054
rect 392982 393818 429626 394054
rect 429862 393818 429946 394054
rect 430182 393818 466826 394054
rect 467062 393818 467146 394054
rect 467382 393818 504026 394054
rect 504262 393818 504346 394054
rect 504582 393818 541226 394054
rect 541462 393818 541546 394054
rect 541782 393818 578426 394054
rect 578662 393818 578746 394054
rect 578982 393818 582820 394054
rect 1104 393734 582820 393818
rect 1104 393498 20426 393734
rect 20662 393498 20746 393734
rect 20982 393498 57626 393734
rect 57862 393498 57946 393734
rect 58182 393498 94826 393734
rect 95062 393498 95146 393734
rect 95382 393498 132026 393734
rect 132262 393498 132346 393734
rect 132582 393498 169226 393734
rect 169462 393498 169546 393734
rect 169782 393498 206426 393734
rect 206662 393498 206746 393734
rect 206982 393498 243626 393734
rect 243862 393498 243946 393734
rect 244182 393498 280826 393734
rect 281062 393498 281146 393734
rect 281382 393498 318026 393734
rect 318262 393498 318346 393734
rect 318582 393498 355226 393734
rect 355462 393498 355546 393734
rect 355782 393498 392426 393734
rect 392662 393498 392746 393734
rect 392982 393498 429626 393734
rect 429862 393498 429946 393734
rect 430182 393498 466826 393734
rect 467062 393498 467146 393734
rect 467382 393498 504026 393734
rect 504262 393498 504346 393734
rect 504582 393498 541226 393734
rect 541462 393498 541546 393734
rect 541782 393498 578426 393734
rect 578662 393498 578746 393734
rect 578982 393498 582820 393734
rect 1104 393466 582820 393498
rect 1104 390334 582820 390366
rect 1104 390098 16706 390334
rect 16942 390098 17026 390334
rect 17262 390098 53906 390334
rect 54142 390098 54226 390334
rect 54462 390098 91106 390334
rect 91342 390098 91426 390334
rect 91662 390098 128306 390334
rect 128542 390098 128626 390334
rect 128862 390098 165506 390334
rect 165742 390098 165826 390334
rect 166062 390098 202706 390334
rect 202942 390098 203026 390334
rect 203262 390098 239906 390334
rect 240142 390098 240226 390334
rect 240462 390098 277106 390334
rect 277342 390098 277426 390334
rect 277662 390098 314306 390334
rect 314542 390098 314626 390334
rect 314862 390098 351506 390334
rect 351742 390098 351826 390334
rect 352062 390098 388706 390334
rect 388942 390098 389026 390334
rect 389262 390098 425906 390334
rect 426142 390098 426226 390334
rect 426462 390098 463106 390334
rect 463342 390098 463426 390334
rect 463662 390098 500306 390334
rect 500542 390098 500626 390334
rect 500862 390098 537506 390334
rect 537742 390098 537826 390334
rect 538062 390098 574706 390334
rect 574942 390098 575026 390334
rect 575262 390098 582820 390334
rect 1104 390014 582820 390098
rect 1104 389778 16706 390014
rect 16942 389778 17026 390014
rect 17262 389778 53906 390014
rect 54142 389778 54226 390014
rect 54462 389778 91106 390014
rect 91342 389778 91426 390014
rect 91662 389778 128306 390014
rect 128542 389778 128626 390014
rect 128862 389778 165506 390014
rect 165742 389778 165826 390014
rect 166062 389778 202706 390014
rect 202942 389778 203026 390014
rect 203262 389778 239906 390014
rect 240142 389778 240226 390014
rect 240462 389778 277106 390014
rect 277342 389778 277426 390014
rect 277662 389778 314306 390014
rect 314542 389778 314626 390014
rect 314862 389778 351506 390014
rect 351742 389778 351826 390014
rect 352062 389778 388706 390014
rect 388942 389778 389026 390014
rect 389262 389778 425906 390014
rect 426142 389778 426226 390014
rect 426462 389778 463106 390014
rect 463342 389778 463426 390014
rect 463662 389778 500306 390014
rect 500542 389778 500626 390014
rect 500862 389778 537506 390014
rect 537742 389778 537826 390014
rect 538062 389778 574706 390014
rect 574942 389778 575026 390014
rect 575262 389778 582820 390014
rect 1104 389746 582820 389778
rect 1104 386614 582820 386646
rect 1104 386378 12986 386614
rect 13222 386378 13306 386614
rect 13542 386378 50186 386614
rect 50422 386378 50506 386614
rect 50742 386378 87386 386614
rect 87622 386378 87706 386614
rect 87942 386378 124586 386614
rect 124822 386378 124906 386614
rect 125142 386378 161786 386614
rect 162022 386378 162106 386614
rect 162342 386378 198986 386614
rect 199222 386378 199306 386614
rect 199542 386378 236186 386614
rect 236422 386378 236506 386614
rect 236742 386378 273386 386614
rect 273622 386378 273706 386614
rect 273942 386378 310586 386614
rect 310822 386378 310906 386614
rect 311142 386378 347786 386614
rect 348022 386378 348106 386614
rect 348342 386378 384986 386614
rect 385222 386378 385306 386614
rect 385542 386378 422186 386614
rect 422422 386378 422506 386614
rect 422742 386378 459386 386614
rect 459622 386378 459706 386614
rect 459942 386378 496586 386614
rect 496822 386378 496906 386614
rect 497142 386378 533786 386614
rect 534022 386378 534106 386614
rect 534342 386378 570986 386614
rect 571222 386378 571306 386614
rect 571542 386378 582820 386614
rect 1104 386294 582820 386378
rect 1104 386058 12986 386294
rect 13222 386058 13306 386294
rect 13542 386058 50186 386294
rect 50422 386058 50506 386294
rect 50742 386058 87386 386294
rect 87622 386058 87706 386294
rect 87942 386058 124586 386294
rect 124822 386058 124906 386294
rect 125142 386058 161786 386294
rect 162022 386058 162106 386294
rect 162342 386058 198986 386294
rect 199222 386058 199306 386294
rect 199542 386058 236186 386294
rect 236422 386058 236506 386294
rect 236742 386058 273386 386294
rect 273622 386058 273706 386294
rect 273942 386058 310586 386294
rect 310822 386058 310906 386294
rect 311142 386058 347786 386294
rect 348022 386058 348106 386294
rect 348342 386058 384986 386294
rect 385222 386058 385306 386294
rect 385542 386058 422186 386294
rect 422422 386058 422506 386294
rect 422742 386058 459386 386294
rect 459622 386058 459706 386294
rect 459942 386058 496586 386294
rect 496822 386058 496906 386294
rect 497142 386058 533786 386294
rect 534022 386058 534106 386294
rect 534342 386058 570986 386294
rect 571222 386058 571306 386294
rect 571542 386058 582820 386294
rect 1104 386026 582820 386058
rect 1104 382894 582820 382926
rect 1104 382658 9266 382894
rect 9502 382658 9586 382894
rect 9822 382658 46466 382894
rect 46702 382658 46786 382894
rect 47022 382658 83666 382894
rect 83902 382658 83986 382894
rect 84222 382658 120866 382894
rect 121102 382658 121186 382894
rect 121422 382658 158066 382894
rect 158302 382658 158386 382894
rect 158622 382658 195266 382894
rect 195502 382658 195586 382894
rect 195822 382658 232466 382894
rect 232702 382658 232786 382894
rect 233022 382658 269666 382894
rect 269902 382658 269986 382894
rect 270222 382658 306866 382894
rect 307102 382658 307186 382894
rect 307422 382658 344066 382894
rect 344302 382658 344386 382894
rect 344622 382658 381266 382894
rect 381502 382658 381586 382894
rect 381822 382658 418466 382894
rect 418702 382658 418786 382894
rect 419022 382658 455666 382894
rect 455902 382658 455986 382894
rect 456222 382658 492866 382894
rect 493102 382658 493186 382894
rect 493422 382658 530066 382894
rect 530302 382658 530386 382894
rect 530622 382658 567266 382894
rect 567502 382658 567586 382894
rect 567822 382658 582820 382894
rect 1104 382574 582820 382658
rect 1104 382338 9266 382574
rect 9502 382338 9586 382574
rect 9822 382338 46466 382574
rect 46702 382338 46786 382574
rect 47022 382338 83666 382574
rect 83902 382338 83986 382574
rect 84222 382338 120866 382574
rect 121102 382338 121186 382574
rect 121422 382338 158066 382574
rect 158302 382338 158386 382574
rect 158622 382338 195266 382574
rect 195502 382338 195586 382574
rect 195822 382338 232466 382574
rect 232702 382338 232786 382574
rect 233022 382338 269666 382574
rect 269902 382338 269986 382574
rect 270222 382338 306866 382574
rect 307102 382338 307186 382574
rect 307422 382338 344066 382574
rect 344302 382338 344386 382574
rect 344622 382338 381266 382574
rect 381502 382338 381586 382574
rect 381822 382338 418466 382574
rect 418702 382338 418786 382574
rect 419022 382338 455666 382574
rect 455902 382338 455986 382574
rect 456222 382338 492866 382574
rect 493102 382338 493186 382574
rect 493422 382338 530066 382574
rect 530302 382338 530386 382574
rect 530622 382338 567266 382574
rect 567502 382338 567586 382574
rect 567822 382338 582820 382574
rect 1104 382306 582820 382338
rect 1104 379174 582820 379206
rect 1104 378938 5546 379174
rect 5782 378938 5866 379174
rect 6102 378938 42746 379174
rect 42982 378938 43066 379174
rect 43302 378938 79946 379174
rect 80182 378938 80266 379174
rect 80502 378938 117146 379174
rect 117382 378938 117466 379174
rect 117702 378938 154346 379174
rect 154582 378938 154666 379174
rect 154902 378938 191546 379174
rect 191782 378938 191866 379174
rect 192102 378938 228746 379174
rect 228982 378938 229066 379174
rect 229302 378938 265946 379174
rect 266182 378938 266266 379174
rect 266502 378938 303146 379174
rect 303382 378938 303466 379174
rect 303702 378938 340346 379174
rect 340582 378938 340666 379174
rect 340902 378938 377546 379174
rect 377782 378938 377866 379174
rect 378102 378938 414746 379174
rect 414982 378938 415066 379174
rect 415302 378938 451946 379174
rect 452182 378938 452266 379174
rect 452502 378938 489146 379174
rect 489382 378938 489466 379174
rect 489702 378938 526346 379174
rect 526582 378938 526666 379174
rect 526902 378938 563546 379174
rect 563782 378938 563866 379174
rect 564102 378938 582820 379174
rect 1104 378854 582820 378938
rect 1104 378618 5546 378854
rect 5782 378618 5866 378854
rect 6102 378618 42746 378854
rect 42982 378618 43066 378854
rect 43302 378618 79946 378854
rect 80182 378618 80266 378854
rect 80502 378618 117146 378854
rect 117382 378618 117466 378854
rect 117702 378618 154346 378854
rect 154582 378618 154666 378854
rect 154902 378618 191546 378854
rect 191782 378618 191866 378854
rect 192102 378618 228746 378854
rect 228982 378618 229066 378854
rect 229302 378618 265946 378854
rect 266182 378618 266266 378854
rect 266502 378618 303146 378854
rect 303382 378618 303466 378854
rect 303702 378618 340346 378854
rect 340582 378618 340666 378854
rect 340902 378618 377546 378854
rect 377782 378618 377866 378854
rect 378102 378618 414746 378854
rect 414982 378618 415066 378854
rect 415302 378618 451946 378854
rect 452182 378618 452266 378854
rect 452502 378618 489146 378854
rect 489382 378618 489466 378854
rect 489702 378618 526346 378854
rect 526582 378618 526666 378854
rect 526902 378618 563546 378854
rect 563782 378618 563866 378854
rect 564102 378618 582820 378854
rect 1104 378586 582820 378618
rect 1104 375454 582820 375486
rect 1104 375218 1826 375454
rect 2062 375218 2146 375454
rect 2382 375218 39026 375454
rect 39262 375218 39346 375454
rect 39582 375218 76226 375454
rect 76462 375218 76546 375454
rect 76782 375218 113426 375454
rect 113662 375218 113746 375454
rect 113982 375218 150626 375454
rect 150862 375218 150946 375454
rect 151182 375218 187826 375454
rect 188062 375218 188146 375454
rect 188382 375218 225026 375454
rect 225262 375218 225346 375454
rect 225582 375218 262226 375454
rect 262462 375218 262546 375454
rect 262782 375218 299426 375454
rect 299662 375218 299746 375454
rect 299982 375218 336626 375454
rect 336862 375218 336946 375454
rect 337182 375218 373826 375454
rect 374062 375218 374146 375454
rect 374382 375218 411026 375454
rect 411262 375218 411346 375454
rect 411582 375218 448226 375454
rect 448462 375218 448546 375454
rect 448782 375218 485426 375454
rect 485662 375218 485746 375454
rect 485982 375218 522626 375454
rect 522862 375218 522946 375454
rect 523182 375218 559826 375454
rect 560062 375218 560146 375454
rect 560382 375218 582820 375454
rect 1104 375134 582820 375218
rect 1104 374898 1826 375134
rect 2062 374898 2146 375134
rect 2382 374898 39026 375134
rect 39262 374898 39346 375134
rect 39582 374898 76226 375134
rect 76462 374898 76546 375134
rect 76782 374898 113426 375134
rect 113662 374898 113746 375134
rect 113982 374898 150626 375134
rect 150862 374898 150946 375134
rect 151182 374898 187826 375134
rect 188062 374898 188146 375134
rect 188382 374898 225026 375134
rect 225262 374898 225346 375134
rect 225582 374898 262226 375134
rect 262462 374898 262546 375134
rect 262782 374898 299426 375134
rect 299662 374898 299746 375134
rect 299982 374898 336626 375134
rect 336862 374898 336946 375134
rect 337182 374898 373826 375134
rect 374062 374898 374146 375134
rect 374382 374898 411026 375134
rect 411262 374898 411346 375134
rect 411582 374898 448226 375134
rect 448462 374898 448546 375134
rect 448782 374898 485426 375134
rect 485662 374898 485746 375134
rect 485982 374898 522626 375134
rect 522862 374898 522946 375134
rect 523182 374898 559826 375134
rect 560062 374898 560146 375134
rect 560382 374898 582820 375134
rect 1104 374866 582820 374898
rect 1104 364294 582820 364326
rect 1104 364058 27866 364294
rect 28102 364058 28186 364294
rect 28422 364058 65066 364294
rect 65302 364058 65386 364294
rect 65622 364058 102266 364294
rect 102502 364058 102586 364294
rect 102822 364058 139466 364294
rect 139702 364058 139786 364294
rect 140022 364058 176666 364294
rect 176902 364058 176986 364294
rect 177222 364058 213866 364294
rect 214102 364058 214186 364294
rect 214422 364058 251066 364294
rect 251302 364058 251386 364294
rect 251622 364058 288266 364294
rect 288502 364058 288586 364294
rect 288822 364058 325466 364294
rect 325702 364058 325786 364294
rect 326022 364058 362666 364294
rect 362902 364058 362986 364294
rect 363222 364058 399866 364294
rect 400102 364058 400186 364294
rect 400422 364058 437066 364294
rect 437302 364058 437386 364294
rect 437622 364058 474266 364294
rect 474502 364058 474586 364294
rect 474822 364058 511466 364294
rect 511702 364058 511786 364294
rect 512022 364058 548666 364294
rect 548902 364058 548986 364294
rect 549222 364058 582820 364294
rect 1104 363974 582820 364058
rect 1104 363738 27866 363974
rect 28102 363738 28186 363974
rect 28422 363738 65066 363974
rect 65302 363738 65386 363974
rect 65622 363738 102266 363974
rect 102502 363738 102586 363974
rect 102822 363738 139466 363974
rect 139702 363738 139786 363974
rect 140022 363738 176666 363974
rect 176902 363738 176986 363974
rect 177222 363738 213866 363974
rect 214102 363738 214186 363974
rect 214422 363738 251066 363974
rect 251302 363738 251386 363974
rect 251622 363738 288266 363974
rect 288502 363738 288586 363974
rect 288822 363738 325466 363974
rect 325702 363738 325786 363974
rect 326022 363738 362666 363974
rect 362902 363738 362986 363974
rect 363222 363738 399866 363974
rect 400102 363738 400186 363974
rect 400422 363738 437066 363974
rect 437302 363738 437386 363974
rect 437622 363738 474266 363974
rect 474502 363738 474586 363974
rect 474822 363738 511466 363974
rect 511702 363738 511786 363974
rect 512022 363738 548666 363974
rect 548902 363738 548986 363974
rect 549222 363738 582820 363974
rect 1104 363706 582820 363738
rect 1104 360574 582820 360606
rect 1104 360338 24146 360574
rect 24382 360338 24466 360574
rect 24702 360338 61346 360574
rect 61582 360338 61666 360574
rect 61902 360338 98546 360574
rect 98782 360338 98866 360574
rect 99102 360338 135746 360574
rect 135982 360338 136066 360574
rect 136302 360338 172946 360574
rect 173182 360338 173266 360574
rect 173502 360338 210146 360574
rect 210382 360338 210466 360574
rect 210702 360338 247346 360574
rect 247582 360338 247666 360574
rect 247902 360338 284546 360574
rect 284782 360338 284866 360574
rect 285102 360338 321746 360574
rect 321982 360338 322066 360574
rect 322302 360338 358946 360574
rect 359182 360338 359266 360574
rect 359502 360338 396146 360574
rect 396382 360338 396466 360574
rect 396702 360338 433346 360574
rect 433582 360338 433666 360574
rect 433902 360338 470546 360574
rect 470782 360338 470866 360574
rect 471102 360338 507746 360574
rect 507982 360338 508066 360574
rect 508302 360338 544946 360574
rect 545182 360338 545266 360574
rect 545502 360338 582146 360574
rect 582382 360338 582466 360574
rect 582702 360338 582820 360574
rect 1104 360254 582820 360338
rect 1104 360018 24146 360254
rect 24382 360018 24466 360254
rect 24702 360018 61346 360254
rect 61582 360018 61666 360254
rect 61902 360018 98546 360254
rect 98782 360018 98866 360254
rect 99102 360018 135746 360254
rect 135982 360018 136066 360254
rect 136302 360018 172946 360254
rect 173182 360018 173266 360254
rect 173502 360018 210146 360254
rect 210382 360018 210466 360254
rect 210702 360018 247346 360254
rect 247582 360018 247666 360254
rect 247902 360018 284546 360254
rect 284782 360018 284866 360254
rect 285102 360018 321746 360254
rect 321982 360018 322066 360254
rect 322302 360018 358946 360254
rect 359182 360018 359266 360254
rect 359502 360018 396146 360254
rect 396382 360018 396466 360254
rect 396702 360018 433346 360254
rect 433582 360018 433666 360254
rect 433902 360018 470546 360254
rect 470782 360018 470866 360254
rect 471102 360018 507746 360254
rect 507982 360018 508066 360254
rect 508302 360018 544946 360254
rect 545182 360018 545266 360254
rect 545502 360018 582146 360254
rect 582382 360018 582466 360254
rect 582702 360018 582820 360254
rect 1104 359986 582820 360018
rect 1104 356854 582820 356886
rect 1104 356618 20426 356854
rect 20662 356618 20746 356854
rect 20982 356618 57626 356854
rect 57862 356618 57946 356854
rect 58182 356618 94826 356854
rect 95062 356618 95146 356854
rect 95382 356618 132026 356854
rect 132262 356618 132346 356854
rect 132582 356618 169226 356854
rect 169462 356618 169546 356854
rect 169782 356618 206426 356854
rect 206662 356618 206746 356854
rect 206982 356618 243626 356854
rect 243862 356618 243946 356854
rect 244182 356618 280826 356854
rect 281062 356618 281146 356854
rect 281382 356618 318026 356854
rect 318262 356618 318346 356854
rect 318582 356618 355226 356854
rect 355462 356618 355546 356854
rect 355782 356618 392426 356854
rect 392662 356618 392746 356854
rect 392982 356618 429626 356854
rect 429862 356618 429946 356854
rect 430182 356618 466826 356854
rect 467062 356618 467146 356854
rect 467382 356618 504026 356854
rect 504262 356618 504346 356854
rect 504582 356618 541226 356854
rect 541462 356618 541546 356854
rect 541782 356618 578426 356854
rect 578662 356618 578746 356854
rect 578982 356618 582820 356854
rect 1104 356534 582820 356618
rect 1104 356298 20426 356534
rect 20662 356298 20746 356534
rect 20982 356298 57626 356534
rect 57862 356298 57946 356534
rect 58182 356298 94826 356534
rect 95062 356298 95146 356534
rect 95382 356298 132026 356534
rect 132262 356298 132346 356534
rect 132582 356298 169226 356534
rect 169462 356298 169546 356534
rect 169782 356298 206426 356534
rect 206662 356298 206746 356534
rect 206982 356298 243626 356534
rect 243862 356298 243946 356534
rect 244182 356298 280826 356534
rect 281062 356298 281146 356534
rect 281382 356298 318026 356534
rect 318262 356298 318346 356534
rect 318582 356298 355226 356534
rect 355462 356298 355546 356534
rect 355782 356298 392426 356534
rect 392662 356298 392746 356534
rect 392982 356298 429626 356534
rect 429862 356298 429946 356534
rect 430182 356298 466826 356534
rect 467062 356298 467146 356534
rect 467382 356298 504026 356534
rect 504262 356298 504346 356534
rect 504582 356298 541226 356534
rect 541462 356298 541546 356534
rect 541782 356298 578426 356534
rect 578662 356298 578746 356534
rect 578982 356298 582820 356534
rect 1104 356266 582820 356298
rect 1104 353134 582820 353166
rect 1104 352898 16706 353134
rect 16942 352898 17026 353134
rect 17262 352898 53906 353134
rect 54142 352898 54226 353134
rect 54462 352898 91106 353134
rect 91342 352898 91426 353134
rect 91662 352898 128306 353134
rect 128542 352898 128626 353134
rect 128862 352898 165506 353134
rect 165742 352898 165826 353134
rect 166062 352898 202706 353134
rect 202942 352898 203026 353134
rect 203262 352898 239906 353134
rect 240142 352898 240226 353134
rect 240462 352898 277106 353134
rect 277342 352898 277426 353134
rect 277662 352898 314306 353134
rect 314542 352898 314626 353134
rect 314862 352898 351506 353134
rect 351742 352898 351826 353134
rect 352062 352898 388706 353134
rect 388942 352898 389026 353134
rect 389262 352898 425906 353134
rect 426142 352898 426226 353134
rect 426462 352898 463106 353134
rect 463342 352898 463426 353134
rect 463662 352898 500306 353134
rect 500542 352898 500626 353134
rect 500862 352898 537506 353134
rect 537742 352898 537826 353134
rect 538062 352898 574706 353134
rect 574942 352898 575026 353134
rect 575262 352898 582820 353134
rect 1104 352814 582820 352898
rect 1104 352578 16706 352814
rect 16942 352578 17026 352814
rect 17262 352578 53906 352814
rect 54142 352578 54226 352814
rect 54462 352578 91106 352814
rect 91342 352578 91426 352814
rect 91662 352578 128306 352814
rect 128542 352578 128626 352814
rect 128862 352578 165506 352814
rect 165742 352578 165826 352814
rect 166062 352578 202706 352814
rect 202942 352578 203026 352814
rect 203262 352578 239906 352814
rect 240142 352578 240226 352814
rect 240462 352578 277106 352814
rect 277342 352578 277426 352814
rect 277662 352578 314306 352814
rect 314542 352578 314626 352814
rect 314862 352578 351506 352814
rect 351742 352578 351826 352814
rect 352062 352578 388706 352814
rect 388942 352578 389026 352814
rect 389262 352578 425906 352814
rect 426142 352578 426226 352814
rect 426462 352578 463106 352814
rect 463342 352578 463426 352814
rect 463662 352578 500306 352814
rect 500542 352578 500626 352814
rect 500862 352578 537506 352814
rect 537742 352578 537826 352814
rect 538062 352578 574706 352814
rect 574942 352578 575026 352814
rect 575262 352578 582820 352814
rect 1104 352546 582820 352578
rect 1104 349414 582820 349446
rect 1104 349178 12986 349414
rect 13222 349178 13306 349414
rect 13542 349178 50186 349414
rect 50422 349178 50506 349414
rect 50742 349178 87386 349414
rect 87622 349178 87706 349414
rect 87942 349178 124586 349414
rect 124822 349178 124906 349414
rect 125142 349178 161786 349414
rect 162022 349178 162106 349414
rect 162342 349178 198986 349414
rect 199222 349178 199306 349414
rect 199542 349178 236186 349414
rect 236422 349178 236506 349414
rect 236742 349178 273386 349414
rect 273622 349178 273706 349414
rect 273942 349178 310586 349414
rect 310822 349178 310906 349414
rect 311142 349178 347786 349414
rect 348022 349178 348106 349414
rect 348342 349178 384986 349414
rect 385222 349178 385306 349414
rect 385542 349178 422186 349414
rect 422422 349178 422506 349414
rect 422742 349178 459386 349414
rect 459622 349178 459706 349414
rect 459942 349178 496586 349414
rect 496822 349178 496906 349414
rect 497142 349178 533786 349414
rect 534022 349178 534106 349414
rect 534342 349178 570986 349414
rect 571222 349178 571306 349414
rect 571542 349178 582820 349414
rect 1104 349094 582820 349178
rect 1104 348858 12986 349094
rect 13222 348858 13306 349094
rect 13542 348858 50186 349094
rect 50422 348858 50506 349094
rect 50742 348858 87386 349094
rect 87622 348858 87706 349094
rect 87942 348858 124586 349094
rect 124822 348858 124906 349094
rect 125142 348858 161786 349094
rect 162022 348858 162106 349094
rect 162342 348858 198986 349094
rect 199222 348858 199306 349094
rect 199542 348858 236186 349094
rect 236422 348858 236506 349094
rect 236742 348858 273386 349094
rect 273622 348858 273706 349094
rect 273942 348858 310586 349094
rect 310822 348858 310906 349094
rect 311142 348858 347786 349094
rect 348022 348858 348106 349094
rect 348342 348858 384986 349094
rect 385222 348858 385306 349094
rect 385542 348858 422186 349094
rect 422422 348858 422506 349094
rect 422742 348858 459386 349094
rect 459622 348858 459706 349094
rect 459942 348858 496586 349094
rect 496822 348858 496906 349094
rect 497142 348858 533786 349094
rect 534022 348858 534106 349094
rect 534342 348858 570986 349094
rect 571222 348858 571306 349094
rect 571542 348858 582820 349094
rect 1104 348826 582820 348858
rect 1104 345694 582820 345726
rect 1104 345458 9266 345694
rect 9502 345458 9586 345694
rect 9822 345458 46466 345694
rect 46702 345458 46786 345694
rect 47022 345458 83666 345694
rect 83902 345458 83986 345694
rect 84222 345458 120866 345694
rect 121102 345458 121186 345694
rect 121422 345458 158066 345694
rect 158302 345458 158386 345694
rect 158622 345458 195266 345694
rect 195502 345458 195586 345694
rect 195822 345458 232466 345694
rect 232702 345458 232786 345694
rect 233022 345458 269666 345694
rect 269902 345458 269986 345694
rect 270222 345458 306866 345694
rect 307102 345458 307186 345694
rect 307422 345458 344066 345694
rect 344302 345458 344386 345694
rect 344622 345458 381266 345694
rect 381502 345458 381586 345694
rect 381822 345458 418466 345694
rect 418702 345458 418786 345694
rect 419022 345458 455666 345694
rect 455902 345458 455986 345694
rect 456222 345458 492866 345694
rect 493102 345458 493186 345694
rect 493422 345458 530066 345694
rect 530302 345458 530386 345694
rect 530622 345458 567266 345694
rect 567502 345458 567586 345694
rect 567822 345458 582820 345694
rect 1104 345374 582820 345458
rect 1104 345138 9266 345374
rect 9502 345138 9586 345374
rect 9822 345138 46466 345374
rect 46702 345138 46786 345374
rect 47022 345138 83666 345374
rect 83902 345138 83986 345374
rect 84222 345138 120866 345374
rect 121102 345138 121186 345374
rect 121422 345138 158066 345374
rect 158302 345138 158386 345374
rect 158622 345138 195266 345374
rect 195502 345138 195586 345374
rect 195822 345138 232466 345374
rect 232702 345138 232786 345374
rect 233022 345138 269666 345374
rect 269902 345138 269986 345374
rect 270222 345138 306866 345374
rect 307102 345138 307186 345374
rect 307422 345138 344066 345374
rect 344302 345138 344386 345374
rect 344622 345138 381266 345374
rect 381502 345138 381586 345374
rect 381822 345138 418466 345374
rect 418702 345138 418786 345374
rect 419022 345138 455666 345374
rect 455902 345138 455986 345374
rect 456222 345138 492866 345374
rect 493102 345138 493186 345374
rect 493422 345138 530066 345374
rect 530302 345138 530386 345374
rect 530622 345138 567266 345374
rect 567502 345138 567586 345374
rect 567822 345138 582820 345374
rect 1104 345106 582820 345138
rect 1104 341974 582820 342006
rect 1104 341738 5546 341974
rect 5782 341738 5866 341974
rect 6102 341738 42746 341974
rect 42982 341738 43066 341974
rect 43302 341738 79946 341974
rect 80182 341738 80266 341974
rect 80502 341738 117146 341974
rect 117382 341738 117466 341974
rect 117702 341738 154346 341974
rect 154582 341738 154666 341974
rect 154902 341738 191546 341974
rect 191782 341738 191866 341974
rect 192102 341738 228746 341974
rect 228982 341738 229066 341974
rect 229302 341738 265946 341974
rect 266182 341738 266266 341974
rect 266502 341738 303146 341974
rect 303382 341738 303466 341974
rect 303702 341738 340346 341974
rect 340582 341738 340666 341974
rect 340902 341738 377546 341974
rect 377782 341738 377866 341974
rect 378102 341738 414746 341974
rect 414982 341738 415066 341974
rect 415302 341738 451946 341974
rect 452182 341738 452266 341974
rect 452502 341738 489146 341974
rect 489382 341738 489466 341974
rect 489702 341738 526346 341974
rect 526582 341738 526666 341974
rect 526902 341738 563546 341974
rect 563782 341738 563866 341974
rect 564102 341738 582820 341974
rect 1104 341654 582820 341738
rect 1104 341418 5546 341654
rect 5782 341418 5866 341654
rect 6102 341418 42746 341654
rect 42982 341418 43066 341654
rect 43302 341418 79946 341654
rect 80182 341418 80266 341654
rect 80502 341418 117146 341654
rect 117382 341418 117466 341654
rect 117702 341418 154346 341654
rect 154582 341418 154666 341654
rect 154902 341418 191546 341654
rect 191782 341418 191866 341654
rect 192102 341418 228746 341654
rect 228982 341418 229066 341654
rect 229302 341418 265946 341654
rect 266182 341418 266266 341654
rect 266502 341418 303146 341654
rect 303382 341418 303466 341654
rect 303702 341418 340346 341654
rect 340582 341418 340666 341654
rect 340902 341418 377546 341654
rect 377782 341418 377866 341654
rect 378102 341418 414746 341654
rect 414982 341418 415066 341654
rect 415302 341418 451946 341654
rect 452182 341418 452266 341654
rect 452502 341418 489146 341654
rect 489382 341418 489466 341654
rect 489702 341418 526346 341654
rect 526582 341418 526666 341654
rect 526902 341418 563546 341654
rect 563782 341418 563866 341654
rect 564102 341418 582820 341654
rect 1104 341386 582820 341418
rect 1104 338254 582820 338286
rect 1104 338018 1826 338254
rect 2062 338018 2146 338254
rect 2382 338018 39026 338254
rect 39262 338018 39346 338254
rect 39582 338018 76226 338254
rect 76462 338018 76546 338254
rect 76782 338018 113426 338254
rect 113662 338018 113746 338254
rect 113982 338018 150626 338254
rect 150862 338018 150946 338254
rect 151182 338018 187826 338254
rect 188062 338018 188146 338254
rect 188382 338018 225026 338254
rect 225262 338018 225346 338254
rect 225582 338018 262226 338254
rect 262462 338018 262546 338254
rect 262782 338018 299426 338254
rect 299662 338018 299746 338254
rect 299982 338018 336626 338254
rect 336862 338018 336946 338254
rect 337182 338018 373826 338254
rect 374062 338018 374146 338254
rect 374382 338018 411026 338254
rect 411262 338018 411346 338254
rect 411582 338018 448226 338254
rect 448462 338018 448546 338254
rect 448782 338018 481952 338254
rect 482188 338018 483884 338254
rect 484120 338018 485816 338254
rect 486052 338018 487748 338254
rect 487984 338018 522626 338254
rect 522862 338018 522946 338254
rect 523182 338018 559826 338254
rect 560062 338018 560146 338254
rect 560382 338018 582820 338254
rect 1104 337934 582820 338018
rect 1104 337698 1826 337934
rect 2062 337698 2146 337934
rect 2382 337698 39026 337934
rect 39262 337698 39346 337934
rect 39582 337698 76226 337934
rect 76462 337698 76546 337934
rect 76782 337698 113426 337934
rect 113662 337698 113746 337934
rect 113982 337698 150626 337934
rect 150862 337698 150946 337934
rect 151182 337698 187826 337934
rect 188062 337698 188146 337934
rect 188382 337698 225026 337934
rect 225262 337698 225346 337934
rect 225582 337698 262226 337934
rect 262462 337698 262546 337934
rect 262782 337698 299426 337934
rect 299662 337698 299746 337934
rect 299982 337698 336626 337934
rect 336862 337698 336946 337934
rect 337182 337698 373826 337934
rect 374062 337698 374146 337934
rect 374382 337698 411026 337934
rect 411262 337698 411346 337934
rect 411582 337698 448226 337934
rect 448462 337698 448546 337934
rect 448782 337698 481952 337934
rect 482188 337698 483884 337934
rect 484120 337698 485816 337934
rect 486052 337698 487748 337934
rect 487984 337698 522626 337934
rect 522862 337698 522946 337934
rect 523182 337698 559826 337934
rect 560062 337698 560146 337934
rect 560382 337698 582820 337934
rect 1104 337666 582820 337698
rect 1104 327094 582820 327126
rect 1104 326858 27866 327094
rect 28102 326858 28186 327094
rect 28422 326858 65066 327094
rect 65302 326858 65386 327094
rect 65622 326858 102266 327094
rect 102502 326858 102586 327094
rect 102822 326858 139466 327094
rect 139702 326858 139786 327094
rect 140022 326858 176666 327094
rect 176902 326858 176986 327094
rect 177222 326858 213866 327094
rect 214102 326858 214186 327094
rect 214422 326858 251066 327094
rect 251302 326858 251386 327094
rect 251622 326858 288266 327094
rect 288502 326858 288586 327094
rect 288822 326858 325466 327094
rect 325702 326858 325786 327094
rect 326022 326858 362666 327094
rect 362902 326858 362986 327094
rect 363222 326858 399866 327094
rect 400102 326858 400186 327094
rect 400422 326858 437066 327094
rect 437302 326858 437386 327094
rect 437622 326858 474266 327094
rect 474502 326858 474586 327094
rect 474822 326858 511466 327094
rect 511702 326858 511786 327094
rect 512022 326858 548666 327094
rect 548902 326858 548986 327094
rect 549222 326858 582820 327094
rect 1104 326774 582820 326858
rect 1104 326538 27866 326774
rect 28102 326538 28186 326774
rect 28422 326538 65066 326774
rect 65302 326538 65386 326774
rect 65622 326538 102266 326774
rect 102502 326538 102586 326774
rect 102822 326538 139466 326774
rect 139702 326538 139786 326774
rect 140022 326538 176666 326774
rect 176902 326538 176986 326774
rect 177222 326538 213866 326774
rect 214102 326538 214186 326774
rect 214422 326538 251066 326774
rect 251302 326538 251386 326774
rect 251622 326538 288266 326774
rect 288502 326538 288586 326774
rect 288822 326538 325466 326774
rect 325702 326538 325786 326774
rect 326022 326538 362666 326774
rect 362902 326538 362986 326774
rect 363222 326538 399866 326774
rect 400102 326538 400186 326774
rect 400422 326538 437066 326774
rect 437302 326538 437386 326774
rect 437622 326538 474266 326774
rect 474502 326538 474586 326774
rect 474822 326538 511466 326774
rect 511702 326538 511786 326774
rect 512022 326538 548666 326774
rect 548902 326538 548986 326774
rect 549222 326538 582820 326774
rect 1104 326506 582820 326538
rect 1104 323374 582820 323406
rect 1104 323138 24146 323374
rect 24382 323138 24466 323374
rect 24702 323138 61346 323374
rect 61582 323138 61666 323374
rect 61902 323138 98546 323374
rect 98782 323138 98866 323374
rect 99102 323138 135746 323374
rect 135982 323138 136066 323374
rect 136302 323138 172946 323374
rect 173182 323138 173266 323374
rect 173502 323138 210146 323374
rect 210382 323138 210466 323374
rect 210702 323138 247346 323374
rect 247582 323138 247666 323374
rect 247902 323138 284546 323374
rect 284782 323138 284866 323374
rect 285102 323138 321746 323374
rect 321982 323138 322066 323374
rect 322302 323138 358946 323374
rect 359182 323138 359266 323374
rect 359502 323138 396146 323374
rect 396382 323138 396466 323374
rect 396702 323138 433346 323374
rect 433582 323138 433666 323374
rect 433902 323138 470546 323374
rect 470782 323138 470866 323374
rect 471102 323138 507746 323374
rect 507982 323138 508066 323374
rect 508302 323138 544946 323374
rect 545182 323138 545266 323374
rect 545502 323138 582146 323374
rect 582382 323138 582466 323374
rect 582702 323138 582820 323374
rect 1104 323054 582820 323138
rect 1104 322818 24146 323054
rect 24382 322818 24466 323054
rect 24702 322818 61346 323054
rect 61582 322818 61666 323054
rect 61902 322818 98546 323054
rect 98782 322818 98866 323054
rect 99102 322818 135746 323054
rect 135982 322818 136066 323054
rect 136302 322818 172946 323054
rect 173182 322818 173266 323054
rect 173502 322818 210146 323054
rect 210382 322818 210466 323054
rect 210702 322818 247346 323054
rect 247582 322818 247666 323054
rect 247902 322818 284546 323054
rect 284782 322818 284866 323054
rect 285102 322818 321746 323054
rect 321982 322818 322066 323054
rect 322302 322818 358946 323054
rect 359182 322818 359266 323054
rect 359502 322818 396146 323054
rect 396382 322818 396466 323054
rect 396702 322818 433346 323054
rect 433582 322818 433666 323054
rect 433902 322818 470546 323054
rect 470782 322818 470866 323054
rect 471102 322818 507746 323054
rect 507982 322818 508066 323054
rect 508302 322818 544946 323054
rect 545182 322818 545266 323054
rect 545502 322818 582146 323054
rect 582382 322818 582466 323054
rect 582702 322818 582820 323054
rect 1104 322786 582820 322818
rect 1104 319654 582820 319686
rect 1104 319418 20426 319654
rect 20662 319418 20746 319654
rect 20982 319418 57626 319654
rect 57862 319418 57946 319654
rect 58182 319418 94826 319654
rect 95062 319418 95146 319654
rect 95382 319418 132026 319654
rect 132262 319418 132346 319654
rect 132582 319418 169226 319654
rect 169462 319418 169546 319654
rect 169782 319418 206426 319654
rect 206662 319418 206746 319654
rect 206982 319418 243626 319654
rect 243862 319418 243946 319654
rect 244182 319418 280826 319654
rect 281062 319418 281146 319654
rect 281382 319418 318026 319654
rect 318262 319418 318346 319654
rect 318582 319418 355226 319654
rect 355462 319418 355546 319654
rect 355782 319418 392426 319654
rect 392662 319418 392746 319654
rect 392982 319418 429626 319654
rect 429862 319418 429946 319654
rect 430182 319418 466826 319654
rect 467062 319418 467146 319654
rect 467382 319418 504026 319654
rect 504262 319418 504346 319654
rect 504582 319418 541226 319654
rect 541462 319418 541546 319654
rect 541782 319418 578426 319654
rect 578662 319418 578746 319654
rect 578982 319418 582820 319654
rect 1104 319334 582820 319418
rect 1104 319098 20426 319334
rect 20662 319098 20746 319334
rect 20982 319098 57626 319334
rect 57862 319098 57946 319334
rect 58182 319098 94826 319334
rect 95062 319098 95146 319334
rect 95382 319098 132026 319334
rect 132262 319098 132346 319334
rect 132582 319098 169226 319334
rect 169462 319098 169546 319334
rect 169782 319098 206426 319334
rect 206662 319098 206746 319334
rect 206982 319098 243626 319334
rect 243862 319098 243946 319334
rect 244182 319098 280826 319334
rect 281062 319098 281146 319334
rect 281382 319098 318026 319334
rect 318262 319098 318346 319334
rect 318582 319098 355226 319334
rect 355462 319098 355546 319334
rect 355782 319098 392426 319334
rect 392662 319098 392746 319334
rect 392982 319098 429626 319334
rect 429862 319098 429946 319334
rect 430182 319098 466826 319334
rect 467062 319098 467146 319334
rect 467382 319098 504026 319334
rect 504262 319098 504346 319334
rect 504582 319098 541226 319334
rect 541462 319098 541546 319334
rect 541782 319098 578426 319334
rect 578662 319098 578746 319334
rect 578982 319098 582820 319334
rect 1104 319066 582820 319098
rect 1104 315934 582820 315966
rect 1104 315698 16706 315934
rect 16942 315698 17026 315934
rect 17262 315698 53906 315934
rect 54142 315698 54226 315934
rect 54462 315698 91106 315934
rect 91342 315698 91426 315934
rect 91662 315698 128306 315934
rect 128542 315698 128626 315934
rect 128862 315698 165506 315934
rect 165742 315698 165826 315934
rect 166062 315698 202706 315934
rect 202942 315698 203026 315934
rect 203262 315698 239906 315934
rect 240142 315698 240226 315934
rect 240462 315698 277106 315934
rect 277342 315698 277426 315934
rect 277662 315698 314306 315934
rect 314542 315698 314626 315934
rect 314862 315698 351506 315934
rect 351742 315698 351826 315934
rect 352062 315698 388706 315934
rect 388942 315698 389026 315934
rect 389262 315698 425906 315934
rect 426142 315698 426226 315934
rect 426462 315698 463106 315934
rect 463342 315698 463426 315934
rect 463662 315698 500306 315934
rect 500542 315698 500626 315934
rect 500862 315698 537506 315934
rect 537742 315698 537826 315934
rect 538062 315698 574706 315934
rect 574942 315698 575026 315934
rect 575262 315698 582820 315934
rect 1104 315614 582820 315698
rect 1104 315378 16706 315614
rect 16942 315378 17026 315614
rect 17262 315378 53906 315614
rect 54142 315378 54226 315614
rect 54462 315378 91106 315614
rect 91342 315378 91426 315614
rect 91662 315378 128306 315614
rect 128542 315378 128626 315614
rect 128862 315378 165506 315614
rect 165742 315378 165826 315614
rect 166062 315378 202706 315614
rect 202942 315378 203026 315614
rect 203262 315378 239906 315614
rect 240142 315378 240226 315614
rect 240462 315378 277106 315614
rect 277342 315378 277426 315614
rect 277662 315378 314306 315614
rect 314542 315378 314626 315614
rect 314862 315378 351506 315614
rect 351742 315378 351826 315614
rect 352062 315378 388706 315614
rect 388942 315378 389026 315614
rect 389262 315378 425906 315614
rect 426142 315378 426226 315614
rect 426462 315378 463106 315614
rect 463342 315378 463426 315614
rect 463662 315378 500306 315614
rect 500542 315378 500626 315614
rect 500862 315378 537506 315614
rect 537742 315378 537826 315614
rect 538062 315378 574706 315614
rect 574942 315378 575026 315614
rect 575262 315378 582820 315614
rect 1104 315346 582820 315378
rect 1104 312214 582820 312246
rect 1104 311978 12986 312214
rect 13222 311978 13306 312214
rect 13542 311978 50186 312214
rect 50422 311978 50506 312214
rect 50742 311978 87386 312214
rect 87622 311978 87706 312214
rect 87942 311978 124586 312214
rect 124822 311978 124906 312214
rect 125142 311978 161786 312214
rect 162022 311978 162106 312214
rect 162342 311978 198986 312214
rect 199222 311978 199306 312214
rect 199542 311978 236186 312214
rect 236422 311978 236506 312214
rect 236742 311978 273386 312214
rect 273622 311978 273706 312214
rect 273942 311978 310586 312214
rect 310822 311978 310906 312214
rect 311142 311978 347786 312214
rect 348022 311978 348106 312214
rect 348342 311978 384986 312214
rect 385222 311978 385306 312214
rect 385542 311978 422186 312214
rect 422422 311978 422506 312214
rect 422742 311978 459386 312214
rect 459622 311978 459706 312214
rect 459942 311978 496586 312214
rect 496822 311978 496906 312214
rect 497142 311978 533786 312214
rect 534022 311978 534106 312214
rect 534342 311978 570986 312214
rect 571222 311978 571306 312214
rect 571542 311978 582820 312214
rect 1104 311894 582820 311978
rect 1104 311658 12986 311894
rect 13222 311658 13306 311894
rect 13542 311658 50186 311894
rect 50422 311658 50506 311894
rect 50742 311658 87386 311894
rect 87622 311658 87706 311894
rect 87942 311658 124586 311894
rect 124822 311658 124906 311894
rect 125142 311658 161786 311894
rect 162022 311658 162106 311894
rect 162342 311658 198986 311894
rect 199222 311658 199306 311894
rect 199542 311658 236186 311894
rect 236422 311658 236506 311894
rect 236742 311658 273386 311894
rect 273622 311658 273706 311894
rect 273942 311658 310586 311894
rect 310822 311658 310906 311894
rect 311142 311658 347786 311894
rect 348022 311658 348106 311894
rect 348342 311658 384986 311894
rect 385222 311658 385306 311894
rect 385542 311658 422186 311894
rect 422422 311658 422506 311894
rect 422742 311658 459386 311894
rect 459622 311658 459706 311894
rect 459942 311658 496586 311894
rect 496822 311658 496906 311894
rect 497142 311658 533786 311894
rect 534022 311658 534106 311894
rect 534342 311658 570986 311894
rect 571222 311658 571306 311894
rect 571542 311658 582820 311894
rect 1104 311626 582820 311658
rect 1104 308494 582820 308526
rect 1104 308258 9266 308494
rect 9502 308258 9586 308494
rect 9822 308258 46466 308494
rect 46702 308258 46786 308494
rect 47022 308258 83666 308494
rect 83902 308258 83986 308494
rect 84222 308258 120866 308494
rect 121102 308258 121186 308494
rect 121422 308258 158066 308494
rect 158302 308258 158386 308494
rect 158622 308258 195266 308494
rect 195502 308258 195586 308494
rect 195822 308258 232466 308494
rect 232702 308258 232786 308494
rect 233022 308258 269666 308494
rect 269902 308258 269986 308494
rect 270222 308258 306866 308494
rect 307102 308258 307186 308494
rect 307422 308258 344066 308494
rect 344302 308258 344386 308494
rect 344622 308258 381266 308494
rect 381502 308258 381586 308494
rect 381822 308258 418466 308494
rect 418702 308258 418786 308494
rect 419022 308258 455666 308494
rect 455902 308258 455986 308494
rect 456222 308258 492866 308494
rect 493102 308258 493186 308494
rect 493422 308258 530066 308494
rect 530302 308258 530386 308494
rect 530622 308258 567266 308494
rect 567502 308258 567586 308494
rect 567822 308258 582820 308494
rect 1104 308174 582820 308258
rect 1104 307938 9266 308174
rect 9502 307938 9586 308174
rect 9822 307938 46466 308174
rect 46702 307938 46786 308174
rect 47022 307938 83666 308174
rect 83902 307938 83986 308174
rect 84222 307938 120866 308174
rect 121102 307938 121186 308174
rect 121422 307938 158066 308174
rect 158302 307938 158386 308174
rect 158622 307938 195266 308174
rect 195502 307938 195586 308174
rect 195822 307938 232466 308174
rect 232702 307938 232786 308174
rect 233022 307938 269666 308174
rect 269902 307938 269986 308174
rect 270222 307938 306866 308174
rect 307102 307938 307186 308174
rect 307422 307938 344066 308174
rect 344302 307938 344386 308174
rect 344622 307938 381266 308174
rect 381502 307938 381586 308174
rect 381822 307938 418466 308174
rect 418702 307938 418786 308174
rect 419022 307938 455666 308174
rect 455902 307938 455986 308174
rect 456222 307938 492866 308174
rect 493102 307938 493186 308174
rect 493422 307938 530066 308174
rect 530302 307938 530386 308174
rect 530622 307938 567266 308174
rect 567502 307938 567586 308174
rect 567822 307938 582820 308174
rect 1104 307906 582820 307938
rect 1104 304774 582820 304806
rect 1104 304538 5546 304774
rect 5782 304538 5866 304774
rect 6102 304538 42746 304774
rect 42982 304538 43066 304774
rect 43302 304538 79946 304774
rect 80182 304538 80266 304774
rect 80502 304538 117146 304774
rect 117382 304538 117466 304774
rect 117702 304538 154346 304774
rect 154582 304538 154666 304774
rect 154902 304538 191546 304774
rect 191782 304538 191866 304774
rect 192102 304538 228746 304774
rect 228982 304538 229066 304774
rect 229302 304538 265946 304774
rect 266182 304538 266266 304774
rect 266502 304538 303146 304774
rect 303382 304538 303466 304774
rect 303702 304538 340346 304774
rect 340582 304538 340666 304774
rect 340902 304538 377546 304774
rect 377782 304538 377866 304774
rect 378102 304538 414746 304774
rect 414982 304538 415066 304774
rect 415302 304538 451946 304774
rect 452182 304538 452266 304774
rect 452502 304538 489146 304774
rect 489382 304538 489466 304774
rect 489702 304538 526346 304774
rect 526582 304538 526666 304774
rect 526902 304538 563546 304774
rect 563782 304538 563866 304774
rect 564102 304538 582820 304774
rect 1104 304454 582820 304538
rect 1104 304218 5546 304454
rect 5782 304218 5866 304454
rect 6102 304218 42746 304454
rect 42982 304218 43066 304454
rect 43302 304218 79946 304454
rect 80182 304218 80266 304454
rect 80502 304218 117146 304454
rect 117382 304218 117466 304454
rect 117702 304218 154346 304454
rect 154582 304218 154666 304454
rect 154902 304218 191546 304454
rect 191782 304218 191866 304454
rect 192102 304218 228746 304454
rect 228982 304218 229066 304454
rect 229302 304218 265946 304454
rect 266182 304218 266266 304454
rect 266502 304218 303146 304454
rect 303382 304218 303466 304454
rect 303702 304218 340346 304454
rect 340582 304218 340666 304454
rect 340902 304218 377546 304454
rect 377782 304218 377866 304454
rect 378102 304218 414746 304454
rect 414982 304218 415066 304454
rect 415302 304218 451946 304454
rect 452182 304218 452266 304454
rect 452502 304218 489146 304454
rect 489382 304218 489466 304454
rect 489702 304218 526346 304454
rect 526582 304218 526666 304454
rect 526902 304218 563546 304454
rect 563782 304218 563866 304454
rect 564102 304218 582820 304454
rect 1104 304186 582820 304218
rect 1104 301054 582820 301086
rect 1104 300818 1826 301054
rect 2062 300818 2146 301054
rect 2382 300818 39026 301054
rect 39262 300818 39346 301054
rect 39582 300818 76226 301054
rect 76462 300818 76546 301054
rect 76782 300818 113426 301054
rect 113662 300818 113746 301054
rect 113982 300818 150626 301054
rect 150862 300818 150946 301054
rect 151182 300818 187826 301054
rect 188062 300818 188146 301054
rect 188382 300818 225026 301054
rect 225262 300818 225346 301054
rect 225582 300818 262226 301054
rect 262462 300818 262546 301054
rect 262782 300818 299426 301054
rect 299662 300818 299746 301054
rect 299982 300818 336626 301054
rect 336862 300818 336946 301054
rect 337182 300818 373826 301054
rect 374062 300818 374146 301054
rect 374382 300818 411026 301054
rect 411262 300818 411346 301054
rect 411582 300818 448226 301054
rect 448462 300818 448546 301054
rect 448782 300818 485426 301054
rect 485662 300818 485746 301054
rect 485982 300818 522626 301054
rect 522862 300818 522946 301054
rect 523182 300818 559826 301054
rect 560062 300818 560146 301054
rect 560382 300818 582820 301054
rect 1104 300734 582820 300818
rect 1104 300498 1826 300734
rect 2062 300498 2146 300734
rect 2382 300498 39026 300734
rect 39262 300498 39346 300734
rect 39582 300498 76226 300734
rect 76462 300498 76546 300734
rect 76782 300498 113426 300734
rect 113662 300498 113746 300734
rect 113982 300498 150626 300734
rect 150862 300498 150946 300734
rect 151182 300498 187826 300734
rect 188062 300498 188146 300734
rect 188382 300498 225026 300734
rect 225262 300498 225346 300734
rect 225582 300498 262226 300734
rect 262462 300498 262546 300734
rect 262782 300498 299426 300734
rect 299662 300498 299746 300734
rect 299982 300498 336626 300734
rect 336862 300498 336946 300734
rect 337182 300498 373826 300734
rect 374062 300498 374146 300734
rect 374382 300498 411026 300734
rect 411262 300498 411346 300734
rect 411582 300498 448226 300734
rect 448462 300498 448546 300734
rect 448782 300498 485426 300734
rect 485662 300498 485746 300734
rect 485982 300498 522626 300734
rect 522862 300498 522946 300734
rect 523182 300498 559826 300734
rect 560062 300498 560146 300734
rect 560382 300498 582820 300734
rect 1104 300466 582820 300498
rect 1104 289894 582820 289926
rect 1104 289658 27866 289894
rect 28102 289658 28186 289894
rect 28422 289658 65066 289894
rect 65302 289658 65386 289894
rect 65622 289658 102266 289894
rect 102502 289658 102586 289894
rect 102822 289658 139466 289894
rect 139702 289658 139786 289894
rect 140022 289658 176666 289894
rect 176902 289658 176986 289894
rect 177222 289658 213866 289894
rect 214102 289658 214186 289894
rect 214422 289658 251066 289894
rect 251302 289658 251386 289894
rect 251622 289658 288266 289894
rect 288502 289658 288586 289894
rect 288822 289658 325466 289894
rect 325702 289658 325786 289894
rect 326022 289658 362666 289894
rect 362902 289658 362986 289894
rect 363222 289658 399866 289894
rect 400102 289658 400186 289894
rect 400422 289658 437066 289894
rect 437302 289658 437386 289894
rect 437622 289658 474266 289894
rect 474502 289658 474586 289894
rect 474822 289658 511466 289894
rect 511702 289658 511786 289894
rect 512022 289658 548666 289894
rect 548902 289658 548986 289894
rect 549222 289658 582820 289894
rect 1104 289574 582820 289658
rect 1104 289338 27866 289574
rect 28102 289338 28186 289574
rect 28422 289338 65066 289574
rect 65302 289338 65386 289574
rect 65622 289338 102266 289574
rect 102502 289338 102586 289574
rect 102822 289338 139466 289574
rect 139702 289338 139786 289574
rect 140022 289338 176666 289574
rect 176902 289338 176986 289574
rect 177222 289338 213866 289574
rect 214102 289338 214186 289574
rect 214422 289338 251066 289574
rect 251302 289338 251386 289574
rect 251622 289338 288266 289574
rect 288502 289338 288586 289574
rect 288822 289338 325466 289574
rect 325702 289338 325786 289574
rect 326022 289338 362666 289574
rect 362902 289338 362986 289574
rect 363222 289338 399866 289574
rect 400102 289338 400186 289574
rect 400422 289338 437066 289574
rect 437302 289338 437386 289574
rect 437622 289338 474266 289574
rect 474502 289338 474586 289574
rect 474822 289338 511466 289574
rect 511702 289338 511786 289574
rect 512022 289338 548666 289574
rect 548902 289338 548986 289574
rect 549222 289338 582820 289574
rect 1104 289306 582820 289338
rect 1104 286174 582820 286206
rect 1104 285938 24146 286174
rect 24382 285938 24466 286174
rect 24702 285938 61346 286174
rect 61582 285938 61666 286174
rect 61902 285938 98546 286174
rect 98782 285938 98866 286174
rect 99102 285938 135746 286174
rect 135982 285938 136066 286174
rect 136302 285938 172946 286174
rect 173182 285938 173266 286174
rect 173502 285938 210146 286174
rect 210382 285938 210466 286174
rect 210702 285938 247346 286174
rect 247582 285938 247666 286174
rect 247902 285938 284546 286174
rect 284782 285938 284866 286174
rect 285102 285938 321746 286174
rect 321982 285938 322066 286174
rect 322302 285938 358946 286174
rect 359182 285938 359266 286174
rect 359502 285938 396146 286174
rect 396382 285938 396466 286174
rect 396702 285938 433346 286174
rect 433582 285938 433666 286174
rect 433902 285938 470546 286174
rect 470782 285938 470866 286174
rect 471102 285938 507746 286174
rect 507982 285938 508066 286174
rect 508302 285938 544946 286174
rect 545182 285938 545266 286174
rect 545502 285938 582146 286174
rect 582382 285938 582466 286174
rect 582702 285938 582820 286174
rect 1104 285854 582820 285938
rect 1104 285618 24146 285854
rect 24382 285618 24466 285854
rect 24702 285618 61346 285854
rect 61582 285618 61666 285854
rect 61902 285618 98546 285854
rect 98782 285618 98866 285854
rect 99102 285618 135746 285854
rect 135982 285618 136066 285854
rect 136302 285618 172946 285854
rect 173182 285618 173266 285854
rect 173502 285618 210146 285854
rect 210382 285618 210466 285854
rect 210702 285618 247346 285854
rect 247582 285618 247666 285854
rect 247902 285618 284546 285854
rect 284782 285618 284866 285854
rect 285102 285618 321746 285854
rect 321982 285618 322066 285854
rect 322302 285618 358946 285854
rect 359182 285618 359266 285854
rect 359502 285618 396146 285854
rect 396382 285618 396466 285854
rect 396702 285618 433346 285854
rect 433582 285618 433666 285854
rect 433902 285618 470546 285854
rect 470782 285618 470866 285854
rect 471102 285618 507746 285854
rect 507982 285618 508066 285854
rect 508302 285618 544946 285854
rect 545182 285618 545266 285854
rect 545502 285618 582146 285854
rect 582382 285618 582466 285854
rect 582702 285618 582820 285854
rect 1104 285586 582820 285618
rect 1104 282454 582820 282486
rect 1104 282218 20426 282454
rect 20662 282218 20746 282454
rect 20982 282218 57626 282454
rect 57862 282218 57946 282454
rect 58182 282218 94826 282454
rect 95062 282218 95146 282454
rect 95382 282218 132026 282454
rect 132262 282218 132346 282454
rect 132582 282218 169226 282454
rect 169462 282218 169546 282454
rect 169782 282218 206426 282454
rect 206662 282218 206746 282454
rect 206982 282218 243626 282454
rect 243862 282218 243946 282454
rect 244182 282218 280826 282454
rect 281062 282218 281146 282454
rect 281382 282218 318026 282454
rect 318262 282218 318346 282454
rect 318582 282218 355226 282454
rect 355462 282218 355546 282454
rect 355782 282218 392426 282454
rect 392662 282218 392746 282454
rect 392982 282218 429626 282454
rect 429862 282218 429946 282454
rect 430182 282218 466826 282454
rect 467062 282218 467146 282454
rect 467382 282218 504026 282454
rect 504262 282218 504346 282454
rect 504582 282218 541226 282454
rect 541462 282218 541546 282454
rect 541782 282218 578426 282454
rect 578662 282218 578746 282454
rect 578982 282218 582820 282454
rect 1104 282134 582820 282218
rect 1104 281898 20426 282134
rect 20662 281898 20746 282134
rect 20982 281898 57626 282134
rect 57862 281898 57946 282134
rect 58182 281898 94826 282134
rect 95062 281898 95146 282134
rect 95382 281898 132026 282134
rect 132262 281898 132346 282134
rect 132582 281898 169226 282134
rect 169462 281898 169546 282134
rect 169782 281898 206426 282134
rect 206662 281898 206746 282134
rect 206982 281898 243626 282134
rect 243862 281898 243946 282134
rect 244182 281898 280826 282134
rect 281062 281898 281146 282134
rect 281382 281898 318026 282134
rect 318262 281898 318346 282134
rect 318582 281898 355226 282134
rect 355462 281898 355546 282134
rect 355782 281898 392426 282134
rect 392662 281898 392746 282134
rect 392982 281898 429626 282134
rect 429862 281898 429946 282134
rect 430182 281898 466826 282134
rect 467062 281898 467146 282134
rect 467382 281898 504026 282134
rect 504262 281898 504346 282134
rect 504582 281898 541226 282134
rect 541462 281898 541546 282134
rect 541782 281898 578426 282134
rect 578662 281898 578746 282134
rect 578982 281898 582820 282134
rect 1104 281866 582820 281898
rect 1104 278734 582820 278766
rect 1104 278498 16706 278734
rect 16942 278498 17026 278734
rect 17262 278498 53906 278734
rect 54142 278498 54226 278734
rect 54462 278498 91106 278734
rect 91342 278498 91426 278734
rect 91662 278498 128306 278734
rect 128542 278498 128626 278734
rect 128862 278498 165506 278734
rect 165742 278498 165826 278734
rect 166062 278498 202706 278734
rect 202942 278498 203026 278734
rect 203262 278498 239906 278734
rect 240142 278498 240226 278734
rect 240462 278498 277106 278734
rect 277342 278498 277426 278734
rect 277662 278498 314306 278734
rect 314542 278498 314626 278734
rect 314862 278498 351506 278734
rect 351742 278498 351826 278734
rect 352062 278498 388706 278734
rect 388942 278498 389026 278734
rect 389262 278498 425906 278734
rect 426142 278498 426226 278734
rect 426462 278498 463106 278734
rect 463342 278498 463426 278734
rect 463662 278498 500306 278734
rect 500542 278498 500626 278734
rect 500862 278498 537506 278734
rect 537742 278498 537826 278734
rect 538062 278498 574706 278734
rect 574942 278498 575026 278734
rect 575262 278498 582820 278734
rect 1104 278414 582820 278498
rect 1104 278178 16706 278414
rect 16942 278178 17026 278414
rect 17262 278178 53906 278414
rect 54142 278178 54226 278414
rect 54462 278178 91106 278414
rect 91342 278178 91426 278414
rect 91662 278178 128306 278414
rect 128542 278178 128626 278414
rect 128862 278178 165506 278414
rect 165742 278178 165826 278414
rect 166062 278178 202706 278414
rect 202942 278178 203026 278414
rect 203262 278178 239906 278414
rect 240142 278178 240226 278414
rect 240462 278178 277106 278414
rect 277342 278178 277426 278414
rect 277662 278178 314306 278414
rect 314542 278178 314626 278414
rect 314862 278178 351506 278414
rect 351742 278178 351826 278414
rect 352062 278178 388706 278414
rect 388942 278178 389026 278414
rect 389262 278178 425906 278414
rect 426142 278178 426226 278414
rect 426462 278178 463106 278414
rect 463342 278178 463426 278414
rect 463662 278178 500306 278414
rect 500542 278178 500626 278414
rect 500862 278178 537506 278414
rect 537742 278178 537826 278414
rect 538062 278178 574706 278414
rect 574942 278178 575026 278414
rect 575262 278178 582820 278414
rect 1104 278146 582820 278178
rect 1104 275014 582820 275046
rect 1104 274778 12986 275014
rect 13222 274778 13306 275014
rect 13542 274778 50186 275014
rect 50422 274778 50506 275014
rect 50742 274778 87386 275014
rect 87622 274778 87706 275014
rect 87942 274778 124586 275014
rect 124822 274778 124906 275014
rect 125142 274778 161786 275014
rect 162022 274778 162106 275014
rect 162342 274778 198986 275014
rect 199222 274778 199306 275014
rect 199542 274778 236186 275014
rect 236422 274778 236506 275014
rect 236742 274778 273386 275014
rect 273622 274778 273706 275014
rect 273942 274778 310586 275014
rect 310822 274778 310906 275014
rect 311142 274778 347786 275014
rect 348022 274778 348106 275014
rect 348342 274778 384986 275014
rect 385222 274778 385306 275014
rect 385542 274778 422186 275014
rect 422422 274778 422506 275014
rect 422742 274778 459386 275014
rect 459622 274778 459706 275014
rect 459942 274778 496586 275014
rect 496822 274778 496906 275014
rect 497142 274778 533786 275014
rect 534022 274778 534106 275014
rect 534342 274778 570986 275014
rect 571222 274778 571306 275014
rect 571542 274778 582820 275014
rect 1104 274694 582820 274778
rect 1104 274458 12986 274694
rect 13222 274458 13306 274694
rect 13542 274458 50186 274694
rect 50422 274458 50506 274694
rect 50742 274458 87386 274694
rect 87622 274458 87706 274694
rect 87942 274458 124586 274694
rect 124822 274458 124906 274694
rect 125142 274458 161786 274694
rect 162022 274458 162106 274694
rect 162342 274458 198986 274694
rect 199222 274458 199306 274694
rect 199542 274458 236186 274694
rect 236422 274458 236506 274694
rect 236742 274458 273386 274694
rect 273622 274458 273706 274694
rect 273942 274458 310586 274694
rect 310822 274458 310906 274694
rect 311142 274458 347786 274694
rect 348022 274458 348106 274694
rect 348342 274458 384986 274694
rect 385222 274458 385306 274694
rect 385542 274458 422186 274694
rect 422422 274458 422506 274694
rect 422742 274458 459386 274694
rect 459622 274458 459706 274694
rect 459942 274458 496586 274694
rect 496822 274458 496906 274694
rect 497142 274458 533786 274694
rect 534022 274458 534106 274694
rect 534342 274458 570986 274694
rect 571222 274458 571306 274694
rect 571542 274458 582820 274694
rect 1104 274426 582820 274458
rect 1104 271294 582820 271326
rect 1104 271058 9266 271294
rect 9502 271058 9586 271294
rect 9822 271058 46466 271294
rect 46702 271058 46786 271294
rect 47022 271058 83666 271294
rect 83902 271058 83986 271294
rect 84222 271058 120866 271294
rect 121102 271058 121186 271294
rect 121422 271058 158066 271294
rect 158302 271058 158386 271294
rect 158622 271058 195266 271294
rect 195502 271058 195586 271294
rect 195822 271058 232466 271294
rect 232702 271058 232786 271294
rect 233022 271058 269666 271294
rect 269902 271058 269986 271294
rect 270222 271058 306866 271294
rect 307102 271058 307186 271294
rect 307422 271058 344066 271294
rect 344302 271058 344386 271294
rect 344622 271058 381266 271294
rect 381502 271058 381586 271294
rect 381822 271058 418466 271294
rect 418702 271058 418786 271294
rect 419022 271058 455666 271294
rect 455902 271058 455986 271294
rect 456222 271058 492866 271294
rect 493102 271058 493186 271294
rect 493422 271058 530066 271294
rect 530302 271058 530386 271294
rect 530622 271058 567266 271294
rect 567502 271058 567586 271294
rect 567822 271058 582820 271294
rect 1104 270974 582820 271058
rect 1104 270738 9266 270974
rect 9502 270738 9586 270974
rect 9822 270738 46466 270974
rect 46702 270738 46786 270974
rect 47022 270738 83666 270974
rect 83902 270738 83986 270974
rect 84222 270738 120866 270974
rect 121102 270738 121186 270974
rect 121422 270738 158066 270974
rect 158302 270738 158386 270974
rect 158622 270738 195266 270974
rect 195502 270738 195586 270974
rect 195822 270738 232466 270974
rect 232702 270738 232786 270974
rect 233022 270738 269666 270974
rect 269902 270738 269986 270974
rect 270222 270738 306866 270974
rect 307102 270738 307186 270974
rect 307422 270738 344066 270974
rect 344302 270738 344386 270974
rect 344622 270738 381266 270974
rect 381502 270738 381586 270974
rect 381822 270738 418466 270974
rect 418702 270738 418786 270974
rect 419022 270738 455666 270974
rect 455902 270738 455986 270974
rect 456222 270738 492866 270974
rect 493102 270738 493186 270974
rect 493422 270738 530066 270974
rect 530302 270738 530386 270974
rect 530622 270738 567266 270974
rect 567502 270738 567586 270974
rect 567822 270738 582820 270974
rect 1104 270706 582820 270738
rect 1104 267574 582820 267606
rect 1104 267338 5546 267574
rect 5782 267338 5866 267574
rect 6102 267338 42746 267574
rect 42982 267338 43066 267574
rect 43302 267338 79946 267574
rect 80182 267338 80266 267574
rect 80502 267338 117146 267574
rect 117382 267338 117466 267574
rect 117702 267338 154346 267574
rect 154582 267338 154666 267574
rect 154902 267338 191546 267574
rect 191782 267338 191866 267574
rect 192102 267338 228746 267574
rect 228982 267338 229066 267574
rect 229302 267338 265946 267574
rect 266182 267338 266266 267574
rect 266502 267338 303146 267574
rect 303382 267338 303466 267574
rect 303702 267338 340346 267574
rect 340582 267338 340666 267574
rect 340902 267338 377546 267574
rect 377782 267338 377866 267574
rect 378102 267338 414746 267574
rect 414982 267338 415066 267574
rect 415302 267338 451946 267574
rect 452182 267338 452266 267574
rect 452502 267338 489146 267574
rect 489382 267338 489466 267574
rect 489702 267338 526346 267574
rect 526582 267338 526666 267574
rect 526902 267338 563546 267574
rect 563782 267338 563866 267574
rect 564102 267338 582820 267574
rect 1104 267254 582820 267338
rect 1104 267018 5546 267254
rect 5782 267018 5866 267254
rect 6102 267018 42746 267254
rect 42982 267018 43066 267254
rect 43302 267018 79946 267254
rect 80182 267018 80266 267254
rect 80502 267018 117146 267254
rect 117382 267018 117466 267254
rect 117702 267018 154346 267254
rect 154582 267018 154666 267254
rect 154902 267018 191546 267254
rect 191782 267018 191866 267254
rect 192102 267018 228746 267254
rect 228982 267018 229066 267254
rect 229302 267018 265946 267254
rect 266182 267018 266266 267254
rect 266502 267018 303146 267254
rect 303382 267018 303466 267254
rect 303702 267018 340346 267254
rect 340582 267018 340666 267254
rect 340902 267018 377546 267254
rect 377782 267018 377866 267254
rect 378102 267018 414746 267254
rect 414982 267018 415066 267254
rect 415302 267018 451946 267254
rect 452182 267018 452266 267254
rect 452502 267018 489146 267254
rect 489382 267018 489466 267254
rect 489702 267018 526346 267254
rect 526582 267018 526666 267254
rect 526902 267018 563546 267254
rect 563782 267018 563866 267254
rect 564102 267018 582820 267254
rect 1104 266986 582820 267018
rect 1104 263854 582820 263886
rect 1104 263618 1826 263854
rect 2062 263618 2146 263854
rect 2382 263618 39026 263854
rect 39262 263618 39346 263854
rect 39582 263618 76226 263854
rect 76462 263618 76546 263854
rect 76782 263618 113426 263854
rect 113662 263618 113746 263854
rect 113982 263618 150626 263854
rect 150862 263618 150946 263854
rect 151182 263618 187826 263854
rect 188062 263618 188146 263854
rect 188382 263618 225026 263854
rect 225262 263618 225346 263854
rect 225582 263618 262226 263854
rect 262462 263618 262546 263854
rect 262782 263618 299426 263854
rect 299662 263618 299746 263854
rect 299982 263618 336626 263854
rect 336862 263618 336946 263854
rect 337182 263618 373826 263854
rect 374062 263618 374146 263854
rect 374382 263618 411026 263854
rect 411262 263618 411346 263854
rect 411582 263618 448226 263854
rect 448462 263618 448546 263854
rect 448782 263618 485426 263854
rect 485662 263618 485746 263854
rect 485982 263618 522626 263854
rect 522862 263618 522946 263854
rect 523182 263618 559826 263854
rect 560062 263618 560146 263854
rect 560382 263618 582820 263854
rect 1104 263534 582820 263618
rect 1104 263298 1826 263534
rect 2062 263298 2146 263534
rect 2382 263298 39026 263534
rect 39262 263298 39346 263534
rect 39582 263298 76226 263534
rect 76462 263298 76546 263534
rect 76782 263298 113426 263534
rect 113662 263298 113746 263534
rect 113982 263298 150626 263534
rect 150862 263298 150946 263534
rect 151182 263298 187826 263534
rect 188062 263298 188146 263534
rect 188382 263298 225026 263534
rect 225262 263298 225346 263534
rect 225582 263298 262226 263534
rect 262462 263298 262546 263534
rect 262782 263298 299426 263534
rect 299662 263298 299746 263534
rect 299982 263298 336626 263534
rect 336862 263298 336946 263534
rect 337182 263298 373826 263534
rect 374062 263298 374146 263534
rect 374382 263298 411026 263534
rect 411262 263298 411346 263534
rect 411582 263298 448226 263534
rect 448462 263298 448546 263534
rect 448782 263298 485426 263534
rect 485662 263298 485746 263534
rect 485982 263298 522626 263534
rect 522862 263298 522946 263534
rect 523182 263298 559826 263534
rect 560062 263298 560146 263534
rect 560382 263298 582820 263534
rect 1104 263266 582820 263298
rect 1104 252694 582820 252726
rect 1104 252458 27866 252694
rect 28102 252458 28186 252694
rect 28422 252458 65066 252694
rect 65302 252458 65386 252694
rect 65622 252458 102266 252694
rect 102502 252458 102586 252694
rect 102822 252458 139466 252694
rect 139702 252458 139786 252694
rect 140022 252458 176666 252694
rect 176902 252458 176986 252694
rect 177222 252458 213866 252694
rect 214102 252458 214186 252694
rect 214422 252458 251066 252694
rect 251302 252458 251386 252694
rect 251622 252458 288266 252694
rect 288502 252458 288586 252694
rect 288822 252458 325466 252694
rect 325702 252458 325786 252694
rect 326022 252458 362666 252694
rect 362902 252458 362986 252694
rect 363222 252458 399866 252694
rect 400102 252458 400186 252694
rect 400422 252458 437066 252694
rect 437302 252458 437386 252694
rect 437622 252458 474266 252694
rect 474502 252458 474586 252694
rect 474822 252458 511466 252694
rect 511702 252458 511786 252694
rect 512022 252458 548666 252694
rect 548902 252458 548986 252694
rect 549222 252458 582820 252694
rect 1104 252374 582820 252458
rect 1104 252138 27866 252374
rect 28102 252138 28186 252374
rect 28422 252138 65066 252374
rect 65302 252138 65386 252374
rect 65622 252138 102266 252374
rect 102502 252138 102586 252374
rect 102822 252138 139466 252374
rect 139702 252138 139786 252374
rect 140022 252138 176666 252374
rect 176902 252138 176986 252374
rect 177222 252138 213866 252374
rect 214102 252138 214186 252374
rect 214422 252138 251066 252374
rect 251302 252138 251386 252374
rect 251622 252138 288266 252374
rect 288502 252138 288586 252374
rect 288822 252138 325466 252374
rect 325702 252138 325786 252374
rect 326022 252138 362666 252374
rect 362902 252138 362986 252374
rect 363222 252138 399866 252374
rect 400102 252138 400186 252374
rect 400422 252138 437066 252374
rect 437302 252138 437386 252374
rect 437622 252138 474266 252374
rect 474502 252138 474586 252374
rect 474822 252138 511466 252374
rect 511702 252138 511786 252374
rect 512022 252138 548666 252374
rect 548902 252138 548986 252374
rect 549222 252138 582820 252374
rect 1104 252106 582820 252138
rect 1104 248974 582820 249006
rect 1104 248738 24146 248974
rect 24382 248738 24466 248974
rect 24702 248738 61346 248974
rect 61582 248738 61666 248974
rect 61902 248738 98546 248974
rect 98782 248738 98866 248974
rect 99102 248738 135746 248974
rect 135982 248738 136066 248974
rect 136302 248738 172946 248974
rect 173182 248738 173266 248974
rect 173502 248738 210146 248974
rect 210382 248738 210466 248974
rect 210702 248738 247346 248974
rect 247582 248738 247666 248974
rect 247902 248738 284546 248974
rect 284782 248738 284866 248974
rect 285102 248738 321746 248974
rect 321982 248738 322066 248974
rect 322302 248738 358946 248974
rect 359182 248738 359266 248974
rect 359502 248738 396146 248974
rect 396382 248738 396466 248974
rect 396702 248738 433346 248974
rect 433582 248738 433666 248974
rect 433902 248738 470546 248974
rect 470782 248738 470866 248974
rect 471102 248738 507746 248974
rect 507982 248738 508066 248974
rect 508302 248738 544946 248974
rect 545182 248738 545266 248974
rect 545502 248738 582146 248974
rect 582382 248738 582466 248974
rect 582702 248738 582820 248974
rect 1104 248654 582820 248738
rect 1104 248418 24146 248654
rect 24382 248418 24466 248654
rect 24702 248418 61346 248654
rect 61582 248418 61666 248654
rect 61902 248418 98546 248654
rect 98782 248418 98866 248654
rect 99102 248418 135746 248654
rect 135982 248418 136066 248654
rect 136302 248418 172946 248654
rect 173182 248418 173266 248654
rect 173502 248418 210146 248654
rect 210382 248418 210466 248654
rect 210702 248418 247346 248654
rect 247582 248418 247666 248654
rect 247902 248418 284546 248654
rect 284782 248418 284866 248654
rect 285102 248418 321746 248654
rect 321982 248418 322066 248654
rect 322302 248418 358946 248654
rect 359182 248418 359266 248654
rect 359502 248418 396146 248654
rect 396382 248418 396466 248654
rect 396702 248418 433346 248654
rect 433582 248418 433666 248654
rect 433902 248418 470546 248654
rect 470782 248418 470866 248654
rect 471102 248418 507746 248654
rect 507982 248418 508066 248654
rect 508302 248418 544946 248654
rect 545182 248418 545266 248654
rect 545502 248418 582146 248654
rect 582382 248418 582466 248654
rect 582702 248418 582820 248654
rect 1104 248386 582820 248418
rect 1104 245254 582820 245286
rect 1104 245018 20426 245254
rect 20662 245018 20746 245254
rect 20982 245018 57626 245254
rect 57862 245018 57946 245254
rect 58182 245018 94826 245254
rect 95062 245018 95146 245254
rect 95382 245018 132026 245254
rect 132262 245018 132346 245254
rect 132582 245018 169226 245254
rect 169462 245018 169546 245254
rect 169782 245018 206426 245254
rect 206662 245018 206746 245254
rect 206982 245018 243626 245254
rect 243862 245018 243946 245254
rect 244182 245018 280826 245254
rect 281062 245018 281146 245254
rect 281382 245018 318026 245254
rect 318262 245018 318346 245254
rect 318582 245018 355226 245254
rect 355462 245018 355546 245254
rect 355782 245018 392426 245254
rect 392662 245018 392746 245254
rect 392982 245018 429626 245254
rect 429862 245018 429946 245254
rect 430182 245018 466826 245254
rect 467062 245018 467146 245254
rect 467382 245018 504026 245254
rect 504262 245018 504346 245254
rect 504582 245018 541226 245254
rect 541462 245018 541546 245254
rect 541782 245018 578426 245254
rect 578662 245018 578746 245254
rect 578982 245018 582820 245254
rect 1104 244934 582820 245018
rect 1104 244698 20426 244934
rect 20662 244698 20746 244934
rect 20982 244698 57626 244934
rect 57862 244698 57946 244934
rect 58182 244698 94826 244934
rect 95062 244698 95146 244934
rect 95382 244698 132026 244934
rect 132262 244698 132346 244934
rect 132582 244698 169226 244934
rect 169462 244698 169546 244934
rect 169782 244698 206426 244934
rect 206662 244698 206746 244934
rect 206982 244698 243626 244934
rect 243862 244698 243946 244934
rect 244182 244698 280826 244934
rect 281062 244698 281146 244934
rect 281382 244698 318026 244934
rect 318262 244698 318346 244934
rect 318582 244698 355226 244934
rect 355462 244698 355546 244934
rect 355782 244698 392426 244934
rect 392662 244698 392746 244934
rect 392982 244698 429626 244934
rect 429862 244698 429946 244934
rect 430182 244698 466826 244934
rect 467062 244698 467146 244934
rect 467382 244698 504026 244934
rect 504262 244698 504346 244934
rect 504582 244698 541226 244934
rect 541462 244698 541546 244934
rect 541782 244698 578426 244934
rect 578662 244698 578746 244934
rect 578982 244698 582820 244934
rect 1104 244666 582820 244698
rect 1104 241534 582820 241566
rect 1104 241298 16706 241534
rect 16942 241298 17026 241534
rect 17262 241298 53906 241534
rect 54142 241298 54226 241534
rect 54462 241298 91106 241534
rect 91342 241298 91426 241534
rect 91662 241298 128306 241534
rect 128542 241298 128626 241534
rect 128862 241298 165506 241534
rect 165742 241298 165826 241534
rect 166062 241298 202706 241534
rect 202942 241298 203026 241534
rect 203262 241298 239906 241534
rect 240142 241298 240226 241534
rect 240462 241298 277106 241534
rect 277342 241298 277426 241534
rect 277662 241298 314306 241534
rect 314542 241298 314626 241534
rect 314862 241298 351506 241534
rect 351742 241298 351826 241534
rect 352062 241298 388706 241534
rect 388942 241298 389026 241534
rect 389262 241298 425906 241534
rect 426142 241298 426226 241534
rect 426462 241298 463106 241534
rect 463342 241298 463426 241534
rect 463662 241298 500306 241534
rect 500542 241298 500626 241534
rect 500862 241298 537506 241534
rect 537742 241298 537826 241534
rect 538062 241298 574706 241534
rect 574942 241298 575026 241534
rect 575262 241298 582820 241534
rect 1104 241214 582820 241298
rect 1104 240978 16706 241214
rect 16942 240978 17026 241214
rect 17262 240978 53906 241214
rect 54142 240978 54226 241214
rect 54462 240978 91106 241214
rect 91342 240978 91426 241214
rect 91662 240978 128306 241214
rect 128542 240978 128626 241214
rect 128862 240978 165506 241214
rect 165742 240978 165826 241214
rect 166062 240978 202706 241214
rect 202942 240978 203026 241214
rect 203262 240978 239906 241214
rect 240142 240978 240226 241214
rect 240462 240978 277106 241214
rect 277342 240978 277426 241214
rect 277662 240978 314306 241214
rect 314542 240978 314626 241214
rect 314862 240978 351506 241214
rect 351742 240978 351826 241214
rect 352062 240978 388706 241214
rect 388942 240978 389026 241214
rect 389262 240978 425906 241214
rect 426142 240978 426226 241214
rect 426462 240978 463106 241214
rect 463342 240978 463426 241214
rect 463662 240978 500306 241214
rect 500542 240978 500626 241214
rect 500862 240978 537506 241214
rect 537742 240978 537826 241214
rect 538062 240978 574706 241214
rect 574942 240978 575026 241214
rect 575262 240978 582820 241214
rect 1104 240946 582820 240978
rect 1104 237814 582820 237846
rect 1104 237578 12986 237814
rect 13222 237578 13306 237814
rect 13542 237578 50186 237814
rect 50422 237578 50506 237814
rect 50742 237578 87386 237814
rect 87622 237578 87706 237814
rect 87942 237578 124586 237814
rect 124822 237578 124906 237814
rect 125142 237578 161786 237814
rect 162022 237578 162106 237814
rect 162342 237578 198986 237814
rect 199222 237578 199306 237814
rect 199542 237578 236186 237814
rect 236422 237578 236506 237814
rect 236742 237578 273386 237814
rect 273622 237578 273706 237814
rect 273942 237578 310586 237814
rect 310822 237578 310906 237814
rect 311142 237578 347786 237814
rect 348022 237578 348106 237814
rect 348342 237578 384986 237814
rect 385222 237578 385306 237814
rect 385542 237578 422186 237814
rect 422422 237578 422506 237814
rect 422742 237578 459386 237814
rect 459622 237578 459706 237814
rect 459942 237578 496586 237814
rect 496822 237578 496906 237814
rect 497142 237578 533786 237814
rect 534022 237578 534106 237814
rect 534342 237578 570986 237814
rect 571222 237578 571306 237814
rect 571542 237578 582820 237814
rect 1104 237494 582820 237578
rect 1104 237258 12986 237494
rect 13222 237258 13306 237494
rect 13542 237258 50186 237494
rect 50422 237258 50506 237494
rect 50742 237258 87386 237494
rect 87622 237258 87706 237494
rect 87942 237258 124586 237494
rect 124822 237258 124906 237494
rect 125142 237258 161786 237494
rect 162022 237258 162106 237494
rect 162342 237258 198986 237494
rect 199222 237258 199306 237494
rect 199542 237258 236186 237494
rect 236422 237258 236506 237494
rect 236742 237258 273386 237494
rect 273622 237258 273706 237494
rect 273942 237258 310586 237494
rect 310822 237258 310906 237494
rect 311142 237258 347786 237494
rect 348022 237258 348106 237494
rect 348342 237258 384986 237494
rect 385222 237258 385306 237494
rect 385542 237258 422186 237494
rect 422422 237258 422506 237494
rect 422742 237258 459386 237494
rect 459622 237258 459706 237494
rect 459942 237258 496586 237494
rect 496822 237258 496906 237494
rect 497142 237258 533786 237494
rect 534022 237258 534106 237494
rect 534342 237258 570986 237494
rect 571222 237258 571306 237494
rect 571542 237258 582820 237494
rect 1104 237226 582820 237258
rect 1104 234094 582820 234126
rect 1104 233858 9266 234094
rect 9502 233858 9586 234094
rect 9822 233858 46466 234094
rect 46702 233858 46786 234094
rect 47022 233858 83666 234094
rect 83902 233858 83986 234094
rect 84222 233858 120866 234094
rect 121102 233858 121186 234094
rect 121422 233858 158066 234094
rect 158302 233858 158386 234094
rect 158622 233858 195266 234094
rect 195502 233858 195586 234094
rect 195822 233858 232466 234094
rect 232702 233858 232786 234094
rect 233022 233858 269666 234094
rect 269902 233858 269986 234094
rect 270222 233858 306866 234094
rect 307102 233858 307186 234094
rect 307422 233858 344066 234094
rect 344302 233858 344386 234094
rect 344622 233858 381266 234094
rect 381502 233858 381586 234094
rect 381822 233858 418466 234094
rect 418702 233858 418786 234094
rect 419022 233858 455666 234094
rect 455902 233858 455986 234094
rect 456222 233858 492866 234094
rect 493102 233858 493186 234094
rect 493422 233858 530066 234094
rect 530302 233858 530386 234094
rect 530622 233858 567266 234094
rect 567502 233858 567586 234094
rect 567822 233858 582820 234094
rect 1104 233774 582820 233858
rect 1104 233538 9266 233774
rect 9502 233538 9586 233774
rect 9822 233538 46466 233774
rect 46702 233538 46786 233774
rect 47022 233538 83666 233774
rect 83902 233538 83986 233774
rect 84222 233538 120866 233774
rect 121102 233538 121186 233774
rect 121422 233538 158066 233774
rect 158302 233538 158386 233774
rect 158622 233538 195266 233774
rect 195502 233538 195586 233774
rect 195822 233538 232466 233774
rect 232702 233538 232786 233774
rect 233022 233538 269666 233774
rect 269902 233538 269986 233774
rect 270222 233538 306866 233774
rect 307102 233538 307186 233774
rect 307422 233538 344066 233774
rect 344302 233538 344386 233774
rect 344622 233538 381266 233774
rect 381502 233538 381586 233774
rect 381822 233538 418466 233774
rect 418702 233538 418786 233774
rect 419022 233538 455666 233774
rect 455902 233538 455986 233774
rect 456222 233538 492866 233774
rect 493102 233538 493186 233774
rect 493422 233538 530066 233774
rect 530302 233538 530386 233774
rect 530622 233538 567266 233774
rect 567502 233538 567586 233774
rect 567822 233538 582820 233774
rect 1104 233506 582820 233538
rect 1104 230374 582820 230406
rect 1104 230138 5546 230374
rect 5782 230138 5866 230374
rect 6102 230138 42746 230374
rect 42982 230138 43066 230374
rect 43302 230138 79946 230374
rect 80182 230138 80266 230374
rect 80502 230138 117146 230374
rect 117382 230138 117466 230374
rect 117702 230138 154346 230374
rect 154582 230138 154666 230374
rect 154902 230138 191546 230374
rect 191782 230138 191866 230374
rect 192102 230138 228746 230374
rect 228982 230138 229066 230374
rect 229302 230138 265946 230374
rect 266182 230138 266266 230374
rect 266502 230138 303146 230374
rect 303382 230138 303466 230374
rect 303702 230138 340346 230374
rect 340582 230138 340666 230374
rect 340902 230138 377546 230374
rect 377782 230138 377866 230374
rect 378102 230138 414746 230374
rect 414982 230138 415066 230374
rect 415302 230138 451946 230374
rect 452182 230138 452266 230374
rect 452502 230138 489146 230374
rect 489382 230138 489466 230374
rect 489702 230138 526346 230374
rect 526582 230138 526666 230374
rect 526902 230138 563546 230374
rect 563782 230138 563866 230374
rect 564102 230138 582820 230374
rect 1104 230054 582820 230138
rect 1104 229818 5546 230054
rect 5782 229818 5866 230054
rect 6102 229818 42746 230054
rect 42982 229818 43066 230054
rect 43302 229818 79946 230054
rect 80182 229818 80266 230054
rect 80502 229818 117146 230054
rect 117382 229818 117466 230054
rect 117702 229818 154346 230054
rect 154582 229818 154666 230054
rect 154902 229818 191546 230054
rect 191782 229818 191866 230054
rect 192102 229818 228746 230054
rect 228982 229818 229066 230054
rect 229302 229818 265946 230054
rect 266182 229818 266266 230054
rect 266502 229818 303146 230054
rect 303382 229818 303466 230054
rect 303702 229818 340346 230054
rect 340582 229818 340666 230054
rect 340902 229818 377546 230054
rect 377782 229818 377866 230054
rect 378102 229818 414746 230054
rect 414982 229818 415066 230054
rect 415302 229818 451946 230054
rect 452182 229818 452266 230054
rect 452502 229818 489146 230054
rect 489382 229818 489466 230054
rect 489702 229818 526346 230054
rect 526582 229818 526666 230054
rect 526902 229818 563546 230054
rect 563782 229818 563866 230054
rect 564102 229818 582820 230054
rect 1104 229786 582820 229818
rect 1104 226654 582820 226686
rect 1104 226418 1826 226654
rect 2062 226418 2146 226654
rect 2382 226418 39026 226654
rect 39262 226418 39346 226654
rect 39582 226418 76226 226654
rect 76462 226418 76546 226654
rect 76782 226418 113426 226654
rect 113662 226418 113746 226654
rect 113982 226418 150626 226654
rect 150862 226418 150946 226654
rect 151182 226418 187826 226654
rect 188062 226418 188146 226654
rect 188382 226418 225026 226654
rect 225262 226418 225346 226654
rect 225582 226418 262226 226654
rect 262462 226418 262546 226654
rect 262782 226418 299426 226654
rect 299662 226418 299746 226654
rect 299982 226418 336626 226654
rect 336862 226418 336946 226654
rect 337182 226418 373826 226654
rect 374062 226418 374146 226654
rect 374382 226418 411026 226654
rect 411262 226418 411346 226654
rect 411582 226418 448226 226654
rect 448462 226418 448546 226654
rect 448782 226418 485426 226654
rect 485662 226418 485746 226654
rect 485982 226418 522626 226654
rect 522862 226418 522946 226654
rect 523182 226418 559826 226654
rect 560062 226418 560146 226654
rect 560382 226418 582820 226654
rect 1104 226334 582820 226418
rect 1104 226098 1826 226334
rect 2062 226098 2146 226334
rect 2382 226098 39026 226334
rect 39262 226098 39346 226334
rect 39582 226098 76226 226334
rect 76462 226098 76546 226334
rect 76782 226098 113426 226334
rect 113662 226098 113746 226334
rect 113982 226098 150626 226334
rect 150862 226098 150946 226334
rect 151182 226098 187826 226334
rect 188062 226098 188146 226334
rect 188382 226098 225026 226334
rect 225262 226098 225346 226334
rect 225582 226098 262226 226334
rect 262462 226098 262546 226334
rect 262782 226098 299426 226334
rect 299662 226098 299746 226334
rect 299982 226098 336626 226334
rect 336862 226098 336946 226334
rect 337182 226098 373826 226334
rect 374062 226098 374146 226334
rect 374382 226098 411026 226334
rect 411262 226098 411346 226334
rect 411582 226098 448226 226334
rect 448462 226098 448546 226334
rect 448782 226098 485426 226334
rect 485662 226098 485746 226334
rect 485982 226098 522626 226334
rect 522862 226098 522946 226334
rect 523182 226098 559826 226334
rect 560062 226098 560146 226334
rect 560382 226098 582820 226334
rect 1104 226066 582820 226098
rect 1104 215494 582820 215526
rect 1104 215258 27866 215494
rect 28102 215258 28186 215494
rect 28422 215258 65066 215494
rect 65302 215258 65386 215494
rect 65622 215258 102266 215494
rect 102502 215258 102586 215494
rect 102822 215258 139466 215494
rect 139702 215258 139786 215494
rect 140022 215258 176666 215494
rect 176902 215258 176986 215494
rect 177222 215258 213866 215494
rect 214102 215258 214186 215494
rect 214422 215258 251066 215494
rect 251302 215258 251386 215494
rect 251622 215258 288266 215494
rect 288502 215258 288586 215494
rect 288822 215258 325466 215494
rect 325702 215258 325786 215494
rect 326022 215258 362666 215494
rect 362902 215258 362986 215494
rect 363222 215258 399866 215494
rect 400102 215258 400186 215494
rect 400422 215258 437066 215494
rect 437302 215258 437386 215494
rect 437622 215258 474266 215494
rect 474502 215258 474586 215494
rect 474822 215258 511466 215494
rect 511702 215258 511786 215494
rect 512022 215258 548666 215494
rect 548902 215258 548986 215494
rect 549222 215258 582820 215494
rect 1104 215174 582820 215258
rect 1104 214938 27866 215174
rect 28102 214938 28186 215174
rect 28422 214938 65066 215174
rect 65302 214938 65386 215174
rect 65622 214938 102266 215174
rect 102502 214938 102586 215174
rect 102822 214938 139466 215174
rect 139702 214938 139786 215174
rect 140022 214938 176666 215174
rect 176902 214938 176986 215174
rect 177222 214938 213866 215174
rect 214102 214938 214186 215174
rect 214422 214938 251066 215174
rect 251302 214938 251386 215174
rect 251622 214938 288266 215174
rect 288502 214938 288586 215174
rect 288822 214938 325466 215174
rect 325702 214938 325786 215174
rect 326022 214938 362666 215174
rect 362902 214938 362986 215174
rect 363222 214938 399866 215174
rect 400102 214938 400186 215174
rect 400422 214938 437066 215174
rect 437302 214938 437386 215174
rect 437622 214938 474266 215174
rect 474502 214938 474586 215174
rect 474822 214938 511466 215174
rect 511702 214938 511786 215174
rect 512022 214938 548666 215174
rect 548902 214938 548986 215174
rect 549222 214938 582820 215174
rect 1104 214906 582820 214938
rect 1104 211774 582820 211806
rect 1104 211538 24146 211774
rect 24382 211538 24466 211774
rect 24702 211538 61346 211774
rect 61582 211538 61666 211774
rect 61902 211538 98546 211774
rect 98782 211538 98866 211774
rect 99102 211538 135746 211774
rect 135982 211538 136066 211774
rect 136302 211538 172946 211774
rect 173182 211538 173266 211774
rect 173502 211538 210146 211774
rect 210382 211538 210466 211774
rect 210702 211538 247346 211774
rect 247582 211538 247666 211774
rect 247902 211538 284546 211774
rect 284782 211538 284866 211774
rect 285102 211538 321746 211774
rect 321982 211538 322066 211774
rect 322302 211538 358946 211774
rect 359182 211538 359266 211774
rect 359502 211538 396146 211774
rect 396382 211538 396466 211774
rect 396702 211538 433346 211774
rect 433582 211538 433666 211774
rect 433902 211538 470546 211774
rect 470782 211538 470866 211774
rect 471102 211538 507746 211774
rect 507982 211538 508066 211774
rect 508302 211538 544946 211774
rect 545182 211538 545266 211774
rect 545502 211538 582146 211774
rect 582382 211538 582466 211774
rect 582702 211538 582820 211774
rect 1104 211454 582820 211538
rect 1104 211218 24146 211454
rect 24382 211218 24466 211454
rect 24702 211218 61346 211454
rect 61582 211218 61666 211454
rect 61902 211218 98546 211454
rect 98782 211218 98866 211454
rect 99102 211218 135746 211454
rect 135982 211218 136066 211454
rect 136302 211218 172946 211454
rect 173182 211218 173266 211454
rect 173502 211218 210146 211454
rect 210382 211218 210466 211454
rect 210702 211218 247346 211454
rect 247582 211218 247666 211454
rect 247902 211218 284546 211454
rect 284782 211218 284866 211454
rect 285102 211218 321746 211454
rect 321982 211218 322066 211454
rect 322302 211218 358946 211454
rect 359182 211218 359266 211454
rect 359502 211218 396146 211454
rect 396382 211218 396466 211454
rect 396702 211218 433346 211454
rect 433582 211218 433666 211454
rect 433902 211218 470546 211454
rect 470782 211218 470866 211454
rect 471102 211218 507746 211454
rect 507982 211218 508066 211454
rect 508302 211218 544946 211454
rect 545182 211218 545266 211454
rect 545502 211218 582146 211454
rect 582382 211218 582466 211454
rect 582702 211218 582820 211454
rect 1104 211186 582820 211218
rect 1104 208054 582820 208086
rect 1104 207818 20426 208054
rect 20662 207818 20746 208054
rect 20982 207818 57626 208054
rect 57862 207818 57946 208054
rect 58182 207818 94826 208054
rect 95062 207818 95146 208054
rect 95382 207818 132026 208054
rect 132262 207818 132346 208054
rect 132582 207818 169226 208054
rect 169462 207818 169546 208054
rect 169782 207818 206426 208054
rect 206662 207818 206746 208054
rect 206982 207818 243626 208054
rect 243862 207818 243946 208054
rect 244182 207818 280826 208054
rect 281062 207818 281146 208054
rect 281382 207818 318026 208054
rect 318262 207818 318346 208054
rect 318582 207818 355226 208054
rect 355462 207818 355546 208054
rect 355782 207818 392426 208054
rect 392662 207818 392746 208054
rect 392982 207818 429626 208054
rect 429862 207818 429946 208054
rect 430182 207818 466826 208054
rect 467062 207818 467146 208054
rect 467382 207818 504026 208054
rect 504262 207818 504346 208054
rect 504582 207818 541226 208054
rect 541462 207818 541546 208054
rect 541782 207818 578426 208054
rect 578662 207818 578746 208054
rect 578982 207818 582820 208054
rect 1104 207734 582820 207818
rect 1104 207498 20426 207734
rect 20662 207498 20746 207734
rect 20982 207498 57626 207734
rect 57862 207498 57946 207734
rect 58182 207498 94826 207734
rect 95062 207498 95146 207734
rect 95382 207498 132026 207734
rect 132262 207498 132346 207734
rect 132582 207498 169226 207734
rect 169462 207498 169546 207734
rect 169782 207498 206426 207734
rect 206662 207498 206746 207734
rect 206982 207498 243626 207734
rect 243862 207498 243946 207734
rect 244182 207498 280826 207734
rect 281062 207498 281146 207734
rect 281382 207498 318026 207734
rect 318262 207498 318346 207734
rect 318582 207498 355226 207734
rect 355462 207498 355546 207734
rect 355782 207498 392426 207734
rect 392662 207498 392746 207734
rect 392982 207498 429626 207734
rect 429862 207498 429946 207734
rect 430182 207498 466826 207734
rect 467062 207498 467146 207734
rect 467382 207498 504026 207734
rect 504262 207498 504346 207734
rect 504582 207498 541226 207734
rect 541462 207498 541546 207734
rect 541782 207498 578426 207734
rect 578662 207498 578746 207734
rect 578982 207498 582820 207734
rect 1104 207466 582820 207498
rect 1104 204334 582820 204366
rect 1104 204098 16706 204334
rect 16942 204098 17026 204334
rect 17262 204098 53906 204334
rect 54142 204098 54226 204334
rect 54462 204098 91106 204334
rect 91342 204098 91426 204334
rect 91662 204098 128306 204334
rect 128542 204098 128626 204334
rect 128862 204098 165506 204334
rect 165742 204098 165826 204334
rect 166062 204098 202706 204334
rect 202942 204098 203026 204334
rect 203262 204098 239906 204334
rect 240142 204098 240226 204334
rect 240462 204098 277106 204334
rect 277342 204098 277426 204334
rect 277662 204098 314306 204334
rect 314542 204098 314626 204334
rect 314862 204098 351506 204334
rect 351742 204098 351826 204334
rect 352062 204098 388706 204334
rect 388942 204098 389026 204334
rect 389262 204098 425906 204334
rect 426142 204098 426226 204334
rect 426462 204098 463106 204334
rect 463342 204098 463426 204334
rect 463662 204098 500306 204334
rect 500542 204098 500626 204334
rect 500862 204098 537506 204334
rect 537742 204098 537826 204334
rect 538062 204098 574706 204334
rect 574942 204098 575026 204334
rect 575262 204098 582820 204334
rect 1104 204014 582820 204098
rect 1104 203778 16706 204014
rect 16942 203778 17026 204014
rect 17262 203778 53906 204014
rect 54142 203778 54226 204014
rect 54462 203778 91106 204014
rect 91342 203778 91426 204014
rect 91662 203778 128306 204014
rect 128542 203778 128626 204014
rect 128862 203778 165506 204014
rect 165742 203778 165826 204014
rect 166062 203778 202706 204014
rect 202942 203778 203026 204014
rect 203262 203778 239906 204014
rect 240142 203778 240226 204014
rect 240462 203778 277106 204014
rect 277342 203778 277426 204014
rect 277662 203778 314306 204014
rect 314542 203778 314626 204014
rect 314862 203778 351506 204014
rect 351742 203778 351826 204014
rect 352062 203778 388706 204014
rect 388942 203778 389026 204014
rect 389262 203778 425906 204014
rect 426142 203778 426226 204014
rect 426462 203778 463106 204014
rect 463342 203778 463426 204014
rect 463662 203778 500306 204014
rect 500542 203778 500626 204014
rect 500862 203778 537506 204014
rect 537742 203778 537826 204014
rect 538062 203778 574706 204014
rect 574942 203778 575026 204014
rect 575262 203778 582820 204014
rect 1104 203746 582820 203778
rect 1104 200614 582820 200646
rect 1104 200378 12986 200614
rect 13222 200378 13306 200614
rect 13542 200378 50186 200614
rect 50422 200378 50506 200614
rect 50742 200378 87386 200614
rect 87622 200378 87706 200614
rect 87942 200378 124586 200614
rect 124822 200378 124906 200614
rect 125142 200378 161786 200614
rect 162022 200378 162106 200614
rect 162342 200378 198986 200614
rect 199222 200378 199306 200614
rect 199542 200378 236186 200614
rect 236422 200378 236506 200614
rect 236742 200378 273386 200614
rect 273622 200378 273706 200614
rect 273942 200378 310586 200614
rect 310822 200378 310906 200614
rect 311142 200378 347786 200614
rect 348022 200378 348106 200614
rect 348342 200378 384986 200614
rect 385222 200378 385306 200614
rect 385542 200378 422186 200614
rect 422422 200378 422506 200614
rect 422742 200378 459386 200614
rect 459622 200378 459706 200614
rect 459942 200378 496586 200614
rect 496822 200378 496906 200614
rect 497142 200378 533786 200614
rect 534022 200378 534106 200614
rect 534342 200378 570986 200614
rect 571222 200378 571306 200614
rect 571542 200378 582820 200614
rect 1104 200294 582820 200378
rect 1104 200058 12986 200294
rect 13222 200058 13306 200294
rect 13542 200058 50186 200294
rect 50422 200058 50506 200294
rect 50742 200058 87386 200294
rect 87622 200058 87706 200294
rect 87942 200058 124586 200294
rect 124822 200058 124906 200294
rect 125142 200058 161786 200294
rect 162022 200058 162106 200294
rect 162342 200058 198986 200294
rect 199222 200058 199306 200294
rect 199542 200058 236186 200294
rect 236422 200058 236506 200294
rect 236742 200058 273386 200294
rect 273622 200058 273706 200294
rect 273942 200058 310586 200294
rect 310822 200058 310906 200294
rect 311142 200058 347786 200294
rect 348022 200058 348106 200294
rect 348342 200058 384986 200294
rect 385222 200058 385306 200294
rect 385542 200058 422186 200294
rect 422422 200058 422506 200294
rect 422742 200058 459386 200294
rect 459622 200058 459706 200294
rect 459942 200058 496586 200294
rect 496822 200058 496906 200294
rect 497142 200058 533786 200294
rect 534022 200058 534106 200294
rect 534342 200058 570986 200294
rect 571222 200058 571306 200294
rect 571542 200058 582820 200294
rect 1104 200026 582820 200058
rect 1104 196894 582820 196926
rect 1104 196658 9266 196894
rect 9502 196658 9586 196894
rect 9822 196658 46466 196894
rect 46702 196658 46786 196894
rect 47022 196658 83666 196894
rect 83902 196658 83986 196894
rect 84222 196658 120866 196894
rect 121102 196658 121186 196894
rect 121422 196658 158066 196894
rect 158302 196658 158386 196894
rect 158622 196658 195266 196894
rect 195502 196658 195586 196894
rect 195822 196658 232466 196894
rect 232702 196658 232786 196894
rect 233022 196658 269666 196894
rect 269902 196658 269986 196894
rect 270222 196658 306866 196894
rect 307102 196658 307186 196894
rect 307422 196658 344066 196894
rect 344302 196658 344386 196894
rect 344622 196658 381266 196894
rect 381502 196658 381586 196894
rect 381822 196658 418466 196894
rect 418702 196658 418786 196894
rect 419022 196658 455666 196894
rect 455902 196658 455986 196894
rect 456222 196658 492866 196894
rect 493102 196658 493186 196894
rect 493422 196658 530066 196894
rect 530302 196658 530386 196894
rect 530622 196658 567266 196894
rect 567502 196658 567586 196894
rect 567822 196658 582820 196894
rect 1104 196574 582820 196658
rect 1104 196338 9266 196574
rect 9502 196338 9586 196574
rect 9822 196338 46466 196574
rect 46702 196338 46786 196574
rect 47022 196338 83666 196574
rect 83902 196338 83986 196574
rect 84222 196338 120866 196574
rect 121102 196338 121186 196574
rect 121422 196338 158066 196574
rect 158302 196338 158386 196574
rect 158622 196338 195266 196574
rect 195502 196338 195586 196574
rect 195822 196338 232466 196574
rect 232702 196338 232786 196574
rect 233022 196338 269666 196574
rect 269902 196338 269986 196574
rect 270222 196338 306866 196574
rect 307102 196338 307186 196574
rect 307422 196338 344066 196574
rect 344302 196338 344386 196574
rect 344622 196338 381266 196574
rect 381502 196338 381586 196574
rect 381822 196338 418466 196574
rect 418702 196338 418786 196574
rect 419022 196338 455666 196574
rect 455902 196338 455986 196574
rect 456222 196338 492866 196574
rect 493102 196338 493186 196574
rect 493422 196338 530066 196574
rect 530302 196338 530386 196574
rect 530622 196338 567266 196574
rect 567502 196338 567586 196574
rect 567822 196338 582820 196574
rect 1104 196306 582820 196338
rect 1104 193174 582820 193206
rect 1104 192938 5546 193174
rect 5782 192938 5866 193174
rect 6102 192938 42746 193174
rect 42982 192938 43066 193174
rect 43302 192938 79946 193174
rect 80182 192938 80266 193174
rect 80502 192938 117146 193174
rect 117382 192938 117466 193174
rect 117702 192938 154346 193174
rect 154582 192938 154666 193174
rect 154902 192938 191546 193174
rect 191782 192938 191866 193174
rect 192102 192938 228746 193174
rect 228982 192938 229066 193174
rect 229302 192938 265946 193174
rect 266182 192938 266266 193174
rect 266502 192938 303146 193174
rect 303382 192938 303466 193174
rect 303702 192938 340346 193174
rect 340582 192938 340666 193174
rect 340902 192938 377546 193174
rect 377782 192938 377866 193174
rect 378102 192938 414746 193174
rect 414982 192938 415066 193174
rect 415302 192938 451946 193174
rect 452182 192938 452266 193174
rect 452502 192938 489146 193174
rect 489382 192938 489466 193174
rect 489702 192938 526346 193174
rect 526582 192938 526666 193174
rect 526902 192938 563546 193174
rect 563782 192938 563866 193174
rect 564102 192938 582820 193174
rect 1104 192854 582820 192938
rect 1104 192618 5546 192854
rect 5782 192618 5866 192854
rect 6102 192618 42746 192854
rect 42982 192618 43066 192854
rect 43302 192618 79946 192854
rect 80182 192618 80266 192854
rect 80502 192618 117146 192854
rect 117382 192618 117466 192854
rect 117702 192618 154346 192854
rect 154582 192618 154666 192854
rect 154902 192618 191546 192854
rect 191782 192618 191866 192854
rect 192102 192618 228746 192854
rect 228982 192618 229066 192854
rect 229302 192618 265946 192854
rect 266182 192618 266266 192854
rect 266502 192618 303146 192854
rect 303382 192618 303466 192854
rect 303702 192618 340346 192854
rect 340582 192618 340666 192854
rect 340902 192618 377546 192854
rect 377782 192618 377866 192854
rect 378102 192618 414746 192854
rect 414982 192618 415066 192854
rect 415302 192618 451946 192854
rect 452182 192618 452266 192854
rect 452502 192618 489146 192854
rect 489382 192618 489466 192854
rect 489702 192618 526346 192854
rect 526582 192618 526666 192854
rect 526902 192618 563546 192854
rect 563782 192618 563866 192854
rect 564102 192618 582820 192854
rect 1104 192586 582820 192618
rect 1104 189454 582820 189486
rect 1104 189218 1826 189454
rect 2062 189218 2146 189454
rect 2382 189218 39026 189454
rect 39262 189218 39346 189454
rect 39582 189218 76226 189454
rect 76462 189218 76546 189454
rect 76782 189218 113426 189454
rect 113662 189218 113746 189454
rect 113982 189218 150626 189454
rect 150862 189218 150946 189454
rect 151182 189218 187826 189454
rect 188062 189218 188146 189454
rect 188382 189218 225026 189454
rect 225262 189218 225346 189454
rect 225582 189218 262226 189454
rect 262462 189218 262546 189454
rect 262782 189218 299426 189454
rect 299662 189218 299746 189454
rect 299982 189218 336626 189454
rect 336862 189218 336946 189454
rect 337182 189218 373826 189454
rect 374062 189218 374146 189454
rect 374382 189218 411026 189454
rect 411262 189218 411346 189454
rect 411582 189218 448226 189454
rect 448462 189218 448546 189454
rect 448782 189218 485426 189454
rect 485662 189218 485746 189454
rect 485982 189218 522626 189454
rect 522862 189218 522946 189454
rect 523182 189218 559826 189454
rect 560062 189218 560146 189454
rect 560382 189218 582820 189454
rect 1104 189134 582820 189218
rect 1104 188898 1826 189134
rect 2062 188898 2146 189134
rect 2382 188898 39026 189134
rect 39262 188898 39346 189134
rect 39582 188898 76226 189134
rect 76462 188898 76546 189134
rect 76782 188898 113426 189134
rect 113662 188898 113746 189134
rect 113982 188898 150626 189134
rect 150862 188898 150946 189134
rect 151182 188898 187826 189134
rect 188062 188898 188146 189134
rect 188382 188898 225026 189134
rect 225262 188898 225346 189134
rect 225582 188898 262226 189134
rect 262462 188898 262546 189134
rect 262782 188898 299426 189134
rect 299662 188898 299746 189134
rect 299982 188898 336626 189134
rect 336862 188898 336946 189134
rect 337182 188898 373826 189134
rect 374062 188898 374146 189134
rect 374382 188898 411026 189134
rect 411262 188898 411346 189134
rect 411582 188898 448226 189134
rect 448462 188898 448546 189134
rect 448782 188898 485426 189134
rect 485662 188898 485746 189134
rect 485982 188898 522626 189134
rect 522862 188898 522946 189134
rect 523182 188898 559826 189134
rect 560062 188898 560146 189134
rect 560382 188898 582820 189134
rect 1104 188866 582820 188898
rect 1104 178294 582820 178326
rect 1104 178058 27866 178294
rect 28102 178058 28186 178294
rect 28422 178058 65066 178294
rect 65302 178058 65386 178294
rect 65622 178058 102266 178294
rect 102502 178058 102586 178294
rect 102822 178058 139466 178294
rect 139702 178058 139786 178294
rect 140022 178058 176666 178294
rect 176902 178058 176986 178294
rect 177222 178058 213866 178294
rect 214102 178058 214186 178294
rect 214422 178058 251066 178294
rect 251302 178058 251386 178294
rect 251622 178058 288266 178294
rect 288502 178058 288586 178294
rect 288822 178058 325466 178294
rect 325702 178058 325786 178294
rect 326022 178058 362666 178294
rect 362902 178058 362986 178294
rect 363222 178058 399866 178294
rect 400102 178058 400186 178294
rect 400422 178058 437066 178294
rect 437302 178058 437386 178294
rect 437622 178058 474266 178294
rect 474502 178058 474586 178294
rect 474822 178058 511466 178294
rect 511702 178058 511786 178294
rect 512022 178058 548666 178294
rect 548902 178058 548986 178294
rect 549222 178058 582820 178294
rect 1104 177974 582820 178058
rect 1104 177738 27866 177974
rect 28102 177738 28186 177974
rect 28422 177738 65066 177974
rect 65302 177738 65386 177974
rect 65622 177738 102266 177974
rect 102502 177738 102586 177974
rect 102822 177738 139466 177974
rect 139702 177738 139786 177974
rect 140022 177738 176666 177974
rect 176902 177738 176986 177974
rect 177222 177738 213866 177974
rect 214102 177738 214186 177974
rect 214422 177738 251066 177974
rect 251302 177738 251386 177974
rect 251622 177738 288266 177974
rect 288502 177738 288586 177974
rect 288822 177738 325466 177974
rect 325702 177738 325786 177974
rect 326022 177738 362666 177974
rect 362902 177738 362986 177974
rect 363222 177738 399866 177974
rect 400102 177738 400186 177974
rect 400422 177738 437066 177974
rect 437302 177738 437386 177974
rect 437622 177738 474266 177974
rect 474502 177738 474586 177974
rect 474822 177738 511466 177974
rect 511702 177738 511786 177974
rect 512022 177738 548666 177974
rect 548902 177738 548986 177974
rect 549222 177738 582820 177974
rect 1104 177706 582820 177738
rect 1104 174574 582820 174606
rect 1104 174338 24146 174574
rect 24382 174338 24466 174574
rect 24702 174338 61346 174574
rect 61582 174338 61666 174574
rect 61902 174338 98546 174574
rect 98782 174338 98866 174574
rect 99102 174338 135746 174574
rect 135982 174338 136066 174574
rect 136302 174338 172946 174574
rect 173182 174338 173266 174574
rect 173502 174338 210146 174574
rect 210382 174338 210466 174574
rect 210702 174338 247346 174574
rect 247582 174338 247666 174574
rect 247902 174338 284546 174574
rect 284782 174338 284866 174574
rect 285102 174338 321746 174574
rect 321982 174338 322066 174574
rect 322302 174338 358946 174574
rect 359182 174338 359266 174574
rect 359502 174338 396146 174574
rect 396382 174338 396466 174574
rect 396702 174338 433346 174574
rect 433582 174338 433666 174574
rect 433902 174338 470546 174574
rect 470782 174338 470866 174574
rect 471102 174338 507746 174574
rect 507982 174338 508066 174574
rect 508302 174338 544946 174574
rect 545182 174338 545266 174574
rect 545502 174338 582146 174574
rect 582382 174338 582466 174574
rect 582702 174338 582820 174574
rect 1104 174254 582820 174338
rect 1104 174018 24146 174254
rect 24382 174018 24466 174254
rect 24702 174018 61346 174254
rect 61582 174018 61666 174254
rect 61902 174018 98546 174254
rect 98782 174018 98866 174254
rect 99102 174018 135746 174254
rect 135982 174018 136066 174254
rect 136302 174018 172946 174254
rect 173182 174018 173266 174254
rect 173502 174018 210146 174254
rect 210382 174018 210466 174254
rect 210702 174018 247346 174254
rect 247582 174018 247666 174254
rect 247902 174018 284546 174254
rect 284782 174018 284866 174254
rect 285102 174018 321746 174254
rect 321982 174018 322066 174254
rect 322302 174018 358946 174254
rect 359182 174018 359266 174254
rect 359502 174018 396146 174254
rect 396382 174018 396466 174254
rect 396702 174018 433346 174254
rect 433582 174018 433666 174254
rect 433902 174018 470546 174254
rect 470782 174018 470866 174254
rect 471102 174018 507746 174254
rect 507982 174018 508066 174254
rect 508302 174018 544946 174254
rect 545182 174018 545266 174254
rect 545502 174018 582146 174254
rect 582382 174018 582466 174254
rect 582702 174018 582820 174254
rect 1104 173986 582820 174018
rect 1104 170854 582820 170886
rect 1104 170618 20426 170854
rect 20662 170618 20746 170854
rect 20982 170618 57626 170854
rect 57862 170618 57946 170854
rect 58182 170618 94826 170854
rect 95062 170618 95146 170854
rect 95382 170618 132026 170854
rect 132262 170618 132346 170854
rect 132582 170618 169226 170854
rect 169462 170618 169546 170854
rect 169782 170618 206426 170854
rect 206662 170618 206746 170854
rect 206982 170618 243626 170854
rect 243862 170618 243946 170854
rect 244182 170618 280826 170854
rect 281062 170618 281146 170854
rect 281382 170618 318026 170854
rect 318262 170618 318346 170854
rect 318582 170618 355226 170854
rect 355462 170618 355546 170854
rect 355782 170618 392426 170854
rect 392662 170618 392746 170854
rect 392982 170618 429626 170854
rect 429862 170618 429946 170854
rect 430182 170618 466826 170854
rect 467062 170618 467146 170854
rect 467382 170618 504026 170854
rect 504262 170618 504346 170854
rect 504582 170618 541226 170854
rect 541462 170618 541546 170854
rect 541782 170618 578426 170854
rect 578662 170618 578746 170854
rect 578982 170618 582820 170854
rect 1104 170534 582820 170618
rect 1104 170298 20426 170534
rect 20662 170298 20746 170534
rect 20982 170298 57626 170534
rect 57862 170298 57946 170534
rect 58182 170298 94826 170534
rect 95062 170298 95146 170534
rect 95382 170298 132026 170534
rect 132262 170298 132346 170534
rect 132582 170298 169226 170534
rect 169462 170298 169546 170534
rect 169782 170298 206426 170534
rect 206662 170298 206746 170534
rect 206982 170298 243626 170534
rect 243862 170298 243946 170534
rect 244182 170298 280826 170534
rect 281062 170298 281146 170534
rect 281382 170298 318026 170534
rect 318262 170298 318346 170534
rect 318582 170298 355226 170534
rect 355462 170298 355546 170534
rect 355782 170298 392426 170534
rect 392662 170298 392746 170534
rect 392982 170298 429626 170534
rect 429862 170298 429946 170534
rect 430182 170298 466826 170534
rect 467062 170298 467146 170534
rect 467382 170298 504026 170534
rect 504262 170298 504346 170534
rect 504582 170298 541226 170534
rect 541462 170298 541546 170534
rect 541782 170298 578426 170534
rect 578662 170298 578746 170534
rect 578982 170298 582820 170534
rect 1104 170266 582820 170298
rect 1104 167134 582820 167166
rect 1104 166898 16706 167134
rect 16942 166898 17026 167134
rect 17262 166898 53906 167134
rect 54142 166898 54226 167134
rect 54462 166898 91106 167134
rect 91342 166898 91426 167134
rect 91662 166898 128306 167134
rect 128542 166898 128626 167134
rect 128862 166898 165506 167134
rect 165742 166898 165826 167134
rect 166062 166898 202706 167134
rect 202942 166898 203026 167134
rect 203262 166898 239906 167134
rect 240142 166898 240226 167134
rect 240462 166898 277106 167134
rect 277342 166898 277426 167134
rect 277662 166898 314306 167134
rect 314542 166898 314626 167134
rect 314862 166898 351506 167134
rect 351742 166898 351826 167134
rect 352062 166898 388706 167134
rect 388942 166898 389026 167134
rect 389262 166898 425906 167134
rect 426142 166898 426226 167134
rect 426462 166898 463106 167134
rect 463342 166898 463426 167134
rect 463662 166898 500306 167134
rect 500542 166898 500626 167134
rect 500862 166898 537506 167134
rect 537742 166898 537826 167134
rect 538062 166898 574706 167134
rect 574942 166898 575026 167134
rect 575262 166898 582820 167134
rect 1104 166814 582820 166898
rect 1104 166578 16706 166814
rect 16942 166578 17026 166814
rect 17262 166578 53906 166814
rect 54142 166578 54226 166814
rect 54462 166578 91106 166814
rect 91342 166578 91426 166814
rect 91662 166578 128306 166814
rect 128542 166578 128626 166814
rect 128862 166578 165506 166814
rect 165742 166578 165826 166814
rect 166062 166578 202706 166814
rect 202942 166578 203026 166814
rect 203262 166578 239906 166814
rect 240142 166578 240226 166814
rect 240462 166578 277106 166814
rect 277342 166578 277426 166814
rect 277662 166578 314306 166814
rect 314542 166578 314626 166814
rect 314862 166578 351506 166814
rect 351742 166578 351826 166814
rect 352062 166578 388706 166814
rect 388942 166578 389026 166814
rect 389262 166578 425906 166814
rect 426142 166578 426226 166814
rect 426462 166578 463106 166814
rect 463342 166578 463426 166814
rect 463662 166578 500306 166814
rect 500542 166578 500626 166814
rect 500862 166578 537506 166814
rect 537742 166578 537826 166814
rect 538062 166578 574706 166814
rect 574942 166578 575026 166814
rect 575262 166578 582820 166814
rect 1104 166546 582820 166578
rect 1104 163414 582820 163446
rect 1104 163178 12986 163414
rect 13222 163178 13306 163414
rect 13542 163178 50186 163414
rect 50422 163178 50506 163414
rect 50742 163178 87386 163414
rect 87622 163178 87706 163414
rect 87942 163178 124586 163414
rect 124822 163178 124906 163414
rect 125142 163178 161786 163414
rect 162022 163178 162106 163414
rect 162342 163178 198986 163414
rect 199222 163178 199306 163414
rect 199542 163178 236186 163414
rect 236422 163178 236506 163414
rect 236742 163178 273386 163414
rect 273622 163178 273706 163414
rect 273942 163178 310586 163414
rect 310822 163178 310906 163414
rect 311142 163178 347786 163414
rect 348022 163178 348106 163414
rect 348342 163178 384986 163414
rect 385222 163178 385306 163414
rect 385542 163178 422186 163414
rect 422422 163178 422506 163414
rect 422742 163178 459386 163414
rect 459622 163178 459706 163414
rect 459942 163178 496586 163414
rect 496822 163178 496906 163414
rect 497142 163178 533786 163414
rect 534022 163178 534106 163414
rect 534342 163178 570986 163414
rect 571222 163178 571306 163414
rect 571542 163178 582820 163414
rect 1104 163094 582820 163178
rect 1104 162858 12986 163094
rect 13222 162858 13306 163094
rect 13542 162858 50186 163094
rect 50422 162858 50506 163094
rect 50742 162858 87386 163094
rect 87622 162858 87706 163094
rect 87942 162858 124586 163094
rect 124822 162858 124906 163094
rect 125142 162858 161786 163094
rect 162022 162858 162106 163094
rect 162342 162858 198986 163094
rect 199222 162858 199306 163094
rect 199542 162858 236186 163094
rect 236422 162858 236506 163094
rect 236742 162858 273386 163094
rect 273622 162858 273706 163094
rect 273942 162858 310586 163094
rect 310822 162858 310906 163094
rect 311142 162858 347786 163094
rect 348022 162858 348106 163094
rect 348342 162858 384986 163094
rect 385222 162858 385306 163094
rect 385542 162858 422186 163094
rect 422422 162858 422506 163094
rect 422742 162858 459386 163094
rect 459622 162858 459706 163094
rect 459942 162858 496586 163094
rect 496822 162858 496906 163094
rect 497142 162858 533786 163094
rect 534022 162858 534106 163094
rect 534342 162858 570986 163094
rect 571222 162858 571306 163094
rect 571542 162858 582820 163094
rect 1104 162826 582820 162858
rect 1104 159694 582820 159726
rect 1104 159458 9266 159694
rect 9502 159458 9586 159694
rect 9822 159458 46466 159694
rect 46702 159458 46786 159694
rect 47022 159458 83666 159694
rect 83902 159458 83986 159694
rect 84222 159458 120866 159694
rect 121102 159458 121186 159694
rect 121422 159458 158066 159694
rect 158302 159458 158386 159694
rect 158622 159458 195266 159694
rect 195502 159458 195586 159694
rect 195822 159458 232466 159694
rect 232702 159458 232786 159694
rect 233022 159458 269666 159694
rect 269902 159458 269986 159694
rect 270222 159458 306866 159694
rect 307102 159458 307186 159694
rect 307422 159458 344066 159694
rect 344302 159458 344386 159694
rect 344622 159458 381266 159694
rect 381502 159458 381586 159694
rect 381822 159458 418466 159694
rect 418702 159458 418786 159694
rect 419022 159458 455666 159694
rect 455902 159458 455986 159694
rect 456222 159458 492866 159694
rect 493102 159458 493186 159694
rect 493422 159458 530066 159694
rect 530302 159458 530386 159694
rect 530622 159458 567266 159694
rect 567502 159458 567586 159694
rect 567822 159458 582820 159694
rect 1104 159374 582820 159458
rect 1104 159138 9266 159374
rect 9502 159138 9586 159374
rect 9822 159138 46466 159374
rect 46702 159138 46786 159374
rect 47022 159138 83666 159374
rect 83902 159138 83986 159374
rect 84222 159138 120866 159374
rect 121102 159138 121186 159374
rect 121422 159138 158066 159374
rect 158302 159138 158386 159374
rect 158622 159138 195266 159374
rect 195502 159138 195586 159374
rect 195822 159138 232466 159374
rect 232702 159138 232786 159374
rect 233022 159138 269666 159374
rect 269902 159138 269986 159374
rect 270222 159138 306866 159374
rect 307102 159138 307186 159374
rect 307422 159138 344066 159374
rect 344302 159138 344386 159374
rect 344622 159138 381266 159374
rect 381502 159138 381586 159374
rect 381822 159138 418466 159374
rect 418702 159138 418786 159374
rect 419022 159138 455666 159374
rect 455902 159138 455986 159374
rect 456222 159138 492866 159374
rect 493102 159138 493186 159374
rect 493422 159138 530066 159374
rect 530302 159138 530386 159374
rect 530622 159138 567266 159374
rect 567502 159138 567586 159374
rect 567822 159138 582820 159374
rect 1104 159106 582820 159138
rect 1104 155974 582820 156006
rect 1104 155738 5546 155974
rect 5782 155738 5866 155974
rect 6102 155738 42746 155974
rect 42982 155738 43066 155974
rect 43302 155738 79946 155974
rect 80182 155738 80266 155974
rect 80502 155738 117146 155974
rect 117382 155738 117466 155974
rect 117702 155738 154346 155974
rect 154582 155738 154666 155974
rect 154902 155738 191546 155974
rect 191782 155738 191866 155974
rect 192102 155738 228746 155974
rect 228982 155738 229066 155974
rect 229302 155738 265946 155974
rect 266182 155738 266266 155974
rect 266502 155738 303146 155974
rect 303382 155738 303466 155974
rect 303702 155738 340346 155974
rect 340582 155738 340666 155974
rect 340902 155738 377546 155974
rect 377782 155738 377866 155974
rect 378102 155738 414746 155974
rect 414982 155738 415066 155974
rect 415302 155738 451946 155974
rect 452182 155738 452266 155974
rect 452502 155738 489146 155974
rect 489382 155738 489466 155974
rect 489702 155738 526346 155974
rect 526582 155738 526666 155974
rect 526902 155738 563546 155974
rect 563782 155738 563866 155974
rect 564102 155738 582820 155974
rect 1104 155654 582820 155738
rect 1104 155418 5546 155654
rect 5782 155418 5866 155654
rect 6102 155418 42746 155654
rect 42982 155418 43066 155654
rect 43302 155418 79946 155654
rect 80182 155418 80266 155654
rect 80502 155418 117146 155654
rect 117382 155418 117466 155654
rect 117702 155418 154346 155654
rect 154582 155418 154666 155654
rect 154902 155418 191546 155654
rect 191782 155418 191866 155654
rect 192102 155418 228746 155654
rect 228982 155418 229066 155654
rect 229302 155418 265946 155654
rect 266182 155418 266266 155654
rect 266502 155418 303146 155654
rect 303382 155418 303466 155654
rect 303702 155418 340346 155654
rect 340582 155418 340666 155654
rect 340902 155418 377546 155654
rect 377782 155418 377866 155654
rect 378102 155418 414746 155654
rect 414982 155418 415066 155654
rect 415302 155418 451946 155654
rect 452182 155418 452266 155654
rect 452502 155418 489146 155654
rect 489382 155418 489466 155654
rect 489702 155418 526346 155654
rect 526582 155418 526666 155654
rect 526902 155418 563546 155654
rect 563782 155418 563866 155654
rect 564102 155418 582820 155654
rect 1104 155386 582820 155418
rect 1104 152254 582820 152286
rect 1104 152018 1826 152254
rect 2062 152018 2146 152254
rect 2382 152018 39026 152254
rect 39262 152018 39346 152254
rect 39582 152018 76226 152254
rect 76462 152018 76546 152254
rect 76782 152018 113426 152254
rect 113662 152018 113746 152254
rect 113982 152018 150626 152254
rect 150862 152018 150946 152254
rect 151182 152018 187826 152254
rect 188062 152018 188146 152254
rect 188382 152018 225026 152254
rect 225262 152018 225346 152254
rect 225582 152018 262226 152254
rect 262462 152018 262546 152254
rect 262782 152018 299426 152254
rect 299662 152018 299746 152254
rect 299982 152018 336626 152254
rect 336862 152018 336946 152254
rect 337182 152018 373826 152254
rect 374062 152018 374146 152254
rect 374382 152018 411026 152254
rect 411262 152018 411346 152254
rect 411582 152018 448226 152254
rect 448462 152018 448546 152254
rect 448782 152018 485426 152254
rect 485662 152018 485746 152254
rect 485982 152018 522626 152254
rect 522862 152018 522946 152254
rect 523182 152018 559826 152254
rect 560062 152018 560146 152254
rect 560382 152018 582820 152254
rect 1104 151934 582820 152018
rect 1104 151698 1826 151934
rect 2062 151698 2146 151934
rect 2382 151698 39026 151934
rect 39262 151698 39346 151934
rect 39582 151698 76226 151934
rect 76462 151698 76546 151934
rect 76782 151698 113426 151934
rect 113662 151698 113746 151934
rect 113982 151698 150626 151934
rect 150862 151698 150946 151934
rect 151182 151698 187826 151934
rect 188062 151698 188146 151934
rect 188382 151698 225026 151934
rect 225262 151698 225346 151934
rect 225582 151698 262226 151934
rect 262462 151698 262546 151934
rect 262782 151698 299426 151934
rect 299662 151698 299746 151934
rect 299982 151698 336626 151934
rect 336862 151698 336946 151934
rect 337182 151698 373826 151934
rect 374062 151698 374146 151934
rect 374382 151698 411026 151934
rect 411262 151698 411346 151934
rect 411582 151698 448226 151934
rect 448462 151698 448546 151934
rect 448782 151698 485426 151934
rect 485662 151698 485746 151934
rect 485982 151698 522626 151934
rect 522862 151698 522946 151934
rect 523182 151698 559826 151934
rect 560062 151698 560146 151934
rect 560382 151698 582820 151934
rect 1104 151666 582820 151698
rect 1104 141094 582820 141126
rect 1104 140858 27866 141094
rect 28102 140858 28186 141094
rect 28422 140858 65066 141094
rect 65302 140858 65386 141094
rect 65622 140858 102266 141094
rect 102502 140858 102586 141094
rect 102822 140858 139466 141094
rect 139702 140858 139786 141094
rect 140022 140858 176666 141094
rect 176902 140858 176986 141094
rect 177222 140858 213866 141094
rect 214102 140858 214186 141094
rect 214422 140858 251066 141094
rect 251302 140858 251386 141094
rect 251622 140858 288266 141094
rect 288502 140858 288586 141094
rect 288822 140858 325466 141094
rect 325702 140858 325786 141094
rect 326022 140858 362666 141094
rect 362902 140858 362986 141094
rect 363222 140858 399866 141094
rect 400102 140858 400186 141094
rect 400422 140858 437066 141094
rect 437302 140858 437386 141094
rect 437622 140858 474266 141094
rect 474502 140858 474586 141094
rect 474822 140858 511466 141094
rect 511702 140858 511786 141094
rect 512022 140858 548666 141094
rect 548902 140858 548986 141094
rect 549222 140858 582820 141094
rect 1104 140774 582820 140858
rect 1104 140538 27866 140774
rect 28102 140538 28186 140774
rect 28422 140538 65066 140774
rect 65302 140538 65386 140774
rect 65622 140538 102266 140774
rect 102502 140538 102586 140774
rect 102822 140538 139466 140774
rect 139702 140538 139786 140774
rect 140022 140538 176666 140774
rect 176902 140538 176986 140774
rect 177222 140538 213866 140774
rect 214102 140538 214186 140774
rect 214422 140538 251066 140774
rect 251302 140538 251386 140774
rect 251622 140538 288266 140774
rect 288502 140538 288586 140774
rect 288822 140538 325466 140774
rect 325702 140538 325786 140774
rect 326022 140538 362666 140774
rect 362902 140538 362986 140774
rect 363222 140538 399866 140774
rect 400102 140538 400186 140774
rect 400422 140538 437066 140774
rect 437302 140538 437386 140774
rect 437622 140538 474266 140774
rect 474502 140538 474586 140774
rect 474822 140538 511466 140774
rect 511702 140538 511786 140774
rect 512022 140538 548666 140774
rect 548902 140538 548986 140774
rect 549222 140538 582820 140774
rect 1104 140506 582820 140538
rect 1104 137374 582820 137406
rect 1104 137138 24146 137374
rect 24382 137138 24466 137374
rect 24702 137138 61346 137374
rect 61582 137138 61666 137374
rect 61902 137138 98546 137374
rect 98782 137138 98866 137374
rect 99102 137138 135746 137374
rect 135982 137138 136066 137374
rect 136302 137138 172946 137374
rect 173182 137138 173266 137374
rect 173502 137138 210146 137374
rect 210382 137138 210466 137374
rect 210702 137138 247346 137374
rect 247582 137138 247666 137374
rect 247902 137138 284546 137374
rect 284782 137138 284866 137374
rect 285102 137138 321746 137374
rect 321982 137138 322066 137374
rect 322302 137138 358946 137374
rect 359182 137138 359266 137374
rect 359502 137138 396146 137374
rect 396382 137138 396466 137374
rect 396702 137138 433346 137374
rect 433582 137138 433666 137374
rect 433902 137138 470546 137374
rect 470782 137138 470866 137374
rect 471102 137138 507746 137374
rect 507982 137138 508066 137374
rect 508302 137138 544946 137374
rect 545182 137138 545266 137374
rect 545502 137138 582146 137374
rect 582382 137138 582466 137374
rect 582702 137138 582820 137374
rect 1104 137054 582820 137138
rect 1104 136818 24146 137054
rect 24382 136818 24466 137054
rect 24702 136818 61346 137054
rect 61582 136818 61666 137054
rect 61902 136818 98546 137054
rect 98782 136818 98866 137054
rect 99102 136818 135746 137054
rect 135982 136818 136066 137054
rect 136302 136818 172946 137054
rect 173182 136818 173266 137054
rect 173502 136818 210146 137054
rect 210382 136818 210466 137054
rect 210702 136818 247346 137054
rect 247582 136818 247666 137054
rect 247902 136818 284546 137054
rect 284782 136818 284866 137054
rect 285102 136818 321746 137054
rect 321982 136818 322066 137054
rect 322302 136818 358946 137054
rect 359182 136818 359266 137054
rect 359502 136818 396146 137054
rect 396382 136818 396466 137054
rect 396702 136818 433346 137054
rect 433582 136818 433666 137054
rect 433902 136818 470546 137054
rect 470782 136818 470866 137054
rect 471102 136818 507746 137054
rect 507982 136818 508066 137054
rect 508302 136818 544946 137054
rect 545182 136818 545266 137054
rect 545502 136818 582146 137054
rect 582382 136818 582466 137054
rect 582702 136818 582820 137054
rect 1104 136786 582820 136818
rect 1104 133654 582820 133686
rect 1104 133418 20426 133654
rect 20662 133418 20746 133654
rect 20982 133418 57626 133654
rect 57862 133418 57946 133654
rect 58182 133418 94826 133654
rect 95062 133418 95146 133654
rect 95382 133418 132026 133654
rect 132262 133418 132346 133654
rect 132582 133418 169226 133654
rect 169462 133418 169546 133654
rect 169782 133418 206426 133654
rect 206662 133418 206746 133654
rect 206982 133418 243626 133654
rect 243862 133418 243946 133654
rect 244182 133418 280826 133654
rect 281062 133418 281146 133654
rect 281382 133418 318026 133654
rect 318262 133418 318346 133654
rect 318582 133418 355226 133654
rect 355462 133418 355546 133654
rect 355782 133418 392426 133654
rect 392662 133418 392746 133654
rect 392982 133418 429626 133654
rect 429862 133418 429946 133654
rect 430182 133418 466826 133654
rect 467062 133418 467146 133654
rect 467382 133418 504026 133654
rect 504262 133418 504346 133654
rect 504582 133418 541226 133654
rect 541462 133418 541546 133654
rect 541782 133418 578426 133654
rect 578662 133418 578746 133654
rect 578982 133418 582820 133654
rect 1104 133334 582820 133418
rect 1104 133098 20426 133334
rect 20662 133098 20746 133334
rect 20982 133098 57626 133334
rect 57862 133098 57946 133334
rect 58182 133098 94826 133334
rect 95062 133098 95146 133334
rect 95382 133098 132026 133334
rect 132262 133098 132346 133334
rect 132582 133098 169226 133334
rect 169462 133098 169546 133334
rect 169782 133098 206426 133334
rect 206662 133098 206746 133334
rect 206982 133098 243626 133334
rect 243862 133098 243946 133334
rect 244182 133098 280826 133334
rect 281062 133098 281146 133334
rect 281382 133098 318026 133334
rect 318262 133098 318346 133334
rect 318582 133098 355226 133334
rect 355462 133098 355546 133334
rect 355782 133098 392426 133334
rect 392662 133098 392746 133334
rect 392982 133098 429626 133334
rect 429862 133098 429946 133334
rect 430182 133098 466826 133334
rect 467062 133098 467146 133334
rect 467382 133098 504026 133334
rect 504262 133098 504346 133334
rect 504582 133098 541226 133334
rect 541462 133098 541546 133334
rect 541782 133098 578426 133334
rect 578662 133098 578746 133334
rect 578982 133098 582820 133334
rect 1104 133066 582820 133098
rect 1104 129934 582820 129966
rect 1104 129698 16706 129934
rect 16942 129698 17026 129934
rect 17262 129698 53906 129934
rect 54142 129698 54226 129934
rect 54462 129698 91106 129934
rect 91342 129698 91426 129934
rect 91662 129698 128306 129934
rect 128542 129698 128626 129934
rect 128862 129698 165506 129934
rect 165742 129698 165826 129934
rect 166062 129698 202706 129934
rect 202942 129698 203026 129934
rect 203262 129698 239906 129934
rect 240142 129698 240226 129934
rect 240462 129698 277106 129934
rect 277342 129698 277426 129934
rect 277662 129698 314306 129934
rect 314542 129698 314626 129934
rect 314862 129698 351506 129934
rect 351742 129698 351826 129934
rect 352062 129698 388706 129934
rect 388942 129698 389026 129934
rect 389262 129698 425906 129934
rect 426142 129698 426226 129934
rect 426462 129698 463106 129934
rect 463342 129698 463426 129934
rect 463662 129698 500306 129934
rect 500542 129698 500626 129934
rect 500862 129698 537506 129934
rect 537742 129698 537826 129934
rect 538062 129698 574706 129934
rect 574942 129698 575026 129934
rect 575262 129698 582820 129934
rect 1104 129614 582820 129698
rect 1104 129378 16706 129614
rect 16942 129378 17026 129614
rect 17262 129378 53906 129614
rect 54142 129378 54226 129614
rect 54462 129378 91106 129614
rect 91342 129378 91426 129614
rect 91662 129378 128306 129614
rect 128542 129378 128626 129614
rect 128862 129378 165506 129614
rect 165742 129378 165826 129614
rect 166062 129378 202706 129614
rect 202942 129378 203026 129614
rect 203262 129378 239906 129614
rect 240142 129378 240226 129614
rect 240462 129378 277106 129614
rect 277342 129378 277426 129614
rect 277662 129378 314306 129614
rect 314542 129378 314626 129614
rect 314862 129378 351506 129614
rect 351742 129378 351826 129614
rect 352062 129378 388706 129614
rect 388942 129378 389026 129614
rect 389262 129378 425906 129614
rect 426142 129378 426226 129614
rect 426462 129378 463106 129614
rect 463342 129378 463426 129614
rect 463662 129378 500306 129614
rect 500542 129378 500626 129614
rect 500862 129378 537506 129614
rect 537742 129378 537826 129614
rect 538062 129378 574706 129614
rect 574942 129378 575026 129614
rect 575262 129378 582820 129614
rect 1104 129346 582820 129378
rect 1104 126214 582820 126246
rect 1104 125978 12986 126214
rect 13222 125978 13306 126214
rect 13542 125978 50186 126214
rect 50422 125978 50506 126214
rect 50742 125978 87386 126214
rect 87622 125978 87706 126214
rect 87942 125978 124586 126214
rect 124822 125978 124906 126214
rect 125142 125978 161786 126214
rect 162022 125978 162106 126214
rect 162342 125978 198986 126214
rect 199222 125978 199306 126214
rect 199542 125978 236186 126214
rect 236422 125978 236506 126214
rect 236742 125978 273386 126214
rect 273622 125978 273706 126214
rect 273942 125978 310586 126214
rect 310822 125978 310906 126214
rect 311142 125978 347786 126214
rect 348022 125978 348106 126214
rect 348342 125978 384986 126214
rect 385222 125978 385306 126214
rect 385542 125978 422186 126214
rect 422422 125978 422506 126214
rect 422742 125978 459386 126214
rect 459622 125978 459706 126214
rect 459942 125978 496586 126214
rect 496822 125978 496906 126214
rect 497142 125978 533786 126214
rect 534022 125978 534106 126214
rect 534342 125978 570986 126214
rect 571222 125978 571306 126214
rect 571542 125978 582820 126214
rect 1104 125894 582820 125978
rect 1104 125658 12986 125894
rect 13222 125658 13306 125894
rect 13542 125658 50186 125894
rect 50422 125658 50506 125894
rect 50742 125658 87386 125894
rect 87622 125658 87706 125894
rect 87942 125658 124586 125894
rect 124822 125658 124906 125894
rect 125142 125658 161786 125894
rect 162022 125658 162106 125894
rect 162342 125658 198986 125894
rect 199222 125658 199306 125894
rect 199542 125658 236186 125894
rect 236422 125658 236506 125894
rect 236742 125658 273386 125894
rect 273622 125658 273706 125894
rect 273942 125658 310586 125894
rect 310822 125658 310906 125894
rect 311142 125658 347786 125894
rect 348022 125658 348106 125894
rect 348342 125658 384986 125894
rect 385222 125658 385306 125894
rect 385542 125658 422186 125894
rect 422422 125658 422506 125894
rect 422742 125658 459386 125894
rect 459622 125658 459706 125894
rect 459942 125658 496586 125894
rect 496822 125658 496906 125894
rect 497142 125658 533786 125894
rect 534022 125658 534106 125894
rect 534342 125658 570986 125894
rect 571222 125658 571306 125894
rect 571542 125658 582820 125894
rect 1104 125626 582820 125658
rect 1104 122494 582820 122526
rect 1104 122258 9266 122494
rect 9502 122258 9586 122494
rect 9822 122258 46466 122494
rect 46702 122258 46786 122494
rect 47022 122258 83666 122494
rect 83902 122258 83986 122494
rect 84222 122258 120866 122494
rect 121102 122258 121186 122494
rect 121422 122258 158066 122494
rect 158302 122258 158386 122494
rect 158622 122258 195266 122494
rect 195502 122258 195586 122494
rect 195822 122258 232466 122494
rect 232702 122258 232786 122494
rect 233022 122258 269666 122494
rect 269902 122258 269986 122494
rect 270222 122258 306866 122494
rect 307102 122258 307186 122494
rect 307422 122258 344066 122494
rect 344302 122258 344386 122494
rect 344622 122258 381266 122494
rect 381502 122258 381586 122494
rect 381822 122258 418466 122494
rect 418702 122258 418786 122494
rect 419022 122258 455666 122494
rect 455902 122258 455986 122494
rect 456222 122258 492866 122494
rect 493102 122258 493186 122494
rect 493422 122258 530066 122494
rect 530302 122258 530386 122494
rect 530622 122258 567266 122494
rect 567502 122258 567586 122494
rect 567822 122258 582820 122494
rect 1104 122174 582820 122258
rect 1104 121938 9266 122174
rect 9502 121938 9586 122174
rect 9822 121938 46466 122174
rect 46702 121938 46786 122174
rect 47022 121938 83666 122174
rect 83902 121938 83986 122174
rect 84222 121938 120866 122174
rect 121102 121938 121186 122174
rect 121422 121938 158066 122174
rect 158302 121938 158386 122174
rect 158622 121938 195266 122174
rect 195502 121938 195586 122174
rect 195822 121938 232466 122174
rect 232702 121938 232786 122174
rect 233022 121938 269666 122174
rect 269902 121938 269986 122174
rect 270222 121938 306866 122174
rect 307102 121938 307186 122174
rect 307422 121938 344066 122174
rect 344302 121938 344386 122174
rect 344622 121938 381266 122174
rect 381502 121938 381586 122174
rect 381822 121938 418466 122174
rect 418702 121938 418786 122174
rect 419022 121938 455666 122174
rect 455902 121938 455986 122174
rect 456222 121938 492866 122174
rect 493102 121938 493186 122174
rect 493422 121938 530066 122174
rect 530302 121938 530386 122174
rect 530622 121938 567266 122174
rect 567502 121938 567586 122174
rect 567822 121938 582820 122174
rect 1104 121906 582820 121938
rect 1104 118774 582820 118806
rect 1104 118538 5546 118774
rect 5782 118538 5866 118774
rect 6102 118538 42746 118774
rect 42982 118538 43066 118774
rect 43302 118538 79946 118774
rect 80182 118538 80266 118774
rect 80502 118538 117146 118774
rect 117382 118538 117466 118774
rect 117702 118538 154346 118774
rect 154582 118538 154666 118774
rect 154902 118538 191546 118774
rect 191782 118538 191866 118774
rect 192102 118538 228746 118774
rect 228982 118538 229066 118774
rect 229302 118538 265946 118774
rect 266182 118538 266266 118774
rect 266502 118538 303146 118774
rect 303382 118538 303466 118774
rect 303702 118538 340346 118774
rect 340582 118538 340666 118774
rect 340902 118538 377546 118774
rect 377782 118538 377866 118774
rect 378102 118538 414746 118774
rect 414982 118538 415066 118774
rect 415302 118538 451946 118774
rect 452182 118538 452266 118774
rect 452502 118538 489146 118774
rect 489382 118538 489466 118774
rect 489702 118538 526346 118774
rect 526582 118538 526666 118774
rect 526902 118538 563546 118774
rect 563782 118538 563866 118774
rect 564102 118538 582820 118774
rect 1104 118454 582820 118538
rect 1104 118218 5546 118454
rect 5782 118218 5866 118454
rect 6102 118218 42746 118454
rect 42982 118218 43066 118454
rect 43302 118218 79946 118454
rect 80182 118218 80266 118454
rect 80502 118218 117146 118454
rect 117382 118218 117466 118454
rect 117702 118218 154346 118454
rect 154582 118218 154666 118454
rect 154902 118218 191546 118454
rect 191782 118218 191866 118454
rect 192102 118218 228746 118454
rect 228982 118218 229066 118454
rect 229302 118218 265946 118454
rect 266182 118218 266266 118454
rect 266502 118218 303146 118454
rect 303382 118218 303466 118454
rect 303702 118218 340346 118454
rect 340582 118218 340666 118454
rect 340902 118218 377546 118454
rect 377782 118218 377866 118454
rect 378102 118218 414746 118454
rect 414982 118218 415066 118454
rect 415302 118218 451946 118454
rect 452182 118218 452266 118454
rect 452502 118218 489146 118454
rect 489382 118218 489466 118454
rect 489702 118218 526346 118454
rect 526582 118218 526666 118454
rect 526902 118218 563546 118454
rect 563782 118218 563866 118454
rect 564102 118218 582820 118454
rect 1104 118186 582820 118218
rect 1104 115054 582820 115086
rect 1104 114818 1826 115054
rect 2062 114818 2146 115054
rect 2382 114818 39026 115054
rect 39262 114818 39346 115054
rect 39582 114818 76226 115054
rect 76462 114818 76546 115054
rect 76782 114818 113426 115054
rect 113662 114818 113746 115054
rect 113982 114818 150626 115054
rect 150862 114818 150946 115054
rect 151182 114818 187826 115054
rect 188062 114818 188146 115054
rect 188382 114818 225026 115054
rect 225262 114818 225346 115054
rect 225582 114818 262226 115054
rect 262462 114818 262546 115054
rect 262782 114818 299426 115054
rect 299662 114818 299746 115054
rect 299982 114818 336626 115054
rect 336862 114818 336946 115054
rect 337182 114818 373826 115054
rect 374062 114818 374146 115054
rect 374382 114818 411026 115054
rect 411262 114818 411346 115054
rect 411582 114818 448226 115054
rect 448462 114818 448546 115054
rect 448782 114818 485426 115054
rect 485662 114818 485746 115054
rect 485982 114818 522626 115054
rect 522862 114818 522946 115054
rect 523182 114818 559826 115054
rect 560062 114818 560146 115054
rect 560382 114818 582820 115054
rect 1104 114734 582820 114818
rect 1104 114498 1826 114734
rect 2062 114498 2146 114734
rect 2382 114498 39026 114734
rect 39262 114498 39346 114734
rect 39582 114498 76226 114734
rect 76462 114498 76546 114734
rect 76782 114498 113426 114734
rect 113662 114498 113746 114734
rect 113982 114498 150626 114734
rect 150862 114498 150946 114734
rect 151182 114498 187826 114734
rect 188062 114498 188146 114734
rect 188382 114498 225026 114734
rect 225262 114498 225346 114734
rect 225582 114498 262226 114734
rect 262462 114498 262546 114734
rect 262782 114498 299426 114734
rect 299662 114498 299746 114734
rect 299982 114498 336626 114734
rect 336862 114498 336946 114734
rect 337182 114498 373826 114734
rect 374062 114498 374146 114734
rect 374382 114498 411026 114734
rect 411262 114498 411346 114734
rect 411582 114498 448226 114734
rect 448462 114498 448546 114734
rect 448782 114498 485426 114734
rect 485662 114498 485746 114734
rect 485982 114498 522626 114734
rect 522862 114498 522946 114734
rect 523182 114498 559826 114734
rect 560062 114498 560146 114734
rect 560382 114498 582820 114734
rect 1104 114466 582820 114498
rect 1104 103894 582820 103926
rect 1104 103658 27866 103894
rect 28102 103658 28186 103894
rect 28422 103658 65066 103894
rect 65302 103658 65386 103894
rect 65622 103658 102266 103894
rect 102502 103658 102586 103894
rect 102822 103658 139466 103894
rect 139702 103658 139786 103894
rect 140022 103658 176666 103894
rect 176902 103658 176986 103894
rect 177222 103658 213866 103894
rect 214102 103658 214186 103894
rect 214422 103658 251066 103894
rect 251302 103658 251386 103894
rect 251622 103658 288266 103894
rect 288502 103658 288586 103894
rect 288822 103658 325466 103894
rect 325702 103658 325786 103894
rect 326022 103658 362666 103894
rect 362902 103658 362986 103894
rect 363222 103658 399866 103894
rect 400102 103658 400186 103894
rect 400422 103658 437066 103894
rect 437302 103658 437386 103894
rect 437622 103658 474266 103894
rect 474502 103658 474586 103894
rect 474822 103658 511466 103894
rect 511702 103658 511786 103894
rect 512022 103658 548666 103894
rect 548902 103658 548986 103894
rect 549222 103658 582820 103894
rect 1104 103574 582820 103658
rect 1104 103338 27866 103574
rect 28102 103338 28186 103574
rect 28422 103338 65066 103574
rect 65302 103338 65386 103574
rect 65622 103338 102266 103574
rect 102502 103338 102586 103574
rect 102822 103338 139466 103574
rect 139702 103338 139786 103574
rect 140022 103338 176666 103574
rect 176902 103338 176986 103574
rect 177222 103338 213866 103574
rect 214102 103338 214186 103574
rect 214422 103338 251066 103574
rect 251302 103338 251386 103574
rect 251622 103338 288266 103574
rect 288502 103338 288586 103574
rect 288822 103338 325466 103574
rect 325702 103338 325786 103574
rect 326022 103338 362666 103574
rect 362902 103338 362986 103574
rect 363222 103338 399866 103574
rect 400102 103338 400186 103574
rect 400422 103338 437066 103574
rect 437302 103338 437386 103574
rect 437622 103338 474266 103574
rect 474502 103338 474586 103574
rect 474822 103338 511466 103574
rect 511702 103338 511786 103574
rect 512022 103338 548666 103574
rect 548902 103338 548986 103574
rect 549222 103338 582820 103574
rect 1104 103306 582820 103338
rect 1104 100174 582820 100206
rect 1104 99938 24146 100174
rect 24382 99938 24466 100174
rect 24702 99938 61346 100174
rect 61582 99938 61666 100174
rect 61902 99938 98546 100174
rect 98782 99938 98866 100174
rect 99102 99938 135746 100174
rect 135982 99938 136066 100174
rect 136302 99938 172946 100174
rect 173182 99938 173266 100174
rect 173502 99938 210146 100174
rect 210382 99938 210466 100174
rect 210702 99938 247346 100174
rect 247582 99938 247666 100174
rect 247902 99938 284546 100174
rect 284782 99938 284866 100174
rect 285102 99938 321746 100174
rect 321982 99938 322066 100174
rect 322302 99938 358946 100174
rect 359182 99938 359266 100174
rect 359502 99938 396146 100174
rect 396382 99938 396466 100174
rect 396702 99938 433346 100174
rect 433582 99938 433666 100174
rect 433902 99938 470546 100174
rect 470782 99938 470866 100174
rect 471102 99938 507746 100174
rect 507982 99938 508066 100174
rect 508302 99938 544946 100174
rect 545182 99938 545266 100174
rect 545502 99938 582146 100174
rect 582382 99938 582466 100174
rect 582702 99938 582820 100174
rect 1104 99854 582820 99938
rect 1104 99618 24146 99854
rect 24382 99618 24466 99854
rect 24702 99618 61346 99854
rect 61582 99618 61666 99854
rect 61902 99618 98546 99854
rect 98782 99618 98866 99854
rect 99102 99618 135746 99854
rect 135982 99618 136066 99854
rect 136302 99618 172946 99854
rect 173182 99618 173266 99854
rect 173502 99618 210146 99854
rect 210382 99618 210466 99854
rect 210702 99618 247346 99854
rect 247582 99618 247666 99854
rect 247902 99618 284546 99854
rect 284782 99618 284866 99854
rect 285102 99618 321746 99854
rect 321982 99618 322066 99854
rect 322302 99618 358946 99854
rect 359182 99618 359266 99854
rect 359502 99618 396146 99854
rect 396382 99618 396466 99854
rect 396702 99618 433346 99854
rect 433582 99618 433666 99854
rect 433902 99618 470546 99854
rect 470782 99618 470866 99854
rect 471102 99618 507746 99854
rect 507982 99618 508066 99854
rect 508302 99618 544946 99854
rect 545182 99618 545266 99854
rect 545502 99618 582146 99854
rect 582382 99618 582466 99854
rect 582702 99618 582820 99854
rect 1104 99586 582820 99618
rect 1104 96454 582820 96486
rect 1104 96218 20426 96454
rect 20662 96218 20746 96454
rect 20982 96218 57626 96454
rect 57862 96218 57946 96454
rect 58182 96218 94826 96454
rect 95062 96218 95146 96454
rect 95382 96218 132026 96454
rect 132262 96218 132346 96454
rect 132582 96218 169226 96454
rect 169462 96218 169546 96454
rect 169782 96218 206426 96454
rect 206662 96218 206746 96454
rect 206982 96218 243626 96454
rect 243862 96218 243946 96454
rect 244182 96218 280826 96454
rect 281062 96218 281146 96454
rect 281382 96218 318026 96454
rect 318262 96218 318346 96454
rect 318582 96218 355226 96454
rect 355462 96218 355546 96454
rect 355782 96218 392426 96454
rect 392662 96218 392746 96454
rect 392982 96218 429626 96454
rect 429862 96218 429946 96454
rect 430182 96218 466826 96454
rect 467062 96218 467146 96454
rect 467382 96218 504026 96454
rect 504262 96218 504346 96454
rect 504582 96218 541226 96454
rect 541462 96218 541546 96454
rect 541782 96218 578426 96454
rect 578662 96218 578746 96454
rect 578982 96218 582820 96454
rect 1104 96134 582820 96218
rect 1104 95898 20426 96134
rect 20662 95898 20746 96134
rect 20982 95898 57626 96134
rect 57862 95898 57946 96134
rect 58182 95898 94826 96134
rect 95062 95898 95146 96134
rect 95382 95898 132026 96134
rect 132262 95898 132346 96134
rect 132582 95898 169226 96134
rect 169462 95898 169546 96134
rect 169782 95898 206426 96134
rect 206662 95898 206746 96134
rect 206982 95898 243626 96134
rect 243862 95898 243946 96134
rect 244182 95898 280826 96134
rect 281062 95898 281146 96134
rect 281382 95898 318026 96134
rect 318262 95898 318346 96134
rect 318582 95898 355226 96134
rect 355462 95898 355546 96134
rect 355782 95898 392426 96134
rect 392662 95898 392746 96134
rect 392982 95898 429626 96134
rect 429862 95898 429946 96134
rect 430182 95898 466826 96134
rect 467062 95898 467146 96134
rect 467382 95898 504026 96134
rect 504262 95898 504346 96134
rect 504582 95898 541226 96134
rect 541462 95898 541546 96134
rect 541782 95898 578426 96134
rect 578662 95898 578746 96134
rect 578982 95898 582820 96134
rect 1104 95866 582820 95898
rect 1104 92734 582820 92766
rect 1104 92498 16706 92734
rect 16942 92498 17026 92734
rect 17262 92498 53906 92734
rect 54142 92498 54226 92734
rect 54462 92498 91106 92734
rect 91342 92498 91426 92734
rect 91662 92498 128306 92734
rect 128542 92498 128626 92734
rect 128862 92498 165506 92734
rect 165742 92498 165826 92734
rect 166062 92498 202706 92734
rect 202942 92498 203026 92734
rect 203262 92498 239906 92734
rect 240142 92498 240226 92734
rect 240462 92498 277106 92734
rect 277342 92498 277426 92734
rect 277662 92498 314306 92734
rect 314542 92498 314626 92734
rect 314862 92498 351506 92734
rect 351742 92498 351826 92734
rect 352062 92498 388706 92734
rect 388942 92498 389026 92734
rect 389262 92498 425906 92734
rect 426142 92498 426226 92734
rect 426462 92498 463106 92734
rect 463342 92498 463426 92734
rect 463662 92498 500306 92734
rect 500542 92498 500626 92734
rect 500862 92498 537506 92734
rect 537742 92498 537826 92734
rect 538062 92498 574706 92734
rect 574942 92498 575026 92734
rect 575262 92498 582820 92734
rect 1104 92414 582820 92498
rect 1104 92178 16706 92414
rect 16942 92178 17026 92414
rect 17262 92178 53906 92414
rect 54142 92178 54226 92414
rect 54462 92178 91106 92414
rect 91342 92178 91426 92414
rect 91662 92178 128306 92414
rect 128542 92178 128626 92414
rect 128862 92178 165506 92414
rect 165742 92178 165826 92414
rect 166062 92178 202706 92414
rect 202942 92178 203026 92414
rect 203262 92178 239906 92414
rect 240142 92178 240226 92414
rect 240462 92178 277106 92414
rect 277342 92178 277426 92414
rect 277662 92178 314306 92414
rect 314542 92178 314626 92414
rect 314862 92178 351506 92414
rect 351742 92178 351826 92414
rect 352062 92178 388706 92414
rect 388942 92178 389026 92414
rect 389262 92178 425906 92414
rect 426142 92178 426226 92414
rect 426462 92178 463106 92414
rect 463342 92178 463426 92414
rect 463662 92178 500306 92414
rect 500542 92178 500626 92414
rect 500862 92178 537506 92414
rect 537742 92178 537826 92414
rect 538062 92178 574706 92414
rect 574942 92178 575026 92414
rect 575262 92178 582820 92414
rect 1104 92146 582820 92178
rect 1104 89014 582820 89046
rect 1104 88778 12986 89014
rect 13222 88778 13306 89014
rect 13542 88778 50186 89014
rect 50422 88778 50506 89014
rect 50742 88778 87386 89014
rect 87622 88778 87706 89014
rect 87942 88778 124586 89014
rect 124822 88778 124906 89014
rect 125142 88778 161786 89014
rect 162022 88778 162106 89014
rect 162342 88778 198986 89014
rect 199222 88778 199306 89014
rect 199542 88778 236186 89014
rect 236422 88778 236506 89014
rect 236742 88778 273386 89014
rect 273622 88778 273706 89014
rect 273942 88778 310586 89014
rect 310822 88778 310906 89014
rect 311142 88778 347786 89014
rect 348022 88778 348106 89014
rect 348342 88778 384986 89014
rect 385222 88778 385306 89014
rect 385542 88778 422186 89014
rect 422422 88778 422506 89014
rect 422742 88778 459386 89014
rect 459622 88778 459706 89014
rect 459942 88778 496586 89014
rect 496822 88778 496906 89014
rect 497142 88778 533786 89014
rect 534022 88778 534106 89014
rect 534342 88778 570986 89014
rect 571222 88778 571306 89014
rect 571542 88778 582820 89014
rect 1104 88694 582820 88778
rect 1104 88458 12986 88694
rect 13222 88458 13306 88694
rect 13542 88458 50186 88694
rect 50422 88458 50506 88694
rect 50742 88458 87386 88694
rect 87622 88458 87706 88694
rect 87942 88458 124586 88694
rect 124822 88458 124906 88694
rect 125142 88458 161786 88694
rect 162022 88458 162106 88694
rect 162342 88458 198986 88694
rect 199222 88458 199306 88694
rect 199542 88458 236186 88694
rect 236422 88458 236506 88694
rect 236742 88458 273386 88694
rect 273622 88458 273706 88694
rect 273942 88458 310586 88694
rect 310822 88458 310906 88694
rect 311142 88458 347786 88694
rect 348022 88458 348106 88694
rect 348342 88458 384986 88694
rect 385222 88458 385306 88694
rect 385542 88458 422186 88694
rect 422422 88458 422506 88694
rect 422742 88458 459386 88694
rect 459622 88458 459706 88694
rect 459942 88458 496586 88694
rect 496822 88458 496906 88694
rect 497142 88458 533786 88694
rect 534022 88458 534106 88694
rect 534342 88458 570986 88694
rect 571222 88458 571306 88694
rect 571542 88458 582820 88694
rect 1104 88426 582820 88458
rect 1104 85294 582820 85326
rect 1104 85058 9266 85294
rect 9502 85058 9586 85294
rect 9822 85058 46466 85294
rect 46702 85058 46786 85294
rect 47022 85058 83666 85294
rect 83902 85058 83986 85294
rect 84222 85058 120866 85294
rect 121102 85058 121186 85294
rect 121422 85058 158066 85294
rect 158302 85058 158386 85294
rect 158622 85058 195266 85294
rect 195502 85058 195586 85294
rect 195822 85058 232466 85294
rect 232702 85058 232786 85294
rect 233022 85058 269666 85294
rect 269902 85058 269986 85294
rect 270222 85058 306866 85294
rect 307102 85058 307186 85294
rect 307422 85058 344066 85294
rect 344302 85058 344386 85294
rect 344622 85058 381266 85294
rect 381502 85058 381586 85294
rect 381822 85058 418466 85294
rect 418702 85058 418786 85294
rect 419022 85058 455666 85294
rect 455902 85058 455986 85294
rect 456222 85058 492866 85294
rect 493102 85058 493186 85294
rect 493422 85058 530066 85294
rect 530302 85058 530386 85294
rect 530622 85058 567266 85294
rect 567502 85058 567586 85294
rect 567822 85058 582820 85294
rect 1104 84974 582820 85058
rect 1104 84738 9266 84974
rect 9502 84738 9586 84974
rect 9822 84738 46466 84974
rect 46702 84738 46786 84974
rect 47022 84738 83666 84974
rect 83902 84738 83986 84974
rect 84222 84738 120866 84974
rect 121102 84738 121186 84974
rect 121422 84738 158066 84974
rect 158302 84738 158386 84974
rect 158622 84738 195266 84974
rect 195502 84738 195586 84974
rect 195822 84738 232466 84974
rect 232702 84738 232786 84974
rect 233022 84738 269666 84974
rect 269902 84738 269986 84974
rect 270222 84738 306866 84974
rect 307102 84738 307186 84974
rect 307422 84738 344066 84974
rect 344302 84738 344386 84974
rect 344622 84738 381266 84974
rect 381502 84738 381586 84974
rect 381822 84738 418466 84974
rect 418702 84738 418786 84974
rect 419022 84738 455666 84974
rect 455902 84738 455986 84974
rect 456222 84738 492866 84974
rect 493102 84738 493186 84974
rect 493422 84738 530066 84974
rect 530302 84738 530386 84974
rect 530622 84738 567266 84974
rect 567502 84738 567586 84974
rect 567822 84738 582820 84974
rect 1104 84706 582820 84738
rect 1104 81574 582820 81606
rect 1104 81338 5546 81574
rect 5782 81338 5866 81574
rect 6102 81338 42746 81574
rect 42982 81338 43066 81574
rect 43302 81338 79946 81574
rect 80182 81338 80266 81574
rect 80502 81338 117146 81574
rect 117382 81338 117466 81574
rect 117702 81338 154346 81574
rect 154582 81338 154666 81574
rect 154902 81338 191546 81574
rect 191782 81338 191866 81574
rect 192102 81338 228746 81574
rect 228982 81338 229066 81574
rect 229302 81338 265946 81574
rect 266182 81338 266266 81574
rect 266502 81338 303146 81574
rect 303382 81338 303466 81574
rect 303702 81338 340346 81574
rect 340582 81338 340666 81574
rect 340902 81338 377546 81574
rect 377782 81338 377866 81574
rect 378102 81338 414746 81574
rect 414982 81338 415066 81574
rect 415302 81338 451946 81574
rect 452182 81338 452266 81574
rect 452502 81338 489146 81574
rect 489382 81338 489466 81574
rect 489702 81338 526346 81574
rect 526582 81338 526666 81574
rect 526902 81338 563546 81574
rect 563782 81338 563866 81574
rect 564102 81338 582820 81574
rect 1104 81254 582820 81338
rect 1104 81018 5546 81254
rect 5782 81018 5866 81254
rect 6102 81018 42746 81254
rect 42982 81018 43066 81254
rect 43302 81018 79946 81254
rect 80182 81018 80266 81254
rect 80502 81018 117146 81254
rect 117382 81018 117466 81254
rect 117702 81018 154346 81254
rect 154582 81018 154666 81254
rect 154902 81018 191546 81254
rect 191782 81018 191866 81254
rect 192102 81018 228746 81254
rect 228982 81018 229066 81254
rect 229302 81018 265946 81254
rect 266182 81018 266266 81254
rect 266502 81018 303146 81254
rect 303382 81018 303466 81254
rect 303702 81018 340346 81254
rect 340582 81018 340666 81254
rect 340902 81018 377546 81254
rect 377782 81018 377866 81254
rect 378102 81018 414746 81254
rect 414982 81018 415066 81254
rect 415302 81018 451946 81254
rect 452182 81018 452266 81254
rect 452502 81018 489146 81254
rect 489382 81018 489466 81254
rect 489702 81018 526346 81254
rect 526582 81018 526666 81254
rect 526902 81018 563546 81254
rect 563782 81018 563866 81254
rect 564102 81018 582820 81254
rect 1104 80986 582820 81018
rect 1104 77854 582820 77886
rect 1104 77618 1826 77854
rect 2062 77618 2146 77854
rect 2382 77618 39026 77854
rect 39262 77618 39346 77854
rect 39582 77618 76226 77854
rect 76462 77618 76546 77854
rect 76782 77618 113426 77854
rect 113662 77618 113746 77854
rect 113982 77618 150626 77854
rect 150862 77618 150946 77854
rect 151182 77618 187826 77854
rect 188062 77618 188146 77854
rect 188382 77618 225026 77854
rect 225262 77618 225346 77854
rect 225582 77618 262226 77854
rect 262462 77618 262546 77854
rect 262782 77618 299426 77854
rect 299662 77618 299746 77854
rect 299982 77618 336626 77854
rect 336862 77618 336946 77854
rect 337182 77618 373826 77854
rect 374062 77618 374146 77854
rect 374382 77618 411026 77854
rect 411262 77618 411346 77854
rect 411582 77618 448226 77854
rect 448462 77618 448546 77854
rect 448782 77618 485426 77854
rect 485662 77618 485746 77854
rect 485982 77618 522626 77854
rect 522862 77618 522946 77854
rect 523182 77618 559826 77854
rect 560062 77618 560146 77854
rect 560382 77618 582820 77854
rect 1104 77534 582820 77618
rect 1104 77298 1826 77534
rect 2062 77298 2146 77534
rect 2382 77298 39026 77534
rect 39262 77298 39346 77534
rect 39582 77298 76226 77534
rect 76462 77298 76546 77534
rect 76782 77298 113426 77534
rect 113662 77298 113746 77534
rect 113982 77298 150626 77534
rect 150862 77298 150946 77534
rect 151182 77298 187826 77534
rect 188062 77298 188146 77534
rect 188382 77298 225026 77534
rect 225262 77298 225346 77534
rect 225582 77298 262226 77534
rect 262462 77298 262546 77534
rect 262782 77298 299426 77534
rect 299662 77298 299746 77534
rect 299982 77298 336626 77534
rect 336862 77298 336946 77534
rect 337182 77298 373826 77534
rect 374062 77298 374146 77534
rect 374382 77298 411026 77534
rect 411262 77298 411346 77534
rect 411582 77298 448226 77534
rect 448462 77298 448546 77534
rect 448782 77298 485426 77534
rect 485662 77298 485746 77534
rect 485982 77298 522626 77534
rect 522862 77298 522946 77534
rect 523182 77298 559826 77534
rect 560062 77298 560146 77534
rect 560382 77298 582820 77534
rect 1104 77266 582820 77298
rect 1104 66694 582820 66726
rect 1104 66458 27866 66694
rect 28102 66458 28186 66694
rect 28422 66458 65066 66694
rect 65302 66458 65386 66694
rect 65622 66458 102266 66694
rect 102502 66458 102586 66694
rect 102822 66458 139466 66694
rect 139702 66458 139786 66694
rect 140022 66458 176666 66694
rect 176902 66458 176986 66694
rect 177222 66458 213866 66694
rect 214102 66458 214186 66694
rect 214422 66458 251066 66694
rect 251302 66458 251386 66694
rect 251622 66458 288266 66694
rect 288502 66458 288586 66694
rect 288822 66458 325466 66694
rect 325702 66458 325786 66694
rect 326022 66458 362666 66694
rect 362902 66458 362986 66694
rect 363222 66458 399866 66694
rect 400102 66458 400186 66694
rect 400422 66458 437066 66694
rect 437302 66458 437386 66694
rect 437622 66458 474266 66694
rect 474502 66458 474586 66694
rect 474822 66458 511466 66694
rect 511702 66458 511786 66694
rect 512022 66458 548666 66694
rect 548902 66458 548986 66694
rect 549222 66458 582820 66694
rect 1104 66374 582820 66458
rect 1104 66138 27866 66374
rect 28102 66138 28186 66374
rect 28422 66138 65066 66374
rect 65302 66138 65386 66374
rect 65622 66138 102266 66374
rect 102502 66138 102586 66374
rect 102822 66138 139466 66374
rect 139702 66138 139786 66374
rect 140022 66138 176666 66374
rect 176902 66138 176986 66374
rect 177222 66138 213866 66374
rect 214102 66138 214186 66374
rect 214422 66138 251066 66374
rect 251302 66138 251386 66374
rect 251622 66138 288266 66374
rect 288502 66138 288586 66374
rect 288822 66138 325466 66374
rect 325702 66138 325786 66374
rect 326022 66138 362666 66374
rect 362902 66138 362986 66374
rect 363222 66138 399866 66374
rect 400102 66138 400186 66374
rect 400422 66138 437066 66374
rect 437302 66138 437386 66374
rect 437622 66138 474266 66374
rect 474502 66138 474586 66374
rect 474822 66138 511466 66374
rect 511702 66138 511786 66374
rect 512022 66138 548666 66374
rect 548902 66138 548986 66374
rect 549222 66138 582820 66374
rect 1104 66106 582820 66138
rect 1104 62974 582820 63006
rect 1104 62738 24146 62974
rect 24382 62738 24466 62974
rect 24702 62738 61346 62974
rect 61582 62738 61666 62974
rect 61902 62738 98546 62974
rect 98782 62738 98866 62974
rect 99102 62738 135746 62974
rect 135982 62738 136066 62974
rect 136302 62738 172946 62974
rect 173182 62738 173266 62974
rect 173502 62738 210146 62974
rect 210382 62738 210466 62974
rect 210702 62738 247346 62974
rect 247582 62738 247666 62974
rect 247902 62738 284546 62974
rect 284782 62738 284866 62974
rect 285102 62738 321746 62974
rect 321982 62738 322066 62974
rect 322302 62738 358946 62974
rect 359182 62738 359266 62974
rect 359502 62738 396146 62974
rect 396382 62738 396466 62974
rect 396702 62738 433346 62974
rect 433582 62738 433666 62974
rect 433902 62738 470546 62974
rect 470782 62738 470866 62974
rect 471102 62738 507746 62974
rect 507982 62738 508066 62974
rect 508302 62738 544946 62974
rect 545182 62738 545266 62974
rect 545502 62738 582146 62974
rect 582382 62738 582466 62974
rect 582702 62738 582820 62974
rect 1104 62654 582820 62738
rect 1104 62418 24146 62654
rect 24382 62418 24466 62654
rect 24702 62418 61346 62654
rect 61582 62418 61666 62654
rect 61902 62418 98546 62654
rect 98782 62418 98866 62654
rect 99102 62418 135746 62654
rect 135982 62418 136066 62654
rect 136302 62418 172946 62654
rect 173182 62418 173266 62654
rect 173502 62418 210146 62654
rect 210382 62418 210466 62654
rect 210702 62418 247346 62654
rect 247582 62418 247666 62654
rect 247902 62418 284546 62654
rect 284782 62418 284866 62654
rect 285102 62418 321746 62654
rect 321982 62418 322066 62654
rect 322302 62418 358946 62654
rect 359182 62418 359266 62654
rect 359502 62418 396146 62654
rect 396382 62418 396466 62654
rect 396702 62418 433346 62654
rect 433582 62418 433666 62654
rect 433902 62418 470546 62654
rect 470782 62418 470866 62654
rect 471102 62418 507746 62654
rect 507982 62418 508066 62654
rect 508302 62418 544946 62654
rect 545182 62418 545266 62654
rect 545502 62418 582146 62654
rect 582382 62418 582466 62654
rect 582702 62418 582820 62654
rect 1104 62386 582820 62418
rect 1104 59254 582820 59286
rect 1104 59018 20426 59254
rect 20662 59018 20746 59254
rect 20982 59018 57626 59254
rect 57862 59018 57946 59254
rect 58182 59018 94826 59254
rect 95062 59018 95146 59254
rect 95382 59018 132026 59254
rect 132262 59018 132346 59254
rect 132582 59018 169226 59254
rect 169462 59018 169546 59254
rect 169782 59018 206426 59254
rect 206662 59018 206746 59254
rect 206982 59018 243626 59254
rect 243862 59018 243946 59254
rect 244182 59018 280826 59254
rect 281062 59018 281146 59254
rect 281382 59018 318026 59254
rect 318262 59018 318346 59254
rect 318582 59018 355226 59254
rect 355462 59018 355546 59254
rect 355782 59018 392426 59254
rect 392662 59018 392746 59254
rect 392982 59018 429626 59254
rect 429862 59018 429946 59254
rect 430182 59018 466826 59254
rect 467062 59018 467146 59254
rect 467382 59018 504026 59254
rect 504262 59018 504346 59254
rect 504582 59018 541226 59254
rect 541462 59018 541546 59254
rect 541782 59018 578426 59254
rect 578662 59018 578746 59254
rect 578982 59018 582820 59254
rect 1104 58934 582820 59018
rect 1104 58698 20426 58934
rect 20662 58698 20746 58934
rect 20982 58698 57626 58934
rect 57862 58698 57946 58934
rect 58182 58698 94826 58934
rect 95062 58698 95146 58934
rect 95382 58698 132026 58934
rect 132262 58698 132346 58934
rect 132582 58698 169226 58934
rect 169462 58698 169546 58934
rect 169782 58698 206426 58934
rect 206662 58698 206746 58934
rect 206982 58698 243626 58934
rect 243862 58698 243946 58934
rect 244182 58698 280826 58934
rect 281062 58698 281146 58934
rect 281382 58698 318026 58934
rect 318262 58698 318346 58934
rect 318582 58698 355226 58934
rect 355462 58698 355546 58934
rect 355782 58698 392426 58934
rect 392662 58698 392746 58934
rect 392982 58698 429626 58934
rect 429862 58698 429946 58934
rect 430182 58698 466826 58934
rect 467062 58698 467146 58934
rect 467382 58698 504026 58934
rect 504262 58698 504346 58934
rect 504582 58698 541226 58934
rect 541462 58698 541546 58934
rect 541782 58698 578426 58934
rect 578662 58698 578746 58934
rect 578982 58698 582820 58934
rect 1104 58666 582820 58698
rect 1104 55534 582820 55566
rect 1104 55298 16706 55534
rect 16942 55298 17026 55534
rect 17262 55298 53906 55534
rect 54142 55298 54226 55534
rect 54462 55298 91106 55534
rect 91342 55298 91426 55534
rect 91662 55298 128306 55534
rect 128542 55298 128626 55534
rect 128862 55298 165506 55534
rect 165742 55298 165826 55534
rect 166062 55298 202706 55534
rect 202942 55298 203026 55534
rect 203262 55298 239906 55534
rect 240142 55298 240226 55534
rect 240462 55298 277106 55534
rect 277342 55298 277426 55534
rect 277662 55298 314306 55534
rect 314542 55298 314626 55534
rect 314862 55298 351506 55534
rect 351742 55298 351826 55534
rect 352062 55298 388706 55534
rect 388942 55298 389026 55534
rect 389262 55298 425906 55534
rect 426142 55298 426226 55534
rect 426462 55298 463106 55534
rect 463342 55298 463426 55534
rect 463662 55298 500306 55534
rect 500542 55298 500626 55534
rect 500862 55298 537506 55534
rect 537742 55298 537826 55534
rect 538062 55298 574706 55534
rect 574942 55298 575026 55534
rect 575262 55298 582820 55534
rect 1104 55214 582820 55298
rect 1104 54978 16706 55214
rect 16942 54978 17026 55214
rect 17262 54978 53906 55214
rect 54142 54978 54226 55214
rect 54462 54978 91106 55214
rect 91342 54978 91426 55214
rect 91662 54978 128306 55214
rect 128542 54978 128626 55214
rect 128862 54978 165506 55214
rect 165742 54978 165826 55214
rect 166062 54978 202706 55214
rect 202942 54978 203026 55214
rect 203262 54978 239906 55214
rect 240142 54978 240226 55214
rect 240462 54978 277106 55214
rect 277342 54978 277426 55214
rect 277662 54978 314306 55214
rect 314542 54978 314626 55214
rect 314862 54978 351506 55214
rect 351742 54978 351826 55214
rect 352062 54978 388706 55214
rect 388942 54978 389026 55214
rect 389262 54978 425906 55214
rect 426142 54978 426226 55214
rect 426462 54978 463106 55214
rect 463342 54978 463426 55214
rect 463662 54978 500306 55214
rect 500542 54978 500626 55214
rect 500862 54978 537506 55214
rect 537742 54978 537826 55214
rect 538062 54978 574706 55214
rect 574942 54978 575026 55214
rect 575262 54978 582820 55214
rect 1104 54946 582820 54978
rect 1104 51814 582820 51846
rect 1104 51578 12986 51814
rect 13222 51578 13306 51814
rect 13542 51578 50186 51814
rect 50422 51578 50506 51814
rect 50742 51578 87386 51814
rect 87622 51578 87706 51814
rect 87942 51578 124586 51814
rect 124822 51578 124906 51814
rect 125142 51578 161786 51814
rect 162022 51578 162106 51814
rect 162342 51578 198986 51814
rect 199222 51578 199306 51814
rect 199542 51578 236186 51814
rect 236422 51578 236506 51814
rect 236742 51578 273386 51814
rect 273622 51578 273706 51814
rect 273942 51578 310586 51814
rect 310822 51578 310906 51814
rect 311142 51578 347786 51814
rect 348022 51578 348106 51814
rect 348342 51578 384986 51814
rect 385222 51578 385306 51814
rect 385542 51578 422186 51814
rect 422422 51578 422506 51814
rect 422742 51578 459386 51814
rect 459622 51578 459706 51814
rect 459942 51578 496586 51814
rect 496822 51578 496906 51814
rect 497142 51578 533786 51814
rect 534022 51578 534106 51814
rect 534342 51578 570986 51814
rect 571222 51578 571306 51814
rect 571542 51578 582820 51814
rect 1104 51494 582820 51578
rect 1104 51258 12986 51494
rect 13222 51258 13306 51494
rect 13542 51258 50186 51494
rect 50422 51258 50506 51494
rect 50742 51258 87386 51494
rect 87622 51258 87706 51494
rect 87942 51258 124586 51494
rect 124822 51258 124906 51494
rect 125142 51258 161786 51494
rect 162022 51258 162106 51494
rect 162342 51258 198986 51494
rect 199222 51258 199306 51494
rect 199542 51258 236186 51494
rect 236422 51258 236506 51494
rect 236742 51258 273386 51494
rect 273622 51258 273706 51494
rect 273942 51258 310586 51494
rect 310822 51258 310906 51494
rect 311142 51258 347786 51494
rect 348022 51258 348106 51494
rect 348342 51258 384986 51494
rect 385222 51258 385306 51494
rect 385542 51258 422186 51494
rect 422422 51258 422506 51494
rect 422742 51258 459386 51494
rect 459622 51258 459706 51494
rect 459942 51258 496586 51494
rect 496822 51258 496906 51494
rect 497142 51258 533786 51494
rect 534022 51258 534106 51494
rect 534342 51258 570986 51494
rect 571222 51258 571306 51494
rect 571542 51258 582820 51494
rect 1104 51226 582820 51258
rect 1104 48094 582820 48126
rect 1104 47858 9266 48094
rect 9502 47858 9586 48094
rect 9822 47858 46466 48094
rect 46702 47858 46786 48094
rect 47022 47858 83666 48094
rect 83902 47858 83986 48094
rect 84222 47858 120866 48094
rect 121102 47858 121186 48094
rect 121422 47858 158066 48094
rect 158302 47858 158386 48094
rect 158622 47858 195266 48094
rect 195502 47858 195586 48094
rect 195822 47858 232466 48094
rect 232702 47858 232786 48094
rect 233022 47858 269666 48094
rect 269902 47858 269986 48094
rect 270222 47858 306866 48094
rect 307102 47858 307186 48094
rect 307422 47858 344066 48094
rect 344302 47858 344386 48094
rect 344622 47858 381266 48094
rect 381502 47858 381586 48094
rect 381822 47858 418466 48094
rect 418702 47858 418786 48094
rect 419022 47858 455666 48094
rect 455902 47858 455986 48094
rect 456222 47858 492866 48094
rect 493102 47858 493186 48094
rect 493422 47858 530066 48094
rect 530302 47858 530386 48094
rect 530622 47858 567266 48094
rect 567502 47858 567586 48094
rect 567822 47858 582820 48094
rect 1104 47774 582820 47858
rect 1104 47538 9266 47774
rect 9502 47538 9586 47774
rect 9822 47538 46466 47774
rect 46702 47538 46786 47774
rect 47022 47538 83666 47774
rect 83902 47538 83986 47774
rect 84222 47538 120866 47774
rect 121102 47538 121186 47774
rect 121422 47538 158066 47774
rect 158302 47538 158386 47774
rect 158622 47538 195266 47774
rect 195502 47538 195586 47774
rect 195822 47538 232466 47774
rect 232702 47538 232786 47774
rect 233022 47538 269666 47774
rect 269902 47538 269986 47774
rect 270222 47538 306866 47774
rect 307102 47538 307186 47774
rect 307422 47538 344066 47774
rect 344302 47538 344386 47774
rect 344622 47538 381266 47774
rect 381502 47538 381586 47774
rect 381822 47538 418466 47774
rect 418702 47538 418786 47774
rect 419022 47538 455666 47774
rect 455902 47538 455986 47774
rect 456222 47538 492866 47774
rect 493102 47538 493186 47774
rect 493422 47538 530066 47774
rect 530302 47538 530386 47774
rect 530622 47538 567266 47774
rect 567502 47538 567586 47774
rect 567822 47538 582820 47774
rect 1104 47506 582820 47538
rect 1104 44374 582820 44406
rect 1104 44138 5546 44374
rect 5782 44138 5866 44374
rect 6102 44138 42746 44374
rect 42982 44138 43066 44374
rect 43302 44138 79946 44374
rect 80182 44138 80266 44374
rect 80502 44138 117146 44374
rect 117382 44138 117466 44374
rect 117702 44138 154346 44374
rect 154582 44138 154666 44374
rect 154902 44138 191546 44374
rect 191782 44138 191866 44374
rect 192102 44138 228746 44374
rect 228982 44138 229066 44374
rect 229302 44138 265946 44374
rect 266182 44138 266266 44374
rect 266502 44138 303146 44374
rect 303382 44138 303466 44374
rect 303702 44138 340346 44374
rect 340582 44138 340666 44374
rect 340902 44138 377546 44374
rect 377782 44138 377866 44374
rect 378102 44138 414746 44374
rect 414982 44138 415066 44374
rect 415302 44138 451946 44374
rect 452182 44138 452266 44374
rect 452502 44138 489146 44374
rect 489382 44138 489466 44374
rect 489702 44138 526346 44374
rect 526582 44138 526666 44374
rect 526902 44138 563546 44374
rect 563782 44138 563866 44374
rect 564102 44138 582820 44374
rect 1104 44054 582820 44138
rect 1104 43818 5546 44054
rect 5782 43818 5866 44054
rect 6102 43818 42746 44054
rect 42982 43818 43066 44054
rect 43302 43818 79946 44054
rect 80182 43818 80266 44054
rect 80502 43818 117146 44054
rect 117382 43818 117466 44054
rect 117702 43818 154346 44054
rect 154582 43818 154666 44054
rect 154902 43818 191546 44054
rect 191782 43818 191866 44054
rect 192102 43818 228746 44054
rect 228982 43818 229066 44054
rect 229302 43818 265946 44054
rect 266182 43818 266266 44054
rect 266502 43818 303146 44054
rect 303382 43818 303466 44054
rect 303702 43818 340346 44054
rect 340582 43818 340666 44054
rect 340902 43818 377546 44054
rect 377782 43818 377866 44054
rect 378102 43818 414746 44054
rect 414982 43818 415066 44054
rect 415302 43818 451946 44054
rect 452182 43818 452266 44054
rect 452502 43818 489146 44054
rect 489382 43818 489466 44054
rect 489702 43818 526346 44054
rect 526582 43818 526666 44054
rect 526902 43818 563546 44054
rect 563782 43818 563866 44054
rect 564102 43818 582820 44054
rect 1104 43786 582820 43818
rect 1104 40654 582820 40686
rect 1104 40418 1826 40654
rect 2062 40418 2146 40654
rect 2382 40418 39026 40654
rect 39262 40418 39346 40654
rect 39582 40418 76226 40654
rect 76462 40418 76546 40654
rect 76782 40418 113426 40654
rect 113662 40418 113746 40654
rect 113982 40418 150626 40654
rect 150862 40418 150946 40654
rect 151182 40418 187826 40654
rect 188062 40418 188146 40654
rect 188382 40418 225026 40654
rect 225262 40418 225346 40654
rect 225582 40418 262226 40654
rect 262462 40418 262546 40654
rect 262782 40418 299426 40654
rect 299662 40418 299746 40654
rect 299982 40418 336626 40654
rect 336862 40418 336946 40654
rect 337182 40418 373826 40654
rect 374062 40418 374146 40654
rect 374382 40418 411026 40654
rect 411262 40418 411346 40654
rect 411582 40418 448226 40654
rect 448462 40418 448546 40654
rect 448782 40418 485426 40654
rect 485662 40418 485746 40654
rect 485982 40418 522626 40654
rect 522862 40418 522946 40654
rect 523182 40418 559826 40654
rect 560062 40418 560146 40654
rect 560382 40418 582820 40654
rect 1104 40334 582820 40418
rect 1104 40098 1826 40334
rect 2062 40098 2146 40334
rect 2382 40098 39026 40334
rect 39262 40098 39346 40334
rect 39582 40098 76226 40334
rect 76462 40098 76546 40334
rect 76782 40098 113426 40334
rect 113662 40098 113746 40334
rect 113982 40098 150626 40334
rect 150862 40098 150946 40334
rect 151182 40098 187826 40334
rect 188062 40098 188146 40334
rect 188382 40098 225026 40334
rect 225262 40098 225346 40334
rect 225582 40098 262226 40334
rect 262462 40098 262546 40334
rect 262782 40098 299426 40334
rect 299662 40098 299746 40334
rect 299982 40098 336626 40334
rect 336862 40098 336946 40334
rect 337182 40098 373826 40334
rect 374062 40098 374146 40334
rect 374382 40098 411026 40334
rect 411262 40098 411346 40334
rect 411582 40098 448226 40334
rect 448462 40098 448546 40334
rect 448782 40098 485426 40334
rect 485662 40098 485746 40334
rect 485982 40098 522626 40334
rect 522862 40098 522946 40334
rect 523182 40098 559826 40334
rect 560062 40098 560146 40334
rect 560382 40098 582820 40334
rect 1104 40066 582820 40098
rect 1104 29494 582820 29526
rect 1104 29258 27866 29494
rect 28102 29258 28186 29494
rect 28422 29258 65066 29494
rect 65302 29258 65386 29494
rect 65622 29258 102266 29494
rect 102502 29258 102586 29494
rect 102822 29258 139466 29494
rect 139702 29258 139786 29494
rect 140022 29258 176666 29494
rect 176902 29258 176986 29494
rect 177222 29258 213866 29494
rect 214102 29258 214186 29494
rect 214422 29258 251066 29494
rect 251302 29258 251386 29494
rect 251622 29258 288266 29494
rect 288502 29258 288586 29494
rect 288822 29258 325466 29494
rect 325702 29258 325786 29494
rect 326022 29258 362666 29494
rect 362902 29258 362986 29494
rect 363222 29258 399866 29494
rect 400102 29258 400186 29494
rect 400422 29258 437066 29494
rect 437302 29258 437386 29494
rect 437622 29258 474266 29494
rect 474502 29258 474586 29494
rect 474822 29258 511466 29494
rect 511702 29258 511786 29494
rect 512022 29258 548666 29494
rect 548902 29258 548986 29494
rect 549222 29258 582820 29494
rect 1104 29174 582820 29258
rect 1104 28938 27866 29174
rect 28102 28938 28186 29174
rect 28422 28938 65066 29174
rect 65302 28938 65386 29174
rect 65622 28938 102266 29174
rect 102502 28938 102586 29174
rect 102822 28938 139466 29174
rect 139702 28938 139786 29174
rect 140022 28938 176666 29174
rect 176902 28938 176986 29174
rect 177222 28938 213866 29174
rect 214102 28938 214186 29174
rect 214422 28938 251066 29174
rect 251302 28938 251386 29174
rect 251622 28938 288266 29174
rect 288502 28938 288586 29174
rect 288822 28938 325466 29174
rect 325702 28938 325786 29174
rect 326022 28938 362666 29174
rect 362902 28938 362986 29174
rect 363222 28938 399866 29174
rect 400102 28938 400186 29174
rect 400422 28938 437066 29174
rect 437302 28938 437386 29174
rect 437622 28938 474266 29174
rect 474502 28938 474586 29174
rect 474822 28938 511466 29174
rect 511702 28938 511786 29174
rect 512022 28938 548666 29174
rect 548902 28938 548986 29174
rect 549222 28938 582820 29174
rect 1104 28906 582820 28938
rect 1104 25774 582820 25806
rect 1104 25538 24146 25774
rect 24382 25538 24466 25774
rect 24702 25538 61346 25774
rect 61582 25538 61666 25774
rect 61902 25538 98546 25774
rect 98782 25538 98866 25774
rect 99102 25538 135746 25774
rect 135982 25538 136066 25774
rect 136302 25538 172946 25774
rect 173182 25538 173266 25774
rect 173502 25538 210146 25774
rect 210382 25538 210466 25774
rect 210702 25538 247346 25774
rect 247582 25538 247666 25774
rect 247902 25538 284546 25774
rect 284782 25538 284866 25774
rect 285102 25538 321746 25774
rect 321982 25538 322066 25774
rect 322302 25538 358946 25774
rect 359182 25538 359266 25774
rect 359502 25538 396146 25774
rect 396382 25538 396466 25774
rect 396702 25538 433346 25774
rect 433582 25538 433666 25774
rect 433902 25538 470546 25774
rect 470782 25538 470866 25774
rect 471102 25538 507746 25774
rect 507982 25538 508066 25774
rect 508302 25538 544946 25774
rect 545182 25538 545266 25774
rect 545502 25538 582146 25774
rect 582382 25538 582466 25774
rect 582702 25538 582820 25774
rect 1104 25454 582820 25538
rect 1104 25218 24146 25454
rect 24382 25218 24466 25454
rect 24702 25218 61346 25454
rect 61582 25218 61666 25454
rect 61902 25218 98546 25454
rect 98782 25218 98866 25454
rect 99102 25218 135746 25454
rect 135982 25218 136066 25454
rect 136302 25218 172946 25454
rect 173182 25218 173266 25454
rect 173502 25218 210146 25454
rect 210382 25218 210466 25454
rect 210702 25218 247346 25454
rect 247582 25218 247666 25454
rect 247902 25218 284546 25454
rect 284782 25218 284866 25454
rect 285102 25218 321746 25454
rect 321982 25218 322066 25454
rect 322302 25218 358946 25454
rect 359182 25218 359266 25454
rect 359502 25218 396146 25454
rect 396382 25218 396466 25454
rect 396702 25218 433346 25454
rect 433582 25218 433666 25454
rect 433902 25218 470546 25454
rect 470782 25218 470866 25454
rect 471102 25218 507746 25454
rect 507982 25218 508066 25454
rect 508302 25218 544946 25454
rect 545182 25218 545266 25454
rect 545502 25218 582146 25454
rect 582382 25218 582466 25454
rect 582702 25218 582820 25454
rect 1104 25186 582820 25218
rect 1104 22054 582820 22086
rect 1104 21818 20426 22054
rect 20662 21818 20746 22054
rect 20982 21818 57626 22054
rect 57862 21818 57946 22054
rect 58182 21818 94826 22054
rect 95062 21818 95146 22054
rect 95382 21818 132026 22054
rect 132262 21818 132346 22054
rect 132582 21818 169226 22054
rect 169462 21818 169546 22054
rect 169782 21818 206426 22054
rect 206662 21818 206746 22054
rect 206982 21818 243626 22054
rect 243862 21818 243946 22054
rect 244182 21818 280826 22054
rect 281062 21818 281146 22054
rect 281382 21818 318026 22054
rect 318262 21818 318346 22054
rect 318582 21818 355226 22054
rect 355462 21818 355546 22054
rect 355782 21818 392426 22054
rect 392662 21818 392746 22054
rect 392982 21818 429626 22054
rect 429862 21818 429946 22054
rect 430182 21818 466826 22054
rect 467062 21818 467146 22054
rect 467382 21818 504026 22054
rect 504262 21818 504346 22054
rect 504582 21818 541226 22054
rect 541462 21818 541546 22054
rect 541782 21818 578426 22054
rect 578662 21818 578746 22054
rect 578982 21818 582820 22054
rect 1104 21734 582820 21818
rect 1104 21498 20426 21734
rect 20662 21498 20746 21734
rect 20982 21498 57626 21734
rect 57862 21498 57946 21734
rect 58182 21498 94826 21734
rect 95062 21498 95146 21734
rect 95382 21498 132026 21734
rect 132262 21498 132346 21734
rect 132582 21498 169226 21734
rect 169462 21498 169546 21734
rect 169782 21498 206426 21734
rect 206662 21498 206746 21734
rect 206982 21498 243626 21734
rect 243862 21498 243946 21734
rect 244182 21498 280826 21734
rect 281062 21498 281146 21734
rect 281382 21498 318026 21734
rect 318262 21498 318346 21734
rect 318582 21498 355226 21734
rect 355462 21498 355546 21734
rect 355782 21498 392426 21734
rect 392662 21498 392746 21734
rect 392982 21498 429626 21734
rect 429862 21498 429946 21734
rect 430182 21498 466826 21734
rect 467062 21498 467146 21734
rect 467382 21498 504026 21734
rect 504262 21498 504346 21734
rect 504582 21498 541226 21734
rect 541462 21498 541546 21734
rect 541782 21498 578426 21734
rect 578662 21498 578746 21734
rect 578982 21498 582820 21734
rect 1104 21466 582820 21498
rect 1104 18334 582820 18366
rect 1104 18098 16706 18334
rect 16942 18098 17026 18334
rect 17262 18098 53906 18334
rect 54142 18098 54226 18334
rect 54462 18098 91106 18334
rect 91342 18098 91426 18334
rect 91662 18098 128306 18334
rect 128542 18098 128626 18334
rect 128862 18098 165506 18334
rect 165742 18098 165826 18334
rect 166062 18098 202706 18334
rect 202942 18098 203026 18334
rect 203262 18098 239906 18334
rect 240142 18098 240226 18334
rect 240462 18098 277106 18334
rect 277342 18098 277426 18334
rect 277662 18098 314306 18334
rect 314542 18098 314626 18334
rect 314862 18098 351506 18334
rect 351742 18098 351826 18334
rect 352062 18098 388706 18334
rect 388942 18098 389026 18334
rect 389262 18098 425906 18334
rect 426142 18098 426226 18334
rect 426462 18098 463106 18334
rect 463342 18098 463426 18334
rect 463662 18098 500306 18334
rect 500542 18098 500626 18334
rect 500862 18098 537506 18334
rect 537742 18098 537826 18334
rect 538062 18098 574706 18334
rect 574942 18098 575026 18334
rect 575262 18098 582820 18334
rect 1104 18014 582820 18098
rect 1104 17778 16706 18014
rect 16942 17778 17026 18014
rect 17262 17778 53906 18014
rect 54142 17778 54226 18014
rect 54462 17778 91106 18014
rect 91342 17778 91426 18014
rect 91662 17778 128306 18014
rect 128542 17778 128626 18014
rect 128862 17778 165506 18014
rect 165742 17778 165826 18014
rect 166062 17778 202706 18014
rect 202942 17778 203026 18014
rect 203262 17778 239906 18014
rect 240142 17778 240226 18014
rect 240462 17778 277106 18014
rect 277342 17778 277426 18014
rect 277662 17778 314306 18014
rect 314542 17778 314626 18014
rect 314862 17778 351506 18014
rect 351742 17778 351826 18014
rect 352062 17778 388706 18014
rect 388942 17778 389026 18014
rect 389262 17778 425906 18014
rect 426142 17778 426226 18014
rect 426462 17778 463106 18014
rect 463342 17778 463426 18014
rect 463662 17778 500306 18014
rect 500542 17778 500626 18014
rect 500862 17778 537506 18014
rect 537742 17778 537826 18014
rect 538062 17778 574706 18014
rect 574942 17778 575026 18014
rect 575262 17778 582820 18014
rect 1104 17746 582820 17778
rect 1104 14614 582820 14646
rect 1104 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 50186 14614
rect 50422 14378 50506 14614
rect 50742 14378 87386 14614
rect 87622 14378 87706 14614
rect 87942 14378 124586 14614
rect 124822 14378 124906 14614
rect 125142 14378 161786 14614
rect 162022 14378 162106 14614
rect 162342 14378 198986 14614
rect 199222 14378 199306 14614
rect 199542 14378 236186 14614
rect 236422 14378 236506 14614
rect 236742 14378 273386 14614
rect 273622 14378 273706 14614
rect 273942 14378 310586 14614
rect 310822 14378 310906 14614
rect 311142 14378 347786 14614
rect 348022 14378 348106 14614
rect 348342 14378 384986 14614
rect 385222 14378 385306 14614
rect 385542 14378 422186 14614
rect 422422 14378 422506 14614
rect 422742 14378 459386 14614
rect 459622 14378 459706 14614
rect 459942 14378 496586 14614
rect 496822 14378 496906 14614
rect 497142 14378 533786 14614
rect 534022 14378 534106 14614
rect 534342 14378 570986 14614
rect 571222 14378 571306 14614
rect 571542 14378 582820 14614
rect 1104 14294 582820 14378
rect 1104 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 50186 14294
rect 50422 14058 50506 14294
rect 50742 14058 87386 14294
rect 87622 14058 87706 14294
rect 87942 14058 124586 14294
rect 124822 14058 124906 14294
rect 125142 14058 161786 14294
rect 162022 14058 162106 14294
rect 162342 14058 198986 14294
rect 199222 14058 199306 14294
rect 199542 14058 236186 14294
rect 236422 14058 236506 14294
rect 236742 14058 273386 14294
rect 273622 14058 273706 14294
rect 273942 14058 310586 14294
rect 310822 14058 310906 14294
rect 311142 14058 347786 14294
rect 348022 14058 348106 14294
rect 348342 14058 384986 14294
rect 385222 14058 385306 14294
rect 385542 14058 422186 14294
rect 422422 14058 422506 14294
rect 422742 14058 459386 14294
rect 459622 14058 459706 14294
rect 459942 14058 496586 14294
rect 496822 14058 496906 14294
rect 497142 14058 533786 14294
rect 534022 14058 534106 14294
rect 534342 14058 570986 14294
rect 571222 14058 571306 14294
rect 571542 14058 582820 14294
rect 1104 14026 582820 14058
rect 1104 10894 582820 10926
rect 1104 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 46466 10894
rect 46702 10658 46786 10894
rect 47022 10658 83666 10894
rect 83902 10658 83986 10894
rect 84222 10658 120866 10894
rect 121102 10658 121186 10894
rect 121422 10658 158066 10894
rect 158302 10658 158386 10894
rect 158622 10658 195266 10894
rect 195502 10658 195586 10894
rect 195822 10658 232466 10894
rect 232702 10658 232786 10894
rect 233022 10658 269666 10894
rect 269902 10658 269986 10894
rect 270222 10658 306866 10894
rect 307102 10658 307186 10894
rect 307422 10658 344066 10894
rect 344302 10658 344386 10894
rect 344622 10658 381266 10894
rect 381502 10658 381586 10894
rect 381822 10658 418466 10894
rect 418702 10658 418786 10894
rect 419022 10658 455666 10894
rect 455902 10658 455986 10894
rect 456222 10658 492866 10894
rect 493102 10658 493186 10894
rect 493422 10658 530066 10894
rect 530302 10658 530386 10894
rect 530622 10658 567266 10894
rect 567502 10658 567586 10894
rect 567822 10658 582820 10894
rect 1104 10574 582820 10658
rect 1104 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 46466 10574
rect 46702 10338 46786 10574
rect 47022 10338 83666 10574
rect 83902 10338 83986 10574
rect 84222 10338 120866 10574
rect 121102 10338 121186 10574
rect 121422 10338 158066 10574
rect 158302 10338 158386 10574
rect 158622 10338 195266 10574
rect 195502 10338 195586 10574
rect 195822 10338 232466 10574
rect 232702 10338 232786 10574
rect 233022 10338 269666 10574
rect 269902 10338 269986 10574
rect 270222 10338 306866 10574
rect 307102 10338 307186 10574
rect 307422 10338 344066 10574
rect 344302 10338 344386 10574
rect 344622 10338 381266 10574
rect 381502 10338 381586 10574
rect 381822 10338 418466 10574
rect 418702 10338 418786 10574
rect 419022 10338 455666 10574
rect 455902 10338 455986 10574
rect 456222 10338 492866 10574
rect 493102 10338 493186 10574
rect 493422 10338 530066 10574
rect 530302 10338 530386 10574
rect 530622 10338 567266 10574
rect 567502 10338 567586 10574
rect 567822 10338 582820 10574
rect 1104 10306 582820 10338
rect 1104 7174 582820 7206
rect 1104 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 42746 7174
rect 42982 6938 43066 7174
rect 43302 6938 79946 7174
rect 80182 6938 80266 7174
rect 80502 6938 117146 7174
rect 117382 6938 117466 7174
rect 117702 6938 154346 7174
rect 154582 6938 154666 7174
rect 154902 6938 191546 7174
rect 191782 6938 191866 7174
rect 192102 6938 228746 7174
rect 228982 6938 229066 7174
rect 229302 6938 265946 7174
rect 266182 6938 266266 7174
rect 266502 6938 303146 7174
rect 303382 6938 303466 7174
rect 303702 6938 340346 7174
rect 340582 6938 340666 7174
rect 340902 6938 377546 7174
rect 377782 6938 377866 7174
rect 378102 6938 414746 7174
rect 414982 6938 415066 7174
rect 415302 6938 451946 7174
rect 452182 6938 452266 7174
rect 452502 6938 489146 7174
rect 489382 6938 489466 7174
rect 489702 6938 526346 7174
rect 526582 6938 526666 7174
rect 526902 6938 563546 7174
rect 563782 6938 563866 7174
rect 564102 6938 582820 7174
rect 1104 6854 582820 6938
rect 1104 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 42746 6854
rect 42982 6618 43066 6854
rect 43302 6618 79946 6854
rect 80182 6618 80266 6854
rect 80502 6618 117146 6854
rect 117382 6618 117466 6854
rect 117702 6618 154346 6854
rect 154582 6618 154666 6854
rect 154902 6618 191546 6854
rect 191782 6618 191866 6854
rect 192102 6618 228746 6854
rect 228982 6618 229066 6854
rect 229302 6618 265946 6854
rect 266182 6618 266266 6854
rect 266502 6618 303146 6854
rect 303382 6618 303466 6854
rect 303702 6618 340346 6854
rect 340582 6618 340666 6854
rect 340902 6618 377546 6854
rect 377782 6618 377866 6854
rect 378102 6618 414746 6854
rect 414982 6618 415066 6854
rect 415302 6618 451946 6854
rect 452182 6618 452266 6854
rect 452502 6618 489146 6854
rect 489382 6618 489466 6854
rect 489702 6618 526346 6854
rect 526582 6618 526666 6854
rect 526902 6618 563546 6854
rect 563782 6618 563866 6854
rect 564102 6618 582820 6854
rect 1104 6586 582820 6618
rect 1104 3454 582820 3486
rect 1104 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 39026 3454
rect 39262 3218 39346 3454
rect 39582 3218 76226 3454
rect 76462 3218 76546 3454
rect 76782 3218 113426 3454
rect 113662 3218 113746 3454
rect 113982 3218 150626 3454
rect 150862 3218 150946 3454
rect 151182 3218 187826 3454
rect 188062 3218 188146 3454
rect 188382 3218 225026 3454
rect 225262 3218 225346 3454
rect 225582 3218 262226 3454
rect 262462 3218 262546 3454
rect 262782 3218 299426 3454
rect 299662 3218 299746 3454
rect 299982 3218 336626 3454
rect 336862 3218 336946 3454
rect 337182 3218 373826 3454
rect 374062 3218 374146 3454
rect 374382 3218 411026 3454
rect 411262 3218 411346 3454
rect 411582 3218 448226 3454
rect 448462 3218 448546 3454
rect 448782 3218 485426 3454
rect 485662 3218 485746 3454
rect 485982 3218 522626 3454
rect 522862 3218 522946 3454
rect 523182 3218 559826 3454
rect 560062 3218 560146 3454
rect 560382 3218 582820 3454
rect 1104 3134 582820 3218
rect 1104 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 39026 3134
rect 39262 2898 39346 3134
rect 39582 2898 76226 3134
rect 76462 2898 76546 3134
rect 76782 2898 113426 3134
rect 113662 2898 113746 3134
rect 113982 2898 150626 3134
rect 150862 2898 150946 3134
rect 151182 2898 187826 3134
rect 188062 2898 188146 3134
rect 188382 2898 225026 3134
rect 225262 2898 225346 3134
rect 225582 2898 262226 3134
rect 262462 2898 262546 3134
rect 262782 2898 299426 3134
rect 299662 2898 299746 3134
rect 299982 2898 336626 3134
rect 336862 2898 336946 3134
rect 337182 2898 373826 3134
rect 374062 2898 374146 3134
rect 374382 2898 411026 3134
rect 411262 2898 411346 3134
rect 411582 2898 448226 3134
rect 448462 2898 448546 3134
rect 448782 2898 485426 3134
rect 485662 2898 485746 3134
rect 485982 2898 522626 3134
rect 522862 2898 522946 3134
rect 523182 2898 559826 3134
rect 560062 2898 560146 3134
rect 560382 2898 582820 3134
rect 1104 2866 582820 2898
use mux16x1_project  mprj
timestamp 0
transform 1 0 480000 0 1 320000
box 0 552 10000 22000
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s 1794 2176 2414 701760 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 38994 2176 39614 701760 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 76194 2176 76814 701760 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 113394 2176 114014 701760 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 150594 2176 151214 701760 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 187794 2176 188414 701760 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 224994 2176 225614 701760 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 262194 2176 262814 701760 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 299394 2176 300014 701760 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 336594 2176 337214 701760 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 373794 2176 374414 701760 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 410994 2176 411614 701760 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 448194 2176 448814 701760 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 485394 2176 486014 319988 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 485394 341772 486014 701760 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 522594 2176 523214 701760 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 559794 2176 560414 701760 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s 1104 2866 582820 3486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s 1104 40066 582820 40686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s 1104 77266 582820 77886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s 1104 114466 582820 115086 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s 1104 151666 582820 152286 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s 1104 188866 582820 189486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s 1104 226066 582820 226686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s 1104 263266 582820 263886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s 1104 300466 582820 301086 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s 1104 337666 582820 338286 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s 1104 374866 582820 375486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s 1104 412066 582820 412686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s 1104 449266 582820 449886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s 1104 486466 582820 487086 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s 1104 523666 582820 524286 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s 1104 560866 582820 561486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s 1104 598066 582820 598686 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s 1104 635266 582820 635886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s 1104 672466 582820 673086 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 9234 2176 9854 701760 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 46434 2176 47054 701760 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 83634 2176 84254 701760 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 120834 2176 121454 701760 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 158034 2176 158654 701760 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 195234 2176 195854 701760 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 232434 2176 233054 701760 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 269634 2176 270254 701760 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 306834 2176 307454 701760 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 344034 2176 344654 701760 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 381234 2176 381854 701760 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 418434 2176 419054 701760 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 455634 2176 456254 701760 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 492834 2176 493454 701760 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 530034 2176 530654 701760 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 567234 2176 567854 701760 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s 1104 10306 582820 10926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s 1104 47506 582820 48126 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s 1104 84706 582820 85326 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s 1104 121906 582820 122526 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s 1104 159106 582820 159726 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s 1104 196306 582820 196926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s 1104 233506 582820 234126 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s 1104 270706 582820 271326 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s 1104 307906 582820 308526 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s 1104 345106 582820 345726 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s 1104 382306 582820 382926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s 1104 419506 582820 420126 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s 1104 456706 582820 457326 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s 1104 493906 582820 494526 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s 1104 531106 582820 531726 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s 1104 568306 582820 568926 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s 1104 605506 582820 606126 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s 1104 642706 582820 643326 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s 1104 679906 582820 680526 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 16674 2176 17294 701760 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 53874 2176 54494 701760 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 91074 2176 91694 701760 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 128274 2176 128894 701760 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 165474 2176 166094 701760 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 202674 2176 203294 701760 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 239874 2176 240494 701760 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 277074 2176 277694 701760 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 314274 2176 314894 701760 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 351474 2176 352094 701760 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 388674 2176 389294 701760 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 425874 2176 426494 701760 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 463074 2176 463694 701760 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 500274 2176 500894 701760 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 537474 2176 538094 701760 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 574674 2176 575294 701760 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s 1104 17746 582820 18366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s 1104 54946 582820 55566 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s 1104 92146 582820 92766 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s 1104 129346 582820 129966 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s 1104 166546 582820 167166 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s 1104 203746 582820 204366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s 1104 240946 582820 241566 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s 1104 278146 582820 278766 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s 1104 315346 582820 315966 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s 1104 352546 582820 353166 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s 1104 389746 582820 390366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s 1104 426946 582820 427566 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s 1104 464146 582820 464766 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s 1104 501346 582820 501966 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s 1104 538546 582820 539166 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s 1104 575746 582820 576366 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s 1104 612946 582820 613566 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s 1104 650146 582820 650766 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s 1104 687346 582820 687966 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 24114 2176 24734 701760 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 61314 2176 61934 701760 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 98514 2176 99134 701760 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 135714 2176 136334 701760 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 172914 2176 173534 701760 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 210114 2176 210734 701760 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 247314 2176 247934 701760 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 284514 2176 285134 701760 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 321714 2176 322334 701760 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 358914 2176 359534 701760 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 396114 2176 396734 701760 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 433314 2176 433934 701760 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 470514 2176 471134 701760 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 507714 2176 508334 701760 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 544914 2176 545534 701760 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 582114 2176 582734 701760 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s 1104 25186 582820 25806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s 1104 62386 582820 63006 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s 1104 99586 582820 100206 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s 1104 136786 582820 137406 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s 1104 173986 582820 174606 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s 1104 211186 582820 211806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s 1104 248386 582820 249006 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s 1104 285586 582820 286206 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s 1104 322786 582820 323406 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s 1104 359986 582820 360606 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s 1104 397186 582820 397806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s 1104 434386 582820 435006 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s 1104 471586 582820 472206 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s 1104 508786 582820 509406 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s 1104 545986 582820 546606 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s 1104 583186 582820 583806 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s 1104 620386 582820 621006 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s 1104 657586 582820 658206 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s 1104 694786 582820 695406 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 20394 2176 21014 701760 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 57594 2176 58214 701760 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 94794 2176 95414 701760 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 131994 2176 132614 701760 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 169194 2176 169814 701760 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 206394 2176 207014 701760 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 243594 2176 244214 701760 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 280794 2176 281414 701760 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 317994 2176 318614 701760 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 355194 2176 355814 701760 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 392394 2176 393014 701760 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 429594 2176 430214 701760 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 466794 2176 467414 701760 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 503994 2176 504614 701760 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 541194 2176 541814 701760 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 578394 2176 579014 701760 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s 1104 21466 582820 22086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s 1104 58666 582820 59286 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s 1104 95866 582820 96486 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s 1104 133066 582820 133686 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s 1104 170266 582820 170886 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s 1104 207466 582820 208086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s 1104 244666 582820 245286 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s 1104 281866 582820 282486 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s 1104 319066 582820 319686 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s 1104 356266 582820 356886 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s 1104 393466 582820 394086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s 1104 430666 582820 431286 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s 1104 467866 582820 468486 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s 1104 505066 582820 505686 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s 1104 542266 582820 542886 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s 1104 579466 582820 580086 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s 1104 616666 582820 617286 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s 1104 653866 582820 654486 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s 1104 691066 582820 691686 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 27834 2176 28454 701760 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 65034 2176 65654 701760 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 102234 2176 102854 701760 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 139434 2176 140054 701760 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 176634 2176 177254 701760 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 213834 2176 214454 701760 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 251034 2176 251654 701760 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 288234 2176 288854 701760 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 325434 2176 326054 701760 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 362634 2176 363254 701760 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 399834 2176 400454 701760 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 437034 2176 437654 701760 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 474234 2176 474854 701760 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 511434 2176 512054 701760 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 548634 2176 549254 701760 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s 1104 28906 582820 29526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s 1104 66106 582820 66726 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s 1104 103306 582820 103926 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s 1104 140506 582820 141126 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s 1104 177706 582820 178326 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s 1104 214906 582820 215526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s 1104 252106 582820 252726 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s 1104 289306 582820 289926 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s 1104 326506 582820 327126 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s 1104 363706 582820 364326 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s 1104 400906 582820 401526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s 1104 438106 582820 438726 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s 1104 475306 582820 475926 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s 1104 512506 582820 513126 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s 1104 549706 582820 550326 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s 1104 586906 582820 587526 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s 1104 624106 582820 624726 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s 1104 661306 582820 661926 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s 1104 698506 582820 699126 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 5514 2176 6134 701760 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 42714 2176 43334 701760 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 79914 2176 80534 701760 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 117114 2176 117734 701760 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 154314 2176 154934 701760 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 191514 2176 192134 701760 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 228714 2176 229334 701760 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 265914 2176 266534 701760 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 303114 2176 303734 701760 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 340314 2176 340934 701760 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 377514 2176 378134 701760 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 414714 2176 415334 701760 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 451914 2176 452534 701760 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 489114 2176 489734 319988 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 489114 341386 489734 701760 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 526314 2176 526934 701760 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 563514 2176 564134 701760 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s 1104 6586 582820 7206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s 1104 43786 582820 44406 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s 1104 80986 582820 81606 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s 1104 118186 582820 118806 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s 1104 155386 582820 156006 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s 1104 192586 582820 193206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s 1104 229786 582820 230406 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s 1104 266986 582820 267606 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s 1104 304186 582820 304806 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s 1104 341386 582820 342006 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s 1104 378586 582820 379206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s 1104 415786 582820 416406 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s 1104 452986 582820 453606 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s 1104 490186 582820 490806 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s 1104 527386 582820 528006 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s 1104 564586 582820 565206 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s 1104 601786 582820 602406 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s 1104 638986 582820 639606 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s 1104 676186 582820 676806 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 12954 2176 13574 701760 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 50154 2176 50774 701760 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 87354 2176 87974 701760 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 124554 2176 125174 701760 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 161754 2176 162374 701760 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 198954 2176 199574 701760 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 236154 2176 236774 701760 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 273354 2176 273974 701760 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 310554 2176 311174 701760 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 347754 2176 348374 701760 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 384954 2176 385574 701760 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 422154 2176 422774 701760 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 459354 2176 459974 701760 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 496554 2176 497174 701760 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 533754 2176 534374 701760 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 570954 2176 571574 701760 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s 1104 14026 582820 14646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s 1104 51226 582820 51846 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s 1104 88426 582820 89046 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s 1104 125626 582820 126246 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s 1104 162826 582820 163446 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s 1104 200026 582820 200646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s 1104 237226 582820 237846 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s 1104 274426 582820 275046 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s 1104 311626 582820 312246 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s 1104 348826 582820 349446 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s 1104 386026 582820 386646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s 1104 423226 582820 423846 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s 1104 460426 582820 461046 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s 1104 497626 582820 498246 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s 1104 534826 582820 535446 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s 1104 572026 582820 572646 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s 1104 609226 582820 609846 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s 1104 646426 582820 647046 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s 1104 683626 582820 684246 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
