magic
tech sky130A
magscale 1 2
timestamp 1708619853
<< error_s >>
rect 3131 2103 3132 2114
rect 3321 2103 3322 2114
rect 3407 2103 3408 2114
rect 4906 2103 4907 2114
rect 5096 2103 5097 2114
rect 5182 2103 5183 2114
rect 5862 2103 5863 2114
rect 6052 2103 6053 2114
rect 6138 2103 6139 2114
rect 6411 2103 6412 2114
rect 6609 2103 6610 2114
rect 8062 2103 8063 2114
rect 8252 2103 8253 2114
rect 8338 2103 8339 2114
rect 9018 2103 9019 2114
rect 9208 2103 9209 2114
rect 9294 2103 9295 2114
rect 9567 2103 9568 2114
rect 9765 2103 9766 2114
rect 11217 2103 11218 2114
rect 11407 2103 11408 2114
rect 11493 2103 11494 2114
rect 12173 2103 12174 2114
rect 12363 2103 12364 2114
rect 12449 2103 12450 2114
rect 12722 2103 12723 2114
rect 12920 2103 12921 2114
rect 14374 2103 14375 2114
rect 14564 2103 14565 2114
rect 14650 2103 14651 2114
rect 15330 2103 15331 2114
rect 15520 2103 15521 2114
rect 15606 2103 15607 2114
rect 15879 2103 15880 2114
rect 16077 2103 16078 2114
rect 17531 2103 17532 2114
rect 17721 2103 17722 2114
rect 17807 2103 17808 2114
rect 18487 2103 18488 2114
rect 18677 2103 18678 2114
rect 18763 2103 18764 2114
rect 19036 2103 19037 2114
rect 19234 2103 19235 2114
rect 3142 2063 3143 2103
rect 3332 2063 3333 2103
rect 3418 2063 3419 2103
rect 4917 2063 4918 2103
rect 5107 2063 5108 2103
rect 5193 2063 5194 2103
rect 5873 2063 5874 2103
rect 6063 2063 6064 2103
rect 6149 2063 6150 2103
rect 6422 2063 6423 2103
rect 6620 2063 6621 2103
rect 8073 2063 8074 2103
rect 8263 2063 8264 2103
rect 8349 2063 8350 2103
rect 9029 2063 9030 2103
rect 9219 2063 9220 2103
rect 9305 2063 9306 2103
rect 9578 2063 9579 2103
rect 9776 2063 9777 2103
rect 11228 2063 11229 2103
rect 11418 2063 11419 2103
rect 11504 2063 11505 2103
rect 12184 2063 12185 2103
rect 12374 2063 12375 2103
rect 12460 2063 12461 2103
rect 12733 2063 12734 2103
rect 12931 2063 12932 2103
rect 14385 2063 14386 2103
rect 14575 2063 14576 2103
rect 14661 2063 14662 2103
rect 15341 2063 15342 2103
rect 15531 2063 15532 2103
rect 15617 2063 15618 2103
rect 15890 2063 15891 2103
rect 16088 2063 16089 2103
rect 17542 2063 17543 2103
rect 17732 2063 17733 2103
rect 17818 2063 17819 2103
rect 18498 2063 18499 2103
rect 18688 2063 18689 2103
rect 18774 2063 18775 2103
rect 19047 2063 19048 2103
rect 19245 2063 19246 2103
rect 6070 1936 6097 1943
rect 9226 1936 9253 1943
rect 12381 1936 12408 1943
rect 15538 1936 15565 1943
rect 18695 1936 18722 1943
rect 6070 1915 6138 1936
rect 9226 1915 9294 1936
rect 12381 1915 12449 1936
rect 15538 1915 15606 1936
rect 18695 1915 18763 1936
rect 6070 1909 6125 1915
rect 9226 1909 9281 1915
rect 12381 1909 12436 1915
rect 15538 1909 15593 1915
rect 18695 1909 18750 1915
rect 6109 1908 6110 1909
rect 9265 1908 9266 1909
rect 12420 1908 12421 1909
rect 15577 1908 15578 1909
rect 18734 1908 18735 1909
rect 6082 1902 6137 1908
rect 9238 1902 9293 1908
rect 12393 1902 12448 1908
rect 15550 1902 15605 1908
rect 18707 1902 18762 1908
rect 6109 1880 6110 1902
rect 9265 1880 9266 1902
rect 12420 1880 12421 1902
rect 15577 1880 15578 1902
rect 18734 1880 18735 1902
rect 4959 1754 4981 1783
rect 4987 1754 5009 1755
rect 8115 1754 8137 1783
rect 8143 1754 8165 1755
rect 11270 1754 11292 1783
rect 11298 1754 11320 1755
rect 14427 1754 14449 1783
rect 14455 1754 14477 1755
rect 17584 1754 17606 1783
rect 17612 1754 17634 1755
rect 13031 1749 13176 1750
rect 3131 1673 3132 1684
rect 3321 1673 3322 1684
rect 3407 1673 3408 1684
rect 4906 1673 4907 1684
rect 5096 1673 5097 1684
rect 5182 1673 5183 1684
rect 5862 1673 5863 1684
rect 6052 1673 6053 1684
rect 6138 1673 6139 1684
rect 6411 1673 6412 1684
rect 6609 1673 6610 1684
rect 8062 1673 8063 1684
rect 8252 1673 8253 1684
rect 8338 1673 8339 1684
rect 9018 1673 9019 1684
rect 9208 1673 9209 1684
rect 9294 1673 9295 1684
rect 9567 1673 9568 1684
rect 9765 1673 9766 1684
rect 11217 1673 11218 1684
rect 11407 1673 11408 1684
rect 11493 1673 11494 1684
rect 12173 1673 12174 1684
rect 12363 1673 12364 1684
rect 12449 1673 12450 1684
rect 12722 1673 12723 1684
rect 12920 1673 12921 1684
rect 14374 1673 14375 1684
rect 14564 1673 14565 1684
rect 14650 1673 14651 1684
rect 15330 1673 15331 1684
rect 15520 1673 15521 1684
rect 15606 1673 15607 1684
rect 15879 1673 15880 1684
rect 16077 1673 16078 1684
rect 17531 1673 17532 1684
rect 17721 1673 17722 1684
rect 17807 1673 17808 1684
rect 18487 1673 18488 1684
rect 18677 1673 18678 1684
rect 18763 1673 18764 1684
rect 19036 1673 19037 1684
rect 19234 1673 19235 1684
rect 3142 1477 3143 1673
rect 3332 1477 3333 1673
rect 3418 1477 3419 1673
rect 4852 1641 4879 1647
rect 4880 1646 4907 1647
rect 4917 1477 4918 1673
rect 5107 1477 5108 1673
rect 5193 1477 5194 1673
rect 5873 1477 5874 1673
rect 6063 1477 6064 1673
rect 6149 1477 6150 1673
rect 6422 1477 6423 1673
rect 6620 1477 6621 1673
rect 8008 1641 8035 1647
rect 8036 1646 8063 1647
rect 8073 1477 8074 1673
rect 8263 1477 8264 1673
rect 8349 1477 8350 1673
rect 9029 1477 9030 1673
rect 9219 1477 9220 1673
rect 9305 1477 9306 1673
rect 9578 1477 9579 1673
rect 9776 1477 9777 1673
rect 11163 1641 11190 1647
rect 11191 1646 11218 1647
rect 11228 1477 11229 1673
rect 11418 1477 11419 1673
rect 11504 1477 11505 1673
rect 12184 1477 12185 1673
rect 12374 1477 12375 1673
rect 12460 1477 12461 1673
rect 12733 1477 12734 1673
rect 12931 1477 12932 1673
rect 14320 1641 14347 1647
rect 14348 1646 14375 1647
rect 14385 1477 14386 1673
rect 14575 1477 14576 1673
rect 14661 1477 14662 1673
rect 15341 1477 15342 1673
rect 15531 1477 15532 1673
rect 15617 1477 15618 1673
rect 15890 1477 15891 1673
rect 16088 1477 16089 1673
rect 17477 1641 17504 1647
rect 17505 1646 17532 1647
rect 17542 1477 17543 1673
rect 17732 1477 17733 1673
rect 17818 1477 17819 1673
rect 18498 1477 18499 1673
rect 18688 1477 18689 1673
rect 18774 1477 18775 1673
rect 19047 1477 19048 1673
rect 19245 1477 19246 1673
rect 3456 1373 3480 1407
rect 5231 1373 5255 1407
rect 6187 1373 6211 1407
rect 8387 1373 8411 1407
rect 9343 1373 9367 1407
rect 11542 1373 11566 1407
rect 12498 1373 12522 1407
rect 14699 1373 14723 1407
rect 15655 1373 15679 1407
rect 17856 1373 17880 1407
rect 18812 1373 18836 1407
rect 6187 1085 6211 1119
rect 9343 1085 9367 1119
rect 12498 1085 12522 1119
rect 15655 1085 15679 1119
rect 18812 1085 18836 1119
rect 4939 1037 5082 1039
rect 8095 1037 8238 1039
rect 11250 1037 11393 1039
rect 14407 1037 14550 1039
rect 17564 1037 17707 1039
rect 3880 1023 3981 1034
rect 4167 1033 4431 1034
rect 4431 1023 4486 1033
rect 4589 1027 4598 1036
rect 4636 1027 4645 1036
rect 4939 1034 5061 1037
rect 4911 1033 4928 1034
rect 4741 1027 4911 1033
rect 3865 1021 3880 1023
rect 3859 1019 3865 1021
rect 4488 1019 4493 1021
rect 3855 1014 3859 1019
rect 4493 1014 4500 1019
rect 4580 1018 4589 1027
rect 4645 1024 4741 1027
rect 5082 1023 5190 1037
rect 4940 1015 4956 1022
rect 4958 1015 4974 1022
rect 4500 1007 4512 1014
rect 4930 1013 4942 1015
rect 4952 1013 4964 1015
rect 4970 1013 4974 1015
rect 5158 1013 5174 1022
rect 5190 1021 5208 1023
rect 5209 1017 5216 1020
rect 5216 1013 5222 1017
rect 5862 1015 5863 1026
rect 6052 1015 6053 1026
rect 6138 1015 6139 1026
rect 6411 1015 6412 1026
rect 6608 1015 6609 1026
rect 7036 1023 7137 1034
rect 7323 1033 7587 1034
rect 7587 1023 7642 1033
rect 7745 1027 7754 1036
rect 7792 1027 7801 1036
rect 8095 1034 8217 1037
rect 8067 1033 8084 1034
rect 7897 1027 8067 1033
rect 7021 1021 7036 1023
rect 7015 1019 7021 1021
rect 7644 1019 7649 1021
rect 4930 1008 4974 1013
rect 5117 1008 5154 1009
rect 5222 1008 5225 1013
rect 4926 1006 4928 1008
rect 4930 1006 5062 1008
rect 3981 1005 4335 1006
rect 3961 1003 3979 1005
rect 4421 1003 4434 1005
rect 4513 1003 4516 1005
rect 4924 1003 5062 1006
rect 3905 1000 3961 1003
rect 3779 992 3791 1000
rect 3801 992 3813 1000
rect 3877 994 3961 1000
rect 4434 994 4444 1003
rect 3877 993 3905 994
rect 3775 989 3777 992
rect 3877 991 3896 993
rect 4445 991 4448 993
rect 3817 988 3821 989
rect 3767 977 3775 988
rect 3778 986 3813 988
rect 3776 977 3778 983
rect 3767 976 3776 977
rect 3775 972 3776 976
rect 3774 971 3775 972
rect 3772 966 3774 969
rect 3647 964 3712 965
rect 3639 956 3647 964
rect 3712 956 3716 964
rect 3638 950 3639 956
rect 3767 954 3775 966
rect 3779 956 3781 986
rect 3810 985 3813 986
rect 3812 979 3813 985
rect 3817 981 3825 988
rect 3821 980 3829 981
rect 3853 980 3854 990
rect 3877 980 3892 991
rect 4151 981 4188 983
rect 3829 979 3835 980
rect 3852 979 3853 980
rect 3877 979 3884 980
rect 3835 969 3897 979
rect 3905 972 3911 978
rect 3951 972 3957 978
rect 4151 977 4177 981
rect 4188 977 4193 981
rect 4448 980 4461 991
rect 4424 979 4438 980
rect 4145 972 4151 977
rect 4193 972 4202 977
rect 4406 972 4424 979
rect 4438 977 4445 979
rect 4516 977 4537 1003
rect 4918 996 5062 1003
rect 5078 1006 5179 1008
rect 5078 996 5190 1006
rect 4879 990 4940 996
rect 4844 987 4879 990
rect 4657 981 4844 987
rect 4930 986 4940 990
rect 4445 972 4460 977
rect 3899 969 3905 972
rect 3906 970 3963 972
rect 4202 971 4203 972
rect 4040 970 4043 971
rect 4061 970 4064 971
rect 4143 970 4144 971
rect 4203 970 4206 971
rect 3906 969 3914 970
rect 3877 968 3914 969
rect 3779 954 3813 956
rect 3768 951 3770 954
rect 3764 938 3768 950
rect 3779 942 3791 950
rect 3804 945 3813 954
rect 3851 952 3852 955
rect 3877 951 3882 968
rect 3899 966 3914 968
rect 3957 966 3963 970
rect 4039 969 4040 970
rect 4064 969 4065 970
rect 4398 969 4406 972
rect 4435 971 4460 972
rect 4469 971 4473 972
rect 4431 970 4435 971
rect 4445 970 4482 971
rect 4430 969 4431 970
rect 4036 967 4039 969
rect 4065 967 4069 969
rect 4206 968 4207 969
rect 4207 967 4210 968
rect 3905 964 3914 966
rect 4032 965 4036 967
rect 4069 965 4073 967
rect 4390 966 4398 969
rect 4428 968 4430 969
rect 4424 967 4428 968
rect 4419 965 4424 967
rect 4445 965 4460 970
rect 4469 969 4473 970
rect 4482 969 4483 970
rect 4539 969 4544 975
rect 4580 971 4589 980
rect 4645 978 4657 981
rect 4645 971 4654 978
rect 4924 972 4940 986
rect 4963 972 4964 996
rect 4969 991 4990 996
rect 4974 990 4990 991
rect 5107 989 5113 996
rect 5159 989 5165 996
rect 5179 990 5190 996
rect 5225 990 5234 1008
rect 4974 972 4990 988
rect 5107 985 5115 989
rect 5113 983 5115 985
rect 5044 977 5051 978
rect 5053 977 5055 978
rect 5023 974 5044 977
rect 5055 974 5064 977
rect 5021 972 5023 974
rect 5064 972 5066 974
rect 4473 965 4478 969
rect 4483 965 4485 968
rect 4544 965 4547 969
rect 4030 964 4032 965
rect 4073 964 4075 965
rect 4385 964 4389 965
rect 4460 964 4463 965
rect 4485 964 4486 965
rect 3905 951 3910 964
rect 3958 955 3977 958
rect 4016 956 4030 964
rect 4075 959 4087 964
rect 4142 959 4143 964
rect 4087 956 4090 959
rect 4210 957 4213 964
rect 4381 962 4385 964
rect 4012 955 4016 956
rect 3814 949 3819 950
rect 3819 948 3824 949
rect 3824 947 3827 948
rect 3829 945 3838 947
rect 3802 942 3804 945
rect 3838 944 3843 945
rect 3843 943 3849 944
rect 3850 943 3851 951
rect 3877 943 3883 951
rect 3801 939 3802 942
rect 3849 938 3883 943
rect 3762 931 3764 937
rect 3799 930 3801 938
rect 3850 932 3851 938
rect 3877 935 3905 938
rect 3877 933 3907 935
rect 3877 931 3908 933
rect 3909 931 3910 951
rect 3977 946 4039 955
rect 4090 952 4095 956
rect 4141 951 4142 956
rect 4213 954 4214 956
rect 4350 950 4381 962
rect 4465 959 4469 962
rect 4480 960 4484 963
rect 4589 962 4598 971
rect 4622 961 4625 963
rect 4636 962 4645 971
rect 4930 970 4964 972
rect 4973 971 4974 972
rect 5020 971 5021 972
rect 4969 970 4974 971
rect 5019 970 5020 971
rect 4930 968 4974 970
rect 5017 969 5019 970
rect 5066 969 5069 972
rect 4926 965 4927 967
rect 4700 961 4709 963
rect 4617 959 4622 961
rect 3995 945 4005 946
rect 4027 945 4028 946
rect 3991 943 3995 945
rect 4039 943 4059 946
rect 4140 943 4141 950
rect 4213 943 4214 950
rect 4348 949 4350 950
rect 4262 943 4268 949
rect 4308 948 4314 949
rect 4345 948 4348 949
rect 4308 947 4345 948
rect 4308 943 4314 947
rect 4400 946 4406 952
rect 4446 946 4452 952
rect 4468 950 4469 959
rect 4615 958 4617 959
rect 4711 958 4717 961
rect 4486 955 4490 958
rect 4554 955 4556 958
rect 4717 956 4720 958
rect 4940 956 4956 968
rect 4958 956 4974 968
rect 5013 965 5017 968
rect 5069 965 5073 969
rect 5113 967 5116 983
rect 5012 964 5013 965
rect 5073 964 5074 965
rect 5011 963 5012 964
rect 5009 961 5011 963
rect 5074 961 5077 964
rect 5115 961 5116 967
rect 5119 967 5120 989
rect 5158 985 5165 989
rect 5186 987 5188 990
rect 5158 983 5159 985
rect 5179 984 5180 986
rect 5119 963 5121 967
rect 5152 963 5153 966
rect 5157 965 5159 983
rect 5188 981 5191 987
rect 5191 979 5192 981
rect 5193 975 5194 977
rect 5194 972 5195 975
rect 5234 973 5242 990
rect 5196 965 5199 969
rect 5119 961 5123 963
rect 5157 962 5158 965
rect 5199 963 5200 965
rect 5005 958 5008 961
rect 5077 959 5080 961
rect 5004 956 5005 958
rect 5080 957 5082 959
rect 4490 946 4500 955
rect 3979 931 3987 943
rect 3991 941 4025 943
rect 3715 924 3716 929
rect 3665 915 3674 924
rect 3712 920 3721 924
rect 3712 915 3726 920
rect 3656 912 3665 915
rect 3656 911 3659 912
rect 3649 908 3658 911
rect 3637 907 3658 908
rect 3637 905 3655 907
rect 3695 905 3701 911
rect 3715 906 3730 915
rect 3755 908 3762 929
rect 3637 900 3649 905
rect 3633 898 3636 900
rect 3637 899 3638 900
rect 3643 899 3649 900
rect 3701 899 3707 905
rect 3714 904 3726 906
rect 3753 904 3755 908
rect 3793 907 3799 929
rect 3850 926 3851 929
rect 3877 928 3938 931
rect 3877 917 3883 928
rect 3905 926 3938 928
rect 3899 925 3938 926
rect 3957 925 3963 926
rect 3899 921 3963 925
rect 3899 920 3985 921
rect 3877 913 3886 917
rect 3905 914 3911 920
rect 3951 914 3957 920
rect 3960 917 3985 920
rect 3969 913 3985 917
rect 3991 913 3993 941
rect 4022 939 4025 941
rect 3877 909 3892 913
rect 3979 909 3993 913
rect 4023 909 4025 939
rect 4029 931 4037 943
rect 4059 934 4122 943
rect 4256 938 4262 943
rect 4274 941 4310 943
rect 4274 938 4279 941
rect 4215 937 4262 938
rect 4276 937 4279 938
rect 4314 937 4320 943
rect 4394 940 4400 946
rect 4452 940 4458 946
rect 4215 936 4258 937
rect 4139 934 4140 936
rect 4161 934 4215 936
rect 4095 922 4110 934
rect 4122 933 4161 934
rect 4139 929 4140 933
rect 4271 929 4274 936
rect 4398 933 4400 934
rect 4396 929 4398 933
rect 3792 904 3793 906
rect 3852 905 3853 909
rect 3712 899 3714 904
rect 3858 903 3864 909
rect 3877 903 3896 909
rect 3904 903 3910 909
rect 3752 899 3753 903
rect 3711 897 3712 899
rect 3751 897 3752 899
rect 3625 884 3633 896
rect 3637 894 3655 896
rect 3710 895 3711 896
rect 3790 895 3792 903
rect 3852 897 3858 903
rect 3877 897 3916 903
rect 3918 897 3930 905
rect 3991 904 4008 909
rect 3999 899 4006 904
rect 4008 903 4012 904
rect 4028 903 4029 905
rect 4095 904 4110 920
rect 4137 906 4139 928
rect 4012 900 4031 903
rect 4136 900 4148 905
rect 4158 900 4170 905
rect 4211 904 4213 928
rect 4262 904 4271 928
rect 4307 904 4310 909
rect 4348 908 4383 910
rect 4394 908 4396 929
rect 4418 909 4419 929
rect 4466 928 4468 944
rect 4500 942 4505 946
rect 4556 942 4568 955
rect 4720 951 4730 956
rect 5003 953 5004 956
rect 4838 952 4875 953
rect 5002 952 5003 953
rect 5082 952 5084 956
rect 5110 955 5116 961
rect 5123 959 5129 961
rect 5130 957 5136 959
rect 5136 956 5139 957
rect 5156 956 5162 961
rect 5200 960 5201 963
rect 5201 958 5202 960
rect 4838 951 4863 952
rect 4875 951 4876 952
rect 5001 951 5002 952
rect 4732 948 4736 951
rect 4803 948 4830 951
rect 4878 948 4885 951
rect 4885 943 4896 948
rect 4931 945 4933 949
rect 4966 947 4967 949
rect 4999 948 5001 951
rect 4896 942 4900 943
rect 4568 939 4569 942
rect 4900 938 4907 942
rect 4510 929 4520 938
rect 4570 931 4576 938
rect 4907 937 4909 938
rect 4909 933 4925 937
rect 4925 932 4930 933
rect 4933 932 4941 944
rect 4930 929 4941 932
rect 4967 929 4971 944
rect 4997 943 4999 948
rect 5084 944 5087 951
rect 5104 949 5110 955
rect 5139 951 5180 956
rect 5202 955 5204 958
rect 5162 949 5168 951
rect 5204 948 5207 955
rect 4996 942 4997 943
rect 5207 942 5210 948
rect 5242 943 5243 973
rect 5350 951 5366 954
rect 5278 943 5301 951
rect 5356 943 5373 951
rect 4995 940 4996 942
rect 4994 939 4995 940
rect 5210 939 5211 942
rect 4993 937 4994 938
rect 4990 933 4993 937
rect 4988 932 4990 933
rect 4986 929 4988 932
rect 5211 931 5212 938
rect 5241 929 5242 942
rect 5270 938 5278 943
rect 5356 938 5380 943
rect 5260 932 5270 938
rect 5253 929 5260 932
rect 4463 917 4465 920
rect 4459 914 4462 916
rect 4457 913 4459 914
rect 4454 911 4457 913
rect 4452 910 4454 911
rect 4338 906 4348 908
rect 4383 906 4400 908
rect 4327 904 4338 906
rect 4261 900 4262 903
rect 4305 900 4307 904
rect 4319 902 4327 904
rect 4315 901 4319 902
rect 4394 900 4396 906
rect 4418 904 4419 906
rect 4486 904 4502 920
rect 4520 910 4542 929
rect 4580 920 4588 927
rect 4588 918 4595 920
rect 4595 914 4611 918
rect 4614 914 4615 929
rect 4933 928 4946 929
rect 4939 927 4946 928
rect 4971 927 4972 928
rect 4985 927 4986 929
rect 5109 927 5110 929
rect 4941 923 4942 926
rect 4946 924 4983 927
rect 4673 921 4704 922
rect 4664 920 4673 921
rect 4704 920 4711 921
rect 4971 920 4972 924
rect 4635 917 4664 920
rect 4711 917 4726 920
rect 4633 916 4635 917
rect 4626 914 4633 916
rect 4726 914 4738 917
rect 4943 915 4944 917
rect 4972 915 4973 920
rect 4977 915 4986 924
rect 5024 915 5033 924
rect 5108 922 5109 927
rect 5107 920 5108 922
rect 5106 918 5107 920
rect 5105 916 5106 918
rect 4968 914 4977 915
rect 4611 911 4977 914
rect 4614 910 4615 911
rect 4617 910 4619 911
rect 4753 910 4761 911
rect 4542 909 4544 910
rect 4419 900 4423 904
rect 4473 900 4486 904
rect 4544 903 4552 909
rect 4613 908 4617 910
rect 4761 906 4779 910
rect 4944 906 4945 909
rect 4974 906 4975 909
rect 4606 904 4611 906
rect 3877 895 3932 897
rect 4006 895 4012 899
rect 4026 898 4027 900
rect 4025 895 4026 897
rect 4031 896 4200 900
rect 4259 897 4261 900
rect 4256 896 4262 897
rect 4302 896 4305 900
rect 4136 895 4137 896
rect 4200 895 4262 896
rect 3625 862 3633 874
rect 3637 865 3639 894
rect 3709 893 3710 894
rect 3750 893 3751 894
rect 3877 893 3934 895
rect 4012 893 4013 895
rect 3704 889 3710 893
rect 3749 889 3750 893
rect 3789 889 3790 893
rect 3845 889 3852 893
rect 3877 892 3942 893
rect 3690 888 3710 889
rect 3690 878 3704 888
rect 3746 879 3749 889
rect 3787 878 3789 889
rect 3842 879 3845 889
rect 3674 866 3690 878
rect 3637 862 3640 865
rect 3671 862 3674 866
rect 3721 859 3730 868
rect 3742 866 3746 878
rect 3786 875 3787 878
rect 3841 875 3842 878
rect 3741 862 3742 866
rect 3636 857 3638 858
rect 3643 857 3649 859
rect 3637 853 3649 857
rect 3701 853 3707 859
rect 3713 857 3721 859
rect 3740 858 3741 862
rect 3782 859 3786 875
rect 3836 859 3841 875
rect 3854 864 3857 892
rect 3904 891 3930 892
rect 3928 861 3930 891
rect 3934 881 3942 892
rect 4013 879 4033 893
rect 4081 879 4095 894
rect 4124 881 4132 893
rect 4136 891 4170 893
rect 3989 876 3990 879
rect 4019 876 4020 879
rect 4033 877 4045 879
rect 4079 877 4081 879
rect 4033 875 4079 877
rect 3904 859 3930 861
rect 3934 859 3942 871
rect 3987 869 3989 875
rect 4017 870 4019 875
rect 3985 862 3987 869
rect 4014 862 4017 869
rect 3984 859 3985 862
rect 4013 859 4014 862
rect 4136 859 4138 891
rect 4168 875 4170 891
rect 4174 881 4182 893
rect 4256 891 4262 895
rect 4300 891 4302 895
rect 4314 891 4320 897
rect 4394 894 4400 900
rect 4423 896 4438 900
rect 4438 895 4439 896
rect 4452 895 4486 900
rect 4552 899 4558 903
rect 4603 902 4606 904
rect 4779 902 4799 906
rect 4870 902 4883 903
rect 4210 881 4211 889
rect 4254 881 4257 891
rect 4262 885 4268 891
rect 4294 881 4300 891
rect 4308 885 4314 891
rect 4397 883 4398 891
rect 4400 888 4406 894
rect 4439 893 4458 895
rect 4169 865 4170 874
rect 4174 872 4175 875
rect 4204 870 4210 880
rect 4249 870 4254 881
rect 4192 866 4204 870
rect 4248 867 4249 870
rect 4287 867 4294 881
rect 4437 872 4440 892
rect 4446 888 4452 893
rect 4470 888 4486 895
rect 4558 894 4569 899
rect 4597 898 4601 900
rect 4594 897 4597 898
rect 4591 895 4594 897
rect 4614 895 4617 900
rect 4799 897 4824 902
rect 4849 900 4867 902
rect 4888 900 4911 902
rect 4847 899 4859 900
rect 4911 899 4920 900
rect 4920 898 4921 899
rect 4945 898 4946 902
rect 4824 895 4829 897
rect 4840 895 4847 898
rect 4569 885 4600 894
rect 4617 893 4619 895
rect 4619 891 4621 893
rect 4829 891 4847 895
rect 4921 894 4928 898
rect 4975 897 4976 902
rect 5033 901 5042 915
rect 5103 911 5104 914
rect 5130 909 5162 913
rect 5097 903 5101 906
rect 5104 903 5110 909
rect 5130 904 5168 909
rect 5199 904 5253 929
rect 5356 922 5382 938
rect 5127 903 5168 904
rect 5084 901 5096 902
rect 5042 899 5046 901
rect 5064 900 5084 901
rect 5058 899 5064 900
rect 5084 895 5086 900
rect 5110 897 5116 903
rect 5144 899 5145 901
rect 4928 891 4934 894
rect 4946 891 4947 895
rect 4559 880 4600 885
rect 4621 888 4694 891
rect 4829 889 4846 891
rect 4621 885 4701 888
rect 4621 881 4694 885
rect 4701 881 4771 885
rect 4832 882 4840 889
rect 4846 887 4851 889
rect 4851 885 4855 887
rect 4934 885 4947 891
rect 4976 887 4978 895
rect 5082 892 5084 895
rect 5081 891 5082 892
rect 4559 876 4575 880
rect 4600 876 4618 880
rect 4621 876 4639 881
rect 4694 876 4799 881
rect 4618 875 4799 876
rect 4825 875 4832 882
rect 4855 876 4877 885
rect 4934 882 4948 885
rect 4947 881 4950 882
rect 4947 878 4948 881
rect 4950 880 4951 881
rect 4951 879 4960 880
rect 4978 879 4980 885
rect 5069 882 5081 891
rect 5063 881 5069 882
rect 5035 880 5051 881
rect 5059 880 5063 881
rect 5128 880 5143 899
rect 5156 897 5162 903
rect 5193 901 5199 904
rect 5207 903 5208 904
rect 5182 895 5193 901
rect 5206 899 5207 901
rect 5179 892 5182 895
rect 5178 891 5179 892
rect 5170 885 5178 891
rect 5007 879 5030 880
rect 4877 875 4880 876
rect 4286 866 4287 867
rect 4191 865 4192 866
rect 4169 862 4191 865
rect 4245 862 4248 866
rect 4170 859 4191 862
rect 4242 859 4248 862
rect 3712 855 3721 857
rect 3637 852 3646 853
rect 3637 850 3647 852
rect 3649 850 3655 853
rect 3647 847 3655 850
rect 3647 842 3651 847
rect 3700 840 3701 853
rect 3710 852 3721 855
rect 3708 851 3710 852
rect 3705 850 3708 851
rect 3712 850 3721 852
rect 3736 845 3740 858
rect 3779 846 3782 858
rect 3832 846 3836 858
rect 3852 851 3858 857
rect 3881 856 3885 859
rect 4175 858 4176 859
rect 3858 845 3864 851
rect 3876 845 3881 856
rect 3910 851 3916 857
rect 3983 855 3984 858
rect 4012 855 4013 858
rect 4242 857 4245 859
rect 4244 856 4245 857
rect 4240 855 4244 856
rect 3904 845 3910 851
rect 3918 847 3930 855
rect 4134 853 4135 855
rect 3732 841 3736 845
rect 3778 841 3779 845
rect 3830 842 3832 845
rect 3730 840 3732 841
rect 3874 840 3876 845
rect 3978 841 3981 850
rect 4008 841 4011 850
rect 4135 841 4137 849
rect 4176 842 4177 849
rect 4237 847 4244 855
rect 4231 845 4238 847
rect 4240 845 4244 847
rect 4274 845 4286 865
rect 4398 859 4400 872
rect 4231 840 4240 845
rect 4271 844 4278 845
rect 4433 844 4437 870
rect 4548 869 4558 875
rect 4611 872 4811 875
rect 4822 872 4825 875
rect 4880 872 4890 875
rect 4896 872 4908 878
rect 4951 875 5030 879
rect 5158 876 5190 885
rect 5203 880 5206 898
rect 5202 876 5203 880
rect 5238 878 5240 904
rect 5356 895 5379 922
rect 5411 895 5412 929
rect 5356 881 5378 895
rect 5390 889 5412 895
rect 4611 871 4619 872
rect 4606 869 4610 871
rect 4546 868 4548 869
rect 4543 866 4546 868
rect 4601 866 4605 868
rect 4694 867 4918 872
rect 4948 871 4949 875
rect 4960 871 5007 875
rect 5121 872 5124 876
rect 5155 875 5190 876
rect 4966 869 5007 871
rect 4972 868 4997 869
rect 4710 866 4918 867
rect 4536 862 4543 866
rect 4591 862 4601 866
rect 4710 863 4920 866
rect 4823 862 4832 863
rect 4906 862 4928 863
rect 4949 862 4950 868
rect 4973 867 4997 868
rect 5113 863 5121 872
rect 5168 869 5169 874
rect 4530 858 4536 862
rect 4832 858 4839 862
rect 4528 857 4530 858
rect 4519 852 4528 857
rect 4839 852 4850 858
rect 4906 854 4920 862
rect 4928 856 4961 862
rect 4980 859 4981 862
rect 5109 857 5113 862
rect 5036 856 5048 857
rect 4961 855 4967 856
rect 4985 855 5007 856
rect 4967 854 5007 855
rect 5028 854 5048 856
rect 4514 850 4519 852
rect 4850 850 4854 852
rect 4479 849 4485 850
rect 4512 849 4514 850
rect 4461 844 4512 849
rect 4525 844 4531 850
rect 4575 845 4578 849
rect 4855 845 4863 849
rect 4906 846 4918 854
rect 5036 852 5068 854
rect 4951 850 4952 852
rect 4981 850 4982 852
rect 5037 847 5068 852
rect 5106 849 5108 856
rect 5106 847 5107 849
rect 4271 840 4275 844
rect 3652 836 3653 840
rect 3653 833 3654 836
rect 3700 832 3702 840
rect 3718 832 3730 840
rect 3777 838 3778 840
rect 3829 838 3830 840
rect 3776 832 3777 838
rect 3828 833 3829 838
rect 3871 832 3874 840
rect 3977 837 3978 840
rect 3976 833 3977 836
rect 4005 834 4007 840
rect 4177 837 4178 840
rect 4138 832 4142 837
rect 4229 832 4238 840
rect 4267 834 4275 840
rect 4267 832 4271 834
rect 3654 817 3662 832
rect 3700 825 3704 832
rect 3716 828 3718 832
rect 3775 828 3776 832
rect 3826 828 3827 832
rect 3702 817 3704 825
rect 3713 819 3716 828
rect 3773 819 3775 828
rect 3824 824 3826 827
rect 3820 820 3826 824
rect 3662 809 3666 817
rect 3704 811 3705 817
rect 3712 815 3713 819
rect 3772 815 3773 819
rect 3820 815 3824 820
rect 3866 819 3871 832
rect 3711 809 3712 814
rect 3770 809 3772 814
rect 3820 809 3822 815
rect 3863 814 3866 818
rect 3916 814 3932 824
rect 3934 814 3950 824
rect 3970 817 3976 832
rect 3859 809 3863 814
rect 3903 809 3910 814
rect 3955 808 3963 814
rect 3968 811 3970 817
rect 3998 811 4005 832
rect 4139 827 4143 832
rect 4178 827 4184 832
rect 3997 809 3998 811
rect 4012 808 4028 824
rect 4128 822 4194 827
rect 4214 824 4229 832
rect 4128 821 4184 822
rect 4119 814 4128 821
rect 4139 818 4143 821
rect 4035 808 4054 809
rect 4060 808 4062 809
rect 3667 804 3668 807
rect 3668 799 3670 803
rect 3705 799 3706 803
rect 3708 800 3711 808
rect 3768 800 3770 808
rect 3670 794 3672 798
rect 3708 794 3710 800
rect 3766 794 3768 798
rect 3673 785 3676 793
rect 3707 790 3709 793
rect 3710 790 3724 794
rect 3707 786 3724 790
rect 3676 775 3681 785
rect 3681 771 3682 775
rect 3708 774 3724 786
rect 3758 790 3766 794
rect 3804 792 3820 808
rect 3854 801 3859 808
rect 3899 801 3903 808
rect 3955 807 3966 808
rect 3996 807 4012 808
rect 4062 807 4063 808
rect 4111 807 4119 814
rect 4142 811 4143 817
rect 4178 811 4184 821
rect 4194 814 4198 821
rect 4212 819 4229 824
rect 4260 819 4267 832
rect 4269 828 4271 832
rect 4400 832 4402 844
rect 4412 840 4424 844
rect 4440 842 4461 844
rect 4431 841 4440 842
rect 4426 840 4433 841
rect 4412 836 4426 840
rect 4212 818 4214 819
rect 4212 815 4213 818
rect 4258 817 4260 819
rect 4257 816 4258 817
rect 4198 812 4202 814
rect 4211 812 4212 813
rect 4257 812 4260 816
rect 4290 812 4302 815
rect 4184 809 4185 811
rect 4139 808 4141 809
rect 4198 808 4209 812
rect 4256 808 4257 812
rect 4290 808 4306 812
rect 4308 808 4324 824
rect 4326 808 4342 824
rect 4400 820 4408 832
rect 4412 831 4428 832
rect 4412 830 4422 831
rect 4344 808 4353 812
rect 4403 810 4404 814
rect 4128 807 4138 808
rect 3955 806 3967 807
rect 3962 804 3967 806
rect 3995 804 4012 807
rect 4063 806 4066 807
rect 3854 792 3858 801
rect 3758 774 3774 790
rect 3804 774 3820 790
rect 3854 787 3870 790
rect 3849 781 3870 787
rect 3890 787 3899 801
rect 3962 792 3966 804
rect 3994 799 3995 803
rect 3992 794 3994 798
rect 3996 792 4012 804
rect 4035 798 4047 806
rect 4066 804 4069 806
rect 4099 804 4128 807
rect 4050 799 4099 804
rect 4100 799 4106 804
rect 4111 799 4119 804
rect 4185 799 4187 804
rect 4196 803 4211 808
rect 4256 806 4261 808
rect 4290 807 4307 808
rect 4312 807 4324 808
rect 3890 785 3901 787
rect 3910 785 3922 791
rect 3962 785 3963 792
rect 3990 788 3992 792
rect 3879 783 3901 785
rect 3911 783 3922 785
rect 3961 783 3966 785
rect 3873 781 3878 783
rect 3843 775 3849 781
rect 3854 774 3870 781
rect 3888 779 3890 783
rect 3895 781 3901 783
rect 3922 781 3926 783
rect 3901 775 3907 781
rect 3910 778 3922 779
rect 3710 771 3714 774
rect 3682 754 3690 771
rect 3714 754 3721 771
rect 3724 758 3740 774
rect 3742 758 3758 774
rect 3820 772 3828 774
rect 3846 772 3854 774
rect 3920 772 3922 778
rect 3926 772 3934 779
rect 3959 778 3961 783
rect 3962 778 3966 783
rect 3959 774 3966 778
rect 3959 772 3961 774
rect 3820 758 3836 772
rect 3838 758 3854 772
rect 3901 757 3964 772
rect 3988 760 3990 786
rect 3996 774 4012 790
rect 4023 782 4031 794
rect 4035 793 4056 794
rect 4094 793 4100 799
rect 4035 792 4053 793
rect 4012 763 4016 767
rect 4023 763 4031 772
rect 4035 763 4037 792
rect 4188 788 4190 796
rect 4196 794 4218 803
rect 4196 792 4211 794
rect 4248 792 4261 806
rect 4286 804 4288 807
rect 4292 806 4306 807
rect 4290 803 4306 806
rect 4342 805 4358 808
rect 4340 803 4358 805
rect 4248 790 4256 792
rect 4278 791 4286 803
rect 4288 801 4324 803
rect 4288 793 4308 801
rect 4321 800 4324 801
rect 4322 793 4324 800
rect 4328 799 4336 803
rect 4340 799 4362 803
rect 4342 794 4362 799
rect 4400 798 4408 810
rect 4412 800 4414 830
rect 4431 826 4433 840
rect 4473 838 4479 844
rect 4531 838 4537 844
rect 4570 841 4575 845
rect 4863 841 4868 845
rect 4862 832 4870 841
rect 4874 834 4876 839
rect 4906 834 4908 846
rect 5166 845 5168 865
rect 5200 863 5202 872
rect 5237 863 5238 872
rect 5356 868 5373 881
rect 5401 868 5406 872
rect 5356 866 5365 868
rect 5356 865 5364 866
rect 5390 865 5398 866
rect 5199 857 5200 862
rect 5197 849 5198 855
rect 4918 844 4926 845
rect 4874 832 4908 834
rect 4912 832 4926 844
rect 4446 826 4447 832
rect 4918 830 4926 832
rect 4557 829 4560 830
rect 4533 827 4568 829
rect 4431 818 4432 826
rect 4529 825 4533 827
rect 4432 800 4435 814
rect 4447 812 4449 825
rect 4500 808 4529 825
rect 4531 814 4533 817
rect 4541 812 4557 827
rect 4536 811 4557 812
rect 4568 824 4728 827
rect 4412 798 4446 800
rect 4432 795 4435 798
rect 4190 778 4193 788
rect 4193 769 4195 778
rect 4196 774 4211 790
rect 4248 774 4262 790
rect 4285 781 4286 788
rect 4195 765 4196 769
rect 4012 762 4037 763
rect 4066 762 4069 763
rect 4012 760 4069 762
rect 4012 758 4028 760
rect 4196 759 4197 763
rect 3690 746 3693 754
rect 3721 748 3726 754
rect 3726 745 3730 748
rect 3920 745 3922 757
rect 3925 745 3959 757
rect 3964 756 3966 757
rect 4073 756 4100 759
rect 4197 757 4198 759
rect 4212 758 4228 772
rect 4230 758 4246 772
rect 4278 769 4286 781
rect 4290 774 4308 793
rect 4342 792 4358 794
rect 4342 774 4358 790
rect 4388 774 4403 790
rect 4405 775 4407 789
rect 4412 786 4424 794
rect 4434 786 4446 794
rect 4448 790 4449 808
rect 4535 805 4545 811
rect 4568 808 4734 824
rect 4796 808 4812 824
rect 4814 808 4830 824
rect 4874 820 4886 828
rect 4896 820 4908 828
rect 4874 810 4876 820
rect 4926 816 4930 830
rect 4952 828 4954 845
rect 4954 819 4955 828
rect 4982 819 4985 845
rect 4987 843 5036 845
rect 5071 843 5073 844
rect 4987 833 5029 843
rect 5107 838 5108 843
rect 5074 827 5075 836
rect 5108 827 5109 836
rect 5165 834 5166 844
rect 5196 843 5197 847
rect 5195 837 5196 843
rect 5024 811 5029 823
rect 5076 817 5077 820
rect 5109 816 5110 820
rect 5164 819 5165 832
rect 5193 827 5195 836
rect 5235 829 5237 862
rect 5348 855 5364 865
rect 5401 864 5405 868
rect 5285 845 5348 855
rect 5393 851 5401 864
rect 5276 844 5285 845
rect 5270 842 5276 844
rect 5260 834 5270 842
rect 5192 821 5193 826
rect 5233 820 5235 827
rect 5077 811 5078 814
rect 5110 811 5111 814
rect 5163 811 5164 818
rect 5177 811 5183 817
rect 5191 816 5192 820
rect 5232 818 5233 820
rect 5240 818 5260 834
rect 5190 814 5191 816
rect 5189 812 5190 814
rect 5223 811 5229 817
rect 5231 813 5240 818
rect 5230 811 5240 813
rect 4986 808 4987 810
rect 5078 808 5079 810
rect 4540 803 4545 805
rect 4665 803 4674 808
rect 4712 803 4721 808
rect 4452 802 4461 803
rect 4450 798 4458 802
rect 4461 799 4476 802
rect 4476 798 4479 799
rect 4473 792 4479 798
rect 4531 792 4537 798
rect 4545 794 4554 803
rect 4656 794 4665 803
rect 4721 794 4730 803
rect 4647 792 4654 793
rect 4479 790 4485 792
rect 4290 772 4324 774
rect 4337 772 4342 774
rect 4435 772 4438 786
rect 4448 774 4454 790
rect 4479 786 4500 790
rect 4525 786 4531 792
rect 4641 791 4647 792
rect 4698 791 4702 793
rect 4734 792 4750 808
rect 4780 792 4796 808
rect 4807 803 4813 808
rect 4807 802 4822 803
rect 4801 796 4807 802
rect 4830 798 4846 808
rect 4853 802 4859 808
rect 4806 791 4807 793
rect 4839 791 4844 798
rect 4859 796 4865 802
rect 4877 800 4878 808
rect 4639 790 4641 791
rect 4638 787 4639 790
rect 4703 789 4705 790
rect 4484 774 4500 786
rect 4551 778 4578 781
rect 4534 774 4551 778
rect 4578 774 4586 778
rect 4290 769 4342 772
rect 4403 769 4409 772
rect 4438 771 4442 772
rect 4290 757 4294 765
rect 4326 758 4342 769
rect 4404 762 4421 769
rect 4438 762 4448 771
rect 4404 758 4420 762
rect 4421 760 4426 762
rect 4430 760 4442 762
rect 4426 759 4442 760
rect 4422 758 4442 759
rect 4500 758 4516 774
rect 4586 772 4589 774
rect 4654 772 4660 778
rect 4663 772 4665 779
rect 4705 772 4706 778
rect 4734 774 4750 790
rect 4780 774 4796 790
rect 4798 779 4807 791
rect 4733 772 4734 774
rect 4589 763 4609 772
rect 4638 767 4639 769
rect 4648 766 4654 772
rect 4706 766 4712 772
rect 4727 763 4734 772
rect 4609 762 4611 763
rect 4611 759 4617 762
rect 3966 751 3987 756
rect 3987 747 4003 751
rect 4035 748 4047 756
rect 4198 754 4199 756
rect 4094 747 4100 753
rect 4125 747 4180 753
rect 4199 750 4200 754
rect 4200 747 4202 748
rect 4209 747 4218 756
rect 4288 747 4294 756
rect 4346 747 4352 753
rect 4353 747 4362 756
rect 4407 751 4410 758
rect 3693 741 3695 745
rect 3730 740 3738 745
rect 3956 742 3957 745
rect 4003 742 4023 747
rect 4023 741 4028 742
rect 4100 741 4106 747
rect 4146 741 4152 747
rect 3922 740 3924 741
rect 3695 737 3697 740
rect 3738 737 3743 740
rect 3912 739 3922 740
rect 3901 738 3922 739
rect 4028 738 4032 741
rect 4153 738 4162 747
rect 4200 745 4209 747
rect 4200 742 4215 745
rect 4200 738 4209 742
rect 4215 740 4219 742
rect 4294 741 4306 747
rect 4340 741 4353 747
rect 4409 744 4410 751
rect 4219 739 4222 740
rect 3743 736 3745 737
rect 3910 736 3929 738
rect 3698 733 3699 736
rect 3745 733 3749 736
rect 3699 727 3702 733
rect 3749 731 3753 733
rect 3753 729 3756 731
rect 3843 729 3849 735
rect 3901 729 3907 735
rect 3910 733 3947 736
rect 3954 733 3955 736
rect 3921 729 3947 733
rect 3950 729 3954 731
rect 3986 729 3987 730
rect 3756 726 3760 729
rect 3702 720 3706 726
rect 3760 720 3770 726
rect 3773 720 3785 724
rect 3849 723 3855 729
rect 3895 723 3901 729
rect 3947 726 3987 729
rect 3947 723 3986 726
rect 4032 725 4049 738
rect 4153 737 4154 738
rect 4222 736 4229 739
rect 4297 738 4306 741
rect 4344 738 4353 741
rect 4403 739 4410 744
rect 4438 742 4442 758
rect 4480 747 4489 756
rect 4545 747 4554 756
rect 4617 754 4628 759
rect 4721 758 4734 763
rect 4796 772 4797 774
rect 4796 769 4805 772
rect 4806 769 4807 779
rect 4796 763 4807 769
rect 4810 763 4812 791
rect 4878 790 4880 791
rect 4876 785 4880 790
rect 4929 790 4930 808
rect 5036 799 5048 804
rect 5080 796 5081 799
rect 5111 796 5112 805
rect 5162 799 5163 808
rect 5171 805 5177 811
rect 5229 808 5235 811
rect 5284 808 5300 824
rect 5873 819 5874 1015
rect 6063 819 6064 1015
rect 6149 819 6150 1015
rect 6422 819 6423 1015
rect 6619 819 6620 1015
rect 7011 1014 7015 1019
rect 7649 1014 7656 1019
rect 7736 1018 7745 1027
rect 7801 1024 7897 1027
rect 8238 1023 8346 1037
rect 8096 1015 8112 1022
rect 8114 1015 8130 1022
rect 7656 1007 7668 1014
rect 8086 1013 8098 1015
rect 8108 1013 8120 1015
rect 8126 1013 8130 1015
rect 8314 1013 8330 1022
rect 8346 1021 8364 1023
rect 8365 1017 8372 1020
rect 8372 1013 8378 1017
rect 9018 1015 9019 1026
rect 9208 1015 9209 1026
rect 9294 1015 9295 1026
rect 9567 1015 9568 1026
rect 9764 1015 9765 1026
rect 10191 1023 10292 1034
rect 10478 1033 10742 1034
rect 10742 1023 10797 1033
rect 10900 1027 10909 1036
rect 10947 1027 10956 1036
rect 11250 1034 11372 1037
rect 11222 1033 11239 1034
rect 11052 1027 11222 1033
rect 10176 1021 10191 1023
rect 10170 1019 10176 1021
rect 10799 1019 10804 1021
rect 8086 1008 8130 1013
rect 8273 1008 8310 1009
rect 8378 1008 8381 1013
rect 8082 1006 8084 1008
rect 8086 1006 8218 1008
rect 7137 1005 7491 1006
rect 7117 1003 7135 1005
rect 7577 1003 7590 1005
rect 7669 1003 7672 1005
rect 8080 1003 8218 1006
rect 7061 1000 7117 1003
rect 6935 992 6947 1000
rect 6957 992 6969 1000
rect 7033 994 7117 1000
rect 7590 994 7600 1003
rect 7033 993 7061 994
rect 6931 989 6933 992
rect 7033 991 7052 993
rect 7601 991 7604 993
rect 6973 988 6977 989
rect 6923 977 6931 988
rect 6934 986 6969 988
rect 6932 977 6934 983
rect 6923 976 6932 977
rect 6931 972 6932 976
rect 6930 971 6931 972
rect 6928 966 6930 969
rect 6803 964 6868 965
rect 6795 956 6803 964
rect 6868 956 6872 964
rect 6794 950 6795 956
rect 6923 954 6931 966
rect 6935 956 6937 986
rect 6966 985 6969 986
rect 6968 979 6969 985
rect 6973 981 6981 988
rect 6977 980 6985 981
rect 7009 980 7010 990
rect 7033 980 7048 991
rect 7307 981 7344 983
rect 6985 979 6991 980
rect 7008 979 7009 980
rect 7033 979 7040 980
rect 6991 969 7053 979
rect 7061 972 7067 978
rect 7107 972 7113 978
rect 7307 977 7333 981
rect 7344 977 7349 981
rect 7604 980 7617 991
rect 7580 979 7594 980
rect 7301 972 7307 977
rect 7349 972 7358 977
rect 7562 972 7580 979
rect 7594 977 7601 979
rect 7672 977 7693 1003
rect 8074 996 8218 1003
rect 8234 1006 8335 1008
rect 8234 996 8346 1006
rect 8035 990 8096 996
rect 8000 987 8035 990
rect 7813 981 8000 987
rect 8086 986 8096 990
rect 7601 972 7616 977
rect 7055 969 7061 972
rect 7062 970 7119 972
rect 7358 971 7359 972
rect 7196 970 7199 971
rect 7217 970 7220 971
rect 7299 970 7300 971
rect 7359 970 7362 971
rect 7062 969 7070 970
rect 7033 968 7070 969
rect 6935 954 6969 956
rect 6924 951 6926 954
rect 6920 938 6924 950
rect 6935 942 6947 950
rect 6960 945 6969 954
rect 7007 952 7008 955
rect 7033 951 7038 968
rect 7055 966 7070 968
rect 7113 966 7119 970
rect 7195 969 7196 970
rect 7220 969 7221 970
rect 7554 969 7562 972
rect 7591 971 7616 972
rect 7625 971 7629 972
rect 7587 970 7591 971
rect 7601 970 7638 971
rect 7586 969 7587 970
rect 7192 967 7195 969
rect 7221 967 7225 969
rect 7362 968 7363 969
rect 7363 967 7366 968
rect 7061 964 7070 966
rect 7188 965 7192 967
rect 7225 965 7229 967
rect 7546 966 7554 969
rect 7584 968 7586 969
rect 7580 967 7584 968
rect 7575 965 7580 967
rect 7601 965 7616 970
rect 7625 969 7629 970
rect 7638 969 7639 970
rect 7695 969 7700 975
rect 7736 971 7745 980
rect 7801 978 7813 981
rect 7801 971 7810 978
rect 8080 972 8096 986
rect 8119 972 8120 996
rect 8125 991 8146 996
rect 8130 990 8146 991
rect 8263 989 8269 996
rect 8315 989 8321 996
rect 8335 990 8346 996
rect 8381 990 8390 1008
rect 8130 972 8146 988
rect 8263 985 8271 989
rect 8269 983 8271 985
rect 8200 977 8207 978
rect 8209 977 8211 978
rect 8179 974 8200 977
rect 8211 974 8220 977
rect 8177 972 8179 974
rect 8220 972 8222 974
rect 7629 965 7634 969
rect 7639 965 7641 968
rect 7700 965 7703 969
rect 7186 964 7188 965
rect 7229 964 7231 965
rect 7541 964 7545 965
rect 7616 964 7619 965
rect 7641 964 7642 965
rect 7061 951 7066 964
rect 7114 955 7133 958
rect 7172 956 7186 964
rect 7231 959 7243 964
rect 7298 959 7299 964
rect 7243 956 7246 959
rect 7366 957 7369 964
rect 7537 962 7541 964
rect 7168 955 7172 956
rect 6970 949 6975 950
rect 6975 948 6980 949
rect 6980 947 6983 948
rect 6985 945 6994 947
rect 6958 942 6960 945
rect 6994 944 6999 945
rect 6999 943 7005 944
rect 7006 943 7007 951
rect 7033 943 7039 951
rect 6957 939 6958 942
rect 7005 938 7039 943
rect 6918 931 6920 937
rect 6955 930 6957 938
rect 7006 932 7007 938
rect 7033 935 7061 938
rect 7033 933 7063 935
rect 7033 931 7064 933
rect 7065 931 7066 951
rect 7133 946 7195 955
rect 7246 952 7251 956
rect 7297 951 7298 956
rect 7369 954 7370 956
rect 7506 950 7537 962
rect 7621 959 7625 962
rect 7636 960 7640 963
rect 7745 962 7754 971
rect 7778 961 7781 963
rect 7792 962 7801 971
rect 8086 970 8120 972
rect 8129 971 8130 972
rect 8176 971 8177 972
rect 8125 970 8130 971
rect 8175 970 8176 971
rect 8086 968 8130 970
rect 8173 969 8175 970
rect 8222 969 8225 972
rect 8082 965 8083 967
rect 7856 961 7865 963
rect 7773 959 7778 961
rect 7151 945 7161 946
rect 7183 945 7184 946
rect 7147 943 7151 945
rect 7195 943 7215 946
rect 7296 943 7297 950
rect 7369 943 7370 950
rect 7504 949 7506 950
rect 7418 943 7424 949
rect 7464 948 7470 949
rect 7501 948 7504 949
rect 7464 947 7501 948
rect 7464 943 7470 947
rect 7556 946 7562 952
rect 7602 946 7608 952
rect 7624 950 7625 959
rect 7771 958 7773 959
rect 7867 958 7873 961
rect 7642 955 7646 958
rect 7710 955 7712 958
rect 7873 956 7876 958
rect 8096 956 8112 968
rect 8114 956 8130 968
rect 8169 965 8173 968
rect 8225 965 8229 969
rect 8269 967 8272 983
rect 8168 964 8169 965
rect 8229 964 8230 965
rect 8167 963 8168 964
rect 8165 961 8167 963
rect 8230 961 8233 964
rect 8271 961 8272 967
rect 8275 967 8276 989
rect 8314 985 8321 989
rect 8342 987 8344 990
rect 8314 983 8315 985
rect 8335 984 8336 986
rect 8275 963 8277 967
rect 8308 963 8309 966
rect 8313 965 8315 983
rect 8344 981 8347 987
rect 8347 979 8348 981
rect 8349 975 8350 977
rect 8350 972 8351 975
rect 8390 973 8398 990
rect 8352 965 8355 969
rect 8275 961 8279 963
rect 8313 962 8314 965
rect 8355 963 8356 965
rect 8161 958 8164 961
rect 8233 959 8236 961
rect 8160 956 8161 958
rect 8236 957 8238 959
rect 7646 946 7656 955
rect 7135 931 7143 943
rect 7147 941 7181 943
rect 6871 924 6872 929
rect 6821 915 6830 924
rect 6868 920 6877 924
rect 6868 915 6882 920
rect 6812 912 6821 915
rect 6812 911 6815 912
rect 6805 908 6814 911
rect 6793 907 6814 908
rect 6793 905 6811 907
rect 6851 905 6857 911
rect 6871 906 6886 915
rect 6911 908 6918 929
rect 6793 900 6805 905
rect 6789 898 6792 900
rect 6793 899 6794 900
rect 6799 899 6805 900
rect 6857 899 6863 905
rect 6870 904 6882 906
rect 6909 904 6911 908
rect 6949 907 6955 929
rect 7006 926 7007 929
rect 7033 928 7094 931
rect 7033 917 7039 928
rect 7061 926 7094 928
rect 7055 925 7094 926
rect 7113 925 7119 926
rect 7055 921 7119 925
rect 7055 920 7141 921
rect 7033 913 7042 917
rect 7061 914 7067 920
rect 7107 914 7113 920
rect 7116 917 7141 920
rect 7125 913 7141 917
rect 7147 913 7149 941
rect 7178 939 7181 941
rect 7033 909 7048 913
rect 7135 909 7149 913
rect 7179 909 7181 939
rect 7185 931 7193 943
rect 7215 934 7278 943
rect 7412 938 7418 943
rect 7430 941 7466 943
rect 7430 938 7435 941
rect 7371 937 7418 938
rect 7432 937 7435 938
rect 7470 937 7476 943
rect 7550 940 7556 946
rect 7608 940 7614 946
rect 7371 936 7414 937
rect 7295 934 7296 936
rect 7317 934 7371 936
rect 7251 922 7266 934
rect 7278 933 7317 934
rect 7295 929 7296 933
rect 7427 929 7430 936
rect 7554 933 7556 934
rect 7552 929 7554 933
rect 6948 904 6949 906
rect 7008 905 7009 909
rect 6868 899 6870 904
rect 7014 903 7020 909
rect 7033 903 7052 909
rect 7060 903 7066 909
rect 6908 899 6909 903
rect 6867 897 6868 899
rect 6907 897 6908 899
rect 6781 884 6789 896
rect 6793 894 6811 896
rect 6866 895 6867 896
rect 6946 895 6948 903
rect 7008 897 7014 903
rect 7033 897 7072 903
rect 7074 897 7086 905
rect 7147 904 7164 909
rect 7155 899 7162 904
rect 7164 903 7168 904
rect 7184 903 7185 905
rect 7251 904 7266 920
rect 7293 906 7295 928
rect 7168 900 7187 903
rect 7292 900 7304 905
rect 7314 900 7326 905
rect 7367 904 7369 928
rect 7418 904 7427 928
rect 7463 904 7466 909
rect 7504 908 7539 910
rect 7550 908 7552 929
rect 7574 909 7575 929
rect 7622 928 7624 944
rect 7656 942 7661 946
rect 7712 942 7724 955
rect 7876 951 7886 956
rect 8159 953 8160 956
rect 7994 952 8031 953
rect 8158 952 8159 953
rect 8238 952 8240 956
rect 8266 955 8272 961
rect 8279 959 8285 961
rect 8286 957 8292 959
rect 8292 956 8295 957
rect 8312 956 8318 961
rect 8356 960 8357 963
rect 8357 958 8358 960
rect 7994 951 8019 952
rect 8031 951 8032 952
rect 8157 951 8158 952
rect 7888 948 7892 951
rect 7959 948 7986 951
rect 8034 948 8041 951
rect 8041 943 8052 948
rect 8087 945 8089 949
rect 8122 947 8123 949
rect 8155 948 8157 951
rect 8052 942 8056 943
rect 7724 939 7725 942
rect 8056 938 8063 942
rect 7666 929 7676 938
rect 7726 931 7732 938
rect 8063 937 8065 938
rect 8065 933 8081 937
rect 8081 932 8086 933
rect 8089 932 8097 944
rect 8086 929 8097 932
rect 8123 929 8127 944
rect 8153 943 8155 948
rect 8240 944 8243 951
rect 8260 949 8266 955
rect 8295 951 8336 956
rect 8358 955 8360 958
rect 8318 949 8324 951
rect 8360 948 8363 955
rect 8152 942 8153 943
rect 8363 942 8366 948
rect 8398 943 8399 973
rect 8506 951 8522 954
rect 8434 943 8457 951
rect 8512 943 8529 951
rect 8151 940 8152 942
rect 8150 939 8151 940
rect 8366 939 8367 942
rect 8149 937 8150 938
rect 8146 933 8149 937
rect 8144 932 8146 933
rect 8142 929 8144 932
rect 8367 931 8368 938
rect 8397 929 8398 942
rect 8426 938 8434 943
rect 8512 938 8536 943
rect 8416 932 8426 938
rect 8409 929 8416 932
rect 7619 917 7621 920
rect 7615 914 7618 916
rect 7613 913 7615 914
rect 7610 911 7613 913
rect 7608 910 7610 911
rect 7494 906 7504 908
rect 7539 906 7556 908
rect 7483 904 7494 906
rect 7417 900 7418 903
rect 7461 900 7463 904
rect 7475 902 7483 904
rect 7471 901 7475 902
rect 7550 900 7552 906
rect 7574 904 7575 906
rect 7642 904 7658 920
rect 7676 910 7698 929
rect 7736 920 7744 927
rect 7744 918 7751 920
rect 7751 914 7767 918
rect 7770 914 7771 929
rect 8089 928 8102 929
rect 8095 927 8102 928
rect 8127 927 8128 928
rect 8141 927 8142 929
rect 8265 927 8266 929
rect 8097 923 8098 926
rect 8102 924 8139 927
rect 7829 921 7860 922
rect 7820 920 7829 921
rect 7860 920 7867 921
rect 8127 920 8128 924
rect 7791 917 7820 920
rect 7867 917 7882 920
rect 7789 916 7791 917
rect 7782 914 7789 916
rect 7882 914 7894 917
rect 8099 915 8100 917
rect 8128 915 8129 920
rect 8133 915 8142 924
rect 8180 915 8189 924
rect 8264 922 8265 927
rect 8263 920 8264 922
rect 8262 918 8263 920
rect 8261 916 8262 918
rect 8124 914 8133 915
rect 7767 911 8133 914
rect 7770 910 7771 911
rect 7773 910 7775 911
rect 7909 910 7917 911
rect 7698 909 7700 910
rect 7575 900 7579 904
rect 7629 900 7642 904
rect 7700 903 7708 909
rect 7769 908 7773 910
rect 7917 906 7935 910
rect 8100 906 8101 909
rect 8130 906 8131 909
rect 7762 904 7767 906
rect 7033 895 7088 897
rect 7162 895 7168 899
rect 7182 898 7183 900
rect 7181 895 7182 897
rect 7187 896 7356 900
rect 7415 897 7417 900
rect 7412 896 7418 897
rect 7458 896 7461 900
rect 7292 895 7293 896
rect 7356 895 7418 896
rect 6781 862 6789 874
rect 6793 865 6795 894
rect 6865 893 6866 894
rect 6906 893 6907 894
rect 7033 893 7090 895
rect 7168 893 7169 895
rect 6860 889 6866 893
rect 6905 889 6906 893
rect 6945 889 6946 893
rect 7001 889 7008 893
rect 7033 892 7098 893
rect 6846 888 6866 889
rect 6846 878 6860 888
rect 6902 879 6905 889
rect 6943 878 6945 889
rect 6998 879 7001 889
rect 6830 866 6846 878
rect 6793 862 6796 865
rect 6827 862 6830 866
rect 6877 859 6886 868
rect 6898 866 6902 878
rect 6942 875 6943 878
rect 6997 875 6998 878
rect 6897 862 6898 866
rect 6792 857 6794 858
rect 6799 857 6805 859
rect 6793 853 6805 857
rect 6857 853 6863 859
rect 6869 857 6877 859
rect 6896 858 6897 862
rect 6938 859 6942 875
rect 6992 859 6997 875
rect 7010 864 7013 892
rect 7060 891 7086 892
rect 7084 861 7086 891
rect 7090 881 7098 892
rect 7169 879 7189 893
rect 7237 879 7251 894
rect 7280 881 7288 893
rect 7292 891 7326 893
rect 7145 876 7146 879
rect 7175 876 7176 879
rect 7189 877 7201 879
rect 7235 877 7237 879
rect 7189 875 7235 877
rect 7060 859 7086 861
rect 7090 859 7098 871
rect 7143 869 7145 875
rect 7173 870 7175 875
rect 7141 862 7143 869
rect 7170 862 7173 869
rect 7140 859 7141 862
rect 7169 859 7170 862
rect 7292 859 7294 891
rect 7324 875 7326 891
rect 7330 881 7338 893
rect 7412 891 7418 895
rect 7456 891 7458 895
rect 7470 891 7476 897
rect 7550 894 7556 900
rect 7579 896 7594 900
rect 7594 895 7595 896
rect 7608 895 7642 900
rect 7708 899 7714 903
rect 7759 902 7762 904
rect 7935 902 7955 906
rect 8026 902 8039 903
rect 7366 881 7367 889
rect 7410 881 7413 891
rect 7418 885 7424 891
rect 7450 881 7456 891
rect 7464 885 7470 891
rect 7553 883 7554 891
rect 7556 888 7562 894
rect 7595 893 7614 895
rect 7325 865 7326 874
rect 7330 872 7331 875
rect 7360 870 7366 880
rect 7405 870 7410 881
rect 7348 866 7360 870
rect 7404 867 7405 870
rect 7443 867 7450 881
rect 7593 872 7596 892
rect 7602 888 7608 893
rect 7626 888 7642 895
rect 7714 894 7725 899
rect 7753 898 7757 900
rect 7750 897 7753 898
rect 7747 895 7750 897
rect 7770 895 7773 900
rect 7955 897 7980 902
rect 8005 900 8023 902
rect 8044 900 8067 902
rect 8003 899 8015 900
rect 8067 899 8076 900
rect 8076 898 8077 899
rect 8101 898 8102 902
rect 7980 895 7985 897
rect 7996 895 8003 898
rect 7725 885 7756 894
rect 7773 893 7775 895
rect 7775 891 7777 893
rect 7985 891 8003 895
rect 8077 894 8084 898
rect 8131 897 8132 902
rect 8189 901 8198 915
rect 8259 911 8260 914
rect 8286 909 8318 913
rect 8253 903 8257 906
rect 8260 903 8266 909
rect 8286 904 8324 909
rect 8355 904 8409 929
rect 8512 922 8538 938
rect 8283 903 8324 904
rect 8240 901 8252 902
rect 8198 899 8202 901
rect 8220 900 8240 901
rect 8214 899 8220 900
rect 8240 895 8242 900
rect 8266 897 8272 903
rect 8300 899 8301 901
rect 8084 891 8090 894
rect 8102 891 8103 895
rect 7715 880 7756 885
rect 7777 888 7850 891
rect 7985 889 8002 891
rect 7777 885 7857 888
rect 7777 881 7850 885
rect 7857 881 7927 885
rect 7988 882 7996 889
rect 8002 887 8007 889
rect 8007 885 8011 887
rect 8090 885 8103 891
rect 8132 887 8134 895
rect 8238 892 8240 895
rect 8237 891 8238 892
rect 7715 876 7731 880
rect 7756 876 7774 880
rect 7777 876 7795 881
rect 7850 876 7955 881
rect 7774 875 7955 876
rect 7981 875 7988 882
rect 8011 876 8033 885
rect 8090 882 8104 885
rect 8103 881 8106 882
rect 8103 878 8104 881
rect 8106 880 8107 881
rect 8107 879 8116 880
rect 8134 879 8136 885
rect 8225 882 8237 891
rect 8219 881 8225 882
rect 8191 880 8207 881
rect 8215 880 8219 881
rect 8284 880 8299 899
rect 8312 897 8318 903
rect 8349 901 8355 904
rect 8363 903 8364 904
rect 8338 895 8349 901
rect 8362 899 8363 901
rect 8335 892 8338 895
rect 8334 891 8335 892
rect 8326 885 8334 891
rect 8163 879 8186 880
rect 8033 875 8036 876
rect 7442 866 7443 867
rect 7347 865 7348 866
rect 7325 862 7347 865
rect 7401 862 7404 866
rect 7326 859 7347 862
rect 7398 859 7404 862
rect 6868 855 6877 857
rect 6793 852 6802 853
rect 6793 850 6803 852
rect 6805 850 6811 853
rect 6803 847 6811 850
rect 6803 842 6807 847
rect 6856 840 6857 853
rect 6866 852 6877 855
rect 6864 851 6866 852
rect 6861 850 6864 851
rect 6868 850 6877 852
rect 6892 845 6896 858
rect 6935 846 6938 858
rect 6988 846 6992 858
rect 7008 851 7014 857
rect 7037 856 7041 859
rect 7331 858 7332 859
rect 7014 845 7020 851
rect 7032 845 7037 856
rect 7066 851 7072 857
rect 7139 855 7140 858
rect 7168 855 7169 858
rect 7398 857 7401 859
rect 7400 856 7401 857
rect 7396 855 7400 856
rect 7060 845 7066 851
rect 7074 847 7086 855
rect 7290 853 7291 855
rect 6888 841 6892 845
rect 6934 841 6935 845
rect 6986 842 6988 845
rect 6886 840 6888 841
rect 7030 840 7032 845
rect 7134 841 7137 850
rect 7164 841 7167 850
rect 7291 841 7293 849
rect 7332 842 7333 849
rect 7393 847 7400 855
rect 7387 845 7394 847
rect 7396 845 7400 847
rect 7430 845 7442 865
rect 7554 859 7556 872
rect 7387 840 7396 845
rect 7427 844 7434 845
rect 7589 844 7593 870
rect 7704 869 7714 875
rect 7767 872 7967 875
rect 7978 872 7981 875
rect 8036 872 8046 875
rect 8052 872 8064 878
rect 8107 875 8186 879
rect 8314 876 8346 885
rect 8359 880 8362 898
rect 8358 876 8359 880
rect 8394 878 8396 904
rect 8512 895 8535 922
rect 8567 895 8568 929
rect 8512 881 8534 895
rect 8546 889 8568 895
rect 7767 871 7775 872
rect 7762 869 7766 871
rect 7702 868 7704 869
rect 7699 866 7702 868
rect 7757 866 7761 868
rect 7850 867 8074 872
rect 8104 871 8105 875
rect 8116 871 8163 875
rect 8277 872 8280 876
rect 8311 875 8346 876
rect 8122 869 8163 871
rect 8128 868 8153 869
rect 7866 866 8074 867
rect 7692 862 7699 866
rect 7747 862 7757 866
rect 7866 863 8076 866
rect 7979 862 7988 863
rect 8062 862 8084 863
rect 8105 862 8106 868
rect 8129 867 8153 868
rect 8269 863 8277 872
rect 8324 869 8325 874
rect 7686 858 7692 862
rect 7988 858 7995 862
rect 7684 857 7686 858
rect 7675 852 7684 857
rect 7995 852 8006 858
rect 8062 854 8076 862
rect 8084 856 8117 862
rect 8136 859 8137 862
rect 8265 857 8269 862
rect 8192 856 8204 857
rect 8117 855 8123 856
rect 8141 855 8163 856
rect 8123 854 8163 855
rect 8184 854 8204 856
rect 7670 850 7675 852
rect 8006 850 8010 852
rect 7635 849 7641 850
rect 7668 849 7670 850
rect 7617 844 7668 849
rect 7681 844 7687 850
rect 7731 845 7734 849
rect 8011 845 8019 849
rect 8062 846 8074 854
rect 8192 852 8224 854
rect 8107 850 8108 852
rect 8137 850 8138 852
rect 8193 847 8224 852
rect 8262 849 8264 856
rect 8262 847 8263 849
rect 7427 840 7431 844
rect 6808 836 6809 840
rect 6809 833 6810 836
rect 6856 832 6858 840
rect 6874 832 6886 840
rect 6933 838 6934 840
rect 6985 838 6986 840
rect 6932 832 6933 838
rect 6984 833 6985 838
rect 7027 832 7030 840
rect 7133 837 7134 840
rect 7132 833 7133 836
rect 7161 834 7163 840
rect 7333 837 7334 840
rect 7294 832 7298 837
rect 7385 832 7394 840
rect 7423 834 7431 840
rect 7423 832 7427 834
rect 6810 817 6818 832
rect 6856 825 6860 832
rect 6872 828 6874 832
rect 6931 828 6932 832
rect 6982 828 6983 832
rect 6858 817 6860 825
rect 6869 819 6872 828
rect 6929 819 6931 828
rect 6980 824 6982 827
rect 6976 820 6982 824
rect 6818 809 6822 817
rect 6860 811 6861 817
rect 6868 815 6869 819
rect 6928 815 6929 819
rect 6976 815 6980 820
rect 7022 819 7027 832
rect 6867 809 6868 814
rect 6926 809 6928 814
rect 6976 809 6978 815
rect 7019 814 7022 818
rect 7072 814 7088 824
rect 7090 814 7106 824
rect 7126 817 7132 832
rect 7015 809 7019 814
rect 7059 809 7066 814
rect 7111 808 7119 814
rect 7124 811 7126 817
rect 7154 811 7161 832
rect 7295 827 7299 832
rect 7334 827 7340 832
rect 7153 809 7154 811
rect 7168 808 7184 824
rect 7284 822 7350 827
rect 7370 824 7385 832
rect 7284 821 7340 822
rect 7275 814 7284 821
rect 7295 818 7299 821
rect 7191 808 7210 809
rect 7216 808 7218 809
rect 5227 805 5235 808
rect 5227 804 5229 805
rect 5230 800 5231 802
rect 5231 797 5233 800
rect 4796 758 4812 763
rect 4861 773 4922 785
rect 4929 779 4942 790
rect 4928 774 4942 779
rect 4972 774 4987 790
rect 4988 777 4990 793
rect 5081 789 5082 793
rect 5112 789 5113 795
rect 4861 759 4926 773
rect 4892 758 4908 759
rect 4910 758 4926 759
rect 4953 758 4954 760
rect 4988 758 5004 774
rect 5082 767 5086 785
rect 5113 779 5114 788
rect 5162 787 5164 794
rect 5227 790 5228 794
rect 5233 791 5236 797
rect 5268 792 5284 808
rect 5318 802 5346 808
rect 6823 804 6824 807
rect 5312 794 5346 802
rect 6824 799 6826 803
rect 6861 799 6862 803
rect 6864 800 6867 808
rect 6924 800 6926 808
rect 6826 794 6828 798
rect 6864 794 6866 800
rect 6922 794 6924 798
rect 5308 791 5310 794
rect 5318 790 5346 794
rect 5164 781 5165 787
rect 5227 782 5244 790
rect 5114 766 5119 779
rect 5166 774 5174 780
rect 5228 776 5244 782
rect 5300 779 5308 790
rect 5297 778 5308 779
rect 5312 788 5346 790
rect 5228 774 5238 776
rect 5174 773 5176 774
rect 5176 772 5177 773
rect 5086 760 5087 766
rect 5119 759 5121 766
rect 5177 765 5190 772
rect 5228 766 5229 772
rect 5244 768 5249 776
rect 5297 770 5306 778
rect 5225 765 5229 766
rect 5171 764 5204 765
rect 5225 764 5235 765
rect 5171 759 5177 764
rect 4721 756 4727 758
rect 4798 757 4812 758
rect 4924 757 4927 758
rect 4806 756 4859 757
rect 4639 754 4640 756
rect 4721 754 4730 756
rect 4403 738 4409 739
rect 4449 738 4455 744
rect 4489 738 4498 747
rect 4536 738 4545 747
rect 4628 746 4642 754
rect 4716 747 4730 754
rect 4801 750 4865 756
rect 4928 750 4943 756
rect 4950 754 4951 756
rect 4992 752 4993 753
rect 4716 746 4721 747
rect 4642 745 4645 746
rect 4715 745 4721 746
rect 4155 734 4156 736
rect 4157 727 4160 733
rect 4229 731 4244 736
rect 4397 732 4403 738
rect 4455 733 4461 738
rect 4509 734 4521 738
rect 4562 734 4578 744
rect 4640 742 4641 745
rect 4645 742 4684 745
rect 4714 743 4715 745
rect 4641 740 4684 742
rect 4645 737 4684 740
rect 4707 739 4714 743
rect 4716 739 4721 745
rect 4807 745 4822 750
rect 4853 747 4862 750
rect 4807 744 4813 745
rect 4853 744 4859 747
rect 4862 742 4876 747
rect 4943 745 4956 750
rect 4992 747 5000 752
rect 5088 751 5089 756
rect 5122 750 5125 756
rect 5177 753 5183 759
rect 5188 758 5204 764
rect 5206 758 5222 764
rect 5229 759 5235 764
rect 5249 762 5252 768
rect 5288 761 5297 770
rect 5223 753 5229 759
rect 5254 756 5256 760
rect 5284 757 5285 758
rect 4942 742 4944 745
rect 4956 742 4962 745
rect 4993 744 5000 747
rect 5089 746 5090 750
rect 5125 744 5127 750
rect 5211 745 5214 747
rect 5002 742 5003 744
rect 5256 743 5264 756
rect 5285 754 5288 757
rect 5300 756 5308 768
rect 5312 758 5314 788
rect 5343 787 5346 788
rect 5350 779 5393 791
rect 6829 785 6832 793
rect 6863 790 6865 793
rect 6866 790 6880 794
rect 6863 786 6880 790
rect 5344 776 5393 779
rect 5344 770 5353 776
rect 5364 774 5380 776
rect 5393 774 5414 776
rect 6832 775 6837 785
rect 5353 764 5362 770
rect 5356 763 5362 764
rect 5380 768 5414 774
rect 6837 771 6838 775
rect 6864 774 6880 786
rect 6914 790 6922 794
rect 6960 792 6976 808
rect 7010 801 7015 808
rect 7055 801 7059 808
rect 7111 807 7122 808
rect 7152 807 7168 808
rect 7218 807 7219 808
rect 7267 807 7275 814
rect 7298 811 7299 817
rect 7334 811 7340 821
rect 7350 814 7354 821
rect 7368 819 7385 824
rect 7416 819 7423 832
rect 7425 828 7427 832
rect 7556 832 7558 844
rect 7568 840 7580 844
rect 7596 842 7617 844
rect 7587 841 7596 842
rect 7582 840 7589 841
rect 7568 836 7582 840
rect 7368 818 7370 819
rect 7368 815 7369 818
rect 7414 817 7416 819
rect 7413 816 7414 817
rect 7354 812 7358 814
rect 7367 812 7368 813
rect 7413 812 7416 816
rect 7446 812 7458 815
rect 7340 809 7341 811
rect 7295 808 7297 809
rect 7354 808 7365 812
rect 7412 808 7413 812
rect 7446 808 7462 812
rect 7464 808 7480 824
rect 7482 808 7498 824
rect 7556 820 7564 832
rect 7568 831 7584 832
rect 7568 830 7578 831
rect 7500 808 7509 812
rect 7559 810 7560 814
rect 7284 807 7294 808
rect 7111 806 7123 807
rect 7118 804 7123 806
rect 7151 804 7168 807
rect 7219 806 7222 807
rect 7010 792 7014 801
rect 6914 774 6930 790
rect 6960 774 6976 790
rect 7010 787 7026 790
rect 7005 781 7026 787
rect 7046 787 7055 801
rect 7118 792 7122 804
rect 7150 799 7151 803
rect 7148 794 7150 798
rect 7152 792 7168 804
rect 7191 798 7203 806
rect 7222 804 7225 806
rect 7255 804 7284 807
rect 7206 799 7255 804
rect 7256 799 7262 804
rect 7267 799 7275 804
rect 7341 799 7343 804
rect 7352 803 7367 808
rect 7412 806 7417 808
rect 7446 807 7463 808
rect 7468 807 7480 808
rect 7046 785 7057 787
rect 7066 785 7078 791
rect 7118 785 7119 792
rect 7146 788 7148 792
rect 7035 783 7057 785
rect 7067 783 7078 785
rect 7117 783 7122 785
rect 7029 781 7034 783
rect 6999 775 7005 781
rect 7010 774 7026 781
rect 7044 779 7046 783
rect 7051 781 7057 783
rect 7078 781 7082 783
rect 7057 775 7063 781
rect 7066 778 7078 779
rect 6866 771 6870 774
rect 5357 759 5360 763
rect 5380 758 5396 768
rect 5414 762 5431 768
rect 5417 758 5423 762
rect 5431 760 5437 762
rect 5437 758 5441 760
rect 5463 758 5469 764
rect 5312 757 5327 758
rect 5312 756 5331 757
rect 5288 750 5293 754
rect 5328 752 5346 756
rect 5363 753 5369 756
rect 5411 753 5417 758
rect 5312 750 5346 752
rect 5369 751 5417 753
rect 5469 752 5475 758
rect 6838 754 6846 771
rect 6870 754 6877 771
rect 6880 758 6896 774
rect 6898 758 6914 774
rect 6976 772 6984 774
rect 7002 772 7010 774
rect 7076 772 7078 778
rect 7082 772 7090 779
rect 7115 778 7117 783
rect 7118 778 7122 783
rect 7115 774 7122 778
rect 7115 772 7117 774
rect 6976 758 6992 772
rect 6994 758 7010 772
rect 7057 757 7120 772
rect 7144 760 7146 786
rect 7152 774 7168 790
rect 7179 782 7187 794
rect 7191 793 7212 794
rect 7250 793 7256 799
rect 7191 792 7209 793
rect 7168 763 7172 767
rect 7179 763 7187 772
rect 7191 763 7193 792
rect 7344 788 7346 796
rect 7352 794 7374 803
rect 7352 792 7367 794
rect 7404 792 7417 806
rect 7442 804 7444 807
rect 7448 806 7462 807
rect 7446 803 7462 806
rect 7498 805 7514 808
rect 7496 803 7514 805
rect 7404 790 7412 792
rect 7434 791 7442 803
rect 7444 801 7480 803
rect 7444 793 7464 801
rect 7477 800 7480 801
rect 7478 793 7480 800
rect 7484 799 7492 803
rect 7496 799 7518 803
rect 7498 794 7518 799
rect 7556 798 7564 810
rect 7568 800 7570 830
rect 7587 826 7589 840
rect 7629 838 7635 844
rect 7687 838 7693 844
rect 7726 841 7731 845
rect 8019 841 8024 845
rect 8018 832 8026 841
rect 8030 834 8032 839
rect 8062 834 8064 846
rect 8322 845 8324 865
rect 8356 863 8358 872
rect 8393 863 8394 872
rect 8512 868 8529 881
rect 8557 868 8562 872
rect 8512 866 8521 868
rect 8512 865 8520 866
rect 8546 865 8554 866
rect 8355 857 8356 862
rect 8353 849 8354 855
rect 8074 844 8082 845
rect 8030 832 8064 834
rect 8068 832 8082 844
rect 7602 826 7603 832
rect 8074 830 8082 832
rect 7713 829 7716 830
rect 7689 827 7724 829
rect 7587 818 7588 826
rect 7685 825 7689 827
rect 7588 800 7591 814
rect 7603 812 7605 825
rect 7656 808 7685 825
rect 7687 814 7689 817
rect 7697 812 7713 827
rect 7692 811 7713 812
rect 7724 824 7884 827
rect 7568 798 7602 800
rect 7588 795 7591 798
rect 7346 778 7349 788
rect 7349 769 7351 778
rect 7352 774 7367 790
rect 7404 774 7418 790
rect 7441 781 7442 788
rect 7351 765 7352 769
rect 7168 762 7193 763
rect 7222 762 7225 763
rect 7168 760 7225 762
rect 7168 758 7184 760
rect 7352 759 7353 763
rect 5293 749 5329 750
rect 5312 744 5324 749
rect 5379 744 5390 749
rect 6846 746 6849 754
rect 6877 748 6882 754
rect 6882 745 6886 748
rect 7076 745 7078 757
rect 7081 745 7115 757
rect 7120 756 7122 757
rect 7229 756 7256 759
rect 7353 757 7354 759
rect 7368 758 7384 772
rect 7386 758 7402 772
rect 7434 769 7442 781
rect 7446 774 7464 793
rect 7498 792 7514 794
rect 7498 774 7514 790
rect 7544 774 7559 790
rect 7561 775 7563 789
rect 7568 786 7580 794
rect 7590 786 7602 794
rect 7604 790 7605 808
rect 7691 805 7701 811
rect 7724 808 7890 824
rect 7952 808 7968 824
rect 7970 808 7986 824
rect 8030 820 8042 828
rect 8052 820 8064 828
rect 8030 810 8032 820
rect 8082 816 8086 830
rect 8108 828 8110 845
rect 8110 819 8111 828
rect 8138 819 8141 845
rect 8143 843 8192 845
rect 8227 843 8229 844
rect 8143 833 8185 843
rect 8263 838 8264 843
rect 8230 827 8231 836
rect 8264 827 8265 836
rect 8321 834 8322 844
rect 8352 843 8353 847
rect 8351 837 8352 843
rect 8180 811 8185 823
rect 8232 817 8233 820
rect 8265 816 8266 820
rect 8320 819 8321 832
rect 8349 827 8351 836
rect 8391 829 8393 862
rect 8504 855 8520 865
rect 8557 864 8561 868
rect 8441 845 8504 855
rect 8549 851 8557 864
rect 8432 844 8441 845
rect 8426 842 8432 844
rect 8416 834 8426 842
rect 8348 821 8349 826
rect 8389 820 8391 827
rect 8233 811 8234 814
rect 8266 811 8267 814
rect 8319 811 8320 818
rect 8333 811 8339 817
rect 8347 816 8348 820
rect 8388 818 8389 820
rect 8396 818 8416 834
rect 8346 814 8347 816
rect 8345 812 8346 814
rect 8379 811 8385 817
rect 8387 813 8396 818
rect 8386 811 8396 813
rect 8142 808 8143 810
rect 8234 808 8235 810
rect 7696 803 7701 805
rect 7821 803 7830 808
rect 7868 803 7877 808
rect 7608 802 7617 803
rect 7606 798 7614 802
rect 7617 799 7632 802
rect 7632 798 7635 799
rect 7629 792 7635 798
rect 7687 792 7693 798
rect 7701 794 7710 803
rect 7812 794 7821 803
rect 7877 794 7886 803
rect 7803 792 7810 793
rect 7635 790 7641 792
rect 7446 772 7480 774
rect 7493 772 7498 774
rect 7591 772 7594 786
rect 7604 774 7610 790
rect 7635 786 7656 790
rect 7681 786 7687 792
rect 7797 791 7803 792
rect 7854 791 7858 793
rect 7890 792 7906 808
rect 7936 792 7952 808
rect 7963 803 7969 808
rect 7963 802 7978 803
rect 7957 796 7963 802
rect 7986 798 8002 808
rect 8009 802 8015 808
rect 7962 791 7963 793
rect 7995 791 8000 798
rect 8015 796 8021 802
rect 8033 800 8034 808
rect 7795 790 7797 791
rect 7794 787 7795 790
rect 7859 789 7861 790
rect 7640 774 7656 786
rect 7707 778 7734 781
rect 7690 774 7707 778
rect 7734 774 7742 778
rect 7446 769 7498 772
rect 7559 769 7565 772
rect 7594 771 7598 772
rect 7446 757 7450 765
rect 7482 758 7498 769
rect 7560 762 7577 769
rect 7594 762 7604 771
rect 7560 758 7576 762
rect 7577 760 7582 762
rect 7586 760 7598 762
rect 7582 759 7598 760
rect 7578 758 7598 759
rect 7656 758 7672 774
rect 7742 772 7745 774
rect 7810 772 7816 778
rect 7819 772 7821 779
rect 7861 772 7862 778
rect 7890 774 7906 790
rect 7936 774 7952 790
rect 7954 779 7963 791
rect 7889 772 7890 774
rect 7745 763 7765 772
rect 7794 767 7795 769
rect 7804 766 7810 772
rect 7862 766 7868 772
rect 7883 763 7890 772
rect 7765 762 7767 763
rect 7767 759 7773 762
rect 7122 751 7143 756
rect 7143 747 7159 751
rect 7191 748 7203 756
rect 7354 754 7355 756
rect 7250 747 7256 753
rect 7281 747 7336 753
rect 7355 750 7356 754
rect 7356 747 7358 748
rect 7365 747 7374 756
rect 7444 747 7450 756
rect 7502 747 7508 753
rect 7509 747 7518 756
rect 7563 751 7566 758
rect 5390 743 5392 744
rect 4876 739 4885 742
rect 4962 741 4964 742
rect 5264 741 5265 743
rect 6849 741 6851 745
rect 4707 738 4721 739
rect 4694 737 4707 738
rect 4714 735 4716 738
rect 4885 735 4896 739
rect 4939 737 4940 739
rect 4896 734 4899 735
rect 4505 733 4587 734
rect 4455 732 4521 733
rect 4498 731 4521 732
rect 4244 726 4256 731
rect 4498 729 4505 731
rect 4509 730 4521 731
rect 4587 729 4590 732
rect 4706 731 4713 734
rect 4899 731 4908 734
rect 4936 733 4938 736
rect 4908 729 4915 731
rect 4931 729 4935 731
rect 4494 728 4498 729
rect 4487 726 4494 728
rect 4524 727 4525 729
rect 4590 728 4592 729
rect 3946 721 4017 723
rect 3770 719 3785 720
rect 3947 719 4017 721
rect 4049 719 4053 725
rect 4160 723 4162 726
rect 3773 716 3785 719
rect 3709 712 3714 716
rect 3786 714 3789 716
rect 3938 712 3946 719
rect 3948 717 3958 719
rect 3982 717 4037 719
rect 3948 712 3952 717
rect 3714 696 3735 712
rect 3779 710 3803 712
rect 3783 705 3803 710
rect 3938 707 3948 712
rect 3945 705 3948 707
rect 3735 695 3737 696
rect 3741 689 3742 692
rect 3739 678 3746 687
rect 3783 680 3785 705
rect 3789 700 3797 705
rect 3803 699 3809 705
rect 3943 701 3945 705
rect 3937 699 3945 701
rect 3809 694 3815 699
rect 3937 695 3943 699
rect 3815 692 3818 694
rect 3751 678 3785 680
rect 3789 678 3797 690
rect 3818 688 3819 692
rect 3931 689 3937 695
rect 3941 692 3942 694
rect 3940 688 3941 691
rect 3950 689 3952 712
rect 3982 712 3992 717
rect 3998 715 4037 717
rect 4013 713 4037 715
rect 4057 713 4058 715
rect 3982 701 3984 712
rect 3992 701 4005 712
rect 4018 708 4037 713
rect 4058 708 4062 713
rect 4162 710 4169 723
rect 4256 722 4286 726
rect 4505 724 4521 726
rect 4256 714 4298 722
rect 4025 701 4037 708
rect 4062 706 4063 708
rect 4169 705 4172 710
rect 4250 709 4299 710
rect 3982 695 3989 701
rect 3982 693 3995 695
rect 3982 689 3984 693
rect 3989 689 3995 693
rect 4000 691 4009 700
rect 4028 696 4037 701
rect 4068 696 4071 701
rect 4031 691 4037 696
rect 3939 685 3940 687
rect 3983 685 3984 689
rect 4001 687 4018 691
rect 4034 689 4037 691
rect 4071 689 4077 696
rect 4172 695 4209 705
rect 4250 702 4264 709
rect 4280 708 4299 709
rect 4296 703 4299 708
rect 4249 699 4250 701
rect 4209 693 4215 695
rect 4247 694 4249 699
rect 4215 692 4220 693
rect 4246 692 4247 694
rect 4036 687 4037 689
rect 4002 686 4018 687
rect 4077 686 4079 689
rect 4220 688 4236 692
rect 4236 687 4238 688
rect 3819 680 3821 685
rect 3938 680 3939 685
rect 4004 682 4007 686
rect 4009 682 4018 686
rect 4010 680 4011 682
rect 3746 676 3747 678
rect 3750 676 3751 678
rect 3937 676 3938 678
rect 4011 677 4012 678
rect 3746 660 3750 676
rect 3786 674 3789 676
rect 3751 666 3763 674
rect 3773 666 3785 674
rect 3821 660 3825 676
rect 3745 654 3746 658
rect 3825 657 3826 660
rect 3745 630 3747 654
rect 3825 630 3826 654
rect 3937 649 3989 663
rect 4010 662 4012 675
rect 4039 672 4051 685
rect 4079 672 4091 686
rect 4241 685 4247 687
rect 4247 683 4255 685
rect 4252 681 4256 683
rect 4252 676 4259 681
rect 4296 678 4298 703
rect 4299 697 4300 702
rect 4302 698 4310 710
rect 4455 694 4483 695
rect 4519 694 4521 724
rect 4525 714 4533 726
rect 4592 712 4594 728
rect 4915 727 4921 729
rect 4928 727 4931 729
rect 4648 720 4654 726
rect 4706 720 4712 726
rect 4912 723 4932 727
rect 4964 723 4985 741
rect 4990 738 5001 740
rect 4912 721 4928 723
rect 4907 720 4912 721
rect 4932 720 4940 723
rect 4654 714 4660 720
rect 4700 714 4706 720
rect 4900 717 4907 720
rect 4940 719 4943 720
rect 4985 719 4990 723
rect 4895 716 4900 717
rect 4943 716 4949 719
rect 4990 716 4994 719
rect 4998 716 5000 738
rect 5001 737 5002 738
rect 5004 737 5012 740
rect 5002 734 5012 737
rect 5004 728 5012 734
rect 5091 733 5092 741
rect 5128 737 5131 741
rect 5092 729 5093 733
rect 5121 729 5133 737
rect 5143 729 5155 737
rect 5218 729 5231 741
rect 5010 726 5013 728
rect 5013 719 5020 726
rect 5093 724 5100 729
rect 5117 727 5120 729
rect 5133 725 5134 729
rect 5140 725 5146 729
rect 5094 723 5100 724
rect 5109 723 5117 725
rect 5121 723 5167 725
rect 5004 716 5012 718
rect 4886 713 4895 716
rect 4881 711 4886 713
rect 4300 693 4301 694
rect 4475 692 4483 694
rect 4487 692 4521 694
rect 4525 692 4533 704
rect 4592 694 4594 710
rect 4865 706 4881 711
rect 4949 706 4960 716
rect 4994 707 5012 716
rect 5020 712 5028 719
rect 5088 717 5094 723
rect 5121 717 5123 723
rect 5146 717 5152 723
rect 5153 719 5167 723
rect 5092 713 5094 714
rect 4976 706 5012 707
rect 5028 706 5036 712
rect 5090 709 5092 713
rect 4849 701 4865 706
rect 4960 705 4967 706
rect 5005 705 5038 706
rect 4960 702 4968 705
rect 4942 701 4976 702
rect 5002 701 5063 705
rect 5153 702 5155 719
rect 5159 713 5167 719
rect 5162 712 5167 713
rect 5231 712 5250 729
rect 5265 715 5299 741
rect 5394 723 5417 741
rect 6886 740 6894 745
rect 7112 742 7113 745
rect 7159 742 7179 747
rect 7179 741 7184 742
rect 7256 741 7262 747
rect 7302 741 7308 747
rect 7078 740 7080 741
rect 6851 737 6853 740
rect 6894 737 6899 740
rect 7068 739 7078 740
rect 7057 738 7078 739
rect 7184 738 7188 741
rect 7309 738 7318 747
rect 7356 745 7365 747
rect 7356 742 7371 745
rect 7356 738 7365 742
rect 7371 740 7375 742
rect 7450 741 7462 747
rect 7496 741 7509 747
rect 7565 744 7566 751
rect 7375 739 7378 740
rect 6899 736 6901 737
rect 7066 736 7085 738
rect 6854 733 6855 736
rect 6901 733 6905 736
rect 6855 727 6858 733
rect 6905 731 6909 733
rect 6909 729 6912 731
rect 6999 729 7005 735
rect 7057 729 7063 735
rect 7066 733 7103 736
rect 7110 733 7111 736
rect 7077 729 7103 733
rect 7106 729 7110 731
rect 7142 729 7143 730
rect 6912 726 6916 729
rect 6858 720 6862 726
rect 6916 720 6926 726
rect 6929 720 6941 724
rect 7005 723 7011 729
rect 7051 723 7057 729
rect 7103 726 7143 729
rect 7103 723 7142 726
rect 7188 725 7205 738
rect 7309 737 7310 738
rect 7378 736 7385 739
rect 7453 738 7462 741
rect 7500 738 7509 741
rect 7559 739 7566 744
rect 7594 742 7598 758
rect 7636 747 7645 756
rect 7701 747 7710 756
rect 7773 754 7784 759
rect 7877 758 7890 763
rect 7952 772 7953 774
rect 7952 769 7961 772
rect 7962 769 7963 779
rect 7952 763 7963 769
rect 7966 763 7968 791
rect 8034 790 8036 791
rect 8032 785 8036 790
rect 8085 790 8086 808
rect 8192 799 8204 804
rect 8236 796 8237 799
rect 8267 796 8268 805
rect 8318 799 8319 808
rect 8327 805 8333 811
rect 8385 808 8391 811
rect 8440 808 8456 824
rect 9029 819 9030 1015
rect 9219 819 9220 1015
rect 9305 819 9306 1015
rect 9578 819 9579 1015
rect 9775 819 9776 1015
rect 10166 1014 10170 1019
rect 10804 1014 10811 1019
rect 10891 1018 10900 1027
rect 10956 1024 11052 1027
rect 11393 1023 11501 1037
rect 11251 1015 11267 1022
rect 11269 1015 11285 1022
rect 10811 1007 10823 1014
rect 11241 1013 11253 1015
rect 11263 1013 11275 1015
rect 11281 1013 11285 1015
rect 11469 1013 11485 1022
rect 11501 1021 11519 1023
rect 11520 1017 11527 1020
rect 11527 1013 11533 1017
rect 12173 1015 12174 1026
rect 12363 1015 12364 1026
rect 12449 1015 12450 1026
rect 12722 1015 12723 1026
rect 12919 1015 12920 1026
rect 13348 1023 13449 1034
rect 13635 1033 13899 1034
rect 13899 1023 13954 1033
rect 14057 1027 14066 1036
rect 14104 1027 14113 1036
rect 14407 1034 14529 1037
rect 14379 1033 14396 1034
rect 14209 1027 14379 1033
rect 13333 1021 13348 1023
rect 13327 1019 13333 1021
rect 13956 1019 13961 1021
rect 11241 1008 11285 1013
rect 11428 1008 11465 1009
rect 11533 1008 11536 1013
rect 11237 1006 11239 1008
rect 11241 1006 11373 1008
rect 10292 1005 10646 1006
rect 10272 1003 10290 1005
rect 10732 1003 10745 1005
rect 10824 1003 10827 1005
rect 11235 1003 11373 1006
rect 10216 1000 10272 1003
rect 10090 992 10102 1000
rect 10112 992 10124 1000
rect 10188 994 10272 1000
rect 10745 994 10755 1003
rect 10188 993 10216 994
rect 10086 989 10088 992
rect 10188 991 10207 993
rect 10756 991 10759 993
rect 10128 988 10132 989
rect 10078 977 10086 988
rect 10089 986 10124 988
rect 10087 977 10089 983
rect 10078 976 10087 977
rect 10086 972 10087 976
rect 10085 971 10086 972
rect 10083 966 10085 969
rect 9958 964 10023 965
rect 9950 956 9958 964
rect 10023 956 10027 964
rect 9949 950 9950 956
rect 10078 954 10086 966
rect 10090 956 10092 986
rect 10121 985 10124 986
rect 10123 979 10124 985
rect 10128 981 10136 988
rect 10132 980 10140 981
rect 10164 980 10165 990
rect 10188 980 10203 991
rect 10462 981 10499 983
rect 10140 979 10146 980
rect 10163 979 10164 980
rect 10188 979 10195 980
rect 10146 969 10208 979
rect 10216 972 10222 978
rect 10262 972 10268 978
rect 10462 977 10488 981
rect 10499 977 10504 981
rect 10759 980 10772 991
rect 10735 979 10749 980
rect 10456 972 10462 977
rect 10504 972 10513 977
rect 10717 972 10735 979
rect 10749 977 10756 979
rect 10827 977 10848 1003
rect 11229 996 11373 1003
rect 11389 1006 11490 1008
rect 11389 996 11501 1006
rect 11190 990 11251 996
rect 11155 987 11190 990
rect 10968 981 11155 987
rect 11241 986 11251 990
rect 10756 972 10771 977
rect 10210 969 10216 972
rect 10217 970 10274 972
rect 10513 971 10514 972
rect 10351 970 10354 971
rect 10372 970 10375 971
rect 10454 970 10455 971
rect 10514 970 10517 971
rect 10217 969 10225 970
rect 10188 968 10225 969
rect 10090 954 10124 956
rect 10079 951 10081 954
rect 10075 938 10079 950
rect 10090 942 10102 950
rect 10115 945 10124 954
rect 10162 952 10163 955
rect 10188 951 10193 968
rect 10210 966 10225 968
rect 10268 966 10274 970
rect 10350 969 10351 970
rect 10375 969 10376 970
rect 10709 969 10717 972
rect 10746 971 10771 972
rect 10780 971 10784 972
rect 10742 970 10746 971
rect 10756 970 10793 971
rect 10741 969 10742 970
rect 10347 967 10350 969
rect 10376 967 10380 969
rect 10517 968 10518 969
rect 10518 967 10521 968
rect 10216 964 10225 966
rect 10343 965 10347 967
rect 10380 965 10384 967
rect 10701 966 10709 969
rect 10739 968 10741 969
rect 10735 967 10739 968
rect 10730 965 10735 967
rect 10756 965 10771 970
rect 10780 969 10784 970
rect 10793 969 10794 970
rect 10850 969 10855 975
rect 10891 971 10900 980
rect 10956 978 10968 981
rect 10956 971 10965 978
rect 11235 972 11251 986
rect 11274 972 11275 996
rect 11280 991 11301 996
rect 11285 990 11301 991
rect 11418 989 11424 996
rect 11470 989 11476 996
rect 11490 990 11501 996
rect 11536 990 11545 1008
rect 11285 972 11301 988
rect 11418 985 11426 989
rect 11424 983 11426 985
rect 11355 977 11362 978
rect 11364 977 11366 978
rect 11334 974 11355 977
rect 11366 974 11375 977
rect 11332 972 11334 974
rect 11375 972 11377 974
rect 10784 965 10789 969
rect 10794 965 10796 968
rect 10855 965 10858 969
rect 10341 964 10343 965
rect 10384 964 10386 965
rect 10696 964 10700 965
rect 10771 964 10774 965
rect 10796 964 10797 965
rect 10216 951 10221 964
rect 10269 955 10288 958
rect 10327 956 10341 964
rect 10386 959 10398 964
rect 10453 959 10454 964
rect 10398 956 10401 959
rect 10521 957 10524 964
rect 10692 962 10696 964
rect 10323 955 10327 956
rect 10125 949 10130 950
rect 10130 948 10135 949
rect 10135 947 10138 948
rect 10140 945 10149 947
rect 10113 942 10115 945
rect 10149 944 10154 945
rect 10154 943 10160 944
rect 10161 943 10162 951
rect 10188 943 10194 951
rect 10112 939 10113 942
rect 10160 938 10194 943
rect 10073 931 10075 937
rect 10110 930 10112 938
rect 10161 932 10162 938
rect 10188 935 10216 938
rect 10188 933 10218 935
rect 10188 931 10219 933
rect 10220 931 10221 951
rect 10288 946 10350 955
rect 10401 952 10406 956
rect 10452 951 10453 956
rect 10524 954 10525 956
rect 10661 950 10692 962
rect 10776 959 10780 962
rect 10791 960 10795 963
rect 10900 962 10909 971
rect 10933 961 10936 963
rect 10947 962 10956 971
rect 11241 970 11275 972
rect 11284 971 11285 972
rect 11331 971 11332 972
rect 11280 970 11285 971
rect 11330 970 11331 971
rect 11241 968 11285 970
rect 11328 969 11330 970
rect 11377 969 11380 972
rect 11237 965 11238 967
rect 11011 961 11020 963
rect 10928 959 10933 961
rect 10306 945 10316 946
rect 10338 945 10339 946
rect 10302 943 10306 945
rect 10350 943 10370 946
rect 10451 943 10452 950
rect 10524 943 10525 950
rect 10659 949 10661 950
rect 10573 943 10579 949
rect 10619 948 10625 949
rect 10656 948 10659 949
rect 10619 947 10656 948
rect 10619 943 10625 947
rect 10711 946 10717 952
rect 10757 946 10763 952
rect 10779 950 10780 959
rect 10926 958 10928 959
rect 11022 958 11028 961
rect 10797 955 10801 958
rect 10865 955 10867 958
rect 11028 956 11031 958
rect 11251 956 11267 968
rect 11269 956 11285 968
rect 11324 965 11328 968
rect 11380 965 11384 969
rect 11424 967 11427 983
rect 11323 964 11324 965
rect 11384 964 11385 965
rect 11322 963 11323 964
rect 11320 961 11322 963
rect 11385 961 11388 964
rect 11426 961 11427 967
rect 11430 967 11431 989
rect 11469 985 11476 989
rect 11497 987 11499 990
rect 11469 983 11470 985
rect 11490 984 11491 986
rect 11430 963 11432 967
rect 11463 963 11464 966
rect 11468 965 11470 983
rect 11499 981 11502 987
rect 11502 979 11503 981
rect 11504 975 11505 977
rect 11505 972 11506 975
rect 11545 973 11553 990
rect 11507 965 11510 969
rect 11430 961 11434 963
rect 11468 962 11469 965
rect 11510 963 11511 965
rect 11316 958 11319 961
rect 11388 959 11391 961
rect 11315 956 11316 958
rect 11391 957 11393 959
rect 10801 946 10811 955
rect 10290 931 10298 943
rect 10302 941 10336 943
rect 10026 924 10027 929
rect 9976 915 9985 924
rect 10023 920 10032 924
rect 10023 915 10037 920
rect 9967 912 9976 915
rect 9967 911 9970 912
rect 9960 908 9969 911
rect 9948 907 9969 908
rect 9948 905 9966 907
rect 10006 905 10012 911
rect 10026 906 10041 915
rect 10066 908 10073 929
rect 9948 900 9960 905
rect 9944 898 9947 900
rect 9948 899 9949 900
rect 9954 899 9960 900
rect 10012 899 10018 905
rect 10025 904 10037 906
rect 10064 904 10066 908
rect 10104 907 10110 929
rect 10161 926 10162 929
rect 10188 928 10249 931
rect 10188 917 10194 928
rect 10216 926 10249 928
rect 10210 925 10249 926
rect 10268 925 10274 926
rect 10210 921 10274 925
rect 10210 920 10296 921
rect 10188 913 10197 917
rect 10216 914 10222 920
rect 10262 914 10268 920
rect 10271 917 10296 920
rect 10280 913 10296 917
rect 10302 913 10304 941
rect 10333 939 10336 941
rect 10188 909 10203 913
rect 10290 909 10304 913
rect 10334 909 10336 939
rect 10340 931 10348 943
rect 10370 934 10433 943
rect 10567 938 10573 943
rect 10585 941 10621 943
rect 10585 938 10590 941
rect 10526 937 10573 938
rect 10587 937 10590 938
rect 10625 937 10631 943
rect 10705 940 10711 946
rect 10763 940 10769 946
rect 10526 936 10569 937
rect 10450 934 10451 936
rect 10472 934 10526 936
rect 10406 922 10421 934
rect 10433 933 10472 934
rect 10450 929 10451 933
rect 10582 929 10585 936
rect 10709 933 10711 934
rect 10707 929 10709 933
rect 10103 904 10104 906
rect 10163 905 10164 909
rect 10023 899 10025 904
rect 10169 903 10175 909
rect 10188 903 10207 909
rect 10215 903 10221 909
rect 10063 899 10064 903
rect 10022 897 10023 899
rect 10062 897 10063 899
rect 9936 884 9944 896
rect 9948 894 9966 896
rect 10021 895 10022 896
rect 10101 895 10103 903
rect 10163 897 10169 903
rect 10188 897 10227 903
rect 10229 897 10241 905
rect 10302 904 10319 909
rect 10310 899 10317 904
rect 10319 903 10323 904
rect 10339 903 10340 905
rect 10406 904 10421 920
rect 10448 906 10450 928
rect 10323 900 10342 903
rect 10447 900 10459 905
rect 10469 900 10481 905
rect 10522 904 10524 928
rect 10573 904 10582 928
rect 10618 904 10621 909
rect 10659 908 10694 910
rect 10705 908 10707 929
rect 10729 909 10730 929
rect 10777 928 10779 944
rect 10811 942 10816 946
rect 10867 942 10879 955
rect 11031 951 11041 956
rect 11314 953 11315 956
rect 11149 952 11186 953
rect 11313 952 11314 953
rect 11393 952 11395 956
rect 11421 955 11427 961
rect 11434 959 11440 961
rect 11441 957 11447 959
rect 11447 956 11450 957
rect 11467 956 11473 961
rect 11511 960 11512 963
rect 11512 958 11513 960
rect 11149 951 11174 952
rect 11186 951 11187 952
rect 11312 951 11313 952
rect 11043 948 11047 951
rect 11114 948 11141 951
rect 11189 948 11196 951
rect 11196 943 11207 948
rect 11242 945 11244 949
rect 11277 947 11278 949
rect 11310 948 11312 951
rect 11207 942 11211 943
rect 10879 939 10880 942
rect 11211 938 11218 942
rect 10821 929 10831 938
rect 10881 931 10887 938
rect 11218 937 11220 938
rect 11220 933 11236 937
rect 11236 932 11241 933
rect 11244 932 11252 944
rect 11241 929 11252 932
rect 11278 929 11282 944
rect 11308 943 11310 948
rect 11395 944 11398 951
rect 11415 949 11421 955
rect 11450 951 11491 956
rect 11513 955 11515 958
rect 11473 949 11479 951
rect 11515 948 11518 955
rect 11307 942 11308 943
rect 11518 942 11521 948
rect 11553 943 11554 973
rect 11661 951 11677 954
rect 11589 943 11612 951
rect 11667 943 11684 951
rect 11306 940 11307 942
rect 11305 939 11306 940
rect 11521 939 11522 942
rect 11304 937 11305 938
rect 11301 933 11304 937
rect 11299 932 11301 933
rect 11297 929 11299 932
rect 11522 931 11523 938
rect 11552 929 11553 942
rect 11581 938 11589 943
rect 11667 938 11691 943
rect 11571 932 11581 938
rect 11564 929 11571 932
rect 10774 917 10776 920
rect 10770 914 10773 916
rect 10768 913 10770 914
rect 10765 911 10768 913
rect 10763 910 10765 911
rect 10649 906 10659 908
rect 10694 906 10711 908
rect 10638 904 10649 906
rect 10572 900 10573 903
rect 10616 900 10618 904
rect 10630 902 10638 904
rect 10626 901 10630 902
rect 10705 900 10707 906
rect 10729 904 10730 906
rect 10797 904 10813 920
rect 10831 910 10853 929
rect 10891 920 10899 927
rect 10899 918 10906 920
rect 10906 914 10922 918
rect 10925 914 10926 929
rect 11244 928 11257 929
rect 11250 927 11257 928
rect 11282 927 11283 928
rect 11296 927 11297 929
rect 11420 927 11421 929
rect 11252 923 11253 926
rect 11257 924 11294 927
rect 10984 921 11015 922
rect 10975 920 10984 921
rect 11015 920 11022 921
rect 11282 920 11283 924
rect 10946 917 10975 920
rect 11022 917 11037 920
rect 10944 916 10946 917
rect 10937 914 10944 916
rect 11037 914 11049 917
rect 11254 915 11255 917
rect 11283 915 11284 920
rect 11288 915 11297 924
rect 11335 915 11344 924
rect 11419 922 11420 927
rect 11418 920 11419 922
rect 11417 918 11418 920
rect 11416 916 11417 918
rect 11279 914 11288 915
rect 10922 911 11288 914
rect 10925 910 10926 911
rect 10928 910 10930 911
rect 11064 910 11072 911
rect 10853 909 10855 910
rect 10730 900 10734 904
rect 10784 900 10797 904
rect 10855 903 10863 909
rect 10924 908 10928 910
rect 11072 906 11090 910
rect 11255 906 11256 909
rect 11285 906 11286 909
rect 10917 904 10922 906
rect 10188 895 10243 897
rect 10317 895 10323 899
rect 10337 898 10338 900
rect 10336 895 10337 897
rect 10342 896 10511 900
rect 10570 897 10572 900
rect 10567 896 10573 897
rect 10613 896 10616 900
rect 10447 895 10448 896
rect 10511 895 10573 896
rect 9936 862 9944 874
rect 9948 865 9950 894
rect 10020 893 10021 894
rect 10061 893 10062 894
rect 10188 893 10245 895
rect 10323 893 10324 895
rect 10015 889 10021 893
rect 10060 889 10061 893
rect 10100 889 10101 893
rect 10156 889 10163 893
rect 10188 892 10253 893
rect 10001 888 10021 889
rect 10001 878 10015 888
rect 10057 879 10060 889
rect 10098 878 10100 889
rect 10153 879 10156 889
rect 9985 866 10001 878
rect 9948 862 9951 865
rect 9982 862 9985 866
rect 10032 859 10041 868
rect 10053 866 10057 878
rect 10097 875 10098 878
rect 10152 875 10153 878
rect 10052 862 10053 866
rect 9947 857 9949 858
rect 9954 857 9960 859
rect 9948 853 9960 857
rect 10012 853 10018 859
rect 10024 857 10032 859
rect 10051 858 10052 862
rect 10093 859 10097 875
rect 10147 859 10152 875
rect 10165 864 10168 892
rect 10215 891 10241 892
rect 10239 861 10241 891
rect 10245 881 10253 892
rect 10324 879 10344 893
rect 10392 879 10406 894
rect 10435 881 10443 893
rect 10447 891 10481 893
rect 10300 876 10301 879
rect 10330 876 10331 879
rect 10344 877 10356 879
rect 10390 877 10392 879
rect 10344 875 10390 877
rect 10215 859 10241 861
rect 10245 859 10253 871
rect 10298 869 10300 875
rect 10328 870 10330 875
rect 10296 862 10298 869
rect 10325 862 10328 869
rect 10295 859 10296 862
rect 10324 859 10325 862
rect 10447 859 10449 891
rect 10479 875 10481 891
rect 10485 881 10493 893
rect 10567 891 10573 895
rect 10611 891 10613 895
rect 10625 891 10631 897
rect 10705 894 10711 900
rect 10734 896 10749 900
rect 10749 895 10750 896
rect 10763 895 10797 900
rect 10863 899 10869 903
rect 10914 902 10917 904
rect 11090 902 11110 906
rect 11181 902 11194 903
rect 10521 881 10522 889
rect 10565 881 10568 891
rect 10573 885 10579 891
rect 10605 881 10611 891
rect 10619 885 10625 891
rect 10708 883 10709 891
rect 10711 888 10717 894
rect 10750 893 10769 895
rect 10480 865 10481 874
rect 10485 872 10486 875
rect 10515 870 10521 880
rect 10560 870 10565 881
rect 10503 866 10515 870
rect 10559 867 10560 870
rect 10598 867 10605 881
rect 10748 872 10751 892
rect 10757 888 10763 893
rect 10781 888 10797 895
rect 10869 894 10880 899
rect 10908 898 10912 900
rect 10905 897 10908 898
rect 10902 895 10905 897
rect 10925 895 10928 900
rect 11110 897 11135 902
rect 11160 900 11178 902
rect 11199 900 11222 902
rect 11158 899 11170 900
rect 11222 899 11231 900
rect 11231 898 11232 899
rect 11256 898 11257 902
rect 11135 895 11140 897
rect 11151 895 11158 898
rect 10880 885 10911 894
rect 10928 893 10930 895
rect 10930 891 10932 893
rect 11140 891 11158 895
rect 11232 894 11239 898
rect 11286 897 11287 902
rect 11344 901 11353 915
rect 11414 911 11415 914
rect 11441 909 11473 913
rect 11408 903 11412 906
rect 11415 903 11421 909
rect 11441 904 11479 909
rect 11510 904 11564 929
rect 11667 922 11693 938
rect 11438 903 11479 904
rect 11395 901 11407 902
rect 11353 899 11357 901
rect 11375 900 11395 901
rect 11369 899 11375 900
rect 11395 895 11397 900
rect 11421 897 11427 903
rect 11455 899 11456 901
rect 11239 891 11245 894
rect 11257 891 11258 895
rect 10870 880 10911 885
rect 10932 888 11005 891
rect 11140 889 11157 891
rect 10932 885 11012 888
rect 10932 881 11005 885
rect 11012 881 11082 885
rect 11143 882 11151 889
rect 11157 887 11162 889
rect 11162 885 11166 887
rect 11245 885 11258 891
rect 11287 887 11289 895
rect 11393 892 11395 895
rect 11392 891 11393 892
rect 10870 876 10886 880
rect 10911 876 10929 880
rect 10932 876 10950 881
rect 11005 876 11110 881
rect 10929 875 11110 876
rect 11136 875 11143 882
rect 11166 876 11188 885
rect 11245 882 11259 885
rect 11258 881 11261 882
rect 11258 878 11259 881
rect 11261 880 11262 881
rect 11262 879 11271 880
rect 11289 879 11291 885
rect 11380 882 11392 891
rect 11374 881 11380 882
rect 11346 880 11362 881
rect 11370 880 11374 881
rect 11439 880 11454 899
rect 11467 897 11473 903
rect 11504 901 11510 904
rect 11518 903 11519 904
rect 11493 895 11504 901
rect 11517 899 11518 901
rect 11490 892 11493 895
rect 11489 891 11490 892
rect 11481 885 11489 891
rect 11318 879 11341 880
rect 11188 875 11191 876
rect 10597 866 10598 867
rect 10502 865 10503 866
rect 10480 862 10502 865
rect 10556 862 10559 866
rect 10481 859 10502 862
rect 10553 859 10559 862
rect 10023 855 10032 857
rect 9948 852 9957 853
rect 9948 850 9958 852
rect 9960 850 9966 853
rect 9958 847 9966 850
rect 9958 842 9962 847
rect 10011 840 10012 853
rect 10021 852 10032 855
rect 10019 851 10021 852
rect 10016 850 10019 851
rect 10023 850 10032 852
rect 10047 845 10051 858
rect 10090 846 10093 858
rect 10143 846 10147 858
rect 10163 851 10169 857
rect 10192 856 10196 859
rect 10486 858 10487 859
rect 10169 845 10175 851
rect 10187 845 10192 856
rect 10221 851 10227 857
rect 10294 855 10295 858
rect 10323 855 10324 858
rect 10553 857 10556 859
rect 10555 856 10556 857
rect 10551 855 10555 856
rect 10215 845 10221 851
rect 10229 847 10241 855
rect 10445 853 10446 855
rect 10043 841 10047 845
rect 10089 841 10090 845
rect 10141 842 10143 845
rect 10041 840 10043 841
rect 10185 840 10187 845
rect 10289 841 10292 850
rect 10319 841 10322 850
rect 10446 841 10448 849
rect 10487 842 10488 849
rect 10548 847 10555 855
rect 10542 845 10549 847
rect 10551 845 10555 847
rect 10585 845 10597 865
rect 10709 859 10711 872
rect 10542 840 10551 845
rect 10582 844 10589 845
rect 10744 844 10748 870
rect 10859 869 10869 875
rect 10922 872 11122 875
rect 11133 872 11136 875
rect 11191 872 11201 875
rect 11207 872 11219 878
rect 11262 875 11341 879
rect 11469 876 11501 885
rect 11514 880 11517 898
rect 11513 876 11514 880
rect 11549 878 11551 904
rect 11667 895 11690 922
rect 11722 895 11723 929
rect 11667 881 11689 895
rect 11701 889 11723 895
rect 10922 871 10930 872
rect 10917 869 10921 871
rect 10857 868 10859 869
rect 10854 866 10857 868
rect 10912 866 10916 868
rect 11005 867 11229 872
rect 11259 871 11260 875
rect 11271 871 11318 875
rect 11432 872 11435 876
rect 11466 875 11501 876
rect 11277 869 11318 871
rect 11283 868 11308 869
rect 11021 866 11229 867
rect 10847 862 10854 866
rect 10902 862 10912 866
rect 11021 863 11231 866
rect 11134 862 11143 863
rect 11217 862 11239 863
rect 11260 862 11261 868
rect 11284 867 11308 868
rect 11424 863 11432 872
rect 11479 869 11480 874
rect 10841 858 10847 862
rect 11143 858 11150 862
rect 10839 857 10841 858
rect 10830 852 10839 857
rect 11150 852 11161 858
rect 11217 854 11231 862
rect 11239 856 11272 862
rect 11291 859 11292 862
rect 11420 857 11424 862
rect 11347 856 11359 857
rect 11272 855 11278 856
rect 11296 855 11318 856
rect 11278 854 11318 855
rect 11339 854 11359 856
rect 10825 850 10830 852
rect 11161 850 11165 852
rect 10790 849 10796 850
rect 10823 849 10825 850
rect 10772 844 10823 849
rect 10836 844 10842 850
rect 10886 845 10889 849
rect 11166 845 11174 849
rect 11217 846 11229 854
rect 11347 852 11379 854
rect 11262 850 11263 852
rect 11292 850 11293 852
rect 11348 847 11379 852
rect 11417 849 11419 856
rect 11417 847 11418 849
rect 10582 840 10586 844
rect 9963 836 9964 840
rect 9964 833 9965 836
rect 10011 832 10013 840
rect 10029 832 10041 840
rect 10088 838 10089 840
rect 10140 838 10141 840
rect 10087 832 10088 838
rect 10139 833 10140 838
rect 10182 832 10185 840
rect 10288 837 10289 840
rect 10287 833 10288 836
rect 10316 834 10318 840
rect 10488 837 10489 840
rect 10449 832 10453 837
rect 10540 832 10549 840
rect 10578 834 10586 840
rect 10578 832 10582 834
rect 9965 817 9973 832
rect 10011 825 10015 832
rect 10027 828 10029 832
rect 10086 828 10087 832
rect 10137 828 10138 832
rect 10013 817 10015 825
rect 10024 819 10027 828
rect 10084 819 10086 828
rect 10135 824 10137 827
rect 10131 820 10137 824
rect 9973 809 9977 817
rect 10015 811 10016 817
rect 10023 815 10024 819
rect 10083 815 10084 819
rect 10131 815 10135 820
rect 10177 819 10182 832
rect 10022 809 10023 814
rect 10081 809 10083 814
rect 10131 809 10133 815
rect 10174 814 10177 818
rect 10227 814 10243 824
rect 10245 814 10261 824
rect 10281 817 10287 832
rect 10170 809 10174 814
rect 10214 809 10221 814
rect 10266 808 10274 814
rect 10279 811 10281 817
rect 10309 811 10316 832
rect 10450 827 10454 832
rect 10489 827 10495 832
rect 10308 809 10309 811
rect 10323 808 10339 824
rect 10439 822 10505 827
rect 10525 824 10540 832
rect 10439 821 10495 822
rect 10430 814 10439 821
rect 10450 818 10454 821
rect 10346 808 10365 809
rect 10371 808 10373 809
rect 8383 805 8391 808
rect 8383 804 8385 805
rect 8386 800 8387 802
rect 8387 797 8389 800
rect 7952 758 7968 763
rect 8017 773 8078 785
rect 8085 779 8098 790
rect 8084 774 8098 779
rect 8128 774 8143 790
rect 8144 777 8146 793
rect 8237 789 8238 793
rect 8268 789 8269 795
rect 8017 759 8082 773
rect 8048 758 8064 759
rect 8066 758 8082 759
rect 8109 758 8110 760
rect 8144 758 8160 774
rect 8238 767 8242 785
rect 8269 779 8270 788
rect 8318 787 8320 794
rect 8383 790 8384 794
rect 8389 791 8392 797
rect 8424 792 8440 808
rect 8474 802 8502 808
rect 9978 804 9979 807
rect 8468 794 8502 802
rect 9979 799 9981 803
rect 10016 799 10017 803
rect 10019 800 10022 808
rect 10079 800 10081 808
rect 9981 794 9983 798
rect 10019 794 10021 800
rect 10077 794 10079 798
rect 8464 791 8466 794
rect 8474 790 8502 794
rect 8320 781 8321 787
rect 8383 782 8400 790
rect 8270 766 8275 779
rect 8322 774 8330 780
rect 8384 776 8400 782
rect 8456 779 8464 790
rect 8453 778 8464 779
rect 8468 788 8502 790
rect 8384 774 8394 776
rect 8330 773 8332 774
rect 8332 772 8333 773
rect 8242 760 8243 766
rect 8275 759 8277 766
rect 8333 765 8346 772
rect 8384 766 8385 772
rect 8400 768 8405 776
rect 8453 770 8462 778
rect 8381 765 8385 766
rect 8327 764 8360 765
rect 8381 764 8391 765
rect 8327 759 8333 764
rect 7877 756 7883 758
rect 7954 757 7968 758
rect 8080 757 8083 758
rect 7962 756 8015 757
rect 7795 754 7796 756
rect 7877 754 7886 756
rect 7559 738 7565 739
rect 7605 738 7611 744
rect 7645 738 7654 747
rect 7692 738 7701 747
rect 7784 746 7798 754
rect 7872 747 7886 754
rect 7957 750 8021 756
rect 8084 750 8099 756
rect 8106 754 8107 756
rect 8148 752 8149 753
rect 7872 746 7877 747
rect 7798 745 7801 746
rect 7871 745 7877 746
rect 7311 734 7312 736
rect 7313 727 7316 733
rect 7385 731 7400 736
rect 7553 732 7559 738
rect 7611 733 7617 738
rect 7665 734 7677 738
rect 7718 734 7734 744
rect 7796 742 7797 745
rect 7801 742 7840 745
rect 7870 743 7871 745
rect 7797 740 7840 742
rect 7801 737 7840 740
rect 7863 739 7870 743
rect 7872 739 7877 745
rect 7963 745 7978 750
rect 8009 747 8018 750
rect 7963 744 7969 745
rect 8009 744 8015 747
rect 8018 742 8032 747
rect 8099 745 8112 750
rect 8148 747 8156 752
rect 8244 751 8245 756
rect 8278 750 8281 756
rect 8333 753 8339 759
rect 8344 758 8360 764
rect 8362 758 8378 764
rect 8385 759 8391 764
rect 8405 762 8408 768
rect 8444 761 8453 770
rect 8379 753 8385 759
rect 8410 756 8412 760
rect 8440 757 8441 758
rect 8098 742 8100 745
rect 8112 742 8118 745
rect 8149 744 8156 747
rect 8245 746 8246 750
rect 8281 744 8283 750
rect 8367 745 8370 747
rect 8158 742 8159 744
rect 8412 743 8420 756
rect 8441 754 8444 757
rect 8456 756 8464 768
rect 8468 758 8470 788
rect 8499 787 8502 788
rect 8506 779 8549 791
rect 9984 785 9987 793
rect 10018 790 10020 793
rect 10021 790 10035 794
rect 10018 786 10035 790
rect 8500 776 8549 779
rect 8500 770 8509 776
rect 8520 774 8536 776
rect 8549 774 8570 776
rect 9987 775 9992 785
rect 8509 764 8518 770
rect 8512 763 8518 764
rect 8536 768 8570 774
rect 9992 771 9993 775
rect 10019 774 10035 786
rect 10069 790 10077 794
rect 10115 792 10131 808
rect 10165 801 10170 808
rect 10210 801 10214 808
rect 10266 807 10277 808
rect 10307 807 10323 808
rect 10373 807 10374 808
rect 10422 807 10430 814
rect 10453 811 10454 817
rect 10489 811 10495 821
rect 10505 814 10509 821
rect 10523 819 10540 824
rect 10571 819 10578 832
rect 10580 828 10582 832
rect 10711 832 10713 844
rect 10723 840 10735 844
rect 10751 842 10772 844
rect 10742 841 10751 842
rect 10737 840 10744 841
rect 10723 836 10737 840
rect 10523 818 10525 819
rect 10523 815 10524 818
rect 10569 817 10571 819
rect 10568 816 10569 817
rect 10509 812 10513 814
rect 10522 812 10523 813
rect 10568 812 10571 816
rect 10601 812 10613 815
rect 10495 809 10496 811
rect 10450 808 10452 809
rect 10509 808 10520 812
rect 10567 808 10568 812
rect 10601 808 10617 812
rect 10619 808 10635 824
rect 10637 808 10653 824
rect 10711 820 10719 832
rect 10723 831 10739 832
rect 10723 830 10733 831
rect 10655 808 10664 812
rect 10714 810 10715 814
rect 10439 807 10449 808
rect 10266 806 10278 807
rect 10273 804 10278 806
rect 10306 804 10323 807
rect 10374 806 10377 807
rect 10165 792 10169 801
rect 10069 774 10085 790
rect 10115 774 10131 790
rect 10165 787 10181 790
rect 10160 781 10181 787
rect 10201 787 10210 801
rect 10273 792 10277 804
rect 10305 799 10306 803
rect 10303 794 10305 798
rect 10307 792 10323 804
rect 10346 798 10358 806
rect 10377 804 10380 806
rect 10410 804 10439 807
rect 10361 799 10410 804
rect 10411 799 10417 804
rect 10422 799 10430 804
rect 10496 799 10498 804
rect 10507 803 10522 808
rect 10567 806 10572 808
rect 10601 807 10618 808
rect 10623 807 10635 808
rect 10201 785 10212 787
rect 10221 785 10233 791
rect 10273 785 10274 792
rect 10301 788 10303 792
rect 10190 783 10212 785
rect 10222 783 10233 785
rect 10272 783 10277 785
rect 10184 781 10189 783
rect 10154 775 10160 781
rect 10165 774 10181 781
rect 10199 779 10201 783
rect 10206 781 10212 783
rect 10233 781 10237 783
rect 10212 775 10218 781
rect 10221 778 10233 779
rect 10021 771 10025 774
rect 8513 759 8516 763
rect 8536 758 8552 768
rect 8570 762 8587 768
rect 8573 758 8579 762
rect 8587 760 8593 762
rect 8593 758 8597 760
rect 8619 758 8625 764
rect 8468 757 8483 758
rect 8468 756 8487 757
rect 8444 750 8449 754
rect 8484 752 8502 756
rect 8519 753 8525 756
rect 8567 753 8573 758
rect 8468 750 8502 752
rect 8525 751 8573 753
rect 8625 752 8631 758
rect 9993 754 10001 771
rect 10025 754 10032 771
rect 10035 758 10051 774
rect 10053 758 10069 774
rect 10131 772 10139 774
rect 10157 772 10165 774
rect 10231 772 10233 778
rect 10237 772 10245 779
rect 10270 778 10272 783
rect 10273 778 10277 783
rect 10270 774 10277 778
rect 10270 772 10272 774
rect 10131 758 10147 772
rect 10149 758 10165 772
rect 10212 757 10275 772
rect 10299 760 10301 786
rect 10307 774 10323 790
rect 10334 782 10342 794
rect 10346 793 10367 794
rect 10405 793 10411 799
rect 10346 792 10364 793
rect 10323 763 10327 767
rect 10334 763 10342 772
rect 10346 763 10348 792
rect 10499 788 10501 796
rect 10507 794 10529 803
rect 10507 792 10522 794
rect 10559 792 10572 806
rect 10597 804 10599 807
rect 10603 806 10617 807
rect 10601 803 10617 806
rect 10653 805 10669 808
rect 10651 803 10669 805
rect 10559 790 10567 792
rect 10589 791 10597 803
rect 10599 801 10635 803
rect 10599 793 10619 801
rect 10632 800 10635 801
rect 10633 793 10635 800
rect 10639 799 10647 803
rect 10651 799 10673 803
rect 10653 794 10673 799
rect 10711 798 10719 810
rect 10723 800 10725 830
rect 10742 826 10744 840
rect 10784 838 10790 844
rect 10842 838 10848 844
rect 10881 841 10886 845
rect 11174 841 11179 845
rect 11173 832 11181 841
rect 11185 834 11187 839
rect 11217 834 11219 846
rect 11477 845 11479 865
rect 11511 863 11513 872
rect 11548 863 11549 872
rect 11667 868 11684 881
rect 11712 868 11717 872
rect 11667 866 11676 868
rect 11667 865 11675 866
rect 11701 865 11709 866
rect 11510 857 11511 862
rect 11508 849 11509 855
rect 11229 844 11237 845
rect 11185 832 11219 834
rect 11223 832 11237 844
rect 10757 826 10758 832
rect 11229 830 11237 832
rect 10868 829 10871 830
rect 10844 827 10879 829
rect 10742 818 10743 826
rect 10840 825 10844 827
rect 10743 800 10746 814
rect 10758 812 10760 825
rect 10811 808 10840 825
rect 10842 814 10844 817
rect 10852 812 10868 827
rect 10847 811 10868 812
rect 10879 824 11039 827
rect 10723 798 10757 800
rect 10743 795 10746 798
rect 10501 778 10504 788
rect 10504 769 10506 778
rect 10507 774 10522 790
rect 10559 774 10573 790
rect 10596 781 10597 788
rect 10506 765 10507 769
rect 10323 762 10348 763
rect 10377 762 10380 763
rect 10323 760 10380 762
rect 10323 758 10339 760
rect 10507 759 10508 763
rect 8449 749 8485 750
rect 8468 744 8480 749
rect 8535 744 8546 749
rect 10001 746 10004 754
rect 10032 748 10037 754
rect 10037 745 10041 748
rect 10231 745 10233 757
rect 10236 745 10270 757
rect 10275 756 10277 757
rect 10384 756 10411 759
rect 10508 757 10509 759
rect 10523 758 10539 772
rect 10541 758 10557 772
rect 10589 769 10597 781
rect 10601 774 10619 793
rect 10653 792 10669 794
rect 10653 774 10669 790
rect 10699 774 10714 790
rect 10716 775 10718 789
rect 10723 786 10735 794
rect 10745 786 10757 794
rect 10759 790 10760 808
rect 10846 805 10856 811
rect 10879 808 11045 824
rect 11107 808 11123 824
rect 11125 808 11141 824
rect 11185 820 11197 828
rect 11207 820 11219 828
rect 11185 810 11187 820
rect 11237 816 11241 830
rect 11263 828 11265 845
rect 11265 819 11266 828
rect 11293 819 11296 845
rect 11298 843 11347 845
rect 11382 843 11384 844
rect 11298 833 11340 843
rect 11418 838 11419 843
rect 11385 827 11386 836
rect 11419 827 11420 836
rect 11476 834 11477 844
rect 11507 843 11508 847
rect 11506 837 11507 843
rect 11335 811 11340 823
rect 11387 817 11388 820
rect 11420 816 11421 820
rect 11475 819 11476 832
rect 11504 827 11506 836
rect 11546 829 11548 862
rect 11659 855 11675 865
rect 11712 864 11716 868
rect 11596 845 11659 855
rect 11704 851 11712 864
rect 11587 844 11596 845
rect 11581 842 11587 844
rect 11571 834 11581 842
rect 11503 821 11504 826
rect 11544 820 11546 827
rect 11388 811 11389 814
rect 11421 811 11422 814
rect 11474 811 11475 818
rect 11488 811 11494 817
rect 11502 816 11503 820
rect 11543 818 11544 820
rect 11551 818 11571 834
rect 11501 814 11502 816
rect 11500 812 11501 814
rect 11534 811 11540 817
rect 11542 813 11551 818
rect 11541 811 11551 813
rect 11297 808 11298 810
rect 11389 808 11390 810
rect 10851 803 10856 805
rect 10976 803 10985 808
rect 11023 803 11032 808
rect 10763 802 10772 803
rect 10761 798 10769 802
rect 10772 799 10787 802
rect 10787 798 10790 799
rect 10784 792 10790 798
rect 10842 792 10848 798
rect 10856 794 10865 803
rect 10967 794 10976 803
rect 11032 794 11041 803
rect 10958 792 10965 793
rect 10790 790 10796 792
rect 10601 772 10635 774
rect 10648 772 10653 774
rect 10746 772 10749 786
rect 10759 774 10765 790
rect 10790 786 10811 790
rect 10836 786 10842 792
rect 10952 791 10958 792
rect 11009 791 11013 793
rect 11045 792 11061 808
rect 11091 792 11107 808
rect 11118 803 11124 808
rect 11118 802 11133 803
rect 11112 796 11118 802
rect 11141 798 11157 808
rect 11164 802 11170 808
rect 11117 791 11118 793
rect 11150 791 11155 798
rect 11170 796 11176 802
rect 11188 800 11189 808
rect 10950 790 10952 791
rect 10949 787 10950 790
rect 11014 789 11016 790
rect 10795 774 10811 786
rect 10862 778 10889 781
rect 10845 774 10862 778
rect 10889 774 10897 778
rect 10601 769 10653 772
rect 10714 769 10720 772
rect 10749 771 10753 772
rect 10601 757 10605 765
rect 10637 758 10653 769
rect 10715 762 10732 769
rect 10749 762 10759 771
rect 10715 758 10731 762
rect 10732 760 10737 762
rect 10741 760 10753 762
rect 10737 759 10753 760
rect 10733 758 10753 759
rect 10811 758 10827 774
rect 10897 772 10900 774
rect 10965 772 10971 778
rect 10974 772 10976 779
rect 11016 772 11017 778
rect 11045 774 11061 790
rect 11091 774 11107 790
rect 11109 779 11118 791
rect 11044 772 11045 774
rect 10900 763 10920 772
rect 10949 767 10950 769
rect 10959 766 10965 772
rect 11017 766 11023 772
rect 11038 763 11045 772
rect 10920 762 10922 763
rect 10922 759 10928 762
rect 10277 751 10298 756
rect 10298 747 10314 751
rect 10346 748 10358 756
rect 10509 754 10510 756
rect 10405 747 10411 753
rect 10436 747 10491 753
rect 10510 750 10511 754
rect 10511 747 10513 748
rect 10520 747 10529 756
rect 10599 747 10605 756
rect 10657 747 10663 753
rect 10664 747 10673 756
rect 10718 751 10721 758
rect 8546 743 8548 744
rect 8032 739 8041 742
rect 8118 741 8120 742
rect 8420 741 8421 743
rect 10004 741 10006 745
rect 7863 738 7877 739
rect 7850 737 7863 738
rect 7870 735 7872 738
rect 8041 735 8052 739
rect 8095 737 8096 739
rect 8052 734 8055 735
rect 7661 733 7743 734
rect 7611 732 7677 733
rect 7654 731 7677 732
rect 7400 726 7412 731
rect 7654 729 7661 731
rect 7665 730 7677 731
rect 7743 729 7746 732
rect 7862 731 7869 734
rect 8055 731 8064 734
rect 8092 733 8094 736
rect 8064 729 8071 731
rect 8087 729 8091 731
rect 7650 728 7654 729
rect 7643 726 7650 728
rect 7680 727 7681 729
rect 7746 728 7748 729
rect 7102 721 7173 723
rect 6926 719 6941 720
rect 7103 719 7173 721
rect 7205 719 7209 725
rect 7316 723 7318 726
rect 6929 716 6941 719
rect 5167 705 5174 712
rect 5253 706 5263 709
rect 5264 706 5276 715
rect 5299 714 5301 715
rect 5301 709 5341 714
rect 5363 709 5375 714
rect 6865 712 6870 716
rect 6942 714 6945 716
rect 7094 712 7102 719
rect 7104 717 7114 719
rect 7138 717 7193 719
rect 7104 712 7108 717
rect 5341 707 5375 709
rect 5341 706 5389 707
rect 5411 706 5417 712
rect 5469 706 5475 712
rect 4838 698 4849 701
rect 4932 698 4940 701
rect 4960 700 4968 701
rect 4301 688 4302 692
rect 4264 676 4298 678
rect 4302 676 4310 688
rect 4397 686 4403 692
rect 4455 686 4461 692
rect 4487 688 4494 692
rect 4603 691 4609 697
rect 4649 691 4655 697
rect 4695 691 4838 698
rect 4910 691 4932 698
rect 4966 692 4968 700
rect 4969 693 4975 698
rect 4988 694 5000 701
rect 4590 688 4592 691
rect 4487 687 4499 688
rect 4403 680 4409 686
rect 4449 680 4455 686
rect 4487 685 4502 687
rect 4509 685 4521 688
rect 4589 687 4590 688
rect 4588 685 4589 687
rect 4597 685 4603 691
rect 4655 685 4661 691
rect 4662 689 4683 691
rect 4905 689 4910 691
rect 4899 687 4905 689
rect 4968 688 4969 692
rect 4977 689 4980 691
rect 4666 685 4701 687
rect 4487 680 4499 685
rect 4502 680 4524 685
rect 4586 683 4588 685
rect 4524 678 4530 680
rect 4530 676 4537 678
rect 4537 675 4542 676
rect 4551 675 4601 683
rect 4654 682 4666 685
rect 4645 680 4654 682
rect 4706 680 4708 685
rect 4889 684 4897 687
rect 4969 686 4970 687
rect 4882 682 4889 684
rect 4875 679 4882 682
rect 4970 680 4972 682
rect 4870 678 4875 679
rect 4972 678 4973 680
rect 4986 678 4993 684
rect 5005 682 5063 701
rect 5090 692 5091 698
rect 5154 692 5155 701
rect 5159 693 5167 703
rect 5174 702 5178 705
rect 5239 702 5264 706
rect 5361 704 5374 706
rect 5162 691 5167 693
rect 5178 692 5189 702
rect 5005 678 5038 682
rect 5063 678 5067 682
rect 5092 679 5093 682
rect 4644 676 4645 678
rect 4864 676 4870 678
rect 4973 676 4974 678
rect 4300 672 4302 675
rect 4542 674 4601 675
rect 4551 672 4601 674
rect 4007 656 4010 662
rect 3931 643 3995 649
rect 4005 648 4007 656
rect 4051 652 4068 672
rect 4091 666 4098 672
rect 4264 666 4276 672
rect 4286 666 4298 672
rect 4528 666 4551 672
rect 4098 664 4304 666
rect 4517 664 4528 666
rect 3937 637 3964 643
rect 3983 637 3989 643
rect 3999 642 4005 647
rect 4009 642 4018 644
rect 4068 643 4076 652
rect 4245 642 4246 660
rect 3747 626 3750 630
rect 3940 626 3964 637
rect 3999 635 4018 642
rect 4077 639 4081 642
rect 4081 636 4086 639
rect 4086 635 4094 636
rect 3999 630 4014 635
rect 4094 631 4130 635
rect 3998 626 4014 630
rect 4130 628 4150 631
rect 4244 630 4246 642
rect 4304 654 4463 664
rect 4475 654 4517 664
rect 4641 663 4644 674
rect 4708 663 4711 676
rect 4859 674 4864 676
rect 4856 673 4859 674
rect 4851 672 4856 673
rect 4845 670 4851 672
rect 4974 670 4977 676
rect 4993 671 5001 678
rect 5038 671 5046 678
rect 5067 676 5069 678
rect 5094 677 5095 687
rect 5146 681 5159 682
rect 5146 679 5155 681
rect 5189 679 5194 692
rect 5239 688 5288 702
rect 5313 698 5359 704
rect 5377 703 5379 706
rect 5389 704 5409 706
rect 5417 704 5436 706
rect 5360 700 5375 702
rect 5305 694 5313 698
rect 5239 687 5264 688
rect 5288 687 5294 688
rect 5296 687 5305 694
rect 5221 678 5239 687
rect 5288 686 5296 687
rect 5294 685 5298 686
rect 5284 677 5291 683
rect 5298 682 5306 685
rect 5306 681 5311 682
rect 5311 680 5316 681
rect 5317 678 5320 679
rect 5088 676 5109 677
rect 5146 676 5152 677
rect 5069 673 5073 676
rect 4826 668 4845 670
rect 4789 664 4826 668
rect 4712 663 4789 664
rect 4603 655 4789 663
rect 4977 660 4990 670
rect 5001 660 5023 671
rect 5046 663 5056 671
rect 5073 663 5077 673
rect 5088 671 5094 676
rect 5095 672 5109 676
rect 5135 671 5152 676
rect 5193 671 5194 676
rect 5204 671 5219 677
rect 5094 665 5100 671
rect 5140 665 5146 671
rect 5184 663 5204 671
rect 5275 669 5284 677
rect 5323 676 5328 678
rect 5329 674 5335 676
rect 4304 652 4475 654
rect 4603 653 4718 655
rect 4304 642 4306 652
rect 4603 651 4715 653
rect 4603 649 4708 651
rect 4603 648 4671 649
rect 4603 645 4655 648
rect 4597 644 4661 645
rect 4575 642 4661 644
rect 4304 634 4310 642
rect 4569 639 4586 642
rect 4597 639 4661 642
rect 4694 641 4706 649
rect 4711 643 4715 651
rect 4551 636 4569 639
rect 4305 630 4310 634
rect 4532 633 4551 636
rect 4603 633 4609 639
rect 4635 636 4641 639
rect 4649 633 4655 639
rect 4713 636 4715 643
rect 4990 642 5036 660
rect 5056 652 5086 663
rect 5066 647 5100 652
rect 5120 647 5121 660
rect 5157 652 5184 663
rect 5193 660 5194 663
rect 5066 646 5137 647
rect 5145 646 5174 652
rect 5066 643 5174 646
rect 5072 642 5077 643
rect 4990 641 5038 642
rect 4517 631 4532 633
rect 4321 630 4361 631
rect 4515 630 4517 631
rect 4160 628 4321 630
rect 4361 628 4390 630
rect 4244 626 4247 628
rect 4303 626 4310 628
rect 3750 618 3758 626
rect 3818 618 3825 625
rect 3758 617 3818 618
rect 3982 610 3998 626
rect 4247 615 4253 626
rect 4300 618 4303 625
rect 4390 622 4451 628
rect 4461 622 4511 630
rect 4711 627 4713 636
rect 4292 615 4300 618
rect 4253 613 4294 615
rect 4635 613 4648 624
rect 4689 616 4711 627
rect 4990 626 5036 641
rect 5040 637 5043 639
rect 5043 636 5045 637
rect 5045 633 5052 636
rect 5072 634 5086 642
rect 5120 634 5121 643
rect 5192 637 5193 653
rect 5234 652 5275 669
rect 5329 668 5337 674
rect 5341 670 5343 672
rect 5373 670 5375 700
rect 5379 690 5387 702
rect 5417 700 5423 704
rect 5463 700 5469 706
rect 5487 693 5498 702
rect 6870 696 6891 712
rect 6935 710 6959 712
rect 6939 705 6959 710
rect 7094 707 7104 712
rect 7101 705 7104 707
rect 6891 695 6893 696
rect 5341 668 5375 670
rect 5379 668 5387 680
rect 5498 678 5501 692
rect 6897 689 6898 692
rect 6895 678 6902 687
rect 6939 680 6941 705
rect 6945 700 6953 705
rect 6959 699 6965 705
rect 7099 701 7101 705
rect 7093 699 7101 701
rect 6965 694 6971 699
rect 7093 695 7099 699
rect 6971 692 6974 694
rect 6907 678 6941 680
rect 6945 678 6953 690
rect 6974 688 6975 692
rect 7087 689 7093 695
rect 7097 692 7098 694
rect 7096 688 7097 691
rect 7106 689 7108 712
rect 7138 712 7148 717
rect 7154 715 7193 717
rect 7169 713 7193 715
rect 7213 713 7214 715
rect 7138 701 7140 712
rect 7148 701 7161 712
rect 7174 708 7193 713
rect 7214 708 7218 713
rect 7318 710 7325 723
rect 7412 722 7442 726
rect 7661 724 7677 726
rect 7412 714 7454 722
rect 7181 701 7193 708
rect 7218 706 7219 708
rect 7325 705 7328 710
rect 7406 709 7455 710
rect 7138 695 7145 701
rect 7138 693 7151 695
rect 7138 689 7140 693
rect 7145 689 7151 693
rect 7156 691 7165 700
rect 7184 696 7193 701
rect 7224 696 7227 701
rect 7187 691 7193 696
rect 7095 685 7096 687
rect 7139 685 7140 689
rect 7157 687 7174 691
rect 7190 689 7193 691
rect 7227 689 7233 696
rect 7328 695 7365 705
rect 7406 702 7420 709
rect 7436 708 7455 709
rect 7452 703 7455 708
rect 7405 699 7406 701
rect 7365 693 7371 695
rect 7403 694 7405 699
rect 7371 692 7376 693
rect 7402 692 7403 694
rect 7192 687 7193 689
rect 7158 686 7174 687
rect 7233 686 7235 689
rect 7376 688 7392 692
rect 7392 687 7394 688
rect 6975 680 6977 685
rect 7094 680 7095 685
rect 7160 682 7163 686
rect 7165 682 7174 686
rect 7166 680 7167 682
rect 5501 676 5502 678
rect 6902 676 6903 678
rect 6906 676 6907 678
rect 7093 676 7094 678
rect 7167 677 7168 678
rect 5337 664 5340 666
rect 5341 656 5353 664
rect 5363 656 5375 664
rect 5502 661 5505 676
rect 5219 646 5234 652
rect 5341 648 5350 656
rect 5504 648 5505 661
rect 6902 660 6906 676
rect 6942 674 6945 676
rect 6907 666 6919 674
rect 6929 666 6941 674
rect 6977 660 6981 676
rect 6901 654 6902 658
rect 6981 657 6982 660
rect 5205 641 5217 646
rect 5196 637 5205 641
rect 5052 631 5058 633
rect 5070 630 5086 634
rect 5061 626 5086 630
rect 5120 626 5122 630
rect 5054 622 5079 626
rect 4649 613 4689 616
rect 4260 610 4276 613
rect 4278 610 4294 613
rect 5054 610 5070 622
rect 5079 619 5087 622
rect 5087 618 5096 619
rect 5122 615 5127 626
rect 5154 620 5196 637
rect 5151 619 5154 620
rect 5145 618 5151 619
rect 5183 618 5190 620
rect 5179 615 5183 618
rect 5127 611 5148 615
rect 5170 611 5179 615
rect 5320 606 5344 629
rect 5350 626 5389 648
rect 5389 621 5398 626
rect 5495 622 5504 643
rect 6901 630 6903 654
rect 6981 630 6982 654
rect 7093 649 7145 663
rect 7166 662 7168 675
rect 7195 672 7207 685
rect 7235 672 7247 686
rect 7397 685 7403 687
rect 7403 683 7411 685
rect 7408 681 7412 683
rect 7408 676 7415 681
rect 7452 678 7454 703
rect 7455 697 7456 702
rect 7458 698 7466 710
rect 7611 694 7639 695
rect 7675 694 7677 724
rect 7681 714 7689 726
rect 7748 712 7750 728
rect 8071 727 8077 729
rect 8084 727 8087 729
rect 7804 720 7810 726
rect 7862 720 7868 726
rect 8068 723 8088 727
rect 8120 723 8141 741
rect 8146 738 8157 740
rect 8068 721 8084 723
rect 8063 720 8068 721
rect 8088 720 8096 723
rect 7810 714 7816 720
rect 7856 714 7862 720
rect 8056 717 8063 720
rect 8096 719 8099 720
rect 8141 719 8146 723
rect 8051 716 8056 717
rect 8099 716 8105 719
rect 8146 716 8150 719
rect 8154 716 8156 738
rect 8157 737 8158 738
rect 8160 737 8168 740
rect 8158 734 8168 737
rect 8160 728 8168 734
rect 8247 733 8248 741
rect 8284 737 8287 741
rect 8248 729 8249 733
rect 8277 729 8289 737
rect 8299 729 8311 737
rect 8374 729 8387 741
rect 8166 726 8169 728
rect 8169 719 8176 726
rect 8249 724 8256 729
rect 8273 727 8276 729
rect 8289 725 8290 729
rect 8296 725 8302 729
rect 8250 723 8256 724
rect 8265 723 8273 725
rect 8277 723 8323 725
rect 8160 716 8168 718
rect 8042 713 8051 716
rect 8037 711 8042 713
rect 7456 693 7457 694
rect 7631 692 7639 694
rect 7643 692 7677 694
rect 7681 692 7689 704
rect 7748 694 7750 710
rect 8021 706 8037 711
rect 8105 706 8116 716
rect 8150 707 8168 716
rect 8176 712 8184 719
rect 8244 717 8250 723
rect 8277 717 8279 723
rect 8302 717 8308 723
rect 8309 719 8323 723
rect 8248 713 8250 714
rect 8132 706 8168 707
rect 8184 706 8192 712
rect 8246 709 8248 713
rect 8005 701 8021 706
rect 8116 705 8123 706
rect 8161 705 8194 706
rect 8116 702 8124 705
rect 8098 701 8132 702
rect 8158 701 8219 705
rect 8309 702 8311 719
rect 8315 713 8323 719
rect 8318 712 8323 713
rect 8387 712 8406 729
rect 8421 715 8455 741
rect 8550 723 8573 741
rect 10041 740 10049 745
rect 10267 742 10268 745
rect 10314 742 10334 747
rect 10334 741 10339 742
rect 10411 741 10417 747
rect 10457 741 10463 747
rect 10233 740 10235 741
rect 10006 737 10008 740
rect 10049 737 10054 740
rect 10223 739 10233 740
rect 10212 738 10233 739
rect 10339 738 10343 741
rect 10464 738 10473 747
rect 10511 745 10520 747
rect 10511 742 10526 745
rect 10511 738 10520 742
rect 10526 740 10530 742
rect 10605 741 10617 747
rect 10651 741 10664 747
rect 10720 744 10721 751
rect 10530 739 10533 740
rect 10054 736 10056 737
rect 10221 736 10240 738
rect 10009 733 10010 736
rect 10056 733 10060 736
rect 10010 727 10013 733
rect 10060 731 10064 733
rect 10064 729 10067 731
rect 10154 729 10160 735
rect 10212 729 10218 735
rect 10221 733 10258 736
rect 10265 733 10266 736
rect 10232 729 10258 733
rect 10261 729 10265 731
rect 10297 729 10298 730
rect 10067 726 10071 729
rect 10013 720 10017 726
rect 10071 720 10081 726
rect 10084 720 10096 724
rect 10160 723 10166 729
rect 10206 723 10212 729
rect 10258 726 10298 729
rect 10258 723 10297 726
rect 10343 725 10360 738
rect 10464 737 10465 738
rect 10533 736 10540 739
rect 10608 738 10617 741
rect 10655 738 10664 741
rect 10714 739 10721 744
rect 10749 742 10753 758
rect 10791 747 10800 756
rect 10856 747 10865 756
rect 10928 754 10939 759
rect 11032 758 11045 763
rect 11107 772 11108 774
rect 11107 769 11116 772
rect 11117 769 11118 779
rect 11107 763 11118 769
rect 11121 763 11123 791
rect 11189 790 11191 791
rect 11187 785 11191 790
rect 11240 790 11241 808
rect 11347 799 11359 804
rect 11391 796 11392 799
rect 11422 796 11423 805
rect 11473 799 11474 808
rect 11482 805 11488 811
rect 11540 808 11546 811
rect 11595 808 11611 824
rect 12184 819 12185 1015
rect 12374 819 12375 1015
rect 12460 819 12461 1015
rect 12733 819 12734 1015
rect 12930 819 12931 1015
rect 13323 1014 13327 1019
rect 13961 1014 13968 1019
rect 14048 1018 14057 1027
rect 14113 1024 14209 1027
rect 14550 1023 14658 1037
rect 14408 1015 14424 1022
rect 14426 1015 14442 1022
rect 13968 1007 13980 1014
rect 14398 1013 14410 1015
rect 14420 1013 14432 1015
rect 14438 1013 14442 1015
rect 14626 1013 14642 1022
rect 14658 1021 14676 1023
rect 14677 1017 14684 1020
rect 14684 1013 14690 1017
rect 15330 1015 15331 1026
rect 15520 1015 15521 1026
rect 15606 1015 15607 1026
rect 15879 1015 15880 1026
rect 16076 1015 16077 1026
rect 16505 1023 16606 1034
rect 16792 1033 17056 1034
rect 17056 1023 17111 1033
rect 17214 1027 17223 1036
rect 17261 1027 17270 1036
rect 17564 1034 17686 1037
rect 17536 1033 17553 1034
rect 17366 1027 17536 1033
rect 16490 1021 16505 1023
rect 16484 1019 16490 1021
rect 17113 1019 17118 1021
rect 14398 1008 14442 1013
rect 14585 1008 14622 1009
rect 14690 1008 14693 1013
rect 14394 1006 14396 1008
rect 14398 1006 14530 1008
rect 13449 1005 13803 1006
rect 13429 1003 13447 1005
rect 13889 1003 13902 1005
rect 13981 1003 13984 1005
rect 14392 1003 14530 1006
rect 13373 1000 13429 1003
rect 13247 992 13259 1000
rect 13269 992 13281 1000
rect 13345 994 13429 1000
rect 13902 994 13912 1003
rect 13345 993 13373 994
rect 13243 989 13245 992
rect 13345 991 13364 993
rect 13913 991 13916 993
rect 13285 988 13289 989
rect 13235 977 13243 988
rect 13246 986 13281 988
rect 13244 977 13246 983
rect 13235 976 13244 977
rect 13243 972 13244 976
rect 13242 971 13243 972
rect 13240 966 13242 969
rect 13115 964 13180 965
rect 13107 956 13115 964
rect 13180 956 13184 964
rect 13106 950 13107 956
rect 13235 954 13243 966
rect 13247 956 13249 986
rect 13278 985 13281 986
rect 13280 979 13281 985
rect 13285 981 13293 988
rect 13289 980 13297 981
rect 13321 980 13322 990
rect 13345 980 13360 991
rect 13619 981 13656 983
rect 13297 979 13303 980
rect 13320 979 13321 980
rect 13345 979 13352 980
rect 13303 969 13365 979
rect 13373 972 13379 978
rect 13419 972 13425 978
rect 13619 977 13645 981
rect 13656 977 13661 981
rect 13916 980 13929 991
rect 13892 979 13906 980
rect 13613 972 13619 977
rect 13661 972 13670 977
rect 13874 972 13892 979
rect 13906 977 13913 979
rect 13984 977 14005 1003
rect 14386 996 14530 1003
rect 14546 1006 14647 1008
rect 14546 996 14658 1006
rect 14347 990 14408 996
rect 14312 987 14347 990
rect 14125 981 14312 987
rect 14398 986 14408 990
rect 13913 972 13928 977
rect 13367 969 13373 972
rect 13374 970 13431 972
rect 13670 971 13671 972
rect 13508 970 13511 971
rect 13529 970 13532 971
rect 13611 970 13612 971
rect 13671 970 13674 971
rect 13374 969 13382 970
rect 13345 968 13382 969
rect 13247 954 13281 956
rect 13236 951 13238 954
rect 13232 938 13236 950
rect 13247 942 13259 950
rect 13272 945 13281 954
rect 13319 952 13320 955
rect 13345 951 13350 968
rect 13367 966 13382 968
rect 13425 966 13431 970
rect 13504 967 13508 970
rect 13532 967 13537 970
rect 13674 968 13675 970
rect 13866 969 13874 972
rect 13903 971 13928 972
rect 13937 971 13941 972
rect 13899 970 13903 971
rect 13913 970 13950 971
rect 13675 967 13678 968
rect 13373 964 13382 966
rect 13373 951 13378 964
rect 13426 955 13445 958
rect 13480 955 13504 967
rect 13537 959 13555 967
rect 13610 959 13611 967
rect 13282 949 13287 950
rect 13287 948 13292 949
rect 13292 947 13295 948
rect 13297 945 13306 947
rect 13270 942 13272 945
rect 13306 944 13311 945
rect 13311 943 13317 944
rect 13318 943 13319 951
rect 13345 943 13351 951
rect 13269 939 13270 942
rect 13317 938 13351 943
rect 13230 931 13232 937
rect 13267 930 13269 938
rect 13318 932 13319 938
rect 13345 935 13373 938
rect 13345 933 13375 935
rect 13345 931 13376 933
rect 13377 931 13378 951
rect 13445 946 13507 955
rect 13555 952 13563 959
rect 13609 951 13610 958
rect 13678 954 13682 967
rect 13858 966 13866 969
rect 13896 968 13899 970
rect 13892 967 13896 968
rect 13887 965 13892 967
rect 13913 965 13928 970
rect 13937 969 13941 970
rect 13950 969 13951 970
rect 14007 969 14012 975
rect 14048 971 14057 980
rect 14113 978 14125 981
rect 14113 971 14122 978
rect 14392 972 14408 986
rect 14431 972 14432 996
rect 14437 991 14458 996
rect 14442 990 14458 991
rect 14575 989 14581 996
rect 14627 989 14633 996
rect 14647 990 14658 996
rect 14693 990 14702 1008
rect 14442 972 14458 988
rect 14575 985 14583 989
rect 14581 983 14583 985
rect 14491 974 14519 978
rect 14521 974 14532 978
rect 13941 965 13946 969
rect 13951 965 13953 968
rect 14012 965 14015 969
rect 13853 964 13857 965
rect 13928 964 13931 965
rect 13953 964 13954 965
rect 13849 962 13853 964
rect 13463 945 13473 946
rect 13495 945 13496 946
rect 13459 943 13463 945
rect 13507 943 13527 946
rect 13608 943 13609 950
rect 13681 943 13682 950
rect 13816 949 13849 962
rect 13933 959 13937 962
rect 13948 960 13952 963
rect 14057 962 14066 971
rect 14090 961 14093 963
rect 14104 962 14113 971
rect 14398 970 14432 972
rect 14441 971 14442 972
rect 14488 971 14491 974
rect 14437 970 14442 971
rect 14487 970 14488 971
rect 14398 968 14442 970
rect 14485 969 14487 970
rect 14394 965 14395 967
rect 14168 961 14177 963
rect 14085 959 14090 961
rect 13730 943 13736 949
rect 13776 948 13782 949
rect 13813 948 13816 949
rect 13776 947 13813 948
rect 13776 943 13782 947
rect 13868 946 13874 952
rect 13914 946 13920 952
rect 13936 949 13937 959
rect 14083 958 14085 959
rect 14179 958 14185 961
rect 13954 955 13958 958
rect 14022 955 14024 958
rect 13958 946 13968 955
rect 13447 931 13455 943
rect 13459 941 13493 943
rect 13183 924 13184 929
rect 13133 915 13142 924
rect 13180 920 13189 924
rect 13180 915 13194 920
rect 13124 912 13133 915
rect 13124 911 13127 912
rect 13117 908 13126 911
rect 13105 907 13126 908
rect 13105 905 13123 907
rect 13163 905 13169 911
rect 13183 906 13198 915
rect 13223 908 13230 929
rect 13105 900 13117 905
rect 13101 898 13104 900
rect 13105 899 13106 900
rect 13111 899 13117 900
rect 13169 899 13175 905
rect 13182 904 13194 906
rect 13221 904 13223 908
rect 13261 907 13267 929
rect 13318 926 13319 929
rect 13345 928 13406 931
rect 13345 917 13351 928
rect 13373 926 13406 928
rect 13367 925 13406 926
rect 13425 925 13431 926
rect 13367 921 13431 925
rect 13367 920 13453 921
rect 13345 913 13354 917
rect 13373 914 13379 920
rect 13419 914 13425 920
rect 13428 917 13453 920
rect 13437 913 13453 917
rect 13459 913 13461 941
rect 13490 939 13493 941
rect 13345 909 13360 913
rect 13447 909 13461 913
rect 13491 909 13493 939
rect 13497 931 13505 943
rect 13527 934 13590 943
rect 13724 938 13730 943
rect 13742 941 13778 943
rect 13742 938 13747 941
rect 13683 937 13730 938
rect 13744 937 13747 938
rect 13782 937 13788 943
rect 13862 940 13868 946
rect 13920 940 13926 946
rect 13683 936 13726 937
rect 13607 934 13608 936
rect 13629 934 13683 936
rect 13563 922 13578 934
rect 13590 933 13629 934
rect 13607 929 13608 933
rect 13739 929 13742 936
rect 13866 933 13868 934
rect 13864 929 13866 933
rect 13260 904 13261 906
rect 13320 905 13321 909
rect 13180 899 13182 904
rect 13326 903 13332 909
rect 13345 903 13364 909
rect 13372 903 13378 909
rect 13220 899 13221 903
rect 13179 897 13180 899
rect 13219 897 13220 899
rect 13093 884 13101 896
rect 13105 894 13123 896
rect 13178 895 13179 896
rect 13258 895 13260 903
rect 13320 897 13326 903
rect 13345 897 13384 903
rect 13386 897 13398 905
rect 13459 904 13476 909
rect 13467 899 13474 904
rect 13476 903 13480 904
rect 13496 903 13497 905
rect 13563 904 13578 920
rect 13605 906 13607 928
rect 13480 900 13499 903
rect 13604 900 13616 905
rect 13626 900 13638 905
rect 13679 904 13681 928
rect 13730 904 13739 928
rect 13775 904 13778 909
rect 13816 908 13851 910
rect 13862 908 13864 929
rect 13886 909 13887 929
rect 13934 928 13936 944
rect 13968 942 13973 946
rect 14024 942 14036 955
rect 14185 951 14198 958
rect 14408 956 14424 968
rect 14426 956 14442 968
rect 14481 965 14485 968
rect 14479 963 14481 965
rect 14477 961 14479 963
rect 14532 961 14545 974
rect 14581 967 14584 983
rect 14583 961 14584 967
rect 14587 967 14588 989
rect 14626 985 14633 989
rect 14654 987 14656 990
rect 14626 983 14627 985
rect 14647 984 14648 986
rect 14587 963 14589 967
rect 14620 963 14621 966
rect 14625 965 14627 983
rect 14656 981 14659 987
rect 14659 979 14660 981
rect 14661 975 14662 977
rect 14662 972 14663 975
rect 14702 973 14710 990
rect 14664 965 14667 969
rect 14587 961 14591 963
rect 14625 962 14626 965
rect 14667 963 14668 965
rect 14473 958 14476 961
rect 14545 959 14548 961
rect 14471 953 14473 958
rect 14548 957 14550 959
rect 14306 952 14343 953
rect 14470 952 14471 953
rect 14550 952 14552 957
rect 14578 955 14584 961
rect 14591 959 14597 961
rect 14598 957 14604 959
rect 14624 957 14630 961
rect 14668 960 14669 963
rect 14669 958 14670 960
rect 14604 956 14630 957
rect 14306 951 14331 952
rect 14343 951 14344 952
rect 14200 948 14204 951
rect 14271 948 14298 951
rect 14346 948 14353 951
rect 14398 949 14399 952
rect 14469 951 14470 952
rect 14353 943 14364 948
rect 14399 945 14401 949
rect 14434 947 14435 949
rect 14467 948 14469 951
rect 14364 942 14368 943
rect 14036 939 14037 942
rect 14368 938 14375 942
rect 13978 929 13988 938
rect 14038 931 14044 938
rect 14375 937 14377 938
rect 14377 933 14393 937
rect 14393 932 14398 933
rect 14401 932 14409 944
rect 14398 929 14409 932
rect 14435 929 14439 944
rect 14465 943 14467 948
rect 14552 944 14555 951
rect 14572 949 14578 955
rect 14604 951 14648 956
rect 14670 955 14672 958
rect 14630 949 14636 951
rect 14672 948 14675 955
rect 14464 942 14465 943
rect 14675 942 14678 948
rect 14710 943 14711 973
rect 14818 951 14834 954
rect 14746 943 14769 951
rect 14824 943 14841 951
rect 14463 940 14464 942
rect 14462 939 14463 940
rect 14678 939 14679 942
rect 14461 937 14462 938
rect 14458 933 14461 937
rect 14456 932 14458 933
rect 14454 929 14456 932
rect 14679 931 14680 938
rect 14709 929 14710 942
rect 14738 938 14746 943
rect 14824 938 14848 943
rect 14728 932 14738 938
rect 14721 929 14728 932
rect 13931 917 13933 920
rect 13927 914 13930 916
rect 13925 913 13927 914
rect 13922 911 13925 913
rect 13920 910 13922 911
rect 13806 906 13816 908
rect 13851 906 13868 908
rect 13795 904 13806 906
rect 13729 900 13730 903
rect 13773 900 13775 904
rect 13787 902 13795 904
rect 13783 901 13787 902
rect 13862 900 13864 906
rect 13886 904 13887 906
rect 13954 904 13970 920
rect 13988 910 14010 929
rect 14048 920 14056 927
rect 14056 918 14063 920
rect 14063 914 14079 918
rect 14082 914 14083 929
rect 14401 928 14414 929
rect 14407 927 14414 928
rect 14439 927 14440 928
rect 14453 927 14454 929
rect 14577 927 14578 929
rect 14409 923 14410 926
rect 14414 924 14451 927
rect 14141 921 14172 922
rect 14132 920 14141 921
rect 14172 920 14179 921
rect 14439 920 14440 924
rect 14103 917 14132 920
rect 14179 917 14194 920
rect 14101 916 14103 917
rect 14094 914 14101 916
rect 14194 914 14206 917
rect 14411 915 14412 917
rect 14440 915 14441 920
rect 14445 915 14454 924
rect 14492 915 14501 924
rect 14576 922 14577 927
rect 14575 920 14576 922
rect 14574 918 14575 920
rect 14573 916 14574 918
rect 14436 914 14445 915
rect 14079 911 14445 914
rect 14082 910 14083 911
rect 14085 910 14087 911
rect 14221 910 14229 911
rect 14010 909 14012 910
rect 13887 900 13891 904
rect 13941 900 13954 904
rect 14012 903 14020 909
rect 14081 908 14085 910
rect 14229 906 14247 910
rect 14412 906 14413 909
rect 14442 906 14443 909
rect 14074 904 14079 906
rect 13345 895 13400 897
rect 13474 895 13480 899
rect 13494 898 13495 900
rect 13493 895 13494 897
rect 13499 896 13668 900
rect 13727 897 13729 900
rect 13724 896 13730 897
rect 13770 896 13773 900
rect 13604 895 13605 896
rect 13668 895 13730 896
rect 13093 862 13101 874
rect 13105 865 13107 894
rect 13177 893 13178 894
rect 13218 893 13219 894
rect 13345 893 13402 895
rect 13480 893 13481 895
rect 13172 889 13178 893
rect 13217 889 13218 893
rect 13257 889 13258 893
rect 13313 889 13320 893
rect 13345 892 13410 893
rect 13158 888 13178 889
rect 13158 878 13172 888
rect 13214 879 13217 889
rect 13255 878 13257 889
rect 13310 879 13313 889
rect 13142 866 13158 878
rect 13105 862 13108 865
rect 13139 862 13142 866
rect 13189 859 13198 868
rect 13210 866 13214 878
rect 13254 875 13255 878
rect 13309 875 13310 878
rect 13209 862 13210 866
rect 13104 857 13106 858
rect 13111 857 13117 859
rect 13105 853 13117 857
rect 13169 853 13175 859
rect 13181 857 13189 859
rect 13208 858 13209 862
rect 13250 859 13254 875
rect 13304 859 13309 875
rect 13322 864 13325 892
rect 13372 891 13398 892
rect 13396 861 13398 891
rect 13402 881 13410 892
rect 13481 879 13501 893
rect 13549 879 13563 894
rect 13592 881 13600 893
rect 13604 891 13638 893
rect 13457 876 13458 879
rect 13487 876 13488 879
rect 13501 877 13513 879
rect 13547 877 13549 879
rect 13501 875 13547 877
rect 13372 859 13398 861
rect 13402 859 13410 871
rect 13455 869 13457 875
rect 13485 870 13487 875
rect 13453 862 13455 869
rect 13482 862 13485 869
rect 13452 859 13453 862
rect 13481 859 13482 862
rect 13604 859 13606 891
rect 13636 875 13638 891
rect 13642 881 13650 893
rect 13724 891 13730 895
rect 13768 891 13770 895
rect 13782 891 13788 897
rect 13862 894 13868 900
rect 13891 896 13906 900
rect 13906 895 13907 896
rect 13920 895 13954 900
rect 14020 899 14026 903
rect 14071 902 14074 904
rect 14247 902 14267 906
rect 14338 902 14351 903
rect 13678 881 13679 889
rect 13722 881 13725 891
rect 13730 885 13736 891
rect 13762 881 13768 891
rect 13776 885 13782 891
rect 13865 883 13866 891
rect 13868 888 13874 894
rect 13907 893 13926 895
rect 13637 865 13638 874
rect 13642 872 13643 875
rect 13672 870 13678 880
rect 13717 870 13722 881
rect 13660 866 13672 870
rect 13716 867 13717 870
rect 13755 867 13762 881
rect 13905 872 13908 892
rect 13914 888 13920 893
rect 13938 888 13954 895
rect 14026 894 14037 899
rect 14065 898 14069 900
rect 14062 897 14065 898
rect 14059 895 14062 897
rect 14082 895 14085 900
rect 14267 897 14292 902
rect 14317 900 14335 902
rect 14356 900 14379 902
rect 14315 899 14327 900
rect 14379 899 14388 900
rect 14388 898 14389 899
rect 14413 898 14414 902
rect 14292 895 14297 897
rect 14308 895 14315 898
rect 14037 885 14068 894
rect 14085 893 14087 895
rect 14087 891 14089 893
rect 14297 891 14315 895
rect 14389 894 14396 898
rect 14443 897 14444 902
rect 14501 901 14510 915
rect 14571 911 14572 914
rect 14598 909 14630 913
rect 14565 903 14569 906
rect 14572 903 14578 909
rect 14598 904 14636 909
rect 14667 904 14721 929
rect 14824 922 14850 938
rect 14595 903 14636 904
rect 14552 901 14564 902
rect 14510 899 14514 901
rect 14532 900 14552 901
rect 14526 899 14532 900
rect 14552 895 14554 900
rect 14578 897 14584 903
rect 14612 899 14613 901
rect 14396 891 14402 894
rect 14414 891 14415 895
rect 14027 880 14068 885
rect 14089 888 14162 891
rect 14297 889 14314 891
rect 14089 885 14169 888
rect 14089 881 14162 885
rect 14169 881 14239 885
rect 14300 882 14308 889
rect 14314 887 14319 889
rect 14319 885 14323 887
rect 14402 885 14415 891
rect 14444 887 14446 895
rect 14550 892 14552 895
rect 14549 891 14550 892
rect 14027 876 14043 880
rect 14068 876 14086 880
rect 14089 876 14107 881
rect 14162 876 14267 881
rect 14086 875 14267 876
rect 14293 875 14300 882
rect 14323 876 14345 885
rect 14402 882 14416 885
rect 14415 881 14418 882
rect 14415 878 14416 881
rect 14418 880 14419 881
rect 14419 879 14428 880
rect 14446 879 14448 885
rect 14537 882 14549 891
rect 14531 881 14537 882
rect 14503 880 14519 881
rect 14527 880 14531 881
rect 14596 880 14611 899
rect 14624 897 14630 903
rect 14661 901 14667 904
rect 14675 903 14676 904
rect 14650 895 14661 901
rect 14674 899 14675 901
rect 14647 892 14650 895
rect 14646 891 14647 892
rect 14638 885 14646 891
rect 14475 879 14498 880
rect 14345 875 14348 876
rect 13754 866 13755 867
rect 13659 865 13660 866
rect 13637 862 13659 865
rect 13713 862 13716 866
rect 13638 859 13659 862
rect 13710 859 13716 862
rect 13180 855 13189 857
rect 13105 852 13114 853
rect 13105 850 13115 852
rect 13117 850 13123 853
rect 13115 847 13123 850
rect 13115 842 13119 847
rect 13168 840 13169 853
rect 13178 852 13189 855
rect 13176 851 13178 852
rect 13173 850 13176 851
rect 13180 850 13189 852
rect 13204 845 13208 858
rect 13247 846 13250 858
rect 13300 846 13304 858
rect 13320 851 13326 857
rect 13349 856 13353 859
rect 13643 858 13644 859
rect 13326 845 13332 851
rect 13344 845 13349 856
rect 13378 851 13384 857
rect 13451 855 13452 858
rect 13480 855 13481 858
rect 13710 857 13713 859
rect 13712 856 13713 857
rect 13708 855 13712 856
rect 13372 845 13378 851
rect 13386 847 13398 855
rect 13602 853 13603 855
rect 13200 841 13204 845
rect 13246 841 13247 845
rect 13298 842 13300 845
rect 13198 840 13200 841
rect 13342 840 13344 845
rect 13446 841 13449 850
rect 13476 841 13479 850
rect 13603 841 13605 849
rect 13644 842 13645 849
rect 13705 847 13712 855
rect 13699 845 13706 847
rect 13708 845 13712 847
rect 13742 845 13754 865
rect 13866 859 13868 872
rect 13699 840 13708 845
rect 13739 844 13746 845
rect 13901 844 13905 870
rect 14016 869 14026 875
rect 14079 872 14279 875
rect 14290 872 14293 875
rect 14348 872 14358 875
rect 14364 872 14376 878
rect 14419 875 14498 879
rect 14626 876 14658 885
rect 14671 880 14674 898
rect 14670 876 14671 880
rect 14706 878 14708 904
rect 14824 895 14847 922
rect 14879 895 14880 929
rect 14824 881 14846 895
rect 14858 889 14880 895
rect 14079 871 14087 872
rect 14074 869 14078 871
rect 14014 868 14016 869
rect 14011 866 14014 868
rect 14069 866 14073 868
rect 14162 867 14386 872
rect 14416 871 14417 875
rect 14428 871 14475 875
rect 14589 872 14592 876
rect 14623 875 14658 876
rect 14434 869 14475 871
rect 14440 868 14465 869
rect 14178 866 14386 867
rect 14004 862 14011 866
rect 14059 862 14069 866
rect 14178 863 14388 866
rect 14291 862 14300 863
rect 14374 862 14396 863
rect 14417 862 14418 868
rect 14441 867 14465 868
rect 14581 863 14589 872
rect 14636 869 14637 874
rect 13998 858 14004 862
rect 14300 858 14307 862
rect 13996 857 13998 858
rect 13987 852 13996 857
rect 14307 852 14318 858
rect 14374 854 14388 862
rect 14396 856 14429 862
rect 14448 859 14449 862
rect 14577 857 14581 862
rect 14504 856 14516 857
rect 14429 855 14435 856
rect 14453 855 14475 856
rect 14435 854 14475 855
rect 14496 854 14516 856
rect 13982 850 13987 852
rect 14318 850 14322 852
rect 13947 849 13953 850
rect 13980 849 13982 850
rect 13929 844 13980 849
rect 13993 844 13999 850
rect 14043 845 14046 849
rect 14323 845 14331 849
rect 14374 846 14386 854
rect 14504 852 14536 854
rect 14419 850 14420 852
rect 14449 850 14450 852
rect 14505 847 14536 852
rect 14574 849 14576 856
rect 14574 847 14575 849
rect 13739 840 13743 844
rect 13120 836 13121 840
rect 13121 833 13122 836
rect 13168 832 13170 840
rect 13186 832 13198 840
rect 13245 838 13246 840
rect 13297 838 13298 840
rect 13244 832 13245 838
rect 13296 833 13297 838
rect 13339 832 13342 840
rect 13445 837 13446 840
rect 13444 833 13445 836
rect 13473 834 13475 840
rect 13645 837 13646 840
rect 13606 832 13610 837
rect 13697 832 13706 840
rect 13735 834 13743 840
rect 13735 832 13739 834
rect 13122 817 13130 832
rect 13168 825 13172 832
rect 13184 828 13186 832
rect 13243 828 13244 832
rect 13294 828 13295 832
rect 13170 817 13172 825
rect 13181 819 13184 828
rect 13241 819 13243 828
rect 13292 824 13294 827
rect 13288 820 13294 824
rect 13130 809 13134 817
rect 13172 811 13173 817
rect 13180 815 13181 819
rect 13240 815 13241 819
rect 13288 815 13292 820
rect 13334 819 13339 832
rect 13179 809 13180 814
rect 13238 809 13240 814
rect 13288 809 13290 815
rect 13331 814 13334 818
rect 13384 814 13400 824
rect 13402 814 13418 824
rect 13438 817 13444 832
rect 13327 809 13331 814
rect 13371 809 13378 814
rect 13423 808 13431 814
rect 13436 811 13438 817
rect 13466 811 13473 832
rect 13607 827 13611 832
rect 13646 827 13652 832
rect 13465 809 13466 811
rect 13480 808 13496 824
rect 13596 822 13662 827
rect 13682 824 13697 832
rect 13596 821 13652 822
rect 13587 814 13596 821
rect 13607 818 13611 821
rect 13503 808 13522 809
rect 13528 808 13530 809
rect 11538 805 11546 808
rect 11538 804 11540 805
rect 11541 800 11542 802
rect 11542 797 11544 800
rect 11107 758 11123 763
rect 11172 773 11233 785
rect 11240 779 11253 790
rect 11239 774 11253 779
rect 11283 774 11298 790
rect 11299 777 11301 793
rect 11392 789 11393 793
rect 11423 789 11424 795
rect 11172 759 11237 773
rect 11203 758 11219 759
rect 11221 758 11237 759
rect 11264 758 11265 760
rect 11299 758 11315 774
rect 11393 767 11397 785
rect 11424 779 11425 788
rect 11473 787 11475 794
rect 11538 790 11539 794
rect 11544 791 11547 797
rect 11579 792 11595 808
rect 11629 802 11657 808
rect 13135 804 13136 807
rect 11623 794 11657 802
rect 13136 799 13138 803
rect 13173 799 13174 803
rect 13176 800 13179 808
rect 13236 800 13238 808
rect 13138 794 13140 798
rect 13176 794 13178 800
rect 13234 794 13236 798
rect 11619 791 11621 794
rect 11629 790 11657 794
rect 11475 781 11476 787
rect 11538 782 11555 790
rect 11425 766 11430 779
rect 11477 774 11485 780
rect 11539 776 11555 782
rect 11611 779 11619 790
rect 11608 778 11619 779
rect 11623 788 11657 790
rect 11539 774 11549 776
rect 11485 773 11487 774
rect 11487 772 11488 773
rect 11397 760 11398 766
rect 11430 759 11432 766
rect 11488 765 11501 772
rect 11539 766 11540 772
rect 11555 768 11560 776
rect 11608 770 11617 778
rect 11536 765 11540 766
rect 11482 764 11515 765
rect 11536 764 11546 765
rect 11482 759 11488 764
rect 11032 756 11038 758
rect 11109 757 11123 758
rect 11235 757 11238 758
rect 11117 756 11170 757
rect 10950 754 10951 756
rect 11032 754 11041 756
rect 10714 738 10720 739
rect 10760 738 10766 744
rect 10800 738 10809 747
rect 10847 738 10856 747
rect 10939 746 10953 754
rect 11027 747 11041 754
rect 11112 750 11176 756
rect 11239 750 11254 756
rect 11261 754 11262 756
rect 11303 752 11304 753
rect 11027 746 11032 747
rect 10953 745 10956 746
rect 11026 745 11032 746
rect 10466 734 10467 736
rect 10468 727 10471 733
rect 10540 731 10555 736
rect 10708 732 10714 738
rect 10766 733 10772 738
rect 10820 734 10832 738
rect 10873 734 10889 744
rect 10951 742 10952 745
rect 10956 742 10995 745
rect 11025 743 11026 745
rect 10952 740 10995 742
rect 10956 737 10995 740
rect 11018 739 11025 743
rect 11027 739 11032 745
rect 11118 745 11133 750
rect 11164 747 11173 750
rect 11118 744 11124 745
rect 11164 744 11170 747
rect 11173 742 11187 747
rect 11254 745 11267 750
rect 11303 747 11311 752
rect 11399 751 11400 756
rect 11433 750 11436 756
rect 11488 753 11494 759
rect 11499 758 11515 764
rect 11517 758 11533 764
rect 11540 759 11546 764
rect 11560 762 11563 768
rect 11599 761 11608 770
rect 11534 753 11540 759
rect 11565 756 11567 760
rect 11595 757 11596 758
rect 11253 742 11255 745
rect 11267 742 11273 745
rect 11304 744 11311 747
rect 11400 746 11401 750
rect 11436 744 11438 750
rect 11522 745 11525 747
rect 11313 742 11314 744
rect 11567 743 11575 756
rect 11596 754 11599 757
rect 11611 756 11619 768
rect 11623 758 11625 788
rect 11654 787 11657 788
rect 11661 779 11704 791
rect 13141 785 13144 793
rect 13175 790 13177 793
rect 13178 790 13192 794
rect 13175 786 13192 790
rect 11655 776 11704 779
rect 11655 770 11664 776
rect 11675 774 11691 776
rect 11704 774 11725 776
rect 13144 775 13149 785
rect 11664 764 11673 770
rect 11667 763 11673 764
rect 11691 768 11725 774
rect 13149 771 13150 775
rect 13176 774 13192 786
rect 13226 790 13234 794
rect 13272 792 13288 808
rect 13322 801 13327 808
rect 13367 801 13371 808
rect 13423 807 13434 808
rect 13464 807 13480 808
rect 13530 807 13531 808
rect 13579 807 13587 814
rect 13610 811 13611 817
rect 13646 811 13652 821
rect 13662 814 13666 821
rect 13680 819 13697 824
rect 13728 819 13735 832
rect 13737 828 13739 832
rect 13868 832 13870 844
rect 13880 840 13892 844
rect 13908 842 13929 844
rect 13899 841 13908 842
rect 13894 840 13901 841
rect 13880 836 13894 840
rect 13680 818 13682 819
rect 13680 815 13681 818
rect 13726 817 13728 819
rect 13725 816 13726 817
rect 13666 812 13670 814
rect 13679 812 13680 813
rect 13725 812 13728 816
rect 13758 812 13770 815
rect 13652 809 13653 811
rect 13607 808 13609 809
rect 13666 808 13677 812
rect 13724 808 13725 812
rect 13758 808 13774 812
rect 13776 808 13792 824
rect 13794 808 13810 824
rect 13868 820 13876 832
rect 13880 831 13896 832
rect 13880 830 13890 831
rect 13812 808 13821 812
rect 13871 810 13872 814
rect 13596 807 13606 808
rect 13423 806 13435 807
rect 13430 804 13435 806
rect 13463 804 13480 807
rect 13531 806 13534 807
rect 13322 792 13326 801
rect 13226 774 13242 790
rect 13272 774 13288 790
rect 13322 787 13338 790
rect 13317 781 13338 787
rect 13358 787 13367 801
rect 13430 792 13434 804
rect 13462 799 13463 803
rect 13460 794 13462 798
rect 13464 792 13480 804
rect 13503 798 13515 806
rect 13534 804 13537 806
rect 13567 804 13596 807
rect 13518 799 13567 804
rect 13568 799 13574 804
rect 13579 799 13587 804
rect 13653 799 13655 804
rect 13664 803 13679 808
rect 13724 806 13729 808
rect 13758 807 13775 808
rect 13780 807 13792 808
rect 13358 785 13369 787
rect 13378 785 13390 791
rect 13430 785 13431 792
rect 13458 788 13460 792
rect 13347 783 13369 785
rect 13379 783 13390 785
rect 13429 783 13434 785
rect 13341 781 13346 783
rect 13311 775 13317 781
rect 13322 774 13338 781
rect 13356 779 13358 783
rect 13363 781 13369 783
rect 13390 781 13394 783
rect 13369 775 13375 781
rect 13378 778 13390 779
rect 13178 771 13182 774
rect 11668 759 11671 763
rect 11691 758 11707 768
rect 11725 762 11742 768
rect 11728 758 11734 762
rect 11742 760 11748 762
rect 11748 758 11752 760
rect 11774 758 11780 764
rect 11623 757 11638 758
rect 11623 756 11642 757
rect 11599 750 11604 754
rect 11639 752 11657 756
rect 11674 753 11680 756
rect 11722 753 11728 758
rect 11623 750 11657 752
rect 11680 751 11728 753
rect 11780 752 11786 758
rect 13150 754 13158 771
rect 13182 754 13189 771
rect 13192 758 13208 774
rect 13210 758 13226 774
rect 13288 772 13296 774
rect 13314 772 13322 774
rect 13388 772 13390 778
rect 13394 772 13402 779
rect 13427 778 13429 783
rect 13430 778 13434 783
rect 13427 774 13434 778
rect 13427 772 13429 774
rect 13288 758 13304 772
rect 13306 758 13322 772
rect 13369 757 13432 772
rect 13456 760 13458 786
rect 13464 774 13480 790
rect 13491 782 13499 794
rect 13503 793 13524 794
rect 13562 793 13568 799
rect 13503 792 13521 793
rect 13480 763 13484 767
rect 13491 763 13499 772
rect 13503 763 13505 792
rect 13656 788 13658 796
rect 13664 794 13686 803
rect 13664 792 13679 794
rect 13716 792 13729 806
rect 13754 804 13756 807
rect 13760 806 13774 807
rect 13758 803 13774 806
rect 13810 805 13826 808
rect 13808 803 13826 805
rect 13716 790 13724 792
rect 13746 791 13754 803
rect 13756 801 13792 803
rect 13756 793 13776 801
rect 13789 800 13792 801
rect 13790 793 13792 800
rect 13796 799 13804 803
rect 13808 799 13830 803
rect 13810 794 13830 799
rect 13868 798 13876 810
rect 13880 800 13882 830
rect 13899 826 13901 840
rect 13941 838 13947 844
rect 13999 838 14005 844
rect 14038 841 14043 845
rect 14331 841 14336 845
rect 14330 832 14338 841
rect 14342 834 14344 839
rect 14374 834 14376 846
rect 14634 845 14636 865
rect 14668 863 14670 872
rect 14705 863 14706 872
rect 14824 868 14841 881
rect 14869 868 14874 872
rect 14824 866 14833 868
rect 14824 865 14832 866
rect 14858 865 14866 866
rect 14667 857 14668 862
rect 14665 849 14666 855
rect 14386 844 14394 845
rect 14342 832 14376 834
rect 14380 832 14394 844
rect 13914 826 13915 832
rect 14386 830 14394 832
rect 14025 829 14028 830
rect 14001 827 14036 829
rect 13899 818 13900 826
rect 13997 825 14001 827
rect 13900 800 13903 814
rect 13915 812 13917 825
rect 13968 808 13997 825
rect 13999 814 14001 817
rect 14009 812 14025 827
rect 14004 811 14025 812
rect 14036 824 14196 827
rect 13880 798 13914 800
rect 13900 795 13903 798
rect 13658 778 13661 788
rect 13661 769 13663 778
rect 13664 774 13679 790
rect 13716 774 13730 790
rect 13753 781 13754 788
rect 13663 765 13664 769
rect 13480 762 13505 763
rect 13534 762 13537 763
rect 13480 760 13537 762
rect 13480 758 13496 760
rect 13664 759 13665 763
rect 11604 749 11640 750
rect 11623 744 11635 749
rect 11690 744 11701 749
rect 13158 746 13161 754
rect 13189 748 13194 754
rect 13194 745 13198 748
rect 13388 745 13390 757
rect 13393 745 13427 757
rect 13432 756 13434 757
rect 13541 756 13568 759
rect 13665 757 13666 759
rect 13680 758 13696 772
rect 13698 758 13714 772
rect 13746 769 13754 781
rect 13758 774 13776 793
rect 13810 792 13826 794
rect 13810 774 13826 790
rect 13856 774 13871 790
rect 13873 775 13875 789
rect 13880 786 13892 794
rect 13902 786 13914 794
rect 13916 790 13917 808
rect 14003 805 14013 811
rect 14036 808 14202 824
rect 14264 808 14280 824
rect 14282 808 14298 824
rect 14342 820 14354 828
rect 14364 820 14376 828
rect 14342 810 14344 820
rect 14394 816 14398 830
rect 14420 828 14422 845
rect 14422 819 14423 828
rect 14450 819 14453 845
rect 14455 843 14504 845
rect 14539 843 14541 844
rect 14455 833 14497 843
rect 14575 838 14576 843
rect 14542 827 14543 836
rect 14576 827 14577 836
rect 14633 834 14634 844
rect 14664 843 14665 847
rect 14663 837 14664 843
rect 14492 811 14497 823
rect 14544 817 14545 820
rect 14577 816 14578 820
rect 14632 819 14633 832
rect 14661 827 14663 836
rect 14703 829 14705 862
rect 14816 855 14832 865
rect 14869 864 14873 868
rect 14753 845 14816 855
rect 14861 851 14869 864
rect 14744 844 14753 845
rect 14738 842 14744 844
rect 14728 834 14738 842
rect 14660 821 14661 826
rect 14701 820 14703 827
rect 14545 811 14546 814
rect 14578 811 14579 814
rect 14631 811 14632 818
rect 14645 811 14651 817
rect 14659 816 14660 820
rect 14700 818 14701 820
rect 14708 818 14728 834
rect 14658 814 14659 816
rect 14657 812 14658 814
rect 14691 811 14697 817
rect 14699 813 14708 818
rect 14698 811 14708 813
rect 14454 808 14455 810
rect 14546 808 14547 810
rect 14008 803 14013 805
rect 14133 803 14142 808
rect 14180 803 14189 808
rect 13920 802 13929 803
rect 13918 798 13926 802
rect 13929 799 13944 802
rect 13944 798 13947 799
rect 13941 792 13947 798
rect 13999 792 14005 798
rect 14013 794 14022 803
rect 14124 794 14133 803
rect 14189 794 14198 803
rect 14115 792 14122 793
rect 13947 790 13953 792
rect 13758 772 13792 774
rect 13805 772 13810 774
rect 13903 772 13906 786
rect 13916 774 13922 790
rect 13947 786 13968 790
rect 13993 786 13999 792
rect 14109 791 14115 792
rect 14166 791 14170 793
rect 14202 792 14218 808
rect 14248 792 14264 808
rect 14275 803 14281 808
rect 14275 802 14290 803
rect 14269 796 14275 802
rect 14298 798 14314 808
rect 14321 802 14327 808
rect 14274 791 14275 793
rect 14307 791 14312 798
rect 14327 796 14333 802
rect 14345 800 14346 808
rect 14107 790 14109 791
rect 14106 787 14107 790
rect 14171 789 14173 790
rect 13952 774 13968 786
rect 14019 778 14046 781
rect 14002 774 14019 778
rect 14046 774 14054 778
rect 13758 769 13810 772
rect 13871 769 13877 772
rect 13906 771 13910 772
rect 13758 757 13762 765
rect 13794 758 13810 769
rect 13872 762 13889 769
rect 13906 762 13916 771
rect 13872 758 13888 762
rect 13889 760 13894 762
rect 13898 760 13910 762
rect 13894 759 13910 760
rect 13890 758 13910 759
rect 13968 758 13984 774
rect 14054 772 14057 774
rect 14122 772 14128 778
rect 14131 772 14133 779
rect 14173 772 14174 778
rect 14202 774 14218 790
rect 14248 774 14264 790
rect 14266 779 14275 791
rect 14057 763 14077 772
rect 14106 767 14107 769
rect 14116 766 14122 772
rect 14174 766 14180 772
rect 14195 763 14202 774
rect 14077 762 14079 763
rect 14079 759 14085 762
rect 13434 751 13455 756
rect 13455 747 13471 751
rect 13503 748 13515 756
rect 13666 754 13667 756
rect 13562 747 13568 753
rect 13593 747 13648 753
rect 13667 750 13668 754
rect 13668 747 13670 748
rect 13677 747 13686 756
rect 13756 747 13762 756
rect 13814 747 13820 753
rect 13821 747 13830 756
rect 13875 751 13878 758
rect 11701 743 11703 744
rect 11187 739 11196 742
rect 11273 741 11275 742
rect 11575 741 11576 743
rect 13161 741 13163 745
rect 11018 738 11032 739
rect 11005 737 11018 738
rect 11025 735 11027 738
rect 11196 735 11207 739
rect 11250 737 11251 739
rect 11207 734 11210 735
rect 10816 733 10898 734
rect 10766 732 10832 733
rect 10809 731 10832 732
rect 10555 726 10567 731
rect 10809 729 10816 731
rect 10820 730 10832 731
rect 10898 729 10901 732
rect 11017 731 11024 734
rect 11210 731 11219 734
rect 11247 733 11249 736
rect 11219 729 11226 731
rect 11242 729 11246 731
rect 10805 728 10809 729
rect 10798 726 10805 728
rect 10835 727 10836 729
rect 10901 728 10903 729
rect 10257 721 10328 723
rect 10081 719 10096 720
rect 10258 719 10328 721
rect 10360 719 10364 725
rect 10471 723 10473 726
rect 10084 716 10096 719
rect 8323 705 8330 712
rect 8409 706 8419 709
rect 8420 706 8432 715
rect 8455 714 8457 715
rect 8457 709 8497 714
rect 8519 709 8531 714
rect 10020 712 10025 716
rect 10097 714 10100 716
rect 10249 712 10257 719
rect 10259 717 10269 719
rect 10293 717 10348 719
rect 10259 712 10263 717
rect 8497 707 8531 709
rect 8497 706 8545 707
rect 8567 706 8573 712
rect 8625 706 8631 712
rect 7994 698 8005 701
rect 8088 698 8096 701
rect 8116 700 8124 701
rect 7457 688 7458 692
rect 7420 676 7454 678
rect 7458 676 7466 688
rect 7553 686 7559 692
rect 7611 686 7617 692
rect 7643 688 7650 692
rect 7759 691 7765 697
rect 7805 691 7811 697
rect 7851 691 7994 698
rect 8066 691 8088 698
rect 8122 692 8124 700
rect 8125 693 8131 698
rect 8144 694 8156 701
rect 7746 688 7748 691
rect 7643 687 7655 688
rect 7559 680 7565 686
rect 7605 680 7611 686
rect 7643 685 7658 687
rect 7665 685 7677 688
rect 7745 687 7746 688
rect 7744 685 7745 687
rect 7753 685 7759 691
rect 7811 685 7817 691
rect 7818 689 7839 691
rect 8061 689 8066 691
rect 8055 687 8061 689
rect 8124 688 8125 692
rect 8133 689 8136 691
rect 7822 685 7857 687
rect 7643 680 7655 685
rect 7658 680 7680 685
rect 7742 683 7744 685
rect 7680 678 7686 680
rect 7686 676 7693 678
rect 7693 675 7698 676
rect 7707 675 7757 683
rect 7810 682 7822 685
rect 7801 680 7810 682
rect 7862 680 7864 685
rect 8045 684 8053 687
rect 8125 686 8126 687
rect 8038 682 8045 684
rect 8031 679 8038 682
rect 8126 680 8128 682
rect 8026 678 8031 679
rect 8128 678 8129 680
rect 8142 678 8149 684
rect 8161 682 8219 701
rect 8246 692 8247 698
rect 8310 692 8311 701
rect 8315 693 8323 703
rect 8330 702 8334 705
rect 8395 702 8420 706
rect 8517 704 8530 706
rect 8318 691 8323 693
rect 8334 692 8345 702
rect 8161 678 8194 682
rect 8219 678 8223 682
rect 8248 679 8249 682
rect 7800 676 7801 678
rect 8020 676 8026 678
rect 8129 676 8130 678
rect 7456 672 7458 675
rect 7698 674 7757 675
rect 7707 672 7757 674
rect 7163 656 7166 662
rect 7087 643 7151 649
rect 7161 648 7163 656
rect 7207 652 7224 672
rect 7247 666 7254 672
rect 7420 666 7432 672
rect 7442 666 7454 672
rect 7684 666 7707 672
rect 7254 664 7460 666
rect 7673 664 7684 666
rect 7093 637 7120 643
rect 7139 637 7145 643
rect 7155 642 7161 647
rect 7165 642 7174 644
rect 7224 643 7232 652
rect 7401 642 7402 660
rect 6082 623 6109 629
rect 6903 626 6906 630
rect 7096 626 7120 637
rect 7155 635 7174 642
rect 7233 639 7237 642
rect 7237 636 7242 639
rect 7242 635 7250 636
rect 7155 630 7170 635
rect 7250 631 7286 635
rect 7154 626 7170 630
rect 7286 628 7306 631
rect 7400 630 7402 642
rect 7460 654 7619 664
rect 7631 654 7673 664
rect 7797 663 7800 674
rect 7864 663 7867 676
rect 8015 674 8020 676
rect 8012 673 8015 674
rect 8007 672 8012 673
rect 8001 670 8007 672
rect 8130 670 8133 676
rect 8149 671 8157 678
rect 8194 671 8202 678
rect 8223 676 8225 678
rect 8250 677 8251 687
rect 8302 681 8315 682
rect 8302 679 8311 681
rect 8345 679 8350 692
rect 8395 688 8444 702
rect 8469 698 8515 704
rect 8533 703 8535 706
rect 8545 704 8565 706
rect 8573 704 8592 706
rect 8516 700 8531 702
rect 8461 694 8469 698
rect 8395 687 8420 688
rect 8444 687 8450 688
rect 8452 687 8461 694
rect 8377 678 8395 687
rect 8444 686 8452 687
rect 8450 685 8454 686
rect 8440 677 8447 683
rect 8454 682 8462 685
rect 8462 681 8467 682
rect 8467 680 8472 681
rect 8473 678 8476 679
rect 8244 676 8265 677
rect 8302 676 8308 677
rect 8225 673 8229 676
rect 7982 668 8001 670
rect 7945 664 7982 668
rect 7868 663 7945 664
rect 7759 655 7945 663
rect 8133 660 8146 670
rect 8157 660 8179 671
rect 8202 663 8212 671
rect 8229 663 8233 673
rect 8244 671 8250 676
rect 8251 672 8265 676
rect 8291 671 8308 676
rect 8349 671 8350 676
rect 8360 671 8375 677
rect 8250 665 8256 671
rect 8296 665 8302 671
rect 8340 663 8360 671
rect 8431 669 8440 677
rect 8479 676 8484 678
rect 8485 674 8491 676
rect 7460 652 7631 654
rect 7759 653 7874 655
rect 7460 642 7462 652
rect 7759 651 7871 653
rect 7759 649 7864 651
rect 7759 648 7827 649
rect 7759 645 7811 648
rect 7753 644 7817 645
rect 7731 642 7817 644
rect 7460 634 7466 642
rect 7725 639 7742 642
rect 7753 639 7817 642
rect 7850 641 7862 649
rect 7867 643 7871 651
rect 7707 636 7725 639
rect 7461 630 7466 634
rect 7688 633 7707 636
rect 7759 633 7765 639
rect 7791 636 7797 639
rect 7805 633 7811 639
rect 7869 636 7871 643
rect 8146 642 8192 660
rect 8212 652 8242 663
rect 8222 647 8256 652
rect 8276 647 8277 660
rect 8313 652 8340 663
rect 8349 660 8350 663
rect 8222 646 8293 647
rect 8301 646 8330 652
rect 8222 643 8330 646
rect 8228 642 8233 643
rect 8146 641 8194 642
rect 7673 631 7688 633
rect 7477 630 7517 631
rect 7671 630 7673 631
rect 7316 628 7477 630
rect 7517 628 7546 630
rect 7400 626 7403 628
rect 7459 626 7466 628
rect 6110 623 6137 624
rect 5494 621 5495 622
rect 5398 615 5415 621
rect 5490 616 5494 621
rect 6906 618 6914 626
rect 6974 618 6981 625
rect 6914 617 6974 618
rect 5487 615 5490 616
rect 5415 611 5487 615
rect 7138 610 7154 626
rect 7403 615 7409 626
rect 7456 618 7459 625
rect 7546 622 7607 628
rect 7617 622 7667 630
rect 7867 627 7869 636
rect 7448 615 7456 618
rect 7409 613 7450 615
rect 7791 613 7804 624
rect 7845 616 7867 627
rect 8146 626 8192 641
rect 8196 637 8199 639
rect 8199 636 8201 637
rect 8201 633 8208 636
rect 8228 634 8242 642
rect 8276 634 8277 643
rect 8348 637 8349 653
rect 8390 652 8431 669
rect 8485 668 8493 674
rect 8497 670 8499 672
rect 8529 670 8531 700
rect 8535 690 8543 702
rect 8573 700 8579 704
rect 8619 700 8625 706
rect 8643 693 8654 702
rect 10025 696 10046 712
rect 10090 710 10114 712
rect 10094 705 10114 710
rect 10249 707 10259 712
rect 10256 705 10259 707
rect 10046 695 10048 696
rect 8497 668 8531 670
rect 8535 668 8543 680
rect 8654 678 8657 692
rect 10052 689 10053 692
rect 10050 678 10057 687
rect 10094 680 10096 705
rect 10100 700 10108 705
rect 10114 699 10120 705
rect 10254 701 10256 705
rect 10248 699 10256 701
rect 10120 694 10126 699
rect 10248 695 10254 699
rect 10126 692 10129 694
rect 10062 678 10096 680
rect 10100 678 10108 690
rect 10129 688 10130 692
rect 10242 689 10248 695
rect 10252 692 10253 694
rect 10251 688 10252 691
rect 10261 689 10263 712
rect 10293 712 10303 717
rect 10309 715 10348 717
rect 10324 713 10348 715
rect 10368 713 10369 715
rect 10293 701 10295 712
rect 10303 701 10316 712
rect 10329 708 10348 713
rect 10369 708 10373 713
rect 10473 710 10480 723
rect 10567 722 10597 726
rect 10816 724 10832 726
rect 10567 714 10609 722
rect 10336 701 10348 708
rect 10373 706 10374 708
rect 10480 705 10483 710
rect 10561 709 10610 710
rect 10293 695 10300 701
rect 10293 693 10306 695
rect 10293 689 10295 693
rect 10300 689 10306 693
rect 10311 691 10320 700
rect 10339 696 10348 701
rect 10379 696 10382 701
rect 10342 691 10348 696
rect 10250 685 10251 687
rect 10294 685 10295 689
rect 10312 687 10329 691
rect 10345 689 10348 691
rect 10382 689 10388 696
rect 10483 695 10520 705
rect 10561 702 10575 709
rect 10591 708 10610 709
rect 10607 703 10610 708
rect 10560 699 10561 701
rect 10520 693 10526 695
rect 10558 694 10560 699
rect 10526 692 10531 693
rect 10557 692 10558 694
rect 10347 687 10348 689
rect 10313 686 10329 687
rect 10388 686 10390 689
rect 10531 688 10547 692
rect 10547 687 10549 688
rect 10130 680 10132 685
rect 10249 680 10250 685
rect 10315 682 10318 686
rect 10320 682 10329 686
rect 10321 680 10322 682
rect 8657 676 8658 678
rect 10057 676 10058 678
rect 10061 676 10062 678
rect 10248 676 10249 678
rect 10322 677 10323 678
rect 8493 664 8496 666
rect 8497 656 8509 664
rect 8519 656 8531 664
rect 8658 661 8661 676
rect 8375 646 8390 652
rect 8497 648 8506 656
rect 8660 648 8661 661
rect 10057 660 10061 676
rect 10097 674 10100 676
rect 10062 666 10074 674
rect 10084 666 10096 674
rect 10132 660 10136 676
rect 10056 654 10057 658
rect 10136 657 10137 660
rect 8361 641 8373 646
rect 8352 637 8361 641
rect 8208 631 8214 633
rect 8226 630 8242 634
rect 8217 626 8242 630
rect 8276 626 8278 630
rect 8210 622 8235 626
rect 7805 613 7845 616
rect 7416 610 7432 613
rect 7434 610 7450 613
rect 8210 610 8226 622
rect 8235 619 8243 622
rect 8243 618 8252 619
rect 8278 615 8283 626
rect 8310 620 8352 637
rect 8307 619 8310 620
rect 8301 618 8307 619
rect 8339 618 8346 620
rect 8335 615 8339 618
rect 8283 611 8304 615
rect 8326 611 8335 615
rect 8476 606 8500 629
rect 8506 626 8545 648
rect 8545 621 8554 626
rect 8651 622 8660 643
rect 10056 630 10058 654
rect 10136 630 10137 654
rect 10248 649 10300 663
rect 10321 662 10323 675
rect 10350 672 10362 685
rect 10390 672 10402 686
rect 10552 685 10558 687
rect 10558 683 10566 685
rect 10563 681 10567 683
rect 10563 676 10570 681
rect 10607 678 10609 703
rect 10610 697 10611 702
rect 10613 698 10621 710
rect 10766 694 10794 695
rect 10830 694 10832 724
rect 10836 714 10844 726
rect 10903 712 10905 728
rect 11226 727 11232 729
rect 11239 727 11242 729
rect 10959 720 10965 726
rect 11017 720 11023 726
rect 11223 723 11243 727
rect 11275 723 11296 741
rect 11301 738 11312 740
rect 11223 721 11239 723
rect 11218 720 11223 721
rect 11243 720 11251 723
rect 10965 714 10971 720
rect 11011 714 11017 720
rect 11211 717 11218 720
rect 11251 719 11254 720
rect 11296 719 11301 723
rect 11206 716 11211 717
rect 11254 716 11260 719
rect 11301 716 11305 719
rect 11309 716 11311 738
rect 11312 737 11313 738
rect 11315 737 11323 740
rect 11313 734 11323 737
rect 11315 728 11323 734
rect 11402 733 11403 741
rect 11439 737 11442 741
rect 11403 729 11404 733
rect 11432 729 11444 737
rect 11454 729 11466 737
rect 11529 729 11542 741
rect 11321 726 11324 728
rect 11324 719 11331 726
rect 11404 724 11411 729
rect 11428 727 11431 729
rect 11444 725 11445 729
rect 11451 725 11457 729
rect 11405 723 11411 724
rect 11420 723 11428 725
rect 11432 723 11478 725
rect 11315 716 11323 718
rect 11197 713 11206 716
rect 11192 711 11197 713
rect 10611 693 10612 694
rect 10786 692 10794 694
rect 10798 692 10832 694
rect 10836 692 10844 704
rect 10903 694 10905 710
rect 11176 706 11192 711
rect 11260 706 11271 716
rect 11305 707 11323 716
rect 11331 712 11339 719
rect 11399 717 11405 723
rect 11432 717 11434 723
rect 11457 717 11463 723
rect 11464 719 11478 723
rect 11403 713 11405 714
rect 11287 706 11323 707
rect 11339 706 11347 712
rect 11401 709 11403 713
rect 11160 701 11176 706
rect 11271 705 11278 706
rect 11316 705 11349 706
rect 11271 702 11279 705
rect 11253 701 11287 702
rect 11313 701 11374 705
rect 11464 702 11466 719
rect 11470 713 11478 719
rect 11473 712 11478 713
rect 11542 712 11561 729
rect 11576 715 11610 741
rect 11705 723 11728 741
rect 13198 740 13206 745
rect 13424 742 13425 745
rect 13471 742 13491 747
rect 13491 741 13496 742
rect 13568 741 13574 747
rect 13614 741 13620 747
rect 13390 740 13392 741
rect 13163 737 13165 740
rect 13206 737 13211 740
rect 13380 739 13390 740
rect 13369 738 13390 739
rect 13496 738 13500 741
rect 13621 738 13630 747
rect 13668 745 13677 747
rect 13668 742 13683 745
rect 13668 738 13677 742
rect 13683 740 13687 742
rect 13762 741 13774 747
rect 13808 741 13821 747
rect 13877 744 13878 751
rect 13687 739 13690 740
rect 13211 736 13213 737
rect 13378 736 13397 738
rect 13166 733 13167 736
rect 13213 733 13217 736
rect 13167 727 13170 733
rect 13217 731 13221 733
rect 13221 729 13224 731
rect 13311 729 13317 735
rect 13369 729 13375 735
rect 13378 733 13415 736
rect 13422 733 13423 736
rect 13389 729 13415 733
rect 13418 729 13422 731
rect 13454 729 13455 730
rect 13224 726 13228 729
rect 13170 720 13174 726
rect 13228 720 13238 726
rect 13241 720 13253 724
rect 13317 723 13323 729
rect 13363 723 13369 729
rect 13415 726 13455 729
rect 13415 723 13454 726
rect 13500 725 13517 738
rect 13621 737 13622 738
rect 13690 736 13697 739
rect 13765 738 13774 741
rect 13812 738 13821 741
rect 13871 739 13878 744
rect 13906 742 13910 758
rect 13948 747 13957 756
rect 14013 747 14022 756
rect 14085 754 14096 759
rect 14189 758 14202 763
rect 14264 769 14273 774
rect 14274 769 14275 779
rect 14264 763 14275 769
rect 14278 763 14280 791
rect 14346 790 14348 791
rect 14344 785 14348 790
rect 14397 790 14398 808
rect 14504 799 14516 804
rect 14548 796 14549 799
rect 14579 796 14580 805
rect 14630 799 14631 808
rect 14639 805 14645 811
rect 14697 808 14703 811
rect 14752 808 14768 824
rect 15341 819 15342 1015
rect 15531 819 15532 1015
rect 15617 819 15618 1015
rect 15890 819 15891 1015
rect 16087 819 16088 1015
rect 16480 1014 16484 1019
rect 17118 1014 17125 1019
rect 17205 1018 17214 1027
rect 17270 1024 17366 1027
rect 17707 1023 17815 1037
rect 17565 1015 17581 1022
rect 17583 1015 17599 1022
rect 17125 1007 17137 1014
rect 17555 1013 17567 1015
rect 17577 1013 17589 1015
rect 17595 1013 17599 1015
rect 17783 1013 17799 1022
rect 17815 1021 17833 1023
rect 17834 1017 17841 1020
rect 17841 1013 17847 1017
rect 18487 1015 18488 1026
rect 18677 1015 18678 1026
rect 18763 1015 18764 1026
rect 19036 1015 19037 1026
rect 19233 1015 19234 1026
rect 17555 1008 17599 1013
rect 17742 1008 17779 1009
rect 17847 1008 17850 1013
rect 17551 1006 17553 1008
rect 17555 1006 17687 1008
rect 16606 1005 16960 1006
rect 16586 1003 16604 1005
rect 17046 1003 17059 1005
rect 17138 1003 17141 1005
rect 17549 1003 17687 1006
rect 16530 1000 16586 1003
rect 16404 992 16416 1000
rect 16426 992 16438 1000
rect 16502 994 16586 1000
rect 17059 994 17069 1003
rect 16502 993 16530 994
rect 16400 989 16402 992
rect 16502 991 16521 993
rect 17070 991 17073 993
rect 16442 988 16446 989
rect 16392 977 16400 988
rect 16403 986 16438 988
rect 16401 977 16403 983
rect 16392 976 16401 977
rect 16400 972 16401 976
rect 16399 971 16400 972
rect 16397 966 16399 969
rect 16272 964 16337 965
rect 16264 956 16272 964
rect 16337 956 16341 964
rect 16263 950 16264 956
rect 16392 954 16400 966
rect 16404 956 16406 986
rect 16435 985 16438 986
rect 16437 979 16438 985
rect 16442 981 16450 988
rect 16446 980 16454 981
rect 16478 980 16479 990
rect 16502 980 16517 991
rect 16776 981 16813 983
rect 16454 979 16460 980
rect 16477 979 16478 980
rect 16502 979 16509 980
rect 16460 969 16522 979
rect 16530 972 16536 978
rect 16576 972 16582 978
rect 16776 977 16802 981
rect 16813 977 16818 981
rect 17073 980 17086 991
rect 17049 979 17063 980
rect 16770 972 16776 977
rect 16818 972 16827 977
rect 17031 972 17049 979
rect 17063 977 17070 979
rect 17141 977 17162 1003
rect 17543 996 17687 1003
rect 17703 1006 17804 1008
rect 17703 996 17815 1006
rect 17504 990 17565 996
rect 17469 987 17504 990
rect 17282 981 17469 987
rect 17555 986 17565 990
rect 17070 972 17085 977
rect 16524 969 16530 972
rect 16531 970 16588 972
rect 16827 971 16828 972
rect 16665 970 16668 971
rect 16686 970 16689 971
rect 16768 970 16769 971
rect 16828 970 16831 971
rect 16531 969 16539 970
rect 16502 968 16539 969
rect 16404 954 16438 956
rect 16393 951 16395 954
rect 16389 938 16393 950
rect 16404 942 16416 950
rect 16429 945 16438 954
rect 16476 952 16477 955
rect 16502 951 16507 968
rect 16524 966 16539 968
rect 16582 966 16588 970
rect 16661 967 16665 970
rect 16689 967 16694 970
rect 16831 968 16832 970
rect 17023 969 17031 972
rect 17060 971 17085 972
rect 17094 971 17098 972
rect 17056 970 17060 971
rect 17070 970 17107 971
rect 16832 967 16835 968
rect 16530 964 16539 966
rect 16530 951 16535 964
rect 16583 955 16602 958
rect 16637 955 16661 967
rect 16694 959 16712 967
rect 16767 959 16768 967
rect 16439 949 16444 950
rect 16444 948 16449 949
rect 16449 947 16452 948
rect 16454 945 16463 947
rect 16427 942 16429 945
rect 16463 944 16468 945
rect 16468 943 16474 944
rect 16475 943 16476 951
rect 16502 943 16508 951
rect 16426 939 16427 942
rect 16474 938 16508 943
rect 16387 931 16389 937
rect 16424 930 16426 938
rect 16475 932 16476 938
rect 16502 935 16530 938
rect 16502 933 16532 935
rect 16502 931 16533 933
rect 16534 931 16535 951
rect 16602 946 16664 955
rect 16712 952 16720 959
rect 16766 951 16767 958
rect 16835 954 16839 967
rect 17015 966 17023 969
rect 17053 968 17056 970
rect 17049 967 17053 968
rect 17044 965 17049 967
rect 17070 965 17085 970
rect 17094 969 17098 970
rect 17107 969 17108 970
rect 17164 969 17169 975
rect 17205 971 17214 980
rect 17270 978 17282 981
rect 17270 971 17279 978
rect 17549 972 17565 986
rect 17588 972 17589 996
rect 17594 991 17615 996
rect 17599 990 17615 991
rect 17732 989 17738 996
rect 17784 989 17790 996
rect 17804 990 17815 996
rect 17850 990 17859 1008
rect 17599 972 17615 988
rect 17732 985 17740 989
rect 17738 983 17740 985
rect 17648 974 17676 978
rect 17678 974 17689 978
rect 17098 965 17103 969
rect 17108 965 17110 968
rect 17169 965 17172 969
rect 17010 964 17014 965
rect 17085 964 17088 965
rect 17110 964 17111 965
rect 17006 962 17010 964
rect 16620 945 16630 946
rect 16652 945 16653 946
rect 16616 943 16620 945
rect 16664 943 16684 946
rect 16765 943 16766 950
rect 16838 943 16839 950
rect 16973 949 17006 962
rect 17090 959 17094 962
rect 17105 960 17109 963
rect 17214 962 17223 971
rect 17247 961 17250 963
rect 17261 962 17270 971
rect 17555 970 17589 972
rect 17598 971 17599 972
rect 17645 971 17648 974
rect 17594 970 17599 971
rect 17644 970 17645 971
rect 17555 968 17599 970
rect 17642 969 17644 970
rect 17551 965 17552 967
rect 17325 961 17334 963
rect 17242 959 17247 961
rect 16887 943 16893 949
rect 16933 948 16939 949
rect 16970 948 16973 949
rect 16933 947 16970 948
rect 16933 943 16939 947
rect 17025 946 17031 952
rect 17071 946 17077 952
rect 17093 949 17094 959
rect 17240 958 17242 959
rect 17336 958 17342 961
rect 17111 955 17115 958
rect 17179 955 17181 958
rect 17115 946 17125 955
rect 16604 931 16612 943
rect 16616 941 16650 943
rect 16340 924 16341 929
rect 16290 915 16299 924
rect 16337 920 16346 924
rect 16337 915 16351 920
rect 16281 912 16290 915
rect 16281 911 16284 912
rect 16274 908 16283 911
rect 16262 907 16283 908
rect 16262 905 16280 907
rect 16320 905 16326 911
rect 16340 906 16355 915
rect 16380 908 16387 929
rect 16262 900 16274 905
rect 16258 898 16261 900
rect 16262 899 16263 900
rect 16268 899 16274 900
rect 16326 899 16332 905
rect 16339 904 16351 906
rect 16378 904 16380 908
rect 16418 907 16424 929
rect 16475 926 16476 929
rect 16502 928 16563 931
rect 16502 917 16508 928
rect 16530 926 16563 928
rect 16524 925 16563 926
rect 16582 925 16588 926
rect 16524 921 16588 925
rect 16524 920 16610 921
rect 16502 913 16511 917
rect 16530 914 16536 920
rect 16576 914 16582 920
rect 16585 917 16610 920
rect 16594 913 16610 917
rect 16616 913 16618 941
rect 16647 939 16650 941
rect 16502 909 16517 913
rect 16604 909 16618 913
rect 16648 909 16650 939
rect 16654 931 16662 943
rect 16684 934 16747 943
rect 16881 938 16887 943
rect 16899 941 16935 943
rect 16899 938 16904 941
rect 16840 937 16887 938
rect 16901 937 16904 938
rect 16939 937 16945 943
rect 17019 940 17025 946
rect 17077 940 17083 946
rect 16840 936 16883 937
rect 16764 934 16765 936
rect 16786 934 16840 936
rect 16720 922 16735 934
rect 16747 933 16786 934
rect 16764 929 16765 933
rect 16896 929 16899 936
rect 17023 933 17025 934
rect 17021 929 17023 933
rect 16417 904 16418 906
rect 16477 905 16478 909
rect 16337 899 16339 904
rect 16483 903 16489 909
rect 16502 903 16521 909
rect 16529 903 16535 909
rect 16377 899 16378 903
rect 16336 897 16337 899
rect 16376 897 16377 899
rect 16250 884 16258 896
rect 16262 894 16280 896
rect 16335 895 16336 896
rect 16415 895 16417 903
rect 16477 897 16483 903
rect 16502 897 16541 903
rect 16543 897 16555 905
rect 16616 904 16633 909
rect 16624 899 16631 904
rect 16633 903 16637 904
rect 16653 903 16654 905
rect 16720 904 16735 920
rect 16762 906 16764 928
rect 16637 900 16656 903
rect 16761 900 16773 905
rect 16783 900 16795 905
rect 16836 904 16838 928
rect 16887 904 16896 928
rect 16932 904 16935 909
rect 16973 908 17008 910
rect 17019 908 17021 929
rect 17043 909 17044 929
rect 17091 928 17093 944
rect 17125 942 17130 946
rect 17181 942 17193 955
rect 17342 951 17355 958
rect 17565 956 17581 968
rect 17583 956 17599 968
rect 17638 965 17642 968
rect 17636 963 17638 965
rect 17634 961 17636 963
rect 17689 961 17702 974
rect 17738 967 17741 983
rect 17740 961 17741 967
rect 17744 967 17745 989
rect 17783 985 17790 989
rect 17811 987 17813 990
rect 17783 983 17784 985
rect 17804 984 17805 986
rect 17744 963 17746 967
rect 17777 963 17778 966
rect 17782 965 17784 983
rect 17813 981 17816 987
rect 17816 979 17817 981
rect 17818 975 17819 977
rect 17819 972 17820 975
rect 17859 973 17867 990
rect 17821 965 17824 969
rect 17744 961 17748 963
rect 17782 962 17783 965
rect 17824 963 17825 965
rect 17630 958 17633 961
rect 17702 959 17705 961
rect 17628 953 17630 958
rect 17705 957 17707 959
rect 17463 952 17500 953
rect 17627 952 17628 953
rect 17707 952 17709 957
rect 17735 955 17741 961
rect 17748 959 17754 961
rect 17755 957 17761 959
rect 17781 957 17787 961
rect 17825 960 17826 963
rect 17826 958 17827 960
rect 17761 956 17787 957
rect 17463 951 17488 952
rect 17500 951 17501 952
rect 17357 948 17361 951
rect 17428 948 17455 951
rect 17503 948 17510 951
rect 17555 949 17556 952
rect 17626 951 17627 952
rect 17510 943 17521 948
rect 17556 945 17558 949
rect 17591 947 17592 949
rect 17624 948 17626 951
rect 17521 942 17525 943
rect 17193 939 17194 942
rect 17525 938 17532 942
rect 17135 929 17145 938
rect 17195 931 17201 938
rect 17532 937 17534 938
rect 17534 933 17550 937
rect 17550 932 17555 933
rect 17558 932 17566 944
rect 17555 929 17566 932
rect 17592 929 17596 944
rect 17622 943 17624 948
rect 17709 944 17712 951
rect 17729 949 17735 955
rect 17761 951 17805 956
rect 17827 955 17829 958
rect 17787 949 17793 951
rect 17829 948 17832 955
rect 17621 942 17622 943
rect 17832 942 17835 948
rect 17867 943 17868 973
rect 17975 951 17991 954
rect 17903 943 17926 951
rect 17981 943 17998 951
rect 17620 940 17621 942
rect 17619 939 17620 940
rect 17835 939 17836 942
rect 17618 937 17619 938
rect 17615 933 17618 937
rect 17613 932 17615 933
rect 17611 929 17613 932
rect 17836 931 17837 938
rect 17866 929 17867 942
rect 17895 938 17903 943
rect 17981 938 18005 943
rect 17885 932 17895 938
rect 17878 929 17885 932
rect 17088 917 17090 920
rect 17084 914 17087 916
rect 17082 913 17084 914
rect 17079 911 17082 913
rect 17077 910 17079 911
rect 16963 906 16973 908
rect 17008 906 17025 908
rect 16952 904 16963 906
rect 16886 900 16887 903
rect 16930 900 16932 904
rect 16944 902 16952 904
rect 16940 901 16944 902
rect 17019 900 17021 906
rect 17043 904 17044 906
rect 17111 904 17127 920
rect 17145 910 17167 929
rect 17205 920 17213 927
rect 17213 918 17220 920
rect 17220 914 17236 918
rect 17239 914 17240 929
rect 17558 928 17571 929
rect 17564 927 17571 928
rect 17596 927 17597 928
rect 17610 927 17611 929
rect 17734 927 17735 929
rect 17566 923 17567 926
rect 17571 924 17608 927
rect 17298 921 17329 922
rect 17289 920 17298 921
rect 17329 920 17336 921
rect 17596 920 17597 924
rect 17260 917 17289 920
rect 17336 917 17351 920
rect 17258 916 17260 917
rect 17251 914 17258 916
rect 17351 914 17363 917
rect 17568 915 17569 917
rect 17597 915 17598 920
rect 17602 915 17611 924
rect 17649 915 17658 924
rect 17733 922 17734 927
rect 17732 920 17733 922
rect 17731 918 17732 920
rect 17730 916 17731 918
rect 17593 914 17602 915
rect 17236 911 17602 914
rect 17239 910 17240 911
rect 17242 910 17244 911
rect 17378 910 17386 911
rect 17167 909 17169 910
rect 17044 900 17048 904
rect 17098 900 17111 904
rect 17169 903 17177 909
rect 17238 908 17242 910
rect 17386 906 17404 910
rect 17569 906 17570 909
rect 17599 906 17600 909
rect 17231 904 17236 906
rect 16502 895 16557 897
rect 16631 895 16637 899
rect 16651 898 16652 900
rect 16650 895 16651 897
rect 16656 896 16825 900
rect 16884 897 16886 900
rect 16881 896 16887 897
rect 16927 896 16930 900
rect 16761 895 16762 896
rect 16825 895 16887 896
rect 16250 862 16258 874
rect 16262 865 16264 894
rect 16334 893 16335 894
rect 16375 893 16376 894
rect 16502 893 16559 895
rect 16637 893 16638 895
rect 16329 889 16335 893
rect 16374 889 16375 893
rect 16414 889 16415 893
rect 16470 889 16477 893
rect 16502 892 16567 893
rect 16315 888 16335 889
rect 16315 878 16329 888
rect 16371 879 16374 889
rect 16412 878 16414 889
rect 16467 879 16470 889
rect 16299 866 16315 878
rect 16262 862 16265 865
rect 16296 862 16299 866
rect 16346 859 16355 868
rect 16367 866 16371 878
rect 16411 875 16412 878
rect 16466 875 16467 878
rect 16366 862 16367 866
rect 16261 857 16263 858
rect 16268 857 16274 859
rect 16262 853 16274 857
rect 16326 853 16332 859
rect 16338 857 16346 859
rect 16365 858 16366 862
rect 16407 859 16411 875
rect 16461 859 16466 875
rect 16479 864 16482 892
rect 16529 891 16555 892
rect 16553 861 16555 891
rect 16559 881 16567 892
rect 16638 879 16658 893
rect 16706 879 16720 894
rect 16749 881 16757 893
rect 16761 891 16795 893
rect 16614 876 16615 879
rect 16644 876 16645 879
rect 16658 877 16670 879
rect 16704 877 16706 879
rect 16658 875 16704 877
rect 16529 859 16555 861
rect 16559 859 16567 871
rect 16612 869 16614 875
rect 16642 870 16644 875
rect 16610 862 16612 869
rect 16639 862 16642 869
rect 16609 859 16610 862
rect 16638 859 16639 862
rect 16761 859 16763 891
rect 16793 875 16795 891
rect 16799 881 16807 893
rect 16881 891 16887 895
rect 16925 891 16927 895
rect 16939 891 16945 897
rect 17019 894 17025 900
rect 17048 896 17063 900
rect 17063 895 17064 896
rect 17077 895 17111 900
rect 17177 899 17183 903
rect 17228 902 17231 904
rect 17404 902 17424 906
rect 17495 902 17508 903
rect 16835 881 16836 889
rect 16879 881 16882 891
rect 16887 885 16893 891
rect 16919 881 16925 891
rect 16933 885 16939 891
rect 17022 883 17023 891
rect 17025 888 17031 894
rect 17064 893 17083 895
rect 16794 865 16795 874
rect 16799 872 16800 875
rect 16829 870 16835 880
rect 16874 870 16879 881
rect 16817 866 16829 870
rect 16873 867 16874 870
rect 16912 867 16919 881
rect 17062 872 17065 892
rect 17071 888 17077 893
rect 17095 888 17111 895
rect 17183 894 17194 899
rect 17222 898 17226 900
rect 17219 897 17222 898
rect 17216 895 17219 897
rect 17239 895 17242 900
rect 17424 897 17449 902
rect 17474 900 17492 902
rect 17513 900 17536 902
rect 17472 899 17484 900
rect 17536 899 17545 900
rect 17545 898 17546 899
rect 17570 898 17571 902
rect 17449 895 17454 897
rect 17465 895 17472 898
rect 17194 885 17225 894
rect 17242 893 17244 895
rect 17244 891 17246 893
rect 17454 891 17472 895
rect 17546 894 17553 898
rect 17600 897 17601 902
rect 17658 901 17667 915
rect 17728 911 17729 914
rect 17755 909 17787 913
rect 17722 903 17726 906
rect 17729 903 17735 909
rect 17755 904 17793 909
rect 17824 904 17878 929
rect 17981 922 18007 938
rect 17752 903 17793 904
rect 17709 901 17721 902
rect 17667 899 17671 901
rect 17689 900 17709 901
rect 17683 899 17689 900
rect 17709 895 17711 900
rect 17735 897 17741 903
rect 17769 899 17770 901
rect 17553 891 17559 894
rect 17571 891 17572 895
rect 17184 880 17225 885
rect 17246 888 17319 891
rect 17454 889 17471 891
rect 17246 885 17326 888
rect 17246 881 17319 885
rect 17326 881 17396 885
rect 17457 882 17465 889
rect 17471 887 17476 889
rect 17476 885 17480 887
rect 17559 885 17572 891
rect 17601 887 17603 895
rect 17707 892 17709 895
rect 17706 891 17707 892
rect 17184 876 17200 880
rect 17225 876 17243 880
rect 17246 876 17264 881
rect 17319 876 17424 881
rect 17243 875 17424 876
rect 17450 875 17457 882
rect 17480 876 17502 885
rect 17559 882 17573 885
rect 17572 881 17575 882
rect 17572 878 17573 881
rect 17575 880 17576 881
rect 17576 879 17585 880
rect 17603 879 17605 885
rect 17694 882 17706 891
rect 17688 881 17694 882
rect 17660 880 17676 881
rect 17684 880 17688 881
rect 17753 880 17768 899
rect 17781 897 17787 903
rect 17818 901 17824 904
rect 17832 903 17833 904
rect 17807 895 17818 901
rect 17831 899 17832 901
rect 17804 892 17807 895
rect 17803 891 17804 892
rect 17795 885 17803 891
rect 17632 879 17655 880
rect 17502 875 17505 876
rect 16911 866 16912 867
rect 16816 865 16817 866
rect 16794 862 16816 865
rect 16870 862 16873 866
rect 16795 859 16816 862
rect 16867 859 16873 862
rect 16337 855 16346 857
rect 16262 852 16271 853
rect 16262 850 16272 852
rect 16274 850 16280 853
rect 16272 847 16280 850
rect 16272 846 16274 847
rect 16274 842 16276 845
rect 16325 840 16326 853
rect 16335 852 16346 855
rect 16333 851 16335 852
rect 16330 850 16333 851
rect 16337 850 16346 852
rect 16361 845 16365 858
rect 16404 846 16407 858
rect 16457 846 16461 858
rect 16477 851 16483 857
rect 16506 856 16510 859
rect 16800 858 16801 859
rect 16483 845 16489 851
rect 16501 845 16506 856
rect 16535 851 16541 857
rect 16608 855 16609 858
rect 16637 855 16638 858
rect 16867 857 16870 859
rect 16869 856 16870 857
rect 16865 855 16869 856
rect 16529 845 16535 851
rect 16543 847 16555 855
rect 16759 853 16760 855
rect 16357 841 16361 845
rect 16403 841 16404 845
rect 16455 842 16457 845
rect 16355 840 16357 841
rect 16499 840 16501 845
rect 16603 841 16606 850
rect 16633 841 16636 850
rect 16760 841 16762 849
rect 16801 842 16802 849
rect 16862 847 16869 855
rect 16856 845 16863 847
rect 16865 845 16869 847
rect 16899 845 16911 865
rect 17023 859 17025 872
rect 16856 840 16865 845
rect 16896 844 16903 845
rect 17058 844 17062 870
rect 17173 869 17183 875
rect 17236 872 17436 875
rect 17447 872 17450 875
rect 17505 872 17515 875
rect 17521 872 17533 878
rect 17576 875 17655 879
rect 17783 876 17815 885
rect 17828 880 17831 898
rect 17827 876 17828 880
rect 17863 878 17865 904
rect 17981 895 18004 922
rect 18036 895 18037 929
rect 17981 881 18003 895
rect 18015 889 18037 895
rect 17236 871 17244 872
rect 17231 869 17235 871
rect 17171 868 17173 869
rect 17168 866 17171 868
rect 17226 866 17230 868
rect 17319 867 17543 872
rect 17573 871 17574 875
rect 17585 871 17632 875
rect 17746 872 17749 876
rect 17780 875 17815 876
rect 17591 869 17632 871
rect 17597 868 17622 869
rect 17335 866 17543 867
rect 17161 862 17168 866
rect 17216 862 17226 866
rect 17335 863 17545 866
rect 17448 862 17457 863
rect 17531 862 17553 863
rect 17574 862 17575 868
rect 17598 867 17622 868
rect 17738 863 17746 872
rect 17793 869 17794 874
rect 17155 858 17161 862
rect 17457 858 17464 862
rect 17153 857 17155 858
rect 17144 852 17153 857
rect 17464 852 17475 858
rect 17531 854 17545 862
rect 17553 856 17586 862
rect 17605 859 17606 862
rect 17734 857 17738 862
rect 17661 856 17673 857
rect 17586 855 17592 856
rect 17610 855 17632 856
rect 17592 854 17632 855
rect 17653 854 17673 856
rect 17139 850 17144 852
rect 17475 850 17479 852
rect 17104 849 17110 850
rect 17137 849 17139 850
rect 17086 844 17137 849
rect 17150 844 17156 850
rect 17200 845 17203 849
rect 17480 845 17488 849
rect 17531 846 17543 854
rect 17661 852 17693 854
rect 17576 850 17577 852
rect 17606 850 17607 852
rect 17662 847 17693 852
rect 17731 849 17733 856
rect 17731 847 17732 849
rect 16896 840 16900 844
rect 16277 836 16278 840
rect 16278 833 16279 836
rect 16325 832 16327 840
rect 16343 832 16355 840
rect 16402 838 16403 840
rect 16454 838 16455 840
rect 16401 832 16402 838
rect 16453 833 16454 838
rect 16496 832 16499 840
rect 16602 837 16603 840
rect 16601 833 16602 836
rect 16630 834 16632 840
rect 16802 837 16803 840
rect 16763 832 16767 837
rect 16854 832 16863 840
rect 16892 834 16900 840
rect 16892 832 16896 834
rect 16279 817 16287 832
rect 16325 825 16329 832
rect 16341 828 16343 832
rect 16400 828 16401 832
rect 16451 828 16452 832
rect 16327 817 16329 825
rect 16338 819 16341 828
rect 16398 819 16400 828
rect 16449 824 16451 827
rect 16445 820 16451 824
rect 16287 811 16290 817
rect 16329 811 16330 817
rect 16337 815 16338 819
rect 16397 815 16398 819
rect 16445 815 16449 820
rect 16491 819 16496 832
rect 16290 809 16291 811
rect 16336 809 16337 814
rect 16395 809 16397 814
rect 16445 809 16447 815
rect 16488 814 16491 818
rect 16541 814 16557 824
rect 16559 814 16575 824
rect 16595 817 16601 832
rect 16484 809 16488 814
rect 16528 809 16535 814
rect 16580 808 16588 814
rect 16593 811 16595 817
rect 16623 811 16630 832
rect 16764 827 16768 832
rect 16803 827 16809 832
rect 16622 809 16623 811
rect 16637 808 16653 824
rect 16753 822 16819 827
rect 16839 824 16854 832
rect 16753 821 16809 822
rect 16744 814 16753 821
rect 16764 818 16768 821
rect 16660 808 16679 809
rect 16685 808 16687 809
rect 14695 805 14703 808
rect 14695 804 14697 805
rect 14698 800 14699 802
rect 14699 797 14701 800
rect 14264 758 14280 763
rect 14329 773 14390 785
rect 14397 779 14410 790
rect 14396 774 14410 779
rect 14440 774 14455 790
rect 14456 777 14458 793
rect 14549 789 14550 793
rect 14580 789 14581 795
rect 14329 759 14394 773
rect 14360 758 14376 759
rect 14378 758 14394 759
rect 14421 758 14422 760
rect 14456 758 14472 774
rect 14550 767 14554 785
rect 14581 779 14582 788
rect 14630 787 14632 794
rect 14695 790 14696 794
rect 14701 791 14704 797
rect 14736 792 14752 808
rect 14786 802 14814 808
rect 14780 794 14814 802
rect 16293 799 16295 803
rect 16330 799 16331 803
rect 16333 800 16336 808
rect 16393 800 16395 808
rect 16295 794 16297 798
rect 16333 794 16335 800
rect 16391 794 16393 798
rect 14776 791 14778 794
rect 14786 790 14814 794
rect 14632 781 14633 787
rect 14695 782 14712 790
rect 14582 766 14587 779
rect 14634 774 14642 780
rect 14696 776 14712 782
rect 14768 779 14776 790
rect 14765 778 14776 779
rect 14780 788 14814 790
rect 14696 774 14706 776
rect 14642 773 14644 774
rect 14554 760 14555 766
rect 14587 759 14589 766
rect 14644 765 14658 773
rect 14696 766 14697 774
rect 14712 768 14717 776
rect 14765 770 14774 778
rect 14693 765 14697 766
rect 14639 764 14672 765
rect 14693 764 14703 765
rect 14639 759 14645 764
rect 14189 756 14195 758
rect 14266 757 14280 758
rect 14392 757 14395 758
rect 14274 756 14327 757
rect 14107 754 14108 756
rect 14189 754 14198 756
rect 13871 738 13877 739
rect 13917 738 13923 744
rect 13957 738 13966 747
rect 14004 738 14013 747
rect 14096 746 14110 754
rect 14184 747 14198 754
rect 14269 750 14333 756
rect 14396 750 14411 756
rect 14418 754 14419 756
rect 14460 752 14461 753
rect 14184 746 14189 747
rect 14110 745 14113 746
rect 13623 734 13624 736
rect 13625 727 13628 733
rect 13697 731 13712 736
rect 13865 732 13871 738
rect 13923 733 13929 738
rect 13977 734 13989 738
rect 14030 734 14046 744
rect 14108 742 14109 745
rect 14113 742 14152 745
rect 14182 743 14189 746
rect 14275 745 14290 750
rect 14321 747 14330 750
rect 14275 744 14281 745
rect 14321 744 14327 747
rect 14109 740 14152 742
rect 14113 737 14152 740
rect 14175 739 14182 743
rect 14184 739 14189 743
rect 14330 742 14344 747
rect 14411 745 14424 750
rect 14460 747 14468 752
rect 14556 751 14557 756
rect 14590 750 14593 756
rect 14645 753 14651 759
rect 14656 758 14672 764
rect 14674 758 14690 764
rect 14697 759 14703 764
rect 14717 762 14720 768
rect 14756 761 14765 770
rect 14691 753 14697 759
rect 14722 756 14724 760
rect 14752 757 14753 758
rect 14410 742 14412 745
rect 14424 742 14430 745
rect 14461 744 14468 747
rect 14557 746 14558 750
rect 14593 744 14595 750
rect 14679 745 14682 747
rect 14470 742 14471 744
rect 14724 743 14732 756
rect 14753 754 14756 757
rect 14768 756 14776 768
rect 14780 758 14782 788
rect 14811 787 14814 788
rect 14818 779 14861 791
rect 16298 785 16301 793
rect 16332 790 16334 793
rect 16335 790 16349 794
rect 16332 786 16349 790
rect 14812 776 14861 779
rect 16301 777 16305 785
rect 14812 770 14821 776
rect 14832 774 14848 776
rect 14861 774 14882 776
rect 16305 775 16306 777
rect 14821 764 14830 770
rect 14824 763 14830 764
rect 14848 768 14882 774
rect 16306 771 16307 775
rect 16333 774 16349 786
rect 16383 790 16391 794
rect 16429 792 16445 808
rect 16479 801 16484 808
rect 16524 801 16528 808
rect 16580 807 16591 808
rect 16621 807 16637 808
rect 16687 807 16688 808
rect 16736 807 16744 814
rect 16767 811 16768 817
rect 16803 811 16809 821
rect 16819 814 16823 821
rect 16837 819 16854 824
rect 16885 819 16892 832
rect 16894 828 16896 832
rect 17025 832 17027 844
rect 17037 840 17049 844
rect 17065 842 17086 844
rect 17056 841 17065 842
rect 17051 840 17058 841
rect 17037 836 17051 840
rect 16837 818 16839 819
rect 16837 815 16838 818
rect 16883 817 16885 819
rect 16882 816 16883 817
rect 16823 812 16827 814
rect 16836 812 16837 813
rect 16882 812 16885 816
rect 16915 812 16927 815
rect 16809 809 16810 811
rect 16764 808 16766 809
rect 16823 808 16834 812
rect 16881 808 16882 812
rect 16915 808 16931 812
rect 16933 808 16949 824
rect 16951 808 16967 824
rect 17025 820 17033 832
rect 17037 831 17053 832
rect 17037 830 17047 831
rect 16969 808 16978 812
rect 17028 810 17029 814
rect 16753 807 16763 808
rect 16580 806 16592 807
rect 16587 804 16592 806
rect 16620 804 16637 807
rect 16688 806 16691 807
rect 16479 792 16483 801
rect 16383 774 16399 790
rect 16429 774 16445 790
rect 16479 787 16495 790
rect 16474 781 16495 787
rect 16515 787 16524 801
rect 16587 792 16591 804
rect 16619 799 16620 803
rect 16617 794 16619 798
rect 16621 792 16637 804
rect 16660 798 16672 806
rect 16691 804 16694 806
rect 16724 804 16753 807
rect 16675 799 16724 804
rect 16725 799 16731 804
rect 16736 799 16744 804
rect 16810 799 16812 804
rect 16821 803 16836 808
rect 16881 806 16886 808
rect 16915 807 16932 808
rect 16937 807 16949 808
rect 16515 785 16526 787
rect 16535 785 16547 791
rect 16587 785 16588 792
rect 16615 788 16617 792
rect 16504 783 16526 785
rect 16536 783 16547 785
rect 16586 783 16591 785
rect 16498 781 16503 783
rect 16468 775 16474 781
rect 16479 774 16495 781
rect 16513 779 16515 783
rect 16520 781 16526 783
rect 16547 781 16551 783
rect 16526 775 16532 781
rect 16535 778 16547 779
rect 16335 771 16339 774
rect 14825 759 14828 763
rect 14848 758 14864 768
rect 14882 762 14899 768
rect 14885 758 14891 762
rect 14899 760 14905 762
rect 14905 758 14909 760
rect 14931 758 14937 764
rect 14780 757 14795 758
rect 14780 756 14799 757
rect 14756 750 14761 754
rect 14796 752 14814 756
rect 14831 753 14837 756
rect 14879 753 14885 758
rect 14780 750 14814 752
rect 14837 751 14885 753
rect 14937 752 14943 758
rect 16307 754 16315 771
rect 16339 754 16346 771
rect 16349 758 16365 774
rect 16367 758 16383 774
rect 16445 772 16453 774
rect 16471 772 16479 774
rect 16545 772 16547 778
rect 16551 772 16559 779
rect 16584 778 16586 783
rect 16587 778 16591 783
rect 16584 774 16591 778
rect 16584 772 16586 774
rect 16445 758 16461 772
rect 16463 758 16479 772
rect 16526 757 16589 772
rect 16613 760 16615 786
rect 16621 774 16637 790
rect 16648 782 16656 794
rect 16660 793 16681 794
rect 16719 793 16725 799
rect 16660 792 16678 793
rect 16637 763 16641 767
rect 16648 763 16656 772
rect 16660 763 16662 792
rect 16813 788 16815 796
rect 16821 794 16843 803
rect 16821 792 16836 794
rect 16873 792 16886 806
rect 16911 804 16913 807
rect 16917 806 16931 807
rect 16915 803 16931 806
rect 16967 805 16983 808
rect 16965 803 16983 805
rect 16873 790 16881 792
rect 16903 791 16911 803
rect 16913 801 16949 803
rect 16913 793 16933 801
rect 16946 800 16949 801
rect 16947 793 16949 800
rect 16953 799 16961 803
rect 16965 799 16987 803
rect 16967 794 16987 799
rect 17025 798 17033 810
rect 17037 800 17039 830
rect 17056 826 17058 840
rect 17098 838 17104 844
rect 17156 838 17162 844
rect 17195 841 17200 845
rect 17488 841 17493 845
rect 17487 832 17495 841
rect 17499 834 17501 839
rect 17531 834 17533 846
rect 17791 845 17793 865
rect 17825 863 17827 872
rect 17862 863 17863 872
rect 17981 868 17998 881
rect 18026 868 18031 872
rect 17981 866 17990 868
rect 17981 865 17989 866
rect 18015 865 18023 866
rect 17824 857 17825 862
rect 17822 849 17823 855
rect 17543 844 17551 845
rect 17499 832 17533 834
rect 17537 832 17551 844
rect 17071 826 17072 832
rect 17543 830 17551 832
rect 17182 829 17185 830
rect 17158 827 17193 829
rect 17056 818 17057 826
rect 17154 825 17158 827
rect 17057 800 17060 814
rect 17072 812 17074 825
rect 17125 808 17154 825
rect 17156 814 17158 817
rect 17166 812 17182 827
rect 17161 811 17182 812
rect 17193 824 17353 827
rect 17037 798 17071 800
rect 17057 795 17060 798
rect 16815 778 16818 788
rect 16818 769 16820 778
rect 16821 774 16836 790
rect 16873 774 16887 790
rect 16910 781 16911 788
rect 16820 765 16821 769
rect 16637 762 16662 763
rect 16691 762 16694 763
rect 16637 760 16694 762
rect 16637 758 16653 760
rect 16821 759 16822 763
rect 14761 749 14797 750
rect 14780 744 14792 749
rect 14847 744 14858 749
rect 16315 746 16318 754
rect 16346 748 16351 754
rect 16351 745 16355 748
rect 16545 745 16547 757
rect 16550 745 16584 757
rect 16589 756 16591 757
rect 16698 756 16725 759
rect 16822 757 16823 759
rect 16837 758 16853 772
rect 16855 758 16871 772
rect 16903 769 16911 781
rect 16915 774 16933 793
rect 16967 792 16983 794
rect 16967 774 16983 790
rect 17013 774 17028 790
rect 17030 775 17032 789
rect 17037 786 17049 794
rect 17059 786 17071 794
rect 17073 790 17074 808
rect 17160 805 17170 811
rect 17193 808 17359 824
rect 17421 808 17437 824
rect 17439 808 17455 824
rect 17499 820 17511 828
rect 17521 820 17533 828
rect 17499 810 17501 820
rect 17551 816 17555 830
rect 17577 828 17579 845
rect 17579 819 17580 828
rect 17607 819 17610 845
rect 17612 843 17661 845
rect 17696 843 17698 844
rect 17612 833 17654 843
rect 17732 838 17733 843
rect 17699 827 17700 836
rect 17733 827 17734 836
rect 17790 834 17791 844
rect 17821 843 17822 847
rect 17820 837 17821 843
rect 17649 811 17654 823
rect 17701 817 17702 820
rect 17734 816 17735 820
rect 17789 819 17790 832
rect 17818 827 17820 836
rect 17860 829 17862 862
rect 17973 855 17989 865
rect 18026 864 18030 868
rect 17910 845 17973 855
rect 18018 851 18026 864
rect 17901 844 17910 845
rect 17895 842 17901 844
rect 17885 834 17895 842
rect 17817 821 17818 826
rect 17858 820 17860 827
rect 17702 811 17703 814
rect 17735 811 17736 814
rect 17788 811 17789 818
rect 17802 811 17808 817
rect 17816 816 17817 820
rect 17857 818 17858 820
rect 17865 818 17885 834
rect 17815 814 17816 816
rect 17814 812 17815 814
rect 17848 811 17854 817
rect 17856 813 17865 818
rect 17855 811 17865 813
rect 17611 808 17612 810
rect 17703 808 17704 810
rect 17165 803 17170 805
rect 17290 803 17299 808
rect 17337 803 17346 808
rect 17077 802 17086 803
rect 17075 798 17083 802
rect 17086 799 17101 802
rect 17101 798 17104 799
rect 17098 792 17104 798
rect 17156 792 17162 798
rect 17170 794 17179 803
rect 17281 794 17290 803
rect 17346 794 17355 803
rect 17272 792 17279 793
rect 17104 790 17110 792
rect 16915 772 16949 774
rect 16962 772 16967 774
rect 17060 772 17063 786
rect 17073 774 17079 790
rect 17104 786 17125 790
rect 17150 786 17156 792
rect 17266 791 17272 792
rect 17323 791 17327 793
rect 17359 792 17375 808
rect 17405 792 17421 808
rect 17432 803 17438 808
rect 17432 802 17447 803
rect 17426 796 17432 802
rect 17455 798 17471 808
rect 17478 802 17484 808
rect 17431 791 17432 793
rect 17464 791 17469 798
rect 17484 796 17490 802
rect 17502 800 17503 808
rect 17264 790 17266 791
rect 17263 787 17264 790
rect 17328 789 17330 790
rect 17109 774 17125 786
rect 17176 778 17203 781
rect 17159 774 17176 778
rect 17203 774 17211 778
rect 16915 769 16967 772
rect 17028 769 17034 772
rect 17063 771 17067 772
rect 16915 757 16919 765
rect 16951 758 16967 769
rect 17029 762 17046 769
rect 17063 762 17073 771
rect 17029 758 17045 762
rect 17046 760 17051 762
rect 17055 760 17067 762
rect 17051 759 17067 760
rect 17047 758 17067 759
rect 17125 758 17141 774
rect 17211 772 17214 774
rect 17279 772 17285 778
rect 17288 772 17290 779
rect 17330 772 17331 778
rect 17359 774 17375 790
rect 17405 774 17421 790
rect 17423 779 17432 791
rect 17214 763 17234 772
rect 17263 767 17264 769
rect 17273 766 17279 772
rect 17331 766 17337 772
rect 17352 763 17359 774
rect 17234 762 17236 763
rect 17236 759 17242 762
rect 16591 751 16612 756
rect 16612 747 16628 751
rect 16660 748 16672 756
rect 16823 754 16824 756
rect 16719 747 16725 753
rect 16750 747 16805 753
rect 16824 750 16825 754
rect 16825 747 16827 748
rect 16834 747 16843 756
rect 16913 747 16919 756
rect 16971 747 16977 753
rect 16978 747 16987 756
rect 17032 751 17035 758
rect 14858 743 14860 744
rect 14344 739 14353 742
rect 14430 741 14432 742
rect 14732 741 14733 743
rect 16318 741 16320 745
rect 14175 738 14189 739
rect 14162 737 14175 738
rect 14182 735 14184 738
rect 14353 735 14364 739
rect 14407 737 14408 739
rect 14364 734 14367 735
rect 13973 733 14055 734
rect 13923 732 13989 733
rect 13966 731 13989 732
rect 13712 726 13724 731
rect 13966 729 13973 731
rect 13977 730 13989 731
rect 14055 729 14058 732
rect 14174 731 14181 734
rect 14367 731 14376 734
rect 14404 733 14406 736
rect 14376 729 14383 731
rect 14399 729 14403 731
rect 13962 728 13966 729
rect 13955 726 13962 728
rect 13992 727 13993 729
rect 14058 728 14060 729
rect 13414 721 13485 723
rect 13238 719 13253 720
rect 13415 719 13485 721
rect 13517 719 13521 725
rect 13628 723 13630 726
rect 13241 716 13253 719
rect 11478 705 11485 712
rect 11564 706 11574 709
rect 11575 706 11587 715
rect 11610 714 11612 715
rect 11612 709 11652 714
rect 11674 709 11686 714
rect 13177 712 13182 716
rect 13254 714 13257 716
rect 13406 712 13414 719
rect 13416 717 13426 719
rect 13416 712 13420 717
rect 11652 707 11686 709
rect 11652 706 11700 707
rect 11722 706 11728 712
rect 11780 706 11786 712
rect 11149 698 11160 701
rect 11243 698 11251 701
rect 11271 700 11279 701
rect 10612 688 10613 692
rect 10575 676 10609 678
rect 10613 676 10621 688
rect 10708 686 10714 692
rect 10766 686 10772 692
rect 10798 688 10805 692
rect 10914 691 10920 697
rect 10960 691 10966 697
rect 11006 691 11149 698
rect 11221 691 11243 698
rect 11277 692 11279 700
rect 11280 693 11286 698
rect 11299 694 11311 701
rect 10901 688 10903 691
rect 10798 687 10810 688
rect 10714 680 10720 686
rect 10760 680 10766 686
rect 10798 685 10813 687
rect 10820 685 10832 688
rect 10900 687 10901 688
rect 10899 685 10900 687
rect 10908 685 10914 691
rect 10966 685 10972 691
rect 10973 689 10994 691
rect 11216 689 11221 691
rect 11210 687 11216 689
rect 11279 688 11280 692
rect 11288 689 11291 691
rect 10977 685 11012 687
rect 10798 680 10810 685
rect 10813 680 10835 685
rect 10897 683 10899 685
rect 10835 678 10841 680
rect 10841 676 10848 678
rect 10848 675 10853 676
rect 10862 675 10912 683
rect 10965 682 10977 685
rect 10956 680 10965 682
rect 11017 680 11019 685
rect 11200 684 11208 687
rect 11280 686 11281 687
rect 11193 682 11200 684
rect 11186 679 11193 682
rect 11281 680 11283 682
rect 11181 678 11186 679
rect 11283 678 11284 680
rect 11297 678 11304 684
rect 11316 682 11374 701
rect 11401 692 11402 698
rect 11465 692 11466 701
rect 11470 693 11478 703
rect 11485 702 11489 705
rect 11550 702 11575 706
rect 11672 704 11685 706
rect 11473 691 11478 693
rect 11489 692 11500 702
rect 11316 678 11349 682
rect 11374 678 11378 682
rect 11403 679 11404 682
rect 10955 676 10956 678
rect 11175 676 11181 678
rect 11284 676 11285 678
rect 10611 672 10613 675
rect 10853 674 10912 675
rect 10862 672 10912 674
rect 10318 656 10321 662
rect 10242 643 10306 649
rect 10316 648 10318 656
rect 10362 652 10379 672
rect 10402 666 10409 672
rect 10575 666 10587 672
rect 10597 666 10609 672
rect 10839 666 10862 672
rect 10409 664 10615 666
rect 10828 664 10839 666
rect 10248 637 10275 643
rect 10294 637 10300 643
rect 10310 642 10316 647
rect 10320 642 10329 644
rect 10379 643 10387 652
rect 10556 642 10557 660
rect 9238 623 9265 629
rect 10058 626 10061 630
rect 10251 626 10275 637
rect 10310 635 10329 642
rect 10388 639 10392 642
rect 10392 636 10397 639
rect 10397 635 10405 636
rect 10310 630 10325 635
rect 10405 631 10441 635
rect 10309 626 10325 630
rect 10441 628 10461 631
rect 10555 630 10557 642
rect 10615 654 10774 664
rect 10786 654 10828 664
rect 10952 663 10955 674
rect 11019 663 11022 676
rect 11170 674 11175 676
rect 11167 673 11170 674
rect 11162 672 11167 673
rect 11156 670 11162 672
rect 11285 670 11288 676
rect 11304 671 11312 678
rect 11349 671 11357 678
rect 11378 676 11380 678
rect 11405 677 11406 687
rect 11457 681 11470 682
rect 11457 679 11466 681
rect 11500 679 11505 692
rect 11550 688 11599 702
rect 11624 698 11670 704
rect 11688 703 11690 706
rect 11700 704 11720 706
rect 11728 704 11747 706
rect 11671 700 11686 702
rect 11616 694 11624 698
rect 11550 687 11575 688
rect 11599 687 11605 688
rect 11607 687 11616 694
rect 11532 678 11550 687
rect 11599 686 11607 687
rect 11605 685 11609 686
rect 11595 677 11602 683
rect 11609 682 11617 685
rect 11617 681 11622 682
rect 11622 680 11627 681
rect 11628 678 11631 679
rect 11399 676 11420 677
rect 11457 676 11463 677
rect 11380 673 11384 676
rect 11137 668 11156 670
rect 11100 664 11137 668
rect 11023 663 11100 664
rect 10914 655 11100 663
rect 11288 660 11301 670
rect 11312 660 11334 671
rect 11357 663 11367 671
rect 11384 663 11388 673
rect 11399 671 11405 676
rect 11406 672 11420 676
rect 11446 671 11463 676
rect 11504 671 11505 676
rect 11515 671 11530 677
rect 11405 665 11411 671
rect 11451 665 11457 671
rect 11495 663 11515 671
rect 11586 669 11595 677
rect 11634 676 11639 678
rect 11640 674 11646 676
rect 10615 652 10786 654
rect 10914 653 11029 655
rect 10615 642 10617 652
rect 10914 651 11026 653
rect 10914 649 11019 651
rect 10914 648 10982 649
rect 10914 645 10966 648
rect 10908 644 10972 645
rect 10886 642 10972 644
rect 10615 634 10621 642
rect 10880 639 10897 642
rect 10908 639 10972 642
rect 11005 641 11017 649
rect 11022 643 11026 651
rect 10862 636 10880 639
rect 10616 630 10621 634
rect 10843 633 10862 636
rect 10914 633 10920 639
rect 10946 636 10952 639
rect 10960 633 10966 639
rect 11024 636 11026 643
rect 11301 642 11347 660
rect 11367 652 11397 663
rect 11377 647 11411 652
rect 11431 647 11432 660
rect 11468 652 11495 663
rect 11504 660 11505 663
rect 11377 646 11448 647
rect 11456 646 11485 652
rect 11377 643 11485 646
rect 11383 642 11388 643
rect 11301 641 11349 642
rect 10828 631 10843 633
rect 10632 630 10672 631
rect 10826 630 10828 631
rect 10471 628 10632 630
rect 10672 628 10701 630
rect 10555 626 10558 628
rect 10614 626 10621 628
rect 9266 623 9293 624
rect 8650 621 8651 622
rect 8554 615 8571 621
rect 8646 616 8650 621
rect 10061 618 10069 626
rect 10129 618 10136 625
rect 10069 617 10129 618
rect 8643 615 8646 616
rect 8571 611 8643 615
rect 10293 610 10309 626
rect 10558 615 10564 626
rect 10611 618 10614 625
rect 10701 622 10762 628
rect 10772 622 10822 630
rect 11022 627 11024 636
rect 10603 615 10611 618
rect 10564 613 10605 615
rect 10946 613 10959 624
rect 11000 616 11022 627
rect 11301 626 11347 641
rect 11351 637 11354 639
rect 11354 636 11356 637
rect 11356 633 11363 636
rect 11383 634 11397 642
rect 11431 634 11432 643
rect 11503 637 11504 653
rect 11545 652 11586 669
rect 11640 668 11648 674
rect 11652 670 11654 672
rect 11684 670 11686 700
rect 11690 690 11698 702
rect 11728 700 11734 704
rect 11774 700 11780 706
rect 11798 693 11809 702
rect 13182 696 13203 712
rect 13247 710 13271 712
rect 13251 705 13271 710
rect 13406 707 13416 712
rect 13413 705 13416 707
rect 13203 695 13205 696
rect 11652 668 11686 670
rect 11690 668 11698 680
rect 11809 678 11812 692
rect 13209 689 13210 692
rect 13207 678 13214 687
rect 13251 680 13253 705
rect 13257 700 13265 705
rect 13271 699 13277 705
rect 13411 701 13413 705
rect 13405 699 13413 701
rect 13277 694 13283 699
rect 13405 695 13411 699
rect 13283 692 13286 694
rect 13219 678 13253 680
rect 13257 678 13265 690
rect 13286 688 13287 692
rect 13399 689 13405 695
rect 13409 692 13410 694
rect 13408 688 13409 691
rect 13418 689 13420 712
rect 13450 715 13505 719
rect 13450 701 13473 715
rect 13481 713 13505 715
rect 13525 713 13526 715
rect 13486 708 13505 713
rect 13526 708 13530 713
rect 13630 710 13637 723
rect 13724 722 13754 726
rect 13973 724 13989 726
rect 13724 714 13766 722
rect 13493 701 13505 708
rect 13530 706 13531 708
rect 13637 705 13640 710
rect 13718 709 13767 710
rect 13450 695 13457 701
rect 13450 693 13463 695
rect 13450 689 13452 693
rect 13457 689 13463 693
rect 13468 691 13477 700
rect 13496 696 13505 701
rect 13536 696 13539 701
rect 13499 691 13505 696
rect 13407 685 13408 687
rect 13451 685 13452 689
rect 13469 687 13486 691
rect 13502 689 13505 691
rect 13539 689 13545 696
rect 13640 695 13677 705
rect 13718 702 13732 709
rect 13748 708 13767 709
rect 13764 703 13767 708
rect 13717 699 13718 701
rect 13677 693 13683 695
rect 13715 694 13717 699
rect 13683 692 13688 693
rect 13714 692 13715 694
rect 13504 687 13505 689
rect 13470 686 13486 687
rect 13545 686 13547 689
rect 13688 688 13704 692
rect 13704 687 13706 688
rect 13287 680 13289 685
rect 13406 680 13407 685
rect 13472 682 13475 686
rect 13477 682 13486 686
rect 13478 680 13479 682
rect 11812 676 11813 678
rect 13214 676 13215 678
rect 13218 676 13219 678
rect 13405 676 13406 678
rect 13479 677 13480 680
rect 11648 664 11651 666
rect 11652 656 11664 664
rect 11674 656 11686 664
rect 11813 661 11816 676
rect 11530 646 11545 652
rect 11652 648 11661 656
rect 11815 648 11816 661
rect 13214 660 13218 676
rect 13254 674 13257 676
rect 13219 666 13231 674
rect 13241 666 13253 674
rect 13289 660 13293 676
rect 13213 654 13214 658
rect 13293 657 13294 660
rect 11516 641 11528 646
rect 11507 637 11516 641
rect 11363 631 11369 633
rect 11381 630 11397 634
rect 11372 626 11397 630
rect 11431 626 11433 630
rect 11365 622 11390 626
rect 10960 613 11000 616
rect 10571 610 10587 613
rect 10589 610 10605 613
rect 11365 610 11381 622
rect 11390 619 11398 622
rect 11398 618 11407 619
rect 11433 615 11438 626
rect 11465 620 11507 637
rect 11462 619 11465 620
rect 11456 618 11462 619
rect 11494 618 11501 620
rect 11490 615 11494 618
rect 11438 611 11459 615
rect 11481 611 11490 615
rect 11631 606 11655 629
rect 11661 626 11700 648
rect 11700 621 11709 626
rect 11806 622 11815 643
rect 13213 630 13215 654
rect 13293 630 13294 654
rect 13405 649 13457 663
rect 13478 662 13480 675
rect 13507 672 13519 685
rect 13547 672 13559 686
rect 13709 685 13715 687
rect 13715 683 13723 685
rect 13720 681 13724 683
rect 13720 676 13727 681
rect 13764 678 13766 703
rect 13767 697 13768 702
rect 13770 698 13778 710
rect 13923 694 13951 695
rect 13987 694 13989 724
rect 13993 714 14001 726
rect 14060 712 14062 728
rect 14383 727 14389 729
rect 14396 727 14399 729
rect 14116 720 14122 726
rect 14174 720 14180 726
rect 14380 723 14400 727
rect 14432 723 14453 741
rect 14458 738 14469 740
rect 14380 721 14396 723
rect 14375 720 14380 721
rect 14400 720 14408 723
rect 14122 714 14128 720
rect 14168 714 14174 720
rect 14368 717 14375 720
rect 14408 719 14411 720
rect 14453 719 14458 723
rect 14363 716 14368 717
rect 14411 716 14417 719
rect 14458 716 14462 719
rect 14466 716 14468 738
rect 14469 737 14470 738
rect 14472 737 14480 740
rect 14470 734 14480 737
rect 14472 729 14480 734
rect 14559 733 14560 741
rect 14596 737 14599 741
rect 14560 729 14561 733
rect 14589 729 14601 737
rect 14611 729 14623 737
rect 14686 729 14699 741
rect 14472 728 14481 729
rect 14477 726 14481 728
rect 14472 716 14480 718
rect 14354 713 14363 716
rect 14349 711 14354 713
rect 13768 693 13769 694
rect 13943 692 13951 694
rect 13955 692 13989 694
rect 13993 692 14001 704
rect 14060 694 14062 710
rect 14333 706 14349 711
rect 14417 706 14428 716
rect 14462 707 14480 716
rect 14444 706 14480 707
rect 14481 706 14504 726
rect 14561 724 14568 729
rect 14585 727 14588 729
rect 14601 725 14602 729
rect 14608 725 14614 729
rect 14562 723 14568 724
rect 14577 723 14585 725
rect 14589 723 14635 725
rect 14556 717 14562 723
rect 14589 717 14591 723
rect 14614 717 14620 723
rect 14621 717 14635 723
rect 14560 713 14562 714
rect 14558 709 14560 713
rect 14317 701 14333 706
rect 14428 705 14435 706
rect 14473 705 14506 706
rect 14428 702 14436 705
rect 14410 701 14444 702
rect 14470 701 14531 705
rect 14621 702 14623 717
rect 14627 713 14642 717
rect 14630 705 14642 713
rect 14699 712 14718 729
rect 14733 715 14767 741
rect 14862 723 14885 741
rect 16355 740 16363 745
rect 16581 742 16582 745
rect 16628 742 16648 747
rect 16648 741 16653 742
rect 16725 741 16731 747
rect 16771 741 16777 747
rect 16547 740 16549 741
rect 16320 737 16322 740
rect 16363 737 16368 740
rect 16537 739 16547 740
rect 16526 738 16547 739
rect 16653 738 16657 741
rect 16778 738 16787 747
rect 16825 745 16834 747
rect 16825 742 16840 745
rect 16825 738 16834 742
rect 16840 740 16844 742
rect 16919 741 16931 747
rect 16965 741 16978 747
rect 17034 744 17035 751
rect 16844 739 16847 740
rect 16368 736 16370 737
rect 16535 736 16554 738
rect 16323 733 16324 736
rect 16370 733 16374 736
rect 16324 731 16325 733
rect 16374 731 16378 733
rect 16325 727 16327 731
rect 16378 729 16381 731
rect 16468 729 16474 735
rect 16526 729 16532 735
rect 16535 733 16572 736
rect 16579 733 16580 736
rect 16546 729 16572 733
rect 16575 729 16579 731
rect 16611 729 16612 730
rect 16381 726 16385 729
rect 16327 720 16331 726
rect 16385 720 16395 726
rect 16398 720 16410 724
rect 16474 723 16480 729
rect 16520 723 16526 729
rect 16572 726 16612 729
rect 16572 723 16611 726
rect 16657 725 16674 738
rect 16778 737 16779 738
rect 16847 736 16854 739
rect 16922 738 16931 741
rect 16969 738 16978 741
rect 17028 739 17035 744
rect 17063 742 17067 758
rect 17105 747 17114 756
rect 17170 747 17179 756
rect 17242 754 17253 759
rect 17346 758 17359 763
rect 17421 769 17430 774
rect 17431 769 17432 779
rect 17421 763 17432 769
rect 17435 763 17437 791
rect 17503 790 17505 791
rect 17501 785 17505 790
rect 17554 790 17555 808
rect 17661 799 17673 804
rect 17705 796 17706 799
rect 17736 796 17737 805
rect 17787 799 17788 808
rect 17796 805 17802 811
rect 17854 808 17860 811
rect 17909 808 17925 824
rect 18498 819 18499 1015
rect 18688 819 18689 1015
rect 18774 819 18775 1015
rect 19047 819 19048 1015
rect 19244 819 19245 1015
rect 17852 805 17860 808
rect 17852 804 17854 805
rect 17855 800 17856 802
rect 17856 797 17858 800
rect 17421 758 17437 763
rect 17486 773 17547 785
rect 17554 779 17567 790
rect 17553 774 17567 779
rect 17597 774 17612 790
rect 17613 777 17615 793
rect 17706 789 17707 793
rect 17737 789 17738 795
rect 17486 759 17551 773
rect 17517 758 17533 759
rect 17535 758 17551 759
rect 17578 758 17579 760
rect 17613 758 17629 774
rect 17707 767 17711 785
rect 17738 779 17739 788
rect 17787 787 17789 794
rect 17852 790 17853 794
rect 17858 791 17861 797
rect 17893 792 17909 808
rect 17943 802 17971 808
rect 17937 794 17971 802
rect 17933 791 17935 794
rect 17943 790 17971 794
rect 17789 781 17790 787
rect 17852 782 17869 790
rect 17739 766 17744 779
rect 17791 774 17799 780
rect 17853 776 17869 782
rect 17925 779 17933 790
rect 17922 778 17933 779
rect 17937 788 17971 790
rect 17853 774 17863 776
rect 17799 773 17801 774
rect 17711 760 17712 766
rect 17744 759 17746 766
rect 17801 765 17815 773
rect 17853 766 17854 774
rect 17869 768 17874 776
rect 17922 770 17931 778
rect 17850 765 17854 766
rect 17796 764 17829 765
rect 17850 764 17860 765
rect 17796 759 17802 764
rect 17346 756 17352 758
rect 17423 757 17437 758
rect 17549 757 17552 758
rect 17431 756 17484 757
rect 17264 754 17265 756
rect 17346 754 17355 756
rect 17028 738 17034 739
rect 17074 738 17080 744
rect 17114 738 17123 747
rect 17161 738 17170 747
rect 17253 746 17267 754
rect 17341 747 17355 754
rect 17426 750 17490 756
rect 17553 750 17568 756
rect 17575 754 17576 756
rect 17617 752 17618 753
rect 17341 746 17346 747
rect 17267 745 17270 746
rect 16780 734 16781 736
rect 16782 727 16785 733
rect 16854 731 16869 736
rect 17022 732 17028 738
rect 17080 733 17086 738
rect 17134 734 17146 738
rect 17187 734 17203 744
rect 17265 742 17266 745
rect 17270 742 17309 745
rect 17339 743 17346 746
rect 17432 745 17447 750
rect 17478 747 17487 750
rect 17432 744 17438 745
rect 17478 744 17484 747
rect 17266 740 17309 742
rect 17270 737 17309 740
rect 17332 739 17339 743
rect 17341 739 17346 743
rect 17487 742 17501 747
rect 17568 745 17581 750
rect 17617 747 17625 752
rect 17713 751 17714 756
rect 17747 750 17750 756
rect 17802 753 17808 759
rect 17813 758 17829 764
rect 17831 758 17847 764
rect 17854 759 17860 764
rect 17874 762 17877 768
rect 17913 761 17922 770
rect 17848 753 17854 759
rect 17879 756 17881 760
rect 17909 757 17910 758
rect 17567 742 17569 745
rect 17581 742 17587 745
rect 17618 744 17625 747
rect 17714 746 17715 750
rect 17750 744 17752 750
rect 17836 745 17839 747
rect 17627 742 17628 744
rect 17881 743 17889 756
rect 17910 754 17913 757
rect 17925 756 17933 768
rect 17937 758 17939 788
rect 17968 787 17971 788
rect 17975 779 18018 791
rect 17969 776 18018 779
rect 17969 770 17978 776
rect 17989 774 18005 776
rect 18018 774 18039 776
rect 17978 764 17987 770
rect 17981 763 17987 764
rect 18005 768 18039 774
rect 17982 759 17985 763
rect 18005 758 18021 768
rect 18039 762 18056 768
rect 18042 758 18048 762
rect 18056 760 18062 762
rect 18062 758 18066 760
rect 18088 758 18094 764
rect 17937 757 17952 758
rect 17937 756 17956 757
rect 17913 750 17918 754
rect 17953 752 17971 756
rect 17988 753 17994 756
rect 18036 753 18042 758
rect 17937 750 17971 752
rect 17994 751 18042 753
rect 18094 752 18100 758
rect 17918 749 17954 750
rect 17937 744 17949 749
rect 18004 744 18015 749
rect 18015 743 18017 744
rect 17501 739 17510 742
rect 17587 741 17589 742
rect 17889 741 17890 743
rect 17332 738 17346 739
rect 17319 737 17332 738
rect 17339 735 17341 738
rect 17510 735 17521 739
rect 17564 737 17565 739
rect 17521 734 17524 735
rect 17130 733 17212 734
rect 17080 732 17146 733
rect 17123 731 17146 732
rect 16869 726 16881 731
rect 17123 729 17130 731
rect 17134 730 17146 731
rect 17212 729 17215 732
rect 17331 731 17338 734
rect 17524 731 17533 734
rect 17561 733 17563 736
rect 17533 729 17540 731
rect 17556 729 17560 731
rect 17119 728 17123 729
rect 17112 726 17119 728
rect 17149 727 17150 729
rect 17215 728 17217 729
rect 16571 721 16642 723
rect 16395 719 16410 720
rect 16572 719 16642 721
rect 16674 719 16678 725
rect 16785 723 16787 726
rect 16398 716 16410 719
rect 14721 706 14731 709
rect 14732 706 14744 715
rect 14767 714 14769 715
rect 14769 709 14809 714
rect 14831 709 14843 714
rect 16334 712 16339 716
rect 16411 714 16414 716
rect 16563 712 16571 719
rect 16573 717 16583 719
rect 16573 712 16577 717
rect 14809 707 14843 709
rect 14809 706 14857 707
rect 14879 706 14885 712
rect 14937 706 14943 712
rect 14306 698 14317 701
rect 14400 698 14408 701
rect 14428 700 14436 701
rect 13769 688 13770 692
rect 13732 676 13766 678
rect 13770 676 13778 688
rect 13865 686 13871 692
rect 13923 686 13929 692
rect 13955 688 13962 692
rect 14071 691 14077 697
rect 14117 691 14123 697
rect 14163 691 14306 698
rect 14378 691 14400 698
rect 14434 692 14436 700
rect 14437 693 14443 698
rect 14456 694 14468 701
rect 14058 688 14060 691
rect 13955 687 13967 688
rect 13871 680 13877 686
rect 13917 680 13923 686
rect 13955 685 13970 687
rect 13977 685 13989 688
rect 14057 687 14058 688
rect 14056 685 14057 687
rect 14065 685 14071 691
rect 14123 685 14129 691
rect 14130 689 14151 691
rect 14373 689 14378 691
rect 14367 687 14373 689
rect 14436 688 14437 692
rect 14445 689 14448 691
rect 14134 685 14169 687
rect 13955 680 13967 685
rect 13970 680 13992 685
rect 14054 683 14056 685
rect 13992 676 14005 680
rect 14005 675 14010 676
rect 14019 675 14069 683
rect 14122 682 14134 685
rect 14113 680 14122 682
rect 14174 680 14176 685
rect 14357 684 14365 687
rect 14437 686 14438 687
rect 14350 682 14357 684
rect 14112 676 14113 680
rect 14343 679 14350 682
rect 14438 680 14440 682
rect 14338 678 14343 679
rect 14332 676 14338 678
rect 14440 676 14442 680
rect 14454 678 14461 684
rect 14473 682 14531 701
rect 14558 692 14559 698
rect 14622 692 14623 701
rect 14627 693 14635 703
rect 14642 702 14646 705
rect 14707 702 14732 706
rect 14829 704 14842 706
rect 14630 691 14635 693
rect 14646 692 14657 702
rect 14473 678 14506 682
rect 13768 672 13770 675
rect 14010 674 14069 675
rect 14019 672 14069 674
rect 13475 656 13478 662
rect 13399 643 13463 649
rect 13473 648 13475 656
rect 13519 652 13536 672
rect 13559 666 13566 672
rect 13732 666 13744 672
rect 13754 666 13766 672
rect 13996 666 14019 672
rect 13566 664 13772 666
rect 13985 664 13996 666
rect 13405 637 13432 643
rect 13451 637 13457 643
rect 13467 642 13473 647
rect 13477 642 13486 644
rect 13536 643 13544 652
rect 13713 642 13714 660
rect 12393 623 12420 629
rect 13215 626 13218 630
rect 13408 626 13432 637
rect 13467 635 13486 642
rect 13545 639 13549 642
rect 13549 636 13554 639
rect 13554 635 13562 636
rect 13467 630 13482 635
rect 13562 631 13598 635
rect 13466 626 13482 630
rect 13598 628 13618 631
rect 13712 630 13714 642
rect 13772 654 13931 664
rect 13943 654 13985 664
rect 14109 663 14112 674
rect 14176 663 14179 676
rect 14327 674 14332 676
rect 14324 673 14327 674
rect 14319 672 14324 673
rect 14313 670 14319 672
rect 14442 670 14445 676
rect 14461 671 14469 678
rect 14506 671 14514 678
rect 14531 676 14537 682
rect 14560 679 14561 682
rect 14562 677 14563 687
rect 14614 681 14627 682
rect 14614 679 14623 681
rect 14657 679 14662 692
rect 14707 688 14756 702
rect 14781 698 14827 704
rect 14845 703 14847 706
rect 14857 704 14877 706
rect 14885 704 14904 706
rect 14828 700 14843 702
rect 14773 694 14781 698
rect 14707 687 14732 688
rect 14756 687 14762 688
rect 14764 687 14773 694
rect 14689 678 14707 687
rect 14756 686 14764 687
rect 14762 685 14766 686
rect 14752 677 14759 683
rect 14766 682 14774 685
rect 14774 681 14779 682
rect 14779 680 14784 681
rect 14785 678 14788 679
rect 14556 676 14577 677
rect 14614 676 14620 677
rect 14537 673 14541 676
rect 14294 668 14313 670
rect 14257 664 14294 668
rect 14180 663 14257 664
rect 14071 655 14257 663
rect 14445 660 14458 670
rect 14469 660 14491 671
rect 14514 663 14524 671
rect 14541 663 14545 673
rect 14556 671 14562 676
rect 14563 672 14577 676
rect 14603 671 14620 676
rect 14661 671 14662 676
rect 14672 671 14687 677
rect 14562 665 14568 671
rect 14608 665 14614 671
rect 14652 663 14672 671
rect 14743 669 14752 677
rect 14791 676 14796 678
rect 14797 674 14803 676
rect 13772 652 13943 654
rect 14071 653 14186 655
rect 13772 642 13774 652
rect 14071 651 14183 653
rect 14071 649 14176 651
rect 14071 648 14139 649
rect 14071 645 14123 648
rect 14065 644 14129 645
rect 14043 642 14129 644
rect 13772 634 13778 642
rect 14037 639 14054 642
rect 14065 639 14129 642
rect 14162 641 14174 649
rect 14179 643 14183 651
rect 14019 636 14037 639
rect 13773 630 13778 634
rect 14000 633 14019 636
rect 14071 633 14077 639
rect 14103 636 14109 639
rect 14117 633 14123 639
rect 14181 636 14183 643
rect 14458 642 14504 660
rect 14524 652 14554 663
rect 14534 647 14568 652
rect 14588 647 14589 660
rect 14625 652 14652 663
rect 14661 660 14662 663
rect 14534 646 14605 647
rect 14613 646 14642 652
rect 14534 643 14642 646
rect 14540 642 14545 643
rect 14458 641 14506 642
rect 13985 631 14000 633
rect 13789 630 13829 631
rect 13983 630 13985 631
rect 13628 628 13789 630
rect 13829 628 13858 630
rect 13712 626 13715 628
rect 13771 626 13778 628
rect 12421 623 12448 624
rect 11805 621 11806 622
rect 11709 615 11726 621
rect 11801 616 11805 621
rect 13218 618 13226 626
rect 13286 618 13293 625
rect 13226 617 13286 618
rect 11798 615 11801 616
rect 11726 611 11798 615
rect 13450 610 13466 626
rect 13715 615 13721 626
rect 13768 618 13771 625
rect 13858 622 13919 628
rect 13929 622 13979 630
rect 14179 627 14181 636
rect 13760 615 13768 618
rect 13721 613 13762 615
rect 14103 613 14116 624
rect 14157 616 14179 627
rect 14458 626 14504 641
rect 14508 637 14511 639
rect 14511 636 14513 637
rect 14513 633 14520 636
rect 14540 634 14554 642
rect 14588 634 14589 643
rect 14660 637 14661 653
rect 14702 652 14743 669
rect 14797 668 14805 674
rect 14809 670 14811 672
rect 14841 670 14843 700
rect 14847 690 14855 702
rect 14885 700 14891 704
rect 14931 700 14937 706
rect 14955 693 14966 702
rect 16339 696 16360 712
rect 16404 710 16428 712
rect 16408 705 16428 710
rect 16563 707 16573 712
rect 16570 705 16573 707
rect 16360 695 16362 696
rect 14809 668 14843 670
rect 14847 668 14855 680
rect 14966 678 14969 692
rect 16366 689 16367 692
rect 16364 678 16371 687
rect 16408 680 16410 705
rect 16414 700 16422 705
rect 16428 699 16434 705
rect 16568 701 16570 705
rect 16562 699 16570 701
rect 16434 694 16440 699
rect 16562 695 16568 699
rect 16440 692 16443 694
rect 16376 678 16410 680
rect 16414 678 16422 690
rect 16443 688 16444 692
rect 16556 689 16562 695
rect 16566 692 16567 694
rect 16565 688 16566 691
rect 16575 689 16577 712
rect 16607 715 16662 719
rect 16607 701 16630 715
rect 16638 713 16662 715
rect 16682 713 16683 715
rect 16643 708 16662 713
rect 16683 708 16687 713
rect 16787 710 16794 723
rect 16881 722 16911 726
rect 17130 724 17146 726
rect 16881 714 16923 722
rect 16650 701 16662 708
rect 16687 706 16688 708
rect 16794 705 16797 710
rect 16875 709 16924 710
rect 16607 695 16614 701
rect 16607 693 16620 695
rect 16607 689 16609 693
rect 16614 689 16620 693
rect 16625 691 16634 700
rect 16653 696 16662 701
rect 16693 696 16696 701
rect 16656 691 16662 696
rect 16564 685 16565 687
rect 16608 685 16609 689
rect 16626 687 16643 691
rect 16659 689 16662 691
rect 16696 689 16702 696
rect 16797 695 16834 705
rect 16875 702 16889 709
rect 16905 708 16924 709
rect 16921 703 16924 708
rect 16874 699 16875 701
rect 16834 693 16840 695
rect 16872 694 16874 699
rect 16840 692 16845 693
rect 16871 692 16872 694
rect 16661 687 16662 689
rect 16627 686 16643 687
rect 16702 686 16704 689
rect 16845 688 16861 692
rect 16861 687 16863 688
rect 16444 680 16446 685
rect 16563 680 16564 685
rect 16629 682 16632 686
rect 16634 682 16643 686
rect 16635 680 16636 682
rect 14969 676 14970 678
rect 16371 676 16372 678
rect 16375 676 16376 678
rect 16562 676 16563 678
rect 16636 677 16637 680
rect 14805 664 14808 666
rect 14809 656 14821 664
rect 14831 656 14843 664
rect 14970 661 14973 676
rect 14687 646 14702 652
rect 14809 648 14818 656
rect 14972 648 14973 661
rect 16371 660 16375 676
rect 16411 674 16414 676
rect 16376 666 16388 674
rect 16398 666 16410 674
rect 16446 660 16450 676
rect 16370 654 16371 658
rect 16450 657 16451 660
rect 14673 641 14685 646
rect 14664 637 14673 641
rect 14520 631 14526 633
rect 14538 630 14554 634
rect 14529 626 14554 630
rect 14588 626 14590 630
rect 14522 622 14547 626
rect 14117 613 14157 616
rect 13728 610 13744 613
rect 13746 610 13762 613
rect 14522 610 14538 622
rect 14547 619 14555 622
rect 14555 618 14564 619
rect 14590 615 14595 626
rect 14622 620 14664 637
rect 14619 619 14622 620
rect 14613 618 14619 619
rect 14651 618 14658 620
rect 14647 615 14651 618
rect 14595 611 14616 615
rect 14638 611 14647 615
rect 14788 606 14812 629
rect 14818 626 14857 648
rect 14857 621 14866 626
rect 14963 622 14972 643
rect 16370 630 16372 654
rect 16450 630 16451 654
rect 16562 649 16614 663
rect 16635 662 16637 675
rect 16664 672 16676 685
rect 16704 672 16716 686
rect 16866 685 16872 687
rect 16872 683 16880 685
rect 16877 681 16881 683
rect 16877 676 16884 681
rect 16921 678 16923 703
rect 16924 697 16925 702
rect 16927 698 16935 710
rect 17080 694 17108 695
rect 17144 694 17146 724
rect 17150 714 17158 726
rect 17217 712 17219 728
rect 17540 727 17546 729
rect 17553 727 17556 729
rect 17273 720 17279 726
rect 17331 720 17337 726
rect 17537 723 17557 727
rect 17589 723 17610 741
rect 17615 738 17626 740
rect 17537 721 17553 723
rect 17532 720 17537 721
rect 17557 720 17565 723
rect 17279 714 17285 720
rect 17325 714 17331 720
rect 17525 717 17532 720
rect 17565 719 17568 720
rect 17610 719 17615 723
rect 17520 716 17525 717
rect 17568 716 17574 719
rect 17615 716 17619 719
rect 17623 716 17625 738
rect 17626 737 17627 738
rect 17629 737 17637 740
rect 17627 734 17637 737
rect 17629 729 17637 734
rect 17716 733 17717 741
rect 17753 737 17756 741
rect 17717 729 17718 733
rect 17746 729 17758 737
rect 17768 729 17780 737
rect 17843 729 17856 741
rect 17629 728 17638 729
rect 17634 726 17638 728
rect 17629 716 17637 718
rect 17511 713 17520 716
rect 17506 711 17511 713
rect 16925 693 16926 694
rect 17100 692 17108 694
rect 17112 692 17146 694
rect 17150 692 17158 704
rect 17217 694 17219 710
rect 17490 706 17506 711
rect 17574 706 17585 716
rect 17619 707 17637 716
rect 17601 706 17637 707
rect 17638 706 17661 726
rect 17718 724 17725 729
rect 17742 727 17745 729
rect 17758 725 17759 729
rect 17765 725 17771 729
rect 17719 723 17725 724
rect 17734 723 17742 725
rect 17746 723 17792 725
rect 17713 717 17719 723
rect 17746 717 17748 723
rect 17771 717 17777 723
rect 17778 717 17792 723
rect 17717 713 17719 714
rect 17715 709 17717 713
rect 17474 701 17490 706
rect 17585 705 17592 706
rect 17630 705 17663 706
rect 17585 702 17593 705
rect 17567 701 17601 702
rect 17627 701 17688 705
rect 17778 702 17780 717
rect 17784 713 17799 717
rect 17787 705 17799 713
rect 17856 712 17875 729
rect 17890 715 17924 741
rect 18019 723 18042 741
rect 17878 706 17888 709
rect 17889 706 17901 715
rect 17924 714 17926 715
rect 17926 709 17966 714
rect 17988 709 18000 714
rect 17966 707 18000 709
rect 17966 706 18014 707
rect 18036 706 18042 712
rect 18094 706 18100 712
rect 17463 698 17474 701
rect 17557 698 17565 701
rect 17585 700 17593 701
rect 16926 688 16927 692
rect 16889 676 16923 678
rect 16927 676 16935 688
rect 17022 686 17028 692
rect 17080 686 17086 692
rect 17112 688 17119 692
rect 17228 691 17234 697
rect 17274 691 17280 697
rect 17320 691 17463 698
rect 17535 691 17557 698
rect 17591 692 17593 700
rect 17594 693 17600 698
rect 17613 694 17625 701
rect 17215 688 17217 691
rect 17112 687 17124 688
rect 17028 680 17034 686
rect 17074 680 17080 686
rect 17112 685 17127 687
rect 17134 685 17146 688
rect 17214 687 17215 688
rect 17213 685 17214 687
rect 17222 685 17228 691
rect 17280 685 17286 691
rect 17287 689 17308 691
rect 17530 689 17535 691
rect 17524 687 17530 689
rect 17593 688 17594 692
rect 17602 689 17605 691
rect 17291 685 17326 687
rect 17112 680 17124 685
rect 17127 680 17149 685
rect 17211 683 17213 685
rect 17149 676 17162 680
rect 17162 675 17167 676
rect 17176 675 17226 683
rect 17279 682 17291 685
rect 17270 680 17279 682
rect 17331 680 17333 685
rect 17514 684 17522 687
rect 17594 686 17595 687
rect 17507 682 17514 684
rect 17269 676 17270 680
rect 17500 679 17507 682
rect 17595 680 17597 682
rect 17495 678 17500 679
rect 17489 676 17495 678
rect 17597 676 17599 680
rect 17611 678 17618 684
rect 17630 682 17688 701
rect 17715 692 17716 698
rect 17779 692 17780 701
rect 17784 693 17792 703
rect 17799 702 17803 705
rect 17864 702 17889 706
rect 17986 704 17999 706
rect 17787 691 17792 693
rect 17803 692 17814 702
rect 17630 678 17663 682
rect 16925 672 16927 675
rect 17167 674 17226 675
rect 17176 672 17226 674
rect 16632 656 16635 662
rect 16556 643 16620 649
rect 16630 648 16632 656
rect 16676 652 16693 672
rect 16716 666 16723 672
rect 16889 666 16901 672
rect 16911 666 16923 672
rect 17153 666 17176 672
rect 16723 664 16929 666
rect 17142 664 17153 666
rect 16562 637 16589 643
rect 16608 637 16614 643
rect 16624 642 16630 647
rect 16634 642 16643 644
rect 16693 643 16701 652
rect 16870 642 16871 660
rect 15550 623 15577 629
rect 16372 626 16375 630
rect 16565 626 16589 637
rect 16624 635 16643 642
rect 16702 639 16706 642
rect 16706 636 16711 639
rect 16711 635 16719 636
rect 16624 630 16639 635
rect 16719 631 16755 635
rect 16623 626 16639 630
rect 16755 628 16775 631
rect 16869 630 16871 642
rect 16929 654 17088 664
rect 17100 654 17142 664
rect 17266 663 17269 674
rect 17333 663 17336 676
rect 17484 674 17489 676
rect 17481 673 17484 674
rect 17476 672 17481 673
rect 17470 670 17476 672
rect 17599 670 17602 676
rect 17618 671 17626 678
rect 17663 671 17671 678
rect 17688 676 17694 682
rect 17717 679 17718 682
rect 17719 677 17720 687
rect 17771 681 17784 682
rect 17771 679 17780 681
rect 17814 679 17819 692
rect 17864 688 17913 702
rect 17938 698 17984 704
rect 18002 703 18004 706
rect 18014 704 18034 706
rect 18042 704 18061 706
rect 17985 700 18000 702
rect 17930 694 17938 698
rect 17864 687 17889 688
rect 17913 687 17919 688
rect 17921 687 17930 694
rect 17846 678 17864 687
rect 17913 686 17921 687
rect 17919 685 17923 686
rect 17909 677 17916 683
rect 17923 682 17931 685
rect 17931 681 17936 682
rect 17936 680 17941 681
rect 17942 678 17945 679
rect 17713 676 17734 677
rect 17771 676 17777 677
rect 17694 673 17698 676
rect 17451 668 17470 670
rect 17414 664 17451 668
rect 17337 663 17414 664
rect 17228 655 17414 663
rect 17602 660 17615 670
rect 17626 660 17648 671
rect 17671 663 17681 671
rect 17698 663 17702 673
rect 17713 671 17719 676
rect 17720 672 17734 676
rect 17760 671 17777 676
rect 17818 671 17819 676
rect 17829 671 17844 677
rect 17719 665 17725 671
rect 17765 665 17771 671
rect 17809 663 17829 671
rect 17900 669 17909 677
rect 17948 676 17953 678
rect 17954 674 17960 676
rect 16929 652 17100 654
rect 17228 653 17343 655
rect 16929 642 16931 652
rect 17228 651 17340 653
rect 17228 649 17333 651
rect 17228 648 17296 649
rect 17228 645 17280 648
rect 17222 644 17286 645
rect 17200 642 17286 644
rect 16929 634 16935 642
rect 17194 639 17211 642
rect 17222 639 17286 642
rect 17319 641 17331 649
rect 17336 643 17340 651
rect 17176 636 17194 639
rect 16930 630 16935 634
rect 17157 633 17176 636
rect 17228 633 17234 639
rect 17260 636 17266 639
rect 17274 633 17280 639
rect 17338 636 17340 643
rect 17615 642 17661 660
rect 17681 652 17711 663
rect 17691 647 17725 652
rect 17745 647 17746 660
rect 17782 652 17809 663
rect 17818 660 17819 663
rect 17691 646 17762 647
rect 17770 646 17799 652
rect 17691 643 17799 646
rect 17697 642 17702 643
rect 17615 641 17663 642
rect 17142 631 17157 633
rect 16946 630 16986 631
rect 17140 630 17142 631
rect 16785 628 16946 630
rect 16986 628 17015 630
rect 16869 626 16872 628
rect 16928 626 16935 628
rect 15578 623 15605 624
rect 14962 621 14963 622
rect 14866 615 14883 621
rect 14958 616 14962 621
rect 16375 618 16383 626
rect 16443 618 16450 625
rect 16383 617 16443 618
rect 14955 615 14958 616
rect 14883 611 14955 615
rect 16607 610 16623 626
rect 16872 615 16878 626
rect 16925 618 16928 625
rect 17015 622 17076 628
rect 17086 622 17136 630
rect 17336 627 17338 636
rect 16917 615 16925 618
rect 16878 613 16919 615
rect 17260 613 17273 624
rect 17314 616 17336 627
rect 17615 626 17661 641
rect 17665 637 17668 639
rect 17668 636 17670 637
rect 17670 633 17677 636
rect 17697 634 17711 642
rect 17745 634 17746 643
rect 17817 637 17818 653
rect 17859 652 17900 669
rect 17954 668 17962 674
rect 17966 670 17968 672
rect 17998 670 18000 700
rect 18004 690 18012 702
rect 18042 700 18048 704
rect 18088 700 18094 706
rect 18112 693 18123 702
rect 17966 668 18000 670
rect 18004 668 18012 680
rect 18123 678 18126 692
rect 18126 676 18127 678
rect 17962 664 17965 666
rect 17966 656 17978 664
rect 17988 656 18000 664
rect 18127 661 18130 676
rect 17844 646 17859 652
rect 17966 648 17975 656
rect 18129 648 18130 661
rect 17830 641 17842 646
rect 17821 637 17830 641
rect 17677 631 17683 633
rect 17695 630 17711 634
rect 17686 626 17711 630
rect 17745 626 17747 630
rect 17679 622 17704 626
rect 17274 613 17314 616
rect 16885 610 16901 613
rect 16903 610 16919 613
rect 17679 610 17695 622
rect 17704 619 17712 622
rect 17712 618 17721 619
rect 17747 615 17752 626
rect 17779 620 17821 637
rect 17776 619 17779 620
rect 17770 618 17776 619
rect 17808 618 17815 620
rect 17804 615 17808 618
rect 17752 611 17773 615
rect 17795 611 17804 615
rect 17945 606 17969 629
rect 17975 626 18014 648
rect 18014 621 18023 626
rect 18120 622 18129 643
rect 18707 623 18734 629
rect 18735 623 18762 624
rect 18119 621 18120 622
rect 18023 615 18040 621
rect 18115 616 18119 621
rect 18112 615 18115 616
rect 18040 611 18112 615
rect 3676 557 3726 606
rect 3756 557 3822 606
rect 3852 557 3918 606
rect 3948 557 4014 606
rect 4044 557 4094 606
rect 4164 557 4214 606
rect 4244 557 4310 606
rect 4340 557 4406 606
rect 4436 557 4502 606
rect 4532 557 4582 606
rect 4652 557 4702 606
rect 4732 557 4798 606
rect 4828 557 4894 606
rect 4924 557 4990 606
rect 5020 557 5070 606
rect 5140 557 5190 606
rect 5220 557 5286 606
rect 5316 557 5382 606
rect 5412 557 5462 606
rect 6832 557 6882 606
rect 6912 557 6978 606
rect 7008 557 7074 606
rect 7104 557 7170 606
rect 7200 557 7250 606
rect 7320 557 7370 606
rect 7400 557 7466 606
rect 7496 557 7562 606
rect 7592 557 7658 606
rect 7688 557 7738 606
rect 7808 557 7858 606
rect 7888 557 7954 606
rect 7984 557 8050 606
rect 8080 557 8146 606
rect 8176 557 8226 606
rect 8296 557 8346 606
rect 8376 557 8442 606
rect 8472 557 8538 606
rect 8568 557 8618 606
rect 9987 557 10037 606
rect 10067 557 10133 606
rect 10163 557 10229 606
rect 10259 557 10325 606
rect 10355 557 10405 606
rect 10475 557 10525 606
rect 10555 557 10621 606
rect 10651 557 10717 606
rect 10747 557 10813 606
rect 10843 557 10893 606
rect 10963 557 11013 606
rect 11043 557 11109 606
rect 11139 557 11205 606
rect 11235 557 11301 606
rect 11331 557 11381 606
rect 11451 557 11501 606
rect 11531 557 11597 606
rect 11627 557 11693 606
rect 11723 557 11773 606
rect 13144 557 13194 606
rect 13224 557 13290 606
rect 13320 557 13386 606
rect 13416 557 13482 606
rect 13512 557 13562 606
rect 13632 557 13682 606
rect 13712 557 13778 606
rect 13808 557 13874 606
rect 13904 557 13970 606
rect 14000 557 14050 606
rect 14120 557 14170 606
rect 14200 557 14266 606
rect 14296 557 14362 606
rect 14392 557 14458 606
rect 14488 557 14538 606
rect 14608 557 14658 606
rect 14688 557 14754 606
rect 14784 557 14850 606
rect 14880 557 14930 606
rect 16301 557 16351 606
rect 16381 557 16447 606
rect 16477 557 16543 606
rect 16573 557 16639 606
rect 16669 557 16719 606
rect 16789 557 16839 606
rect 16869 557 16935 606
rect 16965 557 17031 606
rect 17061 557 17127 606
rect 17157 557 17207 606
rect 17277 557 17327 606
rect 17357 557 17423 606
rect 17453 557 17519 606
rect 17549 557 17615 606
rect 17645 557 17695 606
rect 17765 557 17815 606
rect 17845 557 17911 606
rect 17941 557 18007 606
rect 18037 557 18087 606
rect 6653 481 6654 487
rect 9809 481 9810 487
rect 12964 481 12965 487
rect 16121 481 16122 487
rect 19278 481 19279 487
rect 6619 441 6654 475
rect 6665 463 6666 475
rect 6665 441 6666 453
rect 9775 441 9810 475
rect 9821 463 9822 475
rect 9821 441 9822 453
rect 12930 441 12965 475
rect 12976 463 12977 475
rect 12976 441 12977 453
rect 16087 441 16122 475
rect 16133 463 16134 475
rect 16133 441 16134 453
rect 19244 441 19279 475
rect 19290 463 19291 475
rect 19290 441 19291 453
rect 5862 429 5863 440
rect 6052 429 6053 440
rect 6138 429 6139 440
rect 6411 429 6412 440
rect 6608 429 6609 440
rect 6642 429 6654 435
rect 9018 429 9019 440
rect 9208 429 9209 440
rect 9294 429 9295 440
rect 9567 429 9568 440
rect 9764 429 9765 440
rect 9798 429 9810 435
rect 12173 429 12174 440
rect 12363 429 12364 440
rect 12449 429 12450 440
rect 12722 429 12723 440
rect 12919 429 12920 440
rect 12953 429 12965 435
rect 15330 429 15331 440
rect 15520 429 15521 440
rect 15606 429 15607 440
rect 15879 429 15880 440
rect 16076 429 16077 440
rect 16110 429 16122 435
rect 18487 429 18488 440
rect 18677 429 18678 440
rect 18763 429 18764 440
rect 19036 429 19037 440
rect 19233 429 19234 440
rect 19267 429 19279 435
rect 5873 389 5874 429
rect 6063 389 6064 429
rect 6149 389 6150 429
rect 6422 389 6423 429
rect 6619 389 6620 429
rect 9029 389 9030 429
rect 9219 389 9220 429
rect 9305 389 9306 429
rect 9578 389 9579 429
rect 9775 389 9776 429
rect 12184 389 12185 429
rect 12374 389 12375 429
rect 12460 389 12461 429
rect 12733 389 12734 429
rect 12930 389 12931 429
rect 15341 389 15342 429
rect 15531 389 15532 429
rect 15617 389 15618 429
rect 15890 389 15891 429
rect 16087 389 16088 429
rect 18498 389 18499 429
rect 18688 389 18689 429
rect 18774 389 18775 429
rect 19047 389 19048 429
rect 19244 389 19245 429
<< nwell >>
rect 3002 1406 4488 1748
rect 13008 1742 13031 1750
rect 4834 1646 4868 1680
rect 7990 1646 8024 1680
rect 11145 1646 11179 1680
rect 14302 1644 14336 1678
rect 17459 1644 17493 1678
rect 3001 1086 19354 1406
rect 3001 1018 4488 1086
rect 3002 820 4488 1018
<< ndiff >>
rect 6620 442 6654 475
rect 9776 442 9810 475
rect 12931 442 12965 475
rect 6623 441 6654 442
rect 9779 441 9810 442
rect 12934 441 12965 442
rect 16088 440 16122 473
rect 19245 440 19279 473
rect 16091 439 16122 440
rect 19248 439 19279 440
<< pdiff >>
rect 4834 1646 4868 1680
rect 7990 1646 8024 1680
rect 11145 1646 11179 1680
rect 14302 1644 14336 1678
rect 17459 1644 17493 1678
<< locali >>
rect 0 2172 19355 2492
rect 3419 1406 3453 1475
rect 12994 1406 13045 1407
rect 1 1086 19354 1406
rect 1 0 19355 320
<< metal1 >>
rect 0 2172 19355 2492
rect 4947 2100 4981 2172
rect 8103 2048 8137 2172
rect 11258 2035 11292 2172
rect 14415 2049 14449 2172
rect 17572 2067 17606 2172
rect 19275 1980 19280 2014
rect 19240 1974 19310 1980
rect 3303 1862 3309 1920
rect 3367 1862 3373 1920
rect 19240 1916 19246 1974
rect 19304 1916 19310 1974
rect 19240 1910 19310 1916
rect 6619 1853 6689 1859
rect 5222 1842 5292 1848
rect 5222 1784 5228 1842
rect 5286 1784 5292 1842
rect 6619 1795 6625 1853
rect 6683 1795 6689 1853
rect 9774 1853 9845 1860
rect 6619 1789 6689 1795
rect 8384 1844 8454 1850
rect 5222 1778 5292 1784
rect 8384 1786 8390 1844
rect 8448 1786 8454 1844
rect 9774 1795 9781 1853
rect 9839 1795 9845 1853
rect 12921 1853 12991 1859
rect 9774 1789 9845 1795
rect 11540 1844 11610 1850
rect 8384 1780 8454 1786
rect 11540 1786 11546 1844
rect 11604 1786 11610 1844
rect 12921 1795 12927 1853
rect 12985 1795 12991 1853
rect 16078 1853 16148 1859
rect 12921 1789 12991 1795
rect 14686 1842 14756 1848
rect 11540 1780 11610 1786
rect 14686 1784 14692 1842
rect 14750 1784 14756 1842
rect 16078 1795 16084 1853
rect 16142 1795 16148 1853
rect 16078 1789 16148 1795
rect 17843 1844 17913 1850
rect 14686 1778 14756 1784
rect 17843 1786 17849 1844
rect 17907 1786 17913 1844
rect 17843 1780 17913 1786
rect 3228 1714 3234 1772
rect 3292 1714 3298 1772
rect 3035 1640 3093 1686
rect 4834 1646 4868 1680
rect 7990 1646 8024 1680
rect 11145 1646 11179 1680
rect 14302 1644 14336 1678
rect 17459 1644 17493 1678
rect 12994 1406 13045 1407
rect 1 1086 19354 1406
rect 6620 441 6654 475
rect 9776 441 9810 475
rect 12931 441 12965 475
rect 16088 439 16122 473
rect 19245 439 19279 473
rect 1 0 19355 320
<< via1 >>
rect 3309 1862 3367 1920
rect 19246 1916 19304 1974
rect 5228 1784 5286 1842
rect 6625 1795 6683 1853
rect 8390 1786 8448 1844
rect 9781 1795 9839 1853
rect 11546 1786 11604 1844
rect 12927 1795 12985 1853
rect 14692 1784 14750 1842
rect 16084 1795 16142 1853
rect 17849 1786 17907 1844
rect 3234 1714 3292 1772
<< metal2 >>
rect 3246 2169 13151 2171
rect 3246 2137 19280 2169
rect 3246 1778 3280 2137
rect 13151 2135 19280 2137
rect 19246 1980 19280 2135
rect 19240 1974 19310 1980
rect 3309 1920 3367 1926
rect 19240 1916 19246 1974
rect 19304 1916 19310 1974
rect 19240 1910 19310 1916
rect 3367 1868 3592 1902
rect 3309 1856 3367 1862
rect 3558 1828 3592 1868
rect 6619 1853 6689 1859
rect 5222 1842 5292 1848
rect 5222 1828 5228 1842
rect 3558 1794 5228 1828
rect 5222 1784 5228 1794
rect 5286 1784 5292 1842
rect 6619 1795 6625 1853
rect 6683 1835 6689 1853
rect 9775 1853 9845 1859
rect 8384 1844 8454 1850
rect 8384 1835 8390 1844
rect 6683 1795 8390 1835
rect 6619 1789 6689 1795
rect 5222 1778 5292 1784
rect 8384 1786 8390 1795
rect 8448 1786 8454 1844
rect 9775 1795 9781 1853
rect 9839 1835 9845 1853
rect 12921 1853 12991 1859
rect 11540 1844 11610 1850
rect 11540 1835 11546 1844
rect 9839 1795 11546 1835
rect 9775 1789 9845 1795
rect 8384 1780 8454 1786
rect 11540 1786 11546 1795
rect 11604 1786 11610 1844
rect 12921 1795 12927 1853
rect 12985 1835 12991 1853
rect 16078 1853 16148 1859
rect 14686 1842 14756 1848
rect 12985 1833 13151 1835
rect 14686 1833 14692 1842
rect 12985 1795 14692 1833
rect 12921 1789 12991 1795
rect 13151 1793 14692 1795
rect 11540 1780 11610 1786
rect 14686 1784 14692 1793
rect 14750 1784 14756 1842
rect 16078 1795 16084 1853
rect 16142 1835 16148 1853
rect 17843 1844 17913 1850
rect 17843 1835 17849 1844
rect 16142 1795 17849 1835
rect 16078 1789 16148 1795
rect 14686 1778 14756 1784
rect 17843 1786 17849 1795
rect 17907 1786 17913 1844
rect 17843 1780 17913 1786
rect 3234 1772 3292 1778
rect 3234 1708 3292 1714
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_0
timestamp 1698882961
transform 1 0 3022 0 -1 2233
box -8 0 552 902
use sky130_osu_single_mpr2aa_8_b0r2  sky130_osu_single_mpr2aa_8_b0r2_0
timestamp 1707510517
transform 1 0 16184 0 1 0
box 0 0 3171 2492
use sky130_osu_single_mpr2aa_8_b0r2  sky130_osu_single_mpr2aa_8_b0r2_1
timestamp 1707510517
transform 1 0 3559 0 1 0
box 0 0 3171 2492
use sky130_osu_single_mpr2aa_8_b0r2  sky130_osu_single_mpr2aa_8_b0r2_2
timestamp 1707510517
transform 1 0 6715 0 1 0
box 0 0 3171 2492
use sky130_osu_single_mpr2aa_8_b0r2  sky130_osu_single_mpr2aa_8_b0r2_3
timestamp 1707510517
transform 1 0 9870 0 1 0
box 0 0 3171 2492
use sky130_osu_single_mpr2aa_8_b0r2  sky130_osu_single_mpr2aa_8_b0r2_4
timestamp 1707510517
transform 1 0 13027 0 1 0
box 0 0 3171 2492
<< labels >>
flabel metal1 s 3035 1640 3093 1686 0 FreeSans 100 0 0 0 start
port 13 nsew signal input
flabel metal1 s 4834 1646 4868 1680 0 FreeSans 100 0 0 0 s1
port 1 nsew signal input
flabel metal1 s 7990 1646 8024 1680 0 FreeSans 100 0 0 0 s2
port 2 nsew signal input
flabel metal1 s 11145 1646 11179 1680 0 FreeSans 100 0 0 0 s3
port 3 nsew signal input
flabel metal1 s 14302 1644 14336 1678 0 FreeSans 100 0 0 0 s4
port 4 nsew signal input
flabel metal1 s 17459 1644 17493 1678 0 FreeSans 100 0 0 0 s5
port 5 nsew signal input
flabel metal1 s 6620 441 6654 475 0 FreeSans 100 0 0 0 X1_Y1
port 6 nsew signal output
flabel metal1 s 9776 441 9810 475 0 FreeSans 100 0 0 0 X2_Y1
port 7 nsew signal output
flabel metal1 s 12931 441 12965 475 0 FreeSans 100 0 0 0 X3_Y1
port 8 nsew signal output
flabel metal1 s 16088 439 16122 473 0 FreeSans 100 0 0 0 X4_Y1
port 9 nsew signal output
flabel metal1 s 19245 439 19279 473 0 FreeSans 100 0 0 0 X5_Y1
port 10 nsew signal output
flabel metal1 s 0 2172 19355 2492 0 FreeSans 100 0 0 0 vssd1
port 14 nsew ground bidirectional
flabel metal1 s 1 1086 19354 1406 0 FreeSans 100 0 0 0 vccd1
port 15 nsew power bidirectional
flabel metal1 s 1 0 19355 320 0 FreeSans 100 0 0 0 vssd1
port 14 nsew ground bidirectional
<< end >>
