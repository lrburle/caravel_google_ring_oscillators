magic
tech sky130A
magscale 1 2
timestamp 1713889922
<< obsli1 >>
rect 468600 153935 578864 451491
<< obsm1 >>
rect 468600 153904 580230 451491
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< obsm2 >>
rect 469022 154022 580226 451491
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
<< obsm3 >>
rect 469026 444988 583520 451491
rect 469026 444588 583440 444988
rect 469026 431796 583520 444588
rect 469026 431396 583440 431796
rect 469026 418468 583520 431396
rect 469026 418068 583440 418468
rect 469026 405140 583520 418068
rect 469026 404740 583440 405140
rect 469026 391948 583520 404740
rect 469026 391548 583440 391948
rect 469026 378620 583520 391548
rect 469026 378220 583440 378620
rect 469026 365292 583520 378220
rect 469026 364892 583440 365292
rect 469026 352100 583520 364892
rect 469026 351700 583440 352100
rect 469026 338772 583520 351700
rect 469026 338372 583440 338772
rect 469026 325444 583520 338372
rect 469026 325044 583440 325444
rect 469026 312252 583520 325044
rect 469026 311852 583440 312252
rect 469026 298924 583520 311852
rect 469026 298524 583440 298924
rect 469026 285596 583520 298524
rect 469026 285196 583440 285596
rect 469026 272404 583520 285196
rect 469026 272004 583440 272404
rect 469026 259076 583520 272004
rect 469026 258676 583440 259076
rect 469026 245748 583520 258676
rect 469026 245348 583440 245748
rect 469026 232556 583520 245348
rect 469026 232156 583440 232556
rect 469026 219228 583520 232156
rect 469026 218828 583440 219228
rect 469026 205900 583520 218828
rect 469026 205500 583440 205900
rect 469026 192708 583520 205500
rect 469026 192308 583440 192708
rect 469026 179380 583520 192308
rect 469026 178980 583440 179380
rect 469026 166052 583520 178980
rect 469026 165652 583440 166052
rect 469026 152860 583520 165652
rect 469026 152460 583440 152860
rect 469026 139532 583520 152460
rect 469026 139132 583440 139532
rect 469026 126204 583520 139132
rect 469026 125804 583440 126204
rect 469026 113012 583520 125804
rect 469026 112612 583440 113012
rect 469026 99684 583520 112612
rect 469026 99284 583440 99684
rect 469026 86356 583520 99284
rect 469026 85956 583440 86356
rect 469026 73164 583520 85956
rect 469026 72764 583440 73164
rect 469026 59836 583520 72764
rect 469026 59436 583440 59836
rect 469026 46508 583520 59436
rect 469026 46108 583440 46508
rect 469026 33316 583520 46108
rect 469026 32916 583440 33316
rect 469026 19988 583520 32916
rect 469026 19588 583440 19988
rect 469026 6796 583520 19588
rect 469026 6564 583440 6796
<< metal4 >>
rect -8726 -7654 -8106 711590
rect -7766 -6694 -7146 710630
rect -6806 -5734 -6186 709670
rect -5846 -4774 -5226 708710
rect -4886 -3814 -4266 707750
rect -3926 -2854 -3306 706790
rect -2966 -1894 -2346 705830
rect -2006 -934 -1386 704870
rect 994 -7654 1614 711590
rect 2234 -7654 2854 711590
rect 3474 -7654 4094 711590
rect 4714 -7654 5334 711590
rect 5954 -7654 6574 711590
rect 7194 -7654 7814 711590
rect 8434 -7654 9054 711590
rect 9674 -7654 10294 711590
rect 36994 -7654 37614 711590
rect 38234 -7654 38854 711590
rect 39474 -7654 40094 711590
rect 40714 -7654 41334 711590
rect 41954 -7654 42574 711590
rect 43194 -7654 43814 711590
rect 44434 -7654 45054 711590
rect 45674 -7654 46294 711590
rect 72994 -7654 73614 711590
rect 74234 -7654 74854 711590
rect 75474 -7654 76094 711590
rect 76714 -7654 77334 711590
rect 77954 -7654 78574 711590
rect 79194 -7654 79814 711590
rect 80434 -7654 81054 711590
rect 81674 -7654 82294 711590
rect 108994 -7654 109614 711590
rect 110234 -7654 110854 711590
rect 111474 -7654 112094 711590
rect 112714 -7654 113334 711590
rect 113954 -7654 114574 711590
rect 115194 -7654 115814 711590
rect 116434 -7654 117054 711590
rect 117674 -7654 118294 711590
rect 144994 -7654 145614 711590
rect 146234 -7654 146854 711590
rect 147474 -7654 148094 711590
rect 148714 -7654 149334 711590
rect 149954 -7654 150574 711590
rect 151194 -7654 151814 711590
rect 152434 -7654 153054 711590
rect 153674 -7654 154294 711590
rect 180994 -7654 181614 711590
rect 182234 -7654 182854 711590
rect 183474 -7654 184094 711590
rect 184714 -7654 185334 711590
rect 185954 -7654 186574 711590
rect 187194 -7654 187814 711590
rect 188434 -7654 189054 711590
rect 189674 -7654 190294 711590
rect 216994 -7654 217614 711590
rect 218234 -7654 218854 711590
rect 219474 -7654 220094 711590
rect 220714 -7654 221334 711590
rect 221954 -7654 222574 711590
rect 223194 -7654 223814 711590
rect 224434 -7654 225054 711590
rect 225674 -7654 226294 711590
rect 252994 -7654 253614 711590
rect 254234 -7654 254854 711590
rect 255474 -7654 256094 711590
rect 256714 -7654 257334 711590
rect 257954 -7654 258574 711590
rect 259194 -7654 259814 711590
rect 260434 -7654 261054 711590
rect 261674 -7654 262294 711590
rect 288994 -7654 289614 711590
rect 290234 -7654 290854 711590
rect 291474 -7654 292094 711590
rect 292714 -7654 293334 711590
rect 293954 -7654 294574 711590
rect 295194 -7654 295814 711590
rect 296434 -7654 297054 711590
rect 297674 -7654 298294 711590
rect 324994 -7654 325614 711590
rect 326234 -7654 326854 711590
rect 327474 -7654 328094 711590
rect 328714 -7654 329334 711590
rect 329954 -7654 330574 711590
rect 331194 -7654 331814 711590
rect 332434 -7654 333054 711590
rect 333674 -7654 334294 711590
rect 360994 -7654 361614 711590
rect 362234 -7654 362854 711590
rect 363474 -7654 364094 711590
rect 364714 -7654 365334 711590
rect 365954 -7654 366574 711590
rect 367194 -7654 367814 711590
rect 368434 -7654 369054 711590
rect 369674 -7654 370294 711590
rect 396994 -7654 397614 711590
rect 398234 -7654 398854 711590
rect 399474 -7654 400094 711590
rect 400714 -7654 401334 711590
rect 401954 -7654 402574 711590
rect 403194 -7654 403814 711590
rect 404434 -7654 405054 711590
rect 405674 -7654 406294 711590
rect 432994 -7654 433614 711590
rect 434234 -7654 434854 711590
rect 435474 -7654 436094 711590
rect 436714 -7654 437334 711590
rect 437954 -7654 438574 711590
rect 439194 -7654 439814 711590
rect 440434 -7654 441054 711590
rect 441674 -7654 442294 711590
rect 468994 -7654 469614 711590
rect 470234 -7654 470854 711590
rect 471474 -7654 472094 711590
rect 472714 359060 473334 711590
rect 473954 359060 474574 711590
rect 475194 359060 475814 711590
rect 476434 359060 477054 711590
rect 477674 359060 478294 711590
rect 472714 268060 473334 354615
rect 473954 268060 474574 354615
rect 475194 268060 475814 354615
rect 476434 268060 477054 354615
rect 477674 268060 478294 354615
rect 472714 -7654 473334 263615
rect 473954 -7654 474574 263615
rect 475194 -7654 475814 263615
rect 476434 -7654 477054 263615
rect 477674 -7654 478294 263615
rect 504994 -7654 505614 711590
rect 506234 -7654 506854 711590
rect 507474 -7654 508094 711590
rect 508714 -7654 509334 711590
rect 509954 -7654 510574 711590
rect 511194 -7654 511814 711590
rect 512434 -7654 513054 711590
rect 513674 -7654 514294 711590
rect 540994 445572 541614 711590
rect 542234 445572 542854 711590
rect 543474 445572 544094 711590
rect 544714 445572 545334 711590
rect 545954 445572 546574 711590
rect 540994 -7654 541614 279788
rect 542234 -7654 542854 279788
rect 543474 -7654 544094 279788
rect 544714 -7654 545334 279788
rect 545954 -7654 546574 279788
rect 547194 -7654 547814 711590
rect 548434 -7654 549054 711590
rect 549674 -7654 550294 711590
rect 576994 -7654 577614 711590
rect 578234 -7654 578854 711590
rect 579474 -7654 580094 711590
rect 580714 -7654 581334 711590
rect 581954 -7654 582574 711590
rect 585310 -934 585930 704870
rect 586270 -1894 586890 705830
rect 587230 -2854 587850 706790
rect 588190 -3814 588810 707750
rect 589150 -4774 589770 708710
rect 590110 -5734 590730 709670
rect 591070 -6694 591690 710630
rect 592030 -7654 592650 711590
<< obsm4 >>
rect 473675 358980 473874 450261
rect 474654 358980 475114 450261
rect 475894 358980 476354 450261
rect 477134 358980 477594 450261
rect 478374 358980 504914 450261
rect 473675 354695 504914 358980
rect 473675 267980 473874 354695
rect 474654 267980 475114 354695
rect 475894 267980 476354 354695
rect 477134 267980 477594 354695
rect 478374 267980 504914 354695
rect 473675 263695 504914 267980
rect 473675 6563 473874 263695
rect 474654 6563 475114 263695
rect 475894 6563 476354 263695
rect 477134 6563 477594 263695
rect 478374 6563 504914 263695
rect 505694 6563 506154 450261
rect 506934 6563 507394 450261
rect 508174 6563 508634 450261
rect 509414 6563 509874 450261
rect 510654 6563 511114 450261
rect 511894 6563 512354 450261
rect 513134 6563 513594 450261
rect 514374 445492 540914 450261
rect 541694 445492 542154 450261
rect 542934 445492 543394 450261
rect 544174 445492 544634 450261
rect 545414 445492 545874 450261
rect 546654 445492 547114 450261
rect 514374 279868 547114 445492
rect 514374 6563 540914 279868
rect 541694 6563 542154 279868
rect 542934 6563 543394 279868
rect 544174 6563 544634 279868
rect 545414 6563 545874 279868
rect 546654 6563 547114 279868
rect 547894 6563 548354 450261
rect 549134 6563 549365 450261
<< metal5 >>
rect -8726 710970 592650 711590
rect -7766 710010 591690 710630
rect -6806 709050 590730 709670
rect -5846 708090 589770 708710
rect -4886 707130 588810 707750
rect -3926 706170 587850 706790
rect -2966 705210 586890 705830
rect -2006 704250 585930 704870
rect -8726 694746 592650 695366
rect -8726 693506 592650 694126
rect -8726 692266 592650 692886
rect -8726 691026 592650 691646
rect -8726 689786 592650 690406
rect -8726 688546 592650 689166
rect -8726 687306 592650 687926
rect -8726 686066 592650 686686
rect -8726 658746 592650 659366
rect -8726 657506 592650 658126
rect -8726 656266 592650 656886
rect -8726 655026 592650 655646
rect -8726 653786 592650 654406
rect -8726 652546 592650 653166
rect -8726 651306 592650 651926
rect -8726 650066 592650 650686
rect -8726 622746 592650 623366
rect -8726 621506 592650 622126
rect -8726 620266 592650 620886
rect -8726 619026 592650 619646
rect -8726 617786 592650 618406
rect -8726 616546 592650 617166
rect -8726 615306 592650 615926
rect -8726 614066 592650 614686
rect -8726 586746 592650 587366
rect -8726 585506 592650 586126
rect -8726 584266 592650 584886
rect -8726 583026 592650 583646
rect -8726 581786 592650 582406
rect -8726 580546 592650 581166
rect -8726 579306 592650 579926
rect -8726 578066 592650 578686
rect -8726 550746 592650 551366
rect -8726 549506 592650 550126
rect -8726 548266 592650 548886
rect -8726 547026 592650 547646
rect -8726 545786 592650 546406
rect -8726 544546 592650 545166
rect -8726 543306 592650 543926
rect -8726 542066 592650 542686
rect -8726 514746 592650 515366
rect -8726 513506 592650 514126
rect -8726 512266 592650 512886
rect -8726 511026 592650 511646
rect -8726 509786 592650 510406
rect -8726 508546 592650 509166
rect -8726 507306 592650 507926
rect -8726 506066 592650 506686
rect -8726 478746 592650 479366
rect -8726 477506 592650 478126
rect -8726 476266 592650 476886
rect -8726 475026 592650 475646
rect -8726 473786 592650 474406
rect -8726 472546 592650 473166
rect -8726 471306 592650 471926
rect -8726 470066 592650 470686
rect -8726 442746 592650 443366
rect -8726 441506 592650 442126
rect -8726 440266 592650 440886
rect -8726 439026 592650 439646
rect -8726 437786 592650 438406
rect -8726 436546 592650 437166
rect -8726 435306 592650 435926
rect -8726 434066 592650 434686
rect -8726 406746 592650 407366
rect -8726 405506 592650 406126
rect -8726 404266 592650 404886
rect -8726 403026 592650 403646
rect -8726 401786 592650 402406
rect -8726 400546 592650 401166
rect -8726 399306 592650 399926
rect -8726 398066 592650 398686
rect -8726 370746 592650 371366
rect -8726 369506 592650 370126
rect -8726 368266 592650 368886
rect -8726 367026 592650 367646
rect -8726 365786 592650 366406
rect -8726 364546 592650 365166
rect -8726 363306 592650 363926
rect -8726 362066 592650 362686
rect -8726 334746 592650 335366
rect -8726 333506 592650 334126
rect -8726 332266 592650 332886
rect -8726 331026 592650 331646
rect -8726 329786 592650 330406
rect -8726 328546 592650 329166
rect -8726 327306 592650 327926
rect -8726 326066 592650 326686
rect -8726 298746 592650 299366
rect -8726 297506 592650 298126
rect -8726 296266 592650 296886
rect -8726 295026 592650 295646
rect -8726 293786 592650 294406
rect -8726 292546 592650 293166
rect -8726 291306 592650 291926
rect -8726 290066 592650 290686
rect -8726 262746 592650 263366
rect -8726 261506 592650 262126
rect -8726 260266 592650 260886
rect -8726 259026 592650 259646
rect -8726 257786 592650 258406
rect -8726 256546 592650 257166
rect -8726 255306 592650 255926
rect -8726 254066 592650 254686
rect -8726 226746 592650 227366
rect -8726 225506 592650 226126
rect -8726 224266 592650 224886
rect -8726 223026 592650 223646
rect -8726 221786 592650 222406
rect -8726 220546 592650 221166
rect -8726 219306 592650 219926
rect -8726 218066 592650 218686
rect -8726 190746 592650 191366
rect -8726 189506 592650 190126
rect -8726 188266 592650 188886
rect -8726 187026 592650 187646
rect -8726 185786 592650 186406
rect -8726 184546 592650 185166
rect -8726 183306 592650 183926
rect -8726 182066 592650 182686
rect -8726 154746 592650 155366
rect -8726 153506 592650 154126
rect -8726 152266 592650 152886
rect -8726 151026 592650 151646
rect -8726 149786 592650 150406
rect -8726 148546 592650 149166
rect -8726 147306 592650 147926
rect -8726 146066 592650 146686
rect -8726 118746 592650 119366
rect -8726 117506 592650 118126
rect -8726 116266 592650 116886
rect -8726 115026 592650 115646
rect -8726 113786 592650 114406
rect -8726 112546 592650 113166
rect -8726 111306 592650 111926
rect -8726 110066 592650 110686
rect -8726 82746 592650 83366
rect -8726 81506 592650 82126
rect -8726 80266 592650 80886
rect -8726 79026 592650 79646
rect -8726 77786 592650 78406
rect -8726 76546 592650 77166
rect -8726 75306 592650 75926
rect -8726 74066 592650 74686
rect -8726 46746 592650 47366
rect -8726 45506 592650 46126
rect -8726 44266 592650 44886
rect -8726 43026 592650 43646
rect -8726 41786 592650 42406
rect -8726 40546 592650 41166
rect -8726 39306 592650 39926
rect -8726 38066 592650 38686
rect -8726 10746 592650 11366
rect -8726 9506 592650 10126
rect -8726 8266 592650 8886
rect -8726 7026 592650 7646
rect -8726 5786 592650 6406
rect -8726 4546 592650 5166
rect -8726 3306 592650 3926
rect -8726 2066 592650 2686
rect -2006 -934 585930 -314
rect -2966 -1894 586890 -1274
rect -3926 -2854 587850 -2234
rect -4886 -3814 588810 -3194
rect -5846 -4774 589770 -4154
rect -6806 -5734 590730 -5114
rect -7766 -6694 591690 -6074
rect -8726 -7654 592650 -7034
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 528 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 531 nsew signal output
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 994 -7654 1614 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 36994 -7654 37614 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 72994 -7654 73614 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 108994 -7654 109614 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 144994 -7654 145614 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 180994 -7654 181614 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 216994 -7654 217614 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 252994 -7654 253614 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 288994 -7654 289614 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 324994 -7654 325614 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 360994 -7654 361614 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 396994 -7654 397614 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 432994 -7654 433614 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 468994 -7654 469614 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 504994 -7654 505614 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 540994 -7654 541614 279788 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 540994 445572 541614 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 576994 -7654 577614 711590 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 2066 592650 2686 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 38066 592650 38686 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 74066 592650 74686 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 110066 592650 110686 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 146066 592650 146686 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 182066 592650 182686 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 218066 592650 218686 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 254066 592650 254686 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 290066 592650 290686 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 326066 592650 326686 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 362066 592650 362686 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 398066 592650 398686 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 434066 592650 434686 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 470066 592650 470686 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 506066 592650 506686 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 542066 592650 542686 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 578066 592650 578686 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 614066 592650 614686 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 650066 592650 650686 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s -8726 686066 592650 686686 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 3474 -7654 4094 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 39474 -7654 40094 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 75474 -7654 76094 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 111474 -7654 112094 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 147474 -7654 148094 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 183474 -7654 184094 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 219474 -7654 220094 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 255474 -7654 256094 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 291474 -7654 292094 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 327474 -7654 328094 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 363474 -7654 364094 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 399474 -7654 400094 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 435474 -7654 436094 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 471474 -7654 472094 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 507474 -7654 508094 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 543474 -7654 544094 279788 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 543474 445572 544094 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 579474 -7654 580094 711590 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 4546 592650 5166 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 40546 592650 41166 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 76546 592650 77166 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 112546 592650 113166 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 148546 592650 149166 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 184546 592650 185166 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 220546 592650 221166 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 256546 592650 257166 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 292546 592650 293166 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 328546 592650 329166 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 364546 592650 365166 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 400546 592650 401166 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 436546 592650 437166 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 472546 592650 473166 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 508546 592650 509166 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 544546 592650 545166 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 580546 592650 581166 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 616546 592650 617166 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 652546 592650 653166 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s -8726 688546 592650 689166 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 5954 -7654 6574 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 41954 -7654 42574 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 77954 -7654 78574 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 113954 -7654 114574 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 149954 -7654 150574 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 185954 -7654 186574 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 221954 -7654 222574 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 257954 -7654 258574 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 293954 -7654 294574 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 329954 -7654 330574 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 365954 -7654 366574 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 401954 -7654 402574 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 437954 -7654 438574 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 473954 -7654 474574 263615 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 473954 268060 474574 354615 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 473954 359060 474574 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 509954 -7654 510574 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 545954 -7654 546574 279788 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 545954 445572 546574 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 581954 -7654 582574 711590 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 7026 592650 7646 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 43026 592650 43646 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 79026 592650 79646 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 115026 592650 115646 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 151026 592650 151646 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 187026 592650 187646 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 223026 592650 223646 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 259026 592650 259646 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 295026 592650 295646 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 331026 592650 331646 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 367026 592650 367646 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 403026 592650 403646 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 439026 592650 439646 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 475026 592650 475646 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 511026 592650 511646 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 547026 592650 547646 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 583026 592650 583646 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 619026 592650 619646 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 655026 592650 655646 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s -8726 691026 592650 691646 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 8434 -7654 9054 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 44434 -7654 45054 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 80434 -7654 81054 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 116434 -7654 117054 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 152434 -7654 153054 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 188434 -7654 189054 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 224434 -7654 225054 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 260434 -7654 261054 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 296434 -7654 297054 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 332434 -7654 333054 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 368434 -7654 369054 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 404434 -7654 405054 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 440434 -7654 441054 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 476434 -7654 477054 263615 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 476434 268060 477054 354615 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 476434 359060 477054 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 512434 -7654 513054 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 548434 -7654 549054 711590 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 9506 592650 10126 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 45506 592650 46126 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 81506 592650 82126 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 117506 592650 118126 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 153506 592650 154126 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 189506 592650 190126 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 225506 592650 226126 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 261506 592650 262126 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 297506 592650 298126 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 333506 592650 334126 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 369506 592650 370126 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 405506 592650 406126 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 441506 592650 442126 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 477506 592650 478126 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 513506 592650 514126 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 549506 592650 550126 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 585506 592650 586126 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 621506 592650 622126 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 657506 592650 658126 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s -8726 693506 592650 694126 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 7194 -7654 7814 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 43194 -7654 43814 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 79194 -7654 79814 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 115194 -7654 115814 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 151194 -7654 151814 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 187194 -7654 187814 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 223194 -7654 223814 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 259194 -7654 259814 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 295194 -7654 295814 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 331194 -7654 331814 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 367194 -7654 367814 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 403194 -7654 403814 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 439194 -7654 439814 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 475194 -7654 475814 263615 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 475194 268060 475814 354615 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 475194 359060 475814 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 511194 -7654 511814 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 547194 -7654 547814 711590 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 8266 592650 8886 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 44266 592650 44886 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 80266 592650 80886 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 116266 592650 116886 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 152266 592650 152886 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 188266 592650 188886 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 224266 592650 224886 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 260266 592650 260886 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 296266 592650 296886 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 332266 592650 332886 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 368266 592650 368886 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 404266 592650 404886 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 440266 592650 440886 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 476266 592650 476886 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 512266 592650 512886 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 548266 592650 548886 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 584266 592650 584886 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 620266 592650 620886 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 656266 592650 656886 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s -8726 692266 592650 692886 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 9674 -7654 10294 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 45674 -7654 46294 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 81674 -7654 82294 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 117674 -7654 118294 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 153674 -7654 154294 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 189674 -7654 190294 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 225674 -7654 226294 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 261674 -7654 262294 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 297674 -7654 298294 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 333674 -7654 334294 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 369674 -7654 370294 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 405674 -7654 406294 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 441674 -7654 442294 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 477674 -7654 478294 263615 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 477674 268060 478294 354615 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 477674 359060 478294 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 513674 -7654 514294 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 549674 -7654 550294 711590 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 10746 592650 11366 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 46746 592650 47366 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 82746 592650 83366 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 118746 592650 119366 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 154746 592650 155366 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 190746 592650 191366 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 226746 592650 227366 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 262746 592650 263366 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 298746 592650 299366 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 334746 592650 335366 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 370746 592650 371366 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 406746 592650 407366 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 442746 592650 443366 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 478746 592650 479366 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 514746 592650 515366 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 550746 592650 551366 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 586746 592650 587366 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 622746 592650 623366 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 658746 592650 659366 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s -8726 694746 592650 695366 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 2234 -7654 2854 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 38234 -7654 38854 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 74234 -7654 74854 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 110234 -7654 110854 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 146234 -7654 146854 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 182234 -7654 182854 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 218234 -7654 218854 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 254234 -7654 254854 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 290234 -7654 290854 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 326234 -7654 326854 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 362234 -7654 362854 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 398234 -7654 398854 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 434234 -7654 434854 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 470234 -7654 470854 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 506234 -7654 506854 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 542234 -7654 542854 279788 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 542234 445572 542854 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 578234 -7654 578854 711590 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 3306 592650 3926 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 39306 592650 39926 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 75306 592650 75926 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 111306 592650 111926 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 147306 592650 147926 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 183306 592650 183926 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 219306 592650 219926 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 255306 592650 255926 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 291306 592650 291926 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 327306 592650 327926 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 363306 592650 363926 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 399306 592650 399926 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 435306 592650 435926 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 471306 592650 471926 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 507306 592650 507926 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 543306 592650 543926 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 579306 592650 579926 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 615306 592650 615926 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 651306 592650 651926 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s -8726 687306 592650 687926 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 4714 -7654 5334 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 40714 -7654 41334 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 76714 -7654 77334 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 112714 -7654 113334 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 148714 -7654 149334 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 184714 -7654 185334 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 220714 -7654 221334 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 256714 -7654 257334 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 292714 -7654 293334 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 328714 -7654 329334 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 364714 -7654 365334 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 400714 -7654 401334 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 436714 -7654 437334 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 472714 -7654 473334 263615 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 472714 268060 473334 354615 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 472714 359060 473334 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 508714 -7654 509334 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 544714 -7654 545334 279788 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 544714 445572 545334 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 580714 -7654 581334 711590 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 5786 592650 6406 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 41786 592650 42406 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 77786 592650 78406 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 113786 592650 114406 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 149786 592650 150406 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 185786 592650 186406 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 221786 592650 222406 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 257786 592650 258406 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 293786 592650 294406 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 329786 592650 330406 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 365786 592650 366406 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 401786 592650 402406 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 437786 592650 438406 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 473786 592650 474406 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 509786 592650 510406 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 545786 592650 546406 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 581786 592650 582406 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 617786 592650 618406 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 653786 592650 654406 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s -8726 689786 592650 690406 6 vssd2
port 539 nsew ground bidirectional
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 540 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 541 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 542 nsew signal output
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 543 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 544 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 545 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 546 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 547 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 548 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 549 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 550 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 551 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 552 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 553 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 554 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 555 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 556 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 557 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 558 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 559 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 560 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 561 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 562 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 563 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 564 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 565 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 566 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 567 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 568 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 569 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 570 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 571 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 572 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 573 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 574 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 575 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 576 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 577 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 578 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 579 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 580 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 581 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 582 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 583 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 584 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 585 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 586 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 587 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 588 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 589 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 590 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 591 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 592 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 593 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 594 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 595 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 596 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 597 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 598 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 599 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 600 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 601 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 602 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 603 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 604 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 605 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 606 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 607 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 608 nsew signal output
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 609 nsew signal output
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 610 nsew signal output
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 611 nsew signal output
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 612 nsew signal output
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 613 nsew signal output
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 614 nsew signal output
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 615 nsew signal output
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 616 nsew signal output
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 617 nsew signal output
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 618 nsew signal output
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 619 nsew signal output
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 620 nsew signal output
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 621 nsew signal output
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 622 nsew signal output
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 623 nsew signal output
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 624 nsew signal output
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 625 nsew signal output
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 626 nsew signal output
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 627 nsew signal output
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 628 nsew signal output
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 629 nsew signal output
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 630 nsew signal output
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 631 nsew signal output
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 632 nsew signal output
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 633 nsew signal output
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 634 nsew signal output
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 635 nsew signal output
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 636 nsew signal output
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 637 nsew signal output
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 638 nsew signal output
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 639 nsew signal output
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 640 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 641 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 642 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 643 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 644 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 645 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2564114
string GDS_FILE /import/yukari1/lrburle/google_ring_oscillator/caravel/openlane/user_project_wrapper/runs/24_04_23_11_29/results/signoff/user_project_wrapper.magic.gds
string GDS_START 1159662
<< end >>

