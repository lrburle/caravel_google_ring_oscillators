magic
tech sky130A
magscale 1 2
timestamp 1713888380
<< nwell >>
rect 0 1626 702 1748
rect 2147 1645 2337 1748
rect 0 1406 706 1626
rect 2147 1406 2342 1645
rect 2364 1630 2429 1695
rect 0 1405 716 1406
rect 0 1085 764 1405
rect 2130 1380 2352 1406
rect 2130 1376 2914 1380
rect 3273 1376 3318 1748
rect 2130 1193 3318 1376
rect 2104 1086 3318 1193
rect 0 865 706 1085
rect 2120 1058 2342 1086
rect 1697 1029 2342 1058
rect 2120 943 2342 1029
rect 2121 924 2342 943
rect 2101 921 2342 924
rect 2121 901 2342 921
rect 0 861 707 865
rect 2120 861 2342 901
rect 0 743 702 861
rect 2179 744 2342 861
rect 3124 772 3154 807
rect 3273 744 3318 1086
rect 0 742 595 743
<< ndiff >>
rect 3209 442 3244 476
<< psubdiff >>
rect 2367 2172 2379 2206
rect 2505 2172 2580 2206
<< locali >>
rect 1 2177 3318 2491
rect 1 2171 793 2177
rect 743 1700 793 2171
rect 848 1700 903 2177
rect 958 1700 1013 2177
rect 1068 1700 1123 2177
rect 1178 1700 1233 2177
rect 1288 1700 1343 2177
rect 1398 1700 1453 2177
rect 1508 1700 1563 2177
rect 1618 1700 1673 2177
rect 1728 1700 1783 2177
rect 1838 1700 1893 2177
rect 1948 1700 2003 2177
rect 2058 2171 3318 2177
rect 2058 1700 2127 2171
rect 2893 1868 2971 1895
rect 2847 1861 2971 1868
rect 3042 1720 3152 1754
rect 743 1672 2127 1700
rect 3045 1688 3046 1720
rect 743 1671 757 1672
rect 2123 1671 2127 1672
rect 3210 1461 3244 1495
rect 1 1085 764 1405
rect 2130 1380 2352 1406
rect 2130 1376 2914 1380
rect 3282 1376 3318 1406
rect 2130 1193 3318 1376
rect 2104 1086 3318 1193
rect 3210 997 3244 1031
rect 3044 716 3169 750
rect 2847 624 2971 642
rect 693 590 757 619
rect 2123 618 2162 619
rect 2098 615 2162 618
rect 2123 590 2162 615
rect 693 589 963 590
rect 693 586 855 589
rect 693 585 795 586
rect 693 320 745 585
rect 803 320 855 586
rect 907 585 963 589
rect 1014 587 1175 590
rect 1014 585 1071 587
rect 1123 585 1175 587
rect 1224 585 1279 590
rect 1327 585 1383 590
rect 1431 585 1487 590
rect 1535 585 1591 590
rect 911 320 963 585
rect 1019 320 1067 585
rect 1127 320 1175 585
rect 1231 320 1279 585
rect 1335 320 1383 585
rect 1439 320 1487 585
rect 1543 320 1591 585
rect 1639 320 1687 590
rect 1735 320 1783 590
rect 1831 320 1879 590
rect 1927 320 1975 590
rect 2023 320 2071 590
rect 2119 320 2162 590
rect 2893 608 2971 624
rect 1 0 3318 320
<< viali >>
rect 2847 1868 2893 1914
rect 3209 1742 3243 1776
rect 2847 578 2893 624
rect 3210 442 3244 476
<< metal1 >>
rect 1 2177 3318 2491
rect 1 2171 793 2177
rect 289 1720 323 2171
rect 388 1926 462 1935
rect 388 1870 397 1926
rect 453 1870 462 1926
rect 388 1861 462 1870
rect 488 1783 494 1839
rect 550 1783 556 1839
rect 743 1700 793 2171
rect 848 1700 903 2177
rect 958 1700 1013 2177
rect 1068 1700 1123 2177
rect 1178 1700 1233 2177
rect 1288 1700 1343 2177
rect 1398 1700 1453 2177
rect 1508 1700 1563 2177
rect 1618 1700 1673 2177
rect 1728 1700 1783 2177
rect 1838 1700 1893 2177
rect 1948 1700 2003 2177
rect 2058 2171 3318 2177
rect 2058 1700 2127 2171
rect 2835 1915 2905 1920
rect 2687 1914 2905 1915
rect 2687 1908 2847 1914
rect 2699 1902 2847 1908
rect 2653 1881 2847 1902
rect 2653 1868 2699 1881
rect 2835 1868 2847 1881
rect 2893 1868 2905 1914
rect 2835 1862 2905 1868
rect 2732 1846 2797 1853
rect 2732 1794 2739 1846
rect 2791 1794 2797 1846
rect 2732 1788 2797 1794
rect 2572 1772 2636 1778
rect 2572 1720 2578 1772
rect 2630 1720 2636 1772
rect 2572 1713 2636 1720
rect 116 1634 122 1690
rect 178 1680 184 1690
rect 178 1673 185 1680
rect 578 1673 584 1691
rect 178 1646 584 1673
rect 178 1634 184 1646
rect 185 1638 584 1646
rect 578 1635 584 1638
rect 640 1635 646 1691
rect 743 1672 2127 1700
rect 743 1665 757 1672
rect 1036 1467 1064 1672
rect 2114 1665 2127 1672
rect 2364 1688 2429 1695
rect 2364 1636 2371 1688
rect 2423 1636 2429 1688
rect 2364 1630 2429 1636
rect 1 1085 764 1405
rect 2130 1380 2352 1406
rect 2130 1376 2914 1380
rect 3282 1376 3318 1406
rect 2130 1193 3318 1376
rect 2104 1086 3318 1193
rect 2363 1044 2428 1051
rect 2363 992 2370 1044
rect 2422 992 2428 1044
rect 2363 986 2428 992
rect 2121 954 2186 961
rect 2121 924 2128 954
rect 2101 921 2128 924
rect 1933 902 2128 921
rect 2180 902 2186 954
rect 1933 896 2186 902
rect 1933 893 2129 896
rect 2378 846 2414 986
rect 2572 790 2636 796
rect 2572 772 2578 790
rect 2509 738 2578 772
rect 2630 738 2636 790
rect 2572 732 2636 738
rect 2238 716 2303 723
rect 2238 664 2245 716
rect 2297 698 2303 716
rect 2727 716 2797 722
rect 2297 664 2722 698
rect 2238 658 2303 664
rect 2727 658 2733 716
rect 2791 658 2797 716
rect 2727 652 2797 658
rect 693 590 757 625
rect 2123 590 2162 625
rect 2835 624 2905 630
rect 2653 623 2687 624
rect 2699 623 2847 624
rect 2653 590 2847 623
rect 693 589 963 590
rect 693 586 855 589
rect 693 585 795 586
rect 693 320 745 585
rect 803 320 855 586
rect 907 585 963 589
rect 1014 587 1175 590
rect 1014 585 1071 587
rect 1123 585 1175 587
rect 1224 585 1279 590
rect 1327 585 1383 590
rect 1431 585 1487 590
rect 1535 585 1591 590
rect 911 320 963 585
rect 1019 320 1067 585
rect 1127 320 1175 585
rect 1231 320 1279 585
rect 1335 320 1383 585
rect 1439 320 1487 585
rect 1543 320 1591 585
rect 1639 320 1687 590
rect 1735 320 1783 590
rect 1831 320 1879 590
rect 1927 320 1975 590
rect 2023 320 2071 590
rect 2119 320 2162 590
rect 2835 578 2847 590
rect 2893 578 2905 624
rect 2835 572 2905 578
rect 1 0 3318 320
<< via1 >>
rect 397 1870 453 1926
rect 494 1783 550 1839
rect 2739 1794 2791 1846
rect 2578 1720 2630 1772
rect 122 1634 178 1690
rect 584 1635 640 1691
rect 2371 1636 2423 1688
rect 2370 992 2422 1044
rect 2128 902 2180 954
rect 2578 738 2630 790
rect 2245 664 2297 716
rect 2733 658 2791 716
<< metal2 >>
rect 505 1944 2541 1978
rect 388 1926 462 1935
rect 388 1870 397 1926
rect 453 1870 462 1926
rect 388 1861 462 1870
rect 505 1845 539 1944
rect 595 1863 2412 1897
rect 494 1839 550 1845
rect 494 1777 550 1783
rect 122 1690 178 1699
rect 595 1697 629 1863
rect 122 1625 178 1634
rect 584 1691 640 1697
rect 2377 1695 2412 1863
rect 2509 1840 2541 1944
rect 2732 1846 2797 1853
rect 2732 1840 2739 1846
rect 2509 1806 2739 1840
rect 584 1629 640 1635
rect 2364 1688 2429 1695
rect 2364 1636 2371 1688
rect 2423 1636 2429 1688
rect 2364 1630 2429 1636
rect 2377 1051 2412 1630
rect 2363 1044 2428 1051
rect 2363 992 2370 1044
rect 2422 992 2428 1044
rect 2363 986 2428 992
rect 2121 954 2186 961
rect 2121 902 2128 954
rect 2180 939 2186 954
rect 2180 902 2287 939
rect 2121 896 2186 902
rect 2253 723 2287 902
rect 2509 772 2541 1806
rect 2732 1794 2739 1806
rect 2791 1794 2797 1846
rect 2732 1788 2797 1794
rect 2572 1772 2636 1778
rect 2572 1720 2578 1772
rect 2630 1720 2636 1772
rect 2572 1713 2636 1720
rect 2578 1666 2612 1713
rect 2578 1631 2613 1666
rect 2578 1596 2773 1631
rect 2572 790 2636 796
rect 2572 772 2578 790
rect 2509 738 2578 772
rect 2630 738 2636 790
rect 2572 732 2636 738
rect 2238 716 2303 723
rect 2738 722 2773 1596
rect 2238 664 2245 716
rect 2297 664 2303 716
rect 2238 658 2303 664
rect 2727 716 2797 722
rect 2727 658 2733 716
rect 2791 658 2797 716
rect 2727 652 2797 658
<< via2 >>
rect 397 1870 453 1926
rect 122 1634 178 1690
<< metal3 >>
rect 116 1690 184 2491
rect 388 1926 462 1935
rect 388 1870 397 1926
rect 453 1923 462 1926
rect 453 1870 1434 1923
rect 388 1863 1434 1870
rect 388 1861 462 1863
rect 116 1634 122 1690
rect 178 1634 184 1690
rect 116 1625 184 1634
rect 1358 1485 1418 1863
rect 1232 1482 1420 1485
rect 1232 1479 1608 1482
rect 1232 1422 1621 1479
rect 1232 1078 1292 1422
rect 1519 1419 1621 1422
rect 1425 1276 1432 1280
rect 1425 1216 1491 1276
rect 1232 1012 1763 1078
rect 1703 1011 1763 1012
rect 1703 810 1763 872
rect 1699 805 1763 810
use scs130hd_mpr2ca_8  scs130hd_mpr2ca_8_0
timestamp 1713475024
transform 1 0 744 0 1 601
box -38 -60 1418 1148
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_1
timestamp 1713887963
transform 1 0 2891 0 1 260
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_2
timestamp 1713887963
transform 1 0 3089 0 1 260
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_3
timestamp 1713887963
transform 1 0 3089 0 -1 2232
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_4
timestamp 1713887963
transform 1 0 2891 0 -1 2232
box -10 0 199 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_0
timestamp 1713481735
transform 1 0 2342 0 1 260
box -10 0 552 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_1
timestamp 1713481735
transform 1 0 97 0 -1 2231
box -10 0 552 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_2
timestamp 1713481735
transform 1 0 2342 0 -1 2232
box -10 0 552 902
<< labels >>
rlabel via1 2397 1019 2397 1019 1 sel
port 8 n
rlabel metal1 60 291 60 291 1 vssd1
port 5 n
rlabel metal1 63 1349 63 1349 1 vccd1
port 6 n
rlabel via1 536 1810 536 1810 1 in
port 9 n
rlabel metal1 49 2199 49 2199 1 vssd1
port 5 n
rlabel viali 3210 442 3244 476 1 Y1
port 11 n
rlabel viali 3209 1742 3243 1776 1 Y0
port 10 n
<< end >>
