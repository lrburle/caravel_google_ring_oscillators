magic
tech sky130A
magscale 1 2
timestamp 1713455153
<< nwell >>
rect 3041 1446 4334 1748
rect 10236 1747 10281 1749
rect 13550 1747 13586 1750
rect 7071 1635 7127 1691
rect 10388 1636 10444 1692
rect 13705 1637 13761 1693
rect 17021 1637 17077 1693
rect 3041 1407 4335 1446
rect 3041 1085 4393 1407
rect 5762 1086 7715 1406
rect 9079 1086 11032 1406
rect 12396 1086 14349 1406
rect 15713 1086 17666 1406
rect 19029 1086 20217 1406
rect 3041 941 4335 1085
rect 6830 987 6888 1045
rect 10147 987 10205 1045
rect 13464 988 13522 1046
rect 16781 989 16839 1047
rect 20097 989 20155 1047
rect 3042 861 4335 941
rect 3042 743 4334 861
<< ndiff >>
rect 6841 442 6878 476
rect 10158 442 10196 476
rect 13475 443 13512 477
rect 16792 444 16829 478
rect 20108 444 20146 478
rect 13478 442 13511 443
rect 16795 442 16828 444
rect 20111 442 20146 444
<< pdiff >>
rect 3119 1645 3153 1679
rect 3754 1635 3810 1691
rect 7071 1635 7127 1691
rect 10388 1636 10444 1692
rect 13705 1637 13761 1693
rect 17021 1637 17077 1693
<< locali >>
rect 0 2172 20217 2492
rect 3480 1405 3514 1477
rect 0 1085 4393 1405
rect 5762 1086 7715 1406
rect 9079 1086 11032 1406
rect 12396 1102 14349 1406
rect 12367 1086 14349 1102
rect 15713 1096 17666 1406
rect 15682 1086 17666 1096
rect 19029 1094 20217 1406
rect 19000 1086 20217 1094
rect 0 0 20217 320
<< viali >>
rect 3119 1645 3153 1679
rect 6842 442 6876 476
rect 10159 442 10193 476
rect 13476 443 13510 477
rect 16793 444 16827 478
rect 20109 444 20143 478
<< metal1 >>
rect 0 2172 20217 2492
rect 20141 1982 20143 2014
rect 20102 1975 20167 1982
rect 20102 1923 20109 1975
rect 20161 1923 20167 1975
rect 3378 1862 3384 1918
rect 3440 1862 3446 1918
rect 20102 1917 20167 1923
rect 6842 1847 6907 1854
rect 6842 1795 6849 1847
rect 6901 1795 6907 1847
rect 6842 1789 6907 1795
rect 10159 1847 10224 1854
rect 10159 1795 10166 1847
rect 10218 1795 10224 1847
rect 13476 1848 13541 1855
rect 10760 1839 10816 1846
rect 10159 1789 10224 1795
rect 10748 1777 10822 1811
rect 13476 1796 13483 1848
rect 13535 1796 13541 1848
rect 13476 1790 13541 1796
rect 16793 1849 16858 1856
rect 16793 1797 16800 1849
rect 16852 1797 16858 1849
rect 16793 1791 16858 1797
rect 3301 1714 3307 1770
rect 3363 1714 3369 1770
rect 3108 1679 3166 1686
rect 3108 1645 3119 1679
rect 3153 1645 3166 1679
rect 3108 1640 3166 1645
rect 0 1085 4393 1405
rect 5762 1086 7715 1406
rect 9079 1086 11032 1406
rect 12396 1086 14349 1406
rect 15713 1086 17666 1406
rect 19029 1086 20217 1406
rect 13475 442 13511 443
rect 16792 442 16828 444
rect 20108 442 20146 444
rect 0 0 20217 320
<< via1 >>
rect 20109 1923 20161 1975
rect 3384 1862 3440 1918
rect 6849 1795 6901 1847
rect 10166 1795 10218 1847
rect 13483 1796 13535 1848
rect 16800 1797 16852 1849
rect 3307 1714 3363 1770
rect 3754 1635 3810 1691
rect 7071 1635 7127 1691
rect 10388 1636 10444 1692
rect 13705 1637 13761 1693
rect 17021 1637 17077 1693
rect 6830 987 6888 1045
rect 10147 987 10205 1045
rect 13464 988 13522 1046
rect 16781 989 16839 1047
rect 20097 989 20155 1047
<< metal2 >>
rect 3315 2013 20143 2047
rect 3315 1776 3349 2013
rect 20109 1982 20143 2013
rect 20102 1975 20167 1982
rect 3384 1918 3440 1924
rect 3440 1869 3622 1903
rect 3384 1856 3440 1862
rect 3588 1828 3622 1869
rect 17354 1858 17362 1932
rect 20102 1923 20109 1975
rect 20161 1923 20167 1975
rect 20102 1917 20167 1923
rect 10654 1856 10728 1858
rect 13971 1856 14045 1858
rect 6842 1847 6907 1854
rect 3588 1794 4152 1828
rect 6842 1795 6849 1847
rect 6901 1829 6907 1847
rect 10159 1847 10224 1854
rect 6901 1828 7052 1829
rect 6901 1795 7455 1828
rect 6842 1789 6907 1795
rect 7052 1794 7455 1795
rect 10159 1795 10166 1847
rect 10218 1829 10224 1847
rect 13476 1848 13541 1855
rect 10218 1828 10415 1829
rect 10218 1795 10780 1828
rect 10159 1789 10224 1795
rect 10415 1794 10780 1795
rect 13476 1796 13483 1848
rect 13535 1830 13541 1848
rect 14088 1845 14101 1858
rect 17288 1856 17362 1858
rect 14077 1839 14101 1845
rect 16793 1849 16858 1856
rect 13535 1828 13661 1830
rect 13535 1796 14077 1828
rect 13476 1790 13541 1796
rect 13661 1794 14077 1796
rect 16793 1797 16800 1849
rect 16852 1831 16858 1849
rect 16852 1828 16968 1831
rect 16852 1797 17393 1828
rect 16793 1791 16858 1797
rect 16968 1794 17393 1797
rect 14077 1781 14101 1783
rect 3307 1770 3363 1776
rect 3307 1708 3363 1714
<< via2 >>
rect 3754 1635 3810 1691
rect 7071 1635 7127 1691
rect 10388 1636 10444 1692
rect 13705 1637 13761 1693
rect 17021 1637 17077 1693
rect 6830 987 6888 1045
rect 10147 987 10205 1045
rect 13464 988 13522 1046
rect 16781 989 16839 1047
rect 20097 989 20155 1047
<< metal3 >>
rect 3748 1691 3816 2492
rect 7065 1691 7133 2492
rect 10382 1692 10450 2493
rect 13699 1693 13767 2494
rect 17015 1693 17083 2494
rect 6821 0 6897 987
rect 10138 0 10214 987
rect 13455 1 13531 988
rect 16772 2 16848 989
rect 20088 2 20164 989
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_0
timestamp 1713287902
transform 1 0 3083 0 -1 2231
box -10 0 552 902
use sky130_osu_single_mpr2ca_8_b0r2  sky130_osu_single_mpr2ca_8_b0r2_0
timestamp 1713454653
transform 1 0 16899 0 1 2
box 0 0 3318 2492
use sky130_osu_single_mpr2ca_8_b0r2  sky130_osu_single_mpr2ca_8_b0r2_1
timestamp 1713454653
transform 1 0 3632 0 1 0
box 0 0 3318 2492
use sky130_osu_single_mpr2ca_8_b0r2  sky130_osu_single_mpr2ca_8_b0r2_2
timestamp 1713454653
transform 1 0 6949 0 1 0
box 0 0 3318 2492
use sky130_osu_single_mpr2ca_8_b0r2  sky130_osu_single_mpr2ca_8_b0r2_3
timestamp 1713454653
transform 1 0 10266 0 1 1
box 0 0 3318 2492
use sky130_osu_single_mpr2ca_8_b0r2  sky130_osu_single_mpr2ca_8_b0r2_4
timestamp 1713454653
transform 1 0 13583 0 1 2
box 0 0 3318 2492
<< labels >>
flabel metal1 s 3108 1640 3166 1686 0 FreeSans 100 0 0 0 start
port 13 nsew signal input
flabel viali s 6842 442 6876 476 0 FreeSans 100 0 0 0 X1_Y1
port 10 se signal output
flabel viali s 10159 442 10193 476 0 FreeSans 100 0 0 0 X2_Y1
port 9 se signal output
flabel metal1 s 9079 1086 11032 1406 0 FreeSans 100 0 0 0 vccd1
port 14 nsew power bidirectional
flabel metal1 s 12396 1086 14349 1406 0 FreeSans 100 0 0 0 vccd1
port 14 nsew power bidirectional
flabel metal1 s 15713 1086 17666 1406 0 FreeSans 100 0 0 0 vccd1
port 14 nsew power bidirectional
flabel metal1 s 19029 1086 20217 1406 0 FreeSans 100 0 0 0 vccd1
port 14 nsew power bidirectional
flabel metal1 s 5762 1086 7715 1406 0 FreeSans 100 0 0 0 vccd1
port 14 nsew power bidirectional
flabel metal1 s 0 2172 20217 2492 0 FreeSans 100 0 0 0 vssd1
port 15 nsew ground bidirectional
flabel metal1 s 0 0 20217 320 0 FreeSans 100 0 0 0 vssd1
port 15 nsew ground bidirectional
flabel metal1 s 0 1085 4393 1405 0 FreeSans 100 0 0 0 vccd1
port 14 nsew power bidirectional
flabel metal1 s 13716 1647 13750 1681 0 FreeSans 100 0 0 0 s4
port 4 nw signal input
flabel metal1 s 17032 1647 17066 1681 0 FreeSans 100 0 0 0 s5
port 5 nw signal input
flabel metal1 s 10399 1646 10433 1680 0 FreeSans 100 0 0 0 s3
port 3 nw signal input
flabel metal1 s 7082 1645 7116 1679 0 FreeSans 100 0 0 0 s2
port 2 nw signal input
flabel metal1 s 3765 1645 3799 1679 0 FreeSans 100 0 0 0 s1
port 1 nw signal input
flabel viali s 13476 443 13510 477 0 FreeSans 100 0 0 0 X3_Y1
port 8 se signal output
flabel viali s 16793 444 16827 478 0 FreeSans 100 0 0 0 X4_Y1
port 7 se signal output
flabel viali s 20109 444 20143 478 0 FreeSans 100 0 0 0 X5_Y1
port 6 se signal output
<< end >>
