magic
tech sky130A
magscale 1 2
timestamp 1708620448
<< error_s >>
rect 3151 2133 3152 2144
rect 3341 2133 3342 2144
rect 3427 2133 3428 2144
rect 5357 2133 5358 2144
rect 5547 2133 5548 2144
rect 5633 2133 5634 2144
rect 6309 2133 6310 2144
rect 6499 2133 6500 2144
rect 6585 2133 6586 2144
rect 6858 2133 6859 2144
rect 7056 2133 7057 2144
rect 8942 2133 8943 2144
rect 9132 2133 9133 2144
rect 9218 2133 9219 2144
rect 9894 2133 9895 2144
rect 10084 2133 10085 2144
rect 10170 2133 10171 2144
rect 10443 2133 10444 2144
rect 10641 2133 10642 2144
rect 12527 2133 12528 2144
rect 12717 2133 12718 2144
rect 12803 2133 12804 2144
rect 13479 2133 13480 2144
rect 13669 2133 13670 2144
rect 13755 2133 13756 2144
rect 14028 2133 14029 2144
rect 14226 2133 14227 2144
rect 16112 2133 16113 2144
rect 16302 2133 16303 2144
rect 16388 2133 16389 2144
rect 17064 2133 17065 2144
rect 17254 2133 17255 2144
rect 17340 2133 17341 2144
rect 17613 2133 17614 2144
rect 17811 2133 17812 2144
rect 19697 2133 19698 2144
rect 19887 2133 19888 2144
rect 19973 2133 19974 2144
rect 20649 2133 20650 2144
rect 20839 2133 20840 2144
rect 20925 2133 20926 2144
rect 21198 2133 21199 2144
rect 21396 2133 21397 2144
rect 3162 2093 3163 2133
rect 3352 2093 3353 2133
rect 3438 2093 3439 2133
rect 5368 2093 5369 2133
rect 5558 2093 5559 2133
rect 5644 2093 5645 2133
rect 6320 2093 6321 2133
rect 6510 2093 6511 2133
rect 6596 2093 6597 2133
rect 6869 2093 6870 2133
rect 7067 2093 7068 2133
rect 8953 2093 8954 2133
rect 9143 2093 9144 2133
rect 9229 2093 9230 2133
rect 9905 2093 9906 2133
rect 10095 2093 10096 2133
rect 10181 2093 10182 2133
rect 10454 2093 10455 2133
rect 10652 2093 10653 2133
rect 12538 2093 12539 2133
rect 12728 2093 12729 2133
rect 12814 2093 12815 2133
rect 13490 2093 13491 2133
rect 13680 2093 13681 2133
rect 13766 2093 13767 2133
rect 14039 2093 14040 2133
rect 14237 2093 14238 2133
rect 16123 2093 16124 2133
rect 16313 2093 16314 2133
rect 16399 2093 16400 2133
rect 17075 2093 17076 2133
rect 17265 2093 17266 2133
rect 17351 2093 17352 2133
rect 17624 2093 17625 2133
rect 17822 2093 17823 2133
rect 19708 2093 19709 2133
rect 19898 2093 19899 2133
rect 19984 2093 19985 2133
rect 20660 2093 20661 2133
rect 20850 2093 20851 2133
rect 20936 2093 20937 2133
rect 21209 2093 21210 2133
rect 21407 2093 21408 2133
rect 6517 1966 6544 1973
rect 10102 1966 10129 1973
rect 13687 1966 13714 1973
rect 17272 1966 17299 1973
rect 20857 1966 20884 1973
rect 6517 1945 6585 1966
rect 10102 1945 10170 1966
rect 13687 1945 13755 1966
rect 17272 1945 17340 1966
rect 20857 1945 20925 1966
rect 6517 1939 6572 1945
rect 10102 1939 10157 1945
rect 13687 1939 13742 1945
rect 17272 1939 17327 1945
rect 20857 1939 20912 1945
rect 6556 1938 6557 1939
rect 10141 1938 10142 1939
rect 13726 1938 13727 1939
rect 17311 1938 17312 1939
rect 20896 1938 20897 1939
rect 6529 1932 6584 1938
rect 10114 1932 10169 1938
rect 13699 1932 13754 1938
rect 17284 1932 17339 1938
rect 20869 1932 20924 1938
rect 6556 1910 6557 1932
rect 10141 1910 10142 1932
rect 13726 1910 13727 1932
rect 17311 1910 17312 1932
rect 20896 1910 20897 1932
rect 3151 1703 3152 1714
rect 3341 1703 3342 1714
rect 3427 1703 3428 1714
rect 5357 1703 5358 1714
rect 5547 1703 5548 1714
rect 5633 1703 5634 1714
rect 6309 1703 6310 1714
rect 6499 1703 6500 1714
rect 6585 1703 6586 1714
rect 6858 1703 6859 1714
rect 7056 1703 7057 1714
rect 8942 1703 8943 1714
rect 9132 1703 9133 1714
rect 9218 1703 9219 1714
rect 9894 1703 9895 1714
rect 10084 1703 10085 1714
rect 10170 1703 10171 1714
rect 10443 1703 10444 1714
rect 10641 1703 10642 1714
rect 12527 1703 12528 1714
rect 12717 1703 12718 1714
rect 12803 1703 12804 1714
rect 13479 1703 13480 1714
rect 13669 1703 13670 1714
rect 13755 1703 13756 1714
rect 14028 1703 14029 1714
rect 14226 1703 14227 1714
rect 16112 1703 16113 1714
rect 16302 1703 16303 1714
rect 16388 1703 16389 1714
rect 17064 1703 17065 1714
rect 17254 1703 17255 1714
rect 17340 1703 17341 1714
rect 17613 1703 17614 1714
rect 17811 1703 17812 1714
rect 19697 1703 19698 1714
rect 19887 1703 19888 1714
rect 19973 1703 19974 1714
rect 20649 1703 20650 1714
rect 20839 1703 20840 1714
rect 20925 1703 20926 1714
rect 21198 1703 21199 1714
rect 21396 1703 21397 1714
rect 3162 1507 3163 1703
rect 3352 1507 3353 1703
rect 3438 1507 3439 1703
rect 5306 1671 5330 1677
rect 5334 1676 5358 1677
rect 5368 1507 5369 1703
rect 5558 1507 5559 1703
rect 5644 1507 5645 1703
rect 6320 1507 6321 1703
rect 6510 1507 6511 1703
rect 6596 1507 6597 1703
rect 6869 1507 6870 1703
rect 7067 1507 7068 1703
rect 8891 1671 8915 1677
rect 8919 1676 8943 1677
rect 8953 1507 8954 1703
rect 9143 1507 9144 1703
rect 9229 1507 9230 1703
rect 9905 1507 9906 1703
rect 10095 1507 10096 1703
rect 10181 1507 10182 1703
rect 10454 1507 10455 1703
rect 10652 1507 10653 1703
rect 12476 1671 12500 1677
rect 12504 1676 12528 1677
rect 12538 1507 12539 1703
rect 12728 1507 12729 1703
rect 12814 1507 12815 1703
rect 13490 1507 13491 1703
rect 13680 1507 13681 1703
rect 13766 1507 13767 1703
rect 14039 1507 14040 1703
rect 14237 1507 14238 1703
rect 16061 1671 16085 1677
rect 16089 1676 16113 1677
rect 16123 1507 16124 1703
rect 16313 1507 16314 1703
rect 16399 1507 16400 1703
rect 17075 1507 17076 1703
rect 17265 1507 17266 1703
rect 17351 1507 17352 1703
rect 17624 1507 17625 1703
rect 17822 1507 17823 1703
rect 19646 1671 19670 1677
rect 19674 1676 19698 1677
rect 19708 1507 19709 1703
rect 19898 1507 19899 1703
rect 19984 1507 19985 1703
rect 20660 1507 20661 1703
rect 20850 1507 20851 1703
rect 20936 1507 20937 1703
rect 21209 1507 21210 1703
rect 21407 1507 21408 1703
rect 3476 1403 3500 1437
rect 5682 1403 5706 1437
rect 6634 1403 6658 1437
rect 9267 1403 9291 1437
rect 10219 1403 10243 1437
rect 12852 1403 12876 1437
rect 13804 1403 13828 1437
rect 16437 1403 16461 1437
rect 17389 1403 17413 1437
rect 20022 1403 20046 1437
rect 20974 1403 20998 1437
rect 6634 1085 6658 1119
rect 10219 1085 10243 1119
rect 13804 1085 13828 1119
rect 17389 1085 17413 1119
rect 20974 1085 20998 1119
rect 3723 1057 3732 1066
rect 3770 1057 3779 1066
rect 5034 1057 5043 1066
rect 5379 1057 5388 1066
rect 5426 1057 5435 1066
rect 5579 1057 5588 1066
rect 5626 1057 5635 1066
rect 7308 1057 7317 1066
rect 7355 1057 7364 1066
rect 8619 1057 8628 1066
rect 8964 1057 8973 1066
rect 9011 1057 9020 1066
rect 9164 1057 9173 1066
rect 9211 1057 9220 1066
rect 10893 1057 10902 1066
rect 10940 1057 10949 1066
rect 12204 1057 12213 1066
rect 12549 1057 12558 1066
rect 12596 1057 12605 1066
rect 12749 1057 12758 1066
rect 12796 1057 12805 1066
rect 14478 1057 14487 1066
rect 14525 1057 14534 1066
rect 15789 1057 15798 1066
rect 16134 1057 16143 1066
rect 16181 1057 16190 1066
rect 16334 1057 16343 1066
rect 16381 1057 16390 1066
rect 18063 1057 18072 1066
rect 18110 1057 18119 1066
rect 19374 1057 19383 1066
rect 19719 1057 19728 1066
rect 19766 1057 19775 1066
rect 19919 1057 19928 1066
rect 19966 1057 19975 1066
rect 3714 1048 3723 1057
rect 3779 1048 3788 1057
rect 4693 1038 4699 1044
rect 4739 1038 4745 1044
rect 5001 1043 5013 1051
rect 5023 1043 5035 1051
rect 5043 1048 5052 1057
rect 5102 1051 5118 1052
rect 4997 1040 4999 1043
rect 5037 1040 5039 1043
rect 5096 1039 5107 1051
rect 5370 1048 5379 1057
rect 5435 1051 5444 1057
rect 5376 1045 5379 1047
rect 5383 1045 5389 1051
rect 5429 1048 5444 1051
rect 5570 1048 5579 1057
rect 5635 1050 5644 1057
rect 5429 1045 5435 1048
rect 4687 1032 4693 1038
rect 4745 1032 4751 1038
rect 4978 1031 4984 1037
rect 4989 1031 4997 1039
rect 5000 1037 5035 1039
rect 5000 1036 5001 1037
rect 5033 1036 5035 1037
rect 3720 1026 3723 1030
rect 3706 1023 3745 1026
rect 4747 1023 4786 1028
rect 4972 1025 4978 1031
rect 4998 1026 5000 1035
rect 5001 1031 5002 1036
rect 4997 1024 4998 1026
rect 3703 1022 3706 1023
rect 3703 1015 3715 1022
rect 3720 1020 3723 1023
rect 3719 1016 3720 1019
rect 3703 1013 3719 1015
rect 3725 1013 3737 1022
rect 3745 1020 3774 1023
rect 3774 1014 3778 1020
rect 4514 1018 4566 1020
rect 4786 1018 4800 1023
rect 4996 1020 4997 1023
rect 4486 1016 4566 1018
rect 4486 1015 4537 1016
rect 3778 1013 3779 1014
rect 4461 1013 4486 1015
rect 4508 1014 4514 1015
rect 4537 1014 4542 1015
rect 3699 1011 3703 1013
rect 3715 1010 3719 1013
rect 4427 1011 4457 1013
rect 4503 1012 4508 1014
rect 3691 998 3699 1010
rect 3698 988 3699 998
rect 3703 1007 3737 1010
rect 3703 1003 3705 1007
rect 3703 996 3704 1003
rect 3715 1001 3719 1007
rect 3734 1005 3737 1007
rect 3740 1004 3749 1010
rect 3702 994 3704 996
rect 3701 988 3707 994
rect 3712 988 3715 1001
rect 3695 982 3701 988
rect 3698 976 3699 982
rect 3702 962 3703 988
rect 3735 982 3737 1004
rect 3741 998 3749 1004
rect 3779 1001 3788 1010
rect 4310 1005 4324 1007
rect 4336 1005 4427 1011
rect 4499 1007 4503 1012
rect 4310 1004 4336 1005
rect 4310 1003 4324 1004
rect 4304 1002 4324 1003
rect 4345 1002 4350 1005
rect 4495 1002 4499 1007
rect 4542 1005 4559 1014
rect 4559 1004 4561 1005
rect 3747 988 3753 994
rect 3770 992 3779 1001
rect 4295 997 4319 1002
rect 4350 997 4356 1002
rect 4494 1001 4495 1002
rect 4566 1001 4583 1016
rect 4800 1015 4807 1018
rect 4995 1016 4996 1020
rect 4807 1014 4810 1015
rect 4810 1005 4832 1014
rect 4993 1012 4995 1016
rect 5033 1014 5037 1036
rect 5039 1027 5047 1039
rect 5305 1037 5317 1045
rect 5366 1041 5376 1045
rect 5377 1041 5383 1045
rect 5341 1037 5383 1041
rect 5435 1039 5441 1045
rect 5588 1044 5594 1050
rect 5634 1048 5644 1050
rect 7299 1048 7308 1057
rect 7364 1048 7373 1057
rect 5597 1044 5609 1048
rect 5619 1044 5631 1048
rect 5634 1044 5640 1048
rect 5582 1038 5588 1044
rect 5640 1038 5646 1044
rect 8278 1038 8284 1044
rect 8324 1038 8330 1044
rect 8586 1043 8598 1051
rect 8608 1043 8620 1051
rect 8628 1048 8637 1057
rect 8687 1051 8703 1052
rect 8582 1040 8584 1043
rect 8622 1040 8624 1043
rect 8681 1039 8692 1051
rect 8955 1048 8964 1057
rect 9020 1051 9029 1057
rect 8961 1045 8964 1047
rect 8968 1045 8974 1051
rect 9014 1048 9029 1051
rect 9155 1048 9164 1057
rect 9220 1050 9229 1057
rect 9014 1045 9020 1048
rect 5086 1020 5096 1036
rect 5117 1034 5129 1037
rect 5311 1036 5317 1037
rect 5363 1036 5366 1037
rect 5111 1033 5131 1034
rect 5305 1033 5311 1036
rect 5347 1033 5377 1036
rect 5111 1031 5117 1033
rect 5131 1031 5161 1033
rect 5108 1025 5111 1031
rect 5105 1022 5111 1025
rect 5163 1024 5184 1031
rect 5211 1024 5217 1030
rect 4832 1004 4835 1005
rect 4692 1001 4693 1004
rect 3753 982 3759 988
rect 3770 986 3774 992
rect 4282 989 4295 997
rect 4304 993 4319 997
rect 3768 974 3769 979
rect 3926 976 3942 984
rect 4109 976 4125 989
rect 4192 979 4209 989
rect 4268 981 4282 989
rect 4262 979 4268 981
rect 4209 978 4262 979
rect 4293 977 4301 989
rect 4305 987 4310 989
rect 4356 987 4369 997
rect 3926 974 3983 976
rect 3764 957 3768 972
rect 3926 968 3971 974
rect 3983 968 3987 974
rect 3702 944 3709 957
rect 3763 953 3764 956
rect 3762 949 3763 952
rect 3765 944 3779 953
rect 3910 952 3926 968
rect 3987 961 3992 968
rect 4174 952 4180 958
rect 4220 952 4226 958
rect 4293 956 4301 967
rect 4305 958 4307 987
rect 4555 984 4557 1001
rect 4561 999 4583 1001
rect 4561 989 4569 999
rect 4687 992 4692 1001
rect 4835 996 4856 1004
rect 4990 1002 4993 1011
rect 5033 1007 5035 1014
rect 5024 1005 5035 1007
rect 5039 1010 5047 1017
rect 5039 1005 5052 1010
rect 5037 1004 5038 1005
rect 5038 1001 5039 1002
rect 5043 1001 5052 1005
rect 5086 1002 5096 1018
rect 5105 1015 5108 1022
rect 5159 1018 5165 1024
rect 5217 1018 5223 1024
rect 5293 1021 5301 1033
rect 5305 1031 5339 1033
rect 5305 1030 5311 1031
rect 5305 1029 5308 1030
rect 5105 1014 5107 1015
rect 5105 1013 5109 1014
rect 5107 1001 5109 1013
rect 4745 995 4778 996
rect 4856 995 4858 996
rect 4780 993 4786 995
rect 4687 986 4693 992
rect 4745 987 4751 992
rect 4786 991 4790 993
rect 4858 991 4868 995
rect 4988 991 4990 999
rect 5030 993 5043 1001
rect 5105 998 5109 1001
rect 5293 999 5301 1011
rect 5305 1002 5307 1029
rect 5585 1024 5588 1036
rect 5640 1032 5643 1036
rect 8272 1032 8278 1038
rect 8330 1032 8336 1038
rect 5593 1018 5597 1032
rect 5640 1021 5656 1032
rect 8563 1031 8569 1037
rect 8574 1031 8582 1039
rect 8585 1037 8620 1039
rect 8585 1036 8586 1037
rect 8618 1036 8620 1037
rect 7305 1026 7308 1030
rect 5656 1018 5672 1021
rect 5382 1007 5383 1008
rect 5383 1005 5384 1006
rect 5305 1001 5308 1002
rect 5351 1001 5379 1002
rect 5305 999 5317 1001
rect 5351 1000 5377 1001
rect 5035 992 5043 993
rect 5096 991 5100 996
rect 5105 991 5110 998
rect 5305 995 5309 999
rect 5351 998 5373 1000
rect 5379 999 5383 1001
rect 5351 996 5366 998
rect 5305 993 5311 995
rect 5351 994 5367 996
rect 5377 995 5383 999
rect 5386 997 5391 1003
rect 5435 1001 5444 1010
rect 5570 1001 5579 1010
rect 5579 1000 5585 1001
rect 4414 981 4430 984
rect 4432 981 4448 984
rect 4408 978 4428 981
rect 4549 979 4561 984
rect 4685 979 4686 983
rect 4693 980 4699 986
rect 4703 983 4771 987
rect 4790 986 4802 991
rect 4452 974 4453 978
rect 4410 972 4502 974
rect 4549 972 4569 979
rect 4684 974 4685 979
rect 4703 977 4729 983
rect 4739 980 4745 983
rect 4771 977 4784 983
rect 4802 978 4823 986
rect 4868 978 4902 991
rect 5034 988 5035 990
rect 4972 979 4978 985
rect 4988 983 4989 987
rect 5031 985 5034 986
rect 4683 972 4684 974
rect 4721 972 4729 977
rect 4314 963 4410 972
rect 4452 969 4453 972
rect 4411 963 4423 965
rect 4314 960 4411 963
rect 4305 957 4309 958
rect 4314 957 4410 960
rect 4305 956 4314 957
rect 4288 955 4312 956
rect 4316 955 4339 956
rect 4288 953 4307 955
rect 4356 954 4371 957
rect 4281 952 4288 953
rect 4301 952 4302 953
rect 3917 944 3926 952
rect 4168 946 4174 952
rect 4226 946 4232 952
rect 4262 949 4281 952
rect 4349 951 4356 954
rect 4305 950 4316 951
rect 4347 950 4349 951
rect 4240 946 4262 949
rect 4232 945 4254 946
rect 3695 936 3701 942
rect 3709 939 3721 944
rect 3757 942 3765 944
rect 3753 939 3765 942
rect 3915 939 3917 944
rect 4305 943 4317 950
rect 3920 940 3926 941
rect 3920 939 3962 940
rect 3966 939 3972 941
rect 3701 930 3707 936
rect 3721 934 3734 939
rect 3749 936 3759 939
rect 3747 934 3757 936
rect 3913 935 3915 939
rect 3920 936 3931 939
rect 3920 935 3926 936
rect 3962 935 3972 939
rect 3913 934 3920 935
rect 3740 929 3743 934
rect 3747 930 3753 934
rect 3738 926 3740 929
rect 3736 923 3738 926
rect 3910 925 3913 934
rect 3914 929 3920 934
rect 3972 929 3978 935
rect 3979 933 3991 941
rect 4052 934 4058 940
rect 4098 934 4104 940
rect 4368 939 4369 954
rect 4398 952 4408 957
rect 4407 939 4408 952
rect 4453 952 4464 968
rect 4425 942 4433 944
rect 4453 943 4456 952
rect 4494 947 4495 968
rect 4502 965 4574 972
rect 4498 963 4574 965
rect 4502 956 4574 963
rect 4583 962 4584 968
rect 4577 956 4584 962
rect 4623 956 4629 962
rect 4678 956 4683 972
rect 4545 955 4586 956
rect 4571 950 4586 955
rect 4629 950 4635 956
rect 4460 942 4506 944
rect 4415 940 4425 942
rect 4506 940 4514 942
rect 4413 939 4415 940
rect 4514 939 4517 940
rect 3993 932 3995 933
rect 3966 927 3991 929
rect 3908 924 3910 925
rect 3731 914 3736 923
rect 3824 922 3854 924
rect 3904 922 3908 924
rect 3729 907 3731 914
rect 3697 895 3698 905
rect 3727 896 3729 907
rect 3800 906 3824 922
rect 3854 916 3904 922
rect 3989 915 3991 927
rect 3995 917 4003 929
rect 4040 926 4052 934
rect 4104 928 4110 934
rect 4226 926 4229 930
rect 4355 927 4413 939
rect 4456 938 4457 939
rect 4425 930 4437 938
rect 4447 930 4459 938
rect 4350 926 4355 927
rect 4109 922 4111 924
rect 3989 906 3992 915
rect 4028 910 4036 922
rect 4040 920 4058 922
rect 3726 891 3727 895
rect 3725 888 3726 891
rect 3787 886 3800 906
rect 3989 902 3991 906
rect 3974 897 3991 902
rect 3966 896 3991 897
rect 3965 895 3991 896
rect 3995 895 4003 907
rect 3914 886 3920 889
rect 3962 886 3991 895
rect 3994 892 3995 894
rect 4028 888 4036 900
rect 4040 890 4042 920
rect 4111 916 4118 922
rect 4118 914 4121 916
rect 4229 914 4243 926
rect 4336 923 4350 926
rect 4359 924 4368 927
rect 4457 926 4459 930
rect 4517 927 4564 939
rect 4577 935 4586 950
rect 4676 949 4678 956
rect 4694 952 4703 968
rect 4712 955 4721 972
rect 4784 968 4801 977
rect 4823 968 4862 978
rect 4675 946 4676 949
rect 4579 934 4580 935
rect 4629 933 4635 936
rect 4564 926 4569 927
rect 4577 926 4579 933
rect 4635 930 4642 933
rect 4652 930 4664 938
rect 4672 937 4674 942
rect 4694 937 4703 950
rect 4709 946 4712 955
rect 4754 954 4783 964
rect 4801 963 4862 968
rect 4801 957 4823 963
rect 4862 960 4872 963
rect 4747 945 4783 954
rect 4794 952 4803 954
rect 4706 937 4708 942
rect 4665 926 4672 937
rect 4694 934 4706 937
rect 4738 936 4747 945
rect 4754 944 4783 945
rect 4784 945 4803 952
rect 4823 950 4844 957
rect 4872 956 4882 960
rect 4902 956 4959 978
rect 4978 973 4984 979
rect 4989 977 4990 983
rect 5030 979 5036 985
rect 4990 972 4991 977
rect 5024 974 5030 979
rect 5031 974 5034 979
rect 5024 973 5031 974
rect 5030 972 5031 973
rect 4988 968 4991 972
rect 5039 971 5041 991
rect 5100 985 5106 991
rect 5111 988 5112 990
rect 5113 986 5116 987
rect 5116 985 5121 986
rect 5100 984 5156 985
rect 5305 984 5316 993
rect 5351 990 5363 994
rect 5377 993 5391 995
rect 5435 993 5441 999
rect 5579 998 5586 1000
rect 5588 998 5597 1018
rect 5672 1015 5685 1018
rect 6309 1015 6310 1026
rect 6499 1015 6500 1026
rect 6585 1015 6586 1026
rect 6858 1015 6859 1026
rect 7055 1015 7056 1026
rect 7291 1023 7330 1026
rect 8332 1023 8371 1028
rect 8557 1025 8563 1031
rect 8583 1026 8585 1035
rect 8586 1031 8587 1036
rect 8582 1024 8583 1026
rect 7288 1022 7291 1023
rect 7288 1015 7300 1022
rect 7305 1020 7308 1023
rect 7304 1016 7305 1019
rect 5685 1001 5749 1015
rect 5749 998 5759 1001
rect 5379 992 5389 993
rect 5426 992 5435 993
rect 5579 992 5597 998
rect 5640 992 5646 998
rect 5759 992 5804 998
rect 5899 994 5917 995
rect 5887 992 5899 994
rect 5351 986 5369 990
rect 5383 987 5389 992
rect 5429 987 5435 992
rect 5588 991 5594 992
rect 5588 989 5595 991
rect 5596 990 5597 992
rect 5626 991 5629 992
rect 5588 986 5594 989
rect 5596 987 5600 988
rect 5615 987 5626 991
rect 5631 986 5640 992
rect 5759 988 5887 992
rect 5100 983 5165 984
rect 5309 983 5317 984
rect 5117 981 5165 983
rect 5117 979 5129 981
rect 5311 978 5327 983
rect 5332 981 5333 984
rect 5159 972 5165 978
rect 5217 972 5223 978
rect 4988 967 4993 968
rect 5029 967 5030 971
rect 4979 958 4993 967
rect 4882 954 4887 956
rect 4959 955 4978 956
rect 4979 955 4991 958
rect 4887 951 4894 954
rect 4959 951 4991 955
rect 4993 951 4994 957
rect 4894 950 4896 951
rect 4784 944 4796 945
rect 4754 943 4761 944
rect 4803 943 4812 945
rect 4754 942 4759 943
rect 4754 941 4756 942
rect 4754 940 4800 941
rect 4801 940 4812 943
rect 4750 939 4755 940
rect 4762 939 4796 940
rect 4750 938 4796 939
rect 4750 937 4762 938
rect 4699 926 4706 934
rect 4749 931 4762 937
rect 4793 936 4796 938
rect 4800 937 4812 940
rect 4844 943 4914 950
rect 4959 949 4979 951
rect 4982 949 4996 950
rect 4972 948 4996 949
rect 4972 946 4979 948
rect 4982 945 4999 948
rect 5024 946 5029 967
rect 5041 951 5043 968
rect 5165 966 5171 972
rect 5174 967 5177 972
rect 5043 949 5048 950
rect 4844 942 4917 943
rect 4844 939 4914 942
rect 4917 939 4926 942
rect 4982 939 4996 945
rect 4999 943 5009 945
rect 5038 943 5048 949
rect 5177 948 5184 967
rect 5211 966 5223 972
rect 5316 968 5327 978
rect 5351 980 5370 986
rect 5351 973 5388 980
rect 5512 976 5528 984
rect 5590 982 5593 986
rect 5589 976 5590 981
rect 5333 968 5336 972
rect 5217 945 5223 966
rect 5327 953 5339 968
rect 5355 965 5388 973
rect 5472 968 5475 976
rect 5513 975 5528 976
rect 5588 970 5589 975
rect 5631 969 5634 986
rect 5643 972 5744 977
rect 5744 969 5755 972
rect 5786 969 5887 988
rect 5917 980 5939 994
rect 5333 951 5336 953
rect 5339 951 5341 953
rect 4914 937 4946 939
rect 4794 931 4796 936
rect 4807 931 4813 937
rect 4914 934 4978 937
rect 4982 934 4998 939
rect 5009 934 5073 943
rect 5341 942 5361 951
rect 5370 948 5388 965
rect 5468 957 5472 968
rect 5463 955 5468 957
rect 5425 950 5426 953
rect 5186 939 5193 942
rect 5210 939 5250 942
rect 5174 936 5210 939
rect 5157 934 5174 936
rect 4750 930 4762 931
rect 4327 921 4336 923
rect 4315 920 4327 921
rect 4354 920 4359 924
rect 4268 915 4354 920
rect 4256 914 4268 915
rect 4296 914 4315 915
rect 4413 914 4421 926
rect 4425 924 4459 926
rect 4121 913 4251 914
rect 4229 909 4243 913
rect 4285 911 4296 914
rect 4278 907 4284 911
rect 4168 900 4174 906
rect 4174 894 4180 900
rect 4202 892 4215 900
rect 4245 892 4256 907
rect 4270 900 4275 904
rect 4407 901 4416 913
rect 4425 901 4427 924
rect 4040 888 4058 890
rect 4202 889 4211 892
rect 4215 891 4217 892
rect 4257 889 4259 891
rect 4267 889 4276 898
rect 4416 892 4427 901
rect 4457 892 4459 924
rect 4463 914 4471 926
rect 4569 924 4579 926
rect 4636 924 4664 926
rect 4665 924 4676 926
rect 4569 923 4577 924
rect 4574 921 4577 923
rect 4629 921 4630 924
rect 4662 921 4676 924
rect 4495 907 4509 921
rect 4564 910 4574 921
rect 4628 917 4629 921
rect 4564 907 4577 910
rect 4627 907 4628 916
rect 4662 915 4664 921
rect 4665 915 4676 921
rect 4699 924 4707 926
rect 4699 915 4706 924
rect 4707 921 4711 924
rect 4710 918 4716 921
rect 4711 916 4716 918
rect 4662 911 4665 915
rect 4667 914 4676 915
rect 4667 912 4668 914
rect 4509 906 4564 907
rect 4571 904 4577 907
rect 4626 904 4627 906
rect 4629 904 4635 910
rect 4662 906 4664 911
rect 4668 907 4670 912
rect 4670 906 4671 907
rect 4661 904 4664 906
rect 4671 904 4672 906
rect 4577 898 4583 904
rect 4619 902 4622 904
rect 4623 902 4629 904
rect 4618 898 4629 902
rect 4660 901 4661 904
rect 4618 892 4625 898
rect 4659 897 4660 900
rect 4657 894 4659 895
rect 4662 894 4664 904
rect 4630 892 4664 894
rect 4668 901 4676 904
rect 4668 892 4682 901
rect 4657 891 4659 892
rect 4682 890 4685 892
rect 3783 879 3787 885
rect 3909 879 3962 886
rect 3972 883 3978 886
rect 3979 883 3991 886
rect 4046 884 4052 888
rect 3780 875 3783 879
rect 3879 875 3909 879
rect 3920 877 3926 879
rect 3725 871 3726 875
rect 3777 870 3780 874
rect 3841 870 3879 875
rect 3839 869 3841 870
rect 3776 868 3777 869
rect 3837 868 3839 869
rect 3928 868 3930 879
rect 3963 868 3964 879
rect 3966 877 3972 883
rect 4040 882 4052 884
rect 4104 882 4110 888
rect 4040 876 4058 882
rect 4098 876 4104 882
rect 4211 880 4220 889
rect 4257 888 4267 889
rect 4655 888 4657 889
rect 4258 887 4267 888
rect 4258 880 4278 887
rect 4460 885 4461 888
rect 4421 882 4422 884
rect 4630 880 4642 888
rect 4652 882 4664 888
rect 4685 884 4687 890
rect 4689 885 4699 915
rect 4716 912 4729 916
rect 4729 907 4741 912
rect 4744 906 4746 907
rect 4755 906 4762 930
rect 4807 928 4808 931
rect 4930 919 4978 934
rect 4998 932 5073 934
rect 5090 933 5141 934
rect 5143 933 5154 934
rect 5090 932 5151 933
rect 4998 930 5090 932
rect 4746 904 4751 906
rect 4755 904 4807 906
rect 4751 901 4807 904
rect 4755 899 4807 901
rect 4738 889 4747 898
rect 4755 896 4824 899
rect 4755 891 4812 896
rect 4824 892 4849 896
rect 4946 894 4954 919
rect 4978 916 4985 919
rect 4998 918 5014 930
rect 5016 918 5032 930
rect 5137 929 5152 932
rect 5133 927 5137 929
rect 5117 922 5133 927
rect 5143 926 5152 929
rect 5186 926 5193 936
rect 5146 920 5151 922
rect 4964 900 4968 916
rect 4985 914 5016 916
rect 5017 914 5019 918
rect 4985 909 5017 914
rect 5008 907 5025 909
rect 5008 902 5017 907
rect 5025 906 5029 907
rect 4968 896 4969 899
rect 4988 898 5008 902
rect 4749 889 4813 891
rect 4849 890 4861 892
rect 4945 890 4946 893
rect 4747 885 4813 889
rect 4651 880 4664 882
rect 4221 875 4224 880
rect 4265 879 4278 880
rect 3763 864 3776 868
rect 3831 864 3837 868
rect 3757 862 3763 864
rect 3828 862 3831 864
rect 3754 858 3757 862
rect 3821 857 3828 862
rect 3753 856 3754 857
rect 3820 856 3821 857
rect 3752 849 3753 856
rect 3817 849 3820 856
rect 3751 841 3752 849
rect 3819 838 3828 842
rect 3866 838 3875 842
rect 3878 838 3894 854
rect 3896 838 3912 854
rect 3930 838 3934 867
rect 3961 847 3963 867
rect 4224 860 4231 875
rect 4263 873 4278 875
rect 3974 849 3988 854
rect 4070 842 4074 856
rect 3747 804 3751 838
rect 3816 833 3828 838
rect 3862 833 3878 838
rect 3912 837 3928 838
rect 3919 834 3928 837
rect 3810 832 3823 833
rect 3862 832 3884 833
rect 3808 831 3817 832
rect 3808 811 3810 831
rect 3811 826 3817 831
rect 3807 810 3810 811
rect 3808 804 3810 810
rect 3816 820 3817 826
rect 3849 824 3884 832
rect 3849 823 3878 824
rect 3849 822 3897 823
rect 3923 822 3928 834
rect 3849 820 3869 822
rect 3878 820 3897 822
rect 3816 804 3832 820
rect 3862 804 3878 820
rect 3922 812 3923 817
rect 3751 799 3764 804
rect 3781 799 3816 804
rect 3764 797 3781 799
rect 3800 788 3817 799
rect 3878 797 3881 803
rect 3878 795 3882 797
rect 3878 788 3888 795
rect 3808 786 3817 788
rect 3882 786 3888 788
rect 3933 786 3934 828
rect 3958 822 3971 838
rect 4104 833 4108 838
rect 4126 837 4138 845
rect 4192 838 4208 854
rect 4231 842 4240 860
rect 4232 841 4240 842
rect 4244 845 4245 862
rect 4244 843 4248 845
rect 4276 844 4278 873
rect 4279 869 4290 875
rect 4282 863 4290 869
rect 4286 859 4289 863
rect 4422 860 4426 879
rect 4459 866 4460 880
rect 4541 867 4547 873
rect 4587 867 4593 873
rect 4651 870 4655 880
rect 4684 870 4689 884
rect 4747 880 4761 885
rect 4755 871 4761 880
rect 4797 880 4807 885
rect 4797 870 4798 880
rect 4801 879 4807 880
rect 4861 879 4928 890
rect 4944 885 4945 889
rect 4943 881 4944 885
rect 4929 875 4933 879
rect 4933 872 4936 875
rect 4940 871 4943 881
rect 4969 879 4973 896
rect 4983 891 4988 898
rect 5029 892 5086 906
rect 5086 891 5089 892
rect 4980 881 4982 889
rect 5089 888 5103 891
rect 5149 890 5151 920
rect 5155 910 5163 922
rect 5193 914 5198 926
rect 5198 902 5203 914
rect 5223 910 5230 939
rect 5250 936 5256 939
rect 5256 934 5260 936
rect 5337 935 5338 942
rect 5361 939 5367 942
rect 5367 936 5373 939
rect 5260 933 5261 934
rect 5261 927 5264 933
rect 5264 922 5267 927
rect 5267 919 5269 922
rect 5269 916 5270 919
rect 5120 888 5151 890
rect 5155 888 5163 900
rect 5203 899 5204 902
rect 5230 900 5232 910
rect 5270 902 5277 916
rect 5338 910 5342 935
rect 5373 934 5377 936
rect 5388 935 5389 942
rect 5375 933 5381 934
rect 5375 932 5383 933
rect 5389 932 5390 935
rect 5425 934 5440 950
rect 5463 948 5475 955
rect 5462 947 5475 948
rect 5485 947 5497 955
rect 5528 952 5544 968
rect 5459 945 5468 947
rect 5458 943 5459 945
rect 5462 943 5468 945
rect 5501 943 5502 945
rect 5508 943 5514 948
rect 5451 942 5458 943
rect 5462 942 5497 943
rect 5501 942 5514 943
rect 5451 937 5462 942
rect 5463 941 5497 942
rect 5449 934 5455 937
rect 5456 936 5462 937
rect 5496 936 5497 941
rect 5514 936 5520 942
rect 5528 934 5544 950
rect 5581 939 5588 968
rect 5634 956 5635 968
rect 5639 965 5640 969
rect 5755 968 5774 969
rect 5782 968 5786 969
rect 5746 964 5782 968
rect 5832 965 5836 969
rect 5580 934 5581 938
rect 5445 932 5449 934
rect 5383 931 5424 932
rect 5389 918 5406 931
rect 5408 926 5424 931
rect 5442 930 5445 932
rect 5435 926 5442 930
rect 5527 927 5528 931
rect 5579 927 5580 932
rect 5408 918 5435 926
rect 5526 920 5528 927
rect 5578 922 5579 927
rect 5589 922 5597 934
rect 5601 922 5603 956
rect 5639 951 5640 964
rect 5746 960 5794 964
rect 5737 954 5746 960
rect 5634 945 5635 951
rect 5640 936 5641 945
rect 5729 939 5737 954
rect 5775 949 5794 960
rect 5794 948 5796 949
rect 5836 948 5841 965
rect 5939 961 5942 980
rect 5942 954 5943 960
rect 5796 945 5800 948
rect 5841 945 5842 948
rect 5726 936 5729 939
rect 5641 928 5647 934
rect 5642 922 5647 928
rect 5721 928 5733 936
rect 5743 928 5755 936
rect 5800 934 5815 945
rect 5842 934 5846 945
rect 5943 941 5946 954
rect 5945 939 5946 941
rect 5943 934 5945 939
rect 5815 932 5816 934
rect 5816 928 5817 930
rect 5846 929 5848 934
rect 5721 924 5726 928
rect 5759 926 5760 928
rect 5761 924 5764 925
rect 5525 919 5528 920
rect 5389 905 5390 918
rect 5417 916 5435 918
rect 5524 918 5528 919
rect 5524 916 5525 918
rect 5577 916 5578 919
rect 5597 916 5598 921
rect 5411 912 5417 916
rect 5520 909 5524 916
rect 5576 909 5577 916
rect 5598 912 5600 916
rect 5628 913 5635 922
rect 5642 916 5643 922
rect 5621 911 5628 913
rect 5639 911 5643 916
rect 5709 912 5717 924
rect 5721 922 5755 924
rect 5721 921 5724 922
rect 5601 910 5639 911
rect 5390 902 5391 904
rect 5277 899 5279 902
rect 5232 894 5233 899
rect 5279 896 5280 899
rect 5103 885 5114 888
rect 5117 885 5156 888
rect 5114 884 5156 885
rect 4973 872 4975 879
rect 4975 870 4976 872
rect 4977 871 4980 881
rect 5117 879 5156 884
rect 5205 881 5207 889
rect 5139 876 5151 879
rect 5156 874 5178 879
rect 5207 874 5208 881
rect 5192 872 5197 874
rect 4626 868 4627 869
rect 4650 867 4651 870
rect 4535 861 4541 867
rect 4593 861 4599 867
rect 4648 860 4650 867
rect 4289 854 4293 858
rect 4289 853 4304 854
rect 4275 843 4278 844
rect 4244 841 4278 843
rect 4282 841 4290 853
rect 4293 850 4304 853
rect 4426 852 4427 858
rect 4460 854 4461 858
rect 4295 845 4304 850
rect 4298 840 4304 845
rect 4061 831 4138 833
rect 3961 820 3966 822
rect 3958 804 3971 820
rect 3961 787 3966 804
rect 3974 788 3990 799
rect 3810 780 3817 786
rect 3875 785 3888 786
rect 3875 783 3922 785
rect 3850 780 3897 783
rect 3810 777 3823 780
rect 3863 777 3869 780
rect 3875 779 3897 780
rect 3875 777 3884 779
rect 4061 777 4119 831
rect 4136 799 4138 831
rect 4142 821 4150 833
rect 4208 822 4224 838
rect 4278 837 4282 840
rect 4302 838 4304 840
rect 4326 838 4332 844
rect 4372 839 4378 844
rect 4368 838 4380 839
rect 4427 838 4430 850
rect 4462 841 4478 854
rect 4533 852 4541 858
rect 4531 850 4541 852
rect 4645 851 4648 860
rect 4594 848 4604 850
rect 4604 846 4610 848
rect 4643 847 4645 851
rect 4521 845 4529 846
rect 4531 845 4535 846
rect 4461 840 4478 841
rect 4461 838 4465 840
rect 4244 829 4256 837
rect 4266 829 4278 837
rect 4304 832 4384 838
rect 4430 832 4431 837
rect 4244 828 4245 829
rect 4245 818 4247 828
rect 4304 822 4320 832
rect 4326 831 4380 832
rect 4326 827 4378 831
rect 4247 814 4249 818
rect 4249 809 4250 812
rect 4250 805 4251 809
rect 4251 799 4252 803
rect 4252 792 4254 799
rect 4326 793 4346 827
rect 4372 825 4380 827
rect 4378 794 4380 825
rect 4384 815 4392 827
rect 4372 793 4380 794
rect 4384 793 4392 805
rect 4408 804 4416 820
rect 4431 814 4434 829
rect 4446 822 4465 838
rect 4499 833 4508 842
rect 4521 841 4531 845
rect 4533 844 4535 845
rect 4610 844 4617 846
rect 4533 841 4541 844
rect 4617 843 4621 844
rect 4621 842 4626 843
rect 4642 842 4643 844
rect 4638 841 4649 842
rect 4674 841 4684 869
rect 4689 866 4690 869
rect 4690 854 4693 865
rect 4761 860 4766 870
rect 4937 869 4940 870
rect 4936 865 4940 869
rect 4937 860 4940 865
rect 4967 866 4977 870
rect 5197 866 5214 872
rect 5233 871 5237 890
rect 5280 888 5284 896
rect 5388 890 5391 896
rect 5397 891 5408 908
rect 5463 903 5475 909
rect 5575 908 5576 909
rect 5504 903 5520 908
rect 5574 903 5575 908
rect 5621 903 5628 910
rect 5475 902 5504 903
rect 5573 896 5574 899
rect 5456 890 5462 896
rect 5514 890 5520 896
rect 5284 874 5292 888
rect 5386 885 5388 889
rect 5394 886 5397 890
rect 4766 854 4767 860
rect 4936 854 4939 860
rect 4690 852 4696 854
rect 4693 846 4696 852
rect 4758 849 4774 854
rect 4757 848 4771 849
rect 4776 848 4792 854
rect 4694 841 4696 846
rect 4754 845 4757 848
rect 4771 845 4792 848
rect 4749 841 4754 845
rect 4782 842 4794 845
rect 4521 838 4535 841
rect 4641 839 4642 841
rect 4649 840 4684 841
rect 4695 840 4696 841
rect 4747 840 4749 841
rect 4674 839 4722 840
rect 4745 838 4747 840
rect 4761 839 4773 842
rect 4854 841 4870 854
rect 4872 841 4888 854
rect 4934 847 4936 853
rect 4937 852 4939 854
rect 4967 852 4985 866
rect 5208 863 5223 866
rect 4794 840 4795 841
rect 4847 840 4848 841
rect 4766 838 4773 839
rect 4515 834 4529 838
rect 4515 833 4526 834
rect 4490 824 4499 833
rect 4461 820 4465 822
rect 4446 814 4465 820
rect 4434 809 4435 812
rect 4435 799 4437 808
rect 4446 804 4462 814
rect 4521 812 4529 824
rect 4533 814 4535 838
rect 4638 832 4641 838
rect 4593 815 4599 821
rect 4627 818 4645 832
rect 4633 815 4634 818
rect 4587 814 4593 815
rect 4632 814 4633 815
rect 4533 812 4567 814
rect 4576 812 4635 814
rect 4645 813 4651 818
rect 4646 812 4652 813
rect 4465 808 4466 812
rect 4557 809 4567 812
rect 4571 810 4576 812
rect 4548 808 4557 809
rect 4560 808 4566 809
rect 4568 808 4571 810
rect 4587 809 4593 812
rect 4466 804 4467 808
rect 4533 805 4545 808
rect 4548 805 4567 808
rect 4533 804 4546 805
rect 4462 794 4470 804
rect 4493 800 4545 804
rect 4555 800 4567 805
rect 4623 800 4632 811
rect 4635 810 4643 812
rect 4646 810 4657 812
rect 4665 811 4674 838
rect 4696 822 4712 838
rect 4736 832 4744 838
rect 4643 809 4657 810
rect 4659 809 4665 810
rect 4643 808 4665 809
rect 4696 808 4712 820
rect 4765 811 4767 838
rect 4768 837 4773 838
rect 4770 836 4773 837
rect 4795 838 4796 840
rect 4846 838 4847 840
rect 4771 834 4775 836
rect 4776 832 4777 834
rect 4795 832 4808 838
rect 4769 828 4773 830
rect 4646 804 4712 808
rect 4655 800 4696 804
rect 4736 801 4737 804
rect 4462 793 4472 794
rect 4326 792 4378 793
rect 4462 792 4474 793
rect 4254 789 4260 792
rect 4260 784 4267 789
rect 4320 788 4400 792
rect 4438 790 4439 792
rect 4462 789 4483 792
rect 4462 788 4477 789
rect 4320 786 4384 788
rect 4472 786 4477 788
rect 4483 787 4488 789
rect 4488 786 4492 787
rect 4493 786 4544 800
rect 4556 793 4560 800
rect 4618 793 4623 799
rect 4555 790 4556 793
rect 4616 790 4618 793
rect 4267 783 4268 784
rect 4303 783 4304 785
rect 4269 779 4275 783
rect 4300 779 4303 783
rect 4326 780 4332 786
rect 4368 781 4380 786
rect 4488 785 4499 786
rect 4490 783 4499 785
rect 4490 782 4502 783
rect 4372 780 4378 781
rect 4438 779 4439 781
rect 4275 777 4280 779
rect 4299 777 4300 779
rect 3697 755 3698 775
rect 3726 772 3727 775
rect 3817 774 3856 777
rect 3863 774 3875 777
rect 3727 759 3735 772
rect 3819 768 3856 774
rect 3866 768 3875 774
rect 3932 768 3933 777
rect 3727 755 3738 759
rect 3698 749 3699 755
rect 3735 753 3738 755
rect 3736 750 3741 753
rect 3710 747 3739 748
rect 3742 747 3743 749
rect 3692 713 3699 725
rect 3704 716 3705 747
rect 3733 745 3738 747
rect 3737 716 3738 745
rect 3739 738 3750 747
rect 3966 740 3970 777
rect 4275 776 4299 777
rect 4436 775 4438 779
rect 4490 777 4499 782
rect 4505 779 4508 781
rect 4508 777 4527 779
rect 4555 777 4564 786
rect 4586 782 4592 788
rect 4613 786 4616 790
rect 4632 782 4638 788
rect 4650 786 4659 800
rect 4662 788 4678 800
rect 4680 796 4716 800
rect 4737 798 4739 801
rect 4764 800 4765 810
rect 4771 798 4773 828
rect 4777 818 4785 830
rect 4794 822 4808 832
rect 4838 836 4846 838
rect 4900 837 4904 841
rect 4932 839 4934 847
rect 4967 838 4977 852
rect 4985 848 4988 852
rect 5115 842 5121 844
rect 5115 838 5129 842
rect 5161 838 5167 844
rect 5168 838 5184 854
rect 5208 838 5214 863
rect 5223 853 5226 863
rect 5226 846 5228 852
rect 5228 838 5231 845
rect 4838 822 4845 836
rect 4862 826 4874 832
rect 4859 825 4918 826
rect 4922 825 4932 838
rect 4859 823 4867 825
rect 4918 823 4932 825
rect 4939 823 4942 838
rect 4794 820 4797 822
rect 4858 821 4859 823
rect 4737 796 4773 798
rect 4777 796 4785 808
rect 4794 804 4808 820
rect 4850 816 4858 820
rect 4862 818 4869 820
rect 4850 808 4856 816
rect 4862 814 4863 818
rect 4922 816 4947 823
rect 4956 816 4967 837
rect 4988 822 5000 838
rect 5109 832 5115 838
rect 5113 830 5115 832
rect 5117 830 5150 838
rect 5167 832 5173 838
rect 5184 832 5200 838
rect 5214 832 5215 838
rect 5167 830 5200 832
rect 5231 830 5234 838
rect 5237 830 5249 870
rect 5292 863 5297 874
rect 5339 871 5342 885
rect 5376 881 5386 885
rect 5462 884 5468 890
rect 5472 887 5473 890
rect 5482 886 5489 890
rect 5473 883 5476 885
rect 5479 884 5481 885
rect 5508 884 5514 890
rect 5571 888 5573 896
rect 5473 882 5478 883
rect 5374 874 5392 881
rect 5357 870 5374 874
rect 5376 870 5386 874
rect 5297 859 5299 863
rect 5323 838 5339 870
rect 5357 866 5376 870
rect 5355 863 5357 866
rect 5353 859 5355 863
rect 5369 859 5376 866
rect 5351 856 5353 859
rect 5349 854 5351 856
rect 5342 851 5351 854
rect 5342 845 5349 851
rect 5342 839 5346 845
rect 5342 838 5343 839
rect 5299 830 5300 838
rect 5323 830 5342 838
rect 5356 830 5369 859
rect 5386 846 5393 858
rect 5398 848 5399 880
rect 5465 876 5471 879
rect 5462 874 5465 876
rect 5453 869 5462 874
rect 5473 870 5476 882
rect 5510 870 5513 884
rect 5570 881 5571 888
rect 5569 874 5570 881
rect 5446 860 5447 863
rect 5476 860 5478 870
rect 5510 862 5524 870
rect 5566 863 5569 874
rect 5441 848 5446 860
rect 5398 847 5403 848
rect 5398 846 5432 847
rect 5439 846 5444 848
rect 5393 844 5394 846
rect 5438 844 5439 846
rect 5435 842 5437 843
rect 5398 834 5410 841
rect 5420 834 5432 841
rect 5478 830 5489 859
rect 5513 830 5524 862
rect 5565 856 5566 859
rect 5603 856 5621 903
rect 5709 890 5717 902
rect 5721 890 5723 921
rect 5754 920 5755 922
rect 5761 912 5767 924
rect 5817 913 5819 925
rect 5848 924 5864 928
rect 5934 925 5943 934
rect 5926 924 5934 925
rect 5848 913 5926 924
rect 5761 911 5764 912
rect 5764 903 5769 910
rect 5802 905 5864 913
rect 5796 903 5802 905
rect 5755 890 5796 903
rect 5764 888 5769 890
rect 5819 889 5821 905
rect 5717 886 5720 888
rect 5769 886 5770 888
rect 5821 885 5822 888
rect 5720 884 5722 885
rect 5721 883 5723 884
rect 5721 879 5724 883
rect 5770 880 5771 882
rect 5721 878 5725 879
rect 5724 876 5725 878
rect 5771 876 5772 880
rect 5822 876 5823 879
rect 5848 878 5864 905
rect 5725 869 5728 874
rect 5728 863 5730 869
rect 5663 861 5664 862
rect 5730 860 5731 863
rect 5542 851 5558 854
rect 5562 851 5565 856
rect 5601 851 5603 856
rect 5644 854 5656 855
rect 5542 845 5562 851
rect 5599 846 5601 851
rect 5638 847 5656 854
rect 5666 849 5678 855
rect 5666 847 5715 849
rect 5731 848 5735 860
rect 5638 845 5654 847
rect 5667 846 5715 847
rect 5660 845 5667 846
rect 5687 845 5715 846
rect 5542 843 5548 845
rect 5598 843 5599 845
rect 5638 843 5660 845
rect 5715 843 5729 845
rect 5735 844 5736 847
rect 5752 843 5768 854
rect 5540 839 5543 843
rect 5596 839 5598 843
rect 5632 842 5637 843
rect 5632 840 5636 842
rect 5638 841 5678 843
rect 5625 839 5635 840
rect 5638 839 5644 841
rect 5619 838 5624 839
rect 5638 838 5639 839
rect 5526 830 5540 838
rect 5593 836 5596 838
rect 5615 837 5619 838
rect 5606 836 5612 837
rect 5593 834 5606 836
rect 5583 833 5587 834
rect 5577 832 5583 833
rect 5564 830 5577 832
rect 5593 831 5596 834
rect 5105 827 5113 830
rect 5117 828 5120 830
rect 5104 821 5114 827
rect 4793 802 4794 804
rect 4795 800 4797 804
rect 4922 801 4932 816
rect 4934 812 4942 816
rect 4934 804 4943 812
rect 4947 807 4979 816
rect 4988 807 5000 820
rect 5080 807 5104 821
rect 5105 818 5113 821
rect 4943 801 4944 803
rect 4956 801 4967 807
rect 4979 804 5000 807
rect 4680 788 4696 796
rect 4716 795 4721 796
rect 4721 793 4732 795
rect 4739 794 4746 796
rect 4746 793 4752 794
rect 4763 793 4764 796
rect 4732 792 4737 793
rect 4752 792 4772 793
rect 4775 792 4777 795
rect 4792 794 4793 796
rect 4752 786 4773 792
rect 4789 789 4792 793
rect 4774 788 4792 789
rect 4774 786 4789 788
rect 4845 786 4846 788
rect 4850 786 4856 798
rect 4904 789 4905 801
rect 4919 790 4922 800
rect 4944 797 4972 801
rect 4979 797 4998 804
rect 5068 800 5080 807
rect 5066 799 5068 800
rect 4944 796 4998 797
rect 5059 796 5066 799
rect 5105 796 5113 808
rect 5117 796 5119 828
rect 5185 822 5414 830
rect 5185 820 5187 822
rect 5188 820 5414 822
rect 5185 814 5414 820
rect 5442 814 5564 830
rect 5587 818 5593 831
rect 5622 822 5638 838
rect 5585 815 5592 818
rect 5185 812 5442 814
rect 5187 804 5200 812
rect 5217 807 5219 812
rect 5187 803 5188 804
rect 5188 801 5189 802
rect 5185 796 5188 801
rect 5218 800 5219 807
rect 5230 804 5242 812
rect 5242 803 5243 804
rect 5247 803 5249 808
rect 5266 803 5345 812
rect 5243 802 5345 803
rect 5246 799 5262 802
rect 4863 787 4864 788
rect 4862 786 4868 787
rect 4644 782 4650 786
rect 4761 784 4773 786
rect 4435 772 4436 774
rect 4499 772 4527 777
rect 4428 759 4435 772
rect 4499 768 4508 772
rect 4546 768 4555 777
rect 4580 776 4586 782
rect 4638 776 4650 782
rect 4762 776 4763 781
rect 4638 766 4642 773
rect 4794 772 4795 786
rect 4846 783 4847 786
rect 4857 784 4859 785
rect 4903 784 4904 788
rect 4918 787 4919 790
rect 4944 789 4988 796
rect 4998 795 5000 796
rect 5000 792 5007 795
rect 5057 793 5059 796
rect 5156 795 5184 796
rect 5007 789 5011 792
rect 4944 788 4966 789
rect 4968 788 4984 789
rect 5011 788 5013 789
rect 5053 788 5057 793
rect 5168 792 5184 795
rect 5214 793 5218 799
rect 4925 787 4932 788
rect 4940 787 4954 788
rect 5013 787 5016 788
rect 4917 786 4925 787
rect 4912 785 4925 786
rect 4944 785 4954 787
rect 5109 786 5115 792
rect 5167 791 5184 792
rect 5211 791 5214 793
rect 5167 789 5223 791
rect 5244 789 5262 799
rect 5167 788 5184 789
rect 5211 788 5214 789
rect 5223 788 5262 789
rect 5264 788 5345 802
rect 5356 800 5369 812
rect 5432 804 5433 807
rect 5167 786 5173 788
rect 5210 786 5211 788
rect 4909 784 4918 785
rect 4847 780 4859 783
rect 4862 780 4863 781
rect 4871 780 4909 784
rect 4847 779 4906 780
rect 4862 774 4874 779
rect 4793 763 4795 772
rect 4912 763 4918 784
rect 4944 784 4958 785
rect 4418 756 4435 759
rect 4759 756 4762 763
rect 4418 755 4428 756
rect 4418 754 4425 755
rect 4758 754 4759 756
rect 4418 753 4422 754
rect 4407 749 4449 753
rect 4407 748 4434 749
rect 4405 747 4407 748
rect 4449 747 4452 749
rect 4391 745 4405 747
rect 3923 738 3929 740
rect 3966 739 3975 740
rect 3743 735 3761 738
rect 3750 725 3761 735
rect 3923 734 3935 738
rect 3969 734 3975 739
rect 4358 738 4391 745
rect 4352 737 4357 738
rect 3917 728 3923 734
rect 3975 729 3981 734
rect 4329 733 4352 737
rect 4406 735 4414 747
rect 4418 746 4423 747
rect 4323 731 4329 733
rect 4317 729 4319 731
rect 3939 728 4070 729
rect 3923 726 3939 728
rect 3975 727 4278 728
rect 4305 727 4311 729
rect 4316 728 4317 729
rect 4070 726 4071 727
rect 4278 726 4311 727
rect 4314 726 4316 728
rect 3704 714 3708 716
rect 3735 714 3738 716
rect 3704 713 3738 714
rect 3743 713 3761 725
rect 3911 714 3919 726
rect 3923 724 3929 726
rect 3699 711 3700 713
rect 3700 708 3705 711
rect 3738 708 3743 711
rect 3704 707 3716 708
rect 3703 701 3716 707
rect 3726 701 3738 708
rect 3750 707 3761 713
rect 3703 694 3705 701
rect 3761 690 3768 707
rect 3911 692 3919 704
rect 3923 694 3925 724
rect 4072 719 4076 726
rect 4278 723 4313 726
rect 4351 723 4357 729
rect 4076 708 4083 719
rect 4299 717 4305 723
rect 4306 719 4313 723
rect 4357 719 4363 723
rect 4406 719 4414 725
rect 4418 719 4420 746
rect 4747 744 4753 750
rect 4755 744 4758 754
rect 4793 750 4794 763
rect 4899 757 4905 762
rect 4911 757 4912 762
rect 4944 758 4954 784
rect 4958 783 4962 784
rect 5017 783 5023 786
rect 5052 783 5053 786
rect 5115 784 5129 786
rect 5115 783 5121 784
rect 5153 783 5157 784
rect 5024 781 5026 782
rect 5026 780 5029 781
rect 5042 780 5052 783
rect 4971 775 4977 779
rect 4977 772 4982 775
rect 5029 772 5052 780
rect 4983 766 5007 772
rect 5042 769 5074 772
rect 5080 769 5153 783
rect 5161 780 5167 786
rect 5168 784 5169 785
rect 5209 784 5210 786
rect 5244 783 5247 788
rect 5253 787 5345 788
rect 5317 786 5345 787
rect 5294 785 5345 786
rect 5353 785 5356 799
rect 5431 797 5432 801
rect 5478 800 5489 814
rect 5513 804 5524 814
rect 5526 804 5542 814
rect 5579 807 5592 815
rect 5576 805 5592 807
rect 5622 805 5638 820
rect 5676 811 5678 841
rect 5682 831 5690 843
rect 5729 838 5769 843
rect 5772 842 5779 874
rect 5814 840 5822 852
rect 5826 842 5828 874
rect 5858 857 5863 874
rect 5858 842 5860 857
rect 5863 852 5864 856
rect 5826 840 5860 842
rect 5864 840 5872 852
rect 5779 838 5780 840
rect 5866 838 5868 840
rect 5769 837 5784 838
rect 5826 837 5827 838
rect 5778 836 5784 837
rect 5823 836 5825 837
rect 5660 809 5678 811
rect 5682 809 5690 821
rect 5739 805 5749 836
rect 5778 832 5793 836
rect 5781 808 5793 832
rect 5826 828 5838 836
rect 5848 828 5860 836
rect 5866 828 5880 838
rect 5827 820 5829 828
rect 5780 807 5793 808
rect 5565 804 5678 805
rect 5542 803 5678 804
rect 5430 791 5431 796
rect 5429 788 5430 791
rect 5489 789 5492 799
rect 5524 794 5532 800
rect 5542 795 5558 803
rect 5560 799 5678 803
rect 5749 801 5753 805
rect 5779 804 5793 807
rect 5814 815 5829 820
rect 5868 822 5880 828
rect 5868 820 5870 822
rect 5814 804 5830 815
rect 5868 805 5880 820
rect 6320 819 6321 1015
rect 6510 819 6511 1015
rect 6596 819 6597 1015
rect 6869 819 6870 1015
rect 7066 819 7067 1015
rect 7288 1013 7304 1015
rect 7310 1013 7322 1022
rect 7330 1020 7359 1023
rect 7359 1014 7363 1020
rect 8099 1018 8151 1020
rect 8371 1018 8385 1023
rect 8581 1020 8582 1023
rect 8071 1016 8151 1018
rect 8071 1015 8122 1016
rect 7363 1013 7364 1014
rect 8046 1013 8071 1015
rect 8093 1014 8099 1015
rect 8122 1014 8127 1015
rect 7284 1011 7288 1013
rect 7300 1010 7304 1013
rect 8012 1011 8042 1013
rect 8088 1012 8093 1014
rect 7276 998 7284 1010
rect 7283 988 7284 998
rect 7288 1007 7322 1010
rect 7288 1003 7290 1007
rect 7288 996 7289 1003
rect 7300 1001 7304 1007
rect 7319 1005 7322 1007
rect 7325 1004 7334 1010
rect 7287 994 7289 996
rect 7286 988 7292 994
rect 7297 988 7300 1001
rect 7280 982 7286 988
rect 7283 976 7284 982
rect 7287 962 7288 988
rect 7320 982 7322 1004
rect 7326 998 7334 1004
rect 7364 1001 7373 1010
rect 7895 1005 7909 1007
rect 7921 1005 8012 1011
rect 8084 1007 8088 1012
rect 7895 1004 7921 1005
rect 7895 1003 7909 1004
rect 7889 1002 7909 1003
rect 7930 1002 7935 1005
rect 8080 1002 8084 1007
rect 8127 1005 8144 1014
rect 8144 1004 8146 1005
rect 7332 988 7338 994
rect 7355 992 7364 1001
rect 7880 997 7904 1002
rect 7935 997 7941 1002
rect 8079 1001 8080 1002
rect 8151 1001 8168 1016
rect 8385 1015 8392 1018
rect 8580 1016 8581 1020
rect 8392 1014 8395 1015
rect 8395 1005 8417 1014
rect 8578 1012 8580 1016
rect 8618 1014 8622 1036
rect 8624 1027 8632 1039
rect 8890 1037 8902 1045
rect 8951 1041 8961 1045
rect 8962 1041 8968 1045
rect 8926 1037 8968 1041
rect 9020 1039 9026 1045
rect 9173 1044 9179 1050
rect 9219 1048 9229 1050
rect 10884 1048 10893 1057
rect 10949 1048 10958 1057
rect 9182 1044 9194 1048
rect 9204 1044 9216 1048
rect 9219 1044 9225 1048
rect 9167 1038 9173 1044
rect 9225 1038 9231 1044
rect 11863 1038 11869 1044
rect 11909 1038 11915 1044
rect 12171 1043 12183 1051
rect 12193 1043 12205 1051
rect 12213 1048 12222 1057
rect 12272 1051 12288 1052
rect 12167 1040 12169 1043
rect 12207 1040 12209 1043
rect 12266 1039 12277 1051
rect 12540 1048 12549 1057
rect 12605 1051 12614 1057
rect 12546 1045 12549 1047
rect 12553 1045 12559 1051
rect 12599 1048 12614 1051
rect 12740 1048 12749 1057
rect 12805 1050 12814 1057
rect 12599 1045 12605 1048
rect 8671 1020 8681 1036
rect 8702 1034 8714 1037
rect 8896 1036 8902 1037
rect 8948 1036 8951 1037
rect 8696 1033 8716 1034
rect 8890 1033 8896 1036
rect 8932 1033 8962 1036
rect 8696 1031 8702 1033
rect 8716 1031 8746 1033
rect 8693 1025 8696 1031
rect 8690 1022 8696 1025
rect 8748 1024 8769 1031
rect 8796 1024 8802 1030
rect 8417 1004 8420 1005
rect 8277 1001 8278 1004
rect 7338 982 7344 988
rect 7355 986 7359 992
rect 7867 989 7880 997
rect 7889 993 7904 997
rect 7353 974 7354 979
rect 7511 976 7527 984
rect 7694 976 7710 989
rect 7777 979 7794 989
rect 7853 981 7867 989
rect 7847 979 7853 981
rect 7794 978 7847 979
rect 7878 977 7886 989
rect 7890 987 7895 989
rect 7941 987 7954 997
rect 7511 974 7568 976
rect 7349 957 7353 972
rect 7511 968 7556 974
rect 7568 968 7572 974
rect 7287 944 7294 957
rect 7348 953 7349 956
rect 7347 949 7348 952
rect 7350 944 7364 953
rect 7495 952 7511 968
rect 7572 961 7577 968
rect 7759 952 7765 958
rect 7805 952 7811 958
rect 7878 956 7886 967
rect 7890 958 7892 987
rect 8140 984 8142 1001
rect 8146 999 8168 1001
rect 8146 989 8154 999
rect 8272 992 8277 1001
rect 8420 996 8441 1004
rect 8575 1002 8578 1011
rect 8618 1007 8620 1014
rect 8609 1005 8620 1007
rect 8624 1010 8632 1017
rect 8624 1005 8637 1010
rect 8622 1004 8623 1005
rect 8623 1001 8624 1002
rect 8628 1001 8637 1005
rect 8671 1002 8681 1018
rect 8690 1015 8693 1022
rect 8744 1018 8750 1024
rect 8802 1018 8808 1024
rect 8878 1021 8886 1033
rect 8890 1031 8924 1033
rect 8890 1030 8896 1031
rect 8890 1029 8893 1030
rect 8690 1014 8692 1015
rect 8690 1013 8694 1014
rect 8692 1001 8694 1013
rect 8330 995 8363 996
rect 8441 995 8443 996
rect 8365 993 8371 995
rect 8272 986 8278 992
rect 8330 987 8336 992
rect 8371 991 8375 993
rect 8443 991 8453 995
rect 8573 991 8575 999
rect 8615 993 8628 1001
rect 8690 998 8694 1001
rect 8878 999 8886 1011
rect 8890 1002 8892 1029
rect 9170 1024 9173 1036
rect 9225 1032 9228 1036
rect 11857 1032 11863 1038
rect 11915 1032 11921 1038
rect 9178 1018 9182 1032
rect 9225 1021 9241 1032
rect 12148 1031 12154 1037
rect 12159 1031 12167 1039
rect 12170 1037 12205 1039
rect 12170 1036 12171 1037
rect 12203 1036 12205 1037
rect 10890 1026 10893 1030
rect 9241 1018 9257 1021
rect 8967 1007 8968 1008
rect 8968 1005 8969 1006
rect 8890 1001 8893 1002
rect 8936 1001 8964 1002
rect 8890 999 8902 1001
rect 8936 1000 8962 1001
rect 8620 992 8628 993
rect 8681 991 8685 996
rect 8690 991 8695 998
rect 8890 995 8894 999
rect 8936 998 8958 1000
rect 8964 999 8968 1001
rect 8936 996 8951 998
rect 8890 993 8896 995
rect 8936 994 8952 996
rect 8962 995 8968 999
rect 8971 997 8976 1003
rect 9020 1001 9029 1010
rect 9155 1001 9164 1010
rect 9164 1000 9170 1001
rect 7999 981 8015 984
rect 8017 981 8033 984
rect 7993 978 8013 981
rect 8134 979 8146 984
rect 8270 979 8271 983
rect 8278 980 8284 986
rect 8288 983 8356 987
rect 8375 986 8387 991
rect 8037 974 8038 978
rect 7995 972 8087 974
rect 8134 972 8154 979
rect 8269 974 8270 979
rect 8288 977 8314 983
rect 8324 980 8330 983
rect 8356 977 8369 983
rect 8387 978 8408 986
rect 8453 978 8487 991
rect 8619 988 8620 990
rect 8557 979 8563 985
rect 8573 983 8574 987
rect 8616 985 8619 986
rect 8268 972 8269 974
rect 8306 972 8314 977
rect 7899 963 7995 972
rect 8037 969 8038 972
rect 7996 963 8008 965
rect 7899 960 7996 963
rect 7890 957 7894 958
rect 7899 957 7995 960
rect 7890 956 7899 957
rect 7873 955 7897 956
rect 7901 955 7924 956
rect 7873 953 7892 955
rect 7941 954 7956 957
rect 7866 952 7873 953
rect 7886 952 7887 953
rect 7502 944 7511 952
rect 7753 946 7759 952
rect 7811 946 7817 952
rect 7847 949 7866 952
rect 7934 951 7941 954
rect 7890 950 7901 951
rect 7932 950 7934 951
rect 7825 946 7847 949
rect 7817 945 7839 946
rect 7280 936 7286 942
rect 7294 939 7306 944
rect 7342 942 7350 944
rect 7338 939 7350 942
rect 7500 939 7502 944
rect 7890 943 7902 950
rect 7505 940 7511 941
rect 7505 939 7547 940
rect 7551 939 7557 941
rect 7286 930 7292 936
rect 7306 934 7319 939
rect 7334 936 7344 939
rect 7332 934 7342 936
rect 7498 935 7500 939
rect 7505 936 7516 939
rect 7505 935 7511 936
rect 7547 935 7557 939
rect 7498 934 7505 935
rect 7325 929 7328 934
rect 7332 930 7338 934
rect 7323 926 7325 929
rect 7321 923 7323 926
rect 7495 925 7498 934
rect 7499 929 7505 934
rect 7557 929 7563 935
rect 7564 933 7576 941
rect 7637 934 7643 940
rect 7683 934 7689 940
rect 7953 939 7954 954
rect 7983 952 7993 957
rect 7992 939 7993 952
rect 8038 952 8049 968
rect 8010 942 8018 944
rect 8038 943 8041 952
rect 8079 947 8080 968
rect 8087 965 8159 972
rect 8083 963 8159 965
rect 8087 956 8159 963
rect 8168 962 8169 968
rect 8162 956 8169 962
rect 8208 956 8214 962
rect 8263 956 8268 972
rect 8130 955 8171 956
rect 8156 950 8171 955
rect 8214 950 8220 956
rect 8045 942 8091 944
rect 8000 940 8010 942
rect 8091 940 8099 942
rect 7998 939 8000 940
rect 8099 939 8102 940
rect 7578 932 7580 933
rect 7551 927 7576 929
rect 7493 924 7495 925
rect 7316 914 7321 923
rect 7409 922 7439 924
rect 7489 922 7493 924
rect 7314 907 7316 914
rect 7282 895 7283 905
rect 7312 896 7314 907
rect 7385 906 7409 922
rect 7439 916 7489 922
rect 7574 915 7576 927
rect 7580 917 7588 929
rect 7625 926 7637 934
rect 7689 928 7695 934
rect 7811 926 7814 930
rect 7940 927 7998 939
rect 8041 938 8042 939
rect 8010 930 8022 938
rect 8032 930 8044 938
rect 7935 926 7940 927
rect 7694 922 7696 924
rect 7574 906 7577 915
rect 7613 910 7621 922
rect 7625 920 7643 922
rect 7311 891 7312 895
rect 7310 888 7311 891
rect 7372 886 7385 906
rect 7574 902 7576 906
rect 7559 897 7576 902
rect 7551 896 7576 897
rect 7550 895 7576 896
rect 7580 895 7588 907
rect 7499 886 7505 889
rect 7547 886 7576 895
rect 7579 892 7580 894
rect 7613 888 7621 900
rect 7625 890 7627 920
rect 7696 916 7703 922
rect 7703 914 7706 916
rect 7814 914 7828 926
rect 7921 923 7935 926
rect 7944 924 7953 927
rect 8042 926 8044 930
rect 8102 927 8149 939
rect 8162 935 8171 950
rect 8261 949 8263 956
rect 8279 952 8288 968
rect 8297 955 8306 972
rect 8369 968 8386 977
rect 8408 968 8447 978
rect 8260 946 8261 949
rect 8164 934 8165 935
rect 8214 933 8220 936
rect 8149 926 8154 927
rect 8162 926 8164 933
rect 8220 930 8227 933
rect 8237 930 8249 938
rect 8257 937 8259 942
rect 8279 937 8288 950
rect 8294 946 8297 955
rect 8339 954 8368 964
rect 8386 963 8447 968
rect 8386 957 8408 963
rect 8447 960 8457 963
rect 8332 945 8368 954
rect 8379 952 8388 954
rect 8291 937 8293 942
rect 8250 926 8257 937
rect 8279 934 8291 937
rect 8323 936 8332 945
rect 8339 944 8368 945
rect 8369 945 8388 952
rect 8408 950 8429 957
rect 8457 956 8467 960
rect 8487 956 8544 978
rect 8563 973 8569 979
rect 8574 977 8575 983
rect 8615 979 8621 985
rect 8575 972 8576 977
rect 8609 974 8615 979
rect 8616 974 8619 979
rect 8609 973 8616 974
rect 8615 972 8616 973
rect 8573 968 8576 972
rect 8624 971 8626 991
rect 8685 985 8691 991
rect 8696 988 8697 990
rect 8698 986 8701 987
rect 8701 985 8706 986
rect 8685 984 8741 985
rect 8890 984 8901 993
rect 8936 990 8948 994
rect 8962 993 8976 995
rect 9020 993 9026 999
rect 9164 998 9171 1000
rect 9173 998 9182 1018
rect 9257 1015 9270 1018
rect 9894 1015 9895 1026
rect 10084 1015 10085 1026
rect 10170 1015 10171 1026
rect 10443 1015 10444 1026
rect 10640 1015 10641 1026
rect 10876 1023 10915 1026
rect 11917 1023 11956 1028
rect 12142 1025 12148 1031
rect 12168 1026 12170 1035
rect 12171 1031 12172 1036
rect 12167 1024 12168 1026
rect 10873 1022 10876 1023
rect 10873 1015 10885 1022
rect 10890 1020 10893 1023
rect 10889 1016 10890 1019
rect 9270 1001 9334 1015
rect 9334 998 9344 1001
rect 8964 992 8974 993
rect 9011 992 9020 993
rect 9164 992 9182 998
rect 9225 992 9231 998
rect 9344 992 9389 998
rect 9484 994 9502 995
rect 9472 992 9484 994
rect 8936 986 8954 990
rect 8968 987 8974 992
rect 9014 987 9020 992
rect 9173 991 9179 992
rect 9173 989 9180 991
rect 9181 990 9182 992
rect 9211 991 9214 992
rect 9173 986 9179 989
rect 9181 987 9185 988
rect 9200 987 9211 991
rect 9216 986 9225 992
rect 9344 988 9472 992
rect 8685 983 8750 984
rect 8894 983 8902 984
rect 8702 981 8750 983
rect 8702 979 8714 981
rect 8896 978 8912 983
rect 8917 981 8918 984
rect 8744 972 8750 978
rect 8802 972 8808 978
rect 8573 967 8578 968
rect 8614 967 8615 971
rect 8564 958 8578 967
rect 8467 954 8472 956
rect 8544 955 8563 956
rect 8564 955 8576 958
rect 8472 951 8479 954
rect 8544 951 8576 955
rect 8578 951 8579 957
rect 8479 950 8481 951
rect 8369 944 8381 945
rect 8339 943 8346 944
rect 8388 943 8397 945
rect 8339 942 8344 943
rect 8339 941 8341 942
rect 8339 940 8385 941
rect 8386 940 8397 943
rect 8335 939 8340 940
rect 8347 939 8381 940
rect 8335 938 8381 939
rect 8335 937 8347 938
rect 8284 926 8291 934
rect 8334 931 8347 937
rect 8378 936 8381 938
rect 8385 937 8397 940
rect 8429 943 8499 950
rect 8544 949 8564 951
rect 8567 949 8581 950
rect 8557 948 8581 949
rect 8557 946 8564 948
rect 8567 945 8584 948
rect 8609 946 8614 967
rect 8626 951 8628 968
rect 8750 966 8756 972
rect 8759 967 8762 972
rect 8628 949 8633 950
rect 8429 942 8502 943
rect 8429 939 8499 942
rect 8502 939 8511 942
rect 8567 939 8581 945
rect 8584 943 8594 945
rect 8623 943 8633 949
rect 8762 948 8769 967
rect 8796 966 8808 972
rect 8901 968 8912 978
rect 8936 980 8955 986
rect 8936 973 8973 980
rect 9097 976 9113 984
rect 9175 982 9178 986
rect 9174 976 9175 981
rect 8918 968 8921 972
rect 8802 945 8808 966
rect 8912 953 8924 968
rect 8940 965 8973 973
rect 9057 968 9060 976
rect 9098 975 9113 976
rect 9173 970 9174 975
rect 9216 969 9219 986
rect 9228 972 9329 977
rect 9329 969 9340 972
rect 9371 969 9472 988
rect 9502 980 9524 994
rect 8918 951 8921 953
rect 8924 951 8926 953
rect 8499 937 8531 939
rect 8379 931 8381 936
rect 8392 931 8398 937
rect 8499 934 8563 937
rect 8567 934 8583 939
rect 8594 934 8658 943
rect 8926 942 8946 951
rect 8955 948 8973 965
rect 9053 957 9057 968
rect 9048 955 9053 957
rect 9010 950 9011 953
rect 8771 939 8778 942
rect 8795 939 8835 942
rect 8759 936 8795 939
rect 8742 934 8759 936
rect 8335 930 8347 931
rect 7912 921 7921 923
rect 7900 920 7912 921
rect 7939 920 7944 924
rect 7853 915 7939 920
rect 7841 914 7853 915
rect 7881 914 7900 915
rect 7998 914 8006 926
rect 8010 924 8044 926
rect 7706 913 7836 914
rect 7814 909 7828 913
rect 7870 911 7881 914
rect 7863 907 7869 911
rect 7753 900 7759 906
rect 7759 894 7765 900
rect 7787 892 7800 900
rect 7830 892 7841 907
rect 7855 900 7860 904
rect 7992 901 8001 913
rect 8010 901 8012 924
rect 7625 888 7643 890
rect 7787 889 7796 892
rect 7800 891 7802 892
rect 7842 889 7844 891
rect 7852 889 7861 898
rect 8001 892 8012 901
rect 8042 892 8044 924
rect 8048 914 8056 926
rect 8154 924 8164 926
rect 8221 924 8249 926
rect 8250 924 8261 926
rect 8154 923 8162 924
rect 8159 921 8162 923
rect 8214 921 8215 924
rect 8247 921 8261 924
rect 8080 907 8094 921
rect 8149 910 8159 921
rect 8213 917 8214 921
rect 8149 907 8162 910
rect 8212 907 8213 916
rect 8247 915 8249 921
rect 8250 915 8261 921
rect 8284 924 8292 926
rect 8284 915 8291 924
rect 8292 921 8296 924
rect 8295 918 8301 921
rect 8296 916 8301 918
rect 8247 911 8250 915
rect 8252 914 8261 915
rect 8252 912 8253 914
rect 8094 906 8149 907
rect 8156 904 8162 907
rect 8211 904 8212 906
rect 8214 904 8220 910
rect 8247 906 8249 911
rect 8253 907 8255 912
rect 8255 906 8256 907
rect 8246 904 8249 906
rect 8256 904 8257 906
rect 8162 898 8168 904
rect 8204 902 8207 904
rect 8208 902 8214 904
rect 8203 898 8214 902
rect 8245 901 8246 904
rect 8203 892 8210 898
rect 8244 897 8245 900
rect 8242 894 8244 895
rect 8247 894 8249 904
rect 8215 892 8249 894
rect 8253 901 8261 904
rect 8253 892 8267 901
rect 8242 891 8244 892
rect 8267 890 8270 892
rect 7368 879 7372 885
rect 7494 879 7547 886
rect 7557 883 7563 886
rect 7564 883 7576 886
rect 7631 884 7637 888
rect 7365 875 7368 879
rect 7464 875 7494 879
rect 7505 877 7511 879
rect 7310 871 7311 875
rect 7362 870 7365 874
rect 7426 870 7464 875
rect 7424 869 7426 870
rect 7361 868 7362 869
rect 7422 868 7424 869
rect 7513 868 7515 879
rect 7548 868 7549 879
rect 7551 877 7557 883
rect 7625 882 7637 884
rect 7689 882 7695 888
rect 7625 876 7643 882
rect 7683 876 7689 882
rect 7796 880 7805 889
rect 7842 888 7852 889
rect 8240 888 8242 889
rect 7843 887 7852 888
rect 7843 880 7863 887
rect 8045 885 8046 888
rect 8006 882 8007 884
rect 8215 880 8227 888
rect 8237 882 8249 888
rect 8270 884 8272 890
rect 8274 885 8284 915
rect 8301 912 8314 916
rect 8314 907 8326 912
rect 8329 906 8331 907
rect 8340 906 8347 930
rect 8392 928 8393 931
rect 8515 919 8563 934
rect 8583 932 8658 934
rect 8675 933 8726 934
rect 8728 933 8739 934
rect 8675 932 8736 933
rect 8583 930 8675 932
rect 8331 904 8336 906
rect 8340 904 8392 906
rect 8336 901 8392 904
rect 8340 899 8392 901
rect 8323 889 8332 898
rect 8340 896 8409 899
rect 8340 891 8397 896
rect 8409 892 8434 896
rect 8531 894 8539 919
rect 8563 916 8570 919
rect 8583 918 8599 930
rect 8601 918 8617 930
rect 8722 929 8737 932
rect 8718 927 8722 929
rect 8702 922 8718 927
rect 8728 926 8737 929
rect 8771 926 8778 936
rect 8731 920 8736 922
rect 8549 900 8553 916
rect 8570 914 8601 916
rect 8602 914 8604 918
rect 8570 909 8602 914
rect 8593 907 8610 909
rect 8593 902 8602 907
rect 8610 906 8614 907
rect 8553 896 8554 899
rect 8573 898 8593 902
rect 8334 889 8398 891
rect 8434 890 8446 892
rect 8530 890 8531 893
rect 8332 885 8398 889
rect 8236 880 8249 882
rect 7806 875 7809 880
rect 7850 879 7863 880
rect 7348 864 7361 868
rect 7416 864 7422 868
rect 7342 862 7348 864
rect 7413 862 7416 864
rect 7339 858 7342 862
rect 7406 857 7413 862
rect 7338 856 7339 857
rect 7405 856 7406 857
rect 7337 849 7338 856
rect 7402 849 7405 856
rect 7336 841 7337 849
rect 7404 838 7413 842
rect 7451 838 7460 842
rect 7463 838 7479 854
rect 7481 838 7497 854
rect 7515 838 7519 867
rect 7546 847 7548 867
rect 7809 860 7816 875
rect 7848 873 7863 875
rect 7559 849 7573 854
rect 7655 842 7659 856
rect 5870 804 5880 805
rect 7332 804 7336 838
rect 7401 833 7413 838
rect 7447 833 7463 838
rect 7497 837 7513 838
rect 7504 834 7513 837
rect 7395 832 7408 833
rect 7447 832 7469 833
rect 7393 831 7402 832
rect 7393 811 7395 831
rect 7396 826 7402 831
rect 7392 810 7395 811
rect 7393 804 7395 810
rect 7401 820 7402 826
rect 7434 824 7469 832
rect 7434 823 7463 824
rect 7434 822 7482 823
rect 7508 822 7513 834
rect 7434 820 7454 822
rect 7463 820 7482 822
rect 7401 804 7417 820
rect 7447 804 7463 820
rect 7507 812 7508 817
rect 5778 803 5779 804
rect 5777 801 5778 802
rect 5725 799 5768 801
rect 5560 796 5725 799
rect 5560 795 5666 796
rect 5749 795 5768 799
rect 5542 794 5576 795
rect 5524 792 5558 794
rect 5503 789 5532 792
rect 5418 785 5429 788
rect 5478 787 5503 789
rect 5465 786 5478 787
rect 5461 785 5465 786
rect 5320 784 5323 785
rect 5341 784 5429 785
rect 5341 783 5418 784
rect 5434 783 5461 785
rect 5489 784 5492 787
rect 5163 779 5164 780
rect 5201 769 5209 783
rect 5243 778 5244 783
rect 5319 781 5320 783
rect 5342 782 5344 783
rect 5318 778 5319 781
rect 5344 780 5347 782
rect 5352 781 5353 783
rect 5410 782 5434 783
rect 5399 779 5410 782
rect 5347 778 5350 779
rect 4899 756 4917 757
rect 4945 756 4951 758
rect 4893 750 4957 756
rect 4982 753 5012 766
rect 5042 763 5080 769
rect 5198 763 5201 769
rect 5042 759 5074 763
rect 5041 756 5042 758
rect 4982 750 5018 753
rect 5039 752 5041 756
rect 5043 755 5074 759
rect 5071 754 5073 755
rect 5074 754 5077 755
rect 5193 754 5198 763
rect 5070 752 5071 754
rect 5077 751 5082 754
rect 5192 752 5193 754
rect 4793 744 4799 750
rect 4899 745 4951 750
rect 4703 742 4747 744
rect 4552 741 4586 742
rect 4703 741 4709 742
rect 4515 740 4552 741
rect 4492 739 4515 740
rect 4489 737 4492 739
rect 4741 738 4747 742
rect 4799 738 4805 744
rect 4464 723 4489 737
rect 4580 730 4586 736
rect 4638 731 4644 736
rect 4893 733 4905 745
rect 4939 735 4944 745
rect 4669 731 4705 733
rect 4586 724 4592 730
rect 4610 729 4669 731
rect 4705 729 4711 731
rect 4608 726 4610 729
rect 4459 720 4464 723
rect 4357 717 4439 719
rect 4360 716 4439 717
rect 4456 716 4464 720
rect 4406 713 4414 716
rect 4418 715 4420 716
rect 4439 715 4468 716
rect 4418 713 4452 715
rect 4449 709 4452 713
rect 4456 713 4464 715
rect 4468 714 4496 715
rect 4456 711 4459 713
rect 4453 709 4456 711
rect 4496 710 4510 714
rect 4602 713 4608 726
rect 4632 724 4638 729
rect 4711 726 4722 729
rect 4899 726 4905 733
rect 4701 722 4703 723
rect 4722 722 4733 726
rect 4898 723 4905 726
rect 4733 721 4735 722
rect 4735 720 4739 721
rect 4083 707 4084 708
rect 4305 707 4306 708
rect 4418 701 4430 709
rect 4440 701 4452 709
rect 4510 705 4516 710
rect 4600 708 4602 713
rect 4599 707 4600 708
rect 4516 703 4527 705
rect 4144 697 4278 700
rect 4444 698 4448 701
rect 4527 699 4540 703
rect 4540 698 4545 699
rect 4020 695 4144 697
rect 4278 695 4284 697
rect 3923 692 3929 694
rect 3998 692 4020 695
rect 4284 692 4290 695
rect 3705 688 3706 690
rect 3919 688 3921 691
rect 3922 688 3923 690
rect 3975 689 3998 692
rect 4290 689 4296 692
rect 4428 690 4444 698
rect 4545 694 4561 698
rect 4561 692 4577 694
rect 4577 691 4586 692
rect 4592 691 4599 706
rect 4693 693 4701 698
rect 4705 693 4707 720
rect 4893 711 4905 723
rect 4944 711 4946 726
rect 4982 723 5012 750
rect 5038 749 5039 751
rect 5082 750 5084 751
rect 5022 746 5024 747
rect 5036 745 5038 749
rect 5025 737 5039 745
rect 5067 744 5069 749
rect 5087 747 5090 749
rect 5090 746 5092 747
rect 5092 743 5096 746
rect 5116 743 5128 749
rect 5187 744 5190 749
rect 5222 744 5243 778
rect 5309 756 5318 778
rect 5347 776 5352 778
rect 5353 776 5399 779
rect 5492 778 5493 781
rect 5347 775 5399 776
rect 5347 756 5352 775
rect 5493 772 5497 778
rect 5493 756 5500 772
rect 5524 756 5532 789
rect 5542 788 5558 792
rect 5560 788 5576 794
rect 5638 788 5654 795
rect 5752 788 5768 795
rect 5755 787 5756 788
rect 5756 783 5757 785
rect 5758 772 5761 779
rect 5781 778 5793 804
rect 5830 799 5831 802
rect 5830 796 5832 799
rect 5868 796 5870 800
rect 7336 799 7349 804
rect 7366 799 7401 804
rect 7349 797 7366 799
rect 5830 791 5838 796
rect 5865 791 5868 796
rect 5830 788 5846 791
rect 5848 788 5864 791
rect 7385 788 7402 799
rect 7463 797 7466 803
rect 7463 795 7467 797
rect 7463 788 7473 795
rect 7393 786 7402 788
rect 7467 786 7473 788
rect 7518 786 7519 828
rect 7543 822 7556 838
rect 7689 833 7693 838
rect 7711 837 7723 845
rect 7777 838 7793 854
rect 7816 842 7825 860
rect 7817 841 7825 842
rect 7829 845 7830 862
rect 7829 843 7833 845
rect 7861 844 7863 873
rect 7864 869 7875 875
rect 7867 863 7875 869
rect 7871 859 7874 863
rect 8007 860 8011 879
rect 8044 866 8045 880
rect 8126 867 8132 873
rect 8172 867 8178 873
rect 8236 870 8240 880
rect 8269 870 8274 884
rect 8332 880 8346 885
rect 8340 871 8346 880
rect 8382 880 8392 885
rect 8382 870 8383 880
rect 8386 879 8392 880
rect 8446 879 8513 890
rect 8529 885 8530 889
rect 8528 881 8529 885
rect 8514 875 8518 879
rect 8518 872 8521 875
rect 8525 871 8528 881
rect 8554 879 8558 896
rect 8568 891 8573 898
rect 8614 892 8671 906
rect 8671 891 8674 892
rect 8565 881 8567 889
rect 8674 888 8688 891
rect 8734 890 8736 920
rect 8740 910 8748 922
rect 8778 914 8783 926
rect 8783 902 8788 914
rect 8808 910 8815 939
rect 8835 936 8841 939
rect 8841 934 8845 936
rect 8922 935 8923 942
rect 8946 939 8952 942
rect 8952 936 8958 939
rect 8845 933 8846 934
rect 8846 927 8849 933
rect 8849 922 8852 927
rect 8852 919 8854 922
rect 8854 916 8855 919
rect 8705 888 8736 890
rect 8740 888 8748 900
rect 8788 899 8789 902
rect 8815 900 8817 910
rect 8855 902 8862 916
rect 8923 910 8927 935
rect 8958 934 8962 936
rect 8973 935 8974 942
rect 8960 933 8966 934
rect 8960 932 8968 933
rect 8974 932 8975 935
rect 9010 934 9025 950
rect 9048 948 9060 955
rect 9047 947 9060 948
rect 9070 947 9082 955
rect 9113 952 9129 968
rect 9044 945 9053 947
rect 9043 943 9044 945
rect 9047 943 9053 945
rect 9086 943 9087 945
rect 9093 943 9099 948
rect 9036 942 9043 943
rect 9047 942 9082 943
rect 9086 942 9099 943
rect 9036 937 9047 942
rect 9048 941 9082 942
rect 9034 934 9040 937
rect 9041 936 9047 937
rect 9081 936 9082 941
rect 9099 936 9105 942
rect 9113 934 9129 950
rect 9166 939 9173 968
rect 9219 956 9220 968
rect 9224 965 9225 969
rect 9340 968 9359 969
rect 9367 968 9371 969
rect 9331 964 9367 968
rect 9417 965 9421 969
rect 9165 934 9166 938
rect 9030 932 9034 934
rect 8968 931 9009 932
rect 8974 918 8991 931
rect 8993 926 9009 931
rect 9027 930 9030 932
rect 9020 926 9027 930
rect 9112 927 9113 931
rect 9164 927 9165 932
rect 8993 918 9020 926
rect 9111 920 9113 927
rect 9163 922 9164 927
rect 9174 922 9182 934
rect 9186 922 9188 956
rect 9224 951 9225 964
rect 9331 960 9379 964
rect 9322 954 9331 960
rect 9219 945 9220 951
rect 9225 936 9226 945
rect 9314 939 9322 954
rect 9360 949 9379 960
rect 9379 948 9381 949
rect 9421 948 9426 965
rect 9524 961 9527 980
rect 9527 954 9528 960
rect 9381 945 9385 948
rect 9426 945 9427 948
rect 9311 936 9314 939
rect 9226 928 9232 934
rect 9227 922 9232 928
rect 9306 928 9318 936
rect 9328 928 9340 936
rect 9385 934 9400 945
rect 9427 934 9431 945
rect 9528 941 9531 954
rect 9530 939 9531 941
rect 9528 934 9530 939
rect 9400 932 9401 934
rect 9401 928 9402 930
rect 9431 929 9433 934
rect 9306 924 9311 928
rect 9344 926 9345 928
rect 9346 924 9349 925
rect 9110 919 9113 920
rect 8974 905 8975 918
rect 9002 916 9020 918
rect 9109 918 9113 919
rect 9109 916 9110 918
rect 9162 916 9163 919
rect 9182 916 9183 921
rect 8996 912 9002 916
rect 9105 909 9109 916
rect 9161 909 9162 916
rect 9183 912 9185 916
rect 9213 913 9220 922
rect 9227 916 9228 922
rect 9206 911 9213 913
rect 9224 911 9228 916
rect 9294 912 9302 924
rect 9306 922 9340 924
rect 9306 921 9309 922
rect 9186 910 9224 911
rect 8975 902 8976 904
rect 8862 899 8864 902
rect 8817 894 8818 899
rect 8864 896 8865 899
rect 8688 885 8699 888
rect 8702 885 8741 888
rect 8699 884 8741 885
rect 8558 872 8560 879
rect 8560 870 8561 872
rect 8562 871 8565 881
rect 8702 879 8741 884
rect 8790 881 8792 889
rect 8724 876 8736 879
rect 8741 874 8763 879
rect 8792 874 8793 881
rect 8777 872 8782 874
rect 8211 868 8212 869
rect 8235 867 8236 870
rect 8120 861 8126 867
rect 8178 861 8184 867
rect 8233 860 8235 867
rect 7874 854 7878 858
rect 7874 853 7889 854
rect 7860 843 7863 844
rect 7829 841 7863 843
rect 7867 841 7875 853
rect 7878 850 7889 853
rect 8011 852 8012 858
rect 8045 854 8046 858
rect 7880 845 7889 850
rect 7883 840 7889 845
rect 7646 831 7723 833
rect 7546 820 7551 822
rect 7543 804 7556 820
rect 7546 787 7551 804
rect 7559 788 7575 799
rect 7395 780 7402 786
rect 7460 785 7473 786
rect 7460 783 7507 785
rect 7435 780 7482 783
rect 5304 745 5309 756
rect 5344 744 5347 756
rect 5497 750 5500 756
rect 5497 744 5504 750
rect 5532 744 5534 756
rect 5562 751 5574 759
rect 5584 751 5596 759
rect 5761 755 5766 772
rect 5793 770 5797 778
rect 7395 777 7408 780
rect 7448 777 7454 780
rect 7460 779 7482 780
rect 7460 777 7469 779
rect 7646 777 7704 831
rect 7721 799 7723 831
rect 7727 821 7735 833
rect 7793 822 7809 838
rect 7863 837 7867 840
rect 7887 838 7889 840
rect 7911 838 7917 844
rect 7957 839 7963 844
rect 7953 838 7965 839
rect 8012 838 8015 850
rect 8047 841 8063 854
rect 8118 852 8126 858
rect 8116 850 8126 852
rect 8230 851 8233 860
rect 8179 848 8189 850
rect 8189 846 8195 848
rect 8228 847 8230 851
rect 8106 845 8114 846
rect 8116 845 8120 846
rect 8046 840 8063 841
rect 8046 838 8050 840
rect 7829 829 7841 837
rect 7851 829 7863 837
rect 7889 832 7969 838
rect 8015 832 8016 837
rect 7829 828 7830 829
rect 7830 818 7832 828
rect 7889 822 7905 832
rect 7911 831 7965 832
rect 7911 827 7963 831
rect 7832 814 7834 818
rect 7834 809 7835 812
rect 7835 805 7836 809
rect 7836 799 7837 803
rect 7837 792 7839 799
rect 7911 793 7931 827
rect 7957 825 7965 827
rect 7963 794 7965 825
rect 7969 815 7977 827
rect 7957 793 7965 794
rect 7969 793 7977 805
rect 7993 804 8001 820
rect 8016 814 8019 829
rect 8031 822 8050 838
rect 8084 833 8093 842
rect 8106 841 8116 845
rect 8118 844 8120 845
rect 8195 844 8202 846
rect 8118 841 8126 844
rect 8202 843 8206 844
rect 8206 842 8211 843
rect 8227 842 8228 844
rect 8223 841 8234 842
rect 8259 841 8269 869
rect 8274 866 8275 869
rect 8275 854 8278 865
rect 8346 860 8351 870
rect 8522 869 8525 870
rect 8521 865 8525 869
rect 8522 860 8525 865
rect 8552 866 8562 870
rect 8782 866 8799 872
rect 8818 871 8822 890
rect 8865 888 8869 896
rect 8973 890 8976 896
rect 8982 891 8993 908
rect 9048 903 9060 909
rect 9160 908 9161 909
rect 9089 903 9105 908
rect 9159 903 9160 908
rect 9206 903 9213 910
rect 9060 902 9089 903
rect 9158 896 9159 899
rect 9041 890 9047 896
rect 9099 890 9105 896
rect 8869 874 8877 888
rect 8971 885 8973 889
rect 8979 886 8982 890
rect 8351 854 8352 860
rect 8521 854 8524 860
rect 8275 852 8281 854
rect 8278 846 8281 852
rect 8343 849 8359 854
rect 8342 848 8356 849
rect 8361 848 8377 854
rect 8279 841 8281 846
rect 8339 845 8342 848
rect 8356 845 8377 848
rect 8334 841 8339 845
rect 8367 842 8379 845
rect 8106 838 8120 841
rect 8226 839 8227 841
rect 8234 840 8269 841
rect 8280 840 8281 841
rect 8332 840 8334 841
rect 8259 839 8307 840
rect 8330 838 8332 840
rect 8346 839 8358 842
rect 8439 841 8455 854
rect 8457 841 8473 854
rect 8519 847 8521 853
rect 8522 852 8524 854
rect 8552 852 8570 866
rect 8793 863 8808 866
rect 8379 840 8380 841
rect 8432 840 8433 841
rect 8351 838 8358 839
rect 8100 834 8114 838
rect 8100 833 8111 834
rect 8075 824 8084 833
rect 8046 820 8050 822
rect 8031 814 8050 820
rect 8019 809 8020 812
rect 8020 799 8022 808
rect 8031 804 8047 814
rect 8106 812 8114 824
rect 8118 814 8120 838
rect 8223 832 8226 838
rect 8178 815 8184 821
rect 8212 818 8230 832
rect 8218 815 8219 818
rect 8172 814 8178 815
rect 8217 814 8218 815
rect 8118 812 8152 814
rect 8161 812 8220 814
rect 8230 813 8236 818
rect 8231 812 8237 813
rect 8050 808 8051 812
rect 8142 809 8152 812
rect 8156 810 8161 812
rect 8133 808 8142 809
rect 8145 808 8151 809
rect 8153 808 8156 810
rect 8172 809 8178 812
rect 8051 804 8052 808
rect 8118 805 8130 808
rect 8133 805 8152 808
rect 8118 804 8131 805
rect 8047 794 8055 804
rect 8078 800 8130 804
rect 8140 800 8152 805
rect 8208 800 8217 811
rect 8220 810 8228 812
rect 8231 810 8242 812
rect 8250 811 8259 838
rect 8281 822 8297 838
rect 8321 832 8329 838
rect 8228 809 8242 810
rect 8244 809 8250 810
rect 8228 808 8250 809
rect 8281 808 8297 820
rect 8350 811 8352 838
rect 8353 837 8358 838
rect 8355 836 8358 837
rect 8380 838 8381 840
rect 8431 838 8432 840
rect 8356 834 8360 836
rect 8361 832 8362 834
rect 8380 832 8393 838
rect 8354 828 8358 830
rect 8231 804 8297 808
rect 8240 800 8281 804
rect 8321 801 8322 804
rect 8047 793 8057 794
rect 7911 792 7963 793
rect 8047 792 8059 793
rect 7839 789 7845 792
rect 7845 784 7852 789
rect 7905 788 7985 792
rect 8023 790 8024 792
rect 8047 789 8068 792
rect 8047 788 8062 789
rect 7905 786 7969 788
rect 8057 786 8062 788
rect 8068 787 8073 789
rect 8073 786 8077 787
rect 8078 786 8129 800
rect 8141 793 8145 800
rect 8203 793 8208 799
rect 8140 790 8141 793
rect 8201 790 8203 793
rect 7852 783 7853 784
rect 7888 783 7889 785
rect 7854 779 7860 783
rect 7885 779 7888 783
rect 7911 780 7917 786
rect 7953 781 7965 786
rect 8073 785 8084 786
rect 8075 783 8084 785
rect 8075 782 8087 783
rect 7957 780 7963 781
rect 8023 779 8024 781
rect 7860 777 7865 779
rect 7884 777 7885 779
rect 5544 747 5550 750
rect 5598 749 5600 750
rect 5553 747 5557 749
rect 5544 746 5553 747
rect 5543 744 5551 746
rect 5562 745 5598 747
rect 5600 745 5608 747
rect 5065 738 5067 743
rect 5096 741 5128 743
rect 5124 740 5129 741
rect 5131 737 5134 739
rect 5184 738 5187 744
rect 5219 739 5222 744
rect 5302 740 5304 744
rect 5319 740 5331 742
rect 5032 734 5033 737
rect 5039 734 5043 737
rect 5031 732 5032 734
rect 5043 732 5047 734
rect 5063 732 5065 737
rect 5093 736 5094 737
rect 5123 734 5133 737
rect 5134 734 5140 737
rect 5146 734 5152 737
rect 5128 732 5133 734
rect 5028 725 5031 731
rect 5047 729 5051 732
rect 5061 729 5063 731
rect 5027 722 5028 724
rect 5023 711 5027 721
rect 5051 712 5079 729
rect 5092 726 5093 731
rect 5133 727 5137 732
rect 5139 731 5152 734
rect 5177 732 5181 734
rect 5175 731 5177 732
rect 5192 731 5198 737
rect 5282 734 5288 740
rect 5300 734 5301 736
rect 5319 734 5334 740
rect 5343 738 5344 742
rect 5492 738 5498 744
rect 5550 738 5556 744
rect 5562 743 5564 745
rect 5342 734 5343 737
rect 5215 732 5216 734
rect 5276 732 5340 734
rect 5137 726 5139 727
rect 5140 726 5146 731
rect 4894 710 4898 711
rect 4899 710 4951 711
rect 4893 706 4957 710
rect 4888 704 4957 706
rect 5020 704 5023 711
rect 4747 698 4753 699
rect 4761 698 4799 699
rect 4741 695 4753 698
rect 4757 695 4805 698
rect 4741 693 4747 695
rect 4757 693 4795 695
rect 4799 693 4805 695
rect 4693 692 4805 693
rect 4693 691 4787 692
rect 4296 688 4299 689
rect 4303 688 4305 690
rect 3706 669 3716 688
rect 3917 682 3923 688
rect 3975 682 3981 688
rect 4299 686 4305 688
rect 3922 680 3935 682
rect 3922 676 3929 680
rect 3969 676 3975 682
rect 4303 677 4305 686
rect 4405 681 4428 690
rect 4586 689 4608 691
rect 4693 689 4783 691
rect 4405 679 4475 681
rect 3716 658 3726 669
rect 3718 656 3732 658
rect 3768 656 3784 672
rect 3922 668 3923 676
rect 4299 671 4305 677
rect 4357 678 4428 679
rect 4357 676 4421 678
rect 4475 676 4484 679
rect 4357 671 4363 676
rect 3922 656 3934 668
rect 4302 665 4311 671
rect 4351 665 4357 671
rect 4302 662 4305 665
rect 4386 662 4405 676
rect 4484 675 4488 676
rect 4488 672 4490 675
rect 4492 667 4493 669
rect 4302 658 4304 662
rect 4382 659 4386 662
rect 4493 660 4508 667
rect 4592 662 4598 689
rect 4608 686 4643 689
rect 4693 686 4777 689
rect 4793 686 4799 692
rect 4888 690 4893 704
rect 4899 699 4917 704
rect 4899 698 4905 699
rect 4945 698 4951 704
rect 5018 699 5020 704
rect 4946 696 4947 698
rect 5016 695 5018 698
rect 5052 695 5060 712
rect 5080 709 5083 711
rect 5088 709 5092 726
rect 5139 717 5149 726
rect 5198 725 5204 731
rect 5211 725 5215 732
rect 5276 730 5334 732
rect 5335 730 5340 732
rect 5341 730 5342 732
rect 5276 728 5332 730
rect 5209 722 5210 724
rect 5149 709 5151 717
rect 5203 711 5209 721
rect 5083 708 5085 709
rect 5082 707 5086 708
rect 5082 703 5088 707
rect 5094 705 5095 707
rect 5094 703 5111 705
rect 5013 694 5016 695
rect 5009 692 5013 694
rect 5007 691 5009 692
rect 4643 684 4662 686
rect 4701 684 4765 686
rect 4662 683 4670 684
rect 4670 681 4691 683
rect 4701 681 4760 684
rect 4691 679 4760 681
rect 4884 679 4888 689
rect 4947 686 4949 690
rect 5003 689 5007 691
rect 4999 688 5003 689
rect 5049 688 5052 695
rect 5085 690 5088 703
rect 5091 699 5093 700
rect 5094 696 5118 699
rect 5094 691 5106 696
rect 5118 693 5132 696
rect 5151 693 5153 706
rect 5198 702 5203 711
rect 5282 696 5297 728
rect 5329 726 5332 728
rect 5335 726 5343 730
rect 5329 724 5331 726
rect 5330 700 5331 724
rect 5332 718 5343 726
rect 5332 714 5336 718
rect 5332 710 5335 714
rect 5338 712 5340 718
rect 5594 715 5596 745
rect 5598 742 5608 745
rect 5768 743 5770 749
rect 5778 743 5784 749
rect 5797 746 5820 770
rect 7282 755 7283 775
rect 7311 772 7312 775
rect 7402 774 7441 777
rect 7448 774 7460 777
rect 7312 759 7320 772
rect 7404 768 7441 774
rect 7451 768 7460 774
rect 7517 768 7518 777
rect 7312 755 7323 759
rect 7283 749 7284 755
rect 7320 753 7323 755
rect 7321 750 7326 753
rect 5824 743 5830 749
rect 7295 747 7324 748
rect 7327 747 7328 749
rect 5772 742 5778 743
rect 5600 738 5608 742
rect 5600 735 5618 738
rect 5608 731 5618 735
rect 5770 731 5778 742
rect 5783 738 5784 742
rect 5816 739 5822 742
rect 5781 731 5783 738
rect 5817 737 5822 739
rect 5830 737 5836 743
rect 5568 714 5596 715
rect 5563 713 5596 714
rect 5600 713 5608 725
rect 5618 721 5624 731
rect 5770 721 5781 731
rect 5762 720 5781 721
rect 5762 712 5771 720
rect 5337 710 5338 711
rect 5335 707 5339 710
rect 5597 709 5600 711
rect 5571 708 5574 709
rect 5334 702 5339 707
rect 5559 706 5569 708
rect 5550 704 5559 706
rect 5329 696 5331 699
rect 5132 692 5198 693
rect 5138 691 5198 692
rect 4972 686 4999 688
rect 5048 686 5049 688
rect 4947 684 4979 686
rect 4937 683 4979 684
rect 4910 681 4979 683
rect 4892 679 4979 681
rect 5045 679 5048 684
rect 4701 678 4760 679
rect 4704 677 4739 678
rect 4865 677 4979 679
rect 4704 676 4736 677
rect 4738 676 4739 677
rect 4705 674 4717 676
rect 4719 675 4738 676
rect 4843 675 4865 677
rect 4871 676 4979 677
rect 4884 675 4888 676
rect 4719 671 4746 675
rect 4795 671 4843 675
rect 4719 670 4757 671
rect 4784 670 4827 671
rect 4719 664 4827 670
rect 4721 662 4731 664
rect 4884 662 4885 675
rect 4949 672 4951 675
rect 5042 673 5045 679
rect 4598 660 4599 662
rect 4380 658 4382 659
rect 4082 656 4084 657
rect 4302 656 4303 658
rect 4378 656 4380 658
rect 3734 640 3750 656
rect 3752 640 3768 656
rect 3935 653 3937 656
rect 4075 653 4081 656
rect 4304 653 4307 656
rect 4374 653 4378 656
rect 3937 651 3939 653
rect 4074 652 4075 653
rect 4372 652 4374 653
rect 4508 652 4620 660
rect 4712 658 4721 662
rect 4949 659 4952 672
rect 5081 666 5085 689
rect 5144 685 5198 691
rect 5282 688 5334 696
rect 5335 692 5339 702
rect 5492 693 5498 698
rect 5550 693 5556 698
rect 5492 692 5556 693
rect 5339 688 5341 690
rect 5140 679 5204 685
rect 5276 682 5341 688
rect 5498 686 5504 692
rect 5544 686 5550 692
rect 5562 690 5563 706
rect 5584 701 5596 709
rect 5775 707 5781 720
rect 5818 717 5822 737
rect 5774 706 5775 707
rect 5770 697 5774 706
rect 5822 697 5824 717
rect 6585 703 6607 722
rect 7277 713 7284 725
rect 7289 716 7290 747
rect 7318 745 7323 747
rect 7322 716 7323 745
rect 7324 738 7335 747
rect 7551 740 7555 777
rect 7860 776 7884 777
rect 8021 775 8023 779
rect 8075 777 8084 782
rect 8090 779 8093 781
rect 8093 777 8112 779
rect 8140 777 8149 786
rect 8171 782 8177 788
rect 8198 786 8201 790
rect 8217 782 8223 788
rect 8235 786 8244 800
rect 8247 788 8263 800
rect 8265 796 8301 800
rect 8322 798 8324 801
rect 8349 800 8350 810
rect 8356 798 8358 828
rect 8362 818 8370 830
rect 8379 822 8393 832
rect 8423 836 8431 838
rect 8485 837 8489 841
rect 8517 839 8519 847
rect 8552 838 8562 852
rect 8570 848 8573 852
rect 8700 842 8706 844
rect 8700 838 8714 842
rect 8746 838 8752 844
rect 8753 838 8769 854
rect 8793 838 8799 863
rect 8808 853 8811 863
rect 8811 846 8813 852
rect 8813 838 8816 845
rect 8423 822 8430 836
rect 8447 826 8459 832
rect 8444 825 8503 826
rect 8507 825 8517 838
rect 8444 823 8452 825
rect 8503 823 8517 825
rect 8524 823 8527 838
rect 8379 820 8382 822
rect 8443 821 8444 823
rect 8322 796 8358 798
rect 8362 796 8370 808
rect 8379 804 8393 820
rect 8435 816 8443 820
rect 8447 818 8454 820
rect 8435 808 8441 816
rect 8447 814 8448 818
rect 8507 816 8532 823
rect 8541 816 8552 837
rect 8573 822 8585 838
rect 8694 832 8700 838
rect 8698 830 8700 832
rect 8702 830 8735 838
rect 8752 832 8758 838
rect 8769 832 8785 838
rect 8799 832 8800 838
rect 8752 830 8785 832
rect 8816 830 8819 838
rect 8822 830 8834 870
rect 8877 863 8882 874
rect 8924 871 8927 885
rect 8961 881 8971 885
rect 9047 884 9053 890
rect 9057 887 9058 890
rect 9067 886 9074 890
rect 9058 883 9061 885
rect 9064 884 9066 885
rect 9093 884 9099 890
rect 9156 888 9158 896
rect 9058 882 9063 883
rect 8959 874 8977 881
rect 8942 870 8959 874
rect 8961 870 8971 874
rect 8882 859 8884 863
rect 8908 838 8924 870
rect 8942 866 8961 870
rect 8940 863 8942 866
rect 8938 859 8940 863
rect 8954 859 8961 866
rect 8936 856 8938 859
rect 8934 854 8936 856
rect 8927 851 8936 854
rect 8927 845 8934 851
rect 8927 839 8931 845
rect 8927 838 8928 839
rect 8884 830 8885 838
rect 8908 830 8927 838
rect 8941 830 8954 859
rect 8971 846 8978 858
rect 8983 848 8984 880
rect 9050 876 9056 879
rect 9047 874 9050 876
rect 9038 869 9047 874
rect 9058 870 9061 882
rect 9095 870 9098 884
rect 9155 881 9156 888
rect 9154 874 9155 881
rect 9031 860 9032 863
rect 9061 860 9063 870
rect 9095 862 9109 870
rect 9151 863 9154 874
rect 9026 848 9031 860
rect 8983 847 8988 848
rect 8983 846 9017 847
rect 9024 846 9029 848
rect 8978 844 8979 846
rect 9023 844 9024 846
rect 9020 842 9022 843
rect 8983 834 8995 841
rect 9005 834 9017 841
rect 9063 830 9074 859
rect 9098 830 9109 862
rect 9150 856 9151 859
rect 9188 856 9206 903
rect 9294 890 9302 902
rect 9306 890 9308 921
rect 9339 920 9340 922
rect 9346 912 9352 924
rect 9402 913 9404 925
rect 9433 924 9449 928
rect 9519 925 9528 934
rect 9511 924 9519 925
rect 9433 913 9511 924
rect 9346 911 9349 912
rect 9349 903 9354 910
rect 9387 905 9449 913
rect 9381 903 9387 905
rect 9340 890 9381 903
rect 9349 888 9354 890
rect 9404 889 9406 905
rect 9302 886 9305 888
rect 9354 886 9355 888
rect 9406 885 9407 888
rect 9305 884 9307 885
rect 9306 883 9308 884
rect 9306 879 9309 883
rect 9355 880 9356 882
rect 9306 878 9310 879
rect 9309 876 9310 878
rect 9356 876 9357 880
rect 9407 876 9408 879
rect 9433 878 9449 905
rect 9310 869 9313 874
rect 9313 863 9315 869
rect 9248 861 9249 862
rect 9315 860 9316 863
rect 9127 851 9143 854
rect 9147 851 9150 856
rect 9186 851 9188 856
rect 9229 854 9241 855
rect 9127 845 9147 851
rect 9184 846 9186 851
rect 9223 847 9241 854
rect 9251 849 9263 855
rect 9251 847 9300 849
rect 9316 848 9320 860
rect 9223 845 9239 847
rect 9252 846 9300 847
rect 9245 845 9252 846
rect 9272 845 9300 846
rect 9127 843 9133 845
rect 9183 843 9184 845
rect 9223 843 9245 845
rect 9300 843 9314 845
rect 9320 844 9321 847
rect 9337 843 9353 854
rect 9125 839 9128 843
rect 9181 839 9183 843
rect 9217 842 9222 843
rect 9217 840 9221 842
rect 9223 841 9263 843
rect 9210 839 9220 840
rect 9223 839 9229 841
rect 9204 838 9209 839
rect 9223 838 9224 839
rect 9111 830 9125 838
rect 9178 836 9181 838
rect 9200 837 9204 838
rect 9191 836 9197 837
rect 9178 834 9191 836
rect 9168 833 9172 834
rect 9162 832 9168 833
rect 9149 830 9162 832
rect 9178 831 9181 834
rect 8690 827 8698 830
rect 8702 828 8705 830
rect 8689 821 8699 827
rect 8378 802 8379 804
rect 8380 800 8382 804
rect 8507 801 8517 816
rect 8519 812 8527 816
rect 8519 804 8528 812
rect 8532 807 8564 816
rect 8573 807 8585 820
rect 8665 807 8689 821
rect 8690 818 8698 821
rect 8528 801 8529 803
rect 8541 801 8552 807
rect 8564 804 8585 807
rect 8265 788 8281 796
rect 8301 795 8306 796
rect 8306 793 8317 795
rect 8324 794 8331 796
rect 8331 793 8337 794
rect 8348 793 8349 796
rect 8317 792 8322 793
rect 8337 792 8357 793
rect 8360 792 8362 795
rect 8377 794 8378 796
rect 8337 786 8358 792
rect 8374 789 8377 793
rect 8359 788 8377 789
rect 8359 786 8374 788
rect 8430 786 8431 788
rect 8435 786 8441 798
rect 8489 789 8490 801
rect 8504 790 8507 800
rect 8529 797 8557 801
rect 8564 797 8583 804
rect 8653 800 8665 807
rect 8651 799 8653 800
rect 8529 796 8583 797
rect 8644 796 8651 799
rect 8690 796 8698 808
rect 8702 796 8704 828
rect 8770 822 8999 830
rect 8770 820 8772 822
rect 8773 820 8999 822
rect 8770 814 8999 820
rect 9027 814 9149 830
rect 9172 818 9178 831
rect 9207 822 9223 838
rect 9170 815 9177 818
rect 8770 812 9027 814
rect 8772 804 8785 812
rect 8802 807 8804 812
rect 8772 803 8773 804
rect 8773 801 8774 802
rect 8770 796 8773 801
rect 8803 800 8804 807
rect 8815 804 8827 812
rect 8827 803 8828 804
rect 8832 803 8834 808
rect 8851 803 8930 812
rect 8828 802 8930 803
rect 8831 799 8847 802
rect 8448 787 8449 788
rect 8447 786 8453 787
rect 8229 782 8235 786
rect 8346 784 8358 786
rect 8020 772 8021 774
rect 8084 772 8112 777
rect 8013 759 8020 772
rect 8084 768 8093 772
rect 8131 768 8140 777
rect 8165 776 8171 782
rect 8223 776 8235 782
rect 8347 776 8348 781
rect 8223 766 8227 773
rect 8379 772 8380 786
rect 8431 783 8432 786
rect 8442 784 8444 785
rect 8488 784 8489 788
rect 8503 787 8504 790
rect 8529 789 8573 796
rect 8583 795 8585 796
rect 8585 792 8592 795
rect 8642 793 8644 796
rect 8741 795 8769 796
rect 8592 789 8596 792
rect 8529 788 8551 789
rect 8553 788 8569 789
rect 8596 788 8598 789
rect 8638 788 8642 793
rect 8753 792 8769 795
rect 8799 793 8803 799
rect 8510 787 8517 788
rect 8525 787 8539 788
rect 8598 787 8601 788
rect 8502 786 8510 787
rect 8497 785 8510 786
rect 8529 785 8539 787
rect 8694 786 8700 792
rect 8752 791 8769 792
rect 8796 791 8799 793
rect 8752 789 8808 791
rect 8829 789 8847 799
rect 8752 788 8769 789
rect 8796 788 8799 789
rect 8808 788 8847 789
rect 8849 788 8930 802
rect 8941 800 8954 812
rect 9017 804 9018 807
rect 8752 786 8758 788
rect 8795 786 8796 788
rect 8494 784 8503 785
rect 8432 780 8444 783
rect 8447 780 8448 781
rect 8456 780 8494 784
rect 8432 779 8491 780
rect 8447 774 8459 779
rect 8378 763 8380 772
rect 8497 763 8503 784
rect 8529 784 8543 785
rect 8003 756 8020 759
rect 8344 756 8347 763
rect 8003 755 8013 756
rect 8003 754 8010 755
rect 8343 754 8344 756
rect 8003 753 8007 754
rect 7992 749 8034 753
rect 7992 748 8019 749
rect 7990 747 7992 748
rect 8034 747 8037 749
rect 7976 745 7990 747
rect 7508 738 7514 740
rect 7551 739 7560 740
rect 7328 735 7346 738
rect 7335 725 7346 735
rect 7508 734 7520 738
rect 7554 734 7560 739
rect 7943 738 7976 745
rect 7937 737 7942 738
rect 7502 728 7508 734
rect 7560 729 7566 734
rect 7914 733 7937 737
rect 7991 735 7999 747
rect 8003 746 8008 747
rect 7908 731 7914 733
rect 7902 729 7904 731
rect 7524 728 7655 729
rect 7508 726 7524 728
rect 7560 727 7863 728
rect 7890 727 7896 729
rect 7901 728 7902 729
rect 7655 726 7656 727
rect 7863 726 7896 727
rect 7899 726 7901 728
rect 7289 714 7293 716
rect 7320 714 7323 716
rect 7289 713 7323 714
rect 7328 713 7346 725
rect 7496 714 7504 726
rect 7508 724 7514 726
rect 7284 711 7285 713
rect 7285 708 7290 711
rect 7323 708 7328 711
rect 7289 707 7301 708
rect 6556 697 6579 698
rect 6584 697 6607 703
rect 7288 701 7301 707
rect 7311 701 7323 708
rect 7335 707 7346 713
rect 5770 693 5778 697
rect 5830 693 5836 697
rect 7288 694 7290 701
rect 5770 691 5836 693
rect 5770 690 5774 691
rect 5563 686 5565 690
rect 5144 673 5152 679
rect 5192 673 5198 679
rect 5282 676 5288 682
rect 5328 676 5334 682
rect 5144 666 5151 673
rect 5284 672 5287 676
rect 4708 656 4712 658
rect 4885 656 4886 658
rect 4950 657 4952 659
rect 4948 656 4952 657
rect 4703 653 4708 656
rect 4886 653 4889 656
rect 4947 653 4948 656
rect 4982 654 5012 663
rect 5016 654 5029 660
rect 5081 659 5083 666
rect 5144 665 5152 666
rect 4698 652 4699 653
rect 4946 652 4947 653
rect 4979 652 5016 654
rect 5083 653 5085 659
rect 5141 656 5152 665
rect 5278 660 5287 672
rect 5340 672 5341 682
rect 5278 656 5284 660
rect 5340 656 5344 672
rect 5556 660 5565 686
rect 5764 674 5770 690
rect 5778 685 5784 691
rect 5824 685 5830 691
rect 7346 690 7353 707
rect 7496 692 7504 704
rect 7508 694 7510 724
rect 7657 719 7661 726
rect 7863 723 7898 726
rect 7936 723 7942 729
rect 7661 708 7668 719
rect 7884 717 7890 723
rect 7891 719 7898 723
rect 7942 719 7948 723
rect 7991 719 7999 725
rect 8003 719 8005 746
rect 8332 744 8338 750
rect 8340 744 8343 754
rect 8378 750 8379 763
rect 8484 757 8490 762
rect 8496 757 8497 762
rect 8529 758 8539 784
rect 8543 783 8547 784
rect 8602 783 8608 786
rect 8637 783 8638 786
rect 8700 784 8714 786
rect 8700 783 8706 784
rect 8738 783 8742 784
rect 8609 781 8611 782
rect 8611 780 8614 781
rect 8627 780 8637 783
rect 8556 775 8562 779
rect 8562 772 8567 775
rect 8614 772 8637 780
rect 8568 766 8592 772
rect 8627 769 8659 772
rect 8665 769 8738 783
rect 8746 780 8752 786
rect 8753 784 8754 785
rect 8794 784 8795 786
rect 8829 783 8832 788
rect 8838 787 8930 788
rect 8902 786 8930 787
rect 8879 785 8930 786
rect 8938 785 8941 799
rect 9016 797 9017 801
rect 9063 800 9074 814
rect 9098 804 9109 814
rect 9111 804 9127 814
rect 9164 807 9177 815
rect 9161 805 9177 807
rect 9207 805 9223 820
rect 9261 811 9263 841
rect 9267 831 9275 843
rect 9314 838 9354 843
rect 9357 842 9364 874
rect 9399 840 9407 852
rect 9411 842 9413 874
rect 9443 857 9448 874
rect 9443 842 9445 857
rect 9448 852 9449 856
rect 9411 840 9445 842
rect 9449 840 9457 852
rect 9364 838 9365 840
rect 9451 838 9453 840
rect 9354 837 9369 838
rect 9411 837 9412 838
rect 9363 836 9369 837
rect 9408 836 9410 837
rect 9245 809 9263 811
rect 9267 809 9275 821
rect 9324 805 9334 836
rect 9363 832 9378 836
rect 9366 808 9378 832
rect 9411 828 9423 836
rect 9433 828 9445 836
rect 9451 828 9465 838
rect 9412 820 9414 828
rect 9365 807 9378 808
rect 9150 804 9263 805
rect 9127 803 9263 804
rect 9015 791 9016 796
rect 9014 788 9015 791
rect 9074 789 9077 799
rect 9109 794 9117 800
rect 9127 795 9143 803
rect 9145 799 9263 803
rect 9334 801 9338 805
rect 9364 804 9378 807
rect 9399 815 9414 820
rect 9453 822 9465 828
rect 9453 820 9455 822
rect 9399 804 9415 815
rect 9453 805 9465 820
rect 9905 819 9906 1015
rect 10095 819 10096 1015
rect 10181 819 10182 1015
rect 10454 819 10455 1015
rect 10651 819 10652 1015
rect 10873 1013 10889 1015
rect 10895 1013 10907 1022
rect 10915 1020 10944 1023
rect 10944 1014 10948 1020
rect 11684 1018 11736 1020
rect 11956 1018 11970 1023
rect 12166 1020 12167 1023
rect 11656 1016 11736 1018
rect 11656 1015 11707 1016
rect 10948 1013 10949 1014
rect 11631 1013 11656 1015
rect 11678 1014 11684 1015
rect 11707 1014 11712 1015
rect 10869 1011 10873 1013
rect 10885 1010 10889 1013
rect 11597 1011 11627 1013
rect 11673 1012 11678 1014
rect 10861 998 10869 1010
rect 10868 988 10869 998
rect 10873 1007 10907 1010
rect 10873 1003 10875 1007
rect 10873 996 10874 1003
rect 10885 1001 10889 1007
rect 10904 1005 10907 1007
rect 10910 1004 10919 1010
rect 10872 994 10874 996
rect 10871 988 10877 994
rect 10882 988 10885 1001
rect 10865 982 10871 988
rect 10868 976 10869 982
rect 10872 962 10873 988
rect 10905 982 10907 1004
rect 10911 998 10919 1004
rect 10949 1001 10958 1010
rect 11480 1005 11494 1007
rect 11506 1005 11597 1011
rect 11669 1007 11673 1012
rect 11480 1004 11506 1005
rect 11480 1003 11494 1004
rect 11474 1002 11494 1003
rect 11515 1002 11520 1005
rect 11665 1002 11669 1007
rect 11712 1005 11729 1014
rect 11729 1004 11731 1005
rect 10917 988 10923 994
rect 10940 992 10949 1001
rect 11465 997 11489 1002
rect 11520 997 11526 1002
rect 11664 1001 11665 1002
rect 11736 1001 11753 1016
rect 11970 1015 11977 1018
rect 12165 1016 12166 1020
rect 11977 1014 11980 1015
rect 11980 1005 12002 1014
rect 12163 1012 12165 1016
rect 12203 1014 12207 1036
rect 12209 1027 12217 1039
rect 12475 1037 12487 1045
rect 12536 1041 12546 1045
rect 12547 1041 12553 1045
rect 12511 1037 12553 1041
rect 12605 1039 12611 1045
rect 12758 1044 12764 1050
rect 12804 1048 12814 1050
rect 14469 1048 14478 1057
rect 14534 1048 14543 1057
rect 12767 1044 12779 1048
rect 12789 1044 12801 1048
rect 12804 1044 12810 1048
rect 12752 1038 12758 1044
rect 12810 1038 12816 1044
rect 15448 1038 15454 1044
rect 15494 1038 15500 1044
rect 15756 1043 15768 1051
rect 15778 1043 15790 1051
rect 15798 1048 15807 1057
rect 15857 1051 15873 1052
rect 15752 1040 15754 1043
rect 15792 1040 15794 1043
rect 15851 1039 15862 1051
rect 16125 1048 16134 1057
rect 16190 1051 16199 1057
rect 16131 1045 16134 1047
rect 16138 1045 16144 1051
rect 16184 1048 16199 1051
rect 16325 1048 16334 1057
rect 16390 1050 16399 1057
rect 16184 1045 16190 1048
rect 12256 1020 12266 1036
rect 12287 1034 12299 1037
rect 12481 1036 12487 1037
rect 12533 1036 12536 1037
rect 12281 1033 12301 1034
rect 12475 1033 12481 1036
rect 12517 1033 12547 1036
rect 12281 1031 12287 1033
rect 12301 1031 12331 1033
rect 12278 1025 12281 1031
rect 12275 1022 12281 1025
rect 12333 1024 12354 1031
rect 12381 1024 12387 1030
rect 12002 1004 12005 1005
rect 11862 1001 11863 1004
rect 10923 982 10929 988
rect 10940 986 10944 992
rect 11452 989 11465 997
rect 11474 993 11489 997
rect 10938 974 10939 979
rect 11096 976 11112 984
rect 11279 976 11295 989
rect 11362 979 11379 989
rect 11438 981 11452 989
rect 11432 979 11438 981
rect 11379 978 11432 979
rect 11463 977 11471 989
rect 11475 987 11480 989
rect 11526 987 11539 997
rect 11096 974 11153 976
rect 10934 957 10938 972
rect 11096 968 11141 974
rect 11153 968 11157 974
rect 10872 944 10879 957
rect 10933 953 10934 956
rect 10932 949 10933 952
rect 10935 944 10949 953
rect 11080 952 11096 968
rect 11157 961 11162 968
rect 11344 952 11350 958
rect 11390 952 11396 958
rect 11463 956 11471 967
rect 11475 958 11477 987
rect 11725 984 11727 1001
rect 11731 999 11753 1001
rect 11731 989 11739 999
rect 11857 992 11862 1001
rect 12005 996 12026 1004
rect 12160 1002 12163 1011
rect 12203 1007 12205 1014
rect 12194 1005 12205 1007
rect 12209 1010 12217 1017
rect 12209 1005 12222 1010
rect 12207 1004 12208 1005
rect 12208 1001 12209 1002
rect 12213 1001 12222 1005
rect 12256 1002 12266 1018
rect 12275 1015 12278 1022
rect 12329 1018 12335 1024
rect 12387 1018 12393 1024
rect 12463 1021 12471 1033
rect 12475 1031 12509 1033
rect 12475 1030 12481 1031
rect 12475 1029 12478 1030
rect 12275 1014 12277 1015
rect 12275 1013 12279 1014
rect 12277 1001 12279 1013
rect 11915 995 11948 996
rect 12026 995 12028 996
rect 11950 993 11956 995
rect 11857 986 11863 992
rect 11915 987 11921 992
rect 11956 991 11960 993
rect 12028 991 12038 995
rect 12158 991 12160 999
rect 12200 993 12213 1001
rect 12275 998 12279 1001
rect 12463 999 12471 1011
rect 12475 1002 12477 1029
rect 12755 1024 12758 1036
rect 12810 1032 12813 1036
rect 15442 1032 15448 1038
rect 15500 1032 15506 1038
rect 12763 1018 12767 1032
rect 12810 1021 12826 1032
rect 15733 1031 15739 1037
rect 15744 1031 15752 1039
rect 15755 1037 15790 1039
rect 15755 1036 15756 1037
rect 15788 1036 15790 1037
rect 14475 1026 14478 1030
rect 12826 1018 12842 1021
rect 12552 1007 12553 1008
rect 12553 1005 12554 1006
rect 12475 1001 12478 1002
rect 12521 1001 12549 1002
rect 12475 999 12487 1001
rect 12521 1000 12547 1001
rect 12205 992 12213 993
rect 12266 991 12270 996
rect 12275 991 12280 998
rect 12475 995 12479 999
rect 12521 998 12543 1000
rect 12549 999 12553 1001
rect 12521 996 12536 998
rect 12475 993 12481 995
rect 12521 994 12537 996
rect 12547 995 12553 999
rect 12556 997 12561 1003
rect 12605 1001 12614 1010
rect 12740 1001 12749 1010
rect 12749 1000 12755 1001
rect 11584 981 11600 984
rect 11602 981 11618 984
rect 11578 978 11598 981
rect 11719 979 11731 984
rect 11855 979 11856 983
rect 11863 980 11869 986
rect 11873 983 11941 987
rect 11960 986 11972 991
rect 11622 974 11623 978
rect 11580 972 11672 974
rect 11719 972 11739 979
rect 11854 974 11855 979
rect 11873 977 11899 983
rect 11909 980 11915 983
rect 11941 977 11954 983
rect 11972 978 11993 986
rect 12038 978 12072 991
rect 12204 988 12205 990
rect 12142 979 12148 985
rect 12158 983 12159 987
rect 12201 985 12204 986
rect 11853 972 11854 974
rect 11891 972 11899 977
rect 11484 963 11580 972
rect 11622 969 11623 972
rect 11581 963 11593 965
rect 11484 960 11581 963
rect 11475 957 11479 958
rect 11484 957 11580 960
rect 11475 956 11484 957
rect 11458 955 11482 956
rect 11486 955 11509 956
rect 11458 953 11477 955
rect 11526 954 11541 957
rect 11451 952 11458 953
rect 11471 952 11472 953
rect 11087 944 11096 952
rect 11338 946 11344 952
rect 11396 946 11402 952
rect 11432 949 11451 952
rect 11519 951 11526 954
rect 11475 950 11486 951
rect 11517 950 11519 951
rect 11410 946 11432 949
rect 11402 945 11424 946
rect 10865 936 10871 942
rect 10879 939 10891 944
rect 10927 942 10935 944
rect 10923 939 10935 942
rect 11085 939 11087 944
rect 11475 943 11487 950
rect 11090 940 11096 941
rect 11090 939 11132 940
rect 11136 939 11142 941
rect 10871 930 10877 936
rect 10891 934 10904 939
rect 10919 936 10929 939
rect 10917 934 10927 936
rect 11083 935 11085 939
rect 11090 936 11101 939
rect 11090 935 11096 936
rect 11132 935 11142 939
rect 11083 934 11090 935
rect 10910 929 10913 934
rect 10917 930 10923 934
rect 10908 926 10910 929
rect 10906 923 10908 926
rect 11080 925 11083 934
rect 11084 929 11090 934
rect 11142 929 11148 935
rect 11149 933 11161 941
rect 11222 934 11228 940
rect 11268 934 11274 940
rect 11538 939 11539 954
rect 11568 952 11578 957
rect 11577 939 11578 952
rect 11623 952 11634 968
rect 11595 942 11603 944
rect 11623 943 11626 952
rect 11664 947 11665 968
rect 11672 965 11744 972
rect 11668 963 11744 965
rect 11672 956 11744 963
rect 11753 962 11754 968
rect 11747 956 11754 962
rect 11793 956 11799 962
rect 11848 956 11853 972
rect 11715 955 11756 956
rect 11741 950 11756 955
rect 11799 950 11805 956
rect 11630 942 11676 944
rect 11585 940 11595 942
rect 11676 940 11684 942
rect 11583 939 11585 940
rect 11684 939 11687 940
rect 11163 932 11165 933
rect 11136 927 11161 929
rect 11078 924 11080 925
rect 10901 914 10906 923
rect 10994 922 11024 924
rect 11074 922 11078 924
rect 10899 907 10901 914
rect 10867 895 10868 905
rect 10897 896 10899 907
rect 10970 906 10994 922
rect 11024 916 11074 922
rect 11159 915 11161 927
rect 11165 917 11173 929
rect 11210 926 11222 934
rect 11274 928 11280 934
rect 11396 926 11399 930
rect 11525 927 11583 939
rect 11626 938 11627 939
rect 11595 930 11607 938
rect 11617 930 11629 938
rect 11520 926 11525 927
rect 11279 922 11281 924
rect 11159 906 11162 915
rect 11198 910 11206 922
rect 11210 920 11228 922
rect 10896 891 10897 895
rect 10895 888 10896 891
rect 10957 886 10970 906
rect 11159 902 11161 906
rect 11144 897 11161 902
rect 11136 896 11161 897
rect 11135 895 11161 896
rect 11165 895 11173 907
rect 11084 886 11090 889
rect 11132 886 11161 895
rect 11164 892 11165 894
rect 11198 888 11206 900
rect 11210 890 11212 920
rect 11281 916 11288 922
rect 11288 914 11291 916
rect 11399 914 11413 926
rect 11506 923 11520 926
rect 11529 924 11538 927
rect 11627 926 11629 930
rect 11687 927 11734 939
rect 11747 935 11756 950
rect 11846 949 11848 956
rect 11864 952 11873 968
rect 11882 955 11891 972
rect 11954 968 11971 977
rect 11993 968 12032 978
rect 11845 946 11846 949
rect 11749 934 11750 935
rect 11799 933 11805 936
rect 11734 926 11739 927
rect 11747 926 11749 933
rect 11805 930 11812 933
rect 11822 930 11834 938
rect 11842 937 11844 942
rect 11864 937 11873 950
rect 11879 946 11882 955
rect 11924 954 11953 964
rect 11971 963 12032 968
rect 11971 957 11993 963
rect 12032 960 12042 963
rect 11917 945 11953 954
rect 11964 952 11973 954
rect 11876 937 11878 942
rect 11835 926 11842 937
rect 11864 934 11876 937
rect 11908 936 11917 945
rect 11924 944 11953 945
rect 11954 945 11973 952
rect 11993 950 12014 957
rect 12042 956 12052 960
rect 12072 956 12129 978
rect 12148 973 12154 979
rect 12159 977 12160 983
rect 12200 979 12206 985
rect 12160 972 12161 977
rect 12194 974 12200 979
rect 12201 974 12204 979
rect 12194 973 12201 974
rect 12200 972 12201 973
rect 12158 968 12161 972
rect 12209 971 12211 991
rect 12270 985 12276 991
rect 12281 988 12282 990
rect 12283 986 12286 987
rect 12286 985 12291 986
rect 12270 984 12326 985
rect 12475 984 12486 993
rect 12521 990 12533 994
rect 12547 993 12561 995
rect 12605 993 12611 999
rect 12749 998 12756 1000
rect 12758 998 12767 1018
rect 12842 1015 12855 1018
rect 13479 1015 13480 1026
rect 13669 1015 13670 1026
rect 13755 1015 13756 1026
rect 14028 1015 14029 1026
rect 14225 1015 14226 1026
rect 14461 1023 14500 1026
rect 15502 1023 15541 1028
rect 15727 1025 15733 1031
rect 15753 1026 15755 1035
rect 15756 1031 15757 1036
rect 15752 1024 15753 1026
rect 14458 1022 14461 1023
rect 14458 1015 14470 1022
rect 14475 1020 14478 1023
rect 14474 1016 14475 1019
rect 12855 1001 12919 1015
rect 12919 998 12929 1001
rect 12549 992 12559 993
rect 12596 992 12605 993
rect 12749 992 12767 998
rect 12810 992 12816 998
rect 12929 992 12974 998
rect 13069 994 13087 995
rect 13057 992 13069 994
rect 12521 986 12539 990
rect 12553 987 12559 992
rect 12599 987 12605 992
rect 12758 991 12764 992
rect 12758 989 12765 991
rect 12766 990 12767 992
rect 12796 991 12799 992
rect 12758 986 12764 989
rect 12766 987 12770 988
rect 12785 987 12796 991
rect 12801 986 12810 992
rect 12929 988 13057 992
rect 12270 983 12335 984
rect 12479 983 12487 984
rect 12287 981 12335 983
rect 12287 979 12299 981
rect 12481 978 12497 983
rect 12502 981 12503 984
rect 12329 972 12335 978
rect 12387 972 12393 978
rect 12158 967 12163 968
rect 12199 967 12200 971
rect 12149 958 12163 967
rect 12052 954 12057 956
rect 12129 955 12148 956
rect 12149 955 12161 958
rect 12057 951 12064 954
rect 12129 951 12161 955
rect 12163 951 12164 957
rect 12064 950 12066 951
rect 11954 944 11966 945
rect 11924 943 11931 944
rect 11973 943 11982 945
rect 11924 942 11929 943
rect 11924 941 11926 942
rect 11924 940 11970 941
rect 11971 940 11982 943
rect 11920 939 11925 940
rect 11932 939 11966 940
rect 11920 938 11966 939
rect 11920 937 11932 938
rect 11869 926 11876 934
rect 11919 931 11932 937
rect 11963 936 11966 938
rect 11970 937 11982 940
rect 12014 943 12084 950
rect 12129 949 12149 951
rect 12152 949 12166 950
rect 12142 948 12166 949
rect 12142 946 12149 948
rect 12152 945 12169 948
rect 12194 946 12199 967
rect 12211 951 12213 968
rect 12335 966 12341 972
rect 12344 967 12347 972
rect 12213 949 12218 950
rect 12014 942 12087 943
rect 12014 939 12084 942
rect 12087 939 12096 942
rect 12152 939 12166 945
rect 12169 943 12179 945
rect 12208 943 12218 949
rect 12347 948 12354 967
rect 12381 966 12393 972
rect 12486 968 12497 978
rect 12521 980 12540 986
rect 12521 973 12558 980
rect 12682 976 12698 984
rect 12760 982 12763 986
rect 12759 976 12760 981
rect 12503 968 12506 972
rect 12387 945 12393 966
rect 12497 953 12509 968
rect 12525 965 12558 973
rect 12642 968 12645 976
rect 12683 975 12698 976
rect 12758 970 12759 975
rect 12801 969 12804 986
rect 12813 972 12914 977
rect 12914 969 12925 972
rect 12956 969 13057 988
rect 13087 980 13109 994
rect 12503 951 12506 953
rect 12509 951 12511 953
rect 12084 937 12116 939
rect 11964 931 11966 936
rect 11977 931 11983 937
rect 12084 934 12148 937
rect 12152 934 12168 939
rect 12179 934 12243 943
rect 12511 942 12531 951
rect 12540 948 12558 965
rect 12638 957 12642 968
rect 12633 955 12638 957
rect 12595 950 12596 953
rect 12356 939 12363 942
rect 12380 939 12420 942
rect 12344 936 12380 939
rect 12327 934 12344 936
rect 11920 930 11932 931
rect 11497 921 11506 923
rect 11485 920 11497 921
rect 11524 920 11529 924
rect 11438 915 11524 920
rect 11426 914 11438 915
rect 11466 914 11485 915
rect 11583 914 11591 926
rect 11595 924 11629 926
rect 11291 913 11421 914
rect 11399 909 11413 913
rect 11455 911 11466 914
rect 11448 907 11454 911
rect 11338 900 11344 906
rect 11344 894 11350 900
rect 11372 892 11385 900
rect 11415 892 11426 907
rect 11440 900 11445 904
rect 11577 901 11586 913
rect 11595 901 11597 924
rect 11210 888 11228 890
rect 11372 889 11381 892
rect 11385 891 11387 892
rect 11427 889 11429 891
rect 11437 889 11446 898
rect 11586 892 11597 901
rect 11627 892 11629 924
rect 11633 914 11641 926
rect 11739 924 11749 926
rect 11806 924 11834 926
rect 11835 924 11846 926
rect 11739 923 11747 924
rect 11744 921 11747 923
rect 11799 921 11800 924
rect 11832 921 11846 924
rect 11665 907 11679 921
rect 11734 910 11744 921
rect 11798 917 11799 921
rect 11734 907 11747 910
rect 11797 907 11798 916
rect 11832 915 11834 921
rect 11835 915 11846 921
rect 11869 924 11877 926
rect 11869 915 11876 924
rect 11877 921 11881 924
rect 11880 918 11886 921
rect 11881 916 11886 918
rect 11832 911 11835 915
rect 11837 914 11846 915
rect 11837 912 11838 914
rect 11679 906 11734 907
rect 11741 904 11747 907
rect 11796 904 11797 906
rect 11799 904 11805 910
rect 11832 906 11834 911
rect 11838 907 11840 912
rect 11840 906 11841 907
rect 11831 904 11834 906
rect 11841 904 11842 906
rect 11747 898 11753 904
rect 11789 902 11792 904
rect 11793 902 11799 904
rect 11788 898 11799 902
rect 11830 901 11831 904
rect 11788 892 11795 898
rect 11829 897 11830 900
rect 11827 894 11829 895
rect 11832 894 11834 904
rect 11800 892 11834 894
rect 11838 901 11846 904
rect 11838 892 11852 901
rect 11827 891 11829 892
rect 11852 890 11855 892
rect 10953 879 10957 885
rect 11079 879 11132 886
rect 11142 883 11148 886
rect 11149 883 11161 886
rect 11216 884 11222 888
rect 10950 875 10953 879
rect 11049 875 11079 879
rect 11090 877 11096 879
rect 10895 871 10896 875
rect 10947 870 10950 874
rect 11011 870 11049 875
rect 11009 869 11011 870
rect 10946 868 10947 869
rect 11007 868 11009 869
rect 11098 868 11100 879
rect 11133 868 11134 879
rect 11136 877 11142 883
rect 11210 882 11222 884
rect 11274 882 11280 888
rect 11210 876 11228 882
rect 11268 876 11274 882
rect 11381 880 11390 889
rect 11427 888 11437 889
rect 11825 888 11827 889
rect 11428 887 11437 888
rect 11428 880 11448 887
rect 11630 885 11631 888
rect 11591 882 11592 884
rect 11800 880 11812 888
rect 11822 882 11834 888
rect 11855 884 11857 890
rect 11859 885 11869 915
rect 11886 912 11899 916
rect 11899 907 11911 912
rect 11914 906 11916 907
rect 11925 906 11932 930
rect 11977 928 11978 931
rect 12100 919 12148 934
rect 12168 932 12243 934
rect 12260 933 12311 934
rect 12313 933 12324 934
rect 12260 932 12321 933
rect 12168 930 12260 932
rect 11916 904 11921 906
rect 11925 904 11977 906
rect 11921 901 11977 904
rect 11925 899 11977 901
rect 11908 889 11917 898
rect 11925 896 11994 899
rect 11925 891 11982 896
rect 11994 892 12019 896
rect 12116 894 12124 919
rect 12148 916 12155 919
rect 12168 918 12184 930
rect 12186 918 12202 930
rect 12307 929 12322 932
rect 12303 927 12307 929
rect 12287 922 12303 927
rect 12313 926 12322 929
rect 12356 926 12363 936
rect 12316 920 12321 922
rect 12134 900 12138 916
rect 12155 914 12186 916
rect 12187 914 12189 918
rect 12155 909 12187 914
rect 12178 907 12195 909
rect 12178 902 12187 907
rect 12195 906 12199 907
rect 12138 896 12139 899
rect 12158 898 12178 902
rect 11919 889 11983 891
rect 12019 890 12031 892
rect 12115 890 12116 893
rect 11917 885 11983 889
rect 11821 880 11834 882
rect 11391 875 11394 880
rect 11435 879 11448 880
rect 10933 864 10946 868
rect 11001 864 11007 868
rect 10927 862 10933 864
rect 10998 862 11001 864
rect 10924 858 10927 862
rect 10991 857 10998 862
rect 10923 856 10924 857
rect 10990 856 10991 857
rect 10922 849 10923 856
rect 10987 849 10990 856
rect 10921 841 10922 849
rect 10989 838 10998 842
rect 11036 838 11045 842
rect 11048 838 11064 854
rect 11066 838 11082 854
rect 11100 838 11104 867
rect 11131 847 11133 867
rect 11394 860 11401 875
rect 11433 873 11448 875
rect 11144 849 11158 854
rect 11240 842 11244 856
rect 9455 804 9465 805
rect 10917 804 10921 838
rect 10986 833 10998 838
rect 11032 833 11048 838
rect 11082 837 11098 838
rect 11089 834 11098 837
rect 10980 832 10993 833
rect 11032 832 11054 833
rect 10978 831 10987 832
rect 10978 811 10980 831
rect 10981 826 10987 831
rect 10977 810 10980 811
rect 10978 804 10980 810
rect 10986 820 10987 826
rect 11019 824 11054 832
rect 11019 823 11048 824
rect 11019 822 11067 823
rect 11093 822 11098 834
rect 11019 820 11039 822
rect 11048 820 11067 822
rect 10986 804 11002 820
rect 11032 804 11048 820
rect 11092 812 11093 817
rect 9363 803 9364 804
rect 9362 801 9363 802
rect 9310 799 9353 801
rect 9145 796 9310 799
rect 9145 795 9251 796
rect 9334 795 9353 799
rect 9127 794 9161 795
rect 9109 792 9143 794
rect 9088 789 9117 792
rect 9003 785 9014 788
rect 9063 787 9088 789
rect 9050 786 9063 787
rect 9046 785 9050 786
rect 8905 784 8908 785
rect 8926 784 9014 785
rect 8926 783 9003 784
rect 9019 783 9046 785
rect 9074 784 9077 787
rect 8748 779 8749 780
rect 8786 769 8794 783
rect 8828 778 8829 783
rect 8904 781 8905 783
rect 8927 782 8929 783
rect 8903 778 8904 781
rect 8929 780 8932 782
rect 8937 781 8938 783
rect 8995 782 9019 783
rect 8984 779 8995 782
rect 8932 778 8935 779
rect 8484 756 8502 757
rect 8530 756 8536 758
rect 8478 750 8542 756
rect 8567 753 8597 766
rect 8627 763 8665 769
rect 8783 763 8786 769
rect 8627 759 8659 763
rect 8626 756 8627 758
rect 8567 750 8603 753
rect 8624 752 8626 756
rect 8628 755 8659 759
rect 8656 754 8658 755
rect 8659 754 8662 755
rect 8778 754 8783 763
rect 8655 752 8656 754
rect 8662 751 8667 754
rect 8777 752 8778 754
rect 8378 744 8384 750
rect 8484 745 8536 750
rect 8288 742 8332 744
rect 8137 741 8171 742
rect 8288 741 8294 742
rect 8100 740 8137 741
rect 8077 739 8100 740
rect 8074 737 8077 739
rect 8326 738 8332 742
rect 8384 738 8390 744
rect 8049 723 8074 737
rect 8165 730 8171 736
rect 8223 731 8229 736
rect 8478 733 8490 745
rect 8524 735 8529 745
rect 8254 731 8290 733
rect 8171 724 8177 730
rect 8195 729 8254 731
rect 8290 729 8296 731
rect 8193 726 8195 729
rect 8044 720 8049 723
rect 7942 717 8024 719
rect 7945 716 8024 717
rect 8041 716 8049 720
rect 7991 713 7999 716
rect 8003 715 8005 716
rect 8024 715 8053 716
rect 8003 713 8037 715
rect 8034 709 8037 713
rect 8041 713 8049 715
rect 8053 714 8081 715
rect 8041 711 8044 713
rect 8038 709 8041 711
rect 8081 710 8095 714
rect 8187 713 8193 726
rect 8217 724 8223 729
rect 8296 726 8307 729
rect 8484 726 8490 733
rect 8286 722 8288 723
rect 8307 722 8318 726
rect 8483 723 8490 726
rect 8318 721 8320 722
rect 8320 720 8324 721
rect 7668 707 7669 708
rect 7890 707 7891 708
rect 8003 701 8015 709
rect 8025 701 8037 709
rect 8095 705 8101 710
rect 8185 708 8187 713
rect 8184 707 8185 708
rect 8101 703 8112 705
rect 7729 697 7863 700
rect 8029 698 8033 701
rect 8112 699 8125 703
rect 8125 698 8130 699
rect 7605 695 7729 697
rect 7863 695 7869 697
rect 7508 692 7514 694
rect 7583 692 7605 695
rect 7869 692 7875 695
rect 7290 688 7291 690
rect 7504 688 7506 691
rect 7507 688 7508 690
rect 7560 689 7583 692
rect 7875 689 7881 692
rect 8013 690 8029 698
rect 8130 694 8146 698
rect 8146 692 8162 694
rect 8162 691 8171 692
rect 8177 691 8184 706
rect 8278 693 8286 698
rect 8290 693 8292 720
rect 8478 711 8490 723
rect 8529 711 8531 726
rect 8567 723 8597 750
rect 8623 749 8624 751
rect 8667 750 8669 751
rect 8607 746 8609 747
rect 8621 745 8623 749
rect 8610 737 8624 745
rect 8652 744 8654 749
rect 8672 747 8675 749
rect 8675 746 8677 747
rect 8677 743 8681 746
rect 8701 743 8713 749
rect 8772 744 8775 749
rect 8807 744 8828 778
rect 8894 756 8903 778
rect 8932 776 8937 778
rect 8938 776 8984 779
rect 9077 778 9078 781
rect 8932 775 8984 776
rect 8932 756 8937 775
rect 9078 772 9082 778
rect 9078 756 9085 772
rect 9109 756 9117 789
rect 9127 788 9143 792
rect 9145 788 9161 794
rect 9223 788 9239 795
rect 9337 788 9353 795
rect 9340 787 9341 788
rect 9341 783 9342 785
rect 9343 772 9346 779
rect 9366 778 9378 804
rect 9415 799 9416 802
rect 9415 796 9417 799
rect 9453 796 9455 800
rect 10921 799 10934 804
rect 10951 799 10986 804
rect 10934 797 10951 799
rect 9415 791 9423 796
rect 9450 791 9453 796
rect 9415 788 9431 791
rect 9433 788 9449 791
rect 10970 788 10987 799
rect 11048 797 11051 803
rect 11048 795 11052 797
rect 11048 788 11058 795
rect 10978 786 10987 788
rect 11052 786 11058 788
rect 11103 786 11104 828
rect 11128 822 11141 838
rect 11274 833 11278 838
rect 11296 837 11308 845
rect 11362 838 11378 854
rect 11401 842 11410 860
rect 11402 841 11410 842
rect 11414 845 11415 862
rect 11414 843 11418 845
rect 11446 844 11448 873
rect 11449 869 11460 875
rect 11452 863 11460 869
rect 11456 859 11459 863
rect 11592 860 11596 879
rect 11629 866 11630 880
rect 11711 867 11717 873
rect 11757 867 11763 873
rect 11821 870 11825 880
rect 11854 870 11859 884
rect 11917 880 11931 885
rect 11925 871 11931 880
rect 11967 880 11977 885
rect 11967 870 11968 880
rect 11971 879 11977 880
rect 12031 879 12098 890
rect 12114 885 12115 889
rect 12113 881 12114 885
rect 12099 875 12103 879
rect 12103 872 12106 875
rect 12110 871 12113 881
rect 12139 879 12143 896
rect 12153 891 12158 898
rect 12199 892 12256 906
rect 12256 891 12259 892
rect 12150 881 12152 889
rect 12259 888 12273 891
rect 12319 890 12321 920
rect 12325 910 12333 922
rect 12363 914 12368 926
rect 12368 902 12373 914
rect 12393 910 12400 939
rect 12420 936 12426 939
rect 12426 934 12430 936
rect 12507 935 12508 942
rect 12531 939 12537 942
rect 12537 936 12543 939
rect 12430 933 12431 934
rect 12431 927 12434 933
rect 12434 922 12437 927
rect 12437 919 12439 922
rect 12439 916 12440 919
rect 12290 888 12321 890
rect 12325 888 12333 900
rect 12373 899 12374 902
rect 12400 900 12402 910
rect 12440 902 12447 916
rect 12508 910 12512 935
rect 12543 934 12547 936
rect 12558 935 12559 942
rect 12545 933 12551 934
rect 12545 932 12553 933
rect 12559 932 12560 935
rect 12595 934 12610 950
rect 12633 948 12645 955
rect 12632 947 12645 948
rect 12655 947 12667 955
rect 12698 952 12714 968
rect 12629 945 12638 947
rect 12628 943 12629 945
rect 12632 943 12638 945
rect 12671 943 12672 945
rect 12678 943 12684 948
rect 12621 942 12628 943
rect 12632 942 12667 943
rect 12671 942 12684 943
rect 12621 937 12632 942
rect 12633 941 12667 942
rect 12619 934 12625 937
rect 12626 936 12632 937
rect 12666 936 12667 941
rect 12684 936 12690 942
rect 12698 934 12714 950
rect 12751 939 12758 968
rect 12804 956 12805 968
rect 12809 965 12810 969
rect 12925 968 12944 969
rect 12952 968 12956 969
rect 12916 964 12952 968
rect 13002 965 13006 969
rect 12750 934 12751 938
rect 12615 932 12619 934
rect 12553 931 12594 932
rect 12559 918 12576 931
rect 12578 926 12594 931
rect 12612 930 12615 932
rect 12605 926 12612 930
rect 12697 927 12698 931
rect 12749 927 12750 932
rect 12578 918 12605 926
rect 12696 920 12698 927
rect 12748 922 12749 927
rect 12759 922 12767 934
rect 12771 922 12773 956
rect 12809 951 12810 964
rect 12916 960 12964 964
rect 12907 954 12916 960
rect 12804 945 12805 951
rect 12810 936 12811 945
rect 12899 939 12907 954
rect 12945 949 12964 960
rect 12964 948 12966 949
rect 13006 948 13011 965
rect 13109 961 13112 980
rect 13112 954 13113 960
rect 12966 945 12970 948
rect 13011 945 13012 948
rect 12896 936 12899 939
rect 12811 928 12817 934
rect 12812 922 12817 928
rect 12891 928 12903 936
rect 12913 928 12925 936
rect 12970 934 12985 945
rect 13012 934 13016 945
rect 13113 941 13116 954
rect 13115 939 13116 941
rect 13113 934 13115 939
rect 12985 932 12986 934
rect 12986 928 12987 930
rect 13016 929 13018 934
rect 12891 924 12896 928
rect 12929 926 12930 928
rect 12931 924 12934 925
rect 12695 919 12698 920
rect 12559 905 12560 918
rect 12587 916 12605 918
rect 12694 918 12698 919
rect 12694 916 12695 918
rect 12747 916 12748 919
rect 12767 916 12768 921
rect 12581 912 12587 916
rect 12690 909 12694 916
rect 12746 909 12747 916
rect 12768 912 12770 916
rect 12798 913 12805 922
rect 12812 916 12813 922
rect 12791 911 12798 913
rect 12809 911 12813 916
rect 12879 912 12887 924
rect 12891 922 12925 924
rect 12891 921 12894 922
rect 12771 910 12809 911
rect 12560 902 12561 904
rect 12447 899 12449 902
rect 12402 894 12403 899
rect 12449 896 12450 899
rect 12273 885 12284 888
rect 12287 885 12326 888
rect 12284 884 12326 885
rect 12143 872 12145 879
rect 12145 870 12146 872
rect 12147 871 12150 881
rect 12287 879 12326 884
rect 12375 881 12377 889
rect 12309 876 12321 879
rect 12326 874 12348 879
rect 12377 874 12378 881
rect 12362 872 12367 874
rect 11796 868 11797 869
rect 11820 867 11821 870
rect 11705 861 11711 867
rect 11763 861 11769 867
rect 11818 860 11820 867
rect 11459 854 11463 858
rect 11459 853 11474 854
rect 11445 843 11448 844
rect 11414 841 11448 843
rect 11452 841 11460 853
rect 11463 850 11474 853
rect 11596 852 11597 858
rect 11630 854 11631 858
rect 11465 845 11474 850
rect 11468 840 11474 845
rect 11231 831 11308 833
rect 11131 820 11136 822
rect 11128 804 11141 820
rect 11131 787 11136 804
rect 11144 788 11160 799
rect 10980 780 10987 786
rect 11045 785 11058 786
rect 11045 783 11092 785
rect 11020 780 11067 783
rect 8889 745 8894 756
rect 8929 744 8932 756
rect 9082 750 9085 756
rect 9082 744 9089 750
rect 9117 744 9119 756
rect 9147 751 9159 759
rect 9169 751 9181 759
rect 9346 755 9351 772
rect 9378 770 9382 778
rect 10980 777 10993 780
rect 11033 777 11039 780
rect 11045 779 11067 780
rect 11045 777 11054 779
rect 11231 777 11289 831
rect 11306 799 11308 831
rect 11312 821 11320 833
rect 11378 822 11394 838
rect 11448 837 11452 840
rect 11472 838 11474 840
rect 11496 838 11502 844
rect 11542 839 11548 844
rect 11538 838 11550 839
rect 11597 838 11600 850
rect 11632 841 11648 854
rect 11703 852 11711 858
rect 11701 850 11711 852
rect 11815 851 11818 860
rect 11764 848 11774 850
rect 11774 846 11780 848
rect 11813 847 11815 851
rect 11691 845 11699 846
rect 11701 845 11705 846
rect 11631 840 11648 841
rect 11631 838 11635 840
rect 11414 829 11426 837
rect 11436 829 11448 837
rect 11474 832 11554 838
rect 11600 832 11601 837
rect 11414 828 11415 829
rect 11415 818 11417 828
rect 11474 822 11490 832
rect 11496 831 11550 832
rect 11496 827 11548 831
rect 11417 814 11419 818
rect 11419 809 11420 812
rect 11420 805 11421 809
rect 11421 799 11422 803
rect 11422 792 11424 799
rect 11496 793 11516 827
rect 11542 825 11550 827
rect 11548 794 11550 825
rect 11554 815 11562 827
rect 11542 793 11550 794
rect 11554 793 11562 805
rect 11578 804 11586 820
rect 11601 814 11604 829
rect 11616 822 11635 838
rect 11669 833 11678 842
rect 11691 841 11701 845
rect 11703 844 11705 845
rect 11780 844 11787 846
rect 11703 841 11711 844
rect 11787 843 11791 844
rect 11791 842 11796 843
rect 11812 842 11813 844
rect 11808 841 11819 842
rect 11844 841 11854 869
rect 11859 866 11860 869
rect 11860 854 11863 865
rect 11931 860 11936 870
rect 12107 869 12110 870
rect 12106 865 12110 869
rect 12107 860 12110 865
rect 12137 866 12147 870
rect 12367 866 12384 872
rect 12403 871 12407 890
rect 12450 888 12454 896
rect 12558 890 12561 896
rect 12567 891 12578 908
rect 12633 903 12645 909
rect 12745 908 12746 909
rect 12674 903 12690 908
rect 12744 903 12745 908
rect 12791 903 12798 910
rect 12645 902 12674 903
rect 12743 896 12744 899
rect 12626 890 12632 896
rect 12684 890 12690 896
rect 12454 874 12462 888
rect 12556 885 12558 889
rect 12564 886 12567 890
rect 11936 854 11937 860
rect 12106 854 12109 860
rect 11860 852 11866 854
rect 11863 846 11866 852
rect 11928 849 11944 854
rect 11927 848 11941 849
rect 11946 848 11962 854
rect 11864 841 11866 846
rect 11924 845 11927 848
rect 11941 845 11962 848
rect 11919 841 11924 845
rect 11952 842 11964 845
rect 11691 838 11705 841
rect 11811 839 11812 841
rect 11819 840 11854 841
rect 11865 840 11866 841
rect 11917 840 11919 841
rect 11844 839 11892 840
rect 11915 838 11917 840
rect 11931 839 11943 842
rect 12024 841 12040 854
rect 12042 841 12058 854
rect 12104 847 12106 853
rect 12107 852 12109 854
rect 12137 852 12155 866
rect 12378 863 12393 866
rect 11964 840 11965 841
rect 12017 840 12018 841
rect 11936 838 11943 839
rect 11685 834 11699 838
rect 11685 833 11696 834
rect 11660 824 11669 833
rect 11631 820 11635 822
rect 11616 814 11635 820
rect 11604 809 11605 812
rect 11605 799 11607 808
rect 11616 804 11632 814
rect 11691 812 11699 824
rect 11703 814 11705 838
rect 11808 832 11811 838
rect 11763 815 11769 821
rect 11797 818 11815 832
rect 11803 815 11804 818
rect 11757 814 11763 815
rect 11802 814 11803 815
rect 11703 812 11737 814
rect 11746 812 11805 814
rect 11815 813 11821 818
rect 11816 812 11822 813
rect 11635 808 11636 812
rect 11727 809 11737 812
rect 11741 810 11746 812
rect 11718 808 11727 809
rect 11730 808 11736 809
rect 11738 808 11741 810
rect 11757 809 11763 812
rect 11636 804 11637 808
rect 11703 805 11715 808
rect 11718 805 11737 808
rect 11703 804 11716 805
rect 11632 794 11640 804
rect 11663 800 11715 804
rect 11725 800 11737 805
rect 11793 800 11802 811
rect 11805 810 11813 812
rect 11816 810 11827 812
rect 11835 811 11844 838
rect 11866 822 11882 838
rect 11906 832 11914 838
rect 11813 809 11827 810
rect 11829 809 11835 810
rect 11813 808 11835 809
rect 11866 808 11882 820
rect 11935 811 11937 838
rect 11938 837 11943 838
rect 11940 836 11943 837
rect 11965 838 11966 840
rect 12016 838 12017 840
rect 11941 834 11945 836
rect 11946 832 11947 834
rect 11965 832 11978 838
rect 11939 828 11943 830
rect 11816 804 11882 808
rect 11825 800 11866 804
rect 11906 801 11907 804
rect 11632 793 11642 794
rect 11496 792 11548 793
rect 11632 792 11644 793
rect 11424 789 11430 792
rect 11430 784 11437 789
rect 11490 788 11570 792
rect 11608 790 11609 792
rect 11632 789 11653 792
rect 11632 788 11647 789
rect 11490 786 11554 788
rect 11642 786 11647 788
rect 11653 787 11658 789
rect 11658 786 11662 787
rect 11663 786 11714 800
rect 11726 793 11730 800
rect 11788 793 11793 799
rect 11725 790 11726 793
rect 11786 790 11788 793
rect 11437 783 11438 784
rect 11473 783 11474 785
rect 11439 779 11445 783
rect 11470 779 11473 783
rect 11496 780 11502 786
rect 11538 781 11550 786
rect 11658 785 11669 786
rect 11660 783 11669 785
rect 11660 782 11672 783
rect 11542 780 11548 781
rect 11608 779 11609 781
rect 11445 777 11450 779
rect 11469 777 11470 779
rect 9129 747 9135 750
rect 9183 749 9185 750
rect 9138 747 9142 749
rect 9129 746 9138 747
rect 9128 744 9136 746
rect 9147 745 9183 747
rect 9185 745 9193 747
rect 8650 738 8652 743
rect 8681 741 8713 743
rect 8709 740 8714 741
rect 8716 737 8719 739
rect 8769 738 8772 744
rect 8804 739 8807 744
rect 8887 740 8889 744
rect 8904 740 8916 742
rect 8617 734 8618 737
rect 8624 734 8628 737
rect 8616 732 8617 734
rect 8628 732 8632 734
rect 8648 732 8650 737
rect 8678 736 8679 737
rect 8708 734 8718 737
rect 8719 734 8725 737
rect 8731 734 8737 737
rect 8713 732 8718 734
rect 8613 725 8616 731
rect 8632 729 8636 732
rect 8646 729 8648 731
rect 8612 722 8613 724
rect 8608 711 8612 721
rect 8636 712 8664 729
rect 8677 726 8678 731
rect 8718 727 8722 732
rect 8724 731 8737 734
rect 8762 732 8766 734
rect 8760 731 8762 732
rect 8777 731 8783 737
rect 8867 734 8873 740
rect 8885 734 8886 736
rect 8904 734 8919 740
rect 8928 738 8929 742
rect 9077 738 9083 744
rect 9135 738 9141 744
rect 9147 743 9149 745
rect 8927 734 8928 737
rect 8800 732 8801 734
rect 8861 732 8925 734
rect 8722 726 8724 727
rect 8725 726 8731 731
rect 8479 710 8483 711
rect 8484 710 8536 711
rect 8478 706 8542 710
rect 8473 704 8542 706
rect 8605 704 8608 711
rect 8332 698 8338 699
rect 8346 698 8384 699
rect 8326 695 8338 698
rect 8342 695 8390 698
rect 8326 693 8332 695
rect 8342 693 8380 695
rect 8384 693 8390 695
rect 8278 692 8390 693
rect 8278 691 8372 692
rect 7881 688 7884 689
rect 7888 688 7890 690
rect 5824 674 5827 685
rect 5140 653 5141 655
rect 5283 654 5284 656
rect 4072 651 4074 652
rect 3939 649 4015 651
rect 4067 649 4072 651
rect 4307 649 4311 652
rect 4370 650 4372 652
rect 4360 649 4370 650
rect 4022 648 4066 649
rect 4318 640 4334 649
rect 4335 648 4336 649
rect 4600 647 4602 651
rect 4620 647 4732 652
rect 4614 644 4732 647
rect 4830 644 4979 652
rect 4614 640 4630 644
rect 4732 641 4743 644
rect 4783 641 4830 644
rect 4743 640 4783 641
rect 4920 640 4936 644
rect 4982 636 5012 652
rect 5120 640 5136 653
rect 5283 644 5293 654
rect 5556 652 5569 660
rect 5624 656 5640 672
rect 5762 665 5771 674
rect 5824 667 5836 674
rect 7291 669 7301 688
rect 7502 682 7508 688
rect 7560 682 7566 688
rect 7884 686 7890 688
rect 7507 680 7520 682
rect 7507 676 7514 680
rect 7554 676 7560 682
rect 7888 677 7890 686
rect 7990 681 8013 690
rect 8171 689 8193 691
rect 8278 689 8368 691
rect 7990 679 8060 681
rect 5827 665 5836 667
rect 5764 656 5765 665
rect 5771 656 5780 665
rect 5818 656 5832 665
rect 7301 658 7311 669
rect 7303 656 7317 658
rect 7353 656 7369 672
rect 7507 668 7508 676
rect 7884 671 7890 677
rect 7942 678 8013 679
rect 7942 676 8006 678
rect 8060 676 8069 679
rect 7942 671 7948 676
rect 7507 656 7519 668
rect 7887 665 7896 671
rect 7936 665 7942 671
rect 7887 662 7890 665
rect 7971 662 7990 676
rect 8069 675 8073 676
rect 8073 672 8075 675
rect 8077 667 8078 669
rect 7887 658 7889 662
rect 7967 659 7971 662
rect 8078 660 8093 667
rect 8177 662 8183 689
rect 8193 686 8228 689
rect 8278 686 8362 689
rect 8378 686 8384 692
rect 8473 690 8478 704
rect 8484 699 8502 704
rect 8484 698 8490 699
rect 8530 698 8536 704
rect 8603 699 8605 704
rect 8531 696 8532 698
rect 8601 695 8603 698
rect 8637 695 8645 712
rect 8665 709 8668 711
rect 8673 709 8677 726
rect 8724 717 8734 726
rect 8783 725 8789 731
rect 8796 725 8800 732
rect 8861 730 8919 732
rect 8920 730 8925 732
rect 8926 730 8927 732
rect 8861 728 8917 730
rect 8794 722 8795 724
rect 8734 709 8736 717
rect 8788 711 8794 721
rect 8668 708 8670 709
rect 8667 707 8671 708
rect 8667 703 8673 707
rect 8679 705 8680 707
rect 8679 703 8696 705
rect 8598 694 8601 695
rect 8594 692 8598 694
rect 8592 691 8594 692
rect 8228 684 8247 686
rect 8286 684 8350 686
rect 8247 683 8255 684
rect 8255 681 8276 683
rect 8286 681 8345 684
rect 8276 679 8345 681
rect 8469 679 8473 689
rect 8532 686 8534 690
rect 8588 689 8592 691
rect 8584 688 8588 689
rect 8634 688 8637 695
rect 8670 690 8673 703
rect 8676 699 8678 700
rect 8679 696 8703 699
rect 8679 691 8691 696
rect 8703 693 8717 696
rect 8736 693 8738 706
rect 8783 702 8788 711
rect 8867 696 8882 728
rect 8914 726 8917 728
rect 8920 726 8928 730
rect 8914 724 8916 726
rect 8915 700 8916 724
rect 8917 718 8928 726
rect 8917 714 8921 718
rect 8917 710 8920 714
rect 8923 712 8925 718
rect 9179 715 9181 745
rect 9183 742 9193 745
rect 9353 743 9355 749
rect 9363 743 9369 749
rect 9382 746 9405 770
rect 10867 755 10868 775
rect 10896 772 10897 775
rect 10987 774 11026 777
rect 11033 774 11045 777
rect 10897 759 10905 772
rect 10989 768 11026 774
rect 11036 768 11045 774
rect 11102 768 11103 777
rect 10897 755 10908 759
rect 10868 749 10869 755
rect 10905 753 10908 755
rect 10906 750 10911 753
rect 9409 743 9415 749
rect 10880 747 10909 748
rect 10912 747 10913 749
rect 9357 742 9363 743
rect 9185 738 9193 742
rect 9185 735 9203 738
rect 9193 731 9203 735
rect 9355 731 9363 742
rect 9368 738 9369 742
rect 9401 739 9407 742
rect 9366 731 9368 738
rect 9402 737 9407 739
rect 9415 737 9421 743
rect 9153 714 9181 715
rect 9148 713 9181 714
rect 9185 713 9193 725
rect 9203 721 9209 731
rect 9355 721 9366 731
rect 9347 720 9366 721
rect 9347 712 9356 720
rect 8922 710 8923 711
rect 8920 707 8924 710
rect 9182 709 9185 711
rect 9156 708 9159 709
rect 8919 702 8924 707
rect 9144 706 9154 708
rect 9135 704 9144 706
rect 8914 696 8916 699
rect 8717 692 8783 693
rect 8723 691 8783 692
rect 8557 686 8584 688
rect 8633 686 8634 688
rect 8532 684 8564 686
rect 8522 683 8564 684
rect 8495 681 8564 683
rect 8477 679 8564 681
rect 8630 679 8633 684
rect 8286 678 8345 679
rect 8289 677 8324 678
rect 8450 677 8564 679
rect 8289 676 8321 677
rect 8323 676 8324 677
rect 8290 674 8302 676
rect 8304 675 8323 676
rect 8428 675 8450 677
rect 8456 676 8564 677
rect 8469 675 8473 676
rect 8304 671 8331 675
rect 8380 671 8428 675
rect 8304 670 8342 671
rect 8369 670 8412 671
rect 8304 664 8412 670
rect 8306 662 8316 664
rect 8469 662 8470 675
rect 8534 672 8536 675
rect 8627 673 8630 679
rect 8183 660 8184 662
rect 7965 658 7967 659
rect 7667 656 7669 657
rect 7887 656 7888 658
rect 7963 656 7965 658
rect 5591 652 5624 656
rect 5824 652 5827 656
rect 5571 651 5590 652
rect 5339 645 5340 651
rect 5294 640 5310 644
rect 5312 640 5328 644
rect 5608 640 5624 652
rect 5765 645 5775 652
rect 5819 646 5824 652
rect 5813 645 5819 646
rect 5775 644 5816 645
rect 5800 640 5816 644
rect 7319 640 7335 656
rect 7337 640 7353 656
rect 7520 653 7522 656
rect 7660 653 7666 656
rect 7889 653 7892 656
rect 7959 653 7963 656
rect 7522 651 7524 653
rect 7659 652 7660 653
rect 7957 652 7959 653
rect 8093 652 8205 660
rect 8297 658 8306 662
rect 8534 659 8537 672
rect 8666 666 8670 689
rect 8729 685 8783 691
rect 8867 688 8919 696
rect 8920 692 8924 702
rect 9077 693 9083 698
rect 9135 693 9141 698
rect 9077 692 9141 693
rect 8924 688 8926 690
rect 8725 679 8789 685
rect 8861 682 8926 688
rect 9083 686 9089 692
rect 9129 686 9135 692
rect 9147 690 9148 706
rect 9169 701 9181 709
rect 9360 707 9366 720
rect 9403 717 9407 737
rect 9359 706 9360 707
rect 9355 697 9359 706
rect 9407 697 9409 717
rect 10170 703 10192 722
rect 10862 713 10869 725
rect 10874 716 10875 747
rect 10903 745 10908 747
rect 10907 716 10908 745
rect 10909 738 10920 747
rect 11136 740 11140 777
rect 11445 776 11469 777
rect 11606 775 11608 779
rect 11660 777 11669 782
rect 11675 779 11678 781
rect 11678 777 11697 779
rect 11725 777 11734 786
rect 11756 782 11762 788
rect 11783 786 11786 790
rect 11802 782 11808 788
rect 11820 786 11829 800
rect 11832 788 11848 800
rect 11850 796 11886 800
rect 11907 798 11909 801
rect 11934 800 11935 810
rect 11941 798 11943 828
rect 11947 818 11955 830
rect 11964 822 11978 832
rect 12008 836 12016 838
rect 12070 837 12074 841
rect 12102 839 12104 847
rect 12137 838 12147 852
rect 12155 848 12158 852
rect 12285 842 12291 844
rect 12285 838 12299 842
rect 12331 838 12337 844
rect 12338 838 12354 854
rect 12378 838 12384 863
rect 12393 853 12396 863
rect 12396 846 12398 852
rect 12398 838 12401 845
rect 12008 822 12015 836
rect 12032 826 12044 832
rect 12029 825 12088 826
rect 12092 825 12102 838
rect 12029 823 12037 825
rect 12088 823 12102 825
rect 12109 823 12112 838
rect 11964 820 11967 822
rect 12028 821 12029 823
rect 11907 796 11943 798
rect 11947 796 11955 808
rect 11964 804 11978 820
rect 12020 816 12028 820
rect 12032 818 12039 820
rect 12020 808 12026 816
rect 12032 814 12033 818
rect 12092 816 12117 823
rect 12126 816 12137 837
rect 12158 822 12170 838
rect 12279 832 12285 838
rect 12283 830 12285 832
rect 12287 830 12320 838
rect 12337 832 12343 838
rect 12354 832 12370 838
rect 12384 832 12385 838
rect 12337 830 12370 832
rect 12401 830 12404 838
rect 12407 830 12419 870
rect 12462 863 12467 874
rect 12509 871 12512 885
rect 12546 881 12556 885
rect 12632 884 12638 890
rect 12642 887 12643 890
rect 12652 886 12659 890
rect 12643 883 12646 885
rect 12649 884 12651 885
rect 12678 884 12684 890
rect 12741 888 12743 896
rect 12643 882 12648 883
rect 12544 874 12562 881
rect 12527 870 12544 874
rect 12546 870 12556 874
rect 12467 859 12469 863
rect 12493 838 12509 870
rect 12527 866 12546 870
rect 12525 863 12527 866
rect 12523 859 12525 863
rect 12539 859 12546 866
rect 12521 856 12523 859
rect 12519 854 12521 856
rect 12512 851 12521 854
rect 12512 845 12519 851
rect 12512 839 12516 845
rect 12512 838 12513 839
rect 12469 830 12470 838
rect 12493 830 12512 838
rect 12526 830 12539 859
rect 12556 846 12563 858
rect 12568 848 12569 880
rect 12635 876 12641 879
rect 12632 874 12635 876
rect 12623 869 12632 874
rect 12643 870 12646 882
rect 12680 870 12683 884
rect 12740 881 12741 888
rect 12739 874 12740 881
rect 12616 860 12617 863
rect 12646 860 12648 870
rect 12680 862 12694 870
rect 12736 863 12739 874
rect 12611 848 12616 860
rect 12568 847 12573 848
rect 12568 846 12602 847
rect 12609 846 12614 848
rect 12563 844 12564 846
rect 12608 844 12609 846
rect 12605 842 12607 843
rect 12568 834 12580 841
rect 12590 834 12602 841
rect 12648 830 12659 859
rect 12683 830 12694 862
rect 12735 856 12736 859
rect 12773 856 12791 903
rect 12879 890 12887 902
rect 12891 890 12893 921
rect 12924 920 12925 922
rect 12931 912 12937 924
rect 12987 913 12989 925
rect 13018 924 13034 928
rect 13104 925 13113 934
rect 13096 924 13104 925
rect 13018 913 13096 924
rect 12931 911 12934 912
rect 12934 903 12939 910
rect 12972 905 13034 913
rect 12966 903 12972 905
rect 12925 890 12966 903
rect 12934 888 12939 890
rect 12989 889 12991 905
rect 12887 886 12890 888
rect 12939 886 12940 888
rect 12991 885 12992 888
rect 12890 884 12892 885
rect 12891 883 12893 884
rect 12891 879 12894 883
rect 12940 880 12941 882
rect 12891 878 12895 879
rect 12894 876 12895 878
rect 12941 876 12942 880
rect 12992 876 12993 879
rect 13018 878 13034 905
rect 12895 869 12898 874
rect 12898 863 12900 869
rect 12833 861 12834 862
rect 12900 860 12901 863
rect 12712 851 12728 854
rect 12732 851 12735 856
rect 12771 851 12773 856
rect 12814 854 12826 855
rect 12712 845 12732 851
rect 12769 846 12771 851
rect 12808 847 12826 854
rect 12836 849 12848 855
rect 12836 847 12885 849
rect 12901 848 12905 860
rect 12808 845 12824 847
rect 12837 846 12885 847
rect 12830 845 12837 846
rect 12857 845 12885 846
rect 12712 843 12718 845
rect 12768 843 12769 845
rect 12808 843 12830 845
rect 12885 843 12899 845
rect 12905 844 12906 847
rect 12922 843 12938 854
rect 12710 839 12713 843
rect 12766 839 12768 843
rect 12802 842 12807 843
rect 12802 840 12806 842
rect 12808 841 12848 843
rect 12795 839 12805 840
rect 12808 839 12814 841
rect 12789 838 12794 839
rect 12808 838 12809 839
rect 12696 830 12710 838
rect 12763 836 12766 838
rect 12785 837 12789 838
rect 12776 836 12782 837
rect 12763 834 12776 836
rect 12753 833 12757 834
rect 12747 832 12753 833
rect 12734 830 12747 832
rect 12763 831 12766 834
rect 12275 827 12283 830
rect 12287 828 12290 830
rect 12274 821 12284 827
rect 11963 802 11964 804
rect 11965 800 11967 804
rect 12092 801 12102 816
rect 12104 812 12112 816
rect 12104 804 12113 812
rect 12117 807 12149 816
rect 12158 807 12170 820
rect 12250 807 12274 821
rect 12275 818 12283 821
rect 12113 801 12114 803
rect 12126 801 12137 807
rect 12149 804 12170 807
rect 11850 788 11866 796
rect 11886 795 11891 796
rect 11891 793 11902 795
rect 11909 794 11916 796
rect 11916 793 11922 794
rect 11933 793 11934 796
rect 11902 792 11907 793
rect 11922 792 11942 793
rect 11945 792 11947 795
rect 11962 794 11963 796
rect 11922 786 11943 792
rect 11959 789 11962 793
rect 11944 788 11962 789
rect 11944 786 11959 788
rect 12015 786 12016 788
rect 12020 786 12026 798
rect 12074 789 12075 801
rect 12089 790 12092 800
rect 12114 797 12142 801
rect 12149 797 12168 804
rect 12238 800 12250 807
rect 12236 799 12238 800
rect 12114 796 12168 797
rect 12229 796 12236 799
rect 12275 796 12283 808
rect 12287 796 12289 828
rect 12355 822 12584 830
rect 12355 820 12357 822
rect 12358 820 12584 822
rect 12355 814 12584 820
rect 12612 814 12734 830
rect 12757 818 12763 831
rect 12792 822 12808 838
rect 12755 815 12762 818
rect 12355 812 12612 814
rect 12357 804 12370 812
rect 12387 807 12389 812
rect 12357 803 12358 804
rect 12358 801 12359 802
rect 12355 796 12358 801
rect 12388 800 12389 807
rect 12400 804 12412 812
rect 12412 803 12413 804
rect 12417 803 12419 808
rect 12436 803 12515 812
rect 12413 802 12515 803
rect 12416 799 12432 802
rect 12033 787 12034 788
rect 12032 786 12038 787
rect 11814 782 11820 786
rect 11931 784 11943 786
rect 11605 772 11606 774
rect 11669 772 11697 777
rect 11598 759 11605 772
rect 11669 768 11678 772
rect 11716 768 11725 777
rect 11750 776 11756 782
rect 11808 776 11820 782
rect 11932 776 11933 781
rect 11808 766 11812 773
rect 11964 772 11965 786
rect 12016 783 12017 786
rect 12027 784 12029 785
rect 12073 784 12074 788
rect 12088 787 12089 790
rect 12114 789 12158 796
rect 12168 795 12170 796
rect 12170 792 12177 795
rect 12227 793 12229 796
rect 12326 795 12354 796
rect 12177 789 12181 792
rect 12114 788 12136 789
rect 12138 788 12154 789
rect 12181 788 12183 789
rect 12223 788 12227 793
rect 12338 792 12354 795
rect 12384 793 12388 799
rect 12095 787 12102 788
rect 12110 787 12124 788
rect 12183 787 12186 788
rect 12087 786 12095 787
rect 12082 785 12095 786
rect 12114 785 12124 787
rect 12279 786 12285 792
rect 12337 791 12354 792
rect 12381 791 12384 793
rect 12337 789 12393 791
rect 12414 789 12432 799
rect 12337 788 12354 789
rect 12381 788 12384 789
rect 12393 788 12432 789
rect 12434 788 12515 802
rect 12526 800 12539 812
rect 12602 804 12603 807
rect 12337 786 12343 788
rect 12380 786 12381 788
rect 12079 784 12088 785
rect 12017 780 12029 783
rect 12032 780 12033 781
rect 12041 780 12079 784
rect 12017 779 12076 780
rect 12032 774 12044 779
rect 11963 763 11965 772
rect 12082 763 12088 784
rect 12114 784 12128 785
rect 11588 756 11605 759
rect 11929 756 11932 763
rect 11588 755 11598 756
rect 11588 754 11595 755
rect 11928 754 11929 756
rect 11588 753 11592 754
rect 11577 749 11619 753
rect 11577 748 11604 749
rect 11575 747 11577 748
rect 11619 747 11622 749
rect 11561 745 11575 747
rect 11093 738 11099 740
rect 11136 739 11145 740
rect 10913 735 10931 738
rect 10920 725 10931 735
rect 11093 734 11105 738
rect 11139 734 11145 739
rect 11528 738 11561 745
rect 11522 737 11527 738
rect 11087 728 11093 734
rect 11145 729 11151 734
rect 11499 733 11522 737
rect 11576 735 11584 747
rect 11588 746 11593 747
rect 11493 731 11499 733
rect 11487 729 11489 731
rect 11109 728 11240 729
rect 11093 726 11109 728
rect 11145 727 11448 728
rect 11475 727 11481 729
rect 11486 728 11487 729
rect 11240 726 11241 727
rect 11448 726 11481 727
rect 11484 726 11486 728
rect 10874 714 10878 716
rect 10905 714 10908 716
rect 10874 713 10908 714
rect 10913 713 10931 725
rect 11081 714 11089 726
rect 11093 724 11099 726
rect 10869 711 10870 713
rect 10870 708 10875 711
rect 10908 708 10913 711
rect 10874 707 10886 708
rect 10141 697 10164 698
rect 10169 697 10192 703
rect 10873 701 10886 707
rect 10896 701 10908 708
rect 10920 707 10931 713
rect 9355 693 9363 697
rect 9415 693 9421 697
rect 10873 694 10875 701
rect 9355 691 9421 693
rect 9355 690 9359 691
rect 9148 686 9150 690
rect 8729 673 8737 679
rect 8777 673 8783 679
rect 8867 676 8873 682
rect 8913 676 8919 682
rect 8729 666 8736 673
rect 8869 672 8872 676
rect 8293 656 8297 658
rect 8470 656 8471 658
rect 8535 657 8537 659
rect 8533 656 8537 657
rect 8288 653 8293 656
rect 8471 653 8474 656
rect 8532 653 8533 656
rect 8567 654 8597 663
rect 8601 654 8614 660
rect 8666 659 8668 666
rect 8729 665 8737 666
rect 8283 652 8284 653
rect 8531 652 8532 653
rect 8564 652 8601 654
rect 8668 653 8670 659
rect 8726 656 8737 665
rect 8863 660 8872 672
rect 8925 672 8926 682
rect 8863 656 8869 660
rect 8925 656 8929 672
rect 9141 660 9150 686
rect 9349 674 9355 690
rect 9363 685 9369 691
rect 9409 685 9415 691
rect 10931 690 10938 707
rect 11081 692 11089 704
rect 11093 694 11095 724
rect 11242 719 11246 726
rect 11448 723 11483 726
rect 11521 723 11527 729
rect 11246 708 11253 719
rect 11469 717 11475 723
rect 11476 719 11483 723
rect 11527 719 11533 723
rect 11576 719 11584 725
rect 11588 719 11590 746
rect 11917 744 11923 750
rect 11925 744 11928 754
rect 11963 750 11964 763
rect 12069 757 12075 762
rect 12081 757 12082 762
rect 12114 758 12124 784
rect 12128 783 12132 784
rect 12187 783 12193 786
rect 12222 783 12223 786
rect 12285 784 12299 786
rect 12285 783 12291 784
rect 12323 783 12327 784
rect 12194 781 12196 782
rect 12196 780 12199 781
rect 12212 780 12222 783
rect 12141 775 12147 779
rect 12147 772 12152 775
rect 12199 772 12222 780
rect 12153 766 12177 772
rect 12212 769 12244 772
rect 12250 769 12323 783
rect 12331 780 12337 786
rect 12338 784 12339 785
rect 12379 784 12380 786
rect 12414 783 12417 788
rect 12423 787 12515 788
rect 12487 786 12515 787
rect 12464 785 12515 786
rect 12523 785 12526 799
rect 12601 797 12602 801
rect 12648 800 12659 814
rect 12683 804 12694 814
rect 12696 804 12712 814
rect 12749 807 12762 815
rect 12746 805 12762 807
rect 12792 805 12808 820
rect 12846 811 12848 841
rect 12852 831 12860 843
rect 12899 838 12939 843
rect 12942 842 12949 874
rect 12984 840 12992 852
rect 12996 842 12998 874
rect 13028 857 13033 874
rect 13028 842 13030 857
rect 13033 852 13034 856
rect 12996 840 13030 842
rect 13034 840 13042 852
rect 12949 838 12950 840
rect 13036 838 13038 840
rect 12939 837 12954 838
rect 12996 837 12997 838
rect 12948 836 12954 837
rect 12993 836 12995 837
rect 12830 809 12848 811
rect 12852 809 12860 821
rect 12909 805 12919 836
rect 12948 832 12963 836
rect 12951 808 12963 832
rect 12996 828 13008 836
rect 13018 828 13030 836
rect 13036 828 13050 838
rect 12997 820 12999 828
rect 12950 807 12963 808
rect 12735 804 12848 805
rect 12712 803 12848 804
rect 12600 791 12601 796
rect 12599 788 12600 791
rect 12659 789 12662 799
rect 12694 794 12702 800
rect 12712 795 12728 803
rect 12730 799 12848 803
rect 12919 801 12923 805
rect 12949 804 12963 807
rect 12984 815 12999 820
rect 13038 822 13050 828
rect 13038 820 13040 822
rect 12984 804 13000 815
rect 13038 805 13050 820
rect 13490 819 13491 1015
rect 13680 819 13681 1015
rect 13766 819 13767 1015
rect 14039 819 14040 1015
rect 14236 819 14237 1015
rect 14458 1013 14474 1015
rect 14480 1013 14492 1022
rect 14500 1020 14529 1023
rect 14529 1014 14533 1020
rect 15269 1018 15321 1020
rect 15541 1018 15555 1023
rect 15751 1020 15752 1023
rect 15241 1016 15321 1018
rect 15241 1015 15292 1016
rect 14533 1013 14534 1014
rect 15216 1013 15241 1015
rect 15263 1014 15269 1015
rect 15292 1014 15297 1015
rect 14454 1011 14458 1013
rect 14470 1010 14474 1013
rect 15182 1011 15212 1013
rect 15258 1012 15263 1014
rect 14446 998 14454 1010
rect 14453 988 14454 998
rect 14458 1007 14492 1010
rect 14458 1003 14460 1007
rect 14458 996 14459 1003
rect 14470 1001 14474 1007
rect 14489 1005 14492 1007
rect 14495 1004 14504 1010
rect 14457 994 14459 996
rect 14456 988 14462 994
rect 14467 988 14470 1001
rect 14450 982 14456 988
rect 14453 976 14454 982
rect 14457 962 14458 988
rect 14490 982 14492 1004
rect 14496 998 14504 1004
rect 14534 1001 14543 1010
rect 15065 1005 15079 1007
rect 15091 1005 15182 1011
rect 15254 1007 15258 1012
rect 15065 1004 15091 1005
rect 15065 1003 15079 1004
rect 15059 1002 15079 1003
rect 15100 1002 15105 1005
rect 15250 1002 15254 1007
rect 15297 1005 15314 1014
rect 15314 1004 15316 1005
rect 14502 988 14508 994
rect 14525 992 14534 1001
rect 15050 997 15074 1002
rect 15105 997 15111 1002
rect 15249 1001 15250 1002
rect 15321 1001 15338 1016
rect 15555 1015 15562 1018
rect 15750 1016 15751 1020
rect 15562 1014 15565 1015
rect 15565 1005 15587 1014
rect 15748 1012 15750 1016
rect 15788 1014 15792 1036
rect 15794 1027 15802 1039
rect 16060 1037 16072 1045
rect 16121 1041 16131 1045
rect 16132 1041 16138 1045
rect 16096 1037 16138 1041
rect 16190 1039 16196 1045
rect 16343 1044 16349 1050
rect 16389 1048 16399 1050
rect 18054 1048 18063 1057
rect 18119 1048 18128 1057
rect 16352 1044 16364 1048
rect 16374 1044 16386 1048
rect 16389 1044 16395 1048
rect 16337 1038 16343 1044
rect 16395 1038 16401 1044
rect 19033 1038 19039 1044
rect 19079 1038 19085 1044
rect 19341 1043 19353 1051
rect 19363 1043 19375 1051
rect 19383 1048 19392 1057
rect 19442 1051 19458 1052
rect 19337 1040 19339 1043
rect 19377 1040 19379 1043
rect 19436 1039 19447 1051
rect 19710 1048 19719 1057
rect 19775 1051 19784 1057
rect 19716 1045 19719 1047
rect 19723 1045 19729 1051
rect 19769 1048 19784 1051
rect 19910 1048 19919 1057
rect 19975 1050 19984 1057
rect 19769 1045 19775 1048
rect 15841 1020 15851 1036
rect 15872 1034 15884 1037
rect 16066 1036 16072 1037
rect 16118 1036 16121 1037
rect 15866 1033 15886 1034
rect 16060 1033 16066 1036
rect 16102 1033 16132 1036
rect 15866 1031 15872 1033
rect 15886 1031 15916 1033
rect 15863 1025 15866 1031
rect 15860 1022 15866 1025
rect 15918 1024 15939 1031
rect 15966 1024 15972 1030
rect 15587 1004 15590 1005
rect 15447 1001 15448 1004
rect 14508 982 14514 988
rect 14525 986 14529 992
rect 15037 989 15050 997
rect 15059 993 15074 997
rect 14523 974 14524 979
rect 14681 976 14697 984
rect 14864 976 14880 989
rect 14947 979 14964 989
rect 15023 981 15037 989
rect 15017 979 15023 981
rect 14964 978 15017 979
rect 15048 977 15056 989
rect 15060 987 15065 989
rect 15111 987 15124 997
rect 14681 974 14738 976
rect 14519 957 14523 972
rect 14681 968 14726 974
rect 14738 968 14742 974
rect 14457 944 14464 957
rect 14518 953 14519 956
rect 14517 949 14518 952
rect 14520 944 14534 953
rect 14665 952 14681 968
rect 14742 961 14747 968
rect 14929 952 14935 958
rect 14975 952 14981 958
rect 15048 956 15056 967
rect 15060 958 15062 987
rect 15310 984 15312 1001
rect 15316 999 15338 1001
rect 15316 989 15324 999
rect 15442 992 15447 1001
rect 15590 996 15611 1004
rect 15745 1002 15748 1011
rect 15788 1007 15790 1014
rect 15779 1005 15790 1007
rect 15794 1010 15802 1017
rect 15794 1005 15807 1010
rect 15792 1004 15793 1005
rect 15793 1001 15794 1002
rect 15798 1001 15807 1005
rect 15841 1002 15851 1018
rect 15860 1015 15863 1022
rect 15914 1018 15920 1024
rect 15972 1018 15978 1024
rect 16048 1021 16056 1033
rect 16060 1031 16094 1033
rect 16060 1030 16066 1031
rect 16060 1029 16063 1030
rect 15860 1014 15862 1015
rect 15860 1013 15864 1014
rect 15862 1001 15864 1013
rect 15500 995 15533 996
rect 15611 995 15613 996
rect 15535 993 15541 995
rect 15442 986 15448 992
rect 15500 987 15506 992
rect 15541 991 15545 993
rect 15613 991 15623 995
rect 15743 991 15745 999
rect 15785 993 15798 1001
rect 15860 998 15864 1001
rect 16048 999 16056 1011
rect 16060 1002 16062 1029
rect 16340 1024 16343 1036
rect 16395 1032 16398 1036
rect 19027 1032 19033 1038
rect 19085 1032 19091 1038
rect 16348 1018 16352 1032
rect 16395 1021 16411 1032
rect 19318 1031 19324 1037
rect 19329 1031 19337 1039
rect 19340 1037 19375 1039
rect 19340 1036 19341 1037
rect 19373 1036 19375 1037
rect 18060 1026 18063 1030
rect 16411 1018 16427 1021
rect 16137 1007 16138 1008
rect 16138 1005 16139 1006
rect 16060 1001 16063 1002
rect 16106 1001 16134 1002
rect 16060 999 16072 1001
rect 16106 1000 16132 1001
rect 15790 992 15798 993
rect 15851 991 15855 996
rect 15860 991 15865 998
rect 16060 995 16064 999
rect 16106 998 16128 1000
rect 16134 999 16138 1001
rect 16106 996 16121 998
rect 16060 993 16066 995
rect 16106 994 16122 996
rect 16132 995 16138 999
rect 16141 997 16146 1003
rect 16190 1001 16199 1010
rect 16325 1001 16334 1010
rect 16334 1000 16340 1001
rect 15169 981 15185 984
rect 15187 981 15203 984
rect 15163 978 15183 981
rect 15304 979 15316 984
rect 15440 979 15441 983
rect 15448 980 15454 986
rect 15458 983 15526 987
rect 15545 986 15557 991
rect 15207 974 15208 978
rect 15165 972 15257 974
rect 15304 972 15324 979
rect 15439 974 15440 979
rect 15458 977 15484 983
rect 15494 980 15500 983
rect 15526 977 15539 983
rect 15557 978 15578 986
rect 15623 978 15657 991
rect 15789 988 15790 990
rect 15727 979 15733 985
rect 15743 983 15744 987
rect 15786 985 15789 986
rect 15438 972 15439 974
rect 15476 972 15484 977
rect 15069 963 15165 972
rect 15207 969 15208 972
rect 15166 963 15178 965
rect 15069 960 15166 963
rect 15060 957 15064 958
rect 15069 957 15165 960
rect 15060 956 15069 957
rect 15043 955 15067 956
rect 15071 955 15094 956
rect 15043 953 15062 955
rect 15111 954 15126 957
rect 15036 952 15043 953
rect 15056 952 15057 953
rect 14672 944 14681 952
rect 14923 946 14929 952
rect 14981 946 14987 952
rect 15017 949 15036 952
rect 15104 951 15111 954
rect 15060 950 15071 951
rect 15102 950 15104 951
rect 14995 946 15017 949
rect 14987 945 15009 946
rect 14450 936 14456 942
rect 14464 939 14476 944
rect 14512 942 14520 944
rect 14508 939 14520 942
rect 14670 939 14672 944
rect 15060 943 15072 950
rect 14675 940 14681 941
rect 14675 939 14717 940
rect 14721 939 14727 941
rect 14456 930 14462 936
rect 14476 934 14489 939
rect 14504 936 14514 939
rect 14502 934 14512 936
rect 14668 935 14670 939
rect 14675 936 14686 939
rect 14675 935 14681 936
rect 14717 935 14727 939
rect 14668 934 14675 935
rect 14495 929 14498 934
rect 14502 930 14508 934
rect 14493 926 14495 929
rect 14491 923 14493 926
rect 14665 925 14668 934
rect 14669 929 14675 934
rect 14727 929 14733 935
rect 14734 933 14746 941
rect 14807 934 14813 940
rect 14853 934 14859 940
rect 15123 939 15124 954
rect 15153 952 15163 957
rect 15162 939 15163 952
rect 15208 952 15219 968
rect 15180 942 15188 944
rect 15208 943 15211 952
rect 15249 947 15250 968
rect 15257 965 15329 972
rect 15253 963 15329 965
rect 15257 956 15329 963
rect 15338 962 15339 968
rect 15332 956 15339 962
rect 15378 956 15384 962
rect 15433 956 15438 972
rect 15300 955 15341 956
rect 15326 950 15341 955
rect 15384 950 15390 956
rect 15215 942 15261 944
rect 15170 940 15180 942
rect 15261 940 15269 942
rect 15168 939 15170 940
rect 15269 939 15272 940
rect 14748 932 14750 933
rect 14721 927 14746 929
rect 14663 924 14665 925
rect 14486 914 14491 923
rect 14579 922 14609 924
rect 14659 922 14663 924
rect 14484 907 14486 914
rect 14452 895 14453 905
rect 14482 896 14484 907
rect 14555 906 14579 922
rect 14609 916 14659 922
rect 14744 915 14746 927
rect 14750 917 14758 929
rect 14795 926 14807 934
rect 14859 928 14865 934
rect 14981 926 14984 930
rect 15110 927 15168 939
rect 15211 938 15212 939
rect 15180 930 15192 938
rect 15202 930 15214 938
rect 15105 926 15110 927
rect 14864 922 14866 924
rect 14744 906 14747 915
rect 14783 910 14791 922
rect 14795 920 14813 922
rect 14481 891 14482 895
rect 14480 888 14481 891
rect 14542 886 14555 906
rect 14744 902 14746 906
rect 14729 897 14746 902
rect 14721 896 14746 897
rect 14720 895 14746 896
rect 14750 895 14758 907
rect 14669 886 14675 889
rect 14717 886 14746 895
rect 14749 892 14750 894
rect 14783 888 14791 900
rect 14795 890 14797 920
rect 14866 916 14873 922
rect 14873 914 14876 916
rect 14984 914 14998 926
rect 15091 923 15105 926
rect 15114 924 15123 927
rect 15212 926 15214 930
rect 15272 927 15319 939
rect 15332 935 15341 950
rect 15431 949 15433 956
rect 15449 952 15458 968
rect 15467 955 15476 972
rect 15539 968 15556 977
rect 15578 968 15617 978
rect 15430 946 15431 949
rect 15334 934 15335 935
rect 15384 933 15390 936
rect 15319 926 15324 927
rect 15332 926 15334 933
rect 15390 930 15397 933
rect 15407 930 15419 938
rect 15427 937 15429 942
rect 15449 937 15458 950
rect 15464 946 15467 955
rect 15509 954 15538 964
rect 15556 963 15617 968
rect 15556 957 15578 963
rect 15617 960 15627 963
rect 15502 945 15538 954
rect 15549 952 15558 954
rect 15461 937 15463 942
rect 15420 926 15427 937
rect 15449 934 15461 937
rect 15493 936 15502 945
rect 15509 944 15538 945
rect 15539 945 15558 952
rect 15578 950 15599 957
rect 15627 956 15637 960
rect 15657 956 15714 978
rect 15733 973 15739 979
rect 15744 977 15745 983
rect 15785 979 15791 985
rect 15745 972 15746 977
rect 15779 974 15785 979
rect 15786 974 15789 979
rect 15779 973 15786 974
rect 15785 972 15786 973
rect 15743 968 15746 972
rect 15794 971 15796 991
rect 15855 985 15861 991
rect 15866 988 15867 990
rect 15868 986 15871 987
rect 15871 985 15876 986
rect 15855 984 15911 985
rect 16060 984 16071 993
rect 16106 990 16118 994
rect 16132 993 16146 995
rect 16190 993 16196 999
rect 16334 998 16341 1000
rect 16343 998 16352 1018
rect 16427 1015 16440 1018
rect 17064 1015 17065 1026
rect 17254 1015 17255 1026
rect 17340 1015 17341 1026
rect 17613 1015 17614 1026
rect 17810 1015 17811 1026
rect 18046 1023 18085 1026
rect 19087 1023 19126 1028
rect 19312 1025 19318 1031
rect 19338 1026 19340 1035
rect 19341 1031 19342 1036
rect 19337 1024 19338 1026
rect 18043 1022 18046 1023
rect 18043 1015 18055 1022
rect 18060 1020 18063 1023
rect 18059 1016 18060 1019
rect 16440 1001 16504 1015
rect 16504 998 16514 1001
rect 16134 992 16144 993
rect 16181 992 16190 993
rect 16334 992 16352 998
rect 16395 992 16401 998
rect 16514 992 16559 998
rect 16654 994 16672 995
rect 16642 992 16654 994
rect 16106 986 16124 990
rect 16138 987 16144 992
rect 16184 987 16190 992
rect 16343 991 16349 992
rect 16343 989 16350 991
rect 16351 990 16352 992
rect 16381 991 16384 992
rect 16343 986 16349 989
rect 16351 987 16355 988
rect 16370 987 16381 991
rect 16386 986 16395 992
rect 16514 988 16642 992
rect 15855 983 15920 984
rect 16064 983 16072 984
rect 15872 981 15920 983
rect 15872 979 15884 981
rect 16066 978 16082 983
rect 16087 981 16088 984
rect 15914 972 15920 978
rect 15972 972 15978 978
rect 15743 967 15748 968
rect 15784 967 15785 971
rect 15734 958 15748 967
rect 15637 954 15642 956
rect 15714 955 15733 956
rect 15734 955 15746 958
rect 15642 951 15649 954
rect 15714 951 15746 955
rect 15748 951 15749 957
rect 15649 950 15651 951
rect 15539 944 15551 945
rect 15509 943 15516 944
rect 15558 943 15567 945
rect 15509 942 15514 943
rect 15509 941 15511 942
rect 15509 940 15555 941
rect 15556 940 15567 943
rect 15505 939 15510 940
rect 15517 939 15551 940
rect 15505 938 15551 939
rect 15505 937 15517 938
rect 15454 926 15461 934
rect 15504 931 15517 937
rect 15548 936 15551 938
rect 15555 937 15567 940
rect 15599 943 15669 950
rect 15714 949 15734 951
rect 15737 949 15751 950
rect 15727 948 15751 949
rect 15727 946 15734 948
rect 15737 945 15754 948
rect 15779 946 15784 967
rect 15796 951 15798 968
rect 15920 966 15926 972
rect 15929 967 15932 972
rect 15798 949 15803 950
rect 15599 942 15672 943
rect 15599 939 15669 942
rect 15672 939 15681 942
rect 15737 939 15751 945
rect 15754 943 15764 945
rect 15793 943 15803 949
rect 15932 948 15939 967
rect 15966 966 15978 972
rect 16071 968 16082 978
rect 16106 980 16125 986
rect 16106 973 16143 980
rect 16267 976 16283 984
rect 16345 982 16348 986
rect 16344 976 16345 981
rect 16088 968 16091 972
rect 15972 945 15978 966
rect 16082 953 16094 968
rect 16110 965 16143 973
rect 16227 968 16230 976
rect 16268 975 16283 976
rect 16343 970 16344 975
rect 16386 969 16389 986
rect 16398 972 16499 977
rect 16499 969 16510 972
rect 16541 969 16642 988
rect 16672 980 16694 994
rect 16088 951 16091 953
rect 16094 951 16096 953
rect 15669 937 15701 939
rect 15549 931 15551 936
rect 15562 931 15568 937
rect 15669 934 15733 937
rect 15737 934 15753 939
rect 15764 934 15828 943
rect 16096 942 16116 951
rect 16125 948 16143 965
rect 16223 957 16227 968
rect 16218 955 16223 957
rect 16180 950 16181 953
rect 15941 939 15948 942
rect 15965 939 16005 942
rect 15929 936 15965 939
rect 15912 934 15929 936
rect 15505 930 15517 931
rect 15082 921 15091 923
rect 15070 920 15082 921
rect 15109 920 15114 924
rect 15023 915 15109 920
rect 15011 914 15023 915
rect 15051 914 15070 915
rect 15168 914 15176 926
rect 15180 924 15214 926
rect 14876 913 15006 914
rect 14984 909 14998 913
rect 15040 911 15051 914
rect 15033 907 15039 911
rect 14923 900 14929 906
rect 14929 894 14935 900
rect 14957 892 14970 900
rect 15000 892 15011 907
rect 15025 900 15030 904
rect 15162 901 15171 913
rect 15180 901 15182 924
rect 14795 888 14813 890
rect 14957 889 14966 892
rect 14970 891 14972 892
rect 15012 889 15014 891
rect 15022 889 15031 898
rect 15171 892 15182 901
rect 15212 892 15214 924
rect 15218 914 15226 926
rect 15324 924 15334 926
rect 15391 924 15419 926
rect 15420 924 15431 926
rect 15324 923 15332 924
rect 15329 921 15332 923
rect 15384 921 15385 924
rect 15417 921 15431 924
rect 15250 907 15264 921
rect 15319 910 15329 921
rect 15383 917 15384 921
rect 15319 907 15332 910
rect 15382 907 15383 916
rect 15417 915 15419 921
rect 15420 915 15431 921
rect 15454 924 15462 926
rect 15454 915 15461 924
rect 15462 921 15466 924
rect 15465 918 15471 921
rect 15466 916 15471 918
rect 15417 911 15420 915
rect 15422 914 15431 915
rect 15422 912 15423 914
rect 15264 906 15319 907
rect 15326 904 15332 907
rect 15381 904 15382 906
rect 15384 904 15390 910
rect 15417 906 15419 911
rect 15423 907 15425 912
rect 15425 906 15426 907
rect 15416 904 15419 906
rect 15426 904 15427 906
rect 15332 898 15338 904
rect 15374 902 15377 904
rect 15378 902 15384 904
rect 15373 898 15384 902
rect 15415 901 15416 904
rect 15373 892 15380 898
rect 15414 897 15415 900
rect 15412 894 15414 895
rect 15417 894 15419 904
rect 15385 892 15419 894
rect 15423 901 15431 904
rect 15423 892 15437 901
rect 15412 891 15414 892
rect 15437 890 15440 892
rect 14538 879 14542 885
rect 14664 879 14717 886
rect 14727 883 14733 886
rect 14734 883 14746 886
rect 14801 884 14807 888
rect 14535 875 14538 879
rect 14634 875 14664 879
rect 14675 877 14681 879
rect 14480 871 14481 875
rect 14532 870 14535 874
rect 14596 870 14634 875
rect 14594 869 14596 870
rect 14531 868 14532 869
rect 14592 868 14594 869
rect 14683 868 14685 879
rect 14718 868 14719 879
rect 14721 877 14727 883
rect 14795 882 14807 884
rect 14859 882 14865 888
rect 14795 876 14813 882
rect 14853 876 14859 882
rect 14966 880 14975 889
rect 15012 888 15022 889
rect 15410 888 15412 889
rect 15013 887 15022 888
rect 15013 880 15033 887
rect 15215 885 15216 888
rect 15176 882 15177 884
rect 15385 880 15397 888
rect 15407 882 15419 888
rect 15440 884 15442 890
rect 15444 885 15454 915
rect 15471 912 15484 916
rect 15484 907 15496 912
rect 15499 906 15501 907
rect 15510 906 15517 930
rect 15562 928 15563 931
rect 15685 919 15733 934
rect 15753 932 15828 934
rect 15845 933 15896 934
rect 15898 933 15909 934
rect 15845 932 15906 933
rect 15753 930 15845 932
rect 15501 904 15506 906
rect 15510 904 15562 906
rect 15506 901 15562 904
rect 15510 899 15562 901
rect 15493 889 15502 898
rect 15510 896 15579 899
rect 15510 891 15567 896
rect 15579 892 15604 896
rect 15701 894 15709 919
rect 15733 916 15740 919
rect 15753 918 15769 930
rect 15771 918 15787 930
rect 15892 929 15907 932
rect 15888 927 15892 929
rect 15872 922 15888 927
rect 15898 926 15907 929
rect 15941 926 15948 936
rect 15901 920 15906 922
rect 15719 900 15723 916
rect 15740 914 15771 916
rect 15772 914 15774 918
rect 15740 909 15772 914
rect 15763 907 15780 909
rect 15763 902 15772 907
rect 15780 906 15784 907
rect 15723 896 15724 899
rect 15743 898 15763 902
rect 15504 889 15568 891
rect 15604 890 15616 892
rect 15700 890 15701 893
rect 15502 885 15568 889
rect 15406 880 15419 882
rect 14976 875 14979 880
rect 15020 879 15033 880
rect 14518 864 14531 868
rect 14586 864 14592 868
rect 14512 862 14518 864
rect 14583 862 14586 864
rect 14509 858 14512 862
rect 14576 857 14583 862
rect 14508 856 14509 857
rect 14575 856 14576 857
rect 14507 849 14508 856
rect 14572 849 14575 856
rect 14506 841 14507 849
rect 14574 838 14583 842
rect 14621 838 14630 842
rect 14633 838 14649 854
rect 14651 838 14667 854
rect 14685 838 14689 867
rect 14716 847 14718 867
rect 14979 860 14986 875
rect 15018 873 15033 875
rect 14729 849 14743 854
rect 14825 842 14829 856
rect 13040 804 13050 805
rect 14502 804 14506 838
rect 14571 833 14583 838
rect 14617 833 14633 838
rect 14667 837 14683 838
rect 14674 834 14683 837
rect 14565 832 14578 833
rect 14617 832 14639 833
rect 14563 831 14572 832
rect 14563 811 14565 831
rect 14566 826 14572 831
rect 14562 810 14565 811
rect 14563 804 14565 810
rect 14571 820 14572 826
rect 14604 824 14639 832
rect 14604 823 14633 824
rect 14604 822 14652 823
rect 14678 822 14683 834
rect 14604 820 14624 822
rect 14633 820 14652 822
rect 14571 804 14587 820
rect 14617 804 14633 820
rect 14677 812 14678 817
rect 12948 803 12949 804
rect 12947 801 12948 802
rect 12895 799 12938 801
rect 12730 796 12895 799
rect 12730 795 12836 796
rect 12919 795 12938 799
rect 12712 794 12746 795
rect 12694 792 12728 794
rect 12673 789 12702 792
rect 12588 785 12599 788
rect 12648 787 12673 789
rect 12635 786 12648 787
rect 12631 785 12635 786
rect 12490 784 12493 785
rect 12511 784 12599 785
rect 12511 783 12588 784
rect 12604 783 12631 785
rect 12659 784 12662 787
rect 12333 779 12334 780
rect 12371 769 12379 783
rect 12413 778 12414 783
rect 12489 781 12490 783
rect 12512 782 12514 783
rect 12488 778 12489 781
rect 12514 780 12517 782
rect 12522 781 12523 783
rect 12580 782 12604 783
rect 12569 779 12580 782
rect 12517 778 12520 779
rect 12069 756 12087 757
rect 12115 756 12121 758
rect 12063 750 12127 756
rect 12152 753 12182 766
rect 12212 763 12250 769
rect 12368 763 12371 769
rect 12212 759 12244 763
rect 12211 756 12212 758
rect 12152 750 12188 753
rect 12209 752 12211 756
rect 12213 755 12244 759
rect 12241 754 12243 755
rect 12244 754 12247 755
rect 12363 754 12368 763
rect 12240 752 12241 754
rect 12247 751 12252 754
rect 12362 752 12363 754
rect 11963 744 11969 750
rect 12069 745 12121 750
rect 11873 742 11917 744
rect 11722 741 11756 742
rect 11873 741 11879 742
rect 11685 740 11722 741
rect 11662 739 11685 740
rect 11659 737 11662 739
rect 11911 738 11917 742
rect 11969 738 11975 744
rect 11634 723 11659 737
rect 11750 730 11756 736
rect 11808 731 11814 736
rect 12063 733 12075 745
rect 12109 735 12114 745
rect 11839 731 11875 733
rect 11756 724 11762 730
rect 11780 729 11839 731
rect 11875 729 11881 731
rect 11778 726 11780 729
rect 11629 720 11634 723
rect 11527 717 11609 719
rect 11530 716 11609 717
rect 11626 716 11634 720
rect 11576 713 11584 716
rect 11588 715 11590 716
rect 11609 715 11638 716
rect 11588 713 11622 715
rect 11619 709 11622 713
rect 11626 713 11634 715
rect 11638 714 11666 715
rect 11626 711 11629 713
rect 11623 709 11626 711
rect 11666 710 11680 714
rect 11772 713 11778 726
rect 11802 724 11808 729
rect 11881 726 11892 729
rect 12069 726 12075 733
rect 11871 722 11873 723
rect 11892 722 11903 726
rect 12068 723 12075 726
rect 11903 721 11905 722
rect 11905 720 11909 721
rect 11253 707 11254 708
rect 11475 707 11476 708
rect 11588 701 11600 709
rect 11610 701 11622 709
rect 11680 705 11686 710
rect 11770 708 11772 713
rect 11769 707 11770 708
rect 11686 703 11697 705
rect 11314 697 11448 700
rect 11614 698 11618 701
rect 11697 699 11710 703
rect 11710 698 11715 699
rect 11190 695 11314 697
rect 11448 695 11454 697
rect 11093 692 11099 694
rect 11168 692 11190 695
rect 11454 692 11460 695
rect 10875 688 10876 690
rect 11089 688 11091 691
rect 11092 688 11093 690
rect 11145 689 11168 692
rect 11460 689 11466 692
rect 11598 690 11614 698
rect 11715 694 11731 698
rect 11731 692 11747 694
rect 11747 691 11756 692
rect 11762 691 11769 706
rect 11863 693 11871 698
rect 11875 693 11877 720
rect 12063 711 12075 723
rect 12114 711 12116 726
rect 12152 723 12182 750
rect 12208 749 12209 751
rect 12252 750 12254 751
rect 12192 746 12194 747
rect 12206 745 12208 749
rect 12195 737 12209 745
rect 12237 744 12239 749
rect 12257 747 12260 749
rect 12260 746 12262 747
rect 12262 743 12266 746
rect 12286 743 12298 749
rect 12357 744 12360 749
rect 12392 744 12413 778
rect 12479 756 12488 778
rect 12517 776 12522 778
rect 12523 776 12569 779
rect 12662 778 12663 781
rect 12517 775 12569 776
rect 12517 756 12522 775
rect 12663 772 12667 778
rect 12663 756 12670 772
rect 12694 756 12702 789
rect 12712 788 12728 792
rect 12730 788 12746 794
rect 12808 788 12824 795
rect 12922 788 12938 795
rect 12925 787 12926 788
rect 12926 783 12927 785
rect 12928 772 12931 779
rect 12951 778 12963 804
rect 13000 799 13001 802
rect 13000 796 13002 799
rect 13038 796 13040 800
rect 14506 799 14519 804
rect 14536 799 14571 804
rect 14519 797 14536 799
rect 13000 791 13008 796
rect 13035 791 13038 796
rect 13000 788 13016 791
rect 13018 788 13034 791
rect 14555 788 14572 799
rect 14633 797 14636 803
rect 14633 795 14637 797
rect 14633 788 14643 795
rect 14563 786 14572 788
rect 14637 786 14643 788
rect 14688 786 14689 828
rect 14713 822 14726 838
rect 14859 833 14863 838
rect 14881 837 14893 845
rect 14947 838 14963 854
rect 14986 842 14995 860
rect 14987 841 14995 842
rect 14999 845 15000 862
rect 14999 843 15003 845
rect 15031 844 15033 873
rect 15034 869 15045 875
rect 15037 863 15045 869
rect 15041 859 15044 863
rect 15177 860 15181 879
rect 15214 866 15215 880
rect 15296 867 15302 873
rect 15342 867 15348 873
rect 15406 870 15410 880
rect 15439 870 15444 884
rect 15502 880 15516 885
rect 15510 871 15516 880
rect 15552 880 15562 885
rect 15552 870 15553 880
rect 15556 879 15562 880
rect 15616 879 15683 890
rect 15699 885 15700 889
rect 15698 881 15699 885
rect 15684 875 15688 879
rect 15688 872 15691 875
rect 15695 871 15698 881
rect 15724 879 15728 896
rect 15738 891 15743 898
rect 15784 892 15841 906
rect 15841 891 15844 892
rect 15735 881 15737 889
rect 15844 888 15858 891
rect 15904 890 15906 920
rect 15910 910 15918 922
rect 15948 914 15953 926
rect 15953 902 15958 914
rect 15978 910 15985 939
rect 16005 936 16011 939
rect 16011 934 16015 936
rect 16092 935 16093 942
rect 16116 939 16122 942
rect 16122 936 16128 939
rect 16015 933 16016 934
rect 16016 927 16019 933
rect 16019 922 16022 927
rect 16022 919 16024 922
rect 16024 916 16025 919
rect 15875 888 15906 890
rect 15910 888 15918 900
rect 15958 899 15959 902
rect 15985 900 15987 910
rect 16025 902 16032 916
rect 16093 910 16097 935
rect 16128 934 16132 936
rect 16143 935 16144 942
rect 16130 933 16136 934
rect 16130 932 16138 933
rect 16144 932 16145 935
rect 16180 934 16195 950
rect 16218 948 16230 955
rect 16217 947 16230 948
rect 16240 947 16252 955
rect 16283 952 16299 968
rect 16214 945 16223 947
rect 16213 943 16214 945
rect 16217 943 16223 945
rect 16256 943 16257 945
rect 16263 943 16269 948
rect 16206 942 16213 943
rect 16217 942 16252 943
rect 16256 942 16269 943
rect 16206 937 16217 942
rect 16218 941 16252 942
rect 16204 934 16210 937
rect 16211 936 16217 937
rect 16251 936 16252 941
rect 16269 936 16275 942
rect 16283 934 16299 950
rect 16336 939 16343 968
rect 16389 956 16390 968
rect 16394 965 16395 969
rect 16510 968 16529 969
rect 16537 968 16541 969
rect 16501 964 16537 968
rect 16587 965 16591 969
rect 16335 934 16336 938
rect 16200 932 16204 934
rect 16138 931 16179 932
rect 16144 918 16161 931
rect 16163 926 16179 931
rect 16197 930 16200 932
rect 16190 926 16197 930
rect 16282 927 16283 931
rect 16334 927 16335 932
rect 16163 918 16190 926
rect 16281 920 16283 927
rect 16333 922 16334 927
rect 16344 922 16352 934
rect 16356 922 16358 956
rect 16394 951 16395 964
rect 16501 960 16549 964
rect 16492 954 16501 960
rect 16389 945 16390 951
rect 16395 936 16396 945
rect 16484 939 16492 954
rect 16530 949 16549 960
rect 16549 948 16551 949
rect 16591 948 16596 965
rect 16694 961 16697 980
rect 16697 954 16698 960
rect 16551 945 16555 948
rect 16596 945 16597 948
rect 16481 936 16484 939
rect 16396 928 16402 934
rect 16397 922 16402 928
rect 16476 928 16488 936
rect 16498 928 16510 936
rect 16555 934 16570 945
rect 16597 934 16601 945
rect 16698 941 16701 954
rect 16700 939 16701 941
rect 16698 934 16700 939
rect 16570 932 16571 934
rect 16571 928 16572 930
rect 16601 929 16603 934
rect 16476 924 16481 928
rect 16514 926 16515 928
rect 16516 924 16519 925
rect 16280 919 16283 920
rect 16144 905 16145 918
rect 16172 916 16190 918
rect 16279 918 16283 919
rect 16279 916 16280 918
rect 16332 916 16333 919
rect 16352 916 16353 921
rect 16166 912 16172 916
rect 16275 909 16279 916
rect 16331 909 16332 916
rect 16353 912 16355 916
rect 16383 913 16390 922
rect 16397 916 16398 922
rect 16376 911 16383 913
rect 16394 911 16398 916
rect 16464 912 16472 924
rect 16476 922 16510 924
rect 16476 921 16479 922
rect 16356 910 16394 911
rect 16145 902 16146 904
rect 16032 899 16034 902
rect 15987 894 15988 899
rect 16034 896 16035 899
rect 15858 885 15869 888
rect 15872 885 15911 888
rect 15869 884 15911 885
rect 15728 872 15730 879
rect 15730 870 15731 872
rect 15732 871 15735 881
rect 15872 879 15911 884
rect 15960 881 15962 889
rect 15894 876 15906 879
rect 15911 874 15933 879
rect 15962 874 15963 881
rect 15947 872 15952 874
rect 15381 868 15382 869
rect 15405 867 15406 870
rect 15290 861 15296 867
rect 15348 861 15354 867
rect 15403 860 15405 867
rect 15044 854 15048 858
rect 15044 853 15059 854
rect 15030 843 15033 844
rect 14999 841 15033 843
rect 15037 841 15045 853
rect 15048 850 15059 853
rect 15181 852 15182 858
rect 15215 854 15216 858
rect 15050 845 15059 850
rect 15053 840 15059 845
rect 14816 831 14893 833
rect 14716 820 14721 822
rect 14713 804 14726 820
rect 14716 787 14721 804
rect 14729 788 14745 799
rect 14565 780 14572 786
rect 14630 785 14643 786
rect 14630 783 14677 785
rect 14605 780 14652 783
rect 12474 745 12479 756
rect 12514 744 12517 756
rect 12667 750 12670 756
rect 12667 744 12674 750
rect 12702 744 12704 756
rect 12732 751 12744 759
rect 12754 751 12766 759
rect 12931 755 12936 772
rect 12963 770 12967 778
rect 14565 777 14578 780
rect 14618 777 14624 780
rect 14630 779 14652 780
rect 14630 777 14639 779
rect 14816 777 14874 831
rect 14891 799 14893 831
rect 14897 821 14905 833
rect 14963 822 14979 838
rect 15033 837 15037 840
rect 15057 838 15059 840
rect 15081 838 15087 844
rect 15127 839 15133 844
rect 15123 838 15135 839
rect 15182 838 15185 850
rect 15217 841 15233 854
rect 15288 852 15296 858
rect 15286 850 15296 852
rect 15400 851 15403 860
rect 15349 848 15359 850
rect 15359 846 15365 848
rect 15398 847 15400 851
rect 15276 845 15284 846
rect 15286 845 15290 846
rect 15216 840 15233 841
rect 15216 838 15220 840
rect 14999 829 15011 837
rect 15021 829 15033 837
rect 15059 832 15139 838
rect 15185 832 15186 837
rect 14999 828 15000 829
rect 15000 818 15002 828
rect 15059 822 15075 832
rect 15081 831 15135 832
rect 15081 827 15133 831
rect 15002 814 15004 818
rect 15004 809 15005 812
rect 15005 805 15006 809
rect 15006 799 15007 803
rect 15007 792 15009 799
rect 15081 793 15101 827
rect 15127 825 15135 827
rect 15133 794 15135 825
rect 15139 815 15147 827
rect 15127 793 15135 794
rect 15139 793 15147 805
rect 15163 804 15171 820
rect 15186 814 15189 829
rect 15201 822 15220 838
rect 15254 833 15263 842
rect 15276 841 15286 845
rect 15288 844 15290 845
rect 15365 844 15372 846
rect 15288 841 15296 844
rect 15372 843 15376 844
rect 15376 842 15381 843
rect 15397 842 15398 844
rect 15393 841 15404 842
rect 15429 841 15439 869
rect 15444 866 15445 869
rect 15445 854 15448 865
rect 15516 860 15521 870
rect 15692 869 15695 870
rect 15691 865 15695 869
rect 15692 860 15695 865
rect 15722 866 15732 870
rect 15952 866 15969 872
rect 15988 871 15992 890
rect 16035 888 16039 896
rect 16143 890 16146 896
rect 16152 891 16163 908
rect 16218 903 16230 909
rect 16330 908 16331 909
rect 16259 903 16275 908
rect 16329 903 16330 908
rect 16376 903 16383 910
rect 16230 902 16259 903
rect 16328 896 16329 899
rect 16211 890 16217 896
rect 16269 890 16275 896
rect 16039 874 16047 888
rect 16141 885 16143 889
rect 16149 886 16152 890
rect 15521 854 15522 860
rect 15691 854 15694 860
rect 15445 852 15451 854
rect 15448 846 15451 852
rect 15513 849 15529 854
rect 15512 848 15526 849
rect 15531 848 15547 854
rect 15449 841 15451 846
rect 15509 845 15512 848
rect 15526 845 15547 848
rect 15504 841 15509 845
rect 15537 842 15549 845
rect 15276 838 15290 841
rect 15396 839 15397 841
rect 15404 840 15439 841
rect 15450 840 15451 841
rect 15502 840 15504 841
rect 15429 839 15477 840
rect 15500 838 15502 840
rect 15516 839 15528 842
rect 15609 841 15625 854
rect 15627 841 15643 854
rect 15689 847 15691 853
rect 15692 852 15694 854
rect 15722 852 15740 866
rect 15963 863 15978 866
rect 15549 840 15550 841
rect 15602 840 15603 841
rect 15521 838 15528 839
rect 15270 834 15284 838
rect 15270 833 15281 834
rect 15245 824 15254 833
rect 15216 820 15220 822
rect 15201 814 15220 820
rect 15189 809 15190 812
rect 15190 799 15192 808
rect 15201 804 15217 814
rect 15276 812 15284 824
rect 15288 814 15290 838
rect 15393 832 15396 838
rect 15348 815 15354 821
rect 15382 818 15400 832
rect 15388 815 15389 818
rect 15342 814 15348 815
rect 15387 814 15388 815
rect 15288 812 15322 814
rect 15331 812 15390 814
rect 15400 813 15406 818
rect 15401 812 15407 813
rect 15220 808 15221 812
rect 15312 809 15322 812
rect 15326 810 15331 812
rect 15303 808 15312 809
rect 15315 808 15321 809
rect 15323 808 15326 810
rect 15342 809 15348 812
rect 15221 804 15222 808
rect 15288 805 15300 808
rect 15303 805 15322 808
rect 15288 804 15301 805
rect 15217 794 15225 804
rect 15248 800 15300 804
rect 15310 800 15322 805
rect 15378 800 15387 811
rect 15390 810 15398 812
rect 15401 810 15412 812
rect 15420 811 15429 838
rect 15451 822 15467 838
rect 15491 832 15499 838
rect 15398 809 15412 810
rect 15414 809 15420 810
rect 15398 808 15420 809
rect 15451 808 15467 820
rect 15520 811 15522 838
rect 15523 837 15528 838
rect 15525 836 15528 837
rect 15550 838 15551 840
rect 15601 838 15602 840
rect 15526 834 15530 836
rect 15531 832 15532 834
rect 15550 832 15563 838
rect 15524 828 15528 830
rect 15401 804 15467 808
rect 15410 800 15451 804
rect 15491 801 15492 804
rect 15217 793 15227 794
rect 15081 792 15133 793
rect 15217 792 15229 793
rect 15009 789 15015 792
rect 15015 784 15022 789
rect 15075 788 15155 792
rect 15193 790 15194 792
rect 15217 789 15238 792
rect 15217 788 15232 789
rect 15075 786 15139 788
rect 15227 786 15232 788
rect 15238 787 15243 789
rect 15243 786 15247 787
rect 15248 786 15299 800
rect 15311 793 15315 800
rect 15373 793 15378 799
rect 15310 790 15311 793
rect 15371 790 15373 793
rect 15022 783 15023 784
rect 15058 783 15059 785
rect 15024 779 15030 783
rect 15055 779 15058 783
rect 15081 780 15087 786
rect 15123 781 15135 786
rect 15243 785 15254 786
rect 15245 783 15254 785
rect 15245 782 15257 783
rect 15127 780 15133 781
rect 15193 779 15194 781
rect 15030 777 15035 779
rect 15054 777 15055 779
rect 12714 747 12720 750
rect 12768 749 12770 750
rect 12723 747 12727 749
rect 12714 746 12723 747
rect 12713 744 12721 746
rect 12732 745 12768 747
rect 12770 745 12778 747
rect 12235 738 12237 743
rect 12266 741 12298 743
rect 12294 740 12299 741
rect 12301 737 12304 739
rect 12354 738 12357 744
rect 12389 739 12392 744
rect 12472 740 12474 744
rect 12489 740 12501 742
rect 12202 734 12203 737
rect 12209 734 12213 737
rect 12201 732 12202 734
rect 12213 732 12217 734
rect 12233 732 12235 737
rect 12263 736 12264 737
rect 12293 734 12303 737
rect 12304 734 12310 737
rect 12316 734 12322 737
rect 12298 732 12303 734
rect 12198 725 12201 731
rect 12217 729 12221 732
rect 12231 729 12233 731
rect 12197 722 12198 724
rect 12193 711 12197 721
rect 12221 712 12249 729
rect 12262 726 12263 731
rect 12303 727 12307 732
rect 12309 731 12322 734
rect 12347 732 12351 734
rect 12345 731 12347 732
rect 12362 731 12368 737
rect 12452 734 12458 740
rect 12470 734 12471 736
rect 12489 734 12504 740
rect 12513 738 12514 742
rect 12662 738 12668 744
rect 12720 738 12726 744
rect 12732 743 12734 745
rect 12512 734 12513 737
rect 12385 732 12386 734
rect 12446 732 12510 734
rect 12307 726 12309 727
rect 12310 726 12316 731
rect 12064 710 12068 711
rect 12069 710 12121 711
rect 12063 706 12127 710
rect 12058 704 12127 706
rect 12190 704 12193 711
rect 11917 698 11923 699
rect 11931 698 11969 699
rect 11911 695 11923 698
rect 11927 695 11975 698
rect 11911 693 11917 695
rect 11927 693 11965 695
rect 11969 693 11975 695
rect 11863 692 11975 693
rect 11863 691 11957 692
rect 11466 688 11469 689
rect 11473 688 11475 690
rect 9409 674 9412 685
rect 8725 653 8726 655
rect 8868 654 8869 656
rect 7657 651 7659 652
rect 7524 649 7600 651
rect 7652 649 7657 651
rect 7892 649 7896 652
rect 7955 650 7957 652
rect 7945 649 7955 650
rect 7607 648 7651 649
rect 7903 640 7919 649
rect 7920 648 7921 649
rect 8185 647 8187 651
rect 8205 647 8317 652
rect 8199 644 8317 647
rect 8415 644 8564 652
rect 8199 640 8215 644
rect 8317 641 8328 644
rect 8368 641 8415 644
rect 8328 640 8368 641
rect 8505 640 8521 644
rect 5313 639 5314 640
rect 8567 636 8597 652
rect 8705 640 8721 653
rect 8868 644 8878 654
rect 9141 652 9154 660
rect 9209 656 9225 672
rect 9347 665 9356 674
rect 9409 667 9421 674
rect 10876 669 10886 688
rect 11087 682 11093 688
rect 11145 682 11151 688
rect 11469 686 11475 688
rect 11092 680 11105 682
rect 11092 676 11099 680
rect 11139 676 11145 682
rect 11473 677 11475 686
rect 11575 681 11598 690
rect 11756 689 11778 691
rect 11863 689 11953 691
rect 11575 679 11645 681
rect 9412 665 9421 667
rect 9349 656 9350 665
rect 9356 656 9365 665
rect 9403 656 9417 665
rect 10886 658 10896 669
rect 10888 656 10902 658
rect 10938 656 10954 672
rect 11092 668 11093 676
rect 11469 671 11475 677
rect 11527 678 11598 679
rect 11527 676 11591 678
rect 11645 676 11654 679
rect 11527 671 11533 676
rect 11092 656 11104 668
rect 11472 665 11481 671
rect 11521 665 11527 671
rect 11472 662 11475 665
rect 11556 662 11575 676
rect 11654 675 11658 676
rect 11658 672 11660 675
rect 11662 667 11663 669
rect 11472 658 11474 662
rect 11552 659 11556 662
rect 11663 660 11678 667
rect 11762 662 11768 689
rect 11778 686 11813 689
rect 11863 686 11947 689
rect 11963 686 11969 692
rect 12058 690 12063 704
rect 12069 699 12087 704
rect 12069 698 12075 699
rect 12115 698 12121 704
rect 12188 699 12190 704
rect 12116 696 12117 698
rect 12186 695 12188 698
rect 12222 695 12230 712
rect 12250 709 12253 711
rect 12258 709 12262 726
rect 12309 717 12319 726
rect 12368 725 12374 731
rect 12381 725 12385 732
rect 12446 730 12504 732
rect 12505 730 12510 732
rect 12511 730 12512 732
rect 12446 728 12502 730
rect 12379 722 12380 724
rect 12319 709 12321 717
rect 12373 711 12379 721
rect 12253 708 12255 709
rect 12252 707 12256 708
rect 12252 703 12258 707
rect 12264 705 12265 707
rect 12264 703 12281 705
rect 12183 694 12186 695
rect 12179 692 12183 694
rect 12177 691 12179 692
rect 11813 684 11832 686
rect 11871 684 11935 686
rect 11832 683 11840 684
rect 11840 681 11861 683
rect 11871 681 11930 684
rect 11861 679 11930 681
rect 12054 679 12058 689
rect 12117 686 12119 690
rect 12173 689 12177 691
rect 12169 688 12173 689
rect 12219 688 12222 695
rect 12255 690 12258 703
rect 12261 699 12263 700
rect 12264 696 12288 699
rect 12264 691 12276 696
rect 12288 693 12302 696
rect 12321 693 12323 706
rect 12368 702 12373 711
rect 12452 696 12467 728
rect 12499 726 12502 728
rect 12505 726 12513 730
rect 12499 724 12501 726
rect 12500 700 12501 724
rect 12502 718 12513 726
rect 12502 714 12506 718
rect 12502 710 12505 714
rect 12508 712 12510 718
rect 12764 715 12766 745
rect 12768 742 12778 745
rect 12938 743 12940 749
rect 12948 743 12954 749
rect 12967 746 12990 770
rect 14452 755 14453 775
rect 14481 772 14482 775
rect 14572 774 14611 777
rect 14618 774 14630 777
rect 14482 759 14490 772
rect 14574 768 14611 774
rect 14621 768 14630 774
rect 14687 768 14688 777
rect 14482 755 14493 759
rect 14453 749 14454 755
rect 14490 753 14493 755
rect 14491 750 14496 753
rect 12994 743 13000 749
rect 14465 747 14494 748
rect 14497 747 14498 749
rect 12942 742 12948 743
rect 12770 738 12778 742
rect 12770 735 12788 738
rect 12778 731 12788 735
rect 12940 731 12948 742
rect 12953 738 12954 742
rect 12986 739 12992 742
rect 12951 731 12953 738
rect 12987 737 12992 739
rect 13000 737 13006 743
rect 12738 714 12766 715
rect 12733 713 12766 714
rect 12770 713 12778 725
rect 12788 721 12794 731
rect 12940 721 12951 731
rect 12932 720 12951 721
rect 12932 712 12941 720
rect 12507 710 12508 711
rect 12505 707 12509 710
rect 12767 709 12770 711
rect 12741 708 12744 709
rect 12504 702 12509 707
rect 12729 706 12739 708
rect 12720 704 12729 706
rect 12499 696 12501 699
rect 12302 692 12368 693
rect 12308 691 12368 692
rect 12142 686 12169 688
rect 12218 686 12219 688
rect 12117 684 12149 686
rect 12107 683 12149 684
rect 12080 681 12149 683
rect 12062 679 12149 681
rect 12215 679 12218 684
rect 11871 678 11930 679
rect 11874 677 11909 678
rect 12035 677 12149 679
rect 11874 676 11906 677
rect 11908 676 11909 677
rect 11875 674 11887 676
rect 11889 675 11908 676
rect 12013 675 12035 677
rect 12041 676 12149 677
rect 12054 675 12058 676
rect 11889 671 11916 675
rect 11965 671 12013 675
rect 11889 670 11927 671
rect 11954 670 11997 671
rect 11889 664 11997 670
rect 11891 662 11901 664
rect 12054 662 12055 675
rect 12119 672 12121 675
rect 12212 673 12215 679
rect 11768 660 11769 662
rect 11550 658 11552 659
rect 11252 656 11254 657
rect 11472 656 11473 658
rect 11548 656 11550 658
rect 9176 652 9209 656
rect 9409 652 9412 656
rect 9156 651 9175 652
rect 8924 645 8925 651
rect 8879 640 8895 644
rect 8897 640 8913 644
rect 9193 640 9209 652
rect 9350 645 9360 652
rect 9404 646 9409 652
rect 9398 645 9404 646
rect 9360 644 9401 645
rect 9385 640 9401 644
rect 10904 640 10920 656
rect 10922 640 10938 656
rect 11105 653 11107 656
rect 11245 653 11251 656
rect 11474 653 11477 656
rect 11544 653 11548 656
rect 11107 651 11109 653
rect 11244 652 11245 653
rect 11542 652 11544 653
rect 11678 652 11790 660
rect 11882 658 11891 662
rect 12119 659 12122 672
rect 12251 666 12255 689
rect 12314 685 12368 691
rect 12452 688 12504 696
rect 12505 692 12509 702
rect 12662 693 12668 698
rect 12720 693 12726 698
rect 12662 692 12726 693
rect 12509 688 12511 690
rect 12310 679 12374 685
rect 12446 682 12511 688
rect 12668 686 12674 692
rect 12714 686 12720 692
rect 12732 690 12733 706
rect 12754 701 12766 709
rect 12945 707 12951 720
rect 12988 717 12992 737
rect 12944 706 12945 707
rect 12940 697 12944 706
rect 12992 697 12994 717
rect 13755 703 13777 722
rect 14447 713 14454 725
rect 14459 716 14460 747
rect 14488 745 14493 747
rect 14492 716 14493 745
rect 14494 738 14505 747
rect 14721 740 14725 777
rect 15030 776 15054 777
rect 15191 775 15193 779
rect 15245 777 15254 782
rect 15260 779 15263 781
rect 15263 777 15282 779
rect 15310 777 15319 786
rect 15341 782 15347 788
rect 15368 786 15371 790
rect 15387 782 15393 788
rect 15405 786 15414 800
rect 15417 788 15433 800
rect 15435 796 15471 800
rect 15492 798 15494 801
rect 15519 800 15520 810
rect 15526 798 15528 828
rect 15532 818 15540 830
rect 15549 822 15563 832
rect 15593 836 15601 838
rect 15655 837 15659 841
rect 15687 839 15689 847
rect 15722 838 15732 852
rect 15740 848 15743 852
rect 15870 842 15876 844
rect 15870 838 15884 842
rect 15916 838 15922 844
rect 15923 838 15939 854
rect 15963 838 15969 863
rect 15978 853 15981 863
rect 15981 846 15983 852
rect 15983 838 15986 845
rect 15593 822 15600 836
rect 15617 826 15629 832
rect 15614 825 15673 826
rect 15677 825 15687 838
rect 15614 823 15622 825
rect 15673 823 15687 825
rect 15694 823 15697 838
rect 15549 820 15552 822
rect 15613 821 15614 823
rect 15492 796 15528 798
rect 15532 796 15540 808
rect 15549 804 15563 820
rect 15605 816 15613 820
rect 15617 818 15624 820
rect 15605 808 15611 816
rect 15617 814 15618 818
rect 15677 816 15702 823
rect 15711 816 15722 837
rect 15743 822 15755 838
rect 15864 832 15870 838
rect 15868 830 15870 832
rect 15872 830 15905 838
rect 15922 832 15928 838
rect 15939 832 15955 838
rect 15969 832 15970 838
rect 15922 830 15955 832
rect 15986 830 15989 838
rect 15992 830 16004 870
rect 16047 863 16052 874
rect 16094 871 16097 885
rect 16131 881 16141 885
rect 16217 884 16223 890
rect 16227 887 16228 890
rect 16237 886 16244 890
rect 16228 883 16231 885
rect 16234 884 16236 885
rect 16263 884 16269 890
rect 16326 888 16328 896
rect 16228 882 16233 883
rect 16129 874 16147 881
rect 16112 870 16129 874
rect 16131 870 16141 874
rect 16052 859 16054 863
rect 16078 838 16094 870
rect 16112 866 16131 870
rect 16110 863 16112 866
rect 16108 859 16110 863
rect 16124 859 16131 866
rect 16106 856 16108 859
rect 16104 854 16106 856
rect 16097 851 16106 854
rect 16097 845 16104 851
rect 16097 839 16101 845
rect 16097 838 16098 839
rect 16054 830 16055 838
rect 16078 830 16097 838
rect 16111 830 16124 859
rect 16141 846 16148 858
rect 16153 848 16154 880
rect 16220 876 16226 879
rect 16217 874 16220 876
rect 16208 869 16217 874
rect 16228 870 16231 882
rect 16265 870 16268 884
rect 16325 881 16326 888
rect 16324 874 16325 881
rect 16201 860 16202 863
rect 16231 860 16233 870
rect 16265 862 16279 870
rect 16321 863 16324 874
rect 16196 848 16201 860
rect 16153 847 16158 848
rect 16153 846 16187 847
rect 16194 846 16199 848
rect 16148 844 16149 846
rect 16193 844 16194 846
rect 16190 842 16192 843
rect 16153 834 16165 841
rect 16175 834 16187 841
rect 16233 830 16244 859
rect 16268 830 16279 862
rect 16320 856 16321 859
rect 16358 856 16376 903
rect 16464 890 16472 902
rect 16476 890 16478 921
rect 16509 920 16510 922
rect 16516 912 16522 924
rect 16572 913 16574 925
rect 16603 924 16619 928
rect 16689 925 16698 934
rect 16681 924 16689 925
rect 16603 913 16681 924
rect 16516 911 16519 912
rect 16519 903 16524 910
rect 16557 905 16619 913
rect 16551 903 16557 905
rect 16510 890 16551 903
rect 16519 888 16524 890
rect 16574 889 16576 905
rect 16472 886 16475 888
rect 16524 886 16525 888
rect 16576 885 16577 888
rect 16475 884 16477 885
rect 16476 883 16478 884
rect 16476 879 16479 883
rect 16525 880 16526 882
rect 16476 878 16480 879
rect 16479 876 16480 878
rect 16526 876 16527 880
rect 16577 876 16578 879
rect 16603 878 16619 905
rect 16480 869 16483 874
rect 16483 863 16485 869
rect 16418 861 16419 862
rect 16485 860 16486 863
rect 16297 851 16313 854
rect 16317 851 16320 856
rect 16356 851 16358 856
rect 16399 854 16411 855
rect 16297 845 16317 851
rect 16354 846 16356 851
rect 16393 847 16411 854
rect 16421 849 16433 855
rect 16421 847 16470 849
rect 16486 848 16490 860
rect 16393 845 16409 847
rect 16422 846 16470 847
rect 16415 845 16422 846
rect 16442 845 16470 846
rect 16297 843 16303 845
rect 16353 843 16354 845
rect 16393 843 16415 845
rect 16470 843 16484 845
rect 16490 844 16491 847
rect 16507 843 16523 854
rect 16295 839 16298 843
rect 16351 839 16353 843
rect 16387 842 16392 843
rect 16387 840 16391 842
rect 16393 841 16433 843
rect 16380 839 16390 840
rect 16393 839 16399 841
rect 16374 838 16379 839
rect 16393 838 16394 839
rect 16281 830 16295 838
rect 16348 836 16351 838
rect 16370 837 16374 838
rect 16361 836 16367 837
rect 16348 834 16361 836
rect 16338 833 16342 834
rect 16332 832 16338 833
rect 16319 830 16332 832
rect 16348 831 16351 834
rect 15860 827 15868 830
rect 15872 828 15875 830
rect 15859 821 15869 827
rect 15548 802 15549 804
rect 15550 800 15552 804
rect 15677 801 15687 816
rect 15689 812 15697 816
rect 15689 804 15698 812
rect 15702 807 15734 816
rect 15743 807 15755 820
rect 15835 807 15859 821
rect 15860 818 15868 821
rect 15698 801 15699 803
rect 15711 801 15722 807
rect 15734 804 15755 807
rect 15435 788 15451 796
rect 15471 795 15476 796
rect 15476 793 15487 795
rect 15494 794 15501 796
rect 15501 793 15507 794
rect 15518 793 15519 796
rect 15487 792 15492 793
rect 15507 792 15527 793
rect 15530 792 15532 795
rect 15547 794 15548 796
rect 15507 786 15528 792
rect 15544 789 15547 793
rect 15529 788 15547 789
rect 15529 786 15544 788
rect 15600 786 15601 788
rect 15605 786 15611 798
rect 15659 789 15660 801
rect 15674 790 15677 800
rect 15699 797 15727 801
rect 15734 797 15753 804
rect 15823 800 15835 807
rect 15821 799 15823 800
rect 15699 796 15753 797
rect 15814 796 15821 799
rect 15860 796 15868 808
rect 15872 796 15874 828
rect 15940 822 16169 830
rect 15940 820 15942 822
rect 15943 820 16169 822
rect 15940 814 16169 820
rect 16197 814 16319 830
rect 16342 818 16348 831
rect 16377 822 16393 838
rect 16340 815 16347 818
rect 15940 812 16197 814
rect 15942 804 15955 812
rect 15972 807 15974 812
rect 15942 803 15943 804
rect 15943 801 15944 802
rect 15940 796 15943 801
rect 15973 800 15974 807
rect 15985 804 15997 812
rect 15997 803 15998 804
rect 16002 803 16004 808
rect 16021 803 16100 812
rect 15998 802 16100 803
rect 16001 799 16017 802
rect 15618 787 15619 788
rect 15617 786 15623 787
rect 15399 782 15405 786
rect 15516 784 15528 786
rect 15190 772 15191 774
rect 15254 772 15282 777
rect 15183 759 15190 772
rect 15254 768 15263 772
rect 15301 768 15310 777
rect 15335 776 15341 782
rect 15393 776 15405 782
rect 15517 776 15518 781
rect 15393 766 15397 773
rect 15549 772 15550 786
rect 15601 783 15602 786
rect 15612 784 15614 785
rect 15658 784 15659 788
rect 15673 787 15674 790
rect 15699 789 15743 796
rect 15753 795 15755 796
rect 15755 792 15762 795
rect 15812 793 15814 796
rect 15911 795 15939 796
rect 15762 789 15766 792
rect 15699 788 15721 789
rect 15723 788 15739 789
rect 15766 788 15768 789
rect 15808 788 15812 793
rect 15923 792 15939 795
rect 15969 793 15973 799
rect 15680 787 15687 788
rect 15695 787 15709 788
rect 15768 787 15771 788
rect 15672 786 15680 787
rect 15667 785 15680 786
rect 15699 785 15709 787
rect 15864 786 15870 792
rect 15922 791 15939 792
rect 15966 791 15969 793
rect 15922 789 15978 791
rect 15999 789 16017 799
rect 15922 788 15939 789
rect 15966 788 15969 789
rect 15978 788 16017 789
rect 16019 788 16100 802
rect 16111 800 16124 812
rect 16187 804 16188 807
rect 15922 786 15928 788
rect 15965 786 15966 788
rect 15664 784 15673 785
rect 15602 780 15614 783
rect 15617 780 15618 781
rect 15626 780 15664 784
rect 15602 779 15661 780
rect 15617 774 15629 779
rect 15548 763 15550 772
rect 15667 763 15673 784
rect 15699 784 15713 785
rect 15173 756 15190 759
rect 15514 756 15517 763
rect 15173 755 15183 756
rect 15173 754 15180 755
rect 15513 754 15514 756
rect 15173 753 15177 754
rect 15162 749 15204 753
rect 15162 748 15189 749
rect 15160 747 15162 748
rect 15204 747 15207 749
rect 15146 745 15160 747
rect 14678 738 14684 740
rect 14721 739 14730 740
rect 14498 735 14516 738
rect 14505 725 14516 735
rect 14678 734 14690 738
rect 14724 734 14730 739
rect 15113 738 15146 745
rect 15107 737 15112 738
rect 14672 728 14678 734
rect 14730 729 14736 734
rect 15084 733 15107 737
rect 15161 735 15169 747
rect 15173 746 15178 747
rect 15078 731 15084 733
rect 15072 729 15074 731
rect 14694 728 14825 729
rect 14678 726 14694 728
rect 14730 727 15033 728
rect 15060 727 15066 729
rect 15071 728 15072 729
rect 14825 726 14826 727
rect 15033 726 15066 727
rect 15069 726 15071 728
rect 14459 714 14463 716
rect 14490 714 14493 716
rect 14459 713 14493 714
rect 14498 713 14516 725
rect 14666 714 14674 726
rect 14678 724 14684 726
rect 14454 711 14455 713
rect 14455 708 14460 711
rect 14493 708 14498 711
rect 14459 707 14471 708
rect 13726 697 13749 698
rect 13754 697 13777 703
rect 14458 701 14471 707
rect 14481 701 14493 708
rect 14505 707 14516 713
rect 12940 693 12948 697
rect 13000 693 13006 697
rect 14458 694 14460 701
rect 12940 691 13006 693
rect 12940 690 12944 691
rect 12733 686 12735 690
rect 12314 673 12322 679
rect 12362 673 12368 679
rect 12452 676 12458 682
rect 12498 676 12504 682
rect 12314 666 12321 673
rect 12454 672 12457 676
rect 11878 656 11882 658
rect 12055 656 12056 658
rect 12120 657 12122 659
rect 12118 656 12122 657
rect 11873 653 11878 656
rect 12056 653 12059 656
rect 12117 653 12118 656
rect 12152 654 12182 663
rect 12186 654 12199 660
rect 12251 659 12253 666
rect 12314 665 12322 666
rect 11868 652 11869 653
rect 12116 652 12117 653
rect 12149 652 12186 654
rect 12253 653 12255 659
rect 12311 656 12322 665
rect 12448 660 12457 672
rect 12510 672 12511 682
rect 12448 656 12454 660
rect 12510 656 12514 672
rect 12726 660 12735 686
rect 12934 674 12940 690
rect 12948 685 12954 691
rect 12994 685 13000 691
rect 14516 690 14523 707
rect 14666 692 14674 704
rect 14678 694 14680 724
rect 14827 719 14831 726
rect 15033 723 15068 726
rect 15106 723 15112 729
rect 14831 708 14838 719
rect 15054 717 15060 723
rect 15061 719 15068 723
rect 15112 719 15118 723
rect 15161 719 15169 725
rect 15173 719 15175 746
rect 15502 744 15508 750
rect 15510 744 15513 754
rect 15548 750 15549 763
rect 15654 757 15660 762
rect 15666 757 15667 762
rect 15699 758 15709 784
rect 15713 783 15717 784
rect 15772 783 15778 786
rect 15807 783 15808 786
rect 15870 784 15884 786
rect 15870 783 15876 784
rect 15908 783 15912 784
rect 15779 781 15781 782
rect 15781 780 15784 781
rect 15797 780 15807 783
rect 15726 775 15732 779
rect 15732 772 15737 775
rect 15784 772 15807 780
rect 15738 766 15762 772
rect 15797 769 15829 772
rect 15835 769 15908 783
rect 15916 780 15922 786
rect 15923 784 15924 785
rect 15964 784 15965 786
rect 15999 783 16002 788
rect 16008 787 16100 788
rect 16072 786 16100 787
rect 16049 785 16100 786
rect 16108 785 16111 799
rect 16186 797 16187 801
rect 16233 800 16244 814
rect 16268 804 16279 814
rect 16281 804 16297 814
rect 16334 807 16347 815
rect 16331 805 16347 807
rect 16377 805 16393 820
rect 16431 811 16433 841
rect 16437 831 16445 843
rect 16484 838 16524 843
rect 16527 842 16534 874
rect 16569 840 16577 852
rect 16581 842 16583 874
rect 16613 857 16618 874
rect 16613 842 16615 857
rect 16618 852 16619 856
rect 16581 840 16615 842
rect 16619 840 16627 852
rect 16534 838 16535 840
rect 16621 838 16623 840
rect 16524 837 16539 838
rect 16581 837 16582 838
rect 16533 836 16539 837
rect 16578 836 16580 837
rect 16415 809 16433 811
rect 16437 809 16445 821
rect 16494 805 16504 836
rect 16533 832 16548 836
rect 16536 808 16548 832
rect 16581 828 16593 836
rect 16603 828 16615 836
rect 16621 828 16635 838
rect 16582 820 16584 828
rect 16535 807 16548 808
rect 16320 804 16433 805
rect 16297 803 16433 804
rect 16185 791 16186 796
rect 16184 788 16185 791
rect 16244 789 16247 799
rect 16279 794 16287 800
rect 16297 795 16313 803
rect 16315 799 16433 803
rect 16504 801 16508 805
rect 16534 804 16548 807
rect 16569 815 16584 820
rect 16623 822 16635 828
rect 16623 820 16625 822
rect 16569 804 16585 815
rect 16623 805 16635 820
rect 17075 819 17076 1015
rect 17265 819 17266 1015
rect 17351 819 17352 1015
rect 17624 819 17625 1015
rect 17821 819 17822 1015
rect 18043 1013 18059 1015
rect 18065 1013 18077 1022
rect 18085 1020 18114 1023
rect 18114 1014 18118 1020
rect 18854 1018 18906 1020
rect 19126 1018 19140 1023
rect 19336 1020 19337 1023
rect 18826 1016 18906 1018
rect 18826 1015 18877 1016
rect 18118 1013 18119 1014
rect 18801 1013 18826 1015
rect 18848 1014 18854 1015
rect 18877 1014 18882 1015
rect 18039 1011 18043 1013
rect 18055 1010 18059 1013
rect 18767 1011 18797 1013
rect 18843 1012 18848 1014
rect 18031 998 18039 1010
rect 18038 988 18039 998
rect 18043 1007 18077 1010
rect 18043 1003 18045 1007
rect 18043 996 18044 1003
rect 18055 1001 18059 1007
rect 18074 1005 18077 1007
rect 18080 1004 18089 1010
rect 18042 994 18044 996
rect 18041 988 18047 994
rect 18052 988 18055 1001
rect 18035 982 18041 988
rect 18038 977 18039 982
rect 18042 977 18043 988
rect 18075 982 18077 1004
rect 18081 998 18089 1004
rect 18119 1001 18128 1010
rect 18650 1005 18664 1007
rect 18676 1005 18767 1011
rect 18839 1007 18843 1012
rect 18650 1004 18676 1005
rect 18650 1003 18664 1004
rect 18644 1002 18664 1003
rect 18685 1002 18690 1005
rect 18835 1002 18839 1007
rect 18882 1005 18899 1014
rect 18899 1004 18901 1005
rect 18087 988 18093 994
rect 18110 992 18119 1001
rect 18635 997 18659 1002
rect 18690 997 18696 1002
rect 18834 1001 18835 1002
rect 18906 1001 18923 1016
rect 19140 1015 19147 1018
rect 19335 1016 19336 1020
rect 19147 1014 19150 1015
rect 19150 1005 19172 1014
rect 19333 1012 19335 1016
rect 19373 1014 19377 1036
rect 19379 1027 19387 1039
rect 19645 1037 19657 1045
rect 19706 1041 19716 1045
rect 19717 1041 19723 1045
rect 19681 1037 19723 1041
rect 19775 1039 19781 1045
rect 19928 1044 19934 1050
rect 19974 1048 19984 1050
rect 19937 1044 19949 1048
rect 19959 1044 19971 1048
rect 19974 1044 19980 1048
rect 19922 1038 19928 1044
rect 19980 1038 19986 1044
rect 19426 1020 19436 1036
rect 19457 1034 19469 1037
rect 19651 1036 19657 1037
rect 19703 1036 19706 1037
rect 19451 1033 19471 1034
rect 19645 1033 19651 1036
rect 19687 1033 19717 1036
rect 19451 1031 19457 1033
rect 19471 1031 19501 1033
rect 19448 1025 19451 1031
rect 19445 1022 19451 1025
rect 19503 1024 19524 1031
rect 19551 1024 19557 1030
rect 19172 1004 19175 1005
rect 19032 1001 19033 1004
rect 18093 982 18099 988
rect 18110 986 18114 992
rect 18622 989 18635 997
rect 18644 993 18659 997
rect 18042 976 18044 977
rect 18042 962 18043 976
rect 18108 974 18109 979
rect 18266 976 18282 984
rect 18449 976 18465 989
rect 18532 979 18549 989
rect 18608 981 18622 989
rect 18602 979 18608 981
rect 18549 978 18602 979
rect 18633 977 18641 989
rect 18645 987 18650 989
rect 18696 987 18709 997
rect 18266 974 18323 976
rect 18104 957 18108 972
rect 18266 968 18311 974
rect 18323 968 18327 974
rect 18042 944 18049 957
rect 18103 953 18104 956
rect 18102 949 18103 952
rect 18105 944 18119 953
rect 18250 952 18266 968
rect 18327 961 18332 968
rect 18514 952 18520 958
rect 18560 952 18566 958
rect 18633 956 18641 967
rect 18645 958 18647 987
rect 18895 984 18897 1001
rect 18901 999 18923 1001
rect 18901 989 18909 999
rect 19027 992 19032 1001
rect 19175 996 19196 1004
rect 19330 1002 19333 1011
rect 19373 1007 19375 1014
rect 19364 1005 19375 1007
rect 19379 1010 19387 1017
rect 19379 1005 19392 1010
rect 19377 1004 19378 1005
rect 19378 1001 19379 1002
rect 19383 1001 19392 1005
rect 19426 1002 19436 1018
rect 19445 1015 19448 1022
rect 19499 1018 19505 1024
rect 19557 1018 19563 1024
rect 19633 1021 19641 1033
rect 19645 1031 19679 1033
rect 19645 1030 19651 1031
rect 19645 1029 19648 1030
rect 19445 1014 19447 1015
rect 19445 1013 19449 1014
rect 19447 1001 19449 1013
rect 19085 995 19118 996
rect 19196 995 19198 996
rect 19120 993 19126 995
rect 19027 986 19033 992
rect 19085 987 19091 992
rect 19126 991 19130 993
rect 19198 991 19208 995
rect 19328 991 19330 999
rect 19370 993 19383 1001
rect 19445 998 19449 1001
rect 19633 999 19641 1011
rect 19645 1002 19647 1029
rect 19925 1024 19928 1036
rect 19980 1032 19983 1036
rect 19933 1018 19937 1032
rect 19980 1021 19996 1032
rect 19996 1018 20012 1021
rect 19722 1007 19723 1008
rect 19723 1005 19724 1006
rect 19645 1001 19648 1002
rect 19691 1001 19719 1002
rect 19645 999 19657 1001
rect 19691 1000 19717 1001
rect 19375 992 19383 993
rect 19436 991 19440 996
rect 19445 991 19450 998
rect 19645 995 19649 999
rect 19691 998 19713 1000
rect 19719 999 19723 1001
rect 19691 996 19706 998
rect 19645 993 19651 995
rect 19691 994 19707 996
rect 19717 995 19723 999
rect 19726 997 19731 1003
rect 19775 1001 19784 1010
rect 19910 1001 19919 1010
rect 19919 1000 19925 1001
rect 18754 981 18770 984
rect 18772 981 18788 984
rect 18748 978 18768 981
rect 18889 979 18901 984
rect 19025 979 19026 983
rect 19033 980 19039 986
rect 19043 983 19111 987
rect 19130 986 19142 991
rect 18792 974 18793 978
rect 18750 972 18842 974
rect 18889 972 18909 979
rect 19024 974 19025 979
rect 19043 977 19069 983
rect 19079 980 19085 983
rect 19111 977 19124 983
rect 19142 978 19163 986
rect 19208 978 19242 991
rect 19374 988 19375 990
rect 19312 979 19318 985
rect 19328 983 19329 987
rect 19371 985 19374 986
rect 19023 972 19024 974
rect 19061 972 19069 977
rect 18654 963 18750 972
rect 18792 969 18793 972
rect 18751 963 18763 965
rect 18654 960 18751 963
rect 18645 957 18649 958
rect 18654 957 18750 960
rect 18645 956 18654 957
rect 18628 955 18652 956
rect 18656 955 18679 956
rect 18628 953 18647 955
rect 18696 954 18711 957
rect 18621 952 18628 953
rect 18641 952 18642 953
rect 18257 944 18266 952
rect 18508 946 18514 952
rect 18566 946 18572 952
rect 18602 949 18621 952
rect 18689 951 18696 954
rect 18645 950 18656 951
rect 18687 950 18689 951
rect 18580 946 18602 949
rect 18572 945 18594 946
rect 18035 936 18041 942
rect 18049 939 18061 944
rect 18097 942 18105 944
rect 18093 939 18105 942
rect 18255 939 18257 944
rect 18645 943 18657 950
rect 18260 940 18266 941
rect 18260 939 18302 940
rect 18306 939 18312 941
rect 18041 930 18047 936
rect 18061 934 18074 939
rect 18089 936 18099 939
rect 18087 934 18097 936
rect 18253 935 18255 939
rect 18260 936 18271 939
rect 18260 935 18266 936
rect 18302 935 18312 939
rect 18253 934 18260 935
rect 18080 929 18083 934
rect 18087 930 18093 934
rect 18078 926 18080 929
rect 18076 923 18078 926
rect 18250 925 18253 934
rect 18254 929 18260 934
rect 18312 929 18318 935
rect 18319 933 18331 941
rect 18392 934 18398 940
rect 18438 934 18444 940
rect 18708 939 18709 954
rect 18738 952 18748 957
rect 18747 939 18748 952
rect 18793 952 18804 968
rect 18765 942 18773 944
rect 18793 943 18796 952
rect 18834 947 18835 968
rect 18842 965 18914 972
rect 18838 963 18914 965
rect 18842 956 18914 963
rect 18923 962 18924 968
rect 18917 956 18924 962
rect 18963 956 18969 962
rect 19018 956 19023 972
rect 18885 955 18926 956
rect 18911 950 18926 955
rect 18969 950 18975 956
rect 18800 942 18846 944
rect 18755 940 18765 942
rect 18846 940 18854 942
rect 18753 939 18755 940
rect 18854 939 18857 940
rect 18333 932 18335 933
rect 18306 927 18331 929
rect 18248 924 18250 925
rect 18071 914 18076 923
rect 18164 922 18194 924
rect 18244 922 18248 924
rect 18069 907 18071 914
rect 18037 895 18038 905
rect 18067 896 18069 907
rect 18140 906 18164 922
rect 18194 916 18244 922
rect 18329 915 18331 927
rect 18335 917 18343 929
rect 18380 926 18392 934
rect 18444 928 18450 934
rect 18566 926 18569 930
rect 18695 927 18753 939
rect 18796 938 18797 939
rect 18765 930 18777 938
rect 18787 930 18799 938
rect 18690 926 18695 927
rect 18449 922 18451 924
rect 18329 906 18332 915
rect 18368 910 18376 922
rect 18380 920 18398 922
rect 18066 891 18067 895
rect 18065 888 18066 891
rect 18127 886 18140 906
rect 18329 902 18331 906
rect 18314 897 18331 902
rect 18306 896 18331 897
rect 18305 895 18331 896
rect 18335 895 18343 907
rect 18254 886 18260 889
rect 18302 886 18331 895
rect 18334 892 18335 894
rect 18368 888 18376 900
rect 18380 890 18382 920
rect 18451 916 18458 922
rect 18458 914 18461 916
rect 18569 914 18583 926
rect 18676 923 18690 926
rect 18699 924 18708 927
rect 18797 926 18799 930
rect 18857 927 18904 939
rect 18917 935 18926 950
rect 19016 949 19018 956
rect 19034 952 19043 968
rect 19052 955 19061 972
rect 19124 968 19141 977
rect 19163 968 19202 978
rect 19015 946 19016 949
rect 18919 934 18920 935
rect 18969 933 18975 936
rect 18904 926 18909 927
rect 18917 926 18919 933
rect 18975 930 18982 933
rect 18992 930 19004 938
rect 19012 937 19014 942
rect 19034 937 19043 950
rect 19049 946 19052 955
rect 19094 954 19123 964
rect 19141 963 19202 968
rect 19141 957 19163 963
rect 19202 960 19212 963
rect 19087 945 19123 954
rect 19134 952 19143 954
rect 19046 937 19048 942
rect 19005 926 19012 937
rect 19034 934 19046 937
rect 19078 936 19087 945
rect 19094 944 19123 945
rect 19124 945 19143 952
rect 19163 950 19184 957
rect 19212 956 19222 960
rect 19242 956 19299 978
rect 19318 973 19324 979
rect 19329 977 19330 983
rect 19370 979 19376 985
rect 19330 972 19331 977
rect 19364 974 19370 979
rect 19371 974 19374 979
rect 19364 973 19371 974
rect 19370 972 19371 973
rect 19328 968 19331 972
rect 19379 971 19381 991
rect 19440 985 19446 991
rect 19451 988 19452 990
rect 19453 986 19456 987
rect 19456 985 19461 986
rect 19440 984 19496 985
rect 19645 984 19656 993
rect 19691 990 19703 994
rect 19717 993 19731 995
rect 19775 993 19781 999
rect 19919 998 19926 1000
rect 19928 998 19937 1018
rect 20012 1015 20025 1018
rect 20649 1015 20650 1026
rect 20839 1015 20840 1026
rect 20925 1015 20926 1026
rect 21198 1015 21199 1026
rect 21395 1015 21396 1026
rect 20025 1001 20089 1015
rect 20089 998 20099 1001
rect 19719 992 19729 993
rect 19766 992 19775 993
rect 19919 992 19937 998
rect 19980 992 19986 998
rect 20099 992 20144 998
rect 20239 994 20257 995
rect 20227 992 20239 994
rect 19691 986 19709 990
rect 19723 987 19729 992
rect 19769 987 19775 992
rect 19928 991 19934 992
rect 19928 989 19935 991
rect 19936 990 19937 992
rect 19966 991 19969 992
rect 19928 986 19934 989
rect 19936 987 19940 988
rect 19955 987 19966 991
rect 19971 986 19980 992
rect 20099 988 20227 992
rect 19440 983 19505 984
rect 19649 983 19657 984
rect 19457 981 19505 983
rect 19457 979 19469 981
rect 19651 978 19667 983
rect 19672 981 19673 984
rect 19499 972 19505 978
rect 19557 972 19563 978
rect 19328 967 19333 968
rect 19369 967 19370 971
rect 19319 958 19333 967
rect 19222 954 19227 956
rect 19299 955 19318 956
rect 19319 955 19331 958
rect 19227 951 19234 954
rect 19299 951 19331 955
rect 19333 951 19334 957
rect 19234 950 19236 951
rect 19124 944 19136 945
rect 19094 943 19101 944
rect 19143 943 19152 945
rect 19094 942 19099 943
rect 19094 941 19096 942
rect 19094 940 19140 941
rect 19141 940 19152 943
rect 19090 939 19095 940
rect 19102 939 19136 940
rect 19090 938 19136 939
rect 19090 937 19102 938
rect 19039 926 19046 934
rect 19089 931 19102 937
rect 19133 936 19136 938
rect 19140 937 19152 940
rect 19184 943 19254 950
rect 19299 949 19319 951
rect 19322 949 19336 950
rect 19312 948 19336 949
rect 19312 946 19319 948
rect 19322 945 19339 948
rect 19364 946 19369 967
rect 19381 951 19383 968
rect 19505 966 19511 972
rect 19514 967 19517 972
rect 19383 949 19388 950
rect 19184 942 19257 943
rect 19184 939 19254 942
rect 19257 939 19266 942
rect 19322 939 19336 945
rect 19339 943 19349 945
rect 19378 943 19388 949
rect 19517 948 19524 967
rect 19551 966 19563 972
rect 19656 968 19667 978
rect 19691 980 19710 986
rect 19691 973 19728 980
rect 19852 976 19868 984
rect 19930 982 19933 986
rect 19929 976 19930 981
rect 19673 968 19676 972
rect 19557 945 19563 966
rect 19667 953 19679 968
rect 19695 965 19728 973
rect 19812 968 19815 976
rect 19853 975 19868 976
rect 19928 970 19929 975
rect 19971 969 19974 986
rect 19983 972 20084 977
rect 20084 969 20095 972
rect 20126 969 20227 988
rect 20257 980 20279 994
rect 19673 951 19676 953
rect 19679 951 19681 953
rect 19254 937 19286 939
rect 19134 931 19136 936
rect 19147 931 19153 937
rect 19254 934 19318 937
rect 19322 934 19338 939
rect 19349 934 19413 943
rect 19681 942 19701 951
rect 19710 948 19728 965
rect 19808 957 19812 968
rect 19803 955 19808 957
rect 19765 950 19766 953
rect 19526 939 19533 942
rect 19550 939 19590 942
rect 19514 936 19550 939
rect 19497 934 19514 936
rect 19090 930 19102 931
rect 18667 921 18676 923
rect 18655 920 18667 921
rect 18694 920 18699 924
rect 18608 915 18694 920
rect 18596 914 18608 915
rect 18636 914 18655 915
rect 18753 914 18761 926
rect 18765 924 18799 926
rect 18461 913 18591 914
rect 18569 909 18583 913
rect 18625 911 18636 914
rect 18618 907 18624 911
rect 18508 900 18514 906
rect 18514 894 18520 900
rect 18542 892 18555 900
rect 18585 892 18596 907
rect 18610 900 18615 904
rect 18747 901 18756 913
rect 18765 901 18767 924
rect 18380 888 18398 890
rect 18542 889 18551 892
rect 18555 891 18557 892
rect 18597 889 18599 891
rect 18607 889 18616 898
rect 18756 892 18767 901
rect 18797 892 18799 924
rect 18803 914 18811 926
rect 18909 924 18919 926
rect 18976 924 19004 926
rect 19005 924 19016 926
rect 18909 923 18917 924
rect 18914 921 18917 923
rect 18969 921 18970 924
rect 19002 921 19016 924
rect 18835 907 18849 921
rect 18904 910 18914 921
rect 18968 917 18969 921
rect 18904 907 18917 910
rect 18967 907 18968 916
rect 19002 915 19004 921
rect 19005 915 19016 921
rect 19039 924 19047 926
rect 19039 915 19046 924
rect 19047 921 19051 924
rect 19050 918 19056 921
rect 19051 916 19056 918
rect 19002 911 19005 915
rect 19007 914 19016 915
rect 19007 912 19008 914
rect 18849 906 18904 907
rect 18911 904 18917 907
rect 18966 904 18967 906
rect 18969 904 18975 910
rect 19002 906 19004 911
rect 19008 907 19010 912
rect 19010 906 19011 907
rect 19001 904 19004 906
rect 19011 904 19012 906
rect 18917 898 18923 904
rect 18959 902 18962 904
rect 18963 902 18969 904
rect 18958 898 18969 902
rect 19000 901 19001 904
rect 18958 892 18965 898
rect 18999 897 19000 900
rect 18997 894 18999 895
rect 19002 894 19004 904
rect 18970 892 19004 894
rect 19008 901 19016 904
rect 19008 892 19022 901
rect 18997 891 18999 892
rect 19022 890 19025 892
rect 18123 879 18127 885
rect 18249 879 18302 886
rect 18312 883 18318 886
rect 18319 883 18331 886
rect 18386 884 18392 888
rect 18120 875 18123 879
rect 18219 875 18249 879
rect 18260 877 18266 879
rect 18065 871 18066 875
rect 18117 870 18120 874
rect 18181 870 18219 875
rect 18179 869 18181 870
rect 18116 868 18117 869
rect 18177 868 18179 869
rect 18268 868 18270 879
rect 18303 868 18304 879
rect 18306 877 18312 883
rect 18380 882 18392 884
rect 18444 882 18450 888
rect 18380 876 18398 882
rect 18438 876 18444 882
rect 18551 880 18560 889
rect 18597 888 18607 889
rect 18995 888 18997 889
rect 18598 887 18607 888
rect 18598 880 18618 887
rect 18800 885 18801 888
rect 18761 882 18762 884
rect 18970 880 18982 888
rect 18992 882 19004 888
rect 19025 884 19027 890
rect 19029 885 19039 915
rect 19056 912 19069 916
rect 19069 907 19081 912
rect 19084 906 19086 907
rect 19095 906 19102 930
rect 19147 928 19148 931
rect 19270 919 19318 934
rect 19338 932 19413 934
rect 19430 933 19481 934
rect 19483 933 19494 934
rect 19430 932 19491 933
rect 19338 930 19430 932
rect 19086 904 19091 906
rect 19095 904 19147 906
rect 19091 901 19147 904
rect 19095 899 19147 901
rect 19078 889 19087 898
rect 19095 896 19164 899
rect 19095 891 19152 896
rect 19164 892 19189 896
rect 19286 894 19294 919
rect 19318 916 19325 919
rect 19338 918 19354 930
rect 19356 918 19372 930
rect 19477 929 19492 932
rect 19473 927 19477 929
rect 19457 922 19473 927
rect 19483 926 19492 929
rect 19526 926 19533 936
rect 19486 920 19491 922
rect 19304 900 19308 916
rect 19325 914 19356 916
rect 19357 914 19359 918
rect 19325 909 19357 914
rect 19348 907 19365 909
rect 19348 902 19357 907
rect 19365 906 19369 907
rect 19308 896 19309 899
rect 19328 898 19348 902
rect 19089 889 19153 891
rect 19189 890 19201 892
rect 19285 890 19286 893
rect 19087 885 19153 889
rect 18991 880 19004 882
rect 18561 875 18564 880
rect 18605 879 18618 880
rect 18103 864 18116 868
rect 18171 864 18177 868
rect 18097 862 18103 864
rect 18168 862 18171 864
rect 18094 858 18097 862
rect 18161 857 18168 862
rect 18093 856 18094 857
rect 18160 856 18161 857
rect 18092 849 18093 856
rect 18157 849 18160 856
rect 18091 841 18092 849
rect 18159 838 18168 842
rect 18206 838 18215 842
rect 18218 838 18234 854
rect 18236 838 18252 854
rect 18270 838 18274 867
rect 18301 847 18303 867
rect 18564 860 18571 875
rect 18603 873 18618 875
rect 18314 849 18328 854
rect 18410 842 18414 856
rect 16625 804 16635 805
rect 18087 804 18091 838
rect 18156 833 18168 838
rect 18202 833 18218 838
rect 18252 837 18268 838
rect 18259 834 18268 837
rect 18150 832 18163 833
rect 18202 832 18224 833
rect 18148 831 18157 832
rect 18148 811 18150 831
rect 18151 826 18157 831
rect 18147 810 18150 811
rect 18148 804 18150 810
rect 18156 820 18157 826
rect 18189 824 18224 832
rect 18189 823 18218 824
rect 18189 822 18237 823
rect 18263 822 18268 834
rect 18189 820 18209 822
rect 18218 820 18237 822
rect 18156 804 18172 820
rect 18202 804 18218 820
rect 18262 812 18263 817
rect 16533 803 16534 804
rect 16532 801 16533 802
rect 16480 799 16523 801
rect 16315 796 16480 799
rect 16315 795 16421 796
rect 16504 795 16523 799
rect 16297 794 16331 795
rect 16279 792 16313 794
rect 16258 789 16287 792
rect 16173 785 16184 788
rect 16233 787 16258 789
rect 16220 786 16233 787
rect 16216 785 16220 786
rect 16075 784 16078 785
rect 16096 784 16184 785
rect 16096 783 16173 784
rect 16189 783 16216 785
rect 16244 784 16247 787
rect 15918 779 15919 780
rect 15956 769 15964 783
rect 15998 778 15999 783
rect 16074 781 16075 783
rect 16097 782 16099 783
rect 16073 778 16074 781
rect 16099 780 16102 782
rect 16107 781 16108 783
rect 16165 782 16189 783
rect 16154 779 16165 782
rect 16102 778 16105 779
rect 15654 756 15672 757
rect 15700 756 15706 758
rect 15648 750 15712 756
rect 15737 753 15767 766
rect 15797 763 15835 769
rect 15953 763 15956 769
rect 15797 759 15829 763
rect 15796 756 15797 758
rect 15737 750 15773 753
rect 15794 752 15796 756
rect 15798 755 15829 759
rect 15826 754 15828 755
rect 15829 754 15832 755
rect 15948 754 15953 763
rect 15825 752 15826 754
rect 15832 751 15837 754
rect 15947 752 15948 754
rect 15548 744 15554 750
rect 15654 745 15706 750
rect 15458 742 15502 744
rect 15307 741 15341 742
rect 15458 741 15464 742
rect 15270 740 15307 741
rect 15247 739 15270 740
rect 15244 737 15247 739
rect 15496 738 15502 742
rect 15554 738 15560 744
rect 15219 723 15244 737
rect 15335 730 15341 736
rect 15393 731 15399 736
rect 15648 733 15660 745
rect 15694 735 15699 745
rect 15424 731 15460 733
rect 15341 724 15347 730
rect 15365 729 15424 731
rect 15460 729 15466 731
rect 15363 726 15365 729
rect 15214 720 15219 723
rect 15112 717 15194 719
rect 15115 716 15194 717
rect 15211 716 15219 720
rect 15161 713 15169 716
rect 15173 715 15175 716
rect 15194 715 15223 716
rect 15173 713 15207 715
rect 15204 709 15207 713
rect 15211 713 15219 715
rect 15223 714 15251 715
rect 15211 711 15214 713
rect 15208 709 15211 711
rect 15251 710 15265 714
rect 15357 713 15363 726
rect 15387 724 15393 729
rect 15466 726 15477 729
rect 15654 726 15660 733
rect 15456 722 15458 723
rect 15477 722 15488 726
rect 15653 723 15660 726
rect 15488 721 15490 722
rect 15490 720 15494 721
rect 14838 707 14839 708
rect 15060 707 15061 708
rect 15173 701 15185 709
rect 15195 701 15207 709
rect 15265 705 15271 710
rect 15355 708 15357 713
rect 15354 707 15355 708
rect 15271 703 15282 705
rect 14899 697 15033 700
rect 15199 698 15203 701
rect 15282 699 15295 703
rect 15295 698 15300 699
rect 14775 695 14899 697
rect 15033 695 15039 697
rect 14678 692 14684 694
rect 14753 692 14775 695
rect 15039 692 15045 695
rect 14460 688 14461 690
rect 14674 688 14676 691
rect 14677 688 14678 690
rect 14730 689 14753 692
rect 15045 689 15051 692
rect 15183 690 15199 698
rect 15300 694 15316 698
rect 15316 692 15332 694
rect 15332 691 15341 692
rect 15347 691 15354 706
rect 15448 693 15456 698
rect 15460 693 15462 720
rect 15648 711 15660 723
rect 15699 711 15701 726
rect 15737 723 15767 750
rect 15793 749 15794 751
rect 15837 750 15839 751
rect 15777 746 15779 747
rect 15791 745 15793 749
rect 15780 737 15794 745
rect 15822 744 15824 749
rect 15842 747 15845 749
rect 15845 746 15847 747
rect 15847 743 15851 746
rect 15871 743 15883 749
rect 15942 744 15945 749
rect 15977 744 15998 778
rect 16064 756 16073 778
rect 16102 776 16107 778
rect 16108 776 16154 779
rect 16247 778 16248 781
rect 16102 775 16154 776
rect 16102 756 16107 775
rect 16248 772 16252 778
rect 16248 756 16255 772
rect 16279 756 16287 789
rect 16297 788 16313 792
rect 16315 788 16331 794
rect 16393 788 16409 795
rect 16507 788 16523 795
rect 16510 787 16511 788
rect 16511 783 16512 785
rect 16513 772 16516 779
rect 16536 778 16548 804
rect 16585 799 16586 802
rect 16585 796 16587 799
rect 16623 796 16625 800
rect 18091 799 18104 804
rect 18121 799 18156 804
rect 18104 797 18121 799
rect 16585 791 16593 796
rect 16620 791 16623 796
rect 16585 788 16601 791
rect 16603 788 16619 791
rect 18140 788 18157 799
rect 18218 797 18221 803
rect 18218 795 18222 797
rect 18218 788 18228 795
rect 18148 786 18157 788
rect 18222 786 18228 788
rect 18273 786 18274 828
rect 18298 822 18311 838
rect 18444 833 18448 838
rect 18466 837 18478 845
rect 18532 838 18548 854
rect 18571 842 18580 860
rect 18572 841 18580 842
rect 18584 845 18585 862
rect 18584 843 18588 845
rect 18616 844 18618 873
rect 18619 869 18630 875
rect 18622 863 18630 869
rect 18626 859 18629 863
rect 18762 860 18766 879
rect 18799 866 18800 880
rect 18881 867 18887 873
rect 18927 867 18933 873
rect 18991 870 18995 880
rect 19024 870 19029 884
rect 19087 880 19101 885
rect 19095 871 19101 880
rect 19137 880 19147 885
rect 19137 870 19138 880
rect 19141 879 19147 880
rect 19201 879 19268 890
rect 19284 885 19285 889
rect 19283 881 19284 885
rect 19269 875 19273 879
rect 19273 872 19276 875
rect 19280 871 19283 881
rect 19309 879 19313 896
rect 19323 891 19328 898
rect 19369 892 19426 906
rect 19426 891 19429 892
rect 19320 881 19322 889
rect 19429 888 19443 891
rect 19489 890 19491 920
rect 19495 910 19503 922
rect 19533 914 19538 926
rect 19538 902 19543 914
rect 19563 910 19570 939
rect 19590 936 19596 939
rect 19596 934 19600 936
rect 19677 935 19678 942
rect 19701 939 19707 942
rect 19707 936 19713 939
rect 19600 933 19601 934
rect 19601 927 19604 933
rect 19604 922 19607 927
rect 19607 919 19609 922
rect 19609 916 19610 919
rect 19460 888 19491 890
rect 19495 888 19503 900
rect 19543 899 19544 902
rect 19570 900 19572 910
rect 19610 902 19617 916
rect 19678 910 19682 935
rect 19713 934 19717 936
rect 19728 935 19729 942
rect 19715 933 19721 934
rect 19715 932 19723 933
rect 19729 932 19730 935
rect 19765 934 19780 950
rect 19803 948 19815 955
rect 19802 947 19815 948
rect 19825 947 19837 955
rect 19868 952 19884 968
rect 19799 945 19808 947
rect 19798 943 19799 945
rect 19802 943 19808 945
rect 19841 943 19842 945
rect 19848 943 19854 948
rect 19791 942 19798 943
rect 19802 942 19837 943
rect 19841 942 19854 943
rect 19791 937 19802 942
rect 19803 941 19837 942
rect 19789 934 19795 937
rect 19796 936 19802 937
rect 19836 936 19837 941
rect 19854 936 19860 942
rect 19868 934 19884 950
rect 19921 939 19928 968
rect 19974 956 19975 968
rect 19979 965 19980 969
rect 20095 968 20114 969
rect 20122 968 20126 969
rect 20086 964 20122 968
rect 20172 965 20176 969
rect 19920 934 19921 938
rect 19785 932 19789 934
rect 19723 931 19764 932
rect 19729 918 19746 931
rect 19748 926 19764 931
rect 19782 930 19785 932
rect 19775 926 19782 930
rect 19867 927 19868 931
rect 19919 927 19920 932
rect 19748 918 19775 926
rect 19866 920 19868 927
rect 19918 922 19919 927
rect 19929 922 19937 934
rect 19941 922 19943 956
rect 19979 951 19980 964
rect 20086 960 20134 964
rect 20077 954 20086 960
rect 19974 945 19975 951
rect 19980 936 19981 945
rect 20069 939 20077 954
rect 20115 949 20134 960
rect 20134 948 20136 949
rect 20176 948 20181 965
rect 20279 961 20282 980
rect 20282 954 20283 960
rect 20136 945 20140 948
rect 20181 945 20182 948
rect 20066 936 20069 939
rect 19981 928 19987 934
rect 19982 922 19987 928
rect 20061 928 20073 936
rect 20083 928 20095 936
rect 20140 934 20155 945
rect 20182 934 20186 945
rect 20283 941 20286 954
rect 20285 939 20286 941
rect 20283 934 20285 939
rect 20155 932 20156 934
rect 20156 928 20157 930
rect 20186 929 20188 934
rect 20061 924 20066 928
rect 20099 926 20100 928
rect 20101 924 20104 925
rect 19865 919 19868 920
rect 19729 905 19730 918
rect 19757 916 19775 918
rect 19864 918 19868 919
rect 19864 916 19865 918
rect 19917 916 19918 919
rect 19937 916 19938 921
rect 19751 912 19757 916
rect 19860 909 19864 916
rect 19916 909 19917 916
rect 19938 912 19940 916
rect 19968 913 19975 922
rect 19982 916 19983 922
rect 19961 911 19968 913
rect 19979 911 19983 916
rect 20049 912 20057 924
rect 20061 922 20095 924
rect 20061 921 20064 922
rect 19941 910 19979 911
rect 19730 902 19731 904
rect 19617 899 19619 902
rect 19572 894 19573 899
rect 19619 896 19620 899
rect 19443 885 19454 888
rect 19457 885 19496 888
rect 19454 884 19496 885
rect 19313 872 19315 879
rect 19315 870 19316 872
rect 19317 871 19320 881
rect 19457 879 19496 884
rect 19545 881 19547 889
rect 19479 876 19491 879
rect 19496 874 19518 879
rect 19547 874 19548 881
rect 19532 872 19537 874
rect 18966 868 18967 869
rect 18990 867 18991 870
rect 18875 861 18881 867
rect 18933 861 18939 867
rect 18988 860 18990 867
rect 18629 854 18633 858
rect 18629 853 18644 854
rect 18615 843 18618 844
rect 18584 841 18618 843
rect 18622 841 18630 853
rect 18633 850 18644 853
rect 18766 852 18767 858
rect 18800 854 18801 858
rect 18635 845 18644 850
rect 18638 840 18644 845
rect 18401 831 18478 833
rect 18301 820 18306 822
rect 18298 804 18311 820
rect 18301 787 18306 804
rect 18314 788 18330 799
rect 18150 780 18157 786
rect 18215 785 18228 786
rect 18215 783 18262 785
rect 18190 780 18237 783
rect 16059 745 16064 756
rect 16099 744 16102 756
rect 16252 750 16255 756
rect 16252 744 16259 750
rect 16287 744 16289 756
rect 16317 751 16329 759
rect 16339 751 16351 759
rect 16516 755 16521 772
rect 16548 770 16552 778
rect 18150 777 18163 780
rect 18203 777 18209 780
rect 18215 779 18237 780
rect 18215 777 18224 779
rect 18401 777 18459 831
rect 18476 799 18478 831
rect 18482 821 18490 833
rect 18548 822 18564 838
rect 18618 837 18622 840
rect 18642 838 18644 840
rect 18666 838 18672 844
rect 18712 839 18718 844
rect 18708 838 18720 839
rect 18767 838 18770 850
rect 18802 841 18818 854
rect 18873 852 18881 858
rect 18871 850 18881 852
rect 18985 851 18988 860
rect 18934 848 18944 850
rect 18944 846 18950 848
rect 18983 847 18985 851
rect 18861 845 18869 846
rect 18871 845 18875 846
rect 18801 840 18818 841
rect 18801 838 18805 840
rect 18584 829 18596 837
rect 18606 829 18618 837
rect 18644 832 18724 838
rect 18770 832 18771 837
rect 18584 828 18585 829
rect 18585 818 18587 828
rect 18644 822 18660 832
rect 18666 831 18720 832
rect 18666 827 18718 831
rect 18587 814 18589 818
rect 18589 809 18590 812
rect 18590 805 18591 809
rect 18591 799 18592 803
rect 18592 792 18594 799
rect 18666 793 18686 827
rect 18712 825 18720 827
rect 18718 794 18720 825
rect 18724 815 18732 827
rect 18712 793 18720 794
rect 18724 793 18732 805
rect 18748 804 18756 820
rect 18771 814 18774 829
rect 18786 822 18805 838
rect 18839 833 18848 842
rect 18861 841 18871 845
rect 18873 844 18875 845
rect 18950 844 18957 846
rect 18873 841 18881 844
rect 18957 843 18961 844
rect 18961 842 18966 843
rect 18982 842 18983 844
rect 18978 841 18989 842
rect 19014 841 19024 869
rect 19029 866 19030 869
rect 19030 854 19033 865
rect 19101 860 19106 870
rect 19277 869 19280 870
rect 19276 865 19280 869
rect 19277 860 19280 865
rect 19307 866 19317 870
rect 19537 866 19554 872
rect 19573 871 19577 890
rect 19620 888 19624 896
rect 19728 890 19731 896
rect 19737 891 19748 908
rect 19803 903 19815 909
rect 19915 908 19916 909
rect 19844 903 19860 908
rect 19914 903 19915 908
rect 19961 903 19968 910
rect 19815 902 19844 903
rect 19913 896 19914 899
rect 19796 890 19802 896
rect 19854 890 19860 896
rect 19624 874 19632 888
rect 19726 885 19728 889
rect 19734 886 19737 890
rect 19106 854 19107 860
rect 19276 854 19279 860
rect 19030 852 19036 854
rect 19033 846 19036 852
rect 19098 849 19114 854
rect 19097 848 19111 849
rect 19116 848 19132 854
rect 19034 841 19036 846
rect 19094 845 19097 848
rect 19111 845 19132 848
rect 19089 841 19094 845
rect 19122 842 19134 845
rect 18861 838 18875 841
rect 18981 839 18982 841
rect 18989 840 19024 841
rect 19035 840 19036 841
rect 19087 840 19089 841
rect 19014 839 19062 840
rect 19085 838 19087 840
rect 19101 839 19113 842
rect 19194 841 19210 854
rect 19212 841 19228 854
rect 19274 847 19276 853
rect 19277 852 19279 854
rect 19307 852 19325 866
rect 19548 863 19563 866
rect 19134 840 19135 841
rect 19187 840 19188 841
rect 19106 838 19113 839
rect 18855 834 18869 838
rect 18855 833 18866 834
rect 18830 824 18839 833
rect 18801 820 18805 822
rect 18786 814 18805 820
rect 18774 809 18775 812
rect 18775 799 18777 808
rect 18786 804 18802 814
rect 18861 812 18869 824
rect 18873 814 18875 838
rect 18978 832 18981 838
rect 18933 815 18939 821
rect 18967 818 18985 832
rect 18973 815 18974 818
rect 18927 814 18933 815
rect 18972 814 18973 815
rect 18873 812 18907 814
rect 18916 812 18975 814
rect 18985 813 18991 818
rect 18986 812 18992 813
rect 18805 808 18806 812
rect 18897 809 18907 812
rect 18911 810 18916 812
rect 18888 808 18897 809
rect 18900 808 18906 809
rect 18908 808 18911 810
rect 18927 809 18933 812
rect 18806 804 18807 808
rect 18873 805 18885 808
rect 18888 805 18907 808
rect 18873 804 18886 805
rect 18802 794 18810 804
rect 18833 800 18885 804
rect 18895 800 18907 805
rect 18963 800 18972 811
rect 18975 810 18983 812
rect 18986 810 18997 812
rect 19005 811 19014 838
rect 19036 822 19052 838
rect 19076 832 19084 838
rect 18983 809 18997 810
rect 18999 809 19005 810
rect 18983 808 19005 809
rect 19036 808 19052 820
rect 19105 811 19107 838
rect 19108 837 19113 838
rect 19110 836 19113 837
rect 19135 838 19136 840
rect 19186 838 19187 840
rect 19111 834 19115 836
rect 19116 832 19117 834
rect 19135 832 19148 838
rect 19109 828 19113 830
rect 18986 804 19052 808
rect 18995 800 19036 804
rect 19076 801 19077 804
rect 18802 793 18812 794
rect 18666 792 18718 793
rect 18802 792 18814 793
rect 18594 789 18600 792
rect 18600 784 18607 789
rect 18660 788 18740 792
rect 18778 790 18779 792
rect 18802 789 18823 792
rect 18802 788 18817 789
rect 18660 786 18724 788
rect 18812 786 18817 788
rect 18823 787 18828 789
rect 18828 786 18832 787
rect 18833 786 18884 800
rect 18896 793 18900 800
rect 18958 793 18963 799
rect 18895 790 18896 793
rect 18956 790 18958 793
rect 18607 783 18608 784
rect 18643 783 18644 785
rect 18609 779 18615 783
rect 18640 779 18643 783
rect 18666 780 18672 786
rect 18708 781 18720 786
rect 18828 785 18839 786
rect 18830 783 18839 785
rect 18830 782 18842 783
rect 18712 780 18718 781
rect 18778 779 18779 781
rect 18615 777 18620 779
rect 18639 777 18640 779
rect 16299 747 16305 750
rect 16353 749 16355 750
rect 16308 747 16312 749
rect 16299 746 16308 747
rect 16298 744 16306 746
rect 16317 745 16353 747
rect 16355 745 16363 747
rect 15820 738 15822 743
rect 15851 741 15883 743
rect 15879 740 15884 741
rect 15886 737 15889 739
rect 15939 738 15942 744
rect 15974 739 15977 744
rect 16057 740 16059 744
rect 16074 740 16086 742
rect 15787 734 15788 737
rect 15794 734 15798 737
rect 15786 732 15787 734
rect 15798 732 15802 734
rect 15818 732 15820 737
rect 15848 736 15849 737
rect 15878 734 15888 737
rect 15889 734 15895 737
rect 15901 734 15907 737
rect 15883 732 15888 734
rect 15783 725 15786 731
rect 15802 729 15806 732
rect 15816 729 15818 731
rect 15782 722 15783 724
rect 15778 711 15782 721
rect 15806 712 15834 729
rect 15847 726 15848 731
rect 15888 727 15892 732
rect 15894 731 15907 734
rect 15932 732 15936 734
rect 15930 731 15932 732
rect 15947 731 15953 737
rect 16037 734 16043 740
rect 16055 734 16056 736
rect 16074 734 16089 740
rect 16098 738 16099 742
rect 16247 738 16253 744
rect 16305 738 16311 744
rect 16317 743 16319 745
rect 16097 734 16098 737
rect 15970 732 15971 734
rect 16031 732 16095 734
rect 15892 726 15894 727
rect 15895 726 15901 731
rect 15649 710 15653 711
rect 15654 710 15706 711
rect 15648 706 15712 710
rect 15643 704 15712 706
rect 15775 704 15778 711
rect 15502 698 15508 699
rect 15516 698 15554 699
rect 15496 695 15508 698
rect 15512 695 15560 698
rect 15496 693 15502 695
rect 15512 693 15550 695
rect 15554 693 15560 695
rect 15448 692 15560 693
rect 15448 691 15542 692
rect 15051 688 15054 689
rect 15058 688 15060 690
rect 12994 674 12997 685
rect 12310 653 12311 655
rect 12453 654 12454 656
rect 11242 651 11244 652
rect 11109 649 11185 651
rect 11237 649 11242 651
rect 11477 649 11481 652
rect 11540 650 11542 652
rect 11530 649 11540 650
rect 11192 648 11236 649
rect 11488 640 11504 649
rect 11505 648 11506 649
rect 11770 647 11772 651
rect 11790 647 11902 652
rect 11784 644 11902 647
rect 12000 644 12149 652
rect 11784 640 11800 644
rect 11902 641 11913 644
rect 11953 641 12000 644
rect 11913 640 11953 641
rect 12090 640 12106 644
rect 8898 639 8899 640
rect 12152 636 12182 652
rect 12290 640 12306 653
rect 12453 644 12463 654
rect 12726 652 12739 660
rect 12794 656 12810 672
rect 12932 665 12941 674
rect 12994 667 13006 674
rect 14461 669 14471 688
rect 14672 682 14678 688
rect 14730 682 14736 688
rect 15054 686 15060 688
rect 14677 680 14690 682
rect 14677 676 14684 680
rect 14724 676 14730 682
rect 15058 677 15060 686
rect 15160 681 15183 690
rect 15341 689 15363 691
rect 15448 689 15538 691
rect 15160 679 15230 681
rect 12997 665 13006 667
rect 12934 656 12935 665
rect 12941 656 12950 665
rect 12988 656 13002 665
rect 14471 658 14481 669
rect 14473 656 14487 658
rect 14523 656 14539 672
rect 14677 668 14678 676
rect 15054 671 15060 677
rect 15112 678 15183 679
rect 15112 676 15176 678
rect 15230 676 15239 679
rect 15112 671 15118 676
rect 14677 656 14689 668
rect 15057 665 15066 671
rect 15106 665 15112 671
rect 15057 662 15060 665
rect 15141 662 15160 676
rect 15239 675 15243 676
rect 15243 672 15245 675
rect 15247 667 15248 669
rect 15057 658 15059 662
rect 15137 659 15141 662
rect 15248 660 15263 667
rect 15347 662 15353 689
rect 15363 686 15398 689
rect 15448 686 15532 689
rect 15548 686 15554 692
rect 15643 690 15648 704
rect 15654 699 15672 704
rect 15654 698 15660 699
rect 15700 698 15706 704
rect 15773 699 15775 704
rect 15701 696 15702 698
rect 15771 695 15773 698
rect 15807 695 15815 712
rect 15835 709 15838 711
rect 15843 709 15847 726
rect 15894 717 15904 726
rect 15953 725 15959 731
rect 15966 725 15970 732
rect 16031 730 16089 732
rect 16090 730 16095 732
rect 16096 730 16097 732
rect 16031 728 16087 730
rect 15964 722 15965 724
rect 15904 709 15906 717
rect 15958 711 15964 721
rect 15838 708 15840 709
rect 15837 707 15841 708
rect 15837 703 15843 707
rect 15849 705 15850 707
rect 15849 703 15866 705
rect 15768 694 15771 695
rect 15764 692 15768 694
rect 15762 691 15764 692
rect 15398 684 15417 686
rect 15456 684 15520 686
rect 15417 683 15425 684
rect 15425 681 15446 683
rect 15456 681 15515 684
rect 15446 679 15515 681
rect 15639 679 15643 689
rect 15702 686 15704 690
rect 15758 689 15762 691
rect 15754 688 15758 689
rect 15804 688 15807 695
rect 15840 690 15843 703
rect 15846 699 15848 700
rect 15849 696 15873 699
rect 15849 691 15861 696
rect 15873 693 15887 696
rect 15906 693 15908 706
rect 15953 702 15958 711
rect 16037 696 16052 728
rect 16084 726 16087 728
rect 16090 726 16098 730
rect 16084 724 16086 726
rect 16085 700 16086 724
rect 16087 718 16098 726
rect 16087 714 16091 718
rect 16087 710 16090 714
rect 16093 712 16095 718
rect 16349 715 16351 745
rect 16353 742 16363 745
rect 16523 743 16525 749
rect 16533 743 16539 749
rect 16552 746 16575 770
rect 18037 755 18038 775
rect 18066 772 18067 775
rect 18157 774 18196 777
rect 18203 774 18215 777
rect 18067 759 18075 772
rect 18159 768 18196 774
rect 18206 768 18215 774
rect 18272 768 18273 777
rect 18067 755 18078 759
rect 18038 749 18039 755
rect 18075 753 18078 755
rect 18076 750 18081 753
rect 16579 743 16585 749
rect 18050 747 18079 748
rect 18082 747 18083 749
rect 16527 742 16533 743
rect 16355 738 16363 742
rect 16355 735 16373 738
rect 16363 731 16373 735
rect 16525 731 16533 742
rect 16538 738 16539 742
rect 16571 739 16577 742
rect 16536 731 16538 738
rect 16572 737 16577 739
rect 16585 737 16591 743
rect 16323 714 16351 715
rect 16318 713 16351 714
rect 16355 713 16363 725
rect 16373 721 16379 731
rect 16525 721 16536 731
rect 16517 720 16536 721
rect 16517 712 16526 720
rect 16092 710 16093 711
rect 16090 707 16094 710
rect 16352 709 16355 711
rect 16326 708 16329 709
rect 16089 702 16094 707
rect 16314 706 16324 708
rect 16305 704 16314 706
rect 16084 696 16086 699
rect 15887 692 15953 693
rect 15893 691 15953 692
rect 15727 686 15754 688
rect 15803 686 15804 688
rect 15702 684 15734 686
rect 15692 683 15734 684
rect 15665 681 15734 683
rect 15647 679 15734 681
rect 15800 679 15803 684
rect 15456 678 15515 679
rect 15459 677 15494 678
rect 15620 677 15734 679
rect 15459 676 15491 677
rect 15493 676 15494 677
rect 15460 674 15472 676
rect 15474 675 15493 676
rect 15598 675 15620 677
rect 15626 676 15734 677
rect 15639 675 15643 676
rect 15474 671 15501 675
rect 15550 671 15598 675
rect 15474 670 15512 671
rect 15539 670 15582 671
rect 15474 664 15582 670
rect 15476 662 15486 664
rect 15639 662 15640 675
rect 15704 672 15706 675
rect 15797 673 15800 679
rect 15353 660 15354 662
rect 15135 658 15137 659
rect 14837 656 14839 657
rect 15057 656 15058 658
rect 15133 656 15135 658
rect 12761 652 12794 656
rect 12994 652 12997 656
rect 12741 651 12760 652
rect 12509 645 12510 651
rect 12464 640 12480 644
rect 12482 640 12498 644
rect 12778 640 12794 652
rect 12935 645 12945 652
rect 12989 646 12994 652
rect 12983 645 12989 646
rect 12945 644 12986 645
rect 12970 640 12986 644
rect 14489 640 14505 656
rect 14507 640 14523 656
rect 14690 653 14692 656
rect 14830 653 14836 656
rect 15059 653 15062 656
rect 15129 653 15133 656
rect 14692 651 14694 653
rect 14829 652 14830 653
rect 15127 652 15129 653
rect 15263 652 15375 660
rect 15467 658 15476 662
rect 15704 659 15707 672
rect 15836 666 15840 689
rect 15899 685 15953 691
rect 16037 688 16089 696
rect 16090 692 16094 702
rect 16247 693 16253 698
rect 16305 693 16311 698
rect 16247 692 16311 693
rect 16094 688 16096 690
rect 15895 679 15959 685
rect 16031 682 16096 688
rect 16253 686 16259 692
rect 16299 686 16305 692
rect 16317 690 16318 706
rect 16339 701 16351 709
rect 16530 707 16536 720
rect 16573 717 16577 737
rect 16529 706 16530 707
rect 16525 697 16529 706
rect 16577 697 16579 717
rect 17340 703 17362 722
rect 18032 713 18039 725
rect 18044 716 18045 747
rect 18073 745 18078 747
rect 18077 716 18078 745
rect 18079 738 18090 747
rect 18306 740 18310 777
rect 18615 776 18639 777
rect 18776 775 18778 779
rect 18830 777 18839 782
rect 18845 779 18848 781
rect 18848 777 18867 779
rect 18895 777 18904 786
rect 18926 782 18932 788
rect 18953 786 18956 790
rect 18972 782 18978 788
rect 18990 786 18999 800
rect 19002 788 19018 800
rect 19020 796 19056 800
rect 19077 798 19079 801
rect 19104 800 19105 810
rect 19111 798 19113 828
rect 19117 818 19125 830
rect 19134 822 19148 832
rect 19178 836 19186 838
rect 19240 837 19244 841
rect 19272 839 19274 847
rect 19307 838 19317 852
rect 19325 848 19328 852
rect 19455 842 19461 844
rect 19455 838 19469 842
rect 19501 838 19507 844
rect 19508 838 19524 854
rect 19548 838 19554 863
rect 19563 853 19566 863
rect 19566 846 19568 852
rect 19568 838 19571 845
rect 19178 822 19185 836
rect 19202 826 19214 832
rect 19199 825 19258 826
rect 19262 825 19272 838
rect 19199 823 19207 825
rect 19258 823 19272 825
rect 19279 823 19282 838
rect 19134 820 19137 822
rect 19198 821 19199 823
rect 19077 796 19113 798
rect 19117 796 19125 808
rect 19134 804 19148 820
rect 19190 816 19198 820
rect 19202 818 19209 820
rect 19190 808 19196 816
rect 19202 814 19203 818
rect 19262 816 19287 823
rect 19296 816 19307 837
rect 19328 822 19340 838
rect 19449 832 19455 838
rect 19453 830 19455 832
rect 19457 830 19490 838
rect 19507 832 19513 838
rect 19524 832 19540 838
rect 19554 832 19555 838
rect 19507 830 19540 832
rect 19571 830 19574 838
rect 19577 830 19589 870
rect 19632 863 19637 874
rect 19679 871 19682 885
rect 19716 881 19726 885
rect 19802 884 19808 890
rect 19812 887 19813 890
rect 19822 886 19829 890
rect 19813 883 19816 885
rect 19819 884 19821 885
rect 19848 884 19854 890
rect 19911 888 19913 896
rect 19813 882 19818 883
rect 19714 874 19732 881
rect 19697 870 19714 874
rect 19716 870 19726 874
rect 19637 859 19639 863
rect 19663 838 19679 870
rect 19697 866 19716 870
rect 19695 863 19697 866
rect 19693 859 19695 863
rect 19709 859 19716 866
rect 19691 856 19693 859
rect 19689 854 19691 856
rect 19682 851 19691 854
rect 19682 845 19689 851
rect 19682 839 19686 845
rect 19682 838 19683 839
rect 19639 830 19640 838
rect 19663 830 19682 838
rect 19696 830 19709 859
rect 19726 846 19733 858
rect 19738 848 19739 880
rect 19805 876 19811 879
rect 19802 874 19805 876
rect 19793 869 19802 874
rect 19813 870 19816 882
rect 19850 870 19853 884
rect 19910 881 19911 888
rect 19909 874 19910 881
rect 19786 860 19787 863
rect 19816 860 19818 870
rect 19850 862 19864 870
rect 19906 863 19909 874
rect 19781 848 19786 860
rect 19738 847 19743 848
rect 19738 846 19772 847
rect 19779 846 19784 848
rect 19733 844 19734 846
rect 19778 844 19779 846
rect 19775 842 19777 843
rect 19738 834 19750 841
rect 19760 834 19772 841
rect 19818 830 19829 859
rect 19853 830 19864 862
rect 19905 856 19906 859
rect 19943 856 19961 903
rect 20049 890 20057 902
rect 20061 890 20063 921
rect 20094 920 20095 922
rect 20101 912 20107 924
rect 20157 913 20159 925
rect 20188 924 20204 928
rect 20274 925 20283 934
rect 20266 924 20274 925
rect 20188 913 20266 924
rect 20101 911 20104 912
rect 20104 903 20109 910
rect 20142 905 20204 913
rect 20136 903 20142 905
rect 20095 890 20136 903
rect 20104 888 20109 890
rect 20159 889 20161 905
rect 20057 886 20060 888
rect 20109 886 20110 888
rect 20161 885 20162 888
rect 20060 884 20062 885
rect 20061 883 20063 884
rect 20061 879 20064 883
rect 20110 880 20111 882
rect 20061 878 20065 879
rect 20064 876 20065 878
rect 20111 876 20112 880
rect 20162 876 20163 879
rect 20188 878 20204 905
rect 20065 869 20068 874
rect 20068 863 20070 869
rect 20003 861 20004 862
rect 20070 860 20071 863
rect 19882 851 19898 854
rect 19902 851 19905 856
rect 19941 851 19943 856
rect 19984 854 19996 855
rect 19882 845 19902 851
rect 19939 846 19941 851
rect 19978 847 19996 854
rect 20006 849 20018 855
rect 20006 847 20055 849
rect 20071 848 20075 860
rect 19978 845 19994 847
rect 20007 846 20055 847
rect 20000 845 20007 846
rect 20027 845 20055 846
rect 19882 843 19888 845
rect 19938 843 19939 845
rect 19978 843 20000 845
rect 20055 843 20069 845
rect 20075 844 20076 847
rect 20092 843 20108 854
rect 19880 839 19883 843
rect 19936 839 19938 843
rect 19972 842 19977 843
rect 19972 840 19976 842
rect 19978 841 20018 843
rect 19965 839 19975 840
rect 19978 839 19984 841
rect 19959 838 19964 839
rect 19978 838 19979 839
rect 19866 830 19880 838
rect 19933 836 19936 838
rect 19955 837 19959 838
rect 19946 836 19952 837
rect 19933 834 19946 836
rect 19923 833 19927 834
rect 19917 832 19923 833
rect 19904 830 19917 832
rect 19933 831 19936 834
rect 19445 827 19453 830
rect 19457 828 19460 830
rect 19444 821 19454 827
rect 19133 802 19134 804
rect 19135 800 19137 804
rect 19262 801 19272 816
rect 19274 812 19282 816
rect 19274 804 19283 812
rect 19287 807 19319 816
rect 19328 807 19340 820
rect 19420 807 19444 821
rect 19445 818 19453 821
rect 19283 801 19284 803
rect 19296 801 19307 807
rect 19319 804 19340 807
rect 19020 788 19036 796
rect 19056 795 19061 796
rect 19061 793 19072 795
rect 19079 794 19086 796
rect 19086 793 19092 794
rect 19103 793 19104 796
rect 19072 792 19077 793
rect 19092 792 19112 793
rect 19115 792 19117 795
rect 19132 794 19133 796
rect 19092 786 19113 792
rect 19129 789 19132 793
rect 19114 788 19132 789
rect 19114 786 19129 788
rect 19185 786 19186 788
rect 19190 786 19196 798
rect 19244 789 19245 801
rect 19259 790 19262 800
rect 19284 797 19312 801
rect 19319 797 19338 804
rect 19408 800 19420 807
rect 19406 799 19408 800
rect 19284 796 19338 797
rect 19399 796 19406 799
rect 19445 796 19453 808
rect 19457 796 19459 828
rect 19525 822 19754 830
rect 19525 820 19527 822
rect 19528 820 19754 822
rect 19525 814 19754 820
rect 19782 814 19904 830
rect 19927 818 19933 831
rect 19962 822 19978 838
rect 19925 815 19932 818
rect 19525 812 19782 814
rect 19527 804 19540 812
rect 19557 807 19559 812
rect 19527 803 19528 804
rect 19528 801 19529 802
rect 19525 796 19528 801
rect 19558 800 19559 807
rect 19570 804 19582 812
rect 19582 803 19583 804
rect 19587 803 19589 808
rect 19606 803 19685 812
rect 19583 802 19685 803
rect 19586 799 19602 802
rect 19203 787 19204 788
rect 19202 786 19208 787
rect 18984 782 18990 786
rect 19101 784 19113 786
rect 18775 772 18776 774
rect 18839 772 18867 777
rect 18768 759 18775 772
rect 18839 768 18848 772
rect 18886 768 18895 777
rect 18920 776 18926 782
rect 18978 776 18990 782
rect 19102 776 19103 781
rect 18978 766 18982 773
rect 19134 772 19135 786
rect 19186 783 19187 786
rect 19197 784 19199 785
rect 19243 784 19244 788
rect 19258 787 19259 790
rect 19284 789 19328 796
rect 19338 795 19340 796
rect 19340 792 19347 795
rect 19397 793 19399 796
rect 19496 795 19524 796
rect 19347 789 19351 792
rect 19284 788 19306 789
rect 19308 788 19324 789
rect 19351 788 19353 789
rect 19393 788 19397 793
rect 19508 792 19524 795
rect 19554 793 19558 799
rect 19265 787 19272 788
rect 19280 787 19294 788
rect 19353 787 19356 788
rect 19257 786 19265 787
rect 19252 785 19265 786
rect 19284 785 19294 787
rect 19449 786 19455 792
rect 19507 791 19524 792
rect 19551 791 19554 793
rect 19507 789 19563 791
rect 19584 789 19602 799
rect 19507 788 19524 789
rect 19551 788 19554 789
rect 19563 788 19602 789
rect 19604 788 19685 802
rect 19696 800 19709 812
rect 19772 804 19773 807
rect 19507 786 19513 788
rect 19550 786 19551 788
rect 19249 784 19258 785
rect 19187 780 19199 783
rect 19202 780 19203 781
rect 19211 780 19249 784
rect 19187 779 19246 780
rect 19202 774 19214 779
rect 19133 763 19135 772
rect 19252 763 19258 784
rect 19284 784 19298 785
rect 18758 756 18775 759
rect 19099 756 19102 763
rect 18758 755 18768 756
rect 18758 754 18765 755
rect 19098 754 19099 756
rect 18758 753 18762 754
rect 18747 749 18789 753
rect 18747 748 18774 749
rect 18745 747 18747 748
rect 18789 747 18792 749
rect 18731 745 18745 747
rect 18263 738 18269 740
rect 18306 739 18315 740
rect 18083 735 18101 738
rect 18090 725 18101 735
rect 18263 734 18275 738
rect 18309 734 18315 739
rect 18698 738 18731 745
rect 18692 737 18697 738
rect 18257 728 18263 734
rect 18315 729 18321 734
rect 18669 733 18692 737
rect 18746 735 18754 747
rect 18758 746 18763 747
rect 18663 731 18669 733
rect 18657 729 18659 731
rect 18279 728 18410 729
rect 18263 726 18279 728
rect 18315 727 18618 728
rect 18645 727 18651 729
rect 18656 728 18657 729
rect 18410 726 18411 727
rect 18618 726 18651 727
rect 18654 726 18656 728
rect 18044 714 18048 716
rect 18075 714 18078 716
rect 18044 713 18078 714
rect 18083 713 18101 725
rect 18251 714 18259 726
rect 18263 724 18269 726
rect 18039 711 18040 713
rect 18040 708 18045 711
rect 18078 708 18083 711
rect 18044 707 18056 708
rect 17311 697 17334 698
rect 17339 697 17362 703
rect 18043 701 18056 707
rect 18066 701 18078 708
rect 18090 707 18101 713
rect 16525 693 16533 697
rect 16585 693 16591 697
rect 18043 694 18045 701
rect 16525 691 16591 693
rect 16525 690 16529 691
rect 16318 686 16320 690
rect 15899 673 15907 679
rect 15947 673 15953 679
rect 16037 676 16043 682
rect 16083 676 16089 682
rect 15899 666 15906 673
rect 16039 672 16042 676
rect 15463 656 15467 658
rect 15640 656 15641 658
rect 15705 657 15707 659
rect 15703 656 15707 657
rect 15458 653 15463 656
rect 15641 653 15644 656
rect 15702 653 15703 656
rect 15737 654 15767 663
rect 15771 654 15784 660
rect 15836 659 15838 666
rect 15899 665 15907 666
rect 15453 652 15454 653
rect 15701 652 15702 653
rect 15734 652 15771 654
rect 15838 653 15840 659
rect 15896 656 15907 665
rect 16033 660 16042 672
rect 16095 672 16096 682
rect 16033 656 16039 660
rect 16095 656 16099 672
rect 16311 660 16320 686
rect 16519 674 16525 690
rect 16533 685 16539 691
rect 16579 685 16585 691
rect 18101 690 18108 707
rect 18251 692 18259 704
rect 18263 694 18265 724
rect 18412 719 18416 726
rect 18618 723 18653 726
rect 18691 723 18697 729
rect 18416 708 18423 719
rect 18639 717 18645 723
rect 18646 719 18653 723
rect 18697 719 18703 723
rect 18746 719 18754 725
rect 18758 719 18760 746
rect 19087 744 19093 750
rect 19095 744 19098 754
rect 19133 750 19134 763
rect 19239 757 19245 762
rect 19251 757 19252 762
rect 19284 758 19294 784
rect 19298 783 19302 784
rect 19357 783 19363 786
rect 19392 783 19393 786
rect 19455 784 19469 786
rect 19455 783 19461 784
rect 19493 783 19497 784
rect 19364 781 19366 782
rect 19366 780 19369 781
rect 19382 780 19392 783
rect 19311 775 19317 779
rect 19317 772 19322 775
rect 19369 772 19392 780
rect 19323 766 19347 772
rect 19382 769 19414 772
rect 19420 769 19493 783
rect 19501 780 19507 786
rect 19508 784 19509 785
rect 19549 784 19550 786
rect 19584 783 19587 788
rect 19593 787 19685 788
rect 19657 786 19685 787
rect 19634 785 19685 786
rect 19693 785 19696 799
rect 19771 797 19772 801
rect 19818 800 19829 814
rect 19853 804 19864 814
rect 19866 804 19882 814
rect 19919 807 19932 815
rect 19916 805 19932 807
rect 19962 805 19978 820
rect 20016 811 20018 841
rect 20022 831 20030 843
rect 20069 838 20109 843
rect 20112 842 20119 874
rect 20154 840 20162 852
rect 20166 842 20168 874
rect 20198 857 20203 874
rect 20198 842 20200 857
rect 20203 852 20204 856
rect 20166 840 20200 842
rect 20204 840 20212 852
rect 20119 838 20120 840
rect 20206 838 20208 840
rect 20109 837 20124 838
rect 20166 837 20167 838
rect 20118 836 20124 837
rect 20163 836 20165 837
rect 20000 809 20018 811
rect 20022 809 20030 821
rect 20079 805 20089 836
rect 20118 832 20133 836
rect 20121 808 20133 832
rect 20166 828 20178 836
rect 20188 828 20200 836
rect 20206 828 20220 838
rect 20167 820 20169 828
rect 20160 818 20169 820
rect 20120 807 20133 808
rect 19905 804 20018 805
rect 19882 803 20018 804
rect 19770 791 19771 796
rect 19769 788 19770 791
rect 19829 789 19832 799
rect 19864 794 19872 800
rect 19882 795 19898 803
rect 19900 799 20018 803
rect 20089 801 20093 805
rect 20119 804 20133 807
rect 20154 815 20169 818
rect 20208 822 20220 828
rect 20208 820 20210 822
rect 20154 804 20170 815
rect 20208 805 20220 820
rect 20660 819 20661 1015
rect 20850 819 20851 1015
rect 20936 819 20937 1015
rect 21209 819 21210 1015
rect 21406 819 21407 1015
rect 20210 804 20220 805
rect 20118 803 20119 804
rect 20117 801 20118 802
rect 20065 799 20108 801
rect 19900 796 20065 799
rect 19900 795 20006 796
rect 20089 795 20108 799
rect 19882 794 19916 795
rect 19864 792 19898 794
rect 19843 789 19872 792
rect 19758 785 19769 788
rect 19818 787 19843 789
rect 19805 786 19818 787
rect 19801 785 19805 786
rect 19660 784 19663 785
rect 19681 784 19769 785
rect 19681 783 19758 784
rect 19774 783 19801 785
rect 19829 784 19832 787
rect 19503 779 19504 780
rect 19541 769 19549 783
rect 19583 778 19584 783
rect 19659 781 19660 783
rect 19682 782 19684 783
rect 19658 778 19659 781
rect 19684 780 19687 782
rect 19692 781 19693 783
rect 19750 782 19774 783
rect 19739 779 19750 782
rect 19687 778 19690 779
rect 19239 756 19257 757
rect 19285 756 19291 758
rect 19233 750 19297 756
rect 19322 753 19352 766
rect 19382 763 19420 769
rect 19538 763 19541 769
rect 19382 759 19414 763
rect 19381 756 19382 758
rect 19322 750 19358 753
rect 19379 752 19381 756
rect 19383 755 19414 759
rect 19411 754 19413 755
rect 19414 754 19417 755
rect 19533 754 19538 763
rect 19410 752 19411 754
rect 19417 751 19422 754
rect 19532 752 19533 754
rect 19133 744 19139 750
rect 19239 745 19291 750
rect 19043 742 19087 744
rect 18892 741 18926 742
rect 19043 741 19049 742
rect 18855 740 18892 741
rect 18832 739 18855 740
rect 18829 737 18832 739
rect 19081 738 19087 742
rect 19139 738 19145 744
rect 18804 723 18829 737
rect 18920 730 18926 736
rect 18978 731 18984 736
rect 19233 733 19245 745
rect 19279 735 19284 745
rect 19009 731 19045 733
rect 18926 724 18932 730
rect 18950 729 19009 731
rect 19045 729 19051 731
rect 18948 726 18950 729
rect 18799 720 18804 723
rect 18697 717 18779 719
rect 18700 716 18779 717
rect 18796 716 18804 720
rect 18746 713 18754 716
rect 18758 715 18760 716
rect 18779 715 18808 716
rect 18758 713 18792 715
rect 18789 709 18792 713
rect 18796 713 18804 715
rect 18808 714 18836 715
rect 18796 711 18799 713
rect 18793 709 18796 711
rect 18836 710 18850 714
rect 18942 713 18948 726
rect 18972 724 18978 729
rect 19051 726 19062 729
rect 19239 726 19245 733
rect 19041 722 19043 723
rect 19062 722 19073 726
rect 19238 723 19245 726
rect 19073 721 19075 722
rect 19075 720 19079 721
rect 18423 707 18424 708
rect 18645 707 18646 708
rect 18758 701 18770 709
rect 18780 701 18792 709
rect 18850 705 18856 710
rect 18940 708 18942 713
rect 18939 707 18940 708
rect 18856 703 18867 705
rect 18484 697 18618 700
rect 18784 698 18788 701
rect 18867 699 18880 703
rect 18880 698 18885 699
rect 18360 695 18484 697
rect 18618 695 18624 697
rect 18263 692 18269 694
rect 18338 692 18360 695
rect 18624 692 18630 695
rect 18045 688 18046 690
rect 18259 688 18261 691
rect 18262 688 18263 690
rect 18315 689 18338 692
rect 18630 689 18636 692
rect 18768 690 18784 698
rect 18885 694 18901 698
rect 18901 692 18917 694
rect 18917 691 18926 692
rect 18932 691 18939 706
rect 19033 693 19041 698
rect 19045 693 19047 720
rect 19233 711 19245 723
rect 19284 711 19286 726
rect 19322 723 19352 750
rect 19378 749 19379 751
rect 19422 750 19424 751
rect 19362 746 19364 747
rect 19376 745 19378 749
rect 19365 737 19379 745
rect 19407 744 19409 749
rect 19427 747 19430 749
rect 19430 746 19432 747
rect 19432 743 19436 746
rect 19456 743 19468 749
rect 19527 744 19530 749
rect 19562 744 19583 778
rect 19649 756 19658 778
rect 19687 776 19692 778
rect 19693 776 19739 779
rect 19832 778 19833 781
rect 19687 775 19739 776
rect 19687 756 19692 775
rect 19833 772 19837 778
rect 19833 756 19840 772
rect 19864 756 19872 789
rect 19882 788 19898 792
rect 19900 788 19916 794
rect 19978 788 19994 795
rect 20092 788 20108 795
rect 20095 787 20096 788
rect 20096 783 20097 785
rect 20098 772 20101 779
rect 20121 778 20133 804
rect 20170 799 20171 802
rect 20170 796 20172 799
rect 20208 796 20210 800
rect 20170 791 20178 796
rect 20205 791 20208 796
rect 20170 788 20186 791
rect 20188 788 20204 791
rect 19644 745 19649 756
rect 19684 744 19687 756
rect 19837 750 19840 756
rect 19837 744 19844 750
rect 19872 744 19874 756
rect 19902 751 19914 759
rect 19924 751 19936 759
rect 20101 755 20106 772
rect 20133 770 20137 778
rect 19884 747 19890 750
rect 19938 749 19940 750
rect 19893 747 19897 749
rect 19884 746 19893 747
rect 19883 744 19891 746
rect 19902 745 19938 747
rect 19940 745 19948 747
rect 19405 738 19407 743
rect 19436 741 19468 743
rect 19464 740 19469 741
rect 19471 737 19474 739
rect 19524 738 19527 744
rect 19559 739 19562 744
rect 19642 740 19644 744
rect 19659 740 19671 742
rect 19372 734 19373 737
rect 19379 734 19383 737
rect 19371 732 19372 734
rect 19383 732 19387 734
rect 19403 732 19405 737
rect 19433 736 19434 737
rect 19463 734 19473 737
rect 19474 734 19480 737
rect 19486 734 19492 737
rect 19468 732 19473 734
rect 19368 725 19371 731
rect 19387 729 19391 732
rect 19401 729 19403 731
rect 19367 722 19368 724
rect 19363 711 19367 721
rect 19391 712 19419 729
rect 19432 726 19433 731
rect 19473 727 19477 732
rect 19479 731 19492 734
rect 19517 732 19521 734
rect 19515 731 19517 732
rect 19532 731 19538 737
rect 19622 734 19628 740
rect 19640 734 19641 736
rect 19659 734 19674 740
rect 19683 738 19684 742
rect 19832 738 19838 744
rect 19890 738 19896 744
rect 19902 743 19904 745
rect 19682 734 19683 737
rect 19555 732 19556 734
rect 19616 732 19680 734
rect 19477 726 19479 727
rect 19480 726 19486 731
rect 19234 710 19238 711
rect 19239 710 19291 711
rect 19233 706 19297 710
rect 19228 704 19297 706
rect 19360 704 19363 711
rect 19087 698 19093 699
rect 19101 698 19139 699
rect 19081 695 19093 698
rect 19097 695 19145 698
rect 19081 693 19087 695
rect 19097 693 19135 695
rect 19139 693 19145 695
rect 19033 692 19145 693
rect 19033 691 19127 692
rect 18636 688 18639 689
rect 18643 688 18645 690
rect 16579 674 16582 685
rect 15895 653 15896 655
rect 16038 654 16039 656
rect 14827 651 14829 652
rect 14694 649 14770 651
rect 14822 649 14827 651
rect 15062 649 15066 652
rect 15125 650 15127 652
rect 15115 649 15125 650
rect 14777 648 14821 649
rect 15073 640 15089 649
rect 15090 648 15091 649
rect 15355 647 15357 651
rect 15375 647 15487 652
rect 15369 644 15487 647
rect 15585 644 15734 652
rect 15369 640 15385 644
rect 15487 641 15498 644
rect 15538 641 15585 644
rect 15498 640 15538 641
rect 15675 640 15691 644
rect 12483 639 12484 640
rect 15737 636 15767 652
rect 15875 640 15891 653
rect 16038 644 16048 654
rect 16311 652 16324 660
rect 16379 656 16395 672
rect 16517 665 16526 674
rect 16579 667 16591 674
rect 18046 669 18056 688
rect 18257 682 18263 688
rect 18315 682 18321 688
rect 18639 686 18645 688
rect 18262 680 18275 682
rect 18262 676 18269 680
rect 18309 676 18315 682
rect 18643 677 18645 686
rect 18745 681 18768 690
rect 18926 689 18948 691
rect 19033 689 19123 691
rect 18745 679 18815 681
rect 16582 665 16591 667
rect 16519 656 16520 665
rect 16526 656 16535 665
rect 16573 656 16587 665
rect 18056 658 18066 669
rect 18058 656 18072 658
rect 18108 656 18124 672
rect 18262 668 18263 676
rect 18639 671 18645 677
rect 18697 678 18768 679
rect 18697 676 18761 678
rect 18815 676 18824 679
rect 18697 671 18703 676
rect 18262 656 18274 668
rect 18642 665 18651 671
rect 18691 665 18697 671
rect 18642 662 18645 665
rect 18726 662 18745 676
rect 18824 675 18828 676
rect 18828 672 18830 675
rect 18832 667 18833 669
rect 18642 658 18644 662
rect 18722 659 18726 662
rect 18833 660 18848 667
rect 18932 662 18938 689
rect 18948 686 18983 689
rect 19033 686 19117 689
rect 19133 686 19139 692
rect 19228 690 19233 704
rect 19239 699 19257 704
rect 19239 698 19245 699
rect 19285 698 19291 704
rect 19358 699 19360 704
rect 19286 696 19287 698
rect 19356 695 19358 698
rect 19392 695 19400 712
rect 19420 709 19423 711
rect 19428 709 19432 726
rect 19479 717 19489 726
rect 19538 725 19544 731
rect 19551 725 19555 732
rect 19616 730 19674 732
rect 19675 730 19680 732
rect 19681 730 19682 732
rect 19616 728 19672 730
rect 19549 722 19550 724
rect 19489 709 19491 717
rect 19543 711 19549 721
rect 19423 708 19425 709
rect 19422 707 19426 708
rect 19422 703 19428 707
rect 19434 705 19435 707
rect 19434 703 19451 705
rect 19353 694 19356 695
rect 19349 692 19353 694
rect 19347 691 19349 692
rect 18983 684 19002 686
rect 19041 684 19105 686
rect 19002 683 19010 684
rect 19010 681 19031 683
rect 19041 681 19100 684
rect 19031 679 19100 681
rect 19224 679 19228 689
rect 19287 686 19289 690
rect 19343 689 19347 691
rect 19339 688 19343 689
rect 19389 688 19392 695
rect 19425 690 19428 703
rect 19431 699 19433 700
rect 19434 696 19458 699
rect 19434 691 19446 696
rect 19458 693 19472 696
rect 19491 693 19493 706
rect 19538 702 19543 711
rect 19622 696 19637 728
rect 19669 726 19672 728
rect 19675 726 19683 730
rect 19669 724 19671 726
rect 19670 700 19671 724
rect 19672 718 19683 726
rect 19672 714 19676 718
rect 19672 710 19675 714
rect 19678 712 19680 718
rect 19934 715 19936 745
rect 19938 742 19948 745
rect 20108 743 20110 749
rect 20118 743 20124 749
rect 20137 746 20160 770
rect 20164 743 20170 749
rect 20112 742 20118 743
rect 19940 738 19948 742
rect 19940 735 19958 738
rect 19948 731 19958 735
rect 20110 731 20118 742
rect 20123 738 20124 742
rect 20156 739 20162 742
rect 20121 731 20123 738
rect 20157 737 20162 739
rect 20170 737 20176 743
rect 19908 714 19936 715
rect 19903 713 19936 714
rect 19940 713 19948 725
rect 19958 721 19964 731
rect 20110 721 20121 731
rect 20102 720 20121 721
rect 20102 712 20111 720
rect 19677 710 19678 711
rect 19675 707 19679 710
rect 19937 709 19940 711
rect 19911 708 19914 709
rect 19674 702 19679 707
rect 19899 706 19909 708
rect 19890 704 19899 706
rect 19669 696 19671 699
rect 19472 692 19538 693
rect 19478 691 19538 692
rect 19312 686 19339 688
rect 19388 686 19389 688
rect 19287 684 19319 686
rect 19277 683 19319 684
rect 19250 681 19319 683
rect 19232 679 19319 681
rect 19385 679 19388 684
rect 19041 678 19100 679
rect 19044 677 19079 678
rect 19205 677 19319 679
rect 19044 676 19076 677
rect 19078 676 19079 677
rect 19045 674 19057 676
rect 19059 675 19078 676
rect 19183 675 19205 677
rect 19211 676 19319 677
rect 19224 675 19228 676
rect 19059 671 19086 675
rect 19135 671 19183 675
rect 19059 670 19097 671
rect 19124 670 19167 671
rect 19059 664 19167 670
rect 19061 662 19071 664
rect 19224 662 19225 675
rect 19289 672 19291 675
rect 19382 673 19385 679
rect 18938 660 18939 662
rect 18720 658 18722 659
rect 18422 656 18424 657
rect 18642 656 18643 658
rect 18718 656 18720 658
rect 16346 652 16379 656
rect 16579 652 16582 656
rect 16326 651 16345 652
rect 16094 645 16095 651
rect 16049 640 16065 644
rect 16067 640 16083 644
rect 16363 640 16379 652
rect 16520 645 16530 652
rect 16574 646 16579 652
rect 16568 645 16574 646
rect 16530 644 16571 645
rect 16555 640 16571 644
rect 18074 640 18090 656
rect 18092 640 18108 656
rect 18275 653 18277 656
rect 18415 653 18421 656
rect 18644 653 18647 656
rect 18714 653 18718 656
rect 18277 651 18279 653
rect 18414 652 18415 653
rect 18712 652 18714 653
rect 18848 652 18960 660
rect 19052 658 19061 662
rect 19289 659 19292 672
rect 19421 666 19425 689
rect 19484 685 19538 691
rect 19622 688 19674 696
rect 19675 692 19679 702
rect 19832 693 19838 698
rect 19890 693 19896 698
rect 19832 692 19896 693
rect 19679 688 19681 690
rect 19480 679 19544 685
rect 19616 682 19681 688
rect 19838 686 19844 692
rect 19884 686 19890 692
rect 19902 690 19903 706
rect 19924 701 19936 709
rect 20115 707 20121 720
rect 20158 717 20162 737
rect 20114 706 20115 707
rect 20110 697 20114 706
rect 20162 697 20164 717
rect 20925 703 20947 722
rect 20896 697 20919 698
rect 20924 697 20947 703
rect 20110 693 20118 697
rect 20170 693 20176 697
rect 20110 691 20176 693
rect 20110 690 20114 691
rect 19903 686 19905 690
rect 19484 673 19492 679
rect 19532 673 19538 679
rect 19622 676 19628 682
rect 19668 676 19674 682
rect 19484 666 19491 673
rect 19624 672 19627 676
rect 19048 656 19052 658
rect 19225 656 19226 658
rect 19290 657 19292 659
rect 19288 656 19292 657
rect 19043 653 19048 656
rect 19226 653 19229 656
rect 19287 653 19288 656
rect 19322 654 19352 663
rect 19356 654 19369 660
rect 19421 659 19423 666
rect 19484 665 19492 666
rect 19038 652 19039 653
rect 19286 652 19287 653
rect 19319 652 19356 654
rect 19423 653 19425 659
rect 19481 656 19492 665
rect 19618 660 19627 672
rect 19680 672 19681 682
rect 19618 656 19624 660
rect 19680 656 19684 672
rect 19896 660 19905 686
rect 20104 674 20110 690
rect 20118 685 20124 691
rect 20164 685 20170 691
rect 20164 674 20167 685
rect 19480 653 19481 655
rect 19623 654 19624 656
rect 18412 651 18414 652
rect 18279 649 18355 651
rect 18407 649 18412 651
rect 18647 649 18651 652
rect 18710 650 18712 652
rect 18700 649 18710 650
rect 18362 648 18406 649
rect 18658 640 18674 649
rect 18675 648 18676 649
rect 18940 647 18942 651
rect 18960 647 19072 652
rect 18954 644 19072 647
rect 19170 644 19319 652
rect 18954 640 18970 644
rect 19072 641 19083 644
rect 19123 641 19170 644
rect 19083 640 19123 641
rect 19260 640 19276 644
rect 16068 639 16069 640
rect 19322 636 19352 652
rect 19460 640 19476 653
rect 19623 644 19633 654
rect 19896 652 19909 660
rect 19964 656 19980 672
rect 20102 665 20111 674
rect 20164 667 20176 674
rect 20167 665 20176 667
rect 20104 656 20105 665
rect 20111 656 20120 665
rect 20158 656 20172 665
rect 19931 652 19964 656
rect 20164 652 20167 656
rect 19911 651 19930 652
rect 19679 645 19680 651
rect 19634 640 19650 644
rect 19652 640 19668 644
rect 19948 640 19964 652
rect 20105 645 20115 652
rect 20159 646 20164 652
rect 20153 645 20159 646
rect 20115 644 20156 645
rect 20140 640 20156 644
rect 19653 639 19654 640
rect 6529 623 6556 629
rect 6557 623 6584 624
rect 10114 623 10141 629
rect 10142 623 10169 624
rect 13699 623 13726 629
rect 13727 623 13754 624
rect 17284 623 17311 629
rect 17312 623 17339 624
rect 20869 623 20896 629
rect 20897 623 20924 624
rect 7100 481 7101 487
rect 10685 481 10686 487
rect 14270 481 14271 487
rect 17855 481 17856 487
rect 21440 481 21441 487
rect 7066 441 7101 475
rect 7112 463 7113 475
rect 7112 441 7113 453
rect 10651 441 10686 475
rect 10697 463 10698 475
rect 10697 441 10698 453
rect 14236 441 14271 475
rect 14282 463 14283 475
rect 14282 441 14283 453
rect 17821 441 17856 475
rect 17867 463 17868 475
rect 17867 441 17868 453
rect 21406 441 21441 475
rect 21452 463 21453 475
rect 21452 441 21453 453
rect 6309 429 6310 440
rect 6499 429 6500 440
rect 6585 429 6586 440
rect 6858 429 6859 440
rect 7055 429 7056 440
rect 7089 429 7101 435
rect 9894 429 9895 440
rect 10084 429 10085 440
rect 10170 429 10171 440
rect 10443 429 10444 440
rect 10640 429 10641 440
rect 10674 429 10686 435
rect 13479 429 13480 440
rect 13669 429 13670 440
rect 13755 429 13756 440
rect 14028 429 14029 440
rect 14225 429 14226 440
rect 14259 429 14271 435
rect 17064 429 17065 440
rect 17254 429 17255 440
rect 17340 429 17341 440
rect 17613 429 17614 440
rect 17810 429 17811 440
rect 17844 429 17856 435
rect 20649 429 20650 440
rect 20839 429 20840 440
rect 20925 429 20926 440
rect 21198 429 21199 440
rect 21395 429 21396 440
rect 21429 429 21441 435
rect 6320 389 6321 429
rect 6510 389 6511 429
rect 6596 389 6597 429
rect 6869 389 6870 429
rect 7066 389 7067 429
rect 9905 389 9906 429
rect 10095 389 10096 429
rect 10181 389 10182 429
rect 10454 389 10455 429
rect 10651 389 10652 429
rect 13490 389 13491 429
rect 13680 389 13681 429
rect 13766 389 13767 429
rect 14039 389 14040 429
rect 14236 389 14237 429
rect 17075 389 17076 429
rect 17265 389 17266 429
rect 17351 389 17352 429
rect 17624 389 17625 429
rect 17821 389 17822 429
rect 20660 389 20661 429
rect 20850 389 20851 429
rect 20936 389 20937 429
rect 21209 389 21210 429
rect 21406 389 21407 429
<< nwell >>
rect 2996 1436 6195 1778
rect 8870 1676 8904 1710
rect 12455 1676 12489 1710
rect 16040 1676 16074 1710
rect 19625 1676 19659 1710
rect 2996 1116 21516 1436
rect 2996 1078 6195 1116
rect 2996 850 4518 1078
<< ndiff >>
rect 7067 441 7101 475
rect 10652 441 10686 475
rect 14237 441 14271 475
rect 17822 441 17856 475
rect 21407 441 21441 475
<< pdiff >>
rect 5285 1676 5319 1710
rect 8870 1676 8904 1710
rect 12455 1676 12489 1710
rect 16040 1676 16074 1710
rect 19625 1676 19659 1710
<< locali >>
rect 6 2289 21517 2522
rect 7 2202 21517 2289
rect 3439 1436 3473 1518
rect 1 1116 21516 1436
rect 3665 487 6047 548
rect 0 0 21516 320
<< metal1 >>
rect 7 2202 21517 2522
rect 21437 2012 21442 2045
rect 21401 2006 21471 2012
rect 3335 1892 3341 1950
rect 3399 1892 3405 1950
rect 21401 1948 21407 2006
rect 21465 1948 21471 2006
rect 21401 1942 21471 1948
rect 7066 1883 7136 1889
rect 5669 1872 5739 1878
rect 5669 1814 5675 1872
rect 5733 1814 5739 1872
rect 7066 1825 7072 1883
rect 7130 1825 7136 1883
rect 10650 1883 10721 1890
rect 7066 1819 7136 1825
rect 9260 1874 9330 1880
rect 5669 1808 5739 1814
rect 9260 1816 9266 1874
rect 9324 1816 9330 1874
rect 10650 1825 10657 1883
rect 10715 1825 10721 1883
rect 14227 1883 14297 1889
rect 10650 1819 10721 1825
rect 12846 1874 12916 1880
rect 9260 1810 9330 1816
rect 12846 1816 12852 1874
rect 12910 1816 12916 1874
rect 14227 1825 14233 1883
rect 14291 1825 14297 1883
rect 17812 1883 17882 1889
rect 14227 1819 14297 1825
rect 16420 1874 16490 1880
rect 12846 1810 12916 1816
rect 16420 1816 16426 1874
rect 16484 1816 16490 1874
rect 17812 1825 17818 1883
rect 17876 1825 17882 1883
rect 17812 1819 17882 1825
rect 20061 1874 20131 1880
rect 16420 1810 16490 1816
rect 20061 1816 20067 1874
rect 20125 1816 20131 1874
rect 20061 1810 20131 1816
rect 3260 1744 3266 1802
rect 3324 1744 3330 1802
rect 3067 1670 3125 1716
rect 5285 1676 5319 1710
rect 8870 1676 8904 1710
rect 12455 1676 12489 1710
rect 16040 1676 16074 1710
rect 19625 1676 19659 1710
rect 1 1116 21516 1436
rect 3665 492 6047 548
rect 7067 441 7101 475
rect 10652 441 10686 475
rect 14237 441 14271 475
rect 17822 441 17856 475
rect 21407 441 21441 475
rect 0 0 21516 320
<< via1 >>
rect 3341 1892 3399 1950
rect 21407 1948 21465 2006
rect 5675 1814 5733 1872
rect 7072 1825 7130 1883
rect 9266 1816 9324 1874
rect 10657 1825 10715 1883
rect 12852 1816 12910 1874
rect 14233 1825 14291 1883
rect 16426 1816 16484 1874
rect 17818 1825 17876 1883
rect 20067 1816 20125 1874
rect 3266 1744 3324 1802
<< metal2 >>
rect 3278 2167 21441 2201
rect 3278 1808 3312 2167
rect 21407 2012 21441 2167
rect 21401 2006 21471 2012
rect 3341 1950 3399 1956
rect 21401 1948 21407 2006
rect 21465 1948 21471 2006
rect 21401 1942 21471 1948
rect 3399 1898 3603 1932
rect 3341 1886 3399 1892
rect 3569 1858 3603 1898
rect 7066 1883 7136 1889
rect 5669 1872 5739 1878
rect 5669 1858 5675 1872
rect 3569 1824 5675 1858
rect 5669 1814 5675 1824
rect 5733 1814 5739 1872
rect 7066 1825 7072 1883
rect 7130 1865 7136 1883
rect 10651 1883 10721 1889
rect 9260 1874 9330 1880
rect 9260 1865 9266 1874
rect 7130 1825 9266 1865
rect 7066 1819 7136 1825
rect 5669 1808 5739 1814
rect 9260 1816 9266 1825
rect 9324 1816 9330 1874
rect 10651 1825 10657 1883
rect 10715 1865 10721 1883
rect 14227 1883 14297 1889
rect 12846 1874 12916 1880
rect 12846 1865 12852 1874
rect 10715 1825 12852 1865
rect 10651 1819 10721 1825
rect 9260 1810 9330 1816
rect 12846 1816 12852 1825
rect 12910 1816 12916 1874
rect 14227 1825 14233 1883
rect 14291 1865 14297 1883
rect 17812 1883 17882 1889
rect 16420 1874 16490 1880
rect 16420 1865 16426 1874
rect 14291 1825 16426 1865
rect 14227 1819 14297 1825
rect 12846 1810 12916 1816
rect 16420 1816 16426 1825
rect 16484 1816 16490 1874
rect 17812 1825 17818 1883
rect 17876 1865 17882 1883
rect 20061 1874 20131 1880
rect 20061 1865 20067 1874
rect 17876 1825 20067 1865
rect 17812 1819 17882 1825
rect 16420 1810 16490 1816
rect 20061 1816 20067 1825
rect 20125 1816 20131 1874
rect 20061 1810 20131 1816
rect 3266 1802 3324 1808
rect 3266 1738 3324 1744
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_0
timestamp 1698882961
transform 1 0 3042 0 -1 2263
box -8 0 552 902
use sky130_osu_single_mpr2at_8_b0r2  sky130_osu_single_mpr2at_8_b0r2_0
timestamp 1708010873
transform 1 0 17930 0 1 0
box 0 0 3587 2522
use sky130_osu_single_mpr2at_8_b0r2  sky130_osu_single_mpr2at_8_b0r2_1
timestamp 1708010873
transform 1 0 3590 0 1 0
box 0 0 3587 2522
use sky130_osu_single_mpr2at_8_b0r2  sky130_osu_single_mpr2at_8_b0r2_2
timestamp 1708010873
transform 1 0 7175 0 1 0
box 0 0 3587 2522
use sky130_osu_single_mpr2at_8_b0r2  sky130_osu_single_mpr2at_8_b0r2_3
timestamp 1708010873
transform 1 0 10760 0 1 0
box 0 0 3587 2522
use sky130_osu_single_mpr2at_8_b0r2  sky130_osu_single_mpr2at_8_b0r2_4
timestamp 1708010873
transform 1 0 14345 0 1 0
box 0 0 3587 2522
<< labels >>
flabel metal1 s 3067 1670 3125 1716 0 FreeSans 100 0 0 0 start
port 13 nsew signal input
flabel metal1 s 5285 1676 5319 1710 0 FreeSans 100 0 0 0 s1
port 1 nsew signal input
flabel metal1 s 8870 1676 8904 1710 0 FreeSans 100 0 0 0 s2
port 2 nsew signal input
flabel metal1 s 12455 1676 12489 1710 0 FreeSans 100 0 0 0 s3
port 3 nsew signal input
flabel metal1 s 16040 1676 16074 1710 0 FreeSans 100 0 0 0 s4
port 4 nsew signal input
flabel metal1 s 19625 1676 19659 1710 0 FreeSans 100 0 0 0 s5
port 5 nsew signal input
flabel metal1 s 7067 441 7101 475 0 FreeSans 100 0 0 0 X1_Y1
port 6 nsew signal output
flabel metal1 s 10652 441 10686 475 0 FreeSans 100 0 0 0 X2_Y1
port 7 nsew signal output
flabel metal1 s 14237 441 14271 475 0 FreeSans 100 0 0 0 X3_Y1
port 8 nsew signal output
flabel metal1 s 17822 441 17856 475 0 FreeSans 100 0 0 0 X4_Y1
port 9 nsew signal output
flabel metal1 s 21407 441 21441 475 0 FreeSans 100 0 0 0 X5_Y1
port 10 nsew signal output
flabel metal1 s 7 2202 21517 2522 0 FreeSans 100 0 0 0 vssd1
port 14 nsew ground bidirectional
flabel metal1 s 1 1116 21516 1436 0 FreeSans 100 0 0 0 vccd1
port 15 nsew power bidirectional
flabel metal1 s 0 0 21516 320 0 FreeSans 100 0 0 0 vssd1
port 14 nsew ground bidirectional
<< end >>
