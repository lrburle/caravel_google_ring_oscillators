magic
tech sky130A
magscale 1 2
timestamp 1713888962
<< nwell >>
rect 3000 1406 5497 1748
rect 8018 1635 8070 1693
rect 11283 1635 11335 1693
rect 14548 1635 14600 1693
rect 17813 1635 17865 1693
rect 3000 1086 19885 1406
rect 3000 1018 5497 1086
rect 3000 820 4486 1018
rect 6705 986 6763 1044
rect 9970 986 10028 1044
rect 13235 986 13293 1044
rect 16500 986 16558 1044
rect 19765 986 19823 1044
<< ndiff >>
rect 6716 442 6751 476
rect 9981 442 10016 476
rect 13246 442 13281 476
rect 16511 442 16546 476
rect 19776 442 19811 476
rect 6719 441 6750 442
rect 9984 441 10015 442
rect 13249 441 13280 442
rect 16514 441 16545 442
rect 19779 441 19810 442
<< pdiff >>
rect 3046 1647 3080 1681
rect 4753 1635 4805 1693
rect 8018 1635 8070 1693
rect 11283 1635 11335 1693
rect 14548 1635 14600 1693
rect 17813 1635 17865 1693
<< locali >>
rect 10 2172 19886 2492
rect 3407 1406 3441 1475
rect 1 1086 19885 1406
rect 0 0 19885 320
<< viali >>
rect 3040 1635 3086 1681
rect 6717 442 6751 476
rect 9982 442 10016 476
rect 13247 442 13281 476
rect 16512 442 16546 476
rect 19777 442 19811 476
<< metal1 >>
rect 10 2172 19886 2492
rect 19805 2008 19812 2011
rect 19771 2001 19824 2008
rect 19771 1982 19836 2001
rect 19771 1976 19841 1982
rect 3303 1863 3309 1921
rect 3367 1863 3373 1921
rect 19771 1918 19777 1976
rect 19835 1918 19841 1976
rect 19771 1912 19841 1918
rect 6715 1852 6785 1858
rect 5318 1842 5388 1848
rect 5318 1784 5324 1842
rect 5382 1784 5388 1842
rect 5318 1778 5388 1784
rect 6715 1794 6721 1852
rect 6779 1794 6785 1852
rect 9979 1853 10050 1860
rect 6715 1788 6785 1794
rect 8416 1843 8486 1849
rect 3228 1714 3234 1772
rect 3292 1714 3298 1772
rect 6715 1767 6775 1788
rect 8416 1785 8422 1843
rect 8480 1785 8486 1843
rect 8416 1779 8486 1785
rect 9979 1795 9986 1853
rect 10044 1795 10050 1853
rect 13236 1852 13306 1858
rect 9979 1789 10050 1795
rect 11681 1844 11751 1850
rect 9979 1768 10040 1789
rect 11681 1786 11687 1844
rect 11745 1786 11751 1844
rect 11681 1780 11751 1786
rect 13236 1794 13242 1852
rect 13300 1794 13306 1852
rect 16501 1852 16571 1858
rect 13236 1788 13306 1794
rect 14946 1843 15016 1849
rect 13236 1768 13305 1788
rect 14946 1785 14952 1843
rect 15010 1785 15016 1843
rect 14946 1779 15016 1785
rect 16501 1794 16507 1852
rect 16565 1794 16571 1852
rect 16501 1788 16571 1794
rect 18212 1843 18282 1849
rect 16501 1769 16570 1788
rect 18212 1785 18218 1843
rect 18276 1785 18282 1843
rect 18212 1779 18282 1785
rect 3035 1681 3093 1686
rect 3035 1640 3040 1681
rect 3086 1640 3093 1681
rect 1 1086 19885 1406
rect 6716 441 6750 442
rect 9981 441 10015 442
rect 13246 441 13280 442
rect 16511 441 16545 442
rect 19776 441 19810 442
rect 0 0 19885 320
<< via1 >>
rect 3309 1863 3367 1921
rect 19777 1918 19835 1976
rect 5324 1784 5382 1842
rect 6721 1794 6779 1852
rect 3234 1714 3292 1772
rect 8422 1785 8480 1843
rect 9986 1795 10044 1853
rect 11687 1786 11745 1844
rect 13242 1794 13300 1852
rect 14952 1785 15010 1843
rect 16507 1794 16565 1852
rect 18218 1785 18276 1843
rect 4753 1635 4805 1693
rect 8018 1635 8070 1693
rect 11283 1635 11335 1693
rect 14548 1635 14600 1693
rect 17813 1635 17865 1693
<< metal2 >>
rect 3246 2137 19811 2171
rect 3246 1778 3280 2137
rect 19777 1982 19811 2137
rect 19771 1976 19841 1982
rect 3309 1921 3367 1927
rect 19771 1918 19777 1976
rect 19835 1918 19841 1976
rect 19771 1912 19841 1918
rect 3367 1902 3384 1903
rect 3367 1867 3566 1902
rect 3309 1857 3367 1863
rect 3531 1829 3566 1867
rect 6715 1852 6785 1858
rect 5318 1842 5388 1848
rect 5318 1829 5324 1842
rect 3531 1794 5324 1829
rect 5318 1784 5324 1794
rect 5382 1784 5388 1842
rect 6715 1794 6721 1852
rect 6779 1834 6785 1852
rect 9980 1853 10050 1859
rect 8416 1843 8486 1849
rect 8416 1834 8422 1843
rect 6779 1794 8422 1834
rect 6715 1788 6785 1794
rect 5318 1778 5388 1784
rect 8416 1785 8422 1794
rect 8480 1785 8486 1843
rect 9980 1795 9986 1853
rect 10044 1835 10050 1853
rect 13236 1852 13306 1858
rect 11681 1844 11751 1850
rect 11681 1835 11687 1844
rect 10044 1795 11687 1835
rect 9980 1789 10050 1795
rect 8416 1779 8486 1785
rect 11681 1786 11687 1795
rect 11745 1786 11751 1844
rect 13236 1794 13242 1852
rect 13300 1834 13306 1852
rect 16501 1852 16571 1858
rect 14946 1843 15016 1849
rect 14946 1834 14952 1843
rect 13300 1794 14952 1834
rect 13236 1788 13306 1794
rect 11681 1780 11751 1786
rect 14946 1785 14952 1794
rect 15010 1785 15016 1843
rect 16501 1794 16507 1852
rect 16565 1834 16571 1852
rect 18212 1843 18282 1849
rect 18212 1834 18218 1843
rect 16565 1794 18218 1834
rect 16501 1788 16571 1794
rect 14946 1779 15016 1785
rect 18212 1785 18218 1794
rect 18276 1785 18282 1843
rect 18212 1779 18282 1785
rect 3234 1772 3292 1778
rect 3234 1708 3292 1714
<< via2 >>
rect 4753 1635 4805 1693
rect 8018 1635 8070 1693
rect 11283 1635 11335 1693
rect 14548 1635 14600 1693
rect 17813 1635 17865 1693
<< metal3 >>
rect 4747 1693 4814 2492
rect 8012 1693 8079 2492
rect 11277 1693 11344 2492
rect 14542 1693 14609 2492
rect 17807 1693 17874 2492
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_0
timestamp 1713481735
transform 1 0 3010 0 -1 2233
box -10 0 552 902
use sky130_osu_single_mpr2ea_8_b0r1  sky130_osu_single_mpr2ea_8_b0r1_0
timestamp 1713888380
transform 1 0 16618 0 1 0
box 0 0 3268 2492
use sky130_osu_single_mpr2ea_8_b0r1  sky130_osu_single_mpr2ea_8_b0r1_1
timestamp 1713888380
transform 1 0 3558 0 1 0
box 0 0 3268 2492
use sky130_osu_single_mpr2ea_8_b0r1  sky130_osu_single_mpr2ea_8_b0r1_2
timestamp 1713888380
transform 1 0 6823 0 1 0
box 0 0 3268 2492
use sky130_osu_single_mpr2ea_8_b0r1  sky130_osu_single_mpr2ea_8_b0r1_3
timestamp 1713888380
transform 1 0 10088 0 1 0
box 0 0 3268 2492
use sky130_osu_single_mpr2ea_8_b0r1  sky130_osu_single_mpr2ea_8_b0r1_4
timestamp 1713888380
transform 1 0 13353 0 1 0
box 0 0 3268 2492
<< labels >>
flabel metal1 s 3035 1640 3093 1686 0 FreeSans 100 0 0 0 start
port 13 nsew signal input
flabel metal1 s 10 2172 19886 2492 0 FreeSans 100 0 0 0 vssd1
port 14 nsew ground bidirectional
flabel metal1 s 1 1086 19885 1406 0 FreeSans 100 0 0 0 vccd1
port 15 nsew power bidirectional
flabel metal1 s 0 0 19885 320 0 FreeSans 100 0 0 0 vssd1
port 14 nsew ground bidirectional
flabel via2 s 8027 1647 8061 1681 0 FreeSans 100 0 0 0 s2
port 2 nw signal input
flabel via2 s 4762 1647 4796 1681 0 FreeSans 100 0 0 0 s1
port 1 nw signal input
flabel via2 s 11292 1647 11326 1681 0 FreeSans 100 0 0 0 s3
port 3 nw signal input
flabel via2 s 14557 1647 14591 1681 0 FreeSans 100 0 0 0 s4
port 4 nw signal input
flabel via2 s 17822 1647 17856 1681 0 FreeSans 100 0 0 0 s5
port 5 nw signal input
flabel viali s 6717 442 6751 476 0 FreeSans 100 0 0 0 X1_Y1
port 6 se signal output
flabel viali s 9982 442 10016 476 0 FreeSans 100 0 0 0 X2_Y1
port 7 se signal output
flabel viali s 13247 442 13281 476 0 FreeSans 100 0 0 0 X3_Y1
port 8 se signal output
flabel viali s 16512 442 16546 476 0 FreeSans 100 0 0 0 X4_Y1
port 9 se signal output
flabel viali s 19777 442 19811 476 0 FreeSans 100 0 0 0 X5_Y1
port 10 se signal output
<< end >>
