VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sky130_osu_ring_oscillator_mpr2aa_8_b0r1
  CLASS BLOCK ;
  ORIGIN 0.005 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2aa_8_b0r1 ;
  SIZE 81.785 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 18.11 0.915 18.28 1.085 ;
        RECT 18.105 0.91 18.275 1.08 ;
        RECT 18.105 2.39 18.275 2.56 ;
      LAYER li1 ;
        RECT 18.11 0.915 18.28 1.085 ;
        RECT 18.105 0.57 18.275 1.08 ;
        RECT 18.105 2.39 18.275 3.86 ;
      LAYER met1 ;
        RECT 18.045 2.36 18.335 2.59 ;
        RECT 18.045 0.88 18.335 1.11 ;
        RECT 18.105 0.88 18.275 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 33.89 0.915 34.06 1.085 ;
        RECT 33.885 0.91 34.055 1.08 ;
        RECT 33.885 2.39 34.055 2.56 ;
      LAYER li1 ;
        RECT 33.89 0.915 34.06 1.085 ;
        RECT 33.885 0.57 34.055 1.08 ;
        RECT 33.885 2.39 34.055 3.86 ;
      LAYER met1 ;
        RECT 33.825 2.36 34.115 2.59 ;
        RECT 33.825 0.88 34.115 1.11 ;
        RECT 33.885 0.88 34.055 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 49.665 0.915 49.835 1.085 ;
        RECT 49.66 0.91 49.83 1.08 ;
        RECT 49.66 2.39 49.83 2.56 ;
      LAYER li1 ;
        RECT 49.665 0.915 49.835 1.085 ;
        RECT 49.66 0.57 49.83 1.08 ;
        RECT 49.66 2.39 49.83 3.86 ;
      LAYER met1 ;
        RECT 49.6 2.36 49.89 2.59 ;
        RECT 49.6 0.88 49.89 1.11 ;
        RECT 49.66 0.88 49.83 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 65.45 0.915 65.62 1.085 ;
        RECT 65.445 0.91 65.615 1.08 ;
        RECT 65.445 2.39 65.615 2.56 ;
      LAYER li1 ;
        RECT 65.45 0.915 65.62 1.085 ;
        RECT 65.445 0.57 65.615 1.08 ;
        RECT 65.445 2.39 65.615 3.86 ;
      LAYER met1 ;
        RECT 65.385 2.36 65.675 2.59 ;
        RECT 65.385 0.88 65.675 1.11 ;
        RECT 65.445 0.88 65.615 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 81.235 0.915 81.405 1.085 ;
        RECT 81.23 0.91 81.4 1.08 ;
        RECT 81.23 2.39 81.4 2.56 ;
      LAYER li1 ;
        RECT 81.235 0.915 81.405 1.085 ;
        RECT 81.23 0.57 81.4 1.08 ;
        RECT 81.23 2.39 81.4 3.86 ;
      LAYER met1 ;
        RECT 81.17 2.36 81.46 2.59 ;
        RECT 81.17 0.88 81.46 1.11 ;
        RECT 81.23 0.88 81.4 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 13.87 5.855 14.22 6.205 ;
        RECT 13.865 2.705 14.215 3.055 ;
        RECT 13.94 2.705 14.115 6.205 ;
      LAYER li1 ;
        RECT 13.955 1.66 14.125 2.935 ;
        RECT 13.955 5.945 14.125 7.22 ;
        RECT 9.175 5.945 9.345 7.22 ;
      LAYER met1 ;
        RECT 13.865 2.765 14.355 2.935 ;
        RECT 13.865 2.705 14.215 3.055 ;
        RECT 9.115 5.945 14.355 6.115 ;
        RECT 13.87 5.855 14.22 6.205 ;
        RECT 9.115 5.915 9.405 6.145 ;
      LAYER via1 ;
        RECT 13.965 2.805 14.115 2.955 ;
        RECT 13.97 5.955 14.12 6.105 ;
      LAYER mcon ;
        RECT 9.175 5.945 9.345 6.115 ;
        RECT 13.955 5.945 14.125 6.115 ;
        RECT 13.955 2.765 14.125 2.935 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 29.65 5.855 30 6.205 ;
        RECT 29.645 2.705 29.995 3.055 ;
        RECT 29.72 2.705 29.895 6.205 ;
      LAYER li1 ;
        RECT 29.735 1.66 29.905 2.935 ;
        RECT 29.735 5.945 29.905 7.22 ;
        RECT 24.955 5.945 25.125 7.22 ;
      LAYER met1 ;
        RECT 29.645 2.765 30.135 2.935 ;
        RECT 29.645 2.705 29.995 3.055 ;
        RECT 24.895 5.945 30.135 6.115 ;
        RECT 29.65 5.855 30 6.205 ;
        RECT 24.895 5.915 25.185 6.145 ;
      LAYER via1 ;
        RECT 29.745 2.805 29.895 2.955 ;
        RECT 29.75 5.955 29.9 6.105 ;
      LAYER mcon ;
        RECT 24.955 5.945 25.125 6.115 ;
        RECT 29.735 5.945 29.905 6.115 ;
        RECT 29.735 2.765 29.905 2.935 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 45.425 5.855 45.775 6.205 ;
        RECT 45.42 2.705 45.77 3.055 ;
        RECT 45.495 2.705 45.67 6.205 ;
      LAYER li1 ;
        RECT 45.51 1.66 45.68 2.935 ;
        RECT 45.51 5.945 45.68 7.22 ;
        RECT 40.73 5.945 40.9 7.22 ;
      LAYER met1 ;
        RECT 45.42 2.765 45.91 2.935 ;
        RECT 45.42 2.705 45.77 3.055 ;
        RECT 40.67 5.945 45.91 6.115 ;
        RECT 45.425 5.855 45.775 6.205 ;
        RECT 40.67 5.915 40.96 6.145 ;
      LAYER via1 ;
        RECT 45.52 2.805 45.67 2.955 ;
        RECT 45.525 5.955 45.675 6.105 ;
      LAYER mcon ;
        RECT 40.73 5.945 40.9 6.115 ;
        RECT 45.51 5.945 45.68 6.115 ;
        RECT 45.51 2.765 45.68 2.935 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 61.21 5.855 61.56 6.205 ;
        RECT 61.205 2.705 61.555 3.055 ;
        RECT 61.28 2.705 61.455 6.205 ;
      LAYER li1 ;
        RECT 61.295 1.66 61.465 2.935 ;
        RECT 61.295 5.945 61.465 7.22 ;
        RECT 56.515 5.945 56.685 7.22 ;
      LAYER met1 ;
        RECT 61.205 2.765 61.695 2.935 ;
        RECT 61.205 2.705 61.555 3.055 ;
        RECT 56.455 5.945 61.695 6.115 ;
        RECT 61.21 5.855 61.56 6.205 ;
        RECT 56.455 5.915 56.745 6.145 ;
      LAYER via1 ;
        RECT 61.305 2.805 61.455 2.955 ;
        RECT 61.31 5.955 61.46 6.105 ;
      LAYER mcon ;
        RECT 56.515 5.945 56.685 6.115 ;
        RECT 61.295 5.945 61.465 6.115 ;
        RECT 61.295 2.765 61.465 2.935 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 76.995 5.855 77.345 6.205 ;
        RECT 76.99 2.705 77.34 3.055 ;
        RECT 77.065 2.705 77.24 6.205 ;
      LAYER li1 ;
        RECT 77.08 1.66 77.25 2.935 ;
        RECT 77.08 5.945 77.25 7.22 ;
        RECT 72.3 5.945 72.47 7.22 ;
      LAYER met1 ;
        RECT 76.99 2.765 77.48 2.935 ;
        RECT 76.99 2.705 77.34 3.055 ;
        RECT 72.24 5.945 77.48 6.115 ;
        RECT 76.995 5.855 77.345 6.205 ;
        RECT 72.24 5.915 72.53 6.145 ;
      LAYER via1 ;
        RECT 77.09 2.805 77.24 2.955 ;
        RECT 77.095 5.955 77.245 6.105 ;
      LAYER mcon ;
        RECT 72.3 5.945 72.47 6.115 ;
        RECT 77.08 5.945 77.25 6.115 ;
        RECT 77.08 2.765 77.25 2.935 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 0.24 5.945 0.41 7.22 ;
      LAYER met1 ;
        RECT 0.18 5.945 0.64 6.115 ;
        RECT 0.18 5.915 0.47 6.145 ;
      LAYER mcon ;
        RECT 0.24 5.945 0.41 6.115 ;
    END
  END start
  OBS
    LAYER met3 ;
      RECT 73.57 7.04 73.94 7.41 ;
      RECT 73.61 6.72 73.945 7.085 ;
      RECT 73.61 6.72 73.995 7.03 ;
      RECT 73.61 6.72 76.4 7.025 ;
      RECT 76.095 2.85 76.4 7.025 ;
      RECT 76.06 2.85 76.43 3.22 ;
      RECT 75.32 0.815 75.625 4.02 ;
      RECT 75.07 2.975 75.625 3.705 ;
      RECT 75.28 0.815 75.65 1.185 ;
      RECT 71.43 1.85 71.76 2.745 ;
      RECT 70.55 2.015 70.88 2.745 ;
      RECT 71.425 1.85 71.795 2.65 ;
      RECT 74.59 1.85 74.92 2.58 ;
      RECT 74.55 1.735 74.73 2.385 ;
      RECT 70.56 1.85 74.92 2.22 ;
      RECT 71.05 3.535 71.38 3.865 ;
      RECT 69.845 3.55 71.38 3.85 ;
      RECT 69.845 2.43 70.145 3.85 ;
      RECT 69.59 2.415 69.92 2.745 ;
      RECT 57.785 7.04 58.155 7.41 ;
      RECT 57.825 6.72 58.16 7.085 ;
      RECT 57.825 6.72 58.21 7.03 ;
      RECT 57.825 6.72 60.615 7.025 ;
      RECT 60.31 2.85 60.615 7.025 ;
      RECT 60.275 2.85 60.645 3.22 ;
      RECT 59.535 0.815 59.84 4.02 ;
      RECT 59.285 2.975 59.84 3.705 ;
      RECT 59.495 0.815 59.865 1.185 ;
      RECT 55.645 1.85 55.975 2.745 ;
      RECT 54.765 2.015 55.095 2.745 ;
      RECT 55.64 1.85 56.01 2.65 ;
      RECT 58.805 1.85 59.135 2.58 ;
      RECT 58.765 1.735 58.945 2.385 ;
      RECT 54.775 1.85 59.135 2.22 ;
      RECT 55.265 3.535 55.595 3.865 ;
      RECT 54.06 3.55 55.595 3.85 ;
      RECT 54.06 2.43 54.36 3.85 ;
      RECT 53.805 2.415 54.135 2.745 ;
      RECT 42 7.04 42.37 7.41 ;
      RECT 42.04 6.72 42.375 7.085 ;
      RECT 42.04 6.72 42.425 7.03 ;
      RECT 42.04 6.72 44.83 7.025 ;
      RECT 44.525 2.85 44.83 7.025 ;
      RECT 44.49 2.85 44.86 3.22 ;
      RECT 43.75 0.815 44.055 4.02 ;
      RECT 43.5 2.975 44.055 3.705 ;
      RECT 43.71 0.815 44.08 1.185 ;
      RECT 39.86 1.85 40.19 2.745 ;
      RECT 38.98 2.015 39.31 2.745 ;
      RECT 39.855 1.85 40.225 2.65 ;
      RECT 43.02 1.85 43.35 2.58 ;
      RECT 42.98 1.735 43.16 2.385 ;
      RECT 38.99 1.85 43.35 2.22 ;
      RECT 39.48 3.535 39.81 3.865 ;
      RECT 38.275 3.55 39.81 3.85 ;
      RECT 38.275 2.43 38.575 3.85 ;
      RECT 38.02 2.415 38.35 2.745 ;
      RECT 26.225 7.04 26.595 7.41 ;
      RECT 26.265 6.72 26.6 7.085 ;
      RECT 26.265 6.72 26.65 7.03 ;
      RECT 26.265 6.72 29.055 7.025 ;
      RECT 28.75 2.85 29.055 7.025 ;
      RECT 28.715 2.85 29.085 3.22 ;
      RECT 27.975 0.815 28.28 4.02 ;
      RECT 27.725 2.975 28.28 3.705 ;
      RECT 27.935 0.815 28.305 1.185 ;
      RECT 24.085 1.85 24.415 2.745 ;
      RECT 23.205 2.015 23.535 2.745 ;
      RECT 24.08 1.85 24.45 2.65 ;
      RECT 27.245 1.85 27.575 2.58 ;
      RECT 27.205 1.735 27.385 2.385 ;
      RECT 23.215 1.85 27.575 2.22 ;
      RECT 23.705 3.535 24.035 3.865 ;
      RECT 22.5 3.55 24.035 3.85 ;
      RECT 22.5 2.43 22.8 3.85 ;
      RECT 22.245 2.415 22.575 2.745 ;
      RECT 10.445 7.04 10.815 7.41 ;
      RECT 10.485 6.72 10.82 7.085 ;
      RECT 10.485 6.72 10.87 7.03 ;
      RECT 10.485 6.72 13.275 7.025 ;
      RECT 12.97 2.85 13.275 7.025 ;
      RECT 12.935 2.85 13.305 3.22 ;
      RECT 12.195 0.815 12.5 4.02 ;
      RECT 11.945 2.975 12.5 3.705 ;
      RECT 12.155 0.815 12.525 1.185 ;
      RECT 8.305 1.85 8.635 2.745 ;
      RECT 7.425 2.015 7.755 2.745 ;
      RECT 8.3 1.85 8.67 2.65 ;
      RECT 11.465 1.85 11.795 2.58 ;
      RECT 11.425 1.735 11.605 2.385 ;
      RECT 7.435 1.85 11.795 2.22 ;
      RECT 7.925 3.535 8.255 3.865 ;
      RECT 6.72 3.55 8.255 3.85 ;
      RECT 6.72 2.43 7.02 3.85 ;
      RECT 6.465 2.415 6.795 2.745 ;
      RECT 0.25 8.5 0.865 8.88 ;
      RECT 0.02 8.51 0.865 8.87 ;
      RECT 0.055 8.5 0.865 8.87 ;
      RECT 72.99 2.575 73.32 3.305 ;
      RECT 68.87 2.415 69.2 3.145 ;
      RECT 67.87 1.855 68.2 2.585 ;
      RECT 66.43 2.575 66.76 3.305 ;
      RECT 57.205 2.575 57.535 3.305 ;
      RECT 53.085 2.415 53.415 3.145 ;
      RECT 52.085 1.855 52.415 2.585 ;
      RECT 50.645 2.575 50.975 3.305 ;
      RECT 41.42 2.575 41.75 3.305 ;
      RECT 37.3 2.415 37.63 3.145 ;
      RECT 36.3 1.855 36.63 2.585 ;
      RECT 34.86 2.575 35.19 3.305 ;
      RECT 25.645 2.575 25.975 3.305 ;
      RECT 21.525 2.415 21.855 3.145 ;
      RECT 20.525 1.855 20.855 2.585 ;
      RECT 19.085 2.575 19.415 3.305 ;
      RECT 9.865 2.575 10.195 3.305 ;
      RECT 5.745 2.415 6.075 3.145 ;
      RECT 4.745 1.855 5.075 2.585 ;
      RECT 3.305 2.575 3.635 3.305 ;
      RECT 0.64 4.26 1.45 4.64 ;
      RECT 0.585 0 1.395 0.38 ;
    LAYER via2 ;
      RECT 76.145 2.935 76.345 3.135 ;
      RECT 75.365 0.9 75.565 1.1 ;
      RECT 75.135 3.04 75.335 3.24 ;
      RECT 74.655 2.315 74.855 2.515 ;
      RECT 73.655 7.125 73.855 7.325 ;
      RECT 73.055 3.04 73.255 3.24 ;
      RECT 71.495 2.48 71.695 2.68 ;
      RECT 71.115 3.6 71.315 3.8 ;
      RECT 70.615 2.48 70.815 2.68 ;
      RECT 69.655 2.48 69.855 2.68 ;
      RECT 68.935 2.48 69.135 2.68 ;
      RECT 67.935 1.92 68.135 2.12 ;
      RECT 66.495 3.04 66.695 3.24 ;
      RECT 60.36 2.935 60.56 3.135 ;
      RECT 59.58 0.9 59.78 1.1 ;
      RECT 59.35 3.04 59.55 3.24 ;
      RECT 58.87 2.315 59.07 2.515 ;
      RECT 57.87 7.125 58.07 7.325 ;
      RECT 57.27 3.04 57.47 3.24 ;
      RECT 55.71 2.48 55.91 2.68 ;
      RECT 55.33 3.6 55.53 3.8 ;
      RECT 54.83 2.48 55.03 2.68 ;
      RECT 53.87 2.48 54.07 2.68 ;
      RECT 53.15 2.48 53.35 2.68 ;
      RECT 52.15 1.92 52.35 2.12 ;
      RECT 50.71 3.04 50.91 3.24 ;
      RECT 44.575 2.935 44.775 3.135 ;
      RECT 43.795 0.9 43.995 1.1 ;
      RECT 43.565 3.04 43.765 3.24 ;
      RECT 43.085 2.315 43.285 2.515 ;
      RECT 42.085 7.125 42.285 7.325 ;
      RECT 41.485 3.04 41.685 3.24 ;
      RECT 39.925 2.48 40.125 2.68 ;
      RECT 39.545 3.6 39.745 3.8 ;
      RECT 39.045 2.48 39.245 2.68 ;
      RECT 38.085 2.48 38.285 2.68 ;
      RECT 37.365 2.48 37.565 2.68 ;
      RECT 36.365 1.92 36.565 2.12 ;
      RECT 34.925 3.04 35.125 3.24 ;
      RECT 28.8 2.935 29 3.135 ;
      RECT 28.02 0.9 28.22 1.1 ;
      RECT 27.79 3.04 27.99 3.24 ;
      RECT 27.31 2.315 27.51 2.515 ;
      RECT 26.31 7.125 26.51 7.325 ;
      RECT 25.71 3.04 25.91 3.24 ;
      RECT 24.15 2.48 24.35 2.68 ;
      RECT 23.77 3.6 23.97 3.8 ;
      RECT 23.27 2.48 23.47 2.68 ;
      RECT 22.31 2.48 22.51 2.68 ;
      RECT 21.59 2.48 21.79 2.68 ;
      RECT 20.59 1.92 20.79 2.12 ;
      RECT 19.15 3.04 19.35 3.24 ;
      RECT 13.02 2.935 13.22 3.135 ;
      RECT 12.24 0.9 12.44 1.1 ;
      RECT 12.01 3.04 12.21 3.24 ;
      RECT 11.53 2.315 11.73 2.515 ;
      RECT 10.53 7.125 10.73 7.325 ;
      RECT 9.93 3.04 10.13 3.24 ;
      RECT 8.37 2.48 8.57 2.68 ;
      RECT 7.99 3.6 8.19 3.8 ;
      RECT 7.49 2.48 7.69 2.68 ;
      RECT 6.53 2.48 6.73 2.68 ;
      RECT 5.81 2.48 6.01 2.68 ;
      RECT 4.81 1.92 5.01 2.12 ;
      RECT 3.37 3.04 3.57 3.24 ;
      RECT 0.925 4.35 1.125 4.55 ;
      RECT 0.87 0.09 1.07 0.29 ;
      RECT 0.34 8.59 0.54 8.79 ;
    LAYER met2 ;
      RECT 1.24 8.4 81.405 8.57 ;
      RECT 81.235 7.275 81.405 8.57 ;
      RECT 1.24 6.255 1.41 8.57 ;
      RECT 81.205 7.275 81.555 7.625 ;
      RECT 1.175 6.255 1.465 6.605 ;
      RECT 78.045 6.22 78.365 6.545 ;
      RECT 78.075 5.695 78.245 6.545 ;
      RECT 78.075 5.695 78.25 6.045 ;
      RECT 78.075 5.695 79.05 5.87 ;
      RECT 78.875 1.965 79.05 5.87 ;
      RECT 78.82 1.965 79.17 2.315 ;
      RECT 78.845 6.655 79.17 6.98 ;
      RECT 77.73 6.745 79.17 6.915 ;
      RECT 77.73 2.395 77.89 6.915 ;
      RECT 78.045 2.365 78.365 2.685 ;
      RECT 77.73 2.395 78.365 2.565 ;
      RECT 67.815 1.92 68.075 2.18 ;
      RECT 67.87 1.88 68.175 2.16 ;
      RECT 67.87 1.42 68.045 2.18 ;
      RECT 76.385 1.34 76.735 1.69 ;
      RECT 67.87 1.42 76.735 1.595 ;
      RECT 76.06 2.85 76.43 3.22 ;
      RECT 76.145 2.235 76.315 3.22 ;
      RECT 72.165 2.455 72.4 2.715 ;
      RECT 75.31 2.235 75.475 2.495 ;
      RECT 75.215 2.225 75.23 2.495 ;
      RECT 75.31 2.235 76.315 2.415 ;
      RECT 73.815 1.795 73.855 1.935 ;
      RECT 75.23 2.23 75.31 2.495 ;
      RECT 75.175 2.225 75.215 2.461 ;
      RECT 75.161 2.225 75.175 2.461 ;
      RECT 75.075 2.23 75.161 2.463 ;
      RECT 75.03 2.237 75.075 2.465 ;
      RECT 75 2.237 75.03 2.467 ;
      RECT 74.975 2.232 75 2.469 ;
      RECT 74.945 2.228 74.975 2.478 ;
      RECT 74.935 2.225 74.945 2.49 ;
      RECT 74.93 2.225 74.935 2.498 ;
      RECT 74.925 2.225 74.93 2.503 ;
      RECT 74.915 2.224 74.925 2.513 ;
      RECT 74.91 2.223 74.915 2.523 ;
      RECT 74.895 2.222 74.91 2.528 ;
      RECT 74.867 2.219 74.895 2.555 ;
      RECT 74.781 2.211 74.867 2.555 ;
      RECT 74.695 2.2 74.781 2.555 ;
      RECT 74.655 2.185 74.695 2.555 ;
      RECT 74.615 2.159 74.655 2.555 ;
      RECT 74.61 2.141 74.615 2.367 ;
      RECT 74.6 2.137 74.61 2.357 ;
      RECT 74.585 2.127 74.6 2.344 ;
      RECT 74.565 2.111 74.585 2.329 ;
      RECT 74.55 2.096 74.565 2.314 ;
      RECT 74.54 2.085 74.55 2.304 ;
      RECT 74.515 2.069 74.54 2.293 ;
      RECT 74.51 2.056 74.515 2.283 ;
      RECT 74.505 2.052 74.51 2.278 ;
      RECT 74.45 2.038 74.505 2.256 ;
      RECT 74.411 2.019 74.45 2.22 ;
      RECT 74.325 1.993 74.411 2.173 ;
      RECT 74.321 1.975 74.325 2.139 ;
      RECT 74.235 1.956 74.321 2.117 ;
      RECT 74.23 1.938 74.235 2.095 ;
      RECT 74.225 1.936 74.23 2.093 ;
      RECT 74.215 1.935 74.225 2.088 ;
      RECT 74.155 1.922 74.215 2.074 ;
      RECT 74.11 1.9 74.155 2.053 ;
      RECT 74.05 1.877 74.11 2.032 ;
      RECT 73.986 1.852 74.05 2.007 ;
      RECT 73.9 1.822 73.986 1.976 ;
      RECT 73.885 1.802 73.9 1.955 ;
      RECT 73.855 1.797 73.885 1.946 ;
      RECT 73.802 1.795 73.815 1.935 ;
      RECT 73.716 1.795 73.802 1.937 ;
      RECT 73.63 1.795 73.716 1.939 ;
      RECT 73.61 1.795 73.63 1.943 ;
      RECT 73.565 1.797 73.61 1.954 ;
      RECT 73.525 1.807 73.565 1.97 ;
      RECT 73.521 1.816 73.525 1.978 ;
      RECT 73.435 1.836 73.521 1.994 ;
      RECT 73.425 1.855 73.435 2.012 ;
      RECT 73.42 1.857 73.425 2.015 ;
      RECT 73.41 1.861 73.42 2.018 ;
      RECT 73.39 1.866 73.41 2.028 ;
      RECT 73.36 1.876 73.39 2.048 ;
      RECT 73.355 1.883 73.36 2.062 ;
      RECT 73.345 1.887 73.355 2.069 ;
      RECT 73.33 1.895 73.345 2.08 ;
      RECT 73.32 1.905 73.33 2.091 ;
      RECT 73.31 1.912 73.32 2.099 ;
      RECT 73.285 1.925 73.31 2.114 ;
      RECT 73.221 1.961 73.285 2.153 ;
      RECT 73.135 2.024 73.221 2.217 ;
      RECT 73.1 2.075 73.135 2.27 ;
      RECT 73.095 2.092 73.1 2.287 ;
      RECT 73.08 2.101 73.095 2.294 ;
      RECT 73.06 2.116 73.08 2.308 ;
      RECT 73.055 2.127 73.06 2.318 ;
      RECT 73.035 2.14 73.055 2.328 ;
      RECT 73.03 2.15 73.035 2.338 ;
      RECT 73.015 2.155 73.03 2.347 ;
      RECT 73.005 2.165 73.015 2.358 ;
      RECT 72.975 2.182 73.005 2.375 ;
      RECT 72.965 2.2 72.975 2.393 ;
      RECT 72.95 2.211 72.965 2.404 ;
      RECT 72.91 2.235 72.95 2.42 ;
      RECT 72.875 2.269 72.91 2.437 ;
      RECT 72.845 2.292 72.875 2.449 ;
      RECT 72.83 2.302 72.845 2.458 ;
      RECT 72.79 2.312 72.83 2.469 ;
      RECT 72.77 2.323 72.79 2.481 ;
      RECT 72.765 2.327 72.77 2.488 ;
      RECT 72.75 2.331 72.765 2.493 ;
      RECT 72.74 2.336 72.75 2.498 ;
      RECT 72.735 2.339 72.74 2.501 ;
      RECT 72.705 2.345 72.735 2.508 ;
      RECT 72.67 2.355 72.705 2.522 ;
      RECT 72.61 2.37 72.67 2.542 ;
      RECT 72.555 2.39 72.61 2.566 ;
      RECT 72.526 2.405 72.555 2.584 ;
      RECT 72.44 2.425 72.526 2.609 ;
      RECT 72.435 2.44 72.44 2.629 ;
      RECT 72.425 2.443 72.435 2.63 ;
      RECT 72.4 2.45 72.425 2.715 ;
      RECT 75.095 2.943 75.375 3.28 ;
      RECT 75.095 2.953 75.38 3.238 ;
      RECT 75.095 2.962 75.385 3.135 ;
      RECT 75.095 2.977 75.39 3.003 ;
      RECT 75.095 2.805 75.355 3.28 ;
      RECT 65.395 6.655 65.745 7.005 ;
      RECT 74.22 6.61 74.57 6.96 ;
      RECT 65.395 6.685 74.57 6.885 ;
      RECT 72.815 3.685 72.825 3.875 ;
      RECT 71.075 3.56 71.355 3.84 ;
      RECT 74.12 2.5 74.125 2.985 ;
      RECT 74.015 2.5 74.075 2.76 ;
      RECT 74.34 3.47 74.345 3.545 ;
      RECT 74.33 3.337 74.34 3.58 ;
      RECT 74.32 3.172 74.33 3.601 ;
      RECT 74.315 3.042 74.32 3.617 ;
      RECT 74.305 2.932 74.315 3.633 ;
      RECT 74.3 2.831 74.305 3.65 ;
      RECT 74.295 2.813 74.3 3.66 ;
      RECT 74.29 2.795 74.295 3.67 ;
      RECT 74.28 2.77 74.29 3.685 ;
      RECT 74.275 2.75 74.28 3.7 ;
      RECT 74.255 2.5 74.275 3.725 ;
      RECT 74.24 2.5 74.255 3.758 ;
      RECT 74.21 2.5 74.24 3.78 ;
      RECT 74.19 2.5 74.21 3.794 ;
      RECT 74.17 2.5 74.19 3.31 ;
      RECT 74.185 3.377 74.19 3.799 ;
      RECT 74.18 3.407 74.185 3.801 ;
      RECT 74.175 3.42 74.18 3.804 ;
      RECT 74.17 3.43 74.175 3.808 ;
      RECT 74.165 2.5 74.17 3.228 ;
      RECT 74.165 3.44 74.17 3.81 ;
      RECT 74.16 2.5 74.165 3.205 ;
      RECT 74.15 3.462 74.165 3.81 ;
      RECT 74.145 2.5 74.16 3.15 ;
      RECT 74.14 3.487 74.15 3.81 ;
      RECT 74.14 2.5 74.145 3.095 ;
      RECT 74.13 2.5 74.14 3.043 ;
      RECT 74.135 3.5 74.14 3.811 ;
      RECT 74.13 3.512 74.135 3.812 ;
      RECT 74.125 2.5 74.13 3.003 ;
      RECT 74.125 3.525 74.13 3.813 ;
      RECT 74.11 3.54 74.125 3.814 ;
      RECT 74.115 2.5 74.12 2.965 ;
      RECT 74.11 2.5 74.115 2.93 ;
      RECT 74.105 2.5 74.11 2.905 ;
      RECT 74.1 3.567 74.11 3.816 ;
      RECT 74.095 2.5 74.105 2.863 ;
      RECT 74.095 3.585 74.1 3.817 ;
      RECT 74.09 2.5 74.095 2.823 ;
      RECT 74.09 3.592 74.095 3.818 ;
      RECT 74.085 2.5 74.09 2.795 ;
      RECT 74.08 3.61 74.09 3.819 ;
      RECT 74.075 2.5 74.085 2.775 ;
      RECT 74.07 3.63 74.08 3.821 ;
      RECT 74.06 3.647 74.07 3.822 ;
      RECT 74.025 3.67 74.06 3.825 ;
      RECT 73.97 3.688 74.025 3.831 ;
      RECT 73.884 3.696 73.97 3.84 ;
      RECT 73.798 3.707 73.884 3.851 ;
      RECT 73.712 3.717 73.798 3.862 ;
      RECT 73.626 3.727 73.712 3.874 ;
      RECT 73.54 3.737 73.626 3.885 ;
      RECT 73.52 3.743 73.54 3.891 ;
      RECT 73.44 3.745 73.52 3.895 ;
      RECT 73.435 3.744 73.44 3.9 ;
      RECT 73.427 3.743 73.435 3.9 ;
      RECT 73.341 3.739 73.427 3.898 ;
      RECT 73.255 3.731 73.341 3.895 ;
      RECT 73.169 3.722 73.255 3.891 ;
      RECT 73.083 3.714 73.169 3.888 ;
      RECT 72.997 3.706 73.083 3.884 ;
      RECT 72.911 3.697 72.997 3.881 ;
      RECT 72.825 3.689 72.911 3.877 ;
      RECT 72.77 3.682 72.815 3.875 ;
      RECT 72.685 3.675 72.77 3.873 ;
      RECT 72.611 3.667 72.685 3.869 ;
      RECT 72.525 3.659 72.611 3.866 ;
      RECT 72.522 3.655 72.525 3.864 ;
      RECT 72.436 3.651 72.522 3.863 ;
      RECT 72.35 3.643 72.436 3.86 ;
      RECT 72.265 3.638 72.35 3.857 ;
      RECT 72.179 3.635 72.265 3.854 ;
      RECT 72.093 3.633 72.179 3.851 ;
      RECT 72.007 3.63 72.093 3.848 ;
      RECT 71.921 3.627 72.007 3.845 ;
      RECT 71.835 3.624 71.921 3.842 ;
      RECT 71.759 3.622 71.835 3.839 ;
      RECT 71.673 3.619 71.759 3.836 ;
      RECT 71.587 3.616 71.673 3.834 ;
      RECT 71.501 3.614 71.587 3.831 ;
      RECT 71.415 3.611 71.501 3.828 ;
      RECT 71.355 3.602 71.415 3.826 ;
      RECT 73.865 3.22 73.94 3.48 ;
      RECT 73.845 3.2 73.85 3.48 ;
      RECT 73.165 2.985 73.27 3.28 ;
      RECT 67.61 2.96 67.68 3.22 ;
      RECT 73.505 2.835 73.51 3.206 ;
      RECT 73.495 2.89 73.5 3.206 ;
      RECT 73.8 2.06 73.86 2.32 ;
      RECT 73.855 3.215 73.865 3.48 ;
      RECT 73.85 3.205 73.855 3.48 ;
      RECT 73.77 3.152 73.845 3.48 ;
      RECT 73.795 2.06 73.8 2.34 ;
      RECT 73.785 2.06 73.795 2.36 ;
      RECT 73.77 2.06 73.785 2.39 ;
      RECT 73.755 2.06 73.77 2.433 ;
      RECT 73.75 3.095 73.77 3.48 ;
      RECT 73.74 2.06 73.755 2.47 ;
      RECT 73.735 3.075 73.75 3.48 ;
      RECT 73.735 2.06 73.74 2.493 ;
      RECT 73.725 2.06 73.735 2.518 ;
      RECT 73.695 3.042 73.735 3.48 ;
      RECT 73.7 2.06 73.725 2.568 ;
      RECT 73.695 2.06 73.7 2.623 ;
      RECT 73.69 2.06 73.695 2.665 ;
      RECT 73.68 3.005 73.695 3.48 ;
      RECT 73.685 2.06 73.69 2.708 ;
      RECT 73.68 2.06 73.685 2.773 ;
      RECT 73.675 2.06 73.68 2.795 ;
      RECT 73.675 2.993 73.68 3.345 ;
      RECT 73.67 2.06 73.675 2.863 ;
      RECT 73.67 2.985 73.675 3.328 ;
      RECT 73.665 2.06 73.67 2.908 ;
      RECT 73.66 2.967 73.67 3.305 ;
      RECT 73.66 2.06 73.665 2.945 ;
      RECT 73.65 2.06 73.66 3.285 ;
      RECT 73.645 2.06 73.65 3.268 ;
      RECT 73.64 2.06 73.645 3.253 ;
      RECT 73.635 2.06 73.64 3.238 ;
      RECT 73.615 2.06 73.635 3.228 ;
      RECT 73.61 2.06 73.615 3.218 ;
      RECT 73.6 2.06 73.61 3.214 ;
      RECT 73.595 2.337 73.6 3.213 ;
      RECT 73.59 2.36 73.595 3.212 ;
      RECT 73.585 2.39 73.59 3.211 ;
      RECT 73.58 2.417 73.585 3.21 ;
      RECT 73.575 2.445 73.58 3.21 ;
      RECT 73.57 2.472 73.575 3.21 ;
      RECT 73.565 2.492 73.57 3.21 ;
      RECT 73.56 2.52 73.565 3.21 ;
      RECT 73.55 2.562 73.56 3.21 ;
      RECT 73.54 2.607 73.55 3.209 ;
      RECT 73.535 2.66 73.54 3.208 ;
      RECT 73.53 2.692 73.535 3.207 ;
      RECT 73.525 2.712 73.53 3.206 ;
      RECT 73.52 2.75 73.525 3.206 ;
      RECT 73.515 2.772 73.52 3.206 ;
      RECT 73.51 2.797 73.515 3.206 ;
      RECT 73.5 2.862 73.505 3.206 ;
      RECT 73.485 2.922 73.495 3.206 ;
      RECT 73.47 2.932 73.485 3.206 ;
      RECT 73.45 2.942 73.47 3.206 ;
      RECT 73.42 2.947 73.45 3.203 ;
      RECT 73.36 2.957 73.42 3.2 ;
      RECT 73.34 2.966 73.36 3.205 ;
      RECT 73.315 2.972 73.34 3.218 ;
      RECT 73.295 2.977 73.315 3.233 ;
      RECT 73.27 2.982 73.295 3.28 ;
      RECT 73.141 2.984 73.165 3.28 ;
      RECT 73.055 2.979 73.141 3.28 ;
      RECT 73.015 2.976 73.055 3.28 ;
      RECT 72.965 2.978 73.015 3.26 ;
      RECT 72.935 2.982 72.965 3.26 ;
      RECT 72.856 2.992 72.935 3.26 ;
      RECT 72.77 3.007 72.856 3.261 ;
      RECT 72.72 3.017 72.77 3.262 ;
      RECT 72.712 3.02 72.72 3.262 ;
      RECT 72.626 3.022 72.712 3.263 ;
      RECT 72.54 3.026 72.626 3.263 ;
      RECT 72.454 3.03 72.54 3.264 ;
      RECT 72.368 3.033 72.454 3.265 ;
      RECT 72.282 3.037 72.368 3.265 ;
      RECT 72.196 3.041 72.282 3.266 ;
      RECT 72.11 3.044 72.196 3.267 ;
      RECT 72.024 3.048 72.11 3.267 ;
      RECT 71.938 3.052 72.024 3.268 ;
      RECT 71.852 3.056 71.938 3.269 ;
      RECT 71.766 3.059 71.852 3.269 ;
      RECT 71.68 3.063 71.766 3.27 ;
      RECT 71.65 3.065 71.68 3.27 ;
      RECT 71.564 3.068 71.65 3.271 ;
      RECT 71.478 3.072 71.564 3.272 ;
      RECT 71.392 3.076 71.478 3.273 ;
      RECT 71.306 3.079 71.392 3.273 ;
      RECT 71.22 3.083 71.306 3.274 ;
      RECT 71.185 3.088 71.22 3.275 ;
      RECT 71.13 3.098 71.185 3.282 ;
      RECT 71.105 3.11 71.13 3.292 ;
      RECT 71.07 3.123 71.105 3.3 ;
      RECT 71.03 3.14 71.07 3.323 ;
      RECT 71.01 3.153 71.03 3.35 ;
      RECT 70.98 3.165 71.01 3.378 ;
      RECT 70.975 3.173 70.98 3.398 ;
      RECT 70.97 3.176 70.975 3.408 ;
      RECT 70.92 3.188 70.97 3.442 ;
      RECT 70.91 3.203 70.92 3.475 ;
      RECT 70.9 3.209 70.91 3.488 ;
      RECT 70.89 3.216 70.9 3.5 ;
      RECT 70.865 3.229 70.89 3.518 ;
      RECT 70.85 3.244 70.865 3.54 ;
      RECT 70.84 3.252 70.85 3.556 ;
      RECT 70.825 3.261 70.84 3.571 ;
      RECT 70.815 3.271 70.825 3.585 ;
      RECT 70.796 3.284 70.815 3.602 ;
      RECT 70.71 3.329 70.796 3.667 ;
      RECT 70.695 3.374 70.71 3.725 ;
      RECT 70.69 3.383 70.695 3.738 ;
      RECT 70.68 3.39 70.69 3.743 ;
      RECT 70.675 3.395 70.68 3.747 ;
      RECT 70.655 3.405 70.675 3.754 ;
      RECT 70.63 3.425 70.655 3.768 ;
      RECT 70.595 3.45 70.63 3.788 ;
      RECT 70.58 3.473 70.595 3.803 ;
      RECT 70.57 3.483 70.58 3.808 ;
      RECT 70.56 3.491 70.57 3.815 ;
      RECT 70.55 3.5 70.56 3.821 ;
      RECT 70.53 3.512 70.55 3.823 ;
      RECT 70.52 3.525 70.53 3.825 ;
      RECT 70.495 3.54 70.52 3.828 ;
      RECT 70.475 3.557 70.495 3.832 ;
      RECT 70.435 3.585 70.475 3.838 ;
      RECT 70.37 3.632 70.435 3.847 ;
      RECT 70.355 3.665 70.37 3.855 ;
      RECT 70.35 3.672 70.355 3.857 ;
      RECT 70.3 3.697 70.35 3.862 ;
      RECT 70.285 3.721 70.3 3.869 ;
      RECT 70.235 3.726 70.285 3.87 ;
      RECT 70.149 3.73 70.235 3.87 ;
      RECT 70.063 3.73 70.149 3.87 ;
      RECT 69.977 3.73 70.063 3.871 ;
      RECT 69.891 3.73 69.977 3.871 ;
      RECT 69.805 3.73 69.891 3.871 ;
      RECT 69.739 3.73 69.805 3.871 ;
      RECT 69.653 3.73 69.739 3.872 ;
      RECT 69.567 3.73 69.653 3.872 ;
      RECT 69.481 3.731 69.567 3.873 ;
      RECT 69.395 3.731 69.481 3.873 ;
      RECT 69.309 3.731 69.395 3.873 ;
      RECT 69.223 3.731 69.309 3.874 ;
      RECT 69.137 3.731 69.223 3.874 ;
      RECT 69.051 3.732 69.137 3.875 ;
      RECT 68.965 3.732 69.051 3.875 ;
      RECT 68.945 3.732 68.965 3.875 ;
      RECT 68.859 3.732 68.945 3.875 ;
      RECT 68.773 3.732 68.859 3.875 ;
      RECT 68.687 3.733 68.773 3.875 ;
      RECT 68.601 3.733 68.687 3.875 ;
      RECT 68.515 3.733 68.601 3.875 ;
      RECT 68.429 3.734 68.515 3.875 ;
      RECT 68.343 3.734 68.429 3.875 ;
      RECT 68.257 3.734 68.343 3.875 ;
      RECT 68.171 3.734 68.257 3.875 ;
      RECT 68.085 3.735 68.171 3.875 ;
      RECT 68.035 3.732 68.085 3.875 ;
      RECT 68.025 3.73 68.035 3.874 ;
      RECT 68.021 3.73 68.025 3.873 ;
      RECT 67.935 3.725 68.021 3.868 ;
      RECT 67.913 3.718 67.935 3.862 ;
      RECT 67.827 3.709 67.913 3.856 ;
      RECT 67.741 3.696 67.827 3.847 ;
      RECT 67.655 3.682 67.741 3.837 ;
      RECT 67.61 3.672 67.655 3.83 ;
      RECT 67.59 2.96 67.61 3.238 ;
      RECT 67.59 3.665 67.61 3.826 ;
      RECT 67.56 2.96 67.59 3.26 ;
      RECT 67.55 3.632 67.59 3.823 ;
      RECT 67.545 2.96 67.56 3.28 ;
      RECT 67.545 3.597 67.55 3.821 ;
      RECT 67.54 2.96 67.545 3.405 ;
      RECT 67.54 3.557 67.545 3.821 ;
      RECT 67.53 2.96 67.54 3.821 ;
      RECT 67.455 2.96 67.53 3.815 ;
      RECT 67.425 2.96 67.455 3.805 ;
      RECT 67.42 2.96 67.425 3.797 ;
      RECT 67.415 3.002 67.42 3.79 ;
      RECT 67.405 3.071 67.415 3.781 ;
      RECT 67.4 3.141 67.405 3.733 ;
      RECT 67.395 3.205 67.4 3.63 ;
      RECT 67.39 3.24 67.395 3.585 ;
      RECT 67.388 3.277 67.39 3.477 ;
      RECT 67.385 3.285 67.388 3.47 ;
      RECT 67.38 3.35 67.385 3.413 ;
      RECT 71.455 2.44 71.735 2.72 ;
      RECT 71.445 2.44 71.735 2.583 ;
      RECT 71.4 2.305 71.66 2.565 ;
      RECT 71.4 2.42 71.715 2.565 ;
      RECT 71.4 2.39 71.71 2.565 ;
      RECT 71.4 2.377 71.7 2.565 ;
      RECT 71.4 2.367 71.695 2.565 ;
      RECT 67.375 2.35 67.635 2.61 ;
      RECT 71.145 1.9 71.405 2.16 ;
      RECT 71.135 1.925 71.405 2.12 ;
      RECT 71.13 1.925 71.135 2.119 ;
      RECT 71.06 1.92 71.13 2.111 ;
      RECT 70.975 1.907 71.06 2.094 ;
      RECT 70.971 1.899 70.975 2.084 ;
      RECT 70.885 1.892 70.971 2.074 ;
      RECT 70.876 1.884 70.885 2.064 ;
      RECT 70.79 1.877 70.876 2.052 ;
      RECT 70.77 1.868 70.79 2.038 ;
      RECT 70.715 1.863 70.77 2.03 ;
      RECT 70.705 1.857 70.715 2.024 ;
      RECT 70.685 1.855 70.705 2.02 ;
      RECT 70.677 1.854 70.685 2.016 ;
      RECT 70.591 1.846 70.677 2.005 ;
      RECT 70.505 1.832 70.591 1.985 ;
      RECT 70.445 1.82 70.505 1.97 ;
      RECT 70.435 1.815 70.445 1.965 ;
      RECT 70.385 1.815 70.435 1.967 ;
      RECT 70.338 1.817 70.385 1.971 ;
      RECT 70.252 1.824 70.338 1.976 ;
      RECT 70.166 1.832 70.252 1.982 ;
      RECT 70.08 1.841 70.166 1.988 ;
      RECT 70.021 1.847 70.08 1.993 ;
      RECT 69.935 1.852 70.021 1.999 ;
      RECT 69.86 1.857 69.935 2.005 ;
      RECT 69.821 1.859 69.86 2.01 ;
      RECT 69.735 1.856 69.821 2.015 ;
      RECT 69.65 1.854 69.735 2.022 ;
      RECT 69.618 1.853 69.65 2.025 ;
      RECT 69.532 1.852 69.618 2.026 ;
      RECT 69.446 1.851 69.532 2.027 ;
      RECT 69.36 1.85 69.446 2.027 ;
      RECT 69.274 1.849 69.36 2.028 ;
      RECT 69.188 1.848 69.274 2.029 ;
      RECT 69.102 1.847 69.188 2.03 ;
      RECT 69.016 1.846 69.102 2.03 ;
      RECT 68.93 1.845 69.016 2.031 ;
      RECT 68.88 1.845 68.93 2.032 ;
      RECT 68.866 1.846 68.88 2.032 ;
      RECT 68.78 1.853 68.866 2.033 ;
      RECT 68.706 1.864 68.78 2.034 ;
      RECT 68.62 1.873 68.706 2.035 ;
      RECT 68.585 1.88 68.62 2.05 ;
      RECT 68.56 1.883 68.585 2.08 ;
      RECT 68.535 1.892 68.56 2.109 ;
      RECT 68.525 1.903 68.535 2.129 ;
      RECT 68.515 1.911 68.525 2.143 ;
      RECT 68.51 1.917 68.515 2.153 ;
      RECT 68.485 1.934 68.51 2.17 ;
      RECT 68.47 1.956 68.485 2.198 ;
      RECT 68.44 1.982 68.47 2.228 ;
      RECT 68.42 2.011 68.44 2.258 ;
      RECT 68.415 2.026 68.42 2.275 ;
      RECT 68.395 2.041 68.415 2.29 ;
      RECT 68.385 2.059 68.395 2.308 ;
      RECT 68.375 2.07 68.385 2.323 ;
      RECT 68.325 2.102 68.375 2.349 ;
      RECT 68.32 2.132 68.325 2.369 ;
      RECT 68.31 2.145 68.32 2.375 ;
      RECT 68.301 2.155 68.31 2.383 ;
      RECT 68.29 2.166 68.301 2.391 ;
      RECT 68.285 2.176 68.29 2.397 ;
      RECT 68.27 2.197 68.285 2.404 ;
      RECT 68.255 2.227 68.27 2.412 ;
      RECT 68.22 2.257 68.255 2.418 ;
      RECT 68.195 2.275 68.22 2.425 ;
      RECT 68.145 2.283 68.195 2.434 ;
      RECT 68.12 2.288 68.145 2.443 ;
      RECT 68.065 2.294 68.12 2.453 ;
      RECT 68.06 2.299 68.065 2.461 ;
      RECT 68.046 2.302 68.06 2.463 ;
      RECT 67.96 2.314 68.046 2.475 ;
      RECT 67.95 2.326 67.96 2.488 ;
      RECT 67.865 2.339 67.95 2.5 ;
      RECT 67.821 2.356 67.865 2.514 ;
      RECT 67.735 2.373 67.821 2.53 ;
      RECT 67.705 2.387 67.735 2.544 ;
      RECT 67.695 2.392 67.705 2.549 ;
      RECT 67.635 2.395 67.695 2.558 ;
      RECT 70.525 2.665 70.785 2.925 ;
      RECT 70.525 2.665 70.805 2.778 ;
      RECT 70.525 2.665 70.83 2.745 ;
      RECT 70.525 2.665 70.835 2.725 ;
      RECT 70.575 2.44 70.855 2.72 ;
      RECT 70.13 3.175 70.39 3.435 ;
      RECT 70.12 3.032 70.315 3.373 ;
      RECT 70.115 3.14 70.33 3.365 ;
      RECT 70.11 3.19 70.39 3.355 ;
      RECT 70.1 3.267 70.39 3.34 ;
      RECT 70.12 3.115 70.33 3.373 ;
      RECT 70.13 2.99 70.315 3.435 ;
      RECT 70.13 2.885 70.295 3.435 ;
      RECT 70.14 2.872 70.295 3.435 ;
      RECT 70.14 2.83 70.285 3.435 ;
      RECT 70.145 2.755 70.285 3.435 ;
      RECT 70.175 2.405 70.285 3.435 ;
      RECT 70.18 2.135 70.305 2.758 ;
      RECT 70.15 2.71 70.305 2.758 ;
      RECT 70.165 2.512 70.285 3.435 ;
      RECT 70.155 2.622 70.305 2.758 ;
      RECT 70.18 2.135 70.32 2.615 ;
      RECT 70.18 2.135 70.34 2.49 ;
      RECT 70.145 2.135 70.405 2.395 ;
      RECT 69.615 2.44 69.895 2.72 ;
      RECT 69.6 2.44 69.895 2.7 ;
      RECT 67.655 3.305 67.915 3.565 ;
      RECT 69.44 3.16 69.7 3.42 ;
      RECT 69.42 3.18 69.7 3.395 ;
      RECT 69.377 3.18 69.42 3.394 ;
      RECT 69.291 3.181 69.377 3.391 ;
      RECT 69.205 3.182 69.291 3.387 ;
      RECT 69.13 3.184 69.205 3.384 ;
      RECT 69.107 3.185 69.13 3.382 ;
      RECT 69.021 3.186 69.107 3.38 ;
      RECT 68.935 3.187 69.021 3.377 ;
      RECT 68.911 3.188 68.935 3.375 ;
      RECT 68.825 3.19 68.911 3.372 ;
      RECT 68.74 3.192 68.825 3.373 ;
      RECT 68.683 3.193 68.74 3.379 ;
      RECT 68.597 3.195 68.683 3.389 ;
      RECT 68.511 3.198 68.597 3.402 ;
      RECT 68.425 3.2 68.511 3.414 ;
      RECT 68.411 3.201 68.425 3.421 ;
      RECT 68.325 3.202 68.411 3.429 ;
      RECT 68.285 3.204 68.325 3.438 ;
      RECT 68.276 3.205 68.285 3.441 ;
      RECT 68.19 3.213 68.276 3.447 ;
      RECT 68.17 3.222 68.19 3.455 ;
      RECT 68.085 3.237 68.17 3.463 ;
      RECT 68.025 3.26 68.085 3.474 ;
      RECT 68.015 3.272 68.025 3.479 ;
      RECT 67.975 3.282 68.015 3.483 ;
      RECT 67.92 3.299 67.975 3.491 ;
      RECT 67.915 3.309 67.92 3.495 ;
      RECT 68.981 2.44 69.04 2.837 ;
      RECT 68.895 2.44 69.1 2.828 ;
      RECT 68.89 2.47 69.1 2.823 ;
      RECT 68.856 2.47 69.1 2.821 ;
      RECT 68.77 2.47 69.1 2.815 ;
      RECT 68.725 2.47 69.12 2.793 ;
      RECT 68.725 2.47 69.14 2.748 ;
      RECT 68.685 2.47 69.14 2.738 ;
      RECT 68.895 2.44 69.175 2.72 ;
      RECT 68.63 2.44 68.89 2.7 ;
      RECT 66.455 3 66.735 3.28 ;
      RECT 66.425 2.962 66.68 3.265 ;
      RECT 66.42 2.963 66.68 3.263 ;
      RECT 66.415 2.964 66.68 3.257 ;
      RECT 66.41 2.967 66.68 3.25 ;
      RECT 66.405 3 66.735 3.243 ;
      RECT 66.375 2.97 66.68 3.23 ;
      RECT 66.375 2.997 66.7 3.23 ;
      RECT 66.375 2.987 66.695 3.23 ;
      RECT 66.375 2.972 66.69 3.23 ;
      RECT 66.455 2.959 66.67 3.28 ;
      RECT 66.541 2.957 66.67 3.28 ;
      RECT 66.627 2.955 66.655 3.28 ;
      RECT 62.26 6.22 62.58 6.545 ;
      RECT 62.29 5.695 62.46 6.545 ;
      RECT 62.29 5.695 62.465 6.045 ;
      RECT 62.29 5.695 63.265 5.87 ;
      RECT 63.09 1.965 63.265 5.87 ;
      RECT 63.035 1.965 63.385 2.315 ;
      RECT 63.06 6.655 63.385 6.98 ;
      RECT 61.945 6.745 63.385 6.915 ;
      RECT 61.945 2.395 62.105 6.915 ;
      RECT 62.26 2.365 62.58 2.685 ;
      RECT 61.945 2.395 62.58 2.565 ;
      RECT 52.03 1.92 52.29 2.18 ;
      RECT 52.085 1.88 52.39 2.16 ;
      RECT 52.085 1.42 52.26 2.18 ;
      RECT 60.6 1.34 60.95 1.69 ;
      RECT 52.085 1.42 60.95 1.595 ;
      RECT 60.275 2.85 60.645 3.22 ;
      RECT 60.36 2.235 60.53 3.22 ;
      RECT 56.38 2.455 56.615 2.715 ;
      RECT 59.525 2.235 59.69 2.495 ;
      RECT 59.43 2.225 59.445 2.495 ;
      RECT 59.525 2.235 60.53 2.415 ;
      RECT 58.03 1.795 58.07 1.935 ;
      RECT 59.445 2.23 59.525 2.495 ;
      RECT 59.39 2.225 59.43 2.461 ;
      RECT 59.376 2.225 59.39 2.461 ;
      RECT 59.29 2.23 59.376 2.463 ;
      RECT 59.245 2.237 59.29 2.465 ;
      RECT 59.215 2.237 59.245 2.467 ;
      RECT 59.19 2.232 59.215 2.469 ;
      RECT 59.16 2.228 59.19 2.478 ;
      RECT 59.15 2.225 59.16 2.49 ;
      RECT 59.145 2.225 59.15 2.498 ;
      RECT 59.14 2.225 59.145 2.503 ;
      RECT 59.13 2.224 59.14 2.513 ;
      RECT 59.125 2.223 59.13 2.523 ;
      RECT 59.11 2.222 59.125 2.528 ;
      RECT 59.082 2.219 59.11 2.555 ;
      RECT 58.996 2.211 59.082 2.555 ;
      RECT 58.91 2.2 58.996 2.555 ;
      RECT 58.87 2.185 58.91 2.555 ;
      RECT 58.83 2.159 58.87 2.555 ;
      RECT 58.825 2.141 58.83 2.367 ;
      RECT 58.815 2.137 58.825 2.357 ;
      RECT 58.8 2.127 58.815 2.344 ;
      RECT 58.78 2.111 58.8 2.329 ;
      RECT 58.765 2.096 58.78 2.314 ;
      RECT 58.755 2.085 58.765 2.304 ;
      RECT 58.73 2.069 58.755 2.293 ;
      RECT 58.725 2.056 58.73 2.283 ;
      RECT 58.72 2.052 58.725 2.278 ;
      RECT 58.665 2.038 58.72 2.256 ;
      RECT 58.626 2.019 58.665 2.22 ;
      RECT 58.54 1.993 58.626 2.173 ;
      RECT 58.536 1.975 58.54 2.139 ;
      RECT 58.45 1.956 58.536 2.117 ;
      RECT 58.445 1.938 58.45 2.095 ;
      RECT 58.44 1.936 58.445 2.093 ;
      RECT 58.43 1.935 58.44 2.088 ;
      RECT 58.37 1.922 58.43 2.074 ;
      RECT 58.325 1.9 58.37 2.053 ;
      RECT 58.265 1.877 58.325 2.032 ;
      RECT 58.201 1.852 58.265 2.007 ;
      RECT 58.115 1.822 58.201 1.976 ;
      RECT 58.1 1.802 58.115 1.955 ;
      RECT 58.07 1.797 58.1 1.946 ;
      RECT 58.017 1.795 58.03 1.935 ;
      RECT 57.931 1.795 58.017 1.937 ;
      RECT 57.845 1.795 57.931 1.939 ;
      RECT 57.825 1.795 57.845 1.943 ;
      RECT 57.78 1.797 57.825 1.954 ;
      RECT 57.74 1.807 57.78 1.97 ;
      RECT 57.736 1.816 57.74 1.978 ;
      RECT 57.65 1.836 57.736 1.994 ;
      RECT 57.64 1.855 57.65 2.012 ;
      RECT 57.635 1.857 57.64 2.015 ;
      RECT 57.625 1.861 57.635 2.018 ;
      RECT 57.605 1.866 57.625 2.028 ;
      RECT 57.575 1.876 57.605 2.048 ;
      RECT 57.57 1.883 57.575 2.062 ;
      RECT 57.56 1.887 57.57 2.069 ;
      RECT 57.545 1.895 57.56 2.08 ;
      RECT 57.535 1.905 57.545 2.091 ;
      RECT 57.525 1.912 57.535 2.099 ;
      RECT 57.5 1.925 57.525 2.114 ;
      RECT 57.436 1.961 57.5 2.153 ;
      RECT 57.35 2.024 57.436 2.217 ;
      RECT 57.315 2.075 57.35 2.27 ;
      RECT 57.31 2.092 57.315 2.287 ;
      RECT 57.295 2.101 57.31 2.294 ;
      RECT 57.275 2.116 57.295 2.308 ;
      RECT 57.27 2.127 57.275 2.318 ;
      RECT 57.25 2.14 57.27 2.328 ;
      RECT 57.245 2.15 57.25 2.338 ;
      RECT 57.23 2.155 57.245 2.347 ;
      RECT 57.22 2.165 57.23 2.358 ;
      RECT 57.19 2.182 57.22 2.375 ;
      RECT 57.18 2.2 57.19 2.393 ;
      RECT 57.165 2.211 57.18 2.404 ;
      RECT 57.125 2.235 57.165 2.42 ;
      RECT 57.09 2.269 57.125 2.437 ;
      RECT 57.06 2.292 57.09 2.449 ;
      RECT 57.045 2.302 57.06 2.458 ;
      RECT 57.005 2.312 57.045 2.469 ;
      RECT 56.985 2.323 57.005 2.481 ;
      RECT 56.98 2.327 56.985 2.488 ;
      RECT 56.965 2.331 56.98 2.493 ;
      RECT 56.955 2.336 56.965 2.498 ;
      RECT 56.95 2.339 56.955 2.501 ;
      RECT 56.92 2.345 56.95 2.508 ;
      RECT 56.885 2.355 56.92 2.522 ;
      RECT 56.825 2.37 56.885 2.542 ;
      RECT 56.77 2.39 56.825 2.566 ;
      RECT 56.741 2.405 56.77 2.584 ;
      RECT 56.655 2.425 56.741 2.609 ;
      RECT 56.65 2.44 56.655 2.629 ;
      RECT 56.64 2.443 56.65 2.63 ;
      RECT 56.615 2.45 56.64 2.715 ;
      RECT 59.31 2.943 59.59 3.28 ;
      RECT 59.31 2.953 59.595 3.238 ;
      RECT 59.31 2.962 59.6 3.135 ;
      RECT 59.31 2.977 59.605 3.003 ;
      RECT 59.31 2.805 59.57 3.28 ;
      RECT 49.61 6.655 49.96 7.005 ;
      RECT 58.435 6.61 58.785 6.96 ;
      RECT 49.61 6.685 58.785 6.885 ;
      RECT 57.03 3.685 57.04 3.875 ;
      RECT 55.29 3.56 55.57 3.84 ;
      RECT 58.335 2.5 58.34 2.985 ;
      RECT 58.23 2.5 58.29 2.76 ;
      RECT 58.555 3.47 58.56 3.545 ;
      RECT 58.545 3.337 58.555 3.58 ;
      RECT 58.535 3.172 58.545 3.601 ;
      RECT 58.53 3.042 58.535 3.617 ;
      RECT 58.52 2.932 58.53 3.633 ;
      RECT 58.515 2.831 58.52 3.65 ;
      RECT 58.51 2.813 58.515 3.66 ;
      RECT 58.505 2.795 58.51 3.67 ;
      RECT 58.495 2.77 58.505 3.685 ;
      RECT 58.49 2.75 58.495 3.7 ;
      RECT 58.47 2.5 58.49 3.725 ;
      RECT 58.455 2.5 58.47 3.758 ;
      RECT 58.425 2.5 58.455 3.78 ;
      RECT 58.405 2.5 58.425 3.794 ;
      RECT 58.385 2.5 58.405 3.31 ;
      RECT 58.4 3.377 58.405 3.799 ;
      RECT 58.395 3.407 58.4 3.801 ;
      RECT 58.39 3.42 58.395 3.804 ;
      RECT 58.385 3.43 58.39 3.808 ;
      RECT 58.38 2.5 58.385 3.228 ;
      RECT 58.38 3.44 58.385 3.81 ;
      RECT 58.375 2.5 58.38 3.205 ;
      RECT 58.365 3.462 58.38 3.81 ;
      RECT 58.36 2.5 58.375 3.15 ;
      RECT 58.355 3.487 58.365 3.81 ;
      RECT 58.355 2.5 58.36 3.095 ;
      RECT 58.345 2.5 58.355 3.043 ;
      RECT 58.35 3.5 58.355 3.811 ;
      RECT 58.345 3.512 58.35 3.812 ;
      RECT 58.34 2.5 58.345 3.003 ;
      RECT 58.34 3.525 58.345 3.813 ;
      RECT 58.325 3.54 58.34 3.814 ;
      RECT 58.33 2.5 58.335 2.965 ;
      RECT 58.325 2.5 58.33 2.93 ;
      RECT 58.32 2.5 58.325 2.905 ;
      RECT 58.315 3.567 58.325 3.816 ;
      RECT 58.31 2.5 58.32 2.863 ;
      RECT 58.31 3.585 58.315 3.817 ;
      RECT 58.305 2.5 58.31 2.823 ;
      RECT 58.305 3.592 58.31 3.818 ;
      RECT 58.3 2.5 58.305 2.795 ;
      RECT 58.295 3.61 58.305 3.819 ;
      RECT 58.29 2.5 58.3 2.775 ;
      RECT 58.285 3.63 58.295 3.821 ;
      RECT 58.275 3.647 58.285 3.822 ;
      RECT 58.24 3.67 58.275 3.825 ;
      RECT 58.185 3.688 58.24 3.831 ;
      RECT 58.099 3.696 58.185 3.84 ;
      RECT 58.013 3.707 58.099 3.851 ;
      RECT 57.927 3.717 58.013 3.862 ;
      RECT 57.841 3.727 57.927 3.874 ;
      RECT 57.755 3.737 57.841 3.885 ;
      RECT 57.735 3.743 57.755 3.891 ;
      RECT 57.655 3.745 57.735 3.895 ;
      RECT 57.65 3.744 57.655 3.9 ;
      RECT 57.642 3.743 57.65 3.9 ;
      RECT 57.556 3.739 57.642 3.898 ;
      RECT 57.47 3.731 57.556 3.895 ;
      RECT 57.384 3.722 57.47 3.891 ;
      RECT 57.298 3.714 57.384 3.888 ;
      RECT 57.212 3.706 57.298 3.884 ;
      RECT 57.126 3.697 57.212 3.881 ;
      RECT 57.04 3.689 57.126 3.877 ;
      RECT 56.985 3.682 57.03 3.875 ;
      RECT 56.9 3.675 56.985 3.873 ;
      RECT 56.826 3.667 56.9 3.869 ;
      RECT 56.74 3.659 56.826 3.866 ;
      RECT 56.737 3.655 56.74 3.864 ;
      RECT 56.651 3.651 56.737 3.863 ;
      RECT 56.565 3.643 56.651 3.86 ;
      RECT 56.48 3.638 56.565 3.857 ;
      RECT 56.394 3.635 56.48 3.854 ;
      RECT 56.308 3.633 56.394 3.851 ;
      RECT 56.222 3.63 56.308 3.848 ;
      RECT 56.136 3.627 56.222 3.845 ;
      RECT 56.05 3.624 56.136 3.842 ;
      RECT 55.974 3.622 56.05 3.839 ;
      RECT 55.888 3.619 55.974 3.836 ;
      RECT 55.802 3.616 55.888 3.834 ;
      RECT 55.716 3.614 55.802 3.831 ;
      RECT 55.63 3.611 55.716 3.828 ;
      RECT 55.57 3.602 55.63 3.826 ;
      RECT 58.08 3.22 58.155 3.48 ;
      RECT 58.06 3.2 58.065 3.48 ;
      RECT 57.38 2.985 57.485 3.28 ;
      RECT 51.825 2.96 51.895 3.22 ;
      RECT 57.72 2.835 57.725 3.206 ;
      RECT 57.71 2.89 57.715 3.206 ;
      RECT 58.015 2.06 58.075 2.32 ;
      RECT 58.07 3.215 58.08 3.48 ;
      RECT 58.065 3.205 58.07 3.48 ;
      RECT 57.985 3.152 58.06 3.48 ;
      RECT 58.01 2.06 58.015 2.34 ;
      RECT 58 2.06 58.01 2.36 ;
      RECT 57.985 2.06 58 2.39 ;
      RECT 57.97 2.06 57.985 2.433 ;
      RECT 57.965 3.095 57.985 3.48 ;
      RECT 57.955 2.06 57.97 2.47 ;
      RECT 57.95 3.075 57.965 3.48 ;
      RECT 57.95 2.06 57.955 2.493 ;
      RECT 57.94 2.06 57.95 2.518 ;
      RECT 57.91 3.042 57.95 3.48 ;
      RECT 57.915 2.06 57.94 2.568 ;
      RECT 57.91 2.06 57.915 2.623 ;
      RECT 57.905 2.06 57.91 2.665 ;
      RECT 57.895 3.005 57.91 3.48 ;
      RECT 57.9 2.06 57.905 2.708 ;
      RECT 57.895 2.06 57.9 2.773 ;
      RECT 57.89 2.06 57.895 2.795 ;
      RECT 57.89 2.993 57.895 3.345 ;
      RECT 57.885 2.06 57.89 2.863 ;
      RECT 57.885 2.985 57.89 3.328 ;
      RECT 57.88 2.06 57.885 2.908 ;
      RECT 57.875 2.967 57.885 3.305 ;
      RECT 57.875 2.06 57.88 2.945 ;
      RECT 57.865 2.06 57.875 3.285 ;
      RECT 57.86 2.06 57.865 3.268 ;
      RECT 57.855 2.06 57.86 3.253 ;
      RECT 57.85 2.06 57.855 3.238 ;
      RECT 57.83 2.06 57.85 3.228 ;
      RECT 57.825 2.06 57.83 3.218 ;
      RECT 57.815 2.06 57.825 3.214 ;
      RECT 57.81 2.337 57.815 3.213 ;
      RECT 57.805 2.36 57.81 3.212 ;
      RECT 57.8 2.39 57.805 3.211 ;
      RECT 57.795 2.417 57.8 3.21 ;
      RECT 57.79 2.445 57.795 3.21 ;
      RECT 57.785 2.472 57.79 3.21 ;
      RECT 57.78 2.492 57.785 3.21 ;
      RECT 57.775 2.52 57.78 3.21 ;
      RECT 57.765 2.562 57.775 3.21 ;
      RECT 57.755 2.607 57.765 3.209 ;
      RECT 57.75 2.66 57.755 3.208 ;
      RECT 57.745 2.692 57.75 3.207 ;
      RECT 57.74 2.712 57.745 3.206 ;
      RECT 57.735 2.75 57.74 3.206 ;
      RECT 57.73 2.772 57.735 3.206 ;
      RECT 57.725 2.797 57.73 3.206 ;
      RECT 57.715 2.862 57.72 3.206 ;
      RECT 57.7 2.922 57.71 3.206 ;
      RECT 57.685 2.932 57.7 3.206 ;
      RECT 57.665 2.942 57.685 3.206 ;
      RECT 57.635 2.947 57.665 3.203 ;
      RECT 57.575 2.957 57.635 3.2 ;
      RECT 57.555 2.966 57.575 3.205 ;
      RECT 57.53 2.972 57.555 3.218 ;
      RECT 57.51 2.977 57.53 3.233 ;
      RECT 57.485 2.982 57.51 3.28 ;
      RECT 57.356 2.984 57.38 3.28 ;
      RECT 57.27 2.979 57.356 3.28 ;
      RECT 57.23 2.976 57.27 3.28 ;
      RECT 57.18 2.978 57.23 3.26 ;
      RECT 57.15 2.982 57.18 3.26 ;
      RECT 57.071 2.992 57.15 3.26 ;
      RECT 56.985 3.007 57.071 3.261 ;
      RECT 56.935 3.017 56.985 3.262 ;
      RECT 56.927 3.02 56.935 3.262 ;
      RECT 56.841 3.022 56.927 3.263 ;
      RECT 56.755 3.026 56.841 3.263 ;
      RECT 56.669 3.03 56.755 3.264 ;
      RECT 56.583 3.033 56.669 3.265 ;
      RECT 56.497 3.037 56.583 3.265 ;
      RECT 56.411 3.041 56.497 3.266 ;
      RECT 56.325 3.044 56.411 3.267 ;
      RECT 56.239 3.048 56.325 3.267 ;
      RECT 56.153 3.052 56.239 3.268 ;
      RECT 56.067 3.056 56.153 3.269 ;
      RECT 55.981 3.059 56.067 3.269 ;
      RECT 55.895 3.063 55.981 3.27 ;
      RECT 55.865 3.065 55.895 3.27 ;
      RECT 55.779 3.068 55.865 3.271 ;
      RECT 55.693 3.072 55.779 3.272 ;
      RECT 55.607 3.076 55.693 3.273 ;
      RECT 55.521 3.079 55.607 3.273 ;
      RECT 55.435 3.083 55.521 3.274 ;
      RECT 55.4 3.088 55.435 3.275 ;
      RECT 55.345 3.098 55.4 3.282 ;
      RECT 55.32 3.11 55.345 3.292 ;
      RECT 55.285 3.123 55.32 3.3 ;
      RECT 55.245 3.14 55.285 3.323 ;
      RECT 55.225 3.153 55.245 3.35 ;
      RECT 55.195 3.165 55.225 3.378 ;
      RECT 55.19 3.173 55.195 3.398 ;
      RECT 55.185 3.176 55.19 3.408 ;
      RECT 55.135 3.188 55.185 3.442 ;
      RECT 55.125 3.203 55.135 3.475 ;
      RECT 55.115 3.209 55.125 3.488 ;
      RECT 55.105 3.216 55.115 3.5 ;
      RECT 55.08 3.229 55.105 3.518 ;
      RECT 55.065 3.244 55.08 3.54 ;
      RECT 55.055 3.252 55.065 3.556 ;
      RECT 55.04 3.261 55.055 3.571 ;
      RECT 55.03 3.271 55.04 3.585 ;
      RECT 55.011 3.284 55.03 3.602 ;
      RECT 54.925 3.329 55.011 3.667 ;
      RECT 54.91 3.374 54.925 3.725 ;
      RECT 54.905 3.383 54.91 3.738 ;
      RECT 54.895 3.39 54.905 3.743 ;
      RECT 54.89 3.395 54.895 3.747 ;
      RECT 54.87 3.405 54.89 3.754 ;
      RECT 54.845 3.425 54.87 3.768 ;
      RECT 54.81 3.45 54.845 3.788 ;
      RECT 54.795 3.473 54.81 3.803 ;
      RECT 54.785 3.483 54.795 3.808 ;
      RECT 54.775 3.491 54.785 3.815 ;
      RECT 54.765 3.5 54.775 3.821 ;
      RECT 54.745 3.512 54.765 3.823 ;
      RECT 54.735 3.525 54.745 3.825 ;
      RECT 54.71 3.54 54.735 3.828 ;
      RECT 54.69 3.557 54.71 3.832 ;
      RECT 54.65 3.585 54.69 3.838 ;
      RECT 54.585 3.632 54.65 3.847 ;
      RECT 54.57 3.665 54.585 3.855 ;
      RECT 54.565 3.672 54.57 3.857 ;
      RECT 54.515 3.697 54.565 3.862 ;
      RECT 54.5 3.721 54.515 3.869 ;
      RECT 54.45 3.726 54.5 3.87 ;
      RECT 54.364 3.73 54.45 3.87 ;
      RECT 54.278 3.73 54.364 3.87 ;
      RECT 54.192 3.73 54.278 3.871 ;
      RECT 54.106 3.73 54.192 3.871 ;
      RECT 54.02 3.73 54.106 3.871 ;
      RECT 53.954 3.73 54.02 3.871 ;
      RECT 53.868 3.73 53.954 3.872 ;
      RECT 53.782 3.73 53.868 3.872 ;
      RECT 53.696 3.731 53.782 3.873 ;
      RECT 53.61 3.731 53.696 3.873 ;
      RECT 53.524 3.731 53.61 3.873 ;
      RECT 53.438 3.731 53.524 3.874 ;
      RECT 53.352 3.731 53.438 3.874 ;
      RECT 53.266 3.732 53.352 3.875 ;
      RECT 53.18 3.732 53.266 3.875 ;
      RECT 53.16 3.732 53.18 3.875 ;
      RECT 53.074 3.732 53.16 3.875 ;
      RECT 52.988 3.732 53.074 3.875 ;
      RECT 52.902 3.733 52.988 3.875 ;
      RECT 52.816 3.733 52.902 3.875 ;
      RECT 52.73 3.733 52.816 3.875 ;
      RECT 52.644 3.734 52.73 3.875 ;
      RECT 52.558 3.734 52.644 3.875 ;
      RECT 52.472 3.734 52.558 3.875 ;
      RECT 52.386 3.734 52.472 3.875 ;
      RECT 52.3 3.735 52.386 3.875 ;
      RECT 52.25 3.732 52.3 3.875 ;
      RECT 52.24 3.73 52.25 3.874 ;
      RECT 52.236 3.73 52.24 3.873 ;
      RECT 52.15 3.725 52.236 3.868 ;
      RECT 52.128 3.718 52.15 3.862 ;
      RECT 52.042 3.709 52.128 3.856 ;
      RECT 51.956 3.696 52.042 3.847 ;
      RECT 51.87 3.682 51.956 3.837 ;
      RECT 51.825 3.672 51.87 3.83 ;
      RECT 51.805 2.96 51.825 3.238 ;
      RECT 51.805 3.665 51.825 3.826 ;
      RECT 51.775 2.96 51.805 3.26 ;
      RECT 51.765 3.632 51.805 3.823 ;
      RECT 51.76 2.96 51.775 3.28 ;
      RECT 51.76 3.597 51.765 3.821 ;
      RECT 51.755 2.96 51.76 3.405 ;
      RECT 51.755 3.557 51.76 3.821 ;
      RECT 51.745 2.96 51.755 3.821 ;
      RECT 51.67 2.96 51.745 3.815 ;
      RECT 51.64 2.96 51.67 3.805 ;
      RECT 51.635 2.96 51.64 3.797 ;
      RECT 51.63 3.002 51.635 3.79 ;
      RECT 51.62 3.071 51.63 3.781 ;
      RECT 51.615 3.141 51.62 3.733 ;
      RECT 51.61 3.205 51.615 3.63 ;
      RECT 51.605 3.24 51.61 3.585 ;
      RECT 51.603 3.277 51.605 3.477 ;
      RECT 51.6 3.285 51.603 3.47 ;
      RECT 51.595 3.35 51.6 3.413 ;
      RECT 55.67 2.44 55.95 2.72 ;
      RECT 55.66 2.44 55.95 2.583 ;
      RECT 55.615 2.305 55.875 2.565 ;
      RECT 55.615 2.42 55.93 2.565 ;
      RECT 55.615 2.39 55.925 2.565 ;
      RECT 55.615 2.377 55.915 2.565 ;
      RECT 55.615 2.367 55.91 2.565 ;
      RECT 51.59 2.35 51.85 2.61 ;
      RECT 55.36 1.9 55.62 2.16 ;
      RECT 55.35 1.925 55.62 2.12 ;
      RECT 55.345 1.925 55.35 2.119 ;
      RECT 55.275 1.92 55.345 2.111 ;
      RECT 55.19 1.907 55.275 2.094 ;
      RECT 55.186 1.899 55.19 2.084 ;
      RECT 55.1 1.892 55.186 2.074 ;
      RECT 55.091 1.884 55.1 2.064 ;
      RECT 55.005 1.877 55.091 2.052 ;
      RECT 54.985 1.868 55.005 2.038 ;
      RECT 54.93 1.863 54.985 2.03 ;
      RECT 54.92 1.857 54.93 2.024 ;
      RECT 54.9 1.855 54.92 2.02 ;
      RECT 54.892 1.854 54.9 2.016 ;
      RECT 54.806 1.846 54.892 2.005 ;
      RECT 54.72 1.832 54.806 1.985 ;
      RECT 54.66 1.82 54.72 1.97 ;
      RECT 54.65 1.815 54.66 1.965 ;
      RECT 54.6 1.815 54.65 1.967 ;
      RECT 54.553 1.817 54.6 1.971 ;
      RECT 54.467 1.824 54.553 1.976 ;
      RECT 54.381 1.832 54.467 1.982 ;
      RECT 54.295 1.841 54.381 1.988 ;
      RECT 54.236 1.847 54.295 1.993 ;
      RECT 54.15 1.852 54.236 1.999 ;
      RECT 54.075 1.857 54.15 2.005 ;
      RECT 54.036 1.859 54.075 2.01 ;
      RECT 53.95 1.856 54.036 2.015 ;
      RECT 53.865 1.854 53.95 2.022 ;
      RECT 53.833 1.853 53.865 2.025 ;
      RECT 53.747 1.852 53.833 2.026 ;
      RECT 53.661 1.851 53.747 2.027 ;
      RECT 53.575 1.85 53.661 2.027 ;
      RECT 53.489 1.849 53.575 2.028 ;
      RECT 53.403 1.848 53.489 2.029 ;
      RECT 53.317 1.847 53.403 2.03 ;
      RECT 53.231 1.846 53.317 2.03 ;
      RECT 53.145 1.845 53.231 2.031 ;
      RECT 53.095 1.845 53.145 2.032 ;
      RECT 53.081 1.846 53.095 2.032 ;
      RECT 52.995 1.853 53.081 2.033 ;
      RECT 52.921 1.864 52.995 2.034 ;
      RECT 52.835 1.873 52.921 2.035 ;
      RECT 52.8 1.88 52.835 2.05 ;
      RECT 52.775 1.883 52.8 2.08 ;
      RECT 52.75 1.892 52.775 2.109 ;
      RECT 52.74 1.903 52.75 2.129 ;
      RECT 52.73 1.911 52.74 2.143 ;
      RECT 52.725 1.917 52.73 2.153 ;
      RECT 52.7 1.934 52.725 2.17 ;
      RECT 52.685 1.956 52.7 2.198 ;
      RECT 52.655 1.982 52.685 2.228 ;
      RECT 52.635 2.011 52.655 2.258 ;
      RECT 52.63 2.026 52.635 2.275 ;
      RECT 52.61 2.041 52.63 2.29 ;
      RECT 52.6 2.059 52.61 2.308 ;
      RECT 52.59 2.07 52.6 2.323 ;
      RECT 52.54 2.102 52.59 2.349 ;
      RECT 52.535 2.132 52.54 2.369 ;
      RECT 52.525 2.145 52.535 2.375 ;
      RECT 52.516 2.155 52.525 2.383 ;
      RECT 52.505 2.166 52.516 2.391 ;
      RECT 52.5 2.176 52.505 2.397 ;
      RECT 52.485 2.197 52.5 2.404 ;
      RECT 52.47 2.227 52.485 2.412 ;
      RECT 52.435 2.257 52.47 2.418 ;
      RECT 52.41 2.275 52.435 2.425 ;
      RECT 52.36 2.283 52.41 2.434 ;
      RECT 52.335 2.288 52.36 2.443 ;
      RECT 52.28 2.294 52.335 2.453 ;
      RECT 52.275 2.299 52.28 2.461 ;
      RECT 52.261 2.302 52.275 2.463 ;
      RECT 52.175 2.314 52.261 2.475 ;
      RECT 52.165 2.326 52.175 2.488 ;
      RECT 52.08 2.339 52.165 2.5 ;
      RECT 52.036 2.356 52.08 2.514 ;
      RECT 51.95 2.373 52.036 2.53 ;
      RECT 51.92 2.387 51.95 2.544 ;
      RECT 51.91 2.392 51.92 2.549 ;
      RECT 51.85 2.395 51.91 2.558 ;
      RECT 54.74 2.665 55 2.925 ;
      RECT 54.74 2.665 55.02 2.778 ;
      RECT 54.74 2.665 55.045 2.745 ;
      RECT 54.74 2.665 55.05 2.725 ;
      RECT 54.79 2.44 55.07 2.72 ;
      RECT 54.345 3.175 54.605 3.435 ;
      RECT 54.335 3.032 54.53 3.373 ;
      RECT 54.33 3.14 54.545 3.365 ;
      RECT 54.325 3.19 54.605 3.355 ;
      RECT 54.315 3.267 54.605 3.34 ;
      RECT 54.335 3.115 54.545 3.373 ;
      RECT 54.345 2.99 54.53 3.435 ;
      RECT 54.345 2.885 54.51 3.435 ;
      RECT 54.355 2.872 54.51 3.435 ;
      RECT 54.355 2.83 54.5 3.435 ;
      RECT 54.36 2.755 54.5 3.435 ;
      RECT 54.39 2.405 54.5 3.435 ;
      RECT 54.395 2.135 54.52 2.758 ;
      RECT 54.365 2.71 54.52 2.758 ;
      RECT 54.38 2.512 54.5 3.435 ;
      RECT 54.37 2.622 54.52 2.758 ;
      RECT 54.395 2.135 54.535 2.615 ;
      RECT 54.395 2.135 54.555 2.49 ;
      RECT 54.36 2.135 54.62 2.395 ;
      RECT 53.83 2.44 54.11 2.72 ;
      RECT 53.815 2.44 54.11 2.7 ;
      RECT 51.87 3.305 52.13 3.565 ;
      RECT 53.655 3.16 53.915 3.42 ;
      RECT 53.635 3.18 53.915 3.395 ;
      RECT 53.592 3.18 53.635 3.394 ;
      RECT 53.506 3.181 53.592 3.391 ;
      RECT 53.42 3.182 53.506 3.387 ;
      RECT 53.345 3.184 53.42 3.384 ;
      RECT 53.322 3.185 53.345 3.382 ;
      RECT 53.236 3.186 53.322 3.38 ;
      RECT 53.15 3.187 53.236 3.377 ;
      RECT 53.126 3.188 53.15 3.375 ;
      RECT 53.04 3.19 53.126 3.372 ;
      RECT 52.955 3.192 53.04 3.373 ;
      RECT 52.898 3.193 52.955 3.379 ;
      RECT 52.812 3.195 52.898 3.389 ;
      RECT 52.726 3.198 52.812 3.402 ;
      RECT 52.64 3.2 52.726 3.414 ;
      RECT 52.626 3.201 52.64 3.421 ;
      RECT 52.54 3.202 52.626 3.429 ;
      RECT 52.5 3.204 52.54 3.438 ;
      RECT 52.491 3.205 52.5 3.441 ;
      RECT 52.405 3.213 52.491 3.447 ;
      RECT 52.385 3.222 52.405 3.455 ;
      RECT 52.3 3.237 52.385 3.463 ;
      RECT 52.24 3.26 52.3 3.474 ;
      RECT 52.23 3.272 52.24 3.479 ;
      RECT 52.19 3.282 52.23 3.483 ;
      RECT 52.135 3.299 52.19 3.491 ;
      RECT 52.13 3.309 52.135 3.495 ;
      RECT 53.196 2.44 53.255 2.837 ;
      RECT 53.11 2.44 53.315 2.828 ;
      RECT 53.105 2.47 53.315 2.823 ;
      RECT 53.071 2.47 53.315 2.821 ;
      RECT 52.985 2.47 53.315 2.815 ;
      RECT 52.94 2.47 53.335 2.793 ;
      RECT 52.94 2.47 53.355 2.748 ;
      RECT 52.9 2.47 53.355 2.738 ;
      RECT 53.11 2.44 53.39 2.72 ;
      RECT 52.845 2.44 53.105 2.7 ;
      RECT 50.67 3 50.95 3.28 ;
      RECT 50.64 2.962 50.895 3.265 ;
      RECT 50.635 2.963 50.895 3.263 ;
      RECT 50.63 2.964 50.895 3.257 ;
      RECT 50.625 2.967 50.895 3.25 ;
      RECT 50.62 3 50.95 3.243 ;
      RECT 50.59 2.97 50.895 3.23 ;
      RECT 50.59 2.997 50.915 3.23 ;
      RECT 50.59 2.987 50.91 3.23 ;
      RECT 50.59 2.972 50.905 3.23 ;
      RECT 50.67 2.959 50.885 3.28 ;
      RECT 50.756 2.957 50.885 3.28 ;
      RECT 50.842 2.955 50.87 3.28 ;
      RECT 46.475 6.22 46.795 6.545 ;
      RECT 46.505 5.695 46.675 6.545 ;
      RECT 46.505 5.695 46.68 6.045 ;
      RECT 46.505 5.695 47.48 5.87 ;
      RECT 47.305 1.965 47.48 5.87 ;
      RECT 47.25 1.965 47.6 2.315 ;
      RECT 47.275 6.655 47.6 6.98 ;
      RECT 46.16 6.745 47.6 6.915 ;
      RECT 46.16 2.395 46.32 6.915 ;
      RECT 46.475 2.365 46.795 2.685 ;
      RECT 46.16 2.395 46.795 2.565 ;
      RECT 36.245 1.92 36.505 2.18 ;
      RECT 36.3 1.88 36.605 2.16 ;
      RECT 36.3 1.42 36.475 2.18 ;
      RECT 44.815 1.34 45.165 1.69 ;
      RECT 36.3 1.42 45.165 1.595 ;
      RECT 44.49 2.85 44.86 3.22 ;
      RECT 44.575 2.235 44.745 3.22 ;
      RECT 40.595 2.455 40.83 2.715 ;
      RECT 43.74 2.235 43.905 2.495 ;
      RECT 43.645 2.225 43.66 2.495 ;
      RECT 43.74 2.235 44.745 2.415 ;
      RECT 42.245 1.795 42.285 1.935 ;
      RECT 43.66 2.23 43.74 2.495 ;
      RECT 43.605 2.225 43.645 2.461 ;
      RECT 43.591 2.225 43.605 2.461 ;
      RECT 43.505 2.23 43.591 2.463 ;
      RECT 43.46 2.237 43.505 2.465 ;
      RECT 43.43 2.237 43.46 2.467 ;
      RECT 43.405 2.232 43.43 2.469 ;
      RECT 43.375 2.228 43.405 2.478 ;
      RECT 43.365 2.225 43.375 2.49 ;
      RECT 43.36 2.225 43.365 2.498 ;
      RECT 43.355 2.225 43.36 2.503 ;
      RECT 43.345 2.224 43.355 2.513 ;
      RECT 43.34 2.223 43.345 2.523 ;
      RECT 43.325 2.222 43.34 2.528 ;
      RECT 43.297 2.219 43.325 2.555 ;
      RECT 43.211 2.211 43.297 2.555 ;
      RECT 43.125 2.2 43.211 2.555 ;
      RECT 43.085 2.185 43.125 2.555 ;
      RECT 43.045 2.159 43.085 2.555 ;
      RECT 43.04 2.141 43.045 2.367 ;
      RECT 43.03 2.137 43.04 2.357 ;
      RECT 43.015 2.127 43.03 2.344 ;
      RECT 42.995 2.111 43.015 2.329 ;
      RECT 42.98 2.096 42.995 2.314 ;
      RECT 42.97 2.085 42.98 2.304 ;
      RECT 42.945 2.069 42.97 2.293 ;
      RECT 42.94 2.056 42.945 2.283 ;
      RECT 42.935 2.052 42.94 2.278 ;
      RECT 42.88 2.038 42.935 2.256 ;
      RECT 42.841 2.019 42.88 2.22 ;
      RECT 42.755 1.993 42.841 2.173 ;
      RECT 42.751 1.975 42.755 2.139 ;
      RECT 42.665 1.956 42.751 2.117 ;
      RECT 42.66 1.938 42.665 2.095 ;
      RECT 42.655 1.936 42.66 2.093 ;
      RECT 42.645 1.935 42.655 2.088 ;
      RECT 42.585 1.922 42.645 2.074 ;
      RECT 42.54 1.9 42.585 2.053 ;
      RECT 42.48 1.877 42.54 2.032 ;
      RECT 42.416 1.852 42.48 2.007 ;
      RECT 42.33 1.822 42.416 1.976 ;
      RECT 42.315 1.802 42.33 1.955 ;
      RECT 42.285 1.797 42.315 1.946 ;
      RECT 42.232 1.795 42.245 1.935 ;
      RECT 42.146 1.795 42.232 1.937 ;
      RECT 42.06 1.795 42.146 1.939 ;
      RECT 42.04 1.795 42.06 1.943 ;
      RECT 41.995 1.797 42.04 1.954 ;
      RECT 41.955 1.807 41.995 1.97 ;
      RECT 41.951 1.816 41.955 1.978 ;
      RECT 41.865 1.836 41.951 1.994 ;
      RECT 41.855 1.855 41.865 2.012 ;
      RECT 41.85 1.857 41.855 2.015 ;
      RECT 41.84 1.861 41.85 2.018 ;
      RECT 41.82 1.866 41.84 2.028 ;
      RECT 41.79 1.876 41.82 2.048 ;
      RECT 41.785 1.883 41.79 2.062 ;
      RECT 41.775 1.887 41.785 2.069 ;
      RECT 41.76 1.895 41.775 2.08 ;
      RECT 41.75 1.905 41.76 2.091 ;
      RECT 41.74 1.912 41.75 2.099 ;
      RECT 41.715 1.925 41.74 2.114 ;
      RECT 41.651 1.961 41.715 2.153 ;
      RECT 41.565 2.024 41.651 2.217 ;
      RECT 41.53 2.075 41.565 2.27 ;
      RECT 41.525 2.092 41.53 2.287 ;
      RECT 41.51 2.101 41.525 2.294 ;
      RECT 41.49 2.116 41.51 2.308 ;
      RECT 41.485 2.127 41.49 2.318 ;
      RECT 41.465 2.14 41.485 2.328 ;
      RECT 41.46 2.15 41.465 2.338 ;
      RECT 41.445 2.155 41.46 2.347 ;
      RECT 41.435 2.165 41.445 2.358 ;
      RECT 41.405 2.182 41.435 2.375 ;
      RECT 41.395 2.2 41.405 2.393 ;
      RECT 41.38 2.211 41.395 2.404 ;
      RECT 41.34 2.235 41.38 2.42 ;
      RECT 41.305 2.269 41.34 2.437 ;
      RECT 41.275 2.292 41.305 2.449 ;
      RECT 41.26 2.302 41.275 2.458 ;
      RECT 41.22 2.312 41.26 2.469 ;
      RECT 41.2 2.323 41.22 2.481 ;
      RECT 41.195 2.327 41.2 2.488 ;
      RECT 41.18 2.331 41.195 2.493 ;
      RECT 41.17 2.336 41.18 2.498 ;
      RECT 41.165 2.339 41.17 2.501 ;
      RECT 41.135 2.345 41.165 2.508 ;
      RECT 41.1 2.355 41.135 2.522 ;
      RECT 41.04 2.37 41.1 2.542 ;
      RECT 40.985 2.39 41.04 2.566 ;
      RECT 40.956 2.405 40.985 2.584 ;
      RECT 40.87 2.425 40.956 2.609 ;
      RECT 40.865 2.44 40.87 2.629 ;
      RECT 40.855 2.443 40.865 2.63 ;
      RECT 40.83 2.45 40.855 2.715 ;
      RECT 43.525 2.943 43.805 3.28 ;
      RECT 43.525 2.953 43.81 3.238 ;
      RECT 43.525 2.962 43.815 3.135 ;
      RECT 43.525 2.977 43.82 3.003 ;
      RECT 43.525 2.805 43.785 3.28 ;
      RECT 33.88 6.66 34.23 7.01 ;
      RECT 42.705 6.615 43.055 6.965 ;
      RECT 33.88 6.69 43.055 6.89 ;
      RECT 41.245 3.685 41.255 3.875 ;
      RECT 39.505 3.56 39.785 3.84 ;
      RECT 42.55 2.5 42.555 2.985 ;
      RECT 42.445 2.5 42.505 2.76 ;
      RECT 42.77 3.47 42.775 3.545 ;
      RECT 42.76 3.337 42.77 3.58 ;
      RECT 42.75 3.172 42.76 3.601 ;
      RECT 42.745 3.042 42.75 3.617 ;
      RECT 42.735 2.932 42.745 3.633 ;
      RECT 42.73 2.831 42.735 3.65 ;
      RECT 42.725 2.813 42.73 3.66 ;
      RECT 42.72 2.795 42.725 3.67 ;
      RECT 42.71 2.77 42.72 3.685 ;
      RECT 42.705 2.75 42.71 3.7 ;
      RECT 42.685 2.5 42.705 3.725 ;
      RECT 42.67 2.5 42.685 3.758 ;
      RECT 42.64 2.5 42.67 3.78 ;
      RECT 42.62 2.5 42.64 3.794 ;
      RECT 42.6 2.5 42.62 3.31 ;
      RECT 42.615 3.377 42.62 3.799 ;
      RECT 42.61 3.407 42.615 3.801 ;
      RECT 42.605 3.42 42.61 3.804 ;
      RECT 42.6 3.43 42.605 3.808 ;
      RECT 42.595 2.5 42.6 3.228 ;
      RECT 42.595 3.44 42.6 3.81 ;
      RECT 42.59 2.5 42.595 3.205 ;
      RECT 42.58 3.462 42.595 3.81 ;
      RECT 42.575 2.5 42.59 3.15 ;
      RECT 42.57 3.487 42.58 3.81 ;
      RECT 42.57 2.5 42.575 3.095 ;
      RECT 42.56 2.5 42.57 3.043 ;
      RECT 42.565 3.5 42.57 3.811 ;
      RECT 42.56 3.512 42.565 3.812 ;
      RECT 42.555 2.5 42.56 3.003 ;
      RECT 42.555 3.525 42.56 3.813 ;
      RECT 42.54 3.54 42.555 3.814 ;
      RECT 42.545 2.5 42.55 2.965 ;
      RECT 42.54 2.5 42.545 2.93 ;
      RECT 42.535 2.5 42.54 2.905 ;
      RECT 42.53 3.567 42.54 3.816 ;
      RECT 42.525 2.5 42.535 2.863 ;
      RECT 42.525 3.585 42.53 3.817 ;
      RECT 42.52 2.5 42.525 2.823 ;
      RECT 42.52 3.592 42.525 3.818 ;
      RECT 42.515 2.5 42.52 2.795 ;
      RECT 42.51 3.61 42.52 3.819 ;
      RECT 42.505 2.5 42.515 2.775 ;
      RECT 42.5 3.63 42.51 3.821 ;
      RECT 42.49 3.647 42.5 3.822 ;
      RECT 42.455 3.67 42.49 3.825 ;
      RECT 42.4 3.688 42.455 3.831 ;
      RECT 42.314 3.696 42.4 3.84 ;
      RECT 42.228 3.707 42.314 3.851 ;
      RECT 42.142 3.717 42.228 3.862 ;
      RECT 42.056 3.727 42.142 3.874 ;
      RECT 41.97 3.737 42.056 3.885 ;
      RECT 41.95 3.743 41.97 3.891 ;
      RECT 41.87 3.745 41.95 3.895 ;
      RECT 41.865 3.744 41.87 3.9 ;
      RECT 41.857 3.743 41.865 3.9 ;
      RECT 41.771 3.739 41.857 3.898 ;
      RECT 41.685 3.731 41.771 3.895 ;
      RECT 41.599 3.722 41.685 3.891 ;
      RECT 41.513 3.714 41.599 3.888 ;
      RECT 41.427 3.706 41.513 3.884 ;
      RECT 41.341 3.697 41.427 3.881 ;
      RECT 41.255 3.689 41.341 3.877 ;
      RECT 41.2 3.682 41.245 3.875 ;
      RECT 41.115 3.675 41.2 3.873 ;
      RECT 41.041 3.667 41.115 3.869 ;
      RECT 40.955 3.659 41.041 3.866 ;
      RECT 40.952 3.655 40.955 3.864 ;
      RECT 40.866 3.651 40.952 3.863 ;
      RECT 40.78 3.643 40.866 3.86 ;
      RECT 40.695 3.638 40.78 3.857 ;
      RECT 40.609 3.635 40.695 3.854 ;
      RECT 40.523 3.633 40.609 3.851 ;
      RECT 40.437 3.63 40.523 3.848 ;
      RECT 40.351 3.627 40.437 3.845 ;
      RECT 40.265 3.624 40.351 3.842 ;
      RECT 40.189 3.622 40.265 3.839 ;
      RECT 40.103 3.619 40.189 3.836 ;
      RECT 40.017 3.616 40.103 3.834 ;
      RECT 39.931 3.614 40.017 3.831 ;
      RECT 39.845 3.611 39.931 3.828 ;
      RECT 39.785 3.602 39.845 3.826 ;
      RECT 42.295 3.22 42.37 3.48 ;
      RECT 42.275 3.2 42.28 3.48 ;
      RECT 41.595 2.985 41.7 3.28 ;
      RECT 36.04 2.96 36.11 3.22 ;
      RECT 41.935 2.835 41.94 3.206 ;
      RECT 41.925 2.89 41.93 3.206 ;
      RECT 42.23 2.06 42.29 2.32 ;
      RECT 42.285 3.215 42.295 3.48 ;
      RECT 42.28 3.205 42.285 3.48 ;
      RECT 42.2 3.152 42.275 3.48 ;
      RECT 42.225 2.06 42.23 2.34 ;
      RECT 42.215 2.06 42.225 2.36 ;
      RECT 42.2 2.06 42.215 2.39 ;
      RECT 42.185 2.06 42.2 2.433 ;
      RECT 42.18 3.095 42.2 3.48 ;
      RECT 42.17 2.06 42.185 2.47 ;
      RECT 42.165 3.075 42.18 3.48 ;
      RECT 42.165 2.06 42.17 2.493 ;
      RECT 42.155 2.06 42.165 2.518 ;
      RECT 42.125 3.042 42.165 3.48 ;
      RECT 42.13 2.06 42.155 2.568 ;
      RECT 42.125 2.06 42.13 2.623 ;
      RECT 42.12 2.06 42.125 2.665 ;
      RECT 42.11 3.005 42.125 3.48 ;
      RECT 42.115 2.06 42.12 2.708 ;
      RECT 42.11 2.06 42.115 2.773 ;
      RECT 42.105 2.06 42.11 2.795 ;
      RECT 42.105 2.993 42.11 3.345 ;
      RECT 42.1 2.06 42.105 2.863 ;
      RECT 42.1 2.985 42.105 3.328 ;
      RECT 42.095 2.06 42.1 2.908 ;
      RECT 42.09 2.967 42.1 3.305 ;
      RECT 42.09 2.06 42.095 2.945 ;
      RECT 42.08 2.06 42.09 3.285 ;
      RECT 42.075 2.06 42.08 3.268 ;
      RECT 42.07 2.06 42.075 3.253 ;
      RECT 42.065 2.06 42.07 3.238 ;
      RECT 42.045 2.06 42.065 3.228 ;
      RECT 42.04 2.06 42.045 3.218 ;
      RECT 42.03 2.06 42.04 3.214 ;
      RECT 42.025 2.337 42.03 3.213 ;
      RECT 42.02 2.36 42.025 3.212 ;
      RECT 42.015 2.39 42.02 3.211 ;
      RECT 42.01 2.417 42.015 3.21 ;
      RECT 42.005 2.445 42.01 3.21 ;
      RECT 42 2.472 42.005 3.21 ;
      RECT 41.995 2.492 42 3.21 ;
      RECT 41.99 2.52 41.995 3.21 ;
      RECT 41.98 2.562 41.99 3.21 ;
      RECT 41.97 2.607 41.98 3.209 ;
      RECT 41.965 2.66 41.97 3.208 ;
      RECT 41.96 2.692 41.965 3.207 ;
      RECT 41.955 2.712 41.96 3.206 ;
      RECT 41.95 2.75 41.955 3.206 ;
      RECT 41.945 2.772 41.95 3.206 ;
      RECT 41.94 2.797 41.945 3.206 ;
      RECT 41.93 2.862 41.935 3.206 ;
      RECT 41.915 2.922 41.925 3.206 ;
      RECT 41.9 2.932 41.915 3.206 ;
      RECT 41.88 2.942 41.9 3.206 ;
      RECT 41.85 2.947 41.88 3.203 ;
      RECT 41.79 2.957 41.85 3.2 ;
      RECT 41.77 2.966 41.79 3.205 ;
      RECT 41.745 2.972 41.77 3.218 ;
      RECT 41.725 2.977 41.745 3.233 ;
      RECT 41.7 2.982 41.725 3.28 ;
      RECT 41.571 2.984 41.595 3.28 ;
      RECT 41.485 2.979 41.571 3.28 ;
      RECT 41.445 2.976 41.485 3.28 ;
      RECT 41.395 2.978 41.445 3.26 ;
      RECT 41.365 2.982 41.395 3.26 ;
      RECT 41.286 2.992 41.365 3.26 ;
      RECT 41.2 3.007 41.286 3.261 ;
      RECT 41.15 3.017 41.2 3.262 ;
      RECT 41.142 3.02 41.15 3.262 ;
      RECT 41.056 3.022 41.142 3.263 ;
      RECT 40.97 3.026 41.056 3.263 ;
      RECT 40.884 3.03 40.97 3.264 ;
      RECT 40.798 3.033 40.884 3.265 ;
      RECT 40.712 3.037 40.798 3.265 ;
      RECT 40.626 3.041 40.712 3.266 ;
      RECT 40.54 3.044 40.626 3.267 ;
      RECT 40.454 3.048 40.54 3.267 ;
      RECT 40.368 3.052 40.454 3.268 ;
      RECT 40.282 3.056 40.368 3.269 ;
      RECT 40.196 3.059 40.282 3.269 ;
      RECT 40.11 3.063 40.196 3.27 ;
      RECT 40.08 3.065 40.11 3.27 ;
      RECT 39.994 3.068 40.08 3.271 ;
      RECT 39.908 3.072 39.994 3.272 ;
      RECT 39.822 3.076 39.908 3.273 ;
      RECT 39.736 3.079 39.822 3.273 ;
      RECT 39.65 3.083 39.736 3.274 ;
      RECT 39.615 3.088 39.65 3.275 ;
      RECT 39.56 3.098 39.615 3.282 ;
      RECT 39.535 3.11 39.56 3.292 ;
      RECT 39.5 3.123 39.535 3.3 ;
      RECT 39.46 3.14 39.5 3.323 ;
      RECT 39.44 3.153 39.46 3.35 ;
      RECT 39.41 3.165 39.44 3.378 ;
      RECT 39.405 3.173 39.41 3.398 ;
      RECT 39.4 3.176 39.405 3.408 ;
      RECT 39.35 3.188 39.4 3.442 ;
      RECT 39.34 3.203 39.35 3.475 ;
      RECT 39.33 3.209 39.34 3.488 ;
      RECT 39.32 3.216 39.33 3.5 ;
      RECT 39.295 3.229 39.32 3.518 ;
      RECT 39.28 3.244 39.295 3.54 ;
      RECT 39.27 3.252 39.28 3.556 ;
      RECT 39.255 3.261 39.27 3.571 ;
      RECT 39.245 3.271 39.255 3.585 ;
      RECT 39.226 3.284 39.245 3.602 ;
      RECT 39.14 3.329 39.226 3.667 ;
      RECT 39.125 3.374 39.14 3.725 ;
      RECT 39.12 3.383 39.125 3.738 ;
      RECT 39.11 3.39 39.12 3.743 ;
      RECT 39.105 3.395 39.11 3.747 ;
      RECT 39.085 3.405 39.105 3.754 ;
      RECT 39.06 3.425 39.085 3.768 ;
      RECT 39.025 3.45 39.06 3.788 ;
      RECT 39.01 3.473 39.025 3.803 ;
      RECT 39 3.483 39.01 3.808 ;
      RECT 38.99 3.491 39 3.815 ;
      RECT 38.98 3.5 38.99 3.821 ;
      RECT 38.96 3.512 38.98 3.823 ;
      RECT 38.95 3.525 38.96 3.825 ;
      RECT 38.925 3.54 38.95 3.828 ;
      RECT 38.905 3.557 38.925 3.832 ;
      RECT 38.865 3.585 38.905 3.838 ;
      RECT 38.8 3.632 38.865 3.847 ;
      RECT 38.785 3.665 38.8 3.855 ;
      RECT 38.78 3.672 38.785 3.857 ;
      RECT 38.73 3.697 38.78 3.862 ;
      RECT 38.715 3.721 38.73 3.869 ;
      RECT 38.665 3.726 38.715 3.87 ;
      RECT 38.579 3.73 38.665 3.87 ;
      RECT 38.493 3.73 38.579 3.87 ;
      RECT 38.407 3.73 38.493 3.871 ;
      RECT 38.321 3.73 38.407 3.871 ;
      RECT 38.235 3.73 38.321 3.871 ;
      RECT 38.169 3.73 38.235 3.871 ;
      RECT 38.083 3.73 38.169 3.872 ;
      RECT 37.997 3.73 38.083 3.872 ;
      RECT 37.911 3.731 37.997 3.873 ;
      RECT 37.825 3.731 37.911 3.873 ;
      RECT 37.739 3.731 37.825 3.873 ;
      RECT 37.653 3.731 37.739 3.874 ;
      RECT 37.567 3.731 37.653 3.874 ;
      RECT 37.481 3.732 37.567 3.875 ;
      RECT 37.395 3.732 37.481 3.875 ;
      RECT 37.375 3.732 37.395 3.875 ;
      RECT 37.289 3.732 37.375 3.875 ;
      RECT 37.203 3.732 37.289 3.875 ;
      RECT 37.117 3.733 37.203 3.875 ;
      RECT 37.031 3.733 37.117 3.875 ;
      RECT 36.945 3.733 37.031 3.875 ;
      RECT 36.859 3.734 36.945 3.875 ;
      RECT 36.773 3.734 36.859 3.875 ;
      RECT 36.687 3.734 36.773 3.875 ;
      RECT 36.601 3.734 36.687 3.875 ;
      RECT 36.515 3.735 36.601 3.875 ;
      RECT 36.465 3.732 36.515 3.875 ;
      RECT 36.455 3.73 36.465 3.874 ;
      RECT 36.451 3.73 36.455 3.873 ;
      RECT 36.365 3.725 36.451 3.868 ;
      RECT 36.343 3.718 36.365 3.862 ;
      RECT 36.257 3.709 36.343 3.856 ;
      RECT 36.171 3.696 36.257 3.847 ;
      RECT 36.085 3.682 36.171 3.837 ;
      RECT 36.04 3.672 36.085 3.83 ;
      RECT 36.02 2.96 36.04 3.238 ;
      RECT 36.02 3.665 36.04 3.826 ;
      RECT 35.99 2.96 36.02 3.26 ;
      RECT 35.98 3.632 36.02 3.823 ;
      RECT 35.975 2.96 35.99 3.28 ;
      RECT 35.975 3.597 35.98 3.821 ;
      RECT 35.97 2.96 35.975 3.405 ;
      RECT 35.97 3.557 35.975 3.821 ;
      RECT 35.96 2.96 35.97 3.821 ;
      RECT 35.885 2.96 35.96 3.815 ;
      RECT 35.855 2.96 35.885 3.805 ;
      RECT 35.85 2.96 35.855 3.797 ;
      RECT 35.845 3.002 35.85 3.79 ;
      RECT 35.835 3.071 35.845 3.781 ;
      RECT 35.83 3.141 35.835 3.733 ;
      RECT 35.825 3.205 35.83 3.63 ;
      RECT 35.82 3.24 35.825 3.585 ;
      RECT 35.818 3.277 35.82 3.477 ;
      RECT 35.815 3.285 35.818 3.47 ;
      RECT 35.81 3.35 35.815 3.413 ;
      RECT 39.885 2.44 40.165 2.72 ;
      RECT 39.875 2.44 40.165 2.583 ;
      RECT 39.83 2.305 40.09 2.565 ;
      RECT 39.83 2.42 40.145 2.565 ;
      RECT 39.83 2.39 40.14 2.565 ;
      RECT 39.83 2.377 40.13 2.565 ;
      RECT 39.83 2.367 40.125 2.565 ;
      RECT 35.805 2.35 36.065 2.61 ;
      RECT 39.575 1.9 39.835 2.16 ;
      RECT 39.565 1.925 39.835 2.12 ;
      RECT 39.56 1.925 39.565 2.119 ;
      RECT 39.49 1.92 39.56 2.111 ;
      RECT 39.405 1.907 39.49 2.094 ;
      RECT 39.401 1.899 39.405 2.084 ;
      RECT 39.315 1.892 39.401 2.074 ;
      RECT 39.306 1.884 39.315 2.064 ;
      RECT 39.22 1.877 39.306 2.052 ;
      RECT 39.2 1.868 39.22 2.038 ;
      RECT 39.145 1.863 39.2 2.03 ;
      RECT 39.135 1.857 39.145 2.024 ;
      RECT 39.115 1.855 39.135 2.02 ;
      RECT 39.107 1.854 39.115 2.016 ;
      RECT 39.021 1.846 39.107 2.005 ;
      RECT 38.935 1.832 39.021 1.985 ;
      RECT 38.875 1.82 38.935 1.97 ;
      RECT 38.865 1.815 38.875 1.965 ;
      RECT 38.815 1.815 38.865 1.967 ;
      RECT 38.768 1.817 38.815 1.971 ;
      RECT 38.682 1.824 38.768 1.976 ;
      RECT 38.596 1.832 38.682 1.982 ;
      RECT 38.51 1.841 38.596 1.988 ;
      RECT 38.451 1.847 38.51 1.993 ;
      RECT 38.365 1.852 38.451 1.999 ;
      RECT 38.29 1.857 38.365 2.005 ;
      RECT 38.251 1.859 38.29 2.01 ;
      RECT 38.165 1.856 38.251 2.015 ;
      RECT 38.08 1.854 38.165 2.022 ;
      RECT 38.048 1.853 38.08 2.025 ;
      RECT 37.962 1.852 38.048 2.026 ;
      RECT 37.876 1.851 37.962 2.027 ;
      RECT 37.79 1.85 37.876 2.027 ;
      RECT 37.704 1.849 37.79 2.028 ;
      RECT 37.618 1.848 37.704 2.029 ;
      RECT 37.532 1.847 37.618 2.03 ;
      RECT 37.446 1.846 37.532 2.03 ;
      RECT 37.36 1.845 37.446 2.031 ;
      RECT 37.31 1.845 37.36 2.032 ;
      RECT 37.296 1.846 37.31 2.032 ;
      RECT 37.21 1.853 37.296 2.033 ;
      RECT 37.136 1.864 37.21 2.034 ;
      RECT 37.05 1.873 37.136 2.035 ;
      RECT 37.015 1.88 37.05 2.05 ;
      RECT 36.99 1.883 37.015 2.08 ;
      RECT 36.965 1.892 36.99 2.109 ;
      RECT 36.955 1.903 36.965 2.129 ;
      RECT 36.945 1.911 36.955 2.143 ;
      RECT 36.94 1.917 36.945 2.153 ;
      RECT 36.915 1.934 36.94 2.17 ;
      RECT 36.9 1.956 36.915 2.198 ;
      RECT 36.87 1.982 36.9 2.228 ;
      RECT 36.85 2.011 36.87 2.258 ;
      RECT 36.845 2.026 36.85 2.275 ;
      RECT 36.825 2.041 36.845 2.29 ;
      RECT 36.815 2.059 36.825 2.308 ;
      RECT 36.805 2.07 36.815 2.323 ;
      RECT 36.755 2.102 36.805 2.349 ;
      RECT 36.75 2.132 36.755 2.369 ;
      RECT 36.74 2.145 36.75 2.375 ;
      RECT 36.731 2.155 36.74 2.383 ;
      RECT 36.72 2.166 36.731 2.391 ;
      RECT 36.715 2.176 36.72 2.397 ;
      RECT 36.7 2.197 36.715 2.404 ;
      RECT 36.685 2.227 36.7 2.412 ;
      RECT 36.65 2.257 36.685 2.418 ;
      RECT 36.625 2.275 36.65 2.425 ;
      RECT 36.575 2.283 36.625 2.434 ;
      RECT 36.55 2.288 36.575 2.443 ;
      RECT 36.495 2.294 36.55 2.453 ;
      RECT 36.49 2.299 36.495 2.461 ;
      RECT 36.476 2.302 36.49 2.463 ;
      RECT 36.39 2.314 36.476 2.475 ;
      RECT 36.38 2.326 36.39 2.488 ;
      RECT 36.295 2.339 36.38 2.5 ;
      RECT 36.251 2.356 36.295 2.514 ;
      RECT 36.165 2.373 36.251 2.53 ;
      RECT 36.135 2.387 36.165 2.544 ;
      RECT 36.125 2.392 36.135 2.549 ;
      RECT 36.065 2.395 36.125 2.558 ;
      RECT 38.955 2.665 39.215 2.925 ;
      RECT 38.955 2.665 39.235 2.778 ;
      RECT 38.955 2.665 39.26 2.745 ;
      RECT 38.955 2.665 39.265 2.725 ;
      RECT 39.005 2.44 39.285 2.72 ;
      RECT 38.56 3.175 38.82 3.435 ;
      RECT 38.55 3.032 38.745 3.373 ;
      RECT 38.545 3.14 38.76 3.365 ;
      RECT 38.54 3.19 38.82 3.355 ;
      RECT 38.53 3.267 38.82 3.34 ;
      RECT 38.55 3.115 38.76 3.373 ;
      RECT 38.56 2.99 38.745 3.435 ;
      RECT 38.56 2.885 38.725 3.435 ;
      RECT 38.57 2.872 38.725 3.435 ;
      RECT 38.57 2.83 38.715 3.435 ;
      RECT 38.575 2.755 38.715 3.435 ;
      RECT 38.605 2.405 38.715 3.435 ;
      RECT 38.61 2.135 38.735 2.758 ;
      RECT 38.58 2.71 38.735 2.758 ;
      RECT 38.595 2.512 38.715 3.435 ;
      RECT 38.585 2.622 38.735 2.758 ;
      RECT 38.61 2.135 38.75 2.615 ;
      RECT 38.61 2.135 38.77 2.49 ;
      RECT 38.575 2.135 38.835 2.395 ;
      RECT 38.045 2.44 38.325 2.72 ;
      RECT 38.03 2.44 38.325 2.7 ;
      RECT 36.085 3.305 36.345 3.565 ;
      RECT 37.87 3.16 38.13 3.42 ;
      RECT 37.85 3.18 38.13 3.395 ;
      RECT 37.807 3.18 37.85 3.394 ;
      RECT 37.721 3.181 37.807 3.391 ;
      RECT 37.635 3.182 37.721 3.387 ;
      RECT 37.56 3.184 37.635 3.384 ;
      RECT 37.537 3.185 37.56 3.382 ;
      RECT 37.451 3.186 37.537 3.38 ;
      RECT 37.365 3.187 37.451 3.377 ;
      RECT 37.341 3.188 37.365 3.375 ;
      RECT 37.255 3.19 37.341 3.372 ;
      RECT 37.17 3.192 37.255 3.373 ;
      RECT 37.113 3.193 37.17 3.379 ;
      RECT 37.027 3.195 37.113 3.389 ;
      RECT 36.941 3.198 37.027 3.402 ;
      RECT 36.855 3.2 36.941 3.414 ;
      RECT 36.841 3.201 36.855 3.421 ;
      RECT 36.755 3.202 36.841 3.429 ;
      RECT 36.715 3.204 36.755 3.438 ;
      RECT 36.706 3.205 36.715 3.441 ;
      RECT 36.62 3.213 36.706 3.447 ;
      RECT 36.6 3.222 36.62 3.455 ;
      RECT 36.515 3.237 36.6 3.463 ;
      RECT 36.455 3.26 36.515 3.474 ;
      RECT 36.445 3.272 36.455 3.479 ;
      RECT 36.405 3.282 36.445 3.483 ;
      RECT 36.35 3.299 36.405 3.491 ;
      RECT 36.345 3.309 36.35 3.495 ;
      RECT 37.411 2.44 37.47 2.837 ;
      RECT 37.325 2.44 37.53 2.828 ;
      RECT 37.32 2.47 37.53 2.823 ;
      RECT 37.286 2.47 37.53 2.821 ;
      RECT 37.2 2.47 37.53 2.815 ;
      RECT 37.155 2.47 37.55 2.793 ;
      RECT 37.155 2.47 37.57 2.748 ;
      RECT 37.115 2.47 37.57 2.738 ;
      RECT 37.325 2.44 37.605 2.72 ;
      RECT 37.06 2.44 37.32 2.7 ;
      RECT 34.885 3 35.165 3.28 ;
      RECT 34.855 2.962 35.11 3.265 ;
      RECT 34.85 2.963 35.11 3.263 ;
      RECT 34.845 2.964 35.11 3.257 ;
      RECT 34.84 2.967 35.11 3.25 ;
      RECT 34.835 3 35.165 3.243 ;
      RECT 34.805 2.97 35.11 3.23 ;
      RECT 34.805 2.997 35.13 3.23 ;
      RECT 34.805 2.987 35.125 3.23 ;
      RECT 34.805 2.972 35.12 3.23 ;
      RECT 34.885 2.959 35.1 3.28 ;
      RECT 34.971 2.957 35.1 3.28 ;
      RECT 35.057 2.955 35.085 3.28 ;
      RECT 30.7 6.22 31.02 6.545 ;
      RECT 30.73 5.695 30.9 6.545 ;
      RECT 30.73 5.695 30.905 6.045 ;
      RECT 30.73 5.695 31.705 5.87 ;
      RECT 31.53 1.965 31.705 5.87 ;
      RECT 31.475 1.965 31.825 2.315 ;
      RECT 31.5 6.655 31.825 6.98 ;
      RECT 30.385 6.745 31.825 6.915 ;
      RECT 30.385 2.395 30.545 6.915 ;
      RECT 30.7 2.365 31.02 2.685 ;
      RECT 30.385 2.395 31.02 2.565 ;
      RECT 20.47 1.92 20.73 2.18 ;
      RECT 20.525 1.88 20.83 2.16 ;
      RECT 20.525 1.42 20.7 2.18 ;
      RECT 29.04 1.34 29.39 1.69 ;
      RECT 20.525 1.42 29.39 1.595 ;
      RECT 28.715 2.85 29.085 3.22 ;
      RECT 28.8 2.235 28.97 3.22 ;
      RECT 24.82 2.455 25.055 2.715 ;
      RECT 27.965 2.235 28.13 2.495 ;
      RECT 27.87 2.225 27.885 2.495 ;
      RECT 27.965 2.235 28.97 2.415 ;
      RECT 26.47 1.795 26.51 1.935 ;
      RECT 27.885 2.23 27.965 2.495 ;
      RECT 27.83 2.225 27.87 2.461 ;
      RECT 27.816 2.225 27.83 2.461 ;
      RECT 27.73 2.23 27.816 2.463 ;
      RECT 27.685 2.237 27.73 2.465 ;
      RECT 27.655 2.237 27.685 2.467 ;
      RECT 27.63 2.232 27.655 2.469 ;
      RECT 27.6 2.228 27.63 2.478 ;
      RECT 27.59 2.225 27.6 2.49 ;
      RECT 27.585 2.225 27.59 2.498 ;
      RECT 27.58 2.225 27.585 2.503 ;
      RECT 27.57 2.224 27.58 2.513 ;
      RECT 27.565 2.223 27.57 2.523 ;
      RECT 27.55 2.222 27.565 2.528 ;
      RECT 27.522 2.219 27.55 2.555 ;
      RECT 27.436 2.211 27.522 2.555 ;
      RECT 27.35 2.2 27.436 2.555 ;
      RECT 27.31 2.185 27.35 2.555 ;
      RECT 27.27 2.159 27.31 2.555 ;
      RECT 27.265 2.141 27.27 2.367 ;
      RECT 27.255 2.137 27.265 2.357 ;
      RECT 27.24 2.127 27.255 2.344 ;
      RECT 27.22 2.111 27.24 2.329 ;
      RECT 27.205 2.096 27.22 2.314 ;
      RECT 27.195 2.085 27.205 2.304 ;
      RECT 27.17 2.069 27.195 2.293 ;
      RECT 27.165 2.056 27.17 2.283 ;
      RECT 27.16 2.052 27.165 2.278 ;
      RECT 27.105 2.038 27.16 2.256 ;
      RECT 27.066 2.019 27.105 2.22 ;
      RECT 26.98 1.993 27.066 2.173 ;
      RECT 26.976 1.975 26.98 2.139 ;
      RECT 26.89 1.956 26.976 2.117 ;
      RECT 26.885 1.938 26.89 2.095 ;
      RECT 26.88 1.936 26.885 2.093 ;
      RECT 26.87 1.935 26.88 2.088 ;
      RECT 26.81 1.922 26.87 2.074 ;
      RECT 26.765 1.9 26.81 2.053 ;
      RECT 26.705 1.877 26.765 2.032 ;
      RECT 26.641 1.852 26.705 2.007 ;
      RECT 26.555 1.822 26.641 1.976 ;
      RECT 26.54 1.802 26.555 1.955 ;
      RECT 26.51 1.797 26.54 1.946 ;
      RECT 26.457 1.795 26.47 1.935 ;
      RECT 26.371 1.795 26.457 1.937 ;
      RECT 26.285 1.795 26.371 1.939 ;
      RECT 26.265 1.795 26.285 1.943 ;
      RECT 26.22 1.797 26.265 1.954 ;
      RECT 26.18 1.807 26.22 1.97 ;
      RECT 26.176 1.816 26.18 1.978 ;
      RECT 26.09 1.836 26.176 1.994 ;
      RECT 26.08 1.855 26.09 2.012 ;
      RECT 26.075 1.857 26.08 2.015 ;
      RECT 26.065 1.861 26.075 2.018 ;
      RECT 26.045 1.866 26.065 2.028 ;
      RECT 26.015 1.876 26.045 2.048 ;
      RECT 26.01 1.883 26.015 2.062 ;
      RECT 26 1.887 26.01 2.069 ;
      RECT 25.985 1.895 26 2.08 ;
      RECT 25.975 1.905 25.985 2.091 ;
      RECT 25.965 1.912 25.975 2.099 ;
      RECT 25.94 1.925 25.965 2.114 ;
      RECT 25.876 1.961 25.94 2.153 ;
      RECT 25.79 2.024 25.876 2.217 ;
      RECT 25.755 2.075 25.79 2.27 ;
      RECT 25.75 2.092 25.755 2.287 ;
      RECT 25.735 2.101 25.75 2.294 ;
      RECT 25.715 2.116 25.735 2.308 ;
      RECT 25.71 2.127 25.715 2.318 ;
      RECT 25.69 2.14 25.71 2.328 ;
      RECT 25.685 2.15 25.69 2.338 ;
      RECT 25.67 2.155 25.685 2.347 ;
      RECT 25.66 2.165 25.67 2.358 ;
      RECT 25.63 2.182 25.66 2.375 ;
      RECT 25.62 2.2 25.63 2.393 ;
      RECT 25.605 2.211 25.62 2.404 ;
      RECT 25.565 2.235 25.605 2.42 ;
      RECT 25.53 2.269 25.565 2.437 ;
      RECT 25.5 2.292 25.53 2.449 ;
      RECT 25.485 2.302 25.5 2.458 ;
      RECT 25.445 2.312 25.485 2.469 ;
      RECT 25.425 2.323 25.445 2.481 ;
      RECT 25.42 2.327 25.425 2.488 ;
      RECT 25.405 2.331 25.42 2.493 ;
      RECT 25.395 2.336 25.405 2.498 ;
      RECT 25.39 2.339 25.395 2.501 ;
      RECT 25.36 2.345 25.39 2.508 ;
      RECT 25.325 2.355 25.36 2.522 ;
      RECT 25.265 2.37 25.325 2.542 ;
      RECT 25.21 2.39 25.265 2.566 ;
      RECT 25.181 2.405 25.21 2.584 ;
      RECT 25.095 2.425 25.181 2.609 ;
      RECT 25.09 2.44 25.095 2.629 ;
      RECT 25.08 2.443 25.09 2.63 ;
      RECT 25.055 2.45 25.08 2.715 ;
      RECT 27.75 2.943 28.03 3.28 ;
      RECT 27.75 2.953 28.035 3.238 ;
      RECT 27.75 2.962 28.04 3.135 ;
      RECT 27.75 2.977 28.045 3.003 ;
      RECT 27.75 2.805 28.01 3.28 ;
      RECT 18.1 6.655 18.45 7.005 ;
      RECT 26.925 6.61 27.275 6.96 ;
      RECT 18.1 6.685 27.275 6.885 ;
      RECT 25.47 3.685 25.48 3.875 ;
      RECT 23.73 3.56 24.01 3.84 ;
      RECT 26.775 2.5 26.78 2.985 ;
      RECT 26.67 2.5 26.73 2.76 ;
      RECT 26.995 3.47 27 3.545 ;
      RECT 26.985 3.337 26.995 3.58 ;
      RECT 26.975 3.172 26.985 3.601 ;
      RECT 26.97 3.042 26.975 3.617 ;
      RECT 26.96 2.932 26.97 3.633 ;
      RECT 26.955 2.831 26.96 3.65 ;
      RECT 26.95 2.813 26.955 3.66 ;
      RECT 26.945 2.795 26.95 3.67 ;
      RECT 26.935 2.77 26.945 3.685 ;
      RECT 26.93 2.75 26.935 3.7 ;
      RECT 26.91 2.5 26.93 3.725 ;
      RECT 26.895 2.5 26.91 3.758 ;
      RECT 26.865 2.5 26.895 3.78 ;
      RECT 26.845 2.5 26.865 3.794 ;
      RECT 26.825 2.5 26.845 3.31 ;
      RECT 26.84 3.377 26.845 3.799 ;
      RECT 26.835 3.407 26.84 3.801 ;
      RECT 26.83 3.42 26.835 3.804 ;
      RECT 26.825 3.43 26.83 3.808 ;
      RECT 26.82 2.5 26.825 3.228 ;
      RECT 26.82 3.44 26.825 3.81 ;
      RECT 26.815 2.5 26.82 3.205 ;
      RECT 26.805 3.462 26.82 3.81 ;
      RECT 26.8 2.5 26.815 3.15 ;
      RECT 26.795 3.487 26.805 3.81 ;
      RECT 26.795 2.5 26.8 3.095 ;
      RECT 26.785 2.5 26.795 3.043 ;
      RECT 26.79 3.5 26.795 3.811 ;
      RECT 26.785 3.512 26.79 3.812 ;
      RECT 26.78 2.5 26.785 3.003 ;
      RECT 26.78 3.525 26.785 3.813 ;
      RECT 26.765 3.54 26.78 3.814 ;
      RECT 26.77 2.5 26.775 2.965 ;
      RECT 26.765 2.5 26.77 2.93 ;
      RECT 26.76 2.5 26.765 2.905 ;
      RECT 26.755 3.567 26.765 3.816 ;
      RECT 26.75 2.5 26.76 2.863 ;
      RECT 26.75 3.585 26.755 3.817 ;
      RECT 26.745 2.5 26.75 2.823 ;
      RECT 26.745 3.592 26.75 3.818 ;
      RECT 26.74 2.5 26.745 2.795 ;
      RECT 26.735 3.61 26.745 3.819 ;
      RECT 26.73 2.5 26.74 2.775 ;
      RECT 26.725 3.63 26.735 3.821 ;
      RECT 26.715 3.647 26.725 3.822 ;
      RECT 26.68 3.67 26.715 3.825 ;
      RECT 26.625 3.688 26.68 3.831 ;
      RECT 26.539 3.696 26.625 3.84 ;
      RECT 26.453 3.707 26.539 3.851 ;
      RECT 26.367 3.717 26.453 3.862 ;
      RECT 26.281 3.727 26.367 3.874 ;
      RECT 26.195 3.737 26.281 3.885 ;
      RECT 26.175 3.743 26.195 3.891 ;
      RECT 26.095 3.745 26.175 3.895 ;
      RECT 26.09 3.744 26.095 3.9 ;
      RECT 26.082 3.743 26.09 3.9 ;
      RECT 25.996 3.739 26.082 3.898 ;
      RECT 25.91 3.731 25.996 3.895 ;
      RECT 25.824 3.722 25.91 3.891 ;
      RECT 25.738 3.714 25.824 3.888 ;
      RECT 25.652 3.706 25.738 3.884 ;
      RECT 25.566 3.697 25.652 3.881 ;
      RECT 25.48 3.689 25.566 3.877 ;
      RECT 25.425 3.682 25.47 3.875 ;
      RECT 25.34 3.675 25.425 3.873 ;
      RECT 25.266 3.667 25.34 3.869 ;
      RECT 25.18 3.659 25.266 3.866 ;
      RECT 25.177 3.655 25.18 3.864 ;
      RECT 25.091 3.651 25.177 3.863 ;
      RECT 25.005 3.643 25.091 3.86 ;
      RECT 24.92 3.638 25.005 3.857 ;
      RECT 24.834 3.635 24.92 3.854 ;
      RECT 24.748 3.633 24.834 3.851 ;
      RECT 24.662 3.63 24.748 3.848 ;
      RECT 24.576 3.627 24.662 3.845 ;
      RECT 24.49 3.624 24.576 3.842 ;
      RECT 24.414 3.622 24.49 3.839 ;
      RECT 24.328 3.619 24.414 3.836 ;
      RECT 24.242 3.616 24.328 3.834 ;
      RECT 24.156 3.614 24.242 3.831 ;
      RECT 24.07 3.611 24.156 3.828 ;
      RECT 24.01 3.602 24.07 3.826 ;
      RECT 26.52 3.22 26.595 3.48 ;
      RECT 26.5 3.2 26.505 3.48 ;
      RECT 25.82 2.985 25.925 3.28 ;
      RECT 20.265 2.96 20.335 3.22 ;
      RECT 26.16 2.835 26.165 3.206 ;
      RECT 26.15 2.89 26.155 3.206 ;
      RECT 26.455 2.06 26.515 2.32 ;
      RECT 26.51 3.215 26.52 3.48 ;
      RECT 26.505 3.205 26.51 3.48 ;
      RECT 26.425 3.152 26.5 3.48 ;
      RECT 26.45 2.06 26.455 2.34 ;
      RECT 26.44 2.06 26.45 2.36 ;
      RECT 26.425 2.06 26.44 2.39 ;
      RECT 26.41 2.06 26.425 2.433 ;
      RECT 26.405 3.095 26.425 3.48 ;
      RECT 26.395 2.06 26.41 2.47 ;
      RECT 26.39 3.075 26.405 3.48 ;
      RECT 26.39 2.06 26.395 2.493 ;
      RECT 26.38 2.06 26.39 2.518 ;
      RECT 26.35 3.042 26.39 3.48 ;
      RECT 26.355 2.06 26.38 2.568 ;
      RECT 26.35 2.06 26.355 2.623 ;
      RECT 26.345 2.06 26.35 2.665 ;
      RECT 26.335 3.005 26.35 3.48 ;
      RECT 26.34 2.06 26.345 2.708 ;
      RECT 26.335 2.06 26.34 2.773 ;
      RECT 26.33 2.06 26.335 2.795 ;
      RECT 26.33 2.993 26.335 3.345 ;
      RECT 26.325 2.06 26.33 2.863 ;
      RECT 26.325 2.985 26.33 3.328 ;
      RECT 26.32 2.06 26.325 2.908 ;
      RECT 26.315 2.967 26.325 3.305 ;
      RECT 26.315 2.06 26.32 2.945 ;
      RECT 26.305 2.06 26.315 3.285 ;
      RECT 26.3 2.06 26.305 3.268 ;
      RECT 26.295 2.06 26.3 3.253 ;
      RECT 26.29 2.06 26.295 3.238 ;
      RECT 26.27 2.06 26.29 3.228 ;
      RECT 26.265 2.06 26.27 3.218 ;
      RECT 26.255 2.06 26.265 3.214 ;
      RECT 26.25 2.337 26.255 3.213 ;
      RECT 26.245 2.36 26.25 3.212 ;
      RECT 26.24 2.39 26.245 3.211 ;
      RECT 26.235 2.417 26.24 3.21 ;
      RECT 26.23 2.445 26.235 3.21 ;
      RECT 26.225 2.472 26.23 3.21 ;
      RECT 26.22 2.492 26.225 3.21 ;
      RECT 26.215 2.52 26.22 3.21 ;
      RECT 26.205 2.562 26.215 3.21 ;
      RECT 26.195 2.607 26.205 3.209 ;
      RECT 26.19 2.66 26.195 3.208 ;
      RECT 26.185 2.692 26.19 3.207 ;
      RECT 26.18 2.712 26.185 3.206 ;
      RECT 26.175 2.75 26.18 3.206 ;
      RECT 26.17 2.772 26.175 3.206 ;
      RECT 26.165 2.797 26.17 3.206 ;
      RECT 26.155 2.862 26.16 3.206 ;
      RECT 26.14 2.922 26.15 3.206 ;
      RECT 26.125 2.932 26.14 3.206 ;
      RECT 26.105 2.942 26.125 3.206 ;
      RECT 26.075 2.947 26.105 3.203 ;
      RECT 26.015 2.957 26.075 3.2 ;
      RECT 25.995 2.966 26.015 3.205 ;
      RECT 25.97 2.972 25.995 3.218 ;
      RECT 25.95 2.977 25.97 3.233 ;
      RECT 25.925 2.982 25.95 3.28 ;
      RECT 25.796 2.984 25.82 3.28 ;
      RECT 25.71 2.979 25.796 3.28 ;
      RECT 25.67 2.976 25.71 3.28 ;
      RECT 25.62 2.978 25.67 3.26 ;
      RECT 25.59 2.982 25.62 3.26 ;
      RECT 25.511 2.992 25.59 3.26 ;
      RECT 25.425 3.007 25.511 3.261 ;
      RECT 25.375 3.017 25.425 3.262 ;
      RECT 25.367 3.02 25.375 3.262 ;
      RECT 25.281 3.022 25.367 3.263 ;
      RECT 25.195 3.026 25.281 3.263 ;
      RECT 25.109 3.03 25.195 3.264 ;
      RECT 25.023 3.033 25.109 3.265 ;
      RECT 24.937 3.037 25.023 3.265 ;
      RECT 24.851 3.041 24.937 3.266 ;
      RECT 24.765 3.044 24.851 3.267 ;
      RECT 24.679 3.048 24.765 3.267 ;
      RECT 24.593 3.052 24.679 3.268 ;
      RECT 24.507 3.056 24.593 3.269 ;
      RECT 24.421 3.059 24.507 3.269 ;
      RECT 24.335 3.063 24.421 3.27 ;
      RECT 24.305 3.065 24.335 3.27 ;
      RECT 24.219 3.068 24.305 3.271 ;
      RECT 24.133 3.072 24.219 3.272 ;
      RECT 24.047 3.076 24.133 3.273 ;
      RECT 23.961 3.079 24.047 3.273 ;
      RECT 23.875 3.083 23.961 3.274 ;
      RECT 23.84 3.088 23.875 3.275 ;
      RECT 23.785 3.098 23.84 3.282 ;
      RECT 23.76 3.11 23.785 3.292 ;
      RECT 23.725 3.123 23.76 3.3 ;
      RECT 23.685 3.14 23.725 3.323 ;
      RECT 23.665 3.153 23.685 3.35 ;
      RECT 23.635 3.165 23.665 3.378 ;
      RECT 23.63 3.173 23.635 3.398 ;
      RECT 23.625 3.176 23.63 3.408 ;
      RECT 23.575 3.188 23.625 3.442 ;
      RECT 23.565 3.203 23.575 3.475 ;
      RECT 23.555 3.209 23.565 3.488 ;
      RECT 23.545 3.216 23.555 3.5 ;
      RECT 23.52 3.229 23.545 3.518 ;
      RECT 23.505 3.244 23.52 3.54 ;
      RECT 23.495 3.252 23.505 3.556 ;
      RECT 23.48 3.261 23.495 3.571 ;
      RECT 23.47 3.271 23.48 3.585 ;
      RECT 23.451 3.284 23.47 3.602 ;
      RECT 23.365 3.329 23.451 3.667 ;
      RECT 23.35 3.374 23.365 3.725 ;
      RECT 23.345 3.383 23.35 3.738 ;
      RECT 23.335 3.39 23.345 3.743 ;
      RECT 23.33 3.395 23.335 3.747 ;
      RECT 23.31 3.405 23.33 3.754 ;
      RECT 23.285 3.425 23.31 3.768 ;
      RECT 23.25 3.45 23.285 3.788 ;
      RECT 23.235 3.473 23.25 3.803 ;
      RECT 23.225 3.483 23.235 3.808 ;
      RECT 23.215 3.491 23.225 3.815 ;
      RECT 23.205 3.5 23.215 3.821 ;
      RECT 23.185 3.512 23.205 3.823 ;
      RECT 23.175 3.525 23.185 3.825 ;
      RECT 23.15 3.54 23.175 3.828 ;
      RECT 23.13 3.557 23.15 3.832 ;
      RECT 23.09 3.585 23.13 3.838 ;
      RECT 23.025 3.632 23.09 3.847 ;
      RECT 23.01 3.665 23.025 3.855 ;
      RECT 23.005 3.672 23.01 3.857 ;
      RECT 22.955 3.697 23.005 3.862 ;
      RECT 22.94 3.721 22.955 3.869 ;
      RECT 22.89 3.726 22.94 3.87 ;
      RECT 22.804 3.73 22.89 3.87 ;
      RECT 22.718 3.73 22.804 3.87 ;
      RECT 22.632 3.73 22.718 3.871 ;
      RECT 22.546 3.73 22.632 3.871 ;
      RECT 22.46 3.73 22.546 3.871 ;
      RECT 22.394 3.73 22.46 3.871 ;
      RECT 22.308 3.73 22.394 3.872 ;
      RECT 22.222 3.73 22.308 3.872 ;
      RECT 22.136 3.731 22.222 3.873 ;
      RECT 22.05 3.731 22.136 3.873 ;
      RECT 21.964 3.731 22.05 3.873 ;
      RECT 21.878 3.731 21.964 3.874 ;
      RECT 21.792 3.731 21.878 3.874 ;
      RECT 21.706 3.732 21.792 3.875 ;
      RECT 21.62 3.732 21.706 3.875 ;
      RECT 21.6 3.732 21.62 3.875 ;
      RECT 21.514 3.732 21.6 3.875 ;
      RECT 21.428 3.732 21.514 3.875 ;
      RECT 21.342 3.733 21.428 3.875 ;
      RECT 21.256 3.733 21.342 3.875 ;
      RECT 21.17 3.733 21.256 3.875 ;
      RECT 21.084 3.734 21.17 3.875 ;
      RECT 20.998 3.734 21.084 3.875 ;
      RECT 20.912 3.734 20.998 3.875 ;
      RECT 20.826 3.734 20.912 3.875 ;
      RECT 20.74 3.735 20.826 3.875 ;
      RECT 20.69 3.732 20.74 3.875 ;
      RECT 20.68 3.73 20.69 3.874 ;
      RECT 20.676 3.73 20.68 3.873 ;
      RECT 20.59 3.725 20.676 3.868 ;
      RECT 20.568 3.718 20.59 3.862 ;
      RECT 20.482 3.709 20.568 3.856 ;
      RECT 20.396 3.696 20.482 3.847 ;
      RECT 20.31 3.682 20.396 3.837 ;
      RECT 20.265 3.672 20.31 3.83 ;
      RECT 20.245 2.96 20.265 3.238 ;
      RECT 20.245 3.665 20.265 3.826 ;
      RECT 20.215 2.96 20.245 3.26 ;
      RECT 20.205 3.632 20.245 3.823 ;
      RECT 20.2 2.96 20.215 3.28 ;
      RECT 20.2 3.597 20.205 3.821 ;
      RECT 20.195 2.96 20.2 3.405 ;
      RECT 20.195 3.557 20.2 3.821 ;
      RECT 20.185 2.96 20.195 3.821 ;
      RECT 20.11 2.96 20.185 3.815 ;
      RECT 20.08 2.96 20.11 3.805 ;
      RECT 20.075 2.96 20.08 3.797 ;
      RECT 20.07 3.002 20.075 3.79 ;
      RECT 20.06 3.071 20.07 3.781 ;
      RECT 20.055 3.141 20.06 3.733 ;
      RECT 20.05 3.205 20.055 3.63 ;
      RECT 20.045 3.24 20.05 3.585 ;
      RECT 20.043 3.277 20.045 3.477 ;
      RECT 20.04 3.285 20.043 3.47 ;
      RECT 20.035 3.35 20.04 3.413 ;
      RECT 24.11 2.44 24.39 2.72 ;
      RECT 24.1 2.44 24.39 2.583 ;
      RECT 24.055 2.305 24.315 2.565 ;
      RECT 24.055 2.42 24.37 2.565 ;
      RECT 24.055 2.39 24.365 2.565 ;
      RECT 24.055 2.377 24.355 2.565 ;
      RECT 24.055 2.367 24.35 2.565 ;
      RECT 20.03 2.35 20.29 2.61 ;
      RECT 23.8 1.9 24.06 2.16 ;
      RECT 23.79 1.925 24.06 2.12 ;
      RECT 23.785 1.925 23.79 2.119 ;
      RECT 23.715 1.92 23.785 2.111 ;
      RECT 23.63 1.907 23.715 2.094 ;
      RECT 23.626 1.899 23.63 2.084 ;
      RECT 23.54 1.892 23.626 2.074 ;
      RECT 23.531 1.884 23.54 2.064 ;
      RECT 23.445 1.877 23.531 2.052 ;
      RECT 23.425 1.868 23.445 2.038 ;
      RECT 23.37 1.863 23.425 2.03 ;
      RECT 23.36 1.857 23.37 2.024 ;
      RECT 23.34 1.855 23.36 2.02 ;
      RECT 23.332 1.854 23.34 2.016 ;
      RECT 23.246 1.846 23.332 2.005 ;
      RECT 23.16 1.832 23.246 1.985 ;
      RECT 23.1 1.82 23.16 1.97 ;
      RECT 23.09 1.815 23.1 1.965 ;
      RECT 23.04 1.815 23.09 1.967 ;
      RECT 22.993 1.817 23.04 1.971 ;
      RECT 22.907 1.824 22.993 1.976 ;
      RECT 22.821 1.832 22.907 1.982 ;
      RECT 22.735 1.841 22.821 1.988 ;
      RECT 22.676 1.847 22.735 1.993 ;
      RECT 22.59 1.852 22.676 1.999 ;
      RECT 22.515 1.857 22.59 2.005 ;
      RECT 22.476 1.859 22.515 2.01 ;
      RECT 22.39 1.856 22.476 2.015 ;
      RECT 22.305 1.854 22.39 2.022 ;
      RECT 22.273 1.853 22.305 2.025 ;
      RECT 22.187 1.852 22.273 2.026 ;
      RECT 22.101 1.851 22.187 2.027 ;
      RECT 22.015 1.85 22.101 2.027 ;
      RECT 21.929 1.849 22.015 2.028 ;
      RECT 21.843 1.848 21.929 2.029 ;
      RECT 21.757 1.847 21.843 2.03 ;
      RECT 21.671 1.846 21.757 2.03 ;
      RECT 21.585 1.845 21.671 2.031 ;
      RECT 21.535 1.845 21.585 2.032 ;
      RECT 21.521 1.846 21.535 2.032 ;
      RECT 21.435 1.853 21.521 2.033 ;
      RECT 21.361 1.864 21.435 2.034 ;
      RECT 21.275 1.873 21.361 2.035 ;
      RECT 21.24 1.88 21.275 2.05 ;
      RECT 21.215 1.883 21.24 2.08 ;
      RECT 21.19 1.892 21.215 2.109 ;
      RECT 21.18 1.903 21.19 2.129 ;
      RECT 21.17 1.911 21.18 2.143 ;
      RECT 21.165 1.917 21.17 2.153 ;
      RECT 21.14 1.934 21.165 2.17 ;
      RECT 21.125 1.956 21.14 2.198 ;
      RECT 21.095 1.982 21.125 2.228 ;
      RECT 21.075 2.011 21.095 2.258 ;
      RECT 21.07 2.026 21.075 2.275 ;
      RECT 21.05 2.041 21.07 2.29 ;
      RECT 21.04 2.059 21.05 2.308 ;
      RECT 21.03 2.07 21.04 2.323 ;
      RECT 20.98 2.102 21.03 2.349 ;
      RECT 20.975 2.132 20.98 2.369 ;
      RECT 20.965 2.145 20.975 2.375 ;
      RECT 20.956 2.155 20.965 2.383 ;
      RECT 20.945 2.166 20.956 2.391 ;
      RECT 20.94 2.176 20.945 2.397 ;
      RECT 20.925 2.197 20.94 2.404 ;
      RECT 20.91 2.227 20.925 2.412 ;
      RECT 20.875 2.257 20.91 2.418 ;
      RECT 20.85 2.275 20.875 2.425 ;
      RECT 20.8 2.283 20.85 2.434 ;
      RECT 20.775 2.288 20.8 2.443 ;
      RECT 20.72 2.294 20.775 2.453 ;
      RECT 20.715 2.299 20.72 2.461 ;
      RECT 20.701 2.302 20.715 2.463 ;
      RECT 20.615 2.314 20.701 2.475 ;
      RECT 20.605 2.326 20.615 2.488 ;
      RECT 20.52 2.339 20.605 2.5 ;
      RECT 20.476 2.356 20.52 2.514 ;
      RECT 20.39 2.373 20.476 2.53 ;
      RECT 20.36 2.387 20.39 2.544 ;
      RECT 20.35 2.392 20.36 2.549 ;
      RECT 20.29 2.395 20.35 2.558 ;
      RECT 23.18 2.665 23.44 2.925 ;
      RECT 23.18 2.665 23.46 2.778 ;
      RECT 23.18 2.665 23.485 2.745 ;
      RECT 23.18 2.665 23.49 2.725 ;
      RECT 23.23 2.44 23.51 2.72 ;
      RECT 22.785 3.175 23.045 3.435 ;
      RECT 22.775 3.032 22.97 3.373 ;
      RECT 22.77 3.14 22.985 3.365 ;
      RECT 22.765 3.19 23.045 3.355 ;
      RECT 22.755 3.267 23.045 3.34 ;
      RECT 22.775 3.115 22.985 3.373 ;
      RECT 22.785 2.99 22.97 3.435 ;
      RECT 22.785 2.885 22.95 3.435 ;
      RECT 22.795 2.872 22.95 3.435 ;
      RECT 22.795 2.83 22.94 3.435 ;
      RECT 22.8 2.755 22.94 3.435 ;
      RECT 22.83 2.405 22.94 3.435 ;
      RECT 22.835 2.135 22.96 2.758 ;
      RECT 22.805 2.71 22.96 2.758 ;
      RECT 22.82 2.512 22.94 3.435 ;
      RECT 22.81 2.622 22.96 2.758 ;
      RECT 22.835 2.135 22.975 2.615 ;
      RECT 22.835 2.135 22.995 2.49 ;
      RECT 22.8 2.135 23.06 2.395 ;
      RECT 22.27 2.44 22.55 2.72 ;
      RECT 22.255 2.44 22.55 2.7 ;
      RECT 20.31 3.305 20.57 3.565 ;
      RECT 22.095 3.16 22.355 3.42 ;
      RECT 22.075 3.18 22.355 3.395 ;
      RECT 22.032 3.18 22.075 3.394 ;
      RECT 21.946 3.181 22.032 3.391 ;
      RECT 21.86 3.182 21.946 3.387 ;
      RECT 21.785 3.184 21.86 3.384 ;
      RECT 21.762 3.185 21.785 3.382 ;
      RECT 21.676 3.186 21.762 3.38 ;
      RECT 21.59 3.187 21.676 3.377 ;
      RECT 21.566 3.188 21.59 3.375 ;
      RECT 21.48 3.19 21.566 3.372 ;
      RECT 21.395 3.192 21.48 3.373 ;
      RECT 21.338 3.193 21.395 3.379 ;
      RECT 21.252 3.195 21.338 3.389 ;
      RECT 21.166 3.198 21.252 3.402 ;
      RECT 21.08 3.2 21.166 3.414 ;
      RECT 21.066 3.201 21.08 3.421 ;
      RECT 20.98 3.202 21.066 3.429 ;
      RECT 20.94 3.204 20.98 3.438 ;
      RECT 20.931 3.205 20.94 3.441 ;
      RECT 20.845 3.213 20.931 3.447 ;
      RECT 20.825 3.222 20.845 3.455 ;
      RECT 20.74 3.237 20.825 3.463 ;
      RECT 20.68 3.26 20.74 3.474 ;
      RECT 20.67 3.272 20.68 3.479 ;
      RECT 20.63 3.282 20.67 3.483 ;
      RECT 20.575 3.299 20.63 3.491 ;
      RECT 20.57 3.309 20.575 3.495 ;
      RECT 21.636 2.44 21.695 2.837 ;
      RECT 21.55 2.44 21.755 2.828 ;
      RECT 21.545 2.47 21.755 2.823 ;
      RECT 21.511 2.47 21.755 2.821 ;
      RECT 21.425 2.47 21.755 2.815 ;
      RECT 21.38 2.47 21.775 2.793 ;
      RECT 21.38 2.47 21.795 2.748 ;
      RECT 21.34 2.47 21.795 2.738 ;
      RECT 21.55 2.44 21.83 2.72 ;
      RECT 21.285 2.44 21.545 2.7 ;
      RECT 19.11 3 19.39 3.28 ;
      RECT 19.08 2.962 19.335 3.265 ;
      RECT 19.075 2.963 19.335 3.263 ;
      RECT 19.07 2.964 19.335 3.257 ;
      RECT 19.065 2.967 19.335 3.25 ;
      RECT 19.06 3 19.39 3.243 ;
      RECT 19.03 2.97 19.335 3.23 ;
      RECT 19.03 2.997 19.355 3.23 ;
      RECT 19.03 2.987 19.35 3.23 ;
      RECT 19.03 2.972 19.345 3.23 ;
      RECT 19.11 2.959 19.325 3.28 ;
      RECT 19.196 2.957 19.325 3.28 ;
      RECT 19.282 2.955 19.31 3.28 ;
      RECT 14.92 6.22 15.24 6.545 ;
      RECT 14.95 5.695 15.12 6.545 ;
      RECT 14.95 5.695 15.125 6.045 ;
      RECT 14.95 5.695 15.925 5.87 ;
      RECT 15.75 1.965 15.925 5.87 ;
      RECT 15.695 1.965 16.045 2.315 ;
      RECT 15.72 6.655 16.045 6.98 ;
      RECT 14.605 6.745 16.045 6.915 ;
      RECT 14.605 2.395 14.765 6.915 ;
      RECT 14.92 2.365 15.24 2.685 ;
      RECT 14.605 2.395 15.24 2.565 ;
      RECT 4.69 1.92 4.95 2.18 ;
      RECT 4.745 1.88 5.05 2.16 ;
      RECT 4.745 1.42 4.92 2.18 ;
      RECT 13.26 1.34 13.61 1.69 ;
      RECT 4.745 1.42 13.61 1.595 ;
      RECT 12.935 2.85 13.305 3.22 ;
      RECT 13.02 2.235 13.19 3.22 ;
      RECT 9.04 2.455 9.275 2.715 ;
      RECT 12.185 2.235 12.35 2.495 ;
      RECT 12.09 2.225 12.105 2.495 ;
      RECT 12.185 2.235 13.19 2.415 ;
      RECT 10.69 1.795 10.73 1.935 ;
      RECT 12.105 2.23 12.185 2.495 ;
      RECT 12.05 2.225 12.09 2.461 ;
      RECT 12.036 2.225 12.05 2.461 ;
      RECT 11.95 2.23 12.036 2.463 ;
      RECT 11.905 2.237 11.95 2.465 ;
      RECT 11.875 2.237 11.905 2.467 ;
      RECT 11.85 2.232 11.875 2.469 ;
      RECT 11.82 2.228 11.85 2.478 ;
      RECT 11.81 2.225 11.82 2.49 ;
      RECT 11.805 2.225 11.81 2.498 ;
      RECT 11.8 2.225 11.805 2.503 ;
      RECT 11.79 2.224 11.8 2.513 ;
      RECT 11.785 2.223 11.79 2.523 ;
      RECT 11.77 2.222 11.785 2.528 ;
      RECT 11.742 2.219 11.77 2.555 ;
      RECT 11.656 2.211 11.742 2.555 ;
      RECT 11.57 2.2 11.656 2.555 ;
      RECT 11.53 2.185 11.57 2.555 ;
      RECT 11.49 2.159 11.53 2.555 ;
      RECT 11.485 2.141 11.49 2.367 ;
      RECT 11.475 2.137 11.485 2.357 ;
      RECT 11.46 2.127 11.475 2.344 ;
      RECT 11.44 2.111 11.46 2.329 ;
      RECT 11.425 2.096 11.44 2.314 ;
      RECT 11.415 2.085 11.425 2.304 ;
      RECT 11.39 2.069 11.415 2.293 ;
      RECT 11.385 2.056 11.39 2.283 ;
      RECT 11.38 2.052 11.385 2.278 ;
      RECT 11.325 2.038 11.38 2.256 ;
      RECT 11.286 2.019 11.325 2.22 ;
      RECT 11.2 1.993 11.286 2.173 ;
      RECT 11.196 1.975 11.2 2.139 ;
      RECT 11.11 1.956 11.196 2.117 ;
      RECT 11.105 1.938 11.11 2.095 ;
      RECT 11.1 1.936 11.105 2.093 ;
      RECT 11.09 1.935 11.1 2.088 ;
      RECT 11.03 1.922 11.09 2.074 ;
      RECT 10.985 1.9 11.03 2.053 ;
      RECT 10.925 1.877 10.985 2.032 ;
      RECT 10.861 1.852 10.925 2.007 ;
      RECT 10.775 1.822 10.861 1.976 ;
      RECT 10.76 1.802 10.775 1.955 ;
      RECT 10.73 1.797 10.76 1.946 ;
      RECT 10.677 1.795 10.69 1.935 ;
      RECT 10.591 1.795 10.677 1.937 ;
      RECT 10.505 1.795 10.591 1.939 ;
      RECT 10.485 1.795 10.505 1.943 ;
      RECT 10.44 1.797 10.485 1.954 ;
      RECT 10.4 1.807 10.44 1.97 ;
      RECT 10.396 1.816 10.4 1.978 ;
      RECT 10.31 1.836 10.396 1.994 ;
      RECT 10.3 1.855 10.31 2.012 ;
      RECT 10.295 1.857 10.3 2.015 ;
      RECT 10.285 1.861 10.295 2.018 ;
      RECT 10.265 1.866 10.285 2.028 ;
      RECT 10.235 1.876 10.265 2.048 ;
      RECT 10.23 1.883 10.235 2.062 ;
      RECT 10.22 1.887 10.23 2.069 ;
      RECT 10.205 1.895 10.22 2.08 ;
      RECT 10.195 1.905 10.205 2.091 ;
      RECT 10.185 1.912 10.195 2.099 ;
      RECT 10.16 1.925 10.185 2.114 ;
      RECT 10.096 1.961 10.16 2.153 ;
      RECT 10.01 2.024 10.096 2.217 ;
      RECT 9.975 2.075 10.01 2.27 ;
      RECT 9.97 2.092 9.975 2.287 ;
      RECT 9.955 2.101 9.97 2.294 ;
      RECT 9.935 2.116 9.955 2.308 ;
      RECT 9.93 2.127 9.935 2.318 ;
      RECT 9.91 2.14 9.93 2.328 ;
      RECT 9.905 2.15 9.91 2.338 ;
      RECT 9.89 2.155 9.905 2.347 ;
      RECT 9.88 2.165 9.89 2.358 ;
      RECT 9.85 2.182 9.88 2.375 ;
      RECT 9.84 2.2 9.85 2.393 ;
      RECT 9.825 2.211 9.84 2.404 ;
      RECT 9.785 2.235 9.825 2.42 ;
      RECT 9.75 2.269 9.785 2.437 ;
      RECT 9.72 2.292 9.75 2.449 ;
      RECT 9.705 2.302 9.72 2.458 ;
      RECT 9.665 2.312 9.705 2.469 ;
      RECT 9.645 2.323 9.665 2.481 ;
      RECT 9.64 2.327 9.645 2.488 ;
      RECT 9.625 2.331 9.64 2.493 ;
      RECT 9.615 2.336 9.625 2.498 ;
      RECT 9.61 2.339 9.615 2.501 ;
      RECT 9.58 2.345 9.61 2.508 ;
      RECT 9.545 2.355 9.58 2.522 ;
      RECT 9.485 2.37 9.545 2.542 ;
      RECT 9.43 2.39 9.485 2.566 ;
      RECT 9.401 2.405 9.43 2.584 ;
      RECT 9.315 2.425 9.401 2.609 ;
      RECT 9.31 2.44 9.315 2.629 ;
      RECT 9.3 2.443 9.31 2.63 ;
      RECT 9.275 2.45 9.3 2.715 ;
      RECT 11.97 2.943 12.25 3.28 ;
      RECT 11.97 2.953 12.255 3.238 ;
      RECT 11.97 2.962 12.26 3.135 ;
      RECT 11.97 2.977 12.265 3.003 ;
      RECT 11.97 2.805 12.23 3.28 ;
      RECT 1.55 6.995 1.84 7.345 ;
      RECT 1.55 7.085 2.955 7.255 ;
      RECT 2.785 6.685 2.955 7.255 ;
      RECT 11.115 6.605 11.465 6.955 ;
      RECT 2.785 6.685 11.465 6.855 ;
      RECT 9.69 3.685 9.7 3.875 ;
      RECT 7.95 3.56 8.23 3.84 ;
      RECT 10.995 2.5 11 2.985 ;
      RECT 10.89 2.5 10.95 2.76 ;
      RECT 11.215 3.47 11.22 3.545 ;
      RECT 11.205 3.337 11.215 3.58 ;
      RECT 11.195 3.172 11.205 3.601 ;
      RECT 11.19 3.042 11.195 3.617 ;
      RECT 11.18 2.932 11.19 3.633 ;
      RECT 11.175 2.831 11.18 3.65 ;
      RECT 11.17 2.813 11.175 3.66 ;
      RECT 11.165 2.795 11.17 3.67 ;
      RECT 11.155 2.77 11.165 3.685 ;
      RECT 11.15 2.75 11.155 3.7 ;
      RECT 11.13 2.5 11.15 3.725 ;
      RECT 11.115 2.5 11.13 3.758 ;
      RECT 11.085 2.5 11.115 3.78 ;
      RECT 11.065 2.5 11.085 3.794 ;
      RECT 11.045 2.5 11.065 3.31 ;
      RECT 11.06 3.377 11.065 3.799 ;
      RECT 11.055 3.407 11.06 3.801 ;
      RECT 11.05 3.42 11.055 3.804 ;
      RECT 11.045 3.43 11.05 3.808 ;
      RECT 11.04 2.5 11.045 3.228 ;
      RECT 11.04 3.44 11.045 3.81 ;
      RECT 11.035 2.5 11.04 3.205 ;
      RECT 11.025 3.462 11.04 3.81 ;
      RECT 11.02 2.5 11.035 3.15 ;
      RECT 11.015 3.487 11.025 3.81 ;
      RECT 11.015 2.5 11.02 3.095 ;
      RECT 11.005 2.5 11.015 3.043 ;
      RECT 11.01 3.5 11.015 3.811 ;
      RECT 11.005 3.512 11.01 3.812 ;
      RECT 11 2.5 11.005 3.003 ;
      RECT 11 3.525 11.005 3.813 ;
      RECT 10.985 3.54 11 3.814 ;
      RECT 10.99 2.5 10.995 2.965 ;
      RECT 10.985 2.5 10.99 2.93 ;
      RECT 10.98 2.5 10.985 2.905 ;
      RECT 10.975 3.567 10.985 3.816 ;
      RECT 10.97 2.5 10.98 2.863 ;
      RECT 10.97 3.585 10.975 3.817 ;
      RECT 10.965 2.5 10.97 2.823 ;
      RECT 10.965 3.592 10.97 3.818 ;
      RECT 10.96 2.5 10.965 2.795 ;
      RECT 10.955 3.61 10.965 3.819 ;
      RECT 10.95 2.5 10.96 2.775 ;
      RECT 10.945 3.63 10.955 3.821 ;
      RECT 10.935 3.647 10.945 3.822 ;
      RECT 10.9 3.67 10.935 3.825 ;
      RECT 10.845 3.688 10.9 3.831 ;
      RECT 10.759 3.696 10.845 3.84 ;
      RECT 10.673 3.707 10.759 3.851 ;
      RECT 10.587 3.717 10.673 3.862 ;
      RECT 10.501 3.727 10.587 3.874 ;
      RECT 10.415 3.737 10.501 3.885 ;
      RECT 10.395 3.743 10.415 3.891 ;
      RECT 10.315 3.745 10.395 3.895 ;
      RECT 10.31 3.744 10.315 3.9 ;
      RECT 10.302 3.743 10.31 3.9 ;
      RECT 10.216 3.739 10.302 3.898 ;
      RECT 10.13 3.731 10.216 3.895 ;
      RECT 10.044 3.722 10.13 3.891 ;
      RECT 9.958 3.714 10.044 3.888 ;
      RECT 9.872 3.706 9.958 3.884 ;
      RECT 9.786 3.697 9.872 3.881 ;
      RECT 9.7 3.689 9.786 3.877 ;
      RECT 9.645 3.682 9.69 3.875 ;
      RECT 9.56 3.675 9.645 3.873 ;
      RECT 9.486 3.667 9.56 3.869 ;
      RECT 9.4 3.659 9.486 3.866 ;
      RECT 9.397 3.655 9.4 3.864 ;
      RECT 9.311 3.651 9.397 3.863 ;
      RECT 9.225 3.643 9.311 3.86 ;
      RECT 9.14 3.638 9.225 3.857 ;
      RECT 9.054 3.635 9.14 3.854 ;
      RECT 8.968 3.633 9.054 3.851 ;
      RECT 8.882 3.63 8.968 3.848 ;
      RECT 8.796 3.627 8.882 3.845 ;
      RECT 8.71 3.624 8.796 3.842 ;
      RECT 8.634 3.622 8.71 3.839 ;
      RECT 8.548 3.619 8.634 3.836 ;
      RECT 8.462 3.616 8.548 3.834 ;
      RECT 8.376 3.614 8.462 3.831 ;
      RECT 8.29 3.611 8.376 3.828 ;
      RECT 8.23 3.602 8.29 3.826 ;
      RECT 10.74 3.22 10.815 3.48 ;
      RECT 10.72 3.2 10.725 3.48 ;
      RECT 10.04 2.985 10.145 3.28 ;
      RECT 4.485 2.96 4.555 3.22 ;
      RECT 10.38 2.835 10.385 3.206 ;
      RECT 10.37 2.89 10.375 3.206 ;
      RECT 10.675 2.06 10.735 2.32 ;
      RECT 10.73 3.215 10.74 3.48 ;
      RECT 10.725 3.205 10.73 3.48 ;
      RECT 10.645 3.152 10.72 3.48 ;
      RECT 10.67 2.06 10.675 2.34 ;
      RECT 10.66 2.06 10.67 2.36 ;
      RECT 10.645 2.06 10.66 2.39 ;
      RECT 10.63 2.06 10.645 2.433 ;
      RECT 10.625 3.095 10.645 3.48 ;
      RECT 10.615 2.06 10.63 2.47 ;
      RECT 10.61 3.075 10.625 3.48 ;
      RECT 10.61 2.06 10.615 2.493 ;
      RECT 10.6 2.06 10.61 2.518 ;
      RECT 10.57 3.042 10.61 3.48 ;
      RECT 10.575 2.06 10.6 2.568 ;
      RECT 10.57 2.06 10.575 2.623 ;
      RECT 10.565 2.06 10.57 2.665 ;
      RECT 10.555 3.005 10.57 3.48 ;
      RECT 10.56 2.06 10.565 2.708 ;
      RECT 10.555 2.06 10.56 2.773 ;
      RECT 10.55 2.06 10.555 2.795 ;
      RECT 10.55 2.993 10.555 3.345 ;
      RECT 10.545 2.06 10.55 2.863 ;
      RECT 10.545 2.985 10.55 3.328 ;
      RECT 10.54 2.06 10.545 2.908 ;
      RECT 10.535 2.967 10.545 3.305 ;
      RECT 10.535 2.06 10.54 2.945 ;
      RECT 10.525 2.06 10.535 3.285 ;
      RECT 10.52 2.06 10.525 3.268 ;
      RECT 10.515 2.06 10.52 3.253 ;
      RECT 10.51 2.06 10.515 3.238 ;
      RECT 10.49 2.06 10.51 3.228 ;
      RECT 10.485 2.06 10.49 3.218 ;
      RECT 10.475 2.06 10.485 3.214 ;
      RECT 10.47 2.337 10.475 3.213 ;
      RECT 10.465 2.36 10.47 3.212 ;
      RECT 10.46 2.39 10.465 3.211 ;
      RECT 10.455 2.417 10.46 3.21 ;
      RECT 10.45 2.445 10.455 3.21 ;
      RECT 10.445 2.472 10.45 3.21 ;
      RECT 10.44 2.492 10.445 3.21 ;
      RECT 10.435 2.52 10.44 3.21 ;
      RECT 10.425 2.562 10.435 3.21 ;
      RECT 10.415 2.607 10.425 3.209 ;
      RECT 10.41 2.66 10.415 3.208 ;
      RECT 10.405 2.692 10.41 3.207 ;
      RECT 10.4 2.712 10.405 3.206 ;
      RECT 10.395 2.75 10.4 3.206 ;
      RECT 10.39 2.772 10.395 3.206 ;
      RECT 10.385 2.797 10.39 3.206 ;
      RECT 10.375 2.862 10.38 3.206 ;
      RECT 10.36 2.922 10.37 3.206 ;
      RECT 10.345 2.932 10.36 3.206 ;
      RECT 10.325 2.942 10.345 3.206 ;
      RECT 10.295 2.947 10.325 3.203 ;
      RECT 10.235 2.957 10.295 3.2 ;
      RECT 10.215 2.966 10.235 3.205 ;
      RECT 10.19 2.972 10.215 3.218 ;
      RECT 10.17 2.977 10.19 3.233 ;
      RECT 10.145 2.982 10.17 3.28 ;
      RECT 10.016 2.984 10.04 3.28 ;
      RECT 9.93 2.979 10.016 3.28 ;
      RECT 9.89 2.976 9.93 3.28 ;
      RECT 9.84 2.978 9.89 3.26 ;
      RECT 9.81 2.982 9.84 3.26 ;
      RECT 9.731 2.992 9.81 3.26 ;
      RECT 9.645 3.007 9.731 3.261 ;
      RECT 9.595 3.017 9.645 3.262 ;
      RECT 9.587 3.02 9.595 3.262 ;
      RECT 9.501 3.022 9.587 3.263 ;
      RECT 9.415 3.026 9.501 3.263 ;
      RECT 9.329 3.03 9.415 3.264 ;
      RECT 9.243 3.033 9.329 3.265 ;
      RECT 9.157 3.037 9.243 3.265 ;
      RECT 9.071 3.041 9.157 3.266 ;
      RECT 8.985 3.044 9.071 3.267 ;
      RECT 8.899 3.048 8.985 3.267 ;
      RECT 8.813 3.052 8.899 3.268 ;
      RECT 8.727 3.056 8.813 3.269 ;
      RECT 8.641 3.059 8.727 3.269 ;
      RECT 8.555 3.063 8.641 3.27 ;
      RECT 8.525 3.065 8.555 3.27 ;
      RECT 8.439 3.068 8.525 3.271 ;
      RECT 8.353 3.072 8.439 3.272 ;
      RECT 8.267 3.076 8.353 3.273 ;
      RECT 8.181 3.079 8.267 3.273 ;
      RECT 8.095 3.083 8.181 3.274 ;
      RECT 8.06 3.088 8.095 3.275 ;
      RECT 8.005 3.098 8.06 3.282 ;
      RECT 7.98 3.11 8.005 3.292 ;
      RECT 7.945 3.123 7.98 3.3 ;
      RECT 7.905 3.14 7.945 3.323 ;
      RECT 7.885 3.153 7.905 3.35 ;
      RECT 7.855 3.165 7.885 3.378 ;
      RECT 7.85 3.173 7.855 3.398 ;
      RECT 7.845 3.176 7.85 3.408 ;
      RECT 7.795 3.188 7.845 3.442 ;
      RECT 7.785 3.203 7.795 3.475 ;
      RECT 7.775 3.209 7.785 3.488 ;
      RECT 7.765 3.216 7.775 3.5 ;
      RECT 7.74 3.229 7.765 3.518 ;
      RECT 7.725 3.244 7.74 3.54 ;
      RECT 7.715 3.252 7.725 3.556 ;
      RECT 7.7 3.261 7.715 3.571 ;
      RECT 7.69 3.271 7.7 3.585 ;
      RECT 7.671 3.284 7.69 3.602 ;
      RECT 7.585 3.329 7.671 3.667 ;
      RECT 7.57 3.374 7.585 3.725 ;
      RECT 7.565 3.383 7.57 3.738 ;
      RECT 7.555 3.39 7.565 3.743 ;
      RECT 7.55 3.395 7.555 3.747 ;
      RECT 7.53 3.405 7.55 3.754 ;
      RECT 7.505 3.425 7.53 3.768 ;
      RECT 7.47 3.45 7.505 3.788 ;
      RECT 7.455 3.473 7.47 3.803 ;
      RECT 7.445 3.483 7.455 3.808 ;
      RECT 7.435 3.491 7.445 3.815 ;
      RECT 7.425 3.5 7.435 3.821 ;
      RECT 7.405 3.512 7.425 3.823 ;
      RECT 7.395 3.525 7.405 3.825 ;
      RECT 7.37 3.54 7.395 3.828 ;
      RECT 7.35 3.557 7.37 3.832 ;
      RECT 7.31 3.585 7.35 3.838 ;
      RECT 7.245 3.632 7.31 3.847 ;
      RECT 7.23 3.665 7.245 3.855 ;
      RECT 7.225 3.672 7.23 3.857 ;
      RECT 7.175 3.697 7.225 3.862 ;
      RECT 7.16 3.721 7.175 3.869 ;
      RECT 7.11 3.726 7.16 3.87 ;
      RECT 7.024 3.73 7.11 3.87 ;
      RECT 6.938 3.73 7.024 3.87 ;
      RECT 6.852 3.73 6.938 3.871 ;
      RECT 6.766 3.73 6.852 3.871 ;
      RECT 6.68 3.73 6.766 3.871 ;
      RECT 6.614 3.73 6.68 3.871 ;
      RECT 6.528 3.73 6.614 3.872 ;
      RECT 6.442 3.73 6.528 3.872 ;
      RECT 6.356 3.731 6.442 3.873 ;
      RECT 6.27 3.731 6.356 3.873 ;
      RECT 6.184 3.731 6.27 3.873 ;
      RECT 6.098 3.731 6.184 3.874 ;
      RECT 6.012 3.731 6.098 3.874 ;
      RECT 5.926 3.732 6.012 3.875 ;
      RECT 5.84 3.732 5.926 3.875 ;
      RECT 5.82 3.732 5.84 3.875 ;
      RECT 5.734 3.732 5.82 3.875 ;
      RECT 5.648 3.732 5.734 3.875 ;
      RECT 5.562 3.733 5.648 3.875 ;
      RECT 5.476 3.733 5.562 3.875 ;
      RECT 5.39 3.733 5.476 3.875 ;
      RECT 5.304 3.734 5.39 3.875 ;
      RECT 5.218 3.734 5.304 3.875 ;
      RECT 5.132 3.734 5.218 3.875 ;
      RECT 5.046 3.734 5.132 3.875 ;
      RECT 4.96 3.735 5.046 3.875 ;
      RECT 4.91 3.732 4.96 3.875 ;
      RECT 4.9 3.73 4.91 3.874 ;
      RECT 4.896 3.73 4.9 3.873 ;
      RECT 4.81 3.725 4.896 3.868 ;
      RECT 4.788 3.718 4.81 3.862 ;
      RECT 4.702 3.709 4.788 3.856 ;
      RECT 4.616 3.696 4.702 3.847 ;
      RECT 4.53 3.682 4.616 3.837 ;
      RECT 4.485 3.672 4.53 3.83 ;
      RECT 4.465 2.96 4.485 3.238 ;
      RECT 4.465 3.665 4.485 3.826 ;
      RECT 4.435 2.96 4.465 3.26 ;
      RECT 4.425 3.632 4.465 3.823 ;
      RECT 4.42 2.96 4.435 3.28 ;
      RECT 4.42 3.597 4.425 3.821 ;
      RECT 4.415 2.96 4.42 3.405 ;
      RECT 4.415 3.557 4.42 3.821 ;
      RECT 4.405 2.96 4.415 3.821 ;
      RECT 4.33 2.96 4.405 3.815 ;
      RECT 4.3 2.96 4.33 3.805 ;
      RECT 4.295 2.96 4.3 3.797 ;
      RECT 4.29 3.002 4.295 3.79 ;
      RECT 4.28 3.071 4.29 3.781 ;
      RECT 4.275 3.141 4.28 3.733 ;
      RECT 4.27 3.205 4.275 3.63 ;
      RECT 4.265 3.24 4.27 3.585 ;
      RECT 4.263 3.277 4.265 3.477 ;
      RECT 4.26 3.285 4.263 3.47 ;
      RECT 4.255 3.35 4.26 3.413 ;
      RECT 8.33 2.44 8.61 2.72 ;
      RECT 8.32 2.44 8.61 2.583 ;
      RECT 8.275 2.305 8.535 2.565 ;
      RECT 8.275 2.42 8.59 2.565 ;
      RECT 8.275 2.39 8.585 2.565 ;
      RECT 8.275 2.377 8.575 2.565 ;
      RECT 8.275 2.367 8.57 2.565 ;
      RECT 4.25 2.35 4.51 2.61 ;
      RECT 8.02 1.9 8.28 2.16 ;
      RECT 8.01 1.925 8.28 2.12 ;
      RECT 8.005 1.925 8.01 2.119 ;
      RECT 7.935 1.92 8.005 2.111 ;
      RECT 7.85 1.907 7.935 2.094 ;
      RECT 7.846 1.899 7.85 2.084 ;
      RECT 7.76 1.892 7.846 2.074 ;
      RECT 7.751 1.884 7.76 2.064 ;
      RECT 7.665 1.877 7.751 2.052 ;
      RECT 7.645 1.868 7.665 2.038 ;
      RECT 7.59 1.863 7.645 2.03 ;
      RECT 7.58 1.857 7.59 2.024 ;
      RECT 7.56 1.855 7.58 2.02 ;
      RECT 7.552 1.854 7.56 2.016 ;
      RECT 7.466 1.846 7.552 2.005 ;
      RECT 7.38 1.832 7.466 1.985 ;
      RECT 7.32 1.82 7.38 1.97 ;
      RECT 7.31 1.815 7.32 1.965 ;
      RECT 7.26 1.815 7.31 1.967 ;
      RECT 7.213 1.817 7.26 1.971 ;
      RECT 7.127 1.824 7.213 1.976 ;
      RECT 7.041 1.832 7.127 1.982 ;
      RECT 6.955 1.841 7.041 1.988 ;
      RECT 6.896 1.847 6.955 1.993 ;
      RECT 6.81 1.852 6.896 1.999 ;
      RECT 6.735 1.857 6.81 2.005 ;
      RECT 6.696 1.859 6.735 2.01 ;
      RECT 6.61 1.856 6.696 2.015 ;
      RECT 6.525 1.854 6.61 2.022 ;
      RECT 6.493 1.853 6.525 2.025 ;
      RECT 6.407 1.852 6.493 2.026 ;
      RECT 6.321 1.851 6.407 2.027 ;
      RECT 6.235 1.85 6.321 2.027 ;
      RECT 6.149 1.849 6.235 2.028 ;
      RECT 6.063 1.848 6.149 2.029 ;
      RECT 5.977 1.847 6.063 2.03 ;
      RECT 5.891 1.846 5.977 2.03 ;
      RECT 5.805 1.845 5.891 2.031 ;
      RECT 5.755 1.845 5.805 2.032 ;
      RECT 5.741 1.846 5.755 2.032 ;
      RECT 5.655 1.853 5.741 2.033 ;
      RECT 5.581 1.864 5.655 2.034 ;
      RECT 5.495 1.873 5.581 2.035 ;
      RECT 5.46 1.88 5.495 2.05 ;
      RECT 5.435 1.883 5.46 2.08 ;
      RECT 5.41 1.892 5.435 2.109 ;
      RECT 5.4 1.903 5.41 2.129 ;
      RECT 5.39 1.911 5.4 2.143 ;
      RECT 5.385 1.917 5.39 2.153 ;
      RECT 5.36 1.934 5.385 2.17 ;
      RECT 5.345 1.956 5.36 2.198 ;
      RECT 5.315 1.982 5.345 2.228 ;
      RECT 5.295 2.011 5.315 2.258 ;
      RECT 5.29 2.026 5.295 2.275 ;
      RECT 5.27 2.041 5.29 2.29 ;
      RECT 5.26 2.059 5.27 2.308 ;
      RECT 5.25 2.07 5.26 2.323 ;
      RECT 5.2 2.102 5.25 2.349 ;
      RECT 5.195 2.132 5.2 2.369 ;
      RECT 5.185 2.145 5.195 2.375 ;
      RECT 5.176 2.155 5.185 2.383 ;
      RECT 5.165 2.166 5.176 2.391 ;
      RECT 5.16 2.176 5.165 2.397 ;
      RECT 5.145 2.197 5.16 2.404 ;
      RECT 5.13 2.227 5.145 2.412 ;
      RECT 5.095 2.257 5.13 2.418 ;
      RECT 5.07 2.275 5.095 2.425 ;
      RECT 5.02 2.283 5.07 2.434 ;
      RECT 4.995 2.288 5.02 2.443 ;
      RECT 4.94 2.294 4.995 2.453 ;
      RECT 4.935 2.299 4.94 2.461 ;
      RECT 4.921 2.302 4.935 2.463 ;
      RECT 4.835 2.314 4.921 2.475 ;
      RECT 4.825 2.326 4.835 2.488 ;
      RECT 4.74 2.339 4.825 2.5 ;
      RECT 4.696 2.356 4.74 2.514 ;
      RECT 4.61 2.373 4.696 2.53 ;
      RECT 4.58 2.387 4.61 2.544 ;
      RECT 4.57 2.392 4.58 2.549 ;
      RECT 4.51 2.395 4.57 2.558 ;
      RECT 7.4 2.665 7.66 2.925 ;
      RECT 7.4 2.665 7.68 2.778 ;
      RECT 7.4 2.665 7.705 2.745 ;
      RECT 7.4 2.665 7.71 2.725 ;
      RECT 7.45 2.44 7.73 2.72 ;
      RECT 7.005 3.175 7.265 3.435 ;
      RECT 6.995 3.032 7.19 3.373 ;
      RECT 6.99 3.14 7.205 3.365 ;
      RECT 6.985 3.19 7.265 3.355 ;
      RECT 6.975 3.267 7.265 3.34 ;
      RECT 6.995 3.115 7.205 3.373 ;
      RECT 7.005 2.99 7.19 3.435 ;
      RECT 7.005 2.885 7.17 3.435 ;
      RECT 7.015 2.872 7.17 3.435 ;
      RECT 7.015 2.83 7.16 3.435 ;
      RECT 7.02 2.755 7.16 3.435 ;
      RECT 7.05 2.405 7.16 3.435 ;
      RECT 7.055 2.135 7.18 2.758 ;
      RECT 7.025 2.71 7.18 2.758 ;
      RECT 7.04 2.512 7.16 3.435 ;
      RECT 7.03 2.622 7.18 2.758 ;
      RECT 7.055 2.135 7.195 2.615 ;
      RECT 7.055 2.135 7.215 2.49 ;
      RECT 7.02 2.135 7.28 2.395 ;
      RECT 6.49 2.44 6.77 2.72 ;
      RECT 6.475 2.44 6.77 2.7 ;
      RECT 4.53 3.305 4.79 3.565 ;
      RECT 6.315 3.16 6.575 3.42 ;
      RECT 6.295 3.18 6.575 3.395 ;
      RECT 6.252 3.18 6.295 3.394 ;
      RECT 6.166 3.181 6.252 3.391 ;
      RECT 6.08 3.182 6.166 3.387 ;
      RECT 6.005 3.184 6.08 3.384 ;
      RECT 5.982 3.185 6.005 3.382 ;
      RECT 5.896 3.186 5.982 3.38 ;
      RECT 5.81 3.187 5.896 3.377 ;
      RECT 5.786 3.188 5.81 3.375 ;
      RECT 5.7 3.19 5.786 3.372 ;
      RECT 5.615 3.192 5.7 3.373 ;
      RECT 5.558 3.193 5.615 3.379 ;
      RECT 5.472 3.195 5.558 3.389 ;
      RECT 5.386 3.198 5.472 3.402 ;
      RECT 5.3 3.2 5.386 3.414 ;
      RECT 5.286 3.201 5.3 3.421 ;
      RECT 5.2 3.202 5.286 3.429 ;
      RECT 5.16 3.204 5.2 3.438 ;
      RECT 5.151 3.205 5.16 3.441 ;
      RECT 5.065 3.213 5.151 3.447 ;
      RECT 5.045 3.222 5.065 3.455 ;
      RECT 4.96 3.237 5.045 3.463 ;
      RECT 4.9 3.26 4.96 3.474 ;
      RECT 4.89 3.272 4.9 3.479 ;
      RECT 4.85 3.282 4.89 3.483 ;
      RECT 4.795 3.299 4.85 3.491 ;
      RECT 4.79 3.309 4.795 3.495 ;
      RECT 5.856 2.44 5.915 2.837 ;
      RECT 5.77 2.44 5.975 2.828 ;
      RECT 5.765 2.47 5.975 2.823 ;
      RECT 5.731 2.47 5.975 2.821 ;
      RECT 5.645 2.47 5.975 2.815 ;
      RECT 5.6 2.47 5.995 2.793 ;
      RECT 5.6 2.47 6.015 2.748 ;
      RECT 5.56 2.47 6.015 2.738 ;
      RECT 5.77 2.44 6.05 2.72 ;
      RECT 5.505 2.44 5.765 2.7 ;
      RECT 3.33 3 3.61 3.28 ;
      RECT 3.3 2.962 3.555 3.265 ;
      RECT 3.295 2.963 3.555 3.263 ;
      RECT 3.29 2.964 3.555 3.257 ;
      RECT 3.285 2.967 3.555 3.25 ;
      RECT 3.28 3 3.61 3.243 ;
      RECT 3.25 2.97 3.555 3.23 ;
      RECT 3.25 2.997 3.575 3.23 ;
      RECT 3.25 2.987 3.57 3.23 ;
      RECT 3.25 2.972 3.565 3.23 ;
      RECT 3.33 2.959 3.545 3.28 ;
      RECT 3.416 2.957 3.545 3.28 ;
      RECT 3.502 2.955 3.53 3.28 ;
      RECT 75.28 0.815 75.65 1.185 ;
      RECT 73.57 7.04 73.94 7.41 ;
      RECT 59.495 0.815 59.865 1.185 ;
      RECT 57.785 7.04 58.155 7.41 ;
      RECT 43.71 0.815 44.08 1.185 ;
      RECT 42 7.04 42.37 7.41 ;
      RECT 27.935 0.815 28.305 1.185 ;
      RECT 26.225 7.04 26.595 7.41 ;
      RECT 12.155 0.815 12.525 1.185 ;
      RECT 10.445 7.04 10.815 7.41 ;
      RECT 0.835 4.26 1.215 4.64 ;
      RECT 0.78 0 1.16 0.38 ;
      RECT 0.25 8.5 0.63 8.88 ;
    LAYER via1 ;
      RECT 81.305 7.375 81.455 7.525 ;
      RECT 78.935 6.74 79.085 6.89 ;
      RECT 78.92 2.065 79.07 2.215 ;
      RECT 78.13 2.45 78.28 2.6 ;
      RECT 78.13 6.325 78.28 6.475 ;
      RECT 76.485 1.44 76.635 1.59 ;
      RECT 76.17 2.96 76.32 3.11 ;
      RECT 75.39 0.925 75.54 1.075 ;
      RECT 75.27 2.29 75.42 2.44 ;
      RECT 75.15 2.86 75.3 3.01 ;
      RECT 74.32 6.71 74.47 6.86 ;
      RECT 74.07 2.555 74.22 2.705 ;
      RECT 73.735 3.275 73.885 3.425 ;
      RECT 73.68 7.15 73.83 7.3 ;
      RECT 73.655 2.115 73.805 2.265 ;
      RECT 72.22 2.51 72.37 2.66 ;
      RECT 71.455 2.36 71.605 2.51 ;
      RECT 71.2 1.955 71.35 2.105 ;
      RECT 70.58 2.72 70.73 2.87 ;
      RECT 70.2 2.19 70.35 2.34 ;
      RECT 70.185 3.23 70.335 3.38 ;
      RECT 69.655 2.495 69.805 2.645 ;
      RECT 69.495 3.215 69.645 3.365 ;
      RECT 68.685 2.495 68.835 2.645 ;
      RECT 67.87 1.975 68.02 2.125 ;
      RECT 67.71 3.36 67.86 3.51 ;
      RECT 67.475 3.015 67.625 3.165 ;
      RECT 67.43 2.405 67.58 2.555 ;
      RECT 66.43 3.025 66.58 3.175 ;
      RECT 65.495 6.755 65.645 6.905 ;
      RECT 63.15 6.74 63.3 6.89 ;
      RECT 63.135 2.065 63.285 2.215 ;
      RECT 62.345 2.45 62.495 2.6 ;
      RECT 62.345 6.325 62.495 6.475 ;
      RECT 60.7 1.44 60.85 1.59 ;
      RECT 60.385 2.96 60.535 3.11 ;
      RECT 59.605 0.925 59.755 1.075 ;
      RECT 59.485 2.29 59.635 2.44 ;
      RECT 59.365 2.86 59.515 3.01 ;
      RECT 58.535 6.71 58.685 6.86 ;
      RECT 58.285 2.555 58.435 2.705 ;
      RECT 57.95 3.275 58.1 3.425 ;
      RECT 57.895 7.15 58.045 7.3 ;
      RECT 57.87 2.115 58.02 2.265 ;
      RECT 56.435 2.51 56.585 2.66 ;
      RECT 55.67 2.36 55.82 2.51 ;
      RECT 55.415 1.955 55.565 2.105 ;
      RECT 54.795 2.72 54.945 2.87 ;
      RECT 54.415 2.19 54.565 2.34 ;
      RECT 54.4 3.23 54.55 3.38 ;
      RECT 53.87 2.495 54.02 2.645 ;
      RECT 53.71 3.215 53.86 3.365 ;
      RECT 52.9 2.495 53.05 2.645 ;
      RECT 52.085 1.975 52.235 2.125 ;
      RECT 51.925 3.36 52.075 3.51 ;
      RECT 51.69 3.015 51.84 3.165 ;
      RECT 51.645 2.405 51.795 2.555 ;
      RECT 50.645 3.025 50.795 3.175 ;
      RECT 49.71 6.755 49.86 6.905 ;
      RECT 47.365 6.74 47.515 6.89 ;
      RECT 47.35 2.065 47.5 2.215 ;
      RECT 46.56 2.45 46.71 2.6 ;
      RECT 46.56 6.325 46.71 6.475 ;
      RECT 44.915 1.44 45.065 1.59 ;
      RECT 44.6 2.96 44.75 3.11 ;
      RECT 43.82 0.925 43.97 1.075 ;
      RECT 43.7 2.29 43.85 2.44 ;
      RECT 43.58 2.86 43.73 3.01 ;
      RECT 42.805 6.715 42.955 6.865 ;
      RECT 42.5 2.555 42.65 2.705 ;
      RECT 42.165 3.275 42.315 3.425 ;
      RECT 42.11 7.15 42.26 7.3 ;
      RECT 42.085 2.115 42.235 2.265 ;
      RECT 40.65 2.51 40.8 2.66 ;
      RECT 39.885 2.36 40.035 2.51 ;
      RECT 39.63 1.955 39.78 2.105 ;
      RECT 39.01 2.72 39.16 2.87 ;
      RECT 38.63 2.19 38.78 2.34 ;
      RECT 38.615 3.23 38.765 3.38 ;
      RECT 38.085 2.495 38.235 2.645 ;
      RECT 37.925 3.215 38.075 3.365 ;
      RECT 37.115 2.495 37.265 2.645 ;
      RECT 36.3 1.975 36.45 2.125 ;
      RECT 36.14 3.36 36.29 3.51 ;
      RECT 35.905 3.015 36.055 3.165 ;
      RECT 35.86 2.405 36.01 2.555 ;
      RECT 34.86 3.025 35.01 3.175 ;
      RECT 33.98 6.76 34.13 6.91 ;
      RECT 31.59 6.74 31.74 6.89 ;
      RECT 31.575 2.065 31.725 2.215 ;
      RECT 30.785 2.45 30.935 2.6 ;
      RECT 30.785 6.325 30.935 6.475 ;
      RECT 29.14 1.44 29.29 1.59 ;
      RECT 28.825 2.96 28.975 3.11 ;
      RECT 28.045 0.925 28.195 1.075 ;
      RECT 27.925 2.29 28.075 2.44 ;
      RECT 27.805 2.86 27.955 3.01 ;
      RECT 27.025 6.71 27.175 6.86 ;
      RECT 26.725 2.555 26.875 2.705 ;
      RECT 26.39 3.275 26.54 3.425 ;
      RECT 26.335 7.15 26.485 7.3 ;
      RECT 26.31 2.115 26.46 2.265 ;
      RECT 24.875 2.51 25.025 2.66 ;
      RECT 24.11 2.36 24.26 2.51 ;
      RECT 23.855 1.955 24.005 2.105 ;
      RECT 23.235 2.72 23.385 2.87 ;
      RECT 22.855 2.19 23.005 2.34 ;
      RECT 22.84 3.23 22.99 3.38 ;
      RECT 22.31 2.495 22.46 2.645 ;
      RECT 22.15 3.215 22.3 3.365 ;
      RECT 21.34 2.495 21.49 2.645 ;
      RECT 20.525 1.975 20.675 2.125 ;
      RECT 20.365 3.36 20.515 3.51 ;
      RECT 20.13 3.015 20.28 3.165 ;
      RECT 20.085 2.405 20.235 2.555 ;
      RECT 19.085 3.025 19.235 3.175 ;
      RECT 18.2 6.755 18.35 6.905 ;
      RECT 15.81 6.74 15.96 6.89 ;
      RECT 15.795 2.065 15.945 2.215 ;
      RECT 15.005 2.45 15.155 2.6 ;
      RECT 15.005 6.325 15.155 6.475 ;
      RECT 13.36 1.44 13.51 1.59 ;
      RECT 13.045 2.96 13.195 3.11 ;
      RECT 12.265 0.925 12.415 1.075 ;
      RECT 12.145 2.29 12.295 2.44 ;
      RECT 12.025 2.86 12.175 3.01 ;
      RECT 11.215 6.705 11.365 6.855 ;
      RECT 10.945 2.555 11.095 2.705 ;
      RECT 10.61 3.275 10.76 3.425 ;
      RECT 10.555 7.15 10.705 7.3 ;
      RECT 10.53 2.115 10.68 2.265 ;
      RECT 9.095 2.51 9.245 2.66 ;
      RECT 8.33 2.36 8.48 2.51 ;
      RECT 8.075 1.955 8.225 2.105 ;
      RECT 7.455 2.72 7.605 2.87 ;
      RECT 7.075 2.19 7.225 2.34 ;
      RECT 7.06 3.23 7.21 3.38 ;
      RECT 6.53 2.495 6.68 2.645 ;
      RECT 6.37 3.215 6.52 3.365 ;
      RECT 5.56 2.495 5.71 2.645 ;
      RECT 4.745 1.975 4.895 2.125 ;
      RECT 4.585 3.36 4.735 3.51 ;
      RECT 4.35 3.015 4.5 3.165 ;
      RECT 4.305 2.405 4.455 2.555 ;
      RECT 3.305 3.025 3.455 3.175 ;
      RECT 1.62 7.095 1.77 7.245 ;
      RECT 1.245 6.355 1.395 6.505 ;
      RECT 0.95 4.365 1.1 4.515 ;
      RECT 0.895 0.115 1.045 0.265 ;
      RECT 0.365 8.615 0.515 8.765 ;
    LAYER met1 ;
      RECT -0.005 8.575 81.78 8.88 ;
      RECT 72.865 6.315 73.035 8.88 ;
      RECT 57.08 6.315 57.25 8.88 ;
      RECT 41.295 6.315 41.465 8.88 ;
      RECT 25.52 6.315 25.69 8.88 ;
      RECT 9.74 6.315 9.91 8.88 ;
      RECT 0.25 8.5 0.63 8.88 ;
      RECT 73.235 6.285 73.525 6.515 ;
      RECT 57.45 6.285 57.74 6.515 ;
      RECT 41.665 6.285 41.955 6.515 ;
      RECT 25.89 6.285 26.18 6.515 ;
      RECT 10.11 6.285 10.4 6.515 ;
      RECT 72.865 6.315 73.525 6.485 ;
      RECT 57.08 6.315 57.74 6.485 ;
      RECT 41.295 6.315 41.955 6.485 ;
      RECT 25.52 6.315 26.18 6.485 ;
      RECT 9.74 6.315 10.4 6.485 ;
      RECT 66.18 1.26 75.84 1.74 ;
      RECT 50.395 1.26 60.055 1.74 ;
      RECT 34.61 1.26 44.27 1.74 ;
      RECT 18.835 1.26 28.495 1.74 ;
      RECT 3.055 1.26 12.715 1.74 ;
      RECT 66.18 1.26 75.895 1.59 ;
      RECT 50.395 1.26 60.11 1.59 ;
      RECT 34.61 1.26 44.325 1.59 ;
      RECT 18.835 1.26 28.55 1.59 ;
      RECT 3.055 1.26 12.77 1.59 ;
      RECT 66.295 0 76.01 1.585 ;
      RECT 50.51 0 60.225 1.585 ;
      RECT 34.725 0 44.44 1.585 ;
      RECT 18.95 0 28.665 1.585 ;
      RECT 3.17 0 12.885 1.585 ;
      RECT 0.795 0 1.145 0.335 ;
      RECT 0.585 0 1.395 0.315 ;
      RECT 0 0 81.775 0.305 ;
      RECT 79.64 4.13 81.62 4.75 ;
      RECT 63.855 4.13 65.835 4.75 ;
      RECT 48.07 4.13 50.05 4.75 ;
      RECT 32.295 4.13 34.275 4.75 ;
      RECT 16.515 4.13 18.495 4.75 ;
      RECT 0 4.135 81.775 4.745 ;
      RECT 66.18 3.98 75.84 4.745 ;
      RECT 50.395 3.98 60.055 4.745 ;
      RECT 34.61 3.98 44.27 4.745 ;
      RECT 18.835 3.98 28.495 4.745 ;
      RECT 3.055 3.98 12.715 4.745 ;
      RECT 81.17 7.77 81.46 8 ;
      RECT 81.23 6.29 81.4 8 ;
      RECT 81.205 7.275 81.555 7.625 ;
      RECT 81.17 6.29 81.46 6.52 ;
      RECT 80.765 2.395 80.87 2.965 ;
      RECT 80.765 2.73 81.09 2.96 ;
      RECT 80.765 2.76 81.26 2.93 ;
      RECT 80.765 2.395 80.955 2.96 ;
      RECT 80.18 2.36 80.47 2.59 ;
      RECT 80.18 2.395 80.955 2.565 ;
      RECT 80.24 0.88 80.41 2.59 ;
      RECT 80.18 0.88 80.47 1.11 ;
      RECT 80.18 7.77 80.47 8 ;
      RECT 80.24 6.29 80.41 8 ;
      RECT 80.18 6.29 80.47 6.52 ;
      RECT 80.18 6.325 81.035 6.485 ;
      RECT 80.865 5.92 81.035 6.485 ;
      RECT 80.18 6.32 80.575 6.485 ;
      RECT 80.8 5.92 81.09 6.15 ;
      RECT 80.8 5.95 81.26 6.12 ;
      RECT 79.81 2.73 80.1 2.96 ;
      RECT 79.81 2.76 80.27 2.93 ;
      RECT 79.875 1.655 80.04 2.96 ;
      RECT 78.39 1.625 78.68 1.855 ;
      RECT 78.39 1.655 80.04 1.825 ;
      RECT 78.45 0.885 78.62 1.855 ;
      RECT 78.39 0.885 78.68 1.115 ;
      RECT 78.39 7.765 78.68 7.995 ;
      RECT 78.45 7.025 78.62 7.995 ;
      RECT 78.45 7.12 80.04 7.29 ;
      RECT 79.87 5.92 80.04 7.29 ;
      RECT 78.39 7.025 78.68 7.255 ;
      RECT 79.81 5.92 80.1 6.15 ;
      RECT 79.81 5.95 80.27 6.12 ;
      RECT 78.82 1.965 79.17 2.315 ;
      RECT 76.485 2.025 79.17 2.195 ;
      RECT 76.485 1.34 76.655 2.195 ;
      RECT 76.385 1.34 76.735 1.69 ;
      RECT 78.845 6.655 79.17 6.98 ;
      RECT 74.22 6.61 74.57 6.96 ;
      RECT 78.82 6.655 79.17 6.885 ;
      RECT 74.04 6.655 74.57 6.885 ;
      RECT 73.87 6.685 79.17 6.855 ;
      RECT 78.045 2.365 78.365 2.685 ;
      RECT 78.015 2.365 78.365 2.595 ;
      RECT 77.845 2.395 78.365 2.565 ;
      RECT 78.045 6.255 78.365 6.545 ;
      RECT 78.015 6.285 78.365 6.515 ;
      RECT 77.845 6.315 78.365 6.485 ;
      RECT 74.68 2.465 74.865 2.675 ;
      RECT 74.67 2.47 74.88 2.668 ;
      RECT 74.67 2.47 74.966 2.645 ;
      RECT 74.67 2.47 75.025 2.62 ;
      RECT 74.67 2.47 75.08 2.6 ;
      RECT 74.67 2.47 75.09 2.588 ;
      RECT 74.67 2.47 75.285 2.527 ;
      RECT 74.67 2.47 75.315 2.51 ;
      RECT 74.67 2.47 75.335 2.5 ;
      RECT 75.215 2.235 75.475 2.495 ;
      RECT 75.2 2.325 75.215 2.542 ;
      RECT 74.735 2.457 75.475 2.495 ;
      RECT 75.186 2.336 75.2 2.548 ;
      RECT 74.775 2.45 75.475 2.495 ;
      RECT 75.1 2.376 75.186 2.567 ;
      RECT 75.025 2.437 75.475 2.495 ;
      RECT 75.095 2.412 75.1 2.584 ;
      RECT 75.08 2.422 75.475 2.495 ;
      RECT 75.09 2.417 75.095 2.586 ;
      RECT 75.385 2.922 75.39 3.014 ;
      RECT 75.38 2.9 75.385 3.031 ;
      RECT 75.375 2.89 75.38 3.043 ;
      RECT 75.365 2.881 75.375 3.053 ;
      RECT 75.36 2.876 75.365 3.061 ;
      RECT 75.355 2.735 75.36 3.064 ;
      RECT 75.321 2.735 75.355 3.075 ;
      RECT 75.235 2.735 75.321 3.11 ;
      RECT 75.155 2.735 75.235 3.158 ;
      RECT 75.126 2.735 75.155 3.182 ;
      RECT 75.04 2.735 75.126 3.188 ;
      RECT 75.035 2.919 75.04 3.193 ;
      RECT 75 2.93 75.035 3.196 ;
      RECT 74.975 2.945 75 3.2 ;
      RECT 74.961 2.954 74.975 3.202 ;
      RECT 74.875 2.981 74.961 3.208 ;
      RECT 74.81 3.022 74.875 3.217 ;
      RECT 74.795 3.042 74.81 3.222 ;
      RECT 74.765 3.052 74.795 3.225 ;
      RECT 74.76 3.062 74.765 3.228 ;
      RECT 74.73 3.067 74.76 3.23 ;
      RECT 74.71 3.072 74.73 3.234 ;
      RECT 74.625 3.075 74.71 3.241 ;
      RECT 74.61 3.072 74.625 3.247 ;
      RECT 74.6 3.069 74.61 3.249 ;
      RECT 74.58 3.066 74.6 3.251 ;
      RECT 74.56 3.062 74.58 3.252 ;
      RECT 74.545 3.058 74.56 3.254 ;
      RECT 74.535 3.055 74.545 3.255 ;
      RECT 74.495 3.049 74.535 3.253 ;
      RECT 74.485 3.044 74.495 3.251 ;
      RECT 74.47 3.041 74.485 3.247 ;
      RECT 74.445 3.036 74.47 3.24 ;
      RECT 74.395 3.027 74.445 3.228 ;
      RECT 74.325 3.013 74.395 3.21 ;
      RECT 74.267 2.998 74.325 3.192 ;
      RECT 74.181 2.981 74.267 3.172 ;
      RECT 74.095 2.96 74.181 3.147 ;
      RECT 74.045 2.945 74.095 3.128 ;
      RECT 74.041 2.939 74.045 3.12 ;
      RECT 73.955 2.929 74.041 3.107 ;
      RECT 73.92 2.914 73.955 3.09 ;
      RECT 73.905 2.907 73.92 3.083 ;
      RECT 73.845 2.895 73.905 3.071 ;
      RECT 73.825 2.882 73.845 3.059 ;
      RECT 73.785 2.873 73.825 3.051 ;
      RECT 73.78 2.865 73.785 3.044 ;
      RECT 73.7 2.855 73.78 3.03 ;
      RECT 73.685 2.842 73.7 3.015 ;
      RECT 73.68 2.84 73.685 3.013 ;
      RECT 73.601 2.828 73.68 3 ;
      RECT 73.515 2.803 73.601 2.975 ;
      RECT 73.5 2.772 73.515 2.96 ;
      RECT 73.485 2.747 73.5 2.956 ;
      RECT 73.47 2.74 73.485 2.952 ;
      RECT 73.295 2.745 73.3 2.948 ;
      RECT 73.29 2.75 73.295 2.943 ;
      RECT 73.3 2.74 73.47 2.95 ;
      RECT 74.015 2.5 74.12 2.76 ;
      RECT 74.83 2.025 74.835 2.25 ;
      RECT 74.96 2.025 75.015 2.235 ;
      RECT 75.015 2.03 75.025 2.228 ;
      RECT 74.921 2.025 74.96 2.238 ;
      RECT 74.835 2.025 74.921 2.245 ;
      RECT 74.815 2.03 74.83 2.251 ;
      RECT 74.805 2.07 74.815 2.253 ;
      RECT 74.775 2.08 74.805 2.255 ;
      RECT 74.77 2.085 74.775 2.257 ;
      RECT 74.745 2.09 74.77 2.259 ;
      RECT 74.73 2.095 74.745 2.261 ;
      RECT 74.715 2.097 74.73 2.263 ;
      RECT 74.71 2.102 74.715 2.265 ;
      RECT 74.66 2.11 74.71 2.268 ;
      RECT 74.635 2.119 74.66 2.273 ;
      RECT 74.625 2.126 74.635 2.278 ;
      RECT 74.62 2.129 74.625 2.282 ;
      RECT 74.6 2.132 74.62 2.291 ;
      RECT 74.57 2.14 74.6 2.311 ;
      RECT 74.541 2.153 74.57 2.333 ;
      RECT 74.455 2.187 74.541 2.377 ;
      RECT 74.45 2.213 74.455 2.415 ;
      RECT 74.445 2.217 74.45 2.424 ;
      RECT 74.41 2.23 74.445 2.457 ;
      RECT 74.4 2.244 74.41 2.495 ;
      RECT 74.395 2.248 74.4 2.508 ;
      RECT 74.39 2.252 74.395 2.513 ;
      RECT 74.38 2.26 74.39 2.525 ;
      RECT 74.375 2.267 74.38 2.54 ;
      RECT 74.35 2.28 74.375 2.565 ;
      RECT 74.31 2.309 74.35 2.62 ;
      RECT 74.295 2.334 74.31 2.675 ;
      RECT 74.285 2.345 74.295 2.698 ;
      RECT 74.28 2.352 74.285 2.71 ;
      RECT 74.275 2.356 74.28 2.718 ;
      RECT 74.22 2.384 74.275 2.76 ;
      RECT 74.2 2.42 74.22 2.76 ;
      RECT 74.185 2.435 74.2 2.76 ;
      RECT 74.13 2.467 74.185 2.76 ;
      RECT 74.12 2.497 74.13 2.76 ;
      RECT 73.73 2.112 73.915 2.35 ;
      RECT 73.715 2.114 73.925 2.345 ;
      RECT 73.6 2.06 73.86 2.32 ;
      RECT 73.595 2.097 73.86 2.274 ;
      RECT 73.59 2.107 73.86 2.271 ;
      RECT 73.585 2.147 73.925 2.265 ;
      RECT 73.58 2.18 73.925 2.255 ;
      RECT 73.59 2.122 73.94 2.193 ;
      RECT 73.887 3.22 73.9 3.75 ;
      RECT 73.801 3.22 73.9 3.749 ;
      RECT 73.801 3.22 73.905 3.748 ;
      RECT 73.715 3.22 73.905 3.746 ;
      RECT 73.71 3.22 73.905 3.743 ;
      RECT 73.71 3.22 73.915 3.741 ;
      RECT 73.705 3.512 73.915 3.738 ;
      RECT 73.705 3.522 73.92 3.735 ;
      RECT 73.705 3.59 73.925 3.731 ;
      RECT 73.695 3.595 73.925 3.73 ;
      RECT 73.695 3.687 73.93 3.727 ;
      RECT 73.68 3.22 73.94 3.48 ;
      RECT 73.61 7.765 73.9 7.995 ;
      RECT 73.67 7.025 73.84 7.995 ;
      RECT 73.585 7.055 73.925 7.4 ;
      RECT 73.61 7.025 73.9 7.4 ;
      RECT 72.91 2.21 72.955 3.745 ;
      RECT 73.11 2.21 73.14 2.425 ;
      RECT 71.485 1.95 71.605 2.16 ;
      RECT 71.145 1.9 71.405 2.16 ;
      RECT 71.145 1.945 71.44 2.15 ;
      RECT 73.15 2.226 73.155 2.28 ;
      RECT 73.145 2.219 73.15 2.413 ;
      RECT 73.14 2.213 73.145 2.42 ;
      RECT 73.095 2.21 73.11 2.433 ;
      RECT 73.09 2.21 73.095 2.455 ;
      RECT 73.085 2.21 73.09 2.503 ;
      RECT 73.08 2.21 73.085 2.523 ;
      RECT 73.07 2.21 73.08 2.63 ;
      RECT 73.065 2.21 73.07 2.693 ;
      RECT 73.06 2.21 73.065 2.75 ;
      RECT 73.055 2.21 73.06 2.758 ;
      RECT 73.04 2.21 73.055 2.865 ;
      RECT 73.03 2.21 73.04 3 ;
      RECT 73.02 2.21 73.03 3.11 ;
      RECT 73.01 2.21 73.02 3.167 ;
      RECT 73.005 2.21 73.01 3.207 ;
      RECT 73 2.21 73.005 3.243 ;
      RECT 72.99 2.21 73 3.283 ;
      RECT 72.985 2.21 72.99 3.325 ;
      RECT 72.965 2.21 72.985 3.39 ;
      RECT 72.97 3.535 72.975 3.715 ;
      RECT 72.965 3.517 72.97 3.723 ;
      RECT 72.96 2.21 72.965 3.453 ;
      RECT 72.96 3.497 72.965 3.73 ;
      RECT 72.955 2.21 72.96 3.74 ;
      RECT 72.9 2.21 72.91 2.51 ;
      RECT 72.905 2.757 72.91 3.745 ;
      RECT 72.9 2.822 72.905 3.745 ;
      RECT 72.895 2.211 72.9 2.5 ;
      RECT 72.89 2.887 72.9 3.745 ;
      RECT 72.885 2.212 72.895 2.49 ;
      RECT 72.875 3 72.89 3.745 ;
      RECT 72.88 2.213 72.885 2.48 ;
      RECT 72.86 2.214 72.88 2.458 ;
      RECT 72.865 3.097 72.875 3.745 ;
      RECT 72.86 3.172 72.865 3.745 ;
      RECT 72.85 2.213 72.86 2.435 ;
      RECT 72.855 3.215 72.86 3.745 ;
      RECT 72.85 3.242 72.855 3.745 ;
      RECT 72.84 2.211 72.85 2.423 ;
      RECT 72.845 3.285 72.85 3.745 ;
      RECT 72.84 3.312 72.845 3.745 ;
      RECT 72.83 2.21 72.84 2.41 ;
      RECT 72.835 3.327 72.84 3.745 ;
      RECT 72.795 3.385 72.835 3.745 ;
      RECT 72.825 2.209 72.83 2.395 ;
      RECT 72.82 2.207 72.825 2.388 ;
      RECT 72.81 2.204 72.82 2.378 ;
      RECT 72.805 2.201 72.81 2.363 ;
      RECT 72.79 2.197 72.805 2.356 ;
      RECT 72.785 3.44 72.795 3.745 ;
      RECT 72.785 2.194 72.79 2.351 ;
      RECT 72.77 2.19 72.785 2.345 ;
      RECT 72.78 3.457 72.785 3.745 ;
      RECT 72.77 3.52 72.78 3.745 ;
      RECT 72.69 2.175 72.77 2.325 ;
      RECT 72.765 3.527 72.77 3.74 ;
      RECT 72.76 3.535 72.765 3.73 ;
      RECT 72.68 2.161 72.69 2.309 ;
      RECT 72.665 2.157 72.68 2.307 ;
      RECT 72.655 2.152 72.665 2.303 ;
      RECT 72.63 2.145 72.655 2.295 ;
      RECT 72.625 2.14 72.63 2.29 ;
      RECT 72.615 2.14 72.625 2.288 ;
      RECT 72.605 2.138 72.615 2.286 ;
      RECT 72.575 2.13 72.605 2.28 ;
      RECT 72.56 2.122 72.575 2.273 ;
      RECT 72.54 2.117 72.56 2.266 ;
      RECT 72.535 2.113 72.54 2.261 ;
      RECT 72.505 2.106 72.535 2.255 ;
      RECT 72.48 2.097 72.505 2.245 ;
      RECT 72.45 2.09 72.48 2.237 ;
      RECT 72.425 2.08 72.45 2.228 ;
      RECT 72.41 2.072 72.425 2.222 ;
      RECT 72.385 2.067 72.41 2.217 ;
      RECT 72.375 2.063 72.385 2.212 ;
      RECT 72.355 2.058 72.375 2.207 ;
      RECT 72.32 2.053 72.355 2.2 ;
      RECT 72.26 2.048 72.32 2.193 ;
      RECT 72.247 2.044 72.26 2.191 ;
      RECT 72.161 2.039 72.247 2.188 ;
      RECT 72.075 2.029 72.161 2.184 ;
      RECT 72.034 2.022 72.075 2.181 ;
      RECT 71.948 2.015 72.034 2.178 ;
      RECT 71.862 2.005 71.948 2.174 ;
      RECT 71.776 1.995 71.862 2.169 ;
      RECT 71.69 1.985 71.776 2.165 ;
      RECT 71.68 1.97 71.69 2.163 ;
      RECT 71.67 1.955 71.68 2.163 ;
      RECT 71.605 1.95 71.67 2.162 ;
      RECT 71.44 1.947 71.485 2.155 ;
      RECT 72.685 2.852 72.69 3.043 ;
      RECT 72.68 2.847 72.685 3.05 ;
      RECT 72.666 2.845 72.68 3.056 ;
      RECT 72.58 2.845 72.666 3.058 ;
      RECT 72.576 2.845 72.58 3.061 ;
      RECT 72.49 2.845 72.576 3.079 ;
      RECT 72.48 2.85 72.49 3.098 ;
      RECT 72.47 2.905 72.48 3.102 ;
      RECT 72.445 2.92 72.47 3.109 ;
      RECT 72.405 2.94 72.445 3.122 ;
      RECT 72.4 2.952 72.405 3.132 ;
      RECT 72.385 2.958 72.4 3.137 ;
      RECT 72.38 2.963 72.385 3.141 ;
      RECT 72.36 2.97 72.38 3.146 ;
      RECT 72.29 2.995 72.36 3.163 ;
      RECT 72.25 3.023 72.29 3.183 ;
      RECT 72.245 3.033 72.25 3.191 ;
      RECT 72.225 3.04 72.245 3.193 ;
      RECT 72.22 3.047 72.225 3.196 ;
      RECT 72.19 3.055 72.22 3.199 ;
      RECT 72.185 3.06 72.19 3.203 ;
      RECT 72.111 3.064 72.185 3.211 ;
      RECT 72.025 3.073 72.111 3.227 ;
      RECT 72.021 3.078 72.025 3.236 ;
      RECT 71.935 3.083 72.021 3.246 ;
      RECT 71.895 3.091 71.935 3.258 ;
      RECT 71.845 3.097 71.895 3.265 ;
      RECT 71.76 3.106 71.845 3.28 ;
      RECT 71.685 3.117 71.76 3.298 ;
      RECT 71.65 3.124 71.685 3.308 ;
      RECT 71.575 3.132 71.65 3.313 ;
      RECT 71.52 3.141 71.575 3.313 ;
      RECT 71.495 3.146 71.52 3.311 ;
      RECT 71.485 3.149 71.495 3.309 ;
      RECT 71.45 3.151 71.485 3.307 ;
      RECT 71.42 3.153 71.45 3.303 ;
      RECT 71.375 3.152 71.42 3.299 ;
      RECT 71.355 3.147 71.375 3.296 ;
      RECT 71.305 3.132 71.355 3.293 ;
      RECT 71.295 3.117 71.305 3.288 ;
      RECT 71.245 3.102 71.295 3.278 ;
      RECT 71.195 3.077 71.245 3.258 ;
      RECT 71.185 3.062 71.195 3.24 ;
      RECT 71.18 3.06 71.185 3.234 ;
      RECT 71.16 3.055 71.18 3.229 ;
      RECT 71.155 3.047 71.16 3.223 ;
      RECT 71.14 3.041 71.155 3.216 ;
      RECT 71.135 3.036 71.14 3.208 ;
      RECT 71.115 3.031 71.135 3.2 ;
      RECT 71.1 3.024 71.115 3.193 ;
      RECT 71.085 3.018 71.1 3.184 ;
      RECT 71.08 3.012 71.085 3.177 ;
      RECT 71.035 2.987 71.08 3.163 ;
      RECT 71.02 2.957 71.035 3.145 ;
      RECT 71.005 2.94 71.02 3.136 ;
      RECT 70.98 2.92 71.005 3.124 ;
      RECT 70.94 2.89 70.98 3.104 ;
      RECT 70.93 2.86 70.94 3.089 ;
      RECT 70.915 2.85 70.93 3.082 ;
      RECT 70.86 2.815 70.915 3.061 ;
      RECT 70.845 2.778 70.86 3.04 ;
      RECT 70.835 2.765 70.845 3.032 ;
      RECT 70.785 2.735 70.835 3.014 ;
      RECT 70.77 2.665 70.785 2.995 ;
      RECT 70.725 2.665 70.77 2.978 ;
      RECT 70.7 2.665 70.725 2.96 ;
      RECT 70.69 2.665 70.7 2.953 ;
      RECT 70.611 2.665 70.69 2.946 ;
      RECT 70.525 2.665 70.611 2.938 ;
      RECT 70.51 2.697 70.525 2.933 ;
      RECT 70.435 2.707 70.51 2.929 ;
      RECT 70.415 2.717 70.435 2.924 ;
      RECT 70.39 2.717 70.415 2.921 ;
      RECT 70.38 2.707 70.39 2.92 ;
      RECT 70.37 2.68 70.38 2.919 ;
      RECT 70.33 2.675 70.37 2.917 ;
      RECT 70.285 2.675 70.33 2.913 ;
      RECT 70.26 2.675 70.285 2.908 ;
      RECT 70.21 2.675 70.26 2.895 ;
      RECT 70.17 2.68 70.18 2.88 ;
      RECT 70.18 2.675 70.21 2.885 ;
      RECT 72.165 2.455 72.425 2.715 ;
      RECT 72.16 2.477 72.425 2.673 ;
      RECT 71.4 2.305 71.62 2.67 ;
      RECT 71.382 2.392 71.62 2.669 ;
      RECT 71.365 2.397 71.62 2.666 ;
      RECT 71.365 2.397 71.64 2.665 ;
      RECT 71.335 2.407 71.64 2.663 ;
      RECT 71.33 2.422 71.64 2.659 ;
      RECT 71.33 2.422 71.645 2.658 ;
      RECT 71.325 2.48 71.645 2.656 ;
      RECT 71.325 2.48 71.655 2.653 ;
      RECT 71.32 2.545 71.655 2.648 ;
      RECT 71.4 2.305 71.66 2.565 ;
      RECT 70.145 2.135 70.405 2.395 ;
      RECT 70.145 2.178 70.491 2.369 ;
      RECT 70.145 2.178 70.535 2.368 ;
      RECT 70.145 2.178 70.555 2.366 ;
      RECT 70.145 2.178 70.655 2.365 ;
      RECT 70.145 2.178 70.675 2.363 ;
      RECT 70.145 2.178 70.685 2.358 ;
      RECT 70.555 2.145 70.745 2.355 ;
      RECT 70.555 2.147 70.75 2.353 ;
      RECT 70.545 2.152 70.755 2.345 ;
      RECT 70.491 2.176 70.755 2.345 ;
      RECT 70.535 2.17 70.545 2.367 ;
      RECT 70.545 2.15 70.75 2.353 ;
      RECT 69.5 3.21 69.705 3.44 ;
      RECT 69.44 3.16 69.495 3.42 ;
      RECT 69.5 3.16 69.7 3.44 ;
      RECT 70.47 3.475 70.475 3.502 ;
      RECT 70.46 3.385 70.47 3.507 ;
      RECT 70.455 3.307 70.46 3.513 ;
      RECT 70.445 3.297 70.455 3.52 ;
      RECT 70.44 3.287 70.445 3.526 ;
      RECT 70.43 3.282 70.44 3.528 ;
      RECT 70.415 3.274 70.43 3.536 ;
      RECT 70.4 3.265 70.415 3.548 ;
      RECT 70.39 3.257 70.4 3.558 ;
      RECT 70.355 3.175 70.39 3.576 ;
      RECT 70.32 3.175 70.355 3.595 ;
      RECT 70.305 3.175 70.32 3.603 ;
      RECT 70.25 3.175 70.305 3.603 ;
      RECT 70.216 3.175 70.25 3.594 ;
      RECT 70.13 3.175 70.216 3.57 ;
      RECT 70.12 3.235 70.13 3.552 ;
      RECT 70.08 3.237 70.12 3.543 ;
      RECT 70.075 3.239 70.08 3.533 ;
      RECT 70.055 3.241 70.075 3.528 ;
      RECT 70.045 3.244 70.055 3.523 ;
      RECT 70.035 3.245 70.045 3.518 ;
      RECT 70.011 3.246 70.035 3.51 ;
      RECT 69.925 3.251 70.011 3.488 ;
      RECT 69.87 3.25 69.925 3.461 ;
      RECT 69.855 3.243 69.87 3.448 ;
      RECT 69.82 3.238 69.855 3.444 ;
      RECT 69.765 3.23 69.82 3.443 ;
      RECT 69.705 3.217 69.765 3.441 ;
      RECT 69.495 3.16 69.5 3.428 ;
      RECT 69.57 2.53 69.755 2.74 ;
      RECT 69.56 2.535 69.77 2.733 ;
      RECT 69.6 2.44 69.86 2.7 ;
      RECT 69.555 2.597 69.86 2.623 ;
      RECT 68.9 2.39 68.905 3.19 ;
      RECT 68.845 2.44 68.875 3.19 ;
      RECT 68.835 2.44 68.84 2.75 ;
      RECT 68.82 2.44 68.825 2.745 ;
      RECT 68.365 2.485 68.38 2.7 ;
      RECT 68.295 2.485 68.38 2.695 ;
      RECT 69.56 2.065 69.63 2.275 ;
      RECT 69.63 2.072 69.64 2.27 ;
      RECT 69.526 2.065 69.56 2.282 ;
      RECT 69.44 2.065 69.526 2.306 ;
      RECT 69.43 2.07 69.44 2.325 ;
      RECT 69.425 2.082 69.43 2.328 ;
      RECT 69.41 2.097 69.425 2.332 ;
      RECT 69.405 2.115 69.41 2.336 ;
      RECT 69.365 2.125 69.405 2.345 ;
      RECT 69.35 2.132 69.365 2.357 ;
      RECT 69.335 2.137 69.35 2.362 ;
      RECT 69.32 2.14 69.335 2.367 ;
      RECT 69.31 2.142 69.32 2.371 ;
      RECT 69.275 2.149 69.31 2.379 ;
      RECT 69.24 2.157 69.275 2.393 ;
      RECT 69.23 2.163 69.24 2.402 ;
      RECT 69.225 2.165 69.23 2.404 ;
      RECT 69.205 2.168 69.225 2.41 ;
      RECT 69.175 2.175 69.205 2.421 ;
      RECT 69.165 2.181 69.175 2.428 ;
      RECT 69.14 2.184 69.165 2.435 ;
      RECT 69.13 2.188 69.14 2.443 ;
      RECT 69.125 2.189 69.13 2.465 ;
      RECT 69.12 2.19 69.125 2.48 ;
      RECT 69.115 2.191 69.12 2.495 ;
      RECT 69.11 2.192 69.115 2.51 ;
      RECT 69.105 2.193 69.11 2.54 ;
      RECT 69.095 2.195 69.105 2.573 ;
      RECT 69.08 2.199 69.095 2.62 ;
      RECT 69.07 2.202 69.08 2.665 ;
      RECT 69.065 2.205 69.07 2.693 ;
      RECT 69.055 2.207 69.065 2.72 ;
      RECT 69.05 2.21 69.055 2.755 ;
      RECT 69.02 2.215 69.05 2.813 ;
      RECT 69.015 2.22 69.02 2.898 ;
      RECT 69.01 2.222 69.015 2.933 ;
      RECT 69.005 2.224 69.01 3.015 ;
      RECT 69 2.226 69.005 3.103 ;
      RECT 68.99 2.228 69 3.185 ;
      RECT 68.975 2.242 68.99 3.19 ;
      RECT 68.94 2.287 68.975 3.19 ;
      RECT 68.93 2.327 68.94 3.19 ;
      RECT 68.915 2.355 68.93 3.19 ;
      RECT 68.91 2.372 68.915 3.19 ;
      RECT 68.905 2.38 68.91 3.19 ;
      RECT 68.895 2.395 68.9 3.19 ;
      RECT 68.89 2.402 68.895 3.19 ;
      RECT 68.88 2.422 68.89 3.19 ;
      RECT 68.875 2.435 68.88 3.19 ;
      RECT 68.84 2.44 68.845 2.775 ;
      RECT 68.825 2.83 68.845 3.19 ;
      RECT 68.825 2.44 68.835 2.748 ;
      RECT 68.82 2.87 68.825 3.19 ;
      RECT 68.77 2.44 68.82 2.743 ;
      RECT 68.815 2.907 68.82 3.19 ;
      RECT 68.805 2.93 68.815 3.19 ;
      RECT 68.8 2.975 68.805 3.19 ;
      RECT 68.79 2.985 68.8 3.183 ;
      RECT 68.716 2.44 68.77 2.737 ;
      RECT 68.63 2.44 68.716 2.73 ;
      RECT 68.581 2.487 68.63 2.723 ;
      RECT 68.495 2.495 68.581 2.716 ;
      RECT 68.48 2.492 68.495 2.711 ;
      RECT 68.466 2.485 68.48 2.71 ;
      RECT 68.38 2.485 68.466 2.705 ;
      RECT 68.285 2.49 68.295 2.69 ;
      RECT 67.875 1.92 67.89 2.32 ;
      RECT 68.07 1.92 68.075 2.18 ;
      RECT 67.815 1.92 67.86 2.18 ;
      RECT 68.27 3.225 68.275 3.43 ;
      RECT 68.265 3.215 68.27 3.435 ;
      RECT 68.26 3.202 68.265 3.44 ;
      RECT 68.255 3.182 68.26 3.44 ;
      RECT 68.23 3.135 68.255 3.44 ;
      RECT 68.195 3.05 68.23 3.44 ;
      RECT 68.19 2.987 68.195 3.44 ;
      RECT 68.185 2.972 68.19 3.44 ;
      RECT 68.17 2.932 68.185 3.44 ;
      RECT 68.165 2.907 68.17 3.44 ;
      RECT 68.155 2.89 68.165 3.44 ;
      RECT 68.12 2.812 68.155 3.44 ;
      RECT 68.115 2.755 68.12 3.44 ;
      RECT 68.11 2.742 68.115 3.44 ;
      RECT 68.1 2.72 68.11 3.44 ;
      RECT 68.09 2.685 68.1 3.44 ;
      RECT 68.08 2.655 68.09 3.44 ;
      RECT 68.07 2.57 68.08 3.083 ;
      RECT 68.077 3.215 68.08 3.44 ;
      RECT 68.075 3.225 68.077 3.44 ;
      RECT 68.065 3.235 68.075 3.435 ;
      RECT 68.06 1.92 68.07 2.315 ;
      RECT 68.065 2.447 68.07 3.058 ;
      RECT 68.06 2.345 68.065 3.041 ;
      RECT 68.05 1.92 68.06 3.017 ;
      RECT 68.045 1.92 68.05 2.988 ;
      RECT 68.04 1.92 68.045 2.978 ;
      RECT 68.02 1.92 68.04 2.94 ;
      RECT 68.015 1.92 68.02 2.898 ;
      RECT 68.01 1.92 68.015 2.878 ;
      RECT 67.98 1.92 68.01 2.828 ;
      RECT 67.97 1.92 67.98 2.775 ;
      RECT 67.965 1.92 67.97 2.748 ;
      RECT 67.96 1.92 67.965 2.733 ;
      RECT 67.95 1.92 67.96 2.71 ;
      RECT 67.94 1.92 67.95 2.685 ;
      RECT 67.935 1.92 67.94 2.625 ;
      RECT 67.925 1.92 67.935 2.563 ;
      RECT 67.92 1.92 67.925 2.483 ;
      RECT 67.915 1.92 67.92 2.448 ;
      RECT 67.91 1.92 67.915 2.423 ;
      RECT 67.905 1.92 67.91 2.408 ;
      RECT 67.9 1.92 67.905 2.378 ;
      RECT 67.895 1.92 67.9 2.355 ;
      RECT 67.89 1.92 67.895 2.328 ;
      RECT 67.86 1.92 67.875 2.315 ;
      RECT 67.015 3.455 67.2 3.665 ;
      RECT 67.005 3.46 67.215 3.658 ;
      RECT 67.005 3.46 67.235 3.63 ;
      RECT 67.005 3.46 67.25 3.609 ;
      RECT 67.005 3.46 67.265 3.607 ;
      RECT 67.005 3.46 67.275 3.606 ;
      RECT 67.005 3.46 67.305 3.603 ;
      RECT 67.655 3.305 67.915 3.565 ;
      RECT 67.615 3.352 67.915 3.548 ;
      RECT 67.606 3.36 67.615 3.551 ;
      RECT 67.2 3.453 67.915 3.548 ;
      RECT 67.52 3.378 67.606 3.558 ;
      RECT 67.215 3.45 67.915 3.548 ;
      RECT 67.461 3.4 67.52 3.57 ;
      RECT 67.235 3.446 67.915 3.548 ;
      RECT 67.375 3.412 67.461 3.581 ;
      RECT 67.25 3.442 67.915 3.548 ;
      RECT 67.32 3.425 67.375 3.593 ;
      RECT 67.265 3.44 67.915 3.548 ;
      RECT 67.305 3.431 67.32 3.599 ;
      RECT 67.275 3.436 67.915 3.548 ;
      RECT 67.42 2.96 67.68 3.22 ;
      RECT 67.42 2.98 67.79 3.19 ;
      RECT 67.42 2.985 67.8 3.185 ;
      RECT 67.611 2.399 67.69 2.63 ;
      RECT 67.525 2.402 67.74 2.625 ;
      RECT 67.52 2.402 67.74 2.62 ;
      RECT 67.52 2.407 67.75 2.618 ;
      RECT 67.495 2.407 67.75 2.615 ;
      RECT 67.495 2.415 67.76 2.613 ;
      RECT 67.375 2.35 67.635 2.61 ;
      RECT 67.375 2.397 67.685 2.61 ;
      RECT 66.63 2.97 66.635 3.23 ;
      RECT 66.46 2.74 66.465 3.23 ;
      RECT 66.345 2.98 66.35 3.205 ;
      RECT 67.055 2.075 67.06 2.285 ;
      RECT 67.06 2.08 67.075 2.28 ;
      RECT 66.995 2.075 67.055 2.293 ;
      RECT 66.98 2.075 66.995 2.303 ;
      RECT 66.93 2.075 66.98 2.32 ;
      RECT 66.91 2.075 66.93 2.343 ;
      RECT 66.895 2.075 66.91 2.355 ;
      RECT 66.875 2.075 66.895 2.365 ;
      RECT 66.865 2.08 66.875 2.374 ;
      RECT 66.86 2.09 66.865 2.379 ;
      RECT 66.855 2.102 66.86 2.383 ;
      RECT 66.845 2.125 66.855 2.388 ;
      RECT 66.84 2.14 66.845 2.392 ;
      RECT 66.835 2.157 66.84 2.395 ;
      RECT 66.83 2.165 66.835 2.398 ;
      RECT 66.82 2.17 66.83 2.402 ;
      RECT 66.815 2.177 66.82 2.407 ;
      RECT 66.805 2.182 66.815 2.411 ;
      RECT 66.78 2.194 66.805 2.422 ;
      RECT 66.76 2.211 66.78 2.438 ;
      RECT 66.735 2.228 66.76 2.46 ;
      RECT 66.7 2.251 66.735 2.518 ;
      RECT 66.68 2.273 66.7 2.58 ;
      RECT 66.675 2.283 66.68 2.615 ;
      RECT 66.665 2.29 66.675 2.653 ;
      RECT 66.66 2.297 66.665 2.673 ;
      RECT 66.655 2.308 66.66 2.71 ;
      RECT 66.65 2.316 66.655 2.775 ;
      RECT 66.64 2.327 66.65 2.828 ;
      RECT 66.635 2.345 66.64 2.898 ;
      RECT 66.63 2.355 66.635 2.935 ;
      RECT 66.625 2.365 66.63 3.23 ;
      RECT 66.62 2.377 66.625 3.23 ;
      RECT 66.615 2.387 66.62 3.23 ;
      RECT 66.605 2.397 66.615 3.23 ;
      RECT 66.595 2.42 66.605 3.23 ;
      RECT 66.58 2.455 66.595 3.23 ;
      RECT 66.54 2.517 66.58 3.23 ;
      RECT 66.535 2.57 66.54 3.23 ;
      RECT 66.51 2.605 66.535 3.23 ;
      RECT 66.495 2.65 66.51 3.23 ;
      RECT 66.49 2.672 66.495 3.23 ;
      RECT 66.48 2.685 66.49 3.23 ;
      RECT 66.47 2.71 66.48 3.23 ;
      RECT 66.465 2.732 66.47 3.23 ;
      RECT 66.44 2.77 66.46 3.23 ;
      RECT 66.4 2.827 66.44 3.23 ;
      RECT 66.395 2.877 66.4 3.23 ;
      RECT 66.39 2.895 66.395 3.23 ;
      RECT 66.385 2.907 66.39 3.23 ;
      RECT 66.375 2.925 66.385 3.23 ;
      RECT 66.365 2.945 66.375 3.205 ;
      RECT 66.36 2.962 66.365 3.205 ;
      RECT 66.35 2.975 66.36 3.205 ;
      RECT 66.32 2.985 66.345 3.205 ;
      RECT 66.31 2.992 66.32 3.205 ;
      RECT 66.295 3.002 66.31 3.2 ;
      RECT 65.385 7.77 65.675 8 ;
      RECT 65.445 6.29 65.615 8 ;
      RECT 65.395 6.655 65.745 7.005 ;
      RECT 65.385 6.29 65.675 6.52 ;
      RECT 64.98 2.395 65.085 2.965 ;
      RECT 64.98 2.73 65.305 2.96 ;
      RECT 64.98 2.76 65.475 2.93 ;
      RECT 64.98 2.395 65.17 2.96 ;
      RECT 64.395 2.36 64.685 2.59 ;
      RECT 64.395 2.395 65.17 2.565 ;
      RECT 64.455 0.88 64.625 2.59 ;
      RECT 64.395 0.88 64.685 1.11 ;
      RECT 64.395 7.77 64.685 8 ;
      RECT 64.455 6.29 64.625 8 ;
      RECT 64.395 6.29 64.685 6.52 ;
      RECT 64.395 6.325 65.25 6.485 ;
      RECT 65.08 5.92 65.25 6.485 ;
      RECT 64.395 6.32 64.79 6.485 ;
      RECT 65.015 5.92 65.305 6.15 ;
      RECT 65.015 5.95 65.475 6.12 ;
      RECT 64.025 2.73 64.315 2.96 ;
      RECT 64.025 2.76 64.485 2.93 ;
      RECT 64.09 1.655 64.255 2.96 ;
      RECT 62.605 1.625 62.895 1.855 ;
      RECT 62.605 1.655 64.255 1.825 ;
      RECT 62.665 0.885 62.835 1.855 ;
      RECT 62.605 0.885 62.895 1.115 ;
      RECT 62.605 7.765 62.895 7.995 ;
      RECT 62.665 7.025 62.835 7.995 ;
      RECT 62.665 7.12 64.255 7.29 ;
      RECT 64.085 5.92 64.255 7.29 ;
      RECT 62.605 7.025 62.895 7.255 ;
      RECT 64.025 5.92 64.315 6.15 ;
      RECT 64.025 5.95 64.485 6.12 ;
      RECT 63.035 1.965 63.385 2.315 ;
      RECT 60.7 2.025 63.385 2.195 ;
      RECT 60.7 1.34 60.87 2.195 ;
      RECT 60.6 1.34 60.95 1.69 ;
      RECT 63.06 6.655 63.385 6.98 ;
      RECT 58.435 6.61 58.785 6.96 ;
      RECT 63.035 6.655 63.385 6.885 ;
      RECT 58.255 6.655 58.785 6.885 ;
      RECT 58.085 6.685 63.385 6.855 ;
      RECT 62.26 2.365 62.58 2.685 ;
      RECT 62.23 2.365 62.58 2.595 ;
      RECT 62.06 2.395 62.58 2.565 ;
      RECT 62.26 6.255 62.58 6.545 ;
      RECT 62.23 6.285 62.58 6.515 ;
      RECT 62.06 6.315 62.58 6.485 ;
      RECT 58.895 2.465 59.08 2.675 ;
      RECT 58.885 2.47 59.095 2.668 ;
      RECT 58.885 2.47 59.181 2.645 ;
      RECT 58.885 2.47 59.24 2.62 ;
      RECT 58.885 2.47 59.295 2.6 ;
      RECT 58.885 2.47 59.305 2.588 ;
      RECT 58.885 2.47 59.5 2.527 ;
      RECT 58.885 2.47 59.53 2.51 ;
      RECT 58.885 2.47 59.55 2.5 ;
      RECT 59.43 2.235 59.69 2.495 ;
      RECT 59.415 2.325 59.43 2.542 ;
      RECT 58.95 2.457 59.69 2.495 ;
      RECT 59.401 2.336 59.415 2.548 ;
      RECT 58.99 2.45 59.69 2.495 ;
      RECT 59.315 2.376 59.401 2.567 ;
      RECT 59.24 2.437 59.69 2.495 ;
      RECT 59.31 2.412 59.315 2.584 ;
      RECT 59.295 2.422 59.69 2.495 ;
      RECT 59.305 2.417 59.31 2.586 ;
      RECT 59.6 2.922 59.605 3.014 ;
      RECT 59.595 2.9 59.6 3.031 ;
      RECT 59.59 2.89 59.595 3.043 ;
      RECT 59.58 2.881 59.59 3.053 ;
      RECT 59.575 2.876 59.58 3.061 ;
      RECT 59.57 2.735 59.575 3.064 ;
      RECT 59.536 2.735 59.57 3.075 ;
      RECT 59.45 2.735 59.536 3.11 ;
      RECT 59.37 2.735 59.45 3.158 ;
      RECT 59.341 2.735 59.37 3.182 ;
      RECT 59.255 2.735 59.341 3.188 ;
      RECT 59.25 2.919 59.255 3.193 ;
      RECT 59.215 2.93 59.25 3.196 ;
      RECT 59.19 2.945 59.215 3.2 ;
      RECT 59.176 2.954 59.19 3.202 ;
      RECT 59.09 2.981 59.176 3.208 ;
      RECT 59.025 3.022 59.09 3.217 ;
      RECT 59.01 3.042 59.025 3.222 ;
      RECT 58.98 3.052 59.01 3.225 ;
      RECT 58.975 3.062 58.98 3.228 ;
      RECT 58.945 3.067 58.975 3.23 ;
      RECT 58.925 3.072 58.945 3.234 ;
      RECT 58.84 3.075 58.925 3.241 ;
      RECT 58.825 3.072 58.84 3.247 ;
      RECT 58.815 3.069 58.825 3.249 ;
      RECT 58.795 3.066 58.815 3.251 ;
      RECT 58.775 3.062 58.795 3.252 ;
      RECT 58.76 3.058 58.775 3.254 ;
      RECT 58.75 3.055 58.76 3.255 ;
      RECT 58.71 3.049 58.75 3.253 ;
      RECT 58.7 3.044 58.71 3.251 ;
      RECT 58.685 3.041 58.7 3.247 ;
      RECT 58.66 3.036 58.685 3.24 ;
      RECT 58.61 3.027 58.66 3.228 ;
      RECT 58.54 3.013 58.61 3.21 ;
      RECT 58.482 2.998 58.54 3.192 ;
      RECT 58.396 2.981 58.482 3.172 ;
      RECT 58.31 2.96 58.396 3.147 ;
      RECT 58.26 2.945 58.31 3.128 ;
      RECT 58.256 2.939 58.26 3.12 ;
      RECT 58.17 2.929 58.256 3.107 ;
      RECT 58.135 2.914 58.17 3.09 ;
      RECT 58.12 2.907 58.135 3.083 ;
      RECT 58.06 2.895 58.12 3.071 ;
      RECT 58.04 2.882 58.06 3.059 ;
      RECT 58 2.873 58.04 3.051 ;
      RECT 57.995 2.865 58 3.044 ;
      RECT 57.915 2.855 57.995 3.03 ;
      RECT 57.9 2.842 57.915 3.015 ;
      RECT 57.895 2.84 57.9 3.013 ;
      RECT 57.816 2.828 57.895 3 ;
      RECT 57.73 2.803 57.816 2.975 ;
      RECT 57.715 2.772 57.73 2.96 ;
      RECT 57.7 2.747 57.715 2.956 ;
      RECT 57.685 2.74 57.7 2.952 ;
      RECT 57.51 2.745 57.515 2.948 ;
      RECT 57.505 2.75 57.51 2.943 ;
      RECT 57.515 2.74 57.685 2.95 ;
      RECT 58.23 2.5 58.335 2.76 ;
      RECT 59.045 2.025 59.05 2.25 ;
      RECT 59.175 2.025 59.23 2.235 ;
      RECT 59.23 2.03 59.24 2.228 ;
      RECT 59.136 2.025 59.175 2.238 ;
      RECT 59.05 2.025 59.136 2.245 ;
      RECT 59.03 2.03 59.045 2.251 ;
      RECT 59.02 2.07 59.03 2.253 ;
      RECT 58.99 2.08 59.02 2.255 ;
      RECT 58.985 2.085 58.99 2.257 ;
      RECT 58.96 2.09 58.985 2.259 ;
      RECT 58.945 2.095 58.96 2.261 ;
      RECT 58.93 2.097 58.945 2.263 ;
      RECT 58.925 2.102 58.93 2.265 ;
      RECT 58.875 2.11 58.925 2.268 ;
      RECT 58.85 2.119 58.875 2.273 ;
      RECT 58.84 2.126 58.85 2.278 ;
      RECT 58.835 2.129 58.84 2.282 ;
      RECT 58.815 2.132 58.835 2.291 ;
      RECT 58.785 2.14 58.815 2.311 ;
      RECT 58.756 2.153 58.785 2.333 ;
      RECT 58.67 2.187 58.756 2.377 ;
      RECT 58.665 2.213 58.67 2.415 ;
      RECT 58.66 2.217 58.665 2.424 ;
      RECT 58.625 2.23 58.66 2.457 ;
      RECT 58.615 2.244 58.625 2.495 ;
      RECT 58.61 2.248 58.615 2.508 ;
      RECT 58.605 2.252 58.61 2.513 ;
      RECT 58.595 2.26 58.605 2.525 ;
      RECT 58.59 2.267 58.595 2.54 ;
      RECT 58.565 2.28 58.59 2.565 ;
      RECT 58.525 2.309 58.565 2.62 ;
      RECT 58.51 2.334 58.525 2.675 ;
      RECT 58.5 2.345 58.51 2.698 ;
      RECT 58.495 2.352 58.5 2.71 ;
      RECT 58.49 2.356 58.495 2.718 ;
      RECT 58.435 2.384 58.49 2.76 ;
      RECT 58.415 2.42 58.435 2.76 ;
      RECT 58.4 2.435 58.415 2.76 ;
      RECT 58.345 2.467 58.4 2.76 ;
      RECT 58.335 2.497 58.345 2.76 ;
      RECT 57.945 2.112 58.13 2.35 ;
      RECT 57.93 2.114 58.14 2.345 ;
      RECT 57.815 2.06 58.075 2.32 ;
      RECT 57.81 2.097 58.075 2.274 ;
      RECT 57.805 2.107 58.075 2.271 ;
      RECT 57.8 2.147 58.14 2.265 ;
      RECT 57.795 2.18 58.14 2.255 ;
      RECT 57.805 2.122 58.155 2.193 ;
      RECT 58.102 3.22 58.115 3.75 ;
      RECT 58.016 3.22 58.115 3.749 ;
      RECT 58.016 3.22 58.12 3.748 ;
      RECT 57.93 3.22 58.12 3.746 ;
      RECT 57.925 3.22 58.12 3.743 ;
      RECT 57.925 3.22 58.13 3.741 ;
      RECT 57.92 3.512 58.13 3.738 ;
      RECT 57.92 3.522 58.135 3.735 ;
      RECT 57.92 3.59 58.14 3.731 ;
      RECT 57.91 3.595 58.14 3.73 ;
      RECT 57.91 3.687 58.145 3.727 ;
      RECT 57.895 3.22 58.155 3.48 ;
      RECT 57.825 7.765 58.115 7.995 ;
      RECT 57.885 7.025 58.055 7.995 ;
      RECT 57.8 7.055 58.14 7.4 ;
      RECT 57.825 7.025 58.115 7.4 ;
      RECT 57.125 2.21 57.17 3.745 ;
      RECT 57.325 2.21 57.355 2.425 ;
      RECT 55.7 1.95 55.82 2.16 ;
      RECT 55.36 1.9 55.62 2.16 ;
      RECT 55.36 1.945 55.655 2.15 ;
      RECT 57.365 2.226 57.37 2.28 ;
      RECT 57.36 2.219 57.365 2.413 ;
      RECT 57.355 2.213 57.36 2.42 ;
      RECT 57.31 2.21 57.325 2.433 ;
      RECT 57.305 2.21 57.31 2.455 ;
      RECT 57.3 2.21 57.305 2.503 ;
      RECT 57.295 2.21 57.3 2.523 ;
      RECT 57.285 2.21 57.295 2.63 ;
      RECT 57.28 2.21 57.285 2.693 ;
      RECT 57.275 2.21 57.28 2.75 ;
      RECT 57.27 2.21 57.275 2.758 ;
      RECT 57.255 2.21 57.27 2.865 ;
      RECT 57.245 2.21 57.255 3 ;
      RECT 57.235 2.21 57.245 3.11 ;
      RECT 57.225 2.21 57.235 3.167 ;
      RECT 57.22 2.21 57.225 3.207 ;
      RECT 57.215 2.21 57.22 3.243 ;
      RECT 57.205 2.21 57.215 3.283 ;
      RECT 57.2 2.21 57.205 3.325 ;
      RECT 57.18 2.21 57.2 3.39 ;
      RECT 57.185 3.535 57.19 3.715 ;
      RECT 57.18 3.517 57.185 3.723 ;
      RECT 57.175 2.21 57.18 3.453 ;
      RECT 57.175 3.497 57.18 3.73 ;
      RECT 57.17 2.21 57.175 3.74 ;
      RECT 57.115 2.21 57.125 2.51 ;
      RECT 57.12 2.757 57.125 3.745 ;
      RECT 57.115 2.822 57.12 3.745 ;
      RECT 57.11 2.211 57.115 2.5 ;
      RECT 57.105 2.887 57.115 3.745 ;
      RECT 57.1 2.212 57.11 2.49 ;
      RECT 57.09 3 57.105 3.745 ;
      RECT 57.095 2.213 57.1 2.48 ;
      RECT 57.075 2.214 57.095 2.458 ;
      RECT 57.08 3.097 57.09 3.745 ;
      RECT 57.075 3.172 57.08 3.745 ;
      RECT 57.065 2.213 57.075 2.435 ;
      RECT 57.07 3.215 57.075 3.745 ;
      RECT 57.065 3.242 57.07 3.745 ;
      RECT 57.055 2.211 57.065 2.423 ;
      RECT 57.06 3.285 57.065 3.745 ;
      RECT 57.055 3.312 57.06 3.745 ;
      RECT 57.045 2.21 57.055 2.41 ;
      RECT 57.05 3.327 57.055 3.745 ;
      RECT 57.01 3.385 57.05 3.745 ;
      RECT 57.04 2.209 57.045 2.395 ;
      RECT 57.035 2.207 57.04 2.388 ;
      RECT 57.025 2.204 57.035 2.378 ;
      RECT 57.02 2.201 57.025 2.363 ;
      RECT 57.005 2.197 57.02 2.356 ;
      RECT 57 3.44 57.01 3.745 ;
      RECT 57 2.194 57.005 2.351 ;
      RECT 56.985 2.19 57 2.345 ;
      RECT 56.995 3.457 57 3.745 ;
      RECT 56.985 3.52 56.995 3.745 ;
      RECT 56.905 2.175 56.985 2.325 ;
      RECT 56.98 3.527 56.985 3.74 ;
      RECT 56.975 3.535 56.98 3.73 ;
      RECT 56.895 2.161 56.905 2.309 ;
      RECT 56.88 2.157 56.895 2.307 ;
      RECT 56.87 2.152 56.88 2.303 ;
      RECT 56.845 2.145 56.87 2.295 ;
      RECT 56.84 2.14 56.845 2.29 ;
      RECT 56.83 2.14 56.84 2.288 ;
      RECT 56.82 2.138 56.83 2.286 ;
      RECT 56.79 2.13 56.82 2.28 ;
      RECT 56.775 2.122 56.79 2.273 ;
      RECT 56.755 2.117 56.775 2.266 ;
      RECT 56.75 2.113 56.755 2.261 ;
      RECT 56.72 2.106 56.75 2.255 ;
      RECT 56.695 2.097 56.72 2.245 ;
      RECT 56.665 2.09 56.695 2.237 ;
      RECT 56.64 2.08 56.665 2.228 ;
      RECT 56.625 2.072 56.64 2.222 ;
      RECT 56.6 2.067 56.625 2.217 ;
      RECT 56.59 2.063 56.6 2.212 ;
      RECT 56.57 2.058 56.59 2.207 ;
      RECT 56.535 2.053 56.57 2.2 ;
      RECT 56.475 2.048 56.535 2.193 ;
      RECT 56.462 2.044 56.475 2.191 ;
      RECT 56.376 2.039 56.462 2.188 ;
      RECT 56.29 2.029 56.376 2.184 ;
      RECT 56.249 2.022 56.29 2.181 ;
      RECT 56.163 2.015 56.249 2.178 ;
      RECT 56.077 2.005 56.163 2.174 ;
      RECT 55.991 1.995 56.077 2.169 ;
      RECT 55.905 1.985 55.991 2.165 ;
      RECT 55.895 1.97 55.905 2.163 ;
      RECT 55.885 1.955 55.895 2.163 ;
      RECT 55.82 1.95 55.885 2.162 ;
      RECT 55.655 1.947 55.7 2.155 ;
      RECT 56.9 2.852 56.905 3.043 ;
      RECT 56.895 2.847 56.9 3.05 ;
      RECT 56.881 2.845 56.895 3.056 ;
      RECT 56.795 2.845 56.881 3.058 ;
      RECT 56.791 2.845 56.795 3.061 ;
      RECT 56.705 2.845 56.791 3.079 ;
      RECT 56.695 2.85 56.705 3.098 ;
      RECT 56.685 2.905 56.695 3.102 ;
      RECT 56.66 2.92 56.685 3.109 ;
      RECT 56.62 2.94 56.66 3.122 ;
      RECT 56.615 2.952 56.62 3.132 ;
      RECT 56.6 2.958 56.615 3.137 ;
      RECT 56.595 2.963 56.6 3.141 ;
      RECT 56.575 2.97 56.595 3.146 ;
      RECT 56.505 2.995 56.575 3.163 ;
      RECT 56.465 3.023 56.505 3.183 ;
      RECT 56.46 3.033 56.465 3.191 ;
      RECT 56.44 3.04 56.46 3.193 ;
      RECT 56.435 3.047 56.44 3.196 ;
      RECT 56.405 3.055 56.435 3.199 ;
      RECT 56.4 3.06 56.405 3.203 ;
      RECT 56.326 3.064 56.4 3.211 ;
      RECT 56.24 3.073 56.326 3.227 ;
      RECT 56.236 3.078 56.24 3.236 ;
      RECT 56.15 3.083 56.236 3.246 ;
      RECT 56.11 3.091 56.15 3.258 ;
      RECT 56.06 3.097 56.11 3.265 ;
      RECT 55.975 3.106 56.06 3.28 ;
      RECT 55.9 3.117 55.975 3.298 ;
      RECT 55.865 3.124 55.9 3.308 ;
      RECT 55.79 3.132 55.865 3.313 ;
      RECT 55.735 3.141 55.79 3.313 ;
      RECT 55.71 3.146 55.735 3.311 ;
      RECT 55.7 3.149 55.71 3.309 ;
      RECT 55.665 3.151 55.7 3.307 ;
      RECT 55.635 3.153 55.665 3.303 ;
      RECT 55.59 3.152 55.635 3.299 ;
      RECT 55.57 3.147 55.59 3.296 ;
      RECT 55.52 3.132 55.57 3.293 ;
      RECT 55.51 3.117 55.52 3.288 ;
      RECT 55.46 3.102 55.51 3.278 ;
      RECT 55.41 3.077 55.46 3.258 ;
      RECT 55.4 3.062 55.41 3.24 ;
      RECT 55.395 3.06 55.4 3.234 ;
      RECT 55.375 3.055 55.395 3.229 ;
      RECT 55.37 3.047 55.375 3.223 ;
      RECT 55.355 3.041 55.37 3.216 ;
      RECT 55.35 3.036 55.355 3.208 ;
      RECT 55.33 3.031 55.35 3.2 ;
      RECT 55.315 3.024 55.33 3.193 ;
      RECT 55.3 3.018 55.315 3.184 ;
      RECT 55.295 3.012 55.3 3.177 ;
      RECT 55.25 2.987 55.295 3.163 ;
      RECT 55.235 2.957 55.25 3.145 ;
      RECT 55.22 2.94 55.235 3.136 ;
      RECT 55.195 2.92 55.22 3.124 ;
      RECT 55.155 2.89 55.195 3.104 ;
      RECT 55.145 2.86 55.155 3.089 ;
      RECT 55.13 2.85 55.145 3.082 ;
      RECT 55.075 2.815 55.13 3.061 ;
      RECT 55.06 2.778 55.075 3.04 ;
      RECT 55.05 2.765 55.06 3.032 ;
      RECT 55 2.735 55.05 3.014 ;
      RECT 54.985 2.665 55 2.995 ;
      RECT 54.94 2.665 54.985 2.978 ;
      RECT 54.915 2.665 54.94 2.96 ;
      RECT 54.905 2.665 54.915 2.953 ;
      RECT 54.826 2.665 54.905 2.946 ;
      RECT 54.74 2.665 54.826 2.938 ;
      RECT 54.725 2.697 54.74 2.933 ;
      RECT 54.65 2.707 54.725 2.929 ;
      RECT 54.63 2.717 54.65 2.924 ;
      RECT 54.605 2.717 54.63 2.921 ;
      RECT 54.595 2.707 54.605 2.92 ;
      RECT 54.585 2.68 54.595 2.919 ;
      RECT 54.545 2.675 54.585 2.917 ;
      RECT 54.5 2.675 54.545 2.913 ;
      RECT 54.475 2.675 54.5 2.908 ;
      RECT 54.425 2.675 54.475 2.895 ;
      RECT 54.385 2.68 54.395 2.88 ;
      RECT 54.395 2.675 54.425 2.885 ;
      RECT 56.38 2.455 56.64 2.715 ;
      RECT 56.375 2.477 56.64 2.673 ;
      RECT 55.615 2.305 55.835 2.67 ;
      RECT 55.597 2.392 55.835 2.669 ;
      RECT 55.58 2.397 55.835 2.666 ;
      RECT 55.58 2.397 55.855 2.665 ;
      RECT 55.55 2.407 55.855 2.663 ;
      RECT 55.545 2.422 55.855 2.659 ;
      RECT 55.545 2.422 55.86 2.658 ;
      RECT 55.54 2.48 55.86 2.656 ;
      RECT 55.54 2.48 55.87 2.653 ;
      RECT 55.535 2.545 55.87 2.648 ;
      RECT 55.615 2.305 55.875 2.565 ;
      RECT 54.36 2.135 54.62 2.395 ;
      RECT 54.36 2.178 54.706 2.369 ;
      RECT 54.36 2.178 54.75 2.368 ;
      RECT 54.36 2.178 54.77 2.366 ;
      RECT 54.36 2.178 54.87 2.365 ;
      RECT 54.36 2.178 54.89 2.363 ;
      RECT 54.36 2.178 54.9 2.358 ;
      RECT 54.77 2.145 54.96 2.355 ;
      RECT 54.77 2.147 54.965 2.353 ;
      RECT 54.76 2.152 54.97 2.345 ;
      RECT 54.706 2.176 54.97 2.345 ;
      RECT 54.75 2.17 54.76 2.367 ;
      RECT 54.76 2.15 54.965 2.353 ;
      RECT 53.715 3.21 53.92 3.44 ;
      RECT 53.655 3.16 53.71 3.42 ;
      RECT 53.715 3.16 53.915 3.44 ;
      RECT 54.685 3.475 54.69 3.502 ;
      RECT 54.675 3.385 54.685 3.507 ;
      RECT 54.67 3.307 54.675 3.513 ;
      RECT 54.66 3.297 54.67 3.52 ;
      RECT 54.655 3.287 54.66 3.526 ;
      RECT 54.645 3.282 54.655 3.528 ;
      RECT 54.63 3.274 54.645 3.536 ;
      RECT 54.615 3.265 54.63 3.548 ;
      RECT 54.605 3.257 54.615 3.558 ;
      RECT 54.57 3.175 54.605 3.576 ;
      RECT 54.535 3.175 54.57 3.595 ;
      RECT 54.52 3.175 54.535 3.603 ;
      RECT 54.465 3.175 54.52 3.603 ;
      RECT 54.431 3.175 54.465 3.594 ;
      RECT 54.345 3.175 54.431 3.57 ;
      RECT 54.335 3.235 54.345 3.552 ;
      RECT 54.295 3.237 54.335 3.543 ;
      RECT 54.29 3.239 54.295 3.533 ;
      RECT 54.27 3.241 54.29 3.528 ;
      RECT 54.26 3.244 54.27 3.523 ;
      RECT 54.25 3.245 54.26 3.518 ;
      RECT 54.226 3.246 54.25 3.51 ;
      RECT 54.14 3.251 54.226 3.488 ;
      RECT 54.085 3.25 54.14 3.461 ;
      RECT 54.07 3.243 54.085 3.448 ;
      RECT 54.035 3.238 54.07 3.444 ;
      RECT 53.98 3.23 54.035 3.443 ;
      RECT 53.92 3.217 53.98 3.441 ;
      RECT 53.71 3.16 53.715 3.428 ;
      RECT 53.785 2.53 53.97 2.74 ;
      RECT 53.775 2.535 53.985 2.733 ;
      RECT 53.815 2.44 54.075 2.7 ;
      RECT 53.77 2.597 54.075 2.623 ;
      RECT 53.115 2.39 53.12 3.19 ;
      RECT 53.06 2.44 53.09 3.19 ;
      RECT 53.05 2.44 53.055 2.75 ;
      RECT 53.035 2.44 53.04 2.745 ;
      RECT 52.58 2.485 52.595 2.7 ;
      RECT 52.51 2.485 52.595 2.695 ;
      RECT 53.775 2.065 53.845 2.275 ;
      RECT 53.845 2.072 53.855 2.27 ;
      RECT 53.741 2.065 53.775 2.282 ;
      RECT 53.655 2.065 53.741 2.306 ;
      RECT 53.645 2.07 53.655 2.325 ;
      RECT 53.64 2.082 53.645 2.328 ;
      RECT 53.625 2.097 53.64 2.332 ;
      RECT 53.62 2.115 53.625 2.336 ;
      RECT 53.58 2.125 53.62 2.345 ;
      RECT 53.565 2.132 53.58 2.357 ;
      RECT 53.55 2.137 53.565 2.362 ;
      RECT 53.535 2.14 53.55 2.367 ;
      RECT 53.525 2.142 53.535 2.371 ;
      RECT 53.49 2.149 53.525 2.379 ;
      RECT 53.455 2.157 53.49 2.393 ;
      RECT 53.445 2.163 53.455 2.402 ;
      RECT 53.44 2.165 53.445 2.404 ;
      RECT 53.42 2.168 53.44 2.41 ;
      RECT 53.39 2.175 53.42 2.421 ;
      RECT 53.38 2.181 53.39 2.428 ;
      RECT 53.355 2.184 53.38 2.435 ;
      RECT 53.345 2.188 53.355 2.443 ;
      RECT 53.34 2.189 53.345 2.465 ;
      RECT 53.335 2.19 53.34 2.48 ;
      RECT 53.33 2.191 53.335 2.495 ;
      RECT 53.325 2.192 53.33 2.51 ;
      RECT 53.32 2.193 53.325 2.54 ;
      RECT 53.31 2.195 53.32 2.573 ;
      RECT 53.295 2.199 53.31 2.62 ;
      RECT 53.285 2.202 53.295 2.665 ;
      RECT 53.28 2.205 53.285 2.693 ;
      RECT 53.27 2.207 53.28 2.72 ;
      RECT 53.265 2.21 53.27 2.755 ;
      RECT 53.235 2.215 53.265 2.813 ;
      RECT 53.23 2.22 53.235 2.898 ;
      RECT 53.225 2.222 53.23 2.933 ;
      RECT 53.22 2.224 53.225 3.015 ;
      RECT 53.215 2.226 53.22 3.103 ;
      RECT 53.205 2.228 53.215 3.185 ;
      RECT 53.19 2.242 53.205 3.19 ;
      RECT 53.155 2.287 53.19 3.19 ;
      RECT 53.145 2.327 53.155 3.19 ;
      RECT 53.13 2.355 53.145 3.19 ;
      RECT 53.125 2.372 53.13 3.19 ;
      RECT 53.12 2.38 53.125 3.19 ;
      RECT 53.11 2.395 53.115 3.19 ;
      RECT 53.105 2.402 53.11 3.19 ;
      RECT 53.095 2.422 53.105 3.19 ;
      RECT 53.09 2.435 53.095 3.19 ;
      RECT 53.055 2.44 53.06 2.775 ;
      RECT 53.04 2.83 53.06 3.19 ;
      RECT 53.04 2.44 53.05 2.748 ;
      RECT 53.035 2.87 53.04 3.19 ;
      RECT 52.985 2.44 53.035 2.743 ;
      RECT 53.03 2.907 53.035 3.19 ;
      RECT 53.02 2.93 53.03 3.19 ;
      RECT 53.015 2.975 53.02 3.19 ;
      RECT 53.005 2.985 53.015 3.183 ;
      RECT 52.931 2.44 52.985 2.737 ;
      RECT 52.845 2.44 52.931 2.73 ;
      RECT 52.796 2.487 52.845 2.723 ;
      RECT 52.71 2.495 52.796 2.716 ;
      RECT 52.695 2.492 52.71 2.711 ;
      RECT 52.681 2.485 52.695 2.71 ;
      RECT 52.595 2.485 52.681 2.705 ;
      RECT 52.5 2.49 52.51 2.69 ;
      RECT 52.09 1.92 52.105 2.32 ;
      RECT 52.285 1.92 52.29 2.18 ;
      RECT 52.03 1.92 52.075 2.18 ;
      RECT 52.485 3.225 52.49 3.43 ;
      RECT 52.48 3.215 52.485 3.435 ;
      RECT 52.475 3.202 52.48 3.44 ;
      RECT 52.47 3.182 52.475 3.44 ;
      RECT 52.445 3.135 52.47 3.44 ;
      RECT 52.41 3.05 52.445 3.44 ;
      RECT 52.405 2.987 52.41 3.44 ;
      RECT 52.4 2.972 52.405 3.44 ;
      RECT 52.385 2.932 52.4 3.44 ;
      RECT 52.38 2.907 52.385 3.44 ;
      RECT 52.37 2.89 52.38 3.44 ;
      RECT 52.335 2.812 52.37 3.44 ;
      RECT 52.33 2.755 52.335 3.44 ;
      RECT 52.325 2.742 52.33 3.44 ;
      RECT 52.315 2.72 52.325 3.44 ;
      RECT 52.305 2.685 52.315 3.44 ;
      RECT 52.295 2.655 52.305 3.44 ;
      RECT 52.285 2.57 52.295 3.083 ;
      RECT 52.292 3.215 52.295 3.44 ;
      RECT 52.29 3.225 52.292 3.44 ;
      RECT 52.28 3.235 52.29 3.435 ;
      RECT 52.275 1.92 52.285 2.315 ;
      RECT 52.28 2.447 52.285 3.058 ;
      RECT 52.275 2.345 52.28 3.041 ;
      RECT 52.265 1.92 52.275 3.017 ;
      RECT 52.26 1.92 52.265 2.988 ;
      RECT 52.255 1.92 52.26 2.978 ;
      RECT 52.235 1.92 52.255 2.94 ;
      RECT 52.23 1.92 52.235 2.898 ;
      RECT 52.225 1.92 52.23 2.878 ;
      RECT 52.195 1.92 52.225 2.828 ;
      RECT 52.185 1.92 52.195 2.775 ;
      RECT 52.18 1.92 52.185 2.748 ;
      RECT 52.175 1.92 52.18 2.733 ;
      RECT 52.165 1.92 52.175 2.71 ;
      RECT 52.155 1.92 52.165 2.685 ;
      RECT 52.15 1.92 52.155 2.625 ;
      RECT 52.14 1.92 52.15 2.563 ;
      RECT 52.135 1.92 52.14 2.483 ;
      RECT 52.13 1.92 52.135 2.448 ;
      RECT 52.125 1.92 52.13 2.423 ;
      RECT 52.12 1.92 52.125 2.408 ;
      RECT 52.115 1.92 52.12 2.378 ;
      RECT 52.11 1.92 52.115 2.355 ;
      RECT 52.105 1.92 52.11 2.328 ;
      RECT 52.075 1.92 52.09 2.315 ;
      RECT 51.23 3.455 51.415 3.665 ;
      RECT 51.22 3.46 51.43 3.658 ;
      RECT 51.22 3.46 51.45 3.63 ;
      RECT 51.22 3.46 51.465 3.609 ;
      RECT 51.22 3.46 51.48 3.607 ;
      RECT 51.22 3.46 51.49 3.606 ;
      RECT 51.22 3.46 51.52 3.603 ;
      RECT 51.87 3.305 52.13 3.565 ;
      RECT 51.83 3.352 52.13 3.548 ;
      RECT 51.821 3.36 51.83 3.551 ;
      RECT 51.415 3.453 52.13 3.548 ;
      RECT 51.735 3.378 51.821 3.558 ;
      RECT 51.43 3.45 52.13 3.548 ;
      RECT 51.676 3.4 51.735 3.57 ;
      RECT 51.45 3.446 52.13 3.548 ;
      RECT 51.59 3.412 51.676 3.581 ;
      RECT 51.465 3.442 52.13 3.548 ;
      RECT 51.535 3.425 51.59 3.593 ;
      RECT 51.48 3.44 52.13 3.548 ;
      RECT 51.52 3.431 51.535 3.599 ;
      RECT 51.49 3.436 52.13 3.548 ;
      RECT 51.635 2.96 51.895 3.22 ;
      RECT 51.635 2.98 52.005 3.19 ;
      RECT 51.635 2.985 52.015 3.185 ;
      RECT 51.826 2.399 51.905 2.63 ;
      RECT 51.74 2.402 51.955 2.625 ;
      RECT 51.735 2.402 51.955 2.62 ;
      RECT 51.735 2.407 51.965 2.618 ;
      RECT 51.71 2.407 51.965 2.615 ;
      RECT 51.71 2.415 51.975 2.613 ;
      RECT 51.59 2.35 51.85 2.61 ;
      RECT 51.59 2.397 51.9 2.61 ;
      RECT 50.845 2.97 50.85 3.23 ;
      RECT 50.675 2.74 50.68 3.23 ;
      RECT 50.56 2.98 50.565 3.205 ;
      RECT 51.27 2.075 51.275 2.285 ;
      RECT 51.275 2.08 51.29 2.28 ;
      RECT 51.21 2.075 51.27 2.293 ;
      RECT 51.195 2.075 51.21 2.303 ;
      RECT 51.145 2.075 51.195 2.32 ;
      RECT 51.125 2.075 51.145 2.343 ;
      RECT 51.11 2.075 51.125 2.355 ;
      RECT 51.09 2.075 51.11 2.365 ;
      RECT 51.08 2.08 51.09 2.374 ;
      RECT 51.075 2.09 51.08 2.379 ;
      RECT 51.07 2.102 51.075 2.383 ;
      RECT 51.06 2.125 51.07 2.388 ;
      RECT 51.055 2.14 51.06 2.392 ;
      RECT 51.05 2.157 51.055 2.395 ;
      RECT 51.045 2.165 51.05 2.398 ;
      RECT 51.035 2.17 51.045 2.402 ;
      RECT 51.03 2.177 51.035 2.407 ;
      RECT 51.02 2.182 51.03 2.411 ;
      RECT 50.995 2.194 51.02 2.422 ;
      RECT 50.975 2.211 50.995 2.438 ;
      RECT 50.95 2.228 50.975 2.46 ;
      RECT 50.915 2.251 50.95 2.518 ;
      RECT 50.895 2.273 50.915 2.58 ;
      RECT 50.89 2.283 50.895 2.615 ;
      RECT 50.88 2.29 50.89 2.653 ;
      RECT 50.875 2.297 50.88 2.673 ;
      RECT 50.87 2.308 50.875 2.71 ;
      RECT 50.865 2.316 50.87 2.775 ;
      RECT 50.855 2.327 50.865 2.828 ;
      RECT 50.85 2.345 50.855 2.898 ;
      RECT 50.845 2.355 50.85 2.935 ;
      RECT 50.84 2.365 50.845 3.23 ;
      RECT 50.835 2.377 50.84 3.23 ;
      RECT 50.83 2.387 50.835 3.23 ;
      RECT 50.82 2.397 50.83 3.23 ;
      RECT 50.81 2.42 50.82 3.23 ;
      RECT 50.795 2.455 50.81 3.23 ;
      RECT 50.755 2.517 50.795 3.23 ;
      RECT 50.75 2.57 50.755 3.23 ;
      RECT 50.725 2.605 50.75 3.23 ;
      RECT 50.71 2.65 50.725 3.23 ;
      RECT 50.705 2.672 50.71 3.23 ;
      RECT 50.695 2.685 50.705 3.23 ;
      RECT 50.685 2.71 50.695 3.23 ;
      RECT 50.68 2.732 50.685 3.23 ;
      RECT 50.655 2.77 50.675 3.23 ;
      RECT 50.615 2.827 50.655 3.23 ;
      RECT 50.61 2.877 50.615 3.23 ;
      RECT 50.605 2.895 50.61 3.23 ;
      RECT 50.6 2.907 50.605 3.23 ;
      RECT 50.59 2.925 50.6 3.23 ;
      RECT 50.58 2.945 50.59 3.205 ;
      RECT 50.575 2.962 50.58 3.205 ;
      RECT 50.565 2.975 50.575 3.205 ;
      RECT 50.535 2.985 50.56 3.205 ;
      RECT 50.525 2.992 50.535 3.205 ;
      RECT 50.51 3.002 50.525 3.2 ;
      RECT 49.6 7.77 49.89 8 ;
      RECT 49.66 6.29 49.83 8 ;
      RECT 49.61 6.655 49.96 7.005 ;
      RECT 49.6 6.29 49.89 6.52 ;
      RECT 49.195 2.395 49.3 2.965 ;
      RECT 49.195 2.73 49.52 2.96 ;
      RECT 49.195 2.76 49.69 2.93 ;
      RECT 49.195 2.395 49.385 2.96 ;
      RECT 48.61 2.36 48.9 2.59 ;
      RECT 48.61 2.395 49.385 2.565 ;
      RECT 48.67 0.88 48.84 2.59 ;
      RECT 48.61 0.88 48.9 1.11 ;
      RECT 48.61 7.77 48.9 8 ;
      RECT 48.67 6.29 48.84 8 ;
      RECT 48.61 6.29 48.9 6.52 ;
      RECT 48.61 6.325 49.465 6.485 ;
      RECT 49.295 5.92 49.465 6.485 ;
      RECT 48.61 6.32 49.005 6.485 ;
      RECT 49.23 5.92 49.52 6.15 ;
      RECT 49.23 5.95 49.69 6.12 ;
      RECT 48.24 2.73 48.53 2.96 ;
      RECT 48.24 2.76 48.7 2.93 ;
      RECT 48.305 1.655 48.47 2.96 ;
      RECT 46.82 1.625 47.11 1.855 ;
      RECT 46.82 1.655 48.47 1.825 ;
      RECT 46.88 0.885 47.05 1.855 ;
      RECT 46.82 0.885 47.11 1.115 ;
      RECT 46.82 7.765 47.11 7.995 ;
      RECT 46.88 7.025 47.05 7.995 ;
      RECT 46.88 7.12 48.47 7.29 ;
      RECT 48.3 5.92 48.47 7.29 ;
      RECT 46.82 7.025 47.11 7.255 ;
      RECT 48.24 5.92 48.53 6.15 ;
      RECT 48.24 5.95 48.7 6.12 ;
      RECT 47.25 1.965 47.6 2.315 ;
      RECT 44.915 2.025 47.6 2.195 ;
      RECT 44.915 1.34 45.085 2.195 ;
      RECT 44.815 1.34 45.165 1.69 ;
      RECT 47.275 6.655 47.6 6.98 ;
      RECT 42.705 6.615 43.055 6.965 ;
      RECT 47.25 6.655 47.6 6.885 ;
      RECT 42.47 6.655 43.055 6.885 ;
      RECT 42.3 6.685 47.6 6.855 ;
      RECT 46.475 2.365 46.795 2.685 ;
      RECT 46.445 2.365 46.795 2.595 ;
      RECT 46.275 2.395 46.795 2.565 ;
      RECT 46.475 6.255 46.795 6.545 ;
      RECT 46.445 6.285 46.795 6.515 ;
      RECT 46.275 6.315 46.795 6.485 ;
      RECT 43.11 2.465 43.295 2.675 ;
      RECT 43.1 2.47 43.31 2.668 ;
      RECT 43.1 2.47 43.396 2.645 ;
      RECT 43.1 2.47 43.455 2.62 ;
      RECT 43.1 2.47 43.51 2.6 ;
      RECT 43.1 2.47 43.52 2.588 ;
      RECT 43.1 2.47 43.715 2.527 ;
      RECT 43.1 2.47 43.745 2.51 ;
      RECT 43.1 2.47 43.765 2.5 ;
      RECT 43.645 2.235 43.905 2.495 ;
      RECT 43.63 2.325 43.645 2.542 ;
      RECT 43.165 2.457 43.905 2.495 ;
      RECT 43.616 2.336 43.63 2.548 ;
      RECT 43.205 2.45 43.905 2.495 ;
      RECT 43.53 2.376 43.616 2.567 ;
      RECT 43.455 2.437 43.905 2.495 ;
      RECT 43.525 2.412 43.53 2.584 ;
      RECT 43.51 2.422 43.905 2.495 ;
      RECT 43.52 2.417 43.525 2.586 ;
      RECT 43.815 2.922 43.82 3.014 ;
      RECT 43.81 2.9 43.815 3.031 ;
      RECT 43.805 2.89 43.81 3.043 ;
      RECT 43.795 2.881 43.805 3.053 ;
      RECT 43.79 2.876 43.795 3.061 ;
      RECT 43.785 2.735 43.79 3.064 ;
      RECT 43.751 2.735 43.785 3.075 ;
      RECT 43.665 2.735 43.751 3.11 ;
      RECT 43.585 2.735 43.665 3.158 ;
      RECT 43.556 2.735 43.585 3.182 ;
      RECT 43.47 2.735 43.556 3.188 ;
      RECT 43.465 2.919 43.47 3.193 ;
      RECT 43.43 2.93 43.465 3.196 ;
      RECT 43.405 2.945 43.43 3.2 ;
      RECT 43.391 2.954 43.405 3.202 ;
      RECT 43.305 2.981 43.391 3.208 ;
      RECT 43.24 3.022 43.305 3.217 ;
      RECT 43.225 3.042 43.24 3.222 ;
      RECT 43.195 3.052 43.225 3.225 ;
      RECT 43.19 3.062 43.195 3.228 ;
      RECT 43.16 3.067 43.19 3.23 ;
      RECT 43.14 3.072 43.16 3.234 ;
      RECT 43.055 3.075 43.14 3.241 ;
      RECT 43.04 3.072 43.055 3.247 ;
      RECT 43.03 3.069 43.04 3.249 ;
      RECT 43.01 3.066 43.03 3.251 ;
      RECT 42.99 3.062 43.01 3.252 ;
      RECT 42.975 3.058 42.99 3.254 ;
      RECT 42.965 3.055 42.975 3.255 ;
      RECT 42.925 3.049 42.965 3.253 ;
      RECT 42.915 3.044 42.925 3.251 ;
      RECT 42.9 3.041 42.915 3.247 ;
      RECT 42.875 3.036 42.9 3.24 ;
      RECT 42.825 3.027 42.875 3.228 ;
      RECT 42.755 3.013 42.825 3.21 ;
      RECT 42.697 2.998 42.755 3.192 ;
      RECT 42.611 2.981 42.697 3.172 ;
      RECT 42.525 2.96 42.611 3.147 ;
      RECT 42.475 2.945 42.525 3.128 ;
      RECT 42.471 2.939 42.475 3.12 ;
      RECT 42.385 2.929 42.471 3.107 ;
      RECT 42.35 2.914 42.385 3.09 ;
      RECT 42.335 2.907 42.35 3.083 ;
      RECT 42.275 2.895 42.335 3.071 ;
      RECT 42.255 2.882 42.275 3.059 ;
      RECT 42.215 2.873 42.255 3.051 ;
      RECT 42.21 2.865 42.215 3.044 ;
      RECT 42.13 2.855 42.21 3.03 ;
      RECT 42.115 2.842 42.13 3.015 ;
      RECT 42.11 2.84 42.115 3.013 ;
      RECT 42.031 2.828 42.11 3 ;
      RECT 41.945 2.803 42.031 2.975 ;
      RECT 41.93 2.772 41.945 2.96 ;
      RECT 41.915 2.747 41.93 2.956 ;
      RECT 41.9 2.74 41.915 2.952 ;
      RECT 41.725 2.745 41.73 2.948 ;
      RECT 41.72 2.75 41.725 2.943 ;
      RECT 41.73 2.74 41.9 2.95 ;
      RECT 42.445 2.5 42.55 2.76 ;
      RECT 43.26 2.025 43.265 2.25 ;
      RECT 43.39 2.025 43.445 2.235 ;
      RECT 43.445 2.03 43.455 2.228 ;
      RECT 43.351 2.025 43.39 2.238 ;
      RECT 43.265 2.025 43.351 2.245 ;
      RECT 43.245 2.03 43.26 2.251 ;
      RECT 43.235 2.07 43.245 2.253 ;
      RECT 43.205 2.08 43.235 2.255 ;
      RECT 43.2 2.085 43.205 2.257 ;
      RECT 43.175 2.09 43.2 2.259 ;
      RECT 43.16 2.095 43.175 2.261 ;
      RECT 43.145 2.097 43.16 2.263 ;
      RECT 43.14 2.102 43.145 2.265 ;
      RECT 43.09 2.11 43.14 2.268 ;
      RECT 43.065 2.119 43.09 2.273 ;
      RECT 43.055 2.126 43.065 2.278 ;
      RECT 43.05 2.129 43.055 2.282 ;
      RECT 43.03 2.132 43.05 2.291 ;
      RECT 43 2.14 43.03 2.311 ;
      RECT 42.971 2.153 43 2.333 ;
      RECT 42.885 2.187 42.971 2.377 ;
      RECT 42.88 2.213 42.885 2.415 ;
      RECT 42.875 2.217 42.88 2.424 ;
      RECT 42.84 2.23 42.875 2.457 ;
      RECT 42.83 2.244 42.84 2.495 ;
      RECT 42.825 2.248 42.83 2.508 ;
      RECT 42.82 2.252 42.825 2.513 ;
      RECT 42.81 2.26 42.82 2.525 ;
      RECT 42.805 2.267 42.81 2.54 ;
      RECT 42.78 2.28 42.805 2.565 ;
      RECT 42.74 2.309 42.78 2.62 ;
      RECT 42.725 2.334 42.74 2.675 ;
      RECT 42.715 2.345 42.725 2.698 ;
      RECT 42.71 2.352 42.715 2.71 ;
      RECT 42.705 2.356 42.71 2.718 ;
      RECT 42.65 2.384 42.705 2.76 ;
      RECT 42.63 2.42 42.65 2.76 ;
      RECT 42.615 2.435 42.63 2.76 ;
      RECT 42.56 2.467 42.615 2.76 ;
      RECT 42.55 2.497 42.56 2.76 ;
      RECT 42.16 2.112 42.345 2.35 ;
      RECT 42.145 2.114 42.355 2.345 ;
      RECT 42.03 2.06 42.29 2.32 ;
      RECT 42.025 2.097 42.29 2.274 ;
      RECT 42.02 2.107 42.29 2.271 ;
      RECT 42.015 2.147 42.355 2.265 ;
      RECT 42.01 2.18 42.355 2.255 ;
      RECT 42.02 2.122 42.37 2.193 ;
      RECT 42.317 3.22 42.33 3.75 ;
      RECT 42.231 3.22 42.33 3.749 ;
      RECT 42.231 3.22 42.335 3.748 ;
      RECT 42.145 3.22 42.335 3.746 ;
      RECT 42.14 3.22 42.335 3.743 ;
      RECT 42.14 3.22 42.345 3.741 ;
      RECT 42.135 3.512 42.345 3.738 ;
      RECT 42.135 3.522 42.35 3.735 ;
      RECT 42.135 3.59 42.355 3.731 ;
      RECT 42.125 3.595 42.355 3.73 ;
      RECT 42.125 3.687 42.36 3.727 ;
      RECT 42.11 3.22 42.37 3.48 ;
      RECT 42.04 7.765 42.33 7.995 ;
      RECT 42.1 7.025 42.27 7.995 ;
      RECT 42.015 7.055 42.355 7.4 ;
      RECT 42.04 7.025 42.33 7.4 ;
      RECT 41.34 2.21 41.385 3.745 ;
      RECT 41.54 2.21 41.57 2.425 ;
      RECT 39.915 1.95 40.035 2.16 ;
      RECT 39.575 1.9 39.835 2.16 ;
      RECT 39.575 1.945 39.87 2.15 ;
      RECT 41.58 2.226 41.585 2.28 ;
      RECT 41.575 2.219 41.58 2.413 ;
      RECT 41.57 2.213 41.575 2.42 ;
      RECT 41.525 2.21 41.54 2.433 ;
      RECT 41.52 2.21 41.525 2.455 ;
      RECT 41.515 2.21 41.52 2.503 ;
      RECT 41.51 2.21 41.515 2.523 ;
      RECT 41.5 2.21 41.51 2.63 ;
      RECT 41.495 2.21 41.5 2.693 ;
      RECT 41.49 2.21 41.495 2.75 ;
      RECT 41.485 2.21 41.49 2.758 ;
      RECT 41.47 2.21 41.485 2.865 ;
      RECT 41.46 2.21 41.47 3 ;
      RECT 41.45 2.21 41.46 3.11 ;
      RECT 41.44 2.21 41.45 3.167 ;
      RECT 41.435 2.21 41.44 3.207 ;
      RECT 41.43 2.21 41.435 3.243 ;
      RECT 41.42 2.21 41.43 3.283 ;
      RECT 41.415 2.21 41.42 3.325 ;
      RECT 41.395 2.21 41.415 3.39 ;
      RECT 41.4 3.535 41.405 3.715 ;
      RECT 41.395 3.517 41.4 3.723 ;
      RECT 41.39 2.21 41.395 3.453 ;
      RECT 41.39 3.497 41.395 3.73 ;
      RECT 41.385 2.21 41.39 3.74 ;
      RECT 41.33 2.21 41.34 2.51 ;
      RECT 41.335 2.757 41.34 3.745 ;
      RECT 41.33 2.822 41.335 3.745 ;
      RECT 41.325 2.211 41.33 2.5 ;
      RECT 41.32 2.887 41.33 3.745 ;
      RECT 41.315 2.212 41.325 2.49 ;
      RECT 41.305 3 41.32 3.745 ;
      RECT 41.31 2.213 41.315 2.48 ;
      RECT 41.29 2.214 41.31 2.458 ;
      RECT 41.295 3.097 41.305 3.745 ;
      RECT 41.29 3.172 41.295 3.745 ;
      RECT 41.28 2.213 41.29 2.435 ;
      RECT 41.285 3.215 41.29 3.745 ;
      RECT 41.28 3.242 41.285 3.745 ;
      RECT 41.27 2.211 41.28 2.423 ;
      RECT 41.275 3.285 41.28 3.745 ;
      RECT 41.27 3.312 41.275 3.745 ;
      RECT 41.26 2.21 41.27 2.41 ;
      RECT 41.265 3.327 41.27 3.745 ;
      RECT 41.225 3.385 41.265 3.745 ;
      RECT 41.255 2.209 41.26 2.395 ;
      RECT 41.25 2.207 41.255 2.388 ;
      RECT 41.24 2.204 41.25 2.378 ;
      RECT 41.235 2.201 41.24 2.363 ;
      RECT 41.22 2.197 41.235 2.356 ;
      RECT 41.215 3.44 41.225 3.745 ;
      RECT 41.215 2.194 41.22 2.351 ;
      RECT 41.2 2.19 41.215 2.345 ;
      RECT 41.21 3.457 41.215 3.745 ;
      RECT 41.2 3.52 41.21 3.745 ;
      RECT 41.12 2.175 41.2 2.325 ;
      RECT 41.195 3.527 41.2 3.74 ;
      RECT 41.19 3.535 41.195 3.73 ;
      RECT 41.11 2.161 41.12 2.309 ;
      RECT 41.095 2.157 41.11 2.307 ;
      RECT 41.085 2.152 41.095 2.303 ;
      RECT 41.06 2.145 41.085 2.295 ;
      RECT 41.055 2.14 41.06 2.29 ;
      RECT 41.045 2.14 41.055 2.288 ;
      RECT 41.035 2.138 41.045 2.286 ;
      RECT 41.005 2.13 41.035 2.28 ;
      RECT 40.99 2.122 41.005 2.273 ;
      RECT 40.97 2.117 40.99 2.266 ;
      RECT 40.965 2.113 40.97 2.261 ;
      RECT 40.935 2.106 40.965 2.255 ;
      RECT 40.91 2.097 40.935 2.245 ;
      RECT 40.88 2.09 40.91 2.237 ;
      RECT 40.855 2.08 40.88 2.228 ;
      RECT 40.84 2.072 40.855 2.222 ;
      RECT 40.815 2.067 40.84 2.217 ;
      RECT 40.805 2.063 40.815 2.212 ;
      RECT 40.785 2.058 40.805 2.207 ;
      RECT 40.75 2.053 40.785 2.2 ;
      RECT 40.69 2.048 40.75 2.193 ;
      RECT 40.677 2.044 40.69 2.191 ;
      RECT 40.591 2.039 40.677 2.188 ;
      RECT 40.505 2.029 40.591 2.184 ;
      RECT 40.464 2.022 40.505 2.181 ;
      RECT 40.378 2.015 40.464 2.178 ;
      RECT 40.292 2.005 40.378 2.174 ;
      RECT 40.206 1.995 40.292 2.169 ;
      RECT 40.12 1.985 40.206 2.165 ;
      RECT 40.11 1.97 40.12 2.163 ;
      RECT 40.1 1.955 40.11 2.163 ;
      RECT 40.035 1.95 40.1 2.162 ;
      RECT 39.87 1.947 39.915 2.155 ;
      RECT 41.115 2.852 41.12 3.043 ;
      RECT 41.11 2.847 41.115 3.05 ;
      RECT 41.096 2.845 41.11 3.056 ;
      RECT 41.01 2.845 41.096 3.058 ;
      RECT 41.006 2.845 41.01 3.061 ;
      RECT 40.92 2.845 41.006 3.079 ;
      RECT 40.91 2.85 40.92 3.098 ;
      RECT 40.9 2.905 40.91 3.102 ;
      RECT 40.875 2.92 40.9 3.109 ;
      RECT 40.835 2.94 40.875 3.122 ;
      RECT 40.83 2.952 40.835 3.132 ;
      RECT 40.815 2.958 40.83 3.137 ;
      RECT 40.81 2.963 40.815 3.141 ;
      RECT 40.79 2.97 40.81 3.146 ;
      RECT 40.72 2.995 40.79 3.163 ;
      RECT 40.68 3.023 40.72 3.183 ;
      RECT 40.675 3.033 40.68 3.191 ;
      RECT 40.655 3.04 40.675 3.193 ;
      RECT 40.65 3.047 40.655 3.196 ;
      RECT 40.62 3.055 40.65 3.199 ;
      RECT 40.615 3.06 40.62 3.203 ;
      RECT 40.541 3.064 40.615 3.211 ;
      RECT 40.455 3.073 40.541 3.227 ;
      RECT 40.451 3.078 40.455 3.236 ;
      RECT 40.365 3.083 40.451 3.246 ;
      RECT 40.325 3.091 40.365 3.258 ;
      RECT 40.275 3.097 40.325 3.265 ;
      RECT 40.19 3.106 40.275 3.28 ;
      RECT 40.115 3.117 40.19 3.298 ;
      RECT 40.08 3.124 40.115 3.308 ;
      RECT 40.005 3.132 40.08 3.313 ;
      RECT 39.95 3.141 40.005 3.313 ;
      RECT 39.925 3.146 39.95 3.311 ;
      RECT 39.915 3.149 39.925 3.309 ;
      RECT 39.88 3.151 39.915 3.307 ;
      RECT 39.85 3.153 39.88 3.303 ;
      RECT 39.805 3.152 39.85 3.299 ;
      RECT 39.785 3.147 39.805 3.296 ;
      RECT 39.735 3.132 39.785 3.293 ;
      RECT 39.725 3.117 39.735 3.288 ;
      RECT 39.675 3.102 39.725 3.278 ;
      RECT 39.625 3.077 39.675 3.258 ;
      RECT 39.615 3.062 39.625 3.24 ;
      RECT 39.61 3.06 39.615 3.234 ;
      RECT 39.59 3.055 39.61 3.229 ;
      RECT 39.585 3.047 39.59 3.223 ;
      RECT 39.57 3.041 39.585 3.216 ;
      RECT 39.565 3.036 39.57 3.208 ;
      RECT 39.545 3.031 39.565 3.2 ;
      RECT 39.53 3.024 39.545 3.193 ;
      RECT 39.515 3.018 39.53 3.184 ;
      RECT 39.51 3.012 39.515 3.177 ;
      RECT 39.465 2.987 39.51 3.163 ;
      RECT 39.45 2.957 39.465 3.145 ;
      RECT 39.435 2.94 39.45 3.136 ;
      RECT 39.41 2.92 39.435 3.124 ;
      RECT 39.37 2.89 39.41 3.104 ;
      RECT 39.36 2.86 39.37 3.089 ;
      RECT 39.345 2.85 39.36 3.082 ;
      RECT 39.29 2.815 39.345 3.061 ;
      RECT 39.275 2.778 39.29 3.04 ;
      RECT 39.265 2.765 39.275 3.032 ;
      RECT 39.215 2.735 39.265 3.014 ;
      RECT 39.2 2.665 39.215 2.995 ;
      RECT 39.155 2.665 39.2 2.978 ;
      RECT 39.13 2.665 39.155 2.96 ;
      RECT 39.12 2.665 39.13 2.953 ;
      RECT 39.041 2.665 39.12 2.946 ;
      RECT 38.955 2.665 39.041 2.938 ;
      RECT 38.94 2.697 38.955 2.933 ;
      RECT 38.865 2.707 38.94 2.929 ;
      RECT 38.845 2.717 38.865 2.924 ;
      RECT 38.82 2.717 38.845 2.921 ;
      RECT 38.81 2.707 38.82 2.92 ;
      RECT 38.8 2.68 38.81 2.919 ;
      RECT 38.76 2.675 38.8 2.917 ;
      RECT 38.715 2.675 38.76 2.913 ;
      RECT 38.69 2.675 38.715 2.908 ;
      RECT 38.64 2.675 38.69 2.895 ;
      RECT 38.6 2.68 38.61 2.88 ;
      RECT 38.61 2.675 38.64 2.885 ;
      RECT 40.595 2.455 40.855 2.715 ;
      RECT 40.59 2.477 40.855 2.673 ;
      RECT 39.83 2.305 40.05 2.67 ;
      RECT 39.812 2.392 40.05 2.669 ;
      RECT 39.795 2.397 40.05 2.666 ;
      RECT 39.795 2.397 40.07 2.665 ;
      RECT 39.765 2.407 40.07 2.663 ;
      RECT 39.76 2.422 40.07 2.659 ;
      RECT 39.76 2.422 40.075 2.658 ;
      RECT 39.755 2.48 40.075 2.656 ;
      RECT 39.755 2.48 40.085 2.653 ;
      RECT 39.75 2.545 40.085 2.648 ;
      RECT 39.83 2.305 40.09 2.565 ;
      RECT 38.575 2.135 38.835 2.395 ;
      RECT 38.575 2.178 38.921 2.369 ;
      RECT 38.575 2.178 38.965 2.368 ;
      RECT 38.575 2.178 38.985 2.366 ;
      RECT 38.575 2.178 39.085 2.365 ;
      RECT 38.575 2.178 39.105 2.363 ;
      RECT 38.575 2.178 39.115 2.358 ;
      RECT 38.985 2.145 39.175 2.355 ;
      RECT 38.985 2.147 39.18 2.353 ;
      RECT 38.975 2.152 39.185 2.345 ;
      RECT 38.921 2.176 39.185 2.345 ;
      RECT 38.965 2.17 38.975 2.367 ;
      RECT 38.975 2.15 39.18 2.353 ;
      RECT 37.93 3.21 38.135 3.44 ;
      RECT 37.87 3.16 37.925 3.42 ;
      RECT 37.93 3.16 38.13 3.44 ;
      RECT 38.9 3.475 38.905 3.502 ;
      RECT 38.89 3.385 38.9 3.507 ;
      RECT 38.885 3.307 38.89 3.513 ;
      RECT 38.875 3.297 38.885 3.52 ;
      RECT 38.87 3.287 38.875 3.526 ;
      RECT 38.86 3.282 38.87 3.528 ;
      RECT 38.845 3.274 38.86 3.536 ;
      RECT 38.83 3.265 38.845 3.548 ;
      RECT 38.82 3.257 38.83 3.558 ;
      RECT 38.785 3.175 38.82 3.576 ;
      RECT 38.75 3.175 38.785 3.595 ;
      RECT 38.735 3.175 38.75 3.603 ;
      RECT 38.68 3.175 38.735 3.603 ;
      RECT 38.646 3.175 38.68 3.594 ;
      RECT 38.56 3.175 38.646 3.57 ;
      RECT 38.55 3.235 38.56 3.552 ;
      RECT 38.51 3.237 38.55 3.543 ;
      RECT 38.505 3.239 38.51 3.533 ;
      RECT 38.485 3.241 38.505 3.528 ;
      RECT 38.475 3.244 38.485 3.523 ;
      RECT 38.465 3.245 38.475 3.518 ;
      RECT 38.441 3.246 38.465 3.51 ;
      RECT 38.355 3.251 38.441 3.488 ;
      RECT 38.3 3.25 38.355 3.461 ;
      RECT 38.285 3.243 38.3 3.448 ;
      RECT 38.25 3.238 38.285 3.444 ;
      RECT 38.195 3.23 38.25 3.443 ;
      RECT 38.135 3.217 38.195 3.441 ;
      RECT 37.925 3.16 37.93 3.428 ;
      RECT 38 2.53 38.185 2.74 ;
      RECT 37.99 2.535 38.2 2.733 ;
      RECT 38.03 2.44 38.29 2.7 ;
      RECT 37.985 2.597 38.29 2.623 ;
      RECT 37.33 2.39 37.335 3.19 ;
      RECT 37.275 2.44 37.305 3.19 ;
      RECT 37.265 2.44 37.27 2.75 ;
      RECT 37.25 2.44 37.255 2.745 ;
      RECT 36.795 2.485 36.81 2.7 ;
      RECT 36.725 2.485 36.81 2.695 ;
      RECT 37.99 2.065 38.06 2.275 ;
      RECT 38.06 2.072 38.07 2.27 ;
      RECT 37.956 2.065 37.99 2.282 ;
      RECT 37.87 2.065 37.956 2.306 ;
      RECT 37.86 2.07 37.87 2.325 ;
      RECT 37.855 2.082 37.86 2.328 ;
      RECT 37.84 2.097 37.855 2.332 ;
      RECT 37.835 2.115 37.84 2.336 ;
      RECT 37.795 2.125 37.835 2.345 ;
      RECT 37.78 2.132 37.795 2.357 ;
      RECT 37.765 2.137 37.78 2.362 ;
      RECT 37.75 2.14 37.765 2.367 ;
      RECT 37.74 2.142 37.75 2.371 ;
      RECT 37.705 2.149 37.74 2.379 ;
      RECT 37.67 2.157 37.705 2.393 ;
      RECT 37.66 2.163 37.67 2.402 ;
      RECT 37.655 2.165 37.66 2.404 ;
      RECT 37.635 2.168 37.655 2.41 ;
      RECT 37.605 2.175 37.635 2.421 ;
      RECT 37.595 2.181 37.605 2.428 ;
      RECT 37.57 2.184 37.595 2.435 ;
      RECT 37.56 2.188 37.57 2.443 ;
      RECT 37.555 2.189 37.56 2.465 ;
      RECT 37.55 2.19 37.555 2.48 ;
      RECT 37.545 2.191 37.55 2.495 ;
      RECT 37.54 2.192 37.545 2.51 ;
      RECT 37.535 2.193 37.54 2.54 ;
      RECT 37.525 2.195 37.535 2.573 ;
      RECT 37.51 2.199 37.525 2.62 ;
      RECT 37.5 2.202 37.51 2.665 ;
      RECT 37.495 2.205 37.5 2.693 ;
      RECT 37.485 2.207 37.495 2.72 ;
      RECT 37.48 2.21 37.485 2.755 ;
      RECT 37.45 2.215 37.48 2.813 ;
      RECT 37.445 2.22 37.45 2.898 ;
      RECT 37.44 2.222 37.445 2.933 ;
      RECT 37.435 2.224 37.44 3.015 ;
      RECT 37.43 2.226 37.435 3.103 ;
      RECT 37.42 2.228 37.43 3.185 ;
      RECT 37.405 2.242 37.42 3.19 ;
      RECT 37.37 2.287 37.405 3.19 ;
      RECT 37.36 2.327 37.37 3.19 ;
      RECT 37.345 2.355 37.36 3.19 ;
      RECT 37.34 2.372 37.345 3.19 ;
      RECT 37.335 2.38 37.34 3.19 ;
      RECT 37.325 2.395 37.33 3.19 ;
      RECT 37.32 2.402 37.325 3.19 ;
      RECT 37.31 2.422 37.32 3.19 ;
      RECT 37.305 2.435 37.31 3.19 ;
      RECT 37.27 2.44 37.275 2.775 ;
      RECT 37.255 2.83 37.275 3.19 ;
      RECT 37.255 2.44 37.265 2.748 ;
      RECT 37.25 2.87 37.255 3.19 ;
      RECT 37.2 2.44 37.25 2.743 ;
      RECT 37.245 2.907 37.25 3.19 ;
      RECT 37.235 2.93 37.245 3.19 ;
      RECT 37.23 2.975 37.235 3.19 ;
      RECT 37.22 2.985 37.23 3.183 ;
      RECT 37.146 2.44 37.2 2.737 ;
      RECT 37.06 2.44 37.146 2.73 ;
      RECT 37.011 2.487 37.06 2.723 ;
      RECT 36.925 2.495 37.011 2.716 ;
      RECT 36.91 2.492 36.925 2.711 ;
      RECT 36.896 2.485 36.91 2.71 ;
      RECT 36.81 2.485 36.896 2.705 ;
      RECT 36.715 2.49 36.725 2.69 ;
      RECT 36.305 1.92 36.32 2.32 ;
      RECT 36.5 1.92 36.505 2.18 ;
      RECT 36.245 1.92 36.29 2.18 ;
      RECT 36.7 3.225 36.705 3.43 ;
      RECT 36.695 3.215 36.7 3.435 ;
      RECT 36.69 3.202 36.695 3.44 ;
      RECT 36.685 3.182 36.69 3.44 ;
      RECT 36.66 3.135 36.685 3.44 ;
      RECT 36.625 3.05 36.66 3.44 ;
      RECT 36.62 2.987 36.625 3.44 ;
      RECT 36.615 2.972 36.62 3.44 ;
      RECT 36.6 2.932 36.615 3.44 ;
      RECT 36.595 2.907 36.6 3.44 ;
      RECT 36.585 2.89 36.595 3.44 ;
      RECT 36.55 2.812 36.585 3.44 ;
      RECT 36.545 2.755 36.55 3.44 ;
      RECT 36.54 2.742 36.545 3.44 ;
      RECT 36.53 2.72 36.54 3.44 ;
      RECT 36.52 2.685 36.53 3.44 ;
      RECT 36.51 2.655 36.52 3.44 ;
      RECT 36.5 2.57 36.51 3.083 ;
      RECT 36.507 3.215 36.51 3.44 ;
      RECT 36.505 3.225 36.507 3.44 ;
      RECT 36.495 3.235 36.505 3.435 ;
      RECT 36.49 1.92 36.5 2.315 ;
      RECT 36.495 2.447 36.5 3.058 ;
      RECT 36.49 2.345 36.495 3.041 ;
      RECT 36.48 1.92 36.49 3.017 ;
      RECT 36.475 1.92 36.48 2.988 ;
      RECT 36.47 1.92 36.475 2.978 ;
      RECT 36.45 1.92 36.47 2.94 ;
      RECT 36.445 1.92 36.45 2.898 ;
      RECT 36.44 1.92 36.445 2.878 ;
      RECT 36.41 1.92 36.44 2.828 ;
      RECT 36.4 1.92 36.41 2.775 ;
      RECT 36.395 1.92 36.4 2.748 ;
      RECT 36.39 1.92 36.395 2.733 ;
      RECT 36.38 1.92 36.39 2.71 ;
      RECT 36.37 1.92 36.38 2.685 ;
      RECT 36.365 1.92 36.37 2.625 ;
      RECT 36.355 1.92 36.365 2.563 ;
      RECT 36.35 1.92 36.355 2.483 ;
      RECT 36.345 1.92 36.35 2.448 ;
      RECT 36.34 1.92 36.345 2.423 ;
      RECT 36.335 1.92 36.34 2.408 ;
      RECT 36.33 1.92 36.335 2.378 ;
      RECT 36.325 1.92 36.33 2.355 ;
      RECT 36.32 1.92 36.325 2.328 ;
      RECT 36.29 1.92 36.305 2.315 ;
      RECT 35.445 3.455 35.63 3.665 ;
      RECT 35.435 3.46 35.645 3.658 ;
      RECT 35.435 3.46 35.665 3.63 ;
      RECT 35.435 3.46 35.68 3.609 ;
      RECT 35.435 3.46 35.695 3.607 ;
      RECT 35.435 3.46 35.705 3.606 ;
      RECT 35.435 3.46 35.735 3.603 ;
      RECT 36.085 3.305 36.345 3.565 ;
      RECT 36.045 3.352 36.345 3.548 ;
      RECT 36.036 3.36 36.045 3.551 ;
      RECT 35.63 3.453 36.345 3.548 ;
      RECT 35.95 3.378 36.036 3.558 ;
      RECT 35.645 3.45 36.345 3.548 ;
      RECT 35.891 3.4 35.95 3.57 ;
      RECT 35.665 3.446 36.345 3.548 ;
      RECT 35.805 3.412 35.891 3.581 ;
      RECT 35.68 3.442 36.345 3.548 ;
      RECT 35.75 3.425 35.805 3.593 ;
      RECT 35.695 3.44 36.345 3.548 ;
      RECT 35.735 3.431 35.75 3.599 ;
      RECT 35.705 3.436 36.345 3.548 ;
      RECT 35.85 2.96 36.11 3.22 ;
      RECT 35.85 2.98 36.22 3.19 ;
      RECT 35.85 2.985 36.23 3.185 ;
      RECT 36.041 2.399 36.12 2.63 ;
      RECT 35.955 2.402 36.17 2.625 ;
      RECT 35.95 2.402 36.17 2.62 ;
      RECT 35.95 2.407 36.18 2.618 ;
      RECT 35.925 2.407 36.18 2.615 ;
      RECT 35.925 2.415 36.19 2.613 ;
      RECT 35.805 2.35 36.065 2.61 ;
      RECT 35.805 2.397 36.115 2.61 ;
      RECT 35.06 2.97 35.065 3.23 ;
      RECT 34.89 2.74 34.895 3.23 ;
      RECT 34.775 2.98 34.78 3.205 ;
      RECT 35.485 2.075 35.49 2.285 ;
      RECT 35.49 2.08 35.505 2.28 ;
      RECT 35.425 2.075 35.485 2.293 ;
      RECT 35.41 2.075 35.425 2.303 ;
      RECT 35.36 2.075 35.41 2.32 ;
      RECT 35.34 2.075 35.36 2.343 ;
      RECT 35.325 2.075 35.34 2.355 ;
      RECT 35.305 2.075 35.325 2.365 ;
      RECT 35.295 2.08 35.305 2.374 ;
      RECT 35.29 2.09 35.295 2.379 ;
      RECT 35.285 2.102 35.29 2.383 ;
      RECT 35.275 2.125 35.285 2.388 ;
      RECT 35.27 2.14 35.275 2.392 ;
      RECT 35.265 2.157 35.27 2.395 ;
      RECT 35.26 2.165 35.265 2.398 ;
      RECT 35.25 2.17 35.26 2.402 ;
      RECT 35.245 2.177 35.25 2.407 ;
      RECT 35.235 2.182 35.245 2.411 ;
      RECT 35.21 2.194 35.235 2.422 ;
      RECT 35.19 2.211 35.21 2.438 ;
      RECT 35.165 2.228 35.19 2.46 ;
      RECT 35.13 2.251 35.165 2.518 ;
      RECT 35.11 2.273 35.13 2.58 ;
      RECT 35.105 2.283 35.11 2.615 ;
      RECT 35.095 2.29 35.105 2.653 ;
      RECT 35.09 2.297 35.095 2.673 ;
      RECT 35.085 2.308 35.09 2.71 ;
      RECT 35.08 2.316 35.085 2.775 ;
      RECT 35.07 2.327 35.08 2.828 ;
      RECT 35.065 2.345 35.07 2.898 ;
      RECT 35.06 2.355 35.065 2.935 ;
      RECT 35.055 2.365 35.06 3.23 ;
      RECT 35.05 2.377 35.055 3.23 ;
      RECT 35.045 2.387 35.05 3.23 ;
      RECT 35.035 2.397 35.045 3.23 ;
      RECT 35.025 2.42 35.035 3.23 ;
      RECT 35.01 2.455 35.025 3.23 ;
      RECT 34.97 2.517 35.01 3.23 ;
      RECT 34.965 2.57 34.97 3.23 ;
      RECT 34.94 2.605 34.965 3.23 ;
      RECT 34.925 2.65 34.94 3.23 ;
      RECT 34.92 2.672 34.925 3.23 ;
      RECT 34.91 2.685 34.92 3.23 ;
      RECT 34.9 2.71 34.91 3.23 ;
      RECT 34.895 2.732 34.9 3.23 ;
      RECT 34.87 2.77 34.89 3.23 ;
      RECT 34.83 2.827 34.87 3.23 ;
      RECT 34.825 2.877 34.83 3.23 ;
      RECT 34.82 2.895 34.825 3.23 ;
      RECT 34.815 2.907 34.82 3.23 ;
      RECT 34.805 2.925 34.815 3.23 ;
      RECT 34.795 2.945 34.805 3.205 ;
      RECT 34.79 2.962 34.795 3.205 ;
      RECT 34.78 2.975 34.79 3.205 ;
      RECT 34.75 2.985 34.775 3.205 ;
      RECT 34.74 2.992 34.75 3.205 ;
      RECT 34.725 3.002 34.74 3.2 ;
      RECT 33.825 7.77 34.115 8 ;
      RECT 33.885 6.29 34.055 8 ;
      RECT 33.875 6.66 34.23 7.015 ;
      RECT 33.825 6.29 34.115 6.52 ;
      RECT 33.42 2.395 33.525 2.965 ;
      RECT 33.42 2.73 33.745 2.96 ;
      RECT 33.42 2.76 33.915 2.93 ;
      RECT 33.42 2.395 33.61 2.96 ;
      RECT 32.835 2.36 33.125 2.59 ;
      RECT 32.835 2.395 33.61 2.565 ;
      RECT 32.895 0.88 33.065 2.59 ;
      RECT 32.835 0.88 33.125 1.11 ;
      RECT 32.835 7.77 33.125 8 ;
      RECT 32.895 6.29 33.065 8 ;
      RECT 32.835 6.29 33.125 6.52 ;
      RECT 32.835 6.325 33.69 6.485 ;
      RECT 33.52 5.92 33.69 6.485 ;
      RECT 32.835 6.32 33.23 6.485 ;
      RECT 33.455 5.92 33.745 6.15 ;
      RECT 33.455 5.95 33.915 6.12 ;
      RECT 32.465 2.73 32.755 2.96 ;
      RECT 32.465 2.76 32.925 2.93 ;
      RECT 32.53 1.655 32.695 2.96 ;
      RECT 31.045 1.625 31.335 1.855 ;
      RECT 31.045 1.655 32.695 1.825 ;
      RECT 31.105 0.885 31.275 1.855 ;
      RECT 31.045 0.885 31.335 1.115 ;
      RECT 31.045 7.765 31.335 7.995 ;
      RECT 31.105 7.025 31.275 7.995 ;
      RECT 31.105 7.12 32.695 7.29 ;
      RECT 32.525 5.92 32.695 7.29 ;
      RECT 31.045 7.025 31.335 7.255 ;
      RECT 32.465 5.92 32.755 6.15 ;
      RECT 32.465 5.95 32.925 6.12 ;
      RECT 31.475 1.965 31.825 2.315 ;
      RECT 29.14 2.025 31.825 2.195 ;
      RECT 29.14 1.34 29.31 2.195 ;
      RECT 29.04 1.34 29.39 1.69 ;
      RECT 31.5 6.655 31.825 6.98 ;
      RECT 26.925 6.61 27.275 6.96 ;
      RECT 31.475 6.655 31.825 6.885 ;
      RECT 26.695 6.655 27.275 6.885 ;
      RECT 26.525 6.685 31.825 6.855 ;
      RECT 30.7 2.365 31.02 2.685 ;
      RECT 30.67 2.365 31.02 2.595 ;
      RECT 30.5 2.395 31.02 2.565 ;
      RECT 30.7 6.255 31.02 6.545 ;
      RECT 30.67 6.285 31.02 6.515 ;
      RECT 30.5 6.315 31.02 6.485 ;
      RECT 27.335 2.465 27.52 2.675 ;
      RECT 27.325 2.47 27.535 2.668 ;
      RECT 27.325 2.47 27.621 2.645 ;
      RECT 27.325 2.47 27.68 2.62 ;
      RECT 27.325 2.47 27.735 2.6 ;
      RECT 27.325 2.47 27.745 2.588 ;
      RECT 27.325 2.47 27.94 2.527 ;
      RECT 27.325 2.47 27.97 2.51 ;
      RECT 27.325 2.47 27.99 2.5 ;
      RECT 27.87 2.235 28.13 2.495 ;
      RECT 27.855 2.325 27.87 2.542 ;
      RECT 27.39 2.457 28.13 2.495 ;
      RECT 27.841 2.336 27.855 2.548 ;
      RECT 27.43 2.45 28.13 2.495 ;
      RECT 27.755 2.376 27.841 2.567 ;
      RECT 27.68 2.437 28.13 2.495 ;
      RECT 27.75 2.412 27.755 2.584 ;
      RECT 27.735 2.422 28.13 2.495 ;
      RECT 27.745 2.417 27.75 2.586 ;
      RECT 28.04 2.922 28.045 3.014 ;
      RECT 28.035 2.9 28.04 3.031 ;
      RECT 28.03 2.89 28.035 3.043 ;
      RECT 28.02 2.881 28.03 3.053 ;
      RECT 28.015 2.876 28.02 3.061 ;
      RECT 28.01 2.735 28.015 3.064 ;
      RECT 27.976 2.735 28.01 3.075 ;
      RECT 27.89 2.735 27.976 3.11 ;
      RECT 27.81 2.735 27.89 3.158 ;
      RECT 27.781 2.735 27.81 3.182 ;
      RECT 27.695 2.735 27.781 3.188 ;
      RECT 27.69 2.919 27.695 3.193 ;
      RECT 27.655 2.93 27.69 3.196 ;
      RECT 27.63 2.945 27.655 3.2 ;
      RECT 27.616 2.954 27.63 3.202 ;
      RECT 27.53 2.981 27.616 3.208 ;
      RECT 27.465 3.022 27.53 3.217 ;
      RECT 27.45 3.042 27.465 3.222 ;
      RECT 27.42 3.052 27.45 3.225 ;
      RECT 27.415 3.062 27.42 3.228 ;
      RECT 27.385 3.067 27.415 3.23 ;
      RECT 27.365 3.072 27.385 3.234 ;
      RECT 27.28 3.075 27.365 3.241 ;
      RECT 27.265 3.072 27.28 3.247 ;
      RECT 27.255 3.069 27.265 3.249 ;
      RECT 27.235 3.066 27.255 3.251 ;
      RECT 27.215 3.062 27.235 3.252 ;
      RECT 27.2 3.058 27.215 3.254 ;
      RECT 27.19 3.055 27.2 3.255 ;
      RECT 27.15 3.049 27.19 3.253 ;
      RECT 27.14 3.044 27.15 3.251 ;
      RECT 27.125 3.041 27.14 3.247 ;
      RECT 27.1 3.036 27.125 3.24 ;
      RECT 27.05 3.027 27.1 3.228 ;
      RECT 26.98 3.013 27.05 3.21 ;
      RECT 26.922 2.998 26.98 3.192 ;
      RECT 26.836 2.981 26.922 3.172 ;
      RECT 26.75 2.96 26.836 3.147 ;
      RECT 26.7 2.945 26.75 3.128 ;
      RECT 26.696 2.939 26.7 3.12 ;
      RECT 26.61 2.929 26.696 3.107 ;
      RECT 26.575 2.914 26.61 3.09 ;
      RECT 26.56 2.907 26.575 3.083 ;
      RECT 26.5 2.895 26.56 3.071 ;
      RECT 26.48 2.882 26.5 3.059 ;
      RECT 26.44 2.873 26.48 3.051 ;
      RECT 26.435 2.865 26.44 3.044 ;
      RECT 26.355 2.855 26.435 3.03 ;
      RECT 26.34 2.842 26.355 3.015 ;
      RECT 26.335 2.84 26.34 3.013 ;
      RECT 26.256 2.828 26.335 3 ;
      RECT 26.17 2.803 26.256 2.975 ;
      RECT 26.155 2.772 26.17 2.96 ;
      RECT 26.14 2.747 26.155 2.956 ;
      RECT 26.125 2.74 26.14 2.952 ;
      RECT 25.95 2.745 25.955 2.948 ;
      RECT 25.945 2.75 25.95 2.943 ;
      RECT 25.955 2.74 26.125 2.95 ;
      RECT 26.67 2.5 26.775 2.76 ;
      RECT 27.485 2.025 27.49 2.25 ;
      RECT 27.615 2.025 27.67 2.235 ;
      RECT 27.67 2.03 27.68 2.228 ;
      RECT 27.576 2.025 27.615 2.238 ;
      RECT 27.49 2.025 27.576 2.245 ;
      RECT 27.47 2.03 27.485 2.251 ;
      RECT 27.46 2.07 27.47 2.253 ;
      RECT 27.43 2.08 27.46 2.255 ;
      RECT 27.425 2.085 27.43 2.257 ;
      RECT 27.4 2.09 27.425 2.259 ;
      RECT 27.385 2.095 27.4 2.261 ;
      RECT 27.37 2.097 27.385 2.263 ;
      RECT 27.365 2.102 27.37 2.265 ;
      RECT 27.315 2.11 27.365 2.268 ;
      RECT 27.29 2.119 27.315 2.273 ;
      RECT 27.28 2.126 27.29 2.278 ;
      RECT 27.275 2.129 27.28 2.282 ;
      RECT 27.255 2.132 27.275 2.291 ;
      RECT 27.225 2.14 27.255 2.311 ;
      RECT 27.196 2.153 27.225 2.333 ;
      RECT 27.11 2.187 27.196 2.377 ;
      RECT 27.105 2.213 27.11 2.415 ;
      RECT 27.1 2.217 27.105 2.424 ;
      RECT 27.065 2.23 27.1 2.457 ;
      RECT 27.055 2.244 27.065 2.495 ;
      RECT 27.05 2.248 27.055 2.508 ;
      RECT 27.045 2.252 27.05 2.513 ;
      RECT 27.035 2.26 27.045 2.525 ;
      RECT 27.03 2.267 27.035 2.54 ;
      RECT 27.005 2.28 27.03 2.565 ;
      RECT 26.965 2.309 27.005 2.62 ;
      RECT 26.95 2.334 26.965 2.675 ;
      RECT 26.94 2.345 26.95 2.698 ;
      RECT 26.935 2.352 26.94 2.71 ;
      RECT 26.93 2.356 26.935 2.718 ;
      RECT 26.875 2.384 26.93 2.76 ;
      RECT 26.855 2.42 26.875 2.76 ;
      RECT 26.84 2.435 26.855 2.76 ;
      RECT 26.785 2.467 26.84 2.76 ;
      RECT 26.775 2.497 26.785 2.76 ;
      RECT 26.385 2.112 26.57 2.35 ;
      RECT 26.37 2.114 26.58 2.345 ;
      RECT 26.255 2.06 26.515 2.32 ;
      RECT 26.25 2.097 26.515 2.274 ;
      RECT 26.245 2.107 26.515 2.271 ;
      RECT 26.24 2.147 26.58 2.265 ;
      RECT 26.235 2.18 26.58 2.255 ;
      RECT 26.245 2.122 26.595 2.193 ;
      RECT 26.542 3.22 26.555 3.75 ;
      RECT 26.456 3.22 26.555 3.749 ;
      RECT 26.456 3.22 26.56 3.748 ;
      RECT 26.37 3.22 26.56 3.746 ;
      RECT 26.365 3.22 26.56 3.743 ;
      RECT 26.365 3.22 26.57 3.741 ;
      RECT 26.36 3.512 26.57 3.738 ;
      RECT 26.36 3.522 26.575 3.735 ;
      RECT 26.36 3.59 26.58 3.731 ;
      RECT 26.35 3.595 26.58 3.73 ;
      RECT 26.35 3.687 26.585 3.727 ;
      RECT 26.335 3.22 26.595 3.48 ;
      RECT 26.265 7.765 26.555 7.995 ;
      RECT 26.325 7.025 26.495 7.995 ;
      RECT 26.24 7.055 26.58 7.4 ;
      RECT 26.265 7.025 26.555 7.4 ;
      RECT 25.565 2.21 25.61 3.745 ;
      RECT 25.765 2.21 25.795 2.425 ;
      RECT 24.14 1.95 24.26 2.16 ;
      RECT 23.8 1.9 24.06 2.16 ;
      RECT 23.8 1.945 24.095 2.15 ;
      RECT 25.805 2.226 25.81 2.28 ;
      RECT 25.8 2.219 25.805 2.413 ;
      RECT 25.795 2.213 25.8 2.42 ;
      RECT 25.75 2.21 25.765 2.433 ;
      RECT 25.745 2.21 25.75 2.455 ;
      RECT 25.74 2.21 25.745 2.503 ;
      RECT 25.735 2.21 25.74 2.523 ;
      RECT 25.725 2.21 25.735 2.63 ;
      RECT 25.72 2.21 25.725 2.693 ;
      RECT 25.715 2.21 25.72 2.75 ;
      RECT 25.71 2.21 25.715 2.758 ;
      RECT 25.695 2.21 25.71 2.865 ;
      RECT 25.685 2.21 25.695 3 ;
      RECT 25.675 2.21 25.685 3.11 ;
      RECT 25.665 2.21 25.675 3.167 ;
      RECT 25.66 2.21 25.665 3.207 ;
      RECT 25.655 2.21 25.66 3.243 ;
      RECT 25.645 2.21 25.655 3.283 ;
      RECT 25.64 2.21 25.645 3.325 ;
      RECT 25.62 2.21 25.64 3.39 ;
      RECT 25.625 3.535 25.63 3.715 ;
      RECT 25.62 3.517 25.625 3.723 ;
      RECT 25.615 2.21 25.62 3.453 ;
      RECT 25.615 3.497 25.62 3.73 ;
      RECT 25.61 2.21 25.615 3.74 ;
      RECT 25.555 2.21 25.565 2.51 ;
      RECT 25.56 2.757 25.565 3.745 ;
      RECT 25.555 2.822 25.56 3.745 ;
      RECT 25.55 2.211 25.555 2.5 ;
      RECT 25.545 2.887 25.555 3.745 ;
      RECT 25.54 2.212 25.55 2.49 ;
      RECT 25.53 3 25.545 3.745 ;
      RECT 25.535 2.213 25.54 2.48 ;
      RECT 25.515 2.214 25.535 2.458 ;
      RECT 25.52 3.097 25.53 3.745 ;
      RECT 25.515 3.172 25.52 3.745 ;
      RECT 25.505 2.213 25.515 2.435 ;
      RECT 25.51 3.215 25.515 3.745 ;
      RECT 25.505 3.242 25.51 3.745 ;
      RECT 25.495 2.211 25.505 2.423 ;
      RECT 25.5 3.285 25.505 3.745 ;
      RECT 25.495 3.312 25.5 3.745 ;
      RECT 25.485 2.21 25.495 2.41 ;
      RECT 25.49 3.327 25.495 3.745 ;
      RECT 25.45 3.385 25.49 3.745 ;
      RECT 25.48 2.209 25.485 2.395 ;
      RECT 25.475 2.207 25.48 2.388 ;
      RECT 25.465 2.204 25.475 2.378 ;
      RECT 25.46 2.201 25.465 2.363 ;
      RECT 25.445 2.197 25.46 2.356 ;
      RECT 25.44 3.44 25.45 3.745 ;
      RECT 25.44 2.194 25.445 2.351 ;
      RECT 25.425 2.19 25.44 2.345 ;
      RECT 25.435 3.457 25.44 3.745 ;
      RECT 25.425 3.52 25.435 3.745 ;
      RECT 25.345 2.175 25.425 2.325 ;
      RECT 25.42 3.527 25.425 3.74 ;
      RECT 25.415 3.535 25.42 3.73 ;
      RECT 25.335 2.161 25.345 2.309 ;
      RECT 25.32 2.157 25.335 2.307 ;
      RECT 25.31 2.152 25.32 2.303 ;
      RECT 25.285 2.145 25.31 2.295 ;
      RECT 25.28 2.14 25.285 2.29 ;
      RECT 25.27 2.14 25.28 2.288 ;
      RECT 25.26 2.138 25.27 2.286 ;
      RECT 25.23 2.13 25.26 2.28 ;
      RECT 25.215 2.122 25.23 2.273 ;
      RECT 25.195 2.117 25.215 2.266 ;
      RECT 25.19 2.113 25.195 2.261 ;
      RECT 25.16 2.106 25.19 2.255 ;
      RECT 25.135 2.097 25.16 2.245 ;
      RECT 25.105 2.09 25.135 2.237 ;
      RECT 25.08 2.08 25.105 2.228 ;
      RECT 25.065 2.072 25.08 2.222 ;
      RECT 25.04 2.067 25.065 2.217 ;
      RECT 25.03 2.063 25.04 2.212 ;
      RECT 25.01 2.058 25.03 2.207 ;
      RECT 24.975 2.053 25.01 2.2 ;
      RECT 24.915 2.048 24.975 2.193 ;
      RECT 24.902 2.044 24.915 2.191 ;
      RECT 24.816 2.039 24.902 2.188 ;
      RECT 24.73 2.029 24.816 2.184 ;
      RECT 24.689 2.022 24.73 2.181 ;
      RECT 24.603 2.015 24.689 2.178 ;
      RECT 24.517 2.005 24.603 2.174 ;
      RECT 24.431 1.995 24.517 2.169 ;
      RECT 24.345 1.985 24.431 2.165 ;
      RECT 24.335 1.97 24.345 2.163 ;
      RECT 24.325 1.955 24.335 2.163 ;
      RECT 24.26 1.95 24.325 2.162 ;
      RECT 24.095 1.947 24.14 2.155 ;
      RECT 25.34 2.852 25.345 3.043 ;
      RECT 25.335 2.847 25.34 3.05 ;
      RECT 25.321 2.845 25.335 3.056 ;
      RECT 25.235 2.845 25.321 3.058 ;
      RECT 25.231 2.845 25.235 3.061 ;
      RECT 25.145 2.845 25.231 3.079 ;
      RECT 25.135 2.85 25.145 3.098 ;
      RECT 25.125 2.905 25.135 3.102 ;
      RECT 25.1 2.92 25.125 3.109 ;
      RECT 25.06 2.94 25.1 3.122 ;
      RECT 25.055 2.952 25.06 3.132 ;
      RECT 25.04 2.958 25.055 3.137 ;
      RECT 25.035 2.963 25.04 3.141 ;
      RECT 25.015 2.97 25.035 3.146 ;
      RECT 24.945 2.995 25.015 3.163 ;
      RECT 24.905 3.023 24.945 3.183 ;
      RECT 24.9 3.033 24.905 3.191 ;
      RECT 24.88 3.04 24.9 3.193 ;
      RECT 24.875 3.047 24.88 3.196 ;
      RECT 24.845 3.055 24.875 3.199 ;
      RECT 24.84 3.06 24.845 3.203 ;
      RECT 24.766 3.064 24.84 3.211 ;
      RECT 24.68 3.073 24.766 3.227 ;
      RECT 24.676 3.078 24.68 3.236 ;
      RECT 24.59 3.083 24.676 3.246 ;
      RECT 24.55 3.091 24.59 3.258 ;
      RECT 24.5 3.097 24.55 3.265 ;
      RECT 24.415 3.106 24.5 3.28 ;
      RECT 24.34 3.117 24.415 3.298 ;
      RECT 24.305 3.124 24.34 3.308 ;
      RECT 24.23 3.132 24.305 3.313 ;
      RECT 24.175 3.141 24.23 3.313 ;
      RECT 24.15 3.146 24.175 3.311 ;
      RECT 24.14 3.149 24.15 3.309 ;
      RECT 24.105 3.151 24.14 3.307 ;
      RECT 24.075 3.153 24.105 3.303 ;
      RECT 24.03 3.152 24.075 3.299 ;
      RECT 24.01 3.147 24.03 3.296 ;
      RECT 23.96 3.132 24.01 3.293 ;
      RECT 23.95 3.117 23.96 3.288 ;
      RECT 23.9 3.102 23.95 3.278 ;
      RECT 23.85 3.077 23.9 3.258 ;
      RECT 23.84 3.062 23.85 3.24 ;
      RECT 23.835 3.06 23.84 3.234 ;
      RECT 23.815 3.055 23.835 3.229 ;
      RECT 23.81 3.047 23.815 3.223 ;
      RECT 23.795 3.041 23.81 3.216 ;
      RECT 23.79 3.036 23.795 3.208 ;
      RECT 23.77 3.031 23.79 3.2 ;
      RECT 23.755 3.024 23.77 3.193 ;
      RECT 23.74 3.018 23.755 3.184 ;
      RECT 23.735 3.012 23.74 3.177 ;
      RECT 23.69 2.987 23.735 3.163 ;
      RECT 23.675 2.957 23.69 3.145 ;
      RECT 23.66 2.94 23.675 3.136 ;
      RECT 23.635 2.92 23.66 3.124 ;
      RECT 23.595 2.89 23.635 3.104 ;
      RECT 23.585 2.86 23.595 3.089 ;
      RECT 23.57 2.85 23.585 3.082 ;
      RECT 23.515 2.815 23.57 3.061 ;
      RECT 23.5 2.778 23.515 3.04 ;
      RECT 23.49 2.765 23.5 3.032 ;
      RECT 23.44 2.735 23.49 3.014 ;
      RECT 23.425 2.665 23.44 2.995 ;
      RECT 23.38 2.665 23.425 2.978 ;
      RECT 23.355 2.665 23.38 2.96 ;
      RECT 23.345 2.665 23.355 2.953 ;
      RECT 23.266 2.665 23.345 2.946 ;
      RECT 23.18 2.665 23.266 2.938 ;
      RECT 23.165 2.697 23.18 2.933 ;
      RECT 23.09 2.707 23.165 2.929 ;
      RECT 23.07 2.717 23.09 2.924 ;
      RECT 23.045 2.717 23.07 2.921 ;
      RECT 23.035 2.707 23.045 2.92 ;
      RECT 23.025 2.68 23.035 2.919 ;
      RECT 22.985 2.675 23.025 2.917 ;
      RECT 22.94 2.675 22.985 2.913 ;
      RECT 22.915 2.675 22.94 2.908 ;
      RECT 22.865 2.675 22.915 2.895 ;
      RECT 22.825 2.68 22.835 2.88 ;
      RECT 22.835 2.675 22.865 2.885 ;
      RECT 24.82 2.455 25.08 2.715 ;
      RECT 24.815 2.477 25.08 2.673 ;
      RECT 24.055 2.305 24.275 2.67 ;
      RECT 24.037 2.392 24.275 2.669 ;
      RECT 24.02 2.397 24.275 2.666 ;
      RECT 24.02 2.397 24.295 2.665 ;
      RECT 23.99 2.407 24.295 2.663 ;
      RECT 23.985 2.422 24.295 2.659 ;
      RECT 23.985 2.422 24.3 2.658 ;
      RECT 23.98 2.48 24.3 2.656 ;
      RECT 23.98 2.48 24.31 2.653 ;
      RECT 23.975 2.545 24.31 2.648 ;
      RECT 24.055 2.305 24.315 2.565 ;
      RECT 22.8 2.135 23.06 2.395 ;
      RECT 22.8 2.178 23.146 2.369 ;
      RECT 22.8 2.178 23.19 2.368 ;
      RECT 22.8 2.178 23.21 2.366 ;
      RECT 22.8 2.178 23.31 2.365 ;
      RECT 22.8 2.178 23.33 2.363 ;
      RECT 22.8 2.178 23.34 2.358 ;
      RECT 23.21 2.145 23.4 2.355 ;
      RECT 23.21 2.147 23.405 2.353 ;
      RECT 23.2 2.152 23.41 2.345 ;
      RECT 23.146 2.176 23.41 2.345 ;
      RECT 23.19 2.17 23.2 2.367 ;
      RECT 23.2 2.15 23.405 2.353 ;
      RECT 22.155 3.21 22.36 3.44 ;
      RECT 22.095 3.16 22.15 3.42 ;
      RECT 22.155 3.16 22.355 3.44 ;
      RECT 23.125 3.475 23.13 3.502 ;
      RECT 23.115 3.385 23.125 3.507 ;
      RECT 23.11 3.307 23.115 3.513 ;
      RECT 23.1 3.297 23.11 3.52 ;
      RECT 23.095 3.287 23.1 3.526 ;
      RECT 23.085 3.282 23.095 3.528 ;
      RECT 23.07 3.274 23.085 3.536 ;
      RECT 23.055 3.265 23.07 3.548 ;
      RECT 23.045 3.257 23.055 3.558 ;
      RECT 23.01 3.175 23.045 3.576 ;
      RECT 22.975 3.175 23.01 3.595 ;
      RECT 22.96 3.175 22.975 3.603 ;
      RECT 22.905 3.175 22.96 3.603 ;
      RECT 22.871 3.175 22.905 3.594 ;
      RECT 22.785 3.175 22.871 3.57 ;
      RECT 22.775 3.235 22.785 3.552 ;
      RECT 22.735 3.237 22.775 3.543 ;
      RECT 22.73 3.239 22.735 3.533 ;
      RECT 22.71 3.241 22.73 3.528 ;
      RECT 22.7 3.244 22.71 3.523 ;
      RECT 22.69 3.245 22.7 3.518 ;
      RECT 22.666 3.246 22.69 3.51 ;
      RECT 22.58 3.251 22.666 3.488 ;
      RECT 22.525 3.25 22.58 3.461 ;
      RECT 22.51 3.243 22.525 3.448 ;
      RECT 22.475 3.238 22.51 3.444 ;
      RECT 22.42 3.23 22.475 3.443 ;
      RECT 22.36 3.217 22.42 3.441 ;
      RECT 22.15 3.16 22.155 3.428 ;
      RECT 22.225 2.53 22.41 2.74 ;
      RECT 22.215 2.535 22.425 2.733 ;
      RECT 22.255 2.44 22.515 2.7 ;
      RECT 22.21 2.597 22.515 2.623 ;
      RECT 21.555 2.39 21.56 3.19 ;
      RECT 21.5 2.44 21.53 3.19 ;
      RECT 21.49 2.44 21.495 2.75 ;
      RECT 21.475 2.44 21.48 2.745 ;
      RECT 21.02 2.485 21.035 2.7 ;
      RECT 20.95 2.485 21.035 2.695 ;
      RECT 22.215 2.065 22.285 2.275 ;
      RECT 22.285 2.072 22.295 2.27 ;
      RECT 22.181 2.065 22.215 2.282 ;
      RECT 22.095 2.065 22.181 2.306 ;
      RECT 22.085 2.07 22.095 2.325 ;
      RECT 22.08 2.082 22.085 2.328 ;
      RECT 22.065 2.097 22.08 2.332 ;
      RECT 22.06 2.115 22.065 2.336 ;
      RECT 22.02 2.125 22.06 2.345 ;
      RECT 22.005 2.132 22.02 2.357 ;
      RECT 21.99 2.137 22.005 2.362 ;
      RECT 21.975 2.14 21.99 2.367 ;
      RECT 21.965 2.142 21.975 2.371 ;
      RECT 21.93 2.149 21.965 2.379 ;
      RECT 21.895 2.157 21.93 2.393 ;
      RECT 21.885 2.163 21.895 2.402 ;
      RECT 21.88 2.165 21.885 2.404 ;
      RECT 21.86 2.168 21.88 2.41 ;
      RECT 21.83 2.175 21.86 2.421 ;
      RECT 21.82 2.181 21.83 2.428 ;
      RECT 21.795 2.184 21.82 2.435 ;
      RECT 21.785 2.188 21.795 2.443 ;
      RECT 21.78 2.189 21.785 2.465 ;
      RECT 21.775 2.19 21.78 2.48 ;
      RECT 21.77 2.191 21.775 2.495 ;
      RECT 21.765 2.192 21.77 2.51 ;
      RECT 21.76 2.193 21.765 2.54 ;
      RECT 21.75 2.195 21.76 2.573 ;
      RECT 21.735 2.199 21.75 2.62 ;
      RECT 21.725 2.202 21.735 2.665 ;
      RECT 21.72 2.205 21.725 2.693 ;
      RECT 21.71 2.207 21.72 2.72 ;
      RECT 21.705 2.21 21.71 2.755 ;
      RECT 21.675 2.215 21.705 2.813 ;
      RECT 21.67 2.22 21.675 2.898 ;
      RECT 21.665 2.222 21.67 2.933 ;
      RECT 21.66 2.224 21.665 3.015 ;
      RECT 21.655 2.226 21.66 3.103 ;
      RECT 21.645 2.228 21.655 3.185 ;
      RECT 21.63 2.242 21.645 3.19 ;
      RECT 21.595 2.287 21.63 3.19 ;
      RECT 21.585 2.327 21.595 3.19 ;
      RECT 21.57 2.355 21.585 3.19 ;
      RECT 21.565 2.372 21.57 3.19 ;
      RECT 21.56 2.38 21.565 3.19 ;
      RECT 21.55 2.395 21.555 3.19 ;
      RECT 21.545 2.402 21.55 3.19 ;
      RECT 21.535 2.422 21.545 3.19 ;
      RECT 21.53 2.435 21.535 3.19 ;
      RECT 21.495 2.44 21.5 2.775 ;
      RECT 21.48 2.83 21.5 3.19 ;
      RECT 21.48 2.44 21.49 2.748 ;
      RECT 21.475 2.87 21.48 3.19 ;
      RECT 21.425 2.44 21.475 2.743 ;
      RECT 21.47 2.907 21.475 3.19 ;
      RECT 21.46 2.93 21.47 3.19 ;
      RECT 21.455 2.975 21.46 3.19 ;
      RECT 21.445 2.985 21.455 3.183 ;
      RECT 21.371 2.44 21.425 2.737 ;
      RECT 21.285 2.44 21.371 2.73 ;
      RECT 21.236 2.487 21.285 2.723 ;
      RECT 21.15 2.495 21.236 2.716 ;
      RECT 21.135 2.492 21.15 2.711 ;
      RECT 21.121 2.485 21.135 2.71 ;
      RECT 21.035 2.485 21.121 2.705 ;
      RECT 20.94 2.49 20.95 2.69 ;
      RECT 20.53 1.92 20.545 2.32 ;
      RECT 20.725 1.92 20.73 2.18 ;
      RECT 20.47 1.92 20.515 2.18 ;
      RECT 20.925 3.225 20.93 3.43 ;
      RECT 20.92 3.215 20.925 3.435 ;
      RECT 20.915 3.202 20.92 3.44 ;
      RECT 20.91 3.182 20.915 3.44 ;
      RECT 20.885 3.135 20.91 3.44 ;
      RECT 20.85 3.05 20.885 3.44 ;
      RECT 20.845 2.987 20.85 3.44 ;
      RECT 20.84 2.972 20.845 3.44 ;
      RECT 20.825 2.932 20.84 3.44 ;
      RECT 20.82 2.907 20.825 3.44 ;
      RECT 20.81 2.89 20.82 3.44 ;
      RECT 20.775 2.812 20.81 3.44 ;
      RECT 20.77 2.755 20.775 3.44 ;
      RECT 20.765 2.742 20.77 3.44 ;
      RECT 20.755 2.72 20.765 3.44 ;
      RECT 20.745 2.685 20.755 3.44 ;
      RECT 20.735 2.655 20.745 3.44 ;
      RECT 20.725 2.57 20.735 3.083 ;
      RECT 20.732 3.215 20.735 3.44 ;
      RECT 20.73 3.225 20.732 3.44 ;
      RECT 20.72 3.235 20.73 3.435 ;
      RECT 20.715 1.92 20.725 2.315 ;
      RECT 20.72 2.447 20.725 3.058 ;
      RECT 20.715 2.345 20.72 3.041 ;
      RECT 20.705 1.92 20.715 3.017 ;
      RECT 20.7 1.92 20.705 2.988 ;
      RECT 20.695 1.92 20.7 2.978 ;
      RECT 20.675 1.92 20.695 2.94 ;
      RECT 20.67 1.92 20.675 2.898 ;
      RECT 20.665 1.92 20.67 2.878 ;
      RECT 20.635 1.92 20.665 2.828 ;
      RECT 20.625 1.92 20.635 2.775 ;
      RECT 20.62 1.92 20.625 2.748 ;
      RECT 20.615 1.92 20.62 2.733 ;
      RECT 20.605 1.92 20.615 2.71 ;
      RECT 20.595 1.92 20.605 2.685 ;
      RECT 20.59 1.92 20.595 2.625 ;
      RECT 20.58 1.92 20.59 2.563 ;
      RECT 20.575 1.92 20.58 2.483 ;
      RECT 20.57 1.92 20.575 2.448 ;
      RECT 20.565 1.92 20.57 2.423 ;
      RECT 20.56 1.92 20.565 2.408 ;
      RECT 20.555 1.92 20.56 2.378 ;
      RECT 20.55 1.92 20.555 2.355 ;
      RECT 20.545 1.92 20.55 2.328 ;
      RECT 20.515 1.92 20.53 2.315 ;
      RECT 19.67 3.455 19.855 3.665 ;
      RECT 19.66 3.46 19.87 3.658 ;
      RECT 19.66 3.46 19.89 3.63 ;
      RECT 19.66 3.46 19.905 3.609 ;
      RECT 19.66 3.46 19.92 3.607 ;
      RECT 19.66 3.46 19.93 3.606 ;
      RECT 19.66 3.46 19.96 3.603 ;
      RECT 20.31 3.305 20.57 3.565 ;
      RECT 20.27 3.352 20.57 3.548 ;
      RECT 20.261 3.36 20.27 3.551 ;
      RECT 19.855 3.453 20.57 3.548 ;
      RECT 20.175 3.378 20.261 3.558 ;
      RECT 19.87 3.45 20.57 3.548 ;
      RECT 20.116 3.4 20.175 3.57 ;
      RECT 19.89 3.446 20.57 3.548 ;
      RECT 20.03 3.412 20.116 3.581 ;
      RECT 19.905 3.442 20.57 3.548 ;
      RECT 19.975 3.425 20.03 3.593 ;
      RECT 19.92 3.44 20.57 3.548 ;
      RECT 19.96 3.431 19.975 3.599 ;
      RECT 19.93 3.436 20.57 3.548 ;
      RECT 20.075 2.96 20.335 3.22 ;
      RECT 20.075 2.98 20.445 3.19 ;
      RECT 20.075 2.985 20.455 3.185 ;
      RECT 20.266 2.399 20.345 2.63 ;
      RECT 20.18 2.402 20.395 2.625 ;
      RECT 20.175 2.402 20.395 2.62 ;
      RECT 20.175 2.407 20.405 2.618 ;
      RECT 20.15 2.407 20.405 2.615 ;
      RECT 20.15 2.415 20.415 2.613 ;
      RECT 20.03 2.35 20.29 2.61 ;
      RECT 20.03 2.397 20.34 2.61 ;
      RECT 19.285 2.97 19.29 3.23 ;
      RECT 19.115 2.74 19.12 3.23 ;
      RECT 19 2.98 19.005 3.205 ;
      RECT 19.71 2.075 19.715 2.285 ;
      RECT 19.715 2.08 19.73 2.28 ;
      RECT 19.65 2.075 19.71 2.293 ;
      RECT 19.635 2.075 19.65 2.303 ;
      RECT 19.585 2.075 19.635 2.32 ;
      RECT 19.565 2.075 19.585 2.343 ;
      RECT 19.55 2.075 19.565 2.355 ;
      RECT 19.53 2.075 19.55 2.365 ;
      RECT 19.52 2.08 19.53 2.374 ;
      RECT 19.515 2.09 19.52 2.379 ;
      RECT 19.51 2.102 19.515 2.383 ;
      RECT 19.5 2.125 19.51 2.388 ;
      RECT 19.495 2.14 19.5 2.392 ;
      RECT 19.49 2.157 19.495 2.395 ;
      RECT 19.485 2.165 19.49 2.398 ;
      RECT 19.475 2.17 19.485 2.402 ;
      RECT 19.47 2.177 19.475 2.407 ;
      RECT 19.46 2.182 19.47 2.411 ;
      RECT 19.435 2.194 19.46 2.422 ;
      RECT 19.415 2.211 19.435 2.438 ;
      RECT 19.39 2.228 19.415 2.46 ;
      RECT 19.355 2.251 19.39 2.518 ;
      RECT 19.335 2.273 19.355 2.58 ;
      RECT 19.33 2.283 19.335 2.615 ;
      RECT 19.32 2.29 19.33 2.653 ;
      RECT 19.315 2.297 19.32 2.673 ;
      RECT 19.31 2.308 19.315 2.71 ;
      RECT 19.305 2.316 19.31 2.775 ;
      RECT 19.295 2.327 19.305 2.828 ;
      RECT 19.29 2.345 19.295 2.898 ;
      RECT 19.285 2.355 19.29 2.935 ;
      RECT 19.28 2.365 19.285 3.23 ;
      RECT 19.275 2.377 19.28 3.23 ;
      RECT 19.27 2.387 19.275 3.23 ;
      RECT 19.26 2.397 19.27 3.23 ;
      RECT 19.25 2.42 19.26 3.23 ;
      RECT 19.235 2.455 19.25 3.23 ;
      RECT 19.195 2.517 19.235 3.23 ;
      RECT 19.19 2.57 19.195 3.23 ;
      RECT 19.165 2.605 19.19 3.23 ;
      RECT 19.15 2.65 19.165 3.23 ;
      RECT 19.145 2.672 19.15 3.23 ;
      RECT 19.135 2.685 19.145 3.23 ;
      RECT 19.125 2.71 19.135 3.23 ;
      RECT 19.12 2.732 19.125 3.23 ;
      RECT 19.095 2.77 19.115 3.23 ;
      RECT 19.055 2.827 19.095 3.23 ;
      RECT 19.05 2.877 19.055 3.23 ;
      RECT 19.045 2.895 19.05 3.23 ;
      RECT 19.04 2.907 19.045 3.23 ;
      RECT 19.03 2.925 19.04 3.23 ;
      RECT 19.02 2.945 19.03 3.205 ;
      RECT 19.015 2.962 19.02 3.205 ;
      RECT 19.005 2.975 19.015 3.205 ;
      RECT 18.975 2.985 19 3.205 ;
      RECT 18.965 2.992 18.975 3.205 ;
      RECT 18.95 3.002 18.965 3.2 ;
      RECT 18.045 7.77 18.335 8 ;
      RECT 18.105 6.29 18.275 8 ;
      RECT 18.1 6.655 18.45 7.005 ;
      RECT 18.045 6.29 18.335 6.52 ;
      RECT 17.64 2.395 17.745 2.965 ;
      RECT 17.64 2.73 17.965 2.96 ;
      RECT 17.64 2.76 18.135 2.93 ;
      RECT 17.64 2.395 17.83 2.96 ;
      RECT 17.055 2.36 17.345 2.59 ;
      RECT 17.055 2.395 17.83 2.565 ;
      RECT 17.115 0.88 17.285 2.59 ;
      RECT 17.055 0.88 17.345 1.11 ;
      RECT 17.055 7.77 17.345 8 ;
      RECT 17.115 6.29 17.285 8 ;
      RECT 17.055 6.29 17.345 6.52 ;
      RECT 17.055 6.325 17.91 6.485 ;
      RECT 17.74 5.92 17.91 6.485 ;
      RECT 17.055 6.32 17.45 6.485 ;
      RECT 17.675 5.92 17.965 6.15 ;
      RECT 17.675 5.95 18.135 6.12 ;
      RECT 16.685 2.73 16.975 2.96 ;
      RECT 16.685 2.76 17.145 2.93 ;
      RECT 16.75 1.655 16.915 2.96 ;
      RECT 15.265 1.625 15.555 1.855 ;
      RECT 15.265 1.655 16.915 1.825 ;
      RECT 15.325 0.885 15.495 1.855 ;
      RECT 15.265 0.885 15.555 1.115 ;
      RECT 15.265 7.765 15.555 7.995 ;
      RECT 15.325 7.025 15.495 7.995 ;
      RECT 15.325 7.12 16.915 7.29 ;
      RECT 16.745 5.92 16.915 7.29 ;
      RECT 15.265 7.025 15.555 7.255 ;
      RECT 16.685 5.92 16.975 6.15 ;
      RECT 16.685 5.95 17.145 6.12 ;
      RECT 15.695 1.965 16.045 2.315 ;
      RECT 13.36 2.025 16.045 2.195 ;
      RECT 13.36 1.34 13.53 2.195 ;
      RECT 13.26 1.34 13.61 1.69 ;
      RECT 15.72 6.655 16.045 6.98 ;
      RECT 11.115 6.605 11.465 6.955 ;
      RECT 15.695 6.655 16.045 6.885 ;
      RECT 10.915 6.655 11.465 6.885 ;
      RECT 10.745 6.685 16.045 6.855 ;
      RECT 14.92 2.365 15.24 2.685 ;
      RECT 14.89 2.365 15.24 2.595 ;
      RECT 14.72 2.395 15.24 2.565 ;
      RECT 14.92 6.255 15.24 6.545 ;
      RECT 14.89 6.285 15.24 6.515 ;
      RECT 14.72 6.315 15.24 6.485 ;
      RECT 11.555 2.465 11.74 2.675 ;
      RECT 11.545 2.47 11.755 2.668 ;
      RECT 11.545 2.47 11.841 2.645 ;
      RECT 11.545 2.47 11.9 2.62 ;
      RECT 11.545 2.47 11.955 2.6 ;
      RECT 11.545 2.47 11.965 2.588 ;
      RECT 11.545 2.47 12.16 2.527 ;
      RECT 11.545 2.47 12.19 2.51 ;
      RECT 11.545 2.47 12.21 2.5 ;
      RECT 12.09 2.235 12.35 2.495 ;
      RECT 12.075 2.325 12.09 2.542 ;
      RECT 11.61 2.457 12.35 2.495 ;
      RECT 12.061 2.336 12.075 2.548 ;
      RECT 11.65 2.45 12.35 2.495 ;
      RECT 11.975 2.376 12.061 2.567 ;
      RECT 11.9 2.437 12.35 2.495 ;
      RECT 11.97 2.412 11.975 2.584 ;
      RECT 11.955 2.422 12.35 2.495 ;
      RECT 11.965 2.417 11.97 2.586 ;
      RECT 12.26 2.922 12.265 3.014 ;
      RECT 12.255 2.9 12.26 3.031 ;
      RECT 12.25 2.89 12.255 3.043 ;
      RECT 12.24 2.881 12.25 3.053 ;
      RECT 12.235 2.876 12.24 3.061 ;
      RECT 12.23 2.735 12.235 3.064 ;
      RECT 12.196 2.735 12.23 3.075 ;
      RECT 12.11 2.735 12.196 3.11 ;
      RECT 12.03 2.735 12.11 3.158 ;
      RECT 12.001 2.735 12.03 3.182 ;
      RECT 11.915 2.735 12.001 3.188 ;
      RECT 11.91 2.919 11.915 3.193 ;
      RECT 11.875 2.93 11.91 3.196 ;
      RECT 11.85 2.945 11.875 3.2 ;
      RECT 11.836 2.954 11.85 3.202 ;
      RECT 11.75 2.981 11.836 3.208 ;
      RECT 11.685 3.022 11.75 3.217 ;
      RECT 11.67 3.042 11.685 3.222 ;
      RECT 11.64 3.052 11.67 3.225 ;
      RECT 11.635 3.062 11.64 3.228 ;
      RECT 11.605 3.067 11.635 3.23 ;
      RECT 11.585 3.072 11.605 3.234 ;
      RECT 11.5 3.075 11.585 3.241 ;
      RECT 11.485 3.072 11.5 3.247 ;
      RECT 11.475 3.069 11.485 3.249 ;
      RECT 11.455 3.066 11.475 3.251 ;
      RECT 11.435 3.062 11.455 3.252 ;
      RECT 11.42 3.058 11.435 3.254 ;
      RECT 11.41 3.055 11.42 3.255 ;
      RECT 11.37 3.049 11.41 3.253 ;
      RECT 11.36 3.044 11.37 3.251 ;
      RECT 11.345 3.041 11.36 3.247 ;
      RECT 11.32 3.036 11.345 3.24 ;
      RECT 11.27 3.027 11.32 3.228 ;
      RECT 11.2 3.013 11.27 3.21 ;
      RECT 11.142 2.998 11.2 3.192 ;
      RECT 11.056 2.981 11.142 3.172 ;
      RECT 10.97 2.96 11.056 3.147 ;
      RECT 10.92 2.945 10.97 3.128 ;
      RECT 10.916 2.939 10.92 3.12 ;
      RECT 10.83 2.929 10.916 3.107 ;
      RECT 10.795 2.914 10.83 3.09 ;
      RECT 10.78 2.907 10.795 3.083 ;
      RECT 10.72 2.895 10.78 3.071 ;
      RECT 10.7 2.882 10.72 3.059 ;
      RECT 10.66 2.873 10.7 3.051 ;
      RECT 10.655 2.865 10.66 3.044 ;
      RECT 10.575 2.855 10.655 3.03 ;
      RECT 10.56 2.842 10.575 3.015 ;
      RECT 10.555 2.84 10.56 3.013 ;
      RECT 10.476 2.828 10.555 3 ;
      RECT 10.39 2.803 10.476 2.975 ;
      RECT 10.375 2.772 10.39 2.96 ;
      RECT 10.36 2.747 10.375 2.956 ;
      RECT 10.345 2.74 10.36 2.952 ;
      RECT 10.17 2.745 10.175 2.948 ;
      RECT 10.165 2.75 10.17 2.943 ;
      RECT 10.175 2.74 10.345 2.95 ;
      RECT 10.89 2.5 10.995 2.76 ;
      RECT 11.705 2.025 11.71 2.25 ;
      RECT 11.835 2.025 11.89 2.235 ;
      RECT 11.89 2.03 11.9 2.228 ;
      RECT 11.796 2.025 11.835 2.238 ;
      RECT 11.71 2.025 11.796 2.245 ;
      RECT 11.69 2.03 11.705 2.251 ;
      RECT 11.68 2.07 11.69 2.253 ;
      RECT 11.65 2.08 11.68 2.255 ;
      RECT 11.645 2.085 11.65 2.257 ;
      RECT 11.62 2.09 11.645 2.259 ;
      RECT 11.605 2.095 11.62 2.261 ;
      RECT 11.59 2.097 11.605 2.263 ;
      RECT 11.585 2.102 11.59 2.265 ;
      RECT 11.535 2.11 11.585 2.268 ;
      RECT 11.51 2.119 11.535 2.273 ;
      RECT 11.5 2.126 11.51 2.278 ;
      RECT 11.495 2.129 11.5 2.282 ;
      RECT 11.475 2.132 11.495 2.291 ;
      RECT 11.445 2.14 11.475 2.311 ;
      RECT 11.416 2.153 11.445 2.333 ;
      RECT 11.33 2.187 11.416 2.377 ;
      RECT 11.325 2.213 11.33 2.415 ;
      RECT 11.32 2.217 11.325 2.424 ;
      RECT 11.285 2.23 11.32 2.457 ;
      RECT 11.275 2.244 11.285 2.495 ;
      RECT 11.27 2.248 11.275 2.508 ;
      RECT 11.265 2.252 11.27 2.513 ;
      RECT 11.255 2.26 11.265 2.525 ;
      RECT 11.25 2.267 11.255 2.54 ;
      RECT 11.225 2.28 11.25 2.565 ;
      RECT 11.185 2.309 11.225 2.62 ;
      RECT 11.17 2.334 11.185 2.675 ;
      RECT 11.16 2.345 11.17 2.698 ;
      RECT 11.155 2.352 11.16 2.71 ;
      RECT 11.15 2.356 11.155 2.718 ;
      RECT 11.095 2.384 11.15 2.76 ;
      RECT 11.075 2.42 11.095 2.76 ;
      RECT 11.06 2.435 11.075 2.76 ;
      RECT 11.005 2.467 11.06 2.76 ;
      RECT 10.995 2.497 11.005 2.76 ;
      RECT 10.605 2.112 10.79 2.35 ;
      RECT 10.59 2.114 10.8 2.345 ;
      RECT 10.475 2.06 10.735 2.32 ;
      RECT 10.47 2.097 10.735 2.274 ;
      RECT 10.465 2.107 10.735 2.271 ;
      RECT 10.46 2.147 10.8 2.265 ;
      RECT 10.455 2.18 10.8 2.255 ;
      RECT 10.465 2.122 10.815 2.193 ;
      RECT 10.762 3.22 10.775 3.75 ;
      RECT 10.676 3.22 10.775 3.749 ;
      RECT 10.676 3.22 10.78 3.748 ;
      RECT 10.59 3.22 10.78 3.746 ;
      RECT 10.585 3.22 10.78 3.743 ;
      RECT 10.585 3.22 10.79 3.741 ;
      RECT 10.58 3.512 10.79 3.738 ;
      RECT 10.58 3.522 10.795 3.735 ;
      RECT 10.58 3.59 10.8 3.731 ;
      RECT 10.57 3.595 10.8 3.73 ;
      RECT 10.57 3.687 10.805 3.727 ;
      RECT 10.555 3.22 10.815 3.48 ;
      RECT 10.485 7.765 10.775 7.995 ;
      RECT 10.545 7.025 10.715 7.995 ;
      RECT 10.46 7.055 10.8 7.4 ;
      RECT 10.485 7.025 10.775 7.4 ;
      RECT 9.785 2.21 9.83 3.745 ;
      RECT 9.985 2.21 10.015 2.425 ;
      RECT 8.36 1.95 8.48 2.16 ;
      RECT 8.02 1.9 8.28 2.16 ;
      RECT 8.02 1.945 8.315 2.15 ;
      RECT 10.025 2.226 10.03 2.28 ;
      RECT 10.02 2.219 10.025 2.413 ;
      RECT 10.015 2.213 10.02 2.42 ;
      RECT 9.97 2.21 9.985 2.433 ;
      RECT 9.965 2.21 9.97 2.455 ;
      RECT 9.96 2.21 9.965 2.503 ;
      RECT 9.955 2.21 9.96 2.523 ;
      RECT 9.945 2.21 9.955 2.63 ;
      RECT 9.94 2.21 9.945 2.693 ;
      RECT 9.935 2.21 9.94 2.75 ;
      RECT 9.93 2.21 9.935 2.758 ;
      RECT 9.915 2.21 9.93 2.865 ;
      RECT 9.905 2.21 9.915 3 ;
      RECT 9.895 2.21 9.905 3.11 ;
      RECT 9.885 2.21 9.895 3.167 ;
      RECT 9.88 2.21 9.885 3.207 ;
      RECT 9.875 2.21 9.88 3.243 ;
      RECT 9.865 2.21 9.875 3.283 ;
      RECT 9.86 2.21 9.865 3.325 ;
      RECT 9.84 2.21 9.86 3.39 ;
      RECT 9.845 3.535 9.85 3.715 ;
      RECT 9.84 3.517 9.845 3.723 ;
      RECT 9.835 2.21 9.84 3.453 ;
      RECT 9.835 3.497 9.84 3.73 ;
      RECT 9.83 2.21 9.835 3.74 ;
      RECT 9.775 2.21 9.785 2.51 ;
      RECT 9.78 2.757 9.785 3.745 ;
      RECT 9.775 2.822 9.78 3.745 ;
      RECT 9.77 2.211 9.775 2.5 ;
      RECT 9.765 2.887 9.775 3.745 ;
      RECT 9.76 2.212 9.77 2.49 ;
      RECT 9.75 3 9.765 3.745 ;
      RECT 9.755 2.213 9.76 2.48 ;
      RECT 9.735 2.214 9.755 2.458 ;
      RECT 9.74 3.097 9.75 3.745 ;
      RECT 9.735 3.172 9.74 3.745 ;
      RECT 9.725 2.213 9.735 2.435 ;
      RECT 9.73 3.215 9.735 3.745 ;
      RECT 9.725 3.242 9.73 3.745 ;
      RECT 9.715 2.211 9.725 2.423 ;
      RECT 9.72 3.285 9.725 3.745 ;
      RECT 9.715 3.312 9.72 3.745 ;
      RECT 9.705 2.21 9.715 2.41 ;
      RECT 9.71 3.327 9.715 3.745 ;
      RECT 9.67 3.385 9.71 3.745 ;
      RECT 9.7 2.209 9.705 2.395 ;
      RECT 9.695 2.207 9.7 2.388 ;
      RECT 9.685 2.204 9.695 2.378 ;
      RECT 9.68 2.201 9.685 2.363 ;
      RECT 9.665 2.197 9.68 2.356 ;
      RECT 9.66 3.44 9.67 3.745 ;
      RECT 9.66 2.194 9.665 2.351 ;
      RECT 9.645 2.19 9.66 2.345 ;
      RECT 9.655 3.457 9.66 3.745 ;
      RECT 9.645 3.52 9.655 3.745 ;
      RECT 9.565 2.175 9.645 2.325 ;
      RECT 9.64 3.527 9.645 3.74 ;
      RECT 9.635 3.535 9.64 3.73 ;
      RECT 9.555 2.161 9.565 2.309 ;
      RECT 9.54 2.157 9.555 2.307 ;
      RECT 9.53 2.152 9.54 2.303 ;
      RECT 9.505 2.145 9.53 2.295 ;
      RECT 9.5 2.14 9.505 2.29 ;
      RECT 9.49 2.14 9.5 2.288 ;
      RECT 9.48 2.138 9.49 2.286 ;
      RECT 9.45 2.13 9.48 2.28 ;
      RECT 9.435 2.122 9.45 2.273 ;
      RECT 9.415 2.117 9.435 2.266 ;
      RECT 9.41 2.113 9.415 2.261 ;
      RECT 9.38 2.106 9.41 2.255 ;
      RECT 9.355 2.097 9.38 2.245 ;
      RECT 9.325 2.09 9.355 2.237 ;
      RECT 9.3 2.08 9.325 2.228 ;
      RECT 9.285 2.072 9.3 2.222 ;
      RECT 9.26 2.067 9.285 2.217 ;
      RECT 9.25 2.063 9.26 2.212 ;
      RECT 9.23 2.058 9.25 2.207 ;
      RECT 9.195 2.053 9.23 2.2 ;
      RECT 9.135 2.048 9.195 2.193 ;
      RECT 9.122 2.044 9.135 2.191 ;
      RECT 9.036 2.039 9.122 2.188 ;
      RECT 8.95 2.029 9.036 2.184 ;
      RECT 8.909 2.022 8.95 2.181 ;
      RECT 8.823 2.015 8.909 2.178 ;
      RECT 8.737 2.005 8.823 2.174 ;
      RECT 8.651 1.995 8.737 2.169 ;
      RECT 8.565 1.985 8.651 2.165 ;
      RECT 8.555 1.97 8.565 2.163 ;
      RECT 8.545 1.955 8.555 2.163 ;
      RECT 8.48 1.95 8.545 2.162 ;
      RECT 8.315 1.947 8.36 2.155 ;
      RECT 9.56 2.852 9.565 3.043 ;
      RECT 9.555 2.847 9.56 3.05 ;
      RECT 9.541 2.845 9.555 3.056 ;
      RECT 9.455 2.845 9.541 3.058 ;
      RECT 9.451 2.845 9.455 3.061 ;
      RECT 9.365 2.845 9.451 3.079 ;
      RECT 9.355 2.85 9.365 3.098 ;
      RECT 9.345 2.905 9.355 3.102 ;
      RECT 9.32 2.92 9.345 3.109 ;
      RECT 9.28 2.94 9.32 3.122 ;
      RECT 9.275 2.952 9.28 3.132 ;
      RECT 9.26 2.958 9.275 3.137 ;
      RECT 9.255 2.963 9.26 3.141 ;
      RECT 9.235 2.97 9.255 3.146 ;
      RECT 9.165 2.995 9.235 3.163 ;
      RECT 9.125 3.023 9.165 3.183 ;
      RECT 9.12 3.033 9.125 3.191 ;
      RECT 9.1 3.04 9.12 3.193 ;
      RECT 9.095 3.047 9.1 3.196 ;
      RECT 9.065 3.055 9.095 3.199 ;
      RECT 9.06 3.06 9.065 3.203 ;
      RECT 8.986 3.064 9.06 3.211 ;
      RECT 8.9 3.073 8.986 3.227 ;
      RECT 8.896 3.078 8.9 3.236 ;
      RECT 8.81 3.083 8.896 3.246 ;
      RECT 8.77 3.091 8.81 3.258 ;
      RECT 8.72 3.097 8.77 3.265 ;
      RECT 8.635 3.106 8.72 3.28 ;
      RECT 8.56 3.117 8.635 3.298 ;
      RECT 8.525 3.124 8.56 3.308 ;
      RECT 8.45 3.132 8.525 3.313 ;
      RECT 8.395 3.141 8.45 3.313 ;
      RECT 8.37 3.146 8.395 3.311 ;
      RECT 8.36 3.149 8.37 3.309 ;
      RECT 8.325 3.151 8.36 3.307 ;
      RECT 8.295 3.153 8.325 3.303 ;
      RECT 8.25 3.152 8.295 3.299 ;
      RECT 8.23 3.147 8.25 3.296 ;
      RECT 8.18 3.132 8.23 3.293 ;
      RECT 8.17 3.117 8.18 3.288 ;
      RECT 8.12 3.102 8.17 3.278 ;
      RECT 8.07 3.077 8.12 3.258 ;
      RECT 8.06 3.062 8.07 3.24 ;
      RECT 8.055 3.06 8.06 3.234 ;
      RECT 8.035 3.055 8.055 3.229 ;
      RECT 8.03 3.047 8.035 3.223 ;
      RECT 8.015 3.041 8.03 3.216 ;
      RECT 8.01 3.036 8.015 3.208 ;
      RECT 7.99 3.031 8.01 3.2 ;
      RECT 7.975 3.024 7.99 3.193 ;
      RECT 7.96 3.018 7.975 3.184 ;
      RECT 7.955 3.012 7.96 3.177 ;
      RECT 7.91 2.987 7.955 3.163 ;
      RECT 7.895 2.957 7.91 3.145 ;
      RECT 7.88 2.94 7.895 3.136 ;
      RECT 7.855 2.92 7.88 3.124 ;
      RECT 7.815 2.89 7.855 3.104 ;
      RECT 7.805 2.86 7.815 3.089 ;
      RECT 7.79 2.85 7.805 3.082 ;
      RECT 7.735 2.815 7.79 3.061 ;
      RECT 7.72 2.778 7.735 3.04 ;
      RECT 7.71 2.765 7.72 3.032 ;
      RECT 7.66 2.735 7.71 3.014 ;
      RECT 7.645 2.665 7.66 2.995 ;
      RECT 7.6 2.665 7.645 2.978 ;
      RECT 7.575 2.665 7.6 2.96 ;
      RECT 7.565 2.665 7.575 2.953 ;
      RECT 7.486 2.665 7.565 2.946 ;
      RECT 7.4 2.665 7.486 2.938 ;
      RECT 7.385 2.697 7.4 2.933 ;
      RECT 7.31 2.707 7.385 2.929 ;
      RECT 7.29 2.717 7.31 2.924 ;
      RECT 7.265 2.717 7.29 2.921 ;
      RECT 7.255 2.707 7.265 2.92 ;
      RECT 7.245 2.68 7.255 2.919 ;
      RECT 7.205 2.675 7.245 2.917 ;
      RECT 7.16 2.675 7.205 2.913 ;
      RECT 7.135 2.675 7.16 2.908 ;
      RECT 7.085 2.675 7.135 2.895 ;
      RECT 7.045 2.68 7.055 2.88 ;
      RECT 7.055 2.675 7.085 2.885 ;
      RECT 9.04 2.455 9.3 2.715 ;
      RECT 9.035 2.477 9.3 2.673 ;
      RECT 8.275 2.305 8.495 2.67 ;
      RECT 8.257 2.392 8.495 2.669 ;
      RECT 8.24 2.397 8.495 2.666 ;
      RECT 8.24 2.397 8.515 2.665 ;
      RECT 8.21 2.407 8.515 2.663 ;
      RECT 8.205 2.422 8.515 2.659 ;
      RECT 8.205 2.422 8.52 2.658 ;
      RECT 8.2 2.48 8.52 2.656 ;
      RECT 8.2 2.48 8.53 2.653 ;
      RECT 8.195 2.545 8.53 2.648 ;
      RECT 8.275 2.305 8.535 2.565 ;
      RECT 7.02 2.135 7.28 2.395 ;
      RECT 7.02 2.178 7.366 2.369 ;
      RECT 7.02 2.178 7.41 2.368 ;
      RECT 7.02 2.178 7.43 2.366 ;
      RECT 7.02 2.178 7.53 2.365 ;
      RECT 7.02 2.178 7.55 2.363 ;
      RECT 7.02 2.178 7.56 2.358 ;
      RECT 7.43 2.145 7.62 2.355 ;
      RECT 7.43 2.147 7.625 2.353 ;
      RECT 7.42 2.152 7.63 2.345 ;
      RECT 7.366 2.176 7.63 2.345 ;
      RECT 7.41 2.17 7.42 2.367 ;
      RECT 7.42 2.15 7.625 2.353 ;
      RECT 6.375 3.21 6.58 3.44 ;
      RECT 6.315 3.16 6.37 3.42 ;
      RECT 6.375 3.16 6.575 3.44 ;
      RECT 7.345 3.475 7.35 3.502 ;
      RECT 7.335 3.385 7.345 3.507 ;
      RECT 7.33 3.307 7.335 3.513 ;
      RECT 7.32 3.297 7.33 3.52 ;
      RECT 7.315 3.287 7.32 3.526 ;
      RECT 7.305 3.282 7.315 3.528 ;
      RECT 7.29 3.274 7.305 3.536 ;
      RECT 7.275 3.265 7.29 3.548 ;
      RECT 7.265 3.257 7.275 3.558 ;
      RECT 7.23 3.175 7.265 3.576 ;
      RECT 7.195 3.175 7.23 3.595 ;
      RECT 7.18 3.175 7.195 3.603 ;
      RECT 7.125 3.175 7.18 3.603 ;
      RECT 7.091 3.175 7.125 3.594 ;
      RECT 7.005 3.175 7.091 3.57 ;
      RECT 6.995 3.235 7.005 3.552 ;
      RECT 6.955 3.237 6.995 3.543 ;
      RECT 6.95 3.239 6.955 3.533 ;
      RECT 6.93 3.241 6.95 3.528 ;
      RECT 6.92 3.244 6.93 3.523 ;
      RECT 6.91 3.245 6.92 3.518 ;
      RECT 6.886 3.246 6.91 3.51 ;
      RECT 6.8 3.251 6.886 3.488 ;
      RECT 6.745 3.25 6.8 3.461 ;
      RECT 6.73 3.243 6.745 3.448 ;
      RECT 6.695 3.238 6.73 3.444 ;
      RECT 6.64 3.23 6.695 3.443 ;
      RECT 6.58 3.217 6.64 3.441 ;
      RECT 6.37 3.16 6.375 3.428 ;
      RECT 6.445 2.53 6.63 2.74 ;
      RECT 6.435 2.535 6.645 2.733 ;
      RECT 6.475 2.44 6.735 2.7 ;
      RECT 6.43 2.597 6.735 2.623 ;
      RECT 5.775 2.39 5.78 3.19 ;
      RECT 5.72 2.44 5.75 3.19 ;
      RECT 5.71 2.44 5.715 2.75 ;
      RECT 5.695 2.44 5.7 2.745 ;
      RECT 5.24 2.485 5.255 2.7 ;
      RECT 5.17 2.485 5.255 2.695 ;
      RECT 6.435 2.065 6.505 2.275 ;
      RECT 6.505 2.072 6.515 2.27 ;
      RECT 6.401 2.065 6.435 2.282 ;
      RECT 6.315 2.065 6.401 2.306 ;
      RECT 6.305 2.07 6.315 2.325 ;
      RECT 6.3 2.082 6.305 2.328 ;
      RECT 6.285 2.097 6.3 2.332 ;
      RECT 6.28 2.115 6.285 2.336 ;
      RECT 6.24 2.125 6.28 2.345 ;
      RECT 6.225 2.132 6.24 2.357 ;
      RECT 6.21 2.137 6.225 2.362 ;
      RECT 6.195 2.14 6.21 2.367 ;
      RECT 6.185 2.142 6.195 2.371 ;
      RECT 6.15 2.149 6.185 2.379 ;
      RECT 6.115 2.157 6.15 2.393 ;
      RECT 6.105 2.163 6.115 2.402 ;
      RECT 6.1 2.165 6.105 2.404 ;
      RECT 6.08 2.168 6.1 2.41 ;
      RECT 6.05 2.175 6.08 2.421 ;
      RECT 6.04 2.181 6.05 2.428 ;
      RECT 6.015 2.184 6.04 2.435 ;
      RECT 6.005 2.188 6.015 2.443 ;
      RECT 6 2.189 6.005 2.465 ;
      RECT 5.995 2.19 6 2.48 ;
      RECT 5.99 2.191 5.995 2.495 ;
      RECT 5.985 2.192 5.99 2.51 ;
      RECT 5.98 2.193 5.985 2.54 ;
      RECT 5.97 2.195 5.98 2.573 ;
      RECT 5.955 2.199 5.97 2.62 ;
      RECT 5.945 2.202 5.955 2.665 ;
      RECT 5.94 2.205 5.945 2.693 ;
      RECT 5.93 2.207 5.94 2.72 ;
      RECT 5.925 2.21 5.93 2.755 ;
      RECT 5.895 2.215 5.925 2.813 ;
      RECT 5.89 2.22 5.895 2.898 ;
      RECT 5.885 2.222 5.89 2.933 ;
      RECT 5.88 2.224 5.885 3.015 ;
      RECT 5.875 2.226 5.88 3.103 ;
      RECT 5.865 2.228 5.875 3.185 ;
      RECT 5.85 2.242 5.865 3.19 ;
      RECT 5.815 2.287 5.85 3.19 ;
      RECT 5.805 2.327 5.815 3.19 ;
      RECT 5.79 2.355 5.805 3.19 ;
      RECT 5.785 2.372 5.79 3.19 ;
      RECT 5.78 2.38 5.785 3.19 ;
      RECT 5.77 2.395 5.775 3.19 ;
      RECT 5.765 2.402 5.77 3.19 ;
      RECT 5.755 2.422 5.765 3.19 ;
      RECT 5.75 2.435 5.755 3.19 ;
      RECT 5.715 2.44 5.72 2.775 ;
      RECT 5.7 2.83 5.72 3.19 ;
      RECT 5.7 2.44 5.71 2.748 ;
      RECT 5.695 2.87 5.7 3.19 ;
      RECT 5.645 2.44 5.695 2.743 ;
      RECT 5.69 2.907 5.695 3.19 ;
      RECT 5.68 2.93 5.69 3.19 ;
      RECT 5.675 2.975 5.68 3.19 ;
      RECT 5.665 2.985 5.675 3.183 ;
      RECT 5.591 2.44 5.645 2.737 ;
      RECT 5.505 2.44 5.591 2.73 ;
      RECT 5.456 2.487 5.505 2.723 ;
      RECT 5.37 2.495 5.456 2.716 ;
      RECT 5.355 2.492 5.37 2.711 ;
      RECT 5.341 2.485 5.355 2.71 ;
      RECT 5.255 2.485 5.341 2.705 ;
      RECT 5.16 2.49 5.17 2.69 ;
      RECT 4.75 1.92 4.765 2.32 ;
      RECT 4.945 1.92 4.95 2.18 ;
      RECT 4.69 1.92 4.735 2.18 ;
      RECT 5.145 3.225 5.15 3.43 ;
      RECT 5.14 3.215 5.145 3.435 ;
      RECT 5.135 3.202 5.14 3.44 ;
      RECT 5.13 3.182 5.135 3.44 ;
      RECT 5.105 3.135 5.13 3.44 ;
      RECT 5.07 3.05 5.105 3.44 ;
      RECT 5.065 2.987 5.07 3.44 ;
      RECT 5.06 2.972 5.065 3.44 ;
      RECT 5.045 2.932 5.06 3.44 ;
      RECT 5.04 2.907 5.045 3.44 ;
      RECT 5.03 2.89 5.04 3.44 ;
      RECT 4.995 2.812 5.03 3.44 ;
      RECT 4.99 2.755 4.995 3.44 ;
      RECT 4.985 2.742 4.99 3.44 ;
      RECT 4.975 2.72 4.985 3.44 ;
      RECT 4.965 2.685 4.975 3.44 ;
      RECT 4.955 2.655 4.965 3.44 ;
      RECT 4.945 2.57 4.955 3.083 ;
      RECT 4.952 3.215 4.955 3.44 ;
      RECT 4.95 3.225 4.952 3.44 ;
      RECT 4.94 3.235 4.95 3.435 ;
      RECT 4.935 1.92 4.945 2.315 ;
      RECT 4.94 2.447 4.945 3.058 ;
      RECT 4.935 2.345 4.94 3.041 ;
      RECT 4.925 1.92 4.935 3.017 ;
      RECT 4.92 1.92 4.925 2.988 ;
      RECT 4.915 1.92 4.92 2.978 ;
      RECT 4.895 1.92 4.915 2.94 ;
      RECT 4.89 1.92 4.895 2.898 ;
      RECT 4.885 1.92 4.89 2.878 ;
      RECT 4.855 1.92 4.885 2.828 ;
      RECT 4.845 1.92 4.855 2.775 ;
      RECT 4.84 1.92 4.845 2.748 ;
      RECT 4.835 1.92 4.84 2.733 ;
      RECT 4.825 1.92 4.835 2.71 ;
      RECT 4.815 1.92 4.825 2.685 ;
      RECT 4.81 1.92 4.815 2.625 ;
      RECT 4.8 1.92 4.81 2.563 ;
      RECT 4.795 1.92 4.8 2.483 ;
      RECT 4.79 1.92 4.795 2.448 ;
      RECT 4.785 1.92 4.79 2.423 ;
      RECT 4.78 1.92 4.785 2.408 ;
      RECT 4.775 1.92 4.78 2.378 ;
      RECT 4.77 1.92 4.775 2.355 ;
      RECT 4.765 1.92 4.77 2.328 ;
      RECT 4.735 1.92 4.75 2.315 ;
      RECT 3.89 3.455 4.075 3.665 ;
      RECT 3.88 3.46 4.09 3.658 ;
      RECT 3.88 3.46 4.11 3.63 ;
      RECT 3.88 3.46 4.125 3.609 ;
      RECT 3.88 3.46 4.14 3.607 ;
      RECT 3.88 3.46 4.15 3.606 ;
      RECT 3.88 3.46 4.18 3.603 ;
      RECT 4.53 3.305 4.79 3.565 ;
      RECT 4.49 3.352 4.79 3.548 ;
      RECT 4.481 3.36 4.49 3.551 ;
      RECT 4.075 3.453 4.79 3.548 ;
      RECT 4.395 3.378 4.481 3.558 ;
      RECT 4.09 3.45 4.79 3.548 ;
      RECT 4.336 3.4 4.395 3.57 ;
      RECT 4.11 3.446 4.79 3.548 ;
      RECT 4.25 3.412 4.336 3.581 ;
      RECT 4.125 3.442 4.79 3.548 ;
      RECT 4.195 3.425 4.25 3.593 ;
      RECT 4.14 3.44 4.79 3.548 ;
      RECT 4.18 3.431 4.195 3.599 ;
      RECT 4.15 3.436 4.79 3.548 ;
      RECT 4.295 2.96 4.555 3.22 ;
      RECT 4.295 2.98 4.665 3.19 ;
      RECT 4.295 2.985 4.675 3.185 ;
      RECT 4.486 2.399 4.565 2.63 ;
      RECT 4.4 2.402 4.615 2.625 ;
      RECT 4.395 2.402 4.615 2.62 ;
      RECT 4.395 2.407 4.625 2.618 ;
      RECT 4.37 2.407 4.625 2.615 ;
      RECT 4.37 2.415 4.635 2.613 ;
      RECT 4.25 2.35 4.51 2.61 ;
      RECT 4.25 2.397 4.56 2.61 ;
      RECT 3.505 2.97 3.51 3.23 ;
      RECT 3.335 2.74 3.34 3.23 ;
      RECT 3.22 2.98 3.225 3.205 ;
      RECT 3.93 2.075 3.935 2.285 ;
      RECT 3.935 2.08 3.95 2.28 ;
      RECT 3.87 2.075 3.93 2.293 ;
      RECT 3.855 2.075 3.87 2.303 ;
      RECT 3.805 2.075 3.855 2.32 ;
      RECT 3.785 2.075 3.805 2.343 ;
      RECT 3.77 2.075 3.785 2.355 ;
      RECT 3.75 2.075 3.77 2.365 ;
      RECT 3.74 2.08 3.75 2.374 ;
      RECT 3.735 2.09 3.74 2.379 ;
      RECT 3.73 2.102 3.735 2.383 ;
      RECT 3.72 2.125 3.73 2.388 ;
      RECT 3.715 2.14 3.72 2.392 ;
      RECT 3.71 2.157 3.715 2.395 ;
      RECT 3.705 2.165 3.71 2.398 ;
      RECT 3.695 2.17 3.705 2.402 ;
      RECT 3.69 2.177 3.695 2.407 ;
      RECT 3.68 2.182 3.69 2.411 ;
      RECT 3.655 2.194 3.68 2.422 ;
      RECT 3.635 2.211 3.655 2.438 ;
      RECT 3.61 2.228 3.635 2.46 ;
      RECT 3.575 2.251 3.61 2.518 ;
      RECT 3.555 2.273 3.575 2.58 ;
      RECT 3.55 2.283 3.555 2.615 ;
      RECT 3.54 2.29 3.55 2.653 ;
      RECT 3.535 2.297 3.54 2.673 ;
      RECT 3.53 2.308 3.535 2.71 ;
      RECT 3.525 2.316 3.53 2.775 ;
      RECT 3.515 2.327 3.525 2.828 ;
      RECT 3.51 2.345 3.515 2.898 ;
      RECT 3.505 2.355 3.51 2.935 ;
      RECT 3.5 2.365 3.505 3.23 ;
      RECT 3.495 2.377 3.5 3.23 ;
      RECT 3.49 2.387 3.495 3.23 ;
      RECT 3.48 2.397 3.49 3.23 ;
      RECT 3.47 2.42 3.48 3.23 ;
      RECT 3.455 2.455 3.47 3.23 ;
      RECT 3.415 2.517 3.455 3.23 ;
      RECT 3.41 2.57 3.415 3.23 ;
      RECT 3.385 2.605 3.41 3.23 ;
      RECT 3.37 2.65 3.385 3.23 ;
      RECT 3.365 2.672 3.37 3.23 ;
      RECT 3.355 2.685 3.365 3.23 ;
      RECT 3.345 2.71 3.355 3.23 ;
      RECT 3.34 2.732 3.345 3.23 ;
      RECT 3.315 2.77 3.335 3.23 ;
      RECT 3.275 2.827 3.315 3.23 ;
      RECT 3.27 2.877 3.275 3.23 ;
      RECT 3.265 2.895 3.27 3.23 ;
      RECT 3.26 2.907 3.265 3.23 ;
      RECT 3.25 2.925 3.26 3.23 ;
      RECT 3.24 2.945 3.25 3.205 ;
      RECT 3.235 2.962 3.24 3.205 ;
      RECT 3.225 2.975 3.235 3.205 ;
      RECT 3.195 2.985 3.22 3.205 ;
      RECT 3.185 2.992 3.195 3.205 ;
      RECT 3.17 3.002 3.185 3.2 ;
      RECT 1.98 6.655 2.27 6.885 ;
      RECT 1.81 6.685 2.27 6.855 ;
      RECT 1.55 7.765 1.84 7.995 ;
      RECT 1.61 7.025 1.78 7.995 ;
      RECT 1.52 7.025 1.87 7.315 ;
      RECT 1.145 6.285 1.495 6.575 ;
      RECT 1.005 6.315 1.495 6.485 ;
      RECT 76.06 2.85 76.43 3.22 ;
      RECT 60.275 2.85 60.645 3.22 ;
      RECT 44.49 2.85 44.86 3.22 ;
      RECT 28.715 2.85 29.085 3.22 ;
      RECT 12.935 2.85 13.305 3.22 ;
    LAYER mcon ;
      RECT 81.23 6.32 81.4 6.49 ;
      RECT 81.235 6.315 81.405 6.485 ;
      RECT 65.445 6.32 65.615 6.49 ;
      RECT 65.45 6.315 65.62 6.485 ;
      RECT 49.66 6.32 49.83 6.49 ;
      RECT 49.665 6.315 49.835 6.485 ;
      RECT 33.885 6.32 34.055 6.49 ;
      RECT 33.89 6.315 34.06 6.485 ;
      RECT 18.105 6.32 18.275 6.49 ;
      RECT 18.11 6.315 18.28 6.485 ;
      RECT 0.355 8.64 0.525 8.81 ;
      RECT 0.31 8.605 0.48 8.775 ;
      RECT 81.23 7.8 81.4 7.97 ;
      RECT 80.88 0.1 81.05 0.27 ;
      RECT 80.88 4.16 81.05 4.33 ;
      RECT 80.88 4.55 81.05 4.72 ;
      RECT 80.88 8.61 81.05 8.78 ;
      RECT 80.86 2.76 81.03 2.93 ;
      RECT 80.86 5.95 81.03 6.12 ;
      RECT 80.24 0.91 80.41 1.08 ;
      RECT 80.24 2.39 80.41 2.56 ;
      RECT 80.24 6.32 80.41 6.49 ;
      RECT 80.24 7.8 80.41 7.97 ;
      RECT 79.89 0.1 80.06 0.27 ;
      RECT 79.89 4.16 80.06 4.33 ;
      RECT 79.89 4.55 80.06 4.72 ;
      RECT 79.89 8.61 80.06 8.78 ;
      RECT 79.87 2.76 80.04 2.93 ;
      RECT 79.87 5.95 80.04 6.12 ;
      RECT 79.19 0.105 79.36 0.275 ;
      RECT 79.19 4.165 79.36 4.335 ;
      RECT 79.19 4.545 79.36 4.715 ;
      RECT 79.19 8.605 79.36 8.775 ;
      RECT 78.88 2.025 79.05 2.195 ;
      RECT 78.88 6.685 79.05 6.855 ;
      RECT 78.51 0.105 78.68 0.275 ;
      RECT 78.51 8.605 78.68 8.775 ;
      RECT 78.45 0.915 78.62 1.085 ;
      RECT 78.45 1.655 78.62 1.825 ;
      RECT 78.45 7.055 78.62 7.225 ;
      RECT 78.45 7.795 78.62 7.965 ;
      RECT 78.075 2.395 78.245 2.565 ;
      RECT 78.075 6.315 78.245 6.485 ;
      RECT 77.83 0.105 78 0.275 ;
      RECT 77.83 8.605 78 8.775 ;
      RECT 77.15 0.105 77.32 0.275 ;
      RECT 77.15 8.605 77.32 8.775 ;
      RECT 75.525 1.415 75.695 1.585 ;
      RECT 75.525 4.135 75.695 4.305 ;
      RECT 75.155 2.875 75.325 3.045 ;
      RECT 75.065 1.415 75.235 1.585 ;
      RECT 75.065 4.135 75.235 4.305 ;
      RECT 74.835 2.045 75.005 2.215 ;
      RECT 74.69 2.485 74.86 2.655 ;
      RECT 74.605 1.415 74.775 1.585 ;
      RECT 74.605 4.135 74.775 4.305 ;
      RECT 74.41 4.545 74.58 4.715 ;
      RECT 74.41 8.605 74.58 8.775 ;
      RECT 74.145 1.415 74.315 1.585 ;
      RECT 74.145 4.135 74.315 4.305 ;
      RECT 74.1 6.685 74.27 6.855 ;
      RECT 74.08 2.525 74.25 2.695 ;
      RECT 73.735 2.16 73.905 2.33 ;
      RECT 73.73 8.605 73.9 8.775 ;
      RECT 73.725 3.52 73.895 3.69 ;
      RECT 73.685 1.415 73.855 1.585 ;
      RECT 73.685 4.135 73.855 4.305 ;
      RECT 73.67 7.055 73.84 7.225 ;
      RECT 73.67 7.795 73.84 7.965 ;
      RECT 73.31 2.76 73.48 2.93 ;
      RECT 73.295 6.315 73.465 6.485 ;
      RECT 73.225 1.415 73.395 1.585 ;
      RECT 73.225 4.135 73.395 4.305 ;
      RECT 73.05 8.605 73.22 8.775 ;
      RECT 72.96 2.235 73.13 2.405 ;
      RECT 72.78 3.55 72.95 3.72 ;
      RECT 72.765 1.415 72.935 1.585 ;
      RECT 72.765 4.135 72.935 4.305 ;
      RECT 72.5 2.865 72.67 3.035 ;
      RECT 72.37 8.605 72.54 8.775 ;
      RECT 72.305 1.415 72.475 1.585 ;
      RECT 72.305 4.135 72.475 4.305 ;
      RECT 72.18 2.49 72.35 2.66 ;
      RECT 71.845 1.415 72.015 1.585 ;
      RECT 71.845 4.135 72.015 4.305 ;
      RECT 71.49 1.97 71.66 2.14 ;
      RECT 71.415 2.44 71.585 2.61 ;
      RECT 71.385 1.415 71.555 1.585 ;
      RECT 71.385 4.135 71.555 4.305 ;
      RECT 70.925 1.415 71.095 1.585 ;
      RECT 70.925 4.135 71.095 4.305 ;
      RECT 70.565 2.165 70.735 2.335 ;
      RECT 70.465 1.415 70.635 1.585 ;
      RECT 70.465 4.135 70.635 4.305 ;
      RECT 70.225 3.36 70.395 3.53 ;
      RECT 70.19 2.695 70.36 2.865 ;
      RECT 70.005 1.415 70.175 1.585 ;
      RECT 70.005 4.135 70.175 4.305 ;
      RECT 69.58 2.55 69.75 2.72 ;
      RECT 69.545 1.415 69.715 1.585 ;
      RECT 69.545 4.135 69.715 4.305 ;
      RECT 69.51 3.25 69.68 3.42 ;
      RECT 69.45 2.085 69.62 2.255 ;
      RECT 69.085 1.415 69.255 1.585 ;
      RECT 69.085 4.135 69.255 4.305 ;
      RECT 68.81 3 68.98 3.17 ;
      RECT 68.625 1.415 68.795 1.585 ;
      RECT 68.625 4.135 68.795 4.305 ;
      RECT 68.305 2.505 68.475 2.675 ;
      RECT 68.165 1.415 68.335 1.585 ;
      RECT 68.165 4.135 68.335 4.305 ;
      RECT 68.085 3.25 68.255 3.42 ;
      RECT 67.88 2.13 68.05 2.3 ;
      RECT 67.705 1.415 67.875 1.585 ;
      RECT 67.705 4.135 67.875 4.305 ;
      RECT 67.61 3 67.78 3.17 ;
      RECT 67.57 2.43 67.74 2.6 ;
      RECT 67.245 1.415 67.415 1.585 ;
      RECT 67.245 4.135 67.415 4.305 ;
      RECT 67.025 3.475 67.195 3.645 ;
      RECT 66.885 2.095 67.055 2.265 ;
      RECT 66.785 1.415 66.955 1.585 ;
      RECT 66.785 4.135 66.955 4.305 ;
      RECT 66.325 1.415 66.495 1.585 ;
      RECT 66.325 4.135 66.495 4.305 ;
      RECT 66.315 3.015 66.485 3.185 ;
      RECT 65.445 7.8 65.615 7.97 ;
      RECT 65.095 0.1 65.265 0.27 ;
      RECT 65.095 4.16 65.265 4.33 ;
      RECT 65.095 4.55 65.265 4.72 ;
      RECT 65.095 8.61 65.265 8.78 ;
      RECT 65.075 2.76 65.245 2.93 ;
      RECT 65.075 5.95 65.245 6.12 ;
      RECT 64.455 0.91 64.625 1.08 ;
      RECT 64.455 2.39 64.625 2.56 ;
      RECT 64.455 6.32 64.625 6.49 ;
      RECT 64.455 7.8 64.625 7.97 ;
      RECT 64.105 0.1 64.275 0.27 ;
      RECT 64.105 4.16 64.275 4.33 ;
      RECT 64.105 4.55 64.275 4.72 ;
      RECT 64.105 8.61 64.275 8.78 ;
      RECT 64.085 2.76 64.255 2.93 ;
      RECT 64.085 5.95 64.255 6.12 ;
      RECT 63.405 0.105 63.575 0.275 ;
      RECT 63.405 4.165 63.575 4.335 ;
      RECT 63.405 4.545 63.575 4.715 ;
      RECT 63.405 8.605 63.575 8.775 ;
      RECT 63.095 2.025 63.265 2.195 ;
      RECT 63.095 6.685 63.265 6.855 ;
      RECT 62.725 0.105 62.895 0.275 ;
      RECT 62.725 8.605 62.895 8.775 ;
      RECT 62.665 0.915 62.835 1.085 ;
      RECT 62.665 1.655 62.835 1.825 ;
      RECT 62.665 7.055 62.835 7.225 ;
      RECT 62.665 7.795 62.835 7.965 ;
      RECT 62.29 2.395 62.46 2.565 ;
      RECT 62.29 6.315 62.46 6.485 ;
      RECT 62.045 0.105 62.215 0.275 ;
      RECT 62.045 8.605 62.215 8.775 ;
      RECT 61.365 0.105 61.535 0.275 ;
      RECT 61.365 8.605 61.535 8.775 ;
      RECT 59.74 1.415 59.91 1.585 ;
      RECT 59.74 4.135 59.91 4.305 ;
      RECT 59.37 2.875 59.54 3.045 ;
      RECT 59.28 1.415 59.45 1.585 ;
      RECT 59.28 4.135 59.45 4.305 ;
      RECT 59.05 2.045 59.22 2.215 ;
      RECT 58.905 2.485 59.075 2.655 ;
      RECT 58.82 1.415 58.99 1.585 ;
      RECT 58.82 4.135 58.99 4.305 ;
      RECT 58.625 4.545 58.795 4.715 ;
      RECT 58.625 8.605 58.795 8.775 ;
      RECT 58.36 1.415 58.53 1.585 ;
      RECT 58.36 4.135 58.53 4.305 ;
      RECT 58.315 6.685 58.485 6.855 ;
      RECT 58.295 2.525 58.465 2.695 ;
      RECT 57.95 2.16 58.12 2.33 ;
      RECT 57.945 8.605 58.115 8.775 ;
      RECT 57.94 3.52 58.11 3.69 ;
      RECT 57.9 1.415 58.07 1.585 ;
      RECT 57.9 4.135 58.07 4.305 ;
      RECT 57.885 7.055 58.055 7.225 ;
      RECT 57.885 7.795 58.055 7.965 ;
      RECT 57.525 2.76 57.695 2.93 ;
      RECT 57.51 6.315 57.68 6.485 ;
      RECT 57.44 1.415 57.61 1.585 ;
      RECT 57.44 4.135 57.61 4.305 ;
      RECT 57.265 8.605 57.435 8.775 ;
      RECT 57.175 2.235 57.345 2.405 ;
      RECT 56.995 3.55 57.165 3.72 ;
      RECT 56.98 1.415 57.15 1.585 ;
      RECT 56.98 4.135 57.15 4.305 ;
      RECT 56.715 2.865 56.885 3.035 ;
      RECT 56.585 8.605 56.755 8.775 ;
      RECT 56.52 1.415 56.69 1.585 ;
      RECT 56.52 4.135 56.69 4.305 ;
      RECT 56.395 2.49 56.565 2.66 ;
      RECT 56.06 1.415 56.23 1.585 ;
      RECT 56.06 4.135 56.23 4.305 ;
      RECT 55.705 1.97 55.875 2.14 ;
      RECT 55.63 2.44 55.8 2.61 ;
      RECT 55.6 1.415 55.77 1.585 ;
      RECT 55.6 4.135 55.77 4.305 ;
      RECT 55.14 1.415 55.31 1.585 ;
      RECT 55.14 4.135 55.31 4.305 ;
      RECT 54.78 2.165 54.95 2.335 ;
      RECT 54.68 1.415 54.85 1.585 ;
      RECT 54.68 4.135 54.85 4.305 ;
      RECT 54.44 3.36 54.61 3.53 ;
      RECT 54.405 2.695 54.575 2.865 ;
      RECT 54.22 1.415 54.39 1.585 ;
      RECT 54.22 4.135 54.39 4.305 ;
      RECT 53.795 2.55 53.965 2.72 ;
      RECT 53.76 1.415 53.93 1.585 ;
      RECT 53.76 4.135 53.93 4.305 ;
      RECT 53.725 3.25 53.895 3.42 ;
      RECT 53.665 2.085 53.835 2.255 ;
      RECT 53.3 1.415 53.47 1.585 ;
      RECT 53.3 4.135 53.47 4.305 ;
      RECT 53.025 3 53.195 3.17 ;
      RECT 52.84 1.415 53.01 1.585 ;
      RECT 52.84 4.135 53.01 4.305 ;
      RECT 52.52 2.505 52.69 2.675 ;
      RECT 52.38 1.415 52.55 1.585 ;
      RECT 52.38 4.135 52.55 4.305 ;
      RECT 52.3 3.25 52.47 3.42 ;
      RECT 52.095 2.13 52.265 2.3 ;
      RECT 51.92 1.415 52.09 1.585 ;
      RECT 51.92 4.135 52.09 4.305 ;
      RECT 51.825 3 51.995 3.17 ;
      RECT 51.785 2.43 51.955 2.6 ;
      RECT 51.46 1.415 51.63 1.585 ;
      RECT 51.46 4.135 51.63 4.305 ;
      RECT 51.24 3.475 51.41 3.645 ;
      RECT 51.1 2.095 51.27 2.265 ;
      RECT 51 1.415 51.17 1.585 ;
      RECT 51 4.135 51.17 4.305 ;
      RECT 50.54 1.415 50.71 1.585 ;
      RECT 50.54 4.135 50.71 4.305 ;
      RECT 50.53 3.015 50.7 3.185 ;
      RECT 49.66 7.8 49.83 7.97 ;
      RECT 49.31 0.1 49.48 0.27 ;
      RECT 49.31 4.16 49.48 4.33 ;
      RECT 49.31 4.55 49.48 4.72 ;
      RECT 49.31 8.61 49.48 8.78 ;
      RECT 49.29 2.76 49.46 2.93 ;
      RECT 49.29 5.95 49.46 6.12 ;
      RECT 48.67 0.91 48.84 1.08 ;
      RECT 48.67 2.39 48.84 2.56 ;
      RECT 48.67 6.32 48.84 6.49 ;
      RECT 48.67 7.8 48.84 7.97 ;
      RECT 48.32 0.1 48.49 0.27 ;
      RECT 48.32 4.16 48.49 4.33 ;
      RECT 48.32 4.55 48.49 4.72 ;
      RECT 48.32 8.61 48.49 8.78 ;
      RECT 48.3 2.76 48.47 2.93 ;
      RECT 48.3 5.95 48.47 6.12 ;
      RECT 47.62 0.105 47.79 0.275 ;
      RECT 47.62 4.165 47.79 4.335 ;
      RECT 47.62 4.545 47.79 4.715 ;
      RECT 47.62 8.605 47.79 8.775 ;
      RECT 47.31 2.025 47.48 2.195 ;
      RECT 47.31 6.685 47.48 6.855 ;
      RECT 46.94 0.105 47.11 0.275 ;
      RECT 46.94 8.605 47.11 8.775 ;
      RECT 46.88 0.915 47.05 1.085 ;
      RECT 46.88 1.655 47.05 1.825 ;
      RECT 46.88 7.055 47.05 7.225 ;
      RECT 46.88 7.795 47.05 7.965 ;
      RECT 46.505 2.395 46.675 2.565 ;
      RECT 46.505 6.315 46.675 6.485 ;
      RECT 46.26 0.105 46.43 0.275 ;
      RECT 46.26 8.605 46.43 8.775 ;
      RECT 45.58 0.105 45.75 0.275 ;
      RECT 45.58 8.605 45.75 8.775 ;
      RECT 43.955 1.415 44.125 1.585 ;
      RECT 43.955 4.135 44.125 4.305 ;
      RECT 43.585 2.875 43.755 3.045 ;
      RECT 43.495 1.415 43.665 1.585 ;
      RECT 43.495 4.135 43.665 4.305 ;
      RECT 43.265 2.045 43.435 2.215 ;
      RECT 43.12 2.485 43.29 2.655 ;
      RECT 43.035 1.415 43.205 1.585 ;
      RECT 43.035 4.135 43.205 4.305 ;
      RECT 42.84 4.545 43.01 4.715 ;
      RECT 42.84 8.605 43.01 8.775 ;
      RECT 42.575 1.415 42.745 1.585 ;
      RECT 42.575 4.135 42.745 4.305 ;
      RECT 42.53 6.685 42.7 6.855 ;
      RECT 42.51 2.525 42.68 2.695 ;
      RECT 42.165 2.16 42.335 2.33 ;
      RECT 42.16 8.605 42.33 8.775 ;
      RECT 42.155 3.52 42.325 3.69 ;
      RECT 42.115 1.415 42.285 1.585 ;
      RECT 42.115 4.135 42.285 4.305 ;
      RECT 42.1 7.055 42.27 7.225 ;
      RECT 42.1 7.795 42.27 7.965 ;
      RECT 41.74 2.76 41.91 2.93 ;
      RECT 41.725 6.315 41.895 6.485 ;
      RECT 41.655 1.415 41.825 1.585 ;
      RECT 41.655 4.135 41.825 4.305 ;
      RECT 41.48 8.605 41.65 8.775 ;
      RECT 41.39 2.235 41.56 2.405 ;
      RECT 41.21 3.55 41.38 3.72 ;
      RECT 41.195 1.415 41.365 1.585 ;
      RECT 41.195 4.135 41.365 4.305 ;
      RECT 40.93 2.865 41.1 3.035 ;
      RECT 40.8 8.605 40.97 8.775 ;
      RECT 40.735 1.415 40.905 1.585 ;
      RECT 40.735 4.135 40.905 4.305 ;
      RECT 40.61 2.49 40.78 2.66 ;
      RECT 40.275 1.415 40.445 1.585 ;
      RECT 40.275 4.135 40.445 4.305 ;
      RECT 39.92 1.97 40.09 2.14 ;
      RECT 39.845 2.44 40.015 2.61 ;
      RECT 39.815 1.415 39.985 1.585 ;
      RECT 39.815 4.135 39.985 4.305 ;
      RECT 39.355 1.415 39.525 1.585 ;
      RECT 39.355 4.135 39.525 4.305 ;
      RECT 38.995 2.165 39.165 2.335 ;
      RECT 38.895 1.415 39.065 1.585 ;
      RECT 38.895 4.135 39.065 4.305 ;
      RECT 38.655 3.36 38.825 3.53 ;
      RECT 38.62 2.695 38.79 2.865 ;
      RECT 38.435 1.415 38.605 1.585 ;
      RECT 38.435 4.135 38.605 4.305 ;
      RECT 38.01 2.55 38.18 2.72 ;
      RECT 37.975 1.415 38.145 1.585 ;
      RECT 37.975 4.135 38.145 4.305 ;
      RECT 37.94 3.25 38.11 3.42 ;
      RECT 37.88 2.085 38.05 2.255 ;
      RECT 37.515 1.415 37.685 1.585 ;
      RECT 37.515 4.135 37.685 4.305 ;
      RECT 37.24 3 37.41 3.17 ;
      RECT 37.055 1.415 37.225 1.585 ;
      RECT 37.055 4.135 37.225 4.305 ;
      RECT 36.735 2.505 36.905 2.675 ;
      RECT 36.595 1.415 36.765 1.585 ;
      RECT 36.595 4.135 36.765 4.305 ;
      RECT 36.515 3.25 36.685 3.42 ;
      RECT 36.31 2.13 36.48 2.3 ;
      RECT 36.135 1.415 36.305 1.585 ;
      RECT 36.135 4.135 36.305 4.305 ;
      RECT 36.04 3 36.21 3.17 ;
      RECT 36 2.43 36.17 2.6 ;
      RECT 35.675 1.415 35.845 1.585 ;
      RECT 35.675 4.135 35.845 4.305 ;
      RECT 35.455 3.475 35.625 3.645 ;
      RECT 35.315 2.095 35.485 2.265 ;
      RECT 35.215 1.415 35.385 1.585 ;
      RECT 35.215 4.135 35.385 4.305 ;
      RECT 34.755 1.415 34.925 1.585 ;
      RECT 34.755 4.135 34.925 4.305 ;
      RECT 34.745 3.015 34.915 3.185 ;
      RECT 33.885 7.8 34.055 7.97 ;
      RECT 33.535 0.1 33.705 0.27 ;
      RECT 33.535 4.16 33.705 4.33 ;
      RECT 33.535 4.55 33.705 4.72 ;
      RECT 33.535 8.61 33.705 8.78 ;
      RECT 33.515 2.76 33.685 2.93 ;
      RECT 33.515 5.95 33.685 6.12 ;
      RECT 32.895 0.91 33.065 1.08 ;
      RECT 32.895 2.39 33.065 2.56 ;
      RECT 32.895 6.32 33.065 6.49 ;
      RECT 32.895 7.8 33.065 7.97 ;
      RECT 32.545 0.1 32.715 0.27 ;
      RECT 32.545 4.16 32.715 4.33 ;
      RECT 32.545 4.55 32.715 4.72 ;
      RECT 32.545 8.61 32.715 8.78 ;
      RECT 32.525 2.76 32.695 2.93 ;
      RECT 32.525 5.95 32.695 6.12 ;
      RECT 31.845 0.105 32.015 0.275 ;
      RECT 31.845 4.165 32.015 4.335 ;
      RECT 31.845 4.545 32.015 4.715 ;
      RECT 31.845 8.605 32.015 8.775 ;
      RECT 31.535 2.025 31.705 2.195 ;
      RECT 31.535 6.685 31.705 6.855 ;
      RECT 31.165 0.105 31.335 0.275 ;
      RECT 31.165 8.605 31.335 8.775 ;
      RECT 31.105 0.915 31.275 1.085 ;
      RECT 31.105 1.655 31.275 1.825 ;
      RECT 31.105 7.055 31.275 7.225 ;
      RECT 31.105 7.795 31.275 7.965 ;
      RECT 30.73 2.395 30.9 2.565 ;
      RECT 30.73 6.315 30.9 6.485 ;
      RECT 30.485 0.105 30.655 0.275 ;
      RECT 30.485 8.605 30.655 8.775 ;
      RECT 29.805 0.105 29.975 0.275 ;
      RECT 29.805 8.605 29.975 8.775 ;
      RECT 28.18 1.415 28.35 1.585 ;
      RECT 28.18 4.135 28.35 4.305 ;
      RECT 27.81 2.875 27.98 3.045 ;
      RECT 27.72 1.415 27.89 1.585 ;
      RECT 27.72 4.135 27.89 4.305 ;
      RECT 27.49 2.045 27.66 2.215 ;
      RECT 27.345 2.485 27.515 2.655 ;
      RECT 27.26 1.415 27.43 1.585 ;
      RECT 27.26 4.135 27.43 4.305 ;
      RECT 27.065 4.545 27.235 4.715 ;
      RECT 27.065 8.605 27.235 8.775 ;
      RECT 26.8 1.415 26.97 1.585 ;
      RECT 26.8 4.135 26.97 4.305 ;
      RECT 26.755 6.685 26.925 6.855 ;
      RECT 26.735 2.525 26.905 2.695 ;
      RECT 26.39 2.16 26.56 2.33 ;
      RECT 26.385 8.605 26.555 8.775 ;
      RECT 26.38 3.52 26.55 3.69 ;
      RECT 26.34 1.415 26.51 1.585 ;
      RECT 26.34 4.135 26.51 4.305 ;
      RECT 26.325 7.055 26.495 7.225 ;
      RECT 26.325 7.795 26.495 7.965 ;
      RECT 25.965 2.76 26.135 2.93 ;
      RECT 25.95 6.315 26.12 6.485 ;
      RECT 25.88 1.415 26.05 1.585 ;
      RECT 25.88 4.135 26.05 4.305 ;
      RECT 25.705 8.605 25.875 8.775 ;
      RECT 25.615 2.235 25.785 2.405 ;
      RECT 25.435 3.55 25.605 3.72 ;
      RECT 25.42 1.415 25.59 1.585 ;
      RECT 25.42 4.135 25.59 4.305 ;
      RECT 25.155 2.865 25.325 3.035 ;
      RECT 25.025 8.605 25.195 8.775 ;
      RECT 24.96 1.415 25.13 1.585 ;
      RECT 24.96 4.135 25.13 4.305 ;
      RECT 24.835 2.49 25.005 2.66 ;
      RECT 24.5 1.415 24.67 1.585 ;
      RECT 24.5 4.135 24.67 4.305 ;
      RECT 24.145 1.97 24.315 2.14 ;
      RECT 24.07 2.44 24.24 2.61 ;
      RECT 24.04 1.415 24.21 1.585 ;
      RECT 24.04 4.135 24.21 4.305 ;
      RECT 23.58 1.415 23.75 1.585 ;
      RECT 23.58 4.135 23.75 4.305 ;
      RECT 23.22 2.165 23.39 2.335 ;
      RECT 23.12 1.415 23.29 1.585 ;
      RECT 23.12 4.135 23.29 4.305 ;
      RECT 22.88 3.36 23.05 3.53 ;
      RECT 22.845 2.695 23.015 2.865 ;
      RECT 22.66 1.415 22.83 1.585 ;
      RECT 22.66 4.135 22.83 4.305 ;
      RECT 22.235 2.55 22.405 2.72 ;
      RECT 22.2 1.415 22.37 1.585 ;
      RECT 22.2 4.135 22.37 4.305 ;
      RECT 22.165 3.25 22.335 3.42 ;
      RECT 22.105 2.085 22.275 2.255 ;
      RECT 21.74 1.415 21.91 1.585 ;
      RECT 21.74 4.135 21.91 4.305 ;
      RECT 21.465 3 21.635 3.17 ;
      RECT 21.28 1.415 21.45 1.585 ;
      RECT 21.28 4.135 21.45 4.305 ;
      RECT 20.96 2.505 21.13 2.675 ;
      RECT 20.82 1.415 20.99 1.585 ;
      RECT 20.82 4.135 20.99 4.305 ;
      RECT 20.74 3.25 20.91 3.42 ;
      RECT 20.535 2.13 20.705 2.3 ;
      RECT 20.36 1.415 20.53 1.585 ;
      RECT 20.36 4.135 20.53 4.305 ;
      RECT 20.265 3 20.435 3.17 ;
      RECT 20.225 2.43 20.395 2.6 ;
      RECT 19.9 1.415 20.07 1.585 ;
      RECT 19.9 4.135 20.07 4.305 ;
      RECT 19.68 3.475 19.85 3.645 ;
      RECT 19.54 2.095 19.71 2.265 ;
      RECT 19.44 1.415 19.61 1.585 ;
      RECT 19.44 4.135 19.61 4.305 ;
      RECT 18.98 1.415 19.15 1.585 ;
      RECT 18.98 4.135 19.15 4.305 ;
      RECT 18.97 3.015 19.14 3.185 ;
      RECT 18.105 7.8 18.275 7.97 ;
      RECT 17.755 0.1 17.925 0.27 ;
      RECT 17.755 4.16 17.925 4.33 ;
      RECT 17.755 4.55 17.925 4.72 ;
      RECT 17.755 8.61 17.925 8.78 ;
      RECT 17.735 2.76 17.905 2.93 ;
      RECT 17.735 5.95 17.905 6.12 ;
      RECT 17.115 0.91 17.285 1.08 ;
      RECT 17.115 2.39 17.285 2.56 ;
      RECT 17.115 6.32 17.285 6.49 ;
      RECT 17.115 7.8 17.285 7.97 ;
      RECT 16.765 0.1 16.935 0.27 ;
      RECT 16.765 4.16 16.935 4.33 ;
      RECT 16.765 4.55 16.935 4.72 ;
      RECT 16.765 8.61 16.935 8.78 ;
      RECT 16.745 2.76 16.915 2.93 ;
      RECT 16.745 5.95 16.915 6.12 ;
      RECT 16.065 0.105 16.235 0.275 ;
      RECT 16.065 4.165 16.235 4.335 ;
      RECT 16.065 4.545 16.235 4.715 ;
      RECT 16.065 8.605 16.235 8.775 ;
      RECT 15.755 2.025 15.925 2.195 ;
      RECT 15.755 6.685 15.925 6.855 ;
      RECT 15.385 0.105 15.555 0.275 ;
      RECT 15.385 8.605 15.555 8.775 ;
      RECT 15.325 0.915 15.495 1.085 ;
      RECT 15.325 1.655 15.495 1.825 ;
      RECT 15.325 7.055 15.495 7.225 ;
      RECT 15.325 7.795 15.495 7.965 ;
      RECT 14.95 2.395 15.12 2.565 ;
      RECT 14.95 6.315 15.12 6.485 ;
      RECT 14.705 0.105 14.875 0.275 ;
      RECT 14.705 8.605 14.875 8.775 ;
      RECT 14.025 0.105 14.195 0.275 ;
      RECT 14.025 8.605 14.195 8.775 ;
      RECT 12.4 1.415 12.57 1.585 ;
      RECT 12.4 4.135 12.57 4.305 ;
      RECT 12.03 2.875 12.2 3.045 ;
      RECT 11.94 1.415 12.11 1.585 ;
      RECT 11.94 4.135 12.11 4.305 ;
      RECT 11.71 2.045 11.88 2.215 ;
      RECT 11.565 2.485 11.735 2.655 ;
      RECT 11.48 1.415 11.65 1.585 ;
      RECT 11.48 4.135 11.65 4.305 ;
      RECT 11.285 4.545 11.455 4.715 ;
      RECT 11.285 8.605 11.455 8.775 ;
      RECT 11.02 1.415 11.19 1.585 ;
      RECT 11.02 4.135 11.19 4.305 ;
      RECT 10.975 6.685 11.145 6.855 ;
      RECT 10.955 2.525 11.125 2.695 ;
      RECT 10.61 2.16 10.78 2.33 ;
      RECT 10.605 8.605 10.775 8.775 ;
      RECT 10.6 3.52 10.77 3.69 ;
      RECT 10.56 1.415 10.73 1.585 ;
      RECT 10.56 4.135 10.73 4.305 ;
      RECT 10.545 7.055 10.715 7.225 ;
      RECT 10.545 7.795 10.715 7.965 ;
      RECT 10.185 2.76 10.355 2.93 ;
      RECT 10.17 6.315 10.34 6.485 ;
      RECT 10.1 1.415 10.27 1.585 ;
      RECT 10.1 4.135 10.27 4.305 ;
      RECT 9.925 8.605 10.095 8.775 ;
      RECT 9.835 2.235 10.005 2.405 ;
      RECT 9.655 3.55 9.825 3.72 ;
      RECT 9.64 1.415 9.81 1.585 ;
      RECT 9.64 4.135 9.81 4.305 ;
      RECT 9.375 2.865 9.545 3.035 ;
      RECT 9.245 8.605 9.415 8.775 ;
      RECT 9.18 1.415 9.35 1.585 ;
      RECT 9.18 4.135 9.35 4.305 ;
      RECT 9.055 2.49 9.225 2.66 ;
      RECT 8.72 1.415 8.89 1.585 ;
      RECT 8.72 4.135 8.89 4.305 ;
      RECT 8.365 1.97 8.535 2.14 ;
      RECT 8.29 2.44 8.46 2.61 ;
      RECT 8.26 1.415 8.43 1.585 ;
      RECT 8.26 4.135 8.43 4.305 ;
      RECT 7.8 1.415 7.97 1.585 ;
      RECT 7.8 4.135 7.97 4.305 ;
      RECT 7.44 2.165 7.61 2.335 ;
      RECT 7.34 1.415 7.51 1.585 ;
      RECT 7.34 4.135 7.51 4.305 ;
      RECT 7.1 3.36 7.27 3.53 ;
      RECT 7.065 2.695 7.235 2.865 ;
      RECT 6.88 1.415 7.05 1.585 ;
      RECT 6.88 4.135 7.05 4.305 ;
      RECT 6.455 2.55 6.625 2.72 ;
      RECT 6.42 1.415 6.59 1.585 ;
      RECT 6.42 4.135 6.59 4.305 ;
      RECT 6.385 3.25 6.555 3.42 ;
      RECT 6.325 2.085 6.495 2.255 ;
      RECT 5.96 1.415 6.13 1.585 ;
      RECT 5.96 4.135 6.13 4.305 ;
      RECT 5.685 3 5.855 3.17 ;
      RECT 5.5 1.415 5.67 1.585 ;
      RECT 5.5 4.135 5.67 4.305 ;
      RECT 5.18 2.505 5.35 2.675 ;
      RECT 5.04 1.415 5.21 1.585 ;
      RECT 5.04 4.135 5.21 4.305 ;
      RECT 4.96 3.25 5.13 3.42 ;
      RECT 4.755 2.13 4.925 2.3 ;
      RECT 4.58 1.415 4.75 1.585 ;
      RECT 4.58 4.135 4.75 4.305 ;
      RECT 4.485 3 4.655 3.17 ;
      RECT 4.445 2.43 4.615 2.6 ;
      RECT 4.12 1.415 4.29 1.585 ;
      RECT 4.12 4.135 4.29 4.305 ;
      RECT 3.9 3.475 4.07 3.645 ;
      RECT 3.76 2.095 3.93 2.265 ;
      RECT 3.66 1.415 3.83 1.585 ;
      RECT 3.66 4.135 3.83 4.305 ;
      RECT 3.2 1.415 3.37 1.585 ;
      RECT 3.2 4.135 3.37 4.305 ;
      RECT 3.19 3.015 3.36 3.185 ;
      RECT 2.35 4.545 2.52 4.715 ;
      RECT 2.35 8.605 2.52 8.775 ;
      RECT 2.04 6.685 2.21 6.855 ;
      RECT 1.67 8.605 1.84 8.775 ;
      RECT 1.61 7.055 1.78 7.225 ;
      RECT 1.61 7.795 1.78 7.965 ;
      RECT 1.235 6.315 1.405 6.485 ;
      RECT 0.99 8.605 1.16 8.775 ;
      RECT 0.94 4.335 1.11 4.505 ;
      RECT 0.885 0.075 1.055 0.245 ;
    LAYER li1 ;
      RECT 74.31 0 74.48 2.085 ;
      RECT 72.35 0 72.52 2.085 ;
      RECT 69.91 0 70.08 2.085 ;
      RECT 68.95 0 69.12 2.085 ;
      RECT 68.43 0 68.6 2.085 ;
      RECT 67.47 0 67.64 2.085 ;
      RECT 66.51 0 66.68 2.085 ;
      RECT 58.525 0 58.695 2.085 ;
      RECT 56.565 0 56.735 2.085 ;
      RECT 54.125 0 54.295 2.085 ;
      RECT 53.165 0 53.335 2.085 ;
      RECT 52.645 0 52.815 2.085 ;
      RECT 51.685 0 51.855 2.085 ;
      RECT 50.725 0 50.895 2.085 ;
      RECT 42.74 0 42.91 2.085 ;
      RECT 40.78 0 40.95 2.085 ;
      RECT 38.34 0 38.51 2.085 ;
      RECT 37.38 0 37.55 2.085 ;
      RECT 36.86 0 37.03 2.085 ;
      RECT 35.9 0 36.07 2.085 ;
      RECT 34.94 0 35.11 2.085 ;
      RECT 26.965 0 27.135 2.085 ;
      RECT 25.005 0 25.175 2.085 ;
      RECT 22.565 0 22.735 2.085 ;
      RECT 21.605 0 21.775 2.085 ;
      RECT 21.085 0 21.255 2.085 ;
      RECT 20.125 0 20.295 2.085 ;
      RECT 19.165 0 19.335 2.085 ;
      RECT 11.185 0 11.355 2.085 ;
      RECT 9.225 0 9.395 2.085 ;
      RECT 6.785 0 6.955 2.085 ;
      RECT 5.825 0 5.995 2.085 ;
      RECT 5.305 0 5.475 2.085 ;
      RECT 4.345 0 4.515 2.085 ;
      RECT 3.385 0 3.555 2.085 ;
      RECT 66.295 0 75.895 1.59 ;
      RECT 50.51 0 60.11 1.59 ;
      RECT 34.725 0 44.325 1.59 ;
      RECT 18.95 0 28.55 1.59 ;
      RECT 3.17 0 12.77 1.59 ;
      RECT 66.18 1.415 76.01 1.585 ;
      RECT 66.295 0 76.01 1.585 ;
      RECT 50.395 1.415 60.225 1.585 ;
      RECT 50.51 0 60.225 1.585 ;
      RECT 34.61 1.415 44.44 1.585 ;
      RECT 34.725 0 44.44 1.585 ;
      RECT 18.835 1.415 28.665 1.585 ;
      RECT 18.95 0 28.665 1.585 ;
      RECT 3.055 1.415 12.885 1.585 ;
      RECT 3.17 0 12.885 1.585 ;
      RECT 77.07 0 77.24 0.935 ;
      RECT 61.285 0 61.455 0.935 ;
      RECT 45.5 0 45.67 0.935 ;
      RECT 29.725 0 29.895 0.935 ;
      RECT 13.945 0 14.115 0.935 ;
      RECT 80.8 0 80.97 0.93 ;
      RECT 79.81 0 79.98 0.93 ;
      RECT 65.015 0 65.185 0.93 ;
      RECT 64.025 0 64.195 0.93 ;
      RECT 49.23 0 49.4 0.93 ;
      RECT 48.24 0 48.41 0.93 ;
      RECT 33.455 0 33.625 0.93 ;
      RECT 32.465 0 32.635 0.93 ;
      RECT 17.675 0 17.845 0.93 ;
      RECT 16.685 0 16.855 0.93 ;
      RECT 0.885 0 1.055 0.365 ;
      RECT 0.585 0 1.395 0.315 ;
      RECT 81.595 0 81.775 0.305 ;
      RECT 65.81 0 79.645 0.305 ;
      RECT 50.025 0 63.86 0.305 ;
      RECT 34.25 0 48.075 0.305 ;
      RECT 18.47 0 32.3 0.305 ;
      RECT 0 0 16.52 0.305 ;
      RECT 0 0 81.775 0.3 ;
      RECT 2.04 4.135 2.21 8.305 ;
      RECT 80.8 3.4 80.97 5.48 ;
      RECT 79.81 3.4 79.98 5.48 ;
      RECT 65.015 3.4 65.185 5.48 ;
      RECT 64.025 3.4 64.195 5.48 ;
      RECT 49.23 3.4 49.4 5.48 ;
      RECT 48.24 3.4 48.41 5.48 ;
      RECT 33.455 3.4 33.625 5.48 ;
      RECT 32.465 3.4 32.635 5.48 ;
      RECT 17.675 3.4 17.845 5.48 ;
      RECT 16.685 3.4 16.855 5.48 ;
      RECT 77.07 3.405 77.24 5.475 ;
      RECT 72.29 4.135 72.46 5.475 ;
      RECT 61.285 3.405 61.455 5.475 ;
      RECT 56.505 4.135 56.675 5.475 ;
      RECT 45.5 3.405 45.67 5.475 ;
      RECT 40.72 4.135 40.89 5.475 ;
      RECT 29.725 3.405 29.895 5.475 ;
      RECT 24.945 4.135 25.115 5.475 ;
      RECT 13.945 3.405 14.115 5.475 ;
      RECT 9.165 4.135 9.335 5.475 ;
      RECT 0.23 4.135 0.4 5.475 ;
      RECT 79.64 4.13 81.62 4.75 ;
      RECT 63.855 4.13 65.835 4.75 ;
      RECT 48.07 4.13 50.05 4.75 ;
      RECT 32.295 4.13 34.275 4.75 ;
      RECT 16.515 4.13 18.495 4.75 ;
      RECT 0 4.135 81.775 4.745 ;
      RECT 75.27 3.635 75.44 4.745 ;
      RECT 74.31 3.635 74.48 4.745 ;
      RECT 71.87 3.635 72.04 4.745 ;
      RECT 70.87 3.635 71.04 4.745 ;
      RECT 69.91 3.635 70.08 4.745 ;
      RECT 67.47 3.635 67.64 4.745 ;
      RECT 59.485 3.635 59.655 4.745 ;
      RECT 58.525 3.635 58.695 4.745 ;
      RECT 56.085 3.635 56.255 4.745 ;
      RECT 55.085 3.635 55.255 4.745 ;
      RECT 54.125 3.635 54.295 4.745 ;
      RECT 51.685 3.635 51.855 4.745 ;
      RECT 43.7 3.635 43.87 4.745 ;
      RECT 42.74 3.635 42.91 4.745 ;
      RECT 40.3 3.635 40.47 4.745 ;
      RECT 39.3 3.635 39.47 4.745 ;
      RECT 38.34 3.635 38.51 4.745 ;
      RECT 35.9 3.635 36.07 4.745 ;
      RECT 27.925 3.635 28.095 4.745 ;
      RECT 26.965 3.635 27.135 4.745 ;
      RECT 24.525 3.635 24.695 4.745 ;
      RECT 23.525 3.635 23.695 4.745 ;
      RECT 22.565 3.635 22.735 4.745 ;
      RECT 20.125 3.635 20.295 4.745 ;
      RECT 12.145 3.635 12.315 4.745 ;
      RECT 11.185 3.635 11.355 4.745 ;
      RECT 8.745 3.635 8.915 4.745 ;
      RECT 7.745 3.635 7.915 4.745 ;
      RECT 6.785 3.635 6.955 4.745 ;
      RECT 4.345 3.635 4.515 4.745 ;
      RECT -0.005 8.58 81.775 8.88 ;
      RECT 81.595 8.575 81.775 8.88 ;
      RECT 80.8 7.95 80.97 8.88 ;
      RECT 79.81 7.95 79.98 8.88 ;
      RECT 65.81 8.575 79.645 8.88 ;
      RECT 65.015 7.95 65.185 8.88 ;
      RECT 64.025 7.95 64.195 8.88 ;
      RECT 50.025 8.575 63.86 8.88 ;
      RECT 49.23 7.95 49.4 8.88 ;
      RECT 48.24 7.95 48.41 8.88 ;
      RECT 34.25 8.575 48.075 8.88 ;
      RECT 33.455 7.95 33.625 8.88 ;
      RECT 32.465 7.95 32.635 8.88 ;
      RECT 18.47 8.575 32.3 8.88 ;
      RECT 17.675 7.95 17.845 8.88 ;
      RECT 16.685 7.95 16.855 8.88 ;
      RECT -0.005 8.575 16.52 8.88 ;
      RECT 77.07 7.945 77.24 8.88 ;
      RECT 72.29 7.945 72.46 8.88 ;
      RECT 61.285 7.945 61.455 8.88 ;
      RECT 56.505 7.945 56.675 8.88 ;
      RECT 45.5 7.945 45.67 8.88 ;
      RECT 40.72 7.945 40.89 8.88 ;
      RECT 29.725 7.945 29.895 8.88 ;
      RECT 24.945 7.945 25.115 8.88 ;
      RECT 13.945 7.945 14.115 8.88 ;
      RECT 9.165 7.945 9.335 8.88 ;
      RECT 0.23 7.945 0.4 8.88 ;
      RECT 81.23 5.02 81.4 6.49 ;
      RECT 81.23 6.315 81.405 6.485 ;
      RECT 80.86 1.74 81.03 2.93 ;
      RECT 80.86 1.74 81.33 1.91 ;
      RECT 80.86 6.97 81.33 7.14 ;
      RECT 80.86 5.95 81.03 7.14 ;
      RECT 79.87 1.74 80.04 2.93 ;
      RECT 79.87 1.74 80.34 1.91 ;
      RECT 79.87 6.97 80.34 7.14 ;
      RECT 79.87 5.95 80.04 7.14 ;
      RECT 78.02 2.635 78.19 3.865 ;
      RECT 78.075 0.855 78.245 2.805 ;
      RECT 78.02 0.575 78.19 1.025 ;
      RECT 78.02 7.855 78.19 8.305 ;
      RECT 78.075 6.075 78.245 8.025 ;
      RECT 78.02 5.015 78.19 6.245 ;
      RECT 77.5 0.575 77.67 3.865 ;
      RECT 77.5 2.075 77.905 2.405 ;
      RECT 77.5 1.235 77.905 1.565 ;
      RECT 77.5 5.015 77.67 8.305 ;
      RECT 77.5 7.315 77.905 7.645 ;
      RECT 77.5 6.475 77.905 6.805 ;
      RECT 74.835 1.975 75.565 2.215 ;
      RECT 75.377 1.77 75.565 2.215 ;
      RECT 75.205 1.782 75.58 2.209 ;
      RECT 75.12 1.797 75.6 2.194 ;
      RECT 75.12 1.812 75.605 2.184 ;
      RECT 75.075 1.832 75.62 2.176 ;
      RECT 75.052 1.867 75.635 2.13 ;
      RECT 74.966 1.89 75.64 2.09 ;
      RECT 74.966 1.908 75.65 2.06 ;
      RECT 74.835 1.977 75.655 2.023 ;
      RECT 74.88 1.92 75.65 2.06 ;
      RECT 74.966 1.872 75.635 2.13 ;
      RECT 75.052 1.841 75.62 2.176 ;
      RECT 75.075 1.822 75.605 2.184 ;
      RECT 75.12 1.795 75.58 2.209 ;
      RECT 75.205 1.777 75.565 2.215 ;
      RECT 75.291 1.771 75.565 2.215 ;
      RECT 75.377 1.766 75.51 2.215 ;
      RECT 75.463 1.761 75.51 2.215 ;
      RECT 75.155 2.659 75.325 3.045 ;
      RECT 75.15 2.659 75.325 3.04 ;
      RECT 75.125 2.659 75.325 3.005 ;
      RECT 75.125 2.687 75.335 2.995 ;
      RECT 75.105 2.687 75.335 2.955 ;
      RECT 75.1 2.687 75.335 2.928 ;
      RECT 75.1 2.705 75.34 2.92 ;
      RECT 75.045 2.705 75.34 2.855 ;
      RECT 75.045 2.722 75.35 2.838 ;
      RECT 75.035 2.722 75.35 2.778 ;
      RECT 75.035 2.739 75.355 2.775 ;
      RECT 75.03 2.575 75.2 2.753 ;
      RECT 75.03 2.609 75.286 2.753 ;
      RECT 75.025 3.375 75.03 3.388 ;
      RECT 75.02 3.27 75.025 3.393 ;
      RECT 74.995 3.13 75.02 3.408 ;
      RECT 74.96 3.081 74.995 3.44 ;
      RECT 74.955 3.049 74.96 3.46 ;
      RECT 74.95 3.04 74.955 3.46 ;
      RECT 74.87 3.005 74.95 3.46 ;
      RECT 74.807 2.975 74.87 3.46 ;
      RECT 74.721 2.963 74.807 3.46 ;
      RECT 74.635 2.949 74.721 3.46 ;
      RECT 74.555 2.936 74.635 3.446 ;
      RECT 74.52 2.928 74.555 3.426 ;
      RECT 74.51 2.925 74.52 3.417 ;
      RECT 74.48 2.92 74.51 3.404 ;
      RECT 74.43 2.895 74.48 3.38 ;
      RECT 74.416 2.869 74.43 3.362 ;
      RECT 74.33 2.829 74.416 3.338 ;
      RECT 74.285 2.777 74.33 3.307 ;
      RECT 74.275 2.752 74.285 3.294 ;
      RECT 74.27 2.533 74.275 2.555 ;
      RECT 74.265 2.735 74.275 3.29 ;
      RECT 74.265 2.531 74.27 2.645 ;
      RECT 74.255 2.527 74.265 3.286 ;
      RECT 74.211 2.525 74.255 3.274 ;
      RECT 74.125 2.525 74.211 3.245 ;
      RECT 74.095 2.525 74.125 3.218 ;
      RECT 74.08 2.525 74.095 3.206 ;
      RECT 74.04 2.537 74.08 3.191 ;
      RECT 74.02 2.556 74.04 3.17 ;
      RECT 74.01 2.566 74.02 3.154 ;
      RECT 74 2.572 74.01 3.143 ;
      RECT 73.98 2.582 74 3.126 ;
      RECT 73.975 2.591 73.98 3.113 ;
      RECT 73.97 2.595 73.975 3.063 ;
      RECT 73.96 2.601 73.97 2.98 ;
      RECT 73.955 2.605 73.96 2.894 ;
      RECT 73.95 2.625 73.955 2.831 ;
      RECT 73.945 2.648 73.95 2.778 ;
      RECT 73.94 2.666 73.945 2.723 ;
      RECT 74.55 2.485 74.72 2.745 ;
      RECT 74.72 2.45 74.765 2.731 ;
      RECT 74.681 2.452 74.77 2.714 ;
      RECT 74.57 2.469 74.856 2.685 ;
      RECT 74.57 2.484 74.86 2.657 ;
      RECT 74.57 2.465 74.77 2.714 ;
      RECT 74.595 2.453 74.72 2.745 ;
      RECT 74.681 2.451 74.765 2.731 ;
      RECT 73.735 1.84 73.905 2.33 ;
      RECT 73.735 1.84 73.94 2.31 ;
      RECT 73.87 1.76 73.98 2.27 ;
      RECT 73.851 1.764 74 2.24 ;
      RECT 73.765 1.772 74.02 2.223 ;
      RECT 73.765 1.778 74.025 2.213 ;
      RECT 73.765 1.787 74.045 2.201 ;
      RECT 73.74 1.812 74.075 2.179 ;
      RECT 73.74 1.832 74.08 2.159 ;
      RECT 73.735 1.845 74.09 2.139 ;
      RECT 73.735 1.912 74.095 2.12 ;
      RECT 73.735 2.045 74.1 2.107 ;
      RECT 73.73 1.85 74.09 1.94 ;
      RECT 73.74 1.807 74.045 2.201 ;
      RECT 73.851 1.762 73.98 2.27 ;
      RECT 73.725 3.515 74.025 3.77 ;
      RECT 73.81 3.481 74.025 3.77 ;
      RECT 73.81 3.484 74.03 3.63 ;
      RECT 73.745 3.505 74.03 3.63 ;
      RECT 73.78 3.495 74.025 3.77 ;
      RECT 73.775 3.5 74.03 3.63 ;
      RECT 73.81 3.479 74.011 3.77 ;
      RECT 73.896 3.47 74.011 3.77 ;
      RECT 73.896 3.464 73.925 3.77 ;
      RECT 73.385 3.105 73.395 3.595 ;
      RECT 73.045 3.04 73.055 3.34 ;
      RECT 73.56 3.212 73.565 3.431 ;
      RECT 73.55 3.192 73.56 3.448 ;
      RECT 73.54 3.172 73.55 3.478 ;
      RECT 73.535 3.162 73.54 3.493 ;
      RECT 73.53 3.158 73.535 3.498 ;
      RECT 73.515 3.15 73.53 3.505 ;
      RECT 73.475 3.13 73.515 3.53 ;
      RECT 73.45 3.112 73.475 3.563 ;
      RECT 73.445 3.11 73.45 3.576 ;
      RECT 73.425 3.107 73.445 3.58 ;
      RECT 73.395 3.105 73.425 3.59 ;
      RECT 73.325 3.107 73.385 3.591 ;
      RECT 73.305 3.107 73.325 3.585 ;
      RECT 73.28 3.105 73.305 3.582 ;
      RECT 73.245 3.1 73.28 3.578 ;
      RECT 73.225 3.094 73.245 3.565 ;
      RECT 73.215 3.091 73.225 3.553 ;
      RECT 73.195 3.088 73.215 3.538 ;
      RECT 73.175 3.084 73.195 3.52 ;
      RECT 73.17 3.081 73.175 3.51 ;
      RECT 73.165 3.08 73.17 3.508 ;
      RECT 73.155 3.077 73.165 3.5 ;
      RECT 73.145 3.071 73.155 3.483 ;
      RECT 73.135 3.065 73.145 3.465 ;
      RECT 73.125 3.059 73.135 3.453 ;
      RECT 73.115 3.053 73.125 3.433 ;
      RECT 73.11 3.049 73.115 3.418 ;
      RECT 73.105 3.047 73.11 3.41 ;
      RECT 73.1 3.045 73.105 3.403 ;
      RECT 73.095 3.043 73.1 3.393 ;
      RECT 73.09 3.041 73.095 3.387 ;
      RECT 73.08 3.04 73.09 3.377 ;
      RECT 73.07 3.04 73.08 3.368 ;
      RECT 73.055 3.04 73.07 3.353 ;
      RECT 73.015 3.04 73.045 3.337 ;
      RECT 72.995 3.042 73.015 3.332 ;
      RECT 72.99 3.047 72.995 3.33 ;
      RECT 72.96 3.055 72.99 3.328 ;
      RECT 72.93 3.07 72.96 3.327 ;
      RECT 72.885 3.092 72.93 3.332 ;
      RECT 72.88 3.107 72.885 3.336 ;
      RECT 72.865 3.112 72.88 3.338 ;
      RECT 72.86 3.116 72.865 3.34 ;
      RECT 72.8 3.139 72.86 3.349 ;
      RECT 72.78 3.165 72.8 3.362 ;
      RECT 72.77 3.172 72.78 3.366 ;
      RECT 72.755 3.179 72.77 3.369 ;
      RECT 72.735 3.189 72.755 3.372 ;
      RECT 72.73 3.197 72.735 3.375 ;
      RECT 72.685 3.202 72.73 3.382 ;
      RECT 72.675 3.205 72.685 3.389 ;
      RECT 72.665 3.205 72.675 3.393 ;
      RECT 72.63 3.207 72.665 3.405 ;
      RECT 72.61 3.21 72.63 3.418 ;
      RECT 72.57 3.213 72.61 3.429 ;
      RECT 72.555 3.215 72.57 3.442 ;
      RECT 72.545 3.215 72.555 3.447 ;
      RECT 72.52 3.216 72.545 3.455 ;
      RECT 72.51 3.218 72.52 3.46 ;
      RECT 72.505 3.219 72.51 3.463 ;
      RECT 72.48 3.217 72.505 3.466 ;
      RECT 72.465 3.215 72.48 3.467 ;
      RECT 72.445 3.212 72.465 3.469 ;
      RECT 72.425 3.207 72.445 3.469 ;
      RECT 72.365 3.202 72.425 3.466 ;
      RECT 72.33 3.177 72.365 3.462 ;
      RECT 72.32 3.154 72.33 3.46 ;
      RECT 72.29 3.131 72.32 3.46 ;
      RECT 72.28 3.11 72.29 3.46 ;
      RECT 72.255 3.092 72.28 3.458 ;
      RECT 72.24 3.07 72.255 3.455 ;
      RECT 72.225 3.052 72.24 3.453 ;
      RECT 72.205 3.042 72.225 3.451 ;
      RECT 72.19 3.037 72.205 3.45 ;
      RECT 72.175 3.035 72.19 3.449 ;
      RECT 72.145 3.036 72.175 3.447 ;
      RECT 72.125 3.039 72.145 3.445 ;
      RECT 72.068 3.043 72.125 3.445 ;
      RECT 71.982 3.052 72.068 3.445 ;
      RECT 71.896 3.063 71.982 3.445 ;
      RECT 71.81 3.074 71.896 3.445 ;
      RECT 71.79 3.081 71.81 3.453 ;
      RECT 71.78 3.084 71.79 3.46 ;
      RECT 71.715 3.089 71.78 3.478 ;
      RECT 71.685 3.096 71.715 3.503 ;
      RECT 71.675 3.099 71.685 3.51 ;
      RECT 71.63 3.103 71.675 3.515 ;
      RECT 71.6 3.108 71.63 3.52 ;
      RECT 71.599 3.11 71.6 3.52 ;
      RECT 71.513 3.116 71.599 3.52 ;
      RECT 71.427 3.127 71.513 3.52 ;
      RECT 71.341 3.139 71.427 3.52 ;
      RECT 71.255 3.15 71.341 3.52 ;
      RECT 71.24 3.157 71.255 3.515 ;
      RECT 71.235 3.159 71.24 3.509 ;
      RECT 71.215 3.17 71.235 3.504 ;
      RECT 71.205 3.188 71.215 3.498 ;
      RECT 71.2 3.2 71.205 3.298 ;
      RECT 73.495 1.953 73.515 2.04 ;
      RECT 73.49 1.888 73.495 2.072 ;
      RECT 73.48 1.855 73.49 2.077 ;
      RECT 73.475 1.835 73.48 2.083 ;
      RECT 73.445 1.835 73.475 2.1 ;
      RECT 73.396 1.835 73.445 2.136 ;
      RECT 73.31 1.835 73.396 2.194 ;
      RECT 73.281 1.845 73.31 2.243 ;
      RECT 73.195 1.887 73.281 2.296 ;
      RECT 73.175 1.925 73.195 2.343 ;
      RECT 73.15 1.942 73.175 2.363 ;
      RECT 73.14 1.956 73.15 2.383 ;
      RECT 73.135 1.962 73.14 2.393 ;
      RECT 73.13 1.966 73.135 2.4 ;
      RECT 73.08 1.986 73.13 2.405 ;
      RECT 73.015 2.03 73.08 2.405 ;
      RECT 72.99 2.08 73.015 2.405 ;
      RECT 72.98 2.11 72.99 2.405 ;
      RECT 72.975 2.137 72.98 2.405 ;
      RECT 72.97 2.155 72.975 2.405 ;
      RECT 72.96 2.197 72.97 2.405 ;
      RECT 73.31 2.755 73.48 2.93 ;
      RECT 73.25 2.583 73.31 2.918 ;
      RECT 73.24 2.576 73.25 2.901 ;
      RECT 73.195 2.755 73.48 2.881 ;
      RECT 73.176 2.755 73.48 2.859 ;
      RECT 73.09 2.755 73.48 2.824 ;
      RECT 73.07 2.575 73.24 2.78 ;
      RECT 73.07 2.722 73.475 2.78 ;
      RECT 73.07 2.67 73.45 2.78 ;
      RECT 73.07 2.625 73.415 2.78 ;
      RECT 73.07 2.607 73.38 2.78 ;
      RECT 73.07 2.597 73.375 2.78 ;
      RECT 73.24 7.855 73.41 8.305 ;
      RECT 73.295 6.075 73.465 8.025 ;
      RECT 73.24 5.015 73.41 6.245 ;
      RECT 72.72 5.015 72.89 8.305 ;
      RECT 72.72 7.315 73.125 7.645 ;
      RECT 72.72 6.475 73.125 6.805 ;
      RECT 72.79 3.555 72.98 3.78 ;
      RECT 72.78 3.556 72.985 3.775 ;
      RECT 72.78 3.558 72.995 3.755 ;
      RECT 72.78 3.562 73 3.74 ;
      RECT 72.78 3.549 72.95 3.775 ;
      RECT 72.78 3.552 72.975 3.775 ;
      RECT 72.79 3.548 72.95 3.78 ;
      RECT 72.876 3.546 72.95 3.78 ;
      RECT 72.5 2.797 72.67 3.035 ;
      RECT 72.5 2.797 72.756 2.949 ;
      RECT 72.5 2.797 72.76 2.859 ;
      RECT 72.55 2.57 72.77 2.838 ;
      RECT 72.545 2.587 72.775 2.811 ;
      RECT 72.51 2.745 72.775 2.811 ;
      RECT 72.53 2.595 72.67 3.035 ;
      RECT 72.52 2.677 72.78 2.794 ;
      RECT 72.515 2.725 72.78 2.794 ;
      RECT 72.52 2.635 72.775 2.811 ;
      RECT 72.545 2.572 72.77 2.838 ;
      RECT 72.11 2.547 72.28 2.745 ;
      RECT 72.11 2.547 72.325 2.72 ;
      RECT 72.18 2.49 72.35 2.678 ;
      RECT 72.155 2.505 72.35 2.678 ;
      RECT 71.77 2.551 71.8 2.745 ;
      RECT 71.765 2.523 71.77 2.745 ;
      RECT 71.735 2.497 71.765 2.747 ;
      RECT 71.71 2.455 71.735 2.75 ;
      RECT 71.7 2.427 71.71 2.752 ;
      RECT 71.665 2.407 71.7 2.754 ;
      RECT 71.6 2.392 71.665 2.76 ;
      RECT 71.55 2.39 71.6 2.766 ;
      RECT 71.527 2.392 71.55 2.771 ;
      RECT 71.441 2.403 71.527 2.777 ;
      RECT 71.355 2.421 71.441 2.787 ;
      RECT 71.34 2.432 71.355 2.793 ;
      RECT 71.27 2.455 71.34 2.799 ;
      RECT 71.215 2.487 71.27 2.807 ;
      RECT 71.175 2.51 71.215 2.813 ;
      RECT 71.161 2.523 71.175 2.816 ;
      RECT 71.075 2.545 71.161 2.822 ;
      RECT 71.06 2.57 71.075 2.828 ;
      RECT 71.02 2.585 71.06 2.832 ;
      RECT 70.97 2.6 71.02 2.837 ;
      RECT 70.945 2.607 70.97 2.841 ;
      RECT 70.885 2.602 70.945 2.845 ;
      RECT 70.87 2.593 70.885 2.849 ;
      RECT 70.8 2.583 70.87 2.845 ;
      RECT 70.775 2.575 70.795 2.835 ;
      RECT 70.716 2.575 70.775 2.813 ;
      RECT 70.63 2.575 70.716 2.77 ;
      RECT 70.795 2.575 70.8 2.84 ;
      RECT 71.49 1.806 71.66 2.14 ;
      RECT 71.46 1.806 71.66 2.135 ;
      RECT 71.4 1.773 71.46 2.123 ;
      RECT 71.4 1.829 71.67 2.118 ;
      RECT 71.375 1.829 71.67 2.112 ;
      RECT 71.37 1.77 71.4 2.109 ;
      RECT 71.355 1.776 71.49 2.107 ;
      RECT 71.35 1.784 71.575 2.095 ;
      RECT 71.35 1.836 71.685 2.048 ;
      RECT 71.335 1.792 71.575 2.043 ;
      RECT 71.335 1.862 71.695 1.984 ;
      RECT 71.305 1.812 71.66 1.945 ;
      RECT 71.305 1.902 71.705 1.941 ;
      RECT 71.355 1.781 71.575 2.107 ;
      RECT 70.695 2.111 70.75 2.375 ;
      RECT 70.695 2.111 70.815 2.374 ;
      RECT 70.695 2.111 70.84 2.373 ;
      RECT 70.695 2.111 70.905 2.372 ;
      RECT 70.84 2.077 70.92 2.371 ;
      RECT 70.655 2.121 71.065 2.37 ;
      RECT 70.695 2.118 71.065 2.37 ;
      RECT 70.655 2.126 71.07 2.363 ;
      RECT 70.64 2.128 71.07 2.362 ;
      RECT 70.64 2.135 71.075 2.358 ;
      RECT 70.62 2.134 71.07 2.354 ;
      RECT 70.62 2.142 71.08 2.353 ;
      RECT 70.615 2.139 71.075 2.349 ;
      RECT 70.615 2.152 71.09 2.348 ;
      RECT 70.6 2.142 71.08 2.347 ;
      RECT 70.565 2.155 71.09 2.34 ;
      RECT 70.75 2.11 71.06 2.37 ;
      RECT 70.75 2.095 71.01 2.37 ;
      RECT 70.815 2.082 70.945 2.37 ;
      RECT 70.36 3.171 70.375 3.564 ;
      RECT 70.325 3.176 70.375 3.563 ;
      RECT 70.36 3.175 70.42 3.562 ;
      RECT 70.305 3.186 70.42 3.561 ;
      RECT 70.32 3.182 70.42 3.561 ;
      RECT 70.285 3.192 70.495 3.558 ;
      RECT 70.285 3.211 70.54 3.556 ;
      RECT 70.285 3.218 70.545 3.553 ;
      RECT 70.27 3.195 70.495 3.55 ;
      RECT 70.25 3.2 70.495 3.543 ;
      RECT 70.245 3.204 70.495 3.539 ;
      RECT 70.245 3.221 70.555 3.538 ;
      RECT 70.225 3.215 70.54 3.534 ;
      RECT 70.225 3.224 70.56 3.528 ;
      RECT 70.22 3.23 70.56 3.3 ;
      RECT 70.285 3.19 70.42 3.558 ;
      RECT 70.16 2.553 70.36 2.865 ;
      RECT 70.235 2.531 70.36 2.865 ;
      RECT 70.175 2.55 70.365 2.85 ;
      RECT 70.145 2.561 70.365 2.848 ;
      RECT 70.16 2.556 70.37 2.814 ;
      RECT 70.145 2.66 70.375 2.781 ;
      RECT 70.175 2.532 70.36 2.865 ;
      RECT 70.235 2.51 70.335 2.865 ;
      RECT 70.26 2.507 70.335 2.865 ;
      RECT 70.26 2.502 70.28 2.865 ;
      RECT 69.665 2.57 69.84 2.745 ;
      RECT 69.66 2.57 69.84 2.743 ;
      RECT 69.635 2.57 69.84 2.738 ;
      RECT 69.58 2.55 69.75 2.728 ;
      RECT 69.58 2.557 69.815 2.728 ;
      RECT 69.665 3.237 69.68 3.42 ;
      RECT 69.655 3.215 69.665 3.42 ;
      RECT 69.64 3.195 69.655 3.42 ;
      RECT 69.63 3.17 69.64 3.42 ;
      RECT 69.6 3.135 69.63 3.42 ;
      RECT 69.565 3.075 69.6 3.42 ;
      RECT 69.56 3.037 69.565 3.42 ;
      RECT 69.51 2.988 69.56 3.42 ;
      RECT 69.5 2.938 69.51 3.408 ;
      RECT 69.485 2.917 69.5 3.368 ;
      RECT 69.465 2.885 69.485 3.318 ;
      RECT 69.44 2.841 69.465 3.258 ;
      RECT 69.435 2.813 69.44 3.213 ;
      RECT 69.43 2.804 69.435 3.199 ;
      RECT 69.425 2.797 69.43 3.186 ;
      RECT 69.42 2.792 69.425 3.175 ;
      RECT 69.415 2.777 69.42 3.165 ;
      RECT 69.41 2.755 69.415 3.152 ;
      RECT 69.4 2.715 69.41 3.127 ;
      RECT 69.375 2.645 69.4 3.083 ;
      RECT 69.37 2.585 69.375 3.048 ;
      RECT 69.355 2.565 69.37 3.015 ;
      RECT 69.35 2.565 69.355 2.99 ;
      RECT 69.32 2.565 69.35 2.945 ;
      RECT 69.275 2.565 69.32 2.885 ;
      RECT 69.2 2.565 69.275 2.833 ;
      RECT 69.195 2.565 69.2 2.798 ;
      RECT 69.19 2.565 69.195 2.788 ;
      RECT 69.185 2.565 69.19 2.768 ;
      RECT 69.45 1.785 69.62 2.255 ;
      RECT 69.395 1.778 69.59 2.239 ;
      RECT 69.395 1.792 69.625 2.238 ;
      RECT 69.38 1.793 69.625 2.219 ;
      RECT 69.375 1.811 69.625 2.205 ;
      RECT 69.38 1.794 69.63 2.203 ;
      RECT 69.365 1.825 69.63 2.188 ;
      RECT 69.38 1.8 69.635 2.173 ;
      RECT 69.36 1.84 69.635 2.17 ;
      RECT 69.375 1.812 69.64 2.155 ;
      RECT 69.375 1.824 69.645 2.135 ;
      RECT 69.36 1.84 69.65 2.118 ;
      RECT 69.36 1.85 69.655 1.973 ;
      RECT 69.355 1.85 69.655 1.93 ;
      RECT 69.355 1.865 69.66 1.908 ;
      RECT 69.45 1.775 69.59 2.255 ;
      RECT 69.45 1.773 69.56 2.255 ;
      RECT 69.536 1.77 69.56 2.255 ;
      RECT 69.195 3.437 69.2 3.483 ;
      RECT 69.185 3.285 69.195 3.507 ;
      RECT 69.18 3.13 69.185 3.532 ;
      RECT 69.165 3.092 69.18 3.543 ;
      RECT 69.16 3.075 69.165 3.55 ;
      RECT 69.15 3.063 69.16 3.557 ;
      RECT 69.145 3.054 69.15 3.559 ;
      RECT 69.14 3.052 69.145 3.563 ;
      RECT 69.095 3.043 69.14 3.578 ;
      RECT 69.09 3.035 69.095 3.592 ;
      RECT 69.085 3.032 69.09 3.596 ;
      RECT 69.07 3.027 69.085 3.604 ;
      RECT 69.015 3.017 69.07 3.615 ;
      RECT 68.98 3.005 69.015 3.616 ;
      RECT 68.971 3 68.98 3.61 ;
      RECT 68.885 3 68.971 3.6 ;
      RECT 68.855 3 68.885 3.578 ;
      RECT 68.845 3 68.85 3.558 ;
      RECT 68.84 3 68.845 3.52 ;
      RECT 68.835 3 68.84 3.478 ;
      RECT 68.83 3 68.835 3.438 ;
      RECT 68.825 3 68.83 3.368 ;
      RECT 68.815 3 68.825 3.29 ;
      RECT 68.81 3 68.815 3.19 ;
      RECT 68.85 3 68.855 3.56 ;
      RECT 68.345 3.082 68.435 3.56 ;
      RECT 68.33 3.085 68.45 3.558 ;
      RECT 68.345 3.084 68.45 3.558 ;
      RECT 68.31 3.091 68.475 3.548 ;
      RECT 68.33 3.085 68.475 3.548 ;
      RECT 68.295 3.097 68.475 3.536 ;
      RECT 68.33 3.088 68.525 3.529 ;
      RECT 68.281 3.105 68.525 3.527 ;
      RECT 68.31 3.095 68.535 3.515 ;
      RECT 68.281 3.116 68.565 3.506 ;
      RECT 68.195 3.14 68.565 3.5 ;
      RECT 68.195 3.153 68.605 3.483 ;
      RECT 68.19 3.175 68.605 3.476 ;
      RECT 68.16 3.19 68.605 3.466 ;
      RECT 68.155 3.201 68.605 3.456 ;
      RECT 68.125 3.214 68.605 3.447 ;
      RECT 68.11 3.232 68.605 3.436 ;
      RECT 68.085 3.245 68.605 3.426 ;
      RECT 68.345 3.081 68.355 3.56 ;
      RECT 68.391 2.505 68.43 2.75 ;
      RECT 68.305 2.505 68.44 2.748 ;
      RECT 68.19 2.53 68.44 2.745 ;
      RECT 68.19 2.53 68.445 2.743 ;
      RECT 68.19 2.53 68.46 2.738 ;
      RECT 68.296 2.505 68.475 2.718 ;
      RECT 68.21 2.513 68.475 2.718 ;
      RECT 67.88 1.865 68.05 2.3 ;
      RECT 67.87 1.899 68.05 2.283 ;
      RECT 67.95 1.835 68.12 2.27 ;
      RECT 67.855 1.91 68.12 2.248 ;
      RECT 67.95 1.845 68.125 2.238 ;
      RECT 67.88 1.897 68.155 2.223 ;
      RECT 67.84 1.923 68.155 2.208 ;
      RECT 67.84 1.965 68.165 2.188 ;
      RECT 67.835 1.99 68.17 2.17 ;
      RECT 67.835 2 68.175 2.155 ;
      RECT 67.83 1.937 68.155 2.153 ;
      RECT 67.83 2.01 68.18 2.138 ;
      RECT 67.825 1.947 68.155 2.135 ;
      RECT 67.82 2.031 68.185 2.118 ;
      RECT 67.82 2.063 68.19 2.098 ;
      RECT 67.815 1.977 68.165 2.09 ;
      RECT 67.82 1.962 68.155 2.118 ;
      RECT 67.835 1.932 68.155 2.17 ;
      RECT 67.68 2.519 67.905 2.775 ;
      RECT 67.68 2.552 67.925 2.765 ;
      RECT 67.645 2.552 67.925 2.763 ;
      RECT 67.645 2.565 67.93 2.753 ;
      RECT 67.645 2.585 67.94 2.745 ;
      RECT 67.645 2.682 67.945 2.738 ;
      RECT 67.625 2.43 67.755 2.728 ;
      RECT 67.58 2.585 67.94 2.67 ;
      RECT 67.57 2.43 67.755 2.615 ;
      RECT 67.57 2.462 67.841 2.615 ;
      RECT 67.535 2.992 67.555 3.17 ;
      RECT 67.5 2.945 67.535 3.17 ;
      RECT 67.485 2.885 67.5 3.17 ;
      RECT 67.46 2.832 67.485 3.17 ;
      RECT 67.445 2.785 67.46 3.17 ;
      RECT 67.425 2.762 67.445 3.17 ;
      RECT 67.4 2.727 67.425 3.17 ;
      RECT 67.39 2.573 67.4 3.17 ;
      RECT 67.36 2.568 67.39 3.161 ;
      RECT 67.355 2.565 67.36 3.151 ;
      RECT 67.34 2.565 67.355 3.125 ;
      RECT 67.335 2.565 67.34 3.088 ;
      RECT 67.31 2.565 67.335 3.04 ;
      RECT 67.29 2.565 67.31 2.965 ;
      RECT 67.28 2.565 67.29 2.925 ;
      RECT 67.275 2.565 67.28 2.9 ;
      RECT 67.27 2.565 67.275 2.883 ;
      RECT 67.265 2.565 67.27 2.865 ;
      RECT 67.26 2.566 67.265 2.855 ;
      RECT 67.25 2.568 67.26 2.823 ;
      RECT 67.24 2.57 67.25 2.79 ;
      RECT 67.23 2.573 67.24 2.763 ;
      RECT 67.555 3 67.78 3.17 ;
      RECT 66.885 1.812 67.055 2.265 ;
      RECT 66.885 1.812 67.145 2.231 ;
      RECT 66.885 1.812 67.175 2.215 ;
      RECT 66.885 1.812 67.205 2.188 ;
      RECT 67.141 1.79 67.22 2.17 ;
      RECT 66.92 1.797 67.225 2.155 ;
      RECT 66.92 1.805 67.235 2.118 ;
      RECT 66.88 1.832 67.235 2.09 ;
      RECT 66.865 1.845 67.235 2.055 ;
      RECT 66.885 1.82 67.255 2.045 ;
      RECT 66.86 1.885 67.255 2.015 ;
      RECT 66.86 1.915 67.26 1.998 ;
      RECT 66.855 1.945 67.26 1.985 ;
      RECT 66.92 1.794 67.22 2.17 ;
      RECT 67.055 1.791 67.141 2.249 ;
      RECT 67.006 1.792 67.22 2.17 ;
      RECT 67.15 3.452 67.195 3.645 ;
      RECT 67.14 3.422 67.15 3.645 ;
      RECT 67.135 3.407 67.14 3.645 ;
      RECT 67.095 3.317 67.135 3.645 ;
      RECT 67.09 3.23 67.095 3.645 ;
      RECT 67.08 3.2 67.09 3.645 ;
      RECT 67.075 3.16 67.08 3.645 ;
      RECT 67.065 3.122 67.075 3.645 ;
      RECT 67.06 3.087 67.065 3.645 ;
      RECT 67.04 3.04 67.06 3.645 ;
      RECT 67.025 2.965 67.04 3.645 ;
      RECT 67.02 2.92 67.025 3.64 ;
      RECT 67.015 2.9 67.02 3.613 ;
      RECT 67.01 2.88 67.015 3.598 ;
      RECT 67.005 2.855 67.01 3.578 ;
      RECT 67 2.833 67.005 3.563 ;
      RECT 66.995 2.811 67 3.545 ;
      RECT 66.99 2.79 66.995 3.535 ;
      RECT 66.98 2.762 66.99 3.505 ;
      RECT 66.97 2.725 66.98 3.473 ;
      RECT 66.96 2.685 66.97 3.44 ;
      RECT 66.95 2.663 66.96 3.41 ;
      RECT 66.92 2.615 66.95 3.342 ;
      RECT 66.905 2.575 66.92 3.269 ;
      RECT 66.895 2.575 66.905 3.235 ;
      RECT 66.89 2.575 66.895 3.21 ;
      RECT 66.885 2.575 66.89 3.195 ;
      RECT 66.88 2.575 66.885 3.173 ;
      RECT 66.875 2.575 66.88 3.16 ;
      RECT 66.86 2.575 66.875 3.125 ;
      RECT 66.84 2.575 66.86 3.065 ;
      RECT 66.83 2.575 66.84 3.015 ;
      RECT 66.81 2.575 66.83 2.963 ;
      RECT 66.79 2.575 66.81 2.92 ;
      RECT 66.78 2.575 66.79 2.908 ;
      RECT 66.75 2.575 66.78 2.895 ;
      RECT 66.72 2.596 66.75 2.875 ;
      RECT 66.71 2.624 66.72 2.855 ;
      RECT 66.695 2.641 66.71 2.823 ;
      RECT 66.69 2.655 66.695 2.79 ;
      RECT 66.685 2.663 66.69 2.763 ;
      RECT 66.68 2.671 66.685 2.725 ;
      RECT 66.685 3.195 66.69 3.53 ;
      RECT 66.65 3.182 66.685 3.529 ;
      RECT 66.58 3.122 66.65 3.528 ;
      RECT 66.5 3.065 66.58 3.527 ;
      RECT 66.365 3.025 66.5 3.526 ;
      RECT 66.365 3.212 66.7 3.515 ;
      RECT 66.325 3.212 66.7 3.505 ;
      RECT 66.325 3.23 66.705 3.5 ;
      RECT 66.325 3.32 66.71 3.49 ;
      RECT 66.32 3.015 66.485 3.47 ;
      RECT 66.315 3.015 66.485 3.213 ;
      RECT 66.315 3.172 66.68 3.213 ;
      RECT 66.315 3.16 66.675 3.213 ;
      RECT 65.445 5.02 65.615 6.49 ;
      RECT 65.445 6.315 65.62 6.485 ;
      RECT 65.075 1.74 65.245 2.93 ;
      RECT 65.075 1.74 65.545 1.91 ;
      RECT 65.075 6.97 65.545 7.14 ;
      RECT 65.075 5.95 65.245 7.14 ;
      RECT 64.085 1.74 64.255 2.93 ;
      RECT 64.085 1.74 64.555 1.91 ;
      RECT 64.085 6.97 64.555 7.14 ;
      RECT 64.085 5.95 64.255 7.14 ;
      RECT 62.235 2.635 62.405 3.865 ;
      RECT 62.29 0.855 62.46 2.805 ;
      RECT 62.235 0.575 62.405 1.025 ;
      RECT 62.235 7.855 62.405 8.305 ;
      RECT 62.29 6.075 62.46 8.025 ;
      RECT 62.235 5.015 62.405 6.245 ;
      RECT 61.715 0.575 61.885 3.865 ;
      RECT 61.715 2.075 62.12 2.405 ;
      RECT 61.715 1.235 62.12 1.565 ;
      RECT 61.715 5.015 61.885 8.305 ;
      RECT 61.715 7.315 62.12 7.645 ;
      RECT 61.715 6.475 62.12 6.805 ;
      RECT 59.05 1.975 59.78 2.215 ;
      RECT 59.592 1.77 59.78 2.215 ;
      RECT 59.42 1.782 59.795 2.209 ;
      RECT 59.335 1.797 59.815 2.194 ;
      RECT 59.335 1.812 59.82 2.184 ;
      RECT 59.29 1.832 59.835 2.176 ;
      RECT 59.267 1.867 59.85 2.13 ;
      RECT 59.181 1.89 59.855 2.09 ;
      RECT 59.181 1.908 59.865 2.06 ;
      RECT 59.05 1.977 59.87 2.023 ;
      RECT 59.095 1.92 59.865 2.06 ;
      RECT 59.181 1.872 59.85 2.13 ;
      RECT 59.267 1.841 59.835 2.176 ;
      RECT 59.29 1.822 59.82 2.184 ;
      RECT 59.335 1.795 59.795 2.209 ;
      RECT 59.42 1.777 59.78 2.215 ;
      RECT 59.506 1.771 59.78 2.215 ;
      RECT 59.592 1.766 59.725 2.215 ;
      RECT 59.678 1.761 59.725 2.215 ;
      RECT 59.37 2.659 59.54 3.045 ;
      RECT 59.365 2.659 59.54 3.04 ;
      RECT 59.34 2.659 59.54 3.005 ;
      RECT 59.34 2.687 59.55 2.995 ;
      RECT 59.32 2.687 59.55 2.955 ;
      RECT 59.315 2.687 59.55 2.928 ;
      RECT 59.315 2.705 59.555 2.92 ;
      RECT 59.26 2.705 59.555 2.855 ;
      RECT 59.26 2.722 59.565 2.838 ;
      RECT 59.25 2.722 59.565 2.778 ;
      RECT 59.25 2.739 59.57 2.775 ;
      RECT 59.245 2.575 59.415 2.753 ;
      RECT 59.245 2.609 59.501 2.753 ;
      RECT 59.24 3.375 59.245 3.388 ;
      RECT 59.235 3.27 59.24 3.393 ;
      RECT 59.21 3.13 59.235 3.408 ;
      RECT 59.175 3.081 59.21 3.44 ;
      RECT 59.17 3.049 59.175 3.46 ;
      RECT 59.165 3.04 59.17 3.46 ;
      RECT 59.085 3.005 59.165 3.46 ;
      RECT 59.022 2.975 59.085 3.46 ;
      RECT 58.936 2.963 59.022 3.46 ;
      RECT 58.85 2.949 58.936 3.46 ;
      RECT 58.77 2.936 58.85 3.446 ;
      RECT 58.735 2.928 58.77 3.426 ;
      RECT 58.725 2.925 58.735 3.417 ;
      RECT 58.695 2.92 58.725 3.404 ;
      RECT 58.645 2.895 58.695 3.38 ;
      RECT 58.631 2.869 58.645 3.362 ;
      RECT 58.545 2.829 58.631 3.338 ;
      RECT 58.5 2.777 58.545 3.307 ;
      RECT 58.49 2.752 58.5 3.294 ;
      RECT 58.485 2.533 58.49 2.555 ;
      RECT 58.48 2.735 58.49 3.29 ;
      RECT 58.48 2.531 58.485 2.645 ;
      RECT 58.47 2.527 58.48 3.286 ;
      RECT 58.426 2.525 58.47 3.274 ;
      RECT 58.34 2.525 58.426 3.245 ;
      RECT 58.31 2.525 58.34 3.218 ;
      RECT 58.295 2.525 58.31 3.206 ;
      RECT 58.255 2.537 58.295 3.191 ;
      RECT 58.235 2.556 58.255 3.17 ;
      RECT 58.225 2.566 58.235 3.154 ;
      RECT 58.215 2.572 58.225 3.143 ;
      RECT 58.195 2.582 58.215 3.126 ;
      RECT 58.19 2.591 58.195 3.113 ;
      RECT 58.185 2.595 58.19 3.063 ;
      RECT 58.175 2.601 58.185 2.98 ;
      RECT 58.17 2.605 58.175 2.894 ;
      RECT 58.165 2.625 58.17 2.831 ;
      RECT 58.16 2.648 58.165 2.778 ;
      RECT 58.155 2.666 58.16 2.723 ;
      RECT 58.765 2.485 58.935 2.745 ;
      RECT 58.935 2.45 58.98 2.731 ;
      RECT 58.896 2.452 58.985 2.714 ;
      RECT 58.785 2.469 59.071 2.685 ;
      RECT 58.785 2.484 59.075 2.657 ;
      RECT 58.785 2.465 58.985 2.714 ;
      RECT 58.81 2.453 58.935 2.745 ;
      RECT 58.896 2.451 58.98 2.731 ;
      RECT 57.95 1.84 58.12 2.33 ;
      RECT 57.95 1.84 58.155 2.31 ;
      RECT 58.085 1.76 58.195 2.27 ;
      RECT 58.066 1.764 58.215 2.24 ;
      RECT 57.98 1.772 58.235 2.223 ;
      RECT 57.98 1.778 58.24 2.213 ;
      RECT 57.98 1.787 58.26 2.201 ;
      RECT 57.955 1.812 58.29 2.179 ;
      RECT 57.955 1.832 58.295 2.159 ;
      RECT 57.95 1.845 58.305 2.139 ;
      RECT 57.95 1.912 58.31 2.12 ;
      RECT 57.95 2.045 58.315 2.107 ;
      RECT 57.945 1.85 58.305 1.94 ;
      RECT 57.955 1.807 58.26 2.201 ;
      RECT 58.066 1.762 58.195 2.27 ;
      RECT 57.94 3.515 58.24 3.77 ;
      RECT 58.025 3.481 58.24 3.77 ;
      RECT 58.025 3.484 58.245 3.63 ;
      RECT 57.96 3.505 58.245 3.63 ;
      RECT 57.995 3.495 58.24 3.77 ;
      RECT 57.99 3.5 58.245 3.63 ;
      RECT 58.025 3.479 58.226 3.77 ;
      RECT 58.111 3.47 58.226 3.77 ;
      RECT 58.111 3.464 58.14 3.77 ;
      RECT 57.6 3.105 57.61 3.595 ;
      RECT 57.26 3.04 57.27 3.34 ;
      RECT 57.775 3.212 57.78 3.431 ;
      RECT 57.765 3.192 57.775 3.448 ;
      RECT 57.755 3.172 57.765 3.478 ;
      RECT 57.75 3.162 57.755 3.493 ;
      RECT 57.745 3.158 57.75 3.498 ;
      RECT 57.73 3.15 57.745 3.505 ;
      RECT 57.69 3.13 57.73 3.53 ;
      RECT 57.665 3.112 57.69 3.563 ;
      RECT 57.66 3.11 57.665 3.576 ;
      RECT 57.64 3.107 57.66 3.58 ;
      RECT 57.61 3.105 57.64 3.59 ;
      RECT 57.54 3.107 57.6 3.591 ;
      RECT 57.52 3.107 57.54 3.585 ;
      RECT 57.495 3.105 57.52 3.582 ;
      RECT 57.46 3.1 57.495 3.578 ;
      RECT 57.44 3.094 57.46 3.565 ;
      RECT 57.43 3.091 57.44 3.553 ;
      RECT 57.41 3.088 57.43 3.538 ;
      RECT 57.39 3.084 57.41 3.52 ;
      RECT 57.385 3.081 57.39 3.51 ;
      RECT 57.38 3.08 57.385 3.508 ;
      RECT 57.37 3.077 57.38 3.5 ;
      RECT 57.36 3.071 57.37 3.483 ;
      RECT 57.35 3.065 57.36 3.465 ;
      RECT 57.34 3.059 57.35 3.453 ;
      RECT 57.33 3.053 57.34 3.433 ;
      RECT 57.325 3.049 57.33 3.418 ;
      RECT 57.32 3.047 57.325 3.41 ;
      RECT 57.315 3.045 57.32 3.403 ;
      RECT 57.31 3.043 57.315 3.393 ;
      RECT 57.305 3.041 57.31 3.387 ;
      RECT 57.295 3.04 57.305 3.377 ;
      RECT 57.285 3.04 57.295 3.368 ;
      RECT 57.27 3.04 57.285 3.353 ;
      RECT 57.23 3.04 57.26 3.337 ;
      RECT 57.21 3.042 57.23 3.332 ;
      RECT 57.205 3.047 57.21 3.33 ;
      RECT 57.175 3.055 57.205 3.328 ;
      RECT 57.145 3.07 57.175 3.327 ;
      RECT 57.1 3.092 57.145 3.332 ;
      RECT 57.095 3.107 57.1 3.336 ;
      RECT 57.08 3.112 57.095 3.338 ;
      RECT 57.075 3.116 57.08 3.34 ;
      RECT 57.015 3.139 57.075 3.349 ;
      RECT 56.995 3.165 57.015 3.362 ;
      RECT 56.985 3.172 56.995 3.366 ;
      RECT 56.97 3.179 56.985 3.369 ;
      RECT 56.95 3.189 56.97 3.372 ;
      RECT 56.945 3.197 56.95 3.375 ;
      RECT 56.9 3.202 56.945 3.382 ;
      RECT 56.89 3.205 56.9 3.389 ;
      RECT 56.88 3.205 56.89 3.393 ;
      RECT 56.845 3.207 56.88 3.405 ;
      RECT 56.825 3.21 56.845 3.418 ;
      RECT 56.785 3.213 56.825 3.429 ;
      RECT 56.77 3.215 56.785 3.442 ;
      RECT 56.76 3.215 56.77 3.447 ;
      RECT 56.735 3.216 56.76 3.455 ;
      RECT 56.725 3.218 56.735 3.46 ;
      RECT 56.72 3.219 56.725 3.463 ;
      RECT 56.695 3.217 56.72 3.466 ;
      RECT 56.68 3.215 56.695 3.467 ;
      RECT 56.66 3.212 56.68 3.469 ;
      RECT 56.64 3.207 56.66 3.469 ;
      RECT 56.58 3.202 56.64 3.466 ;
      RECT 56.545 3.177 56.58 3.462 ;
      RECT 56.535 3.154 56.545 3.46 ;
      RECT 56.505 3.131 56.535 3.46 ;
      RECT 56.495 3.11 56.505 3.46 ;
      RECT 56.47 3.092 56.495 3.458 ;
      RECT 56.455 3.07 56.47 3.455 ;
      RECT 56.44 3.052 56.455 3.453 ;
      RECT 56.42 3.042 56.44 3.451 ;
      RECT 56.405 3.037 56.42 3.45 ;
      RECT 56.39 3.035 56.405 3.449 ;
      RECT 56.36 3.036 56.39 3.447 ;
      RECT 56.34 3.039 56.36 3.445 ;
      RECT 56.283 3.043 56.34 3.445 ;
      RECT 56.197 3.052 56.283 3.445 ;
      RECT 56.111 3.063 56.197 3.445 ;
      RECT 56.025 3.074 56.111 3.445 ;
      RECT 56.005 3.081 56.025 3.453 ;
      RECT 55.995 3.084 56.005 3.46 ;
      RECT 55.93 3.089 55.995 3.478 ;
      RECT 55.9 3.096 55.93 3.503 ;
      RECT 55.89 3.099 55.9 3.51 ;
      RECT 55.845 3.103 55.89 3.515 ;
      RECT 55.815 3.108 55.845 3.52 ;
      RECT 55.814 3.11 55.815 3.52 ;
      RECT 55.728 3.116 55.814 3.52 ;
      RECT 55.642 3.127 55.728 3.52 ;
      RECT 55.556 3.139 55.642 3.52 ;
      RECT 55.47 3.15 55.556 3.52 ;
      RECT 55.455 3.157 55.47 3.515 ;
      RECT 55.45 3.159 55.455 3.509 ;
      RECT 55.43 3.17 55.45 3.504 ;
      RECT 55.42 3.188 55.43 3.498 ;
      RECT 55.415 3.2 55.42 3.298 ;
      RECT 57.71 1.953 57.73 2.04 ;
      RECT 57.705 1.888 57.71 2.072 ;
      RECT 57.695 1.855 57.705 2.077 ;
      RECT 57.69 1.835 57.695 2.083 ;
      RECT 57.66 1.835 57.69 2.1 ;
      RECT 57.611 1.835 57.66 2.136 ;
      RECT 57.525 1.835 57.611 2.194 ;
      RECT 57.496 1.845 57.525 2.243 ;
      RECT 57.41 1.887 57.496 2.296 ;
      RECT 57.39 1.925 57.41 2.343 ;
      RECT 57.365 1.942 57.39 2.363 ;
      RECT 57.355 1.956 57.365 2.383 ;
      RECT 57.35 1.962 57.355 2.393 ;
      RECT 57.345 1.966 57.35 2.4 ;
      RECT 57.295 1.986 57.345 2.405 ;
      RECT 57.23 2.03 57.295 2.405 ;
      RECT 57.205 2.08 57.23 2.405 ;
      RECT 57.195 2.11 57.205 2.405 ;
      RECT 57.19 2.137 57.195 2.405 ;
      RECT 57.185 2.155 57.19 2.405 ;
      RECT 57.175 2.197 57.185 2.405 ;
      RECT 57.525 2.755 57.695 2.93 ;
      RECT 57.465 2.583 57.525 2.918 ;
      RECT 57.455 2.576 57.465 2.901 ;
      RECT 57.41 2.755 57.695 2.881 ;
      RECT 57.391 2.755 57.695 2.859 ;
      RECT 57.305 2.755 57.695 2.824 ;
      RECT 57.285 2.575 57.455 2.78 ;
      RECT 57.285 2.722 57.69 2.78 ;
      RECT 57.285 2.67 57.665 2.78 ;
      RECT 57.285 2.625 57.63 2.78 ;
      RECT 57.285 2.607 57.595 2.78 ;
      RECT 57.285 2.597 57.59 2.78 ;
      RECT 57.455 7.855 57.625 8.305 ;
      RECT 57.51 6.075 57.68 8.025 ;
      RECT 57.455 5.015 57.625 6.245 ;
      RECT 56.935 5.015 57.105 8.305 ;
      RECT 56.935 7.315 57.34 7.645 ;
      RECT 56.935 6.475 57.34 6.805 ;
      RECT 57.005 3.555 57.195 3.78 ;
      RECT 56.995 3.556 57.2 3.775 ;
      RECT 56.995 3.558 57.21 3.755 ;
      RECT 56.995 3.562 57.215 3.74 ;
      RECT 56.995 3.549 57.165 3.775 ;
      RECT 56.995 3.552 57.19 3.775 ;
      RECT 57.005 3.548 57.165 3.78 ;
      RECT 57.091 3.546 57.165 3.78 ;
      RECT 56.715 2.797 56.885 3.035 ;
      RECT 56.715 2.797 56.971 2.949 ;
      RECT 56.715 2.797 56.975 2.859 ;
      RECT 56.765 2.57 56.985 2.838 ;
      RECT 56.76 2.587 56.99 2.811 ;
      RECT 56.725 2.745 56.99 2.811 ;
      RECT 56.745 2.595 56.885 3.035 ;
      RECT 56.735 2.677 56.995 2.794 ;
      RECT 56.73 2.725 56.995 2.794 ;
      RECT 56.735 2.635 56.99 2.811 ;
      RECT 56.76 2.572 56.985 2.838 ;
      RECT 56.325 2.547 56.495 2.745 ;
      RECT 56.325 2.547 56.54 2.72 ;
      RECT 56.395 2.49 56.565 2.678 ;
      RECT 56.37 2.505 56.565 2.678 ;
      RECT 55.985 2.551 56.015 2.745 ;
      RECT 55.98 2.523 55.985 2.745 ;
      RECT 55.95 2.497 55.98 2.747 ;
      RECT 55.925 2.455 55.95 2.75 ;
      RECT 55.915 2.427 55.925 2.752 ;
      RECT 55.88 2.407 55.915 2.754 ;
      RECT 55.815 2.392 55.88 2.76 ;
      RECT 55.765 2.39 55.815 2.766 ;
      RECT 55.742 2.392 55.765 2.771 ;
      RECT 55.656 2.403 55.742 2.777 ;
      RECT 55.57 2.421 55.656 2.787 ;
      RECT 55.555 2.432 55.57 2.793 ;
      RECT 55.485 2.455 55.555 2.799 ;
      RECT 55.43 2.487 55.485 2.807 ;
      RECT 55.39 2.51 55.43 2.813 ;
      RECT 55.376 2.523 55.39 2.816 ;
      RECT 55.29 2.545 55.376 2.822 ;
      RECT 55.275 2.57 55.29 2.828 ;
      RECT 55.235 2.585 55.275 2.832 ;
      RECT 55.185 2.6 55.235 2.837 ;
      RECT 55.16 2.607 55.185 2.841 ;
      RECT 55.1 2.602 55.16 2.845 ;
      RECT 55.085 2.593 55.1 2.849 ;
      RECT 55.015 2.583 55.085 2.845 ;
      RECT 54.99 2.575 55.01 2.835 ;
      RECT 54.931 2.575 54.99 2.813 ;
      RECT 54.845 2.575 54.931 2.77 ;
      RECT 55.01 2.575 55.015 2.84 ;
      RECT 55.705 1.806 55.875 2.14 ;
      RECT 55.675 1.806 55.875 2.135 ;
      RECT 55.615 1.773 55.675 2.123 ;
      RECT 55.615 1.829 55.885 2.118 ;
      RECT 55.59 1.829 55.885 2.112 ;
      RECT 55.585 1.77 55.615 2.109 ;
      RECT 55.57 1.776 55.705 2.107 ;
      RECT 55.565 1.784 55.79 2.095 ;
      RECT 55.565 1.836 55.9 2.048 ;
      RECT 55.55 1.792 55.79 2.043 ;
      RECT 55.55 1.862 55.91 1.984 ;
      RECT 55.52 1.812 55.875 1.945 ;
      RECT 55.52 1.902 55.92 1.941 ;
      RECT 55.57 1.781 55.79 2.107 ;
      RECT 54.91 2.111 54.965 2.375 ;
      RECT 54.91 2.111 55.03 2.374 ;
      RECT 54.91 2.111 55.055 2.373 ;
      RECT 54.91 2.111 55.12 2.372 ;
      RECT 55.055 2.077 55.135 2.371 ;
      RECT 54.87 2.121 55.28 2.37 ;
      RECT 54.91 2.118 55.28 2.37 ;
      RECT 54.87 2.126 55.285 2.363 ;
      RECT 54.855 2.128 55.285 2.362 ;
      RECT 54.855 2.135 55.29 2.358 ;
      RECT 54.835 2.134 55.285 2.354 ;
      RECT 54.835 2.142 55.295 2.353 ;
      RECT 54.83 2.139 55.29 2.349 ;
      RECT 54.83 2.152 55.305 2.348 ;
      RECT 54.815 2.142 55.295 2.347 ;
      RECT 54.78 2.155 55.305 2.34 ;
      RECT 54.965 2.11 55.275 2.37 ;
      RECT 54.965 2.095 55.225 2.37 ;
      RECT 55.03 2.082 55.16 2.37 ;
      RECT 54.575 3.171 54.59 3.564 ;
      RECT 54.54 3.176 54.59 3.563 ;
      RECT 54.575 3.175 54.635 3.562 ;
      RECT 54.52 3.186 54.635 3.561 ;
      RECT 54.535 3.182 54.635 3.561 ;
      RECT 54.5 3.192 54.71 3.558 ;
      RECT 54.5 3.211 54.755 3.556 ;
      RECT 54.5 3.218 54.76 3.553 ;
      RECT 54.485 3.195 54.71 3.55 ;
      RECT 54.465 3.2 54.71 3.543 ;
      RECT 54.46 3.204 54.71 3.539 ;
      RECT 54.46 3.221 54.77 3.538 ;
      RECT 54.44 3.215 54.755 3.534 ;
      RECT 54.44 3.224 54.775 3.528 ;
      RECT 54.435 3.23 54.775 3.3 ;
      RECT 54.5 3.19 54.635 3.558 ;
      RECT 54.375 2.553 54.575 2.865 ;
      RECT 54.45 2.531 54.575 2.865 ;
      RECT 54.39 2.55 54.58 2.85 ;
      RECT 54.36 2.561 54.58 2.848 ;
      RECT 54.375 2.556 54.585 2.814 ;
      RECT 54.36 2.66 54.59 2.781 ;
      RECT 54.39 2.532 54.575 2.865 ;
      RECT 54.45 2.51 54.55 2.865 ;
      RECT 54.475 2.507 54.55 2.865 ;
      RECT 54.475 2.502 54.495 2.865 ;
      RECT 53.88 2.57 54.055 2.745 ;
      RECT 53.875 2.57 54.055 2.743 ;
      RECT 53.85 2.57 54.055 2.738 ;
      RECT 53.795 2.55 53.965 2.728 ;
      RECT 53.795 2.557 54.03 2.728 ;
      RECT 53.88 3.237 53.895 3.42 ;
      RECT 53.87 3.215 53.88 3.42 ;
      RECT 53.855 3.195 53.87 3.42 ;
      RECT 53.845 3.17 53.855 3.42 ;
      RECT 53.815 3.135 53.845 3.42 ;
      RECT 53.78 3.075 53.815 3.42 ;
      RECT 53.775 3.037 53.78 3.42 ;
      RECT 53.725 2.988 53.775 3.42 ;
      RECT 53.715 2.938 53.725 3.408 ;
      RECT 53.7 2.917 53.715 3.368 ;
      RECT 53.68 2.885 53.7 3.318 ;
      RECT 53.655 2.841 53.68 3.258 ;
      RECT 53.65 2.813 53.655 3.213 ;
      RECT 53.645 2.804 53.65 3.199 ;
      RECT 53.64 2.797 53.645 3.186 ;
      RECT 53.635 2.792 53.64 3.175 ;
      RECT 53.63 2.777 53.635 3.165 ;
      RECT 53.625 2.755 53.63 3.152 ;
      RECT 53.615 2.715 53.625 3.127 ;
      RECT 53.59 2.645 53.615 3.083 ;
      RECT 53.585 2.585 53.59 3.048 ;
      RECT 53.57 2.565 53.585 3.015 ;
      RECT 53.565 2.565 53.57 2.99 ;
      RECT 53.535 2.565 53.565 2.945 ;
      RECT 53.49 2.565 53.535 2.885 ;
      RECT 53.415 2.565 53.49 2.833 ;
      RECT 53.41 2.565 53.415 2.798 ;
      RECT 53.405 2.565 53.41 2.788 ;
      RECT 53.4 2.565 53.405 2.768 ;
      RECT 53.665 1.785 53.835 2.255 ;
      RECT 53.61 1.778 53.805 2.239 ;
      RECT 53.61 1.792 53.84 2.238 ;
      RECT 53.595 1.793 53.84 2.219 ;
      RECT 53.59 1.811 53.84 2.205 ;
      RECT 53.595 1.794 53.845 2.203 ;
      RECT 53.58 1.825 53.845 2.188 ;
      RECT 53.595 1.8 53.85 2.173 ;
      RECT 53.575 1.84 53.85 2.17 ;
      RECT 53.59 1.812 53.855 2.155 ;
      RECT 53.59 1.824 53.86 2.135 ;
      RECT 53.575 1.84 53.865 2.118 ;
      RECT 53.575 1.85 53.87 1.973 ;
      RECT 53.57 1.85 53.87 1.93 ;
      RECT 53.57 1.865 53.875 1.908 ;
      RECT 53.665 1.775 53.805 2.255 ;
      RECT 53.665 1.773 53.775 2.255 ;
      RECT 53.751 1.77 53.775 2.255 ;
      RECT 53.41 3.437 53.415 3.483 ;
      RECT 53.4 3.285 53.41 3.507 ;
      RECT 53.395 3.13 53.4 3.532 ;
      RECT 53.38 3.092 53.395 3.543 ;
      RECT 53.375 3.075 53.38 3.55 ;
      RECT 53.365 3.063 53.375 3.557 ;
      RECT 53.36 3.054 53.365 3.559 ;
      RECT 53.355 3.052 53.36 3.563 ;
      RECT 53.31 3.043 53.355 3.578 ;
      RECT 53.305 3.035 53.31 3.592 ;
      RECT 53.3 3.032 53.305 3.596 ;
      RECT 53.285 3.027 53.3 3.604 ;
      RECT 53.23 3.017 53.285 3.615 ;
      RECT 53.195 3.005 53.23 3.616 ;
      RECT 53.186 3 53.195 3.61 ;
      RECT 53.1 3 53.186 3.6 ;
      RECT 53.07 3 53.1 3.578 ;
      RECT 53.06 3 53.065 3.558 ;
      RECT 53.055 3 53.06 3.52 ;
      RECT 53.05 3 53.055 3.478 ;
      RECT 53.045 3 53.05 3.438 ;
      RECT 53.04 3 53.045 3.368 ;
      RECT 53.03 3 53.04 3.29 ;
      RECT 53.025 3 53.03 3.19 ;
      RECT 53.065 3 53.07 3.56 ;
      RECT 52.56 3.082 52.65 3.56 ;
      RECT 52.545 3.085 52.665 3.558 ;
      RECT 52.56 3.084 52.665 3.558 ;
      RECT 52.525 3.091 52.69 3.548 ;
      RECT 52.545 3.085 52.69 3.548 ;
      RECT 52.51 3.097 52.69 3.536 ;
      RECT 52.545 3.088 52.74 3.529 ;
      RECT 52.496 3.105 52.74 3.527 ;
      RECT 52.525 3.095 52.75 3.515 ;
      RECT 52.496 3.116 52.78 3.506 ;
      RECT 52.41 3.14 52.78 3.5 ;
      RECT 52.41 3.153 52.82 3.483 ;
      RECT 52.405 3.175 52.82 3.476 ;
      RECT 52.375 3.19 52.82 3.466 ;
      RECT 52.37 3.201 52.82 3.456 ;
      RECT 52.34 3.214 52.82 3.447 ;
      RECT 52.325 3.232 52.82 3.436 ;
      RECT 52.3 3.245 52.82 3.426 ;
      RECT 52.56 3.081 52.57 3.56 ;
      RECT 52.606 2.505 52.645 2.75 ;
      RECT 52.52 2.505 52.655 2.748 ;
      RECT 52.405 2.53 52.655 2.745 ;
      RECT 52.405 2.53 52.66 2.743 ;
      RECT 52.405 2.53 52.675 2.738 ;
      RECT 52.511 2.505 52.69 2.718 ;
      RECT 52.425 2.513 52.69 2.718 ;
      RECT 52.095 1.865 52.265 2.3 ;
      RECT 52.085 1.899 52.265 2.283 ;
      RECT 52.165 1.835 52.335 2.27 ;
      RECT 52.07 1.91 52.335 2.248 ;
      RECT 52.165 1.845 52.34 2.238 ;
      RECT 52.095 1.897 52.37 2.223 ;
      RECT 52.055 1.923 52.37 2.208 ;
      RECT 52.055 1.965 52.38 2.188 ;
      RECT 52.05 1.99 52.385 2.17 ;
      RECT 52.05 2 52.39 2.155 ;
      RECT 52.045 1.937 52.37 2.153 ;
      RECT 52.045 2.01 52.395 2.138 ;
      RECT 52.04 1.947 52.37 2.135 ;
      RECT 52.035 2.031 52.4 2.118 ;
      RECT 52.035 2.063 52.405 2.098 ;
      RECT 52.03 1.977 52.38 2.09 ;
      RECT 52.035 1.962 52.37 2.118 ;
      RECT 52.05 1.932 52.37 2.17 ;
      RECT 51.895 2.519 52.12 2.775 ;
      RECT 51.895 2.552 52.14 2.765 ;
      RECT 51.86 2.552 52.14 2.763 ;
      RECT 51.86 2.565 52.145 2.753 ;
      RECT 51.86 2.585 52.155 2.745 ;
      RECT 51.86 2.682 52.16 2.738 ;
      RECT 51.84 2.43 51.97 2.728 ;
      RECT 51.795 2.585 52.155 2.67 ;
      RECT 51.785 2.43 51.97 2.615 ;
      RECT 51.785 2.462 52.056 2.615 ;
      RECT 51.75 2.992 51.77 3.17 ;
      RECT 51.715 2.945 51.75 3.17 ;
      RECT 51.7 2.885 51.715 3.17 ;
      RECT 51.675 2.832 51.7 3.17 ;
      RECT 51.66 2.785 51.675 3.17 ;
      RECT 51.64 2.762 51.66 3.17 ;
      RECT 51.615 2.727 51.64 3.17 ;
      RECT 51.605 2.573 51.615 3.17 ;
      RECT 51.575 2.568 51.605 3.161 ;
      RECT 51.57 2.565 51.575 3.151 ;
      RECT 51.555 2.565 51.57 3.125 ;
      RECT 51.55 2.565 51.555 3.088 ;
      RECT 51.525 2.565 51.55 3.04 ;
      RECT 51.505 2.565 51.525 2.965 ;
      RECT 51.495 2.565 51.505 2.925 ;
      RECT 51.49 2.565 51.495 2.9 ;
      RECT 51.485 2.565 51.49 2.883 ;
      RECT 51.48 2.565 51.485 2.865 ;
      RECT 51.475 2.566 51.48 2.855 ;
      RECT 51.465 2.568 51.475 2.823 ;
      RECT 51.455 2.57 51.465 2.79 ;
      RECT 51.445 2.573 51.455 2.763 ;
      RECT 51.77 3 51.995 3.17 ;
      RECT 51.1 1.812 51.27 2.265 ;
      RECT 51.1 1.812 51.36 2.231 ;
      RECT 51.1 1.812 51.39 2.215 ;
      RECT 51.1 1.812 51.42 2.188 ;
      RECT 51.356 1.79 51.435 2.17 ;
      RECT 51.135 1.797 51.44 2.155 ;
      RECT 51.135 1.805 51.45 2.118 ;
      RECT 51.095 1.832 51.45 2.09 ;
      RECT 51.08 1.845 51.45 2.055 ;
      RECT 51.1 1.82 51.47 2.045 ;
      RECT 51.075 1.885 51.47 2.015 ;
      RECT 51.075 1.915 51.475 1.998 ;
      RECT 51.07 1.945 51.475 1.985 ;
      RECT 51.135 1.794 51.435 2.17 ;
      RECT 51.27 1.791 51.356 2.249 ;
      RECT 51.221 1.792 51.435 2.17 ;
      RECT 51.365 3.452 51.41 3.645 ;
      RECT 51.355 3.422 51.365 3.645 ;
      RECT 51.35 3.407 51.355 3.645 ;
      RECT 51.31 3.317 51.35 3.645 ;
      RECT 51.305 3.23 51.31 3.645 ;
      RECT 51.295 3.2 51.305 3.645 ;
      RECT 51.29 3.16 51.295 3.645 ;
      RECT 51.28 3.122 51.29 3.645 ;
      RECT 51.275 3.087 51.28 3.645 ;
      RECT 51.255 3.04 51.275 3.645 ;
      RECT 51.24 2.965 51.255 3.645 ;
      RECT 51.235 2.92 51.24 3.64 ;
      RECT 51.23 2.9 51.235 3.613 ;
      RECT 51.225 2.88 51.23 3.598 ;
      RECT 51.22 2.855 51.225 3.578 ;
      RECT 51.215 2.833 51.22 3.563 ;
      RECT 51.21 2.811 51.215 3.545 ;
      RECT 51.205 2.79 51.21 3.535 ;
      RECT 51.195 2.762 51.205 3.505 ;
      RECT 51.185 2.725 51.195 3.473 ;
      RECT 51.175 2.685 51.185 3.44 ;
      RECT 51.165 2.663 51.175 3.41 ;
      RECT 51.135 2.615 51.165 3.342 ;
      RECT 51.12 2.575 51.135 3.269 ;
      RECT 51.11 2.575 51.12 3.235 ;
      RECT 51.105 2.575 51.11 3.21 ;
      RECT 51.1 2.575 51.105 3.195 ;
      RECT 51.095 2.575 51.1 3.173 ;
      RECT 51.09 2.575 51.095 3.16 ;
      RECT 51.075 2.575 51.09 3.125 ;
      RECT 51.055 2.575 51.075 3.065 ;
      RECT 51.045 2.575 51.055 3.015 ;
      RECT 51.025 2.575 51.045 2.963 ;
      RECT 51.005 2.575 51.025 2.92 ;
      RECT 50.995 2.575 51.005 2.908 ;
      RECT 50.965 2.575 50.995 2.895 ;
      RECT 50.935 2.596 50.965 2.875 ;
      RECT 50.925 2.624 50.935 2.855 ;
      RECT 50.91 2.641 50.925 2.823 ;
      RECT 50.905 2.655 50.91 2.79 ;
      RECT 50.9 2.663 50.905 2.763 ;
      RECT 50.895 2.671 50.9 2.725 ;
      RECT 50.9 3.195 50.905 3.53 ;
      RECT 50.865 3.182 50.9 3.529 ;
      RECT 50.795 3.122 50.865 3.528 ;
      RECT 50.715 3.065 50.795 3.527 ;
      RECT 50.58 3.025 50.715 3.526 ;
      RECT 50.58 3.212 50.915 3.515 ;
      RECT 50.54 3.212 50.915 3.505 ;
      RECT 50.54 3.23 50.92 3.5 ;
      RECT 50.54 3.32 50.925 3.49 ;
      RECT 50.535 3.015 50.7 3.47 ;
      RECT 50.53 3.015 50.7 3.213 ;
      RECT 50.53 3.172 50.895 3.213 ;
      RECT 50.53 3.16 50.89 3.213 ;
      RECT 49.66 5.02 49.83 6.49 ;
      RECT 49.66 6.315 49.835 6.485 ;
      RECT 49.29 1.74 49.46 2.93 ;
      RECT 49.29 1.74 49.76 1.91 ;
      RECT 49.29 6.97 49.76 7.14 ;
      RECT 49.29 5.95 49.46 7.14 ;
      RECT 48.3 1.74 48.47 2.93 ;
      RECT 48.3 1.74 48.77 1.91 ;
      RECT 48.3 6.97 48.77 7.14 ;
      RECT 48.3 5.95 48.47 7.14 ;
      RECT 46.45 2.635 46.62 3.865 ;
      RECT 46.505 0.855 46.675 2.805 ;
      RECT 46.45 0.575 46.62 1.025 ;
      RECT 46.45 7.855 46.62 8.305 ;
      RECT 46.505 6.075 46.675 8.025 ;
      RECT 46.45 5.015 46.62 6.245 ;
      RECT 45.93 0.575 46.1 3.865 ;
      RECT 45.93 2.075 46.335 2.405 ;
      RECT 45.93 1.235 46.335 1.565 ;
      RECT 45.93 5.015 46.1 8.305 ;
      RECT 45.93 7.315 46.335 7.645 ;
      RECT 45.93 6.475 46.335 6.805 ;
      RECT 43.265 1.975 43.995 2.215 ;
      RECT 43.807 1.77 43.995 2.215 ;
      RECT 43.635 1.782 44.01 2.209 ;
      RECT 43.55 1.797 44.03 2.194 ;
      RECT 43.55 1.812 44.035 2.184 ;
      RECT 43.505 1.832 44.05 2.176 ;
      RECT 43.482 1.867 44.065 2.13 ;
      RECT 43.396 1.89 44.07 2.09 ;
      RECT 43.396 1.908 44.08 2.06 ;
      RECT 43.265 1.977 44.085 2.023 ;
      RECT 43.31 1.92 44.08 2.06 ;
      RECT 43.396 1.872 44.065 2.13 ;
      RECT 43.482 1.841 44.05 2.176 ;
      RECT 43.505 1.822 44.035 2.184 ;
      RECT 43.55 1.795 44.01 2.209 ;
      RECT 43.635 1.777 43.995 2.215 ;
      RECT 43.721 1.771 43.995 2.215 ;
      RECT 43.807 1.766 43.94 2.215 ;
      RECT 43.893 1.761 43.94 2.215 ;
      RECT 43.585 2.659 43.755 3.045 ;
      RECT 43.58 2.659 43.755 3.04 ;
      RECT 43.555 2.659 43.755 3.005 ;
      RECT 43.555 2.687 43.765 2.995 ;
      RECT 43.535 2.687 43.765 2.955 ;
      RECT 43.53 2.687 43.765 2.928 ;
      RECT 43.53 2.705 43.77 2.92 ;
      RECT 43.475 2.705 43.77 2.855 ;
      RECT 43.475 2.722 43.78 2.838 ;
      RECT 43.465 2.722 43.78 2.778 ;
      RECT 43.465 2.739 43.785 2.775 ;
      RECT 43.46 2.575 43.63 2.753 ;
      RECT 43.46 2.609 43.716 2.753 ;
      RECT 43.455 3.375 43.46 3.388 ;
      RECT 43.45 3.27 43.455 3.393 ;
      RECT 43.425 3.13 43.45 3.408 ;
      RECT 43.39 3.081 43.425 3.44 ;
      RECT 43.385 3.049 43.39 3.46 ;
      RECT 43.38 3.04 43.385 3.46 ;
      RECT 43.3 3.005 43.38 3.46 ;
      RECT 43.237 2.975 43.3 3.46 ;
      RECT 43.151 2.963 43.237 3.46 ;
      RECT 43.065 2.949 43.151 3.46 ;
      RECT 42.985 2.936 43.065 3.446 ;
      RECT 42.95 2.928 42.985 3.426 ;
      RECT 42.94 2.925 42.95 3.417 ;
      RECT 42.91 2.92 42.94 3.404 ;
      RECT 42.86 2.895 42.91 3.38 ;
      RECT 42.846 2.869 42.86 3.362 ;
      RECT 42.76 2.829 42.846 3.338 ;
      RECT 42.715 2.777 42.76 3.307 ;
      RECT 42.705 2.752 42.715 3.294 ;
      RECT 42.7 2.533 42.705 2.555 ;
      RECT 42.695 2.735 42.705 3.29 ;
      RECT 42.695 2.531 42.7 2.645 ;
      RECT 42.685 2.527 42.695 3.286 ;
      RECT 42.641 2.525 42.685 3.274 ;
      RECT 42.555 2.525 42.641 3.245 ;
      RECT 42.525 2.525 42.555 3.218 ;
      RECT 42.51 2.525 42.525 3.206 ;
      RECT 42.47 2.537 42.51 3.191 ;
      RECT 42.45 2.556 42.47 3.17 ;
      RECT 42.44 2.566 42.45 3.154 ;
      RECT 42.43 2.572 42.44 3.143 ;
      RECT 42.41 2.582 42.43 3.126 ;
      RECT 42.405 2.591 42.41 3.113 ;
      RECT 42.4 2.595 42.405 3.063 ;
      RECT 42.39 2.601 42.4 2.98 ;
      RECT 42.385 2.605 42.39 2.894 ;
      RECT 42.38 2.625 42.385 2.831 ;
      RECT 42.375 2.648 42.38 2.778 ;
      RECT 42.37 2.666 42.375 2.723 ;
      RECT 42.98 2.485 43.15 2.745 ;
      RECT 43.15 2.45 43.195 2.731 ;
      RECT 43.111 2.452 43.2 2.714 ;
      RECT 43 2.469 43.286 2.685 ;
      RECT 43 2.484 43.29 2.657 ;
      RECT 43 2.465 43.2 2.714 ;
      RECT 43.025 2.453 43.15 2.745 ;
      RECT 43.111 2.451 43.195 2.731 ;
      RECT 42.165 1.84 42.335 2.33 ;
      RECT 42.165 1.84 42.37 2.31 ;
      RECT 42.3 1.76 42.41 2.27 ;
      RECT 42.281 1.764 42.43 2.24 ;
      RECT 42.195 1.772 42.45 2.223 ;
      RECT 42.195 1.778 42.455 2.213 ;
      RECT 42.195 1.787 42.475 2.201 ;
      RECT 42.17 1.812 42.505 2.179 ;
      RECT 42.17 1.832 42.51 2.159 ;
      RECT 42.165 1.845 42.52 2.139 ;
      RECT 42.165 1.912 42.525 2.12 ;
      RECT 42.165 2.045 42.53 2.107 ;
      RECT 42.16 1.85 42.52 1.94 ;
      RECT 42.17 1.807 42.475 2.201 ;
      RECT 42.281 1.762 42.41 2.27 ;
      RECT 42.155 3.515 42.455 3.77 ;
      RECT 42.24 3.481 42.455 3.77 ;
      RECT 42.24 3.484 42.46 3.63 ;
      RECT 42.175 3.505 42.46 3.63 ;
      RECT 42.21 3.495 42.455 3.77 ;
      RECT 42.205 3.5 42.46 3.63 ;
      RECT 42.24 3.479 42.441 3.77 ;
      RECT 42.326 3.47 42.441 3.77 ;
      RECT 42.326 3.464 42.355 3.77 ;
      RECT 41.815 3.105 41.825 3.595 ;
      RECT 41.475 3.04 41.485 3.34 ;
      RECT 41.99 3.212 41.995 3.431 ;
      RECT 41.98 3.192 41.99 3.448 ;
      RECT 41.97 3.172 41.98 3.478 ;
      RECT 41.965 3.162 41.97 3.493 ;
      RECT 41.96 3.158 41.965 3.498 ;
      RECT 41.945 3.15 41.96 3.505 ;
      RECT 41.905 3.13 41.945 3.53 ;
      RECT 41.88 3.112 41.905 3.563 ;
      RECT 41.875 3.11 41.88 3.576 ;
      RECT 41.855 3.107 41.875 3.58 ;
      RECT 41.825 3.105 41.855 3.59 ;
      RECT 41.755 3.107 41.815 3.591 ;
      RECT 41.735 3.107 41.755 3.585 ;
      RECT 41.71 3.105 41.735 3.582 ;
      RECT 41.675 3.1 41.71 3.578 ;
      RECT 41.655 3.094 41.675 3.565 ;
      RECT 41.645 3.091 41.655 3.553 ;
      RECT 41.625 3.088 41.645 3.538 ;
      RECT 41.605 3.084 41.625 3.52 ;
      RECT 41.6 3.081 41.605 3.51 ;
      RECT 41.595 3.08 41.6 3.508 ;
      RECT 41.585 3.077 41.595 3.5 ;
      RECT 41.575 3.071 41.585 3.483 ;
      RECT 41.565 3.065 41.575 3.465 ;
      RECT 41.555 3.059 41.565 3.453 ;
      RECT 41.545 3.053 41.555 3.433 ;
      RECT 41.54 3.049 41.545 3.418 ;
      RECT 41.535 3.047 41.54 3.41 ;
      RECT 41.53 3.045 41.535 3.403 ;
      RECT 41.525 3.043 41.53 3.393 ;
      RECT 41.52 3.041 41.525 3.387 ;
      RECT 41.51 3.04 41.52 3.377 ;
      RECT 41.5 3.04 41.51 3.368 ;
      RECT 41.485 3.04 41.5 3.353 ;
      RECT 41.445 3.04 41.475 3.337 ;
      RECT 41.425 3.042 41.445 3.332 ;
      RECT 41.42 3.047 41.425 3.33 ;
      RECT 41.39 3.055 41.42 3.328 ;
      RECT 41.36 3.07 41.39 3.327 ;
      RECT 41.315 3.092 41.36 3.332 ;
      RECT 41.31 3.107 41.315 3.336 ;
      RECT 41.295 3.112 41.31 3.338 ;
      RECT 41.29 3.116 41.295 3.34 ;
      RECT 41.23 3.139 41.29 3.349 ;
      RECT 41.21 3.165 41.23 3.362 ;
      RECT 41.2 3.172 41.21 3.366 ;
      RECT 41.185 3.179 41.2 3.369 ;
      RECT 41.165 3.189 41.185 3.372 ;
      RECT 41.16 3.197 41.165 3.375 ;
      RECT 41.115 3.202 41.16 3.382 ;
      RECT 41.105 3.205 41.115 3.389 ;
      RECT 41.095 3.205 41.105 3.393 ;
      RECT 41.06 3.207 41.095 3.405 ;
      RECT 41.04 3.21 41.06 3.418 ;
      RECT 41 3.213 41.04 3.429 ;
      RECT 40.985 3.215 41 3.442 ;
      RECT 40.975 3.215 40.985 3.447 ;
      RECT 40.95 3.216 40.975 3.455 ;
      RECT 40.94 3.218 40.95 3.46 ;
      RECT 40.935 3.219 40.94 3.463 ;
      RECT 40.91 3.217 40.935 3.466 ;
      RECT 40.895 3.215 40.91 3.467 ;
      RECT 40.875 3.212 40.895 3.469 ;
      RECT 40.855 3.207 40.875 3.469 ;
      RECT 40.795 3.202 40.855 3.466 ;
      RECT 40.76 3.177 40.795 3.462 ;
      RECT 40.75 3.154 40.76 3.46 ;
      RECT 40.72 3.131 40.75 3.46 ;
      RECT 40.71 3.11 40.72 3.46 ;
      RECT 40.685 3.092 40.71 3.458 ;
      RECT 40.67 3.07 40.685 3.455 ;
      RECT 40.655 3.052 40.67 3.453 ;
      RECT 40.635 3.042 40.655 3.451 ;
      RECT 40.62 3.037 40.635 3.45 ;
      RECT 40.605 3.035 40.62 3.449 ;
      RECT 40.575 3.036 40.605 3.447 ;
      RECT 40.555 3.039 40.575 3.445 ;
      RECT 40.498 3.043 40.555 3.445 ;
      RECT 40.412 3.052 40.498 3.445 ;
      RECT 40.326 3.063 40.412 3.445 ;
      RECT 40.24 3.074 40.326 3.445 ;
      RECT 40.22 3.081 40.24 3.453 ;
      RECT 40.21 3.084 40.22 3.46 ;
      RECT 40.145 3.089 40.21 3.478 ;
      RECT 40.115 3.096 40.145 3.503 ;
      RECT 40.105 3.099 40.115 3.51 ;
      RECT 40.06 3.103 40.105 3.515 ;
      RECT 40.03 3.108 40.06 3.52 ;
      RECT 40.029 3.11 40.03 3.52 ;
      RECT 39.943 3.116 40.029 3.52 ;
      RECT 39.857 3.127 39.943 3.52 ;
      RECT 39.771 3.139 39.857 3.52 ;
      RECT 39.685 3.15 39.771 3.52 ;
      RECT 39.67 3.157 39.685 3.515 ;
      RECT 39.665 3.159 39.67 3.509 ;
      RECT 39.645 3.17 39.665 3.504 ;
      RECT 39.635 3.188 39.645 3.498 ;
      RECT 39.63 3.2 39.635 3.298 ;
      RECT 41.925 1.953 41.945 2.04 ;
      RECT 41.92 1.888 41.925 2.072 ;
      RECT 41.91 1.855 41.92 2.077 ;
      RECT 41.905 1.835 41.91 2.083 ;
      RECT 41.875 1.835 41.905 2.1 ;
      RECT 41.826 1.835 41.875 2.136 ;
      RECT 41.74 1.835 41.826 2.194 ;
      RECT 41.711 1.845 41.74 2.243 ;
      RECT 41.625 1.887 41.711 2.296 ;
      RECT 41.605 1.925 41.625 2.343 ;
      RECT 41.58 1.942 41.605 2.363 ;
      RECT 41.57 1.956 41.58 2.383 ;
      RECT 41.565 1.962 41.57 2.393 ;
      RECT 41.56 1.966 41.565 2.4 ;
      RECT 41.51 1.986 41.56 2.405 ;
      RECT 41.445 2.03 41.51 2.405 ;
      RECT 41.42 2.08 41.445 2.405 ;
      RECT 41.41 2.11 41.42 2.405 ;
      RECT 41.405 2.137 41.41 2.405 ;
      RECT 41.4 2.155 41.405 2.405 ;
      RECT 41.39 2.197 41.4 2.405 ;
      RECT 41.74 2.755 41.91 2.93 ;
      RECT 41.68 2.583 41.74 2.918 ;
      RECT 41.67 2.576 41.68 2.901 ;
      RECT 41.625 2.755 41.91 2.881 ;
      RECT 41.606 2.755 41.91 2.859 ;
      RECT 41.52 2.755 41.91 2.824 ;
      RECT 41.5 2.575 41.67 2.78 ;
      RECT 41.5 2.722 41.905 2.78 ;
      RECT 41.5 2.67 41.88 2.78 ;
      RECT 41.5 2.625 41.845 2.78 ;
      RECT 41.5 2.607 41.81 2.78 ;
      RECT 41.5 2.597 41.805 2.78 ;
      RECT 41.67 7.855 41.84 8.305 ;
      RECT 41.725 6.075 41.895 8.025 ;
      RECT 41.67 5.015 41.84 6.245 ;
      RECT 41.15 5.015 41.32 8.305 ;
      RECT 41.15 7.315 41.555 7.645 ;
      RECT 41.15 6.475 41.555 6.805 ;
      RECT 41.22 3.555 41.41 3.78 ;
      RECT 41.21 3.556 41.415 3.775 ;
      RECT 41.21 3.558 41.425 3.755 ;
      RECT 41.21 3.562 41.43 3.74 ;
      RECT 41.21 3.549 41.38 3.775 ;
      RECT 41.21 3.552 41.405 3.775 ;
      RECT 41.22 3.548 41.38 3.78 ;
      RECT 41.306 3.546 41.38 3.78 ;
      RECT 40.93 2.797 41.1 3.035 ;
      RECT 40.93 2.797 41.186 2.949 ;
      RECT 40.93 2.797 41.19 2.859 ;
      RECT 40.98 2.57 41.2 2.838 ;
      RECT 40.975 2.587 41.205 2.811 ;
      RECT 40.94 2.745 41.205 2.811 ;
      RECT 40.96 2.595 41.1 3.035 ;
      RECT 40.95 2.677 41.21 2.794 ;
      RECT 40.945 2.725 41.21 2.794 ;
      RECT 40.95 2.635 41.205 2.811 ;
      RECT 40.975 2.572 41.2 2.838 ;
      RECT 40.54 2.547 40.71 2.745 ;
      RECT 40.54 2.547 40.755 2.72 ;
      RECT 40.61 2.49 40.78 2.678 ;
      RECT 40.585 2.505 40.78 2.678 ;
      RECT 40.2 2.551 40.23 2.745 ;
      RECT 40.195 2.523 40.2 2.745 ;
      RECT 40.165 2.497 40.195 2.747 ;
      RECT 40.14 2.455 40.165 2.75 ;
      RECT 40.13 2.427 40.14 2.752 ;
      RECT 40.095 2.407 40.13 2.754 ;
      RECT 40.03 2.392 40.095 2.76 ;
      RECT 39.98 2.39 40.03 2.766 ;
      RECT 39.957 2.392 39.98 2.771 ;
      RECT 39.871 2.403 39.957 2.777 ;
      RECT 39.785 2.421 39.871 2.787 ;
      RECT 39.77 2.432 39.785 2.793 ;
      RECT 39.7 2.455 39.77 2.799 ;
      RECT 39.645 2.487 39.7 2.807 ;
      RECT 39.605 2.51 39.645 2.813 ;
      RECT 39.591 2.523 39.605 2.816 ;
      RECT 39.505 2.545 39.591 2.822 ;
      RECT 39.49 2.57 39.505 2.828 ;
      RECT 39.45 2.585 39.49 2.832 ;
      RECT 39.4 2.6 39.45 2.837 ;
      RECT 39.375 2.607 39.4 2.841 ;
      RECT 39.315 2.602 39.375 2.845 ;
      RECT 39.3 2.593 39.315 2.849 ;
      RECT 39.23 2.583 39.3 2.845 ;
      RECT 39.205 2.575 39.225 2.835 ;
      RECT 39.146 2.575 39.205 2.813 ;
      RECT 39.06 2.575 39.146 2.77 ;
      RECT 39.225 2.575 39.23 2.84 ;
      RECT 39.92 1.806 40.09 2.14 ;
      RECT 39.89 1.806 40.09 2.135 ;
      RECT 39.83 1.773 39.89 2.123 ;
      RECT 39.83 1.829 40.1 2.118 ;
      RECT 39.805 1.829 40.1 2.112 ;
      RECT 39.8 1.77 39.83 2.109 ;
      RECT 39.785 1.776 39.92 2.107 ;
      RECT 39.78 1.784 40.005 2.095 ;
      RECT 39.78 1.836 40.115 2.048 ;
      RECT 39.765 1.792 40.005 2.043 ;
      RECT 39.765 1.862 40.125 1.984 ;
      RECT 39.735 1.812 40.09 1.945 ;
      RECT 39.735 1.902 40.135 1.941 ;
      RECT 39.785 1.781 40.005 2.107 ;
      RECT 39.125 2.111 39.18 2.375 ;
      RECT 39.125 2.111 39.245 2.374 ;
      RECT 39.125 2.111 39.27 2.373 ;
      RECT 39.125 2.111 39.335 2.372 ;
      RECT 39.27 2.077 39.35 2.371 ;
      RECT 39.085 2.121 39.495 2.37 ;
      RECT 39.125 2.118 39.495 2.37 ;
      RECT 39.085 2.126 39.5 2.363 ;
      RECT 39.07 2.128 39.5 2.362 ;
      RECT 39.07 2.135 39.505 2.358 ;
      RECT 39.05 2.134 39.5 2.354 ;
      RECT 39.05 2.142 39.51 2.353 ;
      RECT 39.045 2.139 39.505 2.349 ;
      RECT 39.045 2.152 39.52 2.348 ;
      RECT 39.03 2.142 39.51 2.347 ;
      RECT 38.995 2.155 39.52 2.34 ;
      RECT 39.18 2.11 39.49 2.37 ;
      RECT 39.18 2.095 39.44 2.37 ;
      RECT 39.245 2.082 39.375 2.37 ;
      RECT 38.79 3.171 38.805 3.564 ;
      RECT 38.755 3.176 38.805 3.563 ;
      RECT 38.79 3.175 38.85 3.562 ;
      RECT 38.735 3.186 38.85 3.561 ;
      RECT 38.75 3.182 38.85 3.561 ;
      RECT 38.715 3.192 38.925 3.558 ;
      RECT 38.715 3.211 38.97 3.556 ;
      RECT 38.715 3.218 38.975 3.553 ;
      RECT 38.7 3.195 38.925 3.55 ;
      RECT 38.68 3.2 38.925 3.543 ;
      RECT 38.675 3.204 38.925 3.539 ;
      RECT 38.675 3.221 38.985 3.538 ;
      RECT 38.655 3.215 38.97 3.534 ;
      RECT 38.655 3.224 38.99 3.528 ;
      RECT 38.65 3.23 38.99 3.3 ;
      RECT 38.715 3.19 38.85 3.558 ;
      RECT 38.59 2.553 38.79 2.865 ;
      RECT 38.665 2.531 38.79 2.865 ;
      RECT 38.605 2.55 38.795 2.85 ;
      RECT 38.575 2.561 38.795 2.848 ;
      RECT 38.59 2.556 38.8 2.814 ;
      RECT 38.575 2.66 38.805 2.781 ;
      RECT 38.605 2.532 38.79 2.865 ;
      RECT 38.665 2.51 38.765 2.865 ;
      RECT 38.69 2.507 38.765 2.865 ;
      RECT 38.69 2.502 38.71 2.865 ;
      RECT 38.095 2.57 38.27 2.745 ;
      RECT 38.09 2.57 38.27 2.743 ;
      RECT 38.065 2.57 38.27 2.738 ;
      RECT 38.01 2.55 38.18 2.728 ;
      RECT 38.01 2.557 38.245 2.728 ;
      RECT 38.095 3.237 38.11 3.42 ;
      RECT 38.085 3.215 38.095 3.42 ;
      RECT 38.07 3.195 38.085 3.42 ;
      RECT 38.06 3.17 38.07 3.42 ;
      RECT 38.03 3.135 38.06 3.42 ;
      RECT 37.995 3.075 38.03 3.42 ;
      RECT 37.99 3.037 37.995 3.42 ;
      RECT 37.94 2.988 37.99 3.42 ;
      RECT 37.93 2.938 37.94 3.408 ;
      RECT 37.915 2.917 37.93 3.368 ;
      RECT 37.895 2.885 37.915 3.318 ;
      RECT 37.87 2.841 37.895 3.258 ;
      RECT 37.865 2.813 37.87 3.213 ;
      RECT 37.86 2.804 37.865 3.199 ;
      RECT 37.855 2.797 37.86 3.186 ;
      RECT 37.85 2.792 37.855 3.175 ;
      RECT 37.845 2.777 37.85 3.165 ;
      RECT 37.84 2.755 37.845 3.152 ;
      RECT 37.83 2.715 37.84 3.127 ;
      RECT 37.805 2.645 37.83 3.083 ;
      RECT 37.8 2.585 37.805 3.048 ;
      RECT 37.785 2.565 37.8 3.015 ;
      RECT 37.78 2.565 37.785 2.99 ;
      RECT 37.75 2.565 37.78 2.945 ;
      RECT 37.705 2.565 37.75 2.885 ;
      RECT 37.63 2.565 37.705 2.833 ;
      RECT 37.625 2.565 37.63 2.798 ;
      RECT 37.62 2.565 37.625 2.788 ;
      RECT 37.615 2.565 37.62 2.768 ;
      RECT 37.88 1.785 38.05 2.255 ;
      RECT 37.825 1.778 38.02 2.239 ;
      RECT 37.825 1.792 38.055 2.238 ;
      RECT 37.81 1.793 38.055 2.219 ;
      RECT 37.805 1.811 38.055 2.205 ;
      RECT 37.81 1.794 38.06 2.203 ;
      RECT 37.795 1.825 38.06 2.188 ;
      RECT 37.81 1.8 38.065 2.173 ;
      RECT 37.79 1.84 38.065 2.17 ;
      RECT 37.805 1.812 38.07 2.155 ;
      RECT 37.805 1.824 38.075 2.135 ;
      RECT 37.79 1.84 38.08 2.118 ;
      RECT 37.79 1.85 38.085 1.973 ;
      RECT 37.785 1.85 38.085 1.93 ;
      RECT 37.785 1.865 38.09 1.908 ;
      RECT 37.88 1.775 38.02 2.255 ;
      RECT 37.88 1.773 37.99 2.255 ;
      RECT 37.966 1.77 37.99 2.255 ;
      RECT 37.625 3.437 37.63 3.483 ;
      RECT 37.615 3.285 37.625 3.507 ;
      RECT 37.61 3.13 37.615 3.532 ;
      RECT 37.595 3.092 37.61 3.543 ;
      RECT 37.59 3.075 37.595 3.55 ;
      RECT 37.58 3.063 37.59 3.557 ;
      RECT 37.575 3.054 37.58 3.559 ;
      RECT 37.57 3.052 37.575 3.563 ;
      RECT 37.525 3.043 37.57 3.578 ;
      RECT 37.52 3.035 37.525 3.592 ;
      RECT 37.515 3.032 37.52 3.596 ;
      RECT 37.5 3.027 37.515 3.604 ;
      RECT 37.445 3.017 37.5 3.615 ;
      RECT 37.41 3.005 37.445 3.616 ;
      RECT 37.401 3 37.41 3.61 ;
      RECT 37.315 3 37.401 3.6 ;
      RECT 37.285 3 37.315 3.578 ;
      RECT 37.275 3 37.28 3.558 ;
      RECT 37.27 3 37.275 3.52 ;
      RECT 37.265 3 37.27 3.478 ;
      RECT 37.26 3 37.265 3.438 ;
      RECT 37.255 3 37.26 3.368 ;
      RECT 37.245 3 37.255 3.29 ;
      RECT 37.24 3 37.245 3.19 ;
      RECT 37.28 3 37.285 3.56 ;
      RECT 36.775 3.082 36.865 3.56 ;
      RECT 36.76 3.085 36.88 3.558 ;
      RECT 36.775 3.084 36.88 3.558 ;
      RECT 36.74 3.091 36.905 3.548 ;
      RECT 36.76 3.085 36.905 3.548 ;
      RECT 36.725 3.097 36.905 3.536 ;
      RECT 36.76 3.088 36.955 3.529 ;
      RECT 36.711 3.105 36.955 3.527 ;
      RECT 36.74 3.095 36.965 3.515 ;
      RECT 36.711 3.116 36.995 3.506 ;
      RECT 36.625 3.14 36.995 3.5 ;
      RECT 36.625 3.153 37.035 3.483 ;
      RECT 36.62 3.175 37.035 3.476 ;
      RECT 36.59 3.19 37.035 3.466 ;
      RECT 36.585 3.201 37.035 3.456 ;
      RECT 36.555 3.214 37.035 3.447 ;
      RECT 36.54 3.232 37.035 3.436 ;
      RECT 36.515 3.245 37.035 3.426 ;
      RECT 36.775 3.081 36.785 3.56 ;
      RECT 36.821 2.505 36.86 2.75 ;
      RECT 36.735 2.505 36.87 2.748 ;
      RECT 36.62 2.53 36.87 2.745 ;
      RECT 36.62 2.53 36.875 2.743 ;
      RECT 36.62 2.53 36.89 2.738 ;
      RECT 36.726 2.505 36.905 2.718 ;
      RECT 36.64 2.513 36.905 2.718 ;
      RECT 36.31 1.865 36.48 2.3 ;
      RECT 36.3 1.899 36.48 2.283 ;
      RECT 36.38 1.835 36.55 2.27 ;
      RECT 36.285 1.91 36.55 2.248 ;
      RECT 36.38 1.845 36.555 2.238 ;
      RECT 36.31 1.897 36.585 2.223 ;
      RECT 36.27 1.923 36.585 2.208 ;
      RECT 36.27 1.965 36.595 2.188 ;
      RECT 36.265 1.99 36.6 2.17 ;
      RECT 36.265 2 36.605 2.155 ;
      RECT 36.26 1.937 36.585 2.153 ;
      RECT 36.26 2.01 36.61 2.138 ;
      RECT 36.255 1.947 36.585 2.135 ;
      RECT 36.25 2.031 36.615 2.118 ;
      RECT 36.25 2.063 36.62 2.098 ;
      RECT 36.245 1.977 36.595 2.09 ;
      RECT 36.25 1.962 36.585 2.118 ;
      RECT 36.265 1.932 36.585 2.17 ;
      RECT 36.11 2.519 36.335 2.775 ;
      RECT 36.11 2.552 36.355 2.765 ;
      RECT 36.075 2.552 36.355 2.763 ;
      RECT 36.075 2.565 36.36 2.753 ;
      RECT 36.075 2.585 36.37 2.745 ;
      RECT 36.075 2.682 36.375 2.738 ;
      RECT 36.055 2.43 36.185 2.728 ;
      RECT 36.01 2.585 36.37 2.67 ;
      RECT 36 2.43 36.185 2.615 ;
      RECT 36 2.462 36.271 2.615 ;
      RECT 35.965 2.992 35.985 3.17 ;
      RECT 35.93 2.945 35.965 3.17 ;
      RECT 35.915 2.885 35.93 3.17 ;
      RECT 35.89 2.832 35.915 3.17 ;
      RECT 35.875 2.785 35.89 3.17 ;
      RECT 35.855 2.762 35.875 3.17 ;
      RECT 35.83 2.727 35.855 3.17 ;
      RECT 35.82 2.573 35.83 3.17 ;
      RECT 35.79 2.568 35.82 3.161 ;
      RECT 35.785 2.565 35.79 3.151 ;
      RECT 35.77 2.565 35.785 3.125 ;
      RECT 35.765 2.565 35.77 3.088 ;
      RECT 35.74 2.565 35.765 3.04 ;
      RECT 35.72 2.565 35.74 2.965 ;
      RECT 35.71 2.565 35.72 2.925 ;
      RECT 35.705 2.565 35.71 2.9 ;
      RECT 35.7 2.565 35.705 2.883 ;
      RECT 35.695 2.565 35.7 2.865 ;
      RECT 35.69 2.566 35.695 2.855 ;
      RECT 35.68 2.568 35.69 2.823 ;
      RECT 35.67 2.57 35.68 2.79 ;
      RECT 35.66 2.573 35.67 2.763 ;
      RECT 35.985 3 36.21 3.17 ;
      RECT 35.315 1.812 35.485 2.265 ;
      RECT 35.315 1.812 35.575 2.231 ;
      RECT 35.315 1.812 35.605 2.215 ;
      RECT 35.315 1.812 35.635 2.188 ;
      RECT 35.571 1.79 35.65 2.17 ;
      RECT 35.35 1.797 35.655 2.155 ;
      RECT 35.35 1.805 35.665 2.118 ;
      RECT 35.31 1.832 35.665 2.09 ;
      RECT 35.295 1.845 35.665 2.055 ;
      RECT 35.315 1.82 35.685 2.045 ;
      RECT 35.29 1.885 35.685 2.015 ;
      RECT 35.29 1.915 35.69 1.998 ;
      RECT 35.285 1.945 35.69 1.985 ;
      RECT 35.35 1.794 35.65 2.17 ;
      RECT 35.485 1.791 35.571 2.249 ;
      RECT 35.436 1.792 35.65 2.17 ;
      RECT 35.58 3.452 35.625 3.645 ;
      RECT 35.57 3.422 35.58 3.645 ;
      RECT 35.565 3.407 35.57 3.645 ;
      RECT 35.525 3.317 35.565 3.645 ;
      RECT 35.52 3.23 35.525 3.645 ;
      RECT 35.51 3.2 35.52 3.645 ;
      RECT 35.505 3.16 35.51 3.645 ;
      RECT 35.495 3.122 35.505 3.645 ;
      RECT 35.49 3.087 35.495 3.645 ;
      RECT 35.47 3.04 35.49 3.645 ;
      RECT 35.455 2.965 35.47 3.645 ;
      RECT 35.45 2.92 35.455 3.64 ;
      RECT 35.445 2.9 35.45 3.613 ;
      RECT 35.44 2.88 35.445 3.598 ;
      RECT 35.435 2.855 35.44 3.578 ;
      RECT 35.43 2.833 35.435 3.563 ;
      RECT 35.425 2.811 35.43 3.545 ;
      RECT 35.42 2.79 35.425 3.535 ;
      RECT 35.41 2.762 35.42 3.505 ;
      RECT 35.4 2.725 35.41 3.473 ;
      RECT 35.39 2.685 35.4 3.44 ;
      RECT 35.38 2.663 35.39 3.41 ;
      RECT 35.35 2.615 35.38 3.342 ;
      RECT 35.335 2.575 35.35 3.269 ;
      RECT 35.325 2.575 35.335 3.235 ;
      RECT 35.32 2.575 35.325 3.21 ;
      RECT 35.315 2.575 35.32 3.195 ;
      RECT 35.31 2.575 35.315 3.173 ;
      RECT 35.305 2.575 35.31 3.16 ;
      RECT 35.29 2.575 35.305 3.125 ;
      RECT 35.27 2.575 35.29 3.065 ;
      RECT 35.26 2.575 35.27 3.015 ;
      RECT 35.24 2.575 35.26 2.963 ;
      RECT 35.22 2.575 35.24 2.92 ;
      RECT 35.21 2.575 35.22 2.908 ;
      RECT 35.18 2.575 35.21 2.895 ;
      RECT 35.15 2.596 35.18 2.875 ;
      RECT 35.14 2.624 35.15 2.855 ;
      RECT 35.125 2.641 35.14 2.823 ;
      RECT 35.12 2.655 35.125 2.79 ;
      RECT 35.115 2.663 35.12 2.763 ;
      RECT 35.11 2.671 35.115 2.725 ;
      RECT 35.115 3.195 35.12 3.53 ;
      RECT 35.08 3.182 35.115 3.529 ;
      RECT 35.01 3.122 35.08 3.528 ;
      RECT 34.93 3.065 35.01 3.527 ;
      RECT 34.795 3.025 34.93 3.526 ;
      RECT 34.795 3.212 35.13 3.515 ;
      RECT 34.755 3.212 35.13 3.505 ;
      RECT 34.755 3.23 35.135 3.5 ;
      RECT 34.755 3.32 35.14 3.49 ;
      RECT 34.75 3.015 34.915 3.47 ;
      RECT 34.745 3.015 34.915 3.213 ;
      RECT 34.745 3.172 35.11 3.213 ;
      RECT 34.745 3.16 35.105 3.213 ;
      RECT 33.885 5.02 34.055 6.49 ;
      RECT 33.885 6.315 34.06 6.485 ;
      RECT 33.515 1.74 33.685 2.93 ;
      RECT 33.515 1.74 33.985 1.91 ;
      RECT 33.515 6.97 33.985 7.14 ;
      RECT 33.515 5.95 33.685 7.14 ;
      RECT 32.525 1.74 32.695 2.93 ;
      RECT 32.525 1.74 32.995 1.91 ;
      RECT 32.525 6.97 32.995 7.14 ;
      RECT 32.525 5.95 32.695 7.14 ;
      RECT 30.675 2.635 30.845 3.865 ;
      RECT 30.73 0.855 30.9 2.805 ;
      RECT 30.675 0.575 30.845 1.025 ;
      RECT 30.675 7.855 30.845 8.305 ;
      RECT 30.73 6.075 30.9 8.025 ;
      RECT 30.675 5.015 30.845 6.245 ;
      RECT 30.155 0.575 30.325 3.865 ;
      RECT 30.155 2.075 30.56 2.405 ;
      RECT 30.155 1.235 30.56 1.565 ;
      RECT 30.155 5.015 30.325 8.305 ;
      RECT 30.155 7.315 30.56 7.645 ;
      RECT 30.155 6.475 30.56 6.805 ;
      RECT 27.49 1.975 28.22 2.215 ;
      RECT 28.032 1.77 28.22 2.215 ;
      RECT 27.86 1.782 28.235 2.209 ;
      RECT 27.775 1.797 28.255 2.194 ;
      RECT 27.775 1.812 28.26 2.184 ;
      RECT 27.73 1.832 28.275 2.176 ;
      RECT 27.707 1.867 28.29 2.13 ;
      RECT 27.621 1.89 28.295 2.09 ;
      RECT 27.621 1.908 28.305 2.06 ;
      RECT 27.49 1.977 28.31 2.023 ;
      RECT 27.535 1.92 28.305 2.06 ;
      RECT 27.621 1.872 28.29 2.13 ;
      RECT 27.707 1.841 28.275 2.176 ;
      RECT 27.73 1.822 28.26 2.184 ;
      RECT 27.775 1.795 28.235 2.209 ;
      RECT 27.86 1.777 28.22 2.215 ;
      RECT 27.946 1.771 28.22 2.215 ;
      RECT 28.032 1.766 28.165 2.215 ;
      RECT 28.118 1.761 28.165 2.215 ;
      RECT 27.81 2.659 27.98 3.045 ;
      RECT 27.805 2.659 27.98 3.04 ;
      RECT 27.78 2.659 27.98 3.005 ;
      RECT 27.78 2.687 27.99 2.995 ;
      RECT 27.76 2.687 27.99 2.955 ;
      RECT 27.755 2.687 27.99 2.928 ;
      RECT 27.755 2.705 27.995 2.92 ;
      RECT 27.7 2.705 27.995 2.855 ;
      RECT 27.7 2.722 28.005 2.838 ;
      RECT 27.69 2.722 28.005 2.778 ;
      RECT 27.69 2.739 28.01 2.775 ;
      RECT 27.685 2.575 27.855 2.753 ;
      RECT 27.685 2.609 27.941 2.753 ;
      RECT 27.68 3.375 27.685 3.388 ;
      RECT 27.675 3.27 27.68 3.393 ;
      RECT 27.65 3.13 27.675 3.408 ;
      RECT 27.615 3.081 27.65 3.44 ;
      RECT 27.61 3.049 27.615 3.46 ;
      RECT 27.605 3.04 27.61 3.46 ;
      RECT 27.525 3.005 27.605 3.46 ;
      RECT 27.462 2.975 27.525 3.46 ;
      RECT 27.376 2.963 27.462 3.46 ;
      RECT 27.29 2.949 27.376 3.46 ;
      RECT 27.21 2.936 27.29 3.446 ;
      RECT 27.175 2.928 27.21 3.426 ;
      RECT 27.165 2.925 27.175 3.417 ;
      RECT 27.135 2.92 27.165 3.404 ;
      RECT 27.085 2.895 27.135 3.38 ;
      RECT 27.071 2.869 27.085 3.362 ;
      RECT 26.985 2.829 27.071 3.338 ;
      RECT 26.94 2.777 26.985 3.307 ;
      RECT 26.93 2.752 26.94 3.294 ;
      RECT 26.925 2.533 26.93 2.555 ;
      RECT 26.92 2.735 26.93 3.29 ;
      RECT 26.92 2.531 26.925 2.645 ;
      RECT 26.91 2.527 26.92 3.286 ;
      RECT 26.866 2.525 26.91 3.274 ;
      RECT 26.78 2.525 26.866 3.245 ;
      RECT 26.75 2.525 26.78 3.218 ;
      RECT 26.735 2.525 26.75 3.206 ;
      RECT 26.695 2.537 26.735 3.191 ;
      RECT 26.675 2.556 26.695 3.17 ;
      RECT 26.665 2.566 26.675 3.154 ;
      RECT 26.655 2.572 26.665 3.143 ;
      RECT 26.635 2.582 26.655 3.126 ;
      RECT 26.63 2.591 26.635 3.113 ;
      RECT 26.625 2.595 26.63 3.063 ;
      RECT 26.615 2.601 26.625 2.98 ;
      RECT 26.61 2.605 26.615 2.894 ;
      RECT 26.605 2.625 26.61 2.831 ;
      RECT 26.6 2.648 26.605 2.778 ;
      RECT 26.595 2.666 26.6 2.723 ;
      RECT 27.205 2.485 27.375 2.745 ;
      RECT 27.375 2.45 27.42 2.731 ;
      RECT 27.336 2.452 27.425 2.714 ;
      RECT 27.225 2.469 27.511 2.685 ;
      RECT 27.225 2.484 27.515 2.657 ;
      RECT 27.225 2.465 27.425 2.714 ;
      RECT 27.25 2.453 27.375 2.745 ;
      RECT 27.336 2.451 27.42 2.731 ;
      RECT 26.39 1.84 26.56 2.33 ;
      RECT 26.39 1.84 26.595 2.31 ;
      RECT 26.525 1.76 26.635 2.27 ;
      RECT 26.506 1.764 26.655 2.24 ;
      RECT 26.42 1.772 26.675 2.223 ;
      RECT 26.42 1.778 26.68 2.213 ;
      RECT 26.42 1.787 26.7 2.201 ;
      RECT 26.395 1.812 26.73 2.179 ;
      RECT 26.395 1.832 26.735 2.159 ;
      RECT 26.39 1.845 26.745 2.139 ;
      RECT 26.39 1.912 26.75 2.12 ;
      RECT 26.39 2.045 26.755 2.107 ;
      RECT 26.385 1.85 26.745 1.94 ;
      RECT 26.395 1.807 26.7 2.201 ;
      RECT 26.506 1.762 26.635 2.27 ;
      RECT 26.38 3.515 26.68 3.77 ;
      RECT 26.465 3.481 26.68 3.77 ;
      RECT 26.465 3.484 26.685 3.63 ;
      RECT 26.4 3.505 26.685 3.63 ;
      RECT 26.435 3.495 26.68 3.77 ;
      RECT 26.43 3.5 26.685 3.63 ;
      RECT 26.465 3.479 26.666 3.77 ;
      RECT 26.551 3.47 26.666 3.77 ;
      RECT 26.551 3.464 26.58 3.77 ;
      RECT 26.04 3.105 26.05 3.595 ;
      RECT 25.7 3.04 25.71 3.34 ;
      RECT 26.215 3.212 26.22 3.431 ;
      RECT 26.205 3.192 26.215 3.448 ;
      RECT 26.195 3.172 26.205 3.478 ;
      RECT 26.19 3.162 26.195 3.493 ;
      RECT 26.185 3.158 26.19 3.498 ;
      RECT 26.17 3.15 26.185 3.505 ;
      RECT 26.13 3.13 26.17 3.53 ;
      RECT 26.105 3.112 26.13 3.563 ;
      RECT 26.1 3.11 26.105 3.576 ;
      RECT 26.08 3.107 26.1 3.58 ;
      RECT 26.05 3.105 26.08 3.59 ;
      RECT 25.98 3.107 26.04 3.591 ;
      RECT 25.96 3.107 25.98 3.585 ;
      RECT 25.935 3.105 25.96 3.582 ;
      RECT 25.9 3.1 25.935 3.578 ;
      RECT 25.88 3.094 25.9 3.565 ;
      RECT 25.87 3.091 25.88 3.553 ;
      RECT 25.85 3.088 25.87 3.538 ;
      RECT 25.83 3.084 25.85 3.52 ;
      RECT 25.825 3.081 25.83 3.51 ;
      RECT 25.82 3.08 25.825 3.508 ;
      RECT 25.81 3.077 25.82 3.5 ;
      RECT 25.8 3.071 25.81 3.483 ;
      RECT 25.79 3.065 25.8 3.465 ;
      RECT 25.78 3.059 25.79 3.453 ;
      RECT 25.77 3.053 25.78 3.433 ;
      RECT 25.765 3.049 25.77 3.418 ;
      RECT 25.76 3.047 25.765 3.41 ;
      RECT 25.755 3.045 25.76 3.403 ;
      RECT 25.75 3.043 25.755 3.393 ;
      RECT 25.745 3.041 25.75 3.387 ;
      RECT 25.735 3.04 25.745 3.377 ;
      RECT 25.725 3.04 25.735 3.368 ;
      RECT 25.71 3.04 25.725 3.353 ;
      RECT 25.67 3.04 25.7 3.337 ;
      RECT 25.65 3.042 25.67 3.332 ;
      RECT 25.645 3.047 25.65 3.33 ;
      RECT 25.615 3.055 25.645 3.328 ;
      RECT 25.585 3.07 25.615 3.327 ;
      RECT 25.54 3.092 25.585 3.332 ;
      RECT 25.535 3.107 25.54 3.336 ;
      RECT 25.52 3.112 25.535 3.338 ;
      RECT 25.515 3.116 25.52 3.34 ;
      RECT 25.455 3.139 25.515 3.349 ;
      RECT 25.435 3.165 25.455 3.362 ;
      RECT 25.425 3.172 25.435 3.366 ;
      RECT 25.41 3.179 25.425 3.369 ;
      RECT 25.39 3.189 25.41 3.372 ;
      RECT 25.385 3.197 25.39 3.375 ;
      RECT 25.34 3.202 25.385 3.382 ;
      RECT 25.33 3.205 25.34 3.389 ;
      RECT 25.32 3.205 25.33 3.393 ;
      RECT 25.285 3.207 25.32 3.405 ;
      RECT 25.265 3.21 25.285 3.418 ;
      RECT 25.225 3.213 25.265 3.429 ;
      RECT 25.21 3.215 25.225 3.442 ;
      RECT 25.2 3.215 25.21 3.447 ;
      RECT 25.175 3.216 25.2 3.455 ;
      RECT 25.165 3.218 25.175 3.46 ;
      RECT 25.16 3.219 25.165 3.463 ;
      RECT 25.135 3.217 25.16 3.466 ;
      RECT 25.12 3.215 25.135 3.467 ;
      RECT 25.1 3.212 25.12 3.469 ;
      RECT 25.08 3.207 25.1 3.469 ;
      RECT 25.02 3.202 25.08 3.466 ;
      RECT 24.985 3.177 25.02 3.462 ;
      RECT 24.975 3.154 24.985 3.46 ;
      RECT 24.945 3.131 24.975 3.46 ;
      RECT 24.935 3.11 24.945 3.46 ;
      RECT 24.91 3.092 24.935 3.458 ;
      RECT 24.895 3.07 24.91 3.455 ;
      RECT 24.88 3.052 24.895 3.453 ;
      RECT 24.86 3.042 24.88 3.451 ;
      RECT 24.845 3.037 24.86 3.45 ;
      RECT 24.83 3.035 24.845 3.449 ;
      RECT 24.8 3.036 24.83 3.447 ;
      RECT 24.78 3.039 24.8 3.445 ;
      RECT 24.723 3.043 24.78 3.445 ;
      RECT 24.637 3.052 24.723 3.445 ;
      RECT 24.551 3.063 24.637 3.445 ;
      RECT 24.465 3.074 24.551 3.445 ;
      RECT 24.445 3.081 24.465 3.453 ;
      RECT 24.435 3.084 24.445 3.46 ;
      RECT 24.37 3.089 24.435 3.478 ;
      RECT 24.34 3.096 24.37 3.503 ;
      RECT 24.33 3.099 24.34 3.51 ;
      RECT 24.285 3.103 24.33 3.515 ;
      RECT 24.255 3.108 24.285 3.52 ;
      RECT 24.254 3.11 24.255 3.52 ;
      RECT 24.168 3.116 24.254 3.52 ;
      RECT 24.082 3.127 24.168 3.52 ;
      RECT 23.996 3.139 24.082 3.52 ;
      RECT 23.91 3.15 23.996 3.52 ;
      RECT 23.895 3.157 23.91 3.515 ;
      RECT 23.89 3.159 23.895 3.509 ;
      RECT 23.87 3.17 23.89 3.504 ;
      RECT 23.86 3.188 23.87 3.498 ;
      RECT 23.855 3.2 23.86 3.298 ;
      RECT 26.15 1.953 26.17 2.04 ;
      RECT 26.145 1.888 26.15 2.072 ;
      RECT 26.135 1.855 26.145 2.077 ;
      RECT 26.13 1.835 26.135 2.083 ;
      RECT 26.1 1.835 26.13 2.1 ;
      RECT 26.051 1.835 26.1 2.136 ;
      RECT 25.965 1.835 26.051 2.194 ;
      RECT 25.936 1.845 25.965 2.243 ;
      RECT 25.85 1.887 25.936 2.296 ;
      RECT 25.83 1.925 25.85 2.343 ;
      RECT 25.805 1.942 25.83 2.363 ;
      RECT 25.795 1.956 25.805 2.383 ;
      RECT 25.79 1.962 25.795 2.393 ;
      RECT 25.785 1.966 25.79 2.4 ;
      RECT 25.735 1.986 25.785 2.405 ;
      RECT 25.67 2.03 25.735 2.405 ;
      RECT 25.645 2.08 25.67 2.405 ;
      RECT 25.635 2.11 25.645 2.405 ;
      RECT 25.63 2.137 25.635 2.405 ;
      RECT 25.625 2.155 25.63 2.405 ;
      RECT 25.615 2.197 25.625 2.405 ;
      RECT 25.965 2.755 26.135 2.93 ;
      RECT 25.905 2.583 25.965 2.918 ;
      RECT 25.895 2.576 25.905 2.901 ;
      RECT 25.85 2.755 26.135 2.881 ;
      RECT 25.831 2.755 26.135 2.859 ;
      RECT 25.745 2.755 26.135 2.824 ;
      RECT 25.725 2.575 25.895 2.78 ;
      RECT 25.725 2.722 26.13 2.78 ;
      RECT 25.725 2.67 26.105 2.78 ;
      RECT 25.725 2.625 26.07 2.78 ;
      RECT 25.725 2.607 26.035 2.78 ;
      RECT 25.725 2.597 26.03 2.78 ;
      RECT 25.895 7.855 26.065 8.305 ;
      RECT 25.95 6.075 26.12 8.025 ;
      RECT 25.895 5.015 26.065 6.245 ;
      RECT 25.375 5.015 25.545 8.305 ;
      RECT 25.375 7.315 25.78 7.645 ;
      RECT 25.375 6.475 25.78 6.805 ;
      RECT 25.445 3.555 25.635 3.78 ;
      RECT 25.435 3.556 25.64 3.775 ;
      RECT 25.435 3.558 25.65 3.755 ;
      RECT 25.435 3.562 25.655 3.74 ;
      RECT 25.435 3.549 25.605 3.775 ;
      RECT 25.435 3.552 25.63 3.775 ;
      RECT 25.445 3.548 25.605 3.78 ;
      RECT 25.531 3.546 25.605 3.78 ;
      RECT 25.155 2.797 25.325 3.035 ;
      RECT 25.155 2.797 25.411 2.949 ;
      RECT 25.155 2.797 25.415 2.859 ;
      RECT 25.205 2.57 25.425 2.838 ;
      RECT 25.2 2.587 25.43 2.811 ;
      RECT 25.165 2.745 25.43 2.811 ;
      RECT 25.185 2.595 25.325 3.035 ;
      RECT 25.175 2.677 25.435 2.794 ;
      RECT 25.17 2.725 25.435 2.794 ;
      RECT 25.175 2.635 25.43 2.811 ;
      RECT 25.2 2.572 25.425 2.838 ;
      RECT 24.765 2.547 24.935 2.745 ;
      RECT 24.765 2.547 24.98 2.72 ;
      RECT 24.835 2.49 25.005 2.678 ;
      RECT 24.81 2.505 25.005 2.678 ;
      RECT 24.425 2.551 24.455 2.745 ;
      RECT 24.42 2.523 24.425 2.745 ;
      RECT 24.39 2.497 24.42 2.747 ;
      RECT 24.365 2.455 24.39 2.75 ;
      RECT 24.355 2.427 24.365 2.752 ;
      RECT 24.32 2.407 24.355 2.754 ;
      RECT 24.255 2.392 24.32 2.76 ;
      RECT 24.205 2.39 24.255 2.766 ;
      RECT 24.182 2.392 24.205 2.771 ;
      RECT 24.096 2.403 24.182 2.777 ;
      RECT 24.01 2.421 24.096 2.787 ;
      RECT 23.995 2.432 24.01 2.793 ;
      RECT 23.925 2.455 23.995 2.799 ;
      RECT 23.87 2.487 23.925 2.807 ;
      RECT 23.83 2.51 23.87 2.813 ;
      RECT 23.816 2.523 23.83 2.816 ;
      RECT 23.73 2.545 23.816 2.822 ;
      RECT 23.715 2.57 23.73 2.828 ;
      RECT 23.675 2.585 23.715 2.832 ;
      RECT 23.625 2.6 23.675 2.837 ;
      RECT 23.6 2.607 23.625 2.841 ;
      RECT 23.54 2.602 23.6 2.845 ;
      RECT 23.525 2.593 23.54 2.849 ;
      RECT 23.455 2.583 23.525 2.845 ;
      RECT 23.43 2.575 23.45 2.835 ;
      RECT 23.371 2.575 23.43 2.813 ;
      RECT 23.285 2.575 23.371 2.77 ;
      RECT 23.45 2.575 23.455 2.84 ;
      RECT 24.145 1.806 24.315 2.14 ;
      RECT 24.115 1.806 24.315 2.135 ;
      RECT 24.055 1.773 24.115 2.123 ;
      RECT 24.055 1.829 24.325 2.118 ;
      RECT 24.03 1.829 24.325 2.112 ;
      RECT 24.025 1.77 24.055 2.109 ;
      RECT 24.01 1.776 24.145 2.107 ;
      RECT 24.005 1.784 24.23 2.095 ;
      RECT 24.005 1.836 24.34 2.048 ;
      RECT 23.99 1.792 24.23 2.043 ;
      RECT 23.99 1.862 24.35 1.984 ;
      RECT 23.96 1.812 24.315 1.945 ;
      RECT 23.96 1.902 24.36 1.941 ;
      RECT 24.01 1.781 24.23 2.107 ;
      RECT 23.35 2.111 23.405 2.375 ;
      RECT 23.35 2.111 23.47 2.374 ;
      RECT 23.35 2.111 23.495 2.373 ;
      RECT 23.35 2.111 23.56 2.372 ;
      RECT 23.495 2.077 23.575 2.371 ;
      RECT 23.31 2.121 23.72 2.37 ;
      RECT 23.35 2.118 23.72 2.37 ;
      RECT 23.31 2.126 23.725 2.363 ;
      RECT 23.295 2.128 23.725 2.362 ;
      RECT 23.295 2.135 23.73 2.358 ;
      RECT 23.275 2.134 23.725 2.354 ;
      RECT 23.275 2.142 23.735 2.353 ;
      RECT 23.27 2.139 23.73 2.349 ;
      RECT 23.27 2.152 23.745 2.348 ;
      RECT 23.255 2.142 23.735 2.347 ;
      RECT 23.22 2.155 23.745 2.34 ;
      RECT 23.405 2.11 23.715 2.37 ;
      RECT 23.405 2.095 23.665 2.37 ;
      RECT 23.47 2.082 23.6 2.37 ;
      RECT 23.015 3.171 23.03 3.564 ;
      RECT 22.98 3.176 23.03 3.563 ;
      RECT 23.015 3.175 23.075 3.562 ;
      RECT 22.96 3.186 23.075 3.561 ;
      RECT 22.975 3.182 23.075 3.561 ;
      RECT 22.94 3.192 23.15 3.558 ;
      RECT 22.94 3.211 23.195 3.556 ;
      RECT 22.94 3.218 23.2 3.553 ;
      RECT 22.925 3.195 23.15 3.55 ;
      RECT 22.905 3.2 23.15 3.543 ;
      RECT 22.9 3.204 23.15 3.539 ;
      RECT 22.9 3.221 23.21 3.538 ;
      RECT 22.88 3.215 23.195 3.534 ;
      RECT 22.88 3.224 23.215 3.528 ;
      RECT 22.875 3.23 23.215 3.3 ;
      RECT 22.94 3.19 23.075 3.558 ;
      RECT 22.815 2.553 23.015 2.865 ;
      RECT 22.89 2.531 23.015 2.865 ;
      RECT 22.83 2.55 23.02 2.85 ;
      RECT 22.8 2.561 23.02 2.848 ;
      RECT 22.815 2.556 23.025 2.814 ;
      RECT 22.8 2.66 23.03 2.781 ;
      RECT 22.83 2.532 23.015 2.865 ;
      RECT 22.89 2.51 22.99 2.865 ;
      RECT 22.915 2.507 22.99 2.865 ;
      RECT 22.915 2.502 22.935 2.865 ;
      RECT 22.32 2.57 22.495 2.745 ;
      RECT 22.315 2.57 22.495 2.743 ;
      RECT 22.29 2.57 22.495 2.738 ;
      RECT 22.235 2.55 22.405 2.728 ;
      RECT 22.235 2.557 22.47 2.728 ;
      RECT 22.32 3.237 22.335 3.42 ;
      RECT 22.31 3.215 22.32 3.42 ;
      RECT 22.295 3.195 22.31 3.42 ;
      RECT 22.285 3.17 22.295 3.42 ;
      RECT 22.255 3.135 22.285 3.42 ;
      RECT 22.22 3.075 22.255 3.42 ;
      RECT 22.215 3.037 22.22 3.42 ;
      RECT 22.165 2.988 22.215 3.42 ;
      RECT 22.155 2.938 22.165 3.408 ;
      RECT 22.14 2.917 22.155 3.368 ;
      RECT 22.12 2.885 22.14 3.318 ;
      RECT 22.095 2.841 22.12 3.258 ;
      RECT 22.09 2.813 22.095 3.213 ;
      RECT 22.085 2.804 22.09 3.199 ;
      RECT 22.08 2.797 22.085 3.186 ;
      RECT 22.075 2.792 22.08 3.175 ;
      RECT 22.07 2.777 22.075 3.165 ;
      RECT 22.065 2.755 22.07 3.152 ;
      RECT 22.055 2.715 22.065 3.127 ;
      RECT 22.03 2.645 22.055 3.083 ;
      RECT 22.025 2.585 22.03 3.048 ;
      RECT 22.01 2.565 22.025 3.015 ;
      RECT 22.005 2.565 22.01 2.99 ;
      RECT 21.975 2.565 22.005 2.945 ;
      RECT 21.93 2.565 21.975 2.885 ;
      RECT 21.855 2.565 21.93 2.833 ;
      RECT 21.85 2.565 21.855 2.798 ;
      RECT 21.845 2.565 21.85 2.788 ;
      RECT 21.84 2.565 21.845 2.768 ;
      RECT 22.105 1.785 22.275 2.255 ;
      RECT 22.05 1.778 22.245 2.239 ;
      RECT 22.05 1.792 22.28 2.238 ;
      RECT 22.035 1.793 22.28 2.219 ;
      RECT 22.03 1.811 22.28 2.205 ;
      RECT 22.035 1.794 22.285 2.203 ;
      RECT 22.02 1.825 22.285 2.188 ;
      RECT 22.035 1.8 22.29 2.173 ;
      RECT 22.015 1.84 22.29 2.17 ;
      RECT 22.03 1.812 22.295 2.155 ;
      RECT 22.03 1.824 22.3 2.135 ;
      RECT 22.015 1.84 22.305 2.118 ;
      RECT 22.015 1.85 22.31 1.973 ;
      RECT 22.01 1.85 22.31 1.93 ;
      RECT 22.01 1.865 22.315 1.908 ;
      RECT 22.105 1.775 22.245 2.255 ;
      RECT 22.105 1.773 22.215 2.255 ;
      RECT 22.191 1.77 22.215 2.255 ;
      RECT 21.85 3.437 21.855 3.483 ;
      RECT 21.84 3.285 21.85 3.507 ;
      RECT 21.835 3.13 21.84 3.532 ;
      RECT 21.82 3.092 21.835 3.543 ;
      RECT 21.815 3.075 21.82 3.55 ;
      RECT 21.805 3.063 21.815 3.557 ;
      RECT 21.8 3.054 21.805 3.559 ;
      RECT 21.795 3.052 21.8 3.563 ;
      RECT 21.75 3.043 21.795 3.578 ;
      RECT 21.745 3.035 21.75 3.592 ;
      RECT 21.74 3.032 21.745 3.596 ;
      RECT 21.725 3.027 21.74 3.604 ;
      RECT 21.67 3.017 21.725 3.615 ;
      RECT 21.635 3.005 21.67 3.616 ;
      RECT 21.626 3 21.635 3.61 ;
      RECT 21.54 3 21.626 3.6 ;
      RECT 21.51 3 21.54 3.578 ;
      RECT 21.5 3 21.505 3.558 ;
      RECT 21.495 3 21.5 3.52 ;
      RECT 21.49 3 21.495 3.478 ;
      RECT 21.485 3 21.49 3.438 ;
      RECT 21.48 3 21.485 3.368 ;
      RECT 21.47 3 21.48 3.29 ;
      RECT 21.465 3 21.47 3.19 ;
      RECT 21.505 3 21.51 3.56 ;
      RECT 21 3.082 21.09 3.56 ;
      RECT 20.985 3.085 21.105 3.558 ;
      RECT 21 3.084 21.105 3.558 ;
      RECT 20.965 3.091 21.13 3.548 ;
      RECT 20.985 3.085 21.13 3.548 ;
      RECT 20.95 3.097 21.13 3.536 ;
      RECT 20.985 3.088 21.18 3.529 ;
      RECT 20.936 3.105 21.18 3.527 ;
      RECT 20.965 3.095 21.19 3.515 ;
      RECT 20.936 3.116 21.22 3.506 ;
      RECT 20.85 3.14 21.22 3.5 ;
      RECT 20.85 3.153 21.26 3.483 ;
      RECT 20.845 3.175 21.26 3.476 ;
      RECT 20.815 3.19 21.26 3.466 ;
      RECT 20.81 3.201 21.26 3.456 ;
      RECT 20.78 3.214 21.26 3.447 ;
      RECT 20.765 3.232 21.26 3.436 ;
      RECT 20.74 3.245 21.26 3.426 ;
      RECT 21 3.081 21.01 3.56 ;
      RECT 21.046 2.505 21.085 2.75 ;
      RECT 20.96 2.505 21.095 2.748 ;
      RECT 20.845 2.53 21.095 2.745 ;
      RECT 20.845 2.53 21.1 2.743 ;
      RECT 20.845 2.53 21.115 2.738 ;
      RECT 20.951 2.505 21.13 2.718 ;
      RECT 20.865 2.513 21.13 2.718 ;
      RECT 20.535 1.865 20.705 2.3 ;
      RECT 20.525 1.899 20.705 2.283 ;
      RECT 20.605 1.835 20.775 2.27 ;
      RECT 20.51 1.91 20.775 2.248 ;
      RECT 20.605 1.845 20.78 2.238 ;
      RECT 20.535 1.897 20.81 2.223 ;
      RECT 20.495 1.923 20.81 2.208 ;
      RECT 20.495 1.965 20.82 2.188 ;
      RECT 20.49 1.99 20.825 2.17 ;
      RECT 20.49 2 20.83 2.155 ;
      RECT 20.485 1.937 20.81 2.153 ;
      RECT 20.485 2.01 20.835 2.138 ;
      RECT 20.48 1.947 20.81 2.135 ;
      RECT 20.475 2.031 20.84 2.118 ;
      RECT 20.475 2.063 20.845 2.098 ;
      RECT 20.47 1.977 20.82 2.09 ;
      RECT 20.475 1.962 20.81 2.118 ;
      RECT 20.49 1.932 20.81 2.17 ;
      RECT 20.335 2.519 20.56 2.775 ;
      RECT 20.335 2.552 20.58 2.765 ;
      RECT 20.3 2.552 20.58 2.763 ;
      RECT 20.3 2.565 20.585 2.753 ;
      RECT 20.3 2.585 20.595 2.745 ;
      RECT 20.3 2.682 20.6 2.738 ;
      RECT 20.28 2.43 20.41 2.728 ;
      RECT 20.235 2.585 20.595 2.67 ;
      RECT 20.225 2.43 20.41 2.615 ;
      RECT 20.225 2.462 20.496 2.615 ;
      RECT 20.19 2.992 20.21 3.17 ;
      RECT 20.155 2.945 20.19 3.17 ;
      RECT 20.14 2.885 20.155 3.17 ;
      RECT 20.115 2.832 20.14 3.17 ;
      RECT 20.1 2.785 20.115 3.17 ;
      RECT 20.08 2.762 20.1 3.17 ;
      RECT 20.055 2.727 20.08 3.17 ;
      RECT 20.045 2.573 20.055 3.17 ;
      RECT 20.015 2.568 20.045 3.161 ;
      RECT 20.01 2.565 20.015 3.151 ;
      RECT 19.995 2.565 20.01 3.125 ;
      RECT 19.99 2.565 19.995 3.088 ;
      RECT 19.965 2.565 19.99 3.04 ;
      RECT 19.945 2.565 19.965 2.965 ;
      RECT 19.935 2.565 19.945 2.925 ;
      RECT 19.93 2.565 19.935 2.9 ;
      RECT 19.925 2.565 19.93 2.883 ;
      RECT 19.92 2.565 19.925 2.865 ;
      RECT 19.915 2.566 19.92 2.855 ;
      RECT 19.905 2.568 19.915 2.823 ;
      RECT 19.895 2.57 19.905 2.79 ;
      RECT 19.885 2.573 19.895 2.763 ;
      RECT 20.21 3 20.435 3.17 ;
      RECT 19.54 1.812 19.71 2.265 ;
      RECT 19.54 1.812 19.8 2.231 ;
      RECT 19.54 1.812 19.83 2.215 ;
      RECT 19.54 1.812 19.86 2.188 ;
      RECT 19.796 1.79 19.875 2.17 ;
      RECT 19.575 1.797 19.88 2.155 ;
      RECT 19.575 1.805 19.89 2.118 ;
      RECT 19.535 1.832 19.89 2.09 ;
      RECT 19.52 1.845 19.89 2.055 ;
      RECT 19.54 1.82 19.91 2.045 ;
      RECT 19.515 1.885 19.91 2.015 ;
      RECT 19.515 1.915 19.915 1.998 ;
      RECT 19.51 1.945 19.915 1.985 ;
      RECT 19.575 1.794 19.875 2.17 ;
      RECT 19.71 1.791 19.796 2.249 ;
      RECT 19.661 1.792 19.875 2.17 ;
      RECT 19.805 3.452 19.85 3.645 ;
      RECT 19.795 3.422 19.805 3.645 ;
      RECT 19.79 3.407 19.795 3.645 ;
      RECT 19.75 3.317 19.79 3.645 ;
      RECT 19.745 3.23 19.75 3.645 ;
      RECT 19.735 3.2 19.745 3.645 ;
      RECT 19.73 3.16 19.735 3.645 ;
      RECT 19.72 3.122 19.73 3.645 ;
      RECT 19.715 3.087 19.72 3.645 ;
      RECT 19.695 3.04 19.715 3.645 ;
      RECT 19.68 2.965 19.695 3.645 ;
      RECT 19.675 2.92 19.68 3.64 ;
      RECT 19.67 2.9 19.675 3.613 ;
      RECT 19.665 2.88 19.67 3.598 ;
      RECT 19.66 2.855 19.665 3.578 ;
      RECT 19.655 2.833 19.66 3.563 ;
      RECT 19.65 2.811 19.655 3.545 ;
      RECT 19.645 2.79 19.65 3.535 ;
      RECT 19.635 2.762 19.645 3.505 ;
      RECT 19.625 2.725 19.635 3.473 ;
      RECT 19.615 2.685 19.625 3.44 ;
      RECT 19.605 2.663 19.615 3.41 ;
      RECT 19.575 2.615 19.605 3.342 ;
      RECT 19.56 2.575 19.575 3.269 ;
      RECT 19.55 2.575 19.56 3.235 ;
      RECT 19.545 2.575 19.55 3.21 ;
      RECT 19.54 2.575 19.545 3.195 ;
      RECT 19.535 2.575 19.54 3.173 ;
      RECT 19.53 2.575 19.535 3.16 ;
      RECT 19.515 2.575 19.53 3.125 ;
      RECT 19.495 2.575 19.515 3.065 ;
      RECT 19.485 2.575 19.495 3.015 ;
      RECT 19.465 2.575 19.485 2.963 ;
      RECT 19.445 2.575 19.465 2.92 ;
      RECT 19.435 2.575 19.445 2.908 ;
      RECT 19.405 2.575 19.435 2.895 ;
      RECT 19.375 2.596 19.405 2.875 ;
      RECT 19.365 2.624 19.375 2.855 ;
      RECT 19.35 2.641 19.365 2.823 ;
      RECT 19.345 2.655 19.35 2.79 ;
      RECT 19.34 2.663 19.345 2.763 ;
      RECT 19.335 2.671 19.34 2.725 ;
      RECT 19.34 3.195 19.345 3.53 ;
      RECT 19.305 3.182 19.34 3.529 ;
      RECT 19.235 3.122 19.305 3.528 ;
      RECT 19.155 3.065 19.235 3.527 ;
      RECT 19.02 3.025 19.155 3.526 ;
      RECT 19.02 3.212 19.355 3.515 ;
      RECT 18.98 3.212 19.355 3.505 ;
      RECT 18.98 3.23 19.36 3.5 ;
      RECT 18.98 3.32 19.365 3.49 ;
      RECT 18.975 3.015 19.14 3.47 ;
      RECT 18.97 3.015 19.14 3.213 ;
      RECT 18.97 3.172 19.335 3.213 ;
      RECT 18.97 3.16 19.33 3.213 ;
      RECT 18.105 5.02 18.275 6.49 ;
      RECT 18.105 6.315 18.28 6.485 ;
      RECT 17.735 1.74 17.905 2.93 ;
      RECT 17.735 1.74 18.205 1.91 ;
      RECT 17.735 6.97 18.205 7.14 ;
      RECT 17.735 5.95 17.905 7.14 ;
      RECT 16.745 1.74 16.915 2.93 ;
      RECT 16.745 1.74 17.215 1.91 ;
      RECT 16.745 6.97 17.215 7.14 ;
      RECT 16.745 5.95 16.915 7.14 ;
      RECT 14.895 2.635 15.065 3.865 ;
      RECT 14.95 0.855 15.12 2.805 ;
      RECT 14.895 0.575 15.065 1.025 ;
      RECT 14.895 7.855 15.065 8.305 ;
      RECT 14.95 6.075 15.12 8.025 ;
      RECT 14.895 5.015 15.065 6.245 ;
      RECT 14.375 0.575 14.545 3.865 ;
      RECT 14.375 2.075 14.78 2.405 ;
      RECT 14.375 1.235 14.78 1.565 ;
      RECT 14.375 5.015 14.545 8.305 ;
      RECT 14.375 7.315 14.78 7.645 ;
      RECT 14.375 6.475 14.78 6.805 ;
      RECT 11.71 1.975 12.44 2.215 ;
      RECT 12.252 1.77 12.44 2.215 ;
      RECT 12.08 1.782 12.455 2.209 ;
      RECT 11.995 1.797 12.475 2.194 ;
      RECT 11.995 1.812 12.48 2.184 ;
      RECT 11.95 1.832 12.495 2.176 ;
      RECT 11.927 1.867 12.51 2.13 ;
      RECT 11.841 1.89 12.515 2.09 ;
      RECT 11.841 1.908 12.525 2.06 ;
      RECT 11.71 1.977 12.53 2.023 ;
      RECT 11.755 1.92 12.525 2.06 ;
      RECT 11.841 1.872 12.51 2.13 ;
      RECT 11.927 1.841 12.495 2.176 ;
      RECT 11.95 1.822 12.48 2.184 ;
      RECT 11.995 1.795 12.455 2.209 ;
      RECT 12.08 1.777 12.44 2.215 ;
      RECT 12.166 1.771 12.44 2.215 ;
      RECT 12.252 1.766 12.385 2.215 ;
      RECT 12.338 1.761 12.385 2.215 ;
      RECT 12.03 2.659 12.2 3.045 ;
      RECT 12.025 2.659 12.2 3.04 ;
      RECT 12 2.659 12.2 3.005 ;
      RECT 12 2.687 12.21 2.995 ;
      RECT 11.98 2.687 12.21 2.955 ;
      RECT 11.975 2.687 12.21 2.928 ;
      RECT 11.975 2.705 12.215 2.92 ;
      RECT 11.92 2.705 12.215 2.855 ;
      RECT 11.92 2.722 12.225 2.838 ;
      RECT 11.91 2.722 12.225 2.778 ;
      RECT 11.91 2.739 12.23 2.775 ;
      RECT 11.905 2.575 12.075 2.753 ;
      RECT 11.905 2.609 12.161 2.753 ;
      RECT 11.9 3.375 11.905 3.388 ;
      RECT 11.895 3.27 11.9 3.393 ;
      RECT 11.87 3.13 11.895 3.408 ;
      RECT 11.835 3.081 11.87 3.44 ;
      RECT 11.83 3.049 11.835 3.46 ;
      RECT 11.825 3.04 11.83 3.46 ;
      RECT 11.745 3.005 11.825 3.46 ;
      RECT 11.682 2.975 11.745 3.46 ;
      RECT 11.596 2.963 11.682 3.46 ;
      RECT 11.51 2.949 11.596 3.46 ;
      RECT 11.43 2.936 11.51 3.446 ;
      RECT 11.395 2.928 11.43 3.426 ;
      RECT 11.385 2.925 11.395 3.417 ;
      RECT 11.355 2.92 11.385 3.404 ;
      RECT 11.305 2.895 11.355 3.38 ;
      RECT 11.291 2.869 11.305 3.362 ;
      RECT 11.205 2.829 11.291 3.338 ;
      RECT 11.16 2.777 11.205 3.307 ;
      RECT 11.15 2.752 11.16 3.294 ;
      RECT 11.145 2.533 11.15 2.555 ;
      RECT 11.14 2.735 11.15 3.29 ;
      RECT 11.14 2.531 11.145 2.645 ;
      RECT 11.13 2.527 11.14 3.286 ;
      RECT 11.086 2.525 11.13 3.274 ;
      RECT 11 2.525 11.086 3.245 ;
      RECT 10.97 2.525 11 3.218 ;
      RECT 10.955 2.525 10.97 3.206 ;
      RECT 10.915 2.537 10.955 3.191 ;
      RECT 10.895 2.556 10.915 3.17 ;
      RECT 10.885 2.566 10.895 3.154 ;
      RECT 10.875 2.572 10.885 3.143 ;
      RECT 10.855 2.582 10.875 3.126 ;
      RECT 10.85 2.591 10.855 3.113 ;
      RECT 10.845 2.595 10.85 3.063 ;
      RECT 10.835 2.601 10.845 2.98 ;
      RECT 10.83 2.605 10.835 2.894 ;
      RECT 10.825 2.625 10.83 2.831 ;
      RECT 10.82 2.648 10.825 2.778 ;
      RECT 10.815 2.666 10.82 2.723 ;
      RECT 11.425 2.485 11.595 2.745 ;
      RECT 11.595 2.45 11.64 2.731 ;
      RECT 11.556 2.452 11.645 2.714 ;
      RECT 11.445 2.469 11.731 2.685 ;
      RECT 11.445 2.484 11.735 2.657 ;
      RECT 11.445 2.465 11.645 2.714 ;
      RECT 11.47 2.453 11.595 2.745 ;
      RECT 11.556 2.451 11.64 2.731 ;
      RECT 10.61 1.84 10.78 2.33 ;
      RECT 10.61 1.84 10.815 2.31 ;
      RECT 10.745 1.76 10.855 2.27 ;
      RECT 10.726 1.764 10.875 2.24 ;
      RECT 10.64 1.772 10.895 2.223 ;
      RECT 10.64 1.778 10.9 2.213 ;
      RECT 10.64 1.787 10.92 2.201 ;
      RECT 10.615 1.812 10.95 2.179 ;
      RECT 10.615 1.832 10.955 2.159 ;
      RECT 10.61 1.845 10.965 2.139 ;
      RECT 10.61 1.912 10.97 2.12 ;
      RECT 10.61 2.045 10.975 2.107 ;
      RECT 10.605 1.85 10.965 1.94 ;
      RECT 10.615 1.807 10.92 2.201 ;
      RECT 10.726 1.762 10.855 2.27 ;
      RECT 10.6 3.515 10.9 3.77 ;
      RECT 10.685 3.481 10.9 3.77 ;
      RECT 10.685 3.484 10.905 3.63 ;
      RECT 10.62 3.505 10.905 3.63 ;
      RECT 10.655 3.495 10.9 3.77 ;
      RECT 10.65 3.5 10.905 3.63 ;
      RECT 10.685 3.479 10.886 3.77 ;
      RECT 10.771 3.47 10.886 3.77 ;
      RECT 10.771 3.464 10.8 3.77 ;
      RECT 10.26 3.105 10.27 3.595 ;
      RECT 9.92 3.04 9.93 3.34 ;
      RECT 10.435 3.212 10.44 3.431 ;
      RECT 10.425 3.192 10.435 3.448 ;
      RECT 10.415 3.172 10.425 3.478 ;
      RECT 10.41 3.162 10.415 3.493 ;
      RECT 10.405 3.158 10.41 3.498 ;
      RECT 10.39 3.15 10.405 3.505 ;
      RECT 10.35 3.13 10.39 3.53 ;
      RECT 10.325 3.112 10.35 3.563 ;
      RECT 10.32 3.11 10.325 3.576 ;
      RECT 10.3 3.107 10.32 3.58 ;
      RECT 10.27 3.105 10.3 3.59 ;
      RECT 10.2 3.107 10.26 3.591 ;
      RECT 10.18 3.107 10.2 3.585 ;
      RECT 10.155 3.105 10.18 3.582 ;
      RECT 10.12 3.1 10.155 3.578 ;
      RECT 10.1 3.094 10.12 3.565 ;
      RECT 10.09 3.091 10.1 3.553 ;
      RECT 10.07 3.088 10.09 3.538 ;
      RECT 10.05 3.084 10.07 3.52 ;
      RECT 10.045 3.081 10.05 3.51 ;
      RECT 10.04 3.08 10.045 3.508 ;
      RECT 10.03 3.077 10.04 3.5 ;
      RECT 10.02 3.071 10.03 3.483 ;
      RECT 10.01 3.065 10.02 3.465 ;
      RECT 10 3.059 10.01 3.453 ;
      RECT 9.99 3.053 10 3.433 ;
      RECT 9.985 3.049 9.99 3.418 ;
      RECT 9.98 3.047 9.985 3.41 ;
      RECT 9.975 3.045 9.98 3.403 ;
      RECT 9.97 3.043 9.975 3.393 ;
      RECT 9.965 3.041 9.97 3.387 ;
      RECT 9.955 3.04 9.965 3.377 ;
      RECT 9.945 3.04 9.955 3.368 ;
      RECT 9.93 3.04 9.945 3.353 ;
      RECT 9.89 3.04 9.92 3.337 ;
      RECT 9.87 3.042 9.89 3.332 ;
      RECT 9.865 3.047 9.87 3.33 ;
      RECT 9.835 3.055 9.865 3.328 ;
      RECT 9.805 3.07 9.835 3.327 ;
      RECT 9.76 3.092 9.805 3.332 ;
      RECT 9.755 3.107 9.76 3.336 ;
      RECT 9.74 3.112 9.755 3.338 ;
      RECT 9.735 3.116 9.74 3.34 ;
      RECT 9.675 3.139 9.735 3.349 ;
      RECT 9.655 3.165 9.675 3.362 ;
      RECT 9.645 3.172 9.655 3.366 ;
      RECT 9.63 3.179 9.645 3.369 ;
      RECT 9.61 3.189 9.63 3.372 ;
      RECT 9.605 3.197 9.61 3.375 ;
      RECT 9.56 3.202 9.605 3.382 ;
      RECT 9.55 3.205 9.56 3.389 ;
      RECT 9.54 3.205 9.55 3.393 ;
      RECT 9.505 3.207 9.54 3.405 ;
      RECT 9.485 3.21 9.505 3.418 ;
      RECT 9.445 3.213 9.485 3.429 ;
      RECT 9.43 3.215 9.445 3.442 ;
      RECT 9.42 3.215 9.43 3.447 ;
      RECT 9.395 3.216 9.42 3.455 ;
      RECT 9.385 3.218 9.395 3.46 ;
      RECT 9.38 3.219 9.385 3.463 ;
      RECT 9.355 3.217 9.38 3.466 ;
      RECT 9.34 3.215 9.355 3.467 ;
      RECT 9.32 3.212 9.34 3.469 ;
      RECT 9.3 3.207 9.32 3.469 ;
      RECT 9.24 3.202 9.3 3.466 ;
      RECT 9.205 3.177 9.24 3.462 ;
      RECT 9.195 3.154 9.205 3.46 ;
      RECT 9.165 3.131 9.195 3.46 ;
      RECT 9.155 3.11 9.165 3.46 ;
      RECT 9.13 3.092 9.155 3.458 ;
      RECT 9.115 3.07 9.13 3.455 ;
      RECT 9.1 3.052 9.115 3.453 ;
      RECT 9.08 3.042 9.1 3.451 ;
      RECT 9.065 3.037 9.08 3.45 ;
      RECT 9.05 3.035 9.065 3.449 ;
      RECT 9.02 3.036 9.05 3.447 ;
      RECT 9 3.039 9.02 3.445 ;
      RECT 8.943 3.043 9 3.445 ;
      RECT 8.857 3.052 8.943 3.445 ;
      RECT 8.771 3.063 8.857 3.445 ;
      RECT 8.685 3.074 8.771 3.445 ;
      RECT 8.665 3.081 8.685 3.453 ;
      RECT 8.655 3.084 8.665 3.46 ;
      RECT 8.59 3.089 8.655 3.478 ;
      RECT 8.56 3.096 8.59 3.503 ;
      RECT 8.55 3.099 8.56 3.51 ;
      RECT 8.505 3.103 8.55 3.515 ;
      RECT 8.475 3.108 8.505 3.52 ;
      RECT 8.474 3.11 8.475 3.52 ;
      RECT 8.388 3.116 8.474 3.52 ;
      RECT 8.302 3.127 8.388 3.52 ;
      RECT 8.216 3.139 8.302 3.52 ;
      RECT 8.13 3.15 8.216 3.52 ;
      RECT 8.115 3.157 8.13 3.515 ;
      RECT 8.11 3.159 8.115 3.509 ;
      RECT 8.09 3.17 8.11 3.504 ;
      RECT 8.08 3.188 8.09 3.498 ;
      RECT 8.075 3.2 8.08 3.298 ;
      RECT 10.37 1.953 10.39 2.04 ;
      RECT 10.365 1.888 10.37 2.072 ;
      RECT 10.355 1.855 10.365 2.077 ;
      RECT 10.35 1.835 10.355 2.083 ;
      RECT 10.32 1.835 10.35 2.1 ;
      RECT 10.271 1.835 10.32 2.136 ;
      RECT 10.185 1.835 10.271 2.194 ;
      RECT 10.156 1.845 10.185 2.243 ;
      RECT 10.07 1.887 10.156 2.296 ;
      RECT 10.05 1.925 10.07 2.343 ;
      RECT 10.025 1.942 10.05 2.363 ;
      RECT 10.015 1.956 10.025 2.383 ;
      RECT 10.01 1.962 10.015 2.393 ;
      RECT 10.005 1.966 10.01 2.4 ;
      RECT 9.955 1.986 10.005 2.405 ;
      RECT 9.89 2.03 9.955 2.405 ;
      RECT 9.865 2.08 9.89 2.405 ;
      RECT 9.855 2.11 9.865 2.405 ;
      RECT 9.85 2.137 9.855 2.405 ;
      RECT 9.845 2.155 9.85 2.405 ;
      RECT 9.835 2.197 9.845 2.405 ;
      RECT 10.185 2.755 10.355 2.93 ;
      RECT 10.125 2.583 10.185 2.918 ;
      RECT 10.115 2.576 10.125 2.901 ;
      RECT 10.07 2.755 10.355 2.881 ;
      RECT 10.051 2.755 10.355 2.859 ;
      RECT 9.965 2.755 10.355 2.824 ;
      RECT 9.945 2.575 10.115 2.78 ;
      RECT 9.945 2.722 10.35 2.78 ;
      RECT 9.945 2.67 10.325 2.78 ;
      RECT 9.945 2.625 10.29 2.78 ;
      RECT 9.945 2.607 10.255 2.78 ;
      RECT 9.945 2.597 10.25 2.78 ;
      RECT 10.115 7.855 10.285 8.305 ;
      RECT 10.17 6.075 10.34 8.025 ;
      RECT 10.115 5.015 10.285 6.245 ;
      RECT 9.595 5.015 9.765 8.305 ;
      RECT 9.595 7.315 10 7.645 ;
      RECT 9.595 6.475 10 6.805 ;
      RECT 9.665 3.555 9.855 3.78 ;
      RECT 9.655 3.556 9.86 3.775 ;
      RECT 9.655 3.558 9.87 3.755 ;
      RECT 9.655 3.562 9.875 3.74 ;
      RECT 9.655 3.549 9.825 3.775 ;
      RECT 9.655 3.552 9.85 3.775 ;
      RECT 9.665 3.548 9.825 3.78 ;
      RECT 9.751 3.546 9.825 3.78 ;
      RECT 9.375 2.797 9.545 3.035 ;
      RECT 9.375 2.797 9.631 2.949 ;
      RECT 9.375 2.797 9.635 2.859 ;
      RECT 9.425 2.57 9.645 2.838 ;
      RECT 9.42 2.587 9.65 2.811 ;
      RECT 9.385 2.745 9.65 2.811 ;
      RECT 9.405 2.595 9.545 3.035 ;
      RECT 9.395 2.677 9.655 2.794 ;
      RECT 9.39 2.725 9.655 2.794 ;
      RECT 9.395 2.635 9.65 2.811 ;
      RECT 9.42 2.572 9.645 2.838 ;
      RECT 8.985 2.547 9.155 2.745 ;
      RECT 8.985 2.547 9.2 2.72 ;
      RECT 9.055 2.49 9.225 2.678 ;
      RECT 9.03 2.505 9.225 2.678 ;
      RECT 8.645 2.551 8.675 2.745 ;
      RECT 8.64 2.523 8.645 2.745 ;
      RECT 8.61 2.497 8.64 2.747 ;
      RECT 8.585 2.455 8.61 2.75 ;
      RECT 8.575 2.427 8.585 2.752 ;
      RECT 8.54 2.407 8.575 2.754 ;
      RECT 8.475 2.392 8.54 2.76 ;
      RECT 8.425 2.39 8.475 2.766 ;
      RECT 8.402 2.392 8.425 2.771 ;
      RECT 8.316 2.403 8.402 2.777 ;
      RECT 8.23 2.421 8.316 2.787 ;
      RECT 8.215 2.432 8.23 2.793 ;
      RECT 8.145 2.455 8.215 2.799 ;
      RECT 8.09 2.487 8.145 2.807 ;
      RECT 8.05 2.51 8.09 2.813 ;
      RECT 8.036 2.523 8.05 2.816 ;
      RECT 7.95 2.545 8.036 2.822 ;
      RECT 7.935 2.57 7.95 2.828 ;
      RECT 7.895 2.585 7.935 2.832 ;
      RECT 7.845 2.6 7.895 2.837 ;
      RECT 7.82 2.607 7.845 2.841 ;
      RECT 7.76 2.602 7.82 2.845 ;
      RECT 7.745 2.593 7.76 2.849 ;
      RECT 7.675 2.583 7.745 2.845 ;
      RECT 7.65 2.575 7.67 2.835 ;
      RECT 7.591 2.575 7.65 2.813 ;
      RECT 7.505 2.575 7.591 2.77 ;
      RECT 7.67 2.575 7.675 2.84 ;
      RECT 8.365 1.806 8.535 2.14 ;
      RECT 8.335 1.806 8.535 2.135 ;
      RECT 8.275 1.773 8.335 2.123 ;
      RECT 8.275 1.829 8.545 2.118 ;
      RECT 8.25 1.829 8.545 2.112 ;
      RECT 8.245 1.77 8.275 2.109 ;
      RECT 8.23 1.776 8.365 2.107 ;
      RECT 8.225 1.784 8.45 2.095 ;
      RECT 8.225 1.836 8.56 2.048 ;
      RECT 8.21 1.792 8.45 2.043 ;
      RECT 8.21 1.862 8.57 1.984 ;
      RECT 8.18 1.812 8.535 1.945 ;
      RECT 8.18 1.902 8.58 1.941 ;
      RECT 8.23 1.781 8.45 2.107 ;
      RECT 7.57 2.111 7.625 2.375 ;
      RECT 7.57 2.111 7.69 2.374 ;
      RECT 7.57 2.111 7.715 2.373 ;
      RECT 7.57 2.111 7.78 2.372 ;
      RECT 7.715 2.077 7.795 2.371 ;
      RECT 7.53 2.121 7.94 2.37 ;
      RECT 7.57 2.118 7.94 2.37 ;
      RECT 7.53 2.126 7.945 2.363 ;
      RECT 7.515 2.128 7.945 2.362 ;
      RECT 7.515 2.135 7.95 2.358 ;
      RECT 7.495 2.134 7.945 2.354 ;
      RECT 7.495 2.142 7.955 2.353 ;
      RECT 7.49 2.139 7.95 2.349 ;
      RECT 7.49 2.152 7.965 2.348 ;
      RECT 7.475 2.142 7.955 2.347 ;
      RECT 7.44 2.155 7.965 2.34 ;
      RECT 7.625 2.11 7.935 2.37 ;
      RECT 7.625 2.095 7.885 2.37 ;
      RECT 7.69 2.082 7.82 2.37 ;
      RECT 7.235 3.171 7.25 3.564 ;
      RECT 7.2 3.176 7.25 3.563 ;
      RECT 7.235 3.175 7.295 3.562 ;
      RECT 7.18 3.186 7.295 3.561 ;
      RECT 7.195 3.182 7.295 3.561 ;
      RECT 7.16 3.192 7.37 3.558 ;
      RECT 7.16 3.211 7.415 3.556 ;
      RECT 7.16 3.218 7.42 3.553 ;
      RECT 7.145 3.195 7.37 3.55 ;
      RECT 7.125 3.2 7.37 3.543 ;
      RECT 7.12 3.204 7.37 3.539 ;
      RECT 7.12 3.221 7.43 3.538 ;
      RECT 7.1 3.215 7.415 3.534 ;
      RECT 7.1 3.224 7.435 3.528 ;
      RECT 7.095 3.23 7.435 3.3 ;
      RECT 7.16 3.19 7.295 3.558 ;
      RECT 7.035 2.553 7.235 2.865 ;
      RECT 7.11 2.531 7.235 2.865 ;
      RECT 7.05 2.55 7.24 2.85 ;
      RECT 7.02 2.561 7.24 2.848 ;
      RECT 7.035 2.556 7.245 2.814 ;
      RECT 7.02 2.66 7.25 2.781 ;
      RECT 7.05 2.532 7.235 2.865 ;
      RECT 7.11 2.51 7.21 2.865 ;
      RECT 7.135 2.507 7.21 2.865 ;
      RECT 7.135 2.502 7.155 2.865 ;
      RECT 6.54 2.57 6.715 2.745 ;
      RECT 6.535 2.57 6.715 2.743 ;
      RECT 6.51 2.57 6.715 2.738 ;
      RECT 6.455 2.55 6.625 2.728 ;
      RECT 6.455 2.557 6.69 2.728 ;
      RECT 6.54 3.237 6.555 3.42 ;
      RECT 6.53 3.215 6.54 3.42 ;
      RECT 6.515 3.195 6.53 3.42 ;
      RECT 6.505 3.17 6.515 3.42 ;
      RECT 6.475 3.135 6.505 3.42 ;
      RECT 6.44 3.075 6.475 3.42 ;
      RECT 6.435 3.037 6.44 3.42 ;
      RECT 6.385 2.988 6.435 3.42 ;
      RECT 6.375 2.938 6.385 3.408 ;
      RECT 6.36 2.917 6.375 3.368 ;
      RECT 6.34 2.885 6.36 3.318 ;
      RECT 6.315 2.841 6.34 3.258 ;
      RECT 6.31 2.813 6.315 3.213 ;
      RECT 6.305 2.804 6.31 3.199 ;
      RECT 6.3 2.797 6.305 3.186 ;
      RECT 6.295 2.792 6.3 3.175 ;
      RECT 6.29 2.777 6.295 3.165 ;
      RECT 6.285 2.755 6.29 3.152 ;
      RECT 6.275 2.715 6.285 3.127 ;
      RECT 6.25 2.645 6.275 3.083 ;
      RECT 6.245 2.585 6.25 3.048 ;
      RECT 6.23 2.565 6.245 3.015 ;
      RECT 6.225 2.565 6.23 2.99 ;
      RECT 6.195 2.565 6.225 2.945 ;
      RECT 6.15 2.565 6.195 2.885 ;
      RECT 6.075 2.565 6.15 2.833 ;
      RECT 6.07 2.565 6.075 2.798 ;
      RECT 6.065 2.565 6.07 2.788 ;
      RECT 6.06 2.565 6.065 2.768 ;
      RECT 6.325 1.785 6.495 2.255 ;
      RECT 6.27 1.778 6.465 2.239 ;
      RECT 6.27 1.792 6.5 2.238 ;
      RECT 6.255 1.793 6.5 2.219 ;
      RECT 6.25 1.811 6.5 2.205 ;
      RECT 6.255 1.794 6.505 2.203 ;
      RECT 6.24 1.825 6.505 2.188 ;
      RECT 6.255 1.8 6.51 2.173 ;
      RECT 6.235 1.84 6.51 2.17 ;
      RECT 6.25 1.812 6.515 2.155 ;
      RECT 6.25 1.824 6.52 2.135 ;
      RECT 6.235 1.84 6.525 2.118 ;
      RECT 6.235 1.85 6.53 1.973 ;
      RECT 6.23 1.85 6.53 1.93 ;
      RECT 6.23 1.865 6.535 1.908 ;
      RECT 6.325 1.775 6.465 2.255 ;
      RECT 6.325 1.773 6.435 2.255 ;
      RECT 6.411 1.77 6.435 2.255 ;
      RECT 6.07 3.437 6.075 3.483 ;
      RECT 6.06 3.285 6.07 3.507 ;
      RECT 6.055 3.13 6.06 3.532 ;
      RECT 6.04 3.092 6.055 3.543 ;
      RECT 6.035 3.075 6.04 3.55 ;
      RECT 6.025 3.063 6.035 3.557 ;
      RECT 6.02 3.054 6.025 3.559 ;
      RECT 6.015 3.052 6.02 3.563 ;
      RECT 5.97 3.043 6.015 3.578 ;
      RECT 5.965 3.035 5.97 3.592 ;
      RECT 5.96 3.032 5.965 3.596 ;
      RECT 5.945 3.027 5.96 3.604 ;
      RECT 5.89 3.017 5.945 3.615 ;
      RECT 5.855 3.005 5.89 3.616 ;
      RECT 5.846 3 5.855 3.61 ;
      RECT 5.76 3 5.846 3.6 ;
      RECT 5.73 3 5.76 3.578 ;
      RECT 5.72 3 5.725 3.558 ;
      RECT 5.715 3 5.72 3.52 ;
      RECT 5.71 3 5.715 3.478 ;
      RECT 5.705 3 5.71 3.438 ;
      RECT 5.7 3 5.705 3.368 ;
      RECT 5.69 3 5.7 3.29 ;
      RECT 5.685 3 5.69 3.19 ;
      RECT 5.725 3 5.73 3.56 ;
      RECT 5.22 3.082 5.31 3.56 ;
      RECT 5.205 3.085 5.325 3.558 ;
      RECT 5.22 3.084 5.325 3.558 ;
      RECT 5.185 3.091 5.35 3.548 ;
      RECT 5.205 3.085 5.35 3.548 ;
      RECT 5.17 3.097 5.35 3.536 ;
      RECT 5.205 3.088 5.4 3.529 ;
      RECT 5.156 3.105 5.4 3.527 ;
      RECT 5.185 3.095 5.41 3.515 ;
      RECT 5.156 3.116 5.44 3.506 ;
      RECT 5.07 3.14 5.44 3.5 ;
      RECT 5.07 3.153 5.48 3.483 ;
      RECT 5.065 3.175 5.48 3.476 ;
      RECT 5.035 3.19 5.48 3.466 ;
      RECT 5.03 3.201 5.48 3.456 ;
      RECT 5 3.214 5.48 3.447 ;
      RECT 4.985 3.232 5.48 3.436 ;
      RECT 4.96 3.245 5.48 3.426 ;
      RECT 5.22 3.081 5.23 3.56 ;
      RECT 5.266 2.505 5.305 2.75 ;
      RECT 5.18 2.505 5.315 2.748 ;
      RECT 5.065 2.53 5.315 2.745 ;
      RECT 5.065 2.53 5.32 2.743 ;
      RECT 5.065 2.53 5.335 2.738 ;
      RECT 5.171 2.505 5.35 2.718 ;
      RECT 5.085 2.513 5.35 2.718 ;
      RECT 4.755 1.865 4.925 2.3 ;
      RECT 4.745 1.899 4.925 2.283 ;
      RECT 4.825 1.835 4.995 2.27 ;
      RECT 4.73 1.91 4.995 2.248 ;
      RECT 4.825 1.845 5 2.238 ;
      RECT 4.755 1.897 5.03 2.223 ;
      RECT 4.715 1.923 5.03 2.208 ;
      RECT 4.715 1.965 5.04 2.188 ;
      RECT 4.71 1.99 5.045 2.17 ;
      RECT 4.71 2 5.05 2.155 ;
      RECT 4.705 1.937 5.03 2.153 ;
      RECT 4.705 2.01 5.055 2.138 ;
      RECT 4.7 1.947 5.03 2.135 ;
      RECT 4.695 2.031 5.06 2.118 ;
      RECT 4.695 2.063 5.065 2.098 ;
      RECT 4.69 1.977 5.04 2.09 ;
      RECT 4.695 1.962 5.03 2.118 ;
      RECT 4.71 1.932 5.03 2.17 ;
      RECT 4.555 2.519 4.78 2.775 ;
      RECT 4.555 2.552 4.8 2.765 ;
      RECT 4.52 2.552 4.8 2.763 ;
      RECT 4.52 2.565 4.805 2.753 ;
      RECT 4.52 2.585 4.815 2.745 ;
      RECT 4.52 2.682 4.82 2.738 ;
      RECT 4.5 2.43 4.63 2.728 ;
      RECT 4.455 2.585 4.815 2.67 ;
      RECT 4.445 2.43 4.63 2.615 ;
      RECT 4.445 2.462 4.716 2.615 ;
      RECT 4.41 2.992 4.43 3.17 ;
      RECT 4.375 2.945 4.41 3.17 ;
      RECT 4.36 2.885 4.375 3.17 ;
      RECT 4.335 2.832 4.36 3.17 ;
      RECT 4.32 2.785 4.335 3.17 ;
      RECT 4.3 2.762 4.32 3.17 ;
      RECT 4.275 2.727 4.3 3.17 ;
      RECT 4.265 2.573 4.275 3.17 ;
      RECT 4.235 2.568 4.265 3.161 ;
      RECT 4.23 2.565 4.235 3.151 ;
      RECT 4.215 2.565 4.23 3.125 ;
      RECT 4.21 2.565 4.215 3.088 ;
      RECT 4.185 2.565 4.21 3.04 ;
      RECT 4.165 2.565 4.185 2.965 ;
      RECT 4.155 2.565 4.165 2.925 ;
      RECT 4.15 2.565 4.155 2.9 ;
      RECT 4.145 2.565 4.15 2.883 ;
      RECT 4.14 2.565 4.145 2.865 ;
      RECT 4.135 2.566 4.14 2.855 ;
      RECT 4.125 2.568 4.135 2.823 ;
      RECT 4.115 2.57 4.125 2.79 ;
      RECT 4.105 2.573 4.115 2.763 ;
      RECT 4.43 3 4.655 3.17 ;
      RECT 3.76 1.812 3.93 2.265 ;
      RECT 3.76 1.812 4.02 2.231 ;
      RECT 3.76 1.812 4.05 2.215 ;
      RECT 3.76 1.812 4.08 2.188 ;
      RECT 4.016 1.79 4.095 2.17 ;
      RECT 3.795 1.797 4.1 2.155 ;
      RECT 3.795 1.805 4.11 2.118 ;
      RECT 3.755 1.832 4.11 2.09 ;
      RECT 3.74 1.845 4.11 2.055 ;
      RECT 3.76 1.82 4.13 2.045 ;
      RECT 3.735 1.885 4.13 2.015 ;
      RECT 3.735 1.915 4.135 1.998 ;
      RECT 3.73 1.945 4.135 1.985 ;
      RECT 3.795 1.794 4.095 2.17 ;
      RECT 3.93 1.791 4.016 2.249 ;
      RECT 3.881 1.792 4.095 2.17 ;
      RECT 4.025 3.452 4.07 3.645 ;
      RECT 4.015 3.422 4.025 3.645 ;
      RECT 4.01 3.407 4.015 3.645 ;
      RECT 3.97 3.317 4.01 3.645 ;
      RECT 3.965 3.23 3.97 3.645 ;
      RECT 3.955 3.2 3.965 3.645 ;
      RECT 3.95 3.16 3.955 3.645 ;
      RECT 3.94 3.122 3.95 3.645 ;
      RECT 3.935 3.087 3.94 3.645 ;
      RECT 3.915 3.04 3.935 3.645 ;
      RECT 3.9 2.965 3.915 3.645 ;
      RECT 3.895 2.92 3.9 3.64 ;
      RECT 3.89 2.9 3.895 3.613 ;
      RECT 3.885 2.88 3.89 3.598 ;
      RECT 3.88 2.855 3.885 3.578 ;
      RECT 3.875 2.833 3.88 3.563 ;
      RECT 3.87 2.811 3.875 3.545 ;
      RECT 3.865 2.79 3.87 3.535 ;
      RECT 3.855 2.762 3.865 3.505 ;
      RECT 3.845 2.725 3.855 3.473 ;
      RECT 3.835 2.685 3.845 3.44 ;
      RECT 3.825 2.663 3.835 3.41 ;
      RECT 3.795 2.615 3.825 3.342 ;
      RECT 3.78 2.575 3.795 3.269 ;
      RECT 3.77 2.575 3.78 3.235 ;
      RECT 3.765 2.575 3.77 3.21 ;
      RECT 3.76 2.575 3.765 3.195 ;
      RECT 3.755 2.575 3.76 3.173 ;
      RECT 3.75 2.575 3.755 3.16 ;
      RECT 3.735 2.575 3.75 3.125 ;
      RECT 3.715 2.575 3.735 3.065 ;
      RECT 3.705 2.575 3.715 3.015 ;
      RECT 3.685 2.575 3.705 2.963 ;
      RECT 3.665 2.575 3.685 2.92 ;
      RECT 3.655 2.575 3.665 2.908 ;
      RECT 3.625 2.575 3.655 2.895 ;
      RECT 3.595 2.596 3.625 2.875 ;
      RECT 3.585 2.624 3.595 2.855 ;
      RECT 3.57 2.641 3.585 2.823 ;
      RECT 3.565 2.655 3.57 2.79 ;
      RECT 3.56 2.663 3.565 2.763 ;
      RECT 3.555 2.671 3.56 2.725 ;
      RECT 3.56 3.195 3.565 3.53 ;
      RECT 3.525 3.182 3.56 3.529 ;
      RECT 3.455 3.122 3.525 3.528 ;
      RECT 3.375 3.065 3.455 3.527 ;
      RECT 3.24 3.025 3.375 3.526 ;
      RECT 3.24 3.212 3.575 3.515 ;
      RECT 3.2 3.212 3.575 3.505 ;
      RECT 3.2 3.23 3.58 3.5 ;
      RECT 3.2 3.32 3.585 3.49 ;
      RECT 3.195 3.015 3.36 3.47 ;
      RECT 3.19 3.015 3.36 3.213 ;
      RECT 3.19 3.172 3.555 3.213 ;
      RECT 3.19 3.16 3.55 3.213 ;
      RECT 1.18 7.855 1.35 8.305 ;
      RECT 1.235 6.075 1.405 8.025 ;
      RECT 1.18 5.015 1.35 6.245 ;
      RECT 0.66 5.015 0.83 8.305 ;
      RECT 0.66 7.315 1.065 7.645 ;
      RECT 0.66 6.475 1.065 6.805 ;
      RECT 81.23 7.8 81.4 8.31 ;
      RECT 80.24 0.57 80.41 1.08 ;
      RECT 80.24 2.39 80.41 3.86 ;
      RECT 80.24 5.02 80.41 6.49 ;
      RECT 80.24 7.8 80.41 8.31 ;
      RECT 78.88 0.575 79.05 3.865 ;
      RECT 78.88 5.015 79.05 8.305 ;
      RECT 78.45 0.575 78.62 1.085 ;
      RECT 78.45 1.655 78.62 3.865 ;
      RECT 78.45 5.015 78.62 7.225 ;
      RECT 78.45 7.795 78.62 8.305 ;
      RECT 76.06 2.85 76.43 3.22 ;
      RECT 74.1 5.015 74.27 8.305 ;
      RECT 73.67 5.015 73.84 7.225 ;
      RECT 73.67 7.795 73.84 8.305 ;
      RECT 65.445 7.8 65.615 8.31 ;
      RECT 64.455 0.57 64.625 1.08 ;
      RECT 64.455 2.39 64.625 3.86 ;
      RECT 64.455 5.02 64.625 6.49 ;
      RECT 64.455 7.8 64.625 8.31 ;
      RECT 63.095 0.575 63.265 3.865 ;
      RECT 63.095 5.015 63.265 8.305 ;
      RECT 62.665 0.575 62.835 1.085 ;
      RECT 62.665 1.655 62.835 3.865 ;
      RECT 62.665 5.015 62.835 7.225 ;
      RECT 62.665 7.795 62.835 8.305 ;
      RECT 60.275 2.85 60.645 3.22 ;
      RECT 58.315 5.015 58.485 8.305 ;
      RECT 57.885 5.015 58.055 7.225 ;
      RECT 57.885 7.795 58.055 8.305 ;
      RECT 49.66 7.8 49.83 8.31 ;
      RECT 48.67 0.57 48.84 1.08 ;
      RECT 48.67 2.39 48.84 3.86 ;
      RECT 48.67 5.02 48.84 6.49 ;
      RECT 48.67 7.8 48.84 8.31 ;
      RECT 47.31 0.575 47.48 3.865 ;
      RECT 47.31 5.015 47.48 8.305 ;
      RECT 46.88 0.575 47.05 1.085 ;
      RECT 46.88 1.655 47.05 3.865 ;
      RECT 46.88 5.015 47.05 7.225 ;
      RECT 46.88 7.795 47.05 8.305 ;
      RECT 44.49 2.85 44.86 3.22 ;
      RECT 42.53 5.015 42.7 8.305 ;
      RECT 42.1 5.015 42.27 7.225 ;
      RECT 42.1 7.795 42.27 8.305 ;
      RECT 33.885 7.8 34.055 8.31 ;
      RECT 32.895 0.57 33.065 1.08 ;
      RECT 32.895 2.39 33.065 3.86 ;
      RECT 32.895 5.02 33.065 6.49 ;
      RECT 32.895 7.8 33.065 8.31 ;
      RECT 31.535 0.575 31.705 3.865 ;
      RECT 31.535 5.015 31.705 8.305 ;
      RECT 31.105 0.575 31.275 1.085 ;
      RECT 31.105 1.655 31.275 3.865 ;
      RECT 31.105 5.015 31.275 7.225 ;
      RECT 31.105 7.795 31.275 8.305 ;
      RECT 28.715 2.85 29.085 3.22 ;
      RECT 26.755 5.015 26.925 8.305 ;
      RECT 26.325 5.015 26.495 7.225 ;
      RECT 26.325 7.795 26.495 8.305 ;
      RECT 18.105 7.8 18.275 8.31 ;
      RECT 17.115 0.57 17.285 1.08 ;
      RECT 17.115 2.39 17.285 3.86 ;
      RECT 17.115 5.02 17.285 6.49 ;
      RECT 17.115 7.8 17.285 8.31 ;
      RECT 15.755 0.575 15.925 3.865 ;
      RECT 15.755 5.015 15.925 8.305 ;
      RECT 15.325 0.575 15.495 1.085 ;
      RECT 15.325 1.655 15.495 3.865 ;
      RECT 15.325 5.015 15.495 7.225 ;
      RECT 15.325 7.795 15.495 8.305 ;
      RECT 12.935 2.85 13.305 3.22 ;
      RECT 10.975 5.015 11.145 8.305 ;
      RECT 10.545 5.015 10.715 7.225 ;
      RECT 10.545 7.795 10.715 8.305 ;
      RECT 1.61 5.015 1.78 7.225 ;
      RECT 1.61 7.795 1.78 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2aa_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2aa_8_b0r2
  CLASS BLOCK ;
  ORIGIN -1.485 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2aa_8_b0r2 ;
  SIZE 81.765 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 19.585 0.915 19.755 1.085 ;
        RECT 19.58 0.91 19.75 1.08 ;
        RECT 19.58 2.39 19.75 2.56 ;
      LAYER li1 ;
        RECT 19.585 0.915 19.755 1.085 ;
        RECT 19.58 0.57 19.75 1.08 ;
        RECT 19.58 2.39 19.75 3.86 ;
      LAYER met1 ;
        RECT 19.52 2.36 19.81 2.59 ;
        RECT 19.52 0.88 19.81 1.11 ;
        RECT 19.58 0.88 19.75 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 35.365 0.915 35.535 1.085 ;
        RECT 35.36 0.91 35.53 1.08 ;
        RECT 35.36 2.39 35.53 2.56 ;
      LAYER li1 ;
        RECT 35.365 0.915 35.535 1.085 ;
        RECT 35.36 0.57 35.53 1.08 ;
        RECT 35.36 2.39 35.53 3.86 ;
      LAYER met1 ;
        RECT 35.3 2.36 35.59 2.59 ;
        RECT 35.3 0.88 35.59 1.11 ;
        RECT 35.36 0.88 35.53 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 51.14 0.915 51.31 1.085 ;
        RECT 51.135 0.91 51.305 1.08 ;
        RECT 51.135 2.39 51.305 2.56 ;
      LAYER li1 ;
        RECT 51.14 0.915 51.31 1.085 ;
        RECT 51.135 0.57 51.305 1.08 ;
        RECT 51.135 2.39 51.305 3.86 ;
      LAYER met1 ;
        RECT 51.075 2.36 51.365 2.59 ;
        RECT 51.075 0.88 51.365 1.11 ;
        RECT 51.135 0.88 51.305 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 66.925 0.915 67.095 1.085 ;
        RECT 66.92 0.91 67.09 1.08 ;
        RECT 66.92 2.39 67.09 2.56 ;
      LAYER li1 ;
        RECT 66.925 0.915 67.095 1.085 ;
        RECT 66.92 0.57 67.09 1.08 ;
        RECT 66.92 2.39 67.09 3.86 ;
      LAYER met1 ;
        RECT 66.86 2.36 67.15 2.59 ;
        RECT 66.86 0.88 67.15 1.11 ;
        RECT 66.92 0.88 67.09 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 82.71 0.915 82.88 1.085 ;
        RECT 82.705 0.91 82.875 1.08 ;
        RECT 82.705 2.39 82.875 2.56 ;
      LAYER li1 ;
        RECT 82.71 0.915 82.88 1.085 ;
        RECT 82.705 0.57 82.875 1.08 ;
        RECT 82.705 2.39 82.875 3.86 ;
      LAYER met1 ;
        RECT 82.645 2.36 82.935 2.59 ;
        RECT 82.645 0.88 82.935 1.11 ;
        RECT 82.705 0.88 82.875 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 15.345 5.855 15.695 6.205 ;
        RECT 15.34 2.705 15.69 3.055 ;
        RECT 15.415 2.705 15.59 6.205 ;
      LAYER li1 ;
        RECT 15.43 1.66 15.6 2.935 ;
        RECT 15.43 5.945 15.6 7.22 ;
        RECT 10.65 5.945 10.82 7.22 ;
      LAYER met1 ;
        RECT 15.34 2.765 15.83 2.935 ;
        RECT 15.34 2.705 15.69 3.055 ;
        RECT 10.59 5.945 15.83 6.115 ;
        RECT 15.345 5.855 15.695 6.205 ;
        RECT 10.59 5.915 10.88 6.145 ;
      LAYER via1 ;
        RECT 15.44 2.805 15.59 2.955 ;
        RECT 15.445 5.955 15.595 6.105 ;
      LAYER mcon ;
        RECT 10.65 5.945 10.82 6.115 ;
        RECT 15.43 5.945 15.6 6.115 ;
        RECT 15.43 2.765 15.6 2.935 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 31.125 5.855 31.475 6.205 ;
        RECT 31.12 2.705 31.47 3.055 ;
        RECT 31.195 2.705 31.37 6.205 ;
      LAYER li1 ;
        RECT 31.21 1.66 31.38 2.935 ;
        RECT 31.21 5.945 31.38 7.22 ;
        RECT 26.43 5.945 26.6 7.22 ;
      LAYER met1 ;
        RECT 31.12 2.765 31.61 2.935 ;
        RECT 31.12 2.705 31.47 3.055 ;
        RECT 26.37 5.945 31.61 6.115 ;
        RECT 31.125 5.855 31.475 6.205 ;
        RECT 26.37 5.915 26.66 6.145 ;
      LAYER via1 ;
        RECT 31.22 2.805 31.37 2.955 ;
        RECT 31.225 5.955 31.375 6.105 ;
      LAYER mcon ;
        RECT 26.43 5.945 26.6 6.115 ;
        RECT 31.21 5.945 31.38 6.115 ;
        RECT 31.21 2.765 31.38 2.935 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 46.9 5.855 47.25 6.205 ;
        RECT 46.895 2.705 47.245 3.055 ;
        RECT 46.97 2.705 47.145 6.205 ;
      LAYER li1 ;
        RECT 46.985 1.66 47.155 2.935 ;
        RECT 46.985 5.945 47.155 7.22 ;
        RECT 42.205 5.945 42.375 7.22 ;
      LAYER met1 ;
        RECT 46.895 2.765 47.385 2.935 ;
        RECT 46.895 2.705 47.245 3.055 ;
        RECT 42.145 5.945 47.385 6.115 ;
        RECT 46.9 5.855 47.25 6.205 ;
        RECT 42.145 5.915 42.435 6.145 ;
      LAYER via1 ;
        RECT 46.995 2.805 47.145 2.955 ;
        RECT 47 5.955 47.15 6.105 ;
      LAYER mcon ;
        RECT 42.205 5.945 42.375 6.115 ;
        RECT 46.985 5.945 47.155 6.115 ;
        RECT 46.985 2.765 47.155 2.935 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 62.685 5.855 63.035 6.205 ;
        RECT 62.68 2.705 63.03 3.055 ;
        RECT 62.755 2.705 62.93 6.205 ;
      LAYER li1 ;
        RECT 62.77 1.66 62.94 2.935 ;
        RECT 62.77 5.945 62.94 7.22 ;
        RECT 57.99 5.945 58.16 7.22 ;
      LAYER met1 ;
        RECT 62.68 2.765 63.17 2.935 ;
        RECT 62.68 2.705 63.03 3.055 ;
        RECT 57.93 5.945 63.17 6.115 ;
        RECT 62.685 5.855 63.035 6.205 ;
        RECT 57.93 5.915 58.22 6.145 ;
      LAYER via1 ;
        RECT 62.78 2.805 62.93 2.955 ;
        RECT 62.785 5.955 62.935 6.105 ;
      LAYER mcon ;
        RECT 57.99 5.945 58.16 6.115 ;
        RECT 62.77 5.945 62.94 6.115 ;
        RECT 62.77 2.765 62.94 2.935 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 78.47 5.855 78.82 6.205 ;
        RECT 78.465 2.705 78.815 3.055 ;
        RECT 78.54 2.705 78.715 6.205 ;
      LAYER li1 ;
        RECT 78.555 1.66 78.725 2.935 ;
        RECT 78.555 5.945 78.725 7.22 ;
        RECT 73.775 5.945 73.945 7.22 ;
      LAYER met1 ;
        RECT 78.465 2.765 78.955 2.935 ;
        RECT 78.465 2.705 78.815 3.055 ;
        RECT 73.715 5.945 78.955 6.115 ;
        RECT 78.47 5.855 78.82 6.205 ;
        RECT 73.715 5.915 74.005 6.145 ;
      LAYER via1 ;
        RECT 78.565 2.805 78.715 2.955 ;
        RECT 78.57 5.955 78.72 6.105 ;
      LAYER mcon ;
        RECT 73.775 5.945 73.945 6.115 ;
        RECT 78.555 5.945 78.725 6.115 ;
        RECT 78.555 2.765 78.725 2.935 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 1.715 5.945 1.885 7.22 ;
      LAYER met1 ;
        RECT 1.655 5.945 2.115 6.115 ;
        RECT 1.655 5.915 1.945 6.145 ;
      LAYER mcon ;
        RECT 1.715 5.945 1.885 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.485 4.135 83.25 4.745 ;
        RECT 81.115 4.13 83.095 4.75 ;
        RECT 82.275 3.4 82.445 5.48 ;
        RECT 81.285 3.4 81.455 5.48 ;
        RECT 78.545 3.405 78.715 5.475 ;
        RECT 76.745 3.635 76.915 4.745 ;
        RECT 75.785 3.635 75.955 4.745 ;
        RECT 73.765 4.135 73.935 5.475 ;
        RECT 73.345 3.635 73.515 4.745 ;
        RECT 72.345 3.635 72.515 4.745 ;
        RECT 71.385 3.635 71.555 4.745 ;
        RECT 68.945 3.635 69.115 4.745 ;
        RECT 65.33 4.13 67.31 4.75 ;
        RECT 66.49 3.4 66.66 5.48 ;
        RECT 65.5 3.4 65.67 5.48 ;
        RECT 62.76 3.405 62.93 5.475 ;
        RECT 60.96 3.635 61.13 4.745 ;
        RECT 60 3.635 60.17 4.745 ;
        RECT 57.98 4.135 58.15 5.475 ;
        RECT 57.56 3.635 57.73 4.745 ;
        RECT 56.56 3.635 56.73 4.745 ;
        RECT 55.6 3.635 55.77 4.745 ;
        RECT 53.16 3.635 53.33 4.745 ;
        RECT 49.545 4.13 51.525 4.75 ;
        RECT 50.705 3.4 50.875 5.48 ;
        RECT 49.715 3.4 49.885 5.48 ;
        RECT 46.975 3.405 47.145 5.475 ;
        RECT 45.175 3.635 45.345 4.745 ;
        RECT 44.215 3.635 44.385 4.745 ;
        RECT 42.195 4.135 42.365 5.475 ;
        RECT 41.775 3.635 41.945 4.745 ;
        RECT 40.775 3.635 40.945 4.745 ;
        RECT 39.815 3.635 39.985 4.745 ;
        RECT 37.375 3.635 37.545 4.745 ;
        RECT 33.77 4.13 35.75 4.75 ;
        RECT 34.93 3.4 35.1 5.48 ;
        RECT 33.94 3.4 34.11 5.48 ;
        RECT 31.2 3.405 31.37 5.475 ;
        RECT 29.4 3.635 29.57 4.745 ;
        RECT 28.44 3.635 28.61 4.745 ;
        RECT 26.42 4.135 26.59 5.475 ;
        RECT 26 3.635 26.17 4.745 ;
        RECT 25 3.635 25.17 4.745 ;
        RECT 24.04 3.635 24.21 4.745 ;
        RECT 21.6 3.635 21.77 4.745 ;
        RECT 17.99 4.13 19.97 4.75 ;
        RECT 19.15 3.4 19.32 5.48 ;
        RECT 18.16 3.4 18.33 5.48 ;
        RECT 15.42 3.405 15.59 5.475 ;
        RECT 13.62 3.635 13.79 4.745 ;
        RECT 12.66 3.635 12.83 4.745 ;
        RECT 10.64 4.135 10.81 5.475 ;
        RECT 10.22 3.635 10.39 4.745 ;
        RECT 9.22 3.635 9.39 4.745 ;
        RECT 8.26 3.635 8.43 4.745 ;
        RECT 5.82 3.635 5.99 4.745 ;
        RECT 3.515 4.135 3.685 8.305 ;
        RECT 1.705 4.135 1.875 5.475 ;
      LAYER met1 ;
        RECT 73.34 4.135 83.25 4.745 ;
        RECT 81.115 4.13 83.095 4.75 ;
        RECT 67.655 3.98 77.315 4.74 ;
        RECT 57.555 4.135 72.955 4.745 ;
        RECT 65.33 4.13 67.31 4.75 ;
        RECT 51.87 3.98 61.53 4.74 ;
        RECT 41.77 4.135 57.17 4.745 ;
        RECT 49.545 4.13 51.525 4.75 ;
        RECT 36.085 3.98 45.745 4.74 ;
        RECT 25.995 4.135 41.385 4.745 ;
        RECT 33.77 4.13 35.75 4.75 ;
        RECT 20.31 3.98 29.97 4.74 ;
        RECT 10.215 4.135 25.61 4.745 ;
        RECT 17.99 4.13 19.97 4.75 ;
        RECT 4.53 3.98 14.19 4.74 ;
        RECT 1.485 4.135 9.83 4.745 ;
        RECT 3.455 6.655 3.745 6.885 ;
        RECT 3.285 6.685 3.745 6.855 ;
      LAYER mcon ;
        RECT 3.515 6.685 3.685 6.855 ;
        RECT 3.825 4.545 3.995 4.715 ;
        RECT 4.675 4.135 4.845 4.305 ;
        RECT 5.135 4.135 5.305 4.305 ;
        RECT 5.595 4.135 5.765 4.305 ;
        RECT 6.055 4.135 6.225 4.305 ;
        RECT 6.515 4.135 6.685 4.305 ;
        RECT 6.975 4.135 7.145 4.305 ;
        RECT 7.435 4.135 7.605 4.305 ;
        RECT 7.895 4.135 8.065 4.305 ;
        RECT 8.355 4.135 8.525 4.305 ;
        RECT 8.815 4.135 8.985 4.305 ;
        RECT 9.275 4.135 9.445 4.305 ;
        RECT 9.735 4.135 9.905 4.305 ;
        RECT 10.195 4.135 10.365 4.305 ;
        RECT 10.655 4.135 10.825 4.305 ;
        RECT 11.115 4.135 11.285 4.305 ;
        RECT 11.575 4.135 11.745 4.305 ;
        RECT 12.035 4.135 12.205 4.305 ;
        RECT 12.495 4.135 12.665 4.305 ;
        RECT 12.76 4.545 12.93 4.715 ;
        RECT 12.955 4.135 13.125 4.305 ;
        RECT 13.415 4.135 13.585 4.305 ;
        RECT 13.875 4.135 14.045 4.305 ;
        RECT 17.54 4.545 17.71 4.715 ;
        RECT 17.54 4.165 17.71 4.335 ;
        RECT 18.24 4.55 18.41 4.72 ;
        RECT 18.24 4.16 18.41 4.33 ;
        RECT 19.23 4.55 19.4 4.72 ;
        RECT 19.23 4.16 19.4 4.33 ;
        RECT 20.455 4.135 20.625 4.305 ;
        RECT 20.915 4.135 21.085 4.305 ;
        RECT 21.375 4.135 21.545 4.305 ;
        RECT 21.835 4.135 22.005 4.305 ;
        RECT 22.295 4.135 22.465 4.305 ;
        RECT 22.755 4.135 22.925 4.305 ;
        RECT 23.215 4.135 23.385 4.305 ;
        RECT 23.675 4.135 23.845 4.305 ;
        RECT 24.135 4.135 24.305 4.305 ;
        RECT 24.595 4.135 24.765 4.305 ;
        RECT 25.055 4.135 25.225 4.305 ;
        RECT 25.515 4.135 25.685 4.305 ;
        RECT 25.975 4.135 26.145 4.305 ;
        RECT 26.435 4.135 26.605 4.305 ;
        RECT 26.895 4.135 27.065 4.305 ;
        RECT 27.355 4.135 27.525 4.305 ;
        RECT 27.815 4.135 27.985 4.305 ;
        RECT 28.275 4.135 28.445 4.305 ;
        RECT 28.54 4.545 28.71 4.715 ;
        RECT 28.735 4.135 28.905 4.305 ;
        RECT 29.195 4.135 29.365 4.305 ;
        RECT 29.655 4.135 29.825 4.305 ;
        RECT 33.32 4.545 33.49 4.715 ;
        RECT 33.32 4.165 33.49 4.335 ;
        RECT 34.02 4.55 34.19 4.72 ;
        RECT 34.02 4.16 34.19 4.33 ;
        RECT 35.01 4.55 35.18 4.72 ;
        RECT 35.01 4.16 35.18 4.33 ;
        RECT 36.23 4.135 36.4 4.305 ;
        RECT 36.69 4.135 36.86 4.305 ;
        RECT 37.15 4.135 37.32 4.305 ;
        RECT 37.61 4.135 37.78 4.305 ;
        RECT 38.07 4.135 38.24 4.305 ;
        RECT 38.53 4.135 38.7 4.305 ;
        RECT 38.99 4.135 39.16 4.305 ;
        RECT 39.45 4.135 39.62 4.305 ;
        RECT 39.91 4.135 40.08 4.305 ;
        RECT 40.37 4.135 40.54 4.305 ;
        RECT 40.83 4.135 41 4.305 ;
        RECT 41.29 4.135 41.46 4.305 ;
        RECT 41.75 4.135 41.92 4.305 ;
        RECT 42.21 4.135 42.38 4.305 ;
        RECT 42.67 4.135 42.84 4.305 ;
        RECT 43.13 4.135 43.3 4.305 ;
        RECT 43.59 4.135 43.76 4.305 ;
        RECT 44.05 4.135 44.22 4.305 ;
        RECT 44.315 4.545 44.485 4.715 ;
        RECT 44.51 4.135 44.68 4.305 ;
        RECT 44.97 4.135 45.14 4.305 ;
        RECT 45.43 4.135 45.6 4.305 ;
        RECT 49.095 4.545 49.265 4.715 ;
        RECT 49.095 4.165 49.265 4.335 ;
        RECT 49.795 4.55 49.965 4.72 ;
        RECT 49.795 4.16 49.965 4.33 ;
        RECT 50.785 4.55 50.955 4.72 ;
        RECT 50.785 4.16 50.955 4.33 ;
        RECT 52.015 4.135 52.185 4.305 ;
        RECT 52.475 4.135 52.645 4.305 ;
        RECT 52.935 4.135 53.105 4.305 ;
        RECT 53.395 4.135 53.565 4.305 ;
        RECT 53.855 4.135 54.025 4.305 ;
        RECT 54.315 4.135 54.485 4.305 ;
        RECT 54.775 4.135 54.945 4.305 ;
        RECT 55.235 4.135 55.405 4.305 ;
        RECT 55.695 4.135 55.865 4.305 ;
        RECT 56.155 4.135 56.325 4.305 ;
        RECT 56.615 4.135 56.785 4.305 ;
        RECT 57.075 4.135 57.245 4.305 ;
        RECT 57.535 4.135 57.705 4.305 ;
        RECT 57.995 4.135 58.165 4.305 ;
        RECT 58.455 4.135 58.625 4.305 ;
        RECT 58.915 4.135 59.085 4.305 ;
        RECT 59.375 4.135 59.545 4.305 ;
        RECT 59.835 4.135 60.005 4.305 ;
        RECT 60.1 4.545 60.27 4.715 ;
        RECT 60.295 4.135 60.465 4.305 ;
        RECT 60.755 4.135 60.925 4.305 ;
        RECT 61.215 4.135 61.385 4.305 ;
        RECT 64.88 4.545 65.05 4.715 ;
        RECT 64.88 4.165 65.05 4.335 ;
        RECT 65.58 4.55 65.75 4.72 ;
        RECT 65.58 4.16 65.75 4.33 ;
        RECT 66.57 4.55 66.74 4.72 ;
        RECT 66.57 4.16 66.74 4.33 ;
        RECT 67.8 4.135 67.97 4.305 ;
        RECT 68.26 4.135 68.43 4.305 ;
        RECT 68.72 4.135 68.89 4.305 ;
        RECT 69.18 4.135 69.35 4.305 ;
        RECT 69.64 4.135 69.81 4.305 ;
        RECT 70.1 4.135 70.27 4.305 ;
        RECT 70.56 4.135 70.73 4.305 ;
        RECT 71.02 4.135 71.19 4.305 ;
        RECT 71.48 4.135 71.65 4.305 ;
        RECT 71.94 4.135 72.11 4.305 ;
        RECT 72.4 4.135 72.57 4.305 ;
        RECT 72.86 4.135 73.03 4.305 ;
        RECT 73.32 4.135 73.49 4.305 ;
        RECT 73.78 4.135 73.95 4.305 ;
        RECT 74.24 4.135 74.41 4.305 ;
        RECT 74.7 4.135 74.87 4.305 ;
        RECT 75.16 4.135 75.33 4.305 ;
        RECT 75.62 4.135 75.79 4.305 ;
        RECT 75.885 4.545 76.055 4.715 ;
        RECT 76.08 4.135 76.25 4.305 ;
        RECT 76.54 4.135 76.71 4.305 ;
        RECT 77 4.135 77.17 4.305 ;
        RECT 80.665 4.545 80.835 4.715 ;
        RECT 80.665 4.165 80.835 4.335 ;
        RECT 81.365 4.55 81.535 4.72 ;
        RECT 81.365 4.16 81.535 4.33 ;
        RECT 82.355 4.55 82.525 4.72 ;
        RECT 82.355 4.16 82.525 4.33 ;
    END
  END vccd1
  OBS
    LAYER met3 ;
      RECT 75.045 7.04 75.415 7.41 ;
      RECT 75.085 6.72 75.415 7.41 ;
      RECT 75.085 6.72 77.875 7.025 ;
      RECT 77.57 2.85 77.875 7.025 ;
      RECT 77.535 2.85 77.905 3.22 ;
      RECT 76.795 0.815 77.1 4.02 ;
      RECT 76.545 2.975 77.1 3.705 ;
      RECT 76.755 0.815 77.125 1.185 ;
      RECT 72.905 1.85 73.235 2.745 ;
      RECT 72.025 2.015 72.355 2.745 ;
      RECT 72.9 1.85 73.27 2.65 ;
      RECT 76.065 1.85 76.395 2.58 ;
      RECT 76.025 1.735 76.205 2.385 ;
      RECT 72.035 1.85 76.395 2.22 ;
      RECT 72.525 3.535 72.855 3.865 ;
      RECT 71.32 3.55 72.855 3.85 ;
      RECT 71.32 2.43 71.62 3.85 ;
      RECT 71.065 2.415 71.395 2.745 ;
      RECT 59.26 7.04 59.63 7.41 ;
      RECT 59.3 6.72 59.63 7.41 ;
      RECT 59.3 6.72 62.09 7.025 ;
      RECT 61.785 2.85 62.09 7.025 ;
      RECT 61.75 2.85 62.12 3.22 ;
      RECT 61.01 0.815 61.315 4.02 ;
      RECT 60.76 2.975 61.315 3.705 ;
      RECT 60.97 0.815 61.34 1.185 ;
      RECT 57.12 1.85 57.45 2.745 ;
      RECT 56.24 2.015 56.57 2.745 ;
      RECT 57.115 1.85 57.485 2.65 ;
      RECT 60.28 1.85 60.61 2.58 ;
      RECT 60.24 1.735 60.42 2.385 ;
      RECT 56.25 1.85 60.61 2.22 ;
      RECT 56.74 3.535 57.07 3.865 ;
      RECT 55.535 3.55 57.07 3.85 ;
      RECT 55.535 2.43 55.835 3.85 ;
      RECT 55.28 2.415 55.61 2.745 ;
      RECT 43.475 7.04 43.845 7.41 ;
      RECT 43.515 6.72 43.845 7.41 ;
      RECT 43.515 6.72 46.305 7.025 ;
      RECT 46 2.85 46.305 7.025 ;
      RECT 45.965 2.85 46.335 3.22 ;
      RECT 45.225 0.815 45.53 4.02 ;
      RECT 44.975 2.975 45.53 3.705 ;
      RECT 45.185 0.815 45.555 1.185 ;
      RECT 41.335 1.85 41.665 2.745 ;
      RECT 40.455 2.015 40.785 2.745 ;
      RECT 41.33 1.85 41.7 2.65 ;
      RECT 44.495 1.85 44.825 2.58 ;
      RECT 44.455 1.735 44.635 2.385 ;
      RECT 40.465 1.85 44.825 2.22 ;
      RECT 40.955 3.535 41.285 3.865 ;
      RECT 39.75 3.55 41.285 3.85 ;
      RECT 39.75 2.43 40.05 3.85 ;
      RECT 39.495 2.415 39.825 2.745 ;
      RECT 27.7 7.04 28.07 7.41 ;
      RECT 27.74 6.72 28.07 7.41 ;
      RECT 27.74 6.72 30.53 7.025 ;
      RECT 30.225 2.85 30.53 7.025 ;
      RECT 30.19 2.85 30.56 3.22 ;
      RECT 29.45 0.815 29.755 4.02 ;
      RECT 29.2 2.975 29.755 3.705 ;
      RECT 29.41 0.815 29.78 1.185 ;
      RECT 25.56 1.85 25.89 2.745 ;
      RECT 24.68 2.015 25.01 2.745 ;
      RECT 25.555 1.85 25.925 2.65 ;
      RECT 28.72 1.85 29.05 2.58 ;
      RECT 28.68 1.735 28.86 2.385 ;
      RECT 24.69 1.85 29.05 2.22 ;
      RECT 25.18 3.535 25.51 3.865 ;
      RECT 23.975 3.55 25.51 3.85 ;
      RECT 23.975 2.43 24.275 3.85 ;
      RECT 23.72 2.415 24.05 2.745 ;
      RECT 11.92 7.04 12.29 7.41 ;
      RECT 11.96 6.72 12.29 7.41 ;
      RECT 11.96 6.72 14.75 7.025 ;
      RECT 14.445 2.85 14.75 7.025 ;
      RECT 14.41 2.85 14.78 3.22 ;
      RECT 13.67 0.815 13.975 4.02 ;
      RECT 13.42 2.975 13.975 3.705 ;
      RECT 13.63 0.815 14 1.185 ;
      RECT 9.78 1.85 10.11 2.745 ;
      RECT 8.9 2.015 9.23 2.745 ;
      RECT 9.775 1.85 10.145 2.65 ;
      RECT 12.94 1.85 13.27 2.58 ;
      RECT 12.9 1.735 13.08 2.385 ;
      RECT 8.91 1.85 13.27 2.22 ;
      RECT 9.4 3.535 9.73 3.865 ;
      RECT 8.195 3.55 9.73 3.85 ;
      RECT 8.195 2.43 8.495 3.85 ;
      RECT 7.94 2.415 8.27 2.745 ;
      RECT 74.465 2.575 74.795 3.305 ;
      RECT 70.345 2.415 70.675 3.145 ;
      RECT 69.345 1.855 69.675 2.585 ;
      RECT 67.905 2.575 68.235 3.305 ;
      RECT 58.68 2.575 59.01 3.305 ;
      RECT 54.56 2.415 54.89 3.145 ;
      RECT 53.56 1.855 53.89 2.585 ;
      RECT 52.12 2.575 52.45 3.305 ;
      RECT 42.895 2.575 43.225 3.305 ;
      RECT 38.775 2.415 39.105 3.145 ;
      RECT 37.775 1.855 38.105 2.585 ;
      RECT 36.335 2.575 36.665 3.305 ;
      RECT 27.12 2.575 27.45 3.305 ;
      RECT 23 2.415 23.33 3.145 ;
      RECT 22 1.855 22.33 2.585 ;
      RECT 20.56 2.575 20.89 3.305 ;
      RECT 11.34 2.575 11.67 3.305 ;
      RECT 7.22 2.415 7.55 3.145 ;
      RECT 6.22 1.855 6.55 2.585 ;
      RECT 4.78 2.575 5.11 3.305 ;
    LAYER via2 ;
      RECT 77.62 2.935 77.82 3.135 ;
      RECT 76.84 0.9 77.04 1.1 ;
      RECT 76.61 3.04 76.81 3.24 ;
      RECT 76.13 2.315 76.33 2.515 ;
      RECT 75.13 7.125 75.33 7.325 ;
      RECT 74.53 3.04 74.73 3.24 ;
      RECT 72.97 2.48 73.17 2.68 ;
      RECT 72.59 3.6 72.79 3.8 ;
      RECT 72.09 2.48 72.29 2.68 ;
      RECT 71.13 2.48 71.33 2.68 ;
      RECT 70.41 2.48 70.61 2.68 ;
      RECT 69.41 1.92 69.61 2.12 ;
      RECT 67.97 3.04 68.17 3.24 ;
      RECT 61.835 2.935 62.035 3.135 ;
      RECT 61.055 0.9 61.255 1.1 ;
      RECT 60.825 3.04 61.025 3.24 ;
      RECT 60.345 2.315 60.545 2.515 ;
      RECT 59.345 7.125 59.545 7.325 ;
      RECT 58.745 3.04 58.945 3.24 ;
      RECT 57.185 2.48 57.385 2.68 ;
      RECT 56.805 3.6 57.005 3.8 ;
      RECT 56.305 2.48 56.505 2.68 ;
      RECT 55.345 2.48 55.545 2.68 ;
      RECT 54.625 2.48 54.825 2.68 ;
      RECT 53.625 1.92 53.825 2.12 ;
      RECT 52.185 3.04 52.385 3.24 ;
      RECT 46.05 2.935 46.25 3.135 ;
      RECT 45.27 0.9 45.47 1.1 ;
      RECT 45.04 3.04 45.24 3.24 ;
      RECT 44.56 2.315 44.76 2.515 ;
      RECT 43.56 7.125 43.76 7.325 ;
      RECT 42.96 3.04 43.16 3.24 ;
      RECT 41.4 2.48 41.6 2.68 ;
      RECT 41.02 3.6 41.22 3.8 ;
      RECT 40.52 2.48 40.72 2.68 ;
      RECT 39.56 2.48 39.76 2.68 ;
      RECT 38.84 2.48 39.04 2.68 ;
      RECT 37.84 1.92 38.04 2.12 ;
      RECT 36.4 3.04 36.6 3.24 ;
      RECT 30.275 2.935 30.475 3.135 ;
      RECT 29.495 0.9 29.695 1.1 ;
      RECT 29.265 3.04 29.465 3.24 ;
      RECT 28.785 2.315 28.985 2.515 ;
      RECT 27.785 7.125 27.985 7.325 ;
      RECT 27.185 3.04 27.385 3.24 ;
      RECT 25.625 2.48 25.825 2.68 ;
      RECT 25.245 3.6 25.445 3.8 ;
      RECT 24.745 2.48 24.945 2.68 ;
      RECT 23.785 2.48 23.985 2.68 ;
      RECT 23.065 2.48 23.265 2.68 ;
      RECT 22.065 1.92 22.265 2.12 ;
      RECT 20.625 3.04 20.825 3.24 ;
      RECT 14.495 2.935 14.695 3.135 ;
      RECT 13.715 0.9 13.915 1.1 ;
      RECT 13.485 3.04 13.685 3.24 ;
      RECT 13.005 2.315 13.205 2.515 ;
      RECT 12.005 7.125 12.205 7.325 ;
      RECT 11.405 3.04 11.605 3.24 ;
      RECT 9.845 2.48 10.045 2.68 ;
      RECT 9.465 3.6 9.665 3.8 ;
      RECT 8.965 2.48 9.165 2.68 ;
      RECT 8.005 2.48 8.205 2.68 ;
      RECT 7.285 2.48 7.485 2.68 ;
      RECT 6.285 1.92 6.485 2.12 ;
      RECT 4.845 3.04 5.045 3.24 ;
    LAYER met2 ;
      RECT 2.71 8.4 82.88 8.57 ;
      RECT 82.71 7.275 82.88 8.57 ;
      RECT 2.71 6.255 2.88 8.57 ;
      RECT 82.68 7.275 83.03 7.625 ;
      RECT 2.65 6.255 2.94 6.605 ;
      RECT 79.52 6.22 79.84 6.545 ;
      RECT 79.55 5.695 79.72 6.545 ;
      RECT 79.55 5.695 79.725 6.045 ;
      RECT 79.55 5.695 80.525 5.87 ;
      RECT 80.35 1.965 80.525 5.87 ;
      RECT 80.295 1.965 80.645 2.315 ;
      RECT 80.32 6.655 80.645 6.98 ;
      RECT 79.205 6.745 80.645 6.915 ;
      RECT 79.205 2.395 79.365 6.915 ;
      RECT 79.52 2.365 79.84 2.685 ;
      RECT 79.205 2.395 79.84 2.565 ;
      RECT 67.93 3 68.21 3.28 ;
      RECT 67.9 3 68.21 3.265 ;
      RECT 67.895 3 68.21 3.263 ;
      RECT 67.89 1.33 68.06 3.257 ;
      RECT 67.885 2.967 68.155 3.25 ;
      RECT 67.88 3 68.21 3.243 ;
      RECT 67.85 2.97 68.155 3.23 ;
      RECT 67.85 2.997 68.175 3.23 ;
      RECT 67.85 2.987 68.17 3.23 ;
      RECT 67.85 2.972 68.165 3.23 ;
      RECT 67.89 2.962 68.155 3.257 ;
      RECT 67.89 2.957 68.145 3.257 ;
      RECT 67.89 2.956 68.13 3.257 ;
      RECT 77.86 1.34 78.21 1.69 ;
      RECT 77.855 1.34 78.21 1.595 ;
      RECT 67.89 1.33 78.1 1.5 ;
      RECT 77.535 2.85 77.905 3.22 ;
      RECT 77.62 2.235 77.79 3.22 ;
      RECT 73.64 2.455 73.875 2.715 ;
      RECT 76.785 2.235 76.95 2.495 ;
      RECT 76.69 2.225 76.705 2.495 ;
      RECT 76.785 2.235 77.79 2.415 ;
      RECT 75.29 1.795 75.33 1.935 ;
      RECT 76.705 2.23 76.785 2.495 ;
      RECT 76.65 2.225 76.69 2.461 ;
      RECT 76.636 2.225 76.65 2.461 ;
      RECT 76.55 2.23 76.636 2.463 ;
      RECT 76.505 2.237 76.55 2.465 ;
      RECT 76.475 2.237 76.505 2.467 ;
      RECT 76.45 2.232 76.475 2.469 ;
      RECT 76.42 2.228 76.45 2.478 ;
      RECT 76.41 2.225 76.42 2.49 ;
      RECT 76.405 2.225 76.41 2.498 ;
      RECT 76.4 2.225 76.405 2.503 ;
      RECT 76.39 2.224 76.4 2.513 ;
      RECT 76.385 2.223 76.39 2.523 ;
      RECT 76.37 2.222 76.385 2.528 ;
      RECT 76.342 2.219 76.37 2.555 ;
      RECT 76.256 2.211 76.342 2.555 ;
      RECT 76.17 2.2 76.256 2.555 ;
      RECT 76.13 2.185 76.17 2.555 ;
      RECT 76.09 2.159 76.13 2.555 ;
      RECT 76.085 2.141 76.09 2.367 ;
      RECT 76.075 2.137 76.085 2.357 ;
      RECT 76.06 2.127 76.075 2.344 ;
      RECT 76.04 2.111 76.06 2.329 ;
      RECT 76.025 2.096 76.04 2.314 ;
      RECT 76.015 2.085 76.025 2.304 ;
      RECT 75.99 2.069 76.015 2.293 ;
      RECT 75.985 2.056 75.99 2.283 ;
      RECT 75.98 2.052 75.985 2.278 ;
      RECT 75.925 2.038 75.98 2.256 ;
      RECT 75.886 2.019 75.925 2.22 ;
      RECT 75.8 1.993 75.886 2.173 ;
      RECT 75.796 1.975 75.8 2.139 ;
      RECT 75.71 1.956 75.796 2.117 ;
      RECT 75.705 1.938 75.71 2.095 ;
      RECT 75.7 1.936 75.705 2.093 ;
      RECT 75.69 1.935 75.7 2.088 ;
      RECT 75.63 1.922 75.69 2.074 ;
      RECT 75.585 1.9 75.63 2.053 ;
      RECT 75.525 1.877 75.585 2.032 ;
      RECT 75.461 1.852 75.525 2.007 ;
      RECT 75.375 1.822 75.461 1.976 ;
      RECT 75.36 1.802 75.375 1.955 ;
      RECT 75.33 1.797 75.36 1.946 ;
      RECT 75.277 1.795 75.29 1.935 ;
      RECT 75.191 1.795 75.277 1.937 ;
      RECT 75.105 1.795 75.191 1.939 ;
      RECT 75.085 1.795 75.105 1.943 ;
      RECT 75.04 1.797 75.085 1.954 ;
      RECT 75 1.807 75.04 1.97 ;
      RECT 74.996 1.816 75 1.978 ;
      RECT 74.91 1.836 74.996 1.994 ;
      RECT 74.9 1.855 74.91 2.012 ;
      RECT 74.895 1.857 74.9 2.015 ;
      RECT 74.885 1.861 74.895 2.018 ;
      RECT 74.865 1.866 74.885 2.028 ;
      RECT 74.835 1.876 74.865 2.048 ;
      RECT 74.83 1.883 74.835 2.062 ;
      RECT 74.82 1.887 74.83 2.069 ;
      RECT 74.805 1.895 74.82 2.08 ;
      RECT 74.795 1.905 74.805 2.091 ;
      RECT 74.785 1.912 74.795 2.099 ;
      RECT 74.76 1.925 74.785 2.114 ;
      RECT 74.696 1.961 74.76 2.153 ;
      RECT 74.61 2.024 74.696 2.217 ;
      RECT 74.575 2.075 74.61 2.27 ;
      RECT 74.57 2.092 74.575 2.287 ;
      RECT 74.555 2.101 74.57 2.294 ;
      RECT 74.535 2.116 74.555 2.308 ;
      RECT 74.53 2.127 74.535 2.318 ;
      RECT 74.51 2.14 74.53 2.328 ;
      RECT 74.505 2.15 74.51 2.338 ;
      RECT 74.49 2.155 74.505 2.347 ;
      RECT 74.48 2.165 74.49 2.358 ;
      RECT 74.45 2.182 74.48 2.375 ;
      RECT 74.44 2.2 74.45 2.393 ;
      RECT 74.425 2.211 74.44 2.404 ;
      RECT 74.385 2.235 74.425 2.42 ;
      RECT 74.35 2.269 74.385 2.437 ;
      RECT 74.32 2.292 74.35 2.449 ;
      RECT 74.305 2.302 74.32 2.458 ;
      RECT 74.265 2.312 74.305 2.469 ;
      RECT 74.245 2.323 74.265 2.481 ;
      RECT 74.24 2.327 74.245 2.488 ;
      RECT 74.225 2.331 74.24 2.493 ;
      RECT 74.215 2.336 74.225 2.498 ;
      RECT 74.21 2.339 74.215 2.501 ;
      RECT 74.18 2.345 74.21 2.508 ;
      RECT 74.145 2.355 74.18 2.522 ;
      RECT 74.085 2.37 74.145 2.542 ;
      RECT 74.03 2.39 74.085 2.566 ;
      RECT 74.001 2.405 74.03 2.584 ;
      RECT 73.915 2.425 74.001 2.609 ;
      RECT 73.91 2.44 73.915 2.629 ;
      RECT 73.9 2.443 73.91 2.63 ;
      RECT 73.875 2.45 73.9 2.715 ;
      RECT 76.57 2.943 76.85 3.28 ;
      RECT 76.57 2.953 76.855 3.238 ;
      RECT 76.57 2.962 76.86 3.135 ;
      RECT 76.57 2.977 76.865 3.003 ;
      RECT 76.57 2.805 76.83 3.28 ;
      RECT 66.87 6.655 67.22 7.005 ;
      RECT 75.695 6.61 76.045 6.96 ;
      RECT 66.87 6.685 76.045 6.885 ;
      RECT 74.29 3.685 74.3 3.875 ;
      RECT 72.55 3.56 72.83 3.84 ;
      RECT 75.595 2.5 75.6 2.985 ;
      RECT 75.49 2.5 75.55 2.76 ;
      RECT 75.815 3.47 75.82 3.545 ;
      RECT 75.805 3.337 75.815 3.58 ;
      RECT 75.795 3.172 75.805 3.601 ;
      RECT 75.79 3.042 75.795 3.617 ;
      RECT 75.78 2.932 75.79 3.633 ;
      RECT 75.775 2.831 75.78 3.65 ;
      RECT 75.77 2.813 75.775 3.66 ;
      RECT 75.765 2.795 75.77 3.67 ;
      RECT 75.755 2.77 75.765 3.685 ;
      RECT 75.75 2.75 75.755 3.7 ;
      RECT 75.73 2.5 75.75 3.725 ;
      RECT 75.715 2.5 75.73 3.758 ;
      RECT 75.685 2.5 75.715 3.78 ;
      RECT 75.665 2.5 75.685 3.794 ;
      RECT 75.645 2.5 75.665 3.31 ;
      RECT 75.66 3.377 75.665 3.799 ;
      RECT 75.655 3.407 75.66 3.801 ;
      RECT 75.65 3.42 75.655 3.804 ;
      RECT 75.645 3.43 75.65 3.808 ;
      RECT 75.64 2.5 75.645 3.228 ;
      RECT 75.64 3.44 75.645 3.81 ;
      RECT 75.635 2.5 75.64 3.205 ;
      RECT 75.625 3.462 75.64 3.81 ;
      RECT 75.62 2.5 75.635 3.15 ;
      RECT 75.615 3.487 75.625 3.81 ;
      RECT 75.615 2.5 75.62 3.095 ;
      RECT 75.605 2.5 75.615 3.043 ;
      RECT 75.61 3.5 75.615 3.811 ;
      RECT 75.605 3.512 75.61 3.812 ;
      RECT 75.6 2.5 75.605 3.003 ;
      RECT 75.6 3.525 75.605 3.813 ;
      RECT 75.585 3.54 75.6 3.814 ;
      RECT 75.59 2.5 75.595 2.965 ;
      RECT 75.585 2.5 75.59 2.93 ;
      RECT 75.58 2.5 75.585 2.905 ;
      RECT 75.575 3.567 75.585 3.816 ;
      RECT 75.57 2.5 75.58 2.863 ;
      RECT 75.57 3.585 75.575 3.817 ;
      RECT 75.565 2.5 75.57 2.823 ;
      RECT 75.565 3.592 75.57 3.818 ;
      RECT 75.56 2.5 75.565 2.795 ;
      RECT 75.555 3.61 75.565 3.819 ;
      RECT 75.55 2.5 75.56 2.775 ;
      RECT 75.545 3.63 75.555 3.821 ;
      RECT 75.535 3.647 75.545 3.822 ;
      RECT 75.5 3.67 75.535 3.825 ;
      RECT 75.445 3.688 75.5 3.831 ;
      RECT 75.359 3.696 75.445 3.84 ;
      RECT 75.273 3.707 75.359 3.851 ;
      RECT 75.187 3.717 75.273 3.862 ;
      RECT 75.101 3.727 75.187 3.874 ;
      RECT 75.015 3.737 75.101 3.885 ;
      RECT 74.995 3.743 75.015 3.891 ;
      RECT 74.915 3.745 74.995 3.895 ;
      RECT 74.91 3.744 74.915 3.9 ;
      RECT 74.902 3.743 74.91 3.9 ;
      RECT 74.816 3.739 74.902 3.898 ;
      RECT 74.73 3.731 74.816 3.895 ;
      RECT 74.644 3.722 74.73 3.891 ;
      RECT 74.558 3.714 74.644 3.888 ;
      RECT 74.472 3.706 74.558 3.884 ;
      RECT 74.386 3.697 74.472 3.881 ;
      RECT 74.3 3.689 74.386 3.877 ;
      RECT 74.245 3.682 74.29 3.875 ;
      RECT 74.16 3.675 74.245 3.873 ;
      RECT 74.086 3.667 74.16 3.869 ;
      RECT 74 3.659 74.086 3.866 ;
      RECT 73.997 3.655 74 3.864 ;
      RECT 73.911 3.651 73.997 3.863 ;
      RECT 73.825 3.643 73.911 3.86 ;
      RECT 73.74 3.638 73.825 3.857 ;
      RECT 73.654 3.635 73.74 3.854 ;
      RECT 73.568 3.633 73.654 3.851 ;
      RECT 73.482 3.63 73.568 3.848 ;
      RECT 73.396 3.627 73.482 3.845 ;
      RECT 73.31 3.624 73.396 3.842 ;
      RECT 73.234 3.622 73.31 3.839 ;
      RECT 73.148 3.619 73.234 3.836 ;
      RECT 73.062 3.616 73.148 3.834 ;
      RECT 72.976 3.614 73.062 3.831 ;
      RECT 72.89 3.611 72.976 3.828 ;
      RECT 72.83 3.602 72.89 3.826 ;
      RECT 75.34 3.22 75.415 3.48 ;
      RECT 75.32 3.2 75.325 3.48 ;
      RECT 74.64 2.985 74.745 3.28 ;
      RECT 69.085 2.96 69.155 3.22 ;
      RECT 74.98 2.835 74.985 3.206 ;
      RECT 74.97 2.89 74.975 3.206 ;
      RECT 75.275 2.06 75.335 2.32 ;
      RECT 75.33 3.215 75.34 3.48 ;
      RECT 75.325 3.205 75.33 3.48 ;
      RECT 75.245 3.152 75.32 3.48 ;
      RECT 75.27 2.06 75.275 2.34 ;
      RECT 75.26 2.06 75.27 2.36 ;
      RECT 75.245 2.06 75.26 2.39 ;
      RECT 75.23 2.06 75.245 2.433 ;
      RECT 75.225 3.095 75.245 3.48 ;
      RECT 75.215 2.06 75.23 2.47 ;
      RECT 75.21 3.075 75.225 3.48 ;
      RECT 75.21 2.06 75.215 2.493 ;
      RECT 75.2 2.06 75.21 2.518 ;
      RECT 75.17 3.042 75.21 3.48 ;
      RECT 75.175 2.06 75.2 2.568 ;
      RECT 75.17 2.06 75.175 2.623 ;
      RECT 75.165 2.06 75.17 2.665 ;
      RECT 75.155 3.005 75.17 3.48 ;
      RECT 75.16 2.06 75.165 2.708 ;
      RECT 75.155 2.06 75.16 2.773 ;
      RECT 75.15 2.06 75.155 2.795 ;
      RECT 75.15 2.993 75.155 3.345 ;
      RECT 75.145 2.06 75.15 2.863 ;
      RECT 75.145 2.985 75.15 3.328 ;
      RECT 75.14 2.06 75.145 2.908 ;
      RECT 75.135 2.967 75.145 3.305 ;
      RECT 75.135 2.06 75.14 2.945 ;
      RECT 75.125 2.06 75.135 3.285 ;
      RECT 75.12 2.06 75.125 3.268 ;
      RECT 75.115 2.06 75.12 3.253 ;
      RECT 75.11 2.06 75.115 3.238 ;
      RECT 75.09 2.06 75.11 3.228 ;
      RECT 75.085 2.06 75.09 3.218 ;
      RECT 75.075 2.06 75.085 3.214 ;
      RECT 75.07 2.337 75.075 3.213 ;
      RECT 75.065 2.36 75.07 3.212 ;
      RECT 75.06 2.39 75.065 3.211 ;
      RECT 75.055 2.417 75.06 3.21 ;
      RECT 75.05 2.445 75.055 3.21 ;
      RECT 75.045 2.472 75.05 3.21 ;
      RECT 75.04 2.492 75.045 3.21 ;
      RECT 75.035 2.52 75.04 3.21 ;
      RECT 75.025 2.562 75.035 3.21 ;
      RECT 75.015 2.607 75.025 3.209 ;
      RECT 75.01 2.66 75.015 3.208 ;
      RECT 75.005 2.692 75.01 3.207 ;
      RECT 75 2.712 75.005 3.206 ;
      RECT 74.995 2.75 75 3.206 ;
      RECT 74.99 2.772 74.995 3.206 ;
      RECT 74.985 2.797 74.99 3.206 ;
      RECT 74.975 2.862 74.98 3.206 ;
      RECT 74.96 2.922 74.97 3.206 ;
      RECT 74.945 2.932 74.96 3.206 ;
      RECT 74.925 2.942 74.945 3.206 ;
      RECT 74.895 2.947 74.925 3.203 ;
      RECT 74.835 2.957 74.895 3.2 ;
      RECT 74.815 2.966 74.835 3.205 ;
      RECT 74.79 2.972 74.815 3.218 ;
      RECT 74.77 2.977 74.79 3.233 ;
      RECT 74.745 2.982 74.77 3.28 ;
      RECT 74.616 2.984 74.64 3.28 ;
      RECT 74.53 2.979 74.616 3.28 ;
      RECT 74.49 2.976 74.53 3.28 ;
      RECT 74.44 2.978 74.49 3.26 ;
      RECT 74.41 2.982 74.44 3.26 ;
      RECT 74.331 2.992 74.41 3.26 ;
      RECT 74.245 3.007 74.331 3.261 ;
      RECT 74.195 3.017 74.245 3.262 ;
      RECT 74.187 3.02 74.195 3.262 ;
      RECT 74.101 3.022 74.187 3.263 ;
      RECT 74.015 3.026 74.101 3.263 ;
      RECT 73.929 3.03 74.015 3.264 ;
      RECT 73.843 3.033 73.929 3.265 ;
      RECT 73.757 3.037 73.843 3.265 ;
      RECT 73.671 3.041 73.757 3.266 ;
      RECT 73.585 3.044 73.671 3.267 ;
      RECT 73.499 3.048 73.585 3.267 ;
      RECT 73.413 3.052 73.499 3.268 ;
      RECT 73.327 3.056 73.413 3.269 ;
      RECT 73.241 3.059 73.327 3.269 ;
      RECT 73.155 3.063 73.241 3.27 ;
      RECT 73.125 3.065 73.155 3.27 ;
      RECT 73.039 3.068 73.125 3.271 ;
      RECT 72.953 3.072 73.039 3.272 ;
      RECT 72.867 3.076 72.953 3.273 ;
      RECT 72.781 3.079 72.867 3.273 ;
      RECT 72.695 3.083 72.781 3.274 ;
      RECT 72.66 3.088 72.695 3.275 ;
      RECT 72.605 3.098 72.66 3.282 ;
      RECT 72.58 3.11 72.605 3.292 ;
      RECT 72.545 3.123 72.58 3.3 ;
      RECT 72.505 3.14 72.545 3.323 ;
      RECT 72.485 3.153 72.505 3.35 ;
      RECT 72.455 3.165 72.485 3.378 ;
      RECT 72.45 3.173 72.455 3.398 ;
      RECT 72.445 3.176 72.45 3.408 ;
      RECT 72.395 3.188 72.445 3.442 ;
      RECT 72.385 3.203 72.395 3.475 ;
      RECT 72.375 3.209 72.385 3.488 ;
      RECT 72.365 3.216 72.375 3.5 ;
      RECT 72.34 3.229 72.365 3.518 ;
      RECT 72.325 3.244 72.34 3.54 ;
      RECT 72.315 3.252 72.325 3.556 ;
      RECT 72.3 3.261 72.315 3.571 ;
      RECT 72.29 3.271 72.3 3.585 ;
      RECT 72.271 3.284 72.29 3.602 ;
      RECT 72.185 3.329 72.271 3.667 ;
      RECT 72.17 3.374 72.185 3.725 ;
      RECT 72.165 3.383 72.17 3.738 ;
      RECT 72.155 3.39 72.165 3.743 ;
      RECT 72.15 3.395 72.155 3.747 ;
      RECT 72.13 3.405 72.15 3.754 ;
      RECT 72.105 3.425 72.13 3.768 ;
      RECT 72.07 3.45 72.105 3.788 ;
      RECT 72.055 3.473 72.07 3.803 ;
      RECT 72.045 3.483 72.055 3.808 ;
      RECT 72.035 3.491 72.045 3.815 ;
      RECT 72.025 3.5 72.035 3.821 ;
      RECT 72.005 3.512 72.025 3.823 ;
      RECT 71.995 3.525 72.005 3.825 ;
      RECT 71.97 3.54 71.995 3.828 ;
      RECT 71.95 3.557 71.97 3.832 ;
      RECT 71.91 3.585 71.95 3.838 ;
      RECT 71.845 3.632 71.91 3.847 ;
      RECT 71.83 3.665 71.845 3.855 ;
      RECT 71.825 3.672 71.83 3.857 ;
      RECT 71.775 3.697 71.825 3.862 ;
      RECT 71.76 3.721 71.775 3.869 ;
      RECT 71.71 3.726 71.76 3.87 ;
      RECT 71.624 3.73 71.71 3.87 ;
      RECT 71.538 3.73 71.624 3.87 ;
      RECT 71.452 3.73 71.538 3.871 ;
      RECT 71.366 3.73 71.452 3.871 ;
      RECT 71.28 3.73 71.366 3.871 ;
      RECT 71.214 3.73 71.28 3.871 ;
      RECT 71.128 3.73 71.214 3.872 ;
      RECT 71.042 3.73 71.128 3.872 ;
      RECT 70.956 3.731 71.042 3.873 ;
      RECT 70.87 3.731 70.956 3.873 ;
      RECT 70.784 3.731 70.87 3.873 ;
      RECT 70.698 3.731 70.784 3.874 ;
      RECT 70.612 3.731 70.698 3.874 ;
      RECT 70.526 3.732 70.612 3.875 ;
      RECT 70.44 3.732 70.526 3.875 ;
      RECT 70.42 3.732 70.44 3.875 ;
      RECT 70.334 3.732 70.42 3.875 ;
      RECT 70.248 3.732 70.334 3.875 ;
      RECT 70.162 3.733 70.248 3.875 ;
      RECT 70.076 3.733 70.162 3.875 ;
      RECT 69.99 3.733 70.076 3.875 ;
      RECT 69.904 3.734 69.99 3.875 ;
      RECT 69.818 3.734 69.904 3.875 ;
      RECT 69.732 3.734 69.818 3.875 ;
      RECT 69.646 3.734 69.732 3.875 ;
      RECT 69.56 3.735 69.646 3.875 ;
      RECT 69.51 3.732 69.56 3.875 ;
      RECT 69.5 3.73 69.51 3.874 ;
      RECT 69.496 3.73 69.5 3.873 ;
      RECT 69.41 3.725 69.496 3.868 ;
      RECT 69.388 3.718 69.41 3.862 ;
      RECT 69.302 3.709 69.388 3.856 ;
      RECT 69.216 3.696 69.302 3.847 ;
      RECT 69.13 3.682 69.216 3.837 ;
      RECT 69.085 3.672 69.13 3.83 ;
      RECT 69.065 2.96 69.085 3.238 ;
      RECT 69.065 3.665 69.085 3.826 ;
      RECT 69.035 2.96 69.065 3.26 ;
      RECT 69.025 3.632 69.065 3.823 ;
      RECT 69.02 2.96 69.035 3.28 ;
      RECT 69.02 3.597 69.025 3.821 ;
      RECT 69.015 2.96 69.02 3.405 ;
      RECT 69.015 3.557 69.02 3.821 ;
      RECT 69.005 2.96 69.015 3.821 ;
      RECT 68.93 2.96 69.005 3.815 ;
      RECT 68.9 2.96 68.93 3.805 ;
      RECT 68.895 2.96 68.9 3.797 ;
      RECT 68.89 3.002 68.895 3.79 ;
      RECT 68.88 3.071 68.89 3.781 ;
      RECT 68.875 3.141 68.88 3.733 ;
      RECT 68.87 3.205 68.875 3.63 ;
      RECT 68.865 3.24 68.87 3.585 ;
      RECT 68.863 3.277 68.865 3.477 ;
      RECT 68.86 3.285 68.863 3.47 ;
      RECT 68.855 3.35 68.86 3.413 ;
      RECT 72.93 2.44 73.21 2.72 ;
      RECT 72.92 2.44 73.21 2.583 ;
      RECT 72.875 2.305 73.135 2.565 ;
      RECT 72.875 2.42 73.19 2.565 ;
      RECT 72.875 2.39 73.185 2.565 ;
      RECT 72.875 2.377 73.175 2.565 ;
      RECT 72.875 2.367 73.17 2.565 ;
      RECT 68.85 2.35 69.11 2.61 ;
      RECT 72.62 1.9 72.88 2.16 ;
      RECT 72.61 1.925 72.88 2.12 ;
      RECT 72.605 1.925 72.61 2.119 ;
      RECT 72.535 1.92 72.605 2.111 ;
      RECT 72.45 1.907 72.535 2.094 ;
      RECT 72.446 1.899 72.45 2.084 ;
      RECT 72.36 1.892 72.446 2.074 ;
      RECT 72.351 1.884 72.36 2.064 ;
      RECT 72.265 1.877 72.351 2.052 ;
      RECT 72.245 1.868 72.265 2.038 ;
      RECT 72.19 1.863 72.245 2.03 ;
      RECT 72.18 1.857 72.19 2.024 ;
      RECT 72.16 1.855 72.18 2.02 ;
      RECT 72.152 1.854 72.16 2.016 ;
      RECT 72.066 1.846 72.152 2.005 ;
      RECT 71.98 1.832 72.066 1.985 ;
      RECT 71.92 1.82 71.98 1.97 ;
      RECT 71.91 1.815 71.92 1.965 ;
      RECT 71.86 1.815 71.91 1.967 ;
      RECT 71.813 1.817 71.86 1.971 ;
      RECT 71.727 1.824 71.813 1.976 ;
      RECT 71.641 1.832 71.727 1.982 ;
      RECT 71.555 1.841 71.641 1.988 ;
      RECT 71.496 1.847 71.555 1.993 ;
      RECT 71.41 1.852 71.496 1.999 ;
      RECT 71.335 1.857 71.41 2.005 ;
      RECT 71.296 1.859 71.335 2.01 ;
      RECT 71.21 1.856 71.296 2.015 ;
      RECT 71.125 1.854 71.21 2.022 ;
      RECT 71.093 1.853 71.125 2.025 ;
      RECT 71.007 1.852 71.093 2.026 ;
      RECT 70.921 1.851 71.007 2.027 ;
      RECT 70.835 1.85 70.921 2.027 ;
      RECT 70.749 1.849 70.835 2.028 ;
      RECT 70.663 1.848 70.749 2.029 ;
      RECT 70.577 1.847 70.663 2.03 ;
      RECT 70.491 1.846 70.577 2.03 ;
      RECT 70.405 1.845 70.491 2.031 ;
      RECT 70.355 1.845 70.405 2.032 ;
      RECT 70.341 1.846 70.355 2.032 ;
      RECT 70.255 1.853 70.341 2.033 ;
      RECT 70.181 1.864 70.255 2.034 ;
      RECT 70.095 1.873 70.181 2.035 ;
      RECT 70.06 1.88 70.095 2.05 ;
      RECT 70.035 1.883 70.06 2.08 ;
      RECT 70.01 1.892 70.035 2.109 ;
      RECT 70 1.903 70.01 2.129 ;
      RECT 69.99 1.911 70 2.143 ;
      RECT 69.985 1.917 69.99 2.153 ;
      RECT 69.96 1.934 69.985 2.17 ;
      RECT 69.945 1.956 69.96 2.198 ;
      RECT 69.915 1.982 69.945 2.228 ;
      RECT 69.895 2.011 69.915 2.258 ;
      RECT 69.89 2.026 69.895 2.275 ;
      RECT 69.87 2.041 69.89 2.29 ;
      RECT 69.86 2.059 69.87 2.308 ;
      RECT 69.85 2.07 69.86 2.323 ;
      RECT 69.8 2.102 69.85 2.349 ;
      RECT 69.795 2.132 69.8 2.369 ;
      RECT 69.785 2.145 69.795 2.375 ;
      RECT 69.776 2.155 69.785 2.383 ;
      RECT 69.765 2.166 69.776 2.391 ;
      RECT 69.76 2.176 69.765 2.397 ;
      RECT 69.745 2.197 69.76 2.404 ;
      RECT 69.73 2.227 69.745 2.412 ;
      RECT 69.695 2.257 69.73 2.418 ;
      RECT 69.67 2.275 69.695 2.425 ;
      RECT 69.62 2.283 69.67 2.434 ;
      RECT 69.595 2.288 69.62 2.443 ;
      RECT 69.54 2.294 69.595 2.453 ;
      RECT 69.535 2.299 69.54 2.461 ;
      RECT 69.521 2.302 69.535 2.463 ;
      RECT 69.435 2.314 69.521 2.475 ;
      RECT 69.425 2.326 69.435 2.488 ;
      RECT 69.34 2.339 69.425 2.5 ;
      RECT 69.296 2.356 69.34 2.514 ;
      RECT 69.21 2.373 69.296 2.53 ;
      RECT 69.18 2.387 69.21 2.544 ;
      RECT 69.17 2.392 69.18 2.549 ;
      RECT 69.11 2.395 69.17 2.558 ;
      RECT 72 2.665 72.26 2.925 ;
      RECT 72 2.665 72.28 2.778 ;
      RECT 72 2.665 72.305 2.745 ;
      RECT 72 2.665 72.31 2.725 ;
      RECT 72.05 2.44 72.33 2.72 ;
      RECT 71.605 3.175 71.865 3.435 ;
      RECT 71.595 3.032 71.79 3.373 ;
      RECT 71.59 3.14 71.805 3.365 ;
      RECT 71.585 3.19 71.865 3.355 ;
      RECT 71.575 3.267 71.865 3.34 ;
      RECT 71.595 3.115 71.805 3.373 ;
      RECT 71.605 2.99 71.79 3.435 ;
      RECT 71.605 2.885 71.77 3.435 ;
      RECT 71.615 2.872 71.77 3.435 ;
      RECT 71.615 2.83 71.76 3.435 ;
      RECT 71.62 2.755 71.76 3.435 ;
      RECT 71.65 2.405 71.76 3.435 ;
      RECT 71.655 2.135 71.78 2.758 ;
      RECT 71.625 2.71 71.78 2.758 ;
      RECT 71.64 2.512 71.76 3.435 ;
      RECT 71.63 2.622 71.78 2.758 ;
      RECT 71.655 2.135 71.795 2.615 ;
      RECT 71.655 2.135 71.815 2.49 ;
      RECT 71.62 2.135 71.88 2.395 ;
      RECT 71.09 2.44 71.37 2.72 ;
      RECT 71.075 2.44 71.37 2.7 ;
      RECT 69.13 3.305 69.39 3.565 ;
      RECT 70.915 3.16 71.175 3.42 ;
      RECT 70.895 3.18 71.175 3.395 ;
      RECT 70.852 3.18 70.895 3.394 ;
      RECT 70.766 3.181 70.852 3.391 ;
      RECT 70.68 3.182 70.766 3.387 ;
      RECT 70.605 3.184 70.68 3.384 ;
      RECT 70.582 3.185 70.605 3.382 ;
      RECT 70.496 3.186 70.582 3.38 ;
      RECT 70.41 3.187 70.496 3.377 ;
      RECT 70.386 3.188 70.41 3.375 ;
      RECT 70.3 3.19 70.386 3.372 ;
      RECT 70.215 3.192 70.3 3.373 ;
      RECT 70.158 3.193 70.215 3.379 ;
      RECT 70.072 3.195 70.158 3.389 ;
      RECT 69.986 3.198 70.072 3.402 ;
      RECT 69.9 3.2 69.986 3.414 ;
      RECT 69.886 3.201 69.9 3.421 ;
      RECT 69.8 3.202 69.886 3.429 ;
      RECT 69.76 3.204 69.8 3.438 ;
      RECT 69.751 3.205 69.76 3.441 ;
      RECT 69.665 3.213 69.751 3.447 ;
      RECT 69.645 3.222 69.665 3.455 ;
      RECT 69.56 3.237 69.645 3.463 ;
      RECT 69.5 3.26 69.56 3.474 ;
      RECT 69.49 3.272 69.5 3.479 ;
      RECT 69.45 3.282 69.49 3.483 ;
      RECT 69.395 3.299 69.45 3.491 ;
      RECT 69.39 3.309 69.395 3.495 ;
      RECT 70.456 2.44 70.515 2.837 ;
      RECT 70.37 2.44 70.575 2.828 ;
      RECT 70.365 2.47 70.575 2.823 ;
      RECT 70.331 2.47 70.575 2.821 ;
      RECT 70.245 2.47 70.575 2.815 ;
      RECT 70.2 2.47 70.595 2.793 ;
      RECT 70.2 2.47 70.615 2.748 ;
      RECT 70.16 2.47 70.615 2.738 ;
      RECT 70.37 2.44 70.65 2.72 ;
      RECT 70.105 2.44 70.365 2.7 ;
      RECT 69.29 1.92 69.55 2.18 ;
      RECT 69.37 1.88 69.65 2.16 ;
      RECT 63.735 6.22 64.055 6.545 ;
      RECT 63.765 5.695 63.935 6.545 ;
      RECT 63.765 5.695 63.94 6.045 ;
      RECT 63.765 5.695 64.74 5.87 ;
      RECT 64.565 1.965 64.74 5.87 ;
      RECT 64.51 1.965 64.86 2.315 ;
      RECT 64.535 6.655 64.86 6.98 ;
      RECT 63.42 6.745 64.86 6.915 ;
      RECT 63.42 2.395 63.58 6.915 ;
      RECT 63.735 2.365 64.055 2.685 ;
      RECT 63.42 2.395 64.055 2.565 ;
      RECT 52.145 3 52.425 3.28 ;
      RECT 52.115 3 52.425 3.265 ;
      RECT 52.11 3 52.425 3.263 ;
      RECT 52.105 1.33 52.275 3.257 ;
      RECT 52.1 2.967 52.37 3.25 ;
      RECT 52.095 3 52.425 3.243 ;
      RECT 52.065 2.97 52.37 3.23 ;
      RECT 52.065 2.997 52.39 3.23 ;
      RECT 52.065 2.987 52.385 3.23 ;
      RECT 52.065 2.972 52.38 3.23 ;
      RECT 52.105 2.962 52.37 3.257 ;
      RECT 52.105 2.957 52.36 3.257 ;
      RECT 52.105 2.956 52.345 3.257 ;
      RECT 62.075 1.34 62.425 1.69 ;
      RECT 62.07 1.34 62.425 1.595 ;
      RECT 52.105 1.33 62.315 1.5 ;
      RECT 61.75 2.85 62.12 3.22 ;
      RECT 61.835 2.235 62.005 3.22 ;
      RECT 57.855 2.455 58.09 2.715 ;
      RECT 61 2.235 61.165 2.495 ;
      RECT 60.905 2.225 60.92 2.495 ;
      RECT 61 2.235 62.005 2.415 ;
      RECT 59.505 1.795 59.545 1.935 ;
      RECT 60.92 2.23 61 2.495 ;
      RECT 60.865 2.225 60.905 2.461 ;
      RECT 60.851 2.225 60.865 2.461 ;
      RECT 60.765 2.23 60.851 2.463 ;
      RECT 60.72 2.237 60.765 2.465 ;
      RECT 60.69 2.237 60.72 2.467 ;
      RECT 60.665 2.232 60.69 2.469 ;
      RECT 60.635 2.228 60.665 2.478 ;
      RECT 60.625 2.225 60.635 2.49 ;
      RECT 60.62 2.225 60.625 2.498 ;
      RECT 60.615 2.225 60.62 2.503 ;
      RECT 60.605 2.224 60.615 2.513 ;
      RECT 60.6 2.223 60.605 2.523 ;
      RECT 60.585 2.222 60.6 2.528 ;
      RECT 60.557 2.219 60.585 2.555 ;
      RECT 60.471 2.211 60.557 2.555 ;
      RECT 60.385 2.2 60.471 2.555 ;
      RECT 60.345 2.185 60.385 2.555 ;
      RECT 60.305 2.159 60.345 2.555 ;
      RECT 60.3 2.141 60.305 2.367 ;
      RECT 60.29 2.137 60.3 2.357 ;
      RECT 60.275 2.127 60.29 2.344 ;
      RECT 60.255 2.111 60.275 2.329 ;
      RECT 60.24 2.096 60.255 2.314 ;
      RECT 60.23 2.085 60.24 2.304 ;
      RECT 60.205 2.069 60.23 2.293 ;
      RECT 60.2 2.056 60.205 2.283 ;
      RECT 60.195 2.052 60.2 2.278 ;
      RECT 60.14 2.038 60.195 2.256 ;
      RECT 60.101 2.019 60.14 2.22 ;
      RECT 60.015 1.993 60.101 2.173 ;
      RECT 60.011 1.975 60.015 2.139 ;
      RECT 59.925 1.956 60.011 2.117 ;
      RECT 59.92 1.938 59.925 2.095 ;
      RECT 59.915 1.936 59.92 2.093 ;
      RECT 59.905 1.935 59.915 2.088 ;
      RECT 59.845 1.922 59.905 2.074 ;
      RECT 59.8 1.9 59.845 2.053 ;
      RECT 59.74 1.877 59.8 2.032 ;
      RECT 59.676 1.852 59.74 2.007 ;
      RECT 59.59 1.822 59.676 1.976 ;
      RECT 59.575 1.802 59.59 1.955 ;
      RECT 59.545 1.797 59.575 1.946 ;
      RECT 59.492 1.795 59.505 1.935 ;
      RECT 59.406 1.795 59.492 1.937 ;
      RECT 59.32 1.795 59.406 1.939 ;
      RECT 59.3 1.795 59.32 1.943 ;
      RECT 59.255 1.797 59.3 1.954 ;
      RECT 59.215 1.807 59.255 1.97 ;
      RECT 59.211 1.816 59.215 1.978 ;
      RECT 59.125 1.836 59.211 1.994 ;
      RECT 59.115 1.855 59.125 2.012 ;
      RECT 59.11 1.857 59.115 2.015 ;
      RECT 59.1 1.861 59.11 2.018 ;
      RECT 59.08 1.866 59.1 2.028 ;
      RECT 59.05 1.876 59.08 2.048 ;
      RECT 59.045 1.883 59.05 2.062 ;
      RECT 59.035 1.887 59.045 2.069 ;
      RECT 59.02 1.895 59.035 2.08 ;
      RECT 59.01 1.905 59.02 2.091 ;
      RECT 59 1.912 59.01 2.099 ;
      RECT 58.975 1.925 59 2.114 ;
      RECT 58.911 1.961 58.975 2.153 ;
      RECT 58.825 2.024 58.911 2.217 ;
      RECT 58.79 2.075 58.825 2.27 ;
      RECT 58.785 2.092 58.79 2.287 ;
      RECT 58.77 2.101 58.785 2.294 ;
      RECT 58.75 2.116 58.77 2.308 ;
      RECT 58.745 2.127 58.75 2.318 ;
      RECT 58.725 2.14 58.745 2.328 ;
      RECT 58.72 2.15 58.725 2.338 ;
      RECT 58.705 2.155 58.72 2.347 ;
      RECT 58.695 2.165 58.705 2.358 ;
      RECT 58.665 2.182 58.695 2.375 ;
      RECT 58.655 2.2 58.665 2.393 ;
      RECT 58.64 2.211 58.655 2.404 ;
      RECT 58.6 2.235 58.64 2.42 ;
      RECT 58.565 2.269 58.6 2.437 ;
      RECT 58.535 2.292 58.565 2.449 ;
      RECT 58.52 2.302 58.535 2.458 ;
      RECT 58.48 2.312 58.52 2.469 ;
      RECT 58.46 2.323 58.48 2.481 ;
      RECT 58.455 2.327 58.46 2.488 ;
      RECT 58.44 2.331 58.455 2.493 ;
      RECT 58.43 2.336 58.44 2.498 ;
      RECT 58.425 2.339 58.43 2.501 ;
      RECT 58.395 2.345 58.425 2.508 ;
      RECT 58.36 2.355 58.395 2.522 ;
      RECT 58.3 2.37 58.36 2.542 ;
      RECT 58.245 2.39 58.3 2.566 ;
      RECT 58.216 2.405 58.245 2.584 ;
      RECT 58.13 2.425 58.216 2.609 ;
      RECT 58.125 2.44 58.13 2.629 ;
      RECT 58.115 2.443 58.125 2.63 ;
      RECT 58.09 2.45 58.115 2.715 ;
      RECT 60.785 2.943 61.065 3.28 ;
      RECT 60.785 2.953 61.07 3.238 ;
      RECT 60.785 2.962 61.075 3.135 ;
      RECT 60.785 2.977 61.08 3.003 ;
      RECT 60.785 2.805 61.045 3.28 ;
      RECT 51.085 6.655 51.435 7.005 ;
      RECT 59.91 6.61 60.26 6.96 ;
      RECT 51.085 6.685 60.26 6.885 ;
      RECT 58.505 3.685 58.515 3.875 ;
      RECT 56.765 3.56 57.045 3.84 ;
      RECT 59.81 2.5 59.815 2.985 ;
      RECT 59.705 2.5 59.765 2.76 ;
      RECT 60.03 3.47 60.035 3.545 ;
      RECT 60.02 3.337 60.03 3.58 ;
      RECT 60.01 3.172 60.02 3.601 ;
      RECT 60.005 3.042 60.01 3.617 ;
      RECT 59.995 2.932 60.005 3.633 ;
      RECT 59.99 2.831 59.995 3.65 ;
      RECT 59.985 2.813 59.99 3.66 ;
      RECT 59.98 2.795 59.985 3.67 ;
      RECT 59.97 2.77 59.98 3.685 ;
      RECT 59.965 2.75 59.97 3.7 ;
      RECT 59.945 2.5 59.965 3.725 ;
      RECT 59.93 2.5 59.945 3.758 ;
      RECT 59.9 2.5 59.93 3.78 ;
      RECT 59.88 2.5 59.9 3.794 ;
      RECT 59.86 2.5 59.88 3.31 ;
      RECT 59.875 3.377 59.88 3.799 ;
      RECT 59.87 3.407 59.875 3.801 ;
      RECT 59.865 3.42 59.87 3.804 ;
      RECT 59.86 3.43 59.865 3.808 ;
      RECT 59.855 2.5 59.86 3.228 ;
      RECT 59.855 3.44 59.86 3.81 ;
      RECT 59.85 2.5 59.855 3.205 ;
      RECT 59.84 3.462 59.855 3.81 ;
      RECT 59.835 2.5 59.85 3.15 ;
      RECT 59.83 3.487 59.84 3.81 ;
      RECT 59.83 2.5 59.835 3.095 ;
      RECT 59.82 2.5 59.83 3.043 ;
      RECT 59.825 3.5 59.83 3.811 ;
      RECT 59.82 3.512 59.825 3.812 ;
      RECT 59.815 2.5 59.82 3.003 ;
      RECT 59.815 3.525 59.82 3.813 ;
      RECT 59.8 3.54 59.815 3.814 ;
      RECT 59.805 2.5 59.81 2.965 ;
      RECT 59.8 2.5 59.805 2.93 ;
      RECT 59.795 2.5 59.8 2.905 ;
      RECT 59.79 3.567 59.8 3.816 ;
      RECT 59.785 2.5 59.795 2.863 ;
      RECT 59.785 3.585 59.79 3.817 ;
      RECT 59.78 2.5 59.785 2.823 ;
      RECT 59.78 3.592 59.785 3.818 ;
      RECT 59.775 2.5 59.78 2.795 ;
      RECT 59.77 3.61 59.78 3.819 ;
      RECT 59.765 2.5 59.775 2.775 ;
      RECT 59.76 3.63 59.77 3.821 ;
      RECT 59.75 3.647 59.76 3.822 ;
      RECT 59.715 3.67 59.75 3.825 ;
      RECT 59.66 3.688 59.715 3.831 ;
      RECT 59.574 3.696 59.66 3.84 ;
      RECT 59.488 3.707 59.574 3.851 ;
      RECT 59.402 3.717 59.488 3.862 ;
      RECT 59.316 3.727 59.402 3.874 ;
      RECT 59.23 3.737 59.316 3.885 ;
      RECT 59.21 3.743 59.23 3.891 ;
      RECT 59.13 3.745 59.21 3.895 ;
      RECT 59.125 3.744 59.13 3.9 ;
      RECT 59.117 3.743 59.125 3.9 ;
      RECT 59.031 3.739 59.117 3.898 ;
      RECT 58.945 3.731 59.031 3.895 ;
      RECT 58.859 3.722 58.945 3.891 ;
      RECT 58.773 3.714 58.859 3.888 ;
      RECT 58.687 3.706 58.773 3.884 ;
      RECT 58.601 3.697 58.687 3.881 ;
      RECT 58.515 3.689 58.601 3.877 ;
      RECT 58.46 3.682 58.505 3.875 ;
      RECT 58.375 3.675 58.46 3.873 ;
      RECT 58.301 3.667 58.375 3.869 ;
      RECT 58.215 3.659 58.301 3.866 ;
      RECT 58.212 3.655 58.215 3.864 ;
      RECT 58.126 3.651 58.212 3.863 ;
      RECT 58.04 3.643 58.126 3.86 ;
      RECT 57.955 3.638 58.04 3.857 ;
      RECT 57.869 3.635 57.955 3.854 ;
      RECT 57.783 3.633 57.869 3.851 ;
      RECT 57.697 3.63 57.783 3.848 ;
      RECT 57.611 3.627 57.697 3.845 ;
      RECT 57.525 3.624 57.611 3.842 ;
      RECT 57.449 3.622 57.525 3.839 ;
      RECT 57.363 3.619 57.449 3.836 ;
      RECT 57.277 3.616 57.363 3.834 ;
      RECT 57.191 3.614 57.277 3.831 ;
      RECT 57.105 3.611 57.191 3.828 ;
      RECT 57.045 3.602 57.105 3.826 ;
      RECT 59.555 3.22 59.63 3.48 ;
      RECT 59.535 3.2 59.54 3.48 ;
      RECT 58.855 2.985 58.96 3.28 ;
      RECT 53.3 2.96 53.37 3.22 ;
      RECT 59.195 2.835 59.2 3.206 ;
      RECT 59.185 2.89 59.19 3.206 ;
      RECT 59.49 2.06 59.55 2.32 ;
      RECT 59.545 3.215 59.555 3.48 ;
      RECT 59.54 3.205 59.545 3.48 ;
      RECT 59.46 3.152 59.535 3.48 ;
      RECT 59.485 2.06 59.49 2.34 ;
      RECT 59.475 2.06 59.485 2.36 ;
      RECT 59.46 2.06 59.475 2.39 ;
      RECT 59.445 2.06 59.46 2.433 ;
      RECT 59.44 3.095 59.46 3.48 ;
      RECT 59.43 2.06 59.445 2.47 ;
      RECT 59.425 3.075 59.44 3.48 ;
      RECT 59.425 2.06 59.43 2.493 ;
      RECT 59.415 2.06 59.425 2.518 ;
      RECT 59.385 3.042 59.425 3.48 ;
      RECT 59.39 2.06 59.415 2.568 ;
      RECT 59.385 2.06 59.39 2.623 ;
      RECT 59.38 2.06 59.385 2.665 ;
      RECT 59.37 3.005 59.385 3.48 ;
      RECT 59.375 2.06 59.38 2.708 ;
      RECT 59.37 2.06 59.375 2.773 ;
      RECT 59.365 2.06 59.37 2.795 ;
      RECT 59.365 2.993 59.37 3.345 ;
      RECT 59.36 2.06 59.365 2.863 ;
      RECT 59.36 2.985 59.365 3.328 ;
      RECT 59.355 2.06 59.36 2.908 ;
      RECT 59.35 2.967 59.36 3.305 ;
      RECT 59.35 2.06 59.355 2.945 ;
      RECT 59.34 2.06 59.35 3.285 ;
      RECT 59.335 2.06 59.34 3.268 ;
      RECT 59.33 2.06 59.335 3.253 ;
      RECT 59.325 2.06 59.33 3.238 ;
      RECT 59.305 2.06 59.325 3.228 ;
      RECT 59.3 2.06 59.305 3.218 ;
      RECT 59.29 2.06 59.3 3.214 ;
      RECT 59.285 2.337 59.29 3.213 ;
      RECT 59.28 2.36 59.285 3.212 ;
      RECT 59.275 2.39 59.28 3.211 ;
      RECT 59.27 2.417 59.275 3.21 ;
      RECT 59.265 2.445 59.27 3.21 ;
      RECT 59.26 2.472 59.265 3.21 ;
      RECT 59.255 2.492 59.26 3.21 ;
      RECT 59.25 2.52 59.255 3.21 ;
      RECT 59.24 2.562 59.25 3.21 ;
      RECT 59.23 2.607 59.24 3.209 ;
      RECT 59.225 2.66 59.23 3.208 ;
      RECT 59.22 2.692 59.225 3.207 ;
      RECT 59.215 2.712 59.22 3.206 ;
      RECT 59.21 2.75 59.215 3.206 ;
      RECT 59.205 2.772 59.21 3.206 ;
      RECT 59.2 2.797 59.205 3.206 ;
      RECT 59.19 2.862 59.195 3.206 ;
      RECT 59.175 2.922 59.185 3.206 ;
      RECT 59.16 2.932 59.175 3.206 ;
      RECT 59.14 2.942 59.16 3.206 ;
      RECT 59.11 2.947 59.14 3.203 ;
      RECT 59.05 2.957 59.11 3.2 ;
      RECT 59.03 2.966 59.05 3.205 ;
      RECT 59.005 2.972 59.03 3.218 ;
      RECT 58.985 2.977 59.005 3.233 ;
      RECT 58.96 2.982 58.985 3.28 ;
      RECT 58.831 2.984 58.855 3.28 ;
      RECT 58.745 2.979 58.831 3.28 ;
      RECT 58.705 2.976 58.745 3.28 ;
      RECT 58.655 2.978 58.705 3.26 ;
      RECT 58.625 2.982 58.655 3.26 ;
      RECT 58.546 2.992 58.625 3.26 ;
      RECT 58.46 3.007 58.546 3.261 ;
      RECT 58.41 3.017 58.46 3.262 ;
      RECT 58.402 3.02 58.41 3.262 ;
      RECT 58.316 3.022 58.402 3.263 ;
      RECT 58.23 3.026 58.316 3.263 ;
      RECT 58.144 3.03 58.23 3.264 ;
      RECT 58.058 3.033 58.144 3.265 ;
      RECT 57.972 3.037 58.058 3.265 ;
      RECT 57.886 3.041 57.972 3.266 ;
      RECT 57.8 3.044 57.886 3.267 ;
      RECT 57.714 3.048 57.8 3.267 ;
      RECT 57.628 3.052 57.714 3.268 ;
      RECT 57.542 3.056 57.628 3.269 ;
      RECT 57.456 3.059 57.542 3.269 ;
      RECT 57.37 3.063 57.456 3.27 ;
      RECT 57.34 3.065 57.37 3.27 ;
      RECT 57.254 3.068 57.34 3.271 ;
      RECT 57.168 3.072 57.254 3.272 ;
      RECT 57.082 3.076 57.168 3.273 ;
      RECT 56.996 3.079 57.082 3.273 ;
      RECT 56.91 3.083 56.996 3.274 ;
      RECT 56.875 3.088 56.91 3.275 ;
      RECT 56.82 3.098 56.875 3.282 ;
      RECT 56.795 3.11 56.82 3.292 ;
      RECT 56.76 3.123 56.795 3.3 ;
      RECT 56.72 3.14 56.76 3.323 ;
      RECT 56.7 3.153 56.72 3.35 ;
      RECT 56.67 3.165 56.7 3.378 ;
      RECT 56.665 3.173 56.67 3.398 ;
      RECT 56.66 3.176 56.665 3.408 ;
      RECT 56.61 3.188 56.66 3.442 ;
      RECT 56.6 3.203 56.61 3.475 ;
      RECT 56.59 3.209 56.6 3.488 ;
      RECT 56.58 3.216 56.59 3.5 ;
      RECT 56.555 3.229 56.58 3.518 ;
      RECT 56.54 3.244 56.555 3.54 ;
      RECT 56.53 3.252 56.54 3.556 ;
      RECT 56.515 3.261 56.53 3.571 ;
      RECT 56.505 3.271 56.515 3.585 ;
      RECT 56.486 3.284 56.505 3.602 ;
      RECT 56.4 3.329 56.486 3.667 ;
      RECT 56.385 3.374 56.4 3.725 ;
      RECT 56.38 3.383 56.385 3.738 ;
      RECT 56.37 3.39 56.38 3.743 ;
      RECT 56.365 3.395 56.37 3.747 ;
      RECT 56.345 3.405 56.365 3.754 ;
      RECT 56.32 3.425 56.345 3.768 ;
      RECT 56.285 3.45 56.32 3.788 ;
      RECT 56.27 3.473 56.285 3.803 ;
      RECT 56.26 3.483 56.27 3.808 ;
      RECT 56.25 3.491 56.26 3.815 ;
      RECT 56.24 3.5 56.25 3.821 ;
      RECT 56.22 3.512 56.24 3.823 ;
      RECT 56.21 3.525 56.22 3.825 ;
      RECT 56.185 3.54 56.21 3.828 ;
      RECT 56.165 3.557 56.185 3.832 ;
      RECT 56.125 3.585 56.165 3.838 ;
      RECT 56.06 3.632 56.125 3.847 ;
      RECT 56.045 3.665 56.06 3.855 ;
      RECT 56.04 3.672 56.045 3.857 ;
      RECT 55.99 3.697 56.04 3.862 ;
      RECT 55.975 3.721 55.99 3.869 ;
      RECT 55.925 3.726 55.975 3.87 ;
      RECT 55.839 3.73 55.925 3.87 ;
      RECT 55.753 3.73 55.839 3.87 ;
      RECT 55.667 3.73 55.753 3.871 ;
      RECT 55.581 3.73 55.667 3.871 ;
      RECT 55.495 3.73 55.581 3.871 ;
      RECT 55.429 3.73 55.495 3.871 ;
      RECT 55.343 3.73 55.429 3.872 ;
      RECT 55.257 3.73 55.343 3.872 ;
      RECT 55.171 3.731 55.257 3.873 ;
      RECT 55.085 3.731 55.171 3.873 ;
      RECT 54.999 3.731 55.085 3.873 ;
      RECT 54.913 3.731 54.999 3.874 ;
      RECT 54.827 3.731 54.913 3.874 ;
      RECT 54.741 3.732 54.827 3.875 ;
      RECT 54.655 3.732 54.741 3.875 ;
      RECT 54.635 3.732 54.655 3.875 ;
      RECT 54.549 3.732 54.635 3.875 ;
      RECT 54.463 3.732 54.549 3.875 ;
      RECT 54.377 3.733 54.463 3.875 ;
      RECT 54.291 3.733 54.377 3.875 ;
      RECT 54.205 3.733 54.291 3.875 ;
      RECT 54.119 3.734 54.205 3.875 ;
      RECT 54.033 3.734 54.119 3.875 ;
      RECT 53.947 3.734 54.033 3.875 ;
      RECT 53.861 3.734 53.947 3.875 ;
      RECT 53.775 3.735 53.861 3.875 ;
      RECT 53.725 3.732 53.775 3.875 ;
      RECT 53.715 3.73 53.725 3.874 ;
      RECT 53.711 3.73 53.715 3.873 ;
      RECT 53.625 3.725 53.711 3.868 ;
      RECT 53.603 3.718 53.625 3.862 ;
      RECT 53.517 3.709 53.603 3.856 ;
      RECT 53.431 3.696 53.517 3.847 ;
      RECT 53.345 3.682 53.431 3.837 ;
      RECT 53.3 3.672 53.345 3.83 ;
      RECT 53.28 2.96 53.3 3.238 ;
      RECT 53.28 3.665 53.3 3.826 ;
      RECT 53.25 2.96 53.28 3.26 ;
      RECT 53.24 3.632 53.28 3.823 ;
      RECT 53.235 2.96 53.25 3.28 ;
      RECT 53.235 3.597 53.24 3.821 ;
      RECT 53.23 2.96 53.235 3.405 ;
      RECT 53.23 3.557 53.235 3.821 ;
      RECT 53.22 2.96 53.23 3.821 ;
      RECT 53.145 2.96 53.22 3.815 ;
      RECT 53.115 2.96 53.145 3.805 ;
      RECT 53.11 2.96 53.115 3.797 ;
      RECT 53.105 3.002 53.11 3.79 ;
      RECT 53.095 3.071 53.105 3.781 ;
      RECT 53.09 3.141 53.095 3.733 ;
      RECT 53.085 3.205 53.09 3.63 ;
      RECT 53.08 3.24 53.085 3.585 ;
      RECT 53.078 3.277 53.08 3.477 ;
      RECT 53.075 3.285 53.078 3.47 ;
      RECT 53.07 3.35 53.075 3.413 ;
      RECT 57.145 2.44 57.425 2.72 ;
      RECT 57.135 2.44 57.425 2.583 ;
      RECT 57.09 2.305 57.35 2.565 ;
      RECT 57.09 2.42 57.405 2.565 ;
      RECT 57.09 2.39 57.4 2.565 ;
      RECT 57.09 2.377 57.39 2.565 ;
      RECT 57.09 2.367 57.385 2.565 ;
      RECT 53.065 2.35 53.325 2.61 ;
      RECT 56.835 1.9 57.095 2.16 ;
      RECT 56.825 1.925 57.095 2.12 ;
      RECT 56.82 1.925 56.825 2.119 ;
      RECT 56.75 1.92 56.82 2.111 ;
      RECT 56.665 1.907 56.75 2.094 ;
      RECT 56.661 1.899 56.665 2.084 ;
      RECT 56.575 1.892 56.661 2.074 ;
      RECT 56.566 1.884 56.575 2.064 ;
      RECT 56.48 1.877 56.566 2.052 ;
      RECT 56.46 1.868 56.48 2.038 ;
      RECT 56.405 1.863 56.46 2.03 ;
      RECT 56.395 1.857 56.405 2.024 ;
      RECT 56.375 1.855 56.395 2.02 ;
      RECT 56.367 1.854 56.375 2.016 ;
      RECT 56.281 1.846 56.367 2.005 ;
      RECT 56.195 1.832 56.281 1.985 ;
      RECT 56.135 1.82 56.195 1.97 ;
      RECT 56.125 1.815 56.135 1.965 ;
      RECT 56.075 1.815 56.125 1.967 ;
      RECT 56.028 1.817 56.075 1.971 ;
      RECT 55.942 1.824 56.028 1.976 ;
      RECT 55.856 1.832 55.942 1.982 ;
      RECT 55.77 1.841 55.856 1.988 ;
      RECT 55.711 1.847 55.77 1.993 ;
      RECT 55.625 1.852 55.711 1.999 ;
      RECT 55.55 1.857 55.625 2.005 ;
      RECT 55.511 1.859 55.55 2.01 ;
      RECT 55.425 1.856 55.511 2.015 ;
      RECT 55.34 1.854 55.425 2.022 ;
      RECT 55.308 1.853 55.34 2.025 ;
      RECT 55.222 1.852 55.308 2.026 ;
      RECT 55.136 1.851 55.222 2.027 ;
      RECT 55.05 1.85 55.136 2.027 ;
      RECT 54.964 1.849 55.05 2.028 ;
      RECT 54.878 1.848 54.964 2.029 ;
      RECT 54.792 1.847 54.878 2.03 ;
      RECT 54.706 1.846 54.792 2.03 ;
      RECT 54.62 1.845 54.706 2.031 ;
      RECT 54.57 1.845 54.62 2.032 ;
      RECT 54.556 1.846 54.57 2.032 ;
      RECT 54.47 1.853 54.556 2.033 ;
      RECT 54.396 1.864 54.47 2.034 ;
      RECT 54.31 1.873 54.396 2.035 ;
      RECT 54.275 1.88 54.31 2.05 ;
      RECT 54.25 1.883 54.275 2.08 ;
      RECT 54.225 1.892 54.25 2.109 ;
      RECT 54.215 1.903 54.225 2.129 ;
      RECT 54.205 1.911 54.215 2.143 ;
      RECT 54.2 1.917 54.205 2.153 ;
      RECT 54.175 1.934 54.2 2.17 ;
      RECT 54.16 1.956 54.175 2.198 ;
      RECT 54.13 1.982 54.16 2.228 ;
      RECT 54.11 2.011 54.13 2.258 ;
      RECT 54.105 2.026 54.11 2.275 ;
      RECT 54.085 2.041 54.105 2.29 ;
      RECT 54.075 2.059 54.085 2.308 ;
      RECT 54.065 2.07 54.075 2.323 ;
      RECT 54.015 2.102 54.065 2.349 ;
      RECT 54.01 2.132 54.015 2.369 ;
      RECT 54 2.145 54.01 2.375 ;
      RECT 53.991 2.155 54 2.383 ;
      RECT 53.98 2.166 53.991 2.391 ;
      RECT 53.975 2.176 53.98 2.397 ;
      RECT 53.96 2.197 53.975 2.404 ;
      RECT 53.945 2.227 53.96 2.412 ;
      RECT 53.91 2.257 53.945 2.418 ;
      RECT 53.885 2.275 53.91 2.425 ;
      RECT 53.835 2.283 53.885 2.434 ;
      RECT 53.81 2.288 53.835 2.443 ;
      RECT 53.755 2.294 53.81 2.453 ;
      RECT 53.75 2.299 53.755 2.461 ;
      RECT 53.736 2.302 53.75 2.463 ;
      RECT 53.65 2.314 53.736 2.475 ;
      RECT 53.64 2.326 53.65 2.488 ;
      RECT 53.555 2.339 53.64 2.5 ;
      RECT 53.511 2.356 53.555 2.514 ;
      RECT 53.425 2.373 53.511 2.53 ;
      RECT 53.395 2.387 53.425 2.544 ;
      RECT 53.385 2.392 53.395 2.549 ;
      RECT 53.325 2.395 53.385 2.558 ;
      RECT 56.215 2.665 56.475 2.925 ;
      RECT 56.215 2.665 56.495 2.778 ;
      RECT 56.215 2.665 56.52 2.745 ;
      RECT 56.215 2.665 56.525 2.725 ;
      RECT 56.265 2.44 56.545 2.72 ;
      RECT 55.82 3.175 56.08 3.435 ;
      RECT 55.81 3.032 56.005 3.373 ;
      RECT 55.805 3.14 56.02 3.365 ;
      RECT 55.8 3.19 56.08 3.355 ;
      RECT 55.79 3.267 56.08 3.34 ;
      RECT 55.81 3.115 56.02 3.373 ;
      RECT 55.82 2.99 56.005 3.435 ;
      RECT 55.82 2.885 55.985 3.435 ;
      RECT 55.83 2.872 55.985 3.435 ;
      RECT 55.83 2.83 55.975 3.435 ;
      RECT 55.835 2.755 55.975 3.435 ;
      RECT 55.865 2.405 55.975 3.435 ;
      RECT 55.87 2.135 55.995 2.758 ;
      RECT 55.84 2.71 55.995 2.758 ;
      RECT 55.855 2.512 55.975 3.435 ;
      RECT 55.845 2.622 55.995 2.758 ;
      RECT 55.87 2.135 56.01 2.615 ;
      RECT 55.87 2.135 56.03 2.49 ;
      RECT 55.835 2.135 56.095 2.395 ;
      RECT 55.305 2.44 55.585 2.72 ;
      RECT 55.29 2.44 55.585 2.7 ;
      RECT 53.345 3.305 53.605 3.565 ;
      RECT 55.13 3.16 55.39 3.42 ;
      RECT 55.11 3.18 55.39 3.395 ;
      RECT 55.067 3.18 55.11 3.394 ;
      RECT 54.981 3.181 55.067 3.391 ;
      RECT 54.895 3.182 54.981 3.387 ;
      RECT 54.82 3.184 54.895 3.384 ;
      RECT 54.797 3.185 54.82 3.382 ;
      RECT 54.711 3.186 54.797 3.38 ;
      RECT 54.625 3.187 54.711 3.377 ;
      RECT 54.601 3.188 54.625 3.375 ;
      RECT 54.515 3.19 54.601 3.372 ;
      RECT 54.43 3.192 54.515 3.373 ;
      RECT 54.373 3.193 54.43 3.379 ;
      RECT 54.287 3.195 54.373 3.389 ;
      RECT 54.201 3.198 54.287 3.402 ;
      RECT 54.115 3.2 54.201 3.414 ;
      RECT 54.101 3.201 54.115 3.421 ;
      RECT 54.015 3.202 54.101 3.429 ;
      RECT 53.975 3.204 54.015 3.438 ;
      RECT 53.966 3.205 53.975 3.441 ;
      RECT 53.88 3.213 53.966 3.447 ;
      RECT 53.86 3.222 53.88 3.455 ;
      RECT 53.775 3.237 53.86 3.463 ;
      RECT 53.715 3.26 53.775 3.474 ;
      RECT 53.705 3.272 53.715 3.479 ;
      RECT 53.665 3.282 53.705 3.483 ;
      RECT 53.61 3.299 53.665 3.491 ;
      RECT 53.605 3.309 53.61 3.495 ;
      RECT 54.671 2.44 54.73 2.837 ;
      RECT 54.585 2.44 54.79 2.828 ;
      RECT 54.58 2.47 54.79 2.823 ;
      RECT 54.546 2.47 54.79 2.821 ;
      RECT 54.46 2.47 54.79 2.815 ;
      RECT 54.415 2.47 54.81 2.793 ;
      RECT 54.415 2.47 54.83 2.748 ;
      RECT 54.375 2.47 54.83 2.738 ;
      RECT 54.585 2.44 54.865 2.72 ;
      RECT 54.32 2.44 54.58 2.7 ;
      RECT 53.505 1.92 53.765 2.18 ;
      RECT 53.585 1.88 53.865 2.16 ;
      RECT 47.95 6.22 48.27 6.545 ;
      RECT 47.98 5.695 48.15 6.545 ;
      RECT 47.98 5.695 48.155 6.045 ;
      RECT 47.98 5.695 48.955 5.87 ;
      RECT 48.78 1.965 48.955 5.87 ;
      RECT 48.725 1.965 49.075 2.315 ;
      RECT 48.75 6.655 49.075 6.98 ;
      RECT 47.635 6.745 49.075 6.915 ;
      RECT 47.635 2.395 47.795 6.915 ;
      RECT 47.95 2.365 48.27 2.685 ;
      RECT 47.635 2.395 48.27 2.565 ;
      RECT 36.36 3 36.64 3.28 ;
      RECT 36.33 3 36.64 3.265 ;
      RECT 36.325 3 36.64 3.263 ;
      RECT 36.32 1.33 36.49 3.257 ;
      RECT 36.315 2.967 36.585 3.25 ;
      RECT 36.31 3 36.64 3.243 ;
      RECT 36.28 2.97 36.585 3.23 ;
      RECT 36.28 2.997 36.605 3.23 ;
      RECT 36.28 2.987 36.6 3.23 ;
      RECT 36.28 2.972 36.595 3.23 ;
      RECT 36.32 2.962 36.585 3.257 ;
      RECT 36.32 2.957 36.575 3.257 ;
      RECT 36.32 2.956 36.56 3.257 ;
      RECT 46.29 1.34 46.64 1.69 ;
      RECT 46.285 1.34 46.64 1.595 ;
      RECT 36.32 1.33 46.53 1.5 ;
      RECT 45.965 2.85 46.335 3.22 ;
      RECT 46.05 2.235 46.22 3.22 ;
      RECT 42.07 2.455 42.305 2.715 ;
      RECT 45.215 2.235 45.38 2.495 ;
      RECT 45.12 2.225 45.135 2.495 ;
      RECT 45.215 2.235 46.22 2.415 ;
      RECT 43.72 1.795 43.76 1.935 ;
      RECT 45.135 2.23 45.215 2.495 ;
      RECT 45.08 2.225 45.12 2.461 ;
      RECT 45.066 2.225 45.08 2.461 ;
      RECT 44.98 2.23 45.066 2.463 ;
      RECT 44.935 2.237 44.98 2.465 ;
      RECT 44.905 2.237 44.935 2.467 ;
      RECT 44.88 2.232 44.905 2.469 ;
      RECT 44.85 2.228 44.88 2.478 ;
      RECT 44.84 2.225 44.85 2.49 ;
      RECT 44.835 2.225 44.84 2.498 ;
      RECT 44.83 2.225 44.835 2.503 ;
      RECT 44.82 2.224 44.83 2.513 ;
      RECT 44.815 2.223 44.82 2.523 ;
      RECT 44.8 2.222 44.815 2.528 ;
      RECT 44.772 2.219 44.8 2.555 ;
      RECT 44.686 2.211 44.772 2.555 ;
      RECT 44.6 2.2 44.686 2.555 ;
      RECT 44.56 2.185 44.6 2.555 ;
      RECT 44.52 2.159 44.56 2.555 ;
      RECT 44.515 2.141 44.52 2.367 ;
      RECT 44.505 2.137 44.515 2.357 ;
      RECT 44.49 2.127 44.505 2.344 ;
      RECT 44.47 2.111 44.49 2.329 ;
      RECT 44.455 2.096 44.47 2.314 ;
      RECT 44.445 2.085 44.455 2.304 ;
      RECT 44.42 2.069 44.445 2.293 ;
      RECT 44.415 2.056 44.42 2.283 ;
      RECT 44.41 2.052 44.415 2.278 ;
      RECT 44.355 2.038 44.41 2.256 ;
      RECT 44.316 2.019 44.355 2.22 ;
      RECT 44.23 1.993 44.316 2.173 ;
      RECT 44.226 1.975 44.23 2.139 ;
      RECT 44.14 1.956 44.226 2.117 ;
      RECT 44.135 1.938 44.14 2.095 ;
      RECT 44.13 1.936 44.135 2.093 ;
      RECT 44.12 1.935 44.13 2.088 ;
      RECT 44.06 1.922 44.12 2.074 ;
      RECT 44.015 1.9 44.06 2.053 ;
      RECT 43.955 1.877 44.015 2.032 ;
      RECT 43.891 1.852 43.955 2.007 ;
      RECT 43.805 1.822 43.891 1.976 ;
      RECT 43.79 1.802 43.805 1.955 ;
      RECT 43.76 1.797 43.79 1.946 ;
      RECT 43.707 1.795 43.72 1.935 ;
      RECT 43.621 1.795 43.707 1.937 ;
      RECT 43.535 1.795 43.621 1.939 ;
      RECT 43.515 1.795 43.535 1.943 ;
      RECT 43.47 1.797 43.515 1.954 ;
      RECT 43.43 1.807 43.47 1.97 ;
      RECT 43.426 1.816 43.43 1.978 ;
      RECT 43.34 1.836 43.426 1.994 ;
      RECT 43.33 1.855 43.34 2.012 ;
      RECT 43.325 1.857 43.33 2.015 ;
      RECT 43.315 1.861 43.325 2.018 ;
      RECT 43.295 1.866 43.315 2.028 ;
      RECT 43.265 1.876 43.295 2.048 ;
      RECT 43.26 1.883 43.265 2.062 ;
      RECT 43.25 1.887 43.26 2.069 ;
      RECT 43.235 1.895 43.25 2.08 ;
      RECT 43.225 1.905 43.235 2.091 ;
      RECT 43.215 1.912 43.225 2.099 ;
      RECT 43.19 1.925 43.215 2.114 ;
      RECT 43.126 1.961 43.19 2.153 ;
      RECT 43.04 2.024 43.126 2.217 ;
      RECT 43.005 2.075 43.04 2.27 ;
      RECT 43 2.092 43.005 2.287 ;
      RECT 42.985 2.101 43 2.294 ;
      RECT 42.965 2.116 42.985 2.308 ;
      RECT 42.96 2.127 42.965 2.318 ;
      RECT 42.94 2.14 42.96 2.328 ;
      RECT 42.935 2.15 42.94 2.338 ;
      RECT 42.92 2.155 42.935 2.347 ;
      RECT 42.91 2.165 42.92 2.358 ;
      RECT 42.88 2.182 42.91 2.375 ;
      RECT 42.87 2.2 42.88 2.393 ;
      RECT 42.855 2.211 42.87 2.404 ;
      RECT 42.815 2.235 42.855 2.42 ;
      RECT 42.78 2.269 42.815 2.437 ;
      RECT 42.75 2.292 42.78 2.449 ;
      RECT 42.735 2.302 42.75 2.458 ;
      RECT 42.695 2.312 42.735 2.469 ;
      RECT 42.675 2.323 42.695 2.481 ;
      RECT 42.67 2.327 42.675 2.488 ;
      RECT 42.655 2.331 42.67 2.493 ;
      RECT 42.645 2.336 42.655 2.498 ;
      RECT 42.64 2.339 42.645 2.501 ;
      RECT 42.61 2.345 42.64 2.508 ;
      RECT 42.575 2.355 42.61 2.522 ;
      RECT 42.515 2.37 42.575 2.542 ;
      RECT 42.46 2.39 42.515 2.566 ;
      RECT 42.431 2.405 42.46 2.584 ;
      RECT 42.345 2.425 42.431 2.609 ;
      RECT 42.34 2.44 42.345 2.629 ;
      RECT 42.33 2.443 42.34 2.63 ;
      RECT 42.305 2.45 42.33 2.715 ;
      RECT 45 2.943 45.28 3.28 ;
      RECT 45 2.953 45.285 3.238 ;
      RECT 45 2.962 45.29 3.135 ;
      RECT 45 2.977 45.295 3.003 ;
      RECT 45 2.805 45.26 3.28 ;
      RECT 35.355 6.66 35.705 7.01 ;
      RECT 44.18 6.615 44.53 6.965 ;
      RECT 35.355 6.69 44.53 6.89 ;
      RECT 42.72 3.685 42.73 3.875 ;
      RECT 40.98 3.56 41.26 3.84 ;
      RECT 44.025 2.5 44.03 2.985 ;
      RECT 43.92 2.5 43.98 2.76 ;
      RECT 44.245 3.47 44.25 3.545 ;
      RECT 44.235 3.337 44.245 3.58 ;
      RECT 44.225 3.172 44.235 3.601 ;
      RECT 44.22 3.042 44.225 3.617 ;
      RECT 44.21 2.932 44.22 3.633 ;
      RECT 44.205 2.831 44.21 3.65 ;
      RECT 44.2 2.813 44.205 3.66 ;
      RECT 44.195 2.795 44.2 3.67 ;
      RECT 44.185 2.77 44.195 3.685 ;
      RECT 44.18 2.75 44.185 3.7 ;
      RECT 44.16 2.5 44.18 3.725 ;
      RECT 44.145 2.5 44.16 3.758 ;
      RECT 44.115 2.5 44.145 3.78 ;
      RECT 44.095 2.5 44.115 3.794 ;
      RECT 44.075 2.5 44.095 3.31 ;
      RECT 44.09 3.377 44.095 3.799 ;
      RECT 44.085 3.407 44.09 3.801 ;
      RECT 44.08 3.42 44.085 3.804 ;
      RECT 44.075 3.43 44.08 3.808 ;
      RECT 44.07 2.5 44.075 3.228 ;
      RECT 44.07 3.44 44.075 3.81 ;
      RECT 44.065 2.5 44.07 3.205 ;
      RECT 44.055 3.462 44.07 3.81 ;
      RECT 44.05 2.5 44.065 3.15 ;
      RECT 44.045 3.487 44.055 3.81 ;
      RECT 44.045 2.5 44.05 3.095 ;
      RECT 44.035 2.5 44.045 3.043 ;
      RECT 44.04 3.5 44.045 3.811 ;
      RECT 44.035 3.512 44.04 3.812 ;
      RECT 44.03 2.5 44.035 3.003 ;
      RECT 44.03 3.525 44.035 3.813 ;
      RECT 44.015 3.54 44.03 3.814 ;
      RECT 44.02 2.5 44.025 2.965 ;
      RECT 44.015 2.5 44.02 2.93 ;
      RECT 44.01 2.5 44.015 2.905 ;
      RECT 44.005 3.567 44.015 3.816 ;
      RECT 44 2.5 44.01 2.863 ;
      RECT 44 3.585 44.005 3.817 ;
      RECT 43.995 2.5 44 2.823 ;
      RECT 43.995 3.592 44 3.818 ;
      RECT 43.99 2.5 43.995 2.795 ;
      RECT 43.985 3.61 43.995 3.819 ;
      RECT 43.98 2.5 43.99 2.775 ;
      RECT 43.975 3.63 43.985 3.821 ;
      RECT 43.965 3.647 43.975 3.822 ;
      RECT 43.93 3.67 43.965 3.825 ;
      RECT 43.875 3.688 43.93 3.831 ;
      RECT 43.789 3.696 43.875 3.84 ;
      RECT 43.703 3.707 43.789 3.851 ;
      RECT 43.617 3.717 43.703 3.862 ;
      RECT 43.531 3.727 43.617 3.874 ;
      RECT 43.445 3.737 43.531 3.885 ;
      RECT 43.425 3.743 43.445 3.891 ;
      RECT 43.345 3.745 43.425 3.895 ;
      RECT 43.34 3.744 43.345 3.9 ;
      RECT 43.332 3.743 43.34 3.9 ;
      RECT 43.246 3.739 43.332 3.898 ;
      RECT 43.16 3.731 43.246 3.895 ;
      RECT 43.074 3.722 43.16 3.891 ;
      RECT 42.988 3.714 43.074 3.888 ;
      RECT 42.902 3.706 42.988 3.884 ;
      RECT 42.816 3.697 42.902 3.881 ;
      RECT 42.73 3.689 42.816 3.877 ;
      RECT 42.675 3.682 42.72 3.875 ;
      RECT 42.59 3.675 42.675 3.873 ;
      RECT 42.516 3.667 42.59 3.869 ;
      RECT 42.43 3.659 42.516 3.866 ;
      RECT 42.427 3.655 42.43 3.864 ;
      RECT 42.341 3.651 42.427 3.863 ;
      RECT 42.255 3.643 42.341 3.86 ;
      RECT 42.17 3.638 42.255 3.857 ;
      RECT 42.084 3.635 42.17 3.854 ;
      RECT 41.998 3.633 42.084 3.851 ;
      RECT 41.912 3.63 41.998 3.848 ;
      RECT 41.826 3.627 41.912 3.845 ;
      RECT 41.74 3.624 41.826 3.842 ;
      RECT 41.664 3.622 41.74 3.839 ;
      RECT 41.578 3.619 41.664 3.836 ;
      RECT 41.492 3.616 41.578 3.834 ;
      RECT 41.406 3.614 41.492 3.831 ;
      RECT 41.32 3.611 41.406 3.828 ;
      RECT 41.26 3.602 41.32 3.826 ;
      RECT 43.77 3.22 43.845 3.48 ;
      RECT 43.75 3.2 43.755 3.48 ;
      RECT 43.07 2.985 43.175 3.28 ;
      RECT 37.515 2.96 37.585 3.22 ;
      RECT 43.41 2.835 43.415 3.206 ;
      RECT 43.4 2.89 43.405 3.206 ;
      RECT 43.705 2.06 43.765 2.32 ;
      RECT 43.76 3.215 43.77 3.48 ;
      RECT 43.755 3.205 43.76 3.48 ;
      RECT 43.675 3.152 43.75 3.48 ;
      RECT 43.7 2.06 43.705 2.34 ;
      RECT 43.69 2.06 43.7 2.36 ;
      RECT 43.675 2.06 43.69 2.39 ;
      RECT 43.66 2.06 43.675 2.433 ;
      RECT 43.655 3.095 43.675 3.48 ;
      RECT 43.645 2.06 43.66 2.47 ;
      RECT 43.64 3.075 43.655 3.48 ;
      RECT 43.64 2.06 43.645 2.493 ;
      RECT 43.63 2.06 43.64 2.518 ;
      RECT 43.6 3.042 43.64 3.48 ;
      RECT 43.605 2.06 43.63 2.568 ;
      RECT 43.6 2.06 43.605 2.623 ;
      RECT 43.595 2.06 43.6 2.665 ;
      RECT 43.585 3.005 43.6 3.48 ;
      RECT 43.59 2.06 43.595 2.708 ;
      RECT 43.585 2.06 43.59 2.773 ;
      RECT 43.58 2.06 43.585 2.795 ;
      RECT 43.58 2.993 43.585 3.345 ;
      RECT 43.575 2.06 43.58 2.863 ;
      RECT 43.575 2.985 43.58 3.328 ;
      RECT 43.57 2.06 43.575 2.908 ;
      RECT 43.565 2.967 43.575 3.305 ;
      RECT 43.565 2.06 43.57 2.945 ;
      RECT 43.555 2.06 43.565 3.285 ;
      RECT 43.55 2.06 43.555 3.268 ;
      RECT 43.545 2.06 43.55 3.253 ;
      RECT 43.54 2.06 43.545 3.238 ;
      RECT 43.52 2.06 43.54 3.228 ;
      RECT 43.515 2.06 43.52 3.218 ;
      RECT 43.505 2.06 43.515 3.214 ;
      RECT 43.5 2.337 43.505 3.213 ;
      RECT 43.495 2.36 43.5 3.212 ;
      RECT 43.49 2.39 43.495 3.211 ;
      RECT 43.485 2.417 43.49 3.21 ;
      RECT 43.48 2.445 43.485 3.21 ;
      RECT 43.475 2.472 43.48 3.21 ;
      RECT 43.47 2.492 43.475 3.21 ;
      RECT 43.465 2.52 43.47 3.21 ;
      RECT 43.455 2.562 43.465 3.21 ;
      RECT 43.445 2.607 43.455 3.209 ;
      RECT 43.44 2.66 43.445 3.208 ;
      RECT 43.435 2.692 43.44 3.207 ;
      RECT 43.43 2.712 43.435 3.206 ;
      RECT 43.425 2.75 43.43 3.206 ;
      RECT 43.42 2.772 43.425 3.206 ;
      RECT 43.415 2.797 43.42 3.206 ;
      RECT 43.405 2.862 43.41 3.206 ;
      RECT 43.39 2.922 43.4 3.206 ;
      RECT 43.375 2.932 43.39 3.206 ;
      RECT 43.355 2.942 43.375 3.206 ;
      RECT 43.325 2.947 43.355 3.203 ;
      RECT 43.265 2.957 43.325 3.2 ;
      RECT 43.245 2.966 43.265 3.205 ;
      RECT 43.22 2.972 43.245 3.218 ;
      RECT 43.2 2.977 43.22 3.233 ;
      RECT 43.175 2.982 43.2 3.28 ;
      RECT 43.046 2.984 43.07 3.28 ;
      RECT 42.96 2.979 43.046 3.28 ;
      RECT 42.92 2.976 42.96 3.28 ;
      RECT 42.87 2.978 42.92 3.26 ;
      RECT 42.84 2.982 42.87 3.26 ;
      RECT 42.761 2.992 42.84 3.26 ;
      RECT 42.675 3.007 42.761 3.261 ;
      RECT 42.625 3.017 42.675 3.262 ;
      RECT 42.617 3.02 42.625 3.262 ;
      RECT 42.531 3.022 42.617 3.263 ;
      RECT 42.445 3.026 42.531 3.263 ;
      RECT 42.359 3.03 42.445 3.264 ;
      RECT 42.273 3.033 42.359 3.265 ;
      RECT 42.187 3.037 42.273 3.265 ;
      RECT 42.101 3.041 42.187 3.266 ;
      RECT 42.015 3.044 42.101 3.267 ;
      RECT 41.929 3.048 42.015 3.267 ;
      RECT 41.843 3.052 41.929 3.268 ;
      RECT 41.757 3.056 41.843 3.269 ;
      RECT 41.671 3.059 41.757 3.269 ;
      RECT 41.585 3.063 41.671 3.27 ;
      RECT 41.555 3.065 41.585 3.27 ;
      RECT 41.469 3.068 41.555 3.271 ;
      RECT 41.383 3.072 41.469 3.272 ;
      RECT 41.297 3.076 41.383 3.273 ;
      RECT 41.211 3.079 41.297 3.273 ;
      RECT 41.125 3.083 41.211 3.274 ;
      RECT 41.09 3.088 41.125 3.275 ;
      RECT 41.035 3.098 41.09 3.282 ;
      RECT 41.01 3.11 41.035 3.292 ;
      RECT 40.975 3.123 41.01 3.3 ;
      RECT 40.935 3.14 40.975 3.323 ;
      RECT 40.915 3.153 40.935 3.35 ;
      RECT 40.885 3.165 40.915 3.378 ;
      RECT 40.88 3.173 40.885 3.398 ;
      RECT 40.875 3.176 40.88 3.408 ;
      RECT 40.825 3.188 40.875 3.442 ;
      RECT 40.815 3.203 40.825 3.475 ;
      RECT 40.805 3.209 40.815 3.488 ;
      RECT 40.795 3.216 40.805 3.5 ;
      RECT 40.77 3.229 40.795 3.518 ;
      RECT 40.755 3.244 40.77 3.54 ;
      RECT 40.745 3.252 40.755 3.556 ;
      RECT 40.73 3.261 40.745 3.571 ;
      RECT 40.72 3.271 40.73 3.585 ;
      RECT 40.701 3.284 40.72 3.602 ;
      RECT 40.615 3.329 40.701 3.667 ;
      RECT 40.6 3.374 40.615 3.725 ;
      RECT 40.595 3.383 40.6 3.738 ;
      RECT 40.585 3.39 40.595 3.743 ;
      RECT 40.58 3.395 40.585 3.747 ;
      RECT 40.56 3.405 40.58 3.754 ;
      RECT 40.535 3.425 40.56 3.768 ;
      RECT 40.5 3.45 40.535 3.788 ;
      RECT 40.485 3.473 40.5 3.803 ;
      RECT 40.475 3.483 40.485 3.808 ;
      RECT 40.465 3.491 40.475 3.815 ;
      RECT 40.455 3.5 40.465 3.821 ;
      RECT 40.435 3.512 40.455 3.823 ;
      RECT 40.425 3.525 40.435 3.825 ;
      RECT 40.4 3.54 40.425 3.828 ;
      RECT 40.38 3.557 40.4 3.832 ;
      RECT 40.34 3.585 40.38 3.838 ;
      RECT 40.275 3.632 40.34 3.847 ;
      RECT 40.26 3.665 40.275 3.855 ;
      RECT 40.255 3.672 40.26 3.857 ;
      RECT 40.205 3.697 40.255 3.862 ;
      RECT 40.19 3.721 40.205 3.869 ;
      RECT 40.14 3.726 40.19 3.87 ;
      RECT 40.054 3.73 40.14 3.87 ;
      RECT 39.968 3.73 40.054 3.87 ;
      RECT 39.882 3.73 39.968 3.871 ;
      RECT 39.796 3.73 39.882 3.871 ;
      RECT 39.71 3.73 39.796 3.871 ;
      RECT 39.644 3.73 39.71 3.871 ;
      RECT 39.558 3.73 39.644 3.872 ;
      RECT 39.472 3.73 39.558 3.872 ;
      RECT 39.386 3.731 39.472 3.873 ;
      RECT 39.3 3.731 39.386 3.873 ;
      RECT 39.214 3.731 39.3 3.873 ;
      RECT 39.128 3.731 39.214 3.874 ;
      RECT 39.042 3.731 39.128 3.874 ;
      RECT 38.956 3.732 39.042 3.875 ;
      RECT 38.87 3.732 38.956 3.875 ;
      RECT 38.85 3.732 38.87 3.875 ;
      RECT 38.764 3.732 38.85 3.875 ;
      RECT 38.678 3.732 38.764 3.875 ;
      RECT 38.592 3.733 38.678 3.875 ;
      RECT 38.506 3.733 38.592 3.875 ;
      RECT 38.42 3.733 38.506 3.875 ;
      RECT 38.334 3.734 38.42 3.875 ;
      RECT 38.248 3.734 38.334 3.875 ;
      RECT 38.162 3.734 38.248 3.875 ;
      RECT 38.076 3.734 38.162 3.875 ;
      RECT 37.99 3.735 38.076 3.875 ;
      RECT 37.94 3.732 37.99 3.875 ;
      RECT 37.93 3.73 37.94 3.874 ;
      RECT 37.926 3.73 37.93 3.873 ;
      RECT 37.84 3.725 37.926 3.868 ;
      RECT 37.818 3.718 37.84 3.862 ;
      RECT 37.732 3.709 37.818 3.856 ;
      RECT 37.646 3.696 37.732 3.847 ;
      RECT 37.56 3.682 37.646 3.837 ;
      RECT 37.515 3.672 37.56 3.83 ;
      RECT 37.495 2.96 37.515 3.238 ;
      RECT 37.495 3.665 37.515 3.826 ;
      RECT 37.465 2.96 37.495 3.26 ;
      RECT 37.455 3.632 37.495 3.823 ;
      RECT 37.45 2.96 37.465 3.28 ;
      RECT 37.45 3.597 37.455 3.821 ;
      RECT 37.445 2.96 37.45 3.405 ;
      RECT 37.445 3.557 37.45 3.821 ;
      RECT 37.435 2.96 37.445 3.821 ;
      RECT 37.36 2.96 37.435 3.815 ;
      RECT 37.33 2.96 37.36 3.805 ;
      RECT 37.325 2.96 37.33 3.797 ;
      RECT 37.32 3.002 37.325 3.79 ;
      RECT 37.31 3.071 37.32 3.781 ;
      RECT 37.305 3.141 37.31 3.733 ;
      RECT 37.3 3.205 37.305 3.63 ;
      RECT 37.295 3.24 37.3 3.585 ;
      RECT 37.293 3.277 37.295 3.477 ;
      RECT 37.29 3.285 37.293 3.47 ;
      RECT 37.285 3.35 37.29 3.413 ;
      RECT 41.36 2.44 41.64 2.72 ;
      RECT 41.35 2.44 41.64 2.583 ;
      RECT 41.305 2.305 41.565 2.565 ;
      RECT 41.305 2.42 41.62 2.565 ;
      RECT 41.305 2.39 41.615 2.565 ;
      RECT 41.305 2.377 41.605 2.565 ;
      RECT 41.305 2.367 41.6 2.565 ;
      RECT 37.28 2.35 37.54 2.61 ;
      RECT 41.05 1.9 41.31 2.16 ;
      RECT 41.04 1.925 41.31 2.12 ;
      RECT 41.035 1.925 41.04 2.119 ;
      RECT 40.965 1.92 41.035 2.111 ;
      RECT 40.88 1.907 40.965 2.094 ;
      RECT 40.876 1.899 40.88 2.084 ;
      RECT 40.79 1.892 40.876 2.074 ;
      RECT 40.781 1.884 40.79 2.064 ;
      RECT 40.695 1.877 40.781 2.052 ;
      RECT 40.675 1.868 40.695 2.038 ;
      RECT 40.62 1.863 40.675 2.03 ;
      RECT 40.61 1.857 40.62 2.024 ;
      RECT 40.59 1.855 40.61 2.02 ;
      RECT 40.582 1.854 40.59 2.016 ;
      RECT 40.496 1.846 40.582 2.005 ;
      RECT 40.41 1.832 40.496 1.985 ;
      RECT 40.35 1.82 40.41 1.97 ;
      RECT 40.34 1.815 40.35 1.965 ;
      RECT 40.29 1.815 40.34 1.967 ;
      RECT 40.243 1.817 40.29 1.971 ;
      RECT 40.157 1.824 40.243 1.976 ;
      RECT 40.071 1.832 40.157 1.982 ;
      RECT 39.985 1.841 40.071 1.988 ;
      RECT 39.926 1.847 39.985 1.993 ;
      RECT 39.84 1.852 39.926 1.999 ;
      RECT 39.765 1.857 39.84 2.005 ;
      RECT 39.726 1.859 39.765 2.01 ;
      RECT 39.64 1.856 39.726 2.015 ;
      RECT 39.555 1.854 39.64 2.022 ;
      RECT 39.523 1.853 39.555 2.025 ;
      RECT 39.437 1.852 39.523 2.026 ;
      RECT 39.351 1.851 39.437 2.027 ;
      RECT 39.265 1.85 39.351 2.027 ;
      RECT 39.179 1.849 39.265 2.028 ;
      RECT 39.093 1.848 39.179 2.029 ;
      RECT 39.007 1.847 39.093 2.03 ;
      RECT 38.921 1.846 39.007 2.03 ;
      RECT 38.835 1.845 38.921 2.031 ;
      RECT 38.785 1.845 38.835 2.032 ;
      RECT 38.771 1.846 38.785 2.032 ;
      RECT 38.685 1.853 38.771 2.033 ;
      RECT 38.611 1.864 38.685 2.034 ;
      RECT 38.525 1.873 38.611 2.035 ;
      RECT 38.49 1.88 38.525 2.05 ;
      RECT 38.465 1.883 38.49 2.08 ;
      RECT 38.44 1.892 38.465 2.109 ;
      RECT 38.43 1.903 38.44 2.129 ;
      RECT 38.42 1.911 38.43 2.143 ;
      RECT 38.415 1.917 38.42 2.153 ;
      RECT 38.39 1.934 38.415 2.17 ;
      RECT 38.375 1.956 38.39 2.198 ;
      RECT 38.345 1.982 38.375 2.228 ;
      RECT 38.325 2.011 38.345 2.258 ;
      RECT 38.32 2.026 38.325 2.275 ;
      RECT 38.3 2.041 38.32 2.29 ;
      RECT 38.29 2.059 38.3 2.308 ;
      RECT 38.28 2.07 38.29 2.323 ;
      RECT 38.23 2.102 38.28 2.349 ;
      RECT 38.225 2.132 38.23 2.369 ;
      RECT 38.215 2.145 38.225 2.375 ;
      RECT 38.206 2.155 38.215 2.383 ;
      RECT 38.195 2.166 38.206 2.391 ;
      RECT 38.19 2.176 38.195 2.397 ;
      RECT 38.175 2.197 38.19 2.404 ;
      RECT 38.16 2.227 38.175 2.412 ;
      RECT 38.125 2.257 38.16 2.418 ;
      RECT 38.1 2.275 38.125 2.425 ;
      RECT 38.05 2.283 38.1 2.434 ;
      RECT 38.025 2.288 38.05 2.443 ;
      RECT 37.97 2.294 38.025 2.453 ;
      RECT 37.965 2.299 37.97 2.461 ;
      RECT 37.951 2.302 37.965 2.463 ;
      RECT 37.865 2.314 37.951 2.475 ;
      RECT 37.855 2.326 37.865 2.488 ;
      RECT 37.77 2.339 37.855 2.5 ;
      RECT 37.726 2.356 37.77 2.514 ;
      RECT 37.64 2.373 37.726 2.53 ;
      RECT 37.61 2.387 37.64 2.544 ;
      RECT 37.6 2.392 37.61 2.549 ;
      RECT 37.54 2.395 37.6 2.558 ;
      RECT 40.43 2.665 40.69 2.925 ;
      RECT 40.43 2.665 40.71 2.778 ;
      RECT 40.43 2.665 40.735 2.745 ;
      RECT 40.43 2.665 40.74 2.725 ;
      RECT 40.48 2.44 40.76 2.72 ;
      RECT 40.035 3.175 40.295 3.435 ;
      RECT 40.025 3.032 40.22 3.373 ;
      RECT 40.02 3.14 40.235 3.365 ;
      RECT 40.015 3.19 40.295 3.355 ;
      RECT 40.005 3.267 40.295 3.34 ;
      RECT 40.025 3.115 40.235 3.373 ;
      RECT 40.035 2.99 40.22 3.435 ;
      RECT 40.035 2.885 40.2 3.435 ;
      RECT 40.045 2.872 40.2 3.435 ;
      RECT 40.045 2.83 40.19 3.435 ;
      RECT 40.05 2.755 40.19 3.435 ;
      RECT 40.08 2.405 40.19 3.435 ;
      RECT 40.085 2.135 40.21 2.758 ;
      RECT 40.055 2.71 40.21 2.758 ;
      RECT 40.07 2.512 40.19 3.435 ;
      RECT 40.06 2.622 40.21 2.758 ;
      RECT 40.085 2.135 40.225 2.615 ;
      RECT 40.085 2.135 40.245 2.49 ;
      RECT 40.05 2.135 40.31 2.395 ;
      RECT 39.52 2.44 39.8 2.72 ;
      RECT 39.505 2.44 39.8 2.7 ;
      RECT 37.56 3.305 37.82 3.565 ;
      RECT 39.345 3.16 39.605 3.42 ;
      RECT 39.325 3.18 39.605 3.395 ;
      RECT 39.282 3.18 39.325 3.394 ;
      RECT 39.196 3.181 39.282 3.391 ;
      RECT 39.11 3.182 39.196 3.387 ;
      RECT 39.035 3.184 39.11 3.384 ;
      RECT 39.012 3.185 39.035 3.382 ;
      RECT 38.926 3.186 39.012 3.38 ;
      RECT 38.84 3.187 38.926 3.377 ;
      RECT 38.816 3.188 38.84 3.375 ;
      RECT 38.73 3.19 38.816 3.372 ;
      RECT 38.645 3.192 38.73 3.373 ;
      RECT 38.588 3.193 38.645 3.379 ;
      RECT 38.502 3.195 38.588 3.389 ;
      RECT 38.416 3.198 38.502 3.402 ;
      RECT 38.33 3.2 38.416 3.414 ;
      RECT 38.316 3.201 38.33 3.421 ;
      RECT 38.23 3.202 38.316 3.429 ;
      RECT 38.19 3.204 38.23 3.438 ;
      RECT 38.181 3.205 38.19 3.441 ;
      RECT 38.095 3.213 38.181 3.447 ;
      RECT 38.075 3.222 38.095 3.455 ;
      RECT 37.99 3.237 38.075 3.463 ;
      RECT 37.93 3.26 37.99 3.474 ;
      RECT 37.92 3.272 37.93 3.479 ;
      RECT 37.88 3.282 37.92 3.483 ;
      RECT 37.825 3.299 37.88 3.491 ;
      RECT 37.82 3.309 37.825 3.495 ;
      RECT 38.886 2.44 38.945 2.837 ;
      RECT 38.8 2.44 39.005 2.828 ;
      RECT 38.795 2.47 39.005 2.823 ;
      RECT 38.761 2.47 39.005 2.821 ;
      RECT 38.675 2.47 39.005 2.815 ;
      RECT 38.63 2.47 39.025 2.793 ;
      RECT 38.63 2.47 39.045 2.748 ;
      RECT 38.59 2.47 39.045 2.738 ;
      RECT 38.8 2.44 39.08 2.72 ;
      RECT 38.535 2.44 38.795 2.7 ;
      RECT 37.72 1.92 37.98 2.18 ;
      RECT 37.8 1.88 38.08 2.16 ;
      RECT 32.175 6.22 32.495 6.545 ;
      RECT 32.205 5.695 32.375 6.545 ;
      RECT 32.205 5.695 32.38 6.045 ;
      RECT 32.205 5.695 33.18 5.87 ;
      RECT 33.005 1.965 33.18 5.87 ;
      RECT 32.95 1.965 33.3 2.315 ;
      RECT 32.975 6.655 33.3 6.98 ;
      RECT 31.86 6.745 33.3 6.915 ;
      RECT 31.86 2.395 32.02 6.915 ;
      RECT 32.175 2.365 32.495 2.685 ;
      RECT 31.86 2.395 32.495 2.565 ;
      RECT 20.585 3 20.865 3.28 ;
      RECT 20.555 3 20.865 3.265 ;
      RECT 20.55 3 20.865 3.263 ;
      RECT 20.545 1.33 20.715 3.257 ;
      RECT 20.54 2.967 20.81 3.25 ;
      RECT 20.535 3 20.865 3.243 ;
      RECT 20.505 2.97 20.81 3.23 ;
      RECT 20.505 2.997 20.83 3.23 ;
      RECT 20.505 2.987 20.825 3.23 ;
      RECT 20.505 2.972 20.82 3.23 ;
      RECT 20.545 2.962 20.81 3.257 ;
      RECT 20.545 2.957 20.8 3.257 ;
      RECT 20.545 2.956 20.785 3.257 ;
      RECT 30.515 1.34 30.865 1.69 ;
      RECT 30.51 1.34 30.865 1.595 ;
      RECT 20.545 1.33 30.755 1.5 ;
      RECT 30.19 2.85 30.56 3.22 ;
      RECT 30.275 2.235 30.445 3.22 ;
      RECT 26.295 2.455 26.53 2.715 ;
      RECT 29.44 2.235 29.605 2.495 ;
      RECT 29.345 2.225 29.36 2.495 ;
      RECT 29.44 2.235 30.445 2.415 ;
      RECT 27.945 1.795 27.985 1.935 ;
      RECT 29.36 2.23 29.44 2.495 ;
      RECT 29.305 2.225 29.345 2.461 ;
      RECT 29.291 2.225 29.305 2.461 ;
      RECT 29.205 2.23 29.291 2.463 ;
      RECT 29.16 2.237 29.205 2.465 ;
      RECT 29.13 2.237 29.16 2.467 ;
      RECT 29.105 2.232 29.13 2.469 ;
      RECT 29.075 2.228 29.105 2.478 ;
      RECT 29.065 2.225 29.075 2.49 ;
      RECT 29.06 2.225 29.065 2.498 ;
      RECT 29.055 2.225 29.06 2.503 ;
      RECT 29.045 2.224 29.055 2.513 ;
      RECT 29.04 2.223 29.045 2.523 ;
      RECT 29.025 2.222 29.04 2.528 ;
      RECT 28.997 2.219 29.025 2.555 ;
      RECT 28.911 2.211 28.997 2.555 ;
      RECT 28.825 2.2 28.911 2.555 ;
      RECT 28.785 2.185 28.825 2.555 ;
      RECT 28.745 2.159 28.785 2.555 ;
      RECT 28.74 2.141 28.745 2.367 ;
      RECT 28.73 2.137 28.74 2.357 ;
      RECT 28.715 2.127 28.73 2.344 ;
      RECT 28.695 2.111 28.715 2.329 ;
      RECT 28.68 2.096 28.695 2.314 ;
      RECT 28.67 2.085 28.68 2.304 ;
      RECT 28.645 2.069 28.67 2.293 ;
      RECT 28.64 2.056 28.645 2.283 ;
      RECT 28.635 2.052 28.64 2.278 ;
      RECT 28.58 2.038 28.635 2.256 ;
      RECT 28.541 2.019 28.58 2.22 ;
      RECT 28.455 1.993 28.541 2.173 ;
      RECT 28.451 1.975 28.455 2.139 ;
      RECT 28.365 1.956 28.451 2.117 ;
      RECT 28.36 1.938 28.365 2.095 ;
      RECT 28.355 1.936 28.36 2.093 ;
      RECT 28.345 1.935 28.355 2.088 ;
      RECT 28.285 1.922 28.345 2.074 ;
      RECT 28.24 1.9 28.285 2.053 ;
      RECT 28.18 1.877 28.24 2.032 ;
      RECT 28.116 1.852 28.18 2.007 ;
      RECT 28.03 1.822 28.116 1.976 ;
      RECT 28.015 1.802 28.03 1.955 ;
      RECT 27.985 1.797 28.015 1.946 ;
      RECT 27.932 1.795 27.945 1.935 ;
      RECT 27.846 1.795 27.932 1.937 ;
      RECT 27.76 1.795 27.846 1.939 ;
      RECT 27.74 1.795 27.76 1.943 ;
      RECT 27.695 1.797 27.74 1.954 ;
      RECT 27.655 1.807 27.695 1.97 ;
      RECT 27.651 1.816 27.655 1.978 ;
      RECT 27.565 1.836 27.651 1.994 ;
      RECT 27.555 1.855 27.565 2.012 ;
      RECT 27.55 1.857 27.555 2.015 ;
      RECT 27.54 1.861 27.55 2.018 ;
      RECT 27.52 1.866 27.54 2.028 ;
      RECT 27.49 1.876 27.52 2.048 ;
      RECT 27.485 1.883 27.49 2.062 ;
      RECT 27.475 1.887 27.485 2.069 ;
      RECT 27.46 1.895 27.475 2.08 ;
      RECT 27.45 1.905 27.46 2.091 ;
      RECT 27.44 1.912 27.45 2.099 ;
      RECT 27.415 1.925 27.44 2.114 ;
      RECT 27.351 1.961 27.415 2.153 ;
      RECT 27.265 2.024 27.351 2.217 ;
      RECT 27.23 2.075 27.265 2.27 ;
      RECT 27.225 2.092 27.23 2.287 ;
      RECT 27.21 2.101 27.225 2.294 ;
      RECT 27.19 2.116 27.21 2.308 ;
      RECT 27.185 2.127 27.19 2.318 ;
      RECT 27.165 2.14 27.185 2.328 ;
      RECT 27.16 2.15 27.165 2.338 ;
      RECT 27.145 2.155 27.16 2.347 ;
      RECT 27.135 2.165 27.145 2.358 ;
      RECT 27.105 2.182 27.135 2.375 ;
      RECT 27.095 2.2 27.105 2.393 ;
      RECT 27.08 2.211 27.095 2.404 ;
      RECT 27.04 2.235 27.08 2.42 ;
      RECT 27.005 2.269 27.04 2.437 ;
      RECT 26.975 2.292 27.005 2.449 ;
      RECT 26.96 2.302 26.975 2.458 ;
      RECT 26.92 2.312 26.96 2.469 ;
      RECT 26.9 2.323 26.92 2.481 ;
      RECT 26.895 2.327 26.9 2.488 ;
      RECT 26.88 2.331 26.895 2.493 ;
      RECT 26.87 2.336 26.88 2.498 ;
      RECT 26.865 2.339 26.87 2.501 ;
      RECT 26.835 2.345 26.865 2.508 ;
      RECT 26.8 2.355 26.835 2.522 ;
      RECT 26.74 2.37 26.8 2.542 ;
      RECT 26.685 2.39 26.74 2.566 ;
      RECT 26.656 2.405 26.685 2.584 ;
      RECT 26.57 2.425 26.656 2.609 ;
      RECT 26.565 2.44 26.57 2.629 ;
      RECT 26.555 2.443 26.565 2.63 ;
      RECT 26.53 2.45 26.555 2.715 ;
      RECT 29.225 2.943 29.505 3.28 ;
      RECT 29.225 2.953 29.51 3.238 ;
      RECT 29.225 2.962 29.515 3.135 ;
      RECT 29.225 2.977 29.52 3.003 ;
      RECT 29.225 2.805 29.485 3.28 ;
      RECT 19.575 6.655 19.925 7.005 ;
      RECT 28.4 6.61 28.75 6.96 ;
      RECT 19.575 6.685 28.75 6.885 ;
      RECT 26.945 3.685 26.955 3.875 ;
      RECT 25.205 3.56 25.485 3.84 ;
      RECT 28.25 2.5 28.255 2.985 ;
      RECT 28.145 2.5 28.205 2.76 ;
      RECT 28.47 3.47 28.475 3.545 ;
      RECT 28.46 3.337 28.47 3.58 ;
      RECT 28.45 3.172 28.46 3.601 ;
      RECT 28.445 3.042 28.45 3.617 ;
      RECT 28.435 2.932 28.445 3.633 ;
      RECT 28.43 2.831 28.435 3.65 ;
      RECT 28.425 2.813 28.43 3.66 ;
      RECT 28.42 2.795 28.425 3.67 ;
      RECT 28.41 2.77 28.42 3.685 ;
      RECT 28.405 2.75 28.41 3.7 ;
      RECT 28.385 2.5 28.405 3.725 ;
      RECT 28.37 2.5 28.385 3.758 ;
      RECT 28.34 2.5 28.37 3.78 ;
      RECT 28.32 2.5 28.34 3.794 ;
      RECT 28.3 2.5 28.32 3.31 ;
      RECT 28.315 3.377 28.32 3.799 ;
      RECT 28.31 3.407 28.315 3.801 ;
      RECT 28.305 3.42 28.31 3.804 ;
      RECT 28.3 3.43 28.305 3.808 ;
      RECT 28.295 2.5 28.3 3.228 ;
      RECT 28.295 3.44 28.3 3.81 ;
      RECT 28.29 2.5 28.295 3.205 ;
      RECT 28.28 3.462 28.295 3.81 ;
      RECT 28.275 2.5 28.29 3.15 ;
      RECT 28.27 3.487 28.28 3.81 ;
      RECT 28.27 2.5 28.275 3.095 ;
      RECT 28.26 2.5 28.27 3.043 ;
      RECT 28.265 3.5 28.27 3.811 ;
      RECT 28.26 3.512 28.265 3.812 ;
      RECT 28.255 2.5 28.26 3.003 ;
      RECT 28.255 3.525 28.26 3.813 ;
      RECT 28.24 3.54 28.255 3.814 ;
      RECT 28.245 2.5 28.25 2.965 ;
      RECT 28.24 2.5 28.245 2.93 ;
      RECT 28.235 2.5 28.24 2.905 ;
      RECT 28.23 3.567 28.24 3.816 ;
      RECT 28.225 2.5 28.235 2.863 ;
      RECT 28.225 3.585 28.23 3.817 ;
      RECT 28.22 2.5 28.225 2.823 ;
      RECT 28.22 3.592 28.225 3.818 ;
      RECT 28.215 2.5 28.22 2.795 ;
      RECT 28.21 3.61 28.22 3.819 ;
      RECT 28.205 2.5 28.215 2.775 ;
      RECT 28.2 3.63 28.21 3.821 ;
      RECT 28.19 3.647 28.2 3.822 ;
      RECT 28.155 3.67 28.19 3.825 ;
      RECT 28.1 3.688 28.155 3.831 ;
      RECT 28.014 3.696 28.1 3.84 ;
      RECT 27.928 3.707 28.014 3.851 ;
      RECT 27.842 3.717 27.928 3.862 ;
      RECT 27.756 3.727 27.842 3.874 ;
      RECT 27.67 3.737 27.756 3.885 ;
      RECT 27.65 3.743 27.67 3.891 ;
      RECT 27.57 3.745 27.65 3.895 ;
      RECT 27.565 3.744 27.57 3.9 ;
      RECT 27.557 3.743 27.565 3.9 ;
      RECT 27.471 3.739 27.557 3.898 ;
      RECT 27.385 3.731 27.471 3.895 ;
      RECT 27.299 3.722 27.385 3.891 ;
      RECT 27.213 3.714 27.299 3.888 ;
      RECT 27.127 3.706 27.213 3.884 ;
      RECT 27.041 3.697 27.127 3.881 ;
      RECT 26.955 3.689 27.041 3.877 ;
      RECT 26.9 3.682 26.945 3.875 ;
      RECT 26.815 3.675 26.9 3.873 ;
      RECT 26.741 3.667 26.815 3.869 ;
      RECT 26.655 3.659 26.741 3.866 ;
      RECT 26.652 3.655 26.655 3.864 ;
      RECT 26.566 3.651 26.652 3.863 ;
      RECT 26.48 3.643 26.566 3.86 ;
      RECT 26.395 3.638 26.48 3.857 ;
      RECT 26.309 3.635 26.395 3.854 ;
      RECT 26.223 3.633 26.309 3.851 ;
      RECT 26.137 3.63 26.223 3.848 ;
      RECT 26.051 3.627 26.137 3.845 ;
      RECT 25.965 3.624 26.051 3.842 ;
      RECT 25.889 3.622 25.965 3.839 ;
      RECT 25.803 3.619 25.889 3.836 ;
      RECT 25.717 3.616 25.803 3.834 ;
      RECT 25.631 3.614 25.717 3.831 ;
      RECT 25.545 3.611 25.631 3.828 ;
      RECT 25.485 3.602 25.545 3.826 ;
      RECT 27.995 3.22 28.07 3.48 ;
      RECT 27.975 3.2 27.98 3.48 ;
      RECT 27.295 2.985 27.4 3.28 ;
      RECT 21.74 2.96 21.81 3.22 ;
      RECT 27.635 2.835 27.64 3.206 ;
      RECT 27.625 2.89 27.63 3.206 ;
      RECT 27.93 2.06 27.99 2.32 ;
      RECT 27.985 3.215 27.995 3.48 ;
      RECT 27.98 3.205 27.985 3.48 ;
      RECT 27.9 3.152 27.975 3.48 ;
      RECT 27.925 2.06 27.93 2.34 ;
      RECT 27.915 2.06 27.925 2.36 ;
      RECT 27.9 2.06 27.915 2.39 ;
      RECT 27.885 2.06 27.9 2.433 ;
      RECT 27.88 3.095 27.9 3.48 ;
      RECT 27.87 2.06 27.885 2.47 ;
      RECT 27.865 3.075 27.88 3.48 ;
      RECT 27.865 2.06 27.87 2.493 ;
      RECT 27.855 2.06 27.865 2.518 ;
      RECT 27.825 3.042 27.865 3.48 ;
      RECT 27.83 2.06 27.855 2.568 ;
      RECT 27.825 2.06 27.83 2.623 ;
      RECT 27.82 2.06 27.825 2.665 ;
      RECT 27.81 3.005 27.825 3.48 ;
      RECT 27.815 2.06 27.82 2.708 ;
      RECT 27.81 2.06 27.815 2.773 ;
      RECT 27.805 2.06 27.81 2.795 ;
      RECT 27.805 2.993 27.81 3.345 ;
      RECT 27.8 2.06 27.805 2.863 ;
      RECT 27.8 2.985 27.805 3.328 ;
      RECT 27.795 2.06 27.8 2.908 ;
      RECT 27.79 2.967 27.8 3.305 ;
      RECT 27.79 2.06 27.795 2.945 ;
      RECT 27.78 2.06 27.79 3.285 ;
      RECT 27.775 2.06 27.78 3.268 ;
      RECT 27.77 2.06 27.775 3.253 ;
      RECT 27.765 2.06 27.77 3.238 ;
      RECT 27.745 2.06 27.765 3.228 ;
      RECT 27.74 2.06 27.745 3.218 ;
      RECT 27.73 2.06 27.74 3.214 ;
      RECT 27.725 2.337 27.73 3.213 ;
      RECT 27.72 2.36 27.725 3.212 ;
      RECT 27.715 2.39 27.72 3.211 ;
      RECT 27.71 2.417 27.715 3.21 ;
      RECT 27.705 2.445 27.71 3.21 ;
      RECT 27.7 2.472 27.705 3.21 ;
      RECT 27.695 2.492 27.7 3.21 ;
      RECT 27.69 2.52 27.695 3.21 ;
      RECT 27.68 2.562 27.69 3.21 ;
      RECT 27.67 2.607 27.68 3.209 ;
      RECT 27.665 2.66 27.67 3.208 ;
      RECT 27.66 2.692 27.665 3.207 ;
      RECT 27.655 2.712 27.66 3.206 ;
      RECT 27.65 2.75 27.655 3.206 ;
      RECT 27.645 2.772 27.65 3.206 ;
      RECT 27.64 2.797 27.645 3.206 ;
      RECT 27.63 2.862 27.635 3.206 ;
      RECT 27.615 2.922 27.625 3.206 ;
      RECT 27.6 2.932 27.615 3.206 ;
      RECT 27.58 2.942 27.6 3.206 ;
      RECT 27.55 2.947 27.58 3.203 ;
      RECT 27.49 2.957 27.55 3.2 ;
      RECT 27.47 2.966 27.49 3.205 ;
      RECT 27.445 2.972 27.47 3.218 ;
      RECT 27.425 2.977 27.445 3.233 ;
      RECT 27.4 2.982 27.425 3.28 ;
      RECT 27.271 2.984 27.295 3.28 ;
      RECT 27.185 2.979 27.271 3.28 ;
      RECT 27.145 2.976 27.185 3.28 ;
      RECT 27.095 2.978 27.145 3.26 ;
      RECT 27.065 2.982 27.095 3.26 ;
      RECT 26.986 2.992 27.065 3.26 ;
      RECT 26.9 3.007 26.986 3.261 ;
      RECT 26.85 3.017 26.9 3.262 ;
      RECT 26.842 3.02 26.85 3.262 ;
      RECT 26.756 3.022 26.842 3.263 ;
      RECT 26.67 3.026 26.756 3.263 ;
      RECT 26.584 3.03 26.67 3.264 ;
      RECT 26.498 3.033 26.584 3.265 ;
      RECT 26.412 3.037 26.498 3.265 ;
      RECT 26.326 3.041 26.412 3.266 ;
      RECT 26.24 3.044 26.326 3.267 ;
      RECT 26.154 3.048 26.24 3.267 ;
      RECT 26.068 3.052 26.154 3.268 ;
      RECT 25.982 3.056 26.068 3.269 ;
      RECT 25.896 3.059 25.982 3.269 ;
      RECT 25.81 3.063 25.896 3.27 ;
      RECT 25.78 3.065 25.81 3.27 ;
      RECT 25.694 3.068 25.78 3.271 ;
      RECT 25.608 3.072 25.694 3.272 ;
      RECT 25.522 3.076 25.608 3.273 ;
      RECT 25.436 3.079 25.522 3.273 ;
      RECT 25.35 3.083 25.436 3.274 ;
      RECT 25.315 3.088 25.35 3.275 ;
      RECT 25.26 3.098 25.315 3.282 ;
      RECT 25.235 3.11 25.26 3.292 ;
      RECT 25.2 3.123 25.235 3.3 ;
      RECT 25.16 3.14 25.2 3.323 ;
      RECT 25.14 3.153 25.16 3.35 ;
      RECT 25.11 3.165 25.14 3.378 ;
      RECT 25.105 3.173 25.11 3.398 ;
      RECT 25.1 3.176 25.105 3.408 ;
      RECT 25.05 3.188 25.1 3.442 ;
      RECT 25.04 3.203 25.05 3.475 ;
      RECT 25.03 3.209 25.04 3.488 ;
      RECT 25.02 3.216 25.03 3.5 ;
      RECT 24.995 3.229 25.02 3.518 ;
      RECT 24.98 3.244 24.995 3.54 ;
      RECT 24.97 3.252 24.98 3.556 ;
      RECT 24.955 3.261 24.97 3.571 ;
      RECT 24.945 3.271 24.955 3.585 ;
      RECT 24.926 3.284 24.945 3.602 ;
      RECT 24.84 3.329 24.926 3.667 ;
      RECT 24.825 3.374 24.84 3.725 ;
      RECT 24.82 3.383 24.825 3.738 ;
      RECT 24.81 3.39 24.82 3.743 ;
      RECT 24.805 3.395 24.81 3.747 ;
      RECT 24.785 3.405 24.805 3.754 ;
      RECT 24.76 3.425 24.785 3.768 ;
      RECT 24.725 3.45 24.76 3.788 ;
      RECT 24.71 3.473 24.725 3.803 ;
      RECT 24.7 3.483 24.71 3.808 ;
      RECT 24.69 3.491 24.7 3.815 ;
      RECT 24.68 3.5 24.69 3.821 ;
      RECT 24.66 3.512 24.68 3.823 ;
      RECT 24.65 3.525 24.66 3.825 ;
      RECT 24.625 3.54 24.65 3.828 ;
      RECT 24.605 3.557 24.625 3.832 ;
      RECT 24.565 3.585 24.605 3.838 ;
      RECT 24.5 3.632 24.565 3.847 ;
      RECT 24.485 3.665 24.5 3.855 ;
      RECT 24.48 3.672 24.485 3.857 ;
      RECT 24.43 3.697 24.48 3.862 ;
      RECT 24.415 3.721 24.43 3.869 ;
      RECT 24.365 3.726 24.415 3.87 ;
      RECT 24.279 3.73 24.365 3.87 ;
      RECT 24.193 3.73 24.279 3.87 ;
      RECT 24.107 3.73 24.193 3.871 ;
      RECT 24.021 3.73 24.107 3.871 ;
      RECT 23.935 3.73 24.021 3.871 ;
      RECT 23.869 3.73 23.935 3.871 ;
      RECT 23.783 3.73 23.869 3.872 ;
      RECT 23.697 3.73 23.783 3.872 ;
      RECT 23.611 3.731 23.697 3.873 ;
      RECT 23.525 3.731 23.611 3.873 ;
      RECT 23.439 3.731 23.525 3.873 ;
      RECT 23.353 3.731 23.439 3.874 ;
      RECT 23.267 3.731 23.353 3.874 ;
      RECT 23.181 3.732 23.267 3.875 ;
      RECT 23.095 3.732 23.181 3.875 ;
      RECT 23.075 3.732 23.095 3.875 ;
      RECT 22.989 3.732 23.075 3.875 ;
      RECT 22.903 3.732 22.989 3.875 ;
      RECT 22.817 3.733 22.903 3.875 ;
      RECT 22.731 3.733 22.817 3.875 ;
      RECT 22.645 3.733 22.731 3.875 ;
      RECT 22.559 3.734 22.645 3.875 ;
      RECT 22.473 3.734 22.559 3.875 ;
      RECT 22.387 3.734 22.473 3.875 ;
      RECT 22.301 3.734 22.387 3.875 ;
      RECT 22.215 3.735 22.301 3.875 ;
      RECT 22.165 3.732 22.215 3.875 ;
      RECT 22.155 3.73 22.165 3.874 ;
      RECT 22.151 3.73 22.155 3.873 ;
      RECT 22.065 3.725 22.151 3.868 ;
      RECT 22.043 3.718 22.065 3.862 ;
      RECT 21.957 3.709 22.043 3.856 ;
      RECT 21.871 3.696 21.957 3.847 ;
      RECT 21.785 3.682 21.871 3.837 ;
      RECT 21.74 3.672 21.785 3.83 ;
      RECT 21.72 2.96 21.74 3.238 ;
      RECT 21.72 3.665 21.74 3.826 ;
      RECT 21.69 2.96 21.72 3.26 ;
      RECT 21.68 3.632 21.72 3.823 ;
      RECT 21.675 2.96 21.69 3.28 ;
      RECT 21.675 3.597 21.68 3.821 ;
      RECT 21.67 2.96 21.675 3.405 ;
      RECT 21.67 3.557 21.675 3.821 ;
      RECT 21.66 2.96 21.67 3.821 ;
      RECT 21.585 2.96 21.66 3.815 ;
      RECT 21.555 2.96 21.585 3.805 ;
      RECT 21.55 2.96 21.555 3.797 ;
      RECT 21.545 3.002 21.55 3.79 ;
      RECT 21.535 3.071 21.545 3.781 ;
      RECT 21.53 3.141 21.535 3.733 ;
      RECT 21.525 3.205 21.53 3.63 ;
      RECT 21.52 3.24 21.525 3.585 ;
      RECT 21.518 3.277 21.52 3.477 ;
      RECT 21.515 3.285 21.518 3.47 ;
      RECT 21.51 3.35 21.515 3.413 ;
      RECT 25.585 2.44 25.865 2.72 ;
      RECT 25.575 2.44 25.865 2.583 ;
      RECT 25.53 2.305 25.79 2.565 ;
      RECT 25.53 2.42 25.845 2.565 ;
      RECT 25.53 2.39 25.84 2.565 ;
      RECT 25.53 2.377 25.83 2.565 ;
      RECT 25.53 2.367 25.825 2.565 ;
      RECT 21.505 2.35 21.765 2.61 ;
      RECT 25.275 1.9 25.535 2.16 ;
      RECT 25.265 1.925 25.535 2.12 ;
      RECT 25.26 1.925 25.265 2.119 ;
      RECT 25.19 1.92 25.26 2.111 ;
      RECT 25.105 1.907 25.19 2.094 ;
      RECT 25.101 1.899 25.105 2.084 ;
      RECT 25.015 1.892 25.101 2.074 ;
      RECT 25.006 1.884 25.015 2.064 ;
      RECT 24.92 1.877 25.006 2.052 ;
      RECT 24.9 1.868 24.92 2.038 ;
      RECT 24.845 1.863 24.9 2.03 ;
      RECT 24.835 1.857 24.845 2.024 ;
      RECT 24.815 1.855 24.835 2.02 ;
      RECT 24.807 1.854 24.815 2.016 ;
      RECT 24.721 1.846 24.807 2.005 ;
      RECT 24.635 1.832 24.721 1.985 ;
      RECT 24.575 1.82 24.635 1.97 ;
      RECT 24.565 1.815 24.575 1.965 ;
      RECT 24.515 1.815 24.565 1.967 ;
      RECT 24.468 1.817 24.515 1.971 ;
      RECT 24.382 1.824 24.468 1.976 ;
      RECT 24.296 1.832 24.382 1.982 ;
      RECT 24.21 1.841 24.296 1.988 ;
      RECT 24.151 1.847 24.21 1.993 ;
      RECT 24.065 1.852 24.151 1.999 ;
      RECT 23.99 1.857 24.065 2.005 ;
      RECT 23.951 1.859 23.99 2.01 ;
      RECT 23.865 1.856 23.951 2.015 ;
      RECT 23.78 1.854 23.865 2.022 ;
      RECT 23.748 1.853 23.78 2.025 ;
      RECT 23.662 1.852 23.748 2.026 ;
      RECT 23.576 1.851 23.662 2.027 ;
      RECT 23.49 1.85 23.576 2.027 ;
      RECT 23.404 1.849 23.49 2.028 ;
      RECT 23.318 1.848 23.404 2.029 ;
      RECT 23.232 1.847 23.318 2.03 ;
      RECT 23.146 1.846 23.232 2.03 ;
      RECT 23.06 1.845 23.146 2.031 ;
      RECT 23.01 1.845 23.06 2.032 ;
      RECT 22.996 1.846 23.01 2.032 ;
      RECT 22.91 1.853 22.996 2.033 ;
      RECT 22.836 1.864 22.91 2.034 ;
      RECT 22.75 1.873 22.836 2.035 ;
      RECT 22.715 1.88 22.75 2.05 ;
      RECT 22.69 1.883 22.715 2.08 ;
      RECT 22.665 1.892 22.69 2.109 ;
      RECT 22.655 1.903 22.665 2.129 ;
      RECT 22.645 1.911 22.655 2.143 ;
      RECT 22.64 1.917 22.645 2.153 ;
      RECT 22.615 1.934 22.64 2.17 ;
      RECT 22.6 1.956 22.615 2.198 ;
      RECT 22.57 1.982 22.6 2.228 ;
      RECT 22.55 2.011 22.57 2.258 ;
      RECT 22.545 2.026 22.55 2.275 ;
      RECT 22.525 2.041 22.545 2.29 ;
      RECT 22.515 2.059 22.525 2.308 ;
      RECT 22.505 2.07 22.515 2.323 ;
      RECT 22.455 2.102 22.505 2.349 ;
      RECT 22.45 2.132 22.455 2.369 ;
      RECT 22.44 2.145 22.45 2.375 ;
      RECT 22.431 2.155 22.44 2.383 ;
      RECT 22.42 2.166 22.431 2.391 ;
      RECT 22.415 2.176 22.42 2.397 ;
      RECT 22.4 2.197 22.415 2.404 ;
      RECT 22.385 2.227 22.4 2.412 ;
      RECT 22.35 2.257 22.385 2.418 ;
      RECT 22.325 2.275 22.35 2.425 ;
      RECT 22.275 2.283 22.325 2.434 ;
      RECT 22.25 2.288 22.275 2.443 ;
      RECT 22.195 2.294 22.25 2.453 ;
      RECT 22.19 2.299 22.195 2.461 ;
      RECT 22.176 2.302 22.19 2.463 ;
      RECT 22.09 2.314 22.176 2.475 ;
      RECT 22.08 2.326 22.09 2.488 ;
      RECT 21.995 2.339 22.08 2.5 ;
      RECT 21.951 2.356 21.995 2.514 ;
      RECT 21.865 2.373 21.951 2.53 ;
      RECT 21.835 2.387 21.865 2.544 ;
      RECT 21.825 2.392 21.835 2.549 ;
      RECT 21.765 2.395 21.825 2.558 ;
      RECT 24.655 2.665 24.915 2.925 ;
      RECT 24.655 2.665 24.935 2.778 ;
      RECT 24.655 2.665 24.96 2.745 ;
      RECT 24.655 2.665 24.965 2.725 ;
      RECT 24.705 2.44 24.985 2.72 ;
      RECT 24.26 3.175 24.52 3.435 ;
      RECT 24.25 3.032 24.445 3.373 ;
      RECT 24.245 3.14 24.46 3.365 ;
      RECT 24.24 3.19 24.52 3.355 ;
      RECT 24.23 3.267 24.52 3.34 ;
      RECT 24.25 3.115 24.46 3.373 ;
      RECT 24.26 2.99 24.445 3.435 ;
      RECT 24.26 2.885 24.425 3.435 ;
      RECT 24.27 2.872 24.425 3.435 ;
      RECT 24.27 2.83 24.415 3.435 ;
      RECT 24.275 2.755 24.415 3.435 ;
      RECT 24.305 2.405 24.415 3.435 ;
      RECT 24.31 2.135 24.435 2.758 ;
      RECT 24.28 2.71 24.435 2.758 ;
      RECT 24.295 2.512 24.415 3.435 ;
      RECT 24.285 2.622 24.435 2.758 ;
      RECT 24.31 2.135 24.45 2.615 ;
      RECT 24.31 2.135 24.47 2.49 ;
      RECT 24.275 2.135 24.535 2.395 ;
      RECT 23.745 2.44 24.025 2.72 ;
      RECT 23.73 2.44 24.025 2.7 ;
      RECT 21.785 3.305 22.045 3.565 ;
      RECT 23.57 3.16 23.83 3.42 ;
      RECT 23.55 3.18 23.83 3.395 ;
      RECT 23.507 3.18 23.55 3.394 ;
      RECT 23.421 3.181 23.507 3.391 ;
      RECT 23.335 3.182 23.421 3.387 ;
      RECT 23.26 3.184 23.335 3.384 ;
      RECT 23.237 3.185 23.26 3.382 ;
      RECT 23.151 3.186 23.237 3.38 ;
      RECT 23.065 3.187 23.151 3.377 ;
      RECT 23.041 3.188 23.065 3.375 ;
      RECT 22.955 3.19 23.041 3.372 ;
      RECT 22.87 3.192 22.955 3.373 ;
      RECT 22.813 3.193 22.87 3.379 ;
      RECT 22.727 3.195 22.813 3.389 ;
      RECT 22.641 3.198 22.727 3.402 ;
      RECT 22.555 3.2 22.641 3.414 ;
      RECT 22.541 3.201 22.555 3.421 ;
      RECT 22.455 3.202 22.541 3.429 ;
      RECT 22.415 3.204 22.455 3.438 ;
      RECT 22.406 3.205 22.415 3.441 ;
      RECT 22.32 3.213 22.406 3.447 ;
      RECT 22.3 3.222 22.32 3.455 ;
      RECT 22.215 3.237 22.3 3.463 ;
      RECT 22.155 3.26 22.215 3.474 ;
      RECT 22.145 3.272 22.155 3.479 ;
      RECT 22.105 3.282 22.145 3.483 ;
      RECT 22.05 3.299 22.105 3.491 ;
      RECT 22.045 3.309 22.05 3.495 ;
      RECT 23.111 2.44 23.17 2.837 ;
      RECT 23.025 2.44 23.23 2.828 ;
      RECT 23.02 2.47 23.23 2.823 ;
      RECT 22.986 2.47 23.23 2.821 ;
      RECT 22.9 2.47 23.23 2.815 ;
      RECT 22.855 2.47 23.25 2.793 ;
      RECT 22.855 2.47 23.27 2.748 ;
      RECT 22.815 2.47 23.27 2.738 ;
      RECT 23.025 2.44 23.305 2.72 ;
      RECT 22.76 2.44 23.02 2.7 ;
      RECT 21.945 1.92 22.205 2.18 ;
      RECT 22.025 1.88 22.305 2.16 ;
      RECT 16.395 6.22 16.715 6.545 ;
      RECT 16.425 5.695 16.595 6.545 ;
      RECT 16.425 5.695 16.6 6.045 ;
      RECT 16.425 5.695 17.4 5.87 ;
      RECT 17.225 1.965 17.4 5.87 ;
      RECT 17.17 1.965 17.52 2.315 ;
      RECT 17.195 6.655 17.52 6.98 ;
      RECT 16.08 6.745 17.52 6.915 ;
      RECT 16.08 2.395 16.24 6.915 ;
      RECT 16.395 2.365 16.715 2.685 ;
      RECT 16.08 2.395 16.715 2.565 ;
      RECT 4.805 3 5.085 3.28 ;
      RECT 4.775 3 5.085 3.265 ;
      RECT 4.77 3 5.085 3.263 ;
      RECT 4.765 1.33 4.935 3.257 ;
      RECT 4.76 2.967 5.03 3.25 ;
      RECT 4.755 3 5.085 3.243 ;
      RECT 4.725 2.97 5.03 3.23 ;
      RECT 4.725 2.997 5.05 3.23 ;
      RECT 4.725 2.987 5.045 3.23 ;
      RECT 4.725 2.972 5.04 3.23 ;
      RECT 4.765 2.962 5.03 3.257 ;
      RECT 4.765 2.957 5.02 3.257 ;
      RECT 4.765 2.956 5.005 3.257 ;
      RECT 14.735 1.34 15.085 1.69 ;
      RECT 14.73 1.34 15.085 1.595 ;
      RECT 4.765 1.33 14.975 1.5 ;
      RECT 14.41 2.85 14.78 3.22 ;
      RECT 14.495 2.235 14.665 3.22 ;
      RECT 10.515 2.455 10.75 2.715 ;
      RECT 13.66 2.235 13.825 2.495 ;
      RECT 13.565 2.225 13.58 2.495 ;
      RECT 13.66 2.235 14.665 2.415 ;
      RECT 12.165 1.795 12.205 1.935 ;
      RECT 13.58 2.23 13.66 2.495 ;
      RECT 13.525 2.225 13.565 2.461 ;
      RECT 13.511 2.225 13.525 2.461 ;
      RECT 13.425 2.23 13.511 2.463 ;
      RECT 13.38 2.237 13.425 2.465 ;
      RECT 13.35 2.237 13.38 2.467 ;
      RECT 13.325 2.232 13.35 2.469 ;
      RECT 13.295 2.228 13.325 2.478 ;
      RECT 13.285 2.225 13.295 2.49 ;
      RECT 13.28 2.225 13.285 2.498 ;
      RECT 13.275 2.225 13.28 2.503 ;
      RECT 13.265 2.224 13.275 2.513 ;
      RECT 13.26 2.223 13.265 2.523 ;
      RECT 13.245 2.222 13.26 2.528 ;
      RECT 13.217 2.219 13.245 2.555 ;
      RECT 13.131 2.211 13.217 2.555 ;
      RECT 13.045 2.2 13.131 2.555 ;
      RECT 13.005 2.185 13.045 2.555 ;
      RECT 12.965 2.159 13.005 2.555 ;
      RECT 12.96 2.141 12.965 2.367 ;
      RECT 12.95 2.137 12.96 2.357 ;
      RECT 12.935 2.127 12.95 2.344 ;
      RECT 12.915 2.111 12.935 2.329 ;
      RECT 12.9 2.096 12.915 2.314 ;
      RECT 12.89 2.085 12.9 2.304 ;
      RECT 12.865 2.069 12.89 2.293 ;
      RECT 12.86 2.056 12.865 2.283 ;
      RECT 12.855 2.052 12.86 2.278 ;
      RECT 12.8 2.038 12.855 2.256 ;
      RECT 12.761 2.019 12.8 2.22 ;
      RECT 12.675 1.993 12.761 2.173 ;
      RECT 12.671 1.975 12.675 2.139 ;
      RECT 12.585 1.956 12.671 2.117 ;
      RECT 12.58 1.938 12.585 2.095 ;
      RECT 12.575 1.936 12.58 2.093 ;
      RECT 12.565 1.935 12.575 2.088 ;
      RECT 12.505 1.922 12.565 2.074 ;
      RECT 12.46 1.9 12.505 2.053 ;
      RECT 12.4 1.877 12.46 2.032 ;
      RECT 12.336 1.852 12.4 2.007 ;
      RECT 12.25 1.822 12.336 1.976 ;
      RECT 12.235 1.802 12.25 1.955 ;
      RECT 12.205 1.797 12.235 1.946 ;
      RECT 12.152 1.795 12.165 1.935 ;
      RECT 12.066 1.795 12.152 1.937 ;
      RECT 11.98 1.795 12.066 1.939 ;
      RECT 11.96 1.795 11.98 1.943 ;
      RECT 11.915 1.797 11.96 1.954 ;
      RECT 11.875 1.807 11.915 1.97 ;
      RECT 11.871 1.816 11.875 1.978 ;
      RECT 11.785 1.836 11.871 1.994 ;
      RECT 11.775 1.855 11.785 2.012 ;
      RECT 11.77 1.857 11.775 2.015 ;
      RECT 11.76 1.861 11.77 2.018 ;
      RECT 11.74 1.866 11.76 2.028 ;
      RECT 11.71 1.876 11.74 2.048 ;
      RECT 11.705 1.883 11.71 2.062 ;
      RECT 11.695 1.887 11.705 2.069 ;
      RECT 11.68 1.895 11.695 2.08 ;
      RECT 11.67 1.905 11.68 2.091 ;
      RECT 11.66 1.912 11.67 2.099 ;
      RECT 11.635 1.925 11.66 2.114 ;
      RECT 11.571 1.961 11.635 2.153 ;
      RECT 11.485 2.024 11.571 2.217 ;
      RECT 11.45 2.075 11.485 2.27 ;
      RECT 11.445 2.092 11.45 2.287 ;
      RECT 11.43 2.101 11.445 2.294 ;
      RECT 11.41 2.116 11.43 2.308 ;
      RECT 11.405 2.127 11.41 2.318 ;
      RECT 11.385 2.14 11.405 2.328 ;
      RECT 11.38 2.15 11.385 2.338 ;
      RECT 11.365 2.155 11.38 2.347 ;
      RECT 11.355 2.165 11.365 2.358 ;
      RECT 11.325 2.182 11.355 2.375 ;
      RECT 11.315 2.2 11.325 2.393 ;
      RECT 11.3 2.211 11.315 2.404 ;
      RECT 11.26 2.235 11.3 2.42 ;
      RECT 11.225 2.269 11.26 2.437 ;
      RECT 11.195 2.292 11.225 2.449 ;
      RECT 11.18 2.302 11.195 2.458 ;
      RECT 11.14 2.312 11.18 2.469 ;
      RECT 11.12 2.323 11.14 2.481 ;
      RECT 11.115 2.327 11.12 2.488 ;
      RECT 11.1 2.331 11.115 2.493 ;
      RECT 11.09 2.336 11.1 2.498 ;
      RECT 11.085 2.339 11.09 2.501 ;
      RECT 11.055 2.345 11.085 2.508 ;
      RECT 11.02 2.355 11.055 2.522 ;
      RECT 10.96 2.37 11.02 2.542 ;
      RECT 10.905 2.39 10.96 2.566 ;
      RECT 10.876 2.405 10.905 2.584 ;
      RECT 10.79 2.425 10.876 2.609 ;
      RECT 10.785 2.44 10.79 2.629 ;
      RECT 10.775 2.443 10.785 2.63 ;
      RECT 10.75 2.45 10.775 2.715 ;
      RECT 13.445 2.943 13.725 3.28 ;
      RECT 13.445 2.953 13.73 3.238 ;
      RECT 13.445 2.962 13.735 3.135 ;
      RECT 13.445 2.977 13.74 3.003 ;
      RECT 13.445 2.805 13.705 3.28 ;
      RECT 3.025 6.995 3.315 7.345 ;
      RECT 3.025 7.055 4.44 7.225 ;
      RECT 4.27 6.685 4.44 7.225 ;
      RECT 12.59 6.605 12.94 6.955 ;
      RECT 4.27 6.685 12.94 6.855 ;
      RECT 11.165 3.685 11.175 3.875 ;
      RECT 9.425 3.56 9.705 3.84 ;
      RECT 12.47 2.5 12.475 2.985 ;
      RECT 12.365 2.5 12.425 2.76 ;
      RECT 12.69 3.47 12.695 3.545 ;
      RECT 12.68 3.337 12.69 3.58 ;
      RECT 12.67 3.172 12.68 3.601 ;
      RECT 12.665 3.042 12.67 3.617 ;
      RECT 12.655 2.932 12.665 3.633 ;
      RECT 12.65 2.831 12.655 3.65 ;
      RECT 12.645 2.813 12.65 3.66 ;
      RECT 12.64 2.795 12.645 3.67 ;
      RECT 12.63 2.77 12.64 3.685 ;
      RECT 12.625 2.75 12.63 3.7 ;
      RECT 12.605 2.5 12.625 3.725 ;
      RECT 12.59 2.5 12.605 3.758 ;
      RECT 12.56 2.5 12.59 3.78 ;
      RECT 12.54 2.5 12.56 3.794 ;
      RECT 12.52 2.5 12.54 3.31 ;
      RECT 12.535 3.377 12.54 3.799 ;
      RECT 12.53 3.407 12.535 3.801 ;
      RECT 12.525 3.42 12.53 3.804 ;
      RECT 12.52 3.43 12.525 3.808 ;
      RECT 12.515 2.5 12.52 3.228 ;
      RECT 12.515 3.44 12.52 3.81 ;
      RECT 12.51 2.5 12.515 3.205 ;
      RECT 12.5 3.462 12.515 3.81 ;
      RECT 12.495 2.5 12.51 3.15 ;
      RECT 12.49 3.487 12.5 3.81 ;
      RECT 12.49 2.5 12.495 3.095 ;
      RECT 12.48 2.5 12.49 3.043 ;
      RECT 12.485 3.5 12.49 3.811 ;
      RECT 12.48 3.512 12.485 3.812 ;
      RECT 12.475 2.5 12.48 3.003 ;
      RECT 12.475 3.525 12.48 3.813 ;
      RECT 12.46 3.54 12.475 3.814 ;
      RECT 12.465 2.5 12.47 2.965 ;
      RECT 12.46 2.5 12.465 2.93 ;
      RECT 12.455 2.5 12.46 2.905 ;
      RECT 12.45 3.567 12.46 3.816 ;
      RECT 12.445 2.5 12.455 2.863 ;
      RECT 12.445 3.585 12.45 3.817 ;
      RECT 12.44 2.5 12.445 2.823 ;
      RECT 12.44 3.592 12.445 3.818 ;
      RECT 12.435 2.5 12.44 2.795 ;
      RECT 12.43 3.61 12.44 3.819 ;
      RECT 12.425 2.5 12.435 2.775 ;
      RECT 12.42 3.63 12.43 3.821 ;
      RECT 12.41 3.647 12.42 3.822 ;
      RECT 12.375 3.67 12.41 3.825 ;
      RECT 12.32 3.688 12.375 3.831 ;
      RECT 12.234 3.696 12.32 3.84 ;
      RECT 12.148 3.707 12.234 3.851 ;
      RECT 12.062 3.717 12.148 3.862 ;
      RECT 11.976 3.727 12.062 3.874 ;
      RECT 11.89 3.737 11.976 3.885 ;
      RECT 11.87 3.743 11.89 3.891 ;
      RECT 11.79 3.745 11.87 3.895 ;
      RECT 11.785 3.744 11.79 3.9 ;
      RECT 11.777 3.743 11.785 3.9 ;
      RECT 11.691 3.739 11.777 3.898 ;
      RECT 11.605 3.731 11.691 3.895 ;
      RECT 11.519 3.722 11.605 3.891 ;
      RECT 11.433 3.714 11.519 3.888 ;
      RECT 11.347 3.706 11.433 3.884 ;
      RECT 11.261 3.697 11.347 3.881 ;
      RECT 11.175 3.689 11.261 3.877 ;
      RECT 11.12 3.682 11.165 3.875 ;
      RECT 11.035 3.675 11.12 3.873 ;
      RECT 10.961 3.667 11.035 3.869 ;
      RECT 10.875 3.659 10.961 3.866 ;
      RECT 10.872 3.655 10.875 3.864 ;
      RECT 10.786 3.651 10.872 3.863 ;
      RECT 10.7 3.643 10.786 3.86 ;
      RECT 10.615 3.638 10.7 3.857 ;
      RECT 10.529 3.635 10.615 3.854 ;
      RECT 10.443 3.633 10.529 3.851 ;
      RECT 10.357 3.63 10.443 3.848 ;
      RECT 10.271 3.627 10.357 3.845 ;
      RECT 10.185 3.624 10.271 3.842 ;
      RECT 10.109 3.622 10.185 3.839 ;
      RECT 10.023 3.619 10.109 3.836 ;
      RECT 9.937 3.616 10.023 3.834 ;
      RECT 9.851 3.614 9.937 3.831 ;
      RECT 9.765 3.611 9.851 3.828 ;
      RECT 9.705 3.602 9.765 3.826 ;
      RECT 12.215 3.22 12.29 3.48 ;
      RECT 12.195 3.2 12.2 3.48 ;
      RECT 11.515 2.985 11.62 3.28 ;
      RECT 5.96 2.96 6.03 3.22 ;
      RECT 11.855 2.835 11.86 3.206 ;
      RECT 11.845 2.89 11.85 3.206 ;
      RECT 12.15 2.06 12.21 2.32 ;
      RECT 12.205 3.215 12.215 3.48 ;
      RECT 12.2 3.205 12.205 3.48 ;
      RECT 12.12 3.152 12.195 3.48 ;
      RECT 12.145 2.06 12.15 2.34 ;
      RECT 12.135 2.06 12.145 2.36 ;
      RECT 12.12 2.06 12.135 2.39 ;
      RECT 12.105 2.06 12.12 2.433 ;
      RECT 12.1 3.095 12.12 3.48 ;
      RECT 12.09 2.06 12.105 2.47 ;
      RECT 12.085 3.075 12.1 3.48 ;
      RECT 12.085 2.06 12.09 2.493 ;
      RECT 12.075 2.06 12.085 2.518 ;
      RECT 12.045 3.042 12.085 3.48 ;
      RECT 12.05 2.06 12.075 2.568 ;
      RECT 12.045 2.06 12.05 2.623 ;
      RECT 12.04 2.06 12.045 2.665 ;
      RECT 12.03 3.005 12.045 3.48 ;
      RECT 12.035 2.06 12.04 2.708 ;
      RECT 12.03 2.06 12.035 2.773 ;
      RECT 12.025 2.06 12.03 2.795 ;
      RECT 12.025 2.993 12.03 3.345 ;
      RECT 12.02 2.06 12.025 2.863 ;
      RECT 12.02 2.985 12.025 3.328 ;
      RECT 12.015 2.06 12.02 2.908 ;
      RECT 12.01 2.967 12.02 3.305 ;
      RECT 12.01 2.06 12.015 2.945 ;
      RECT 12 2.06 12.01 3.285 ;
      RECT 11.995 2.06 12 3.268 ;
      RECT 11.99 2.06 11.995 3.253 ;
      RECT 11.985 2.06 11.99 3.238 ;
      RECT 11.965 2.06 11.985 3.228 ;
      RECT 11.96 2.06 11.965 3.218 ;
      RECT 11.95 2.06 11.96 3.214 ;
      RECT 11.945 2.337 11.95 3.213 ;
      RECT 11.94 2.36 11.945 3.212 ;
      RECT 11.935 2.39 11.94 3.211 ;
      RECT 11.93 2.417 11.935 3.21 ;
      RECT 11.925 2.445 11.93 3.21 ;
      RECT 11.92 2.472 11.925 3.21 ;
      RECT 11.915 2.492 11.92 3.21 ;
      RECT 11.91 2.52 11.915 3.21 ;
      RECT 11.9 2.562 11.91 3.21 ;
      RECT 11.89 2.607 11.9 3.209 ;
      RECT 11.885 2.66 11.89 3.208 ;
      RECT 11.88 2.692 11.885 3.207 ;
      RECT 11.875 2.712 11.88 3.206 ;
      RECT 11.87 2.75 11.875 3.206 ;
      RECT 11.865 2.772 11.87 3.206 ;
      RECT 11.86 2.797 11.865 3.206 ;
      RECT 11.85 2.862 11.855 3.206 ;
      RECT 11.835 2.922 11.845 3.206 ;
      RECT 11.82 2.932 11.835 3.206 ;
      RECT 11.8 2.942 11.82 3.206 ;
      RECT 11.77 2.947 11.8 3.203 ;
      RECT 11.71 2.957 11.77 3.2 ;
      RECT 11.69 2.966 11.71 3.205 ;
      RECT 11.665 2.972 11.69 3.218 ;
      RECT 11.645 2.977 11.665 3.233 ;
      RECT 11.62 2.982 11.645 3.28 ;
      RECT 11.491 2.984 11.515 3.28 ;
      RECT 11.405 2.979 11.491 3.28 ;
      RECT 11.365 2.976 11.405 3.28 ;
      RECT 11.315 2.978 11.365 3.26 ;
      RECT 11.285 2.982 11.315 3.26 ;
      RECT 11.206 2.992 11.285 3.26 ;
      RECT 11.12 3.007 11.206 3.261 ;
      RECT 11.07 3.017 11.12 3.262 ;
      RECT 11.062 3.02 11.07 3.262 ;
      RECT 10.976 3.022 11.062 3.263 ;
      RECT 10.89 3.026 10.976 3.263 ;
      RECT 10.804 3.03 10.89 3.264 ;
      RECT 10.718 3.033 10.804 3.265 ;
      RECT 10.632 3.037 10.718 3.265 ;
      RECT 10.546 3.041 10.632 3.266 ;
      RECT 10.46 3.044 10.546 3.267 ;
      RECT 10.374 3.048 10.46 3.267 ;
      RECT 10.288 3.052 10.374 3.268 ;
      RECT 10.202 3.056 10.288 3.269 ;
      RECT 10.116 3.059 10.202 3.269 ;
      RECT 10.03 3.063 10.116 3.27 ;
      RECT 10 3.065 10.03 3.27 ;
      RECT 9.914 3.068 10 3.271 ;
      RECT 9.828 3.072 9.914 3.272 ;
      RECT 9.742 3.076 9.828 3.273 ;
      RECT 9.656 3.079 9.742 3.273 ;
      RECT 9.57 3.083 9.656 3.274 ;
      RECT 9.535 3.088 9.57 3.275 ;
      RECT 9.48 3.098 9.535 3.282 ;
      RECT 9.455 3.11 9.48 3.292 ;
      RECT 9.42 3.123 9.455 3.3 ;
      RECT 9.38 3.14 9.42 3.323 ;
      RECT 9.36 3.153 9.38 3.35 ;
      RECT 9.33 3.165 9.36 3.378 ;
      RECT 9.325 3.173 9.33 3.398 ;
      RECT 9.32 3.176 9.325 3.408 ;
      RECT 9.27 3.188 9.32 3.442 ;
      RECT 9.26 3.203 9.27 3.475 ;
      RECT 9.25 3.209 9.26 3.488 ;
      RECT 9.24 3.216 9.25 3.5 ;
      RECT 9.215 3.229 9.24 3.518 ;
      RECT 9.2 3.244 9.215 3.54 ;
      RECT 9.19 3.252 9.2 3.556 ;
      RECT 9.175 3.261 9.19 3.571 ;
      RECT 9.165 3.271 9.175 3.585 ;
      RECT 9.146 3.284 9.165 3.602 ;
      RECT 9.06 3.329 9.146 3.667 ;
      RECT 9.045 3.374 9.06 3.725 ;
      RECT 9.04 3.383 9.045 3.738 ;
      RECT 9.03 3.39 9.04 3.743 ;
      RECT 9.025 3.395 9.03 3.747 ;
      RECT 9.005 3.405 9.025 3.754 ;
      RECT 8.98 3.425 9.005 3.768 ;
      RECT 8.945 3.45 8.98 3.788 ;
      RECT 8.93 3.473 8.945 3.803 ;
      RECT 8.92 3.483 8.93 3.808 ;
      RECT 8.91 3.491 8.92 3.815 ;
      RECT 8.9 3.5 8.91 3.821 ;
      RECT 8.88 3.512 8.9 3.823 ;
      RECT 8.87 3.525 8.88 3.825 ;
      RECT 8.845 3.54 8.87 3.828 ;
      RECT 8.825 3.557 8.845 3.832 ;
      RECT 8.785 3.585 8.825 3.838 ;
      RECT 8.72 3.632 8.785 3.847 ;
      RECT 8.705 3.665 8.72 3.855 ;
      RECT 8.7 3.672 8.705 3.857 ;
      RECT 8.65 3.697 8.7 3.862 ;
      RECT 8.635 3.721 8.65 3.869 ;
      RECT 8.585 3.726 8.635 3.87 ;
      RECT 8.499 3.73 8.585 3.87 ;
      RECT 8.413 3.73 8.499 3.87 ;
      RECT 8.327 3.73 8.413 3.871 ;
      RECT 8.241 3.73 8.327 3.871 ;
      RECT 8.155 3.73 8.241 3.871 ;
      RECT 8.089 3.73 8.155 3.871 ;
      RECT 8.003 3.73 8.089 3.872 ;
      RECT 7.917 3.73 8.003 3.872 ;
      RECT 7.831 3.731 7.917 3.873 ;
      RECT 7.745 3.731 7.831 3.873 ;
      RECT 7.659 3.731 7.745 3.873 ;
      RECT 7.573 3.731 7.659 3.874 ;
      RECT 7.487 3.731 7.573 3.874 ;
      RECT 7.401 3.732 7.487 3.875 ;
      RECT 7.315 3.732 7.401 3.875 ;
      RECT 7.295 3.732 7.315 3.875 ;
      RECT 7.209 3.732 7.295 3.875 ;
      RECT 7.123 3.732 7.209 3.875 ;
      RECT 7.037 3.733 7.123 3.875 ;
      RECT 6.951 3.733 7.037 3.875 ;
      RECT 6.865 3.733 6.951 3.875 ;
      RECT 6.779 3.734 6.865 3.875 ;
      RECT 6.693 3.734 6.779 3.875 ;
      RECT 6.607 3.734 6.693 3.875 ;
      RECT 6.521 3.734 6.607 3.875 ;
      RECT 6.435 3.735 6.521 3.875 ;
      RECT 6.385 3.732 6.435 3.875 ;
      RECT 6.375 3.73 6.385 3.874 ;
      RECT 6.371 3.73 6.375 3.873 ;
      RECT 6.285 3.725 6.371 3.868 ;
      RECT 6.263 3.718 6.285 3.862 ;
      RECT 6.177 3.709 6.263 3.856 ;
      RECT 6.091 3.696 6.177 3.847 ;
      RECT 6.005 3.682 6.091 3.837 ;
      RECT 5.96 3.672 6.005 3.83 ;
      RECT 5.94 2.96 5.96 3.238 ;
      RECT 5.94 3.665 5.96 3.826 ;
      RECT 5.91 2.96 5.94 3.26 ;
      RECT 5.9 3.632 5.94 3.823 ;
      RECT 5.895 2.96 5.91 3.28 ;
      RECT 5.895 3.597 5.9 3.821 ;
      RECT 5.89 2.96 5.895 3.405 ;
      RECT 5.89 3.557 5.895 3.821 ;
      RECT 5.88 2.96 5.89 3.821 ;
      RECT 5.805 2.96 5.88 3.815 ;
      RECT 5.775 2.96 5.805 3.805 ;
      RECT 5.77 2.96 5.775 3.797 ;
      RECT 5.765 3.002 5.77 3.79 ;
      RECT 5.755 3.071 5.765 3.781 ;
      RECT 5.75 3.141 5.755 3.733 ;
      RECT 5.745 3.205 5.75 3.63 ;
      RECT 5.74 3.24 5.745 3.585 ;
      RECT 5.738 3.277 5.74 3.477 ;
      RECT 5.735 3.285 5.738 3.47 ;
      RECT 5.73 3.35 5.735 3.413 ;
      RECT 9.805 2.44 10.085 2.72 ;
      RECT 9.795 2.44 10.085 2.583 ;
      RECT 9.75 2.305 10.01 2.565 ;
      RECT 9.75 2.42 10.065 2.565 ;
      RECT 9.75 2.39 10.06 2.565 ;
      RECT 9.75 2.377 10.05 2.565 ;
      RECT 9.75 2.367 10.045 2.565 ;
      RECT 5.725 2.35 5.985 2.61 ;
      RECT 9.495 1.9 9.755 2.16 ;
      RECT 9.485 1.925 9.755 2.12 ;
      RECT 9.48 1.925 9.485 2.119 ;
      RECT 9.41 1.92 9.48 2.111 ;
      RECT 9.325 1.907 9.41 2.094 ;
      RECT 9.321 1.899 9.325 2.084 ;
      RECT 9.235 1.892 9.321 2.074 ;
      RECT 9.226 1.884 9.235 2.064 ;
      RECT 9.14 1.877 9.226 2.052 ;
      RECT 9.12 1.868 9.14 2.038 ;
      RECT 9.065 1.863 9.12 2.03 ;
      RECT 9.055 1.857 9.065 2.024 ;
      RECT 9.035 1.855 9.055 2.02 ;
      RECT 9.027 1.854 9.035 2.016 ;
      RECT 8.941 1.846 9.027 2.005 ;
      RECT 8.855 1.832 8.941 1.985 ;
      RECT 8.795 1.82 8.855 1.97 ;
      RECT 8.785 1.815 8.795 1.965 ;
      RECT 8.735 1.815 8.785 1.967 ;
      RECT 8.688 1.817 8.735 1.971 ;
      RECT 8.602 1.824 8.688 1.976 ;
      RECT 8.516 1.832 8.602 1.982 ;
      RECT 8.43 1.841 8.516 1.988 ;
      RECT 8.371 1.847 8.43 1.993 ;
      RECT 8.285 1.852 8.371 1.999 ;
      RECT 8.21 1.857 8.285 2.005 ;
      RECT 8.171 1.859 8.21 2.01 ;
      RECT 8.085 1.856 8.171 2.015 ;
      RECT 8 1.854 8.085 2.022 ;
      RECT 7.968 1.853 8 2.025 ;
      RECT 7.882 1.852 7.968 2.026 ;
      RECT 7.796 1.851 7.882 2.027 ;
      RECT 7.71 1.85 7.796 2.027 ;
      RECT 7.624 1.849 7.71 2.028 ;
      RECT 7.538 1.848 7.624 2.029 ;
      RECT 7.452 1.847 7.538 2.03 ;
      RECT 7.366 1.846 7.452 2.03 ;
      RECT 7.28 1.845 7.366 2.031 ;
      RECT 7.23 1.845 7.28 2.032 ;
      RECT 7.216 1.846 7.23 2.032 ;
      RECT 7.13 1.853 7.216 2.033 ;
      RECT 7.056 1.864 7.13 2.034 ;
      RECT 6.97 1.873 7.056 2.035 ;
      RECT 6.935 1.88 6.97 2.05 ;
      RECT 6.91 1.883 6.935 2.08 ;
      RECT 6.885 1.892 6.91 2.109 ;
      RECT 6.875 1.903 6.885 2.129 ;
      RECT 6.865 1.911 6.875 2.143 ;
      RECT 6.86 1.917 6.865 2.153 ;
      RECT 6.835 1.934 6.86 2.17 ;
      RECT 6.82 1.956 6.835 2.198 ;
      RECT 6.79 1.982 6.82 2.228 ;
      RECT 6.77 2.011 6.79 2.258 ;
      RECT 6.765 2.026 6.77 2.275 ;
      RECT 6.745 2.041 6.765 2.29 ;
      RECT 6.735 2.059 6.745 2.308 ;
      RECT 6.725 2.07 6.735 2.323 ;
      RECT 6.675 2.102 6.725 2.349 ;
      RECT 6.67 2.132 6.675 2.369 ;
      RECT 6.66 2.145 6.67 2.375 ;
      RECT 6.651 2.155 6.66 2.383 ;
      RECT 6.64 2.166 6.651 2.391 ;
      RECT 6.635 2.176 6.64 2.397 ;
      RECT 6.62 2.197 6.635 2.404 ;
      RECT 6.605 2.227 6.62 2.412 ;
      RECT 6.57 2.257 6.605 2.418 ;
      RECT 6.545 2.275 6.57 2.425 ;
      RECT 6.495 2.283 6.545 2.434 ;
      RECT 6.47 2.288 6.495 2.443 ;
      RECT 6.415 2.294 6.47 2.453 ;
      RECT 6.41 2.299 6.415 2.461 ;
      RECT 6.396 2.302 6.41 2.463 ;
      RECT 6.31 2.314 6.396 2.475 ;
      RECT 6.3 2.326 6.31 2.488 ;
      RECT 6.215 2.339 6.3 2.5 ;
      RECT 6.171 2.356 6.215 2.514 ;
      RECT 6.085 2.373 6.171 2.53 ;
      RECT 6.055 2.387 6.085 2.544 ;
      RECT 6.045 2.392 6.055 2.549 ;
      RECT 5.985 2.395 6.045 2.558 ;
      RECT 8.875 2.665 9.135 2.925 ;
      RECT 8.875 2.665 9.155 2.778 ;
      RECT 8.875 2.665 9.18 2.745 ;
      RECT 8.875 2.665 9.185 2.725 ;
      RECT 8.925 2.44 9.205 2.72 ;
      RECT 8.48 3.175 8.74 3.435 ;
      RECT 8.47 3.032 8.665 3.373 ;
      RECT 8.465 3.14 8.68 3.365 ;
      RECT 8.46 3.19 8.74 3.355 ;
      RECT 8.45 3.267 8.74 3.34 ;
      RECT 8.47 3.115 8.68 3.373 ;
      RECT 8.48 2.99 8.665 3.435 ;
      RECT 8.48 2.885 8.645 3.435 ;
      RECT 8.49 2.872 8.645 3.435 ;
      RECT 8.49 2.83 8.635 3.435 ;
      RECT 8.495 2.755 8.635 3.435 ;
      RECT 8.525 2.405 8.635 3.435 ;
      RECT 8.53 2.135 8.655 2.758 ;
      RECT 8.5 2.71 8.655 2.758 ;
      RECT 8.515 2.512 8.635 3.435 ;
      RECT 8.505 2.622 8.655 2.758 ;
      RECT 8.53 2.135 8.67 2.615 ;
      RECT 8.53 2.135 8.69 2.49 ;
      RECT 8.495 2.135 8.755 2.395 ;
      RECT 7.965 2.44 8.245 2.72 ;
      RECT 7.95 2.44 8.245 2.7 ;
      RECT 6.005 3.305 6.265 3.565 ;
      RECT 7.79 3.16 8.05 3.42 ;
      RECT 7.77 3.18 8.05 3.395 ;
      RECT 7.727 3.18 7.77 3.394 ;
      RECT 7.641 3.181 7.727 3.391 ;
      RECT 7.555 3.182 7.641 3.387 ;
      RECT 7.48 3.184 7.555 3.384 ;
      RECT 7.457 3.185 7.48 3.382 ;
      RECT 7.371 3.186 7.457 3.38 ;
      RECT 7.285 3.187 7.371 3.377 ;
      RECT 7.261 3.188 7.285 3.375 ;
      RECT 7.175 3.19 7.261 3.372 ;
      RECT 7.09 3.192 7.175 3.373 ;
      RECT 7.033 3.193 7.09 3.379 ;
      RECT 6.947 3.195 7.033 3.389 ;
      RECT 6.861 3.198 6.947 3.402 ;
      RECT 6.775 3.2 6.861 3.414 ;
      RECT 6.761 3.201 6.775 3.421 ;
      RECT 6.675 3.202 6.761 3.429 ;
      RECT 6.635 3.204 6.675 3.438 ;
      RECT 6.626 3.205 6.635 3.441 ;
      RECT 6.54 3.213 6.626 3.447 ;
      RECT 6.52 3.222 6.54 3.455 ;
      RECT 6.435 3.237 6.52 3.463 ;
      RECT 6.375 3.26 6.435 3.474 ;
      RECT 6.365 3.272 6.375 3.479 ;
      RECT 6.325 3.282 6.365 3.483 ;
      RECT 6.27 3.299 6.325 3.491 ;
      RECT 6.265 3.309 6.27 3.495 ;
      RECT 7.331 2.44 7.39 2.837 ;
      RECT 7.245 2.44 7.45 2.828 ;
      RECT 7.24 2.47 7.45 2.823 ;
      RECT 7.206 2.47 7.45 2.821 ;
      RECT 7.12 2.47 7.45 2.815 ;
      RECT 7.075 2.47 7.47 2.793 ;
      RECT 7.075 2.47 7.49 2.748 ;
      RECT 7.035 2.47 7.49 2.738 ;
      RECT 7.245 2.44 7.525 2.72 ;
      RECT 6.98 2.44 7.24 2.7 ;
      RECT 6.165 1.92 6.425 2.18 ;
      RECT 6.245 1.88 6.525 2.16 ;
      RECT 76.755 0.815 77.125 1.185 ;
      RECT 75.045 7.04 75.415 7.41 ;
      RECT 60.97 0.815 61.34 1.185 ;
      RECT 59.26 7.04 59.63 7.41 ;
      RECT 45.185 0.815 45.555 1.185 ;
      RECT 43.475 7.04 43.845 7.41 ;
      RECT 29.41 0.815 29.78 1.185 ;
      RECT 27.7 7.04 28.07 7.41 ;
      RECT 13.63 0.815 14 1.185 ;
      RECT 11.92 7.04 12.29 7.41 ;
    LAYER via1 ;
      RECT 82.78 7.375 82.93 7.525 ;
      RECT 80.41 6.74 80.56 6.89 ;
      RECT 80.395 2.065 80.545 2.215 ;
      RECT 79.605 2.45 79.755 2.6 ;
      RECT 79.605 6.325 79.755 6.475 ;
      RECT 77.96 1.44 78.11 1.59 ;
      RECT 77.645 2.96 77.795 3.11 ;
      RECT 76.865 0.925 77.015 1.075 ;
      RECT 76.745 2.29 76.895 2.44 ;
      RECT 76.625 2.86 76.775 3.01 ;
      RECT 75.795 6.71 75.945 6.86 ;
      RECT 75.545 2.555 75.695 2.705 ;
      RECT 75.21 3.275 75.36 3.425 ;
      RECT 75.155 7.15 75.305 7.3 ;
      RECT 75.13 2.115 75.28 2.265 ;
      RECT 73.695 2.51 73.845 2.66 ;
      RECT 72.93 2.36 73.08 2.51 ;
      RECT 72.675 1.955 72.825 2.105 ;
      RECT 72.055 2.72 72.205 2.87 ;
      RECT 71.675 2.19 71.825 2.34 ;
      RECT 71.66 3.23 71.81 3.38 ;
      RECT 71.13 2.495 71.28 2.645 ;
      RECT 70.97 3.215 71.12 3.365 ;
      RECT 70.16 2.495 70.31 2.645 ;
      RECT 69.345 1.975 69.495 2.125 ;
      RECT 69.185 3.36 69.335 3.51 ;
      RECT 68.95 3.015 69.1 3.165 ;
      RECT 68.905 2.405 69.055 2.555 ;
      RECT 67.905 3.025 68.055 3.175 ;
      RECT 66.97 6.755 67.12 6.905 ;
      RECT 64.625 6.74 64.775 6.89 ;
      RECT 64.61 2.065 64.76 2.215 ;
      RECT 63.82 2.45 63.97 2.6 ;
      RECT 63.82 6.325 63.97 6.475 ;
      RECT 62.175 1.44 62.325 1.59 ;
      RECT 61.86 2.96 62.01 3.11 ;
      RECT 61.08 0.925 61.23 1.075 ;
      RECT 60.96 2.29 61.11 2.44 ;
      RECT 60.84 2.86 60.99 3.01 ;
      RECT 60.01 6.71 60.16 6.86 ;
      RECT 59.76 2.555 59.91 2.705 ;
      RECT 59.425 3.275 59.575 3.425 ;
      RECT 59.37 7.15 59.52 7.3 ;
      RECT 59.345 2.115 59.495 2.265 ;
      RECT 57.91 2.51 58.06 2.66 ;
      RECT 57.145 2.36 57.295 2.51 ;
      RECT 56.89 1.955 57.04 2.105 ;
      RECT 56.27 2.72 56.42 2.87 ;
      RECT 55.89 2.19 56.04 2.34 ;
      RECT 55.875 3.23 56.025 3.38 ;
      RECT 55.345 2.495 55.495 2.645 ;
      RECT 55.185 3.215 55.335 3.365 ;
      RECT 54.375 2.495 54.525 2.645 ;
      RECT 53.56 1.975 53.71 2.125 ;
      RECT 53.4 3.36 53.55 3.51 ;
      RECT 53.165 3.015 53.315 3.165 ;
      RECT 53.12 2.405 53.27 2.555 ;
      RECT 52.12 3.025 52.27 3.175 ;
      RECT 51.185 6.755 51.335 6.905 ;
      RECT 48.84 6.74 48.99 6.89 ;
      RECT 48.825 2.065 48.975 2.215 ;
      RECT 48.035 2.45 48.185 2.6 ;
      RECT 48.035 6.325 48.185 6.475 ;
      RECT 46.39 1.44 46.54 1.59 ;
      RECT 46.075 2.96 46.225 3.11 ;
      RECT 45.295 0.925 45.445 1.075 ;
      RECT 45.175 2.29 45.325 2.44 ;
      RECT 45.055 2.86 45.205 3.01 ;
      RECT 44.28 6.715 44.43 6.865 ;
      RECT 43.975 2.555 44.125 2.705 ;
      RECT 43.64 3.275 43.79 3.425 ;
      RECT 43.585 7.15 43.735 7.3 ;
      RECT 43.56 2.115 43.71 2.265 ;
      RECT 42.125 2.51 42.275 2.66 ;
      RECT 41.36 2.36 41.51 2.51 ;
      RECT 41.105 1.955 41.255 2.105 ;
      RECT 40.485 2.72 40.635 2.87 ;
      RECT 40.105 2.19 40.255 2.34 ;
      RECT 40.09 3.23 40.24 3.38 ;
      RECT 39.56 2.495 39.71 2.645 ;
      RECT 39.4 3.215 39.55 3.365 ;
      RECT 38.59 2.495 38.74 2.645 ;
      RECT 37.775 1.975 37.925 2.125 ;
      RECT 37.615 3.36 37.765 3.51 ;
      RECT 37.38 3.015 37.53 3.165 ;
      RECT 37.335 2.405 37.485 2.555 ;
      RECT 36.335 3.025 36.485 3.175 ;
      RECT 35.455 6.76 35.605 6.91 ;
      RECT 33.065 6.74 33.215 6.89 ;
      RECT 33.05 2.065 33.2 2.215 ;
      RECT 32.26 2.45 32.41 2.6 ;
      RECT 32.26 6.325 32.41 6.475 ;
      RECT 30.615 1.44 30.765 1.59 ;
      RECT 30.3 2.96 30.45 3.11 ;
      RECT 29.52 0.925 29.67 1.075 ;
      RECT 29.4 2.29 29.55 2.44 ;
      RECT 29.28 2.86 29.43 3.01 ;
      RECT 28.5 6.71 28.65 6.86 ;
      RECT 28.2 2.555 28.35 2.705 ;
      RECT 27.865 3.275 28.015 3.425 ;
      RECT 27.81 7.15 27.96 7.3 ;
      RECT 27.785 2.115 27.935 2.265 ;
      RECT 26.35 2.51 26.5 2.66 ;
      RECT 25.585 2.36 25.735 2.51 ;
      RECT 25.33 1.955 25.48 2.105 ;
      RECT 24.71 2.72 24.86 2.87 ;
      RECT 24.33 2.19 24.48 2.34 ;
      RECT 24.315 3.23 24.465 3.38 ;
      RECT 23.785 2.495 23.935 2.645 ;
      RECT 23.625 3.215 23.775 3.365 ;
      RECT 22.815 2.495 22.965 2.645 ;
      RECT 22 1.975 22.15 2.125 ;
      RECT 21.84 3.36 21.99 3.51 ;
      RECT 21.605 3.015 21.755 3.165 ;
      RECT 21.56 2.405 21.71 2.555 ;
      RECT 20.56 3.025 20.71 3.175 ;
      RECT 19.675 6.755 19.825 6.905 ;
      RECT 17.285 6.74 17.435 6.89 ;
      RECT 17.27 2.065 17.42 2.215 ;
      RECT 16.48 2.45 16.63 2.6 ;
      RECT 16.48 6.325 16.63 6.475 ;
      RECT 14.835 1.44 14.985 1.59 ;
      RECT 14.52 2.96 14.67 3.11 ;
      RECT 13.74 0.925 13.89 1.075 ;
      RECT 13.62 2.29 13.77 2.44 ;
      RECT 13.5 2.86 13.65 3.01 ;
      RECT 12.69 6.705 12.84 6.855 ;
      RECT 12.42 2.555 12.57 2.705 ;
      RECT 12.085 3.275 12.235 3.425 ;
      RECT 12.03 7.15 12.18 7.3 ;
      RECT 12.005 2.115 12.155 2.265 ;
      RECT 10.57 2.51 10.72 2.66 ;
      RECT 9.805 2.36 9.955 2.51 ;
      RECT 9.55 1.955 9.7 2.105 ;
      RECT 8.93 2.72 9.08 2.87 ;
      RECT 8.55 2.19 8.7 2.34 ;
      RECT 8.535 3.23 8.685 3.38 ;
      RECT 8.005 2.495 8.155 2.645 ;
      RECT 7.845 3.215 7.995 3.365 ;
      RECT 7.035 2.495 7.185 2.645 ;
      RECT 6.22 1.975 6.37 2.125 ;
      RECT 6.06 3.36 6.21 3.51 ;
      RECT 5.825 3.015 5.975 3.165 ;
      RECT 5.78 2.405 5.93 2.555 ;
      RECT 4.78 3.025 4.93 3.175 ;
      RECT 3.095 7.095 3.245 7.245 ;
      RECT 2.72 6.355 2.87 6.505 ;
    LAYER met1 ;
      RECT 67.655 1.26 77.315 1.74 ;
      RECT 51.87 1.26 61.53 1.74 ;
      RECT 36.085 1.26 45.745 1.74 ;
      RECT 20.31 1.26 29.97 1.74 ;
      RECT 4.53 1.26 14.19 1.74 ;
      RECT 67.655 1.26 77.37 1.59 ;
      RECT 51.87 1.26 61.585 1.59 ;
      RECT 36.085 1.26 45.8 1.59 ;
      RECT 20.31 1.26 30.025 1.59 ;
      RECT 4.53 1.26 14.245 1.59 ;
      RECT 67.77 0 77.485 1.585 ;
      RECT 51.985 0 61.7 1.585 ;
      RECT 36.2 0 45.915 1.585 ;
      RECT 20.425 0 30.14 1.585 ;
      RECT 4.645 0 14.36 1.585 ;
      RECT 83.07 0 83.25 0.305 ;
      RECT 67.285 0 81.12 0.305 ;
      RECT 51.5 0 65.335 0.305 ;
      RECT 35.725 0 49.55 0.305 ;
      RECT 19.945 0 33.775 0.305 ;
      RECT 1.485 0 17.995 0.305 ;
      RECT 1.485 0 83.25 0.3 ;
      RECT 1.485 8.58 83.25 8.88 ;
      RECT 83.07 8.575 83.25 8.88 ;
      RECT 67.285 8.575 81.12 8.88 ;
      RECT 51.5 8.575 65.335 8.88 ;
      RECT 35.725 8.575 49.55 8.88 ;
      RECT 19.945 8.575 33.775 8.88 ;
      RECT 1.485 8.575 17.995 8.88 ;
      RECT 74.34 6.315 74.51 8.88 ;
      RECT 58.555 6.315 58.725 8.88 ;
      RECT 42.77 6.315 42.94 8.88 ;
      RECT 26.995 6.315 27.165 8.88 ;
      RECT 11.215 6.315 11.385 8.88 ;
      RECT 74.71 6.285 75 6.515 ;
      RECT 58.925 6.285 59.215 6.515 ;
      RECT 43.14 6.285 43.43 6.515 ;
      RECT 27.365 6.285 27.655 6.515 ;
      RECT 11.585 6.285 11.875 6.515 ;
      RECT 74.34 6.315 75 6.485 ;
      RECT 58.555 6.315 59.215 6.485 ;
      RECT 42.77 6.315 43.43 6.485 ;
      RECT 26.995 6.315 27.655 6.485 ;
      RECT 11.215 6.315 11.875 6.485 ;
      RECT 82.645 7.77 82.935 8 ;
      RECT 82.705 6.29 82.875 8 ;
      RECT 82.68 7.275 83.03 7.625 ;
      RECT 82.645 6.29 82.935 6.52 ;
      RECT 82.24 2.395 82.345 2.965 ;
      RECT 82.24 2.73 82.565 2.96 ;
      RECT 82.24 2.76 82.735 2.93 ;
      RECT 82.24 2.395 82.43 2.96 ;
      RECT 81.655 2.36 81.945 2.59 ;
      RECT 81.655 2.395 82.43 2.565 ;
      RECT 81.715 0.88 81.885 2.59 ;
      RECT 81.655 0.88 81.945 1.11 ;
      RECT 81.655 7.77 81.945 8 ;
      RECT 81.715 6.29 81.885 8 ;
      RECT 81.655 6.29 81.945 6.52 ;
      RECT 81.655 6.325 82.51 6.485 ;
      RECT 82.34 5.92 82.51 6.485 ;
      RECT 81.655 6.32 82.05 6.485 ;
      RECT 82.275 5.92 82.565 6.15 ;
      RECT 82.275 5.95 82.735 6.12 ;
      RECT 81.285 2.73 81.575 2.96 ;
      RECT 81.285 2.76 81.745 2.93 ;
      RECT 81.35 1.655 81.515 2.96 ;
      RECT 79.865 1.625 80.155 1.855 ;
      RECT 79.865 1.655 81.515 1.825 ;
      RECT 79.925 0.885 80.095 1.855 ;
      RECT 79.865 0.885 80.155 1.115 ;
      RECT 79.865 7.765 80.155 7.995 ;
      RECT 79.925 7.025 80.095 7.995 ;
      RECT 79.925 7.12 81.515 7.29 ;
      RECT 81.345 5.92 81.515 7.29 ;
      RECT 79.865 7.025 80.155 7.255 ;
      RECT 81.285 5.92 81.575 6.15 ;
      RECT 81.285 5.95 81.745 6.12 ;
      RECT 80.295 1.965 80.645 2.315 ;
      RECT 77.96 2.025 80.645 2.195 ;
      RECT 77.96 1.34 78.13 2.195 ;
      RECT 77.86 1.34 78.21 1.69 ;
      RECT 80.32 6.655 80.645 6.98 ;
      RECT 75.695 6.61 76.045 6.96 ;
      RECT 80.295 6.655 80.645 6.885 ;
      RECT 75.515 6.655 76.045 6.885 ;
      RECT 75.345 6.685 80.645 6.855 ;
      RECT 79.52 2.365 79.84 2.685 ;
      RECT 79.49 2.365 79.84 2.595 ;
      RECT 79.32 2.395 79.84 2.565 ;
      RECT 79.52 6.255 79.84 6.545 ;
      RECT 79.49 6.285 79.84 6.515 ;
      RECT 79.32 6.315 79.84 6.485 ;
      RECT 76.155 2.465 76.34 2.675 ;
      RECT 76.145 2.47 76.355 2.668 ;
      RECT 76.145 2.47 76.441 2.645 ;
      RECT 76.145 2.47 76.5 2.62 ;
      RECT 76.145 2.47 76.555 2.6 ;
      RECT 76.145 2.47 76.565 2.588 ;
      RECT 76.145 2.47 76.76 2.527 ;
      RECT 76.145 2.47 76.79 2.51 ;
      RECT 76.145 2.47 76.81 2.5 ;
      RECT 76.69 2.235 76.95 2.495 ;
      RECT 76.675 2.325 76.69 2.542 ;
      RECT 76.21 2.457 76.95 2.495 ;
      RECT 76.661 2.336 76.675 2.548 ;
      RECT 76.25 2.45 76.95 2.495 ;
      RECT 76.575 2.376 76.661 2.567 ;
      RECT 76.5 2.437 76.95 2.495 ;
      RECT 76.57 2.412 76.575 2.584 ;
      RECT 76.555 2.422 76.95 2.495 ;
      RECT 76.565 2.417 76.57 2.586 ;
      RECT 76.86 2.922 76.865 3.014 ;
      RECT 76.855 2.9 76.86 3.031 ;
      RECT 76.85 2.89 76.855 3.043 ;
      RECT 76.84 2.881 76.85 3.053 ;
      RECT 76.835 2.876 76.84 3.061 ;
      RECT 76.83 2.735 76.835 3.064 ;
      RECT 76.796 2.735 76.83 3.075 ;
      RECT 76.71 2.735 76.796 3.11 ;
      RECT 76.63 2.735 76.71 3.158 ;
      RECT 76.601 2.735 76.63 3.182 ;
      RECT 76.515 2.735 76.601 3.188 ;
      RECT 76.51 2.919 76.515 3.193 ;
      RECT 76.475 2.93 76.51 3.196 ;
      RECT 76.45 2.945 76.475 3.2 ;
      RECT 76.436 2.954 76.45 3.202 ;
      RECT 76.35 2.981 76.436 3.208 ;
      RECT 76.285 3.022 76.35 3.217 ;
      RECT 76.27 3.042 76.285 3.222 ;
      RECT 76.24 3.052 76.27 3.225 ;
      RECT 76.235 3.062 76.24 3.228 ;
      RECT 76.205 3.067 76.235 3.23 ;
      RECT 76.185 3.072 76.205 3.234 ;
      RECT 76.1 3.075 76.185 3.241 ;
      RECT 76.085 3.072 76.1 3.247 ;
      RECT 76.075 3.069 76.085 3.249 ;
      RECT 76.055 3.066 76.075 3.251 ;
      RECT 76.035 3.062 76.055 3.252 ;
      RECT 76.02 3.058 76.035 3.254 ;
      RECT 76.01 3.055 76.02 3.255 ;
      RECT 75.97 3.049 76.01 3.253 ;
      RECT 75.96 3.044 75.97 3.251 ;
      RECT 75.945 3.041 75.96 3.247 ;
      RECT 75.92 3.036 75.945 3.24 ;
      RECT 75.87 3.027 75.92 3.228 ;
      RECT 75.8 3.013 75.87 3.21 ;
      RECT 75.742 2.998 75.8 3.192 ;
      RECT 75.656 2.981 75.742 3.172 ;
      RECT 75.57 2.96 75.656 3.147 ;
      RECT 75.52 2.945 75.57 3.128 ;
      RECT 75.516 2.939 75.52 3.12 ;
      RECT 75.43 2.929 75.516 3.107 ;
      RECT 75.395 2.914 75.43 3.09 ;
      RECT 75.38 2.907 75.395 3.083 ;
      RECT 75.32 2.895 75.38 3.071 ;
      RECT 75.3 2.882 75.32 3.059 ;
      RECT 75.26 2.873 75.3 3.051 ;
      RECT 75.255 2.865 75.26 3.044 ;
      RECT 75.175 2.855 75.255 3.03 ;
      RECT 75.16 2.842 75.175 3.015 ;
      RECT 75.155 2.84 75.16 3.013 ;
      RECT 75.076 2.828 75.155 3 ;
      RECT 74.99 2.803 75.076 2.975 ;
      RECT 74.975 2.772 74.99 2.96 ;
      RECT 74.96 2.747 74.975 2.956 ;
      RECT 74.945 2.74 74.96 2.952 ;
      RECT 74.77 2.745 74.775 2.948 ;
      RECT 74.765 2.75 74.77 2.943 ;
      RECT 74.775 2.74 74.945 2.95 ;
      RECT 75.49 2.5 75.595 2.76 ;
      RECT 76.305 2.025 76.31 2.25 ;
      RECT 76.435 2.025 76.49 2.235 ;
      RECT 76.49 2.03 76.5 2.228 ;
      RECT 76.396 2.025 76.435 2.238 ;
      RECT 76.31 2.025 76.396 2.245 ;
      RECT 76.29 2.03 76.305 2.251 ;
      RECT 76.28 2.07 76.29 2.253 ;
      RECT 76.25 2.08 76.28 2.255 ;
      RECT 76.245 2.085 76.25 2.257 ;
      RECT 76.22 2.09 76.245 2.259 ;
      RECT 76.205 2.095 76.22 2.261 ;
      RECT 76.19 2.097 76.205 2.263 ;
      RECT 76.185 2.102 76.19 2.265 ;
      RECT 76.135 2.11 76.185 2.268 ;
      RECT 76.11 2.119 76.135 2.273 ;
      RECT 76.1 2.126 76.11 2.278 ;
      RECT 76.095 2.129 76.1 2.282 ;
      RECT 76.075 2.132 76.095 2.291 ;
      RECT 76.045 2.14 76.075 2.311 ;
      RECT 76.016 2.153 76.045 2.333 ;
      RECT 75.93 2.187 76.016 2.377 ;
      RECT 75.925 2.213 75.93 2.415 ;
      RECT 75.92 2.217 75.925 2.424 ;
      RECT 75.885 2.23 75.92 2.457 ;
      RECT 75.875 2.244 75.885 2.495 ;
      RECT 75.87 2.248 75.875 2.508 ;
      RECT 75.865 2.252 75.87 2.513 ;
      RECT 75.855 2.26 75.865 2.525 ;
      RECT 75.85 2.267 75.855 2.54 ;
      RECT 75.825 2.28 75.85 2.565 ;
      RECT 75.785 2.309 75.825 2.62 ;
      RECT 75.77 2.334 75.785 2.675 ;
      RECT 75.76 2.345 75.77 2.698 ;
      RECT 75.755 2.352 75.76 2.71 ;
      RECT 75.75 2.356 75.755 2.718 ;
      RECT 75.695 2.384 75.75 2.76 ;
      RECT 75.675 2.42 75.695 2.76 ;
      RECT 75.66 2.435 75.675 2.76 ;
      RECT 75.605 2.467 75.66 2.76 ;
      RECT 75.595 2.497 75.605 2.76 ;
      RECT 75.205 2.112 75.39 2.35 ;
      RECT 75.19 2.114 75.4 2.345 ;
      RECT 75.075 2.06 75.335 2.32 ;
      RECT 75.07 2.097 75.335 2.274 ;
      RECT 75.065 2.107 75.335 2.271 ;
      RECT 75.06 2.147 75.4 2.265 ;
      RECT 75.055 2.18 75.4 2.255 ;
      RECT 75.065 2.122 75.415 2.193 ;
      RECT 75.362 3.22 75.375 3.75 ;
      RECT 75.276 3.22 75.375 3.749 ;
      RECT 75.276 3.22 75.38 3.748 ;
      RECT 75.19 3.22 75.38 3.746 ;
      RECT 75.185 3.22 75.38 3.743 ;
      RECT 75.185 3.22 75.39 3.741 ;
      RECT 75.18 3.512 75.39 3.738 ;
      RECT 75.18 3.522 75.395 3.735 ;
      RECT 75.18 3.59 75.4 3.731 ;
      RECT 75.17 3.595 75.4 3.73 ;
      RECT 75.17 3.687 75.405 3.727 ;
      RECT 75.155 3.22 75.415 3.48 ;
      RECT 75.085 7.765 75.375 7.995 ;
      RECT 75.145 7.025 75.315 7.995 ;
      RECT 75.06 7.055 75.4 7.4 ;
      RECT 75.085 7.025 75.375 7.4 ;
      RECT 74.385 2.21 74.43 3.745 ;
      RECT 74.585 2.21 74.615 2.425 ;
      RECT 72.96 1.95 73.08 2.16 ;
      RECT 72.62 1.9 72.88 2.16 ;
      RECT 72.62 1.945 72.915 2.15 ;
      RECT 74.625 2.226 74.63 2.28 ;
      RECT 74.62 2.219 74.625 2.413 ;
      RECT 74.615 2.213 74.62 2.42 ;
      RECT 74.57 2.21 74.585 2.433 ;
      RECT 74.565 2.21 74.57 2.455 ;
      RECT 74.56 2.21 74.565 2.503 ;
      RECT 74.555 2.21 74.56 2.523 ;
      RECT 74.545 2.21 74.555 2.63 ;
      RECT 74.54 2.21 74.545 2.693 ;
      RECT 74.535 2.21 74.54 2.75 ;
      RECT 74.53 2.21 74.535 2.758 ;
      RECT 74.515 2.21 74.53 2.865 ;
      RECT 74.505 2.21 74.515 3 ;
      RECT 74.495 2.21 74.505 3.11 ;
      RECT 74.485 2.21 74.495 3.167 ;
      RECT 74.48 2.21 74.485 3.207 ;
      RECT 74.475 2.21 74.48 3.243 ;
      RECT 74.465 2.21 74.475 3.283 ;
      RECT 74.46 2.21 74.465 3.325 ;
      RECT 74.44 2.21 74.46 3.39 ;
      RECT 74.445 3.535 74.45 3.715 ;
      RECT 74.44 3.517 74.445 3.723 ;
      RECT 74.435 2.21 74.44 3.453 ;
      RECT 74.435 3.497 74.44 3.73 ;
      RECT 74.43 2.21 74.435 3.74 ;
      RECT 74.375 2.21 74.385 2.51 ;
      RECT 74.38 2.757 74.385 3.745 ;
      RECT 74.375 2.822 74.38 3.745 ;
      RECT 74.37 2.211 74.375 2.5 ;
      RECT 74.365 2.887 74.375 3.745 ;
      RECT 74.36 2.212 74.37 2.49 ;
      RECT 74.35 3 74.365 3.745 ;
      RECT 74.355 2.213 74.36 2.48 ;
      RECT 74.335 2.214 74.355 2.458 ;
      RECT 74.34 3.097 74.35 3.745 ;
      RECT 74.335 3.172 74.34 3.745 ;
      RECT 74.325 2.213 74.335 2.435 ;
      RECT 74.33 3.215 74.335 3.745 ;
      RECT 74.325 3.242 74.33 3.745 ;
      RECT 74.315 2.211 74.325 2.423 ;
      RECT 74.32 3.285 74.325 3.745 ;
      RECT 74.315 3.312 74.32 3.745 ;
      RECT 74.305 2.21 74.315 2.41 ;
      RECT 74.31 3.327 74.315 3.745 ;
      RECT 74.27 3.385 74.31 3.745 ;
      RECT 74.3 2.209 74.305 2.395 ;
      RECT 74.295 2.207 74.3 2.388 ;
      RECT 74.285 2.204 74.295 2.378 ;
      RECT 74.28 2.201 74.285 2.363 ;
      RECT 74.265 2.197 74.28 2.356 ;
      RECT 74.26 3.44 74.27 3.745 ;
      RECT 74.26 2.194 74.265 2.351 ;
      RECT 74.245 2.19 74.26 2.345 ;
      RECT 74.255 3.457 74.26 3.745 ;
      RECT 74.245 3.52 74.255 3.745 ;
      RECT 74.165 2.175 74.245 2.325 ;
      RECT 74.24 3.527 74.245 3.74 ;
      RECT 74.235 3.535 74.24 3.73 ;
      RECT 74.155 2.161 74.165 2.309 ;
      RECT 74.14 2.157 74.155 2.307 ;
      RECT 74.13 2.152 74.14 2.303 ;
      RECT 74.105 2.145 74.13 2.295 ;
      RECT 74.1 2.14 74.105 2.29 ;
      RECT 74.09 2.14 74.1 2.288 ;
      RECT 74.08 2.138 74.09 2.286 ;
      RECT 74.05 2.13 74.08 2.28 ;
      RECT 74.035 2.122 74.05 2.273 ;
      RECT 74.015 2.117 74.035 2.266 ;
      RECT 74.01 2.113 74.015 2.261 ;
      RECT 73.98 2.106 74.01 2.255 ;
      RECT 73.955 2.097 73.98 2.245 ;
      RECT 73.925 2.09 73.955 2.237 ;
      RECT 73.9 2.08 73.925 2.228 ;
      RECT 73.885 2.072 73.9 2.222 ;
      RECT 73.86 2.067 73.885 2.217 ;
      RECT 73.85 2.063 73.86 2.212 ;
      RECT 73.83 2.058 73.85 2.207 ;
      RECT 73.795 2.053 73.83 2.2 ;
      RECT 73.735 2.048 73.795 2.193 ;
      RECT 73.722 2.044 73.735 2.191 ;
      RECT 73.636 2.039 73.722 2.188 ;
      RECT 73.55 2.029 73.636 2.184 ;
      RECT 73.509 2.022 73.55 2.181 ;
      RECT 73.423 2.015 73.509 2.178 ;
      RECT 73.337 2.005 73.423 2.174 ;
      RECT 73.251 1.995 73.337 2.169 ;
      RECT 73.165 1.985 73.251 2.165 ;
      RECT 73.155 1.97 73.165 2.163 ;
      RECT 73.145 1.955 73.155 2.163 ;
      RECT 73.08 1.95 73.145 2.162 ;
      RECT 72.915 1.947 72.96 2.155 ;
      RECT 74.16 2.852 74.165 3.043 ;
      RECT 74.155 2.847 74.16 3.05 ;
      RECT 74.141 2.845 74.155 3.056 ;
      RECT 74.055 2.845 74.141 3.058 ;
      RECT 74.051 2.845 74.055 3.061 ;
      RECT 73.965 2.845 74.051 3.079 ;
      RECT 73.955 2.85 73.965 3.098 ;
      RECT 73.945 2.905 73.955 3.102 ;
      RECT 73.92 2.92 73.945 3.109 ;
      RECT 73.88 2.94 73.92 3.122 ;
      RECT 73.875 2.952 73.88 3.132 ;
      RECT 73.86 2.958 73.875 3.137 ;
      RECT 73.855 2.963 73.86 3.141 ;
      RECT 73.835 2.97 73.855 3.146 ;
      RECT 73.765 2.995 73.835 3.163 ;
      RECT 73.725 3.023 73.765 3.183 ;
      RECT 73.72 3.033 73.725 3.191 ;
      RECT 73.7 3.04 73.72 3.193 ;
      RECT 73.695 3.047 73.7 3.196 ;
      RECT 73.665 3.055 73.695 3.199 ;
      RECT 73.66 3.06 73.665 3.203 ;
      RECT 73.586 3.064 73.66 3.211 ;
      RECT 73.5 3.073 73.586 3.227 ;
      RECT 73.496 3.078 73.5 3.236 ;
      RECT 73.41 3.083 73.496 3.246 ;
      RECT 73.37 3.091 73.41 3.258 ;
      RECT 73.32 3.097 73.37 3.265 ;
      RECT 73.235 3.106 73.32 3.28 ;
      RECT 73.16 3.117 73.235 3.298 ;
      RECT 73.125 3.124 73.16 3.308 ;
      RECT 73.05 3.132 73.125 3.313 ;
      RECT 72.995 3.141 73.05 3.313 ;
      RECT 72.97 3.146 72.995 3.311 ;
      RECT 72.96 3.149 72.97 3.309 ;
      RECT 72.925 3.151 72.96 3.307 ;
      RECT 72.895 3.153 72.925 3.303 ;
      RECT 72.85 3.152 72.895 3.299 ;
      RECT 72.83 3.147 72.85 3.296 ;
      RECT 72.78 3.132 72.83 3.293 ;
      RECT 72.77 3.117 72.78 3.288 ;
      RECT 72.72 3.102 72.77 3.278 ;
      RECT 72.67 3.077 72.72 3.258 ;
      RECT 72.66 3.062 72.67 3.24 ;
      RECT 72.655 3.06 72.66 3.234 ;
      RECT 72.635 3.055 72.655 3.229 ;
      RECT 72.63 3.047 72.635 3.223 ;
      RECT 72.615 3.041 72.63 3.216 ;
      RECT 72.61 3.036 72.615 3.208 ;
      RECT 72.59 3.031 72.61 3.2 ;
      RECT 72.575 3.024 72.59 3.193 ;
      RECT 72.56 3.018 72.575 3.184 ;
      RECT 72.555 3.012 72.56 3.177 ;
      RECT 72.51 2.987 72.555 3.163 ;
      RECT 72.495 2.957 72.51 3.145 ;
      RECT 72.48 2.94 72.495 3.136 ;
      RECT 72.455 2.92 72.48 3.124 ;
      RECT 72.415 2.89 72.455 3.104 ;
      RECT 72.405 2.86 72.415 3.089 ;
      RECT 72.39 2.85 72.405 3.082 ;
      RECT 72.335 2.815 72.39 3.061 ;
      RECT 72.32 2.778 72.335 3.04 ;
      RECT 72.31 2.765 72.32 3.032 ;
      RECT 72.26 2.735 72.31 3.014 ;
      RECT 72.245 2.665 72.26 2.995 ;
      RECT 72.2 2.665 72.245 2.978 ;
      RECT 72.175 2.665 72.2 2.96 ;
      RECT 72.165 2.665 72.175 2.953 ;
      RECT 72.086 2.665 72.165 2.946 ;
      RECT 72 2.665 72.086 2.938 ;
      RECT 71.985 2.697 72 2.933 ;
      RECT 71.91 2.707 71.985 2.929 ;
      RECT 71.89 2.717 71.91 2.924 ;
      RECT 71.865 2.717 71.89 2.921 ;
      RECT 71.855 2.707 71.865 2.92 ;
      RECT 71.845 2.68 71.855 2.919 ;
      RECT 71.805 2.675 71.845 2.917 ;
      RECT 71.76 2.675 71.805 2.913 ;
      RECT 71.735 2.675 71.76 2.908 ;
      RECT 71.685 2.675 71.735 2.895 ;
      RECT 71.645 2.68 71.655 2.88 ;
      RECT 71.655 2.675 71.685 2.885 ;
      RECT 73.64 2.455 73.9 2.715 ;
      RECT 73.635 2.477 73.9 2.673 ;
      RECT 72.875 2.305 73.095 2.67 ;
      RECT 72.857 2.392 73.095 2.669 ;
      RECT 72.84 2.397 73.095 2.666 ;
      RECT 72.84 2.397 73.115 2.665 ;
      RECT 72.81 2.407 73.115 2.663 ;
      RECT 72.805 2.422 73.115 2.659 ;
      RECT 72.805 2.422 73.12 2.658 ;
      RECT 72.8 2.48 73.12 2.656 ;
      RECT 72.8 2.48 73.13 2.653 ;
      RECT 72.795 2.545 73.13 2.648 ;
      RECT 72.875 2.305 73.135 2.565 ;
      RECT 71.62 2.135 71.88 2.395 ;
      RECT 71.62 2.178 71.966 2.369 ;
      RECT 71.62 2.178 72.01 2.368 ;
      RECT 71.62 2.178 72.03 2.366 ;
      RECT 71.62 2.178 72.13 2.365 ;
      RECT 71.62 2.178 72.15 2.363 ;
      RECT 71.62 2.178 72.16 2.358 ;
      RECT 72.03 2.145 72.22 2.355 ;
      RECT 72.03 2.147 72.225 2.353 ;
      RECT 72.02 2.152 72.23 2.345 ;
      RECT 71.966 2.176 72.23 2.345 ;
      RECT 72.01 2.17 72.02 2.367 ;
      RECT 72.02 2.15 72.225 2.353 ;
      RECT 70.975 3.21 71.18 3.44 ;
      RECT 70.915 3.16 70.97 3.42 ;
      RECT 70.975 3.16 71.175 3.44 ;
      RECT 71.945 3.475 71.95 3.502 ;
      RECT 71.935 3.385 71.945 3.507 ;
      RECT 71.93 3.307 71.935 3.513 ;
      RECT 71.92 3.297 71.93 3.52 ;
      RECT 71.915 3.287 71.92 3.526 ;
      RECT 71.905 3.282 71.915 3.528 ;
      RECT 71.89 3.274 71.905 3.536 ;
      RECT 71.875 3.265 71.89 3.548 ;
      RECT 71.865 3.257 71.875 3.558 ;
      RECT 71.83 3.175 71.865 3.576 ;
      RECT 71.795 3.175 71.83 3.595 ;
      RECT 71.78 3.175 71.795 3.603 ;
      RECT 71.725 3.175 71.78 3.603 ;
      RECT 71.691 3.175 71.725 3.594 ;
      RECT 71.605 3.175 71.691 3.57 ;
      RECT 71.595 3.235 71.605 3.552 ;
      RECT 71.555 3.237 71.595 3.543 ;
      RECT 71.55 3.239 71.555 3.533 ;
      RECT 71.53 3.241 71.55 3.528 ;
      RECT 71.52 3.244 71.53 3.523 ;
      RECT 71.51 3.245 71.52 3.518 ;
      RECT 71.486 3.246 71.51 3.51 ;
      RECT 71.4 3.251 71.486 3.488 ;
      RECT 71.345 3.25 71.4 3.461 ;
      RECT 71.33 3.243 71.345 3.448 ;
      RECT 71.295 3.238 71.33 3.444 ;
      RECT 71.24 3.23 71.295 3.443 ;
      RECT 71.18 3.217 71.24 3.441 ;
      RECT 70.97 3.16 70.975 3.428 ;
      RECT 71.045 2.53 71.23 2.74 ;
      RECT 71.035 2.535 71.245 2.733 ;
      RECT 71.075 2.44 71.335 2.7 ;
      RECT 71.03 2.597 71.335 2.623 ;
      RECT 70.375 2.39 70.38 3.19 ;
      RECT 70.32 2.44 70.35 3.19 ;
      RECT 70.31 2.44 70.315 2.75 ;
      RECT 70.295 2.44 70.3 2.745 ;
      RECT 69.84 2.485 69.855 2.7 ;
      RECT 69.77 2.485 69.855 2.695 ;
      RECT 71.035 2.065 71.105 2.275 ;
      RECT 71.105 2.072 71.115 2.27 ;
      RECT 71.001 2.065 71.035 2.282 ;
      RECT 70.915 2.065 71.001 2.306 ;
      RECT 70.905 2.07 70.915 2.325 ;
      RECT 70.9 2.082 70.905 2.328 ;
      RECT 70.885 2.097 70.9 2.332 ;
      RECT 70.88 2.115 70.885 2.336 ;
      RECT 70.84 2.125 70.88 2.345 ;
      RECT 70.825 2.132 70.84 2.357 ;
      RECT 70.81 2.137 70.825 2.362 ;
      RECT 70.795 2.14 70.81 2.367 ;
      RECT 70.785 2.142 70.795 2.371 ;
      RECT 70.75 2.149 70.785 2.379 ;
      RECT 70.715 2.157 70.75 2.393 ;
      RECT 70.705 2.163 70.715 2.402 ;
      RECT 70.7 2.165 70.705 2.404 ;
      RECT 70.68 2.168 70.7 2.41 ;
      RECT 70.65 2.175 70.68 2.421 ;
      RECT 70.64 2.181 70.65 2.428 ;
      RECT 70.615 2.184 70.64 2.435 ;
      RECT 70.605 2.188 70.615 2.443 ;
      RECT 70.6 2.189 70.605 2.465 ;
      RECT 70.595 2.19 70.6 2.48 ;
      RECT 70.59 2.191 70.595 2.495 ;
      RECT 70.585 2.192 70.59 2.51 ;
      RECT 70.58 2.193 70.585 2.54 ;
      RECT 70.57 2.195 70.58 2.573 ;
      RECT 70.555 2.199 70.57 2.62 ;
      RECT 70.545 2.202 70.555 2.665 ;
      RECT 70.54 2.205 70.545 2.693 ;
      RECT 70.53 2.207 70.54 2.72 ;
      RECT 70.525 2.21 70.53 2.755 ;
      RECT 70.495 2.215 70.525 2.813 ;
      RECT 70.49 2.22 70.495 2.898 ;
      RECT 70.485 2.222 70.49 2.933 ;
      RECT 70.48 2.224 70.485 3.015 ;
      RECT 70.475 2.226 70.48 3.103 ;
      RECT 70.465 2.228 70.475 3.185 ;
      RECT 70.45 2.242 70.465 3.19 ;
      RECT 70.415 2.287 70.45 3.19 ;
      RECT 70.405 2.327 70.415 3.19 ;
      RECT 70.39 2.355 70.405 3.19 ;
      RECT 70.385 2.372 70.39 3.19 ;
      RECT 70.38 2.38 70.385 3.19 ;
      RECT 70.37 2.395 70.375 3.19 ;
      RECT 70.365 2.402 70.37 3.19 ;
      RECT 70.355 2.422 70.365 3.19 ;
      RECT 70.35 2.435 70.355 3.19 ;
      RECT 70.315 2.44 70.32 2.775 ;
      RECT 70.3 2.83 70.32 3.19 ;
      RECT 70.3 2.44 70.31 2.748 ;
      RECT 70.295 2.87 70.3 3.19 ;
      RECT 70.245 2.44 70.295 2.743 ;
      RECT 70.29 2.907 70.295 3.19 ;
      RECT 70.28 2.93 70.29 3.19 ;
      RECT 70.275 2.975 70.28 3.19 ;
      RECT 70.265 2.985 70.275 3.183 ;
      RECT 70.191 2.44 70.245 2.737 ;
      RECT 70.105 2.44 70.191 2.73 ;
      RECT 70.056 2.487 70.105 2.723 ;
      RECT 69.97 2.495 70.056 2.716 ;
      RECT 69.955 2.492 69.97 2.711 ;
      RECT 69.941 2.485 69.955 2.71 ;
      RECT 69.855 2.485 69.941 2.705 ;
      RECT 69.76 2.49 69.77 2.69 ;
      RECT 69.35 1.92 69.365 2.32 ;
      RECT 69.545 1.92 69.55 2.18 ;
      RECT 69.29 1.92 69.335 2.18 ;
      RECT 69.745 3.225 69.75 3.43 ;
      RECT 69.74 3.215 69.745 3.435 ;
      RECT 69.735 3.202 69.74 3.44 ;
      RECT 69.73 3.182 69.735 3.44 ;
      RECT 69.705 3.135 69.73 3.44 ;
      RECT 69.67 3.05 69.705 3.44 ;
      RECT 69.665 2.987 69.67 3.44 ;
      RECT 69.66 2.972 69.665 3.44 ;
      RECT 69.645 2.932 69.66 3.44 ;
      RECT 69.64 2.907 69.645 3.44 ;
      RECT 69.63 2.89 69.64 3.44 ;
      RECT 69.595 2.812 69.63 3.44 ;
      RECT 69.59 2.755 69.595 3.44 ;
      RECT 69.585 2.742 69.59 3.44 ;
      RECT 69.575 2.72 69.585 3.44 ;
      RECT 69.565 2.685 69.575 3.44 ;
      RECT 69.555 2.655 69.565 3.44 ;
      RECT 69.545 2.57 69.555 3.083 ;
      RECT 69.552 3.215 69.555 3.44 ;
      RECT 69.55 3.225 69.552 3.44 ;
      RECT 69.54 3.235 69.55 3.435 ;
      RECT 69.535 1.92 69.545 2.315 ;
      RECT 69.54 2.447 69.545 3.058 ;
      RECT 69.535 2.345 69.54 3.041 ;
      RECT 69.525 1.92 69.535 3.017 ;
      RECT 69.52 1.92 69.525 2.988 ;
      RECT 69.515 1.92 69.52 2.978 ;
      RECT 69.495 1.92 69.515 2.94 ;
      RECT 69.49 1.92 69.495 2.898 ;
      RECT 69.485 1.92 69.49 2.878 ;
      RECT 69.455 1.92 69.485 2.828 ;
      RECT 69.445 1.92 69.455 2.775 ;
      RECT 69.44 1.92 69.445 2.748 ;
      RECT 69.435 1.92 69.44 2.733 ;
      RECT 69.425 1.92 69.435 2.71 ;
      RECT 69.415 1.92 69.425 2.685 ;
      RECT 69.41 1.92 69.415 2.625 ;
      RECT 69.4 1.92 69.41 2.563 ;
      RECT 69.395 1.92 69.4 2.483 ;
      RECT 69.39 1.92 69.395 2.448 ;
      RECT 69.385 1.92 69.39 2.423 ;
      RECT 69.38 1.92 69.385 2.408 ;
      RECT 69.375 1.92 69.38 2.378 ;
      RECT 69.37 1.92 69.375 2.355 ;
      RECT 69.365 1.92 69.37 2.328 ;
      RECT 69.335 1.92 69.35 2.315 ;
      RECT 68.49 3.455 68.675 3.665 ;
      RECT 68.48 3.46 68.69 3.658 ;
      RECT 68.48 3.46 68.71 3.63 ;
      RECT 68.48 3.46 68.725 3.609 ;
      RECT 68.48 3.46 68.74 3.607 ;
      RECT 68.48 3.46 68.75 3.606 ;
      RECT 68.48 3.46 68.78 3.603 ;
      RECT 69.13 3.305 69.39 3.565 ;
      RECT 69.09 3.352 69.39 3.548 ;
      RECT 69.081 3.36 69.09 3.551 ;
      RECT 68.675 3.453 69.39 3.548 ;
      RECT 68.995 3.378 69.081 3.558 ;
      RECT 68.69 3.45 69.39 3.548 ;
      RECT 68.936 3.4 68.995 3.57 ;
      RECT 68.71 3.446 69.39 3.548 ;
      RECT 68.85 3.412 68.936 3.581 ;
      RECT 68.725 3.442 69.39 3.548 ;
      RECT 68.795 3.425 68.85 3.593 ;
      RECT 68.74 3.44 69.39 3.548 ;
      RECT 68.78 3.431 68.795 3.599 ;
      RECT 68.75 3.436 69.39 3.548 ;
      RECT 68.895 2.96 69.155 3.22 ;
      RECT 68.895 2.98 69.265 3.19 ;
      RECT 68.895 2.985 69.275 3.185 ;
      RECT 69.086 2.399 69.165 2.63 ;
      RECT 69 2.402 69.215 2.625 ;
      RECT 68.995 2.402 69.215 2.62 ;
      RECT 68.995 2.407 69.225 2.618 ;
      RECT 68.97 2.407 69.225 2.615 ;
      RECT 68.97 2.415 69.235 2.613 ;
      RECT 68.85 2.35 69.11 2.61 ;
      RECT 68.85 2.397 69.16 2.61 ;
      RECT 68.105 2.97 68.11 3.23 ;
      RECT 67.935 2.74 67.94 3.23 ;
      RECT 67.82 2.98 67.825 3.205 ;
      RECT 68.53 2.075 68.535 2.285 ;
      RECT 68.535 2.08 68.55 2.28 ;
      RECT 68.47 2.075 68.53 2.293 ;
      RECT 68.455 2.075 68.47 2.303 ;
      RECT 68.405 2.075 68.455 2.32 ;
      RECT 68.385 2.075 68.405 2.343 ;
      RECT 68.37 2.075 68.385 2.355 ;
      RECT 68.35 2.075 68.37 2.365 ;
      RECT 68.34 2.08 68.35 2.374 ;
      RECT 68.335 2.09 68.34 2.379 ;
      RECT 68.33 2.102 68.335 2.383 ;
      RECT 68.32 2.125 68.33 2.388 ;
      RECT 68.315 2.14 68.32 2.392 ;
      RECT 68.31 2.157 68.315 2.395 ;
      RECT 68.305 2.165 68.31 2.398 ;
      RECT 68.295 2.17 68.305 2.402 ;
      RECT 68.29 2.177 68.295 2.407 ;
      RECT 68.28 2.182 68.29 2.411 ;
      RECT 68.255 2.194 68.28 2.422 ;
      RECT 68.235 2.211 68.255 2.438 ;
      RECT 68.21 2.228 68.235 2.46 ;
      RECT 68.175 2.251 68.21 2.518 ;
      RECT 68.155 2.273 68.175 2.58 ;
      RECT 68.15 2.283 68.155 2.615 ;
      RECT 68.14 2.29 68.15 2.653 ;
      RECT 68.135 2.297 68.14 2.673 ;
      RECT 68.13 2.308 68.135 2.71 ;
      RECT 68.125 2.316 68.13 2.775 ;
      RECT 68.115 2.327 68.125 2.828 ;
      RECT 68.11 2.345 68.115 2.898 ;
      RECT 68.105 2.355 68.11 2.935 ;
      RECT 68.1 2.365 68.105 3.23 ;
      RECT 68.095 2.377 68.1 3.23 ;
      RECT 68.09 2.387 68.095 3.23 ;
      RECT 68.08 2.397 68.09 3.23 ;
      RECT 68.07 2.42 68.08 3.23 ;
      RECT 68.055 2.455 68.07 3.23 ;
      RECT 68.015 2.517 68.055 3.23 ;
      RECT 68.01 2.57 68.015 3.23 ;
      RECT 67.985 2.605 68.01 3.23 ;
      RECT 67.97 2.65 67.985 3.23 ;
      RECT 67.965 2.672 67.97 3.23 ;
      RECT 67.955 2.685 67.965 3.23 ;
      RECT 67.945 2.71 67.955 3.23 ;
      RECT 67.94 2.732 67.945 3.23 ;
      RECT 67.915 2.77 67.935 3.23 ;
      RECT 67.875 2.827 67.915 3.23 ;
      RECT 67.87 2.877 67.875 3.23 ;
      RECT 67.865 2.895 67.87 3.23 ;
      RECT 67.86 2.907 67.865 3.23 ;
      RECT 67.85 2.925 67.86 3.23 ;
      RECT 67.84 2.945 67.85 3.205 ;
      RECT 67.835 2.962 67.84 3.205 ;
      RECT 67.825 2.975 67.835 3.205 ;
      RECT 67.795 2.985 67.82 3.205 ;
      RECT 67.785 2.992 67.795 3.205 ;
      RECT 67.77 3.002 67.785 3.2 ;
      RECT 66.86 7.77 67.15 8 ;
      RECT 66.92 6.29 67.09 8 ;
      RECT 66.87 6.655 67.22 7.005 ;
      RECT 66.86 6.29 67.15 6.52 ;
      RECT 66.455 2.395 66.56 2.965 ;
      RECT 66.455 2.73 66.78 2.96 ;
      RECT 66.455 2.76 66.95 2.93 ;
      RECT 66.455 2.395 66.645 2.96 ;
      RECT 65.87 2.36 66.16 2.59 ;
      RECT 65.87 2.395 66.645 2.565 ;
      RECT 65.93 0.88 66.1 2.59 ;
      RECT 65.87 0.88 66.16 1.11 ;
      RECT 65.87 7.77 66.16 8 ;
      RECT 65.93 6.29 66.1 8 ;
      RECT 65.87 6.29 66.16 6.52 ;
      RECT 65.87 6.325 66.725 6.485 ;
      RECT 66.555 5.92 66.725 6.485 ;
      RECT 65.87 6.32 66.265 6.485 ;
      RECT 66.49 5.92 66.78 6.15 ;
      RECT 66.49 5.95 66.95 6.12 ;
      RECT 65.5 2.73 65.79 2.96 ;
      RECT 65.5 2.76 65.96 2.93 ;
      RECT 65.565 1.655 65.73 2.96 ;
      RECT 64.08 1.625 64.37 1.855 ;
      RECT 64.08 1.655 65.73 1.825 ;
      RECT 64.14 0.885 64.31 1.855 ;
      RECT 64.08 0.885 64.37 1.115 ;
      RECT 64.08 7.765 64.37 7.995 ;
      RECT 64.14 7.025 64.31 7.995 ;
      RECT 64.14 7.12 65.73 7.29 ;
      RECT 65.56 5.92 65.73 7.29 ;
      RECT 64.08 7.025 64.37 7.255 ;
      RECT 65.5 5.92 65.79 6.15 ;
      RECT 65.5 5.95 65.96 6.12 ;
      RECT 64.51 1.965 64.86 2.315 ;
      RECT 62.175 2.025 64.86 2.195 ;
      RECT 62.175 1.34 62.345 2.195 ;
      RECT 62.075 1.34 62.425 1.69 ;
      RECT 64.535 6.655 64.86 6.98 ;
      RECT 59.91 6.61 60.26 6.96 ;
      RECT 64.51 6.655 64.86 6.885 ;
      RECT 59.73 6.655 60.26 6.885 ;
      RECT 59.56 6.685 64.86 6.855 ;
      RECT 63.735 2.365 64.055 2.685 ;
      RECT 63.705 2.365 64.055 2.595 ;
      RECT 63.535 2.395 64.055 2.565 ;
      RECT 63.735 6.255 64.055 6.545 ;
      RECT 63.705 6.285 64.055 6.515 ;
      RECT 63.535 6.315 64.055 6.485 ;
      RECT 60.37 2.465 60.555 2.675 ;
      RECT 60.36 2.47 60.57 2.668 ;
      RECT 60.36 2.47 60.656 2.645 ;
      RECT 60.36 2.47 60.715 2.62 ;
      RECT 60.36 2.47 60.77 2.6 ;
      RECT 60.36 2.47 60.78 2.588 ;
      RECT 60.36 2.47 60.975 2.527 ;
      RECT 60.36 2.47 61.005 2.51 ;
      RECT 60.36 2.47 61.025 2.5 ;
      RECT 60.905 2.235 61.165 2.495 ;
      RECT 60.89 2.325 60.905 2.542 ;
      RECT 60.425 2.457 61.165 2.495 ;
      RECT 60.876 2.336 60.89 2.548 ;
      RECT 60.465 2.45 61.165 2.495 ;
      RECT 60.79 2.376 60.876 2.567 ;
      RECT 60.715 2.437 61.165 2.495 ;
      RECT 60.785 2.412 60.79 2.584 ;
      RECT 60.77 2.422 61.165 2.495 ;
      RECT 60.78 2.417 60.785 2.586 ;
      RECT 61.075 2.922 61.08 3.014 ;
      RECT 61.07 2.9 61.075 3.031 ;
      RECT 61.065 2.89 61.07 3.043 ;
      RECT 61.055 2.881 61.065 3.053 ;
      RECT 61.05 2.876 61.055 3.061 ;
      RECT 61.045 2.735 61.05 3.064 ;
      RECT 61.011 2.735 61.045 3.075 ;
      RECT 60.925 2.735 61.011 3.11 ;
      RECT 60.845 2.735 60.925 3.158 ;
      RECT 60.816 2.735 60.845 3.182 ;
      RECT 60.73 2.735 60.816 3.188 ;
      RECT 60.725 2.919 60.73 3.193 ;
      RECT 60.69 2.93 60.725 3.196 ;
      RECT 60.665 2.945 60.69 3.2 ;
      RECT 60.651 2.954 60.665 3.202 ;
      RECT 60.565 2.981 60.651 3.208 ;
      RECT 60.5 3.022 60.565 3.217 ;
      RECT 60.485 3.042 60.5 3.222 ;
      RECT 60.455 3.052 60.485 3.225 ;
      RECT 60.45 3.062 60.455 3.228 ;
      RECT 60.42 3.067 60.45 3.23 ;
      RECT 60.4 3.072 60.42 3.234 ;
      RECT 60.315 3.075 60.4 3.241 ;
      RECT 60.3 3.072 60.315 3.247 ;
      RECT 60.29 3.069 60.3 3.249 ;
      RECT 60.27 3.066 60.29 3.251 ;
      RECT 60.25 3.062 60.27 3.252 ;
      RECT 60.235 3.058 60.25 3.254 ;
      RECT 60.225 3.055 60.235 3.255 ;
      RECT 60.185 3.049 60.225 3.253 ;
      RECT 60.175 3.044 60.185 3.251 ;
      RECT 60.16 3.041 60.175 3.247 ;
      RECT 60.135 3.036 60.16 3.24 ;
      RECT 60.085 3.027 60.135 3.228 ;
      RECT 60.015 3.013 60.085 3.21 ;
      RECT 59.957 2.998 60.015 3.192 ;
      RECT 59.871 2.981 59.957 3.172 ;
      RECT 59.785 2.96 59.871 3.147 ;
      RECT 59.735 2.945 59.785 3.128 ;
      RECT 59.731 2.939 59.735 3.12 ;
      RECT 59.645 2.929 59.731 3.107 ;
      RECT 59.61 2.914 59.645 3.09 ;
      RECT 59.595 2.907 59.61 3.083 ;
      RECT 59.535 2.895 59.595 3.071 ;
      RECT 59.515 2.882 59.535 3.059 ;
      RECT 59.475 2.873 59.515 3.051 ;
      RECT 59.47 2.865 59.475 3.044 ;
      RECT 59.39 2.855 59.47 3.03 ;
      RECT 59.375 2.842 59.39 3.015 ;
      RECT 59.37 2.84 59.375 3.013 ;
      RECT 59.291 2.828 59.37 3 ;
      RECT 59.205 2.803 59.291 2.975 ;
      RECT 59.19 2.772 59.205 2.96 ;
      RECT 59.175 2.747 59.19 2.956 ;
      RECT 59.16 2.74 59.175 2.952 ;
      RECT 58.985 2.745 58.99 2.948 ;
      RECT 58.98 2.75 58.985 2.943 ;
      RECT 58.99 2.74 59.16 2.95 ;
      RECT 59.705 2.5 59.81 2.76 ;
      RECT 60.52 2.025 60.525 2.25 ;
      RECT 60.65 2.025 60.705 2.235 ;
      RECT 60.705 2.03 60.715 2.228 ;
      RECT 60.611 2.025 60.65 2.238 ;
      RECT 60.525 2.025 60.611 2.245 ;
      RECT 60.505 2.03 60.52 2.251 ;
      RECT 60.495 2.07 60.505 2.253 ;
      RECT 60.465 2.08 60.495 2.255 ;
      RECT 60.46 2.085 60.465 2.257 ;
      RECT 60.435 2.09 60.46 2.259 ;
      RECT 60.42 2.095 60.435 2.261 ;
      RECT 60.405 2.097 60.42 2.263 ;
      RECT 60.4 2.102 60.405 2.265 ;
      RECT 60.35 2.11 60.4 2.268 ;
      RECT 60.325 2.119 60.35 2.273 ;
      RECT 60.315 2.126 60.325 2.278 ;
      RECT 60.31 2.129 60.315 2.282 ;
      RECT 60.29 2.132 60.31 2.291 ;
      RECT 60.26 2.14 60.29 2.311 ;
      RECT 60.231 2.153 60.26 2.333 ;
      RECT 60.145 2.187 60.231 2.377 ;
      RECT 60.14 2.213 60.145 2.415 ;
      RECT 60.135 2.217 60.14 2.424 ;
      RECT 60.1 2.23 60.135 2.457 ;
      RECT 60.09 2.244 60.1 2.495 ;
      RECT 60.085 2.248 60.09 2.508 ;
      RECT 60.08 2.252 60.085 2.513 ;
      RECT 60.07 2.26 60.08 2.525 ;
      RECT 60.065 2.267 60.07 2.54 ;
      RECT 60.04 2.28 60.065 2.565 ;
      RECT 60 2.309 60.04 2.62 ;
      RECT 59.985 2.334 60 2.675 ;
      RECT 59.975 2.345 59.985 2.698 ;
      RECT 59.97 2.352 59.975 2.71 ;
      RECT 59.965 2.356 59.97 2.718 ;
      RECT 59.91 2.384 59.965 2.76 ;
      RECT 59.89 2.42 59.91 2.76 ;
      RECT 59.875 2.435 59.89 2.76 ;
      RECT 59.82 2.467 59.875 2.76 ;
      RECT 59.81 2.497 59.82 2.76 ;
      RECT 59.42 2.112 59.605 2.35 ;
      RECT 59.405 2.114 59.615 2.345 ;
      RECT 59.29 2.06 59.55 2.32 ;
      RECT 59.285 2.097 59.55 2.274 ;
      RECT 59.28 2.107 59.55 2.271 ;
      RECT 59.275 2.147 59.615 2.265 ;
      RECT 59.27 2.18 59.615 2.255 ;
      RECT 59.28 2.122 59.63 2.193 ;
      RECT 59.577 3.22 59.59 3.75 ;
      RECT 59.491 3.22 59.59 3.749 ;
      RECT 59.491 3.22 59.595 3.748 ;
      RECT 59.405 3.22 59.595 3.746 ;
      RECT 59.4 3.22 59.595 3.743 ;
      RECT 59.4 3.22 59.605 3.741 ;
      RECT 59.395 3.512 59.605 3.738 ;
      RECT 59.395 3.522 59.61 3.735 ;
      RECT 59.395 3.59 59.615 3.731 ;
      RECT 59.385 3.595 59.615 3.73 ;
      RECT 59.385 3.687 59.62 3.727 ;
      RECT 59.37 3.22 59.63 3.48 ;
      RECT 59.3 7.765 59.59 7.995 ;
      RECT 59.36 7.025 59.53 7.995 ;
      RECT 59.275 7.055 59.615 7.4 ;
      RECT 59.3 7.025 59.59 7.4 ;
      RECT 58.6 2.21 58.645 3.745 ;
      RECT 58.8 2.21 58.83 2.425 ;
      RECT 57.175 1.95 57.295 2.16 ;
      RECT 56.835 1.9 57.095 2.16 ;
      RECT 56.835 1.945 57.13 2.15 ;
      RECT 58.84 2.226 58.845 2.28 ;
      RECT 58.835 2.219 58.84 2.413 ;
      RECT 58.83 2.213 58.835 2.42 ;
      RECT 58.785 2.21 58.8 2.433 ;
      RECT 58.78 2.21 58.785 2.455 ;
      RECT 58.775 2.21 58.78 2.503 ;
      RECT 58.77 2.21 58.775 2.523 ;
      RECT 58.76 2.21 58.77 2.63 ;
      RECT 58.755 2.21 58.76 2.693 ;
      RECT 58.75 2.21 58.755 2.75 ;
      RECT 58.745 2.21 58.75 2.758 ;
      RECT 58.73 2.21 58.745 2.865 ;
      RECT 58.72 2.21 58.73 3 ;
      RECT 58.71 2.21 58.72 3.11 ;
      RECT 58.7 2.21 58.71 3.167 ;
      RECT 58.695 2.21 58.7 3.207 ;
      RECT 58.69 2.21 58.695 3.243 ;
      RECT 58.68 2.21 58.69 3.283 ;
      RECT 58.675 2.21 58.68 3.325 ;
      RECT 58.655 2.21 58.675 3.39 ;
      RECT 58.66 3.535 58.665 3.715 ;
      RECT 58.655 3.517 58.66 3.723 ;
      RECT 58.65 2.21 58.655 3.453 ;
      RECT 58.65 3.497 58.655 3.73 ;
      RECT 58.645 2.21 58.65 3.74 ;
      RECT 58.59 2.21 58.6 2.51 ;
      RECT 58.595 2.757 58.6 3.745 ;
      RECT 58.59 2.822 58.595 3.745 ;
      RECT 58.585 2.211 58.59 2.5 ;
      RECT 58.58 2.887 58.59 3.745 ;
      RECT 58.575 2.212 58.585 2.49 ;
      RECT 58.565 3 58.58 3.745 ;
      RECT 58.57 2.213 58.575 2.48 ;
      RECT 58.55 2.214 58.57 2.458 ;
      RECT 58.555 3.097 58.565 3.745 ;
      RECT 58.55 3.172 58.555 3.745 ;
      RECT 58.54 2.213 58.55 2.435 ;
      RECT 58.545 3.215 58.55 3.745 ;
      RECT 58.54 3.242 58.545 3.745 ;
      RECT 58.53 2.211 58.54 2.423 ;
      RECT 58.535 3.285 58.54 3.745 ;
      RECT 58.53 3.312 58.535 3.745 ;
      RECT 58.52 2.21 58.53 2.41 ;
      RECT 58.525 3.327 58.53 3.745 ;
      RECT 58.485 3.385 58.525 3.745 ;
      RECT 58.515 2.209 58.52 2.395 ;
      RECT 58.51 2.207 58.515 2.388 ;
      RECT 58.5 2.204 58.51 2.378 ;
      RECT 58.495 2.201 58.5 2.363 ;
      RECT 58.48 2.197 58.495 2.356 ;
      RECT 58.475 3.44 58.485 3.745 ;
      RECT 58.475 2.194 58.48 2.351 ;
      RECT 58.46 2.19 58.475 2.345 ;
      RECT 58.47 3.457 58.475 3.745 ;
      RECT 58.46 3.52 58.47 3.745 ;
      RECT 58.38 2.175 58.46 2.325 ;
      RECT 58.455 3.527 58.46 3.74 ;
      RECT 58.45 3.535 58.455 3.73 ;
      RECT 58.37 2.161 58.38 2.309 ;
      RECT 58.355 2.157 58.37 2.307 ;
      RECT 58.345 2.152 58.355 2.303 ;
      RECT 58.32 2.145 58.345 2.295 ;
      RECT 58.315 2.14 58.32 2.29 ;
      RECT 58.305 2.14 58.315 2.288 ;
      RECT 58.295 2.138 58.305 2.286 ;
      RECT 58.265 2.13 58.295 2.28 ;
      RECT 58.25 2.122 58.265 2.273 ;
      RECT 58.23 2.117 58.25 2.266 ;
      RECT 58.225 2.113 58.23 2.261 ;
      RECT 58.195 2.106 58.225 2.255 ;
      RECT 58.17 2.097 58.195 2.245 ;
      RECT 58.14 2.09 58.17 2.237 ;
      RECT 58.115 2.08 58.14 2.228 ;
      RECT 58.1 2.072 58.115 2.222 ;
      RECT 58.075 2.067 58.1 2.217 ;
      RECT 58.065 2.063 58.075 2.212 ;
      RECT 58.045 2.058 58.065 2.207 ;
      RECT 58.01 2.053 58.045 2.2 ;
      RECT 57.95 2.048 58.01 2.193 ;
      RECT 57.937 2.044 57.95 2.191 ;
      RECT 57.851 2.039 57.937 2.188 ;
      RECT 57.765 2.029 57.851 2.184 ;
      RECT 57.724 2.022 57.765 2.181 ;
      RECT 57.638 2.015 57.724 2.178 ;
      RECT 57.552 2.005 57.638 2.174 ;
      RECT 57.466 1.995 57.552 2.169 ;
      RECT 57.38 1.985 57.466 2.165 ;
      RECT 57.37 1.97 57.38 2.163 ;
      RECT 57.36 1.955 57.37 2.163 ;
      RECT 57.295 1.95 57.36 2.162 ;
      RECT 57.13 1.947 57.175 2.155 ;
      RECT 58.375 2.852 58.38 3.043 ;
      RECT 58.37 2.847 58.375 3.05 ;
      RECT 58.356 2.845 58.37 3.056 ;
      RECT 58.27 2.845 58.356 3.058 ;
      RECT 58.266 2.845 58.27 3.061 ;
      RECT 58.18 2.845 58.266 3.079 ;
      RECT 58.17 2.85 58.18 3.098 ;
      RECT 58.16 2.905 58.17 3.102 ;
      RECT 58.135 2.92 58.16 3.109 ;
      RECT 58.095 2.94 58.135 3.122 ;
      RECT 58.09 2.952 58.095 3.132 ;
      RECT 58.075 2.958 58.09 3.137 ;
      RECT 58.07 2.963 58.075 3.141 ;
      RECT 58.05 2.97 58.07 3.146 ;
      RECT 57.98 2.995 58.05 3.163 ;
      RECT 57.94 3.023 57.98 3.183 ;
      RECT 57.935 3.033 57.94 3.191 ;
      RECT 57.915 3.04 57.935 3.193 ;
      RECT 57.91 3.047 57.915 3.196 ;
      RECT 57.88 3.055 57.91 3.199 ;
      RECT 57.875 3.06 57.88 3.203 ;
      RECT 57.801 3.064 57.875 3.211 ;
      RECT 57.715 3.073 57.801 3.227 ;
      RECT 57.711 3.078 57.715 3.236 ;
      RECT 57.625 3.083 57.711 3.246 ;
      RECT 57.585 3.091 57.625 3.258 ;
      RECT 57.535 3.097 57.585 3.265 ;
      RECT 57.45 3.106 57.535 3.28 ;
      RECT 57.375 3.117 57.45 3.298 ;
      RECT 57.34 3.124 57.375 3.308 ;
      RECT 57.265 3.132 57.34 3.313 ;
      RECT 57.21 3.141 57.265 3.313 ;
      RECT 57.185 3.146 57.21 3.311 ;
      RECT 57.175 3.149 57.185 3.309 ;
      RECT 57.14 3.151 57.175 3.307 ;
      RECT 57.11 3.153 57.14 3.303 ;
      RECT 57.065 3.152 57.11 3.299 ;
      RECT 57.045 3.147 57.065 3.296 ;
      RECT 56.995 3.132 57.045 3.293 ;
      RECT 56.985 3.117 56.995 3.288 ;
      RECT 56.935 3.102 56.985 3.278 ;
      RECT 56.885 3.077 56.935 3.258 ;
      RECT 56.875 3.062 56.885 3.24 ;
      RECT 56.87 3.06 56.875 3.234 ;
      RECT 56.85 3.055 56.87 3.229 ;
      RECT 56.845 3.047 56.85 3.223 ;
      RECT 56.83 3.041 56.845 3.216 ;
      RECT 56.825 3.036 56.83 3.208 ;
      RECT 56.805 3.031 56.825 3.2 ;
      RECT 56.79 3.024 56.805 3.193 ;
      RECT 56.775 3.018 56.79 3.184 ;
      RECT 56.77 3.012 56.775 3.177 ;
      RECT 56.725 2.987 56.77 3.163 ;
      RECT 56.71 2.957 56.725 3.145 ;
      RECT 56.695 2.94 56.71 3.136 ;
      RECT 56.67 2.92 56.695 3.124 ;
      RECT 56.63 2.89 56.67 3.104 ;
      RECT 56.62 2.86 56.63 3.089 ;
      RECT 56.605 2.85 56.62 3.082 ;
      RECT 56.55 2.815 56.605 3.061 ;
      RECT 56.535 2.778 56.55 3.04 ;
      RECT 56.525 2.765 56.535 3.032 ;
      RECT 56.475 2.735 56.525 3.014 ;
      RECT 56.46 2.665 56.475 2.995 ;
      RECT 56.415 2.665 56.46 2.978 ;
      RECT 56.39 2.665 56.415 2.96 ;
      RECT 56.38 2.665 56.39 2.953 ;
      RECT 56.301 2.665 56.38 2.946 ;
      RECT 56.215 2.665 56.301 2.938 ;
      RECT 56.2 2.697 56.215 2.933 ;
      RECT 56.125 2.707 56.2 2.929 ;
      RECT 56.105 2.717 56.125 2.924 ;
      RECT 56.08 2.717 56.105 2.921 ;
      RECT 56.07 2.707 56.08 2.92 ;
      RECT 56.06 2.68 56.07 2.919 ;
      RECT 56.02 2.675 56.06 2.917 ;
      RECT 55.975 2.675 56.02 2.913 ;
      RECT 55.95 2.675 55.975 2.908 ;
      RECT 55.9 2.675 55.95 2.895 ;
      RECT 55.86 2.68 55.87 2.88 ;
      RECT 55.87 2.675 55.9 2.885 ;
      RECT 57.855 2.455 58.115 2.715 ;
      RECT 57.85 2.477 58.115 2.673 ;
      RECT 57.09 2.305 57.31 2.67 ;
      RECT 57.072 2.392 57.31 2.669 ;
      RECT 57.055 2.397 57.31 2.666 ;
      RECT 57.055 2.397 57.33 2.665 ;
      RECT 57.025 2.407 57.33 2.663 ;
      RECT 57.02 2.422 57.33 2.659 ;
      RECT 57.02 2.422 57.335 2.658 ;
      RECT 57.015 2.48 57.335 2.656 ;
      RECT 57.015 2.48 57.345 2.653 ;
      RECT 57.01 2.545 57.345 2.648 ;
      RECT 57.09 2.305 57.35 2.565 ;
      RECT 55.835 2.135 56.095 2.395 ;
      RECT 55.835 2.178 56.181 2.369 ;
      RECT 55.835 2.178 56.225 2.368 ;
      RECT 55.835 2.178 56.245 2.366 ;
      RECT 55.835 2.178 56.345 2.365 ;
      RECT 55.835 2.178 56.365 2.363 ;
      RECT 55.835 2.178 56.375 2.358 ;
      RECT 56.245 2.145 56.435 2.355 ;
      RECT 56.245 2.147 56.44 2.353 ;
      RECT 56.235 2.152 56.445 2.345 ;
      RECT 56.181 2.176 56.445 2.345 ;
      RECT 56.225 2.17 56.235 2.367 ;
      RECT 56.235 2.15 56.44 2.353 ;
      RECT 55.19 3.21 55.395 3.44 ;
      RECT 55.13 3.16 55.185 3.42 ;
      RECT 55.19 3.16 55.39 3.44 ;
      RECT 56.16 3.475 56.165 3.502 ;
      RECT 56.15 3.385 56.16 3.507 ;
      RECT 56.145 3.307 56.15 3.513 ;
      RECT 56.135 3.297 56.145 3.52 ;
      RECT 56.13 3.287 56.135 3.526 ;
      RECT 56.12 3.282 56.13 3.528 ;
      RECT 56.105 3.274 56.12 3.536 ;
      RECT 56.09 3.265 56.105 3.548 ;
      RECT 56.08 3.257 56.09 3.558 ;
      RECT 56.045 3.175 56.08 3.576 ;
      RECT 56.01 3.175 56.045 3.595 ;
      RECT 55.995 3.175 56.01 3.603 ;
      RECT 55.94 3.175 55.995 3.603 ;
      RECT 55.906 3.175 55.94 3.594 ;
      RECT 55.82 3.175 55.906 3.57 ;
      RECT 55.81 3.235 55.82 3.552 ;
      RECT 55.77 3.237 55.81 3.543 ;
      RECT 55.765 3.239 55.77 3.533 ;
      RECT 55.745 3.241 55.765 3.528 ;
      RECT 55.735 3.244 55.745 3.523 ;
      RECT 55.725 3.245 55.735 3.518 ;
      RECT 55.701 3.246 55.725 3.51 ;
      RECT 55.615 3.251 55.701 3.488 ;
      RECT 55.56 3.25 55.615 3.461 ;
      RECT 55.545 3.243 55.56 3.448 ;
      RECT 55.51 3.238 55.545 3.444 ;
      RECT 55.455 3.23 55.51 3.443 ;
      RECT 55.395 3.217 55.455 3.441 ;
      RECT 55.185 3.16 55.19 3.428 ;
      RECT 55.26 2.53 55.445 2.74 ;
      RECT 55.25 2.535 55.46 2.733 ;
      RECT 55.29 2.44 55.55 2.7 ;
      RECT 55.245 2.597 55.55 2.623 ;
      RECT 54.59 2.39 54.595 3.19 ;
      RECT 54.535 2.44 54.565 3.19 ;
      RECT 54.525 2.44 54.53 2.75 ;
      RECT 54.51 2.44 54.515 2.745 ;
      RECT 54.055 2.485 54.07 2.7 ;
      RECT 53.985 2.485 54.07 2.695 ;
      RECT 55.25 2.065 55.32 2.275 ;
      RECT 55.32 2.072 55.33 2.27 ;
      RECT 55.216 2.065 55.25 2.282 ;
      RECT 55.13 2.065 55.216 2.306 ;
      RECT 55.12 2.07 55.13 2.325 ;
      RECT 55.115 2.082 55.12 2.328 ;
      RECT 55.1 2.097 55.115 2.332 ;
      RECT 55.095 2.115 55.1 2.336 ;
      RECT 55.055 2.125 55.095 2.345 ;
      RECT 55.04 2.132 55.055 2.357 ;
      RECT 55.025 2.137 55.04 2.362 ;
      RECT 55.01 2.14 55.025 2.367 ;
      RECT 55 2.142 55.01 2.371 ;
      RECT 54.965 2.149 55 2.379 ;
      RECT 54.93 2.157 54.965 2.393 ;
      RECT 54.92 2.163 54.93 2.402 ;
      RECT 54.915 2.165 54.92 2.404 ;
      RECT 54.895 2.168 54.915 2.41 ;
      RECT 54.865 2.175 54.895 2.421 ;
      RECT 54.855 2.181 54.865 2.428 ;
      RECT 54.83 2.184 54.855 2.435 ;
      RECT 54.82 2.188 54.83 2.443 ;
      RECT 54.815 2.189 54.82 2.465 ;
      RECT 54.81 2.19 54.815 2.48 ;
      RECT 54.805 2.191 54.81 2.495 ;
      RECT 54.8 2.192 54.805 2.51 ;
      RECT 54.795 2.193 54.8 2.54 ;
      RECT 54.785 2.195 54.795 2.573 ;
      RECT 54.77 2.199 54.785 2.62 ;
      RECT 54.76 2.202 54.77 2.665 ;
      RECT 54.755 2.205 54.76 2.693 ;
      RECT 54.745 2.207 54.755 2.72 ;
      RECT 54.74 2.21 54.745 2.755 ;
      RECT 54.71 2.215 54.74 2.813 ;
      RECT 54.705 2.22 54.71 2.898 ;
      RECT 54.7 2.222 54.705 2.933 ;
      RECT 54.695 2.224 54.7 3.015 ;
      RECT 54.69 2.226 54.695 3.103 ;
      RECT 54.68 2.228 54.69 3.185 ;
      RECT 54.665 2.242 54.68 3.19 ;
      RECT 54.63 2.287 54.665 3.19 ;
      RECT 54.62 2.327 54.63 3.19 ;
      RECT 54.605 2.355 54.62 3.19 ;
      RECT 54.6 2.372 54.605 3.19 ;
      RECT 54.595 2.38 54.6 3.19 ;
      RECT 54.585 2.395 54.59 3.19 ;
      RECT 54.58 2.402 54.585 3.19 ;
      RECT 54.57 2.422 54.58 3.19 ;
      RECT 54.565 2.435 54.57 3.19 ;
      RECT 54.53 2.44 54.535 2.775 ;
      RECT 54.515 2.83 54.535 3.19 ;
      RECT 54.515 2.44 54.525 2.748 ;
      RECT 54.51 2.87 54.515 3.19 ;
      RECT 54.46 2.44 54.51 2.743 ;
      RECT 54.505 2.907 54.51 3.19 ;
      RECT 54.495 2.93 54.505 3.19 ;
      RECT 54.49 2.975 54.495 3.19 ;
      RECT 54.48 2.985 54.49 3.183 ;
      RECT 54.406 2.44 54.46 2.737 ;
      RECT 54.32 2.44 54.406 2.73 ;
      RECT 54.271 2.487 54.32 2.723 ;
      RECT 54.185 2.495 54.271 2.716 ;
      RECT 54.17 2.492 54.185 2.711 ;
      RECT 54.156 2.485 54.17 2.71 ;
      RECT 54.07 2.485 54.156 2.705 ;
      RECT 53.975 2.49 53.985 2.69 ;
      RECT 53.565 1.92 53.58 2.32 ;
      RECT 53.76 1.92 53.765 2.18 ;
      RECT 53.505 1.92 53.55 2.18 ;
      RECT 53.96 3.225 53.965 3.43 ;
      RECT 53.955 3.215 53.96 3.435 ;
      RECT 53.95 3.202 53.955 3.44 ;
      RECT 53.945 3.182 53.95 3.44 ;
      RECT 53.92 3.135 53.945 3.44 ;
      RECT 53.885 3.05 53.92 3.44 ;
      RECT 53.88 2.987 53.885 3.44 ;
      RECT 53.875 2.972 53.88 3.44 ;
      RECT 53.86 2.932 53.875 3.44 ;
      RECT 53.855 2.907 53.86 3.44 ;
      RECT 53.845 2.89 53.855 3.44 ;
      RECT 53.81 2.812 53.845 3.44 ;
      RECT 53.805 2.755 53.81 3.44 ;
      RECT 53.8 2.742 53.805 3.44 ;
      RECT 53.79 2.72 53.8 3.44 ;
      RECT 53.78 2.685 53.79 3.44 ;
      RECT 53.77 2.655 53.78 3.44 ;
      RECT 53.76 2.57 53.77 3.083 ;
      RECT 53.767 3.215 53.77 3.44 ;
      RECT 53.765 3.225 53.767 3.44 ;
      RECT 53.755 3.235 53.765 3.435 ;
      RECT 53.75 1.92 53.76 2.315 ;
      RECT 53.755 2.447 53.76 3.058 ;
      RECT 53.75 2.345 53.755 3.041 ;
      RECT 53.74 1.92 53.75 3.017 ;
      RECT 53.735 1.92 53.74 2.988 ;
      RECT 53.73 1.92 53.735 2.978 ;
      RECT 53.71 1.92 53.73 2.94 ;
      RECT 53.705 1.92 53.71 2.898 ;
      RECT 53.7 1.92 53.705 2.878 ;
      RECT 53.67 1.92 53.7 2.828 ;
      RECT 53.66 1.92 53.67 2.775 ;
      RECT 53.655 1.92 53.66 2.748 ;
      RECT 53.65 1.92 53.655 2.733 ;
      RECT 53.64 1.92 53.65 2.71 ;
      RECT 53.63 1.92 53.64 2.685 ;
      RECT 53.625 1.92 53.63 2.625 ;
      RECT 53.615 1.92 53.625 2.563 ;
      RECT 53.61 1.92 53.615 2.483 ;
      RECT 53.605 1.92 53.61 2.448 ;
      RECT 53.6 1.92 53.605 2.423 ;
      RECT 53.595 1.92 53.6 2.408 ;
      RECT 53.59 1.92 53.595 2.378 ;
      RECT 53.585 1.92 53.59 2.355 ;
      RECT 53.58 1.92 53.585 2.328 ;
      RECT 53.55 1.92 53.565 2.315 ;
      RECT 52.705 3.455 52.89 3.665 ;
      RECT 52.695 3.46 52.905 3.658 ;
      RECT 52.695 3.46 52.925 3.63 ;
      RECT 52.695 3.46 52.94 3.609 ;
      RECT 52.695 3.46 52.955 3.607 ;
      RECT 52.695 3.46 52.965 3.606 ;
      RECT 52.695 3.46 52.995 3.603 ;
      RECT 53.345 3.305 53.605 3.565 ;
      RECT 53.305 3.352 53.605 3.548 ;
      RECT 53.296 3.36 53.305 3.551 ;
      RECT 52.89 3.453 53.605 3.548 ;
      RECT 53.21 3.378 53.296 3.558 ;
      RECT 52.905 3.45 53.605 3.548 ;
      RECT 53.151 3.4 53.21 3.57 ;
      RECT 52.925 3.446 53.605 3.548 ;
      RECT 53.065 3.412 53.151 3.581 ;
      RECT 52.94 3.442 53.605 3.548 ;
      RECT 53.01 3.425 53.065 3.593 ;
      RECT 52.955 3.44 53.605 3.548 ;
      RECT 52.995 3.431 53.01 3.599 ;
      RECT 52.965 3.436 53.605 3.548 ;
      RECT 53.11 2.96 53.37 3.22 ;
      RECT 53.11 2.98 53.48 3.19 ;
      RECT 53.11 2.985 53.49 3.185 ;
      RECT 53.301 2.399 53.38 2.63 ;
      RECT 53.215 2.402 53.43 2.625 ;
      RECT 53.21 2.402 53.43 2.62 ;
      RECT 53.21 2.407 53.44 2.618 ;
      RECT 53.185 2.407 53.44 2.615 ;
      RECT 53.185 2.415 53.45 2.613 ;
      RECT 53.065 2.35 53.325 2.61 ;
      RECT 53.065 2.397 53.375 2.61 ;
      RECT 52.32 2.97 52.325 3.23 ;
      RECT 52.15 2.74 52.155 3.23 ;
      RECT 52.035 2.98 52.04 3.205 ;
      RECT 52.745 2.075 52.75 2.285 ;
      RECT 52.75 2.08 52.765 2.28 ;
      RECT 52.685 2.075 52.745 2.293 ;
      RECT 52.67 2.075 52.685 2.303 ;
      RECT 52.62 2.075 52.67 2.32 ;
      RECT 52.6 2.075 52.62 2.343 ;
      RECT 52.585 2.075 52.6 2.355 ;
      RECT 52.565 2.075 52.585 2.365 ;
      RECT 52.555 2.08 52.565 2.374 ;
      RECT 52.55 2.09 52.555 2.379 ;
      RECT 52.545 2.102 52.55 2.383 ;
      RECT 52.535 2.125 52.545 2.388 ;
      RECT 52.53 2.14 52.535 2.392 ;
      RECT 52.525 2.157 52.53 2.395 ;
      RECT 52.52 2.165 52.525 2.398 ;
      RECT 52.51 2.17 52.52 2.402 ;
      RECT 52.505 2.177 52.51 2.407 ;
      RECT 52.495 2.182 52.505 2.411 ;
      RECT 52.47 2.194 52.495 2.422 ;
      RECT 52.45 2.211 52.47 2.438 ;
      RECT 52.425 2.228 52.45 2.46 ;
      RECT 52.39 2.251 52.425 2.518 ;
      RECT 52.37 2.273 52.39 2.58 ;
      RECT 52.365 2.283 52.37 2.615 ;
      RECT 52.355 2.29 52.365 2.653 ;
      RECT 52.35 2.297 52.355 2.673 ;
      RECT 52.345 2.308 52.35 2.71 ;
      RECT 52.34 2.316 52.345 2.775 ;
      RECT 52.33 2.327 52.34 2.828 ;
      RECT 52.325 2.345 52.33 2.898 ;
      RECT 52.32 2.355 52.325 2.935 ;
      RECT 52.315 2.365 52.32 3.23 ;
      RECT 52.31 2.377 52.315 3.23 ;
      RECT 52.305 2.387 52.31 3.23 ;
      RECT 52.295 2.397 52.305 3.23 ;
      RECT 52.285 2.42 52.295 3.23 ;
      RECT 52.27 2.455 52.285 3.23 ;
      RECT 52.23 2.517 52.27 3.23 ;
      RECT 52.225 2.57 52.23 3.23 ;
      RECT 52.2 2.605 52.225 3.23 ;
      RECT 52.185 2.65 52.2 3.23 ;
      RECT 52.18 2.672 52.185 3.23 ;
      RECT 52.17 2.685 52.18 3.23 ;
      RECT 52.16 2.71 52.17 3.23 ;
      RECT 52.155 2.732 52.16 3.23 ;
      RECT 52.13 2.77 52.15 3.23 ;
      RECT 52.09 2.827 52.13 3.23 ;
      RECT 52.085 2.877 52.09 3.23 ;
      RECT 52.08 2.895 52.085 3.23 ;
      RECT 52.075 2.907 52.08 3.23 ;
      RECT 52.065 2.925 52.075 3.23 ;
      RECT 52.055 2.945 52.065 3.205 ;
      RECT 52.05 2.962 52.055 3.205 ;
      RECT 52.04 2.975 52.05 3.205 ;
      RECT 52.01 2.985 52.035 3.205 ;
      RECT 52 2.992 52.01 3.205 ;
      RECT 51.985 3.002 52 3.2 ;
      RECT 51.075 7.77 51.365 8 ;
      RECT 51.135 6.29 51.305 8 ;
      RECT 51.085 6.655 51.435 7.005 ;
      RECT 51.075 6.29 51.365 6.52 ;
      RECT 50.67 2.395 50.775 2.965 ;
      RECT 50.67 2.73 50.995 2.96 ;
      RECT 50.67 2.76 51.165 2.93 ;
      RECT 50.67 2.395 50.86 2.96 ;
      RECT 50.085 2.36 50.375 2.59 ;
      RECT 50.085 2.395 50.86 2.565 ;
      RECT 50.145 0.88 50.315 2.59 ;
      RECT 50.085 0.88 50.375 1.11 ;
      RECT 50.085 7.77 50.375 8 ;
      RECT 50.145 6.29 50.315 8 ;
      RECT 50.085 6.29 50.375 6.52 ;
      RECT 50.085 6.325 50.94 6.485 ;
      RECT 50.77 5.92 50.94 6.485 ;
      RECT 50.085 6.32 50.48 6.485 ;
      RECT 50.705 5.92 50.995 6.15 ;
      RECT 50.705 5.95 51.165 6.12 ;
      RECT 49.715 2.73 50.005 2.96 ;
      RECT 49.715 2.76 50.175 2.93 ;
      RECT 49.78 1.655 49.945 2.96 ;
      RECT 48.295 1.625 48.585 1.855 ;
      RECT 48.295 1.655 49.945 1.825 ;
      RECT 48.355 0.885 48.525 1.855 ;
      RECT 48.295 0.885 48.585 1.115 ;
      RECT 48.295 7.765 48.585 7.995 ;
      RECT 48.355 7.025 48.525 7.995 ;
      RECT 48.355 7.12 49.945 7.29 ;
      RECT 49.775 5.92 49.945 7.29 ;
      RECT 48.295 7.025 48.585 7.255 ;
      RECT 49.715 5.92 50.005 6.15 ;
      RECT 49.715 5.95 50.175 6.12 ;
      RECT 48.725 1.965 49.075 2.315 ;
      RECT 46.39 2.025 49.075 2.195 ;
      RECT 46.39 1.34 46.56 2.195 ;
      RECT 46.29 1.34 46.64 1.69 ;
      RECT 48.75 6.655 49.075 6.98 ;
      RECT 44.18 6.615 44.53 6.965 ;
      RECT 48.725 6.655 49.075 6.885 ;
      RECT 43.945 6.655 44.53 6.885 ;
      RECT 43.775 6.685 49.075 6.855 ;
      RECT 47.95 2.365 48.27 2.685 ;
      RECT 47.92 2.365 48.27 2.595 ;
      RECT 47.75 2.395 48.27 2.565 ;
      RECT 47.95 6.255 48.27 6.545 ;
      RECT 47.92 6.285 48.27 6.515 ;
      RECT 47.75 6.315 48.27 6.485 ;
      RECT 44.585 2.465 44.77 2.675 ;
      RECT 44.575 2.47 44.785 2.668 ;
      RECT 44.575 2.47 44.871 2.645 ;
      RECT 44.575 2.47 44.93 2.62 ;
      RECT 44.575 2.47 44.985 2.6 ;
      RECT 44.575 2.47 44.995 2.588 ;
      RECT 44.575 2.47 45.19 2.527 ;
      RECT 44.575 2.47 45.22 2.51 ;
      RECT 44.575 2.47 45.24 2.5 ;
      RECT 45.12 2.235 45.38 2.495 ;
      RECT 45.105 2.325 45.12 2.542 ;
      RECT 44.64 2.457 45.38 2.495 ;
      RECT 45.091 2.336 45.105 2.548 ;
      RECT 44.68 2.45 45.38 2.495 ;
      RECT 45.005 2.376 45.091 2.567 ;
      RECT 44.93 2.437 45.38 2.495 ;
      RECT 45 2.412 45.005 2.584 ;
      RECT 44.985 2.422 45.38 2.495 ;
      RECT 44.995 2.417 45 2.586 ;
      RECT 45.29 2.922 45.295 3.014 ;
      RECT 45.285 2.9 45.29 3.031 ;
      RECT 45.28 2.89 45.285 3.043 ;
      RECT 45.27 2.881 45.28 3.053 ;
      RECT 45.265 2.876 45.27 3.061 ;
      RECT 45.26 2.735 45.265 3.064 ;
      RECT 45.226 2.735 45.26 3.075 ;
      RECT 45.14 2.735 45.226 3.11 ;
      RECT 45.06 2.735 45.14 3.158 ;
      RECT 45.031 2.735 45.06 3.182 ;
      RECT 44.945 2.735 45.031 3.188 ;
      RECT 44.94 2.919 44.945 3.193 ;
      RECT 44.905 2.93 44.94 3.196 ;
      RECT 44.88 2.945 44.905 3.2 ;
      RECT 44.866 2.954 44.88 3.202 ;
      RECT 44.78 2.981 44.866 3.208 ;
      RECT 44.715 3.022 44.78 3.217 ;
      RECT 44.7 3.042 44.715 3.222 ;
      RECT 44.67 3.052 44.7 3.225 ;
      RECT 44.665 3.062 44.67 3.228 ;
      RECT 44.635 3.067 44.665 3.23 ;
      RECT 44.615 3.072 44.635 3.234 ;
      RECT 44.53 3.075 44.615 3.241 ;
      RECT 44.515 3.072 44.53 3.247 ;
      RECT 44.505 3.069 44.515 3.249 ;
      RECT 44.485 3.066 44.505 3.251 ;
      RECT 44.465 3.062 44.485 3.252 ;
      RECT 44.45 3.058 44.465 3.254 ;
      RECT 44.44 3.055 44.45 3.255 ;
      RECT 44.4 3.049 44.44 3.253 ;
      RECT 44.39 3.044 44.4 3.251 ;
      RECT 44.375 3.041 44.39 3.247 ;
      RECT 44.35 3.036 44.375 3.24 ;
      RECT 44.3 3.027 44.35 3.228 ;
      RECT 44.23 3.013 44.3 3.21 ;
      RECT 44.172 2.998 44.23 3.192 ;
      RECT 44.086 2.981 44.172 3.172 ;
      RECT 44 2.96 44.086 3.147 ;
      RECT 43.95 2.945 44 3.128 ;
      RECT 43.946 2.939 43.95 3.12 ;
      RECT 43.86 2.929 43.946 3.107 ;
      RECT 43.825 2.914 43.86 3.09 ;
      RECT 43.81 2.907 43.825 3.083 ;
      RECT 43.75 2.895 43.81 3.071 ;
      RECT 43.73 2.882 43.75 3.059 ;
      RECT 43.69 2.873 43.73 3.051 ;
      RECT 43.685 2.865 43.69 3.044 ;
      RECT 43.605 2.855 43.685 3.03 ;
      RECT 43.59 2.842 43.605 3.015 ;
      RECT 43.585 2.84 43.59 3.013 ;
      RECT 43.506 2.828 43.585 3 ;
      RECT 43.42 2.803 43.506 2.975 ;
      RECT 43.405 2.772 43.42 2.96 ;
      RECT 43.39 2.747 43.405 2.956 ;
      RECT 43.375 2.74 43.39 2.952 ;
      RECT 43.2 2.745 43.205 2.948 ;
      RECT 43.195 2.75 43.2 2.943 ;
      RECT 43.205 2.74 43.375 2.95 ;
      RECT 43.92 2.5 44.025 2.76 ;
      RECT 44.735 2.025 44.74 2.25 ;
      RECT 44.865 2.025 44.92 2.235 ;
      RECT 44.92 2.03 44.93 2.228 ;
      RECT 44.826 2.025 44.865 2.238 ;
      RECT 44.74 2.025 44.826 2.245 ;
      RECT 44.72 2.03 44.735 2.251 ;
      RECT 44.71 2.07 44.72 2.253 ;
      RECT 44.68 2.08 44.71 2.255 ;
      RECT 44.675 2.085 44.68 2.257 ;
      RECT 44.65 2.09 44.675 2.259 ;
      RECT 44.635 2.095 44.65 2.261 ;
      RECT 44.62 2.097 44.635 2.263 ;
      RECT 44.615 2.102 44.62 2.265 ;
      RECT 44.565 2.11 44.615 2.268 ;
      RECT 44.54 2.119 44.565 2.273 ;
      RECT 44.53 2.126 44.54 2.278 ;
      RECT 44.525 2.129 44.53 2.282 ;
      RECT 44.505 2.132 44.525 2.291 ;
      RECT 44.475 2.14 44.505 2.311 ;
      RECT 44.446 2.153 44.475 2.333 ;
      RECT 44.36 2.187 44.446 2.377 ;
      RECT 44.355 2.213 44.36 2.415 ;
      RECT 44.35 2.217 44.355 2.424 ;
      RECT 44.315 2.23 44.35 2.457 ;
      RECT 44.305 2.244 44.315 2.495 ;
      RECT 44.3 2.248 44.305 2.508 ;
      RECT 44.295 2.252 44.3 2.513 ;
      RECT 44.285 2.26 44.295 2.525 ;
      RECT 44.28 2.267 44.285 2.54 ;
      RECT 44.255 2.28 44.28 2.565 ;
      RECT 44.215 2.309 44.255 2.62 ;
      RECT 44.2 2.334 44.215 2.675 ;
      RECT 44.19 2.345 44.2 2.698 ;
      RECT 44.185 2.352 44.19 2.71 ;
      RECT 44.18 2.356 44.185 2.718 ;
      RECT 44.125 2.384 44.18 2.76 ;
      RECT 44.105 2.42 44.125 2.76 ;
      RECT 44.09 2.435 44.105 2.76 ;
      RECT 44.035 2.467 44.09 2.76 ;
      RECT 44.025 2.497 44.035 2.76 ;
      RECT 43.635 2.112 43.82 2.35 ;
      RECT 43.62 2.114 43.83 2.345 ;
      RECT 43.505 2.06 43.765 2.32 ;
      RECT 43.5 2.097 43.765 2.274 ;
      RECT 43.495 2.107 43.765 2.271 ;
      RECT 43.49 2.147 43.83 2.265 ;
      RECT 43.485 2.18 43.83 2.255 ;
      RECT 43.495 2.122 43.845 2.193 ;
      RECT 43.792 3.22 43.805 3.75 ;
      RECT 43.706 3.22 43.805 3.749 ;
      RECT 43.706 3.22 43.81 3.748 ;
      RECT 43.62 3.22 43.81 3.746 ;
      RECT 43.615 3.22 43.81 3.743 ;
      RECT 43.615 3.22 43.82 3.741 ;
      RECT 43.61 3.512 43.82 3.738 ;
      RECT 43.61 3.522 43.825 3.735 ;
      RECT 43.61 3.59 43.83 3.731 ;
      RECT 43.6 3.595 43.83 3.73 ;
      RECT 43.6 3.687 43.835 3.727 ;
      RECT 43.585 3.22 43.845 3.48 ;
      RECT 43.515 7.765 43.805 7.995 ;
      RECT 43.575 7.025 43.745 7.995 ;
      RECT 43.49 7.055 43.83 7.4 ;
      RECT 43.515 7.025 43.805 7.4 ;
      RECT 42.815 2.21 42.86 3.745 ;
      RECT 43.015 2.21 43.045 2.425 ;
      RECT 41.39 1.95 41.51 2.16 ;
      RECT 41.05 1.9 41.31 2.16 ;
      RECT 41.05 1.945 41.345 2.15 ;
      RECT 43.055 2.226 43.06 2.28 ;
      RECT 43.05 2.219 43.055 2.413 ;
      RECT 43.045 2.213 43.05 2.42 ;
      RECT 43 2.21 43.015 2.433 ;
      RECT 42.995 2.21 43 2.455 ;
      RECT 42.99 2.21 42.995 2.503 ;
      RECT 42.985 2.21 42.99 2.523 ;
      RECT 42.975 2.21 42.985 2.63 ;
      RECT 42.97 2.21 42.975 2.693 ;
      RECT 42.965 2.21 42.97 2.75 ;
      RECT 42.96 2.21 42.965 2.758 ;
      RECT 42.945 2.21 42.96 2.865 ;
      RECT 42.935 2.21 42.945 3 ;
      RECT 42.925 2.21 42.935 3.11 ;
      RECT 42.915 2.21 42.925 3.167 ;
      RECT 42.91 2.21 42.915 3.207 ;
      RECT 42.905 2.21 42.91 3.243 ;
      RECT 42.895 2.21 42.905 3.283 ;
      RECT 42.89 2.21 42.895 3.325 ;
      RECT 42.87 2.21 42.89 3.39 ;
      RECT 42.875 3.535 42.88 3.715 ;
      RECT 42.87 3.517 42.875 3.723 ;
      RECT 42.865 2.21 42.87 3.453 ;
      RECT 42.865 3.497 42.87 3.73 ;
      RECT 42.86 2.21 42.865 3.74 ;
      RECT 42.805 2.21 42.815 2.51 ;
      RECT 42.81 2.757 42.815 3.745 ;
      RECT 42.805 2.822 42.81 3.745 ;
      RECT 42.8 2.211 42.805 2.5 ;
      RECT 42.795 2.887 42.805 3.745 ;
      RECT 42.79 2.212 42.8 2.49 ;
      RECT 42.78 3 42.795 3.745 ;
      RECT 42.785 2.213 42.79 2.48 ;
      RECT 42.765 2.214 42.785 2.458 ;
      RECT 42.77 3.097 42.78 3.745 ;
      RECT 42.765 3.172 42.77 3.745 ;
      RECT 42.755 2.213 42.765 2.435 ;
      RECT 42.76 3.215 42.765 3.745 ;
      RECT 42.755 3.242 42.76 3.745 ;
      RECT 42.745 2.211 42.755 2.423 ;
      RECT 42.75 3.285 42.755 3.745 ;
      RECT 42.745 3.312 42.75 3.745 ;
      RECT 42.735 2.21 42.745 2.41 ;
      RECT 42.74 3.327 42.745 3.745 ;
      RECT 42.7 3.385 42.74 3.745 ;
      RECT 42.73 2.209 42.735 2.395 ;
      RECT 42.725 2.207 42.73 2.388 ;
      RECT 42.715 2.204 42.725 2.378 ;
      RECT 42.71 2.201 42.715 2.363 ;
      RECT 42.695 2.197 42.71 2.356 ;
      RECT 42.69 3.44 42.7 3.745 ;
      RECT 42.69 2.194 42.695 2.351 ;
      RECT 42.675 2.19 42.69 2.345 ;
      RECT 42.685 3.457 42.69 3.745 ;
      RECT 42.675 3.52 42.685 3.745 ;
      RECT 42.595 2.175 42.675 2.325 ;
      RECT 42.67 3.527 42.675 3.74 ;
      RECT 42.665 3.535 42.67 3.73 ;
      RECT 42.585 2.161 42.595 2.309 ;
      RECT 42.57 2.157 42.585 2.307 ;
      RECT 42.56 2.152 42.57 2.303 ;
      RECT 42.535 2.145 42.56 2.295 ;
      RECT 42.53 2.14 42.535 2.29 ;
      RECT 42.52 2.14 42.53 2.288 ;
      RECT 42.51 2.138 42.52 2.286 ;
      RECT 42.48 2.13 42.51 2.28 ;
      RECT 42.465 2.122 42.48 2.273 ;
      RECT 42.445 2.117 42.465 2.266 ;
      RECT 42.44 2.113 42.445 2.261 ;
      RECT 42.41 2.106 42.44 2.255 ;
      RECT 42.385 2.097 42.41 2.245 ;
      RECT 42.355 2.09 42.385 2.237 ;
      RECT 42.33 2.08 42.355 2.228 ;
      RECT 42.315 2.072 42.33 2.222 ;
      RECT 42.29 2.067 42.315 2.217 ;
      RECT 42.28 2.063 42.29 2.212 ;
      RECT 42.26 2.058 42.28 2.207 ;
      RECT 42.225 2.053 42.26 2.2 ;
      RECT 42.165 2.048 42.225 2.193 ;
      RECT 42.152 2.044 42.165 2.191 ;
      RECT 42.066 2.039 42.152 2.188 ;
      RECT 41.98 2.029 42.066 2.184 ;
      RECT 41.939 2.022 41.98 2.181 ;
      RECT 41.853 2.015 41.939 2.178 ;
      RECT 41.767 2.005 41.853 2.174 ;
      RECT 41.681 1.995 41.767 2.169 ;
      RECT 41.595 1.985 41.681 2.165 ;
      RECT 41.585 1.97 41.595 2.163 ;
      RECT 41.575 1.955 41.585 2.163 ;
      RECT 41.51 1.95 41.575 2.162 ;
      RECT 41.345 1.947 41.39 2.155 ;
      RECT 42.59 2.852 42.595 3.043 ;
      RECT 42.585 2.847 42.59 3.05 ;
      RECT 42.571 2.845 42.585 3.056 ;
      RECT 42.485 2.845 42.571 3.058 ;
      RECT 42.481 2.845 42.485 3.061 ;
      RECT 42.395 2.845 42.481 3.079 ;
      RECT 42.385 2.85 42.395 3.098 ;
      RECT 42.375 2.905 42.385 3.102 ;
      RECT 42.35 2.92 42.375 3.109 ;
      RECT 42.31 2.94 42.35 3.122 ;
      RECT 42.305 2.952 42.31 3.132 ;
      RECT 42.29 2.958 42.305 3.137 ;
      RECT 42.285 2.963 42.29 3.141 ;
      RECT 42.265 2.97 42.285 3.146 ;
      RECT 42.195 2.995 42.265 3.163 ;
      RECT 42.155 3.023 42.195 3.183 ;
      RECT 42.15 3.033 42.155 3.191 ;
      RECT 42.13 3.04 42.15 3.193 ;
      RECT 42.125 3.047 42.13 3.196 ;
      RECT 42.095 3.055 42.125 3.199 ;
      RECT 42.09 3.06 42.095 3.203 ;
      RECT 42.016 3.064 42.09 3.211 ;
      RECT 41.93 3.073 42.016 3.227 ;
      RECT 41.926 3.078 41.93 3.236 ;
      RECT 41.84 3.083 41.926 3.246 ;
      RECT 41.8 3.091 41.84 3.258 ;
      RECT 41.75 3.097 41.8 3.265 ;
      RECT 41.665 3.106 41.75 3.28 ;
      RECT 41.59 3.117 41.665 3.298 ;
      RECT 41.555 3.124 41.59 3.308 ;
      RECT 41.48 3.132 41.555 3.313 ;
      RECT 41.425 3.141 41.48 3.313 ;
      RECT 41.4 3.146 41.425 3.311 ;
      RECT 41.39 3.149 41.4 3.309 ;
      RECT 41.355 3.151 41.39 3.307 ;
      RECT 41.325 3.153 41.355 3.303 ;
      RECT 41.28 3.152 41.325 3.299 ;
      RECT 41.26 3.147 41.28 3.296 ;
      RECT 41.21 3.132 41.26 3.293 ;
      RECT 41.2 3.117 41.21 3.288 ;
      RECT 41.15 3.102 41.2 3.278 ;
      RECT 41.1 3.077 41.15 3.258 ;
      RECT 41.09 3.062 41.1 3.24 ;
      RECT 41.085 3.06 41.09 3.234 ;
      RECT 41.065 3.055 41.085 3.229 ;
      RECT 41.06 3.047 41.065 3.223 ;
      RECT 41.045 3.041 41.06 3.216 ;
      RECT 41.04 3.036 41.045 3.208 ;
      RECT 41.02 3.031 41.04 3.2 ;
      RECT 41.005 3.024 41.02 3.193 ;
      RECT 40.99 3.018 41.005 3.184 ;
      RECT 40.985 3.012 40.99 3.177 ;
      RECT 40.94 2.987 40.985 3.163 ;
      RECT 40.925 2.957 40.94 3.145 ;
      RECT 40.91 2.94 40.925 3.136 ;
      RECT 40.885 2.92 40.91 3.124 ;
      RECT 40.845 2.89 40.885 3.104 ;
      RECT 40.835 2.86 40.845 3.089 ;
      RECT 40.82 2.85 40.835 3.082 ;
      RECT 40.765 2.815 40.82 3.061 ;
      RECT 40.75 2.778 40.765 3.04 ;
      RECT 40.74 2.765 40.75 3.032 ;
      RECT 40.69 2.735 40.74 3.014 ;
      RECT 40.675 2.665 40.69 2.995 ;
      RECT 40.63 2.665 40.675 2.978 ;
      RECT 40.605 2.665 40.63 2.96 ;
      RECT 40.595 2.665 40.605 2.953 ;
      RECT 40.516 2.665 40.595 2.946 ;
      RECT 40.43 2.665 40.516 2.938 ;
      RECT 40.415 2.697 40.43 2.933 ;
      RECT 40.34 2.707 40.415 2.929 ;
      RECT 40.32 2.717 40.34 2.924 ;
      RECT 40.295 2.717 40.32 2.921 ;
      RECT 40.285 2.707 40.295 2.92 ;
      RECT 40.275 2.68 40.285 2.919 ;
      RECT 40.235 2.675 40.275 2.917 ;
      RECT 40.19 2.675 40.235 2.913 ;
      RECT 40.165 2.675 40.19 2.908 ;
      RECT 40.115 2.675 40.165 2.895 ;
      RECT 40.075 2.68 40.085 2.88 ;
      RECT 40.085 2.675 40.115 2.885 ;
      RECT 42.07 2.455 42.33 2.715 ;
      RECT 42.065 2.477 42.33 2.673 ;
      RECT 41.305 2.305 41.525 2.67 ;
      RECT 41.287 2.392 41.525 2.669 ;
      RECT 41.27 2.397 41.525 2.666 ;
      RECT 41.27 2.397 41.545 2.665 ;
      RECT 41.24 2.407 41.545 2.663 ;
      RECT 41.235 2.422 41.545 2.659 ;
      RECT 41.235 2.422 41.55 2.658 ;
      RECT 41.23 2.48 41.55 2.656 ;
      RECT 41.23 2.48 41.56 2.653 ;
      RECT 41.225 2.545 41.56 2.648 ;
      RECT 41.305 2.305 41.565 2.565 ;
      RECT 40.05 2.135 40.31 2.395 ;
      RECT 40.05 2.178 40.396 2.369 ;
      RECT 40.05 2.178 40.44 2.368 ;
      RECT 40.05 2.178 40.46 2.366 ;
      RECT 40.05 2.178 40.56 2.365 ;
      RECT 40.05 2.178 40.58 2.363 ;
      RECT 40.05 2.178 40.59 2.358 ;
      RECT 40.46 2.145 40.65 2.355 ;
      RECT 40.46 2.147 40.655 2.353 ;
      RECT 40.45 2.152 40.66 2.345 ;
      RECT 40.396 2.176 40.66 2.345 ;
      RECT 40.44 2.17 40.45 2.367 ;
      RECT 40.45 2.15 40.655 2.353 ;
      RECT 39.405 3.21 39.61 3.44 ;
      RECT 39.345 3.16 39.4 3.42 ;
      RECT 39.405 3.16 39.605 3.44 ;
      RECT 40.375 3.475 40.38 3.502 ;
      RECT 40.365 3.385 40.375 3.507 ;
      RECT 40.36 3.307 40.365 3.513 ;
      RECT 40.35 3.297 40.36 3.52 ;
      RECT 40.345 3.287 40.35 3.526 ;
      RECT 40.335 3.282 40.345 3.528 ;
      RECT 40.32 3.274 40.335 3.536 ;
      RECT 40.305 3.265 40.32 3.548 ;
      RECT 40.295 3.257 40.305 3.558 ;
      RECT 40.26 3.175 40.295 3.576 ;
      RECT 40.225 3.175 40.26 3.595 ;
      RECT 40.21 3.175 40.225 3.603 ;
      RECT 40.155 3.175 40.21 3.603 ;
      RECT 40.121 3.175 40.155 3.594 ;
      RECT 40.035 3.175 40.121 3.57 ;
      RECT 40.025 3.235 40.035 3.552 ;
      RECT 39.985 3.237 40.025 3.543 ;
      RECT 39.98 3.239 39.985 3.533 ;
      RECT 39.96 3.241 39.98 3.528 ;
      RECT 39.95 3.244 39.96 3.523 ;
      RECT 39.94 3.245 39.95 3.518 ;
      RECT 39.916 3.246 39.94 3.51 ;
      RECT 39.83 3.251 39.916 3.488 ;
      RECT 39.775 3.25 39.83 3.461 ;
      RECT 39.76 3.243 39.775 3.448 ;
      RECT 39.725 3.238 39.76 3.444 ;
      RECT 39.67 3.23 39.725 3.443 ;
      RECT 39.61 3.217 39.67 3.441 ;
      RECT 39.4 3.16 39.405 3.428 ;
      RECT 39.475 2.53 39.66 2.74 ;
      RECT 39.465 2.535 39.675 2.733 ;
      RECT 39.505 2.44 39.765 2.7 ;
      RECT 39.46 2.597 39.765 2.623 ;
      RECT 38.805 2.39 38.81 3.19 ;
      RECT 38.75 2.44 38.78 3.19 ;
      RECT 38.74 2.44 38.745 2.75 ;
      RECT 38.725 2.44 38.73 2.745 ;
      RECT 38.27 2.485 38.285 2.7 ;
      RECT 38.2 2.485 38.285 2.695 ;
      RECT 39.465 2.065 39.535 2.275 ;
      RECT 39.535 2.072 39.545 2.27 ;
      RECT 39.431 2.065 39.465 2.282 ;
      RECT 39.345 2.065 39.431 2.306 ;
      RECT 39.335 2.07 39.345 2.325 ;
      RECT 39.33 2.082 39.335 2.328 ;
      RECT 39.315 2.097 39.33 2.332 ;
      RECT 39.31 2.115 39.315 2.336 ;
      RECT 39.27 2.125 39.31 2.345 ;
      RECT 39.255 2.132 39.27 2.357 ;
      RECT 39.24 2.137 39.255 2.362 ;
      RECT 39.225 2.14 39.24 2.367 ;
      RECT 39.215 2.142 39.225 2.371 ;
      RECT 39.18 2.149 39.215 2.379 ;
      RECT 39.145 2.157 39.18 2.393 ;
      RECT 39.135 2.163 39.145 2.402 ;
      RECT 39.13 2.165 39.135 2.404 ;
      RECT 39.11 2.168 39.13 2.41 ;
      RECT 39.08 2.175 39.11 2.421 ;
      RECT 39.07 2.181 39.08 2.428 ;
      RECT 39.045 2.184 39.07 2.435 ;
      RECT 39.035 2.188 39.045 2.443 ;
      RECT 39.03 2.189 39.035 2.465 ;
      RECT 39.025 2.19 39.03 2.48 ;
      RECT 39.02 2.191 39.025 2.495 ;
      RECT 39.015 2.192 39.02 2.51 ;
      RECT 39.01 2.193 39.015 2.54 ;
      RECT 39 2.195 39.01 2.573 ;
      RECT 38.985 2.199 39 2.62 ;
      RECT 38.975 2.202 38.985 2.665 ;
      RECT 38.97 2.205 38.975 2.693 ;
      RECT 38.96 2.207 38.97 2.72 ;
      RECT 38.955 2.21 38.96 2.755 ;
      RECT 38.925 2.215 38.955 2.813 ;
      RECT 38.92 2.22 38.925 2.898 ;
      RECT 38.915 2.222 38.92 2.933 ;
      RECT 38.91 2.224 38.915 3.015 ;
      RECT 38.905 2.226 38.91 3.103 ;
      RECT 38.895 2.228 38.905 3.185 ;
      RECT 38.88 2.242 38.895 3.19 ;
      RECT 38.845 2.287 38.88 3.19 ;
      RECT 38.835 2.327 38.845 3.19 ;
      RECT 38.82 2.355 38.835 3.19 ;
      RECT 38.815 2.372 38.82 3.19 ;
      RECT 38.81 2.38 38.815 3.19 ;
      RECT 38.8 2.395 38.805 3.19 ;
      RECT 38.795 2.402 38.8 3.19 ;
      RECT 38.785 2.422 38.795 3.19 ;
      RECT 38.78 2.435 38.785 3.19 ;
      RECT 38.745 2.44 38.75 2.775 ;
      RECT 38.73 2.83 38.75 3.19 ;
      RECT 38.73 2.44 38.74 2.748 ;
      RECT 38.725 2.87 38.73 3.19 ;
      RECT 38.675 2.44 38.725 2.743 ;
      RECT 38.72 2.907 38.725 3.19 ;
      RECT 38.71 2.93 38.72 3.19 ;
      RECT 38.705 2.975 38.71 3.19 ;
      RECT 38.695 2.985 38.705 3.183 ;
      RECT 38.621 2.44 38.675 2.737 ;
      RECT 38.535 2.44 38.621 2.73 ;
      RECT 38.486 2.487 38.535 2.723 ;
      RECT 38.4 2.495 38.486 2.716 ;
      RECT 38.385 2.492 38.4 2.711 ;
      RECT 38.371 2.485 38.385 2.71 ;
      RECT 38.285 2.485 38.371 2.705 ;
      RECT 38.19 2.49 38.2 2.69 ;
      RECT 37.78 1.92 37.795 2.32 ;
      RECT 37.975 1.92 37.98 2.18 ;
      RECT 37.72 1.92 37.765 2.18 ;
      RECT 38.175 3.225 38.18 3.43 ;
      RECT 38.17 3.215 38.175 3.435 ;
      RECT 38.165 3.202 38.17 3.44 ;
      RECT 38.16 3.182 38.165 3.44 ;
      RECT 38.135 3.135 38.16 3.44 ;
      RECT 38.1 3.05 38.135 3.44 ;
      RECT 38.095 2.987 38.1 3.44 ;
      RECT 38.09 2.972 38.095 3.44 ;
      RECT 38.075 2.932 38.09 3.44 ;
      RECT 38.07 2.907 38.075 3.44 ;
      RECT 38.06 2.89 38.07 3.44 ;
      RECT 38.025 2.812 38.06 3.44 ;
      RECT 38.02 2.755 38.025 3.44 ;
      RECT 38.015 2.742 38.02 3.44 ;
      RECT 38.005 2.72 38.015 3.44 ;
      RECT 37.995 2.685 38.005 3.44 ;
      RECT 37.985 2.655 37.995 3.44 ;
      RECT 37.975 2.57 37.985 3.083 ;
      RECT 37.982 3.215 37.985 3.44 ;
      RECT 37.98 3.225 37.982 3.44 ;
      RECT 37.97 3.235 37.98 3.435 ;
      RECT 37.965 1.92 37.975 2.315 ;
      RECT 37.97 2.447 37.975 3.058 ;
      RECT 37.965 2.345 37.97 3.041 ;
      RECT 37.955 1.92 37.965 3.017 ;
      RECT 37.95 1.92 37.955 2.988 ;
      RECT 37.945 1.92 37.95 2.978 ;
      RECT 37.925 1.92 37.945 2.94 ;
      RECT 37.92 1.92 37.925 2.898 ;
      RECT 37.915 1.92 37.92 2.878 ;
      RECT 37.885 1.92 37.915 2.828 ;
      RECT 37.875 1.92 37.885 2.775 ;
      RECT 37.87 1.92 37.875 2.748 ;
      RECT 37.865 1.92 37.87 2.733 ;
      RECT 37.855 1.92 37.865 2.71 ;
      RECT 37.845 1.92 37.855 2.685 ;
      RECT 37.84 1.92 37.845 2.625 ;
      RECT 37.83 1.92 37.84 2.563 ;
      RECT 37.825 1.92 37.83 2.483 ;
      RECT 37.82 1.92 37.825 2.448 ;
      RECT 37.815 1.92 37.82 2.423 ;
      RECT 37.81 1.92 37.815 2.408 ;
      RECT 37.805 1.92 37.81 2.378 ;
      RECT 37.8 1.92 37.805 2.355 ;
      RECT 37.795 1.92 37.8 2.328 ;
      RECT 37.765 1.92 37.78 2.315 ;
      RECT 36.92 3.455 37.105 3.665 ;
      RECT 36.91 3.46 37.12 3.658 ;
      RECT 36.91 3.46 37.14 3.63 ;
      RECT 36.91 3.46 37.155 3.609 ;
      RECT 36.91 3.46 37.17 3.607 ;
      RECT 36.91 3.46 37.18 3.606 ;
      RECT 36.91 3.46 37.21 3.603 ;
      RECT 37.56 3.305 37.82 3.565 ;
      RECT 37.52 3.352 37.82 3.548 ;
      RECT 37.511 3.36 37.52 3.551 ;
      RECT 37.105 3.453 37.82 3.548 ;
      RECT 37.425 3.378 37.511 3.558 ;
      RECT 37.12 3.45 37.82 3.548 ;
      RECT 37.366 3.4 37.425 3.57 ;
      RECT 37.14 3.446 37.82 3.548 ;
      RECT 37.28 3.412 37.366 3.581 ;
      RECT 37.155 3.442 37.82 3.548 ;
      RECT 37.225 3.425 37.28 3.593 ;
      RECT 37.17 3.44 37.82 3.548 ;
      RECT 37.21 3.431 37.225 3.599 ;
      RECT 37.18 3.436 37.82 3.548 ;
      RECT 37.325 2.96 37.585 3.22 ;
      RECT 37.325 2.98 37.695 3.19 ;
      RECT 37.325 2.985 37.705 3.185 ;
      RECT 37.516 2.399 37.595 2.63 ;
      RECT 37.43 2.402 37.645 2.625 ;
      RECT 37.425 2.402 37.645 2.62 ;
      RECT 37.425 2.407 37.655 2.618 ;
      RECT 37.4 2.407 37.655 2.615 ;
      RECT 37.4 2.415 37.665 2.613 ;
      RECT 37.28 2.35 37.54 2.61 ;
      RECT 37.28 2.397 37.59 2.61 ;
      RECT 36.535 2.97 36.54 3.23 ;
      RECT 36.365 2.74 36.37 3.23 ;
      RECT 36.25 2.98 36.255 3.205 ;
      RECT 36.96 2.075 36.965 2.285 ;
      RECT 36.965 2.08 36.98 2.28 ;
      RECT 36.9 2.075 36.96 2.293 ;
      RECT 36.885 2.075 36.9 2.303 ;
      RECT 36.835 2.075 36.885 2.32 ;
      RECT 36.815 2.075 36.835 2.343 ;
      RECT 36.8 2.075 36.815 2.355 ;
      RECT 36.78 2.075 36.8 2.365 ;
      RECT 36.77 2.08 36.78 2.374 ;
      RECT 36.765 2.09 36.77 2.379 ;
      RECT 36.76 2.102 36.765 2.383 ;
      RECT 36.75 2.125 36.76 2.388 ;
      RECT 36.745 2.14 36.75 2.392 ;
      RECT 36.74 2.157 36.745 2.395 ;
      RECT 36.735 2.165 36.74 2.398 ;
      RECT 36.725 2.17 36.735 2.402 ;
      RECT 36.72 2.177 36.725 2.407 ;
      RECT 36.71 2.182 36.72 2.411 ;
      RECT 36.685 2.194 36.71 2.422 ;
      RECT 36.665 2.211 36.685 2.438 ;
      RECT 36.64 2.228 36.665 2.46 ;
      RECT 36.605 2.251 36.64 2.518 ;
      RECT 36.585 2.273 36.605 2.58 ;
      RECT 36.58 2.283 36.585 2.615 ;
      RECT 36.57 2.29 36.58 2.653 ;
      RECT 36.565 2.297 36.57 2.673 ;
      RECT 36.56 2.308 36.565 2.71 ;
      RECT 36.555 2.316 36.56 2.775 ;
      RECT 36.545 2.327 36.555 2.828 ;
      RECT 36.54 2.345 36.545 2.898 ;
      RECT 36.535 2.355 36.54 2.935 ;
      RECT 36.53 2.365 36.535 3.23 ;
      RECT 36.525 2.377 36.53 3.23 ;
      RECT 36.52 2.387 36.525 3.23 ;
      RECT 36.51 2.397 36.52 3.23 ;
      RECT 36.5 2.42 36.51 3.23 ;
      RECT 36.485 2.455 36.5 3.23 ;
      RECT 36.445 2.517 36.485 3.23 ;
      RECT 36.44 2.57 36.445 3.23 ;
      RECT 36.415 2.605 36.44 3.23 ;
      RECT 36.4 2.65 36.415 3.23 ;
      RECT 36.395 2.672 36.4 3.23 ;
      RECT 36.385 2.685 36.395 3.23 ;
      RECT 36.375 2.71 36.385 3.23 ;
      RECT 36.37 2.732 36.375 3.23 ;
      RECT 36.345 2.77 36.365 3.23 ;
      RECT 36.305 2.827 36.345 3.23 ;
      RECT 36.3 2.877 36.305 3.23 ;
      RECT 36.295 2.895 36.3 3.23 ;
      RECT 36.29 2.907 36.295 3.23 ;
      RECT 36.28 2.925 36.29 3.23 ;
      RECT 36.27 2.945 36.28 3.205 ;
      RECT 36.265 2.962 36.27 3.205 ;
      RECT 36.255 2.975 36.265 3.205 ;
      RECT 36.225 2.985 36.25 3.205 ;
      RECT 36.215 2.992 36.225 3.205 ;
      RECT 36.2 3.002 36.215 3.2 ;
      RECT 35.3 7.77 35.59 8 ;
      RECT 35.36 6.29 35.53 8 ;
      RECT 35.35 6.66 35.705 7.015 ;
      RECT 35.3 6.29 35.59 6.52 ;
      RECT 34.895 2.395 35 2.965 ;
      RECT 34.895 2.73 35.22 2.96 ;
      RECT 34.895 2.76 35.39 2.93 ;
      RECT 34.895 2.395 35.085 2.96 ;
      RECT 34.31 2.36 34.6 2.59 ;
      RECT 34.31 2.395 35.085 2.565 ;
      RECT 34.37 0.88 34.54 2.59 ;
      RECT 34.31 0.88 34.6 1.11 ;
      RECT 34.31 7.77 34.6 8 ;
      RECT 34.37 6.29 34.54 8 ;
      RECT 34.31 6.29 34.6 6.52 ;
      RECT 34.31 6.325 35.165 6.485 ;
      RECT 34.995 5.92 35.165 6.485 ;
      RECT 34.31 6.32 34.705 6.485 ;
      RECT 34.93 5.92 35.22 6.15 ;
      RECT 34.93 5.95 35.39 6.12 ;
      RECT 33.94 2.73 34.23 2.96 ;
      RECT 33.94 2.76 34.4 2.93 ;
      RECT 34.005 1.655 34.17 2.96 ;
      RECT 32.52 1.625 32.81 1.855 ;
      RECT 32.52 1.655 34.17 1.825 ;
      RECT 32.58 0.885 32.75 1.855 ;
      RECT 32.52 0.885 32.81 1.115 ;
      RECT 32.52 7.765 32.81 7.995 ;
      RECT 32.58 7.025 32.75 7.995 ;
      RECT 32.58 7.12 34.17 7.29 ;
      RECT 34 5.92 34.17 7.29 ;
      RECT 32.52 7.025 32.81 7.255 ;
      RECT 33.94 5.92 34.23 6.15 ;
      RECT 33.94 5.95 34.4 6.12 ;
      RECT 32.95 1.965 33.3 2.315 ;
      RECT 30.615 2.025 33.3 2.195 ;
      RECT 30.615 1.34 30.785 2.195 ;
      RECT 30.515 1.34 30.865 1.69 ;
      RECT 32.975 6.655 33.3 6.98 ;
      RECT 28.4 6.61 28.75 6.96 ;
      RECT 32.95 6.655 33.3 6.885 ;
      RECT 28.17 6.655 28.75 6.885 ;
      RECT 28 6.685 33.3 6.855 ;
      RECT 32.175 2.365 32.495 2.685 ;
      RECT 32.145 2.365 32.495 2.595 ;
      RECT 31.975 2.395 32.495 2.565 ;
      RECT 32.175 6.255 32.495 6.545 ;
      RECT 32.145 6.285 32.495 6.515 ;
      RECT 31.975 6.315 32.495 6.485 ;
      RECT 28.81 2.465 28.995 2.675 ;
      RECT 28.8 2.47 29.01 2.668 ;
      RECT 28.8 2.47 29.096 2.645 ;
      RECT 28.8 2.47 29.155 2.62 ;
      RECT 28.8 2.47 29.21 2.6 ;
      RECT 28.8 2.47 29.22 2.588 ;
      RECT 28.8 2.47 29.415 2.527 ;
      RECT 28.8 2.47 29.445 2.51 ;
      RECT 28.8 2.47 29.465 2.5 ;
      RECT 29.345 2.235 29.605 2.495 ;
      RECT 29.33 2.325 29.345 2.542 ;
      RECT 28.865 2.457 29.605 2.495 ;
      RECT 29.316 2.336 29.33 2.548 ;
      RECT 28.905 2.45 29.605 2.495 ;
      RECT 29.23 2.376 29.316 2.567 ;
      RECT 29.155 2.437 29.605 2.495 ;
      RECT 29.225 2.412 29.23 2.584 ;
      RECT 29.21 2.422 29.605 2.495 ;
      RECT 29.22 2.417 29.225 2.586 ;
      RECT 29.515 2.922 29.52 3.014 ;
      RECT 29.51 2.9 29.515 3.031 ;
      RECT 29.505 2.89 29.51 3.043 ;
      RECT 29.495 2.881 29.505 3.053 ;
      RECT 29.49 2.876 29.495 3.061 ;
      RECT 29.485 2.735 29.49 3.064 ;
      RECT 29.451 2.735 29.485 3.075 ;
      RECT 29.365 2.735 29.451 3.11 ;
      RECT 29.285 2.735 29.365 3.158 ;
      RECT 29.256 2.735 29.285 3.182 ;
      RECT 29.17 2.735 29.256 3.188 ;
      RECT 29.165 2.919 29.17 3.193 ;
      RECT 29.13 2.93 29.165 3.196 ;
      RECT 29.105 2.945 29.13 3.2 ;
      RECT 29.091 2.954 29.105 3.202 ;
      RECT 29.005 2.981 29.091 3.208 ;
      RECT 28.94 3.022 29.005 3.217 ;
      RECT 28.925 3.042 28.94 3.222 ;
      RECT 28.895 3.052 28.925 3.225 ;
      RECT 28.89 3.062 28.895 3.228 ;
      RECT 28.86 3.067 28.89 3.23 ;
      RECT 28.84 3.072 28.86 3.234 ;
      RECT 28.755 3.075 28.84 3.241 ;
      RECT 28.74 3.072 28.755 3.247 ;
      RECT 28.73 3.069 28.74 3.249 ;
      RECT 28.71 3.066 28.73 3.251 ;
      RECT 28.69 3.062 28.71 3.252 ;
      RECT 28.675 3.058 28.69 3.254 ;
      RECT 28.665 3.055 28.675 3.255 ;
      RECT 28.625 3.049 28.665 3.253 ;
      RECT 28.615 3.044 28.625 3.251 ;
      RECT 28.6 3.041 28.615 3.247 ;
      RECT 28.575 3.036 28.6 3.24 ;
      RECT 28.525 3.027 28.575 3.228 ;
      RECT 28.455 3.013 28.525 3.21 ;
      RECT 28.397 2.998 28.455 3.192 ;
      RECT 28.311 2.981 28.397 3.172 ;
      RECT 28.225 2.96 28.311 3.147 ;
      RECT 28.175 2.945 28.225 3.128 ;
      RECT 28.171 2.939 28.175 3.12 ;
      RECT 28.085 2.929 28.171 3.107 ;
      RECT 28.05 2.914 28.085 3.09 ;
      RECT 28.035 2.907 28.05 3.083 ;
      RECT 27.975 2.895 28.035 3.071 ;
      RECT 27.955 2.882 27.975 3.059 ;
      RECT 27.915 2.873 27.955 3.051 ;
      RECT 27.91 2.865 27.915 3.044 ;
      RECT 27.83 2.855 27.91 3.03 ;
      RECT 27.815 2.842 27.83 3.015 ;
      RECT 27.81 2.84 27.815 3.013 ;
      RECT 27.731 2.828 27.81 3 ;
      RECT 27.645 2.803 27.731 2.975 ;
      RECT 27.63 2.772 27.645 2.96 ;
      RECT 27.615 2.747 27.63 2.956 ;
      RECT 27.6 2.74 27.615 2.952 ;
      RECT 27.425 2.745 27.43 2.948 ;
      RECT 27.42 2.75 27.425 2.943 ;
      RECT 27.43 2.74 27.6 2.95 ;
      RECT 28.145 2.5 28.25 2.76 ;
      RECT 28.96 2.025 28.965 2.25 ;
      RECT 29.09 2.025 29.145 2.235 ;
      RECT 29.145 2.03 29.155 2.228 ;
      RECT 29.051 2.025 29.09 2.238 ;
      RECT 28.965 2.025 29.051 2.245 ;
      RECT 28.945 2.03 28.96 2.251 ;
      RECT 28.935 2.07 28.945 2.253 ;
      RECT 28.905 2.08 28.935 2.255 ;
      RECT 28.9 2.085 28.905 2.257 ;
      RECT 28.875 2.09 28.9 2.259 ;
      RECT 28.86 2.095 28.875 2.261 ;
      RECT 28.845 2.097 28.86 2.263 ;
      RECT 28.84 2.102 28.845 2.265 ;
      RECT 28.79 2.11 28.84 2.268 ;
      RECT 28.765 2.119 28.79 2.273 ;
      RECT 28.755 2.126 28.765 2.278 ;
      RECT 28.75 2.129 28.755 2.282 ;
      RECT 28.73 2.132 28.75 2.291 ;
      RECT 28.7 2.14 28.73 2.311 ;
      RECT 28.671 2.153 28.7 2.333 ;
      RECT 28.585 2.187 28.671 2.377 ;
      RECT 28.58 2.213 28.585 2.415 ;
      RECT 28.575 2.217 28.58 2.424 ;
      RECT 28.54 2.23 28.575 2.457 ;
      RECT 28.53 2.244 28.54 2.495 ;
      RECT 28.525 2.248 28.53 2.508 ;
      RECT 28.52 2.252 28.525 2.513 ;
      RECT 28.51 2.26 28.52 2.525 ;
      RECT 28.505 2.267 28.51 2.54 ;
      RECT 28.48 2.28 28.505 2.565 ;
      RECT 28.44 2.309 28.48 2.62 ;
      RECT 28.425 2.334 28.44 2.675 ;
      RECT 28.415 2.345 28.425 2.698 ;
      RECT 28.41 2.352 28.415 2.71 ;
      RECT 28.405 2.356 28.41 2.718 ;
      RECT 28.35 2.384 28.405 2.76 ;
      RECT 28.33 2.42 28.35 2.76 ;
      RECT 28.315 2.435 28.33 2.76 ;
      RECT 28.26 2.467 28.315 2.76 ;
      RECT 28.25 2.497 28.26 2.76 ;
      RECT 27.86 2.112 28.045 2.35 ;
      RECT 27.845 2.114 28.055 2.345 ;
      RECT 27.73 2.06 27.99 2.32 ;
      RECT 27.725 2.097 27.99 2.274 ;
      RECT 27.72 2.107 27.99 2.271 ;
      RECT 27.715 2.147 28.055 2.265 ;
      RECT 27.71 2.18 28.055 2.255 ;
      RECT 27.72 2.122 28.07 2.193 ;
      RECT 28.017 3.22 28.03 3.75 ;
      RECT 27.931 3.22 28.03 3.749 ;
      RECT 27.931 3.22 28.035 3.748 ;
      RECT 27.845 3.22 28.035 3.746 ;
      RECT 27.84 3.22 28.035 3.743 ;
      RECT 27.84 3.22 28.045 3.741 ;
      RECT 27.835 3.512 28.045 3.738 ;
      RECT 27.835 3.522 28.05 3.735 ;
      RECT 27.835 3.59 28.055 3.731 ;
      RECT 27.825 3.595 28.055 3.73 ;
      RECT 27.825 3.687 28.06 3.727 ;
      RECT 27.81 3.22 28.07 3.48 ;
      RECT 27.74 7.765 28.03 7.995 ;
      RECT 27.8 7.025 27.97 7.995 ;
      RECT 27.715 7.055 28.055 7.4 ;
      RECT 27.74 7.025 28.03 7.4 ;
      RECT 27.04 2.21 27.085 3.745 ;
      RECT 27.24 2.21 27.27 2.425 ;
      RECT 25.615 1.95 25.735 2.16 ;
      RECT 25.275 1.9 25.535 2.16 ;
      RECT 25.275 1.945 25.57 2.15 ;
      RECT 27.28 2.226 27.285 2.28 ;
      RECT 27.275 2.219 27.28 2.413 ;
      RECT 27.27 2.213 27.275 2.42 ;
      RECT 27.225 2.21 27.24 2.433 ;
      RECT 27.22 2.21 27.225 2.455 ;
      RECT 27.215 2.21 27.22 2.503 ;
      RECT 27.21 2.21 27.215 2.523 ;
      RECT 27.2 2.21 27.21 2.63 ;
      RECT 27.195 2.21 27.2 2.693 ;
      RECT 27.19 2.21 27.195 2.75 ;
      RECT 27.185 2.21 27.19 2.758 ;
      RECT 27.17 2.21 27.185 2.865 ;
      RECT 27.16 2.21 27.17 3 ;
      RECT 27.15 2.21 27.16 3.11 ;
      RECT 27.14 2.21 27.15 3.167 ;
      RECT 27.135 2.21 27.14 3.207 ;
      RECT 27.13 2.21 27.135 3.243 ;
      RECT 27.12 2.21 27.13 3.283 ;
      RECT 27.115 2.21 27.12 3.325 ;
      RECT 27.095 2.21 27.115 3.39 ;
      RECT 27.1 3.535 27.105 3.715 ;
      RECT 27.095 3.517 27.1 3.723 ;
      RECT 27.09 2.21 27.095 3.453 ;
      RECT 27.09 3.497 27.095 3.73 ;
      RECT 27.085 2.21 27.09 3.74 ;
      RECT 27.03 2.21 27.04 2.51 ;
      RECT 27.035 2.757 27.04 3.745 ;
      RECT 27.03 2.822 27.035 3.745 ;
      RECT 27.025 2.211 27.03 2.5 ;
      RECT 27.02 2.887 27.03 3.745 ;
      RECT 27.015 2.212 27.025 2.49 ;
      RECT 27.005 3 27.02 3.745 ;
      RECT 27.01 2.213 27.015 2.48 ;
      RECT 26.99 2.214 27.01 2.458 ;
      RECT 26.995 3.097 27.005 3.745 ;
      RECT 26.99 3.172 26.995 3.745 ;
      RECT 26.98 2.213 26.99 2.435 ;
      RECT 26.985 3.215 26.99 3.745 ;
      RECT 26.98 3.242 26.985 3.745 ;
      RECT 26.97 2.211 26.98 2.423 ;
      RECT 26.975 3.285 26.98 3.745 ;
      RECT 26.97 3.312 26.975 3.745 ;
      RECT 26.96 2.21 26.97 2.41 ;
      RECT 26.965 3.327 26.97 3.745 ;
      RECT 26.925 3.385 26.965 3.745 ;
      RECT 26.955 2.209 26.96 2.395 ;
      RECT 26.95 2.207 26.955 2.388 ;
      RECT 26.94 2.204 26.95 2.378 ;
      RECT 26.935 2.201 26.94 2.363 ;
      RECT 26.92 2.197 26.935 2.356 ;
      RECT 26.915 3.44 26.925 3.745 ;
      RECT 26.915 2.194 26.92 2.351 ;
      RECT 26.9 2.19 26.915 2.345 ;
      RECT 26.91 3.457 26.915 3.745 ;
      RECT 26.9 3.52 26.91 3.745 ;
      RECT 26.82 2.175 26.9 2.325 ;
      RECT 26.895 3.527 26.9 3.74 ;
      RECT 26.89 3.535 26.895 3.73 ;
      RECT 26.81 2.161 26.82 2.309 ;
      RECT 26.795 2.157 26.81 2.307 ;
      RECT 26.785 2.152 26.795 2.303 ;
      RECT 26.76 2.145 26.785 2.295 ;
      RECT 26.755 2.14 26.76 2.29 ;
      RECT 26.745 2.14 26.755 2.288 ;
      RECT 26.735 2.138 26.745 2.286 ;
      RECT 26.705 2.13 26.735 2.28 ;
      RECT 26.69 2.122 26.705 2.273 ;
      RECT 26.67 2.117 26.69 2.266 ;
      RECT 26.665 2.113 26.67 2.261 ;
      RECT 26.635 2.106 26.665 2.255 ;
      RECT 26.61 2.097 26.635 2.245 ;
      RECT 26.58 2.09 26.61 2.237 ;
      RECT 26.555 2.08 26.58 2.228 ;
      RECT 26.54 2.072 26.555 2.222 ;
      RECT 26.515 2.067 26.54 2.217 ;
      RECT 26.505 2.063 26.515 2.212 ;
      RECT 26.485 2.058 26.505 2.207 ;
      RECT 26.45 2.053 26.485 2.2 ;
      RECT 26.39 2.048 26.45 2.193 ;
      RECT 26.377 2.044 26.39 2.191 ;
      RECT 26.291 2.039 26.377 2.188 ;
      RECT 26.205 2.029 26.291 2.184 ;
      RECT 26.164 2.022 26.205 2.181 ;
      RECT 26.078 2.015 26.164 2.178 ;
      RECT 25.992 2.005 26.078 2.174 ;
      RECT 25.906 1.995 25.992 2.169 ;
      RECT 25.82 1.985 25.906 2.165 ;
      RECT 25.81 1.97 25.82 2.163 ;
      RECT 25.8 1.955 25.81 2.163 ;
      RECT 25.735 1.95 25.8 2.162 ;
      RECT 25.57 1.947 25.615 2.155 ;
      RECT 26.815 2.852 26.82 3.043 ;
      RECT 26.81 2.847 26.815 3.05 ;
      RECT 26.796 2.845 26.81 3.056 ;
      RECT 26.71 2.845 26.796 3.058 ;
      RECT 26.706 2.845 26.71 3.061 ;
      RECT 26.62 2.845 26.706 3.079 ;
      RECT 26.61 2.85 26.62 3.098 ;
      RECT 26.6 2.905 26.61 3.102 ;
      RECT 26.575 2.92 26.6 3.109 ;
      RECT 26.535 2.94 26.575 3.122 ;
      RECT 26.53 2.952 26.535 3.132 ;
      RECT 26.515 2.958 26.53 3.137 ;
      RECT 26.51 2.963 26.515 3.141 ;
      RECT 26.49 2.97 26.51 3.146 ;
      RECT 26.42 2.995 26.49 3.163 ;
      RECT 26.38 3.023 26.42 3.183 ;
      RECT 26.375 3.033 26.38 3.191 ;
      RECT 26.355 3.04 26.375 3.193 ;
      RECT 26.35 3.047 26.355 3.196 ;
      RECT 26.32 3.055 26.35 3.199 ;
      RECT 26.315 3.06 26.32 3.203 ;
      RECT 26.241 3.064 26.315 3.211 ;
      RECT 26.155 3.073 26.241 3.227 ;
      RECT 26.151 3.078 26.155 3.236 ;
      RECT 26.065 3.083 26.151 3.246 ;
      RECT 26.025 3.091 26.065 3.258 ;
      RECT 25.975 3.097 26.025 3.265 ;
      RECT 25.89 3.106 25.975 3.28 ;
      RECT 25.815 3.117 25.89 3.298 ;
      RECT 25.78 3.124 25.815 3.308 ;
      RECT 25.705 3.132 25.78 3.313 ;
      RECT 25.65 3.141 25.705 3.313 ;
      RECT 25.625 3.146 25.65 3.311 ;
      RECT 25.615 3.149 25.625 3.309 ;
      RECT 25.58 3.151 25.615 3.307 ;
      RECT 25.55 3.153 25.58 3.303 ;
      RECT 25.505 3.152 25.55 3.299 ;
      RECT 25.485 3.147 25.505 3.296 ;
      RECT 25.435 3.132 25.485 3.293 ;
      RECT 25.425 3.117 25.435 3.288 ;
      RECT 25.375 3.102 25.425 3.278 ;
      RECT 25.325 3.077 25.375 3.258 ;
      RECT 25.315 3.062 25.325 3.24 ;
      RECT 25.31 3.06 25.315 3.234 ;
      RECT 25.29 3.055 25.31 3.229 ;
      RECT 25.285 3.047 25.29 3.223 ;
      RECT 25.27 3.041 25.285 3.216 ;
      RECT 25.265 3.036 25.27 3.208 ;
      RECT 25.245 3.031 25.265 3.2 ;
      RECT 25.23 3.024 25.245 3.193 ;
      RECT 25.215 3.018 25.23 3.184 ;
      RECT 25.21 3.012 25.215 3.177 ;
      RECT 25.165 2.987 25.21 3.163 ;
      RECT 25.15 2.957 25.165 3.145 ;
      RECT 25.135 2.94 25.15 3.136 ;
      RECT 25.11 2.92 25.135 3.124 ;
      RECT 25.07 2.89 25.11 3.104 ;
      RECT 25.06 2.86 25.07 3.089 ;
      RECT 25.045 2.85 25.06 3.082 ;
      RECT 24.99 2.815 25.045 3.061 ;
      RECT 24.975 2.778 24.99 3.04 ;
      RECT 24.965 2.765 24.975 3.032 ;
      RECT 24.915 2.735 24.965 3.014 ;
      RECT 24.9 2.665 24.915 2.995 ;
      RECT 24.855 2.665 24.9 2.978 ;
      RECT 24.83 2.665 24.855 2.96 ;
      RECT 24.82 2.665 24.83 2.953 ;
      RECT 24.741 2.665 24.82 2.946 ;
      RECT 24.655 2.665 24.741 2.938 ;
      RECT 24.64 2.697 24.655 2.933 ;
      RECT 24.565 2.707 24.64 2.929 ;
      RECT 24.545 2.717 24.565 2.924 ;
      RECT 24.52 2.717 24.545 2.921 ;
      RECT 24.51 2.707 24.52 2.92 ;
      RECT 24.5 2.68 24.51 2.919 ;
      RECT 24.46 2.675 24.5 2.917 ;
      RECT 24.415 2.675 24.46 2.913 ;
      RECT 24.39 2.675 24.415 2.908 ;
      RECT 24.34 2.675 24.39 2.895 ;
      RECT 24.3 2.68 24.31 2.88 ;
      RECT 24.31 2.675 24.34 2.885 ;
      RECT 26.295 2.455 26.555 2.715 ;
      RECT 26.29 2.477 26.555 2.673 ;
      RECT 25.53 2.305 25.75 2.67 ;
      RECT 25.512 2.392 25.75 2.669 ;
      RECT 25.495 2.397 25.75 2.666 ;
      RECT 25.495 2.397 25.77 2.665 ;
      RECT 25.465 2.407 25.77 2.663 ;
      RECT 25.46 2.422 25.77 2.659 ;
      RECT 25.46 2.422 25.775 2.658 ;
      RECT 25.455 2.48 25.775 2.656 ;
      RECT 25.455 2.48 25.785 2.653 ;
      RECT 25.45 2.545 25.785 2.648 ;
      RECT 25.53 2.305 25.79 2.565 ;
      RECT 24.275 2.135 24.535 2.395 ;
      RECT 24.275 2.178 24.621 2.369 ;
      RECT 24.275 2.178 24.665 2.368 ;
      RECT 24.275 2.178 24.685 2.366 ;
      RECT 24.275 2.178 24.785 2.365 ;
      RECT 24.275 2.178 24.805 2.363 ;
      RECT 24.275 2.178 24.815 2.358 ;
      RECT 24.685 2.145 24.875 2.355 ;
      RECT 24.685 2.147 24.88 2.353 ;
      RECT 24.675 2.152 24.885 2.345 ;
      RECT 24.621 2.176 24.885 2.345 ;
      RECT 24.665 2.17 24.675 2.367 ;
      RECT 24.675 2.15 24.88 2.353 ;
      RECT 23.63 3.21 23.835 3.44 ;
      RECT 23.57 3.16 23.625 3.42 ;
      RECT 23.63 3.16 23.83 3.44 ;
      RECT 24.6 3.475 24.605 3.502 ;
      RECT 24.59 3.385 24.6 3.507 ;
      RECT 24.585 3.307 24.59 3.513 ;
      RECT 24.575 3.297 24.585 3.52 ;
      RECT 24.57 3.287 24.575 3.526 ;
      RECT 24.56 3.282 24.57 3.528 ;
      RECT 24.545 3.274 24.56 3.536 ;
      RECT 24.53 3.265 24.545 3.548 ;
      RECT 24.52 3.257 24.53 3.558 ;
      RECT 24.485 3.175 24.52 3.576 ;
      RECT 24.45 3.175 24.485 3.595 ;
      RECT 24.435 3.175 24.45 3.603 ;
      RECT 24.38 3.175 24.435 3.603 ;
      RECT 24.346 3.175 24.38 3.594 ;
      RECT 24.26 3.175 24.346 3.57 ;
      RECT 24.25 3.235 24.26 3.552 ;
      RECT 24.21 3.237 24.25 3.543 ;
      RECT 24.205 3.239 24.21 3.533 ;
      RECT 24.185 3.241 24.205 3.528 ;
      RECT 24.175 3.244 24.185 3.523 ;
      RECT 24.165 3.245 24.175 3.518 ;
      RECT 24.141 3.246 24.165 3.51 ;
      RECT 24.055 3.251 24.141 3.488 ;
      RECT 24 3.25 24.055 3.461 ;
      RECT 23.985 3.243 24 3.448 ;
      RECT 23.95 3.238 23.985 3.444 ;
      RECT 23.895 3.23 23.95 3.443 ;
      RECT 23.835 3.217 23.895 3.441 ;
      RECT 23.625 3.16 23.63 3.428 ;
      RECT 23.7 2.53 23.885 2.74 ;
      RECT 23.69 2.535 23.9 2.733 ;
      RECT 23.73 2.44 23.99 2.7 ;
      RECT 23.685 2.597 23.99 2.623 ;
      RECT 23.03 2.39 23.035 3.19 ;
      RECT 22.975 2.44 23.005 3.19 ;
      RECT 22.965 2.44 22.97 2.75 ;
      RECT 22.95 2.44 22.955 2.745 ;
      RECT 22.495 2.485 22.51 2.7 ;
      RECT 22.425 2.485 22.51 2.695 ;
      RECT 23.69 2.065 23.76 2.275 ;
      RECT 23.76 2.072 23.77 2.27 ;
      RECT 23.656 2.065 23.69 2.282 ;
      RECT 23.57 2.065 23.656 2.306 ;
      RECT 23.56 2.07 23.57 2.325 ;
      RECT 23.555 2.082 23.56 2.328 ;
      RECT 23.54 2.097 23.555 2.332 ;
      RECT 23.535 2.115 23.54 2.336 ;
      RECT 23.495 2.125 23.535 2.345 ;
      RECT 23.48 2.132 23.495 2.357 ;
      RECT 23.465 2.137 23.48 2.362 ;
      RECT 23.45 2.14 23.465 2.367 ;
      RECT 23.44 2.142 23.45 2.371 ;
      RECT 23.405 2.149 23.44 2.379 ;
      RECT 23.37 2.157 23.405 2.393 ;
      RECT 23.36 2.163 23.37 2.402 ;
      RECT 23.355 2.165 23.36 2.404 ;
      RECT 23.335 2.168 23.355 2.41 ;
      RECT 23.305 2.175 23.335 2.421 ;
      RECT 23.295 2.181 23.305 2.428 ;
      RECT 23.27 2.184 23.295 2.435 ;
      RECT 23.26 2.188 23.27 2.443 ;
      RECT 23.255 2.189 23.26 2.465 ;
      RECT 23.25 2.19 23.255 2.48 ;
      RECT 23.245 2.191 23.25 2.495 ;
      RECT 23.24 2.192 23.245 2.51 ;
      RECT 23.235 2.193 23.24 2.54 ;
      RECT 23.225 2.195 23.235 2.573 ;
      RECT 23.21 2.199 23.225 2.62 ;
      RECT 23.2 2.202 23.21 2.665 ;
      RECT 23.195 2.205 23.2 2.693 ;
      RECT 23.185 2.207 23.195 2.72 ;
      RECT 23.18 2.21 23.185 2.755 ;
      RECT 23.15 2.215 23.18 2.813 ;
      RECT 23.145 2.22 23.15 2.898 ;
      RECT 23.14 2.222 23.145 2.933 ;
      RECT 23.135 2.224 23.14 3.015 ;
      RECT 23.13 2.226 23.135 3.103 ;
      RECT 23.12 2.228 23.13 3.185 ;
      RECT 23.105 2.242 23.12 3.19 ;
      RECT 23.07 2.287 23.105 3.19 ;
      RECT 23.06 2.327 23.07 3.19 ;
      RECT 23.045 2.355 23.06 3.19 ;
      RECT 23.04 2.372 23.045 3.19 ;
      RECT 23.035 2.38 23.04 3.19 ;
      RECT 23.025 2.395 23.03 3.19 ;
      RECT 23.02 2.402 23.025 3.19 ;
      RECT 23.01 2.422 23.02 3.19 ;
      RECT 23.005 2.435 23.01 3.19 ;
      RECT 22.97 2.44 22.975 2.775 ;
      RECT 22.955 2.83 22.975 3.19 ;
      RECT 22.955 2.44 22.965 2.748 ;
      RECT 22.95 2.87 22.955 3.19 ;
      RECT 22.9 2.44 22.95 2.743 ;
      RECT 22.945 2.907 22.95 3.19 ;
      RECT 22.935 2.93 22.945 3.19 ;
      RECT 22.93 2.975 22.935 3.19 ;
      RECT 22.92 2.985 22.93 3.183 ;
      RECT 22.846 2.44 22.9 2.737 ;
      RECT 22.76 2.44 22.846 2.73 ;
      RECT 22.711 2.487 22.76 2.723 ;
      RECT 22.625 2.495 22.711 2.716 ;
      RECT 22.61 2.492 22.625 2.711 ;
      RECT 22.596 2.485 22.61 2.71 ;
      RECT 22.51 2.485 22.596 2.705 ;
      RECT 22.415 2.49 22.425 2.69 ;
      RECT 22.005 1.92 22.02 2.32 ;
      RECT 22.2 1.92 22.205 2.18 ;
      RECT 21.945 1.92 21.99 2.18 ;
      RECT 22.4 3.225 22.405 3.43 ;
      RECT 22.395 3.215 22.4 3.435 ;
      RECT 22.39 3.202 22.395 3.44 ;
      RECT 22.385 3.182 22.39 3.44 ;
      RECT 22.36 3.135 22.385 3.44 ;
      RECT 22.325 3.05 22.36 3.44 ;
      RECT 22.32 2.987 22.325 3.44 ;
      RECT 22.315 2.972 22.32 3.44 ;
      RECT 22.3 2.932 22.315 3.44 ;
      RECT 22.295 2.907 22.3 3.44 ;
      RECT 22.285 2.89 22.295 3.44 ;
      RECT 22.25 2.812 22.285 3.44 ;
      RECT 22.245 2.755 22.25 3.44 ;
      RECT 22.24 2.742 22.245 3.44 ;
      RECT 22.23 2.72 22.24 3.44 ;
      RECT 22.22 2.685 22.23 3.44 ;
      RECT 22.21 2.655 22.22 3.44 ;
      RECT 22.2 2.57 22.21 3.083 ;
      RECT 22.207 3.215 22.21 3.44 ;
      RECT 22.205 3.225 22.207 3.44 ;
      RECT 22.195 3.235 22.205 3.435 ;
      RECT 22.19 1.92 22.2 2.315 ;
      RECT 22.195 2.447 22.2 3.058 ;
      RECT 22.19 2.345 22.195 3.041 ;
      RECT 22.18 1.92 22.19 3.017 ;
      RECT 22.175 1.92 22.18 2.988 ;
      RECT 22.17 1.92 22.175 2.978 ;
      RECT 22.15 1.92 22.17 2.94 ;
      RECT 22.145 1.92 22.15 2.898 ;
      RECT 22.14 1.92 22.145 2.878 ;
      RECT 22.11 1.92 22.14 2.828 ;
      RECT 22.1 1.92 22.11 2.775 ;
      RECT 22.095 1.92 22.1 2.748 ;
      RECT 22.09 1.92 22.095 2.733 ;
      RECT 22.08 1.92 22.09 2.71 ;
      RECT 22.07 1.92 22.08 2.685 ;
      RECT 22.065 1.92 22.07 2.625 ;
      RECT 22.055 1.92 22.065 2.563 ;
      RECT 22.05 1.92 22.055 2.483 ;
      RECT 22.045 1.92 22.05 2.448 ;
      RECT 22.04 1.92 22.045 2.423 ;
      RECT 22.035 1.92 22.04 2.408 ;
      RECT 22.03 1.92 22.035 2.378 ;
      RECT 22.025 1.92 22.03 2.355 ;
      RECT 22.02 1.92 22.025 2.328 ;
      RECT 21.99 1.92 22.005 2.315 ;
      RECT 21.145 3.455 21.33 3.665 ;
      RECT 21.135 3.46 21.345 3.658 ;
      RECT 21.135 3.46 21.365 3.63 ;
      RECT 21.135 3.46 21.38 3.609 ;
      RECT 21.135 3.46 21.395 3.607 ;
      RECT 21.135 3.46 21.405 3.606 ;
      RECT 21.135 3.46 21.435 3.603 ;
      RECT 21.785 3.305 22.045 3.565 ;
      RECT 21.745 3.352 22.045 3.548 ;
      RECT 21.736 3.36 21.745 3.551 ;
      RECT 21.33 3.453 22.045 3.548 ;
      RECT 21.65 3.378 21.736 3.558 ;
      RECT 21.345 3.45 22.045 3.548 ;
      RECT 21.591 3.4 21.65 3.57 ;
      RECT 21.365 3.446 22.045 3.548 ;
      RECT 21.505 3.412 21.591 3.581 ;
      RECT 21.38 3.442 22.045 3.548 ;
      RECT 21.45 3.425 21.505 3.593 ;
      RECT 21.395 3.44 22.045 3.548 ;
      RECT 21.435 3.431 21.45 3.599 ;
      RECT 21.405 3.436 22.045 3.548 ;
      RECT 21.55 2.96 21.81 3.22 ;
      RECT 21.55 2.98 21.92 3.19 ;
      RECT 21.55 2.985 21.93 3.185 ;
      RECT 21.741 2.399 21.82 2.63 ;
      RECT 21.655 2.402 21.87 2.625 ;
      RECT 21.65 2.402 21.87 2.62 ;
      RECT 21.65 2.407 21.88 2.618 ;
      RECT 21.625 2.407 21.88 2.615 ;
      RECT 21.625 2.415 21.89 2.613 ;
      RECT 21.505 2.35 21.765 2.61 ;
      RECT 21.505 2.397 21.815 2.61 ;
      RECT 20.76 2.97 20.765 3.23 ;
      RECT 20.59 2.74 20.595 3.23 ;
      RECT 20.475 2.98 20.48 3.205 ;
      RECT 21.185 2.075 21.19 2.285 ;
      RECT 21.19 2.08 21.205 2.28 ;
      RECT 21.125 2.075 21.185 2.293 ;
      RECT 21.11 2.075 21.125 2.303 ;
      RECT 21.06 2.075 21.11 2.32 ;
      RECT 21.04 2.075 21.06 2.343 ;
      RECT 21.025 2.075 21.04 2.355 ;
      RECT 21.005 2.075 21.025 2.365 ;
      RECT 20.995 2.08 21.005 2.374 ;
      RECT 20.99 2.09 20.995 2.379 ;
      RECT 20.985 2.102 20.99 2.383 ;
      RECT 20.975 2.125 20.985 2.388 ;
      RECT 20.97 2.14 20.975 2.392 ;
      RECT 20.965 2.157 20.97 2.395 ;
      RECT 20.96 2.165 20.965 2.398 ;
      RECT 20.95 2.17 20.96 2.402 ;
      RECT 20.945 2.177 20.95 2.407 ;
      RECT 20.935 2.182 20.945 2.411 ;
      RECT 20.91 2.194 20.935 2.422 ;
      RECT 20.89 2.211 20.91 2.438 ;
      RECT 20.865 2.228 20.89 2.46 ;
      RECT 20.83 2.251 20.865 2.518 ;
      RECT 20.81 2.273 20.83 2.58 ;
      RECT 20.805 2.283 20.81 2.615 ;
      RECT 20.795 2.29 20.805 2.653 ;
      RECT 20.79 2.297 20.795 2.673 ;
      RECT 20.785 2.308 20.79 2.71 ;
      RECT 20.78 2.316 20.785 2.775 ;
      RECT 20.77 2.327 20.78 2.828 ;
      RECT 20.765 2.345 20.77 2.898 ;
      RECT 20.76 2.355 20.765 2.935 ;
      RECT 20.755 2.365 20.76 3.23 ;
      RECT 20.75 2.377 20.755 3.23 ;
      RECT 20.745 2.387 20.75 3.23 ;
      RECT 20.735 2.397 20.745 3.23 ;
      RECT 20.725 2.42 20.735 3.23 ;
      RECT 20.71 2.455 20.725 3.23 ;
      RECT 20.67 2.517 20.71 3.23 ;
      RECT 20.665 2.57 20.67 3.23 ;
      RECT 20.64 2.605 20.665 3.23 ;
      RECT 20.625 2.65 20.64 3.23 ;
      RECT 20.62 2.672 20.625 3.23 ;
      RECT 20.61 2.685 20.62 3.23 ;
      RECT 20.6 2.71 20.61 3.23 ;
      RECT 20.595 2.732 20.6 3.23 ;
      RECT 20.57 2.77 20.59 3.23 ;
      RECT 20.53 2.827 20.57 3.23 ;
      RECT 20.525 2.877 20.53 3.23 ;
      RECT 20.52 2.895 20.525 3.23 ;
      RECT 20.515 2.907 20.52 3.23 ;
      RECT 20.505 2.925 20.515 3.23 ;
      RECT 20.495 2.945 20.505 3.205 ;
      RECT 20.49 2.962 20.495 3.205 ;
      RECT 20.48 2.975 20.49 3.205 ;
      RECT 20.45 2.985 20.475 3.205 ;
      RECT 20.44 2.992 20.45 3.205 ;
      RECT 20.425 3.002 20.44 3.2 ;
      RECT 19.52 7.77 19.81 8 ;
      RECT 19.58 6.29 19.75 8 ;
      RECT 19.575 6.655 19.925 7.005 ;
      RECT 19.52 6.29 19.81 6.52 ;
      RECT 19.115 2.395 19.22 2.965 ;
      RECT 19.115 2.73 19.44 2.96 ;
      RECT 19.115 2.76 19.61 2.93 ;
      RECT 19.115 2.395 19.305 2.96 ;
      RECT 18.53 2.36 18.82 2.59 ;
      RECT 18.53 2.395 19.305 2.565 ;
      RECT 18.59 0.88 18.76 2.59 ;
      RECT 18.53 0.88 18.82 1.11 ;
      RECT 18.53 7.77 18.82 8 ;
      RECT 18.59 6.29 18.76 8 ;
      RECT 18.53 6.29 18.82 6.52 ;
      RECT 18.53 6.325 19.385 6.485 ;
      RECT 19.215 5.92 19.385 6.485 ;
      RECT 18.53 6.32 18.925 6.485 ;
      RECT 19.15 5.92 19.44 6.15 ;
      RECT 19.15 5.95 19.61 6.12 ;
      RECT 18.16 2.73 18.45 2.96 ;
      RECT 18.16 2.76 18.62 2.93 ;
      RECT 18.225 1.655 18.39 2.96 ;
      RECT 16.74 1.625 17.03 1.855 ;
      RECT 16.74 1.655 18.39 1.825 ;
      RECT 16.8 0.885 16.97 1.855 ;
      RECT 16.74 0.885 17.03 1.115 ;
      RECT 16.74 7.765 17.03 7.995 ;
      RECT 16.8 7.025 16.97 7.995 ;
      RECT 16.8 7.12 18.39 7.29 ;
      RECT 18.22 5.92 18.39 7.29 ;
      RECT 16.74 7.025 17.03 7.255 ;
      RECT 18.16 5.92 18.45 6.15 ;
      RECT 18.16 5.95 18.62 6.12 ;
      RECT 17.17 1.965 17.52 2.315 ;
      RECT 14.835 2.025 17.52 2.195 ;
      RECT 14.835 1.34 15.005 2.195 ;
      RECT 14.735 1.34 15.085 1.69 ;
      RECT 17.195 6.655 17.52 6.98 ;
      RECT 12.59 6.605 12.94 6.955 ;
      RECT 17.17 6.655 17.52 6.885 ;
      RECT 12.39 6.655 12.94 6.885 ;
      RECT 12.22 6.685 17.52 6.855 ;
      RECT 16.395 2.365 16.715 2.685 ;
      RECT 16.365 2.365 16.715 2.595 ;
      RECT 16.195 2.395 16.715 2.565 ;
      RECT 16.395 6.255 16.715 6.545 ;
      RECT 16.365 6.285 16.715 6.515 ;
      RECT 16.195 6.315 16.715 6.485 ;
      RECT 13.03 2.465 13.215 2.675 ;
      RECT 13.02 2.47 13.23 2.668 ;
      RECT 13.02 2.47 13.316 2.645 ;
      RECT 13.02 2.47 13.375 2.62 ;
      RECT 13.02 2.47 13.43 2.6 ;
      RECT 13.02 2.47 13.44 2.588 ;
      RECT 13.02 2.47 13.635 2.527 ;
      RECT 13.02 2.47 13.665 2.51 ;
      RECT 13.02 2.47 13.685 2.5 ;
      RECT 13.565 2.235 13.825 2.495 ;
      RECT 13.55 2.325 13.565 2.542 ;
      RECT 13.085 2.457 13.825 2.495 ;
      RECT 13.536 2.336 13.55 2.548 ;
      RECT 13.125 2.45 13.825 2.495 ;
      RECT 13.45 2.376 13.536 2.567 ;
      RECT 13.375 2.437 13.825 2.495 ;
      RECT 13.445 2.412 13.45 2.584 ;
      RECT 13.43 2.422 13.825 2.495 ;
      RECT 13.44 2.417 13.445 2.586 ;
      RECT 13.735 2.922 13.74 3.014 ;
      RECT 13.73 2.9 13.735 3.031 ;
      RECT 13.725 2.89 13.73 3.043 ;
      RECT 13.715 2.881 13.725 3.053 ;
      RECT 13.71 2.876 13.715 3.061 ;
      RECT 13.705 2.735 13.71 3.064 ;
      RECT 13.671 2.735 13.705 3.075 ;
      RECT 13.585 2.735 13.671 3.11 ;
      RECT 13.505 2.735 13.585 3.158 ;
      RECT 13.476 2.735 13.505 3.182 ;
      RECT 13.39 2.735 13.476 3.188 ;
      RECT 13.385 2.919 13.39 3.193 ;
      RECT 13.35 2.93 13.385 3.196 ;
      RECT 13.325 2.945 13.35 3.2 ;
      RECT 13.311 2.954 13.325 3.202 ;
      RECT 13.225 2.981 13.311 3.208 ;
      RECT 13.16 3.022 13.225 3.217 ;
      RECT 13.145 3.042 13.16 3.222 ;
      RECT 13.115 3.052 13.145 3.225 ;
      RECT 13.11 3.062 13.115 3.228 ;
      RECT 13.08 3.067 13.11 3.23 ;
      RECT 13.06 3.072 13.08 3.234 ;
      RECT 12.975 3.075 13.06 3.241 ;
      RECT 12.96 3.072 12.975 3.247 ;
      RECT 12.95 3.069 12.96 3.249 ;
      RECT 12.93 3.066 12.95 3.251 ;
      RECT 12.91 3.062 12.93 3.252 ;
      RECT 12.895 3.058 12.91 3.254 ;
      RECT 12.885 3.055 12.895 3.255 ;
      RECT 12.845 3.049 12.885 3.253 ;
      RECT 12.835 3.044 12.845 3.251 ;
      RECT 12.82 3.041 12.835 3.247 ;
      RECT 12.795 3.036 12.82 3.24 ;
      RECT 12.745 3.027 12.795 3.228 ;
      RECT 12.675 3.013 12.745 3.21 ;
      RECT 12.617 2.998 12.675 3.192 ;
      RECT 12.531 2.981 12.617 3.172 ;
      RECT 12.445 2.96 12.531 3.147 ;
      RECT 12.395 2.945 12.445 3.128 ;
      RECT 12.391 2.939 12.395 3.12 ;
      RECT 12.305 2.929 12.391 3.107 ;
      RECT 12.27 2.914 12.305 3.09 ;
      RECT 12.255 2.907 12.27 3.083 ;
      RECT 12.195 2.895 12.255 3.071 ;
      RECT 12.175 2.882 12.195 3.059 ;
      RECT 12.135 2.873 12.175 3.051 ;
      RECT 12.13 2.865 12.135 3.044 ;
      RECT 12.05 2.855 12.13 3.03 ;
      RECT 12.035 2.842 12.05 3.015 ;
      RECT 12.03 2.84 12.035 3.013 ;
      RECT 11.951 2.828 12.03 3 ;
      RECT 11.865 2.803 11.951 2.975 ;
      RECT 11.85 2.772 11.865 2.96 ;
      RECT 11.835 2.747 11.85 2.956 ;
      RECT 11.82 2.74 11.835 2.952 ;
      RECT 11.645 2.745 11.65 2.948 ;
      RECT 11.64 2.75 11.645 2.943 ;
      RECT 11.65 2.74 11.82 2.95 ;
      RECT 12.365 2.5 12.47 2.76 ;
      RECT 13.18 2.025 13.185 2.25 ;
      RECT 13.31 2.025 13.365 2.235 ;
      RECT 13.365 2.03 13.375 2.228 ;
      RECT 13.271 2.025 13.31 2.238 ;
      RECT 13.185 2.025 13.271 2.245 ;
      RECT 13.165 2.03 13.18 2.251 ;
      RECT 13.155 2.07 13.165 2.253 ;
      RECT 13.125 2.08 13.155 2.255 ;
      RECT 13.12 2.085 13.125 2.257 ;
      RECT 13.095 2.09 13.12 2.259 ;
      RECT 13.08 2.095 13.095 2.261 ;
      RECT 13.065 2.097 13.08 2.263 ;
      RECT 13.06 2.102 13.065 2.265 ;
      RECT 13.01 2.11 13.06 2.268 ;
      RECT 12.985 2.119 13.01 2.273 ;
      RECT 12.975 2.126 12.985 2.278 ;
      RECT 12.97 2.129 12.975 2.282 ;
      RECT 12.95 2.132 12.97 2.291 ;
      RECT 12.92 2.14 12.95 2.311 ;
      RECT 12.891 2.153 12.92 2.333 ;
      RECT 12.805 2.187 12.891 2.377 ;
      RECT 12.8 2.213 12.805 2.415 ;
      RECT 12.795 2.217 12.8 2.424 ;
      RECT 12.76 2.23 12.795 2.457 ;
      RECT 12.75 2.244 12.76 2.495 ;
      RECT 12.745 2.248 12.75 2.508 ;
      RECT 12.74 2.252 12.745 2.513 ;
      RECT 12.73 2.26 12.74 2.525 ;
      RECT 12.725 2.267 12.73 2.54 ;
      RECT 12.7 2.28 12.725 2.565 ;
      RECT 12.66 2.309 12.7 2.62 ;
      RECT 12.645 2.334 12.66 2.675 ;
      RECT 12.635 2.345 12.645 2.698 ;
      RECT 12.63 2.352 12.635 2.71 ;
      RECT 12.625 2.356 12.63 2.718 ;
      RECT 12.57 2.384 12.625 2.76 ;
      RECT 12.55 2.42 12.57 2.76 ;
      RECT 12.535 2.435 12.55 2.76 ;
      RECT 12.48 2.467 12.535 2.76 ;
      RECT 12.47 2.497 12.48 2.76 ;
      RECT 12.08 2.112 12.265 2.35 ;
      RECT 12.065 2.114 12.275 2.345 ;
      RECT 11.95 2.06 12.21 2.32 ;
      RECT 11.945 2.097 12.21 2.274 ;
      RECT 11.94 2.107 12.21 2.271 ;
      RECT 11.935 2.147 12.275 2.265 ;
      RECT 11.93 2.18 12.275 2.255 ;
      RECT 11.94 2.122 12.29 2.193 ;
      RECT 12.237 3.22 12.25 3.75 ;
      RECT 12.151 3.22 12.25 3.749 ;
      RECT 12.151 3.22 12.255 3.748 ;
      RECT 12.065 3.22 12.255 3.746 ;
      RECT 12.06 3.22 12.255 3.743 ;
      RECT 12.06 3.22 12.265 3.741 ;
      RECT 12.055 3.512 12.265 3.738 ;
      RECT 12.055 3.522 12.27 3.735 ;
      RECT 12.055 3.59 12.275 3.731 ;
      RECT 12.045 3.595 12.275 3.73 ;
      RECT 12.045 3.687 12.28 3.727 ;
      RECT 12.03 3.22 12.29 3.48 ;
      RECT 11.96 7.765 12.25 7.995 ;
      RECT 12.02 7.025 12.19 7.995 ;
      RECT 11.935 7.055 12.275 7.4 ;
      RECT 11.96 7.025 12.25 7.4 ;
      RECT 11.26 2.21 11.305 3.745 ;
      RECT 11.46 2.21 11.49 2.425 ;
      RECT 9.835 1.95 9.955 2.16 ;
      RECT 9.495 1.9 9.755 2.16 ;
      RECT 9.495 1.945 9.79 2.15 ;
      RECT 11.5 2.226 11.505 2.28 ;
      RECT 11.495 2.219 11.5 2.413 ;
      RECT 11.49 2.213 11.495 2.42 ;
      RECT 11.445 2.21 11.46 2.433 ;
      RECT 11.44 2.21 11.445 2.455 ;
      RECT 11.435 2.21 11.44 2.503 ;
      RECT 11.43 2.21 11.435 2.523 ;
      RECT 11.42 2.21 11.43 2.63 ;
      RECT 11.415 2.21 11.42 2.693 ;
      RECT 11.41 2.21 11.415 2.75 ;
      RECT 11.405 2.21 11.41 2.758 ;
      RECT 11.39 2.21 11.405 2.865 ;
      RECT 11.38 2.21 11.39 3 ;
      RECT 11.37 2.21 11.38 3.11 ;
      RECT 11.36 2.21 11.37 3.167 ;
      RECT 11.355 2.21 11.36 3.207 ;
      RECT 11.35 2.21 11.355 3.243 ;
      RECT 11.34 2.21 11.35 3.283 ;
      RECT 11.335 2.21 11.34 3.325 ;
      RECT 11.315 2.21 11.335 3.39 ;
      RECT 11.32 3.535 11.325 3.715 ;
      RECT 11.315 3.517 11.32 3.723 ;
      RECT 11.31 2.21 11.315 3.453 ;
      RECT 11.31 3.497 11.315 3.73 ;
      RECT 11.305 2.21 11.31 3.74 ;
      RECT 11.25 2.21 11.26 2.51 ;
      RECT 11.255 2.757 11.26 3.745 ;
      RECT 11.25 2.822 11.255 3.745 ;
      RECT 11.245 2.211 11.25 2.5 ;
      RECT 11.24 2.887 11.25 3.745 ;
      RECT 11.235 2.212 11.245 2.49 ;
      RECT 11.225 3 11.24 3.745 ;
      RECT 11.23 2.213 11.235 2.48 ;
      RECT 11.21 2.214 11.23 2.458 ;
      RECT 11.215 3.097 11.225 3.745 ;
      RECT 11.21 3.172 11.215 3.745 ;
      RECT 11.2 2.213 11.21 2.435 ;
      RECT 11.205 3.215 11.21 3.745 ;
      RECT 11.2 3.242 11.205 3.745 ;
      RECT 11.19 2.211 11.2 2.423 ;
      RECT 11.195 3.285 11.2 3.745 ;
      RECT 11.19 3.312 11.195 3.745 ;
      RECT 11.18 2.21 11.19 2.41 ;
      RECT 11.185 3.327 11.19 3.745 ;
      RECT 11.145 3.385 11.185 3.745 ;
      RECT 11.175 2.209 11.18 2.395 ;
      RECT 11.17 2.207 11.175 2.388 ;
      RECT 11.16 2.204 11.17 2.378 ;
      RECT 11.155 2.201 11.16 2.363 ;
      RECT 11.14 2.197 11.155 2.356 ;
      RECT 11.135 3.44 11.145 3.745 ;
      RECT 11.135 2.194 11.14 2.351 ;
      RECT 11.12 2.19 11.135 2.345 ;
      RECT 11.13 3.457 11.135 3.745 ;
      RECT 11.12 3.52 11.13 3.745 ;
      RECT 11.04 2.175 11.12 2.325 ;
      RECT 11.115 3.527 11.12 3.74 ;
      RECT 11.11 3.535 11.115 3.73 ;
      RECT 11.03 2.161 11.04 2.309 ;
      RECT 11.015 2.157 11.03 2.307 ;
      RECT 11.005 2.152 11.015 2.303 ;
      RECT 10.98 2.145 11.005 2.295 ;
      RECT 10.975 2.14 10.98 2.29 ;
      RECT 10.965 2.14 10.975 2.288 ;
      RECT 10.955 2.138 10.965 2.286 ;
      RECT 10.925 2.13 10.955 2.28 ;
      RECT 10.91 2.122 10.925 2.273 ;
      RECT 10.89 2.117 10.91 2.266 ;
      RECT 10.885 2.113 10.89 2.261 ;
      RECT 10.855 2.106 10.885 2.255 ;
      RECT 10.83 2.097 10.855 2.245 ;
      RECT 10.8 2.09 10.83 2.237 ;
      RECT 10.775 2.08 10.8 2.228 ;
      RECT 10.76 2.072 10.775 2.222 ;
      RECT 10.735 2.067 10.76 2.217 ;
      RECT 10.725 2.063 10.735 2.212 ;
      RECT 10.705 2.058 10.725 2.207 ;
      RECT 10.67 2.053 10.705 2.2 ;
      RECT 10.61 2.048 10.67 2.193 ;
      RECT 10.597 2.044 10.61 2.191 ;
      RECT 10.511 2.039 10.597 2.188 ;
      RECT 10.425 2.029 10.511 2.184 ;
      RECT 10.384 2.022 10.425 2.181 ;
      RECT 10.298 2.015 10.384 2.178 ;
      RECT 10.212 2.005 10.298 2.174 ;
      RECT 10.126 1.995 10.212 2.169 ;
      RECT 10.04 1.985 10.126 2.165 ;
      RECT 10.03 1.97 10.04 2.163 ;
      RECT 10.02 1.955 10.03 2.163 ;
      RECT 9.955 1.95 10.02 2.162 ;
      RECT 9.79 1.947 9.835 2.155 ;
      RECT 11.035 2.852 11.04 3.043 ;
      RECT 11.03 2.847 11.035 3.05 ;
      RECT 11.016 2.845 11.03 3.056 ;
      RECT 10.93 2.845 11.016 3.058 ;
      RECT 10.926 2.845 10.93 3.061 ;
      RECT 10.84 2.845 10.926 3.079 ;
      RECT 10.83 2.85 10.84 3.098 ;
      RECT 10.82 2.905 10.83 3.102 ;
      RECT 10.795 2.92 10.82 3.109 ;
      RECT 10.755 2.94 10.795 3.122 ;
      RECT 10.75 2.952 10.755 3.132 ;
      RECT 10.735 2.958 10.75 3.137 ;
      RECT 10.73 2.963 10.735 3.141 ;
      RECT 10.71 2.97 10.73 3.146 ;
      RECT 10.64 2.995 10.71 3.163 ;
      RECT 10.6 3.023 10.64 3.183 ;
      RECT 10.595 3.033 10.6 3.191 ;
      RECT 10.575 3.04 10.595 3.193 ;
      RECT 10.57 3.047 10.575 3.196 ;
      RECT 10.54 3.055 10.57 3.199 ;
      RECT 10.535 3.06 10.54 3.203 ;
      RECT 10.461 3.064 10.535 3.211 ;
      RECT 10.375 3.073 10.461 3.227 ;
      RECT 10.371 3.078 10.375 3.236 ;
      RECT 10.285 3.083 10.371 3.246 ;
      RECT 10.245 3.091 10.285 3.258 ;
      RECT 10.195 3.097 10.245 3.265 ;
      RECT 10.11 3.106 10.195 3.28 ;
      RECT 10.035 3.117 10.11 3.298 ;
      RECT 10 3.124 10.035 3.308 ;
      RECT 9.925 3.132 10 3.313 ;
      RECT 9.87 3.141 9.925 3.313 ;
      RECT 9.845 3.146 9.87 3.311 ;
      RECT 9.835 3.149 9.845 3.309 ;
      RECT 9.8 3.151 9.835 3.307 ;
      RECT 9.77 3.153 9.8 3.303 ;
      RECT 9.725 3.152 9.77 3.299 ;
      RECT 9.705 3.147 9.725 3.296 ;
      RECT 9.655 3.132 9.705 3.293 ;
      RECT 9.645 3.117 9.655 3.288 ;
      RECT 9.595 3.102 9.645 3.278 ;
      RECT 9.545 3.077 9.595 3.258 ;
      RECT 9.535 3.062 9.545 3.24 ;
      RECT 9.53 3.06 9.535 3.234 ;
      RECT 9.51 3.055 9.53 3.229 ;
      RECT 9.505 3.047 9.51 3.223 ;
      RECT 9.49 3.041 9.505 3.216 ;
      RECT 9.485 3.036 9.49 3.208 ;
      RECT 9.465 3.031 9.485 3.2 ;
      RECT 9.45 3.024 9.465 3.193 ;
      RECT 9.435 3.018 9.45 3.184 ;
      RECT 9.43 3.012 9.435 3.177 ;
      RECT 9.385 2.987 9.43 3.163 ;
      RECT 9.37 2.957 9.385 3.145 ;
      RECT 9.355 2.94 9.37 3.136 ;
      RECT 9.33 2.92 9.355 3.124 ;
      RECT 9.29 2.89 9.33 3.104 ;
      RECT 9.28 2.86 9.29 3.089 ;
      RECT 9.265 2.85 9.28 3.082 ;
      RECT 9.21 2.815 9.265 3.061 ;
      RECT 9.195 2.778 9.21 3.04 ;
      RECT 9.185 2.765 9.195 3.032 ;
      RECT 9.135 2.735 9.185 3.014 ;
      RECT 9.12 2.665 9.135 2.995 ;
      RECT 9.075 2.665 9.12 2.978 ;
      RECT 9.05 2.665 9.075 2.96 ;
      RECT 9.04 2.665 9.05 2.953 ;
      RECT 8.961 2.665 9.04 2.946 ;
      RECT 8.875 2.665 8.961 2.938 ;
      RECT 8.86 2.697 8.875 2.933 ;
      RECT 8.785 2.707 8.86 2.929 ;
      RECT 8.765 2.717 8.785 2.924 ;
      RECT 8.74 2.717 8.765 2.921 ;
      RECT 8.73 2.707 8.74 2.92 ;
      RECT 8.72 2.68 8.73 2.919 ;
      RECT 8.68 2.675 8.72 2.917 ;
      RECT 8.635 2.675 8.68 2.913 ;
      RECT 8.61 2.675 8.635 2.908 ;
      RECT 8.56 2.675 8.61 2.895 ;
      RECT 8.52 2.68 8.53 2.88 ;
      RECT 8.53 2.675 8.56 2.885 ;
      RECT 10.515 2.455 10.775 2.715 ;
      RECT 10.51 2.477 10.775 2.673 ;
      RECT 9.75 2.305 9.97 2.67 ;
      RECT 9.732 2.392 9.97 2.669 ;
      RECT 9.715 2.397 9.97 2.666 ;
      RECT 9.715 2.397 9.99 2.665 ;
      RECT 9.685 2.407 9.99 2.663 ;
      RECT 9.68 2.422 9.99 2.659 ;
      RECT 9.68 2.422 9.995 2.658 ;
      RECT 9.675 2.48 9.995 2.656 ;
      RECT 9.675 2.48 10.005 2.653 ;
      RECT 9.67 2.545 10.005 2.648 ;
      RECT 9.75 2.305 10.01 2.565 ;
      RECT 8.495 2.135 8.755 2.395 ;
      RECT 8.495 2.178 8.841 2.369 ;
      RECT 8.495 2.178 8.885 2.368 ;
      RECT 8.495 2.178 8.905 2.366 ;
      RECT 8.495 2.178 9.005 2.365 ;
      RECT 8.495 2.178 9.025 2.363 ;
      RECT 8.495 2.178 9.035 2.358 ;
      RECT 8.905 2.145 9.095 2.355 ;
      RECT 8.905 2.147 9.1 2.353 ;
      RECT 8.895 2.152 9.105 2.345 ;
      RECT 8.841 2.176 9.105 2.345 ;
      RECT 8.885 2.17 8.895 2.367 ;
      RECT 8.895 2.15 9.1 2.353 ;
      RECT 7.85 3.21 8.055 3.44 ;
      RECT 7.79 3.16 7.845 3.42 ;
      RECT 7.85 3.16 8.05 3.44 ;
      RECT 8.82 3.475 8.825 3.502 ;
      RECT 8.81 3.385 8.82 3.507 ;
      RECT 8.805 3.307 8.81 3.513 ;
      RECT 8.795 3.297 8.805 3.52 ;
      RECT 8.79 3.287 8.795 3.526 ;
      RECT 8.78 3.282 8.79 3.528 ;
      RECT 8.765 3.274 8.78 3.536 ;
      RECT 8.75 3.265 8.765 3.548 ;
      RECT 8.74 3.257 8.75 3.558 ;
      RECT 8.705 3.175 8.74 3.576 ;
      RECT 8.67 3.175 8.705 3.595 ;
      RECT 8.655 3.175 8.67 3.603 ;
      RECT 8.6 3.175 8.655 3.603 ;
      RECT 8.566 3.175 8.6 3.594 ;
      RECT 8.48 3.175 8.566 3.57 ;
      RECT 8.47 3.235 8.48 3.552 ;
      RECT 8.43 3.237 8.47 3.543 ;
      RECT 8.425 3.239 8.43 3.533 ;
      RECT 8.405 3.241 8.425 3.528 ;
      RECT 8.395 3.244 8.405 3.523 ;
      RECT 8.385 3.245 8.395 3.518 ;
      RECT 8.361 3.246 8.385 3.51 ;
      RECT 8.275 3.251 8.361 3.488 ;
      RECT 8.22 3.25 8.275 3.461 ;
      RECT 8.205 3.243 8.22 3.448 ;
      RECT 8.17 3.238 8.205 3.444 ;
      RECT 8.115 3.23 8.17 3.443 ;
      RECT 8.055 3.217 8.115 3.441 ;
      RECT 7.845 3.16 7.85 3.428 ;
      RECT 7.92 2.53 8.105 2.74 ;
      RECT 7.91 2.535 8.12 2.733 ;
      RECT 7.95 2.44 8.21 2.7 ;
      RECT 7.905 2.597 8.21 2.623 ;
      RECT 7.25 2.39 7.255 3.19 ;
      RECT 7.195 2.44 7.225 3.19 ;
      RECT 7.185 2.44 7.19 2.75 ;
      RECT 7.17 2.44 7.175 2.745 ;
      RECT 6.715 2.485 6.73 2.7 ;
      RECT 6.645 2.485 6.73 2.695 ;
      RECT 7.91 2.065 7.98 2.275 ;
      RECT 7.98 2.072 7.99 2.27 ;
      RECT 7.876 2.065 7.91 2.282 ;
      RECT 7.79 2.065 7.876 2.306 ;
      RECT 7.78 2.07 7.79 2.325 ;
      RECT 7.775 2.082 7.78 2.328 ;
      RECT 7.76 2.097 7.775 2.332 ;
      RECT 7.755 2.115 7.76 2.336 ;
      RECT 7.715 2.125 7.755 2.345 ;
      RECT 7.7 2.132 7.715 2.357 ;
      RECT 7.685 2.137 7.7 2.362 ;
      RECT 7.67 2.14 7.685 2.367 ;
      RECT 7.66 2.142 7.67 2.371 ;
      RECT 7.625 2.149 7.66 2.379 ;
      RECT 7.59 2.157 7.625 2.393 ;
      RECT 7.58 2.163 7.59 2.402 ;
      RECT 7.575 2.165 7.58 2.404 ;
      RECT 7.555 2.168 7.575 2.41 ;
      RECT 7.525 2.175 7.555 2.421 ;
      RECT 7.515 2.181 7.525 2.428 ;
      RECT 7.49 2.184 7.515 2.435 ;
      RECT 7.48 2.188 7.49 2.443 ;
      RECT 7.475 2.189 7.48 2.465 ;
      RECT 7.47 2.19 7.475 2.48 ;
      RECT 7.465 2.191 7.47 2.495 ;
      RECT 7.46 2.192 7.465 2.51 ;
      RECT 7.455 2.193 7.46 2.54 ;
      RECT 7.445 2.195 7.455 2.573 ;
      RECT 7.43 2.199 7.445 2.62 ;
      RECT 7.42 2.202 7.43 2.665 ;
      RECT 7.415 2.205 7.42 2.693 ;
      RECT 7.405 2.207 7.415 2.72 ;
      RECT 7.4 2.21 7.405 2.755 ;
      RECT 7.37 2.215 7.4 2.813 ;
      RECT 7.365 2.22 7.37 2.898 ;
      RECT 7.36 2.222 7.365 2.933 ;
      RECT 7.355 2.224 7.36 3.015 ;
      RECT 7.35 2.226 7.355 3.103 ;
      RECT 7.34 2.228 7.35 3.185 ;
      RECT 7.325 2.242 7.34 3.19 ;
      RECT 7.29 2.287 7.325 3.19 ;
      RECT 7.28 2.327 7.29 3.19 ;
      RECT 7.265 2.355 7.28 3.19 ;
      RECT 7.26 2.372 7.265 3.19 ;
      RECT 7.255 2.38 7.26 3.19 ;
      RECT 7.245 2.395 7.25 3.19 ;
      RECT 7.24 2.402 7.245 3.19 ;
      RECT 7.23 2.422 7.24 3.19 ;
      RECT 7.225 2.435 7.23 3.19 ;
      RECT 7.19 2.44 7.195 2.775 ;
      RECT 7.175 2.83 7.195 3.19 ;
      RECT 7.175 2.44 7.185 2.748 ;
      RECT 7.17 2.87 7.175 3.19 ;
      RECT 7.12 2.44 7.17 2.743 ;
      RECT 7.165 2.907 7.17 3.19 ;
      RECT 7.155 2.93 7.165 3.19 ;
      RECT 7.15 2.975 7.155 3.19 ;
      RECT 7.14 2.985 7.15 3.183 ;
      RECT 7.066 2.44 7.12 2.737 ;
      RECT 6.98 2.44 7.066 2.73 ;
      RECT 6.931 2.487 6.98 2.723 ;
      RECT 6.845 2.495 6.931 2.716 ;
      RECT 6.83 2.492 6.845 2.711 ;
      RECT 6.816 2.485 6.83 2.71 ;
      RECT 6.73 2.485 6.816 2.705 ;
      RECT 6.635 2.49 6.645 2.69 ;
      RECT 6.225 1.92 6.24 2.32 ;
      RECT 6.42 1.92 6.425 2.18 ;
      RECT 6.165 1.92 6.21 2.18 ;
      RECT 6.62 3.225 6.625 3.43 ;
      RECT 6.615 3.215 6.62 3.435 ;
      RECT 6.61 3.202 6.615 3.44 ;
      RECT 6.605 3.182 6.61 3.44 ;
      RECT 6.58 3.135 6.605 3.44 ;
      RECT 6.545 3.05 6.58 3.44 ;
      RECT 6.54 2.987 6.545 3.44 ;
      RECT 6.535 2.972 6.54 3.44 ;
      RECT 6.52 2.932 6.535 3.44 ;
      RECT 6.515 2.907 6.52 3.44 ;
      RECT 6.505 2.89 6.515 3.44 ;
      RECT 6.47 2.812 6.505 3.44 ;
      RECT 6.465 2.755 6.47 3.44 ;
      RECT 6.46 2.742 6.465 3.44 ;
      RECT 6.45 2.72 6.46 3.44 ;
      RECT 6.44 2.685 6.45 3.44 ;
      RECT 6.43 2.655 6.44 3.44 ;
      RECT 6.42 2.57 6.43 3.083 ;
      RECT 6.427 3.215 6.43 3.44 ;
      RECT 6.425 3.225 6.427 3.44 ;
      RECT 6.415 3.235 6.425 3.435 ;
      RECT 6.41 1.92 6.42 2.315 ;
      RECT 6.415 2.447 6.42 3.058 ;
      RECT 6.41 2.345 6.415 3.041 ;
      RECT 6.4 1.92 6.41 3.017 ;
      RECT 6.395 1.92 6.4 2.988 ;
      RECT 6.39 1.92 6.395 2.978 ;
      RECT 6.37 1.92 6.39 2.94 ;
      RECT 6.365 1.92 6.37 2.898 ;
      RECT 6.36 1.92 6.365 2.878 ;
      RECT 6.33 1.92 6.36 2.828 ;
      RECT 6.32 1.92 6.33 2.775 ;
      RECT 6.315 1.92 6.32 2.748 ;
      RECT 6.31 1.92 6.315 2.733 ;
      RECT 6.3 1.92 6.31 2.71 ;
      RECT 6.29 1.92 6.3 2.685 ;
      RECT 6.285 1.92 6.29 2.625 ;
      RECT 6.275 1.92 6.285 2.563 ;
      RECT 6.27 1.92 6.275 2.483 ;
      RECT 6.265 1.92 6.27 2.448 ;
      RECT 6.26 1.92 6.265 2.423 ;
      RECT 6.255 1.92 6.26 2.408 ;
      RECT 6.25 1.92 6.255 2.378 ;
      RECT 6.245 1.92 6.25 2.355 ;
      RECT 6.24 1.92 6.245 2.328 ;
      RECT 6.21 1.92 6.225 2.315 ;
      RECT 5.365 3.455 5.55 3.665 ;
      RECT 5.355 3.46 5.565 3.658 ;
      RECT 5.355 3.46 5.585 3.63 ;
      RECT 5.355 3.46 5.6 3.609 ;
      RECT 5.355 3.46 5.615 3.607 ;
      RECT 5.355 3.46 5.625 3.606 ;
      RECT 5.355 3.46 5.655 3.603 ;
      RECT 6.005 3.305 6.265 3.565 ;
      RECT 5.965 3.352 6.265 3.548 ;
      RECT 5.956 3.36 5.965 3.551 ;
      RECT 5.55 3.453 6.265 3.548 ;
      RECT 5.87 3.378 5.956 3.558 ;
      RECT 5.565 3.45 6.265 3.548 ;
      RECT 5.811 3.4 5.87 3.57 ;
      RECT 5.585 3.446 6.265 3.548 ;
      RECT 5.725 3.412 5.811 3.581 ;
      RECT 5.6 3.442 6.265 3.548 ;
      RECT 5.67 3.425 5.725 3.593 ;
      RECT 5.615 3.44 6.265 3.548 ;
      RECT 5.655 3.431 5.67 3.599 ;
      RECT 5.625 3.436 6.265 3.548 ;
      RECT 5.77 2.96 6.03 3.22 ;
      RECT 5.77 2.98 6.14 3.19 ;
      RECT 5.77 2.985 6.15 3.185 ;
      RECT 5.961 2.399 6.04 2.63 ;
      RECT 5.875 2.402 6.09 2.625 ;
      RECT 5.87 2.402 6.09 2.62 ;
      RECT 5.87 2.407 6.1 2.618 ;
      RECT 5.845 2.407 6.1 2.615 ;
      RECT 5.845 2.415 6.11 2.613 ;
      RECT 5.725 2.35 5.985 2.61 ;
      RECT 5.725 2.397 6.035 2.61 ;
      RECT 4.98 2.97 4.985 3.23 ;
      RECT 4.81 2.74 4.815 3.23 ;
      RECT 4.695 2.98 4.7 3.205 ;
      RECT 5.405 2.075 5.41 2.285 ;
      RECT 5.41 2.08 5.425 2.28 ;
      RECT 5.345 2.075 5.405 2.293 ;
      RECT 5.33 2.075 5.345 2.303 ;
      RECT 5.28 2.075 5.33 2.32 ;
      RECT 5.26 2.075 5.28 2.343 ;
      RECT 5.245 2.075 5.26 2.355 ;
      RECT 5.225 2.075 5.245 2.365 ;
      RECT 5.215 2.08 5.225 2.374 ;
      RECT 5.21 2.09 5.215 2.379 ;
      RECT 5.205 2.102 5.21 2.383 ;
      RECT 5.195 2.125 5.205 2.388 ;
      RECT 5.19 2.14 5.195 2.392 ;
      RECT 5.185 2.157 5.19 2.395 ;
      RECT 5.18 2.165 5.185 2.398 ;
      RECT 5.17 2.17 5.18 2.402 ;
      RECT 5.165 2.177 5.17 2.407 ;
      RECT 5.155 2.182 5.165 2.411 ;
      RECT 5.13 2.194 5.155 2.422 ;
      RECT 5.11 2.211 5.13 2.438 ;
      RECT 5.085 2.228 5.11 2.46 ;
      RECT 5.05 2.251 5.085 2.518 ;
      RECT 5.03 2.273 5.05 2.58 ;
      RECT 5.025 2.283 5.03 2.615 ;
      RECT 5.015 2.29 5.025 2.653 ;
      RECT 5.01 2.297 5.015 2.673 ;
      RECT 5.005 2.308 5.01 2.71 ;
      RECT 5 2.316 5.005 2.775 ;
      RECT 4.99 2.327 5 2.828 ;
      RECT 4.985 2.345 4.99 2.898 ;
      RECT 4.98 2.355 4.985 2.935 ;
      RECT 4.975 2.365 4.98 3.23 ;
      RECT 4.97 2.377 4.975 3.23 ;
      RECT 4.965 2.387 4.97 3.23 ;
      RECT 4.955 2.397 4.965 3.23 ;
      RECT 4.945 2.42 4.955 3.23 ;
      RECT 4.93 2.455 4.945 3.23 ;
      RECT 4.89 2.517 4.93 3.23 ;
      RECT 4.885 2.57 4.89 3.23 ;
      RECT 4.86 2.605 4.885 3.23 ;
      RECT 4.845 2.65 4.86 3.23 ;
      RECT 4.84 2.672 4.845 3.23 ;
      RECT 4.83 2.685 4.84 3.23 ;
      RECT 4.82 2.71 4.83 3.23 ;
      RECT 4.815 2.732 4.82 3.23 ;
      RECT 4.79 2.77 4.81 3.23 ;
      RECT 4.75 2.827 4.79 3.23 ;
      RECT 4.745 2.877 4.75 3.23 ;
      RECT 4.74 2.895 4.745 3.23 ;
      RECT 4.735 2.907 4.74 3.23 ;
      RECT 4.725 2.925 4.735 3.23 ;
      RECT 4.715 2.945 4.725 3.205 ;
      RECT 4.71 2.962 4.715 3.205 ;
      RECT 4.7 2.975 4.71 3.205 ;
      RECT 4.67 2.985 4.695 3.205 ;
      RECT 4.66 2.992 4.67 3.205 ;
      RECT 4.645 3.002 4.66 3.2 ;
      RECT 3.025 7.765 3.315 7.995 ;
      RECT 3.085 7.025 3.255 7.995 ;
      RECT 2.995 7.025 3.345 7.315 ;
      RECT 2.62 6.285 2.97 6.575 ;
      RECT 2.48 6.315 2.97 6.485 ;
      RECT 77.535 2.85 77.905 3.22 ;
      RECT 61.75 2.85 62.12 3.22 ;
      RECT 45.965 2.85 46.335 3.22 ;
      RECT 30.19 2.85 30.56 3.22 ;
      RECT 14.41 2.85 14.78 3.22 ;
    LAYER mcon ;
      RECT 82.705 6.32 82.875 6.49 ;
      RECT 82.71 6.315 82.88 6.485 ;
      RECT 66.92 6.32 67.09 6.49 ;
      RECT 66.925 6.315 67.095 6.485 ;
      RECT 51.135 6.32 51.305 6.49 ;
      RECT 51.14 6.315 51.31 6.485 ;
      RECT 35.36 6.32 35.53 6.49 ;
      RECT 35.365 6.315 35.535 6.485 ;
      RECT 19.58 6.32 19.75 6.49 ;
      RECT 19.585 6.315 19.755 6.485 ;
      RECT 82.705 7.8 82.875 7.97 ;
      RECT 82.355 0.1 82.525 0.27 ;
      RECT 82.355 8.61 82.525 8.78 ;
      RECT 82.335 2.76 82.505 2.93 ;
      RECT 82.335 5.95 82.505 6.12 ;
      RECT 81.715 0.91 81.885 1.08 ;
      RECT 81.715 2.39 81.885 2.56 ;
      RECT 81.715 6.32 81.885 6.49 ;
      RECT 81.715 7.8 81.885 7.97 ;
      RECT 81.365 0.1 81.535 0.27 ;
      RECT 81.365 8.61 81.535 8.78 ;
      RECT 81.345 2.76 81.515 2.93 ;
      RECT 81.345 5.95 81.515 6.12 ;
      RECT 80.665 0.105 80.835 0.275 ;
      RECT 80.665 8.605 80.835 8.775 ;
      RECT 80.355 2.025 80.525 2.195 ;
      RECT 80.355 6.685 80.525 6.855 ;
      RECT 79.985 0.105 80.155 0.275 ;
      RECT 79.985 8.605 80.155 8.775 ;
      RECT 79.925 0.915 80.095 1.085 ;
      RECT 79.925 1.655 80.095 1.825 ;
      RECT 79.925 7.055 80.095 7.225 ;
      RECT 79.925 7.795 80.095 7.965 ;
      RECT 79.55 2.395 79.72 2.565 ;
      RECT 79.55 6.315 79.72 6.485 ;
      RECT 79.305 0.105 79.475 0.275 ;
      RECT 79.305 8.605 79.475 8.775 ;
      RECT 78.625 0.105 78.795 0.275 ;
      RECT 78.625 8.605 78.795 8.775 ;
      RECT 77 1.415 77.17 1.585 ;
      RECT 76.63 2.875 76.8 3.045 ;
      RECT 76.54 1.415 76.71 1.585 ;
      RECT 76.31 2.045 76.48 2.215 ;
      RECT 76.165 2.485 76.335 2.655 ;
      RECT 76.08 1.415 76.25 1.585 ;
      RECT 75.885 8.605 76.055 8.775 ;
      RECT 75.62 1.415 75.79 1.585 ;
      RECT 75.575 6.685 75.745 6.855 ;
      RECT 75.555 2.525 75.725 2.695 ;
      RECT 75.21 2.16 75.38 2.33 ;
      RECT 75.205 8.605 75.375 8.775 ;
      RECT 75.2 3.52 75.37 3.69 ;
      RECT 75.16 1.415 75.33 1.585 ;
      RECT 75.145 7.055 75.315 7.225 ;
      RECT 75.145 7.795 75.315 7.965 ;
      RECT 74.785 2.76 74.955 2.93 ;
      RECT 74.77 6.315 74.94 6.485 ;
      RECT 74.7 1.415 74.87 1.585 ;
      RECT 74.525 8.605 74.695 8.775 ;
      RECT 74.435 2.235 74.605 2.405 ;
      RECT 74.255 3.55 74.425 3.72 ;
      RECT 74.24 1.415 74.41 1.585 ;
      RECT 73.975 2.865 74.145 3.035 ;
      RECT 73.845 8.605 74.015 8.775 ;
      RECT 73.78 1.415 73.95 1.585 ;
      RECT 73.655 2.49 73.825 2.66 ;
      RECT 73.32 1.415 73.49 1.585 ;
      RECT 72.965 1.97 73.135 2.14 ;
      RECT 72.89 2.44 73.06 2.61 ;
      RECT 72.86 1.415 73.03 1.585 ;
      RECT 72.4 1.415 72.57 1.585 ;
      RECT 72.04 2.165 72.21 2.335 ;
      RECT 71.94 1.415 72.11 1.585 ;
      RECT 71.7 3.36 71.87 3.53 ;
      RECT 71.665 2.695 71.835 2.865 ;
      RECT 71.48 1.415 71.65 1.585 ;
      RECT 71.055 2.55 71.225 2.72 ;
      RECT 71.02 1.415 71.19 1.585 ;
      RECT 70.985 3.25 71.155 3.42 ;
      RECT 70.925 2.085 71.095 2.255 ;
      RECT 70.56 1.415 70.73 1.585 ;
      RECT 70.285 3 70.455 3.17 ;
      RECT 70.1 1.415 70.27 1.585 ;
      RECT 69.78 2.505 69.95 2.675 ;
      RECT 69.64 1.415 69.81 1.585 ;
      RECT 69.56 3.25 69.73 3.42 ;
      RECT 69.355 2.13 69.525 2.3 ;
      RECT 69.18 1.415 69.35 1.585 ;
      RECT 69.085 3 69.255 3.17 ;
      RECT 69.045 2.43 69.215 2.6 ;
      RECT 68.72 1.415 68.89 1.585 ;
      RECT 68.5 3.475 68.67 3.645 ;
      RECT 68.36 2.095 68.53 2.265 ;
      RECT 68.26 1.415 68.43 1.585 ;
      RECT 67.8 1.415 67.97 1.585 ;
      RECT 67.79 3.015 67.96 3.185 ;
      RECT 66.92 7.8 67.09 7.97 ;
      RECT 66.57 0.1 66.74 0.27 ;
      RECT 66.57 8.61 66.74 8.78 ;
      RECT 66.55 2.76 66.72 2.93 ;
      RECT 66.55 5.95 66.72 6.12 ;
      RECT 65.93 0.91 66.1 1.08 ;
      RECT 65.93 2.39 66.1 2.56 ;
      RECT 65.93 6.32 66.1 6.49 ;
      RECT 65.93 7.8 66.1 7.97 ;
      RECT 65.58 0.1 65.75 0.27 ;
      RECT 65.58 8.61 65.75 8.78 ;
      RECT 65.56 2.76 65.73 2.93 ;
      RECT 65.56 5.95 65.73 6.12 ;
      RECT 64.88 0.105 65.05 0.275 ;
      RECT 64.88 8.605 65.05 8.775 ;
      RECT 64.57 2.025 64.74 2.195 ;
      RECT 64.57 6.685 64.74 6.855 ;
      RECT 64.2 0.105 64.37 0.275 ;
      RECT 64.2 8.605 64.37 8.775 ;
      RECT 64.14 0.915 64.31 1.085 ;
      RECT 64.14 1.655 64.31 1.825 ;
      RECT 64.14 7.055 64.31 7.225 ;
      RECT 64.14 7.795 64.31 7.965 ;
      RECT 63.765 2.395 63.935 2.565 ;
      RECT 63.765 6.315 63.935 6.485 ;
      RECT 63.52 0.105 63.69 0.275 ;
      RECT 63.52 8.605 63.69 8.775 ;
      RECT 62.84 0.105 63.01 0.275 ;
      RECT 62.84 8.605 63.01 8.775 ;
      RECT 61.215 1.415 61.385 1.585 ;
      RECT 60.845 2.875 61.015 3.045 ;
      RECT 60.755 1.415 60.925 1.585 ;
      RECT 60.525 2.045 60.695 2.215 ;
      RECT 60.38 2.485 60.55 2.655 ;
      RECT 60.295 1.415 60.465 1.585 ;
      RECT 60.1 8.605 60.27 8.775 ;
      RECT 59.835 1.415 60.005 1.585 ;
      RECT 59.79 6.685 59.96 6.855 ;
      RECT 59.77 2.525 59.94 2.695 ;
      RECT 59.425 2.16 59.595 2.33 ;
      RECT 59.42 8.605 59.59 8.775 ;
      RECT 59.415 3.52 59.585 3.69 ;
      RECT 59.375 1.415 59.545 1.585 ;
      RECT 59.36 7.055 59.53 7.225 ;
      RECT 59.36 7.795 59.53 7.965 ;
      RECT 59 2.76 59.17 2.93 ;
      RECT 58.985 6.315 59.155 6.485 ;
      RECT 58.915 1.415 59.085 1.585 ;
      RECT 58.74 8.605 58.91 8.775 ;
      RECT 58.65 2.235 58.82 2.405 ;
      RECT 58.47 3.55 58.64 3.72 ;
      RECT 58.455 1.415 58.625 1.585 ;
      RECT 58.19 2.865 58.36 3.035 ;
      RECT 58.06 8.605 58.23 8.775 ;
      RECT 57.995 1.415 58.165 1.585 ;
      RECT 57.87 2.49 58.04 2.66 ;
      RECT 57.535 1.415 57.705 1.585 ;
      RECT 57.18 1.97 57.35 2.14 ;
      RECT 57.105 2.44 57.275 2.61 ;
      RECT 57.075 1.415 57.245 1.585 ;
      RECT 56.615 1.415 56.785 1.585 ;
      RECT 56.255 2.165 56.425 2.335 ;
      RECT 56.155 1.415 56.325 1.585 ;
      RECT 55.915 3.36 56.085 3.53 ;
      RECT 55.88 2.695 56.05 2.865 ;
      RECT 55.695 1.415 55.865 1.585 ;
      RECT 55.27 2.55 55.44 2.72 ;
      RECT 55.235 1.415 55.405 1.585 ;
      RECT 55.2 3.25 55.37 3.42 ;
      RECT 55.14 2.085 55.31 2.255 ;
      RECT 54.775 1.415 54.945 1.585 ;
      RECT 54.5 3 54.67 3.17 ;
      RECT 54.315 1.415 54.485 1.585 ;
      RECT 53.995 2.505 54.165 2.675 ;
      RECT 53.855 1.415 54.025 1.585 ;
      RECT 53.775 3.25 53.945 3.42 ;
      RECT 53.57 2.13 53.74 2.3 ;
      RECT 53.395 1.415 53.565 1.585 ;
      RECT 53.3 3 53.47 3.17 ;
      RECT 53.26 2.43 53.43 2.6 ;
      RECT 52.935 1.415 53.105 1.585 ;
      RECT 52.715 3.475 52.885 3.645 ;
      RECT 52.575 2.095 52.745 2.265 ;
      RECT 52.475 1.415 52.645 1.585 ;
      RECT 52.015 1.415 52.185 1.585 ;
      RECT 52.005 3.015 52.175 3.185 ;
      RECT 51.135 7.8 51.305 7.97 ;
      RECT 50.785 0.1 50.955 0.27 ;
      RECT 50.785 8.61 50.955 8.78 ;
      RECT 50.765 2.76 50.935 2.93 ;
      RECT 50.765 5.95 50.935 6.12 ;
      RECT 50.145 0.91 50.315 1.08 ;
      RECT 50.145 2.39 50.315 2.56 ;
      RECT 50.145 6.32 50.315 6.49 ;
      RECT 50.145 7.8 50.315 7.97 ;
      RECT 49.795 0.1 49.965 0.27 ;
      RECT 49.795 8.61 49.965 8.78 ;
      RECT 49.775 2.76 49.945 2.93 ;
      RECT 49.775 5.95 49.945 6.12 ;
      RECT 49.095 0.105 49.265 0.275 ;
      RECT 49.095 8.605 49.265 8.775 ;
      RECT 48.785 2.025 48.955 2.195 ;
      RECT 48.785 6.685 48.955 6.855 ;
      RECT 48.415 0.105 48.585 0.275 ;
      RECT 48.415 8.605 48.585 8.775 ;
      RECT 48.355 0.915 48.525 1.085 ;
      RECT 48.355 1.655 48.525 1.825 ;
      RECT 48.355 7.055 48.525 7.225 ;
      RECT 48.355 7.795 48.525 7.965 ;
      RECT 47.98 2.395 48.15 2.565 ;
      RECT 47.98 6.315 48.15 6.485 ;
      RECT 47.735 0.105 47.905 0.275 ;
      RECT 47.735 8.605 47.905 8.775 ;
      RECT 47.055 0.105 47.225 0.275 ;
      RECT 47.055 8.605 47.225 8.775 ;
      RECT 45.43 1.415 45.6 1.585 ;
      RECT 45.06 2.875 45.23 3.045 ;
      RECT 44.97 1.415 45.14 1.585 ;
      RECT 44.74 2.045 44.91 2.215 ;
      RECT 44.595 2.485 44.765 2.655 ;
      RECT 44.51 1.415 44.68 1.585 ;
      RECT 44.315 8.605 44.485 8.775 ;
      RECT 44.05 1.415 44.22 1.585 ;
      RECT 44.005 6.685 44.175 6.855 ;
      RECT 43.985 2.525 44.155 2.695 ;
      RECT 43.64 2.16 43.81 2.33 ;
      RECT 43.635 8.605 43.805 8.775 ;
      RECT 43.63 3.52 43.8 3.69 ;
      RECT 43.59 1.415 43.76 1.585 ;
      RECT 43.575 7.055 43.745 7.225 ;
      RECT 43.575 7.795 43.745 7.965 ;
      RECT 43.215 2.76 43.385 2.93 ;
      RECT 43.2 6.315 43.37 6.485 ;
      RECT 43.13 1.415 43.3 1.585 ;
      RECT 42.955 8.605 43.125 8.775 ;
      RECT 42.865 2.235 43.035 2.405 ;
      RECT 42.685 3.55 42.855 3.72 ;
      RECT 42.67 1.415 42.84 1.585 ;
      RECT 42.405 2.865 42.575 3.035 ;
      RECT 42.275 8.605 42.445 8.775 ;
      RECT 42.21 1.415 42.38 1.585 ;
      RECT 42.085 2.49 42.255 2.66 ;
      RECT 41.75 1.415 41.92 1.585 ;
      RECT 41.395 1.97 41.565 2.14 ;
      RECT 41.32 2.44 41.49 2.61 ;
      RECT 41.29 1.415 41.46 1.585 ;
      RECT 40.83 1.415 41 1.585 ;
      RECT 40.47 2.165 40.64 2.335 ;
      RECT 40.37 1.415 40.54 1.585 ;
      RECT 40.13 3.36 40.3 3.53 ;
      RECT 40.095 2.695 40.265 2.865 ;
      RECT 39.91 1.415 40.08 1.585 ;
      RECT 39.485 2.55 39.655 2.72 ;
      RECT 39.45 1.415 39.62 1.585 ;
      RECT 39.415 3.25 39.585 3.42 ;
      RECT 39.355 2.085 39.525 2.255 ;
      RECT 38.99 1.415 39.16 1.585 ;
      RECT 38.715 3 38.885 3.17 ;
      RECT 38.53 1.415 38.7 1.585 ;
      RECT 38.21 2.505 38.38 2.675 ;
      RECT 38.07 1.415 38.24 1.585 ;
      RECT 37.99 3.25 38.16 3.42 ;
      RECT 37.785 2.13 37.955 2.3 ;
      RECT 37.61 1.415 37.78 1.585 ;
      RECT 37.515 3 37.685 3.17 ;
      RECT 37.475 2.43 37.645 2.6 ;
      RECT 37.15 1.415 37.32 1.585 ;
      RECT 36.93 3.475 37.1 3.645 ;
      RECT 36.79 2.095 36.96 2.265 ;
      RECT 36.69 1.415 36.86 1.585 ;
      RECT 36.23 1.415 36.4 1.585 ;
      RECT 36.22 3.015 36.39 3.185 ;
      RECT 35.36 7.8 35.53 7.97 ;
      RECT 35.01 0.1 35.18 0.27 ;
      RECT 35.01 8.61 35.18 8.78 ;
      RECT 34.99 2.76 35.16 2.93 ;
      RECT 34.99 5.95 35.16 6.12 ;
      RECT 34.37 0.91 34.54 1.08 ;
      RECT 34.37 2.39 34.54 2.56 ;
      RECT 34.37 6.32 34.54 6.49 ;
      RECT 34.37 7.8 34.54 7.97 ;
      RECT 34.02 0.1 34.19 0.27 ;
      RECT 34.02 8.61 34.19 8.78 ;
      RECT 34 2.76 34.17 2.93 ;
      RECT 34 5.95 34.17 6.12 ;
      RECT 33.32 0.105 33.49 0.275 ;
      RECT 33.32 8.605 33.49 8.775 ;
      RECT 33.01 2.025 33.18 2.195 ;
      RECT 33.01 6.685 33.18 6.855 ;
      RECT 32.64 0.105 32.81 0.275 ;
      RECT 32.64 8.605 32.81 8.775 ;
      RECT 32.58 0.915 32.75 1.085 ;
      RECT 32.58 1.655 32.75 1.825 ;
      RECT 32.58 7.055 32.75 7.225 ;
      RECT 32.58 7.795 32.75 7.965 ;
      RECT 32.205 2.395 32.375 2.565 ;
      RECT 32.205 6.315 32.375 6.485 ;
      RECT 31.96 0.105 32.13 0.275 ;
      RECT 31.96 8.605 32.13 8.775 ;
      RECT 31.28 0.105 31.45 0.275 ;
      RECT 31.28 8.605 31.45 8.775 ;
      RECT 29.655 1.415 29.825 1.585 ;
      RECT 29.285 2.875 29.455 3.045 ;
      RECT 29.195 1.415 29.365 1.585 ;
      RECT 28.965 2.045 29.135 2.215 ;
      RECT 28.82 2.485 28.99 2.655 ;
      RECT 28.735 1.415 28.905 1.585 ;
      RECT 28.54 8.605 28.71 8.775 ;
      RECT 28.275 1.415 28.445 1.585 ;
      RECT 28.23 6.685 28.4 6.855 ;
      RECT 28.21 2.525 28.38 2.695 ;
      RECT 27.865 2.16 28.035 2.33 ;
      RECT 27.86 8.605 28.03 8.775 ;
      RECT 27.855 3.52 28.025 3.69 ;
      RECT 27.815 1.415 27.985 1.585 ;
      RECT 27.8 7.055 27.97 7.225 ;
      RECT 27.8 7.795 27.97 7.965 ;
      RECT 27.44 2.76 27.61 2.93 ;
      RECT 27.425 6.315 27.595 6.485 ;
      RECT 27.355 1.415 27.525 1.585 ;
      RECT 27.18 8.605 27.35 8.775 ;
      RECT 27.09 2.235 27.26 2.405 ;
      RECT 26.91 3.55 27.08 3.72 ;
      RECT 26.895 1.415 27.065 1.585 ;
      RECT 26.63 2.865 26.8 3.035 ;
      RECT 26.5 8.605 26.67 8.775 ;
      RECT 26.435 1.415 26.605 1.585 ;
      RECT 26.31 2.49 26.48 2.66 ;
      RECT 25.975 1.415 26.145 1.585 ;
      RECT 25.62 1.97 25.79 2.14 ;
      RECT 25.545 2.44 25.715 2.61 ;
      RECT 25.515 1.415 25.685 1.585 ;
      RECT 25.055 1.415 25.225 1.585 ;
      RECT 24.695 2.165 24.865 2.335 ;
      RECT 24.595 1.415 24.765 1.585 ;
      RECT 24.355 3.36 24.525 3.53 ;
      RECT 24.32 2.695 24.49 2.865 ;
      RECT 24.135 1.415 24.305 1.585 ;
      RECT 23.71 2.55 23.88 2.72 ;
      RECT 23.675 1.415 23.845 1.585 ;
      RECT 23.64 3.25 23.81 3.42 ;
      RECT 23.58 2.085 23.75 2.255 ;
      RECT 23.215 1.415 23.385 1.585 ;
      RECT 22.94 3 23.11 3.17 ;
      RECT 22.755 1.415 22.925 1.585 ;
      RECT 22.435 2.505 22.605 2.675 ;
      RECT 22.295 1.415 22.465 1.585 ;
      RECT 22.215 3.25 22.385 3.42 ;
      RECT 22.01 2.13 22.18 2.3 ;
      RECT 21.835 1.415 22.005 1.585 ;
      RECT 21.74 3 21.91 3.17 ;
      RECT 21.7 2.43 21.87 2.6 ;
      RECT 21.375 1.415 21.545 1.585 ;
      RECT 21.155 3.475 21.325 3.645 ;
      RECT 21.015 2.095 21.185 2.265 ;
      RECT 20.915 1.415 21.085 1.585 ;
      RECT 20.455 1.415 20.625 1.585 ;
      RECT 20.445 3.015 20.615 3.185 ;
      RECT 19.58 7.8 19.75 7.97 ;
      RECT 19.23 0.1 19.4 0.27 ;
      RECT 19.23 8.61 19.4 8.78 ;
      RECT 19.21 2.76 19.38 2.93 ;
      RECT 19.21 5.95 19.38 6.12 ;
      RECT 18.59 0.91 18.76 1.08 ;
      RECT 18.59 2.39 18.76 2.56 ;
      RECT 18.59 6.32 18.76 6.49 ;
      RECT 18.59 7.8 18.76 7.97 ;
      RECT 18.24 0.1 18.41 0.27 ;
      RECT 18.24 8.61 18.41 8.78 ;
      RECT 18.22 2.76 18.39 2.93 ;
      RECT 18.22 5.95 18.39 6.12 ;
      RECT 17.54 0.105 17.71 0.275 ;
      RECT 17.54 8.605 17.71 8.775 ;
      RECT 17.23 2.025 17.4 2.195 ;
      RECT 17.23 6.685 17.4 6.855 ;
      RECT 16.86 0.105 17.03 0.275 ;
      RECT 16.86 8.605 17.03 8.775 ;
      RECT 16.8 0.915 16.97 1.085 ;
      RECT 16.8 1.655 16.97 1.825 ;
      RECT 16.8 7.055 16.97 7.225 ;
      RECT 16.8 7.795 16.97 7.965 ;
      RECT 16.425 2.395 16.595 2.565 ;
      RECT 16.425 6.315 16.595 6.485 ;
      RECT 16.18 0.105 16.35 0.275 ;
      RECT 16.18 8.605 16.35 8.775 ;
      RECT 15.5 0.105 15.67 0.275 ;
      RECT 15.5 8.605 15.67 8.775 ;
      RECT 13.875 1.415 14.045 1.585 ;
      RECT 13.505 2.875 13.675 3.045 ;
      RECT 13.415 1.415 13.585 1.585 ;
      RECT 13.185 2.045 13.355 2.215 ;
      RECT 13.04 2.485 13.21 2.655 ;
      RECT 12.955 1.415 13.125 1.585 ;
      RECT 12.76 8.605 12.93 8.775 ;
      RECT 12.495 1.415 12.665 1.585 ;
      RECT 12.45 6.685 12.62 6.855 ;
      RECT 12.43 2.525 12.6 2.695 ;
      RECT 12.085 2.16 12.255 2.33 ;
      RECT 12.08 8.605 12.25 8.775 ;
      RECT 12.075 3.52 12.245 3.69 ;
      RECT 12.035 1.415 12.205 1.585 ;
      RECT 12.02 7.055 12.19 7.225 ;
      RECT 12.02 7.795 12.19 7.965 ;
      RECT 11.66 2.76 11.83 2.93 ;
      RECT 11.645 6.315 11.815 6.485 ;
      RECT 11.575 1.415 11.745 1.585 ;
      RECT 11.4 8.605 11.57 8.775 ;
      RECT 11.31 2.235 11.48 2.405 ;
      RECT 11.13 3.55 11.3 3.72 ;
      RECT 11.115 1.415 11.285 1.585 ;
      RECT 10.85 2.865 11.02 3.035 ;
      RECT 10.72 8.605 10.89 8.775 ;
      RECT 10.655 1.415 10.825 1.585 ;
      RECT 10.53 2.49 10.7 2.66 ;
      RECT 10.195 1.415 10.365 1.585 ;
      RECT 9.84 1.97 10.01 2.14 ;
      RECT 9.765 2.44 9.935 2.61 ;
      RECT 9.735 1.415 9.905 1.585 ;
      RECT 9.275 1.415 9.445 1.585 ;
      RECT 8.915 2.165 9.085 2.335 ;
      RECT 8.815 1.415 8.985 1.585 ;
      RECT 8.575 3.36 8.745 3.53 ;
      RECT 8.54 2.695 8.71 2.865 ;
      RECT 8.355 1.415 8.525 1.585 ;
      RECT 7.93 2.55 8.1 2.72 ;
      RECT 7.895 1.415 8.065 1.585 ;
      RECT 7.86 3.25 8.03 3.42 ;
      RECT 7.8 2.085 7.97 2.255 ;
      RECT 7.435 1.415 7.605 1.585 ;
      RECT 7.16 3 7.33 3.17 ;
      RECT 6.975 1.415 7.145 1.585 ;
      RECT 6.655 2.505 6.825 2.675 ;
      RECT 6.515 1.415 6.685 1.585 ;
      RECT 6.435 3.25 6.605 3.42 ;
      RECT 6.23 2.13 6.4 2.3 ;
      RECT 6.055 1.415 6.225 1.585 ;
      RECT 5.96 3 6.13 3.17 ;
      RECT 5.92 2.43 6.09 2.6 ;
      RECT 5.595 1.415 5.765 1.585 ;
      RECT 5.375 3.475 5.545 3.645 ;
      RECT 5.235 2.095 5.405 2.265 ;
      RECT 5.135 1.415 5.305 1.585 ;
      RECT 4.675 1.415 4.845 1.585 ;
      RECT 4.665 3.015 4.835 3.185 ;
      RECT 3.825 8.605 3.995 8.775 ;
      RECT 3.145 8.605 3.315 8.775 ;
      RECT 3.085 7.055 3.255 7.225 ;
      RECT 3.085 7.795 3.255 7.965 ;
      RECT 2.71 6.315 2.88 6.485 ;
      RECT 2.465 8.605 2.635 8.775 ;
      RECT 1.785 8.605 1.955 8.775 ;
    LAYER li1 ;
      RECT 75.785 0 75.955 2.085 ;
      RECT 73.825 0 73.995 2.085 ;
      RECT 71.385 0 71.555 2.085 ;
      RECT 70.425 0 70.595 2.085 ;
      RECT 69.905 0 70.075 2.085 ;
      RECT 68.945 0 69.115 2.085 ;
      RECT 67.985 0 68.155 2.085 ;
      RECT 60 0 60.17 2.085 ;
      RECT 58.04 0 58.21 2.085 ;
      RECT 55.6 0 55.77 2.085 ;
      RECT 54.64 0 54.81 2.085 ;
      RECT 54.12 0 54.29 2.085 ;
      RECT 53.16 0 53.33 2.085 ;
      RECT 52.2 0 52.37 2.085 ;
      RECT 44.215 0 44.385 2.085 ;
      RECT 42.255 0 42.425 2.085 ;
      RECT 39.815 0 39.985 2.085 ;
      RECT 38.855 0 39.025 2.085 ;
      RECT 38.335 0 38.505 2.085 ;
      RECT 37.375 0 37.545 2.085 ;
      RECT 36.415 0 36.585 2.085 ;
      RECT 28.44 0 28.61 2.085 ;
      RECT 26.48 0 26.65 2.085 ;
      RECT 24.04 0 24.21 2.085 ;
      RECT 23.08 0 23.25 2.085 ;
      RECT 22.56 0 22.73 2.085 ;
      RECT 21.6 0 21.77 2.085 ;
      RECT 20.64 0 20.81 2.085 ;
      RECT 12.66 0 12.83 2.085 ;
      RECT 10.7 0 10.87 2.085 ;
      RECT 8.26 0 8.43 2.085 ;
      RECT 7.3 0 7.47 2.085 ;
      RECT 6.78 0 6.95 2.085 ;
      RECT 5.82 0 5.99 2.085 ;
      RECT 4.86 0 5.03 2.085 ;
      RECT 67.77 0 77.37 1.59 ;
      RECT 51.985 0 61.585 1.59 ;
      RECT 36.2 0 45.8 1.59 ;
      RECT 20.425 0 30.025 1.59 ;
      RECT 4.645 0 14.245 1.59 ;
      RECT 67.655 1.415 77.485 1.585 ;
      RECT 67.77 0 77.485 1.585 ;
      RECT 51.87 1.415 61.7 1.585 ;
      RECT 51.985 0 61.7 1.585 ;
      RECT 36.085 1.415 45.915 1.585 ;
      RECT 36.2 0 45.915 1.585 ;
      RECT 20.31 1.415 30.14 1.585 ;
      RECT 20.425 0 30.14 1.585 ;
      RECT 4.53 1.415 14.36 1.585 ;
      RECT 4.645 0 14.36 1.585 ;
      RECT 78.545 0 78.715 0.935 ;
      RECT 62.76 0 62.93 0.935 ;
      RECT 46.975 0 47.145 0.935 ;
      RECT 31.2 0 31.37 0.935 ;
      RECT 15.42 0 15.59 0.935 ;
      RECT 82.275 0 82.445 0.93 ;
      RECT 81.285 0 81.455 0.93 ;
      RECT 66.49 0 66.66 0.93 ;
      RECT 65.5 0 65.67 0.93 ;
      RECT 50.705 0 50.875 0.93 ;
      RECT 49.715 0 49.885 0.93 ;
      RECT 34.93 0 35.1 0.93 ;
      RECT 33.94 0 34.11 0.93 ;
      RECT 19.15 0 19.32 0.93 ;
      RECT 18.16 0 18.33 0.93 ;
      RECT 83.07 0 83.25 0.305 ;
      RECT 67.285 0 81.12 0.305 ;
      RECT 51.5 0 65.335 0.305 ;
      RECT 35.725 0 49.55 0.305 ;
      RECT 19.945 0 33.775 0.305 ;
      RECT 1.485 0 17.995 0.305 ;
      RECT 1.485 0 83.25 0.3 ;
      RECT 1.485 8.58 83.25 8.88 ;
      RECT 83.07 8.575 83.25 8.88 ;
      RECT 82.275 7.95 82.445 8.88 ;
      RECT 81.285 7.95 81.455 8.88 ;
      RECT 67.285 8.575 81.12 8.88 ;
      RECT 66.49 7.95 66.66 8.88 ;
      RECT 65.5 7.95 65.67 8.88 ;
      RECT 51.5 8.575 65.335 8.88 ;
      RECT 50.705 7.95 50.875 8.88 ;
      RECT 49.715 7.95 49.885 8.88 ;
      RECT 35.725 8.575 49.55 8.88 ;
      RECT 34.93 7.95 35.1 8.88 ;
      RECT 33.94 7.95 34.11 8.88 ;
      RECT 19.945 8.575 33.775 8.88 ;
      RECT 19.15 7.95 19.32 8.88 ;
      RECT 18.16 7.95 18.33 8.88 ;
      RECT 1.485 8.575 17.995 8.88 ;
      RECT 78.545 7.945 78.715 8.88 ;
      RECT 73.765 7.945 73.935 8.88 ;
      RECT 62.76 7.945 62.93 8.88 ;
      RECT 57.98 7.945 58.15 8.88 ;
      RECT 46.975 7.945 47.145 8.88 ;
      RECT 42.195 7.945 42.365 8.88 ;
      RECT 31.2 7.945 31.37 8.88 ;
      RECT 26.42 7.945 26.59 8.88 ;
      RECT 15.42 7.945 15.59 8.88 ;
      RECT 10.64 7.945 10.81 8.88 ;
      RECT 1.705 7.945 1.875 8.88 ;
      RECT 82.705 5.02 82.875 6.49 ;
      RECT 82.705 6.315 82.88 6.485 ;
      RECT 82.335 1.74 82.505 2.93 ;
      RECT 82.335 1.74 82.805 1.91 ;
      RECT 82.335 6.97 82.805 7.14 ;
      RECT 82.335 5.95 82.505 7.14 ;
      RECT 81.345 1.74 81.515 2.93 ;
      RECT 81.345 1.74 81.815 1.91 ;
      RECT 81.345 6.97 81.815 7.14 ;
      RECT 81.345 5.95 81.515 7.14 ;
      RECT 79.495 2.635 79.665 3.865 ;
      RECT 79.55 0.855 79.72 2.805 ;
      RECT 79.495 0.575 79.665 1.025 ;
      RECT 79.495 7.855 79.665 8.305 ;
      RECT 79.55 6.075 79.72 8.025 ;
      RECT 79.495 5.015 79.665 6.245 ;
      RECT 78.975 0.575 79.145 3.865 ;
      RECT 78.975 2.075 79.38 2.405 ;
      RECT 78.975 1.235 79.38 1.565 ;
      RECT 78.975 5.015 79.145 8.305 ;
      RECT 78.975 7.315 79.38 7.645 ;
      RECT 78.975 6.475 79.38 6.805 ;
      RECT 76.31 1.975 77.04 2.215 ;
      RECT 76.852 1.77 77.04 2.215 ;
      RECT 76.68 1.782 77.055 2.209 ;
      RECT 76.595 1.797 77.075 2.194 ;
      RECT 76.595 1.812 77.08 2.184 ;
      RECT 76.55 1.832 77.095 2.176 ;
      RECT 76.527 1.867 77.11 2.13 ;
      RECT 76.441 1.89 77.115 2.09 ;
      RECT 76.441 1.908 77.125 2.06 ;
      RECT 76.31 1.977 77.13 2.023 ;
      RECT 76.355 1.92 77.125 2.06 ;
      RECT 76.441 1.872 77.11 2.13 ;
      RECT 76.527 1.841 77.095 2.176 ;
      RECT 76.55 1.822 77.08 2.184 ;
      RECT 76.595 1.795 77.055 2.209 ;
      RECT 76.68 1.777 77.04 2.215 ;
      RECT 76.766 1.771 77.04 2.215 ;
      RECT 76.852 1.766 76.985 2.215 ;
      RECT 76.938 1.761 76.985 2.215 ;
      RECT 76.63 2.659 76.8 3.045 ;
      RECT 76.625 2.659 76.8 3.04 ;
      RECT 76.6 2.659 76.8 3.005 ;
      RECT 76.6 2.687 76.81 2.995 ;
      RECT 76.58 2.687 76.81 2.955 ;
      RECT 76.575 2.687 76.81 2.928 ;
      RECT 76.575 2.705 76.815 2.92 ;
      RECT 76.52 2.705 76.815 2.855 ;
      RECT 76.52 2.722 76.825 2.838 ;
      RECT 76.51 2.722 76.825 2.778 ;
      RECT 76.51 2.739 76.83 2.775 ;
      RECT 76.505 2.575 76.675 2.753 ;
      RECT 76.505 2.609 76.761 2.753 ;
      RECT 76.5 3.375 76.505 3.388 ;
      RECT 76.495 3.27 76.5 3.393 ;
      RECT 76.47 3.13 76.495 3.408 ;
      RECT 76.435 3.081 76.47 3.44 ;
      RECT 76.43 3.049 76.435 3.46 ;
      RECT 76.425 3.04 76.43 3.46 ;
      RECT 76.345 3.005 76.425 3.46 ;
      RECT 76.282 2.975 76.345 3.46 ;
      RECT 76.196 2.963 76.282 3.46 ;
      RECT 76.11 2.949 76.196 3.46 ;
      RECT 76.03 2.936 76.11 3.446 ;
      RECT 75.995 2.928 76.03 3.426 ;
      RECT 75.985 2.925 75.995 3.417 ;
      RECT 75.955 2.92 75.985 3.404 ;
      RECT 75.905 2.895 75.955 3.38 ;
      RECT 75.891 2.869 75.905 3.362 ;
      RECT 75.805 2.829 75.891 3.338 ;
      RECT 75.76 2.777 75.805 3.307 ;
      RECT 75.75 2.752 75.76 3.294 ;
      RECT 75.745 2.533 75.75 2.555 ;
      RECT 75.74 2.735 75.75 3.29 ;
      RECT 75.74 2.531 75.745 2.645 ;
      RECT 75.73 2.527 75.74 3.286 ;
      RECT 75.686 2.525 75.73 3.274 ;
      RECT 75.6 2.525 75.686 3.245 ;
      RECT 75.57 2.525 75.6 3.218 ;
      RECT 75.555 2.525 75.57 3.206 ;
      RECT 75.515 2.537 75.555 3.191 ;
      RECT 75.495 2.556 75.515 3.17 ;
      RECT 75.485 2.566 75.495 3.154 ;
      RECT 75.475 2.572 75.485 3.143 ;
      RECT 75.455 2.582 75.475 3.126 ;
      RECT 75.45 2.591 75.455 3.113 ;
      RECT 75.445 2.595 75.45 3.063 ;
      RECT 75.435 2.601 75.445 2.98 ;
      RECT 75.43 2.605 75.435 2.894 ;
      RECT 75.425 2.625 75.43 2.831 ;
      RECT 75.42 2.648 75.425 2.778 ;
      RECT 75.415 2.666 75.42 2.723 ;
      RECT 76.025 2.485 76.195 2.745 ;
      RECT 76.195 2.45 76.24 2.731 ;
      RECT 76.156 2.452 76.245 2.714 ;
      RECT 76.045 2.469 76.331 2.685 ;
      RECT 76.045 2.484 76.335 2.657 ;
      RECT 76.045 2.465 76.245 2.714 ;
      RECT 76.07 2.453 76.195 2.745 ;
      RECT 76.156 2.451 76.24 2.731 ;
      RECT 75.21 1.84 75.38 2.33 ;
      RECT 75.21 1.84 75.415 2.31 ;
      RECT 75.345 1.76 75.455 2.27 ;
      RECT 75.326 1.764 75.475 2.24 ;
      RECT 75.24 1.772 75.495 2.223 ;
      RECT 75.24 1.778 75.5 2.213 ;
      RECT 75.24 1.787 75.52 2.201 ;
      RECT 75.215 1.812 75.55 2.179 ;
      RECT 75.215 1.832 75.555 2.159 ;
      RECT 75.21 1.845 75.565 2.139 ;
      RECT 75.21 1.912 75.57 2.12 ;
      RECT 75.21 2.045 75.575 2.107 ;
      RECT 75.205 1.85 75.565 1.94 ;
      RECT 75.215 1.807 75.52 2.201 ;
      RECT 75.326 1.762 75.455 2.27 ;
      RECT 75.2 3.515 75.5 3.77 ;
      RECT 75.285 3.481 75.5 3.77 ;
      RECT 75.285 3.484 75.505 3.63 ;
      RECT 75.22 3.505 75.505 3.63 ;
      RECT 75.255 3.495 75.5 3.77 ;
      RECT 75.25 3.5 75.505 3.63 ;
      RECT 75.285 3.479 75.486 3.77 ;
      RECT 75.371 3.47 75.486 3.77 ;
      RECT 75.371 3.464 75.4 3.77 ;
      RECT 74.86 3.105 74.87 3.595 ;
      RECT 74.52 3.04 74.53 3.34 ;
      RECT 75.035 3.212 75.04 3.431 ;
      RECT 75.025 3.192 75.035 3.448 ;
      RECT 75.015 3.172 75.025 3.478 ;
      RECT 75.01 3.162 75.015 3.493 ;
      RECT 75.005 3.158 75.01 3.498 ;
      RECT 74.99 3.15 75.005 3.505 ;
      RECT 74.95 3.13 74.99 3.53 ;
      RECT 74.925 3.112 74.95 3.563 ;
      RECT 74.92 3.11 74.925 3.576 ;
      RECT 74.9 3.107 74.92 3.58 ;
      RECT 74.87 3.105 74.9 3.59 ;
      RECT 74.8 3.107 74.86 3.591 ;
      RECT 74.78 3.107 74.8 3.585 ;
      RECT 74.755 3.105 74.78 3.582 ;
      RECT 74.72 3.1 74.755 3.578 ;
      RECT 74.7 3.094 74.72 3.565 ;
      RECT 74.69 3.091 74.7 3.553 ;
      RECT 74.67 3.088 74.69 3.538 ;
      RECT 74.65 3.084 74.67 3.52 ;
      RECT 74.645 3.081 74.65 3.51 ;
      RECT 74.64 3.08 74.645 3.508 ;
      RECT 74.63 3.077 74.64 3.5 ;
      RECT 74.62 3.071 74.63 3.483 ;
      RECT 74.61 3.065 74.62 3.465 ;
      RECT 74.6 3.059 74.61 3.453 ;
      RECT 74.59 3.053 74.6 3.433 ;
      RECT 74.585 3.049 74.59 3.418 ;
      RECT 74.58 3.047 74.585 3.41 ;
      RECT 74.575 3.045 74.58 3.403 ;
      RECT 74.57 3.043 74.575 3.393 ;
      RECT 74.565 3.041 74.57 3.387 ;
      RECT 74.555 3.04 74.565 3.377 ;
      RECT 74.545 3.04 74.555 3.368 ;
      RECT 74.53 3.04 74.545 3.353 ;
      RECT 74.49 3.04 74.52 3.337 ;
      RECT 74.47 3.042 74.49 3.332 ;
      RECT 74.465 3.047 74.47 3.33 ;
      RECT 74.435 3.055 74.465 3.328 ;
      RECT 74.405 3.07 74.435 3.327 ;
      RECT 74.36 3.092 74.405 3.332 ;
      RECT 74.355 3.107 74.36 3.336 ;
      RECT 74.34 3.112 74.355 3.338 ;
      RECT 74.335 3.116 74.34 3.34 ;
      RECT 74.275 3.139 74.335 3.349 ;
      RECT 74.255 3.165 74.275 3.362 ;
      RECT 74.245 3.172 74.255 3.366 ;
      RECT 74.23 3.179 74.245 3.369 ;
      RECT 74.21 3.189 74.23 3.372 ;
      RECT 74.205 3.197 74.21 3.375 ;
      RECT 74.16 3.202 74.205 3.382 ;
      RECT 74.15 3.205 74.16 3.389 ;
      RECT 74.14 3.205 74.15 3.393 ;
      RECT 74.105 3.207 74.14 3.405 ;
      RECT 74.085 3.21 74.105 3.418 ;
      RECT 74.045 3.213 74.085 3.429 ;
      RECT 74.03 3.215 74.045 3.442 ;
      RECT 74.02 3.215 74.03 3.447 ;
      RECT 73.995 3.216 74.02 3.455 ;
      RECT 73.985 3.218 73.995 3.46 ;
      RECT 73.98 3.219 73.985 3.463 ;
      RECT 73.955 3.217 73.98 3.466 ;
      RECT 73.94 3.215 73.955 3.467 ;
      RECT 73.92 3.212 73.94 3.469 ;
      RECT 73.9 3.207 73.92 3.469 ;
      RECT 73.84 3.202 73.9 3.466 ;
      RECT 73.805 3.177 73.84 3.462 ;
      RECT 73.795 3.154 73.805 3.46 ;
      RECT 73.765 3.131 73.795 3.46 ;
      RECT 73.755 3.11 73.765 3.46 ;
      RECT 73.73 3.092 73.755 3.458 ;
      RECT 73.715 3.07 73.73 3.455 ;
      RECT 73.7 3.052 73.715 3.453 ;
      RECT 73.68 3.042 73.7 3.451 ;
      RECT 73.665 3.037 73.68 3.45 ;
      RECT 73.65 3.035 73.665 3.449 ;
      RECT 73.62 3.036 73.65 3.447 ;
      RECT 73.6 3.039 73.62 3.445 ;
      RECT 73.543 3.043 73.6 3.445 ;
      RECT 73.457 3.052 73.543 3.445 ;
      RECT 73.371 3.063 73.457 3.445 ;
      RECT 73.285 3.074 73.371 3.445 ;
      RECT 73.265 3.081 73.285 3.453 ;
      RECT 73.255 3.084 73.265 3.46 ;
      RECT 73.19 3.089 73.255 3.478 ;
      RECT 73.16 3.096 73.19 3.503 ;
      RECT 73.15 3.099 73.16 3.51 ;
      RECT 73.105 3.103 73.15 3.515 ;
      RECT 73.075 3.108 73.105 3.52 ;
      RECT 73.074 3.11 73.075 3.52 ;
      RECT 72.988 3.116 73.074 3.52 ;
      RECT 72.902 3.127 72.988 3.52 ;
      RECT 72.816 3.139 72.902 3.52 ;
      RECT 72.73 3.15 72.816 3.52 ;
      RECT 72.715 3.157 72.73 3.515 ;
      RECT 72.71 3.159 72.715 3.509 ;
      RECT 72.69 3.17 72.71 3.504 ;
      RECT 72.68 3.188 72.69 3.498 ;
      RECT 72.675 3.2 72.68 3.298 ;
      RECT 74.97 1.953 74.99 2.04 ;
      RECT 74.965 1.888 74.97 2.072 ;
      RECT 74.955 1.855 74.965 2.077 ;
      RECT 74.95 1.835 74.955 2.083 ;
      RECT 74.92 1.835 74.95 2.1 ;
      RECT 74.871 1.835 74.92 2.136 ;
      RECT 74.785 1.835 74.871 2.194 ;
      RECT 74.756 1.845 74.785 2.243 ;
      RECT 74.67 1.887 74.756 2.296 ;
      RECT 74.65 1.925 74.67 2.343 ;
      RECT 74.625 1.942 74.65 2.363 ;
      RECT 74.615 1.956 74.625 2.383 ;
      RECT 74.61 1.962 74.615 2.393 ;
      RECT 74.605 1.966 74.61 2.4 ;
      RECT 74.555 1.986 74.605 2.405 ;
      RECT 74.49 2.03 74.555 2.405 ;
      RECT 74.465 2.08 74.49 2.405 ;
      RECT 74.455 2.11 74.465 2.405 ;
      RECT 74.45 2.137 74.455 2.405 ;
      RECT 74.445 2.155 74.45 2.405 ;
      RECT 74.435 2.197 74.445 2.405 ;
      RECT 74.785 2.755 74.955 2.93 ;
      RECT 74.725 2.583 74.785 2.918 ;
      RECT 74.715 2.576 74.725 2.901 ;
      RECT 74.67 2.755 74.955 2.881 ;
      RECT 74.651 2.755 74.955 2.859 ;
      RECT 74.565 2.755 74.955 2.824 ;
      RECT 74.545 2.575 74.715 2.78 ;
      RECT 74.545 2.722 74.95 2.78 ;
      RECT 74.545 2.67 74.925 2.78 ;
      RECT 74.545 2.625 74.89 2.78 ;
      RECT 74.545 2.607 74.855 2.78 ;
      RECT 74.545 2.597 74.85 2.78 ;
      RECT 74.715 7.855 74.885 8.305 ;
      RECT 74.77 6.075 74.94 8.025 ;
      RECT 74.715 5.015 74.885 6.245 ;
      RECT 74.195 5.015 74.365 8.305 ;
      RECT 74.195 7.315 74.6 7.645 ;
      RECT 74.195 6.475 74.6 6.805 ;
      RECT 74.265 3.555 74.455 3.78 ;
      RECT 74.255 3.556 74.46 3.775 ;
      RECT 74.255 3.558 74.47 3.755 ;
      RECT 74.255 3.562 74.475 3.74 ;
      RECT 74.255 3.549 74.425 3.775 ;
      RECT 74.255 3.552 74.45 3.775 ;
      RECT 74.265 3.548 74.425 3.78 ;
      RECT 74.351 3.546 74.425 3.78 ;
      RECT 73.975 2.797 74.145 3.035 ;
      RECT 73.975 2.797 74.231 2.949 ;
      RECT 73.975 2.797 74.235 2.859 ;
      RECT 74.025 2.57 74.245 2.838 ;
      RECT 74.02 2.587 74.25 2.811 ;
      RECT 73.985 2.745 74.25 2.811 ;
      RECT 74.005 2.595 74.145 3.035 ;
      RECT 73.995 2.677 74.255 2.794 ;
      RECT 73.99 2.725 74.255 2.794 ;
      RECT 73.995 2.635 74.25 2.811 ;
      RECT 74.02 2.572 74.245 2.838 ;
      RECT 73.585 2.547 73.755 2.745 ;
      RECT 73.585 2.547 73.8 2.72 ;
      RECT 73.655 2.49 73.825 2.678 ;
      RECT 73.63 2.505 73.825 2.678 ;
      RECT 73.245 2.551 73.275 2.745 ;
      RECT 73.24 2.523 73.245 2.745 ;
      RECT 73.21 2.497 73.24 2.747 ;
      RECT 73.185 2.455 73.21 2.75 ;
      RECT 73.175 2.427 73.185 2.752 ;
      RECT 73.14 2.407 73.175 2.754 ;
      RECT 73.075 2.392 73.14 2.76 ;
      RECT 73.025 2.39 73.075 2.766 ;
      RECT 73.002 2.392 73.025 2.771 ;
      RECT 72.916 2.403 73.002 2.777 ;
      RECT 72.83 2.421 72.916 2.787 ;
      RECT 72.815 2.432 72.83 2.793 ;
      RECT 72.745 2.455 72.815 2.799 ;
      RECT 72.69 2.487 72.745 2.807 ;
      RECT 72.65 2.51 72.69 2.813 ;
      RECT 72.636 2.523 72.65 2.816 ;
      RECT 72.55 2.545 72.636 2.822 ;
      RECT 72.535 2.57 72.55 2.828 ;
      RECT 72.495 2.585 72.535 2.832 ;
      RECT 72.445 2.6 72.495 2.837 ;
      RECT 72.42 2.607 72.445 2.841 ;
      RECT 72.36 2.602 72.42 2.845 ;
      RECT 72.345 2.593 72.36 2.849 ;
      RECT 72.275 2.583 72.345 2.845 ;
      RECT 72.25 2.575 72.27 2.835 ;
      RECT 72.191 2.575 72.25 2.813 ;
      RECT 72.105 2.575 72.191 2.77 ;
      RECT 72.27 2.575 72.275 2.84 ;
      RECT 72.965 1.806 73.135 2.14 ;
      RECT 72.935 1.806 73.135 2.135 ;
      RECT 72.875 1.773 72.935 2.123 ;
      RECT 72.875 1.829 73.145 2.118 ;
      RECT 72.85 1.829 73.145 2.112 ;
      RECT 72.845 1.77 72.875 2.109 ;
      RECT 72.83 1.776 72.965 2.107 ;
      RECT 72.825 1.784 73.05 2.095 ;
      RECT 72.825 1.836 73.16 2.048 ;
      RECT 72.81 1.792 73.05 2.043 ;
      RECT 72.81 1.862 73.17 1.984 ;
      RECT 72.78 1.812 73.135 1.945 ;
      RECT 72.78 1.902 73.18 1.941 ;
      RECT 72.83 1.781 73.05 2.107 ;
      RECT 72.17 2.111 72.225 2.375 ;
      RECT 72.17 2.111 72.29 2.374 ;
      RECT 72.17 2.111 72.315 2.373 ;
      RECT 72.17 2.111 72.38 2.372 ;
      RECT 72.315 2.077 72.395 2.371 ;
      RECT 72.13 2.121 72.54 2.37 ;
      RECT 72.17 2.118 72.54 2.37 ;
      RECT 72.13 2.126 72.545 2.363 ;
      RECT 72.115 2.128 72.545 2.362 ;
      RECT 72.115 2.135 72.55 2.358 ;
      RECT 72.095 2.134 72.545 2.354 ;
      RECT 72.095 2.142 72.555 2.353 ;
      RECT 72.09 2.139 72.55 2.349 ;
      RECT 72.09 2.152 72.565 2.348 ;
      RECT 72.075 2.142 72.555 2.347 ;
      RECT 72.04 2.155 72.565 2.34 ;
      RECT 72.225 2.11 72.535 2.37 ;
      RECT 72.225 2.095 72.485 2.37 ;
      RECT 72.29 2.082 72.42 2.37 ;
      RECT 71.835 3.171 71.85 3.564 ;
      RECT 71.8 3.176 71.85 3.563 ;
      RECT 71.835 3.175 71.895 3.562 ;
      RECT 71.78 3.186 71.895 3.561 ;
      RECT 71.795 3.182 71.895 3.561 ;
      RECT 71.76 3.192 71.97 3.558 ;
      RECT 71.76 3.211 72.015 3.556 ;
      RECT 71.76 3.218 72.02 3.553 ;
      RECT 71.745 3.195 71.97 3.55 ;
      RECT 71.725 3.2 71.97 3.543 ;
      RECT 71.72 3.204 71.97 3.539 ;
      RECT 71.72 3.221 72.03 3.538 ;
      RECT 71.7 3.215 72.015 3.534 ;
      RECT 71.7 3.224 72.035 3.528 ;
      RECT 71.695 3.23 72.035 3.3 ;
      RECT 71.76 3.19 71.895 3.558 ;
      RECT 71.635 2.553 71.835 2.865 ;
      RECT 71.71 2.531 71.835 2.865 ;
      RECT 71.65 2.55 71.84 2.85 ;
      RECT 71.62 2.561 71.84 2.848 ;
      RECT 71.635 2.556 71.845 2.814 ;
      RECT 71.62 2.66 71.85 2.781 ;
      RECT 71.65 2.532 71.835 2.865 ;
      RECT 71.71 2.51 71.81 2.865 ;
      RECT 71.735 2.507 71.81 2.865 ;
      RECT 71.735 2.502 71.755 2.865 ;
      RECT 71.14 2.57 71.315 2.745 ;
      RECT 71.135 2.57 71.315 2.743 ;
      RECT 71.11 2.57 71.315 2.738 ;
      RECT 71.055 2.55 71.225 2.728 ;
      RECT 71.055 2.557 71.29 2.728 ;
      RECT 71.14 3.237 71.155 3.42 ;
      RECT 71.13 3.215 71.14 3.42 ;
      RECT 71.115 3.195 71.13 3.42 ;
      RECT 71.105 3.17 71.115 3.42 ;
      RECT 71.075 3.135 71.105 3.42 ;
      RECT 71.04 3.075 71.075 3.42 ;
      RECT 71.035 3.037 71.04 3.42 ;
      RECT 70.985 2.988 71.035 3.42 ;
      RECT 70.975 2.938 70.985 3.408 ;
      RECT 70.96 2.917 70.975 3.368 ;
      RECT 70.94 2.885 70.96 3.318 ;
      RECT 70.915 2.841 70.94 3.258 ;
      RECT 70.91 2.813 70.915 3.213 ;
      RECT 70.905 2.804 70.91 3.199 ;
      RECT 70.9 2.797 70.905 3.186 ;
      RECT 70.895 2.792 70.9 3.175 ;
      RECT 70.89 2.777 70.895 3.165 ;
      RECT 70.885 2.755 70.89 3.152 ;
      RECT 70.875 2.715 70.885 3.127 ;
      RECT 70.85 2.645 70.875 3.083 ;
      RECT 70.845 2.585 70.85 3.048 ;
      RECT 70.83 2.565 70.845 3.015 ;
      RECT 70.825 2.565 70.83 2.99 ;
      RECT 70.795 2.565 70.825 2.945 ;
      RECT 70.75 2.565 70.795 2.885 ;
      RECT 70.675 2.565 70.75 2.833 ;
      RECT 70.67 2.565 70.675 2.798 ;
      RECT 70.665 2.565 70.67 2.788 ;
      RECT 70.66 2.565 70.665 2.768 ;
      RECT 70.925 1.785 71.095 2.255 ;
      RECT 70.87 1.778 71.065 2.239 ;
      RECT 70.87 1.792 71.1 2.238 ;
      RECT 70.855 1.793 71.1 2.219 ;
      RECT 70.85 1.811 71.1 2.205 ;
      RECT 70.855 1.794 71.105 2.203 ;
      RECT 70.84 1.825 71.105 2.188 ;
      RECT 70.855 1.8 71.11 2.173 ;
      RECT 70.835 1.84 71.11 2.17 ;
      RECT 70.85 1.812 71.115 2.155 ;
      RECT 70.85 1.824 71.12 2.135 ;
      RECT 70.835 1.84 71.125 2.118 ;
      RECT 70.835 1.85 71.13 1.973 ;
      RECT 70.83 1.85 71.13 1.93 ;
      RECT 70.83 1.865 71.135 1.908 ;
      RECT 70.925 1.775 71.065 2.255 ;
      RECT 70.925 1.773 71.035 2.255 ;
      RECT 71.011 1.77 71.035 2.255 ;
      RECT 70.67 3.437 70.675 3.483 ;
      RECT 70.66 3.285 70.67 3.507 ;
      RECT 70.655 3.13 70.66 3.532 ;
      RECT 70.64 3.092 70.655 3.543 ;
      RECT 70.635 3.075 70.64 3.55 ;
      RECT 70.625 3.063 70.635 3.557 ;
      RECT 70.62 3.054 70.625 3.559 ;
      RECT 70.615 3.052 70.62 3.563 ;
      RECT 70.57 3.043 70.615 3.578 ;
      RECT 70.565 3.035 70.57 3.592 ;
      RECT 70.56 3.032 70.565 3.596 ;
      RECT 70.545 3.027 70.56 3.604 ;
      RECT 70.49 3.017 70.545 3.615 ;
      RECT 70.455 3.005 70.49 3.616 ;
      RECT 70.446 3 70.455 3.61 ;
      RECT 70.36 3 70.446 3.6 ;
      RECT 70.33 3 70.36 3.578 ;
      RECT 70.32 3 70.325 3.558 ;
      RECT 70.315 3 70.32 3.52 ;
      RECT 70.31 3 70.315 3.478 ;
      RECT 70.305 3 70.31 3.438 ;
      RECT 70.3 3 70.305 3.368 ;
      RECT 70.29 3 70.3 3.29 ;
      RECT 70.285 3 70.29 3.19 ;
      RECT 70.325 3 70.33 3.56 ;
      RECT 69.82 3.082 69.91 3.56 ;
      RECT 69.805 3.085 69.925 3.558 ;
      RECT 69.82 3.084 69.925 3.558 ;
      RECT 69.785 3.091 69.95 3.548 ;
      RECT 69.805 3.085 69.95 3.548 ;
      RECT 69.77 3.097 69.95 3.536 ;
      RECT 69.805 3.088 70 3.529 ;
      RECT 69.756 3.105 70 3.527 ;
      RECT 69.785 3.095 70.01 3.515 ;
      RECT 69.756 3.116 70.04 3.506 ;
      RECT 69.67 3.14 70.04 3.5 ;
      RECT 69.67 3.153 70.08 3.483 ;
      RECT 69.665 3.175 70.08 3.476 ;
      RECT 69.635 3.19 70.08 3.466 ;
      RECT 69.63 3.201 70.08 3.456 ;
      RECT 69.6 3.214 70.08 3.447 ;
      RECT 69.585 3.232 70.08 3.436 ;
      RECT 69.56 3.245 70.08 3.426 ;
      RECT 69.82 3.081 69.83 3.56 ;
      RECT 69.866 2.505 69.905 2.75 ;
      RECT 69.78 2.505 69.915 2.748 ;
      RECT 69.665 2.53 69.915 2.745 ;
      RECT 69.665 2.53 69.92 2.743 ;
      RECT 69.665 2.53 69.935 2.738 ;
      RECT 69.771 2.505 69.95 2.718 ;
      RECT 69.685 2.513 69.95 2.718 ;
      RECT 69.355 1.865 69.525 2.3 ;
      RECT 69.345 1.899 69.525 2.283 ;
      RECT 69.425 1.835 69.595 2.27 ;
      RECT 69.33 1.91 69.595 2.248 ;
      RECT 69.425 1.845 69.6 2.238 ;
      RECT 69.355 1.897 69.63 2.223 ;
      RECT 69.315 1.923 69.63 2.208 ;
      RECT 69.315 1.965 69.64 2.188 ;
      RECT 69.31 1.99 69.645 2.17 ;
      RECT 69.31 2 69.65 2.155 ;
      RECT 69.305 1.937 69.63 2.153 ;
      RECT 69.305 2.01 69.655 2.138 ;
      RECT 69.3 1.947 69.63 2.135 ;
      RECT 69.295 2.031 69.66 2.118 ;
      RECT 69.295 2.063 69.665 2.098 ;
      RECT 69.29 1.977 69.64 2.09 ;
      RECT 69.295 1.962 69.63 2.118 ;
      RECT 69.31 1.932 69.63 2.17 ;
      RECT 69.155 2.519 69.38 2.775 ;
      RECT 69.155 2.552 69.4 2.765 ;
      RECT 69.12 2.552 69.4 2.763 ;
      RECT 69.12 2.565 69.405 2.753 ;
      RECT 69.12 2.585 69.415 2.745 ;
      RECT 69.12 2.682 69.42 2.738 ;
      RECT 69.1 2.43 69.23 2.728 ;
      RECT 69.055 2.585 69.415 2.67 ;
      RECT 69.045 2.43 69.23 2.615 ;
      RECT 69.045 2.462 69.316 2.615 ;
      RECT 69.01 2.992 69.03 3.17 ;
      RECT 68.975 2.945 69.01 3.17 ;
      RECT 68.96 2.885 68.975 3.17 ;
      RECT 68.935 2.832 68.96 3.17 ;
      RECT 68.92 2.785 68.935 3.17 ;
      RECT 68.9 2.762 68.92 3.17 ;
      RECT 68.875 2.727 68.9 3.17 ;
      RECT 68.865 2.573 68.875 3.17 ;
      RECT 68.835 2.568 68.865 3.161 ;
      RECT 68.83 2.565 68.835 3.151 ;
      RECT 68.815 2.565 68.83 3.125 ;
      RECT 68.81 2.565 68.815 3.088 ;
      RECT 68.785 2.565 68.81 3.04 ;
      RECT 68.765 2.565 68.785 2.965 ;
      RECT 68.755 2.565 68.765 2.925 ;
      RECT 68.75 2.565 68.755 2.9 ;
      RECT 68.745 2.565 68.75 2.883 ;
      RECT 68.74 2.565 68.745 2.865 ;
      RECT 68.735 2.566 68.74 2.855 ;
      RECT 68.725 2.568 68.735 2.823 ;
      RECT 68.715 2.57 68.725 2.79 ;
      RECT 68.705 2.573 68.715 2.763 ;
      RECT 69.03 3 69.255 3.17 ;
      RECT 68.36 1.812 68.53 2.265 ;
      RECT 68.36 1.812 68.62 2.231 ;
      RECT 68.36 1.812 68.65 2.215 ;
      RECT 68.36 1.812 68.68 2.188 ;
      RECT 68.616 1.79 68.695 2.17 ;
      RECT 68.395 1.797 68.7 2.155 ;
      RECT 68.395 1.805 68.71 2.118 ;
      RECT 68.355 1.832 68.71 2.09 ;
      RECT 68.34 1.845 68.71 2.055 ;
      RECT 68.36 1.82 68.73 2.045 ;
      RECT 68.335 1.885 68.73 2.015 ;
      RECT 68.335 1.915 68.735 1.998 ;
      RECT 68.33 1.945 68.735 1.985 ;
      RECT 68.395 1.794 68.695 2.17 ;
      RECT 68.53 1.791 68.616 2.249 ;
      RECT 68.481 1.792 68.695 2.17 ;
      RECT 68.625 3.452 68.67 3.645 ;
      RECT 68.615 3.422 68.625 3.645 ;
      RECT 68.61 3.407 68.615 3.645 ;
      RECT 68.57 3.317 68.61 3.645 ;
      RECT 68.565 3.23 68.57 3.645 ;
      RECT 68.555 3.2 68.565 3.645 ;
      RECT 68.55 3.16 68.555 3.645 ;
      RECT 68.54 3.122 68.55 3.645 ;
      RECT 68.535 3.087 68.54 3.645 ;
      RECT 68.515 3.04 68.535 3.645 ;
      RECT 68.5 2.965 68.515 3.645 ;
      RECT 68.495 2.92 68.5 3.64 ;
      RECT 68.49 2.9 68.495 3.613 ;
      RECT 68.485 2.88 68.49 3.598 ;
      RECT 68.48 2.855 68.485 3.578 ;
      RECT 68.475 2.833 68.48 3.563 ;
      RECT 68.47 2.811 68.475 3.545 ;
      RECT 68.465 2.79 68.47 3.535 ;
      RECT 68.455 2.762 68.465 3.505 ;
      RECT 68.445 2.725 68.455 3.473 ;
      RECT 68.435 2.685 68.445 3.44 ;
      RECT 68.425 2.663 68.435 3.41 ;
      RECT 68.395 2.615 68.425 3.342 ;
      RECT 68.38 2.575 68.395 3.269 ;
      RECT 68.37 2.575 68.38 3.235 ;
      RECT 68.365 2.575 68.37 3.21 ;
      RECT 68.36 2.575 68.365 3.195 ;
      RECT 68.355 2.575 68.36 3.173 ;
      RECT 68.35 2.575 68.355 3.16 ;
      RECT 68.335 2.575 68.35 3.125 ;
      RECT 68.315 2.575 68.335 3.065 ;
      RECT 68.305 2.575 68.315 3.015 ;
      RECT 68.285 2.575 68.305 2.963 ;
      RECT 68.265 2.575 68.285 2.92 ;
      RECT 68.255 2.575 68.265 2.908 ;
      RECT 68.225 2.575 68.255 2.895 ;
      RECT 68.195 2.596 68.225 2.875 ;
      RECT 68.185 2.624 68.195 2.855 ;
      RECT 68.17 2.641 68.185 2.823 ;
      RECT 68.165 2.655 68.17 2.79 ;
      RECT 68.16 2.663 68.165 2.763 ;
      RECT 68.155 2.671 68.16 2.725 ;
      RECT 68.16 3.195 68.165 3.53 ;
      RECT 68.125 3.182 68.16 3.529 ;
      RECT 68.055 3.122 68.125 3.528 ;
      RECT 67.975 3.065 68.055 3.527 ;
      RECT 67.84 3.025 67.975 3.526 ;
      RECT 67.84 3.212 68.175 3.515 ;
      RECT 67.8 3.212 68.175 3.505 ;
      RECT 67.8 3.23 68.18 3.5 ;
      RECT 67.8 3.32 68.185 3.49 ;
      RECT 67.795 3.015 67.96 3.47 ;
      RECT 67.79 3.015 67.96 3.213 ;
      RECT 67.79 3.172 68.155 3.213 ;
      RECT 67.79 3.16 68.15 3.213 ;
      RECT 66.92 5.02 67.09 6.49 ;
      RECT 66.92 6.315 67.095 6.485 ;
      RECT 66.55 1.74 66.72 2.93 ;
      RECT 66.55 1.74 67.02 1.91 ;
      RECT 66.55 6.97 67.02 7.14 ;
      RECT 66.55 5.95 66.72 7.14 ;
      RECT 65.56 1.74 65.73 2.93 ;
      RECT 65.56 1.74 66.03 1.91 ;
      RECT 65.56 6.97 66.03 7.14 ;
      RECT 65.56 5.95 65.73 7.14 ;
      RECT 63.71 2.635 63.88 3.865 ;
      RECT 63.765 0.855 63.935 2.805 ;
      RECT 63.71 0.575 63.88 1.025 ;
      RECT 63.71 7.855 63.88 8.305 ;
      RECT 63.765 6.075 63.935 8.025 ;
      RECT 63.71 5.015 63.88 6.245 ;
      RECT 63.19 0.575 63.36 3.865 ;
      RECT 63.19 2.075 63.595 2.405 ;
      RECT 63.19 1.235 63.595 1.565 ;
      RECT 63.19 5.015 63.36 8.305 ;
      RECT 63.19 7.315 63.595 7.645 ;
      RECT 63.19 6.475 63.595 6.805 ;
      RECT 60.525 1.975 61.255 2.215 ;
      RECT 61.067 1.77 61.255 2.215 ;
      RECT 60.895 1.782 61.27 2.209 ;
      RECT 60.81 1.797 61.29 2.194 ;
      RECT 60.81 1.812 61.295 2.184 ;
      RECT 60.765 1.832 61.31 2.176 ;
      RECT 60.742 1.867 61.325 2.13 ;
      RECT 60.656 1.89 61.33 2.09 ;
      RECT 60.656 1.908 61.34 2.06 ;
      RECT 60.525 1.977 61.345 2.023 ;
      RECT 60.57 1.92 61.34 2.06 ;
      RECT 60.656 1.872 61.325 2.13 ;
      RECT 60.742 1.841 61.31 2.176 ;
      RECT 60.765 1.822 61.295 2.184 ;
      RECT 60.81 1.795 61.27 2.209 ;
      RECT 60.895 1.777 61.255 2.215 ;
      RECT 60.981 1.771 61.255 2.215 ;
      RECT 61.067 1.766 61.2 2.215 ;
      RECT 61.153 1.761 61.2 2.215 ;
      RECT 60.845 2.659 61.015 3.045 ;
      RECT 60.84 2.659 61.015 3.04 ;
      RECT 60.815 2.659 61.015 3.005 ;
      RECT 60.815 2.687 61.025 2.995 ;
      RECT 60.795 2.687 61.025 2.955 ;
      RECT 60.79 2.687 61.025 2.928 ;
      RECT 60.79 2.705 61.03 2.92 ;
      RECT 60.735 2.705 61.03 2.855 ;
      RECT 60.735 2.722 61.04 2.838 ;
      RECT 60.725 2.722 61.04 2.778 ;
      RECT 60.725 2.739 61.045 2.775 ;
      RECT 60.72 2.575 60.89 2.753 ;
      RECT 60.72 2.609 60.976 2.753 ;
      RECT 60.715 3.375 60.72 3.388 ;
      RECT 60.71 3.27 60.715 3.393 ;
      RECT 60.685 3.13 60.71 3.408 ;
      RECT 60.65 3.081 60.685 3.44 ;
      RECT 60.645 3.049 60.65 3.46 ;
      RECT 60.64 3.04 60.645 3.46 ;
      RECT 60.56 3.005 60.64 3.46 ;
      RECT 60.497 2.975 60.56 3.46 ;
      RECT 60.411 2.963 60.497 3.46 ;
      RECT 60.325 2.949 60.411 3.46 ;
      RECT 60.245 2.936 60.325 3.446 ;
      RECT 60.21 2.928 60.245 3.426 ;
      RECT 60.2 2.925 60.21 3.417 ;
      RECT 60.17 2.92 60.2 3.404 ;
      RECT 60.12 2.895 60.17 3.38 ;
      RECT 60.106 2.869 60.12 3.362 ;
      RECT 60.02 2.829 60.106 3.338 ;
      RECT 59.975 2.777 60.02 3.307 ;
      RECT 59.965 2.752 59.975 3.294 ;
      RECT 59.96 2.533 59.965 2.555 ;
      RECT 59.955 2.735 59.965 3.29 ;
      RECT 59.955 2.531 59.96 2.645 ;
      RECT 59.945 2.527 59.955 3.286 ;
      RECT 59.901 2.525 59.945 3.274 ;
      RECT 59.815 2.525 59.901 3.245 ;
      RECT 59.785 2.525 59.815 3.218 ;
      RECT 59.77 2.525 59.785 3.206 ;
      RECT 59.73 2.537 59.77 3.191 ;
      RECT 59.71 2.556 59.73 3.17 ;
      RECT 59.7 2.566 59.71 3.154 ;
      RECT 59.69 2.572 59.7 3.143 ;
      RECT 59.67 2.582 59.69 3.126 ;
      RECT 59.665 2.591 59.67 3.113 ;
      RECT 59.66 2.595 59.665 3.063 ;
      RECT 59.65 2.601 59.66 2.98 ;
      RECT 59.645 2.605 59.65 2.894 ;
      RECT 59.64 2.625 59.645 2.831 ;
      RECT 59.635 2.648 59.64 2.778 ;
      RECT 59.63 2.666 59.635 2.723 ;
      RECT 60.24 2.485 60.41 2.745 ;
      RECT 60.41 2.45 60.455 2.731 ;
      RECT 60.371 2.452 60.46 2.714 ;
      RECT 60.26 2.469 60.546 2.685 ;
      RECT 60.26 2.484 60.55 2.657 ;
      RECT 60.26 2.465 60.46 2.714 ;
      RECT 60.285 2.453 60.41 2.745 ;
      RECT 60.371 2.451 60.455 2.731 ;
      RECT 59.425 1.84 59.595 2.33 ;
      RECT 59.425 1.84 59.63 2.31 ;
      RECT 59.56 1.76 59.67 2.27 ;
      RECT 59.541 1.764 59.69 2.24 ;
      RECT 59.455 1.772 59.71 2.223 ;
      RECT 59.455 1.778 59.715 2.213 ;
      RECT 59.455 1.787 59.735 2.201 ;
      RECT 59.43 1.812 59.765 2.179 ;
      RECT 59.43 1.832 59.77 2.159 ;
      RECT 59.425 1.845 59.78 2.139 ;
      RECT 59.425 1.912 59.785 2.12 ;
      RECT 59.425 2.045 59.79 2.107 ;
      RECT 59.42 1.85 59.78 1.94 ;
      RECT 59.43 1.807 59.735 2.201 ;
      RECT 59.541 1.762 59.67 2.27 ;
      RECT 59.415 3.515 59.715 3.77 ;
      RECT 59.5 3.481 59.715 3.77 ;
      RECT 59.5 3.484 59.72 3.63 ;
      RECT 59.435 3.505 59.72 3.63 ;
      RECT 59.47 3.495 59.715 3.77 ;
      RECT 59.465 3.5 59.72 3.63 ;
      RECT 59.5 3.479 59.701 3.77 ;
      RECT 59.586 3.47 59.701 3.77 ;
      RECT 59.586 3.464 59.615 3.77 ;
      RECT 59.075 3.105 59.085 3.595 ;
      RECT 58.735 3.04 58.745 3.34 ;
      RECT 59.25 3.212 59.255 3.431 ;
      RECT 59.24 3.192 59.25 3.448 ;
      RECT 59.23 3.172 59.24 3.478 ;
      RECT 59.225 3.162 59.23 3.493 ;
      RECT 59.22 3.158 59.225 3.498 ;
      RECT 59.205 3.15 59.22 3.505 ;
      RECT 59.165 3.13 59.205 3.53 ;
      RECT 59.14 3.112 59.165 3.563 ;
      RECT 59.135 3.11 59.14 3.576 ;
      RECT 59.115 3.107 59.135 3.58 ;
      RECT 59.085 3.105 59.115 3.59 ;
      RECT 59.015 3.107 59.075 3.591 ;
      RECT 58.995 3.107 59.015 3.585 ;
      RECT 58.97 3.105 58.995 3.582 ;
      RECT 58.935 3.1 58.97 3.578 ;
      RECT 58.915 3.094 58.935 3.565 ;
      RECT 58.905 3.091 58.915 3.553 ;
      RECT 58.885 3.088 58.905 3.538 ;
      RECT 58.865 3.084 58.885 3.52 ;
      RECT 58.86 3.081 58.865 3.51 ;
      RECT 58.855 3.08 58.86 3.508 ;
      RECT 58.845 3.077 58.855 3.5 ;
      RECT 58.835 3.071 58.845 3.483 ;
      RECT 58.825 3.065 58.835 3.465 ;
      RECT 58.815 3.059 58.825 3.453 ;
      RECT 58.805 3.053 58.815 3.433 ;
      RECT 58.8 3.049 58.805 3.418 ;
      RECT 58.795 3.047 58.8 3.41 ;
      RECT 58.79 3.045 58.795 3.403 ;
      RECT 58.785 3.043 58.79 3.393 ;
      RECT 58.78 3.041 58.785 3.387 ;
      RECT 58.77 3.04 58.78 3.377 ;
      RECT 58.76 3.04 58.77 3.368 ;
      RECT 58.745 3.04 58.76 3.353 ;
      RECT 58.705 3.04 58.735 3.337 ;
      RECT 58.685 3.042 58.705 3.332 ;
      RECT 58.68 3.047 58.685 3.33 ;
      RECT 58.65 3.055 58.68 3.328 ;
      RECT 58.62 3.07 58.65 3.327 ;
      RECT 58.575 3.092 58.62 3.332 ;
      RECT 58.57 3.107 58.575 3.336 ;
      RECT 58.555 3.112 58.57 3.338 ;
      RECT 58.55 3.116 58.555 3.34 ;
      RECT 58.49 3.139 58.55 3.349 ;
      RECT 58.47 3.165 58.49 3.362 ;
      RECT 58.46 3.172 58.47 3.366 ;
      RECT 58.445 3.179 58.46 3.369 ;
      RECT 58.425 3.189 58.445 3.372 ;
      RECT 58.42 3.197 58.425 3.375 ;
      RECT 58.375 3.202 58.42 3.382 ;
      RECT 58.365 3.205 58.375 3.389 ;
      RECT 58.355 3.205 58.365 3.393 ;
      RECT 58.32 3.207 58.355 3.405 ;
      RECT 58.3 3.21 58.32 3.418 ;
      RECT 58.26 3.213 58.3 3.429 ;
      RECT 58.245 3.215 58.26 3.442 ;
      RECT 58.235 3.215 58.245 3.447 ;
      RECT 58.21 3.216 58.235 3.455 ;
      RECT 58.2 3.218 58.21 3.46 ;
      RECT 58.195 3.219 58.2 3.463 ;
      RECT 58.17 3.217 58.195 3.466 ;
      RECT 58.155 3.215 58.17 3.467 ;
      RECT 58.135 3.212 58.155 3.469 ;
      RECT 58.115 3.207 58.135 3.469 ;
      RECT 58.055 3.202 58.115 3.466 ;
      RECT 58.02 3.177 58.055 3.462 ;
      RECT 58.01 3.154 58.02 3.46 ;
      RECT 57.98 3.131 58.01 3.46 ;
      RECT 57.97 3.11 57.98 3.46 ;
      RECT 57.945 3.092 57.97 3.458 ;
      RECT 57.93 3.07 57.945 3.455 ;
      RECT 57.915 3.052 57.93 3.453 ;
      RECT 57.895 3.042 57.915 3.451 ;
      RECT 57.88 3.037 57.895 3.45 ;
      RECT 57.865 3.035 57.88 3.449 ;
      RECT 57.835 3.036 57.865 3.447 ;
      RECT 57.815 3.039 57.835 3.445 ;
      RECT 57.758 3.043 57.815 3.445 ;
      RECT 57.672 3.052 57.758 3.445 ;
      RECT 57.586 3.063 57.672 3.445 ;
      RECT 57.5 3.074 57.586 3.445 ;
      RECT 57.48 3.081 57.5 3.453 ;
      RECT 57.47 3.084 57.48 3.46 ;
      RECT 57.405 3.089 57.47 3.478 ;
      RECT 57.375 3.096 57.405 3.503 ;
      RECT 57.365 3.099 57.375 3.51 ;
      RECT 57.32 3.103 57.365 3.515 ;
      RECT 57.29 3.108 57.32 3.52 ;
      RECT 57.289 3.11 57.29 3.52 ;
      RECT 57.203 3.116 57.289 3.52 ;
      RECT 57.117 3.127 57.203 3.52 ;
      RECT 57.031 3.139 57.117 3.52 ;
      RECT 56.945 3.15 57.031 3.52 ;
      RECT 56.93 3.157 56.945 3.515 ;
      RECT 56.925 3.159 56.93 3.509 ;
      RECT 56.905 3.17 56.925 3.504 ;
      RECT 56.895 3.188 56.905 3.498 ;
      RECT 56.89 3.2 56.895 3.298 ;
      RECT 59.185 1.953 59.205 2.04 ;
      RECT 59.18 1.888 59.185 2.072 ;
      RECT 59.17 1.855 59.18 2.077 ;
      RECT 59.165 1.835 59.17 2.083 ;
      RECT 59.135 1.835 59.165 2.1 ;
      RECT 59.086 1.835 59.135 2.136 ;
      RECT 59 1.835 59.086 2.194 ;
      RECT 58.971 1.845 59 2.243 ;
      RECT 58.885 1.887 58.971 2.296 ;
      RECT 58.865 1.925 58.885 2.343 ;
      RECT 58.84 1.942 58.865 2.363 ;
      RECT 58.83 1.956 58.84 2.383 ;
      RECT 58.825 1.962 58.83 2.393 ;
      RECT 58.82 1.966 58.825 2.4 ;
      RECT 58.77 1.986 58.82 2.405 ;
      RECT 58.705 2.03 58.77 2.405 ;
      RECT 58.68 2.08 58.705 2.405 ;
      RECT 58.67 2.11 58.68 2.405 ;
      RECT 58.665 2.137 58.67 2.405 ;
      RECT 58.66 2.155 58.665 2.405 ;
      RECT 58.65 2.197 58.66 2.405 ;
      RECT 59 2.755 59.17 2.93 ;
      RECT 58.94 2.583 59 2.918 ;
      RECT 58.93 2.576 58.94 2.901 ;
      RECT 58.885 2.755 59.17 2.881 ;
      RECT 58.866 2.755 59.17 2.859 ;
      RECT 58.78 2.755 59.17 2.824 ;
      RECT 58.76 2.575 58.93 2.78 ;
      RECT 58.76 2.722 59.165 2.78 ;
      RECT 58.76 2.67 59.14 2.78 ;
      RECT 58.76 2.625 59.105 2.78 ;
      RECT 58.76 2.607 59.07 2.78 ;
      RECT 58.76 2.597 59.065 2.78 ;
      RECT 58.93 7.855 59.1 8.305 ;
      RECT 58.985 6.075 59.155 8.025 ;
      RECT 58.93 5.015 59.1 6.245 ;
      RECT 58.41 5.015 58.58 8.305 ;
      RECT 58.41 7.315 58.815 7.645 ;
      RECT 58.41 6.475 58.815 6.805 ;
      RECT 58.48 3.555 58.67 3.78 ;
      RECT 58.47 3.556 58.675 3.775 ;
      RECT 58.47 3.558 58.685 3.755 ;
      RECT 58.47 3.562 58.69 3.74 ;
      RECT 58.47 3.549 58.64 3.775 ;
      RECT 58.47 3.552 58.665 3.775 ;
      RECT 58.48 3.548 58.64 3.78 ;
      RECT 58.566 3.546 58.64 3.78 ;
      RECT 58.19 2.797 58.36 3.035 ;
      RECT 58.19 2.797 58.446 2.949 ;
      RECT 58.19 2.797 58.45 2.859 ;
      RECT 58.24 2.57 58.46 2.838 ;
      RECT 58.235 2.587 58.465 2.811 ;
      RECT 58.2 2.745 58.465 2.811 ;
      RECT 58.22 2.595 58.36 3.035 ;
      RECT 58.21 2.677 58.47 2.794 ;
      RECT 58.205 2.725 58.47 2.794 ;
      RECT 58.21 2.635 58.465 2.811 ;
      RECT 58.235 2.572 58.46 2.838 ;
      RECT 57.8 2.547 57.97 2.745 ;
      RECT 57.8 2.547 58.015 2.72 ;
      RECT 57.87 2.49 58.04 2.678 ;
      RECT 57.845 2.505 58.04 2.678 ;
      RECT 57.46 2.551 57.49 2.745 ;
      RECT 57.455 2.523 57.46 2.745 ;
      RECT 57.425 2.497 57.455 2.747 ;
      RECT 57.4 2.455 57.425 2.75 ;
      RECT 57.39 2.427 57.4 2.752 ;
      RECT 57.355 2.407 57.39 2.754 ;
      RECT 57.29 2.392 57.355 2.76 ;
      RECT 57.24 2.39 57.29 2.766 ;
      RECT 57.217 2.392 57.24 2.771 ;
      RECT 57.131 2.403 57.217 2.777 ;
      RECT 57.045 2.421 57.131 2.787 ;
      RECT 57.03 2.432 57.045 2.793 ;
      RECT 56.96 2.455 57.03 2.799 ;
      RECT 56.905 2.487 56.96 2.807 ;
      RECT 56.865 2.51 56.905 2.813 ;
      RECT 56.851 2.523 56.865 2.816 ;
      RECT 56.765 2.545 56.851 2.822 ;
      RECT 56.75 2.57 56.765 2.828 ;
      RECT 56.71 2.585 56.75 2.832 ;
      RECT 56.66 2.6 56.71 2.837 ;
      RECT 56.635 2.607 56.66 2.841 ;
      RECT 56.575 2.602 56.635 2.845 ;
      RECT 56.56 2.593 56.575 2.849 ;
      RECT 56.49 2.583 56.56 2.845 ;
      RECT 56.465 2.575 56.485 2.835 ;
      RECT 56.406 2.575 56.465 2.813 ;
      RECT 56.32 2.575 56.406 2.77 ;
      RECT 56.485 2.575 56.49 2.84 ;
      RECT 57.18 1.806 57.35 2.14 ;
      RECT 57.15 1.806 57.35 2.135 ;
      RECT 57.09 1.773 57.15 2.123 ;
      RECT 57.09 1.829 57.36 2.118 ;
      RECT 57.065 1.829 57.36 2.112 ;
      RECT 57.06 1.77 57.09 2.109 ;
      RECT 57.045 1.776 57.18 2.107 ;
      RECT 57.04 1.784 57.265 2.095 ;
      RECT 57.04 1.836 57.375 2.048 ;
      RECT 57.025 1.792 57.265 2.043 ;
      RECT 57.025 1.862 57.385 1.984 ;
      RECT 56.995 1.812 57.35 1.945 ;
      RECT 56.995 1.902 57.395 1.941 ;
      RECT 57.045 1.781 57.265 2.107 ;
      RECT 56.385 2.111 56.44 2.375 ;
      RECT 56.385 2.111 56.505 2.374 ;
      RECT 56.385 2.111 56.53 2.373 ;
      RECT 56.385 2.111 56.595 2.372 ;
      RECT 56.53 2.077 56.61 2.371 ;
      RECT 56.345 2.121 56.755 2.37 ;
      RECT 56.385 2.118 56.755 2.37 ;
      RECT 56.345 2.126 56.76 2.363 ;
      RECT 56.33 2.128 56.76 2.362 ;
      RECT 56.33 2.135 56.765 2.358 ;
      RECT 56.31 2.134 56.76 2.354 ;
      RECT 56.31 2.142 56.77 2.353 ;
      RECT 56.305 2.139 56.765 2.349 ;
      RECT 56.305 2.152 56.78 2.348 ;
      RECT 56.29 2.142 56.77 2.347 ;
      RECT 56.255 2.155 56.78 2.34 ;
      RECT 56.44 2.11 56.75 2.37 ;
      RECT 56.44 2.095 56.7 2.37 ;
      RECT 56.505 2.082 56.635 2.37 ;
      RECT 56.05 3.171 56.065 3.564 ;
      RECT 56.015 3.176 56.065 3.563 ;
      RECT 56.05 3.175 56.11 3.562 ;
      RECT 55.995 3.186 56.11 3.561 ;
      RECT 56.01 3.182 56.11 3.561 ;
      RECT 55.975 3.192 56.185 3.558 ;
      RECT 55.975 3.211 56.23 3.556 ;
      RECT 55.975 3.218 56.235 3.553 ;
      RECT 55.96 3.195 56.185 3.55 ;
      RECT 55.94 3.2 56.185 3.543 ;
      RECT 55.935 3.204 56.185 3.539 ;
      RECT 55.935 3.221 56.245 3.538 ;
      RECT 55.915 3.215 56.23 3.534 ;
      RECT 55.915 3.224 56.25 3.528 ;
      RECT 55.91 3.23 56.25 3.3 ;
      RECT 55.975 3.19 56.11 3.558 ;
      RECT 55.85 2.553 56.05 2.865 ;
      RECT 55.925 2.531 56.05 2.865 ;
      RECT 55.865 2.55 56.055 2.85 ;
      RECT 55.835 2.561 56.055 2.848 ;
      RECT 55.85 2.556 56.06 2.814 ;
      RECT 55.835 2.66 56.065 2.781 ;
      RECT 55.865 2.532 56.05 2.865 ;
      RECT 55.925 2.51 56.025 2.865 ;
      RECT 55.95 2.507 56.025 2.865 ;
      RECT 55.95 2.502 55.97 2.865 ;
      RECT 55.355 2.57 55.53 2.745 ;
      RECT 55.35 2.57 55.53 2.743 ;
      RECT 55.325 2.57 55.53 2.738 ;
      RECT 55.27 2.55 55.44 2.728 ;
      RECT 55.27 2.557 55.505 2.728 ;
      RECT 55.355 3.237 55.37 3.42 ;
      RECT 55.345 3.215 55.355 3.42 ;
      RECT 55.33 3.195 55.345 3.42 ;
      RECT 55.32 3.17 55.33 3.42 ;
      RECT 55.29 3.135 55.32 3.42 ;
      RECT 55.255 3.075 55.29 3.42 ;
      RECT 55.25 3.037 55.255 3.42 ;
      RECT 55.2 2.988 55.25 3.42 ;
      RECT 55.19 2.938 55.2 3.408 ;
      RECT 55.175 2.917 55.19 3.368 ;
      RECT 55.155 2.885 55.175 3.318 ;
      RECT 55.13 2.841 55.155 3.258 ;
      RECT 55.125 2.813 55.13 3.213 ;
      RECT 55.12 2.804 55.125 3.199 ;
      RECT 55.115 2.797 55.12 3.186 ;
      RECT 55.11 2.792 55.115 3.175 ;
      RECT 55.105 2.777 55.11 3.165 ;
      RECT 55.1 2.755 55.105 3.152 ;
      RECT 55.09 2.715 55.1 3.127 ;
      RECT 55.065 2.645 55.09 3.083 ;
      RECT 55.06 2.585 55.065 3.048 ;
      RECT 55.045 2.565 55.06 3.015 ;
      RECT 55.04 2.565 55.045 2.99 ;
      RECT 55.01 2.565 55.04 2.945 ;
      RECT 54.965 2.565 55.01 2.885 ;
      RECT 54.89 2.565 54.965 2.833 ;
      RECT 54.885 2.565 54.89 2.798 ;
      RECT 54.88 2.565 54.885 2.788 ;
      RECT 54.875 2.565 54.88 2.768 ;
      RECT 55.14 1.785 55.31 2.255 ;
      RECT 55.085 1.778 55.28 2.239 ;
      RECT 55.085 1.792 55.315 2.238 ;
      RECT 55.07 1.793 55.315 2.219 ;
      RECT 55.065 1.811 55.315 2.205 ;
      RECT 55.07 1.794 55.32 2.203 ;
      RECT 55.055 1.825 55.32 2.188 ;
      RECT 55.07 1.8 55.325 2.173 ;
      RECT 55.05 1.84 55.325 2.17 ;
      RECT 55.065 1.812 55.33 2.155 ;
      RECT 55.065 1.824 55.335 2.135 ;
      RECT 55.05 1.84 55.34 2.118 ;
      RECT 55.05 1.85 55.345 1.973 ;
      RECT 55.045 1.85 55.345 1.93 ;
      RECT 55.045 1.865 55.35 1.908 ;
      RECT 55.14 1.775 55.28 2.255 ;
      RECT 55.14 1.773 55.25 2.255 ;
      RECT 55.226 1.77 55.25 2.255 ;
      RECT 54.885 3.437 54.89 3.483 ;
      RECT 54.875 3.285 54.885 3.507 ;
      RECT 54.87 3.13 54.875 3.532 ;
      RECT 54.855 3.092 54.87 3.543 ;
      RECT 54.85 3.075 54.855 3.55 ;
      RECT 54.84 3.063 54.85 3.557 ;
      RECT 54.835 3.054 54.84 3.559 ;
      RECT 54.83 3.052 54.835 3.563 ;
      RECT 54.785 3.043 54.83 3.578 ;
      RECT 54.78 3.035 54.785 3.592 ;
      RECT 54.775 3.032 54.78 3.596 ;
      RECT 54.76 3.027 54.775 3.604 ;
      RECT 54.705 3.017 54.76 3.615 ;
      RECT 54.67 3.005 54.705 3.616 ;
      RECT 54.661 3 54.67 3.61 ;
      RECT 54.575 3 54.661 3.6 ;
      RECT 54.545 3 54.575 3.578 ;
      RECT 54.535 3 54.54 3.558 ;
      RECT 54.53 3 54.535 3.52 ;
      RECT 54.525 3 54.53 3.478 ;
      RECT 54.52 3 54.525 3.438 ;
      RECT 54.515 3 54.52 3.368 ;
      RECT 54.505 3 54.515 3.29 ;
      RECT 54.5 3 54.505 3.19 ;
      RECT 54.54 3 54.545 3.56 ;
      RECT 54.035 3.082 54.125 3.56 ;
      RECT 54.02 3.085 54.14 3.558 ;
      RECT 54.035 3.084 54.14 3.558 ;
      RECT 54 3.091 54.165 3.548 ;
      RECT 54.02 3.085 54.165 3.548 ;
      RECT 53.985 3.097 54.165 3.536 ;
      RECT 54.02 3.088 54.215 3.529 ;
      RECT 53.971 3.105 54.215 3.527 ;
      RECT 54 3.095 54.225 3.515 ;
      RECT 53.971 3.116 54.255 3.506 ;
      RECT 53.885 3.14 54.255 3.5 ;
      RECT 53.885 3.153 54.295 3.483 ;
      RECT 53.88 3.175 54.295 3.476 ;
      RECT 53.85 3.19 54.295 3.466 ;
      RECT 53.845 3.201 54.295 3.456 ;
      RECT 53.815 3.214 54.295 3.447 ;
      RECT 53.8 3.232 54.295 3.436 ;
      RECT 53.775 3.245 54.295 3.426 ;
      RECT 54.035 3.081 54.045 3.56 ;
      RECT 54.081 2.505 54.12 2.75 ;
      RECT 53.995 2.505 54.13 2.748 ;
      RECT 53.88 2.53 54.13 2.745 ;
      RECT 53.88 2.53 54.135 2.743 ;
      RECT 53.88 2.53 54.15 2.738 ;
      RECT 53.986 2.505 54.165 2.718 ;
      RECT 53.9 2.513 54.165 2.718 ;
      RECT 53.57 1.865 53.74 2.3 ;
      RECT 53.56 1.899 53.74 2.283 ;
      RECT 53.64 1.835 53.81 2.27 ;
      RECT 53.545 1.91 53.81 2.248 ;
      RECT 53.64 1.845 53.815 2.238 ;
      RECT 53.57 1.897 53.845 2.223 ;
      RECT 53.53 1.923 53.845 2.208 ;
      RECT 53.53 1.965 53.855 2.188 ;
      RECT 53.525 1.99 53.86 2.17 ;
      RECT 53.525 2 53.865 2.155 ;
      RECT 53.52 1.937 53.845 2.153 ;
      RECT 53.52 2.01 53.87 2.138 ;
      RECT 53.515 1.947 53.845 2.135 ;
      RECT 53.51 2.031 53.875 2.118 ;
      RECT 53.51 2.063 53.88 2.098 ;
      RECT 53.505 1.977 53.855 2.09 ;
      RECT 53.51 1.962 53.845 2.118 ;
      RECT 53.525 1.932 53.845 2.17 ;
      RECT 53.37 2.519 53.595 2.775 ;
      RECT 53.37 2.552 53.615 2.765 ;
      RECT 53.335 2.552 53.615 2.763 ;
      RECT 53.335 2.565 53.62 2.753 ;
      RECT 53.335 2.585 53.63 2.745 ;
      RECT 53.335 2.682 53.635 2.738 ;
      RECT 53.315 2.43 53.445 2.728 ;
      RECT 53.27 2.585 53.63 2.67 ;
      RECT 53.26 2.43 53.445 2.615 ;
      RECT 53.26 2.462 53.531 2.615 ;
      RECT 53.225 2.992 53.245 3.17 ;
      RECT 53.19 2.945 53.225 3.17 ;
      RECT 53.175 2.885 53.19 3.17 ;
      RECT 53.15 2.832 53.175 3.17 ;
      RECT 53.135 2.785 53.15 3.17 ;
      RECT 53.115 2.762 53.135 3.17 ;
      RECT 53.09 2.727 53.115 3.17 ;
      RECT 53.08 2.573 53.09 3.17 ;
      RECT 53.05 2.568 53.08 3.161 ;
      RECT 53.045 2.565 53.05 3.151 ;
      RECT 53.03 2.565 53.045 3.125 ;
      RECT 53.025 2.565 53.03 3.088 ;
      RECT 53 2.565 53.025 3.04 ;
      RECT 52.98 2.565 53 2.965 ;
      RECT 52.97 2.565 52.98 2.925 ;
      RECT 52.965 2.565 52.97 2.9 ;
      RECT 52.96 2.565 52.965 2.883 ;
      RECT 52.955 2.565 52.96 2.865 ;
      RECT 52.95 2.566 52.955 2.855 ;
      RECT 52.94 2.568 52.95 2.823 ;
      RECT 52.93 2.57 52.94 2.79 ;
      RECT 52.92 2.573 52.93 2.763 ;
      RECT 53.245 3 53.47 3.17 ;
      RECT 52.575 1.812 52.745 2.265 ;
      RECT 52.575 1.812 52.835 2.231 ;
      RECT 52.575 1.812 52.865 2.215 ;
      RECT 52.575 1.812 52.895 2.188 ;
      RECT 52.831 1.79 52.91 2.17 ;
      RECT 52.61 1.797 52.915 2.155 ;
      RECT 52.61 1.805 52.925 2.118 ;
      RECT 52.57 1.832 52.925 2.09 ;
      RECT 52.555 1.845 52.925 2.055 ;
      RECT 52.575 1.82 52.945 2.045 ;
      RECT 52.55 1.885 52.945 2.015 ;
      RECT 52.55 1.915 52.95 1.998 ;
      RECT 52.545 1.945 52.95 1.985 ;
      RECT 52.61 1.794 52.91 2.17 ;
      RECT 52.745 1.791 52.831 2.249 ;
      RECT 52.696 1.792 52.91 2.17 ;
      RECT 52.84 3.452 52.885 3.645 ;
      RECT 52.83 3.422 52.84 3.645 ;
      RECT 52.825 3.407 52.83 3.645 ;
      RECT 52.785 3.317 52.825 3.645 ;
      RECT 52.78 3.23 52.785 3.645 ;
      RECT 52.77 3.2 52.78 3.645 ;
      RECT 52.765 3.16 52.77 3.645 ;
      RECT 52.755 3.122 52.765 3.645 ;
      RECT 52.75 3.087 52.755 3.645 ;
      RECT 52.73 3.04 52.75 3.645 ;
      RECT 52.715 2.965 52.73 3.645 ;
      RECT 52.71 2.92 52.715 3.64 ;
      RECT 52.705 2.9 52.71 3.613 ;
      RECT 52.7 2.88 52.705 3.598 ;
      RECT 52.695 2.855 52.7 3.578 ;
      RECT 52.69 2.833 52.695 3.563 ;
      RECT 52.685 2.811 52.69 3.545 ;
      RECT 52.68 2.79 52.685 3.535 ;
      RECT 52.67 2.762 52.68 3.505 ;
      RECT 52.66 2.725 52.67 3.473 ;
      RECT 52.65 2.685 52.66 3.44 ;
      RECT 52.64 2.663 52.65 3.41 ;
      RECT 52.61 2.615 52.64 3.342 ;
      RECT 52.595 2.575 52.61 3.269 ;
      RECT 52.585 2.575 52.595 3.235 ;
      RECT 52.58 2.575 52.585 3.21 ;
      RECT 52.575 2.575 52.58 3.195 ;
      RECT 52.57 2.575 52.575 3.173 ;
      RECT 52.565 2.575 52.57 3.16 ;
      RECT 52.55 2.575 52.565 3.125 ;
      RECT 52.53 2.575 52.55 3.065 ;
      RECT 52.52 2.575 52.53 3.015 ;
      RECT 52.5 2.575 52.52 2.963 ;
      RECT 52.48 2.575 52.5 2.92 ;
      RECT 52.47 2.575 52.48 2.908 ;
      RECT 52.44 2.575 52.47 2.895 ;
      RECT 52.41 2.596 52.44 2.875 ;
      RECT 52.4 2.624 52.41 2.855 ;
      RECT 52.385 2.641 52.4 2.823 ;
      RECT 52.38 2.655 52.385 2.79 ;
      RECT 52.375 2.663 52.38 2.763 ;
      RECT 52.37 2.671 52.375 2.725 ;
      RECT 52.375 3.195 52.38 3.53 ;
      RECT 52.34 3.182 52.375 3.529 ;
      RECT 52.27 3.122 52.34 3.528 ;
      RECT 52.19 3.065 52.27 3.527 ;
      RECT 52.055 3.025 52.19 3.526 ;
      RECT 52.055 3.212 52.39 3.515 ;
      RECT 52.015 3.212 52.39 3.505 ;
      RECT 52.015 3.23 52.395 3.5 ;
      RECT 52.015 3.32 52.4 3.49 ;
      RECT 52.01 3.015 52.175 3.47 ;
      RECT 52.005 3.015 52.175 3.213 ;
      RECT 52.005 3.172 52.37 3.213 ;
      RECT 52.005 3.16 52.365 3.213 ;
      RECT 51.135 5.02 51.305 6.49 ;
      RECT 51.135 6.315 51.31 6.485 ;
      RECT 50.765 1.74 50.935 2.93 ;
      RECT 50.765 1.74 51.235 1.91 ;
      RECT 50.765 6.97 51.235 7.14 ;
      RECT 50.765 5.95 50.935 7.14 ;
      RECT 49.775 1.74 49.945 2.93 ;
      RECT 49.775 1.74 50.245 1.91 ;
      RECT 49.775 6.97 50.245 7.14 ;
      RECT 49.775 5.95 49.945 7.14 ;
      RECT 47.925 2.635 48.095 3.865 ;
      RECT 47.98 0.855 48.15 2.805 ;
      RECT 47.925 0.575 48.095 1.025 ;
      RECT 47.925 7.855 48.095 8.305 ;
      RECT 47.98 6.075 48.15 8.025 ;
      RECT 47.925 5.015 48.095 6.245 ;
      RECT 47.405 0.575 47.575 3.865 ;
      RECT 47.405 2.075 47.81 2.405 ;
      RECT 47.405 1.235 47.81 1.565 ;
      RECT 47.405 5.015 47.575 8.305 ;
      RECT 47.405 7.315 47.81 7.645 ;
      RECT 47.405 6.475 47.81 6.805 ;
      RECT 44.74 1.975 45.47 2.215 ;
      RECT 45.282 1.77 45.47 2.215 ;
      RECT 45.11 1.782 45.485 2.209 ;
      RECT 45.025 1.797 45.505 2.194 ;
      RECT 45.025 1.812 45.51 2.184 ;
      RECT 44.98 1.832 45.525 2.176 ;
      RECT 44.957 1.867 45.54 2.13 ;
      RECT 44.871 1.89 45.545 2.09 ;
      RECT 44.871 1.908 45.555 2.06 ;
      RECT 44.74 1.977 45.56 2.023 ;
      RECT 44.785 1.92 45.555 2.06 ;
      RECT 44.871 1.872 45.54 2.13 ;
      RECT 44.957 1.841 45.525 2.176 ;
      RECT 44.98 1.822 45.51 2.184 ;
      RECT 45.025 1.795 45.485 2.209 ;
      RECT 45.11 1.777 45.47 2.215 ;
      RECT 45.196 1.771 45.47 2.215 ;
      RECT 45.282 1.766 45.415 2.215 ;
      RECT 45.368 1.761 45.415 2.215 ;
      RECT 45.06 2.659 45.23 3.045 ;
      RECT 45.055 2.659 45.23 3.04 ;
      RECT 45.03 2.659 45.23 3.005 ;
      RECT 45.03 2.687 45.24 2.995 ;
      RECT 45.01 2.687 45.24 2.955 ;
      RECT 45.005 2.687 45.24 2.928 ;
      RECT 45.005 2.705 45.245 2.92 ;
      RECT 44.95 2.705 45.245 2.855 ;
      RECT 44.95 2.722 45.255 2.838 ;
      RECT 44.94 2.722 45.255 2.778 ;
      RECT 44.94 2.739 45.26 2.775 ;
      RECT 44.935 2.575 45.105 2.753 ;
      RECT 44.935 2.609 45.191 2.753 ;
      RECT 44.93 3.375 44.935 3.388 ;
      RECT 44.925 3.27 44.93 3.393 ;
      RECT 44.9 3.13 44.925 3.408 ;
      RECT 44.865 3.081 44.9 3.44 ;
      RECT 44.86 3.049 44.865 3.46 ;
      RECT 44.855 3.04 44.86 3.46 ;
      RECT 44.775 3.005 44.855 3.46 ;
      RECT 44.712 2.975 44.775 3.46 ;
      RECT 44.626 2.963 44.712 3.46 ;
      RECT 44.54 2.949 44.626 3.46 ;
      RECT 44.46 2.936 44.54 3.446 ;
      RECT 44.425 2.928 44.46 3.426 ;
      RECT 44.415 2.925 44.425 3.417 ;
      RECT 44.385 2.92 44.415 3.404 ;
      RECT 44.335 2.895 44.385 3.38 ;
      RECT 44.321 2.869 44.335 3.362 ;
      RECT 44.235 2.829 44.321 3.338 ;
      RECT 44.19 2.777 44.235 3.307 ;
      RECT 44.18 2.752 44.19 3.294 ;
      RECT 44.175 2.533 44.18 2.555 ;
      RECT 44.17 2.735 44.18 3.29 ;
      RECT 44.17 2.531 44.175 2.645 ;
      RECT 44.16 2.527 44.17 3.286 ;
      RECT 44.116 2.525 44.16 3.274 ;
      RECT 44.03 2.525 44.116 3.245 ;
      RECT 44 2.525 44.03 3.218 ;
      RECT 43.985 2.525 44 3.206 ;
      RECT 43.945 2.537 43.985 3.191 ;
      RECT 43.925 2.556 43.945 3.17 ;
      RECT 43.915 2.566 43.925 3.154 ;
      RECT 43.905 2.572 43.915 3.143 ;
      RECT 43.885 2.582 43.905 3.126 ;
      RECT 43.88 2.591 43.885 3.113 ;
      RECT 43.875 2.595 43.88 3.063 ;
      RECT 43.865 2.601 43.875 2.98 ;
      RECT 43.86 2.605 43.865 2.894 ;
      RECT 43.855 2.625 43.86 2.831 ;
      RECT 43.85 2.648 43.855 2.778 ;
      RECT 43.845 2.666 43.85 2.723 ;
      RECT 44.455 2.485 44.625 2.745 ;
      RECT 44.625 2.45 44.67 2.731 ;
      RECT 44.586 2.452 44.675 2.714 ;
      RECT 44.475 2.469 44.761 2.685 ;
      RECT 44.475 2.484 44.765 2.657 ;
      RECT 44.475 2.465 44.675 2.714 ;
      RECT 44.5 2.453 44.625 2.745 ;
      RECT 44.586 2.451 44.67 2.731 ;
      RECT 43.64 1.84 43.81 2.33 ;
      RECT 43.64 1.84 43.845 2.31 ;
      RECT 43.775 1.76 43.885 2.27 ;
      RECT 43.756 1.764 43.905 2.24 ;
      RECT 43.67 1.772 43.925 2.223 ;
      RECT 43.67 1.778 43.93 2.213 ;
      RECT 43.67 1.787 43.95 2.201 ;
      RECT 43.645 1.812 43.98 2.179 ;
      RECT 43.645 1.832 43.985 2.159 ;
      RECT 43.64 1.845 43.995 2.139 ;
      RECT 43.64 1.912 44 2.12 ;
      RECT 43.64 2.045 44.005 2.107 ;
      RECT 43.635 1.85 43.995 1.94 ;
      RECT 43.645 1.807 43.95 2.201 ;
      RECT 43.756 1.762 43.885 2.27 ;
      RECT 43.63 3.515 43.93 3.77 ;
      RECT 43.715 3.481 43.93 3.77 ;
      RECT 43.715 3.484 43.935 3.63 ;
      RECT 43.65 3.505 43.935 3.63 ;
      RECT 43.685 3.495 43.93 3.77 ;
      RECT 43.68 3.5 43.935 3.63 ;
      RECT 43.715 3.479 43.916 3.77 ;
      RECT 43.801 3.47 43.916 3.77 ;
      RECT 43.801 3.464 43.83 3.77 ;
      RECT 43.29 3.105 43.3 3.595 ;
      RECT 42.95 3.04 42.96 3.34 ;
      RECT 43.465 3.212 43.47 3.431 ;
      RECT 43.455 3.192 43.465 3.448 ;
      RECT 43.445 3.172 43.455 3.478 ;
      RECT 43.44 3.162 43.445 3.493 ;
      RECT 43.435 3.158 43.44 3.498 ;
      RECT 43.42 3.15 43.435 3.505 ;
      RECT 43.38 3.13 43.42 3.53 ;
      RECT 43.355 3.112 43.38 3.563 ;
      RECT 43.35 3.11 43.355 3.576 ;
      RECT 43.33 3.107 43.35 3.58 ;
      RECT 43.3 3.105 43.33 3.59 ;
      RECT 43.23 3.107 43.29 3.591 ;
      RECT 43.21 3.107 43.23 3.585 ;
      RECT 43.185 3.105 43.21 3.582 ;
      RECT 43.15 3.1 43.185 3.578 ;
      RECT 43.13 3.094 43.15 3.565 ;
      RECT 43.12 3.091 43.13 3.553 ;
      RECT 43.1 3.088 43.12 3.538 ;
      RECT 43.08 3.084 43.1 3.52 ;
      RECT 43.075 3.081 43.08 3.51 ;
      RECT 43.07 3.08 43.075 3.508 ;
      RECT 43.06 3.077 43.07 3.5 ;
      RECT 43.05 3.071 43.06 3.483 ;
      RECT 43.04 3.065 43.05 3.465 ;
      RECT 43.03 3.059 43.04 3.453 ;
      RECT 43.02 3.053 43.03 3.433 ;
      RECT 43.015 3.049 43.02 3.418 ;
      RECT 43.01 3.047 43.015 3.41 ;
      RECT 43.005 3.045 43.01 3.403 ;
      RECT 43 3.043 43.005 3.393 ;
      RECT 42.995 3.041 43 3.387 ;
      RECT 42.985 3.04 42.995 3.377 ;
      RECT 42.975 3.04 42.985 3.368 ;
      RECT 42.96 3.04 42.975 3.353 ;
      RECT 42.92 3.04 42.95 3.337 ;
      RECT 42.9 3.042 42.92 3.332 ;
      RECT 42.895 3.047 42.9 3.33 ;
      RECT 42.865 3.055 42.895 3.328 ;
      RECT 42.835 3.07 42.865 3.327 ;
      RECT 42.79 3.092 42.835 3.332 ;
      RECT 42.785 3.107 42.79 3.336 ;
      RECT 42.77 3.112 42.785 3.338 ;
      RECT 42.765 3.116 42.77 3.34 ;
      RECT 42.705 3.139 42.765 3.349 ;
      RECT 42.685 3.165 42.705 3.362 ;
      RECT 42.675 3.172 42.685 3.366 ;
      RECT 42.66 3.179 42.675 3.369 ;
      RECT 42.64 3.189 42.66 3.372 ;
      RECT 42.635 3.197 42.64 3.375 ;
      RECT 42.59 3.202 42.635 3.382 ;
      RECT 42.58 3.205 42.59 3.389 ;
      RECT 42.57 3.205 42.58 3.393 ;
      RECT 42.535 3.207 42.57 3.405 ;
      RECT 42.515 3.21 42.535 3.418 ;
      RECT 42.475 3.213 42.515 3.429 ;
      RECT 42.46 3.215 42.475 3.442 ;
      RECT 42.45 3.215 42.46 3.447 ;
      RECT 42.425 3.216 42.45 3.455 ;
      RECT 42.415 3.218 42.425 3.46 ;
      RECT 42.41 3.219 42.415 3.463 ;
      RECT 42.385 3.217 42.41 3.466 ;
      RECT 42.37 3.215 42.385 3.467 ;
      RECT 42.35 3.212 42.37 3.469 ;
      RECT 42.33 3.207 42.35 3.469 ;
      RECT 42.27 3.202 42.33 3.466 ;
      RECT 42.235 3.177 42.27 3.462 ;
      RECT 42.225 3.154 42.235 3.46 ;
      RECT 42.195 3.131 42.225 3.46 ;
      RECT 42.185 3.11 42.195 3.46 ;
      RECT 42.16 3.092 42.185 3.458 ;
      RECT 42.145 3.07 42.16 3.455 ;
      RECT 42.13 3.052 42.145 3.453 ;
      RECT 42.11 3.042 42.13 3.451 ;
      RECT 42.095 3.037 42.11 3.45 ;
      RECT 42.08 3.035 42.095 3.449 ;
      RECT 42.05 3.036 42.08 3.447 ;
      RECT 42.03 3.039 42.05 3.445 ;
      RECT 41.973 3.043 42.03 3.445 ;
      RECT 41.887 3.052 41.973 3.445 ;
      RECT 41.801 3.063 41.887 3.445 ;
      RECT 41.715 3.074 41.801 3.445 ;
      RECT 41.695 3.081 41.715 3.453 ;
      RECT 41.685 3.084 41.695 3.46 ;
      RECT 41.62 3.089 41.685 3.478 ;
      RECT 41.59 3.096 41.62 3.503 ;
      RECT 41.58 3.099 41.59 3.51 ;
      RECT 41.535 3.103 41.58 3.515 ;
      RECT 41.505 3.108 41.535 3.52 ;
      RECT 41.504 3.11 41.505 3.52 ;
      RECT 41.418 3.116 41.504 3.52 ;
      RECT 41.332 3.127 41.418 3.52 ;
      RECT 41.246 3.139 41.332 3.52 ;
      RECT 41.16 3.15 41.246 3.52 ;
      RECT 41.145 3.157 41.16 3.515 ;
      RECT 41.14 3.159 41.145 3.509 ;
      RECT 41.12 3.17 41.14 3.504 ;
      RECT 41.11 3.188 41.12 3.498 ;
      RECT 41.105 3.2 41.11 3.298 ;
      RECT 43.4 1.953 43.42 2.04 ;
      RECT 43.395 1.888 43.4 2.072 ;
      RECT 43.385 1.855 43.395 2.077 ;
      RECT 43.38 1.835 43.385 2.083 ;
      RECT 43.35 1.835 43.38 2.1 ;
      RECT 43.301 1.835 43.35 2.136 ;
      RECT 43.215 1.835 43.301 2.194 ;
      RECT 43.186 1.845 43.215 2.243 ;
      RECT 43.1 1.887 43.186 2.296 ;
      RECT 43.08 1.925 43.1 2.343 ;
      RECT 43.055 1.942 43.08 2.363 ;
      RECT 43.045 1.956 43.055 2.383 ;
      RECT 43.04 1.962 43.045 2.393 ;
      RECT 43.035 1.966 43.04 2.4 ;
      RECT 42.985 1.986 43.035 2.405 ;
      RECT 42.92 2.03 42.985 2.405 ;
      RECT 42.895 2.08 42.92 2.405 ;
      RECT 42.885 2.11 42.895 2.405 ;
      RECT 42.88 2.137 42.885 2.405 ;
      RECT 42.875 2.155 42.88 2.405 ;
      RECT 42.865 2.197 42.875 2.405 ;
      RECT 43.215 2.755 43.385 2.93 ;
      RECT 43.155 2.583 43.215 2.918 ;
      RECT 43.145 2.576 43.155 2.901 ;
      RECT 43.1 2.755 43.385 2.881 ;
      RECT 43.081 2.755 43.385 2.859 ;
      RECT 42.995 2.755 43.385 2.824 ;
      RECT 42.975 2.575 43.145 2.78 ;
      RECT 42.975 2.722 43.38 2.78 ;
      RECT 42.975 2.67 43.355 2.78 ;
      RECT 42.975 2.625 43.32 2.78 ;
      RECT 42.975 2.607 43.285 2.78 ;
      RECT 42.975 2.597 43.28 2.78 ;
      RECT 43.145 7.855 43.315 8.305 ;
      RECT 43.2 6.075 43.37 8.025 ;
      RECT 43.145 5.015 43.315 6.245 ;
      RECT 42.625 5.015 42.795 8.305 ;
      RECT 42.625 7.315 43.03 7.645 ;
      RECT 42.625 6.475 43.03 6.805 ;
      RECT 42.695 3.555 42.885 3.78 ;
      RECT 42.685 3.556 42.89 3.775 ;
      RECT 42.685 3.558 42.9 3.755 ;
      RECT 42.685 3.562 42.905 3.74 ;
      RECT 42.685 3.549 42.855 3.775 ;
      RECT 42.685 3.552 42.88 3.775 ;
      RECT 42.695 3.548 42.855 3.78 ;
      RECT 42.781 3.546 42.855 3.78 ;
      RECT 42.405 2.797 42.575 3.035 ;
      RECT 42.405 2.797 42.661 2.949 ;
      RECT 42.405 2.797 42.665 2.859 ;
      RECT 42.455 2.57 42.675 2.838 ;
      RECT 42.45 2.587 42.68 2.811 ;
      RECT 42.415 2.745 42.68 2.811 ;
      RECT 42.435 2.595 42.575 3.035 ;
      RECT 42.425 2.677 42.685 2.794 ;
      RECT 42.42 2.725 42.685 2.794 ;
      RECT 42.425 2.635 42.68 2.811 ;
      RECT 42.45 2.572 42.675 2.838 ;
      RECT 42.015 2.547 42.185 2.745 ;
      RECT 42.015 2.547 42.23 2.72 ;
      RECT 42.085 2.49 42.255 2.678 ;
      RECT 42.06 2.505 42.255 2.678 ;
      RECT 41.675 2.551 41.705 2.745 ;
      RECT 41.67 2.523 41.675 2.745 ;
      RECT 41.64 2.497 41.67 2.747 ;
      RECT 41.615 2.455 41.64 2.75 ;
      RECT 41.605 2.427 41.615 2.752 ;
      RECT 41.57 2.407 41.605 2.754 ;
      RECT 41.505 2.392 41.57 2.76 ;
      RECT 41.455 2.39 41.505 2.766 ;
      RECT 41.432 2.392 41.455 2.771 ;
      RECT 41.346 2.403 41.432 2.777 ;
      RECT 41.26 2.421 41.346 2.787 ;
      RECT 41.245 2.432 41.26 2.793 ;
      RECT 41.175 2.455 41.245 2.799 ;
      RECT 41.12 2.487 41.175 2.807 ;
      RECT 41.08 2.51 41.12 2.813 ;
      RECT 41.066 2.523 41.08 2.816 ;
      RECT 40.98 2.545 41.066 2.822 ;
      RECT 40.965 2.57 40.98 2.828 ;
      RECT 40.925 2.585 40.965 2.832 ;
      RECT 40.875 2.6 40.925 2.837 ;
      RECT 40.85 2.607 40.875 2.841 ;
      RECT 40.79 2.602 40.85 2.845 ;
      RECT 40.775 2.593 40.79 2.849 ;
      RECT 40.705 2.583 40.775 2.845 ;
      RECT 40.68 2.575 40.7 2.835 ;
      RECT 40.621 2.575 40.68 2.813 ;
      RECT 40.535 2.575 40.621 2.77 ;
      RECT 40.7 2.575 40.705 2.84 ;
      RECT 41.395 1.806 41.565 2.14 ;
      RECT 41.365 1.806 41.565 2.135 ;
      RECT 41.305 1.773 41.365 2.123 ;
      RECT 41.305 1.829 41.575 2.118 ;
      RECT 41.28 1.829 41.575 2.112 ;
      RECT 41.275 1.77 41.305 2.109 ;
      RECT 41.26 1.776 41.395 2.107 ;
      RECT 41.255 1.784 41.48 2.095 ;
      RECT 41.255 1.836 41.59 2.048 ;
      RECT 41.24 1.792 41.48 2.043 ;
      RECT 41.24 1.862 41.6 1.984 ;
      RECT 41.21 1.812 41.565 1.945 ;
      RECT 41.21 1.902 41.61 1.941 ;
      RECT 41.26 1.781 41.48 2.107 ;
      RECT 40.6 2.111 40.655 2.375 ;
      RECT 40.6 2.111 40.72 2.374 ;
      RECT 40.6 2.111 40.745 2.373 ;
      RECT 40.6 2.111 40.81 2.372 ;
      RECT 40.745 2.077 40.825 2.371 ;
      RECT 40.56 2.121 40.97 2.37 ;
      RECT 40.6 2.118 40.97 2.37 ;
      RECT 40.56 2.126 40.975 2.363 ;
      RECT 40.545 2.128 40.975 2.362 ;
      RECT 40.545 2.135 40.98 2.358 ;
      RECT 40.525 2.134 40.975 2.354 ;
      RECT 40.525 2.142 40.985 2.353 ;
      RECT 40.52 2.139 40.98 2.349 ;
      RECT 40.52 2.152 40.995 2.348 ;
      RECT 40.505 2.142 40.985 2.347 ;
      RECT 40.47 2.155 40.995 2.34 ;
      RECT 40.655 2.11 40.965 2.37 ;
      RECT 40.655 2.095 40.915 2.37 ;
      RECT 40.72 2.082 40.85 2.37 ;
      RECT 40.265 3.171 40.28 3.564 ;
      RECT 40.23 3.176 40.28 3.563 ;
      RECT 40.265 3.175 40.325 3.562 ;
      RECT 40.21 3.186 40.325 3.561 ;
      RECT 40.225 3.182 40.325 3.561 ;
      RECT 40.19 3.192 40.4 3.558 ;
      RECT 40.19 3.211 40.445 3.556 ;
      RECT 40.19 3.218 40.45 3.553 ;
      RECT 40.175 3.195 40.4 3.55 ;
      RECT 40.155 3.2 40.4 3.543 ;
      RECT 40.15 3.204 40.4 3.539 ;
      RECT 40.15 3.221 40.46 3.538 ;
      RECT 40.13 3.215 40.445 3.534 ;
      RECT 40.13 3.224 40.465 3.528 ;
      RECT 40.125 3.23 40.465 3.3 ;
      RECT 40.19 3.19 40.325 3.558 ;
      RECT 40.065 2.553 40.265 2.865 ;
      RECT 40.14 2.531 40.265 2.865 ;
      RECT 40.08 2.55 40.27 2.85 ;
      RECT 40.05 2.561 40.27 2.848 ;
      RECT 40.065 2.556 40.275 2.814 ;
      RECT 40.05 2.66 40.28 2.781 ;
      RECT 40.08 2.532 40.265 2.865 ;
      RECT 40.14 2.51 40.24 2.865 ;
      RECT 40.165 2.507 40.24 2.865 ;
      RECT 40.165 2.502 40.185 2.865 ;
      RECT 39.57 2.57 39.745 2.745 ;
      RECT 39.565 2.57 39.745 2.743 ;
      RECT 39.54 2.57 39.745 2.738 ;
      RECT 39.485 2.55 39.655 2.728 ;
      RECT 39.485 2.557 39.72 2.728 ;
      RECT 39.57 3.237 39.585 3.42 ;
      RECT 39.56 3.215 39.57 3.42 ;
      RECT 39.545 3.195 39.56 3.42 ;
      RECT 39.535 3.17 39.545 3.42 ;
      RECT 39.505 3.135 39.535 3.42 ;
      RECT 39.47 3.075 39.505 3.42 ;
      RECT 39.465 3.037 39.47 3.42 ;
      RECT 39.415 2.988 39.465 3.42 ;
      RECT 39.405 2.938 39.415 3.408 ;
      RECT 39.39 2.917 39.405 3.368 ;
      RECT 39.37 2.885 39.39 3.318 ;
      RECT 39.345 2.841 39.37 3.258 ;
      RECT 39.34 2.813 39.345 3.213 ;
      RECT 39.335 2.804 39.34 3.199 ;
      RECT 39.33 2.797 39.335 3.186 ;
      RECT 39.325 2.792 39.33 3.175 ;
      RECT 39.32 2.777 39.325 3.165 ;
      RECT 39.315 2.755 39.32 3.152 ;
      RECT 39.305 2.715 39.315 3.127 ;
      RECT 39.28 2.645 39.305 3.083 ;
      RECT 39.275 2.585 39.28 3.048 ;
      RECT 39.26 2.565 39.275 3.015 ;
      RECT 39.255 2.565 39.26 2.99 ;
      RECT 39.225 2.565 39.255 2.945 ;
      RECT 39.18 2.565 39.225 2.885 ;
      RECT 39.105 2.565 39.18 2.833 ;
      RECT 39.1 2.565 39.105 2.798 ;
      RECT 39.095 2.565 39.1 2.788 ;
      RECT 39.09 2.565 39.095 2.768 ;
      RECT 39.355 1.785 39.525 2.255 ;
      RECT 39.3 1.778 39.495 2.239 ;
      RECT 39.3 1.792 39.53 2.238 ;
      RECT 39.285 1.793 39.53 2.219 ;
      RECT 39.28 1.811 39.53 2.205 ;
      RECT 39.285 1.794 39.535 2.203 ;
      RECT 39.27 1.825 39.535 2.188 ;
      RECT 39.285 1.8 39.54 2.173 ;
      RECT 39.265 1.84 39.54 2.17 ;
      RECT 39.28 1.812 39.545 2.155 ;
      RECT 39.28 1.824 39.55 2.135 ;
      RECT 39.265 1.84 39.555 2.118 ;
      RECT 39.265 1.85 39.56 1.973 ;
      RECT 39.26 1.85 39.56 1.93 ;
      RECT 39.26 1.865 39.565 1.908 ;
      RECT 39.355 1.775 39.495 2.255 ;
      RECT 39.355 1.773 39.465 2.255 ;
      RECT 39.441 1.77 39.465 2.255 ;
      RECT 39.1 3.437 39.105 3.483 ;
      RECT 39.09 3.285 39.1 3.507 ;
      RECT 39.085 3.13 39.09 3.532 ;
      RECT 39.07 3.092 39.085 3.543 ;
      RECT 39.065 3.075 39.07 3.55 ;
      RECT 39.055 3.063 39.065 3.557 ;
      RECT 39.05 3.054 39.055 3.559 ;
      RECT 39.045 3.052 39.05 3.563 ;
      RECT 39 3.043 39.045 3.578 ;
      RECT 38.995 3.035 39 3.592 ;
      RECT 38.99 3.032 38.995 3.596 ;
      RECT 38.975 3.027 38.99 3.604 ;
      RECT 38.92 3.017 38.975 3.615 ;
      RECT 38.885 3.005 38.92 3.616 ;
      RECT 38.876 3 38.885 3.61 ;
      RECT 38.79 3 38.876 3.6 ;
      RECT 38.76 3 38.79 3.578 ;
      RECT 38.75 3 38.755 3.558 ;
      RECT 38.745 3 38.75 3.52 ;
      RECT 38.74 3 38.745 3.478 ;
      RECT 38.735 3 38.74 3.438 ;
      RECT 38.73 3 38.735 3.368 ;
      RECT 38.72 3 38.73 3.29 ;
      RECT 38.715 3 38.72 3.19 ;
      RECT 38.755 3 38.76 3.56 ;
      RECT 38.25 3.082 38.34 3.56 ;
      RECT 38.235 3.085 38.355 3.558 ;
      RECT 38.25 3.084 38.355 3.558 ;
      RECT 38.215 3.091 38.38 3.548 ;
      RECT 38.235 3.085 38.38 3.548 ;
      RECT 38.2 3.097 38.38 3.536 ;
      RECT 38.235 3.088 38.43 3.529 ;
      RECT 38.186 3.105 38.43 3.527 ;
      RECT 38.215 3.095 38.44 3.515 ;
      RECT 38.186 3.116 38.47 3.506 ;
      RECT 38.1 3.14 38.47 3.5 ;
      RECT 38.1 3.153 38.51 3.483 ;
      RECT 38.095 3.175 38.51 3.476 ;
      RECT 38.065 3.19 38.51 3.466 ;
      RECT 38.06 3.201 38.51 3.456 ;
      RECT 38.03 3.214 38.51 3.447 ;
      RECT 38.015 3.232 38.51 3.436 ;
      RECT 37.99 3.245 38.51 3.426 ;
      RECT 38.25 3.081 38.26 3.56 ;
      RECT 38.296 2.505 38.335 2.75 ;
      RECT 38.21 2.505 38.345 2.748 ;
      RECT 38.095 2.53 38.345 2.745 ;
      RECT 38.095 2.53 38.35 2.743 ;
      RECT 38.095 2.53 38.365 2.738 ;
      RECT 38.201 2.505 38.38 2.718 ;
      RECT 38.115 2.513 38.38 2.718 ;
      RECT 37.785 1.865 37.955 2.3 ;
      RECT 37.775 1.899 37.955 2.283 ;
      RECT 37.855 1.835 38.025 2.27 ;
      RECT 37.76 1.91 38.025 2.248 ;
      RECT 37.855 1.845 38.03 2.238 ;
      RECT 37.785 1.897 38.06 2.223 ;
      RECT 37.745 1.923 38.06 2.208 ;
      RECT 37.745 1.965 38.07 2.188 ;
      RECT 37.74 1.99 38.075 2.17 ;
      RECT 37.74 2 38.08 2.155 ;
      RECT 37.735 1.937 38.06 2.153 ;
      RECT 37.735 2.01 38.085 2.138 ;
      RECT 37.73 1.947 38.06 2.135 ;
      RECT 37.725 2.031 38.09 2.118 ;
      RECT 37.725 2.063 38.095 2.098 ;
      RECT 37.72 1.977 38.07 2.09 ;
      RECT 37.725 1.962 38.06 2.118 ;
      RECT 37.74 1.932 38.06 2.17 ;
      RECT 37.585 2.519 37.81 2.775 ;
      RECT 37.585 2.552 37.83 2.765 ;
      RECT 37.55 2.552 37.83 2.763 ;
      RECT 37.55 2.565 37.835 2.753 ;
      RECT 37.55 2.585 37.845 2.745 ;
      RECT 37.55 2.682 37.85 2.738 ;
      RECT 37.53 2.43 37.66 2.728 ;
      RECT 37.485 2.585 37.845 2.67 ;
      RECT 37.475 2.43 37.66 2.615 ;
      RECT 37.475 2.462 37.746 2.615 ;
      RECT 37.44 2.992 37.46 3.17 ;
      RECT 37.405 2.945 37.44 3.17 ;
      RECT 37.39 2.885 37.405 3.17 ;
      RECT 37.365 2.832 37.39 3.17 ;
      RECT 37.35 2.785 37.365 3.17 ;
      RECT 37.33 2.762 37.35 3.17 ;
      RECT 37.305 2.727 37.33 3.17 ;
      RECT 37.295 2.573 37.305 3.17 ;
      RECT 37.265 2.568 37.295 3.161 ;
      RECT 37.26 2.565 37.265 3.151 ;
      RECT 37.245 2.565 37.26 3.125 ;
      RECT 37.24 2.565 37.245 3.088 ;
      RECT 37.215 2.565 37.24 3.04 ;
      RECT 37.195 2.565 37.215 2.965 ;
      RECT 37.185 2.565 37.195 2.925 ;
      RECT 37.18 2.565 37.185 2.9 ;
      RECT 37.175 2.565 37.18 2.883 ;
      RECT 37.17 2.565 37.175 2.865 ;
      RECT 37.165 2.566 37.17 2.855 ;
      RECT 37.155 2.568 37.165 2.823 ;
      RECT 37.145 2.57 37.155 2.79 ;
      RECT 37.135 2.573 37.145 2.763 ;
      RECT 37.46 3 37.685 3.17 ;
      RECT 36.79 1.812 36.96 2.265 ;
      RECT 36.79 1.812 37.05 2.231 ;
      RECT 36.79 1.812 37.08 2.215 ;
      RECT 36.79 1.812 37.11 2.188 ;
      RECT 37.046 1.79 37.125 2.17 ;
      RECT 36.825 1.797 37.13 2.155 ;
      RECT 36.825 1.805 37.14 2.118 ;
      RECT 36.785 1.832 37.14 2.09 ;
      RECT 36.77 1.845 37.14 2.055 ;
      RECT 36.79 1.82 37.16 2.045 ;
      RECT 36.765 1.885 37.16 2.015 ;
      RECT 36.765 1.915 37.165 1.998 ;
      RECT 36.76 1.945 37.165 1.985 ;
      RECT 36.825 1.794 37.125 2.17 ;
      RECT 36.96 1.791 37.046 2.249 ;
      RECT 36.911 1.792 37.125 2.17 ;
      RECT 37.055 3.452 37.1 3.645 ;
      RECT 37.045 3.422 37.055 3.645 ;
      RECT 37.04 3.407 37.045 3.645 ;
      RECT 37 3.317 37.04 3.645 ;
      RECT 36.995 3.23 37 3.645 ;
      RECT 36.985 3.2 36.995 3.645 ;
      RECT 36.98 3.16 36.985 3.645 ;
      RECT 36.97 3.122 36.98 3.645 ;
      RECT 36.965 3.087 36.97 3.645 ;
      RECT 36.945 3.04 36.965 3.645 ;
      RECT 36.93 2.965 36.945 3.645 ;
      RECT 36.925 2.92 36.93 3.64 ;
      RECT 36.92 2.9 36.925 3.613 ;
      RECT 36.915 2.88 36.92 3.598 ;
      RECT 36.91 2.855 36.915 3.578 ;
      RECT 36.905 2.833 36.91 3.563 ;
      RECT 36.9 2.811 36.905 3.545 ;
      RECT 36.895 2.79 36.9 3.535 ;
      RECT 36.885 2.762 36.895 3.505 ;
      RECT 36.875 2.725 36.885 3.473 ;
      RECT 36.865 2.685 36.875 3.44 ;
      RECT 36.855 2.663 36.865 3.41 ;
      RECT 36.825 2.615 36.855 3.342 ;
      RECT 36.81 2.575 36.825 3.269 ;
      RECT 36.8 2.575 36.81 3.235 ;
      RECT 36.795 2.575 36.8 3.21 ;
      RECT 36.79 2.575 36.795 3.195 ;
      RECT 36.785 2.575 36.79 3.173 ;
      RECT 36.78 2.575 36.785 3.16 ;
      RECT 36.765 2.575 36.78 3.125 ;
      RECT 36.745 2.575 36.765 3.065 ;
      RECT 36.735 2.575 36.745 3.015 ;
      RECT 36.715 2.575 36.735 2.963 ;
      RECT 36.695 2.575 36.715 2.92 ;
      RECT 36.685 2.575 36.695 2.908 ;
      RECT 36.655 2.575 36.685 2.895 ;
      RECT 36.625 2.596 36.655 2.875 ;
      RECT 36.615 2.624 36.625 2.855 ;
      RECT 36.6 2.641 36.615 2.823 ;
      RECT 36.595 2.655 36.6 2.79 ;
      RECT 36.59 2.663 36.595 2.763 ;
      RECT 36.585 2.671 36.59 2.725 ;
      RECT 36.59 3.195 36.595 3.53 ;
      RECT 36.555 3.182 36.59 3.529 ;
      RECT 36.485 3.122 36.555 3.528 ;
      RECT 36.405 3.065 36.485 3.527 ;
      RECT 36.27 3.025 36.405 3.526 ;
      RECT 36.27 3.212 36.605 3.515 ;
      RECT 36.23 3.212 36.605 3.505 ;
      RECT 36.23 3.23 36.61 3.5 ;
      RECT 36.23 3.32 36.615 3.49 ;
      RECT 36.225 3.015 36.39 3.47 ;
      RECT 36.22 3.015 36.39 3.213 ;
      RECT 36.22 3.172 36.585 3.213 ;
      RECT 36.22 3.16 36.58 3.213 ;
      RECT 35.36 5.02 35.53 6.49 ;
      RECT 35.36 6.315 35.535 6.485 ;
      RECT 34.99 1.74 35.16 2.93 ;
      RECT 34.99 1.74 35.46 1.91 ;
      RECT 34.99 6.97 35.46 7.14 ;
      RECT 34.99 5.95 35.16 7.14 ;
      RECT 34 1.74 34.17 2.93 ;
      RECT 34 1.74 34.47 1.91 ;
      RECT 34 6.97 34.47 7.14 ;
      RECT 34 5.95 34.17 7.14 ;
      RECT 32.15 2.635 32.32 3.865 ;
      RECT 32.205 0.855 32.375 2.805 ;
      RECT 32.15 0.575 32.32 1.025 ;
      RECT 32.15 7.855 32.32 8.305 ;
      RECT 32.205 6.075 32.375 8.025 ;
      RECT 32.15 5.015 32.32 6.245 ;
      RECT 31.63 0.575 31.8 3.865 ;
      RECT 31.63 2.075 32.035 2.405 ;
      RECT 31.63 1.235 32.035 1.565 ;
      RECT 31.63 5.015 31.8 8.305 ;
      RECT 31.63 7.315 32.035 7.645 ;
      RECT 31.63 6.475 32.035 6.805 ;
      RECT 28.965 1.975 29.695 2.215 ;
      RECT 29.507 1.77 29.695 2.215 ;
      RECT 29.335 1.782 29.71 2.209 ;
      RECT 29.25 1.797 29.73 2.194 ;
      RECT 29.25 1.812 29.735 2.184 ;
      RECT 29.205 1.832 29.75 2.176 ;
      RECT 29.182 1.867 29.765 2.13 ;
      RECT 29.096 1.89 29.77 2.09 ;
      RECT 29.096 1.908 29.78 2.06 ;
      RECT 28.965 1.977 29.785 2.023 ;
      RECT 29.01 1.92 29.78 2.06 ;
      RECT 29.096 1.872 29.765 2.13 ;
      RECT 29.182 1.841 29.75 2.176 ;
      RECT 29.205 1.822 29.735 2.184 ;
      RECT 29.25 1.795 29.71 2.209 ;
      RECT 29.335 1.777 29.695 2.215 ;
      RECT 29.421 1.771 29.695 2.215 ;
      RECT 29.507 1.766 29.64 2.215 ;
      RECT 29.593 1.761 29.64 2.215 ;
      RECT 29.285 2.659 29.455 3.045 ;
      RECT 29.28 2.659 29.455 3.04 ;
      RECT 29.255 2.659 29.455 3.005 ;
      RECT 29.255 2.687 29.465 2.995 ;
      RECT 29.235 2.687 29.465 2.955 ;
      RECT 29.23 2.687 29.465 2.928 ;
      RECT 29.23 2.705 29.47 2.92 ;
      RECT 29.175 2.705 29.47 2.855 ;
      RECT 29.175 2.722 29.48 2.838 ;
      RECT 29.165 2.722 29.48 2.778 ;
      RECT 29.165 2.739 29.485 2.775 ;
      RECT 29.16 2.575 29.33 2.753 ;
      RECT 29.16 2.609 29.416 2.753 ;
      RECT 29.155 3.375 29.16 3.388 ;
      RECT 29.15 3.27 29.155 3.393 ;
      RECT 29.125 3.13 29.15 3.408 ;
      RECT 29.09 3.081 29.125 3.44 ;
      RECT 29.085 3.049 29.09 3.46 ;
      RECT 29.08 3.04 29.085 3.46 ;
      RECT 29 3.005 29.08 3.46 ;
      RECT 28.937 2.975 29 3.46 ;
      RECT 28.851 2.963 28.937 3.46 ;
      RECT 28.765 2.949 28.851 3.46 ;
      RECT 28.685 2.936 28.765 3.446 ;
      RECT 28.65 2.928 28.685 3.426 ;
      RECT 28.64 2.925 28.65 3.417 ;
      RECT 28.61 2.92 28.64 3.404 ;
      RECT 28.56 2.895 28.61 3.38 ;
      RECT 28.546 2.869 28.56 3.362 ;
      RECT 28.46 2.829 28.546 3.338 ;
      RECT 28.415 2.777 28.46 3.307 ;
      RECT 28.405 2.752 28.415 3.294 ;
      RECT 28.4 2.533 28.405 2.555 ;
      RECT 28.395 2.735 28.405 3.29 ;
      RECT 28.395 2.531 28.4 2.645 ;
      RECT 28.385 2.527 28.395 3.286 ;
      RECT 28.341 2.525 28.385 3.274 ;
      RECT 28.255 2.525 28.341 3.245 ;
      RECT 28.225 2.525 28.255 3.218 ;
      RECT 28.21 2.525 28.225 3.206 ;
      RECT 28.17 2.537 28.21 3.191 ;
      RECT 28.15 2.556 28.17 3.17 ;
      RECT 28.14 2.566 28.15 3.154 ;
      RECT 28.13 2.572 28.14 3.143 ;
      RECT 28.11 2.582 28.13 3.126 ;
      RECT 28.105 2.591 28.11 3.113 ;
      RECT 28.1 2.595 28.105 3.063 ;
      RECT 28.09 2.601 28.1 2.98 ;
      RECT 28.085 2.605 28.09 2.894 ;
      RECT 28.08 2.625 28.085 2.831 ;
      RECT 28.075 2.648 28.08 2.778 ;
      RECT 28.07 2.666 28.075 2.723 ;
      RECT 28.68 2.485 28.85 2.745 ;
      RECT 28.85 2.45 28.895 2.731 ;
      RECT 28.811 2.452 28.9 2.714 ;
      RECT 28.7 2.469 28.986 2.685 ;
      RECT 28.7 2.484 28.99 2.657 ;
      RECT 28.7 2.465 28.9 2.714 ;
      RECT 28.725 2.453 28.85 2.745 ;
      RECT 28.811 2.451 28.895 2.731 ;
      RECT 27.865 1.84 28.035 2.33 ;
      RECT 27.865 1.84 28.07 2.31 ;
      RECT 28 1.76 28.11 2.27 ;
      RECT 27.981 1.764 28.13 2.24 ;
      RECT 27.895 1.772 28.15 2.223 ;
      RECT 27.895 1.778 28.155 2.213 ;
      RECT 27.895 1.787 28.175 2.201 ;
      RECT 27.87 1.812 28.205 2.179 ;
      RECT 27.87 1.832 28.21 2.159 ;
      RECT 27.865 1.845 28.22 2.139 ;
      RECT 27.865 1.912 28.225 2.12 ;
      RECT 27.865 2.045 28.23 2.107 ;
      RECT 27.86 1.85 28.22 1.94 ;
      RECT 27.87 1.807 28.175 2.201 ;
      RECT 27.981 1.762 28.11 2.27 ;
      RECT 27.855 3.515 28.155 3.77 ;
      RECT 27.94 3.481 28.155 3.77 ;
      RECT 27.94 3.484 28.16 3.63 ;
      RECT 27.875 3.505 28.16 3.63 ;
      RECT 27.91 3.495 28.155 3.77 ;
      RECT 27.905 3.5 28.16 3.63 ;
      RECT 27.94 3.479 28.141 3.77 ;
      RECT 28.026 3.47 28.141 3.77 ;
      RECT 28.026 3.464 28.055 3.77 ;
      RECT 27.515 3.105 27.525 3.595 ;
      RECT 27.175 3.04 27.185 3.34 ;
      RECT 27.69 3.212 27.695 3.431 ;
      RECT 27.68 3.192 27.69 3.448 ;
      RECT 27.67 3.172 27.68 3.478 ;
      RECT 27.665 3.162 27.67 3.493 ;
      RECT 27.66 3.158 27.665 3.498 ;
      RECT 27.645 3.15 27.66 3.505 ;
      RECT 27.605 3.13 27.645 3.53 ;
      RECT 27.58 3.112 27.605 3.563 ;
      RECT 27.575 3.11 27.58 3.576 ;
      RECT 27.555 3.107 27.575 3.58 ;
      RECT 27.525 3.105 27.555 3.59 ;
      RECT 27.455 3.107 27.515 3.591 ;
      RECT 27.435 3.107 27.455 3.585 ;
      RECT 27.41 3.105 27.435 3.582 ;
      RECT 27.375 3.1 27.41 3.578 ;
      RECT 27.355 3.094 27.375 3.565 ;
      RECT 27.345 3.091 27.355 3.553 ;
      RECT 27.325 3.088 27.345 3.538 ;
      RECT 27.305 3.084 27.325 3.52 ;
      RECT 27.3 3.081 27.305 3.51 ;
      RECT 27.295 3.08 27.3 3.508 ;
      RECT 27.285 3.077 27.295 3.5 ;
      RECT 27.275 3.071 27.285 3.483 ;
      RECT 27.265 3.065 27.275 3.465 ;
      RECT 27.255 3.059 27.265 3.453 ;
      RECT 27.245 3.053 27.255 3.433 ;
      RECT 27.24 3.049 27.245 3.418 ;
      RECT 27.235 3.047 27.24 3.41 ;
      RECT 27.23 3.045 27.235 3.403 ;
      RECT 27.225 3.043 27.23 3.393 ;
      RECT 27.22 3.041 27.225 3.387 ;
      RECT 27.21 3.04 27.22 3.377 ;
      RECT 27.2 3.04 27.21 3.368 ;
      RECT 27.185 3.04 27.2 3.353 ;
      RECT 27.145 3.04 27.175 3.337 ;
      RECT 27.125 3.042 27.145 3.332 ;
      RECT 27.12 3.047 27.125 3.33 ;
      RECT 27.09 3.055 27.12 3.328 ;
      RECT 27.06 3.07 27.09 3.327 ;
      RECT 27.015 3.092 27.06 3.332 ;
      RECT 27.01 3.107 27.015 3.336 ;
      RECT 26.995 3.112 27.01 3.338 ;
      RECT 26.99 3.116 26.995 3.34 ;
      RECT 26.93 3.139 26.99 3.349 ;
      RECT 26.91 3.165 26.93 3.362 ;
      RECT 26.9 3.172 26.91 3.366 ;
      RECT 26.885 3.179 26.9 3.369 ;
      RECT 26.865 3.189 26.885 3.372 ;
      RECT 26.86 3.197 26.865 3.375 ;
      RECT 26.815 3.202 26.86 3.382 ;
      RECT 26.805 3.205 26.815 3.389 ;
      RECT 26.795 3.205 26.805 3.393 ;
      RECT 26.76 3.207 26.795 3.405 ;
      RECT 26.74 3.21 26.76 3.418 ;
      RECT 26.7 3.213 26.74 3.429 ;
      RECT 26.685 3.215 26.7 3.442 ;
      RECT 26.675 3.215 26.685 3.447 ;
      RECT 26.65 3.216 26.675 3.455 ;
      RECT 26.64 3.218 26.65 3.46 ;
      RECT 26.635 3.219 26.64 3.463 ;
      RECT 26.61 3.217 26.635 3.466 ;
      RECT 26.595 3.215 26.61 3.467 ;
      RECT 26.575 3.212 26.595 3.469 ;
      RECT 26.555 3.207 26.575 3.469 ;
      RECT 26.495 3.202 26.555 3.466 ;
      RECT 26.46 3.177 26.495 3.462 ;
      RECT 26.45 3.154 26.46 3.46 ;
      RECT 26.42 3.131 26.45 3.46 ;
      RECT 26.41 3.11 26.42 3.46 ;
      RECT 26.385 3.092 26.41 3.458 ;
      RECT 26.37 3.07 26.385 3.455 ;
      RECT 26.355 3.052 26.37 3.453 ;
      RECT 26.335 3.042 26.355 3.451 ;
      RECT 26.32 3.037 26.335 3.45 ;
      RECT 26.305 3.035 26.32 3.449 ;
      RECT 26.275 3.036 26.305 3.447 ;
      RECT 26.255 3.039 26.275 3.445 ;
      RECT 26.198 3.043 26.255 3.445 ;
      RECT 26.112 3.052 26.198 3.445 ;
      RECT 26.026 3.063 26.112 3.445 ;
      RECT 25.94 3.074 26.026 3.445 ;
      RECT 25.92 3.081 25.94 3.453 ;
      RECT 25.91 3.084 25.92 3.46 ;
      RECT 25.845 3.089 25.91 3.478 ;
      RECT 25.815 3.096 25.845 3.503 ;
      RECT 25.805 3.099 25.815 3.51 ;
      RECT 25.76 3.103 25.805 3.515 ;
      RECT 25.73 3.108 25.76 3.52 ;
      RECT 25.729 3.11 25.73 3.52 ;
      RECT 25.643 3.116 25.729 3.52 ;
      RECT 25.557 3.127 25.643 3.52 ;
      RECT 25.471 3.139 25.557 3.52 ;
      RECT 25.385 3.15 25.471 3.52 ;
      RECT 25.37 3.157 25.385 3.515 ;
      RECT 25.365 3.159 25.37 3.509 ;
      RECT 25.345 3.17 25.365 3.504 ;
      RECT 25.335 3.188 25.345 3.498 ;
      RECT 25.33 3.2 25.335 3.298 ;
      RECT 27.625 1.953 27.645 2.04 ;
      RECT 27.62 1.888 27.625 2.072 ;
      RECT 27.61 1.855 27.62 2.077 ;
      RECT 27.605 1.835 27.61 2.083 ;
      RECT 27.575 1.835 27.605 2.1 ;
      RECT 27.526 1.835 27.575 2.136 ;
      RECT 27.44 1.835 27.526 2.194 ;
      RECT 27.411 1.845 27.44 2.243 ;
      RECT 27.325 1.887 27.411 2.296 ;
      RECT 27.305 1.925 27.325 2.343 ;
      RECT 27.28 1.942 27.305 2.363 ;
      RECT 27.27 1.956 27.28 2.383 ;
      RECT 27.265 1.962 27.27 2.393 ;
      RECT 27.26 1.966 27.265 2.4 ;
      RECT 27.21 1.986 27.26 2.405 ;
      RECT 27.145 2.03 27.21 2.405 ;
      RECT 27.12 2.08 27.145 2.405 ;
      RECT 27.11 2.11 27.12 2.405 ;
      RECT 27.105 2.137 27.11 2.405 ;
      RECT 27.1 2.155 27.105 2.405 ;
      RECT 27.09 2.197 27.1 2.405 ;
      RECT 27.44 2.755 27.61 2.93 ;
      RECT 27.38 2.583 27.44 2.918 ;
      RECT 27.37 2.576 27.38 2.901 ;
      RECT 27.325 2.755 27.61 2.881 ;
      RECT 27.306 2.755 27.61 2.859 ;
      RECT 27.22 2.755 27.61 2.824 ;
      RECT 27.2 2.575 27.37 2.78 ;
      RECT 27.2 2.722 27.605 2.78 ;
      RECT 27.2 2.67 27.58 2.78 ;
      RECT 27.2 2.625 27.545 2.78 ;
      RECT 27.2 2.607 27.51 2.78 ;
      RECT 27.2 2.597 27.505 2.78 ;
      RECT 27.37 7.855 27.54 8.305 ;
      RECT 27.425 6.075 27.595 8.025 ;
      RECT 27.37 5.015 27.54 6.245 ;
      RECT 26.85 5.015 27.02 8.305 ;
      RECT 26.85 7.315 27.255 7.645 ;
      RECT 26.85 6.475 27.255 6.805 ;
      RECT 26.92 3.555 27.11 3.78 ;
      RECT 26.91 3.556 27.115 3.775 ;
      RECT 26.91 3.558 27.125 3.755 ;
      RECT 26.91 3.562 27.13 3.74 ;
      RECT 26.91 3.549 27.08 3.775 ;
      RECT 26.91 3.552 27.105 3.775 ;
      RECT 26.92 3.548 27.08 3.78 ;
      RECT 27.006 3.546 27.08 3.78 ;
      RECT 26.63 2.797 26.8 3.035 ;
      RECT 26.63 2.797 26.886 2.949 ;
      RECT 26.63 2.797 26.89 2.859 ;
      RECT 26.68 2.57 26.9 2.838 ;
      RECT 26.675 2.587 26.905 2.811 ;
      RECT 26.64 2.745 26.905 2.811 ;
      RECT 26.66 2.595 26.8 3.035 ;
      RECT 26.65 2.677 26.91 2.794 ;
      RECT 26.645 2.725 26.91 2.794 ;
      RECT 26.65 2.635 26.905 2.811 ;
      RECT 26.675 2.572 26.9 2.838 ;
      RECT 26.24 2.547 26.41 2.745 ;
      RECT 26.24 2.547 26.455 2.72 ;
      RECT 26.31 2.49 26.48 2.678 ;
      RECT 26.285 2.505 26.48 2.678 ;
      RECT 25.9 2.551 25.93 2.745 ;
      RECT 25.895 2.523 25.9 2.745 ;
      RECT 25.865 2.497 25.895 2.747 ;
      RECT 25.84 2.455 25.865 2.75 ;
      RECT 25.83 2.427 25.84 2.752 ;
      RECT 25.795 2.407 25.83 2.754 ;
      RECT 25.73 2.392 25.795 2.76 ;
      RECT 25.68 2.39 25.73 2.766 ;
      RECT 25.657 2.392 25.68 2.771 ;
      RECT 25.571 2.403 25.657 2.777 ;
      RECT 25.485 2.421 25.571 2.787 ;
      RECT 25.47 2.432 25.485 2.793 ;
      RECT 25.4 2.455 25.47 2.799 ;
      RECT 25.345 2.487 25.4 2.807 ;
      RECT 25.305 2.51 25.345 2.813 ;
      RECT 25.291 2.523 25.305 2.816 ;
      RECT 25.205 2.545 25.291 2.822 ;
      RECT 25.19 2.57 25.205 2.828 ;
      RECT 25.15 2.585 25.19 2.832 ;
      RECT 25.1 2.6 25.15 2.837 ;
      RECT 25.075 2.607 25.1 2.841 ;
      RECT 25.015 2.602 25.075 2.845 ;
      RECT 25 2.593 25.015 2.849 ;
      RECT 24.93 2.583 25 2.845 ;
      RECT 24.905 2.575 24.925 2.835 ;
      RECT 24.846 2.575 24.905 2.813 ;
      RECT 24.76 2.575 24.846 2.77 ;
      RECT 24.925 2.575 24.93 2.84 ;
      RECT 25.62 1.806 25.79 2.14 ;
      RECT 25.59 1.806 25.79 2.135 ;
      RECT 25.53 1.773 25.59 2.123 ;
      RECT 25.53 1.829 25.8 2.118 ;
      RECT 25.505 1.829 25.8 2.112 ;
      RECT 25.5 1.77 25.53 2.109 ;
      RECT 25.485 1.776 25.62 2.107 ;
      RECT 25.48 1.784 25.705 2.095 ;
      RECT 25.48 1.836 25.815 2.048 ;
      RECT 25.465 1.792 25.705 2.043 ;
      RECT 25.465 1.862 25.825 1.984 ;
      RECT 25.435 1.812 25.79 1.945 ;
      RECT 25.435 1.902 25.835 1.941 ;
      RECT 25.485 1.781 25.705 2.107 ;
      RECT 24.825 2.111 24.88 2.375 ;
      RECT 24.825 2.111 24.945 2.374 ;
      RECT 24.825 2.111 24.97 2.373 ;
      RECT 24.825 2.111 25.035 2.372 ;
      RECT 24.97 2.077 25.05 2.371 ;
      RECT 24.785 2.121 25.195 2.37 ;
      RECT 24.825 2.118 25.195 2.37 ;
      RECT 24.785 2.126 25.2 2.363 ;
      RECT 24.77 2.128 25.2 2.362 ;
      RECT 24.77 2.135 25.205 2.358 ;
      RECT 24.75 2.134 25.2 2.354 ;
      RECT 24.75 2.142 25.21 2.353 ;
      RECT 24.745 2.139 25.205 2.349 ;
      RECT 24.745 2.152 25.22 2.348 ;
      RECT 24.73 2.142 25.21 2.347 ;
      RECT 24.695 2.155 25.22 2.34 ;
      RECT 24.88 2.11 25.19 2.37 ;
      RECT 24.88 2.095 25.14 2.37 ;
      RECT 24.945 2.082 25.075 2.37 ;
      RECT 24.49 3.171 24.505 3.564 ;
      RECT 24.455 3.176 24.505 3.563 ;
      RECT 24.49 3.175 24.55 3.562 ;
      RECT 24.435 3.186 24.55 3.561 ;
      RECT 24.45 3.182 24.55 3.561 ;
      RECT 24.415 3.192 24.625 3.558 ;
      RECT 24.415 3.211 24.67 3.556 ;
      RECT 24.415 3.218 24.675 3.553 ;
      RECT 24.4 3.195 24.625 3.55 ;
      RECT 24.38 3.2 24.625 3.543 ;
      RECT 24.375 3.204 24.625 3.539 ;
      RECT 24.375 3.221 24.685 3.538 ;
      RECT 24.355 3.215 24.67 3.534 ;
      RECT 24.355 3.224 24.69 3.528 ;
      RECT 24.35 3.23 24.69 3.3 ;
      RECT 24.415 3.19 24.55 3.558 ;
      RECT 24.29 2.553 24.49 2.865 ;
      RECT 24.365 2.531 24.49 2.865 ;
      RECT 24.305 2.55 24.495 2.85 ;
      RECT 24.275 2.561 24.495 2.848 ;
      RECT 24.29 2.556 24.5 2.814 ;
      RECT 24.275 2.66 24.505 2.781 ;
      RECT 24.305 2.532 24.49 2.865 ;
      RECT 24.365 2.51 24.465 2.865 ;
      RECT 24.39 2.507 24.465 2.865 ;
      RECT 24.39 2.502 24.41 2.865 ;
      RECT 23.795 2.57 23.97 2.745 ;
      RECT 23.79 2.57 23.97 2.743 ;
      RECT 23.765 2.57 23.97 2.738 ;
      RECT 23.71 2.55 23.88 2.728 ;
      RECT 23.71 2.557 23.945 2.728 ;
      RECT 23.795 3.237 23.81 3.42 ;
      RECT 23.785 3.215 23.795 3.42 ;
      RECT 23.77 3.195 23.785 3.42 ;
      RECT 23.76 3.17 23.77 3.42 ;
      RECT 23.73 3.135 23.76 3.42 ;
      RECT 23.695 3.075 23.73 3.42 ;
      RECT 23.69 3.037 23.695 3.42 ;
      RECT 23.64 2.988 23.69 3.42 ;
      RECT 23.63 2.938 23.64 3.408 ;
      RECT 23.615 2.917 23.63 3.368 ;
      RECT 23.595 2.885 23.615 3.318 ;
      RECT 23.57 2.841 23.595 3.258 ;
      RECT 23.565 2.813 23.57 3.213 ;
      RECT 23.56 2.804 23.565 3.199 ;
      RECT 23.555 2.797 23.56 3.186 ;
      RECT 23.55 2.792 23.555 3.175 ;
      RECT 23.545 2.777 23.55 3.165 ;
      RECT 23.54 2.755 23.545 3.152 ;
      RECT 23.53 2.715 23.54 3.127 ;
      RECT 23.505 2.645 23.53 3.083 ;
      RECT 23.5 2.585 23.505 3.048 ;
      RECT 23.485 2.565 23.5 3.015 ;
      RECT 23.48 2.565 23.485 2.99 ;
      RECT 23.45 2.565 23.48 2.945 ;
      RECT 23.405 2.565 23.45 2.885 ;
      RECT 23.33 2.565 23.405 2.833 ;
      RECT 23.325 2.565 23.33 2.798 ;
      RECT 23.32 2.565 23.325 2.788 ;
      RECT 23.315 2.565 23.32 2.768 ;
      RECT 23.58 1.785 23.75 2.255 ;
      RECT 23.525 1.778 23.72 2.239 ;
      RECT 23.525 1.792 23.755 2.238 ;
      RECT 23.51 1.793 23.755 2.219 ;
      RECT 23.505 1.811 23.755 2.205 ;
      RECT 23.51 1.794 23.76 2.203 ;
      RECT 23.495 1.825 23.76 2.188 ;
      RECT 23.51 1.8 23.765 2.173 ;
      RECT 23.49 1.84 23.765 2.17 ;
      RECT 23.505 1.812 23.77 2.155 ;
      RECT 23.505 1.824 23.775 2.135 ;
      RECT 23.49 1.84 23.78 2.118 ;
      RECT 23.49 1.85 23.785 1.973 ;
      RECT 23.485 1.85 23.785 1.93 ;
      RECT 23.485 1.865 23.79 1.908 ;
      RECT 23.58 1.775 23.72 2.255 ;
      RECT 23.58 1.773 23.69 2.255 ;
      RECT 23.666 1.77 23.69 2.255 ;
      RECT 23.325 3.437 23.33 3.483 ;
      RECT 23.315 3.285 23.325 3.507 ;
      RECT 23.31 3.13 23.315 3.532 ;
      RECT 23.295 3.092 23.31 3.543 ;
      RECT 23.29 3.075 23.295 3.55 ;
      RECT 23.28 3.063 23.29 3.557 ;
      RECT 23.275 3.054 23.28 3.559 ;
      RECT 23.27 3.052 23.275 3.563 ;
      RECT 23.225 3.043 23.27 3.578 ;
      RECT 23.22 3.035 23.225 3.592 ;
      RECT 23.215 3.032 23.22 3.596 ;
      RECT 23.2 3.027 23.215 3.604 ;
      RECT 23.145 3.017 23.2 3.615 ;
      RECT 23.11 3.005 23.145 3.616 ;
      RECT 23.101 3 23.11 3.61 ;
      RECT 23.015 3 23.101 3.6 ;
      RECT 22.985 3 23.015 3.578 ;
      RECT 22.975 3 22.98 3.558 ;
      RECT 22.97 3 22.975 3.52 ;
      RECT 22.965 3 22.97 3.478 ;
      RECT 22.96 3 22.965 3.438 ;
      RECT 22.955 3 22.96 3.368 ;
      RECT 22.945 3 22.955 3.29 ;
      RECT 22.94 3 22.945 3.19 ;
      RECT 22.98 3 22.985 3.56 ;
      RECT 22.475 3.082 22.565 3.56 ;
      RECT 22.46 3.085 22.58 3.558 ;
      RECT 22.475 3.084 22.58 3.558 ;
      RECT 22.44 3.091 22.605 3.548 ;
      RECT 22.46 3.085 22.605 3.548 ;
      RECT 22.425 3.097 22.605 3.536 ;
      RECT 22.46 3.088 22.655 3.529 ;
      RECT 22.411 3.105 22.655 3.527 ;
      RECT 22.44 3.095 22.665 3.515 ;
      RECT 22.411 3.116 22.695 3.506 ;
      RECT 22.325 3.14 22.695 3.5 ;
      RECT 22.325 3.153 22.735 3.483 ;
      RECT 22.32 3.175 22.735 3.476 ;
      RECT 22.29 3.19 22.735 3.466 ;
      RECT 22.285 3.201 22.735 3.456 ;
      RECT 22.255 3.214 22.735 3.447 ;
      RECT 22.24 3.232 22.735 3.436 ;
      RECT 22.215 3.245 22.735 3.426 ;
      RECT 22.475 3.081 22.485 3.56 ;
      RECT 22.521 2.505 22.56 2.75 ;
      RECT 22.435 2.505 22.57 2.748 ;
      RECT 22.32 2.53 22.57 2.745 ;
      RECT 22.32 2.53 22.575 2.743 ;
      RECT 22.32 2.53 22.59 2.738 ;
      RECT 22.426 2.505 22.605 2.718 ;
      RECT 22.34 2.513 22.605 2.718 ;
      RECT 22.01 1.865 22.18 2.3 ;
      RECT 22 1.899 22.18 2.283 ;
      RECT 22.08 1.835 22.25 2.27 ;
      RECT 21.985 1.91 22.25 2.248 ;
      RECT 22.08 1.845 22.255 2.238 ;
      RECT 22.01 1.897 22.285 2.223 ;
      RECT 21.97 1.923 22.285 2.208 ;
      RECT 21.97 1.965 22.295 2.188 ;
      RECT 21.965 1.99 22.3 2.17 ;
      RECT 21.965 2 22.305 2.155 ;
      RECT 21.96 1.937 22.285 2.153 ;
      RECT 21.96 2.01 22.31 2.138 ;
      RECT 21.955 1.947 22.285 2.135 ;
      RECT 21.95 2.031 22.315 2.118 ;
      RECT 21.95 2.063 22.32 2.098 ;
      RECT 21.945 1.977 22.295 2.09 ;
      RECT 21.95 1.962 22.285 2.118 ;
      RECT 21.965 1.932 22.285 2.17 ;
      RECT 21.81 2.519 22.035 2.775 ;
      RECT 21.81 2.552 22.055 2.765 ;
      RECT 21.775 2.552 22.055 2.763 ;
      RECT 21.775 2.565 22.06 2.753 ;
      RECT 21.775 2.585 22.07 2.745 ;
      RECT 21.775 2.682 22.075 2.738 ;
      RECT 21.755 2.43 21.885 2.728 ;
      RECT 21.71 2.585 22.07 2.67 ;
      RECT 21.7 2.43 21.885 2.615 ;
      RECT 21.7 2.462 21.971 2.615 ;
      RECT 21.665 2.992 21.685 3.17 ;
      RECT 21.63 2.945 21.665 3.17 ;
      RECT 21.615 2.885 21.63 3.17 ;
      RECT 21.59 2.832 21.615 3.17 ;
      RECT 21.575 2.785 21.59 3.17 ;
      RECT 21.555 2.762 21.575 3.17 ;
      RECT 21.53 2.727 21.555 3.17 ;
      RECT 21.52 2.573 21.53 3.17 ;
      RECT 21.49 2.568 21.52 3.161 ;
      RECT 21.485 2.565 21.49 3.151 ;
      RECT 21.47 2.565 21.485 3.125 ;
      RECT 21.465 2.565 21.47 3.088 ;
      RECT 21.44 2.565 21.465 3.04 ;
      RECT 21.42 2.565 21.44 2.965 ;
      RECT 21.41 2.565 21.42 2.925 ;
      RECT 21.405 2.565 21.41 2.9 ;
      RECT 21.4 2.565 21.405 2.883 ;
      RECT 21.395 2.565 21.4 2.865 ;
      RECT 21.39 2.566 21.395 2.855 ;
      RECT 21.38 2.568 21.39 2.823 ;
      RECT 21.37 2.57 21.38 2.79 ;
      RECT 21.36 2.573 21.37 2.763 ;
      RECT 21.685 3 21.91 3.17 ;
      RECT 21.015 1.812 21.185 2.265 ;
      RECT 21.015 1.812 21.275 2.231 ;
      RECT 21.015 1.812 21.305 2.215 ;
      RECT 21.015 1.812 21.335 2.188 ;
      RECT 21.271 1.79 21.35 2.17 ;
      RECT 21.05 1.797 21.355 2.155 ;
      RECT 21.05 1.805 21.365 2.118 ;
      RECT 21.01 1.832 21.365 2.09 ;
      RECT 20.995 1.845 21.365 2.055 ;
      RECT 21.015 1.82 21.385 2.045 ;
      RECT 20.99 1.885 21.385 2.015 ;
      RECT 20.99 1.915 21.39 1.998 ;
      RECT 20.985 1.945 21.39 1.985 ;
      RECT 21.05 1.794 21.35 2.17 ;
      RECT 21.185 1.791 21.271 2.249 ;
      RECT 21.136 1.792 21.35 2.17 ;
      RECT 21.28 3.452 21.325 3.645 ;
      RECT 21.27 3.422 21.28 3.645 ;
      RECT 21.265 3.407 21.27 3.645 ;
      RECT 21.225 3.317 21.265 3.645 ;
      RECT 21.22 3.23 21.225 3.645 ;
      RECT 21.21 3.2 21.22 3.645 ;
      RECT 21.205 3.16 21.21 3.645 ;
      RECT 21.195 3.122 21.205 3.645 ;
      RECT 21.19 3.087 21.195 3.645 ;
      RECT 21.17 3.04 21.19 3.645 ;
      RECT 21.155 2.965 21.17 3.645 ;
      RECT 21.15 2.92 21.155 3.64 ;
      RECT 21.145 2.9 21.15 3.613 ;
      RECT 21.14 2.88 21.145 3.598 ;
      RECT 21.135 2.855 21.14 3.578 ;
      RECT 21.13 2.833 21.135 3.563 ;
      RECT 21.125 2.811 21.13 3.545 ;
      RECT 21.12 2.79 21.125 3.535 ;
      RECT 21.11 2.762 21.12 3.505 ;
      RECT 21.1 2.725 21.11 3.473 ;
      RECT 21.09 2.685 21.1 3.44 ;
      RECT 21.08 2.663 21.09 3.41 ;
      RECT 21.05 2.615 21.08 3.342 ;
      RECT 21.035 2.575 21.05 3.269 ;
      RECT 21.025 2.575 21.035 3.235 ;
      RECT 21.02 2.575 21.025 3.21 ;
      RECT 21.015 2.575 21.02 3.195 ;
      RECT 21.01 2.575 21.015 3.173 ;
      RECT 21.005 2.575 21.01 3.16 ;
      RECT 20.99 2.575 21.005 3.125 ;
      RECT 20.97 2.575 20.99 3.065 ;
      RECT 20.96 2.575 20.97 3.015 ;
      RECT 20.94 2.575 20.96 2.963 ;
      RECT 20.92 2.575 20.94 2.92 ;
      RECT 20.91 2.575 20.92 2.908 ;
      RECT 20.88 2.575 20.91 2.895 ;
      RECT 20.85 2.596 20.88 2.875 ;
      RECT 20.84 2.624 20.85 2.855 ;
      RECT 20.825 2.641 20.84 2.823 ;
      RECT 20.82 2.655 20.825 2.79 ;
      RECT 20.815 2.663 20.82 2.763 ;
      RECT 20.81 2.671 20.815 2.725 ;
      RECT 20.815 3.195 20.82 3.53 ;
      RECT 20.78 3.182 20.815 3.529 ;
      RECT 20.71 3.122 20.78 3.528 ;
      RECT 20.63 3.065 20.71 3.527 ;
      RECT 20.495 3.025 20.63 3.526 ;
      RECT 20.495 3.212 20.83 3.515 ;
      RECT 20.455 3.212 20.83 3.505 ;
      RECT 20.455 3.23 20.835 3.5 ;
      RECT 20.455 3.32 20.84 3.49 ;
      RECT 20.45 3.015 20.615 3.47 ;
      RECT 20.445 3.015 20.615 3.213 ;
      RECT 20.445 3.172 20.81 3.213 ;
      RECT 20.445 3.16 20.805 3.213 ;
      RECT 19.58 5.02 19.75 6.49 ;
      RECT 19.58 6.315 19.755 6.485 ;
      RECT 19.21 1.74 19.38 2.93 ;
      RECT 19.21 1.74 19.68 1.91 ;
      RECT 19.21 6.97 19.68 7.14 ;
      RECT 19.21 5.95 19.38 7.14 ;
      RECT 18.22 1.74 18.39 2.93 ;
      RECT 18.22 1.74 18.69 1.91 ;
      RECT 18.22 6.97 18.69 7.14 ;
      RECT 18.22 5.95 18.39 7.14 ;
      RECT 16.37 2.635 16.54 3.865 ;
      RECT 16.425 0.855 16.595 2.805 ;
      RECT 16.37 0.575 16.54 1.025 ;
      RECT 16.37 7.855 16.54 8.305 ;
      RECT 16.425 6.075 16.595 8.025 ;
      RECT 16.37 5.015 16.54 6.245 ;
      RECT 15.85 0.575 16.02 3.865 ;
      RECT 15.85 2.075 16.255 2.405 ;
      RECT 15.85 1.235 16.255 1.565 ;
      RECT 15.85 5.015 16.02 8.305 ;
      RECT 15.85 7.315 16.255 7.645 ;
      RECT 15.85 6.475 16.255 6.805 ;
      RECT 13.185 1.975 13.915 2.215 ;
      RECT 13.727 1.77 13.915 2.215 ;
      RECT 13.555 1.782 13.93 2.209 ;
      RECT 13.47 1.797 13.95 2.194 ;
      RECT 13.47 1.812 13.955 2.184 ;
      RECT 13.425 1.832 13.97 2.176 ;
      RECT 13.402 1.867 13.985 2.13 ;
      RECT 13.316 1.89 13.99 2.09 ;
      RECT 13.316 1.908 14 2.06 ;
      RECT 13.185 1.977 14.005 2.023 ;
      RECT 13.23 1.92 14 2.06 ;
      RECT 13.316 1.872 13.985 2.13 ;
      RECT 13.402 1.841 13.97 2.176 ;
      RECT 13.425 1.822 13.955 2.184 ;
      RECT 13.47 1.795 13.93 2.209 ;
      RECT 13.555 1.777 13.915 2.215 ;
      RECT 13.641 1.771 13.915 2.215 ;
      RECT 13.727 1.766 13.86 2.215 ;
      RECT 13.813 1.761 13.86 2.215 ;
      RECT 13.505 2.659 13.675 3.045 ;
      RECT 13.5 2.659 13.675 3.04 ;
      RECT 13.475 2.659 13.675 3.005 ;
      RECT 13.475 2.687 13.685 2.995 ;
      RECT 13.455 2.687 13.685 2.955 ;
      RECT 13.45 2.687 13.685 2.928 ;
      RECT 13.45 2.705 13.69 2.92 ;
      RECT 13.395 2.705 13.69 2.855 ;
      RECT 13.395 2.722 13.7 2.838 ;
      RECT 13.385 2.722 13.7 2.778 ;
      RECT 13.385 2.739 13.705 2.775 ;
      RECT 13.38 2.575 13.55 2.753 ;
      RECT 13.38 2.609 13.636 2.753 ;
      RECT 13.375 3.375 13.38 3.388 ;
      RECT 13.37 3.27 13.375 3.393 ;
      RECT 13.345 3.13 13.37 3.408 ;
      RECT 13.31 3.081 13.345 3.44 ;
      RECT 13.305 3.049 13.31 3.46 ;
      RECT 13.3 3.04 13.305 3.46 ;
      RECT 13.22 3.005 13.3 3.46 ;
      RECT 13.157 2.975 13.22 3.46 ;
      RECT 13.071 2.963 13.157 3.46 ;
      RECT 12.985 2.949 13.071 3.46 ;
      RECT 12.905 2.936 12.985 3.446 ;
      RECT 12.87 2.928 12.905 3.426 ;
      RECT 12.86 2.925 12.87 3.417 ;
      RECT 12.83 2.92 12.86 3.404 ;
      RECT 12.78 2.895 12.83 3.38 ;
      RECT 12.766 2.869 12.78 3.362 ;
      RECT 12.68 2.829 12.766 3.338 ;
      RECT 12.635 2.777 12.68 3.307 ;
      RECT 12.625 2.752 12.635 3.294 ;
      RECT 12.62 2.533 12.625 2.555 ;
      RECT 12.615 2.735 12.625 3.29 ;
      RECT 12.615 2.531 12.62 2.645 ;
      RECT 12.605 2.527 12.615 3.286 ;
      RECT 12.561 2.525 12.605 3.274 ;
      RECT 12.475 2.525 12.561 3.245 ;
      RECT 12.445 2.525 12.475 3.218 ;
      RECT 12.43 2.525 12.445 3.206 ;
      RECT 12.39 2.537 12.43 3.191 ;
      RECT 12.37 2.556 12.39 3.17 ;
      RECT 12.36 2.566 12.37 3.154 ;
      RECT 12.35 2.572 12.36 3.143 ;
      RECT 12.33 2.582 12.35 3.126 ;
      RECT 12.325 2.591 12.33 3.113 ;
      RECT 12.32 2.595 12.325 3.063 ;
      RECT 12.31 2.601 12.32 2.98 ;
      RECT 12.305 2.605 12.31 2.894 ;
      RECT 12.3 2.625 12.305 2.831 ;
      RECT 12.295 2.648 12.3 2.778 ;
      RECT 12.29 2.666 12.295 2.723 ;
      RECT 12.9 2.485 13.07 2.745 ;
      RECT 13.07 2.45 13.115 2.731 ;
      RECT 13.031 2.452 13.12 2.714 ;
      RECT 12.92 2.469 13.206 2.685 ;
      RECT 12.92 2.484 13.21 2.657 ;
      RECT 12.92 2.465 13.12 2.714 ;
      RECT 12.945 2.453 13.07 2.745 ;
      RECT 13.031 2.451 13.115 2.731 ;
      RECT 12.085 1.84 12.255 2.33 ;
      RECT 12.085 1.84 12.29 2.31 ;
      RECT 12.22 1.76 12.33 2.27 ;
      RECT 12.201 1.764 12.35 2.24 ;
      RECT 12.115 1.772 12.37 2.223 ;
      RECT 12.115 1.778 12.375 2.213 ;
      RECT 12.115 1.787 12.395 2.201 ;
      RECT 12.09 1.812 12.425 2.179 ;
      RECT 12.09 1.832 12.43 2.159 ;
      RECT 12.085 1.845 12.44 2.139 ;
      RECT 12.085 1.912 12.445 2.12 ;
      RECT 12.085 2.045 12.45 2.107 ;
      RECT 12.08 1.85 12.44 1.94 ;
      RECT 12.09 1.807 12.395 2.201 ;
      RECT 12.201 1.762 12.33 2.27 ;
      RECT 12.075 3.515 12.375 3.77 ;
      RECT 12.16 3.481 12.375 3.77 ;
      RECT 12.16 3.484 12.38 3.63 ;
      RECT 12.095 3.505 12.38 3.63 ;
      RECT 12.13 3.495 12.375 3.77 ;
      RECT 12.125 3.5 12.38 3.63 ;
      RECT 12.16 3.479 12.361 3.77 ;
      RECT 12.246 3.47 12.361 3.77 ;
      RECT 12.246 3.464 12.275 3.77 ;
      RECT 11.735 3.105 11.745 3.595 ;
      RECT 11.395 3.04 11.405 3.34 ;
      RECT 11.91 3.212 11.915 3.431 ;
      RECT 11.9 3.192 11.91 3.448 ;
      RECT 11.89 3.172 11.9 3.478 ;
      RECT 11.885 3.162 11.89 3.493 ;
      RECT 11.88 3.158 11.885 3.498 ;
      RECT 11.865 3.15 11.88 3.505 ;
      RECT 11.825 3.13 11.865 3.53 ;
      RECT 11.8 3.112 11.825 3.563 ;
      RECT 11.795 3.11 11.8 3.576 ;
      RECT 11.775 3.107 11.795 3.58 ;
      RECT 11.745 3.105 11.775 3.59 ;
      RECT 11.675 3.107 11.735 3.591 ;
      RECT 11.655 3.107 11.675 3.585 ;
      RECT 11.63 3.105 11.655 3.582 ;
      RECT 11.595 3.1 11.63 3.578 ;
      RECT 11.575 3.094 11.595 3.565 ;
      RECT 11.565 3.091 11.575 3.553 ;
      RECT 11.545 3.088 11.565 3.538 ;
      RECT 11.525 3.084 11.545 3.52 ;
      RECT 11.52 3.081 11.525 3.51 ;
      RECT 11.515 3.08 11.52 3.508 ;
      RECT 11.505 3.077 11.515 3.5 ;
      RECT 11.495 3.071 11.505 3.483 ;
      RECT 11.485 3.065 11.495 3.465 ;
      RECT 11.475 3.059 11.485 3.453 ;
      RECT 11.465 3.053 11.475 3.433 ;
      RECT 11.46 3.049 11.465 3.418 ;
      RECT 11.455 3.047 11.46 3.41 ;
      RECT 11.45 3.045 11.455 3.403 ;
      RECT 11.445 3.043 11.45 3.393 ;
      RECT 11.44 3.041 11.445 3.387 ;
      RECT 11.43 3.04 11.44 3.377 ;
      RECT 11.42 3.04 11.43 3.368 ;
      RECT 11.405 3.04 11.42 3.353 ;
      RECT 11.365 3.04 11.395 3.337 ;
      RECT 11.345 3.042 11.365 3.332 ;
      RECT 11.34 3.047 11.345 3.33 ;
      RECT 11.31 3.055 11.34 3.328 ;
      RECT 11.28 3.07 11.31 3.327 ;
      RECT 11.235 3.092 11.28 3.332 ;
      RECT 11.23 3.107 11.235 3.336 ;
      RECT 11.215 3.112 11.23 3.338 ;
      RECT 11.21 3.116 11.215 3.34 ;
      RECT 11.15 3.139 11.21 3.349 ;
      RECT 11.13 3.165 11.15 3.362 ;
      RECT 11.12 3.172 11.13 3.366 ;
      RECT 11.105 3.179 11.12 3.369 ;
      RECT 11.085 3.189 11.105 3.372 ;
      RECT 11.08 3.197 11.085 3.375 ;
      RECT 11.035 3.202 11.08 3.382 ;
      RECT 11.025 3.205 11.035 3.389 ;
      RECT 11.015 3.205 11.025 3.393 ;
      RECT 10.98 3.207 11.015 3.405 ;
      RECT 10.96 3.21 10.98 3.418 ;
      RECT 10.92 3.213 10.96 3.429 ;
      RECT 10.905 3.215 10.92 3.442 ;
      RECT 10.895 3.215 10.905 3.447 ;
      RECT 10.87 3.216 10.895 3.455 ;
      RECT 10.86 3.218 10.87 3.46 ;
      RECT 10.855 3.219 10.86 3.463 ;
      RECT 10.83 3.217 10.855 3.466 ;
      RECT 10.815 3.215 10.83 3.467 ;
      RECT 10.795 3.212 10.815 3.469 ;
      RECT 10.775 3.207 10.795 3.469 ;
      RECT 10.715 3.202 10.775 3.466 ;
      RECT 10.68 3.177 10.715 3.462 ;
      RECT 10.67 3.154 10.68 3.46 ;
      RECT 10.64 3.131 10.67 3.46 ;
      RECT 10.63 3.11 10.64 3.46 ;
      RECT 10.605 3.092 10.63 3.458 ;
      RECT 10.59 3.07 10.605 3.455 ;
      RECT 10.575 3.052 10.59 3.453 ;
      RECT 10.555 3.042 10.575 3.451 ;
      RECT 10.54 3.037 10.555 3.45 ;
      RECT 10.525 3.035 10.54 3.449 ;
      RECT 10.495 3.036 10.525 3.447 ;
      RECT 10.475 3.039 10.495 3.445 ;
      RECT 10.418 3.043 10.475 3.445 ;
      RECT 10.332 3.052 10.418 3.445 ;
      RECT 10.246 3.063 10.332 3.445 ;
      RECT 10.16 3.074 10.246 3.445 ;
      RECT 10.14 3.081 10.16 3.453 ;
      RECT 10.13 3.084 10.14 3.46 ;
      RECT 10.065 3.089 10.13 3.478 ;
      RECT 10.035 3.096 10.065 3.503 ;
      RECT 10.025 3.099 10.035 3.51 ;
      RECT 9.98 3.103 10.025 3.515 ;
      RECT 9.95 3.108 9.98 3.52 ;
      RECT 9.949 3.11 9.95 3.52 ;
      RECT 9.863 3.116 9.949 3.52 ;
      RECT 9.777 3.127 9.863 3.52 ;
      RECT 9.691 3.139 9.777 3.52 ;
      RECT 9.605 3.15 9.691 3.52 ;
      RECT 9.59 3.157 9.605 3.515 ;
      RECT 9.585 3.159 9.59 3.509 ;
      RECT 9.565 3.17 9.585 3.504 ;
      RECT 9.555 3.188 9.565 3.498 ;
      RECT 9.55 3.2 9.555 3.298 ;
      RECT 11.845 1.953 11.865 2.04 ;
      RECT 11.84 1.888 11.845 2.072 ;
      RECT 11.83 1.855 11.84 2.077 ;
      RECT 11.825 1.835 11.83 2.083 ;
      RECT 11.795 1.835 11.825 2.1 ;
      RECT 11.746 1.835 11.795 2.136 ;
      RECT 11.66 1.835 11.746 2.194 ;
      RECT 11.631 1.845 11.66 2.243 ;
      RECT 11.545 1.887 11.631 2.296 ;
      RECT 11.525 1.925 11.545 2.343 ;
      RECT 11.5 1.942 11.525 2.363 ;
      RECT 11.49 1.956 11.5 2.383 ;
      RECT 11.485 1.962 11.49 2.393 ;
      RECT 11.48 1.966 11.485 2.4 ;
      RECT 11.43 1.986 11.48 2.405 ;
      RECT 11.365 2.03 11.43 2.405 ;
      RECT 11.34 2.08 11.365 2.405 ;
      RECT 11.33 2.11 11.34 2.405 ;
      RECT 11.325 2.137 11.33 2.405 ;
      RECT 11.32 2.155 11.325 2.405 ;
      RECT 11.31 2.197 11.32 2.405 ;
      RECT 11.66 2.755 11.83 2.93 ;
      RECT 11.6 2.583 11.66 2.918 ;
      RECT 11.59 2.576 11.6 2.901 ;
      RECT 11.545 2.755 11.83 2.881 ;
      RECT 11.526 2.755 11.83 2.859 ;
      RECT 11.44 2.755 11.83 2.824 ;
      RECT 11.42 2.575 11.59 2.78 ;
      RECT 11.42 2.722 11.825 2.78 ;
      RECT 11.42 2.67 11.8 2.78 ;
      RECT 11.42 2.625 11.765 2.78 ;
      RECT 11.42 2.607 11.73 2.78 ;
      RECT 11.42 2.597 11.725 2.78 ;
      RECT 11.59 7.855 11.76 8.305 ;
      RECT 11.645 6.075 11.815 8.025 ;
      RECT 11.59 5.015 11.76 6.245 ;
      RECT 11.07 5.015 11.24 8.305 ;
      RECT 11.07 7.315 11.475 7.645 ;
      RECT 11.07 6.475 11.475 6.805 ;
      RECT 11.14 3.555 11.33 3.78 ;
      RECT 11.13 3.556 11.335 3.775 ;
      RECT 11.13 3.558 11.345 3.755 ;
      RECT 11.13 3.562 11.35 3.74 ;
      RECT 11.13 3.549 11.3 3.775 ;
      RECT 11.13 3.552 11.325 3.775 ;
      RECT 11.14 3.548 11.3 3.78 ;
      RECT 11.226 3.546 11.3 3.78 ;
      RECT 10.85 2.797 11.02 3.035 ;
      RECT 10.85 2.797 11.106 2.949 ;
      RECT 10.85 2.797 11.11 2.859 ;
      RECT 10.9 2.57 11.12 2.838 ;
      RECT 10.895 2.587 11.125 2.811 ;
      RECT 10.86 2.745 11.125 2.811 ;
      RECT 10.88 2.595 11.02 3.035 ;
      RECT 10.87 2.677 11.13 2.794 ;
      RECT 10.865 2.725 11.13 2.794 ;
      RECT 10.87 2.635 11.125 2.811 ;
      RECT 10.895 2.572 11.12 2.838 ;
      RECT 10.46 2.547 10.63 2.745 ;
      RECT 10.46 2.547 10.675 2.72 ;
      RECT 10.53 2.49 10.7 2.678 ;
      RECT 10.505 2.505 10.7 2.678 ;
      RECT 10.12 2.551 10.15 2.745 ;
      RECT 10.115 2.523 10.12 2.745 ;
      RECT 10.085 2.497 10.115 2.747 ;
      RECT 10.06 2.455 10.085 2.75 ;
      RECT 10.05 2.427 10.06 2.752 ;
      RECT 10.015 2.407 10.05 2.754 ;
      RECT 9.95 2.392 10.015 2.76 ;
      RECT 9.9 2.39 9.95 2.766 ;
      RECT 9.877 2.392 9.9 2.771 ;
      RECT 9.791 2.403 9.877 2.777 ;
      RECT 9.705 2.421 9.791 2.787 ;
      RECT 9.69 2.432 9.705 2.793 ;
      RECT 9.62 2.455 9.69 2.799 ;
      RECT 9.565 2.487 9.62 2.807 ;
      RECT 9.525 2.51 9.565 2.813 ;
      RECT 9.511 2.523 9.525 2.816 ;
      RECT 9.425 2.545 9.511 2.822 ;
      RECT 9.41 2.57 9.425 2.828 ;
      RECT 9.37 2.585 9.41 2.832 ;
      RECT 9.32 2.6 9.37 2.837 ;
      RECT 9.295 2.607 9.32 2.841 ;
      RECT 9.235 2.602 9.295 2.845 ;
      RECT 9.22 2.593 9.235 2.849 ;
      RECT 9.15 2.583 9.22 2.845 ;
      RECT 9.125 2.575 9.145 2.835 ;
      RECT 9.066 2.575 9.125 2.813 ;
      RECT 8.98 2.575 9.066 2.77 ;
      RECT 9.145 2.575 9.15 2.84 ;
      RECT 9.84 1.806 10.01 2.14 ;
      RECT 9.81 1.806 10.01 2.135 ;
      RECT 9.75 1.773 9.81 2.123 ;
      RECT 9.75 1.829 10.02 2.118 ;
      RECT 9.725 1.829 10.02 2.112 ;
      RECT 9.72 1.77 9.75 2.109 ;
      RECT 9.705 1.776 9.84 2.107 ;
      RECT 9.7 1.784 9.925 2.095 ;
      RECT 9.7 1.836 10.035 2.048 ;
      RECT 9.685 1.792 9.925 2.043 ;
      RECT 9.685 1.862 10.045 1.984 ;
      RECT 9.655 1.812 10.01 1.945 ;
      RECT 9.655 1.902 10.055 1.941 ;
      RECT 9.705 1.781 9.925 2.107 ;
      RECT 9.045 2.111 9.1 2.375 ;
      RECT 9.045 2.111 9.165 2.374 ;
      RECT 9.045 2.111 9.19 2.373 ;
      RECT 9.045 2.111 9.255 2.372 ;
      RECT 9.19 2.077 9.27 2.371 ;
      RECT 9.005 2.121 9.415 2.37 ;
      RECT 9.045 2.118 9.415 2.37 ;
      RECT 9.005 2.126 9.42 2.363 ;
      RECT 8.99 2.128 9.42 2.362 ;
      RECT 8.99 2.135 9.425 2.358 ;
      RECT 8.97 2.134 9.42 2.354 ;
      RECT 8.97 2.142 9.43 2.353 ;
      RECT 8.965 2.139 9.425 2.349 ;
      RECT 8.965 2.152 9.44 2.348 ;
      RECT 8.95 2.142 9.43 2.347 ;
      RECT 8.915 2.155 9.44 2.34 ;
      RECT 9.1 2.11 9.41 2.37 ;
      RECT 9.1 2.095 9.36 2.37 ;
      RECT 9.165 2.082 9.295 2.37 ;
      RECT 8.71 3.171 8.725 3.564 ;
      RECT 8.675 3.176 8.725 3.563 ;
      RECT 8.71 3.175 8.77 3.562 ;
      RECT 8.655 3.186 8.77 3.561 ;
      RECT 8.67 3.182 8.77 3.561 ;
      RECT 8.635 3.192 8.845 3.558 ;
      RECT 8.635 3.211 8.89 3.556 ;
      RECT 8.635 3.218 8.895 3.553 ;
      RECT 8.62 3.195 8.845 3.55 ;
      RECT 8.6 3.2 8.845 3.543 ;
      RECT 8.595 3.204 8.845 3.539 ;
      RECT 8.595 3.221 8.905 3.538 ;
      RECT 8.575 3.215 8.89 3.534 ;
      RECT 8.575 3.224 8.91 3.528 ;
      RECT 8.57 3.23 8.91 3.3 ;
      RECT 8.635 3.19 8.77 3.558 ;
      RECT 8.51 2.553 8.71 2.865 ;
      RECT 8.585 2.531 8.71 2.865 ;
      RECT 8.525 2.55 8.715 2.85 ;
      RECT 8.495 2.561 8.715 2.848 ;
      RECT 8.51 2.556 8.72 2.814 ;
      RECT 8.495 2.66 8.725 2.781 ;
      RECT 8.525 2.532 8.71 2.865 ;
      RECT 8.585 2.51 8.685 2.865 ;
      RECT 8.61 2.507 8.685 2.865 ;
      RECT 8.61 2.502 8.63 2.865 ;
      RECT 8.015 2.57 8.19 2.745 ;
      RECT 8.01 2.57 8.19 2.743 ;
      RECT 7.985 2.57 8.19 2.738 ;
      RECT 7.93 2.55 8.1 2.728 ;
      RECT 7.93 2.557 8.165 2.728 ;
      RECT 8.015 3.237 8.03 3.42 ;
      RECT 8.005 3.215 8.015 3.42 ;
      RECT 7.99 3.195 8.005 3.42 ;
      RECT 7.98 3.17 7.99 3.42 ;
      RECT 7.95 3.135 7.98 3.42 ;
      RECT 7.915 3.075 7.95 3.42 ;
      RECT 7.91 3.037 7.915 3.42 ;
      RECT 7.86 2.988 7.91 3.42 ;
      RECT 7.85 2.938 7.86 3.408 ;
      RECT 7.835 2.917 7.85 3.368 ;
      RECT 7.815 2.885 7.835 3.318 ;
      RECT 7.79 2.841 7.815 3.258 ;
      RECT 7.785 2.813 7.79 3.213 ;
      RECT 7.78 2.804 7.785 3.199 ;
      RECT 7.775 2.797 7.78 3.186 ;
      RECT 7.77 2.792 7.775 3.175 ;
      RECT 7.765 2.777 7.77 3.165 ;
      RECT 7.76 2.755 7.765 3.152 ;
      RECT 7.75 2.715 7.76 3.127 ;
      RECT 7.725 2.645 7.75 3.083 ;
      RECT 7.72 2.585 7.725 3.048 ;
      RECT 7.705 2.565 7.72 3.015 ;
      RECT 7.7 2.565 7.705 2.99 ;
      RECT 7.67 2.565 7.7 2.945 ;
      RECT 7.625 2.565 7.67 2.885 ;
      RECT 7.55 2.565 7.625 2.833 ;
      RECT 7.545 2.565 7.55 2.798 ;
      RECT 7.54 2.565 7.545 2.788 ;
      RECT 7.535 2.565 7.54 2.768 ;
      RECT 7.8 1.785 7.97 2.255 ;
      RECT 7.745 1.778 7.94 2.239 ;
      RECT 7.745 1.792 7.975 2.238 ;
      RECT 7.73 1.793 7.975 2.219 ;
      RECT 7.725 1.811 7.975 2.205 ;
      RECT 7.73 1.794 7.98 2.203 ;
      RECT 7.715 1.825 7.98 2.188 ;
      RECT 7.73 1.8 7.985 2.173 ;
      RECT 7.71 1.84 7.985 2.17 ;
      RECT 7.725 1.812 7.99 2.155 ;
      RECT 7.725 1.824 7.995 2.135 ;
      RECT 7.71 1.84 8 2.118 ;
      RECT 7.71 1.85 8.005 1.973 ;
      RECT 7.705 1.85 8.005 1.93 ;
      RECT 7.705 1.865 8.01 1.908 ;
      RECT 7.8 1.775 7.94 2.255 ;
      RECT 7.8 1.773 7.91 2.255 ;
      RECT 7.886 1.77 7.91 2.255 ;
      RECT 7.545 3.437 7.55 3.483 ;
      RECT 7.535 3.285 7.545 3.507 ;
      RECT 7.53 3.13 7.535 3.532 ;
      RECT 7.515 3.092 7.53 3.543 ;
      RECT 7.51 3.075 7.515 3.55 ;
      RECT 7.5 3.063 7.51 3.557 ;
      RECT 7.495 3.054 7.5 3.559 ;
      RECT 7.49 3.052 7.495 3.563 ;
      RECT 7.445 3.043 7.49 3.578 ;
      RECT 7.44 3.035 7.445 3.592 ;
      RECT 7.435 3.032 7.44 3.596 ;
      RECT 7.42 3.027 7.435 3.604 ;
      RECT 7.365 3.017 7.42 3.615 ;
      RECT 7.33 3.005 7.365 3.616 ;
      RECT 7.321 3 7.33 3.61 ;
      RECT 7.235 3 7.321 3.6 ;
      RECT 7.205 3 7.235 3.578 ;
      RECT 7.195 3 7.2 3.558 ;
      RECT 7.19 3 7.195 3.52 ;
      RECT 7.185 3 7.19 3.478 ;
      RECT 7.18 3 7.185 3.438 ;
      RECT 7.175 3 7.18 3.368 ;
      RECT 7.165 3 7.175 3.29 ;
      RECT 7.16 3 7.165 3.19 ;
      RECT 7.2 3 7.205 3.56 ;
      RECT 6.695 3.082 6.785 3.56 ;
      RECT 6.68 3.085 6.8 3.558 ;
      RECT 6.695 3.084 6.8 3.558 ;
      RECT 6.66 3.091 6.825 3.548 ;
      RECT 6.68 3.085 6.825 3.548 ;
      RECT 6.645 3.097 6.825 3.536 ;
      RECT 6.68 3.088 6.875 3.529 ;
      RECT 6.631 3.105 6.875 3.527 ;
      RECT 6.66 3.095 6.885 3.515 ;
      RECT 6.631 3.116 6.915 3.506 ;
      RECT 6.545 3.14 6.915 3.5 ;
      RECT 6.545 3.153 6.955 3.483 ;
      RECT 6.54 3.175 6.955 3.476 ;
      RECT 6.51 3.19 6.955 3.466 ;
      RECT 6.505 3.201 6.955 3.456 ;
      RECT 6.475 3.214 6.955 3.447 ;
      RECT 6.46 3.232 6.955 3.436 ;
      RECT 6.435 3.245 6.955 3.426 ;
      RECT 6.695 3.081 6.705 3.56 ;
      RECT 6.741 2.505 6.78 2.75 ;
      RECT 6.655 2.505 6.79 2.748 ;
      RECT 6.54 2.53 6.79 2.745 ;
      RECT 6.54 2.53 6.795 2.743 ;
      RECT 6.54 2.53 6.81 2.738 ;
      RECT 6.646 2.505 6.825 2.718 ;
      RECT 6.56 2.513 6.825 2.718 ;
      RECT 6.23 1.865 6.4 2.3 ;
      RECT 6.22 1.899 6.4 2.283 ;
      RECT 6.3 1.835 6.47 2.27 ;
      RECT 6.205 1.91 6.47 2.248 ;
      RECT 6.3 1.845 6.475 2.238 ;
      RECT 6.23 1.897 6.505 2.223 ;
      RECT 6.19 1.923 6.505 2.208 ;
      RECT 6.19 1.965 6.515 2.188 ;
      RECT 6.185 1.99 6.52 2.17 ;
      RECT 6.185 2 6.525 2.155 ;
      RECT 6.18 1.937 6.505 2.153 ;
      RECT 6.18 2.01 6.53 2.138 ;
      RECT 6.175 1.947 6.505 2.135 ;
      RECT 6.17 2.031 6.535 2.118 ;
      RECT 6.17 2.063 6.54 2.098 ;
      RECT 6.165 1.977 6.515 2.09 ;
      RECT 6.17 1.962 6.505 2.118 ;
      RECT 6.185 1.932 6.505 2.17 ;
      RECT 6.03 2.519 6.255 2.775 ;
      RECT 6.03 2.552 6.275 2.765 ;
      RECT 5.995 2.552 6.275 2.763 ;
      RECT 5.995 2.565 6.28 2.753 ;
      RECT 5.995 2.585 6.29 2.745 ;
      RECT 5.995 2.682 6.295 2.738 ;
      RECT 5.975 2.43 6.105 2.728 ;
      RECT 5.93 2.585 6.29 2.67 ;
      RECT 5.92 2.43 6.105 2.615 ;
      RECT 5.92 2.462 6.191 2.615 ;
      RECT 5.885 2.992 5.905 3.17 ;
      RECT 5.85 2.945 5.885 3.17 ;
      RECT 5.835 2.885 5.85 3.17 ;
      RECT 5.81 2.832 5.835 3.17 ;
      RECT 5.795 2.785 5.81 3.17 ;
      RECT 5.775 2.762 5.795 3.17 ;
      RECT 5.75 2.727 5.775 3.17 ;
      RECT 5.74 2.573 5.75 3.17 ;
      RECT 5.71 2.568 5.74 3.161 ;
      RECT 5.705 2.565 5.71 3.151 ;
      RECT 5.69 2.565 5.705 3.125 ;
      RECT 5.685 2.565 5.69 3.088 ;
      RECT 5.66 2.565 5.685 3.04 ;
      RECT 5.64 2.565 5.66 2.965 ;
      RECT 5.63 2.565 5.64 2.925 ;
      RECT 5.625 2.565 5.63 2.9 ;
      RECT 5.62 2.565 5.625 2.883 ;
      RECT 5.615 2.565 5.62 2.865 ;
      RECT 5.61 2.566 5.615 2.855 ;
      RECT 5.6 2.568 5.61 2.823 ;
      RECT 5.59 2.57 5.6 2.79 ;
      RECT 5.58 2.573 5.59 2.763 ;
      RECT 5.905 3 6.13 3.17 ;
      RECT 5.235 1.812 5.405 2.265 ;
      RECT 5.235 1.812 5.495 2.231 ;
      RECT 5.235 1.812 5.525 2.215 ;
      RECT 5.235 1.812 5.555 2.188 ;
      RECT 5.491 1.79 5.57 2.17 ;
      RECT 5.27 1.797 5.575 2.155 ;
      RECT 5.27 1.805 5.585 2.118 ;
      RECT 5.23 1.832 5.585 2.09 ;
      RECT 5.215 1.845 5.585 2.055 ;
      RECT 5.235 1.82 5.605 2.045 ;
      RECT 5.21 1.885 5.605 2.015 ;
      RECT 5.21 1.915 5.61 1.998 ;
      RECT 5.205 1.945 5.61 1.985 ;
      RECT 5.27 1.794 5.57 2.17 ;
      RECT 5.405 1.791 5.491 2.249 ;
      RECT 5.356 1.792 5.57 2.17 ;
      RECT 5.5 3.452 5.545 3.645 ;
      RECT 5.49 3.422 5.5 3.645 ;
      RECT 5.485 3.407 5.49 3.645 ;
      RECT 5.445 3.317 5.485 3.645 ;
      RECT 5.44 3.23 5.445 3.645 ;
      RECT 5.43 3.2 5.44 3.645 ;
      RECT 5.425 3.16 5.43 3.645 ;
      RECT 5.415 3.122 5.425 3.645 ;
      RECT 5.41 3.087 5.415 3.645 ;
      RECT 5.39 3.04 5.41 3.645 ;
      RECT 5.375 2.965 5.39 3.645 ;
      RECT 5.37 2.92 5.375 3.64 ;
      RECT 5.365 2.9 5.37 3.613 ;
      RECT 5.36 2.88 5.365 3.598 ;
      RECT 5.355 2.855 5.36 3.578 ;
      RECT 5.35 2.833 5.355 3.563 ;
      RECT 5.345 2.811 5.35 3.545 ;
      RECT 5.34 2.79 5.345 3.535 ;
      RECT 5.33 2.762 5.34 3.505 ;
      RECT 5.32 2.725 5.33 3.473 ;
      RECT 5.31 2.685 5.32 3.44 ;
      RECT 5.3 2.663 5.31 3.41 ;
      RECT 5.27 2.615 5.3 3.342 ;
      RECT 5.255 2.575 5.27 3.269 ;
      RECT 5.245 2.575 5.255 3.235 ;
      RECT 5.24 2.575 5.245 3.21 ;
      RECT 5.235 2.575 5.24 3.195 ;
      RECT 5.23 2.575 5.235 3.173 ;
      RECT 5.225 2.575 5.23 3.16 ;
      RECT 5.21 2.575 5.225 3.125 ;
      RECT 5.19 2.575 5.21 3.065 ;
      RECT 5.18 2.575 5.19 3.015 ;
      RECT 5.16 2.575 5.18 2.963 ;
      RECT 5.14 2.575 5.16 2.92 ;
      RECT 5.13 2.575 5.14 2.908 ;
      RECT 5.1 2.575 5.13 2.895 ;
      RECT 5.07 2.596 5.1 2.875 ;
      RECT 5.06 2.624 5.07 2.855 ;
      RECT 5.045 2.641 5.06 2.823 ;
      RECT 5.04 2.655 5.045 2.79 ;
      RECT 5.035 2.663 5.04 2.763 ;
      RECT 5.03 2.671 5.035 2.725 ;
      RECT 5.035 3.195 5.04 3.53 ;
      RECT 5 3.182 5.035 3.529 ;
      RECT 4.93 3.122 5 3.528 ;
      RECT 4.85 3.065 4.93 3.527 ;
      RECT 4.715 3.025 4.85 3.526 ;
      RECT 4.715 3.212 5.05 3.515 ;
      RECT 4.675 3.212 5.05 3.505 ;
      RECT 4.675 3.23 5.055 3.5 ;
      RECT 4.675 3.32 5.06 3.49 ;
      RECT 4.67 3.015 4.835 3.47 ;
      RECT 4.665 3.015 4.835 3.213 ;
      RECT 4.665 3.172 5.03 3.213 ;
      RECT 4.665 3.16 5.025 3.213 ;
      RECT 2.655 7.855 2.825 8.305 ;
      RECT 2.71 6.075 2.88 8.025 ;
      RECT 2.655 5.015 2.825 6.245 ;
      RECT 2.135 5.015 2.305 8.305 ;
      RECT 2.135 7.315 2.54 7.645 ;
      RECT 2.135 6.475 2.54 6.805 ;
      RECT 82.705 7.8 82.875 8.31 ;
      RECT 81.715 0.57 81.885 1.08 ;
      RECT 81.715 2.39 81.885 3.86 ;
      RECT 81.715 5.02 81.885 6.49 ;
      RECT 81.715 7.8 81.885 8.31 ;
      RECT 80.355 0.575 80.525 3.865 ;
      RECT 80.355 5.015 80.525 8.305 ;
      RECT 79.925 0.575 80.095 1.085 ;
      RECT 79.925 1.655 80.095 3.865 ;
      RECT 79.925 5.015 80.095 7.225 ;
      RECT 79.925 7.795 80.095 8.305 ;
      RECT 77.535 2.85 77.905 3.22 ;
      RECT 75.575 5.015 75.745 8.305 ;
      RECT 75.145 5.015 75.315 7.225 ;
      RECT 75.145 7.795 75.315 8.305 ;
      RECT 66.92 7.8 67.09 8.31 ;
      RECT 65.93 0.57 66.1 1.08 ;
      RECT 65.93 2.39 66.1 3.86 ;
      RECT 65.93 5.02 66.1 6.49 ;
      RECT 65.93 7.8 66.1 8.31 ;
      RECT 64.57 0.575 64.74 3.865 ;
      RECT 64.57 5.015 64.74 8.305 ;
      RECT 64.14 0.575 64.31 1.085 ;
      RECT 64.14 1.655 64.31 3.865 ;
      RECT 64.14 5.015 64.31 7.225 ;
      RECT 64.14 7.795 64.31 8.305 ;
      RECT 61.75 2.85 62.12 3.22 ;
      RECT 59.79 5.015 59.96 8.305 ;
      RECT 59.36 5.015 59.53 7.225 ;
      RECT 59.36 7.795 59.53 8.305 ;
      RECT 51.135 7.8 51.305 8.31 ;
      RECT 50.145 0.57 50.315 1.08 ;
      RECT 50.145 2.39 50.315 3.86 ;
      RECT 50.145 5.02 50.315 6.49 ;
      RECT 50.145 7.8 50.315 8.31 ;
      RECT 48.785 0.575 48.955 3.865 ;
      RECT 48.785 5.015 48.955 8.305 ;
      RECT 48.355 0.575 48.525 1.085 ;
      RECT 48.355 1.655 48.525 3.865 ;
      RECT 48.355 5.015 48.525 7.225 ;
      RECT 48.355 7.795 48.525 8.305 ;
      RECT 45.965 2.85 46.335 3.22 ;
      RECT 44.005 5.015 44.175 8.305 ;
      RECT 43.575 5.015 43.745 7.225 ;
      RECT 43.575 7.795 43.745 8.305 ;
      RECT 35.36 7.8 35.53 8.31 ;
      RECT 34.37 0.57 34.54 1.08 ;
      RECT 34.37 2.39 34.54 3.86 ;
      RECT 34.37 5.02 34.54 6.49 ;
      RECT 34.37 7.8 34.54 8.31 ;
      RECT 33.01 0.575 33.18 3.865 ;
      RECT 33.01 5.015 33.18 8.305 ;
      RECT 32.58 0.575 32.75 1.085 ;
      RECT 32.58 1.655 32.75 3.865 ;
      RECT 32.58 5.015 32.75 7.225 ;
      RECT 32.58 7.795 32.75 8.305 ;
      RECT 30.19 2.85 30.56 3.22 ;
      RECT 28.23 5.015 28.4 8.305 ;
      RECT 27.8 5.015 27.97 7.225 ;
      RECT 27.8 7.795 27.97 8.305 ;
      RECT 19.58 7.8 19.75 8.31 ;
      RECT 18.59 0.57 18.76 1.08 ;
      RECT 18.59 2.39 18.76 3.86 ;
      RECT 18.59 5.02 18.76 6.49 ;
      RECT 18.59 7.8 18.76 8.31 ;
      RECT 17.23 0.575 17.4 3.865 ;
      RECT 17.23 5.015 17.4 8.305 ;
      RECT 16.8 0.575 16.97 1.085 ;
      RECT 16.8 1.655 16.97 3.865 ;
      RECT 16.8 5.015 16.97 7.225 ;
      RECT 16.8 7.795 16.97 8.305 ;
      RECT 14.41 2.85 14.78 3.22 ;
      RECT 12.45 5.015 12.62 8.305 ;
      RECT 12.02 5.015 12.19 7.225 ;
      RECT 12.02 7.795 12.19 8.305 ;
      RECT 3.085 5.015 3.255 7.225 ;
      RECT 3.085 7.795 3.255 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2aa_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2at_8_b0r1
  CLASS BLOCK ;
  ORIGIN -1.46 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2at_8_b0r1 ;
  SIZE 92.435 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 21.655 0.915 21.825 1.085 ;
        RECT 21.65 0.91 21.82 1.08 ;
        RECT 21.65 2.39 21.82 2.56 ;
      LAYER li1 ;
        RECT 21.655 0.915 21.825 1.085 ;
        RECT 21.65 0.57 21.82 1.08 ;
        RECT 21.65 2.39 21.82 3.86 ;
      LAYER met1 ;
        RECT 21.59 2.36 21.88 2.59 ;
        RECT 21.59 0.88 21.88 1.11 ;
        RECT 21.65 0.88 21.82 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 39.58 0.915 39.75 1.085 ;
        RECT 39.575 0.91 39.745 1.08 ;
        RECT 39.575 2.39 39.745 2.56 ;
      LAYER li1 ;
        RECT 39.58 0.915 39.75 1.085 ;
        RECT 39.575 0.57 39.745 1.08 ;
        RECT 39.575 2.39 39.745 3.86 ;
      LAYER met1 ;
        RECT 39.515 2.36 39.805 2.59 ;
        RECT 39.515 0.88 39.805 1.11 ;
        RECT 39.575 0.88 39.745 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 57.505 0.915 57.675 1.085 ;
        RECT 57.5 0.91 57.67 1.08 ;
        RECT 57.5 2.39 57.67 2.56 ;
      LAYER li1 ;
        RECT 57.505 0.915 57.675 1.085 ;
        RECT 57.5 0.57 57.67 1.08 ;
        RECT 57.5 2.39 57.67 3.86 ;
      LAYER met1 ;
        RECT 57.44 2.36 57.73 2.59 ;
        RECT 57.44 0.88 57.73 1.11 ;
        RECT 57.5 0.88 57.67 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 75.43 0.915 75.6 1.085 ;
        RECT 75.425 0.91 75.595 1.08 ;
        RECT 75.425 2.39 75.595 2.56 ;
      LAYER li1 ;
        RECT 75.43 0.915 75.6 1.085 ;
        RECT 75.425 0.57 75.595 1.08 ;
        RECT 75.425 2.39 75.595 3.86 ;
      LAYER met1 ;
        RECT 75.365 2.36 75.655 2.59 ;
        RECT 75.365 0.88 75.655 1.11 ;
        RECT 75.425 0.88 75.595 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 93.355 0.915 93.525 1.085 ;
        RECT 93.35 0.91 93.52 1.08 ;
        RECT 93.35 2.39 93.52 2.56 ;
      LAYER li1 ;
        RECT 93.355 0.915 93.525 1.085 ;
        RECT 93.35 0.57 93.52 1.08 ;
        RECT 93.35 2.39 93.52 3.86 ;
      LAYER met1 ;
        RECT 93.29 2.36 93.58 2.59 ;
        RECT 93.29 0.88 93.58 1.11 ;
        RECT 93.35 0.88 93.52 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 17.5 1.66 17.67 2.935 ;
        RECT 17.5 5.945 17.67 7.22 ;
        RECT 12.74 5.945 12.91 7.22 ;
      LAYER met2 ;
        RECT 17.42 2.705 17.77 3.055 ;
        RECT 17.41 5.84 17.76 6.19 ;
        RECT 17.485 2.705 17.66 6.19 ;
      LAYER met1 ;
        RECT 17.42 2.765 17.9 2.935 ;
        RECT 17.42 2.705 17.77 3.055 ;
        RECT 12.68 5.945 17.9 6.115 ;
        RECT 17.41 5.84 17.76 6.19 ;
        RECT 12.68 5.915 12.97 6.145 ;
      LAYER via1 ;
        RECT 17.51 5.94 17.66 6.09 ;
        RECT 17.52 2.805 17.67 2.955 ;
      LAYER mcon ;
        RECT 12.74 5.945 12.91 6.115 ;
        RECT 17.5 5.945 17.67 6.115 ;
        RECT 17.5 2.765 17.67 2.935 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 35.425 1.66 35.595 2.935 ;
        RECT 35.425 5.945 35.595 7.22 ;
        RECT 30.665 5.945 30.835 7.22 ;
      LAYER met2 ;
        RECT 35.345 2.705 35.695 3.055 ;
        RECT 35.335 5.84 35.685 6.19 ;
        RECT 35.41 2.705 35.585 6.19 ;
      LAYER met1 ;
        RECT 35.345 2.765 35.825 2.935 ;
        RECT 35.345 2.705 35.695 3.055 ;
        RECT 30.605 5.945 35.825 6.115 ;
        RECT 35.335 5.84 35.685 6.19 ;
        RECT 30.605 5.915 30.895 6.145 ;
      LAYER via1 ;
        RECT 35.435 5.94 35.585 6.09 ;
        RECT 35.445 2.805 35.595 2.955 ;
      LAYER mcon ;
        RECT 30.665 5.945 30.835 6.115 ;
        RECT 35.425 5.945 35.595 6.115 ;
        RECT 35.425 2.765 35.595 2.935 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 53.35 1.66 53.52 2.935 ;
        RECT 53.35 5.945 53.52 7.22 ;
        RECT 48.59 5.945 48.76 7.22 ;
      LAYER met2 ;
        RECT 53.27 2.705 53.62 3.055 ;
        RECT 53.26 5.84 53.61 6.19 ;
        RECT 53.335 2.705 53.51 6.19 ;
      LAYER met1 ;
        RECT 53.27 2.765 53.75 2.935 ;
        RECT 53.27 2.705 53.62 3.055 ;
        RECT 48.53 5.945 53.75 6.115 ;
        RECT 53.26 5.84 53.61 6.19 ;
        RECT 48.53 5.915 48.82 6.145 ;
      LAYER via1 ;
        RECT 53.36 5.94 53.51 6.09 ;
        RECT 53.37 2.805 53.52 2.955 ;
      LAYER mcon ;
        RECT 48.59 5.945 48.76 6.115 ;
        RECT 53.35 5.945 53.52 6.115 ;
        RECT 53.35 2.765 53.52 2.935 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 71.275 1.66 71.445 2.935 ;
        RECT 71.275 5.945 71.445 7.22 ;
        RECT 66.515 5.945 66.685 7.22 ;
      LAYER met2 ;
        RECT 71.195 2.705 71.545 3.055 ;
        RECT 71.185 5.84 71.535 6.19 ;
        RECT 71.26 2.705 71.435 6.19 ;
      LAYER met1 ;
        RECT 71.195 2.765 71.675 2.935 ;
        RECT 71.195 2.705 71.545 3.055 ;
        RECT 66.455 5.945 71.675 6.115 ;
        RECT 71.185 5.84 71.535 6.19 ;
        RECT 66.455 5.915 66.745 6.145 ;
      LAYER via1 ;
        RECT 71.285 5.94 71.435 6.09 ;
        RECT 71.295 2.805 71.445 2.955 ;
      LAYER mcon ;
        RECT 66.515 5.945 66.685 6.115 ;
        RECT 71.275 5.945 71.445 6.115 ;
        RECT 71.275 2.765 71.445 2.935 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 89.2 1.66 89.37 2.935 ;
        RECT 89.2 5.945 89.37 7.22 ;
        RECT 84.44 5.945 84.61 7.22 ;
      LAYER met2 ;
        RECT 89.12 2.705 89.47 3.055 ;
        RECT 89.11 5.84 89.46 6.19 ;
        RECT 89.185 2.705 89.36 6.19 ;
      LAYER met1 ;
        RECT 89.12 2.765 89.6 2.935 ;
        RECT 89.12 2.705 89.47 3.055 ;
        RECT 84.38 5.945 89.6 6.115 ;
        RECT 89.11 5.84 89.46 6.19 ;
        RECT 84.38 5.915 84.67 6.145 ;
      LAYER via1 ;
        RECT 89.21 5.94 89.36 6.09 ;
        RECT 89.22 2.805 89.37 2.955 ;
      LAYER mcon ;
        RECT 84.44 5.945 84.61 6.115 ;
        RECT 89.2 5.945 89.37 6.115 ;
        RECT 89.2 2.765 89.37 2.935 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 1.71 5.945 1.88 7.22 ;
      LAYER met1 ;
        RECT 1.65 5.945 2.11 6.115 ;
        RECT 1.65 5.915 1.94 6.145 ;
      LAYER mcon ;
        RECT 1.71 5.945 1.88 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.48 4.285 93.895 4.745 ;
        RECT 87.935 4.135 93.895 4.745 ;
        RECT 91.76 4.13 93.74 4.75 ;
        RECT 92.92 3.4 93.09 5.48 ;
        RECT 91.93 3.4 92.1 5.48 ;
        RECT 89.19 3.405 89.36 5.475 ;
        RECT 86.435 3.785 86.605 4.745 ;
        RECT 84.43 4.285 84.6 5.475 ;
        RECT 83.995 3.785 84.165 4.745 ;
        RECT 82.035 3.785 82.205 4.745 ;
        RECT 81.075 3.785 81.245 4.745 ;
        RECT 79.115 3.785 79.285 4.745 ;
        RECT 78.115 3.785 78.285 4.745 ;
        RECT 77.155 3.785 77.325 4.745 ;
        RECT 70.01 4.135 75.97 4.745 ;
        RECT 73.835 4.13 75.815 4.75 ;
        RECT 74.995 3.4 75.165 5.48 ;
        RECT 74.005 3.4 74.175 5.48 ;
        RECT 71.265 3.405 71.435 5.475 ;
        RECT 68.51 3.785 68.68 4.745 ;
        RECT 66.505 4.285 66.675 5.475 ;
        RECT 66.07 3.785 66.24 4.745 ;
        RECT 64.11 3.785 64.28 4.745 ;
        RECT 63.15 3.785 63.32 4.745 ;
        RECT 61.19 3.785 61.36 4.745 ;
        RECT 60.19 3.785 60.36 4.745 ;
        RECT 59.23 3.785 59.4 4.745 ;
        RECT 52.085 4.135 58.045 4.745 ;
        RECT 55.91 4.13 57.89 4.75 ;
        RECT 57.07 3.4 57.24 5.48 ;
        RECT 56.08 3.4 56.25 5.48 ;
        RECT 53.34 3.405 53.51 5.475 ;
        RECT 50.585 3.785 50.755 4.745 ;
        RECT 48.58 4.285 48.75 5.475 ;
        RECT 48.145 3.785 48.315 4.745 ;
        RECT 46.185 3.785 46.355 4.745 ;
        RECT 45.225 3.785 45.395 4.745 ;
        RECT 43.265 3.785 43.435 4.745 ;
        RECT 42.265 3.785 42.435 4.745 ;
        RECT 41.305 3.785 41.475 4.745 ;
        RECT 34.16 4.135 40.12 4.745 ;
        RECT 37.985 4.13 39.965 4.75 ;
        RECT 39.145 3.4 39.315 5.48 ;
        RECT 38.155 3.4 38.325 5.48 ;
        RECT 35.415 3.405 35.585 5.475 ;
        RECT 32.66 3.785 32.83 4.745 ;
        RECT 30.655 4.285 30.825 5.475 ;
        RECT 30.22 3.785 30.39 4.745 ;
        RECT 28.26 3.785 28.43 4.745 ;
        RECT 27.3 3.785 27.47 4.745 ;
        RECT 25.34 3.785 25.51 4.745 ;
        RECT 24.34 3.785 24.51 4.745 ;
        RECT 23.38 3.785 23.55 4.745 ;
        RECT 16.235 4.135 22.195 4.745 ;
        RECT 20.06 4.13 22.04 4.75 ;
        RECT 21.22 3.4 21.39 5.48 ;
        RECT 20.23 3.4 20.4 5.48 ;
        RECT 17.49 3.405 17.66 5.475 ;
        RECT 14.735 3.785 14.905 4.745 ;
        RECT 12.73 4.285 12.9 5.475 ;
        RECT 12.295 3.785 12.465 4.745 ;
        RECT 10.335 3.785 10.505 4.745 ;
        RECT 9.375 3.785 9.545 4.745 ;
        RECT 7.415 3.785 7.585 4.745 ;
        RECT 6.415 3.785 6.585 4.745 ;
        RECT 5.455 3.785 5.625 4.745 ;
        RECT 3.51 4.285 3.68 8.305 ;
        RECT 1.7 4.285 1.87 5.475 ;
      LAYER met1 ;
        RECT 1.48 4.285 93.895 4.745 ;
        RECT 76.345 4.135 93.895 4.745 ;
        RECT 91.76 4.13 93.74 4.75 ;
        RECT 76.345 4.13 88.305 4.745 ;
        RECT 58.42 4.135 75.97 4.745 ;
        RECT 73.835 4.13 75.815 4.75 ;
        RECT 58.42 4.13 70.38 4.745 ;
        RECT 40.495 4.135 58.045 4.745 ;
        RECT 55.91 4.13 57.89 4.75 ;
        RECT 40.495 4.13 52.455 4.745 ;
        RECT 22.57 4.135 40.12 4.745 ;
        RECT 37.985 4.13 39.965 4.75 ;
        RECT 22.57 4.13 34.53 4.745 ;
        RECT 4.645 4.135 22.195 4.745 ;
        RECT 20.06 4.13 22.04 4.75 ;
        RECT 4.645 4.13 16.605 4.745 ;
        RECT 3.45 6.655 3.74 6.885 ;
        RECT 3.28 6.685 3.74 6.855 ;
      LAYER mcon ;
        RECT 3.51 6.685 3.68 6.855 ;
        RECT 3.82 4.545 3.99 4.715 ;
        RECT 4.79 4.285 4.96 4.455 ;
        RECT 5.25 4.285 5.42 4.455 ;
        RECT 5.71 4.285 5.88 4.455 ;
        RECT 6.17 4.285 6.34 4.455 ;
        RECT 6.63 4.285 6.8 4.455 ;
        RECT 7.09 4.285 7.26 4.455 ;
        RECT 7.55 4.285 7.72 4.455 ;
        RECT 8.01 4.285 8.18 4.455 ;
        RECT 8.47 4.285 8.64 4.455 ;
        RECT 8.93 4.285 9.1 4.455 ;
        RECT 9.39 4.285 9.56 4.455 ;
        RECT 9.85 4.285 10.02 4.455 ;
        RECT 10.31 4.285 10.48 4.455 ;
        RECT 10.77 4.285 10.94 4.455 ;
        RECT 11.23 4.285 11.4 4.455 ;
        RECT 11.69 4.285 11.86 4.455 ;
        RECT 12.15 4.285 12.32 4.455 ;
        RECT 12.61 4.285 12.78 4.455 ;
        RECT 13.07 4.285 13.24 4.455 ;
        RECT 13.53 4.285 13.7 4.455 ;
        RECT 13.99 4.285 14.16 4.455 ;
        RECT 14.45 4.285 14.62 4.455 ;
        RECT 14.85 4.545 15.02 4.715 ;
        RECT 14.91 4.285 15.08 4.455 ;
        RECT 15.37 4.285 15.54 4.455 ;
        RECT 15.83 4.285 16 4.455 ;
        RECT 16.29 4.285 16.46 4.455 ;
        RECT 19.61 4.545 19.78 4.715 ;
        RECT 19.61 4.165 19.78 4.335 ;
        RECT 20.31 4.55 20.48 4.72 ;
        RECT 20.31 4.16 20.48 4.33 ;
        RECT 21.3 4.55 21.47 4.72 ;
        RECT 21.3 4.16 21.47 4.33 ;
        RECT 22.715 4.285 22.885 4.455 ;
        RECT 23.175 4.285 23.345 4.455 ;
        RECT 23.635 4.285 23.805 4.455 ;
        RECT 24.095 4.285 24.265 4.455 ;
        RECT 24.555 4.285 24.725 4.455 ;
        RECT 25.015 4.285 25.185 4.455 ;
        RECT 25.475 4.285 25.645 4.455 ;
        RECT 25.935 4.285 26.105 4.455 ;
        RECT 26.395 4.285 26.565 4.455 ;
        RECT 26.855 4.285 27.025 4.455 ;
        RECT 27.315 4.285 27.485 4.455 ;
        RECT 27.775 4.285 27.945 4.455 ;
        RECT 28.235 4.285 28.405 4.455 ;
        RECT 28.695 4.285 28.865 4.455 ;
        RECT 29.155 4.285 29.325 4.455 ;
        RECT 29.615 4.285 29.785 4.455 ;
        RECT 30.075 4.285 30.245 4.455 ;
        RECT 30.535 4.285 30.705 4.455 ;
        RECT 30.995 4.285 31.165 4.455 ;
        RECT 31.455 4.285 31.625 4.455 ;
        RECT 31.915 4.285 32.085 4.455 ;
        RECT 32.375 4.285 32.545 4.455 ;
        RECT 32.775 4.545 32.945 4.715 ;
        RECT 32.835 4.285 33.005 4.455 ;
        RECT 33.295 4.285 33.465 4.455 ;
        RECT 33.755 4.285 33.925 4.455 ;
        RECT 34.215 4.285 34.385 4.455 ;
        RECT 37.535 4.545 37.705 4.715 ;
        RECT 37.535 4.165 37.705 4.335 ;
        RECT 38.235 4.55 38.405 4.72 ;
        RECT 38.235 4.16 38.405 4.33 ;
        RECT 39.225 4.55 39.395 4.72 ;
        RECT 39.225 4.16 39.395 4.33 ;
        RECT 40.64 4.285 40.81 4.455 ;
        RECT 41.1 4.285 41.27 4.455 ;
        RECT 41.56 4.285 41.73 4.455 ;
        RECT 42.02 4.285 42.19 4.455 ;
        RECT 42.48 4.285 42.65 4.455 ;
        RECT 42.94 4.285 43.11 4.455 ;
        RECT 43.4 4.285 43.57 4.455 ;
        RECT 43.86 4.285 44.03 4.455 ;
        RECT 44.32 4.285 44.49 4.455 ;
        RECT 44.78 4.285 44.95 4.455 ;
        RECT 45.24 4.285 45.41 4.455 ;
        RECT 45.7 4.285 45.87 4.455 ;
        RECT 46.16 4.285 46.33 4.455 ;
        RECT 46.62 4.285 46.79 4.455 ;
        RECT 47.08 4.285 47.25 4.455 ;
        RECT 47.54 4.285 47.71 4.455 ;
        RECT 48 4.285 48.17 4.455 ;
        RECT 48.46 4.285 48.63 4.455 ;
        RECT 48.92 4.285 49.09 4.455 ;
        RECT 49.38 4.285 49.55 4.455 ;
        RECT 49.84 4.285 50.01 4.455 ;
        RECT 50.3 4.285 50.47 4.455 ;
        RECT 50.7 4.545 50.87 4.715 ;
        RECT 50.76 4.285 50.93 4.455 ;
        RECT 51.22 4.285 51.39 4.455 ;
        RECT 51.68 4.285 51.85 4.455 ;
        RECT 52.14 4.285 52.31 4.455 ;
        RECT 55.46 4.545 55.63 4.715 ;
        RECT 55.46 4.165 55.63 4.335 ;
        RECT 56.16 4.55 56.33 4.72 ;
        RECT 56.16 4.16 56.33 4.33 ;
        RECT 57.15 4.55 57.32 4.72 ;
        RECT 57.15 4.16 57.32 4.33 ;
        RECT 58.565 4.285 58.735 4.455 ;
        RECT 59.025 4.285 59.195 4.455 ;
        RECT 59.485 4.285 59.655 4.455 ;
        RECT 59.945 4.285 60.115 4.455 ;
        RECT 60.405 4.285 60.575 4.455 ;
        RECT 60.865 4.285 61.035 4.455 ;
        RECT 61.325 4.285 61.495 4.455 ;
        RECT 61.785 4.285 61.955 4.455 ;
        RECT 62.245 4.285 62.415 4.455 ;
        RECT 62.705 4.285 62.875 4.455 ;
        RECT 63.165 4.285 63.335 4.455 ;
        RECT 63.625 4.285 63.795 4.455 ;
        RECT 64.085 4.285 64.255 4.455 ;
        RECT 64.545 4.285 64.715 4.455 ;
        RECT 65.005 4.285 65.175 4.455 ;
        RECT 65.465 4.285 65.635 4.455 ;
        RECT 65.925 4.285 66.095 4.455 ;
        RECT 66.385 4.285 66.555 4.455 ;
        RECT 66.845 4.285 67.015 4.455 ;
        RECT 67.305 4.285 67.475 4.455 ;
        RECT 67.765 4.285 67.935 4.455 ;
        RECT 68.225 4.285 68.395 4.455 ;
        RECT 68.625 4.545 68.795 4.715 ;
        RECT 68.685 4.285 68.855 4.455 ;
        RECT 69.145 4.285 69.315 4.455 ;
        RECT 69.605 4.285 69.775 4.455 ;
        RECT 70.065 4.285 70.235 4.455 ;
        RECT 73.385 4.545 73.555 4.715 ;
        RECT 73.385 4.165 73.555 4.335 ;
        RECT 74.085 4.55 74.255 4.72 ;
        RECT 74.085 4.16 74.255 4.33 ;
        RECT 75.075 4.55 75.245 4.72 ;
        RECT 75.075 4.16 75.245 4.33 ;
        RECT 76.49 4.285 76.66 4.455 ;
        RECT 76.95 4.285 77.12 4.455 ;
        RECT 77.41 4.285 77.58 4.455 ;
        RECT 77.87 4.285 78.04 4.455 ;
        RECT 78.33 4.285 78.5 4.455 ;
        RECT 78.79 4.285 78.96 4.455 ;
        RECT 79.25 4.285 79.42 4.455 ;
        RECT 79.71 4.285 79.88 4.455 ;
        RECT 80.17 4.285 80.34 4.455 ;
        RECT 80.63 4.285 80.8 4.455 ;
        RECT 81.09 4.285 81.26 4.455 ;
        RECT 81.55 4.285 81.72 4.455 ;
        RECT 82.01 4.285 82.18 4.455 ;
        RECT 82.47 4.285 82.64 4.455 ;
        RECT 82.93 4.285 83.1 4.455 ;
        RECT 83.39 4.285 83.56 4.455 ;
        RECT 83.85 4.285 84.02 4.455 ;
        RECT 84.31 4.285 84.48 4.455 ;
        RECT 84.77 4.285 84.94 4.455 ;
        RECT 85.23 4.285 85.4 4.455 ;
        RECT 85.69 4.285 85.86 4.455 ;
        RECT 86.15 4.285 86.32 4.455 ;
        RECT 86.55 4.545 86.72 4.715 ;
        RECT 86.61 4.285 86.78 4.455 ;
        RECT 87.07 4.285 87.24 4.455 ;
        RECT 87.53 4.285 87.7 4.455 ;
        RECT 87.99 4.285 88.16 4.455 ;
        RECT 91.31 4.545 91.48 4.715 ;
        RECT 91.31 4.165 91.48 4.335 ;
        RECT 92.01 4.55 92.18 4.72 ;
        RECT 92.01 4.16 92.18 4.33 ;
        RECT 93 4.55 93.17 4.72 ;
        RECT 93 4.16 93.17 4.33 ;
    END
  END vccd1
  OBS
    LAYER met3 ;
      RECT 85.7 7.055 86.075 7.425 ;
      RECT 85.735 4.925 86.045 7.425 ;
      RECT 85.735 4.925 88.83 5.235 ;
      RECT 88.52 1.125 88.83 5.235 ;
      RECT 88.52 1.14 88.895 1.51 ;
      RECT 85.65 3.685 86.205 4.015 ;
      RECT 85.65 2.02 85.95 4.015 ;
      RECT 81.715 3.125 82.27 3.455 ;
      RECT 81.97 2.02 82.27 3.455 ;
      RECT 82.765 1.885 82.915 2.535 ;
      RECT 81.97 2.02 85.95 2.32 ;
      RECT 80.485 0.96 80.785 3.91 ;
      RECT 80.475 2.565 81.205 2.895 ;
      RECT 80.44 0.96 80.815 1.33 ;
      RECT 79.035 3.125 79.765 3.455 ;
      RECT 79.05 0.96 79.35 3.455 ;
      RECT 76.925 2.565 77.655 2.895 ;
      RECT 77.08 0.93 77.38 2.895 ;
      RECT 79.005 0.96 79.38 1.33 ;
      RECT 77.035 0.93 77.41 1.3 ;
      RECT 77.035 0.97 79.38 1.27 ;
      RECT 67.775 7.055 68.15 7.425 ;
      RECT 67.81 4.925 68.12 7.425 ;
      RECT 67.81 4.925 70.905 5.235 ;
      RECT 70.595 1.125 70.905 5.235 ;
      RECT 70.595 1.14 70.97 1.51 ;
      RECT 67.725 3.685 68.28 4.015 ;
      RECT 67.725 2.02 68.025 4.015 ;
      RECT 63.79 3.125 64.345 3.455 ;
      RECT 64.045 2.02 64.345 3.455 ;
      RECT 64.84 1.885 64.99 2.535 ;
      RECT 64.045 2.02 68.025 2.32 ;
      RECT 62.56 0.96 62.86 3.91 ;
      RECT 62.55 2.565 63.28 2.895 ;
      RECT 62.515 0.96 62.89 1.33 ;
      RECT 61.11 3.125 61.84 3.455 ;
      RECT 61.125 0.96 61.425 3.455 ;
      RECT 59 2.565 59.73 2.895 ;
      RECT 59.155 0.93 59.455 2.895 ;
      RECT 61.08 0.96 61.455 1.33 ;
      RECT 59.11 0.93 59.485 1.3 ;
      RECT 59.11 0.97 61.455 1.27 ;
      RECT 49.85 7.055 50.225 7.425 ;
      RECT 49.885 4.925 50.195 7.425 ;
      RECT 49.885 4.925 52.98 5.235 ;
      RECT 52.67 1.125 52.98 5.235 ;
      RECT 52.67 1.14 53.045 1.51 ;
      RECT 49.8 3.685 50.355 4.015 ;
      RECT 49.8 2.02 50.1 4.015 ;
      RECT 45.865 3.125 46.42 3.455 ;
      RECT 46.12 2.02 46.42 3.455 ;
      RECT 46.915 1.885 47.065 2.535 ;
      RECT 46.12 2.02 50.1 2.32 ;
      RECT 44.635 0.96 44.935 3.91 ;
      RECT 44.625 2.565 45.355 2.895 ;
      RECT 44.59 0.96 44.965 1.33 ;
      RECT 43.185 3.125 43.915 3.455 ;
      RECT 43.2 0.96 43.5 3.455 ;
      RECT 41.075 2.565 41.805 2.895 ;
      RECT 41.23 0.93 41.53 2.895 ;
      RECT 43.155 0.96 43.53 1.33 ;
      RECT 41.185 0.93 41.56 1.3 ;
      RECT 41.185 0.97 43.53 1.27 ;
      RECT 31.925 7.055 32.3 7.425 ;
      RECT 31.96 4.925 32.27 7.425 ;
      RECT 31.96 4.925 35.055 5.235 ;
      RECT 34.745 1.125 35.055 5.235 ;
      RECT 34.745 1.14 35.12 1.51 ;
      RECT 31.875 3.685 32.43 4.015 ;
      RECT 31.875 2.02 32.175 4.015 ;
      RECT 27.94 3.125 28.495 3.455 ;
      RECT 28.195 2.02 28.495 3.455 ;
      RECT 28.99 1.885 29.14 2.535 ;
      RECT 28.195 2.02 32.175 2.32 ;
      RECT 26.71 0.96 27.01 3.91 ;
      RECT 26.7 2.565 27.43 2.895 ;
      RECT 26.665 0.96 27.04 1.33 ;
      RECT 25.26 3.125 25.99 3.455 ;
      RECT 25.275 0.96 25.575 3.455 ;
      RECT 23.15 2.565 23.88 2.895 ;
      RECT 23.305 0.93 23.605 2.895 ;
      RECT 25.23 0.96 25.605 1.33 ;
      RECT 23.26 0.93 23.635 1.3 ;
      RECT 23.26 0.97 25.605 1.27 ;
      RECT 14 7.055 14.375 7.425 ;
      RECT 14.035 4.925 14.345 7.425 ;
      RECT 14.035 4.925 17.13 5.235 ;
      RECT 16.82 1.125 17.13 5.235 ;
      RECT 16.82 1.14 17.195 1.51 ;
      RECT 13.95 3.685 14.505 4.015 ;
      RECT 13.95 2.02 14.25 4.015 ;
      RECT 10.015 3.125 10.57 3.455 ;
      RECT 10.27 2.02 10.57 3.455 ;
      RECT 11.065 1.885 11.215 2.535 ;
      RECT 10.27 2.02 14.25 2.32 ;
      RECT 8.785 0.96 9.085 3.91 ;
      RECT 8.775 2.565 9.505 2.895 ;
      RECT 8.74 0.96 9.115 1.33 ;
      RECT 7.335 3.125 8.065 3.455 ;
      RECT 7.35 0.96 7.65 3.455 ;
      RECT 5.225 2.565 5.955 2.895 ;
      RECT 5.38 0.93 5.68 2.895 ;
      RECT 7.305 0.96 7.68 1.33 ;
      RECT 5.335 0.93 5.71 1.3 ;
      RECT 5.335 0.97 7.68 1.27 ;
      RECT 86.835 2.005 87.565 2.335 ;
      RECT 84.615 3.685 85.345 4.015 ;
      RECT 82.915 3.685 83.645 4.015 ;
      RECT 77.96 2.565 78.69 2.895 ;
      RECT 76.595 3.685 77.325 4.015 ;
      RECT 68.91 2.005 69.64 2.335 ;
      RECT 66.69 3.685 67.42 4.015 ;
      RECT 64.99 3.685 65.72 4.015 ;
      RECT 60.035 2.565 60.765 2.895 ;
      RECT 58.67 3.685 59.4 4.015 ;
      RECT 50.985 2.005 51.715 2.335 ;
      RECT 48.765 3.685 49.495 4.015 ;
      RECT 47.065 3.685 47.795 4.015 ;
      RECT 42.11 2.565 42.84 2.895 ;
      RECT 40.745 3.685 41.475 4.015 ;
      RECT 33.06 2.005 33.79 2.335 ;
      RECT 30.84 3.685 31.57 4.015 ;
      RECT 29.14 3.685 29.87 4.015 ;
      RECT 24.185 2.565 24.915 2.895 ;
      RECT 22.82 3.685 23.55 4.015 ;
      RECT 15.135 2.005 15.865 2.335 ;
      RECT 12.915 3.685 13.645 4.015 ;
      RECT 11.215 3.685 11.945 4.015 ;
      RECT 6.26 2.565 6.99 2.895 ;
      RECT 4.895 3.685 5.625 4.015 ;
    LAYER via2 ;
      RECT 88.61 1.225 88.81 1.425 ;
      RECT 86.9 2.07 87.1 2.27 ;
      RECT 85.94 3.75 86.14 3.95 ;
      RECT 85.79 7.14 85.99 7.34 ;
      RECT 84.94 3.75 85.14 3.95 ;
      RECT 82.98 3.75 83.18 3.95 ;
      RECT 81.78 3.19 81.98 3.39 ;
      RECT 80.54 2.63 80.74 2.83 ;
      RECT 80.53 1.045 80.73 1.245 ;
      RECT 79.1 3.19 79.3 3.39 ;
      RECT 79.095 1.04 79.295 1.24 ;
      RECT 78.36 2.63 78.56 2.83 ;
      RECT 77.14 2.63 77.34 2.83 ;
      RECT 77.125 1.015 77.325 1.215 ;
      RECT 76.66 3.75 76.86 3.95 ;
      RECT 70.685 1.225 70.885 1.425 ;
      RECT 68.975 2.07 69.175 2.27 ;
      RECT 68.015 3.75 68.215 3.95 ;
      RECT 67.865 7.14 68.065 7.34 ;
      RECT 67.015 3.75 67.215 3.95 ;
      RECT 65.055 3.75 65.255 3.95 ;
      RECT 63.855 3.19 64.055 3.39 ;
      RECT 62.615 2.63 62.815 2.83 ;
      RECT 62.605 1.045 62.805 1.245 ;
      RECT 61.175 3.19 61.375 3.39 ;
      RECT 61.17 1.04 61.37 1.24 ;
      RECT 60.435 2.63 60.635 2.83 ;
      RECT 59.215 2.63 59.415 2.83 ;
      RECT 59.2 1.015 59.4 1.215 ;
      RECT 58.735 3.75 58.935 3.95 ;
      RECT 52.76 1.225 52.96 1.425 ;
      RECT 51.05 2.07 51.25 2.27 ;
      RECT 50.09 3.75 50.29 3.95 ;
      RECT 49.94 7.14 50.14 7.34 ;
      RECT 49.09 3.75 49.29 3.95 ;
      RECT 47.13 3.75 47.33 3.95 ;
      RECT 45.93 3.19 46.13 3.39 ;
      RECT 44.69 2.63 44.89 2.83 ;
      RECT 44.68 1.045 44.88 1.245 ;
      RECT 43.25 3.19 43.45 3.39 ;
      RECT 43.245 1.04 43.445 1.24 ;
      RECT 42.51 2.63 42.71 2.83 ;
      RECT 41.29 2.63 41.49 2.83 ;
      RECT 41.275 1.015 41.475 1.215 ;
      RECT 40.81 3.75 41.01 3.95 ;
      RECT 34.835 1.225 35.035 1.425 ;
      RECT 33.125 2.07 33.325 2.27 ;
      RECT 32.165 3.75 32.365 3.95 ;
      RECT 32.015 7.14 32.215 7.34 ;
      RECT 31.165 3.75 31.365 3.95 ;
      RECT 29.205 3.75 29.405 3.95 ;
      RECT 28.005 3.19 28.205 3.39 ;
      RECT 26.765 2.63 26.965 2.83 ;
      RECT 26.755 1.045 26.955 1.245 ;
      RECT 25.325 3.19 25.525 3.39 ;
      RECT 25.32 1.04 25.52 1.24 ;
      RECT 24.585 2.63 24.785 2.83 ;
      RECT 23.365 2.63 23.565 2.83 ;
      RECT 23.35 1.015 23.55 1.215 ;
      RECT 22.885 3.75 23.085 3.95 ;
      RECT 16.91 1.225 17.11 1.425 ;
      RECT 15.2 2.07 15.4 2.27 ;
      RECT 14.24 3.75 14.44 3.95 ;
      RECT 14.09 7.14 14.29 7.34 ;
      RECT 13.24 3.75 13.44 3.95 ;
      RECT 11.28 3.75 11.48 3.95 ;
      RECT 10.08 3.19 10.28 3.39 ;
      RECT 8.84 2.63 9.04 2.83 ;
      RECT 8.83 1.045 9.03 1.245 ;
      RECT 7.4 3.19 7.6 3.39 ;
      RECT 7.395 1.04 7.595 1.24 ;
      RECT 6.66 2.63 6.86 2.83 ;
      RECT 5.44 2.63 5.64 2.83 ;
      RECT 5.425 1.015 5.625 1.215 ;
      RECT 4.96 3.75 5.16 3.95 ;
    LAYER met2 ;
      RECT 2.7 8.4 93.52 8.57 ;
      RECT 93.35 7.275 93.52 8.57 ;
      RECT 2.7 6.255 2.87 8.57 ;
      RECT 93.32 7.275 93.67 7.625 ;
      RECT 2.645 6.255 2.935 6.605 ;
      RECT 90.165 6.225 90.485 6.545 ;
      RECT 90.195 5.695 90.365 6.545 ;
      RECT 90.195 5.695 90.37 6.045 ;
      RECT 90.195 5.695 91.17 5.87 ;
      RECT 90.995 1.965 91.17 5.87 ;
      RECT 90.94 1.965 91.29 2.315 ;
      RECT 90.965 6.655 91.29 6.98 ;
      RECT 89.85 6.745 91.29 6.915 ;
      RECT 89.85 2.395 90.01 6.915 ;
      RECT 90.165 2.365 90.485 2.685 ;
      RECT 89.85 2.395 90.485 2.565 ;
      RECT 88.52 1.14 88.895 1.51 ;
      RECT 80.44 0.96 80.815 1.33 ;
      RECT 79.005 0.96 79.38 1.33 ;
      RECT 79.005 1.08 88.825 1.25 ;
      RECT 84.95 4.36 88.805 4.53 ;
      RECT 88.635 3.425 88.805 4.53 ;
      RECT 84.95 3.67 85.12 4.53 ;
      RECT 84.9 3.71 85.18 3.99 ;
      RECT 84.92 3.67 85.18 3.99 ;
      RECT 84.56 3.625 84.665 3.885 ;
      RECT 88.545 3.43 88.895 3.78 ;
      RECT 84.415 2.115 84.505 2.375 ;
      RECT 84.955 3.18 84.96 3.22 ;
      RECT 84.95 3.17 84.955 3.305 ;
      RECT 84.945 3.16 84.95 3.398 ;
      RECT 84.935 3.14 84.945 3.454 ;
      RECT 84.855 3.068 84.935 3.534 ;
      RECT 84.89 3.712 84.9 3.937 ;
      RECT 84.885 3.709 84.89 3.932 ;
      RECT 84.87 3.706 84.885 3.925 ;
      RECT 84.835 3.7 84.87 3.907 ;
      RECT 84.85 3.003 84.855 3.608 ;
      RECT 84.83 2.954 84.85 3.623 ;
      RECT 84.82 3.687 84.835 3.89 ;
      RECT 84.825 2.896 84.83 3.638 ;
      RECT 84.82 2.874 84.825 3.648 ;
      RECT 84.785 2.784 84.82 3.885 ;
      RECT 84.77 2.662 84.785 3.885 ;
      RECT 84.765 2.615 84.77 3.885 ;
      RECT 84.74 2.54 84.765 3.885 ;
      RECT 84.725 2.455 84.74 3.885 ;
      RECT 84.72 2.402 84.725 3.885 ;
      RECT 84.715 2.382 84.72 3.885 ;
      RECT 84.71 2.357 84.715 3.119 ;
      RECT 84.695 3.317 84.715 3.885 ;
      RECT 84.705 2.335 84.71 3.096 ;
      RECT 84.695 2.287 84.705 3.061 ;
      RECT 84.69 2.25 84.695 3.027 ;
      RECT 84.69 3.397 84.695 3.885 ;
      RECT 84.675 2.227 84.69 2.982 ;
      RECT 84.67 3.495 84.69 3.885 ;
      RECT 84.62 2.115 84.675 2.824 ;
      RECT 84.665 3.617 84.67 3.885 ;
      RECT 84.605 2.115 84.62 2.663 ;
      RECT 84.6 2.115 84.605 2.615 ;
      RECT 84.595 2.115 84.6 2.603 ;
      RECT 84.55 2.115 84.595 2.54 ;
      RECT 84.525 2.115 84.55 2.458 ;
      RECT 84.51 2.115 84.525 2.41 ;
      RECT 84.505 2.115 84.51 2.38 ;
      RECT 86.895 2.16 87.155 2.42 ;
      RECT 86.89 2.16 87.155 2.368 ;
      RECT 86.885 2.16 87.155 2.338 ;
      RECT 86.86 2.03 87.14 2.31 ;
      RECT 75.375 6.655 75.725 7.005 ;
      RECT 86.62 6.61 86.97 6.96 ;
      RECT 75.375 6.685 86.97 6.885 ;
      RECT 85.9 3.71 86.18 3.99 ;
      RECT 85.94 3.665 86.205 3.925 ;
      RECT 85.93 3.7 86.205 3.925 ;
      RECT 85.935 3.685 86.18 3.99 ;
      RECT 85.94 3.662 86.15 3.99 ;
      RECT 85.94 3.66 86.135 3.99 ;
      RECT 85.98 3.65 86.135 3.99 ;
      RECT 85.95 3.655 86.135 3.99 ;
      RECT 85.98 3.647 86.08 3.99 ;
      RECT 86.005 3.64 86.08 3.99 ;
      RECT 85.985 3.642 86.08 3.99 ;
      RECT 85.315 3.155 85.575 3.415 ;
      RECT 85.365 3.147 85.555 3.415 ;
      RECT 85.37 3.067 85.555 3.415 ;
      RECT 85.49 2.455 85.555 3.415 ;
      RECT 85.395 2.852 85.555 3.415 ;
      RECT 85.47 2.54 85.555 3.415 ;
      RECT 85.505 2.165 85.641 2.893 ;
      RECT 85.45 2.662 85.641 2.893 ;
      RECT 85.465 2.602 85.555 3.415 ;
      RECT 85.505 2.165 85.665 2.558 ;
      RECT 85.505 2.165 85.675 2.455 ;
      RECT 85.495 2.165 85.755 2.425 ;
      RECT 83.83 3.565 83.875 3.825 ;
      RECT 83.735 2.1 83.88 2.36 ;
      RECT 84.24 2.722 84.25 2.813 ;
      RECT 84.225 2.66 84.24 2.869 ;
      RECT 84.22 2.607 84.225 2.915 ;
      RECT 84.17 2.554 84.22 3.041 ;
      RECT 84.165 2.509 84.17 3.188 ;
      RECT 84.155 2.497 84.165 3.23 ;
      RECT 84.12 2.461 84.155 3.335 ;
      RECT 84.115 2.429 84.12 3.441 ;
      RECT 84.1 2.411 84.115 3.486 ;
      RECT 84.095 2.394 84.1 2.72 ;
      RECT 84.09 2.775 84.1 3.543 ;
      RECT 84.085 2.38 84.095 2.693 ;
      RECT 84.08 2.83 84.09 3.825 ;
      RECT 84.075 2.366 84.085 2.678 ;
      RECT 84.075 2.88 84.08 3.825 ;
      RECT 84.06 2.343 84.075 2.658 ;
      RECT 84.04 3.002 84.075 3.825 ;
      RECT 84.055 2.325 84.06 2.64 ;
      RECT 84.05 2.317 84.055 2.63 ;
      RECT 84.02 2.285 84.05 2.594 ;
      RECT 84.03 3.13 84.04 3.825 ;
      RECT 84.025 3.157 84.03 3.825 ;
      RECT 84.02 3.207 84.025 3.825 ;
      RECT 84.01 2.251 84.02 2.559 ;
      RECT 83.97 3.275 84.02 3.825 ;
      RECT 83.995 2.228 84.01 2.535 ;
      RECT 83.97 2.1 83.995 2.498 ;
      RECT 83.965 2.1 83.97 2.47 ;
      RECT 83.935 3.375 83.97 3.825 ;
      RECT 83.96 2.1 83.965 2.463 ;
      RECT 83.955 2.1 83.96 2.453 ;
      RECT 83.94 2.1 83.955 2.438 ;
      RECT 83.925 2.1 83.94 2.41 ;
      RECT 83.89 3.48 83.935 3.825 ;
      RECT 83.91 2.1 83.925 2.383 ;
      RECT 83.88 2.1 83.91 2.368 ;
      RECT 83.875 3.552 83.89 3.825 ;
      RECT 83.8 2.635 83.84 2.895 ;
      RECT 83.575 2.582 83.58 2.84 ;
      RECT 79.53 2.06 79.79 2.32 ;
      RECT 79.53 2.085 79.805 2.3 ;
      RECT 81.92 1.91 81.925 2.055 ;
      RECT 83.79 2.63 83.8 2.895 ;
      RECT 83.77 2.622 83.79 2.895 ;
      RECT 83.752 2.618 83.77 2.895 ;
      RECT 83.666 2.607 83.752 2.895 ;
      RECT 83.58 2.59 83.666 2.895 ;
      RECT 83.525 2.577 83.575 2.825 ;
      RECT 83.491 2.569 83.525 2.8 ;
      RECT 83.405 2.558 83.491 2.765 ;
      RECT 83.37 2.535 83.405 2.73 ;
      RECT 83.36 2.497 83.37 2.716 ;
      RECT 83.355 2.47 83.36 2.712 ;
      RECT 83.35 2.457 83.355 2.709 ;
      RECT 83.34 2.437 83.35 2.705 ;
      RECT 83.335 2.412 83.34 2.701 ;
      RECT 83.31 2.367 83.335 2.695 ;
      RECT 83.3 2.308 83.31 2.687 ;
      RECT 83.29 2.276 83.3 2.678 ;
      RECT 83.27 2.228 83.29 2.658 ;
      RECT 83.265 2.188 83.27 2.628 ;
      RECT 83.25 2.162 83.265 2.602 ;
      RECT 83.245 2.14 83.25 2.578 ;
      RECT 83.23 2.112 83.245 2.554 ;
      RECT 83.215 2.085 83.23 2.518 ;
      RECT 83.2 2.062 83.215 2.48 ;
      RECT 83.195 2.052 83.2 2.455 ;
      RECT 83.185 2.045 83.195 2.438 ;
      RECT 83.17 2.032 83.185 2.408 ;
      RECT 83.165 2.022 83.17 2.383 ;
      RECT 83.16 2.017 83.165 2.37 ;
      RECT 83.15 2.01 83.16 2.35 ;
      RECT 83.145 2.003 83.15 2.335 ;
      RECT 83.12 1.996 83.145 2.293 ;
      RECT 83.105 1.986 83.12 2.243 ;
      RECT 83.095 1.981 83.105 2.213 ;
      RECT 83.085 1.977 83.095 2.188 ;
      RECT 83.07 1.974 83.085 2.178 ;
      RECT 83.02 1.971 83.07 2.163 ;
      RECT 83 1.969 83.02 2.148 ;
      RECT 82.951 1.967 83 2.143 ;
      RECT 82.865 1.963 82.951 2.138 ;
      RECT 82.826 1.96 82.865 2.134 ;
      RECT 82.74 1.956 82.826 2.129 ;
      RECT 82.69 1.953 82.74 2.123 ;
      RECT 82.641 1.95 82.69 2.118 ;
      RECT 82.555 1.947 82.641 2.113 ;
      RECT 82.551 1.945 82.555 2.11 ;
      RECT 82.465 1.942 82.551 2.105 ;
      RECT 82.416 1.938 82.465 2.098 ;
      RECT 82.33 1.935 82.416 2.093 ;
      RECT 82.306 1.932 82.33 2.089 ;
      RECT 82.22 1.93 82.306 2.084 ;
      RECT 82.155 1.926 82.22 2.077 ;
      RECT 82.152 1.925 82.155 2.074 ;
      RECT 82.066 1.922 82.152 2.071 ;
      RECT 81.98 1.916 82.066 2.064 ;
      RECT 81.95 1.912 81.98 2.06 ;
      RECT 81.925 1.91 81.95 2.058 ;
      RECT 81.87 1.907 81.92 2.055 ;
      RECT 81.79 1.906 81.87 2.055 ;
      RECT 81.735 1.908 81.79 2.058 ;
      RECT 81.72 1.909 81.735 2.062 ;
      RECT 81.665 1.917 81.72 2.072 ;
      RECT 81.635 1.925 81.665 2.085 ;
      RECT 81.616 1.926 81.635 2.091 ;
      RECT 81.53 1.929 81.616 2.096 ;
      RECT 81.46 1.934 81.53 2.105 ;
      RECT 81.441 1.937 81.46 2.111 ;
      RECT 81.355 1.941 81.441 2.116 ;
      RECT 81.315 1.945 81.355 2.123 ;
      RECT 81.306 1.947 81.315 2.126 ;
      RECT 81.22 1.951 81.306 2.131 ;
      RECT 81.217 1.954 81.22 2.135 ;
      RECT 81.131 1.957 81.217 2.139 ;
      RECT 81.045 1.963 81.131 2.147 ;
      RECT 81.021 1.967 81.045 2.151 ;
      RECT 80.935 1.971 81.021 2.156 ;
      RECT 80.89 1.976 80.935 2.163 ;
      RECT 80.81 1.981 80.89 2.17 ;
      RECT 80.73 1.987 80.81 2.185 ;
      RECT 80.705 1.991 80.73 2.198 ;
      RECT 80.64 1.994 80.705 2.21 ;
      RECT 80.585 1.999 80.64 2.225 ;
      RECT 80.555 2.002 80.585 2.243 ;
      RECT 80.545 2.004 80.555 2.256 ;
      RECT 80.485 2.019 80.545 2.266 ;
      RECT 80.47 2.036 80.485 2.275 ;
      RECT 80.465 2.045 80.47 2.275 ;
      RECT 80.455 2.055 80.465 2.275 ;
      RECT 80.445 2.072 80.455 2.275 ;
      RECT 80.425 2.082 80.445 2.276 ;
      RECT 80.38 2.092 80.425 2.277 ;
      RECT 80.345 2.101 80.38 2.279 ;
      RECT 80.28 2.106 80.345 2.281 ;
      RECT 80.2 2.107 80.28 2.284 ;
      RECT 80.196 2.105 80.2 2.285 ;
      RECT 80.11 2.102 80.196 2.287 ;
      RECT 80.063 2.099 80.11 2.289 ;
      RECT 79.977 2.095 80.063 2.292 ;
      RECT 79.891 2.091 79.977 2.295 ;
      RECT 79.805 2.087 79.891 2.299 ;
      RECT 83.19 3.71 83.22 3.99 ;
      RECT 82.94 3.6 82.96 3.99 ;
      RECT 82.895 3.6 82.96 3.86 ;
      RECT 82.725 2.225 82.76 2.485 ;
      RECT 82.5 2.225 82.56 2.485 ;
      RECT 83.18 3.69 83.19 3.99 ;
      RECT 83.175 3.65 83.18 3.99 ;
      RECT 83.16 3.605 83.175 3.99 ;
      RECT 83.155 3.57 83.16 3.99 ;
      RECT 83.15 3.55 83.155 3.99 ;
      RECT 83.12 3.477 83.15 3.99 ;
      RECT 83.1 3.375 83.12 3.99 ;
      RECT 83.09 3.305 83.1 3.99 ;
      RECT 83.045 3.245 83.09 3.99 ;
      RECT 82.96 3.206 83.045 3.99 ;
      RECT 82.955 3.197 82.96 3.57 ;
      RECT 82.945 3.196 82.955 3.553 ;
      RECT 82.92 3.177 82.945 3.523 ;
      RECT 82.915 3.152 82.92 3.502 ;
      RECT 82.905 3.13 82.915 3.493 ;
      RECT 82.9 3.101 82.905 3.483 ;
      RECT 82.86 3.027 82.9 3.455 ;
      RECT 82.84 2.928 82.86 3.42 ;
      RECT 82.825 2.864 82.84 3.403 ;
      RECT 82.795 2.788 82.825 3.375 ;
      RECT 82.775 2.703 82.795 3.348 ;
      RECT 82.735 2.599 82.775 3.255 ;
      RECT 82.73 2.52 82.735 3.163 ;
      RECT 82.725 2.503 82.73 3.14 ;
      RECT 82.72 2.225 82.725 3.12 ;
      RECT 82.69 2.225 82.72 3.058 ;
      RECT 82.685 2.225 82.69 2.99 ;
      RECT 82.675 2.225 82.685 2.955 ;
      RECT 82.665 2.225 82.675 2.92 ;
      RECT 82.6 2.225 82.665 2.775 ;
      RECT 82.595 2.225 82.6 2.645 ;
      RECT 82.565 2.225 82.595 2.578 ;
      RECT 82.56 2.225 82.565 2.503 ;
      RECT 81.74 3.15 82.02 3.43 ;
      RECT 81.78 3.13 82.04 3.39 ;
      RECT 81.77 3.14 82.04 3.39 ;
      RECT 81.78 3.067 81.995 3.43 ;
      RECT 81.835 2.99 81.99 3.43 ;
      RECT 81.84 2.775 81.99 3.43 ;
      RECT 81.83 2.577 81.98 2.828 ;
      RECT 81.82 2.577 81.98 2.695 ;
      RECT 81.815 2.455 81.975 2.598 ;
      RECT 81.8 2.455 81.975 2.503 ;
      RECT 81.795 2.165 81.97 2.48 ;
      RECT 81.78 2.165 81.97 2.45 ;
      RECT 81.74 2.165 82 2.425 ;
      RECT 81.65 3.635 81.73 3.895 ;
      RECT 81.055 2.355 81.06 2.62 ;
      RECT 80.935 2.355 81.06 2.615 ;
      RECT 81.61 3.6 81.65 3.895 ;
      RECT 81.565 3.522 81.61 3.895 ;
      RECT 81.545 3.45 81.565 3.895 ;
      RECT 81.535 3.402 81.545 3.895 ;
      RECT 81.5 3.335 81.535 3.895 ;
      RECT 81.47 3.235 81.5 3.895 ;
      RECT 81.45 3.16 81.47 3.695 ;
      RECT 81.44 3.11 81.45 3.65 ;
      RECT 81.435 3.087 81.44 3.623 ;
      RECT 81.43 3.072 81.435 3.61 ;
      RECT 81.425 3.057 81.43 3.588 ;
      RECT 81.42 3.042 81.425 3.57 ;
      RECT 81.395 2.997 81.42 3.525 ;
      RECT 81.385 2.945 81.395 3.468 ;
      RECT 81.375 2.915 81.385 3.435 ;
      RECT 81.365 2.88 81.375 3.403 ;
      RECT 81.33 2.812 81.365 3.335 ;
      RECT 81.325 2.751 81.33 3.27 ;
      RECT 81.315 2.739 81.325 3.25 ;
      RECT 81.31 2.727 81.315 3.23 ;
      RECT 81.305 2.719 81.31 3.218 ;
      RECT 81.3 2.711 81.305 3.198 ;
      RECT 81.29 2.699 81.3 3.17 ;
      RECT 81.28 2.683 81.29 3.14 ;
      RECT 81.255 2.655 81.28 3.078 ;
      RECT 81.245 2.626 81.255 3.023 ;
      RECT 81.23 2.605 81.245 2.983 ;
      RECT 81.225 2.589 81.23 2.955 ;
      RECT 81.22 2.577 81.225 2.945 ;
      RECT 81.215 2.572 81.22 2.918 ;
      RECT 81.21 2.565 81.215 2.905 ;
      RECT 81.195 2.548 81.21 2.878 ;
      RECT 81.185 2.355 81.195 2.838 ;
      RECT 81.175 2.355 81.185 2.805 ;
      RECT 81.165 2.355 81.175 2.78 ;
      RECT 81.095 2.355 81.165 2.715 ;
      RECT 81.085 2.355 81.095 2.663 ;
      RECT 81.07 2.355 81.085 2.645 ;
      RECT 81.06 2.355 81.07 2.63 ;
      RECT 80.89 3.225 81.15 3.485 ;
      RECT 79.425 3.26 79.43 3.467 ;
      RECT 79.06 3.15 79.135 3.465 ;
      RECT 78.875 3.205 79.03 3.465 ;
      RECT 79.06 3.15 79.165 3.43 ;
      RECT 80.875 3.322 80.89 3.483 ;
      RECT 80.85 3.33 80.875 3.488 ;
      RECT 80.825 3.337 80.85 3.493 ;
      RECT 80.762 3.348 80.825 3.502 ;
      RECT 80.676 3.367 80.762 3.519 ;
      RECT 80.59 3.389 80.676 3.538 ;
      RECT 80.575 3.402 80.59 3.549 ;
      RECT 80.535 3.41 80.575 3.556 ;
      RECT 80.515 3.415 80.535 3.563 ;
      RECT 80.477 3.416 80.515 3.566 ;
      RECT 80.391 3.419 80.477 3.567 ;
      RECT 80.305 3.423 80.391 3.568 ;
      RECT 80.256 3.425 80.305 3.57 ;
      RECT 80.17 3.425 80.256 3.572 ;
      RECT 80.13 3.42 80.17 3.574 ;
      RECT 80.12 3.414 80.13 3.575 ;
      RECT 80.08 3.409 80.12 3.572 ;
      RECT 80.07 3.402 80.08 3.568 ;
      RECT 80.055 3.398 80.07 3.566 ;
      RECT 80.038 3.394 80.055 3.564 ;
      RECT 79.952 3.384 80.038 3.556 ;
      RECT 79.866 3.366 79.952 3.542 ;
      RECT 79.78 3.349 79.866 3.528 ;
      RECT 79.755 3.337 79.78 3.519 ;
      RECT 79.685 3.327 79.755 3.512 ;
      RECT 79.64 3.315 79.685 3.503 ;
      RECT 79.58 3.302 79.64 3.495 ;
      RECT 79.575 3.294 79.58 3.49 ;
      RECT 79.54 3.289 79.575 3.488 ;
      RECT 79.485 3.28 79.54 3.481 ;
      RECT 79.445 3.269 79.485 3.473 ;
      RECT 79.43 3.262 79.445 3.469 ;
      RECT 79.41 3.255 79.425 3.466 ;
      RECT 79.395 3.245 79.41 3.464 ;
      RECT 79.38 3.232 79.395 3.461 ;
      RECT 79.355 3.215 79.38 3.457 ;
      RECT 79.34 3.197 79.355 3.454 ;
      RECT 79.315 3.15 79.34 3.452 ;
      RECT 79.291 3.15 79.315 3.449 ;
      RECT 79.205 3.15 79.291 3.441 ;
      RECT 79.165 3.15 79.205 3.433 ;
      RECT 79.03 3.197 79.06 3.465 ;
      RECT 80.71 2.78 80.97 3.04 ;
      RECT 80.67 2.78 80.97 2.918 ;
      RECT 80.635 2.78 80.97 2.903 ;
      RECT 80.58 2.78 80.97 2.883 ;
      RECT 80.5 2.59 80.78 2.87 ;
      RECT 80.5 2.772 80.85 2.87 ;
      RECT 80.5 2.715 80.835 2.87 ;
      RECT 80.5 2.662 80.785 2.87 ;
      RECT 78.33 2.59 78.525 3.375 ;
      RECT 78.41 1.205 78.525 3.375 ;
      RECT 78.265 3.115 78.325 3.375 ;
      RECT 79.635 2.635 79.895 2.895 ;
      RECT 78.32 2.59 78.525 2.87 ;
      RECT 79.63 2.645 79.895 2.83 ;
      RECT 79.345 2.62 79.355 2.77 ;
      RECT 78.58 1.205 78.66 1.55 ;
      RECT 78.315 1.205 78.525 1.55 ;
      RECT 79.62 2.645 79.63 2.829 ;
      RECT 79.61 2.644 79.62 2.826 ;
      RECT 79.601 2.643 79.61 2.824 ;
      RECT 79.515 2.639 79.601 2.814 ;
      RECT 79.441 2.631 79.515 2.796 ;
      RECT 79.355 2.624 79.441 2.779 ;
      RECT 79.295 2.62 79.345 2.769 ;
      RECT 79.26 2.619 79.295 2.766 ;
      RECT 79.205 2.619 79.26 2.768 ;
      RECT 79.17 2.619 79.205 2.772 ;
      RECT 79.084 2.618 79.17 2.779 ;
      RECT 78.998 2.617 79.084 2.789 ;
      RECT 78.912 2.616 78.998 2.8 ;
      RECT 78.826 2.616 78.912 2.81 ;
      RECT 78.74 2.615 78.826 2.82 ;
      RECT 78.705 2.615 78.74 2.86 ;
      RECT 78.7 2.615 78.705 2.903 ;
      RECT 78.675 2.615 78.7 2.92 ;
      RECT 78.6 2.615 78.675 2.935 ;
      RECT 78.58 2.59 78.6 2.948 ;
      RECT 78.575 1.205 78.58 2.958 ;
      RECT 78.55 1.205 78.575 3 ;
      RECT 78.525 1.205 78.55 3.078 ;
      RECT 78.325 2.997 78.33 3.375 ;
      RECT 77.66 2.949 77.675 3.405 ;
      RECT 77.655 3.021 77.761 3.403 ;
      RECT 77.675 2.115 77.81 3.401 ;
      RECT 77.66 2.965 77.815 3.4 ;
      RECT 77.66 3.015 77.82 3.398 ;
      RECT 77.645 3.08 77.82 3.397 ;
      RECT 77.655 3.072 77.825 3.394 ;
      RECT 77.635 3.12 77.825 3.389 ;
      RECT 77.635 3.12 77.84 3.386 ;
      RECT 77.63 3.12 77.84 3.383 ;
      RECT 77.605 3.12 77.865 3.38 ;
      RECT 77.675 2.115 77.835 2.768 ;
      RECT 77.67 2.115 77.835 2.74 ;
      RECT 77.665 2.115 77.835 2.568 ;
      RECT 77.665 2.115 77.855 2.508 ;
      RECT 77.62 2.115 77.88 2.375 ;
      RECT 77.1 2.59 77.38 2.87 ;
      RECT 77.09 2.605 77.38 2.865 ;
      RECT 77.045 2.667 77.38 2.863 ;
      RECT 77.12 2.582 77.285 2.87 ;
      RECT 77.12 2.567 77.241 2.87 ;
      RECT 77.155 2.56 77.241 2.87 ;
      RECT 76.62 3.71 76.9 3.99 ;
      RECT 76.58 3.672 76.875 3.783 ;
      RECT 76.565 3.622 76.855 3.678 ;
      RECT 76.51 3.385 76.77 3.645 ;
      RECT 76.51 3.587 76.85 3.645 ;
      RECT 76.51 3.527 76.845 3.645 ;
      RECT 76.51 3.477 76.825 3.645 ;
      RECT 76.51 3.457 76.82 3.645 ;
      RECT 76.51 3.435 76.815 3.645 ;
      RECT 76.51 3.42 76.785 3.645 ;
      RECT 72.24 6.225 72.56 6.545 ;
      RECT 72.27 5.695 72.44 6.545 ;
      RECT 72.27 5.695 72.445 6.045 ;
      RECT 72.27 5.695 73.245 5.87 ;
      RECT 73.07 1.965 73.245 5.87 ;
      RECT 73.015 1.965 73.365 2.315 ;
      RECT 73.04 6.655 73.365 6.98 ;
      RECT 71.925 6.745 73.365 6.915 ;
      RECT 71.925 2.395 72.085 6.915 ;
      RECT 72.24 2.365 72.56 2.685 ;
      RECT 71.925 2.395 72.56 2.565 ;
      RECT 70.595 1.14 70.97 1.51 ;
      RECT 62.515 0.96 62.89 1.33 ;
      RECT 61.08 0.96 61.455 1.33 ;
      RECT 61.08 1.08 70.9 1.25 ;
      RECT 67.025 4.36 70.88 4.53 ;
      RECT 70.71 3.425 70.88 4.53 ;
      RECT 67.025 3.67 67.195 4.53 ;
      RECT 66.975 3.71 67.255 3.99 ;
      RECT 66.995 3.67 67.255 3.99 ;
      RECT 66.635 3.625 66.74 3.885 ;
      RECT 70.62 3.43 70.97 3.78 ;
      RECT 66.49 2.115 66.58 2.375 ;
      RECT 67.03 3.18 67.035 3.22 ;
      RECT 67.025 3.17 67.03 3.305 ;
      RECT 67.02 3.16 67.025 3.398 ;
      RECT 67.01 3.14 67.02 3.454 ;
      RECT 66.93 3.068 67.01 3.534 ;
      RECT 66.965 3.712 66.975 3.937 ;
      RECT 66.96 3.709 66.965 3.932 ;
      RECT 66.945 3.706 66.96 3.925 ;
      RECT 66.91 3.7 66.945 3.907 ;
      RECT 66.925 3.003 66.93 3.608 ;
      RECT 66.905 2.954 66.925 3.623 ;
      RECT 66.895 3.687 66.91 3.89 ;
      RECT 66.9 2.896 66.905 3.638 ;
      RECT 66.895 2.874 66.9 3.648 ;
      RECT 66.86 2.784 66.895 3.885 ;
      RECT 66.845 2.662 66.86 3.885 ;
      RECT 66.84 2.615 66.845 3.885 ;
      RECT 66.815 2.54 66.84 3.885 ;
      RECT 66.8 2.455 66.815 3.885 ;
      RECT 66.795 2.402 66.8 3.885 ;
      RECT 66.79 2.382 66.795 3.885 ;
      RECT 66.785 2.357 66.79 3.119 ;
      RECT 66.77 3.317 66.79 3.885 ;
      RECT 66.78 2.335 66.785 3.096 ;
      RECT 66.77 2.287 66.78 3.061 ;
      RECT 66.765 2.25 66.77 3.027 ;
      RECT 66.765 3.397 66.77 3.885 ;
      RECT 66.75 2.227 66.765 2.982 ;
      RECT 66.745 3.495 66.765 3.885 ;
      RECT 66.695 2.115 66.75 2.824 ;
      RECT 66.74 3.617 66.745 3.885 ;
      RECT 66.68 2.115 66.695 2.663 ;
      RECT 66.675 2.115 66.68 2.615 ;
      RECT 66.67 2.115 66.675 2.603 ;
      RECT 66.625 2.115 66.67 2.54 ;
      RECT 66.6 2.115 66.625 2.458 ;
      RECT 66.585 2.115 66.6 2.41 ;
      RECT 66.58 2.115 66.585 2.38 ;
      RECT 68.97 2.16 69.23 2.42 ;
      RECT 68.965 2.16 69.23 2.368 ;
      RECT 68.96 2.16 69.23 2.338 ;
      RECT 68.935 2.03 69.215 2.31 ;
      RECT 57.45 6.655 57.8 7.005 ;
      RECT 68.415 6.61 68.765 6.96 ;
      RECT 57.45 6.685 68.765 6.885 ;
      RECT 67.975 3.71 68.255 3.99 ;
      RECT 68.015 3.665 68.28 3.925 ;
      RECT 68.005 3.7 68.28 3.925 ;
      RECT 68.01 3.685 68.255 3.99 ;
      RECT 68.015 3.662 68.225 3.99 ;
      RECT 68.015 3.66 68.21 3.99 ;
      RECT 68.055 3.65 68.21 3.99 ;
      RECT 68.025 3.655 68.21 3.99 ;
      RECT 68.055 3.647 68.155 3.99 ;
      RECT 68.08 3.64 68.155 3.99 ;
      RECT 68.06 3.642 68.155 3.99 ;
      RECT 67.39 3.155 67.65 3.415 ;
      RECT 67.44 3.147 67.63 3.415 ;
      RECT 67.445 3.067 67.63 3.415 ;
      RECT 67.565 2.455 67.63 3.415 ;
      RECT 67.47 2.852 67.63 3.415 ;
      RECT 67.545 2.54 67.63 3.415 ;
      RECT 67.58 2.165 67.716 2.893 ;
      RECT 67.525 2.662 67.716 2.893 ;
      RECT 67.54 2.602 67.63 3.415 ;
      RECT 67.58 2.165 67.74 2.558 ;
      RECT 67.58 2.165 67.75 2.455 ;
      RECT 67.57 2.165 67.83 2.425 ;
      RECT 65.905 3.565 65.95 3.825 ;
      RECT 65.81 2.1 65.955 2.36 ;
      RECT 66.315 2.722 66.325 2.813 ;
      RECT 66.3 2.66 66.315 2.869 ;
      RECT 66.295 2.607 66.3 2.915 ;
      RECT 66.245 2.554 66.295 3.041 ;
      RECT 66.24 2.509 66.245 3.188 ;
      RECT 66.23 2.497 66.24 3.23 ;
      RECT 66.195 2.461 66.23 3.335 ;
      RECT 66.19 2.429 66.195 3.441 ;
      RECT 66.175 2.411 66.19 3.486 ;
      RECT 66.17 2.394 66.175 2.72 ;
      RECT 66.165 2.775 66.175 3.543 ;
      RECT 66.16 2.38 66.17 2.693 ;
      RECT 66.155 2.83 66.165 3.825 ;
      RECT 66.15 2.366 66.16 2.678 ;
      RECT 66.15 2.88 66.155 3.825 ;
      RECT 66.135 2.343 66.15 2.658 ;
      RECT 66.115 3.002 66.15 3.825 ;
      RECT 66.13 2.325 66.135 2.64 ;
      RECT 66.125 2.317 66.13 2.63 ;
      RECT 66.095 2.285 66.125 2.594 ;
      RECT 66.105 3.13 66.115 3.825 ;
      RECT 66.1 3.157 66.105 3.825 ;
      RECT 66.095 3.207 66.1 3.825 ;
      RECT 66.085 2.251 66.095 2.559 ;
      RECT 66.045 3.275 66.095 3.825 ;
      RECT 66.07 2.228 66.085 2.535 ;
      RECT 66.045 2.1 66.07 2.498 ;
      RECT 66.04 2.1 66.045 2.47 ;
      RECT 66.01 3.375 66.045 3.825 ;
      RECT 66.035 2.1 66.04 2.463 ;
      RECT 66.03 2.1 66.035 2.453 ;
      RECT 66.015 2.1 66.03 2.438 ;
      RECT 66 2.1 66.015 2.41 ;
      RECT 65.965 3.48 66.01 3.825 ;
      RECT 65.985 2.1 66 2.383 ;
      RECT 65.955 2.1 65.985 2.368 ;
      RECT 65.95 3.552 65.965 3.825 ;
      RECT 65.875 2.635 65.915 2.895 ;
      RECT 65.65 2.582 65.655 2.84 ;
      RECT 61.605 2.06 61.865 2.32 ;
      RECT 61.605 2.085 61.88 2.3 ;
      RECT 63.995 1.91 64 2.055 ;
      RECT 65.865 2.63 65.875 2.895 ;
      RECT 65.845 2.622 65.865 2.895 ;
      RECT 65.827 2.618 65.845 2.895 ;
      RECT 65.741 2.607 65.827 2.895 ;
      RECT 65.655 2.59 65.741 2.895 ;
      RECT 65.6 2.577 65.65 2.825 ;
      RECT 65.566 2.569 65.6 2.8 ;
      RECT 65.48 2.558 65.566 2.765 ;
      RECT 65.445 2.535 65.48 2.73 ;
      RECT 65.435 2.497 65.445 2.716 ;
      RECT 65.43 2.47 65.435 2.712 ;
      RECT 65.425 2.457 65.43 2.709 ;
      RECT 65.415 2.437 65.425 2.705 ;
      RECT 65.41 2.412 65.415 2.701 ;
      RECT 65.385 2.367 65.41 2.695 ;
      RECT 65.375 2.308 65.385 2.687 ;
      RECT 65.365 2.276 65.375 2.678 ;
      RECT 65.345 2.228 65.365 2.658 ;
      RECT 65.34 2.188 65.345 2.628 ;
      RECT 65.325 2.162 65.34 2.602 ;
      RECT 65.32 2.14 65.325 2.578 ;
      RECT 65.305 2.112 65.32 2.554 ;
      RECT 65.29 2.085 65.305 2.518 ;
      RECT 65.275 2.062 65.29 2.48 ;
      RECT 65.27 2.052 65.275 2.455 ;
      RECT 65.26 2.045 65.27 2.438 ;
      RECT 65.245 2.032 65.26 2.408 ;
      RECT 65.24 2.022 65.245 2.383 ;
      RECT 65.235 2.017 65.24 2.37 ;
      RECT 65.225 2.01 65.235 2.35 ;
      RECT 65.22 2.003 65.225 2.335 ;
      RECT 65.195 1.996 65.22 2.293 ;
      RECT 65.18 1.986 65.195 2.243 ;
      RECT 65.17 1.981 65.18 2.213 ;
      RECT 65.16 1.977 65.17 2.188 ;
      RECT 65.145 1.974 65.16 2.178 ;
      RECT 65.095 1.971 65.145 2.163 ;
      RECT 65.075 1.969 65.095 2.148 ;
      RECT 65.026 1.967 65.075 2.143 ;
      RECT 64.94 1.963 65.026 2.138 ;
      RECT 64.901 1.96 64.94 2.134 ;
      RECT 64.815 1.956 64.901 2.129 ;
      RECT 64.765 1.953 64.815 2.123 ;
      RECT 64.716 1.95 64.765 2.118 ;
      RECT 64.63 1.947 64.716 2.113 ;
      RECT 64.626 1.945 64.63 2.11 ;
      RECT 64.54 1.942 64.626 2.105 ;
      RECT 64.491 1.938 64.54 2.098 ;
      RECT 64.405 1.935 64.491 2.093 ;
      RECT 64.381 1.932 64.405 2.089 ;
      RECT 64.295 1.93 64.381 2.084 ;
      RECT 64.23 1.926 64.295 2.077 ;
      RECT 64.227 1.925 64.23 2.074 ;
      RECT 64.141 1.922 64.227 2.071 ;
      RECT 64.055 1.916 64.141 2.064 ;
      RECT 64.025 1.912 64.055 2.06 ;
      RECT 64 1.91 64.025 2.058 ;
      RECT 63.945 1.907 63.995 2.055 ;
      RECT 63.865 1.906 63.945 2.055 ;
      RECT 63.81 1.908 63.865 2.058 ;
      RECT 63.795 1.909 63.81 2.062 ;
      RECT 63.74 1.917 63.795 2.072 ;
      RECT 63.71 1.925 63.74 2.085 ;
      RECT 63.691 1.926 63.71 2.091 ;
      RECT 63.605 1.929 63.691 2.096 ;
      RECT 63.535 1.934 63.605 2.105 ;
      RECT 63.516 1.937 63.535 2.111 ;
      RECT 63.43 1.941 63.516 2.116 ;
      RECT 63.39 1.945 63.43 2.123 ;
      RECT 63.381 1.947 63.39 2.126 ;
      RECT 63.295 1.951 63.381 2.131 ;
      RECT 63.292 1.954 63.295 2.135 ;
      RECT 63.206 1.957 63.292 2.139 ;
      RECT 63.12 1.963 63.206 2.147 ;
      RECT 63.096 1.967 63.12 2.151 ;
      RECT 63.01 1.971 63.096 2.156 ;
      RECT 62.965 1.976 63.01 2.163 ;
      RECT 62.885 1.981 62.965 2.17 ;
      RECT 62.805 1.987 62.885 2.185 ;
      RECT 62.78 1.991 62.805 2.198 ;
      RECT 62.715 1.994 62.78 2.21 ;
      RECT 62.66 1.999 62.715 2.225 ;
      RECT 62.63 2.002 62.66 2.243 ;
      RECT 62.62 2.004 62.63 2.256 ;
      RECT 62.56 2.019 62.62 2.266 ;
      RECT 62.545 2.036 62.56 2.275 ;
      RECT 62.54 2.045 62.545 2.275 ;
      RECT 62.53 2.055 62.54 2.275 ;
      RECT 62.52 2.072 62.53 2.275 ;
      RECT 62.5 2.082 62.52 2.276 ;
      RECT 62.455 2.092 62.5 2.277 ;
      RECT 62.42 2.101 62.455 2.279 ;
      RECT 62.355 2.106 62.42 2.281 ;
      RECT 62.275 2.107 62.355 2.284 ;
      RECT 62.271 2.105 62.275 2.285 ;
      RECT 62.185 2.102 62.271 2.287 ;
      RECT 62.138 2.099 62.185 2.289 ;
      RECT 62.052 2.095 62.138 2.292 ;
      RECT 61.966 2.091 62.052 2.295 ;
      RECT 61.88 2.087 61.966 2.299 ;
      RECT 65.265 3.71 65.295 3.99 ;
      RECT 65.015 3.6 65.035 3.99 ;
      RECT 64.97 3.6 65.035 3.86 ;
      RECT 64.8 2.225 64.835 2.485 ;
      RECT 64.575 2.225 64.635 2.485 ;
      RECT 65.255 3.69 65.265 3.99 ;
      RECT 65.25 3.65 65.255 3.99 ;
      RECT 65.235 3.605 65.25 3.99 ;
      RECT 65.23 3.57 65.235 3.99 ;
      RECT 65.225 3.55 65.23 3.99 ;
      RECT 65.195 3.477 65.225 3.99 ;
      RECT 65.175 3.375 65.195 3.99 ;
      RECT 65.165 3.305 65.175 3.99 ;
      RECT 65.12 3.245 65.165 3.99 ;
      RECT 65.035 3.206 65.12 3.99 ;
      RECT 65.03 3.197 65.035 3.57 ;
      RECT 65.02 3.196 65.03 3.553 ;
      RECT 64.995 3.177 65.02 3.523 ;
      RECT 64.99 3.152 64.995 3.502 ;
      RECT 64.98 3.13 64.99 3.493 ;
      RECT 64.975 3.101 64.98 3.483 ;
      RECT 64.935 3.027 64.975 3.455 ;
      RECT 64.915 2.928 64.935 3.42 ;
      RECT 64.9 2.864 64.915 3.403 ;
      RECT 64.87 2.788 64.9 3.375 ;
      RECT 64.85 2.703 64.87 3.348 ;
      RECT 64.81 2.599 64.85 3.255 ;
      RECT 64.805 2.52 64.81 3.163 ;
      RECT 64.8 2.503 64.805 3.14 ;
      RECT 64.795 2.225 64.8 3.12 ;
      RECT 64.765 2.225 64.795 3.058 ;
      RECT 64.76 2.225 64.765 2.99 ;
      RECT 64.75 2.225 64.76 2.955 ;
      RECT 64.74 2.225 64.75 2.92 ;
      RECT 64.675 2.225 64.74 2.775 ;
      RECT 64.67 2.225 64.675 2.645 ;
      RECT 64.64 2.225 64.67 2.578 ;
      RECT 64.635 2.225 64.64 2.503 ;
      RECT 63.815 3.15 64.095 3.43 ;
      RECT 63.855 3.13 64.115 3.39 ;
      RECT 63.845 3.14 64.115 3.39 ;
      RECT 63.855 3.067 64.07 3.43 ;
      RECT 63.91 2.99 64.065 3.43 ;
      RECT 63.915 2.775 64.065 3.43 ;
      RECT 63.905 2.577 64.055 2.828 ;
      RECT 63.895 2.577 64.055 2.695 ;
      RECT 63.89 2.455 64.05 2.598 ;
      RECT 63.875 2.455 64.05 2.503 ;
      RECT 63.87 2.165 64.045 2.48 ;
      RECT 63.855 2.165 64.045 2.45 ;
      RECT 63.815 2.165 64.075 2.425 ;
      RECT 63.725 3.635 63.805 3.895 ;
      RECT 63.13 2.355 63.135 2.62 ;
      RECT 63.01 2.355 63.135 2.615 ;
      RECT 63.685 3.6 63.725 3.895 ;
      RECT 63.64 3.522 63.685 3.895 ;
      RECT 63.62 3.45 63.64 3.895 ;
      RECT 63.61 3.402 63.62 3.895 ;
      RECT 63.575 3.335 63.61 3.895 ;
      RECT 63.545 3.235 63.575 3.895 ;
      RECT 63.525 3.16 63.545 3.695 ;
      RECT 63.515 3.11 63.525 3.65 ;
      RECT 63.51 3.087 63.515 3.623 ;
      RECT 63.505 3.072 63.51 3.61 ;
      RECT 63.5 3.057 63.505 3.588 ;
      RECT 63.495 3.042 63.5 3.57 ;
      RECT 63.47 2.997 63.495 3.525 ;
      RECT 63.46 2.945 63.47 3.468 ;
      RECT 63.45 2.915 63.46 3.435 ;
      RECT 63.44 2.88 63.45 3.403 ;
      RECT 63.405 2.812 63.44 3.335 ;
      RECT 63.4 2.751 63.405 3.27 ;
      RECT 63.39 2.739 63.4 3.25 ;
      RECT 63.385 2.727 63.39 3.23 ;
      RECT 63.38 2.719 63.385 3.218 ;
      RECT 63.375 2.711 63.38 3.198 ;
      RECT 63.365 2.699 63.375 3.17 ;
      RECT 63.355 2.683 63.365 3.14 ;
      RECT 63.33 2.655 63.355 3.078 ;
      RECT 63.32 2.626 63.33 3.023 ;
      RECT 63.305 2.605 63.32 2.983 ;
      RECT 63.3 2.589 63.305 2.955 ;
      RECT 63.295 2.577 63.3 2.945 ;
      RECT 63.29 2.572 63.295 2.918 ;
      RECT 63.285 2.565 63.29 2.905 ;
      RECT 63.27 2.548 63.285 2.878 ;
      RECT 63.26 2.355 63.27 2.838 ;
      RECT 63.25 2.355 63.26 2.805 ;
      RECT 63.24 2.355 63.25 2.78 ;
      RECT 63.17 2.355 63.24 2.715 ;
      RECT 63.16 2.355 63.17 2.663 ;
      RECT 63.145 2.355 63.16 2.645 ;
      RECT 63.135 2.355 63.145 2.63 ;
      RECT 62.965 3.225 63.225 3.485 ;
      RECT 61.5 3.26 61.505 3.467 ;
      RECT 61.135 3.15 61.21 3.465 ;
      RECT 60.95 3.205 61.105 3.465 ;
      RECT 61.135 3.15 61.24 3.43 ;
      RECT 62.95 3.322 62.965 3.483 ;
      RECT 62.925 3.33 62.95 3.488 ;
      RECT 62.9 3.337 62.925 3.493 ;
      RECT 62.837 3.348 62.9 3.502 ;
      RECT 62.751 3.367 62.837 3.519 ;
      RECT 62.665 3.389 62.751 3.538 ;
      RECT 62.65 3.402 62.665 3.549 ;
      RECT 62.61 3.41 62.65 3.556 ;
      RECT 62.59 3.415 62.61 3.563 ;
      RECT 62.552 3.416 62.59 3.566 ;
      RECT 62.466 3.419 62.552 3.567 ;
      RECT 62.38 3.423 62.466 3.568 ;
      RECT 62.331 3.425 62.38 3.57 ;
      RECT 62.245 3.425 62.331 3.572 ;
      RECT 62.205 3.42 62.245 3.574 ;
      RECT 62.195 3.414 62.205 3.575 ;
      RECT 62.155 3.409 62.195 3.572 ;
      RECT 62.145 3.402 62.155 3.568 ;
      RECT 62.13 3.398 62.145 3.566 ;
      RECT 62.113 3.394 62.13 3.564 ;
      RECT 62.027 3.384 62.113 3.556 ;
      RECT 61.941 3.366 62.027 3.542 ;
      RECT 61.855 3.349 61.941 3.528 ;
      RECT 61.83 3.337 61.855 3.519 ;
      RECT 61.76 3.327 61.83 3.512 ;
      RECT 61.715 3.315 61.76 3.503 ;
      RECT 61.655 3.302 61.715 3.495 ;
      RECT 61.65 3.294 61.655 3.49 ;
      RECT 61.615 3.289 61.65 3.488 ;
      RECT 61.56 3.28 61.615 3.481 ;
      RECT 61.52 3.269 61.56 3.473 ;
      RECT 61.505 3.262 61.52 3.469 ;
      RECT 61.485 3.255 61.5 3.466 ;
      RECT 61.47 3.245 61.485 3.464 ;
      RECT 61.455 3.232 61.47 3.461 ;
      RECT 61.43 3.215 61.455 3.457 ;
      RECT 61.415 3.197 61.43 3.454 ;
      RECT 61.39 3.15 61.415 3.452 ;
      RECT 61.366 3.15 61.39 3.449 ;
      RECT 61.28 3.15 61.366 3.441 ;
      RECT 61.24 3.15 61.28 3.433 ;
      RECT 61.105 3.197 61.135 3.465 ;
      RECT 62.785 2.78 63.045 3.04 ;
      RECT 62.745 2.78 63.045 2.918 ;
      RECT 62.71 2.78 63.045 2.903 ;
      RECT 62.655 2.78 63.045 2.883 ;
      RECT 62.575 2.59 62.855 2.87 ;
      RECT 62.575 2.772 62.925 2.87 ;
      RECT 62.575 2.715 62.91 2.87 ;
      RECT 62.575 2.662 62.86 2.87 ;
      RECT 60.405 2.59 60.6 3.375 ;
      RECT 60.485 1.205 60.6 3.375 ;
      RECT 60.34 3.115 60.4 3.375 ;
      RECT 61.71 2.635 61.97 2.895 ;
      RECT 60.395 2.59 60.6 2.87 ;
      RECT 61.705 2.645 61.97 2.83 ;
      RECT 61.42 2.62 61.43 2.77 ;
      RECT 60.655 1.205 60.735 1.55 ;
      RECT 60.39 1.205 60.6 1.55 ;
      RECT 61.695 2.645 61.705 2.829 ;
      RECT 61.685 2.644 61.695 2.826 ;
      RECT 61.676 2.643 61.685 2.824 ;
      RECT 61.59 2.639 61.676 2.814 ;
      RECT 61.516 2.631 61.59 2.796 ;
      RECT 61.43 2.624 61.516 2.779 ;
      RECT 61.37 2.62 61.42 2.769 ;
      RECT 61.335 2.619 61.37 2.766 ;
      RECT 61.28 2.619 61.335 2.768 ;
      RECT 61.245 2.619 61.28 2.772 ;
      RECT 61.159 2.618 61.245 2.779 ;
      RECT 61.073 2.617 61.159 2.789 ;
      RECT 60.987 2.616 61.073 2.8 ;
      RECT 60.901 2.616 60.987 2.81 ;
      RECT 60.815 2.615 60.901 2.82 ;
      RECT 60.78 2.615 60.815 2.86 ;
      RECT 60.775 2.615 60.78 2.903 ;
      RECT 60.75 2.615 60.775 2.92 ;
      RECT 60.675 2.615 60.75 2.935 ;
      RECT 60.655 2.59 60.675 2.948 ;
      RECT 60.65 1.205 60.655 2.958 ;
      RECT 60.625 1.205 60.65 3 ;
      RECT 60.6 1.205 60.625 3.078 ;
      RECT 60.4 2.997 60.405 3.375 ;
      RECT 59.735 2.949 59.75 3.405 ;
      RECT 59.73 3.021 59.836 3.403 ;
      RECT 59.75 2.115 59.885 3.401 ;
      RECT 59.735 2.965 59.89 3.4 ;
      RECT 59.735 3.015 59.895 3.398 ;
      RECT 59.72 3.08 59.895 3.397 ;
      RECT 59.73 3.072 59.9 3.394 ;
      RECT 59.71 3.12 59.9 3.389 ;
      RECT 59.71 3.12 59.915 3.386 ;
      RECT 59.705 3.12 59.915 3.383 ;
      RECT 59.68 3.12 59.94 3.38 ;
      RECT 59.75 2.115 59.91 2.768 ;
      RECT 59.745 2.115 59.91 2.74 ;
      RECT 59.74 2.115 59.91 2.568 ;
      RECT 59.74 2.115 59.93 2.508 ;
      RECT 59.695 2.115 59.955 2.375 ;
      RECT 59.175 2.59 59.455 2.87 ;
      RECT 59.165 2.605 59.455 2.865 ;
      RECT 59.12 2.667 59.455 2.863 ;
      RECT 59.195 2.582 59.36 2.87 ;
      RECT 59.195 2.567 59.316 2.87 ;
      RECT 59.23 2.56 59.316 2.87 ;
      RECT 58.695 3.71 58.975 3.99 ;
      RECT 58.655 3.672 58.95 3.783 ;
      RECT 58.64 3.622 58.93 3.678 ;
      RECT 58.585 3.385 58.845 3.645 ;
      RECT 58.585 3.587 58.925 3.645 ;
      RECT 58.585 3.527 58.92 3.645 ;
      RECT 58.585 3.477 58.9 3.645 ;
      RECT 58.585 3.457 58.895 3.645 ;
      RECT 58.585 3.435 58.89 3.645 ;
      RECT 58.585 3.42 58.86 3.645 ;
      RECT 54.315 6.225 54.635 6.545 ;
      RECT 54.345 5.695 54.515 6.545 ;
      RECT 54.345 5.695 54.52 6.045 ;
      RECT 54.345 5.695 55.32 5.87 ;
      RECT 55.145 1.965 55.32 5.87 ;
      RECT 55.09 1.965 55.44 2.315 ;
      RECT 55.115 6.655 55.44 6.98 ;
      RECT 54 6.745 55.44 6.915 ;
      RECT 54 2.395 54.16 6.915 ;
      RECT 54.315 2.365 54.635 2.685 ;
      RECT 54 2.395 54.635 2.565 ;
      RECT 52.67 1.14 53.045 1.51 ;
      RECT 44.59 0.96 44.965 1.33 ;
      RECT 43.155 0.96 43.53 1.33 ;
      RECT 43.155 1.08 52.975 1.25 ;
      RECT 49.1 4.36 52.955 4.53 ;
      RECT 52.785 3.425 52.955 4.53 ;
      RECT 49.1 3.67 49.27 4.53 ;
      RECT 49.05 3.71 49.33 3.99 ;
      RECT 49.07 3.67 49.33 3.99 ;
      RECT 48.71 3.625 48.815 3.885 ;
      RECT 52.695 3.43 53.045 3.78 ;
      RECT 48.565 2.115 48.655 2.375 ;
      RECT 49.105 3.18 49.11 3.22 ;
      RECT 49.1 3.17 49.105 3.305 ;
      RECT 49.095 3.16 49.1 3.398 ;
      RECT 49.085 3.14 49.095 3.454 ;
      RECT 49.005 3.068 49.085 3.534 ;
      RECT 49.04 3.712 49.05 3.937 ;
      RECT 49.035 3.709 49.04 3.932 ;
      RECT 49.02 3.706 49.035 3.925 ;
      RECT 48.985 3.7 49.02 3.907 ;
      RECT 49 3.003 49.005 3.608 ;
      RECT 48.98 2.954 49 3.623 ;
      RECT 48.97 3.687 48.985 3.89 ;
      RECT 48.975 2.896 48.98 3.638 ;
      RECT 48.97 2.874 48.975 3.648 ;
      RECT 48.935 2.784 48.97 3.885 ;
      RECT 48.92 2.662 48.935 3.885 ;
      RECT 48.915 2.615 48.92 3.885 ;
      RECT 48.89 2.54 48.915 3.885 ;
      RECT 48.875 2.455 48.89 3.885 ;
      RECT 48.87 2.402 48.875 3.885 ;
      RECT 48.865 2.382 48.87 3.885 ;
      RECT 48.86 2.357 48.865 3.119 ;
      RECT 48.845 3.317 48.865 3.885 ;
      RECT 48.855 2.335 48.86 3.096 ;
      RECT 48.845 2.287 48.855 3.061 ;
      RECT 48.84 2.25 48.845 3.027 ;
      RECT 48.84 3.397 48.845 3.885 ;
      RECT 48.825 2.227 48.84 2.982 ;
      RECT 48.82 3.495 48.84 3.885 ;
      RECT 48.77 2.115 48.825 2.824 ;
      RECT 48.815 3.617 48.82 3.885 ;
      RECT 48.755 2.115 48.77 2.663 ;
      RECT 48.75 2.115 48.755 2.615 ;
      RECT 48.745 2.115 48.75 2.603 ;
      RECT 48.7 2.115 48.745 2.54 ;
      RECT 48.675 2.115 48.7 2.458 ;
      RECT 48.66 2.115 48.675 2.41 ;
      RECT 48.655 2.115 48.66 2.38 ;
      RECT 51.045 2.16 51.305 2.42 ;
      RECT 51.04 2.16 51.305 2.368 ;
      RECT 51.035 2.16 51.305 2.338 ;
      RECT 51.01 2.03 51.29 2.31 ;
      RECT 39.57 6.66 39.92 7.01 ;
      RECT 50.545 6.615 50.895 6.965 ;
      RECT 39.57 6.69 50.895 6.89 ;
      RECT 50.05 3.71 50.33 3.99 ;
      RECT 50.09 3.665 50.355 3.925 ;
      RECT 50.08 3.7 50.355 3.925 ;
      RECT 50.085 3.685 50.33 3.99 ;
      RECT 50.09 3.662 50.3 3.99 ;
      RECT 50.09 3.66 50.285 3.99 ;
      RECT 50.13 3.65 50.285 3.99 ;
      RECT 50.1 3.655 50.285 3.99 ;
      RECT 50.13 3.647 50.23 3.99 ;
      RECT 50.155 3.64 50.23 3.99 ;
      RECT 50.135 3.642 50.23 3.99 ;
      RECT 49.465 3.155 49.725 3.415 ;
      RECT 49.515 3.147 49.705 3.415 ;
      RECT 49.52 3.067 49.705 3.415 ;
      RECT 49.64 2.455 49.705 3.415 ;
      RECT 49.545 2.852 49.705 3.415 ;
      RECT 49.62 2.54 49.705 3.415 ;
      RECT 49.655 2.165 49.791 2.893 ;
      RECT 49.6 2.662 49.791 2.893 ;
      RECT 49.615 2.602 49.705 3.415 ;
      RECT 49.655 2.165 49.815 2.558 ;
      RECT 49.655 2.165 49.825 2.455 ;
      RECT 49.645 2.165 49.905 2.425 ;
      RECT 47.98 3.565 48.025 3.825 ;
      RECT 47.885 2.1 48.03 2.36 ;
      RECT 48.39 2.722 48.4 2.813 ;
      RECT 48.375 2.66 48.39 2.869 ;
      RECT 48.37 2.607 48.375 2.915 ;
      RECT 48.32 2.554 48.37 3.041 ;
      RECT 48.315 2.509 48.32 3.188 ;
      RECT 48.305 2.497 48.315 3.23 ;
      RECT 48.27 2.461 48.305 3.335 ;
      RECT 48.265 2.429 48.27 3.441 ;
      RECT 48.25 2.411 48.265 3.486 ;
      RECT 48.245 2.394 48.25 2.72 ;
      RECT 48.24 2.775 48.25 3.543 ;
      RECT 48.235 2.38 48.245 2.693 ;
      RECT 48.23 2.83 48.24 3.825 ;
      RECT 48.225 2.366 48.235 2.678 ;
      RECT 48.225 2.88 48.23 3.825 ;
      RECT 48.21 2.343 48.225 2.658 ;
      RECT 48.19 3.002 48.225 3.825 ;
      RECT 48.205 2.325 48.21 2.64 ;
      RECT 48.2 2.317 48.205 2.63 ;
      RECT 48.17 2.285 48.2 2.594 ;
      RECT 48.18 3.13 48.19 3.825 ;
      RECT 48.175 3.157 48.18 3.825 ;
      RECT 48.17 3.207 48.175 3.825 ;
      RECT 48.16 2.251 48.17 2.559 ;
      RECT 48.12 3.275 48.17 3.825 ;
      RECT 48.145 2.228 48.16 2.535 ;
      RECT 48.12 2.1 48.145 2.498 ;
      RECT 48.115 2.1 48.12 2.47 ;
      RECT 48.085 3.375 48.12 3.825 ;
      RECT 48.11 2.1 48.115 2.463 ;
      RECT 48.105 2.1 48.11 2.453 ;
      RECT 48.09 2.1 48.105 2.438 ;
      RECT 48.075 2.1 48.09 2.41 ;
      RECT 48.04 3.48 48.085 3.825 ;
      RECT 48.06 2.1 48.075 2.383 ;
      RECT 48.03 2.1 48.06 2.368 ;
      RECT 48.025 3.552 48.04 3.825 ;
      RECT 47.95 2.635 47.99 2.895 ;
      RECT 47.725 2.582 47.73 2.84 ;
      RECT 43.68 2.06 43.94 2.32 ;
      RECT 43.68 2.085 43.955 2.3 ;
      RECT 46.07 1.91 46.075 2.055 ;
      RECT 47.94 2.63 47.95 2.895 ;
      RECT 47.92 2.622 47.94 2.895 ;
      RECT 47.902 2.618 47.92 2.895 ;
      RECT 47.816 2.607 47.902 2.895 ;
      RECT 47.73 2.59 47.816 2.895 ;
      RECT 47.675 2.577 47.725 2.825 ;
      RECT 47.641 2.569 47.675 2.8 ;
      RECT 47.555 2.558 47.641 2.765 ;
      RECT 47.52 2.535 47.555 2.73 ;
      RECT 47.51 2.497 47.52 2.716 ;
      RECT 47.505 2.47 47.51 2.712 ;
      RECT 47.5 2.457 47.505 2.709 ;
      RECT 47.49 2.437 47.5 2.705 ;
      RECT 47.485 2.412 47.49 2.701 ;
      RECT 47.46 2.367 47.485 2.695 ;
      RECT 47.45 2.308 47.46 2.687 ;
      RECT 47.44 2.276 47.45 2.678 ;
      RECT 47.42 2.228 47.44 2.658 ;
      RECT 47.415 2.188 47.42 2.628 ;
      RECT 47.4 2.162 47.415 2.602 ;
      RECT 47.395 2.14 47.4 2.578 ;
      RECT 47.38 2.112 47.395 2.554 ;
      RECT 47.365 2.085 47.38 2.518 ;
      RECT 47.35 2.062 47.365 2.48 ;
      RECT 47.345 2.052 47.35 2.455 ;
      RECT 47.335 2.045 47.345 2.438 ;
      RECT 47.32 2.032 47.335 2.408 ;
      RECT 47.315 2.022 47.32 2.383 ;
      RECT 47.31 2.017 47.315 2.37 ;
      RECT 47.3 2.01 47.31 2.35 ;
      RECT 47.295 2.003 47.3 2.335 ;
      RECT 47.27 1.996 47.295 2.293 ;
      RECT 47.255 1.986 47.27 2.243 ;
      RECT 47.245 1.981 47.255 2.213 ;
      RECT 47.235 1.977 47.245 2.188 ;
      RECT 47.22 1.974 47.235 2.178 ;
      RECT 47.17 1.971 47.22 2.163 ;
      RECT 47.15 1.969 47.17 2.148 ;
      RECT 47.101 1.967 47.15 2.143 ;
      RECT 47.015 1.963 47.101 2.138 ;
      RECT 46.976 1.96 47.015 2.134 ;
      RECT 46.89 1.956 46.976 2.129 ;
      RECT 46.84 1.953 46.89 2.123 ;
      RECT 46.791 1.95 46.84 2.118 ;
      RECT 46.705 1.947 46.791 2.113 ;
      RECT 46.701 1.945 46.705 2.11 ;
      RECT 46.615 1.942 46.701 2.105 ;
      RECT 46.566 1.938 46.615 2.098 ;
      RECT 46.48 1.935 46.566 2.093 ;
      RECT 46.456 1.932 46.48 2.089 ;
      RECT 46.37 1.93 46.456 2.084 ;
      RECT 46.305 1.926 46.37 2.077 ;
      RECT 46.302 1.925 46.305 2.074 ;
      RECT 46.216 1.922 46.302 2.071 ;
      RECT 46.13 1.916 46.216 2.064 ;
      RECT 46.1 1.912 46.13 2.06 ;
      RECT 46.075 1.91 46.1 2.058 ;
      RECT 46.02 1.907 46.07 2.055 ;
      RECT 45.94 1.906 46.02 2.055 ;
      RECT 45.885 1.908 45.94 2.058 ;
      RECT 45.87 1.909 45.885 2.062 ;
      RECT 45.815 1.917 45.87 2.072 ;
      RECT 45.785 1.925 45.815 2.085 ;
      RECT 45.766 1.926 45.785 2.091 ;
      RECT 45.68 1.929 45.766 2.096 ;
      RECT 45.61 1.934 45.68 2.105 ;
      RECT 45.591 1.937 45.61 2.111 ;
      RECT 45.505 1.941 45.591 2.116 ;
      RECT 45.465 1.945 45.505 2.123 ;
      RECT 45.456 1.947 45.465 2.126 ;
      RECT 45.37 1.951 45.456 2.131 ;
      RECT 45.367 1.954 45.37 2.135 ;
      RECT 45.281 1.957 45.367 2.139 ;
      RECT 45.195 1.963 45.281 2.147 ;
      RECT 45.171 1.967 45.195 2.151 ;
      RECT 45.085 1.971 45.171 2.156 ;
      RECT 45.04 1.976 45.085 2.163 ;
      RECT 44.96 1.981 45.04 2.17 ;
      RECT 44.88 1.987 44.96 2.185 ;
      RECT 44.855 1.991 44.88 2.198 ;
      RECT 44.79 1.994 44.855 2.21 ;
      RECT 44.735 1.999 44.79 2.225 ;
      RECT 44.705 2.002 44.735 2.243 ;
      RECT 44.695 2.004 44.705 2.256 ;
      RECT 44.635 2.019 44.695 2.266 ;
      RECT 44.62 2.036 44.635 2.275 ;
      RECT 44.615 2.045 44.62 2.275 ;
      RECT 44.605 2.055 44.615 2.275 ;
      RECT 44.595 2.072 44.605 2.275 ;
      RECT 44.575 2.082 44.595 2.276 ;
      RECT 44.53 2.092 44.575 2.277 ;
      RECT 44.495 2.101 44.53 2.279 ;
      RECT 44.43 2.106 44.495 2.281 ;
      RECT 44.35 2.107 44.43 2.284 ;
      RECT 44.346 2.105 44.35 2.285 ;
      RECT 44.26 2.102 44.346 2.287 ;
      RECT 44.213 2.099 44.26 2.289 ;
      RECT 44.127 2.095 44.213 2.292 ;
      RECT 44.041 2.091 44.127 2.295 ;
      RECT 43.955 2.087 44.041 2.299 ;
      RECT 47.34 3.71 47.37 3.99 ;
      RECT 47.09 3.6 47.11 3.99 ;
      RECT 47.045 3.6 47.11 3.86 ;
      RECT 46.875 2.225 46.91 2.485 ;
      RECT 46.65 2.225 46.71 2.485 ;
      RECT 47.33 3.69 47.34 3.99 ;
      RECT 47.325 3.65 47.33 3.99 ;
      RECT 47.31 3.605 47.325 3.99 ;
      RECT 47.305 3.57 47.31 3.99 ;
      RECT 47.3 3.55 47.305 3.99 ;
      RECT 47.27 3.477 47.3 3.99 ;
      RECT 47.25 3.375 47.27 3.99 ;
      RECT 47.24 3.305 47.25 3.99 ;
      RECT 47.195 3.245 47.24 3.99 ;
      RECT 47.11 3.206 47.195 3.99 ;
      RECT 47.105 3.197 47.11 3.57 ;
      RECT 47.095 3.196 47.105 3.553 ;
      RECT 47.07 3.177 47.095 3.523 ;
      RECT 47.065 3.152 47.07 3.502 ;
      RECT 47.055 3.13 47.065 3.493 ;
      RECT 47.05 3.101 47.055 3.483 ;
      RECT 47.01 3.027 47.05 3.455 ;
      RECT 46.99 2.928 47.01 3.42 ;
      RECT 46.975 2.864 46.99 3.403 ;
      RECT 46.945 2.788 46.975 3.375 ;
      RECT 46.925 2.703 46.945 3.348 ;
      RECT 46.885 2.599 46.925 3.255 ;
      RECT 46.88 2.52 46.885 3.163 ;
      RECT 46.875 2.503 46.88 3.14 ;
      RECT 46.87 2.225 46.875 3.12 ;
      RECT 46.84 2.225 46.87 3.058 ;
      RECT 46.835 2.225 46.84 2.99 ;
      RECT 46.825 2.225 46.835 2.955 ;
      RECT 46.815 2.225 46.825 2.92 ;
      RECT 46.75 2.225 46.815 2.775 ;
      RECT 46.745 2.225 46.75 2.645 ;
      RECT 46.715 2.225 46.745 2.578 ;
      RECT 46.71 2.225 46.715 2.503 ;
      RECT 45.89 3.15 46.17 3.43 ;
      RECT 45.93 3.13 46.19 3.39 ;
      RECT 45.92 3.14 46.19 3.39 ;
      RECT 45.93 3.067 46.145 3.43 ;
      RECT 45.985 2.99 46.14 3.43 ;
      RECT 45.99 2.775 46.14 3.43 ;
      RECT 45.98 2.577 46.13 2.828 ;
      RECT 45.97 2.577 46.13 2.695 ;
      RECT 45.965 2.455 46.125 2.598 ;
      RECT 45.95 2.455 46.125 2.503 ;
      RECT 45.945 2.165 46.12 2.48 ;
      RECT 45.93 2.165 46.12 2.45 ;
      RECT 45.89 2.165 46.15 2.425 ;
      RECT 45.8 3.635 45.88 3.895 ;
      RECT 45.205 2.355 45.21 2.62 ;
      RECT 45.085 2.355 45.21 2.615 ;
      RECT 45.76 3.6 45.8 3.895 ;
      RECT 45.715 3.522 45.76 3.895 ;
      RECT 45.695 3.45 45.715 3.895 ;
      RECT 45.685 3.402 45.695 3.895 ;
      RECT 45.65 3.335 45.685 3.895 ;
      RECT 45.62 3.235 45.65 3.895 ;
      RECT 45.6 3.16 45.62 3.695 ;
      RECT 45.59 3.11 45.6 3.65 ;
      RECT 45.585 3.087 45.59 3.623 ;
      RECT 45.58 3.072 45.585 3.61 ;
      RECT 45.575 3.057 45.58 3.588 ;
      RECT 45.57 3.042 45.575 3.57 ;
      RECT 45.545 2.997 45.57 3.525 ;
      RECT 45.535 2.945 45.545 3.468 ;
      RECT 45.525 2.915 45.535 3.435 ;
      RECT 45.515 2.88 45.525 3.403 ;
      RECT 45.48 2.812 45.515 3.335 ;
      RECT 45.475 2.751 45.48 3.27 ;
      RECT 45.465 2.739 45.475 3.25 ;
      RECT 45.46 2.727 45.465 3.23 ;
      RECT 45.455 2.719 45.46 3.218 ;
      RECT 45.45 2.711 45.455 3.198 ;
      RECT 45.44 2.699 45.45 3.17 ;
      RECT 45.43 2.683 45.44 3.14 ;
      RECT 45.405 2.655 45.43 3.078 ;
      RECT 45.395 2.626 45.405 3.023 ;
      RECT 45.38 2.605 45.395 2.983 ;
      RECT 45.375 2.589 45.38 2.955 ;
      RECT 45.37 2.577 45.375 2.945 ;
      RECT 45.365 2.572 45.37 2.918 ;
      RECT 45.36 2.565 45.365 2.905 ;
      RECT 45.345 2.548 45.36 2.878 ;
      RECT 45.335 2.355 45.345 2.838 ;
      RECT 45.325 2.355 45.335 2.805 ;
      RECT 45.315 2.355 45.325 2.78 ;
      RECT 45.245 2.355 45.315 2.715 ;
      RECT 45.235 2.355 45.245 2.663 ;
      RECT 45.22 2.355 45.235 2.645 ;
      RECT 45.21 2.355 45.22 2.63 ;
      RECT 45.04 3.225 45.3 3.485 ;
      RECT 43.575 3.26 43.58 3.467 ;
      RECT 43.21 3.15 43.285 3.465 ;
      RECT 43.025 3.205 43.18 3.465 ;
      RECT 43.21 3.15 43.315 3.43 ;
      RECT 45.025 3.322 45.04 3.483 ;
      RECT 45 3.33 45.025 3.488 ;
      RECT 44.975 3.337 45 3.493 ;
      RECT 44.912 3.348 44.975 3.502 ;
      RECT 44.826 3.367 44.912 3.519 ;
      RECT 44.74 3.389 44.826 3.538 ;
      RECT 44.725 3.402 44.74 3.549 ;
      RECT 44.685 3.41 44.725 3.556 ;
      RECT 44.665 3.415 44.685 3.563 ;
      RECT 44.627 3.416 44.665 3.566 ;
      RECT 44.541 3.419 44.627 3.567 ;
      RECT 44.455 3.423 44.541 3.568 ;
      RECT 44.406 3.425 44.455 3.57 ;
      RECT 44.32 3.425 44.406 3.572 ;
      RECT 44.28 3.42 44.32 3.574 ;
      RECT 44.27 3.414 44.28 3.575 ;
      RECT 44.23 3.409 44.27 3.572 ;
      RECT 44.22 3.402 44.23 3.568 ;
      RECT 44.205 3.398 44.22 3.566 ;
      RECT 44.188 3.394 44.205 3.564 ;
      RECT 44.102 3.384 44.188 3.556 ;
      RECT 44.016 3.366 44.102 3.542 ;
      RECT 43.93 3.349 44.016 3.528 ;
      RECT 43.905 3.337 43.93 3.519 ;
      RECT 43.835 3.327 43.905 3.512 ;
      RECT 43.79 3.315 43.835 3.503 ;
      RECT 43.73 3.302 43.79 3.495 ;
      RECT 43.725 3.294 43.73 3.49 ;
      RECT 43.69 3.289 43.725 3.488 ;
      RECT 43.635 3.28 43.69 3.481 ;
      RECT 43.595 3.269 43.635 3.473 ;
      RECT 43.58 3.262 43.595 3.469 ;
      RECT 43.56 3.255 43.575 3.466 ;
      RECT 43.545 3.245 43.56 3.464 ;
      RECT 43.53 3.232 43.545 3.461 ;
      RECT 43.505 3.215 43.53 3.457 ;
      RECT 43.49 3.197 43.505 3.454 ;
      RECT 43.465 3.15 43.49 3.452 ;
      RECT 43.441 3.15 43.465 3.449 ;
      RECT 43.355 3.15 43.441 3.441 ;
      RECT 43.315 3.15 43.355 3.433 ;
      RECT 43.18 3.197 43.21 3.465 ;
      RECT 44.86 2.78 45.12 3.04 ;
      RECT 44.82 2.78 45.12 2.918 ;
      RECT 44.785 2.78 45.12 2.903 ;
      RECT 44.73 2.78 45.12 2.883 ;
      RECT 44.65 2.59 44.93 2.87 ;
      RECT 44.65 2.772 45 2.87 ;
      RECT 44.65 2.715 44.985 2.87 ;
      RECT 44.65 2.662 44.935 2.87 ;
      RECT 42.48 2.59 42.675 3.375 ;
      RECT 42.56 1.205 42.675 3.375 ;
      RECT 42.415 3.115 42.475 3.375 ;
      RECT 43.785 2.635 44.045 2.895 ;
      RECT 42.47 2.59 42.675 2.87 ;
      RECT 43.78 2.645 44.045 2.83 ;
      RECT 43.495 2.62 43.505 2.77 ;
      RECT 42.73 1.205 42.81 1.55 ;
      RECT 42.465 1.205 42.675 1.55 ;
      RECT 43.77 2.645 43.78 2.829 ;
      RECT 43.76 2.644 43.77 2.826 ;
      RECT 43.751 2.643 43.76 2.824 ;
      RECT 43.665 2.639 43.751 2.814 ;
      RECT 43.591 2.631 43.665 2.796 ;
      RECT 43.505 2.624 43.591 2.779 ;
      RECT 43.445 2.62 43.495 2.769 ;
      RECT 43.41 2.619 43.445 2.766 ;
      RECT 43.355 2.619 43.41 2.768 ;
      RECT 43.32 2.619 43.355 2.772 ;
      RECT 43.234 2.618 43.32 2.779 ;
      RECT 43.148 2.617 43.234 2.789 ;
      RECT 43.062 2.616 43.148 2.8 ;
      RECT 42.976 2.616 43.062 2.81 ;
      RECT 42.89 2.615 42.976 2.82 ;
      RECT 42.855 2.615 42.89 2.86 ;
      RECT 42.85 2.615 42.855 2.903 ;
      RECT 42.825 2.615 42.85 2.92 ;
      RECT 42.75 2.615 42.825 2.935 ;
      RECT 42.73 2.59 42.75 2.948 ;
      RECT 42.725 1.205 42.73 2.958 ;
      RECT 42.7 1.205 42.725 3 ;
      RECT 42.675 1.205 42.7 3.078 ;
      RECT 42.475 2.997 42.48 3.375 ;
      RECT 41.81 2.949 41.825 3.405 ;
      RECT 41.805 3.021 41.911 3.403 ;
      RECT 41.825 2.115 41.96 3.401 ;
      RECT 41.81 2.965 41.965 3.4 ;
      RECT 41.81 3.015 41.97 3.398 ;
      RECT 41.795 3.08 41.97 3.397 ;
      RECT 41.805 3.072 41.975 3.394 ;
      RECT 41.785 3.12 41.975 3.389 ;
      RECT 41.785 3.12 41.99 3.386 ;
      RECT 41.78 3.12 41.99 3.383 ;
      RECT 41.755 3.12 42.015 3.38 ;
      RECT 41.825 2.115 41.985 2.768 ;
      RECT 41.82 2.115 41.985 2.74 ;
      RECT 41.815 2.115 41.985 2.568 ;
      RECT 41.815 2.115 42.005 2.508 ;
      RECT 41.77 2.115 42.03 2.375 ;
      RECT 41.25 2.59 41.53 2.87 ;
      RECT 41.24 2.605 41.53 2.865 ;
      RECT 41.195 2.667 41.53 2.863 ;
      RECT 41.27 2.582 41.435 2.87 ;
      RECT 41.27 2.567 41.391 2.87 ;
      RECT 41.305 2.56 41.391 2.87 ;
      RECT 40.77 3.71 41.05 3.99 ;
      RECT 40.73 3.672 41.025 3.783 ;
      RECT 40.715 3.622 41.005 3.678 ;
      RECT 40.66 3.385 40.92 3.645 ;
      RECT 40.66 3.587 41 3.645 ;
      RECT 40.66 3.527 40.995 3.645 ;
      RECT 40.66 3.477 40.975 3.645 ;
      RECT 40.66 3.457 40.97 3.645 ;
      RECT 40.66 3.435 40.965 3.645 ;
      RECT 40.66 3.42 40.935 3.645 ;
      RECT 36.39 6.225 36.71 6.545 ;
      RECT 36.42 5.695 36.59 6.545 ;
      RECT 36.42 5.695 36.595 6.045 ;
      RECT 36.42 5.695 37.395 5.87 ;
      RECT 37.22 1.965 37.395 5.87 ;
      RECT 37.165 1.965 37.515 2.315 ;
      RECT 37.19 6.655 37.515 6.98 ;
      RECT 36.075 6.745 37.515 6.915 ;
      RECT 36.075 2.395 36.235 6.915 ;
      RECT 36.39 2.365 36.71 2.685 ;
      RECT 36.075 2.395 36.71 2.565 ;
      RECT 34.745 1.14 35.12 1.51 ;
      RECT 26.665 0.96 27.04 1.33 ;
      RECT 25.23 0.96 25.605 1.33 ;
      RECT 25.23 1.08 35.05 1.25 ;
      RECT 31.175 4.36 35.03 4.53 ;
      RECT 34.86 3.425 35.03 4.53 ;
      RECT 31.175 3.67 31.345 4.53 ;
      RECT 31.125 3.71 31.405 3.99 ;
      RECT 31.145 3.67 31.405 3.99 ;
      RECT 30.785 3.625 30.89 3.885 ;
      RECT 34.77 3.43 35.12 3.78 ;
      RECT 30.64 2.115 30.73 2.375 ;
      RECT 31.18 3.18 31.185 3.22 ;
      RECT 31.175 3.17 31.18 3.305 ;
      RECT 31.17 3.16 31.175 3.398 ;
      RECT 31.16 3.14 31.17 3.454 ;
      RECT 31.08 3.068 31.16 3.534 ;
      RECT 31.115 3.712 31.125 3.937 ;
      RECT 31.11 3.709 31.115 3.932 ;
      RECT 31.095 3.706 31.11 3.925 ;
      RECT 31.06 3.7 31.095 3.907 ;
      RECT 31.075 3.003 31.08 3.608 ;
      RECT 31.055 2.954 31.075 3.623 ;
      RECT 31.045 3.687 31.06 3.89 ;
      RECT 31.05 2.896 31.055 3.638 ;
      RECT 31.045 2.874 31.05 3.648 ;
      RECT 31.01 2.784 31.045 3.885 ;
      RECT 30.995 2.662 31.01 3.885 ;
      RECT 30.99 2.615 30.995 3.885 ;
      RECT 30.965 2.54 30.99 3.885 ;
      RECT 30.95 2.455 30.965 3.885 ;
      RECT 30.945 2.402 30.95 3.885 ;
      RECT 30.94 2.382 30.945 3.885 ;
      RECT 30.935 2.357 30.94 3.119 ;
      RECT 30.92 3.317 30.94 3.885 ;
      RECT 30.93 2.335 30.935 3.096 ;
      RECT 30.92 2.287 30.93 3.061 ;
      RECT 30.915 2.25 30.92 3.027 ;
      RECT 30.915 3.397 30.92 3.885 ;
      RECT 30.9 2.227 30.915 2.982 ;
      RECT 30.895 3.495 30.915 3.885 ;
      RECT 30.845 2.115 30.9 2.824 ;
      RECT 30.89 3.617 30.895 3.885 ;
      RECT 30.83 2.115 30.845 2.663 ;
      RECT 30.825 2.115 30.83 2.615 ;
      RECT 30.82 2.115 30.825 2.603 ;
      RECT 30.775 2.115 30.82 2.54 ;
      RECT 30.75 2.115 30.775 2.458 ;
      RECT 30.735 2.115 30.75 2.41 ;
      RECT 30.73 2.115 30.735 2.38 ;
      RECT 33.12 2.16 33.38 2.42 ;
      RECT 33.115 2.16 33.38 2.368 ;
      RECT 33.11 2.16 33.38 2.338 ;
      RECT 33.085 2.03 33.365 2.31 ;
      RECT 21.645 6.655 21.995 7.005 ;
      RECT 32.615 6.61 32.965 6.96 ;
      RECT 21.645 6.685 32.965 6.885 ;
      RECT 32.125 3.71 32.405 3.99 ;
      RECT 32.165 3.665 32.43 3.925 ;
      RECT 32.155 3.7 32.43 3.925 ;
      RECT 32.16 3.685 32.405 3.99 ;
      RECT 32.165 3.662 32.375 3.99 ;
      RECT 32.165 3.66 32.36 3.99 ;
      RECT 32.205 3.65 32.36 3.99 ;
      RECT 32.175 3.655 32.36 3.99 ;
      RECT 32.205 3.647 32.305 3.99 ;
      RECT 32.23 3.64 32.305 3.99 ;
      RECT 32.21 3.642 32.305 3.99 ;
      RECT 31.54 3.155 31.8 3.415 ;
      RECT 31.59 3.147 31.78 3.415 ;
      RECT 31.595 3.067 31.78 3.415 ;
      RECT 31.715 2.455 31.78 3.415 ;
      RECT 31.62 2.852 31.78 3.415 ;
      RECT 31.695 2.54 31.78 3.415 ;
      RECT 31.73 2.165 31.866 2.893 ;
      RECT 31.675 2.662 31.866 2.893 ;
      RECT 31.69 2.602 31.78 3.415 ;
      RECT 31.73 2.165 31.89 2.558 ;
      RECT 31.73 2.165 31.9 2.455 ;
      RECT 31.72 2.165 31.98 2.425 ;
      RECT 30.055 3.565 30.1 3.825 ;
      RECT 29.96 2.1 30.105 2.36 ;
      RECT 30.465 2.722 30.475 2.813 ;
      RECT 30.45 2.66 30.465 2.869 ;
      RECT 30.445 2.607 30.45 2.915 ;
      RECT 30.395 2.554 30.445 3.041 ;
      RECT 30.39 2.509 30.395 3.188 ;
      RECT 30.38 2.497 30.39 3.23 ;
      RECT 30.345 2.461 30.38 3.335 ;
      RECT 30.34 2.429 30.345 3.441 ;
      RECT 30.325 2.411 30.34 3.486 ;
      RECT 30.32 2.394 30.325 2.72 ;
      RECT 30.315 2.775 30.325 3.543 ;
      RECT 30.31 2.38 30.32 2.693 ;
      RECT 30.305 2.83 30.315 3.825 ;
      RECT 30.3 2.366 30.31 2.678 ;
      RECT 30.3 2.88 30.305 3.825 ;
      RECT 30.285 2.343 30.3 2.658 ;
      RECT 30.265 3.002 30.3 3.825 ;
      RECT 30.28 2.325 30.285 2.64 ;
      RECT 30.275 2.317 30.28 2.63 ;
      RECT 30.245 2.285 30.275 2.594 ;
      RECT 30.255 3.13 30.265 3.825 ;
      RECT 30.25 3.157 30.255 3.825 ;
      RECT 30.245 3.207 30.25 3.825 ;
      RECT 30.235 2.251 30.245 2.559 ;
      RECT 30.195 3.275 30.245 3.825 ;
      RECT 30.22 2.228 30.235 2.535 ;
      RECT 30.195 2.1 30.22 2.498 ;
      RECT 30.19 2.1 30.195 2.47 ;
      RECT 30.16 3.375 30.195 3.825 ;
      RECT 30.185 2.1 30.19 2.463 ;
      RECT 30.18 2.1 30.185 2.453 ;
      RECT 30.165 2.1 30.18 2.438 ;
      RECT 30.15 2.1 30.165 2.41 ;
      RECT 30.115 3.48 30.16 3.825 ;
      RECT 30.135 2.1 30.15 2.383 ;
      RECT 30.105 2.1 30.135 2.368 ;
      RECT 30.1 3.552 30.115 3.825 ;
      RECT 30.025 2.635 30.065 2.895 ;
      RECT 29.8 2.582 29.805 2.84 ;
      RECT 25.755 2.06 26.015 2.32 ;
      RECT 25.755 2.085 26.03 2.3 ;
      RECT 28.145 1.91 28.15 2.055 ;
      RECT 30.015 2.63 30.025 2.895 ;
      RECT 29.995 2.622 30.015 2.895 ;
      RECT 29.977 2.618 29.995 2.895 ;
      RECT 29.891 2.607 29.977 2.895 ;
      RECT 29.805 2.59 29.891 2.895 ;
      RECT 29.75 2.577 29.8 2.825 ;
      RECT 29.716 2.569 29.75 2.8 ;
      RECT 29.63 2.558 29.716 2.765 ;
      RECT 29.595 2.535 29.63 2.73 ;
      RECT 29.585 2.497 29.595 2.716 ;
      RECT 29.58 2.47 29.585 2.712 ;
      RECT 29.575 2.457 29.58 2.709 ;
      RECT 29.565 2.437 29.575 2.705 ;
      RECT 29.56 2.412 29.565 2.701 ;
      RECT 29.535 2.367 29.56 2.695 ;
      RECT 29.525 2.308 29.535 2.687 ;
      RECT 29.515 2.276 29.525 2.678 ;
      RECT 29.495 2.228 29.515 2.658 ;
      RECT 29.49 2.188 29.495 2.628 ;
      RECT 29.475 2.162 29.49 2.602 ;
      RECT 29.47 2.14 29.475 2.578 ;
      RECT 29.455 2.112 29.47 2.554 ;
      RECT 29.44 2.085 29.455 2.518 ;
      RECT 29.425 2.062 29.44 2.48 ;
      RECT 29.42 2.052 29.425 2.455 ;
      RECT 29.41 2.045 29.42 2.438 ;
      RECT 29.395 2.032 29.41 2.408 ;
      RECT 29.39 2.022 29.395 2.383 ;
      RECT 29.385 2.017 29.39 2.37 ;
      RECT 29.375 2.01 29.385 2.35 ;
      RECT 29.37 2.003 29.375 2.335 ;
      RECT 29.345 1.996 29.37 2.293 ;
      RECT 29.33 1.986 29.345 2.243 ;
      RECT 29.32 1.981 29.33 2.213 ;
      RECT 29.31 1.977 29.32 2.188 ;
      RECT 29.295 1.974 29.31 2.178 ;
      RECT 29.245 1.971 29.295 2.163 ;
      RECT 29.225 1.969 29.245 2.148 ;
      RECT 29.176 1.967 29.225 2.143 ;
      RECT 29.09 1.963 29.176 2.138 ;
      RECT 29.051 1.96 29.09 2.134 ;
      RECT 28.965 1.956 29.051 2.129 ;
      RECT 28.915 1.953 28.965 2.123 ;
      RECT 28.866 1.95 28.915 2.118 ;
      RECT 28.78 1.947 28.866 2.113 ;
      RECT 28.776 1.945 28.78 2.11 ;
      RECT 28.69 1.942 28.776 2.105 ;
      RECT 28.641 1.938 28.69 2.098 ;
      RECT 28.555 1.935 28.641 2.093 ;
      RECT 28.531 1.932 28.555 2.089 ;
      RECT 28.445 1.93 28.531 2.084 ;
      RECT 28.38 1.926 28.445 2.077 ;
      RECT 28.377 1.925 28.38 2.074 ;
      RECT 28.291 1.922 28.377 2.071 ;
      RECT 28.205 1.916 28.291 2.064 ;
      RECT 28.175 1.912 28.205 2.06 ;
      RECT 28.15 1.91 28.175 2.058 ;
      RECT 28.095 1.907 28.145 2.055 ;
      RECT 28.015 1.906 28.095 2.055 ;
      RECT 27.96 1.908 28.015 2.058 ;
      RECT 27.945 1.909 27.96 2.062 ;
      RECT 27.89 1.917 27.945 2.072 ;
      RECT 27.86 1.925 27.89 2.085 ;
      RECT 27.841 1.926 27.86 2.091 ;
      RECT 27.755 1.929 27.841 2.096 ;
      RECT 27.685 1.934 27.755 2.105 ;
      RECT 27.666 1.937 27.685 2.111 ;
      RECT 27.58 1.941 27.666 2.116 ;
      RECT 27.54 1.945 27.58 2.123 ;
      RECT 27.531 1.947 27.54 2.126 ;
      RECT 27.445 1.951 27.531 2.131 ;
      RECT 27.442 1.954 27.445 2.135 ;
      RECT 27.356 1.957 27.442 2.139 ;
      RECT 27.27 1.963 27.356 2.147 ;
      RECT 27.246 1.967 27.27 2.151 ;
      RECT 27.16 1.971 27.246 2.156 ;
      RECT 27.115 1.976 27.16 2.163 ;
      RECT 27.035 1.981 27.115 2.17 ;
      RECT 26.955 1.987 27.035 2.185 ;
      RECT 26.93 1.991 26.955 2.198 ;
      RECT 26.865 1.994 26.93 2.21 ;
      RECT 26.81 1.999 26.865 2.225 ;
      RECT 26.78 2.002 26.81 2.243 ;
      RECT 26.77 2.004 26.78 2.256 ;
      RECT 26.71 2.019 26.77 2.266 ;
      RECT 26.695 2.036 26.71 2.275 ;
      RECT 26.69 2.045 26.695 2.275 ;
      RECT 26.68 2.055 26.69 2.275 ;
      RECT 26.67 2.072 26.68 2.275 ;
      RECT 26.65 2.082 26.67 2.276 ;
      RECT 26.605 2.092 26.65 2.277 ;
      RECT 26.57 2.101 26.605 2.279 ;
      RECT 26.505 2.106 26.57 2.281 ;
      RECT 26.425 2.107 26.505 2.284 ;
      RECT 26.421 2.105 26.425 2.285 ;
      RECT 26.335 2.102 26.421 2.287 ;
      RECT 26.288 2.099 26.335 2.289 ;
      RECT 26.202 2.095 26.288 2.292 ;
      RECT 26.116 2.091 26.202 2.295 ;
      RECT 26.03 2.087 26.116 2.299 ;
      RECT 29.415 3.71 29.445 3.99 ;
      RECT 29.165 3.6 29.185 3.99 ;
      RECT 29.12 3.6 29.185 3.86 ;
      RECT 28.95 2.225 28.985 2.485 ;
      RECT 28.725 2.225 28.785 2.485 ;
      RECT 29.405 3.69 29.415 3.99 ;
      RECT 29.4 3.65 29.405 3.99 ;
      RECT 29.385 3.605 29.4 3.99 ;
      RECT 29.38 3.57 29.385 3.99 ;
      RECT 29.375 3.55 29.38 3.99 ;
      RECT 29.345 3.477 29.375 3.99 ;
      RECT 29.325 3.375 29.345 3.99 ;
      RECT 29.315 3.305 29.325 3.99 ;
      RECT 29.27 3.245 29.315 3.99 ;
      RECT 29.185 3.206 29.27 3.99 ;
      RECT 29.18 3.197 29.185 3.57 ;
      RECT 29.17 3.196 29.18 3.553 ;
      RECT 29.145 3.177 29.17 3.523 ;
      RECT 29.14 3.152 29.145 3.502 ;
      RECT 29.13 3.13 29.14 3.493 ;
      RECT 29.125 3.101 29.13 3.483 ;
      RECT 29.085 3.027 29.125 3.455 ;
      RECT 29.065 2.928 29.085 3.42 ;
      RECT 29.05 2.864 29.065 3.403 ;
      RECT 29.02 2.788 29.05 3.375 ;
      RECT 29 2.703 29.02 3.348 ;
      RECT 28.96 2.599 29 3.255 ;
      RECT 28.955 2.52 28.96 3.163 ;
      RECT 28.95 2.503 28.955 3.14 ;
      RECT 28.945 2.225 28.95 3.12 ;
      RECT 28.915 2.225 28.945 3.058 ;
      RECT 28.91 2.225 28.915 2.99 ;
      RECT 28.9 2.225 28.91 2.955 ;
      RECT 28.89 2.225 28.9 2.92 ;
      RECT 28.825 2.225 28.89 2.775 ;
      RECT 28.82 2.225 28.825 2.645 ;
      RECT 28.79 2.225 28.82 2.578 ;
      RECT 28.785 2.225 28.79 2.503 ;
      RECT 27.965 3.15 28.245 3.43 ;
      RECT 28.005 3.13 28.265 3.39 ;
      RECT 27.995 3.14 28.265 3.39 ;
      RECT 28.005 3.067 28.22 3.43 ;
      RECT 28.06 2.99 28.215 3.43 ;
      RECT 28.065 2.775 28.215 3.43 ;
      RECT 28.055 2.577 28.205 2.828 ;
      RECT 28.045 2.577 28.205 2.695 ;
      RECT 28.04 2.455 28.2 2.598 ;
      RECT 28.025 2.455 28.2 2.503 ;
      RECT 28.02 2.165 28.195 2.48 ;
      RECT 28.005 2.165 28.195 2.45 ;
      RECT 27.965 2.165 28.225 2.425 ;
      RECT 27.875 3.635 27.955 3.895 ;
      RECT 27.28 2.355 27.285 2.62 ;
      RECT 27.16 2.355 27.285 2.615 ;
      RECT 27.835 3.6 27.875 3.895 ;
      RECT 27.79 3.522 27.835 3.895 ;
      RECT 27.77 3.45 27.79 3.895 ;
      RECT 27.76 3.402 27.77 3.895 ;
      RECT 27.725 3.335 27.76 3.895 ;
      RECT 27.695 3.235 27.725 3.895 ;
      RECT 27.675 3.16 27.695 3.695 ;
      RECT 27.665 3.11 27.675 3.65 ;
      RECT 27.66 3.087 27.665 3.623 ;
      RECT 27.655 3.072 27.66 3.61 ;
      RECT 27.65 3.057 27.655 3.588 ;
      RECT 27.645 3.042 27.65 3.57 ;
      RECT 27.62 2.997 27.645 3.525 ;
      RECT 27.61 2.945 27.62 3.468 ;
      RECT 27.6 2.915 27.61 3.435 ;
      RECT 27.59 2.88 27.6 3.403 ;
      RECT 27.555 2.812 27.59 3.335 ;
      RECT 27.55 2.751 27.555 3.27 ;
      RECT 27.54 2.739 27.55 3.25 ;
      RECT 27.535 2.727 27.54 3.23 ;
      RECT 27.53 2.719 27.535 3.218 ;
      RECT 27.525 2.711 27.53 3.198 ;
      RECT 27.515 2.699 27.525 3.17 ;
      RECT 27.505 2.683 27.515 3.14 ;
      RECT 27.48 2.655 27.505 3.078 ;
      RECT 27.47 2.626 27.48 3.023 ;
      RECT 27.455 2.605 27.47 2.983 ;
      RECT 27.45 2.589 27.455 2.955 ;
      RECT 27.445 2.577 27.45 2.945 ;
      RECT 27.44 2.572 27.445 2.918 ;
      RECT 27.435 2.565 27.44 2.905 ;
      RECT 27.42 2.548 27.435 2.878 ;
      RECT 27.41 2.355 27.42 2.838 ;
      RECT 27.4 2.355 27.41 2.805 ;
      RECT 27.39 2.355 27.4 2.78 ;
      RECT 27.32 2.355 27.39 2.715 ;
      RECT 27.31 2.355 27.32 2.663 ;
      RECT 27.295 2.355 27.31 2.645 ;
      RECT 27.285 2.355 27.295 2.63 ;
      RECT 27.115 3.225 27.375 3.485 ;
      RECT 25.65 3.26 25.655 3.467 ;
      RECT 25.285 3.15 25.36 3.465 ;
      RECT 25.1 3.205 25.255 3.465 ;
      RECT 25.285 3.15 25.39 3.43 ;
      RECT 27.1 3.322 27.115 3.483 ;
      RECT 27.075 3.33 27.1 3.488 ;
      RECT 27.05 3.337 27.075 3.493 ;
      RECT 26.987 3.348 27.05 3.502 ;
      RECT 26.901 3.367 26.987 3.519 ;
      RECT 26.815 3.389 26.901 3.538 ;
      RECT 26.8 3.402 26.815 3.549 ;
      RECT 26.76 3.41 26.8 3.556 ;
      RECT 26.74 3.415 26.76 3.563 ;
      RECT 26.702 3.416 26.74 3.566 ;
      RECT 26.616 3.419 26.702 3.567 ;
      RECT 26.53 3.423 26.616 3.568 ;
      RECT 26.481 3.425 26.53 3.57 ;
      RECT 26.395 3.425 26.481 3.572 ;
      RECT 26.355 3.42 26.395 3.574 ;
      RECT 26.345 3.414 26.355 3.575 ;
      RECT 26.305 3.409 26.345 3.572 ;
      RECT 26.295 3.402 26.305 3.568 ;
      RECT 26.28 3.398 26.295 3.566 ;
      RECT 26.263 3.394 26.28 3.564 ;
      RECT 26.177 3.384 26.263 3.556 ;
      RECT 26.091 3.366 26.177 3.542 ;
      RECT 26.005 3.349 26.091 3.528 ;
      RECT 25.98 3.337 26.005 3.519 ;
      RECT 25.91 3.327 25.98 3.512 ;
      RECT 25.865 3.315 25.91 3.503 ;
      RECT 25.805 3.302 25.865 3.495 ;
      RECT 25.8 3.294 25.805 3.49 ;
      RECT 25.765 3.289 25.8 3.488 ;
      RECT 25.71 3.28 25.765 3.481 ;
      RECT 25.67 3.269 25.71 3.473 ;
      RECT 25.655 3.262 25.67 3.469 ;
      RECT 25.635 3.255 25.65 3.466 ;
      RECT 25.62 3.245 25.635 3.464 ;
      RECT 25.605 3.232 25.62 3.461 ;
      RECT 25.58 3.215 25.605 3.457 ;
      RECT 25.565 3.197 25.58 3.454 ;
      RECT 25.54 3.15 25.565 3.452 ;
      RECT 25.516 3.15 25.54 3.449 ;
      RECT 25.43 3.15 25.516 3.441 ;
      RECT 25.39 3.15 25.43 3.433 ;
      RECT 25.255 3.197 25.285 3.465 ;
      RECT 26.935 2.78 27.195 3.04 ;
      RECT 26.895 2.78 27.195 2.918 ;
      RECT 26.86 2.78 27.195 2.903 ;
      RECT 26.805 2.78 27.195 2.883 ;
      RECT 26.725 2.59 27.005 2.87 ;
      RECT 26.725 2.772 27.075 2.87 ;
      RECT 26.725 2.715 27.06 2.87 ;
      RECT 26.725 2.662 27.01 2.87 ;
      RECT 24.555 2.59 24.75 3.375 ;
      RECT 24.635 1.205 24.75 3.375 ;
      RECT 24.49 3.115 24.55 3.375 ;
      RECT 25.86 2.635 26.12 2.895 ;
      RECT 24.545 2.59 24.75 2.87 ;
      RECT 25.855 2.645 26.12 2.83 ;
      RECT 25.57 2.62 25.58 2.77 ;
      RECT 24.805 1.205 24.885 1.55 ;
      RECT 24.54 1.205 24.75 1.55 ;
      RECT 25.845 2.645 25.855 2.829 ;
      RECT 25.835 2.644 25.845 2.826 ;
      RECT 25.826 2.643 25.835 2.824 ;
      RECT 25.74 2.639 25.826 2.814 ;
      RECT 25.666 2.631 25.74 2.796 ;
      RECT 25.58 2.624 25.666 2.779 ;
      RECT 25.52 2.62 25.57 2.769 ;
      RECT 25.485 2.619 25.52 2.766 ;
      RECT 25.43 2.619 25.485 2.768 ;
      RECT 25.395 2.619 25.43 2.772 ;
      RECT 25.309 2.618 25.395 2.779 ;
      RECT 25.223 2.617 25.309 2.789 ;
      RECT 25.137 2.616 25.223 2.8 ;
      RECT 25.051 2.616 25.137 2.81 ;
      RECT 24.965 2.615 25.051 2.82 ;
      RECT 24.93 2.615 24.965 2.86 ;
      RECT 24.925 2.615 24.93 2.903 ;
      RECT 24.9 2.615 24.925 2.92 ;
      RECT 24.825 2.615 24.9 2.935 ;
      RECT 24.805 2.59 24.825 2.948 ;
      RECT 24.8 1.205 24.805 2.958 ;
      RECT 24.775 1.205 24.8 3 ;
      RECT 24.75 1.205 24.775 3.078 ;
      RECT 24.55 2.997 24.555 3.375 ;
      RECT 23.885 2.949 23.9 3.405 ;
      RECT 23.88 3.021 23.986 3.403 ;
      RECT 23.9 2.115 24.035 3.401 ;
      RECT 23.885 2.965 24.04 3.4 ;
      RECT 23.885 3.015 24.045 3.398 ;
      RECT 23.87 3.08 24.045 3.397 ;
      RECT 23.88 3.072 24.05 3.394 ;
      RECT 23.86 3.12 24.05 3.389 ;
      RECT 23.86 3.12 24.065 3.386 ;
      RECT 23.855 3.12 24.065 3.383 ;
      RECT 23.83 3.12 24.09 3.38 ;
      RECT 23.9 2.115 24.06 2.768 ;
      RECT 23.895 2.115 24.06 2.74 ;
      RECT 23.89 2.115 24.06 2.568 ;
      RECT 23.89 2.115 24.08 2.508 ;
      RECT 23.845 2.115 24.105 2.375 ;
      RECT 23.325 2.59 23.605 2.87 ;
      RECT 23.315 2.605 23.605 2.865 ;
      RECT 23.27 2.667 23.605 2.863 ;
      RECT 23.345 2.582 23.51 2.87 ;
      RECT 23.345 2.567 23.466 2.87 ;
      RECT 23.38 2.56 23.466 2.87 ;
      RECT 22.845 3.71 23.125 3.99 ;
      RECT 22.805 3.672 23.1 3.783 ;
      RECT 22.79 3.622 23.08 3.678 ;
      RECT 22.735 3.385 22.995 3.645 ;
      RECT 22.735 3.587 23.075 3.645 ;
      RECT 22.735 3.527 23.07 3.645 ;
      RECT 22.735 3.477 23.05 3.645 ;
      RECT 22.735 3.457 23.045 3.645 ;
      RECT 22.735 3.435 23.04 3.645 ;
      RECT 22.735 3.42 23.01 3.645 ;
      RECT 18.465 6.225 18.785 6.545 ;
      RECT 18.495 5.695 18.665 6.545 ;
      RECT 18.495 5.695 18.67 6.045 ;
      RECT 18.495 5.695 19.47 5.87 ;
      RECT 19.295 1.965 19.47 5.87 ;
      RECT 19.24 1.965 19.59 2.315 ;
      RECT 19.265 6.655 19.59 6.98 ;
      RECT 18.15 6.745 19.59 6.915 ;
      RECT 18.15 2.395 18.31 6.915 ;
      RECT 18.465 2.365 18.785 2.685 ;
      RECT 18.15 2.395 18.785 2.565 ;
      RECT 16.82 1.14 17.195 1.51 ;
      RECT 8.74 0.96 9.115 1.33 ;
      RECT 7.305 0.96 7.68 1.33 ;
      RECT 7.305 1.08 17.125 1.25 ;
      RECT 13.25 4.36 17.105 4.53 ;
      RECT 16.935 3.425 17.105 4.53 ;
      RECT 13.25 3.67 13.42 4.53 ;
      RECT 13.2 3.71 13.48 3.99 ;
      RECT 13.22 3.67 13.48 3.99 ;
      RECT 12.86 3.625 12.965 3.885 ;
      RECT 16.845 3.43 17.195 3.78 ;
      RECT 12.715 2.115 12.805 2.375 ;
      RECT 13.255 3.18 13.26 3.22 ;
      RECT 13.25 3.17 13.255 3.305 ;
      RECT 13.245 3.16 13.25 3.398 ;
      RECT 13.235 3.14 13.245 3.454 ;
      RECT 13.155 3.068 13.235 3.534 ;
      RECT 13.19 3.712 13.2 3.937 ;
      RECT 13.185 3.709 13.19 3.932 ;
      RECT 13.17 3.706 13.185 3.925 ;
      RECT 13.135 3.7 13.17 3.907 ;
      RECT 13.15 3.003 13.155 3.608 ;
      RECT 13.13 2.954 13.15 3.623 ;
      RECT 13.12 3.687 13.135 3.89 ;
      RECT 13.125 2.896 13.13 3.638 ;
      RECT 13.12 2.874 13.125 3.648 ;
      RECT 13.085 2.784 13.12 3.885 ;
      RECT 13.07 2.662 13.085 3.885 ;
      RECT 13.065 2.615 13.07 3.885 ;
      RECT 13.04 2.54 13.065 3.885 ;
      RECT 13.025 2.455 13.04 3.885 ;
      RECT 13.02 2.402 13.025 3.885 ;
      RECT 13.015 2.382 13.02 3.885 ;
      RECT 13.01 2.357 13.015 3.119 ;
      RECT 12.995 3.317 13.015 3.885 ;
      RECT 13.005 2.335 13.01 3.096 ;
      RECT 12.995 2.287 13.005 3.061 ;
      RECT 12.99 2.25 12.995 3.027 ;
      RECT 12.99 3.397 12.995 3.885 ;
      RECT 12.975 2.227 12.99 2.982 ;
      RECT 12.97 3.495 12.99 3.885 ;
      RECT 12.92 2.115 12.975 2.824 ;
      RECT 12.965 3.617 12.97 3.885 ;
      RECT 12.905 2.115 12.92 2.663 ;
      RECT 12.9 2.115 12.905 2.615 ;
      RECT 12.895 2.115 12.9 2.603 ;
      RECT 12.85 2.115 12.895 2.54 ;
      RECT 12.825 2.115 12.85 2.458 ;
      RECT 12.81 2.115 12.825 2.41 ;
      RECT 12.805 2.115 12.81 2.38 ;
      RECT 15.195 2.16 15.455 2.42 ;
      RECT 15.19 2.16 15.455 2.368 ;
      RECT 15.185 2.16 15.455 2.338 ;
      RECT 15.16 2.03 15.44 2.31 ;
      RECT 3.02 6.995 3.31 7.345 ;
      RECT 3.02 7.055 4.155 7.225 ;
      RECT 3.985 6.685 4.155 7.225 ;
      RECT 14.71 6.605 14.88 6.96 ;
      RECT 14.66 6.605 15.01 6.955 ;
      RECT 3.985 6.685 15.01 6.855 ;
      RECT 14.2 3.71 14.48 3.99 ;
      RECT 14.24 3.665 14.505 3.925 ;
      RECT 14.23 3.7 14.505 3.925 ;
      RECT 14.235 3.685 14.48 3.99 ;
      RECT 14.24 3.662 14.45 3.99 ;
      RECT 14.24 3.66 14.435 3.99 ;
      RECT 14.28 3.65 14.435 3.99 ;
      RECT 14.25 3.655 14.435 3.99 ;
      RECT 14.28 3.647 14.38 3.99 ;
      RECT 14.305 3.64 14.38 3.99 ;
      RECT 14.285 3.642 14.38 3.99 ;
      RECT 13.615 3.155 13.875 3.415 ;
      RECT 13.665 3.147 13.855 3.415 ;
      RECT 13.67 3.067 13.855 3.415 ;
      RECT 13.79 2.455 13.855 3.415 ;
      RECT 13.695 2.852 13.855 3.415 ;
      RECT 13.77 2.54 13.855 3.415 ;
      RECT 13.805 2.165 13.941 2.893 ;
      RECT 13.75 2.662 13.941 2.893 ;
      RECT 13.765 2.602 13.855 3.415 ;
      RECT 13.805 2.165 13.965 2.558 ;
      RECT 13.805 2.165 13.975 2.455 ;
      RECT 13.795 2.165 14.055 2.425 ;
      RECT 12.13 3.565 12.175 3.825 ;
      RECT 12.035 2.1 12.18 2.36 ;
      RECT 12.54 2.722 12.55 2.813 ;
      RECT 12.525 2.66 12.54 2.869 ;
      RECT 12.52 2.607 12.525 2.915 ;
      RECT 12.47 2.554 12.52 3.041 ;
      RECT 12.465 2.509 12.47 3.188 ;
      RECT 12.455 2.497 12.465 3.23 ;
      RECT 12.42 2.461 12.455 3.335 ;
      RECT 12.415 2.429 12.42 3.441 ;
      RECT 12.4 2.411 12.415 3.486 ;
      RECT 12.395 2.394 12.4 2.72 ;
      RECT 12.39 2.775 12.4 3.543 ;
      RECT 12.385 2.38 12.395 2.693 ;
      RECT 12.38 2.83 12.39 3.825 ;
      RECT 12.375 2.366 12.385 2.678 ;
      RECT 12.375 2.88 12.38 3.825 ;
      RECT 12.36 2.343 12.375 2.658 ;
      RECT 12.34 3.002 12.375 3.825 ;
      RECT 12.355 2.325 12.36 2.64 ;
      RECT 12.35 2.317 12.355 2.63 ;
      RECT 12.32 2.285 12.35 2.594 ;
      RECT 12.33 3.13 12.34 3.825 ;
      RECT 12.325 3.157 12.33 3.825 ;
      RECT 12.32 3.207 12.325 3.825 ;
      RECT 12.31 2.251 12.32 2.559 ;
      RECT 12.27 3.275 12.32 3.825 ;
      RECT 12.295 2.228 12.31 2.535 ;
      RECT 12.27 2.1 12.295 2.498 ;
      RECT 12.265 2.1 12.27 2.47 ;
      RECT 12.235 3.375 12.27 3.825 ;
      RECT 12.26 2.1 12.265 2.463 ;
      RECT 12.255 2.1 12.26 2.453 ;
      RECT 12.24 2.1 12.255 2.438 ;
      RECT 12.225 2.1 12.24 2.41 ;
      RECT 12.19 3.48 12.235 3.825 ;
      RECT 12.21 2.1 12.225 2.383 ;
      RECT 12.18 2.1 12.21 2.368 ;
      RECT 12.175 3.552 12.19 3.825 ;
      RECT 12.1 2.635 12.14 2.895 ;
      RECT 11.875 2.582 11.88 2.84 ;
      RECT 7.83 2.06 8.09 2.32 ;
      RECT 7.83 2.085 8.105 2.3 ;
      RECT 10.22 1.91 10.225 2.055 ;
      RECT 12.09 2.63 12.1 2.895 ;
      RECT 12.07 2.622 12.09 2.895 ;
      RECT 12.052 2.618 12.07 2.895 ;
      RECT 11.966 2.607 12.052 2.895 ;
      RECT 11.88 2.59 11.966 2.895 ;
      RECT 11.825 2.577 11.875 2.825 ;
      RECT 11.791 2.569 11.825 2.8 ;
      RECT 11.705 2.558 11.791 2.765 ;
      RECT 11.67 2.535 11.705 2.73 ;
      RECT 11.66 2.497 11.67 2.716 ;
      RECT 11.655 2.47 11.66 2.712 ;
      RECT 11.65 2.457 11.655 2.709 ;
      RECT 11.64 2.437 11.65 2.705 ;
      RECT 11.635 2.412 11.64 2.701 ;
      RECT 11.61 2.367 11.635 2.695 ;
      RECT 11.6 2.308 11.61 2.687 ;
      RECT 11.59 2.276 11.6 2.678 ;
      RECT 11.57 2.228 11.59 2.658 ;
      RECT 11.565 2.188 11.57 2.628 ;
      RECT 11.55 2.162 11.565 2.602 ;
      RECT 11.545 2.14 11.55 2.578 ;
      RECT 11.53 2.112 11.545 2.554 ;
      RECT 11.515 2.085 11.53 2.518 ;
      RECT 11.5 2.062 11.515 2.48 ;
      RECT 11.495 2.052 11.5 2.455 ;
      RECT 11.485 2.045 11.495 2.438 ;
      RECT 11.47 2.032 11.485 2.408 ;
      RECT 11.465 2.022 11.47 2.383 ;
      RECT 11.46 2.017 11.465 2.37 ;
      RECT 11.45 2.01 11.46 2.35 ;
      RECT 11.445 2.003 11.45 2.335 ;
      RECT 11.42 1.996 11.445 2.293 ;
      RECT 11.405 1.986 11.42 2.243 ;
      RECT 11.395 1.981 11.405 2.213 ;
      RECT 11.385 1.977 11.395 2.188 ;
      RECT 11.37 1.974 11.385 2.178 ;
      RECT 11.32 1.971 11.37 2.163 ;
      RECT 11.3 1.969 11.32 2.148 ;
      RECT 11.251 1.967 11.3 2.143 ;
      RECT 11.165 1.963 11.251 2.138 ;
      RECT 11.126 1.96 11.165 2.134 ;
      RECT 11.04 1.956 11.126 2.129 ;
      RECT 10.99 1.953 11.04 2.123 ;
      RECT 10.941 1.95 10.99 2.118 ;
      RECT 10.855 1.947 10.941 2.113 ;
      RECT 10.851 1.945 10.855 2.11 ;
      RECT 10.765 1.942 10.851 2.105 ;
      RECT 10.716 1.938 10.765 2.098 ;
      RECT 10.63 1.935 10.716 2.093 ;
      RECT 10.606 1.932 10.63 2.089 ;
      RECT 10.52 1.93 10.606 2.084 ;
      RECT 10.455 1.926 10.52 2.077 ;
      RECT 10.452 1.925 10.455 2.074 ;
      RECT 10.366 1.922 10.452 2.071 ;
      RECT 10.28 1.916 10.366 2.064 ;
      RECT 10.25 1.912 10.28 2.06 ;
      RECT 10.225 1.91 10.25 2.058 ;
      RECT 10.17 1.907 10.22 2.055 ;
      RECT 10.09 1.906 10.17 2.055 ;
      RECT 10.035 1.908 10.09 2.058 ;
      RECT 10.02 1.909 10.035 2.062 ;
      RECT 9.965 1.917 10.02 2.072 ;
      RECT 9.935 1.925 9.965 2.085 ;
      RECT 9.916 1.926 9.935 2.091 ;
      RECT 9.83 1.929 9.916 2.096 ;
      RECT 9.76 1.934 9.83 2.105 ;
      RECT 9.741 1.937 9.76 2.111 ;
      RECT 9.655 1.941 9.741 2.116 ;
      RECT 9.615 1.945 9.655 2.123 ;
      RECT 9.606 1.947 9.615 2.126 ;
      RECT 9.52 1.951 9.606 2.131 ;
      RECT 9.517 1.954 9.52 2.135 ;
      RECT 9.431 1.957 9.517 2.139 ;
      RECT 9.345 1.963 9.431 2.147 ;
      RECT 9.321 1.967 9.345 2.151 ;
      RECT 9.235 1.971 9.321 2.156 ;
      RECT 9.19 1.976 9.235 2.163 ;
      RECT 9.11 1.981 9.19 2.17 ;
      RECT 9.03 1.987 9.11 2.185 ;
      RECT 9.005 1.991 9.03 2.198 ;
      RECT 8.94 1.994 9.005 2.21 ;
      RECT 8.885 1.999 8.94 2.225 ;
      RECT 8.855 2.002 8.885 2.243 ;
      RECT 8.845 2.004 8.855 2.256 ;
      RECT 8.785 2.019 8.845 2.266 ;
      RECT 8.77 2.036 8.785 2.275 ;
      RECT 8.765 2.045 8.77 2.275 ;
      RECT 8.755 2.055 8.765 2.275 ;
      RECT 8.745 2.072 8.755 2.275 ;
      RECT 8.725 2.082 8.745 2.276 ;
      RECT 8.68 2.092 8.725 2.277 ;
      RECT 8.645 2.101 8.68 2.279 ;
      RECT 8.58 2.106 8.645 2.281 ;
      RECT 8.5 2.107 8.58 2.284 ;
      RECT 8.496 2.105 8.5 2.285 ;
      RECT 8.41 2.102 8.496 2.287 ;
      RECT 8.363 2.099 8.41 2.289 ;
      RECT 8.277 2.095 8.363 2.292 ;
      RECT 8.191 2.091 8.277 2.295 ;
      RECT 8.105 2.087 8.191 2.299 ;
      RECT 11.49 3.71 11.52 3.99 ;
      RECT 11.24 3.6 11.26 3.99 ;
      RECT 11.195 3.6 11.26 3.86 ;
      RECT 11.025 2.225 11.06 2.485 ;
      RECT 10.8 2.225 10.86 2.485 ;
      RECT 11.48 3.69 11.49 3.99 ;
      RECT 11.475 3.65 11.48 3.99 ;
      RECT 11.46 3.605 11.475 3.99 ;
      RECT 11.455 3.57 11.46 3.99 ;
      RECT 11.45 3.55 11.455 3.99 ;
      RECT 11.42 3.477 11.45 3.99 ;
      RECT 11.4 3.375 11.42 3.99 ;
      RECT 11.39 3.305 11.4 3.99 ;
      RECT 11.345 3.245 11.39 3.99 ;
      RECT 11.26 3.206 11.345 3.99 ;
      RECT 11.255 3.197 11.26 3.57 ;
      RECT 11.245 3.196 11.255 3.553 ;
      RECT 11.22 3.177 11.245 3.523 ;
      RECT 11.215 3.152 11.22 3.502 ;
      RECT 11.205 3.13 11.215 3.493 ;
      RECT 11.2 3.101 11.205 3.483 ;
      RECT 11.16 3.027 11.2 3.455 ;
      RECT 11.14 2.928 11.16 3.42 ;
      RECT 11.125 2.864 11.14 3.403 ;
      RECT 11.095 2.788 11.125 3.375 ;
      RECT 11.075 2.703 11.095 3.348 ;
      RECT 11.035 2.599 11.075 3.255 ;
      RECT 11.03 2.52 11.035 3.163 ;
      RECT 11.025 2.503 11.03 3.14 ;
      RECT 11.02 2.225 11.025 3.12 ;
      RECT 10.99 2.225 11.02 3.058 ;
      RECT 10.985 2.225 10.99 2.99 ;
      RECT 10.975 2.225 10.985 2.955 ;
      RECT 10.965 2.225 10.975 2.92 ;
      RECT 10.9 2.225 10.965 2.775 ;
      RECT 10.895 2.225 10.9 2.645 ;
      RECT 10.865 2.225 10.895 2.578 ;
      RECT 10.86 2.225 10.865 2.503 ;
      RECT 10.04 3.15 10.32 3.43 ;
      RECT 10.08 3.13 10.34 3.39 ;
      RECT 10.07 3.14 10.34 3.39 ;
      RECT 10.08 3.067 10.295 3.43 ;
      RECT 10.135 2.99 10.29 3.43 ;
      RECT 10.14 2.775 10.29 3.43 ;
      RECT 10.13 2.577 10.28 2.828 ;
      RECT 10.12 2.577 10.28 2.695 ;
      RECT 10.115 2.455 10.275 2.598 ;
      RECT 10.1 2.455 10.275 2.503 ;
      RECT 10.095 2.165 10.27 2.48 ;
      RECT 10.08 2.165 10.27 2.45 ;
      RECT 10.04 2.165 10.3 2.425 ;
      RECT 9.95 3.635 10.03 3.895 ;
      RECT 9.355 2.355 9.36 2.62 ;
      RECT 9.235 2.355 9.36 2.615 ;
      RECT 9.91 3.6 9.95 3.895 ;
      RECT 9.865 3.522 9.91 3.895 ;
      RECT 9.845 3.45 9.865 3.895 ;
      RECT 9.835 3.402 9.845 3.895 ;
      RECT 9.8 3.335 9.835 3.895 ;
      RECT 9.77 3.235 9.8 3.895 ;
      RECT 9.75 3.16 9.77 3.695 ;
      RECT 9.74 3.11 9.75 3.65 ;
      RECT 9.735 3.087 9.74 3.623 ;
      RECT 9.73 3.072 9.735 3.61 ;
      RECT 9.725 3.057 9.73 3.588 ;
      RECT 9.72 3.042 9.725 3.57 ;
      RECT 9.695 2.997 9.72 3.525 ;
      RECT 9.685 2.945 9.695 3.468 ;
      RECT 9.675 2.915 9.685 3.435 ;
      RECT 9.665 2.88 9.675 3.403 ;
      RECT 9.63 2.812 9.665 3.335 ;
      RECT 9.625 2.751 9.63 3.27 ;
      RECT 9.615 2.739 9.625 3.25 ;
      RECT 9.61 2.727 9.615 3.23 ;
      RECT 9.605 2.719 9.61 3.218 ;
      RECT 9.6 2.711 9.605 3.198 ;
      RECT 9.59 2.699 9.6 3.17 ;
      RECT 9.58 2.683 9.59 3.14 ;
      RECT 9.555 2.655 9.58 3.078 ;
      RECT 9.545 2.626 9.555 3.023 ;
      RECT 9.53 2.605 9.545 2.983 ;
      RECT 9.525 2.589 9.53 2.955 ;
      RECT 9.52 2.577 9.525 2.945 ;
      RECT 9.515 2.572 9.52 2.918 ;
      RECT 9.51 2.565 9.515 2.905 ;
      RECT 9.495 2.548 9.51 2.878 ;
      RECT 9.485 2.355 9.495 2.838 ;
      RECT 9.475 2.355 9.485 2.805 ;
      RECT 9.465 2.355 9.475 2.78 ;
      RECT 9.395 2.355 9.465 2.715 ;
      RECT 9.385 2.355 9.395 2.663 ;
      RECT 9.37 2.355 9.385 2.645 ;
      RECT 9.36 2.355 9.37 2.63 ;
      RECT 9.19 3.225 9.45 3.485 ;
      RECT 7.725 3.26 7.73 3.467 ;
      RECT 7.36 3.15 7.435 3.465 ;
      RECT 7.175 3.205 7.33 3.465 ;
      RECT 7.36 3.15 7.465 3.43 ;
      RECT 9.175 3.322 9.19 3.483 ;
      RECT 9.15 3.33 9.175 3.488 ;
      RECT 9.125 3.337 9.15 3.493 ;
      RECT 9.062 3.348 9.125 3.502 ;
      RECT 8.976 3.367 9.062 3.519 ;
      RECT 8.89 3.389 8.976 3.538 ;
      RECT 8.875 3.402 8.89 3.549 ;
      RECT 8.835 3.41 8.875 3.556 ;
      RECT 8.815 3.415 8.835 3.563 ;
      RECT 8.777 3.416 8.815 3.566 ;
      RECT 8.691 3.419 8.777 3.567 ;
      RECT 8.605 3.423 8.691 3.568 ;
      RECT 8.556 3.425 8.605 3.57 ;
      RECT 8.47 3.425 8.556 3.572 ;
      RECT 8.43 3.42 8.47 3.574 ;
      RECT 8.42 3.414 8.43 3.575 ;
      RECT 8.38 3.409 8.42 3.572 ;
      RECT 8.37 3.402 8.38 3.568 ;
      RECT 8.355 3.398 8.37 3.566 ;
      RECT 8.338 3.394 8.355 3.564 ;
      RECT 8.252 3.384 8.338 3.556 ;
      RECT 8.166 3.366 8.252 3.542 ;
      RECT 8.08 3.349 8.166 3.528 ;
      RECT 8.055 3.337 8.08 3.519 ;
      RECT 7.985 3.327 8.055 3.512 ;
      RECT 7.94 3.315 7.985 3.503 ;
      RECT 7.88 3.302 7.94 3.495 ;
      RECT 7.875 3.294 7.88 3.49 ;
      RECT 7.84 3.289 7.875 3.488 ;
      RECT 7.785 3.28 7.84 3.481 ;
      RECT 7.745 3.269 7.785 3.473 ;
      RECT 7.73 3.262 7.745 3.469 ;
      RECT 7.71 3.255 7.725 3.466 ;
      RECT 7.695 3.245 7.71 3.464 ;
      RECT 7.68 3.232 7.695 3.461 ;
      RECT 7.655 3.215 7.68 3.457 ;
      RECT 7.64 3.197 7.655 3.454 ;
      RECT 7.615 3.15 7.64 3.452 ;
      RECT 7.591 3.15 7.615 3.449 ;
      RECT 7.505 3.15 7.591 3.441 ;
      RECT 7.465 3.15 7.505 3.433 ;
      RECT 7.33 3.197 7.36 3.465 ;
      RECT 9.01 2.78 9.27 3.04 ;
      RECT 8.97 2.78 9.27 2.918 ;
      RECT 8.935 2.78 9.27 2.903 ;
      RECT 8.88 2.78 9.27 2.883 ;
      RECT 8.8 2.59 9.08 2.87 ;
      RECT 8.8 2.772 9.15 2.87 ;
      RECT 8.8 2.715 9.135 2.87 ;
      RECT 8.8 2.662 9.085 2.87 ;
      RECT 6.63 2.59 6.825 3.375 ;
      RECT 6.71 1.205 6.825 3.375 ;
      RECT 6.565 3.115 6.625 3.375 ;
      RECT 7.935 2.635 8.195 2.895 ;
      RECT 6.62 2.59 6.825 2.87 ;
      RECT 7.93 2.645 8.195 2.83 ;
      RECT 7.645 2.62 7.655 2.77 ;
      RECT 6.88 1.205 6.96 1.55 ;
      RECT 6.615 1.205 6.825 1.55 ;
      RECT 7.92 2.645 7.93 2.829 ;
      RECT 7.91 2.644 7.92 2.826 ;
      RECT 7.901 2.643 7.91 2.824 ;
      RECT 7.815 2.639 7.901 2.814 ;
      RECT 7.741 2.631 7.815 2.796 ;
      RECT 7.655 2.624 7.741 2.779 ;
      RECT 7.595 2.62 7.645 2.769 ;
      RECT 7.56 2.619 7.595 2.766 ;
      RECT 7.505 2.619 7.56 2.768 ;
      RECT 7.47 2.619 7.505 2.772 ;
      RECT 7.384 2.618 7.47 2.779 ;
      RECT 7.298 2.617 7.384 2.789 ;
      RECT 7.212 2.616 7.298 2.8 ;
      RECT 7.126 2.616 7.212 2.81 ;
      RECT 7.04 2.615 7.126 2.82 ;
      RECT 7.005 2.615 7.04 2.86 ;
      RECT 7 2.615 7.005 2.903 ;
      RECT 6.975 2.615 7 2.92 ;
      RECT 6.9 2.615 6.975 2.935 ;
      RECT 6.88 2.59 6.9 2.948 ;
      RECT 6.875 1.205 6.88 2.958 ;
      RECT 6.85 1.205 6.875 3 ;
      RECT 6.825 1.205 6.85 3.078 ;
      RECT 6.625 2.997 6.63 3.375 ;
      RECT 5.96 2.949 5.975 3.405 ;
      RECT 5.955 3.021 6.061 3.403 ;
      RECT 5.975 2.115 6.11 3.401 ;
      RECT 5.96 2.965 6.115 3.4 ;
      RECT 5.96 3.015 6.12 3.398 ;
      RECT 5.945 3.08 6.12 3.397 ;
      RECT 5.955 3.072 6.125 3.394 ;
      RECT 5.935 3.12 6.125 3.389 ;
      RECT 5.935 3.12 6.14 3.386 ;
      RECT 5.93 3.12 6.14 3.383 ;
      RECT 5.905 3.12 6.165 3.38 ;
      RECT 5.975 2.115 6.135 2.768 ;
      RECT 5.97 2.115 6.135 2.74 ;
      RECT 5.965 2.115 6.135 2.568 ;
      RECT 5.965 2.115 6.155 2.508 ;
      RECT 5.92 2.115 6.18 2.375 ;
      RECT 5.4 2.59 5.68 2.87 ;
      RECT 5.39 2.605 5.68 2.865 ;
      RECT 5.345 2.667 5.68 2.863 ;
      RECT 5.42 2.582 5.585 2.87 ;
      RECT 5.42 2.567 5.541 2.87 ;
      RECT 5.455 2.56 5.541 2.87 ;
      RECT 4.92 3.71 5.2 3.99 ;
      RECT 4.88 3.672 5.175 3.783 ;
      RECT 4.865 3.622 5.155 3.678 ;
      RECT 4.81 3.385 5.07 3.645 ;
      RECT 4.81 3.587 5.15 3.645 ;
      RECT 4.81 3.527 5.145 3.645 ;
      RECT 4.81 3.477 5.125 3.645 ;
      RECT 4.81 3.457 5.12 3.645 ;
      RECT 4.81 3.435 5.115 3.645 ;
      RECT 4.81 3.42 5.085 3.645 ;
      RECT 85.7 7.055 86.075 7.425 ;
      RECT 77.035 0.93 77.41 1.3 ;
      RECT 67.775 7.055 68.15 7.425 ;
      RECT 59.11 0.93 59.485 1.3 ;
      RECT 49.85 7.055 50.225 7.425 ;
      RECT 41.185 0.93 41.56 1.3 ;
      RECT 31.925 7.055 32.3 7.425 ;
      RECT 23.26 0.93 23.635 1.3 ;
      RECT 14 7.055 14.375 7.425 ;
      RECT 5.335 0.93 5.71 1.3 ;
    LAYER via1 ;
      RECT 93.42 7.375 93.57 7.525 ;
      RECT 91.055 6.74 91.205 6.89 ;
      RECT 91.04 2.065 91.19 2.215 ;
      RECT 90.25 2.45 90.4 2.6 ;
      RECT 90.25 6.325 90.4 6.475 ;
      RECT 88.645 3.53 88.795 3.68 ;
      RECT 88.635 1.25 88.785 1.4 ;
      RECT 86.95 2.215 87.1 2.365 ;
      RECT 86.72 6.71 86.87 6.86 ;
      RECT 86 3.72 86.15 3.87 ;
      RECT 85.815 7.165 85.965 7.315 ;
      RECT 85.55 2.22 85.7 2.37 ;
      RECT 85.37 3.21 85.52 3.36 ;
      RECT 84.975 3.725 85.125 3.875 ;
      RECT 84.615 3.68 84.765 3.83 ;
      RECT 84.47 2.17 84.62 2.32 ;
      RECT 83.885 3.62 84.035 3.77 ;
      RECT 83.79 2.155 83.94 2.305 ;
      RECT 83.635 2.69 83.785 2.84 ;
      RECT 82.95 3.655 83.1 3.805 ;
      RECT 82.555 2.28 82.705 2.43 ;
      RECT 81.835 3.185 81.985 3.335 ;
      RECT 81.795 2.22 81.945 2.37 ;
      RECT 81.525 3.69 81.675 3.84 ;
      RECT 80.99 2.41 81.14 2.56 ;
      RECT 80.945 3.28 81.095 3.43 ;
      RECT 80.765 2.835 80.915 2.985 ;
      RECT 79.69 2.69 79.84 2.84 ;
      RECT 79.585 2.115 79.735 2.265 ;
      RECT 78.93 3.26 79.08 3.41 ;
      RECT 78.41 1.3 78.56 1.45 ;
      RECT 78.32 3.17 78.47 3.32 ;
      RECT 77.675 2.17 77.825 2.32 ;
      RECT 77.66 3.175 77.81 3.325 ;
      RECT 77.145 2.66 77.295 2.81 ;
      RECT 76.565 3.44 76.715 3.59 ;
      RECT 75.475 6.755 75.625 6.905 ;
      RECT 73.13 6.74 73.28 6.89 ;
      RECT 73.115 2.065 73.265 2.215 ;
      RECT 72.325 2.45 72.475 2.6 ;
      RECT 72.325 6.325 72.475 6.475 ;
      RECT 70.72 3.53 70.87 3.68 ;
      RECT 70.71 1.25 70.86 1.4 ;
      RECT 69.025 2.215 69.175 2.365 ;
      RECT 68.515 6.71 68.665 6.86 ;
      RECT 68.075 3.72 68.225 3.87 ;
      RECT 67.89 7.165 68.04 7.315 ;
      RECT 67.625 2.22 67.775 2.37 ;
      RECT 67.445 3.21 67.595 3.36 ;
      RECT 67.05 3.725 67.2 3.875 ;
      RECT 66.69 3.68 66.84 3.83 ;
      RECT 66.545 2.17 66.695 2.32 ;
      RECT 65.96 3.62 66.11 3.77 ;
      RECT 65.865 2.155 66.015 2.305 ;
      RECT 65.71 2.69 65.86 2.84 ;
      RECT 65.025 3.655 65.175 3.805 ;
      RECT 64.63 2.28 64.78 2.43 ;
      RECT 63.91 3.185 64.06 3.335 ;
      RECT 63.87 2.22 64.02 2.37 ;
      RECT 63.6 3.69 63.75 3.84 ;
      RECT 63.065 2.41 63.215 2.56 ;
      RECT 63.02 3.28 63.17 3.43 ;
      RECT 62.84 2.835 62.99 2.985 ;
      RECT 61.765 2.69 61.915 2.84 ;
      RECT 61.66 2.115 61.81 2.265 ;
      RECT 61.005 3.26 61.155 3.41 ;
      RECT 60.485 1.3 60.635 1.45 ;
      RECT 60.395 3.17 60.545 3.32 ;
      RECT 59.75 2.17 59.9 2.32 ;
      RECT 59.735 3.175 59.885 3.325 ;
      RECT 59.22 2.66 59.37 2.81 ;
      RECT 58.64 3.44 58.79 3.59 ;
      RECT 57.55 6.755 57.7 6.905 ;
      RECT 55.205 6.74 55.355 6.89 ;
      RECT 55.19 2.065 55.34 2.215 ;
      RECT 54.4 2.45 54.55 2.6 ;
      RECT 54.4 6.325 54.55 6.475 ;
      RECT 52.795 3.53 52.945 3.68 ;
      RECT 52.785 1.25 52.935 1.4 ;
      RECT 51.1 2.215 51.25 2.365 ;
      RECT 50.645 6.715 50.795 6.865 ;
      RECT 50.15 3.72 50.3 3.87 ;
      RECT 49.965 7.165 50.115 7.315 ;
      RECT 49.7 2.22 49.85 2.37 ;
      RECT 49.52 3.21 49.67 3.36 ;
      RECT 49.125 3.725 49.275 3.875 ;
      RECT 48.765 3.68 48.915 3.83 ;
      RECT 48.62 2.17 48.77 2.32 ;
      RECT 48.035 3.62 48.185 3.77 ;
      RECT 47.94 2.155 48.09 2.305 ;
      RECT 47.785 2.69 47.935 2.84 ;
      RECT 47.1 3.655 47.25 3.805 ;
      RECT 46.705 2.28 46.855 2.43 ;
      RECT 45.985 3.185 46.135 3.335 ;
      RECT 45.945 2.22 46.095 2.37 ;
      RECT 45.675 3.69 45.825 3.84 ;
      RECT 45.14 2.41 45.29 2.56 ;
      RECT 45.095 3.28 45.245 3.43 ;
      RECT 44.915 2.835 45.065 2.985 ;
      RECT 43.84 2.69 43.99 2.84 ;
      RECT 43.735 2.115 43.885 2.265 ;
      RECT 43.08 3.26 43.23 3.41 ;
      RECT 42.56 1.3 42.71 1.45 ;
      RECT 42.47 3.17 42.62 3.32 ;
      RECT 41.825 2.17 41.975 2.32 ;
      RECT 41.81 3.175 41.96 3.325 ;
      RECT 41.295 2.66 41.445 2.81 ;
      RECT 40.715 3.44 40.865 3.59 ;
      RECT 39.67 6.76 39.82 6.91 ;
      RECT 37.28 6.74 37.43 6.89 ;
      RECT 37.265 2.065 37.415 2.215 ;
      RECT 36.475 2.45 36.625 2.6 ;
      RECT 36.475 6.325 36.625 6.475 ;
      RECT 34.87 3.53 35.02 3.68 ;
      RECT 34.86 1.25 35.01 1.4 ;
      RECT 33.175 2.215 33.325 2.365 ;
      RECT 32.715 6.71 32.865 6.86 ;
      RECT 32.225 3.72 32.375 3.87 ;
      RECT 32.04 7.165 32.19 7.315 ;
      RECT 31.775 2.22 31.925 2.37 ;
      RECT 31.595 3.21 31.745 3.36 ;
      RECT 31.2 3.725 31.35 3.875 ;
      RECT 30.84 3.68 30.99 3.83 ;
      RECT 30.695 2.17 30.845 2.32 ;
      RECT 30.11 3.62 30.26 3.77 ;
      RECT 30.015 2.155 30.165 2.305 ;
      RECT 29.86 2.69 30.01 2.84 ;
      RECT 29.175 3.655 29.325 3.805 ;
      RECT 28.78 2.28 28.93 2.43 ;
      RECT 28.06 3.185 28.21 3.335 ;
      RECT 28.02 2.22 28.17 2.37 ;
      RECT 27.75 3.69 27.9 3.84 ;
      RECT 27.215 2.41 27.365 2.56 ;
      RECT 27.17 3.28 27.32 3.43 ;
      RECT 26.99 2.835 27.14 2.985 ;
      RECT 25.915 2.69 26.065 2.84 ;
      RECT 25.81 2.115 25.96 2.265 ;
      RECT 25.155 3.26 25.305 3.41 ;
      RECT 24.635 1.3 24.785 1.45 ;
      RECT 24.545 3.17 24.695 3.32 ;
      RECT 23.9 2.17 24.05 2.32 ;
      RECT 23.885 3.175 24.035 3.325 ;
      RECT 23.37 2.66 23.52 2.81 ;
      RECT 22.79 3.44 22.94 3.59 ;
      RECT 21.745 6.755 21.895 6.905 ;
      RECT 19.355 6.74 19.505 6.89 ;
      RECT 19.34 2.065 19.49 2.215 ;
      RECT 18.55 2.45 18.7 2.6 ;
      RECT 18.55 6.325 18.7 6.475 ;
      RECT 16.945 3.53 17.095 3.68 ;
      RECT 16.935 1.25 17.085 1.4 ;
      RECT 15.25 2.215 15.4 2.365 ;
      RECT 14.76 6.705 14.91 6.855 ;
      RECT 14.3 3.72 14.45 3.87 ;
      RECT 14.115 7.165 14.265 7.315 ;
      RECT 13.85 2.22 14 2.37 ;
      RECT 13.67 3.21 13.82 3.36 ;
      RECT 13.275 3.725 13.425 3.875 ;
      RECT 12.915 3.68 13.065 3.83 ;
      RECT 12.77 2.17 12.92 2.32 ;
      RECT 12.185 3.62 12.335 3.77 ;
      RECT 12.09 2.155 12.24 2.305 ;
      RECT 11.935 2.69 12.085 2.84 ;
      RECT 11.25 3.655 11.4 3.805 ;
      RECT 10.855 2.28 11.005 2.43 ;
      RECT 10.135 3.185 10.285 3.335 ;
      RECT 10.095 2.22 10.245 2.37 ;
      RECT 9.825 3.69 9.975 3.84 ;
      RECT 9.29 2.41 9.44 2.56 ;
      RECT 9.245 3.28 9.395 3.43 ;
      RECT 9.065 2.835 9.215 2.985 ;
      RECT 7.99 2.69 8.14 2.84 ;
      RECT 7.885 2.115 8.035 2.265 ;
      RECT 7.23 3.26 7.38 3.41 ;
      RECT 6.71 1.3 6.86 1.45 ;
      RECT 6.62 3.17 6.77 3.32 ;
      RECT 5.975 2.17 6.125 2.32 ;
      RECT 5.96 3.175 6.11 3.325 ;
      RECT 5.445 2.66 5.595 2.81 ;
      RECT 4.865 3.44 5.015 3.59 ;
      RECT 3.09 7.095 3.24 7.245 ;
      RECT 2.715 6.355 2.865 6.505 ;
    LAYER met1 ;
      RECT 76.345 1.285 88.305 1.89 ;
      RECT 80.77 0 88.305 1.89 ;
      RECT 58.42 1.285 70.38 1.89 ;
      RECT 62.845 0 70.38 1.89 ;
      RECT 40.495 1.285 52.455 1.89 ;
      RECT 44.92 0 52.455 1.89 ;
      RECT 22.57 1.285 34.53 1.89 ;
      RECT 26.995 0 34.53 1.89 ;
      RECT 4.645 1.285 16.605 1.89 ;
      RECT 9.07 0 16.605 1.89 ;
      RECT 76.34 0 77.085 1.68 ;
      RECT 58.415 0 59.16 1.68 ;
      RECT 40.49 0 41.235 1.68 ;
      RECT 22.565 0 23.31 1.68 ;
      RECT 4.64 0 5.385 1.68 ;
      RECT 79.335 0 80.49 1.89 ;
      RECT 76.34 1.255 79.055 1.68 ;
      RECT 77.365 0 79.055 1.89 ;
      RECT 61.41 0 62.565 1.89 ;
      RECT 58.415 1.255 61.13 1.68 ;
      RECT 59.44 0 61.13 1.89 ;
      RECT 43.485 0 44.64 1.89 ;
      RECT 40.49 1.255 43.205 1.68 ;
      RECT 41.515 0 43.205 1.89 ;
      RECT 25.56 0 26.715 1.89 ;
      RECT 22.565 1.255 25.28 1.68 ;
      RECT 23.59 0 25.28 1.89 ;
      RECT 7.635 0 8.79 1.89 ;
      RECT 4.64 1.255 7.355 1.68 ;
      RECT 5.665 0 7.355 1.89 ;
      RECT 77.365 0 88.305 1.005 ;
      RECT 59.44 0 70.38 1.005 ;
      RECT 41.515 0 52.455 1.005 ;
      RECT 23.59 0 34.53 1.005 ;
      RECT 5.665 0 16.605 1.005 ;
      RECT 76.34 0 88.305 0.975 ;
      RECT 58.415 0 70.38 0.975 ;
      RECT 40.49 0 52.455 0.975 ;
      RECT 22.565 0 34.53 0.975 ;
      RECT 4.64 0 16.605 0.975 ;
      RECT 93.715 0 93.895 0.305 ;
      RECT 75.79 0 91.765 0.305 ;
      RECT 57.865 0 73.84 0.305 ;
      RECT 39.94 0 55.915 0.305 ;
      RECT 22.015 0 37.99 0.305 ;
      RECT 1.48 0 20.065 0.305 ;
      RECT 1.48 0 93.895 0.3 ;
      RECT 1.46 8.58 93.895 8.88 ;
      RECT 93.715 8.575 93.895 8.88 ;
      RECT 75.79 8.575 91.765 8.88 ;
      RECT 57.865 8.575 73.84 8.88 ;
      RECT 39.94 8.575 55.915 8.88 ;
      RECT 22.015 8.575 37.99 8.88 ;
      RECT 1.46 8.575 20.065 8.88 ;
      RECT 85.04 6.315 85.21 8.88 ;
      RECT 67.115 6.315 67.285 8.88 ;
      RECT 49.19 6.315 49.36 8.88 ;
      RECT 31.265 6.315 31.435 8.88 ;
      RECT 13.34 6.315 13.51 8.88 ;
      RECT 85.375 6.285 85.665 6.515 ;
      RECT 67.45 6.285 67.74 6.515 ;
      RECT 49.525 6.285 49.815 6.515 ;
      RECT 31.6 6.285 31.89 6.515 ;
      RECT 13.675 6.285 13.965 6.515 ;
      RECT 85.04 6.315 85.665 6.485 ;
      RECT 67.115 6.315 67.74 6.485 ;
      RECT 49.19 6.315 49.815 6.485 ;
      RECT 31.265 6.315 31.89 6.485 ;
      RECT 13.34 6.315 13.965 6.485 ;
      RECT 93.29 7.77 93.58 8 ;
      RECT 93.35 6.29 93.52 8 ;
      RECT 93.32 7.275 93.67 7.625 ;
      RECT 93.29 6.29 93.58 6.52 ;
      RECT 92.885 2.395 92.99 2.965 ;
      RECT 92.885 2.73 93.21 2.96 ;
      RECT 92.885 2.76 93.38 2.93 ;
      RECT 92.885 2.395 93.075 2.96 ;
      RECT 92.3 2.36 92.59 2.59 ;
      RECT 92.3 2.395 93.075 2.565 ;
      RECT 92.36 0.88 92.53 2.59 ;
      RECT 92.3 0.88 92.59 1.11 ;
      RECT 92.3 7.77 92.59 8 ;
      RECT 92.36 6.29 92.53 8 ;
      RECT 92.3 6.29 92.59 6.52 ;
      RECT 92.3 6.325 93.155 6.485 ;
      RECT 92.985 5.92 93.155 6.485 ;
      RECT 92.3 6.32 92.695 6.485 ;
      RECT 92.92 5.92 93.21 6.15 ;
      RECT 92.92 5.95 93.38 6.12 ;
      RECT 91.93 2.73 92.22 2.96 ;
      RECT 91.93 2.76 92.39 2.93 ;
      RECT 91.995 1.655 92.16 2.96 ;
      RECT 90.51 1.625 90.8 1.855 ;
      RECT 90.51 1.655 92.16 1.825 ;
      RECT 90.57 0.885 90.74 1.855 ;
      RECT 90.51 0.885 90.8 1.115 ;
      RECT 90.51 7.765 90.8 7.995 ;
      RECT 90.57 7.025 90.74 7.995 ;
      RECT 90.57 7.12 92.16 7.29 ;
      RECT 91.99 5.92 92.16 7.29 ;
      RECT 90.51 7.025 90.8 7.255 ;
      RECT 91.93 5.92 92.22 6.15 ;
      RECT 91.93 5.95 92.39 6.12 ;
      RECT 88.545 3.43 88.895 3.78 ;
      RECT 88.635 2.025 88.805 3.78 ;
      RECT 90.94 1.965 91.29 2.315 ;
      RECT 88.635 2.025 90.255 2.2 ;
      RECT 88.635 2.025 91.29 2.195 ;
      RECT 90.965 6.655 91.29 6.98 ;
      RECT 86.62 6.61 86.97 6.96 ;
      RECT 90.94 6.655 91.29 6.885 ;
      RECT 86.18 6.655 86.47 6.885 ;
      RECT 86.01 6.685 91.29 6.855 ;
      RECT 90.165 2.365 90.485 2.685 ;
      RECT 90.135 2.365 90.485 2.595 ;
      RECT 89.965 2.395 90.485 2.565 ;
      RECT 90.165 6.225 90.485 6.545 ;
      RECT 90.135 6.285 90.485 6.515 ;
      RECT 89.965 6.315 90.485 6.485 ;
      RECT 85.945 3.665 85.985 3.925 ;
      RECT 85.985 3.645 85.99 3.655 ;
      RECT 87.315 2.89 87.325 3.111 ;
      RECT 87.245 2.885 87.315 3.236 ;
      RECT 87.235 2.885 87.245 3.363 ;
      RECT 87.21 2.885 87.235 3.41 ;
      RECT 87.185 2.885 87.21 3.488 ;
      RECT 87.165 2.885 87.185 3.558 ;
      RECT 87.14 2.885 87.165 3.598 ;
      RECT 87.13 2.885 87.14 3.618 ;
      RECT 87.12 2.887 87.13 3.626 ;
      RECT 87.115 2.892 87.12 3.083 ;
      RECT 87.115 3.092 87.12 3.627 ;
      RECT 87.11 3.137 87.115 3.628 ;
      RECT 87.1 3.202 87.11 3.629 ;
      RECT 87.09 3.297 87.1 3.631 ;
      RECT 87.085 3.35 87.09 3.633 ;
      RECT 87.08 3.37 87.085 3.634 ;
      RECT 87.025 3.395 87.08 3.64 ;
      RECT 86.985 3.43 87.025 3.649 ;
      RECT 86.975 3.447 86.985 3.654 ;
      RECT 86.966 3.453 86.975 3.656 ;
      RECT 86.88 3.491 86.966 3.667 ;
      RECT 86.875 3.53 86.88 3.677 ;
      RECT 86.8 3.537 86.875 3.687 ;
      RECT 86.78 3.547 86.8 3.698 ;
      RECT 86.75 3.554 86.78 3.706 ;
      RECT 86.725 3.561 86.75 3.713 ;
      RECT 86.701 3.567 86.725 3.718 ;
      RECT 86.615 3.58 86.701 3.73 ;
      RECT 86.537 3.587 86.615 3.748 ;
      RECT 86.451 3.582 86.537 3.766 ;
      RECT 86.365 3.577 86.451 3.786 ;
      RECT 86.285 3.571 86.365 3.803 ;
      RECT 86.22 3.567 86.285 3.832 ;
      RECT 86.215 3.281 86.22 3.305 ;
      RECT 86.205 3.557 86.22 3.86 ;
      RECT 86.21 3.275 86.215 3.345 ;
      RECT 86.205 3.269 86.21 3.415 ;
      RECT 86.2 3.263 86.205 3.493 ;
      RECT 86.2 3.54 86.205 3.925 ;
      RECT 86.192 3.26 86.2 3.925 ;
      RECT 86.106 3.258 86.192 3.925 ;
      RECT 86.02 3.256 86.106 3.925 ;
      RECT 86.01 3.257 86.02 3.925 ;
      RECT 86.005 3.262 86.01 3.925 ;
      RECT 85.995 3.275 86.005 3.925 ;
      RECT 85.99 3.297 85.995 3.925 ;
      RECT 85.985 3.657 85.99 3.925 ;
      RECT 86.615 3.125 86.62 3.345 ;
      RECT 87.12 2.16 87.155 2.42 ;
      RECT 87.105 2.16 87.12 2.428 ;
      RECT 87.076 2.16 87.105 2.45 ;
      RECT 86.99 2.16 87.076 2.51 ;
      RECT 86.97 2.16 86.99 2.575 ;
      RECT 86.91 2.16 86.97 2.74 ;
      RECT 86.905 2.16 86.91 2.888 ;
      RECT 86.9 2.16 86.905 2.9 ;
      RECT 86.895 2.16 86.9 2.926 ;
      RECT 86.865 2.346 86.895 3.006 ;
      RECT 86.86 2.394 86.865 3.095 ;
      RECT 86.855 2.408 86.86 3.11 ;
      RECT 86.85 2.427 86.855 3.14 ;
      RECT 86.845 2.442 86.85 3.156 ;
      RECT 86.84 2.457 86.845 3.178 ;
      RECT 86.835 2.477 86.84 3.2 ;
      RECT 86.825 2.497 86.835 3.233 ;
      RECT 86.81 2.539 86.825 3.295 ;
      RECT 86.805 2.57 86.81 3.335 ;
      RECT 86.8 2.582 86.805 3.34 ;
      RECT 86.795 2.594 86.8 3.345 ;
      RECT 86.79 2.607 86.795 3.345 ;
      RECT 86.785 2.625 86.79 3.345 ;
      RECT 86.78 2.645 86.785 3.345 ;
      RECT 86.775 2.657 86.78 3.345 ;
      RECT 86.77 2.67 86.775 3.345 ;
      RECT 86.75 2.705 86.77 3.345 ;
      RECT 86.7 2.807 86.75 3.345 ;
      RECT 86.695 2.892 86.7 3.345 ;
      RECT 86.69 2.9 86.695 3.345 ;
      RECT 86.685 2.917 86.69 3.345 ;
      RECT 86.68 2.932 86.685 3.345 ;
      RECT 86.645 2.997 86.68 3.345 ;
      RECT 86.63 3.062 86.645 3.345 ;
      RECT 86.625 3.092 86.63 3.345 ;
      RECT 86.62 3.117 86.625 3.345 ;
      RECT 86.605 3.127 86.615 3.345 ;
      RECT 86.59 3.14 86.605 3.338 ;
      RECT 86.335 2.73 86.405 2.94 ;
      RECT 86.125 2.707 86.13 2.9 ;
      RECT 83.58 2.635 83.84 2.895 ;
      RECT 86.415 2.917 86.42 2.92 ;
      RECT 86.405 2.735 86.415 2.935 ;
      RECT 86.306 2.728 86.335 2.94 ;
      RECT 86.22 2.72 86.306 2.94 ;
      RECT 86.205 2.714 86.22 2.938 ;
      RECT 86.185 2.713 86.205 2.925 ;
      RECT 86.18 2.712 86.185 2.908 ;
      RECT 86.13 2.709 86.18 2.903 ;
      RECT 86.1 2.706 86.125 2.898 ;
      RECT 86.08 2.704 86.1 2.893 ;
      RECT 86.065 2.702 86.08 2.89 ;
      RECT 86.035 2.7 86.065 2.888 ;
      RECT 85.97 2.696 86.035 2.88 ;
      RECT 85.94 2.691 85.97 2.875 ;
      RECT 85.92 2.689 85.94 2.873 ;
      RECT 85.89 2.686 85.92 2.868 ;
      RECT 85.83 2.682 85.89 2.86 ;
      RECT 85.825 2.679 85.83 2.855 ;
      RECT 85.755 2.677 85.825 2.85 ;
      RECT 85.726 2.673 85.755 2.843 ;
      RECT 85.64 2.668 85.726 2.835 ;
      RECT 85.606 2.663 85.64 2.827 ;
      RECT 85.52 2.655 85.606 2.819 ;
      RECT 85.481 2.648 85.52 2.811 ;
      RECT 85.395 2.643 85.481 2.803 ;
      RECT 85.33 2.637 85.395 2.793 ;
      RECT 85.31 2.632 85.33 2.788 ;
      RECT 85.301 2.629 85.31 2.787 ;
      RECT 85.215 2.625 85.301 2.781 ;
      RECT 85.175 2.621 85.215 2.773 ;
      RECT 85.155 2.617 85.175 2.771 ;
      RECT 85.095 2.617 85.155 2.768 ;
      RECT 85.075 2.62 85.095 2.766 ;
      RECT 85.054 2.62 85.075 2.766 ;
      RECT 84.968 2.622 85.054 2.77 ;
      RECT 84.882 2.624 84.968 2.776 ;
      RECT 84.796 2.626 84.882 2.783 ;
      RECT 84.71 2.629 84.796 2.789 ;
      RECT 84.676 2.63 84.71 2.794 ;
      RECT 84.59 2.633 84.676 2.799 ;
      RECT 84.561 2.64 84.59 2.804 ;
      RECT 84.475 2.64 84.561 2.809 ;
      RECT 84.442 2.64 84.475 2.814 ;
      RECT 84.356 2.642 84.442 2.819 ;
      RECT 84.27 2.644 84.356 2.826 ;
      RECT 84.206 2.646 84.27 2.832 ;
      RECT 84.12 2.648 84.206 2.838 ;
      RECT 84.117 2.65 84.12 2.841 ;
      RECT 84.031 2.651 84.117 2.845 ;
      RECT 83.945 2.654 84.031 2.852 ;
      RECT 83.926 2.656 83.945 2.856 ;
      RECT 83.84 2.658 83.926 2.861 ;
      RECT 83.57 2.67 83.58 2.865 ;
      RECT 85.75 7.765 86.04 7.995 ;
      RECT 85.81 7.025 85.98 7.995 ;
      RECT 85.7 7.055 86.075 7.425 ;
      RECT 85.75 7.025 86.04 7.425 ;
      RECT 85.805 2.25 85.99 2.46 ;
      RECT 85.8 2.251 85.995 2.458 ;
      RECT 85.795 2.256 86.005 2.453 ;
      RECT 85.79 2.232 85.795 2.45 ;
      RECT 85.76 2.229 85.79 2.443 ;
      RECT 85.755 2.225 85.76 2.434 ;
      RECT 85.72 2.256 86.005 2.429 ;
      RECT 85.495 2.165 85.755 2.425 ;
      RECT 85.795 2.234 85.8 2.453 ;
      RECT 85.8 2.235 85.805 2.458 ;
      RECT 85.495 2.247 85.875 2.425 ;
      RECT 85.495 2.245 85.86 2.425 ;
      RECT 85.495 2.24 85.85 2.425 ;
      RECT 85.45 3.155 85.5 3.44 ;
      RECT 85.395 3.125 85.4 3.44 ;
      RECT 85.365 3.105 85.37 3.44 ;
      RECT 85.515 3.155 85.575 3.415 ;
      RECT 85.51 3.155 85.515 3.423 ;
      RECT 85.5 3.155 85.51 3.435 ;
      RECT 85.415 3.145 85.45 3.44 ;
      RECT 85.41 3.132 85.415 3.44 ;
      RECT 85.4 3.127 85.41 3.44 ;
      RECT 85.38 3.117 85.395 3.44 ;
      RECT 85.37 3.11 85.38 3.44 ;
      RECT 85.36 3.102 85.365 3.44 ;
      RECT 85.33 3.092 85.36 3.44 ;
      RECT 85.315 3.08 85.33 3.44 ;
      RECT 85.3 3.07 85.315 3.435 ;
      RECT 85.28 3.06 85.3 3.41 ;
      RECT 85.27 3.052 85.28 3.387 ;
      RECT 85.24 3.035 85.27 3.377 ;
      RECT 85.235 3.012 85.24 3.368 ;
      RECT 85.23 2.999 85.235 3.366 ;
      RECT 85.215 2.975 85.23 3.36 ;
      RECT 85.21 2.951 85.215 3.354 ;
      RECT 85.2 2.94 85.21 3.349 ;
      RECT 85.195 2.93 85.2 3.345 ;
      RECT 85.19 2.922 85.195 3.342 ;
      RECT 85.18 2.917 85.19 3.338 ;
      RECT 85.175 2.912 85.18 3.334 ;
      RECT 85.09 2.91 85.175 3.309 ;
      RECT 85.06 2.91 85.09 3.275 ;
      RECT 85.045 2.91 85.06 3.258 ;
      RECT 84.99 2.91 85.045 3.203 ;
      RECT 84.985 2.915 84.99 3.152 ;
      RECT 84.975 2.92 84.985 3.142 ;
      RECT 84.97 2.93 84.975 3.128 ;
      RECT 84.92 3.67 85.18 3.93 ;
      RECT 84.84 3.685 85.18 3.906 ;
      RECT 84.82 3.685 85.18 3.901 ;
      RECT 84.796 3.685 85.18 3.899 ;
      RECT 84.71 3.685 85.18 3.894 ;
      RECT 84.56 3.625 84.82 3.89 ;
      RECT 84.515 3.685 85.18 3.885 ;
      RECT 84.51 3.692 85.18 3.88 ;
      RECT 84.525 3.68 84.84 3.89 ;
      RECT 84.415 2.115 84.675 2.375 ;
      RECT 84.415 2.172 84.68 2.368 ;
      RECT 84.415 2.202 84.685 2.3 ;
      RECT 84.475 2.633 84.59 2.635 ;
      RECT 84.561 2.63 84.59 2.635 ;
      RECT 83.585 3.634 83.61 3.874 ;
      RECT 83.57 3.637 83.66 3.868 ;
      RECT 83.565 3.642 83.746 3.863 ;
      RECT 83.56 3.65 83.81 3.861 ;
      RECT 83.56 3.65 83.82 3.86 ;
      RECT 83.555 3.657 83.83 3.853 ;
      RECT 83.555 3.657 83.916 3.842 ;
      RECT 83.55 3.692 83.916 3.838 ;
      RECT 83.55 3.692 83.925 3.827 ;
      RECT 83.83 3.565 84.09 3.825 ;
      RECT 83.54 3.742 84.09 3.823 ;
      RECT 83.81 3.61 83.83 3.858 ;
      RECT 83.746 3.613 83.81 3.862 ;
      RECT 83.66 3.618 83.746 3.867 ;
      RECT 83.59 3.629 84.09 3.825 ;
      RECT 83.61 3.623 83.66 3.872 ;
      RECT 83.735 2.1 83.745 2.362 ;
      RECT 83.725 2.157 83.735 2.365 ;
      RECT 83.7 2.162 83.725 2.371 ;
      RECT 83.675 2.166 83.7 2.383 ;
      RECT 83.665 2.169 83.675 2.393 ;
      RECT 83.66 2.17 83.665 2.398 ;
      RECT 83.655 2.171 83.66 2.403 ;
      RECT 83.65 2.172 83.655 2.405 ;
      RECT 83.625 2.175 83.65 2.408 ;
      RECT 83.595 2.181 83.625 2.411 ;
      RECT 83.53 2.192 83.595 2.414 ;
      RECT 83.485 2.2 83.53 2.418 ;
      RECT 83.47 2.2 83.485 2.426 ;
      RECT 83.465 2.201 83.47 2.433 ;
      RECT 83.46 2.203 83.465 2.436 ;
      RECT 83.455 2.207 83.46 2.439 ;
      RECT 83.445 2.215 83.455 2.443 ;
      RECT 83.44 2.228 83.445 2.448 ;
      RECT 83.435 2.236 83.44 2.45 ;
      RECT 83.43 2.242 83.435 2.45 ;
      RECT 83.425 2.246 83.43 2.453 ;
      RECT 83.42 2.248 83.425 2.456 ;
      RECT 83.415 2.251 83.42 2.459 ;
      RECT 83.405 2.256 83.415 2.463 ;
      RECT 83.4 2.262 83.405 2.468 ;
      RECT 83.39 2.268 83.4 2.472 ;
      RECT 83.375 2.275 83.39 2.478 ;
      RECT 83.346 2.289 83.375 2.488 ;
      RECT 83.26 2.324 83.346 2.52 ;
      RECT 83.24 2.357 83.26 2.549 ;
      RECT 83.22 2.37 83.24 2.56 ;
      RECT 83.2 2.382 83.22 2.571 ;
      RECT 83.15 2.404 83.2 2.591 ;
      RECT 83.135 2.422 83.15 2.608 ;
      RECT 83.13 2.428 83.135 2.611 ;
      RECT 83.125 2.432 83.13 2.614 ;
      RECT 83.12 2.436 83.125 2.618 ;
      RECT 83.115 2.438 83.12 2.621 ;
      RECT 83.105 2.445 83.115 2.624 ;
      RECT 83.1 2.45 83.105 2.628 ;
      RECT 83.095 2.452 83.1 2.631 ;
      RECT 83.09 2.456 83.095 2.634 ;
      RECT 83.085 2.458 83.09 2.638 ;
      RECT 83.07 2.463 83.085 2.643 ;
      RECT 83.065 2.468 83.07 2.646 ;
      RECT 83.06 2.476 83.065 2.649 ;
      RECT 83.055 2.478 83.06 2.652 ;
      RECT 83.05 2.48 83.055 2.655 ;
      RECT 83.04 2.482 83.05 2.661 ;
      RECT 83.005 2.496 83.04 2.673 ;
      RECT 82.995 2.511 83.005 2.683 ;
      RECT 82.92 2.54 82.995 2.707 ;
      RECT 82.915 2.565 82.92 2.73 ;
      RECT 82.9 2.569 82.915 2.736 ;
      RECT 82.89 2.577 82.9 2.741 ;
      RECT 82.86 2.59 82.89 2.745 ;
      RECT 82.85 2.605 82.86 2.75 ;
      RECT 82.84 2.61 82.85 2.753 ;
      RECT 82.835 2.612 82.84 2.755 ;
      RECT 82.82 2.615 82.835 2.758 ;
      RECT 82.815 2.617 82.82 2.761 ;
      RECT 82.795 2.622 82.815 2.765 ;
      RECT 82.765 2.627 82.795 2.773 ;
      RECT 82.74 2.634 82.765 2.781 ;
      RECT 82.735 2.639 82.74 2.786 ;
      RECT 82.705 2.642 82.735 2.79 ;
      RECT 82.665 2.645 82.705 2.8 ;
      RECT 82.63 2.642 82.665 2.812 ;
      RECT 82.62 2.638 82.63 2.819 ;
      RECT 82.595 2.634 82.62 2.825 ;
      RECT 82.59 2.63 82.595 2.83 ;
      RECT 82.55 2.627 82.59 2.83 ;
      RECT 82.535 2.612 82.55 2.831 ;
      RECT 82.512 2.6 82.535 2.831 ;
      RECT 82.426 2.6 82.512 2.832 ;
      RECT 82.34 2.6 82.426 2.834 ;
      RECT 82.32 2.6 82.34 2.831 ;
      RECT 82.315 2.605 82.32 2.826 ;
      RECT 82.31 2.61 82.315 2.824 ;
      RECT 82.3 2.62 82.31 2.822 ;
      RECT 82.295 2.626 82.3 2.815 ;
      RECT 82.29 2.628 82.295 2.8 ;
      RECT 82.285 2.632 82.29 2.79 ;
      RECT 83.745 2.1 83.995 2.36 ;
      RECT 81.47 3.635 81.73 3.895 ;
      RECT 83.765 3.125 83.77 3.335 ;
      RECT 83.77 3.13 83.78 3.33 ;
      RECT 83.72 3.125 83.765 3.35 ;
      RECT 83.71 3.125 83.72 3.37 ;
      RECT 83.691 3.125 83.71 3.375 ;
      RECT 83.605 3.125 83.691 3.372 ;
      RECT 83.575 3.127 83.605 3.37 ;
      RECT 83.52 3.137 83.575 3.368 ;
      RECT 83.455 3.151 83.52 3.366 ;
      RECT 83.45 3.159 83.455 3.365 ;
      RECT 83.435 3.162 83.45 3.363 ;
      RECT 83.37 3.172 83.435 3.359 ;
      RECT 83.322 3.186 83.37 3.36 ;
      RECT 83.236 3.203 83.322 3.374 ;
      RECT 83.15 3.224 83.236 3.391 ;
      RECT 83.13 3.237 83.15 3.401 ;
      RECT 83.085 3.245 83.13 3.408 ;
      RECT 83.05 3.253 83.085 3.416 ;
      RECT 83.016 3.261 83.05 3.424 ;
      RECT 82.93 3.275 83.016 3.436 ;
      RECT 82.895 3.292 82.93 3.448 ;
      RECT 82.886 3.301 82.895 3.452 ;
      RECT 82.8 3.319 82.886 3.469 ;
      RECT 82.741 3.346 82.8 3.496 ;
      RECT 82.655 3.373 82.741 3.524 ;
      RECT 82.635 3.395 82.655 3.544 ;
      RECT 82.575 3.41 82.635 3.56 ;
      RECT 82.565 3.422 82.575 3.573 ;
      RECT 82.56 3.427 82.565 3.576 ;
      RECT 82.55 3.43 82.56 3.579 ;
      RECT 82.545 3.432 82.55 3.582 ;
      RECT 82.515 3.44 82.545 3.589 ;
      RECT 82.5 3.447 82.515 3.597 ;
      RECT 82.49 3.452 82.5 3.601 ;
      RECT 82.485 3.455 82.49 3.604 ;
      RECT 82.475 3.457 82.485 3.607 ;
      RECT 82.44 3.467 82.475 3.616 ;
      RECT 82.365 3.49 82.44 3.638 ;
      RECT 82.345 3.508 82.365 3.656 ;
      RECT 82.315 3.515 82.345 3.666 ;
      RECT 82.295 3.523 82.315 3.676 ;
      RECT 82.285 3.529 82.295 3.683 ;
      RECT 82.266 3.534 82.285 3.689 ;
      RECT 82.18 3.554 82.266 3.709 ;
      RECT 82.165 3.574 82.18 3.728 ;
      RECT 82.12 3.586 82.165 3.739 ;
      RECT 82.055 3.607 82.12 3.762 ;
      RECT 82.015 3.627 82.055 3.783 ;
      RECT 82.005 3.637 82.015 3.793 ;
      RECT 81.955 3.649 82.005 3.804 ;
      RECT 81.935 3.665 81.955 3.816 ;
      RECT 81.905 3.675 81.935 3.822 ;
      RECT 81.895 3.68 81.905 3.824 ;
      RECT 81.826 3.681 81.895 3.83 ;
      RECT 81.74 3.683 81.826 3.84 ;
      RECT 81.73 3.684 81.74 3.845 ;
      RECT 83 3.71 83.19 3.92 ;
      RECT 82.99 3.715 83.2 3.913 ;
      RECT 82.975 3.715 83.2 3.878 ;
      RECT 82.895 3.6 83.155 3.86 ;
      RECT 81.81 3.13 81.995 3.425 ;
      RECT 81.8 3.13 81.995 3.423 ;
      RECT 81.785 3.13 82 3.418 ;
      RECT 81.785 3.13 82.005 3.415 ;
      RECT 81.78 3.13 82.005 3.413 ;
      RECT 81.775 3.385 82.005 3.403 ;
      RECT 81.78 3.13 82.04 3.39 ;
      RECT 81.74 2.165 82 2.425 ;
      RECT 81.55 2.09 81.636 2.423 ;
      RECT 81.525 2.094 81.68 2.419 ;
      RECT 81.636 2.086 81.68 2.419 ;
      RECT 81.636 2.087 81.685 2.418 ;
      RECT 81.55 2.092 81.7 2.417 ;
      RECT 81.525 2.1 81.74 2.416 ;
      RECT 81.52 2.095 81.7 2.411 ;
      RECT 81.51 2.11 81.74 2.318 ;
      RECT 81.51 2.162 81.94 2.318 ;
      RECT 81.51 2.155 81.92 2.318 ;
      RECT 81.51 2.142 81.89 2.318 ;
      RECT 81.51 2.13 81.83 2.318 ;
      RECT 81.51 2.115 81.805 2.318 ;
      RECT 80.71 2.745 80.845 3.04 ;
      RECT 80.97 2.768 80.975 2.955 ;
      RECT 81.69 2.665 81.835 2.9 ;
      RECT 81.85 2.665 81.855 2.89 ;
      RECT 81.885 2.676 81.89 2.87 ;
      RECT 81.88 2.668 81.885 2.875 ;
      RECT 81.86 2.665 81.88 2.88 ;
      RECT 81.855 2.665 81.86 2.888 ;
      RECT 81.845 2.665 81.85 2.893 ;
      RECT 81.835 2.665 81.845 2.898 ;
      RECT 81.665 2.667 81.69 2.9 ;
      RECT 81.615 2.674 81.665 2.9 ;
      RECT 81.61 2.679 81.615 2.9 ;
      RECT 81.571 2.684 81.61 2.901 ;
      RECT 81.485 2.696 81.571 2.902 ;
      RECT 81.476 2.706 81.485 2.902 ;
      RECT 81.39 2.715 81.476 2.904 ;
      RECT 81.366 2.725 81.39 2.906 ;
      RECT 81.28 2.736 81.366 2.907 ;
      RECT 81.25 2.747 81.28 2.909 ;
      RECT 81.22 2.752 81.25 2.911 ;
      RECT 81.195 2.758 81.22 2.914 ;
      RECT 81.18 2.763 81.195 2.915 ;
      RECT 81.135 2.769 81.18 2.915 ;
      RECT 81.13 2.774 81.135 2.916 ;
      RECT 81.11 2.774 81.13 2.918 ;
      RECT 81.09 2.772 81.11 2.923 ;
      RECT 81.055 2.771 81.09 2.93 ;
      RECT 81.025 2.77 81.055 2.94 ;
      RECT 80.975 2.769 81.025 2.95 ;
      RECT 80.885 2.766 80.97 3.04 ;
      RECT 80.86 2.76 80.885 3.04 ;
      RECT 80.845 2.75 80.86 3.04 ;
      RECT 80.66 2.745 80.71 2.96 ;
      RECT 80.65 2.75 80.66 2.95 ;
      RECT 80.89 3.225 81.15 3.485 ;
      RECT 80.89 3.225 81.18 3.378 ;
      RECT 80.89 3.225 81.215 3.363 ;
      RECT 81.145 3.145 81.335 3.355 ;
      RECT 81.135 3.15 81.345 3.348 ;
      RECT 81.1 3.22 81.345 3.348 ;
      RECT 81.13 3.162 81.15 3.485 ;
      RECT 81.115 3.21 81.345 3.348 ;
      RECT 81.12 3.182 81.15 3.485 ;
      RECT 80.2 2.25 80.27 3.355 ;
      RECT 80.935 2.355 81.195 2.615 ;
      RECT 80.515 2.401 80.53 2.61 ;
      RECT 80.851 2.414 80.935 2.565 ;
      RECT 80.765 2.411 80.851 2.565 ;
      RECT 80.726 2.409 80.765 2.565 ;
      RECT 80.64 2.407 80.726 2.565 ;
      RECT 80.58 2.405 80.64 2.576 ;
      RECT 80.545 2.403 80.58 2.594 ;
      RECT 80.53 2.401 80.545 2.605 ;
      RECT 80.5 2.401 80.515 2.618 ;
      RECT 80.49 2.401 80.5 2.623 ;
      RECT 80.465 2.4 80.49 2.628 ;
      RECT 80.45 2.395 80.465 2.634 ;
      RECT 80.445 2.388 80.45 2.639 ;
      RECT 80.42 2.379 80.445 2.645 ;
      RECT 80.375 2.358 80.42 2.658 ;
      RECT 80.365 2.342 80.375 2.668 ;
      RECT 80.35 2.335 80.365 2.678 ;
      RECT 80.34 2.328 80.35 2.695 ;
      RECT 80.335 2.325 80.34 2.725 ;
      RECT 80.33 2.323 80.335 2.755 ;
      RECT 80.325 2.321 80.33 2.792 ;
      RECT 80.31 2.317 80.325 2.859 ;
      RECT 80.31 3.15 80.32 3.35 ;
      RECT 80.305 2.313 80.31 2.985 ;
      RECT 80.305 3.137 80.31 3.355 ;
      RECT 80.3 2.311 80.305 3.07 ;
      RECT 80.3 3.127 80.305 3.355 ;
      RECT 80.285 2.282 80.3 3.355 ;
      RECT 80.27 2.255 80.285 3.355 ;
      RECT 80.195 2.25 80.2 2.605 ;
      RECT 80.195 2.66 80.2 3.355 ;
      RECT 80.18 2.25 80.195 2.583 ;
      RECT 80.19 2.682 80.195 3.355 ;
      RECT 80.18 2.722 80.19 3.355 ;
      RECT 80.145 2.25 80.18 2.525 ;
      RECT 80.175 2.757 80.18 3.355 ;
      RECT 80.16 2.812 80.175 3.355 ;
      RECT 80.155 2.877 80.16 3.355 ;
      RECT 80.14 2.925 80.155 3.355 ;
      RECT 80.115 2.25 80.145 2.48 ;
      RECT 80.135 2.98 80.14 3.355 ;
      RECT 80.12 3.04 80.135 3.355 ;
      RECT 80.115 3.088 80.12 3.353 ;
      RECT 80.11 2.25 80.115 2.473 ;
      RECT 80.11 3.12 80.115 3.348 ;
      RECT 80.085 2.25 80.11 2.465 ;
      RECT 80.075 2.255 80.085 2.455 ;
      RECT 80.29 3.53 80.31 3.77 ;
      RECT 79.52 3.46 79.525 3.67 ;
      RECT 80.8 3.533 80.81 3.728 ;
      RECT 80.795 3.523 80.8 3.731 ;
      RECT 80.715 3.52 80.795 3.754 ;
      RECT 80.711 3.52 80.715 3.776 ;
      RECT 80.625 3.52 80.711 3.786 ;
      RECT 80.61 3.52 80.625 3.794 ;
      RECT 80.581 3.521 80.61 3.792 ;
      RECT 80.495 3.526 80.581 3.788 ;
      RECT 80.482 3.53 80.495 3.784 ;
      RECT 80.396 3.53 80.482 3.78 ;
      RECT 80.31 3.53 80.396 3.774 ;
      RECT 80.226 3.53 80.29 3.768 ;
      RECT 80.14 3.53 80.226 3.763 ;
      RECT 80.12 3.53 80.14 3.759 ;
      RECT 80.06 3.525 80.12 3.756 ;
      RECT 80.032 3.519 80.06 3.753 ;
      RECT 79.946 3.514 80.032 3.749 ;
      RECT 79.86 3.508 79.946 3.743 ;
      RECT 79.785 3.49 79.86 3.738 ;
      RECT 79.75 3.467 79.785 3.734 ;
      RECT 79.74 3.457 79.75 3.733 ;
      RECT 79.685 3.455 79.74 3.732 ;
      RECT 79.61 3.455 79.685 3.728 ;
      RECT 79.6 3.455 79.61 3.723 ;
      RECT 79.585 3.455 79.6 3.715 ;
      RECT 79.535 3.457 79.585 3.693 ;
      RECT 79.525 3.46 79.535 3.673 ;
      RECT 79.515 3.465 79.52 3.668 ;
      RECT 79.51 3.47 79.515 3.663 ;
      RECT 79.635 2.635 79.895 2.895 ;
      RECT 79.635 2.65 79.915 2.86 ;
      RECT 79.635 2.655 79.925 2.855 ;
      RECT 77.62 2.115 77.88 2.375 ;
      RECT 77.61 2.145 77.88 2.355 ;
      RECT 79.53 2.06 79.79 2.32 ;
      RECT 79.525 2.135 79.53 2.321 ;
      RECT 79.5 2.14 79.525 2.323 ;
      RECT 79.485 2.147 79.5 2.326 ;
      RECT 79.425 2.165 79.485 2.331 ;
      RECT 79.395 2.185 79.425 2.338 ;
      RECT 79.37 2.193 79.395 2.343 ;
      RECT 79.345 2.201 79.37 2.345 ;
      RECT 79.327 2.205 79.345 2.344 ;
      RECT 79.241 2.203 79.327 2.344 ;
      RECT 79.155 2.201 79.241 2.344 ;
      RECT 79.069 2.199 79.155 2.343 ;
      RECT 78.983 2.197 79.069 2.343 ;
      RECT 78.897 2.195 78.983 2.343 ;
      RECT 78.811 2.193 78.897 2.343 ;
      RECT 78.725 2.191 78.811 2.342 ;
      RECT 78.707 2.19 78.725 2.342 ;
      RECT 78.621 2.189 78.707 2.342 ;
      RECT 78.535 2.187 78.621 2.342 ;
      RECT 78.449 2.186 78.535 2.341 ;
      RECT 78.363 2.185 78.449 2.341 ;
      RECT 78.277 2.183 78.363 2.341 ;
      RECT 78.191 2.182 78.277 2.341 ;
      RECT 78.105 2.18 78.191 2.34 ;
      RECT 78.081 2.178 78.105 2.34 ;
      RECT 77.995 2.171 78.081 2.34 ;
      RECT 77.966 2.163 77.995 2.34 ;
      RECT 77.88 2.155 77.966 2.34 ;
      RECT 77.6 2.152 77.61 2.35 ;
      RECT 79.105 3.115 79.11 3.465 ;
      RECT 78.875 3.205 79.015 3.465 ;
      RECT 79.35 2.89 79.395 3.1 ;
      RECT 79.405 2.901 79.415 3.095 ;
      RECT 79.395 2.893 79.405 3.1 ;
      RECT 79.33 2.89 79.35 3.105 ;
      RECT 79.3 2.89 79.33 3.128 ;
      RECT 79.29 2.89 79.3 3.153 ;
      RECT 79.285 2.89 79.29 3.163 ;
      RECT 79.23 2.89 79.285 3.203 ;
      RECT 79.225 2.89 79.23 3.243 ;
      RECT 79.22 2.892 79.225 3.248 ;
      RECT 79.205 2.902 79.22 3.259 ;
      RECT 79.16 2.96 79.205 3.295 ;
      RECT 79.15 3.015 79.16 3.329 ;
      RECT 79.135 3.042 79.15 3.345 ;
      RECT 79.125 3.069 79.135 3.465 ;
      RECT 79.11 3.092 79.125 3.465 ;
      RECT 79.1 3.132 79.105 3.465 ;
      RECT 79.095 3.142 79.1 3.465 ;
      RECT 79.09 3.157 79.095 3.465 ;
      RECT 79.08 3.162 79.09 3.465 ;
      RECT 79.015 3.185 79.08 3.465 ;
      RECT 78.515 2.68 78.705 2.89 ;
      RECT 77.09 2.605 77.35 2.865 ;
      RECT 77.44 2.6 77.535 2.81 ;
      RECT 77.415 2.615 77.425 2.81 ;
      RECT 78.705 2.687 78.715 2.885 ;
      RECT 78.505 2.687 78.515 2.885 ;
      RECT 78.49 2.702 78.505 2.875 ;
      RECT 78.485 2.71 78.49 2.868 ;
      RECT 78.475 2.713 78.485 2.865 ;
      RECT 78.44 2.712 78.475 2.863 ;
      RECT 78.411 2.708 78.44 2.86 ;
      RECT 78.325 2.703 78.411 2.857 ;
      RECT 78.265 2.697 78.325 2.853 ;
      RECT 78.236 2.693 78.265 2.85 ;
      RECT 78.15 2.685 78.236 2.847 ;
      RECT 78.141 2.679 78.15 2.845 ;
      RECT 78.055 2.674 78.141 2.843 ;
      RECT 78.032 2.669 78.055 2.84 ;
      RECT 77.946 2.663 78.032 2.837 ;
      RECT 77.86 2.654 77.946 2.832 ;
      RECT 77.85 2.649 77.86 2.83 ;
      RECT 77.831 2.648 77.85 2.829 ;
      RECT 77.745 2.643 77.831 2.825 ;
      RECT 77.725 2.638 77.745 2.821 ;
      RECT 77.665 2.633 77.725 2.818 ;
      RECT 77.64 2.623 77.665 2.816 ;
      RECT 77.635 2.616 77.64 2.815 ;
      RECT 77.625 2.607 77.635 2.814 ;
      RECT 77.621 2.6 77.625 2.814 ;
      RECT 77.535 2.6 77.621 2.812 ;
      RECT 77.425 2.607 77.44 2.81 ;
      RECT 77.41 2.617 77.415 2.81 ;
      RECT 77.39 2.62 77.41 2.807 ;
      RECT 77.36 2.62 77.39 2.803 ;
      RECT 77.35 2.62 77.36 2.803 ;
      RECT 78.265 3.115 78.525 3.375 ;
      RECT 78.195 3.125 78.525 3.335 ;
      RECT 78.185 3.132 78.525 3.33 ;
      RECT 77.605 3.12 77.865 3.38 ;
      RECT 77.605 3.16 77.97 3.37 ;
      RECT 77.605 3.162 77.975 3.369 ;
      RECT 77.605 3.17 77.98 3.366 ;
      RECT 76.53 2.245 76.63 3.77 ;
      RECT 76.72 3.385 76.77 3.645 ;
      RECT 76.715 2.258 76.72 2.445 ;
      RECT 76.71 3.366 76.72 3.645 ;
      RECT 76.71 2.255 76.715 2.453 ;
      RECT 76.695 2.249 76.71 2.46 ;
      RECT 76.705 3.354 76.71 3.728 ;
      RECT 76.695 3.342 76.705 3.765 ;
      RECT 76.685 2.245 76.695 2.467 ;
      RECT 76.685 3.327 76.695 3.77 ;
      RECT 76.68 2.245 76.685 2.475 ;
      RECT 76.66 3.297 76.685 3.77 ;
      RECT 76.64 2.245 76.68 2.523 ;
      RECT 76.65 3.257 76.66 3.77 ;
      RECT 76.64 3.212 76.65 3.77 ;
      RECT 76.635 2.245 76.64 2.593 ;
      RECT 76.635 3.17 76.64 3.77 ;
      RECT 76.63 2.245 76.635 3.07 ;
      RECT 76.63 3.152 76.635 3.77 ;
      RECT 76.52 2.248 76.53 3.77 ;
      RECT 76.505 2.255 76.52 3.766 ;
      RECT 76.5 2.265 76.505 3.761 ;
      RECT 76.495 2.465 76.5 3.653 ;
      RECT 76.49 2.55 76.495 3.205 ;
      RECT 75.365 7.77 75.655 8 ;
      RECT 75.425 6.29 75.595 8 ;
      RECT 75.375 6.655 75.725 7.005 ;
      RECT 75.365 6.29 75.655 6.52 ;
      RECT 74.96 2.395 75.065 2.965 ;
      RECT 74.96 2.73 75.285 2.96 ;
      RECT 74.96 2.76 75.455 2.93 ;
      RECT 74.96 2.395 75.15 2.96 ;
      RECT 74.375 2.36 74.665 2.59 ;
      RECT 74.375 2.395 75.15 2.565 ;
      RECT 74.435 0.88 74.605 2.59 ;
      RECT 74.375 0.88 74.665 1.11 ;
      RECT 74.375 7.77 74.665 8 ;
      RECT 74.435 6.29 74.605 8 ;
      RECT 74.375 6.29 74.665 6.52 ;
      RECT 74.375 6.325 75.23 6.485 ;
      RECT 75.06 5.92 75.23 6.485 ;
      RECT 74.375 6.32 74.77 6.485 ;
      RECT 74.995 5.92 75.285 6.15 ;
      RECT 74.995 5.95 75.455 6.12 ;
      RECT 74.005 2.73 74.295 2.96 ;
      RECT 74.005 2.76 74.465 2.93 ;
      RECT 74.07 1.655 74.235 2.96 ;
      RECT 72.585 1.625 72.875 1.855 ;
      RECT 72.585 1.655 74.235 1.825 ;
      RECT 72.645 0.885 72.815 1.855 ;
      RECT 72.585 0.885 72.875 1.115 ;
      RECT 72.585 7.765 72.875 7.995 ;
      RECT 72.645 7.025 72.815 7.995 ;
      RECT 72.645 7.12 74.235 7.29 ;
      RECT 74.065 5.92 74.235 7.29 ;
      RECT 72.585 7.025 72.875 7.255 ;
      RECT 74.005 5.92 74.295 6.15 ;
      RECT 74.005 5.95 74.465 6.12 ;
      RECT 70.62 3.43 70.97 3.78 ;
      RECT 70.71 2.025 70.88 3.78 ;
      RECT 73.015 1.965 73.365 2.315 ;
      RECT 70.71 2.025 72.33 2.2 ;
      RECT 70.71 2.025 73.365 2.195 ;
      RECT 73.04 6.655 73.365 6.98 ;
      RECT 68.415 6.61 68.765 6.96 ;
      RECT 73.015 6.655 73.365 6.885 ;
      RECT 68.255 6.655 68.765 6.885 ;
      RECT 68.085 6.685 73.365 6.855 ;
      RECT 72.24 2.365 72.56 2.685 ;
      RECT 72.21 2.365 72.56 2.595 ;
      RECT 72.04 2.395 72.56 2.565 ;
      RECT 72.24 6.225 72.56 6.545 ;
      RECT 72.21 6.285 72.56 6.515 ;
      RECT 72.04 6.315 72.56 6.485 ;
      RECT 68.02 3.665 68.06 3.925 ;
      RECT 68.06 3.645 68.065 3.655 ;
      RECT 69.39 2.89 69.4 3.111 ;
      RECT 69.32 2.885 69.39 3.236 ;
      RECT 69.31 2.885 69.32 3.363 ;
      RECT 69.285 2.885 69.31 3.41 ;
      RECT 69.26 2.885 69.285 3.488 ;
      RECT 69.24 2.885 69.26 3.558 ;
      RECT 69.215 2.885 69.24 3.598 ;
      RECT 69.205 2.885 69.215 3.618 ;
      RECT 69.195 2.887 69.205 3.626 ;
      RECT 69.19 2.892 69.195 3.083 ;
      RECT 69.19 3.092 69.195 3.627 ;
      RECT 69.185 3.137 69.19 3.628 ;
      RECT 69.175 3.202 69.185 3.629 ;
      RECT 69.165 3.297 69.175 3.631 ;
      RECT 69.16 3.35 69.165 3.633 ;
      RECT 69.155 3.37 69.16 3.634 ;
      RECT 69.1 3.395 69.155 3.64 ;
      RECT 69.06 3.43 69.1 3.649 ;
      RECT 69.05 3.447 69.06 3.654 ;
      RECT 69.041 3.453 69.05 3.656 ;
      RECT 68.955 3.491 69.041 3.667 ;
      RECT 68.95 3.53 68.955 3.677 ;
      RECT 68.875 3.537 68.95 3.687 ;
      RECT 68.855 3.547 68.875 3.698 ;
      RECT 68.825 3.554 68.855 3.706 ;
      RECT 68.8 3.561 68.825 3.713 ;
      RECT 68.776 3.567 68.8 3.718 ;
      RECT 68.69 3.58 68.776 3.73 ;
      RECT 68.612 3.587 68.69 3.748 ;
      RECT 68.526 3.582 68.612 3.766 ;
      RECT 68.44 3.577 68.526 3.786 ;
      RECT 68.36 3.571 68.44 3.803 ;
      RECT 68.295 3.567 68.36 3.832 ;
      RECT 68.29 3.281 68.295 3.305 ;
      RECT 68.28 3.557 68.295 3.86 ;
      RECT 68.285 3.275 68.29 3.345 ;
      RECT 68.28 3.269 68.285 3.415 ;
      RECT 68.275 3.263 68.28 3.493 ;
      RECT 68.275 3.54 68.28 3.925 ;
      RECT 68.267 3.26 68.275 3.925 ;
      RECT 68.181 3.258 68.267 3.925 ;
      RECT 68.095 3.256 68.181 3.925 ;
      RECT 68.085 3.257 68.095 3.925 ;
      RECT 68.08 3.262 68.085 3.925 ;
      RECT 68.07 3.275 68.08 3.925 ;
      RECT 68.065 3.297 68.07 3.925 ;
      RECT 68.06 3.657 68.065 3.925 ;
      RECT 68.69 3.125 68.695 3.345 ;
      RECT 69.195 2.16 69.23 2.42 ;
      RECT 69.18 2.16 69.195 2.428 ;
      RECT 69.151 2.16 69.18 2.45 ;
      RECT 69.065 2.16 69.151 2.51 ;
      RECT 69.045 2.16 69.065 2.575 ;
      RECT 68.985 2.16 69.045 2.74 ;
      RECT 68.98 2.16 68.985 2.888 ;
      RECT 68.975 2.16 68.98 2.9 ;
      RECT 68.97 2.16 68.975 2.926 ;
      RECT 68.94 2.346 68.97 3.006 ;
      RECT 68.935 2.394 68.94 3.095 ;
      RECT 68.93 2.408 68.935 3.11 ;
      RECT 68.925 2.427 68.93 3.14 ;
      RECT 68.92 2.442 68.925 3.156 ;
      RECT 68.915 2.457 68.92 3.178 ;
      RECT 68.91 2.477 68.915 3.2 ;
      RECT 68.9 2.497 68.91 3.233 ;
      RECT 68.885 2.539 68.9 3.295 ;
      RECT 68.88 2.57 68.885 3.335 ;
      RECT 68.875 2.582 68.88 3.34 ;
      RECT 68.87 2.594 68.875 3.345 ;
      RECT 68.865 2.607 68.87 3.345 ;
      RECT 68.86 2.625 68.865 3.345 ;
      RECT 68.855 2.645 68.86 3.345 ;
      RECT 68.85 2.657 68.855 3.345 ;
      RECT 68.845 2.67 68.85 3.345 ;
      RECT 68.825 2.705 68.845 3.345 ;
      RECT 68.775 2.807 68.825 3.345 ;
      RECT 68.77 2.892 68.775 3.345 ;
      RECT 68.765 2.9 68.77 3.345 ;
      RECT 68.76 2.917 68.765 3.345 ;
      RECT 68.755 2.932 68.76 3.345 ;
      RECT 68.72 2.997 68.755 3.345 ;
      RECT 68.705 3.062 68.72 3.345 ;
      RECT 68.7 3.092 68.705 3.345 ;
      RECT 68.695 3.117 68.7 3.345 ;
      RECT 68.68 3.127 68.69 3.345 ;
      RECT 68.665 3.14 68.68 3.338 ;
      RECT 68.41 2.73 68.48 2.94 ;
      RECT 68.2 2.707 68.205 2.9 ;
      RECT 65.655 2.635 65.915 2.895 ;
      RECT 68.49 2.917 68.495 2.92 ;
      RECT 68.48 2.735 68.49 2.935 ;
      RECT 68.381 2.728 68.41 2.94 ;
      RECT 68.295 2.72 68.381 2.94 ;
      RECT 68.28 2.714 68.295 2.938 ;
      RECT 68.26 2.713 68.28 2.925 ;
      RECT 68.255 2.712 68.26 2.908 ;
      RECT 68.205 2.709 68.255 2.903 ;
      RECT 68.175 2.706 68.2 2.898 ;
      RECT 68.155 2.704 68.175 2.893 ;
      RECT 68.14 2.702 68.155 2.89 ;
      RECT 68.11 2.7 68.14 2.888 ;
      RECT 68.045 2.696 68.11 2.88 ;
      RECT 68.015 2.691 68.045 2.875 ;
      RECT 67.995 2.689 68.015 2.873 ;
      RECT 67.965 2.686 67.995 2.868 ;
      RECT 67.905 2.682 67.965 2.86 ;
      RECT 67.9 2.679 67.905 2.855 ;
      RECT 67.83 2.677 67.9 2.85 ;
      RECT 67.801 2.673 67.83 2.843 ;
      RECT 67.715 2.668 67.801 2.835 ;
      RECT 67.681 2.663 67.715 2.827 ;
      RECT 67.595 2.655 67.681 2.819 ;
      RECT 67.556 2.648 67.595 2.811 ;
      RECT 67.47 2.643 67.556 2.803 ;
      RECT 67.405 2.637 67.47 2.793 ;
      RECT 67.385 2.632 67.405 2.788 ;
      RECT 67.376 2.629 67.385 2.787 ;
      RECT 67.29 2.625 67.376 2.781 ;
      RECT 67.25 2.621 67.29 2.773 ;
      RECT 67.23 2.617 67.25 2.771 ;
      RECT 67.17 2.617 67.23 2.768 ;
      RECT 67.15 2.62 67.17 2.766 ;
      RECT 67.129 2.62 67.15 2.766 ;
      RECT 67.043 2.622 67.129 2.77 ;
      RECT 66.957 2.624 67.043 2.776 ;
      RECT 66.871 2.626 66.957 2.783 ;
      RECT 66.785 2.629 66.871 2.789 ;
      RECT 66.751 2.63 66.785 2.794 ;
      RECT 66.665 2.633 66.751 2.799 ;
      RECT 66.636 2.64 66.665 2.804 ;
      RECT 66.55 2.64 66.636 2.809 ;
      RECT 66.517 2.64 66.55 2.814 ;
      RECT 66.431 2.642 66.517 2.819 ;
      RECT 66.345 2.644 66.431 2.826 ;
      RECT 66.281 2.646 66.345 2.832 ;
      RECT 66.195 2.648 66.281 2.838 ;
      RECT 66.192 2.65 66.195 2.841 ;
      RECT 66.106 2.651 66.192 2.845 ;
      RECT 66.02 2.654 66.106 2.852 ;
      RECT 66.001 2.656 66.02 2.856 ;
      RECT 65.915 2.658 66.001 2.861 ;
      RECT 65.645 2.67 65.655 2.865 ;
      RECT 67.825 7.765 68.115 7.995 ;
      RECT 67.885 7.025 68.055 7.995 ;
      RECT 67.775 7.055 68.15 7.425 ;
      RECT 67.825 7.025 68.115 7.425 ;
      RECT 67.88 2.25 68.065 2.46 ;
      RECT 67.875 2.251 68.07 2.458 ;
      RECT 67.87 2.256 68.08 2.453 ;
      RECT 67.865 2.232 67.87 2.45 ;
      RECT 67.835 2.229 67.865 2.443 ;
      RECT 67.83 2.225 67.835 2.434 ;
      RECT 67.795 2.256 68.08 2.429 ;
      RECT 67.57 2.165 67.83 2.425 ;
      RECT 67.87 2.234 67.875 2.453 ;
      RECT 67.875 2.235 67.88 2.458 ;
      RECT 67.57 2.247 67.95 2.425 ;
      RECT 67.57 2.245 67.935 2.425 ;
      RECT 67.57 2.24 67.925 2.425 ;
      RECT 67.525 3.155 67.575 3.44 ;
      RECT 67.47 3.125 67.475 3.44 ;
      RECT 67.44 3.105 67.445 3.44 ;
      RECT 67.59 3.155 67.65 3.415 ;
      RECT 67.585 3.155 67.59 3.423 ;
      RECT 67.575 3.155 67.585 3.435 ;
      RECT 67.49 3.145 67.525 3.44 ;
      RECT 67.485 3.132 67.49 3.44 ;
      RECT 67.475 3.127 67.485 3.44 ;
      RECT 67.455 3.117 67.47 3.44 ;
      RECT 67.445 3.11 67.455 3.44 ;
      RECT 67.435 3.102 67.44 3.44 ;
      RECT 67.405 3.092 67.435 3.44 ;
      RECT 67.39 3.08 67.405 3.44 ;
      RECT 67.375 3.07 67.39 3.435 ;
      RECT 67.355 3.06 67.375 3.41 ;
      RECT 67.345 3.052 67.355 3.387 ;
      RECT 67.315 3.035 67.345 3.377 ;
      RECT 67.31 3.012 67.315 3.368 ;
      RECT 67.305 2.999 67.31 3.366 ;
      RECT 67.29 2.975 67.305 3.36 ;
      RECT 67.285 2.951 67.29 3.354 ;
      RECT 67.275 2.94 67.285 3.349 ;
      RECT 67.27 2.93 67.275 3.345 ;
      RECT 67.265 2.922 67.27 3.342 ;
      RECT 67.255 2.917 67.265 3.338 ;
      RECT 67.25 2.912 67.255 3.334 ;
      RECT 67.165 2.91 67.25 3.309 ;
      RECT 67.135 2.91 67.165 3.275 ;
      RECT 67.12 2.91 67.135 3.258 ;
      RECT 67.065 2.91 67.12 3.203 ;
      RECT 67.06 2.915 67.065 3.152 ;
      RECT 67.05 2.92 67.06 3.142 ;
      RECT 67.045 2.93 67.05 3.128 ;
      RECT 66.995 3.67 67.255 3.93 ;
      RECT 66.915 3.685 67.255 3.906 ;
      RECT 66.895 3.685 67.255 3.901 ;
      RECT 66.871 3.685 67.255 3.899 ;
      RECT 66.785 3.685 67.255 3.894 ;
      RECT 66.635 3.625 66.895 3.89 ;
      RECT 66.59 3.685 67.255 3.885 ;
      RECT 66.585 3.692 67.255 3.88 ;
      RECT 66.6 3.68 66.915 3.89 ;
      RECT 66.49 2.115 66.75 2.375 ;
      RECT 66.49 2.172 66.755 2.368 ;
      RECT 66.49 2.202 66.76 2.3 ;
      RECT 66.55 2.633 66.665 2.635 ;
      RECT 66.636 2.63 66.665 2.635 ;
      RECT 65.66 3.634 65.685 3.874 ;
      RECT 65.645 3.637 65.735 3.868 ;
      RECT 65.64 3.642 65.821 3.863 ;
      RECT 65.635 3.65 65.885 3.861 ;
      RECT 65.635 3.65 65.895 3.86 ;
      RECT 65.63 3.657 65.905 3.853 ;
      RECT 65.63 3.657 65.991 3.842 ;
      RECT 65.625 3.692 65.991 3.838 ;
      RECT 65.625 3.692 66 3.827 ;
      RECT 65.905 3.565 66.165 3.825 ;
      RECT 65.615 3.742 66.165 3.823 ;
      RECT 65.885 3.61 65.905 3.858 ;
      RECT 65.821 3.613 65.885 3.862 ;
      RECT 65.735 3.618 65.821 3.867 ;
      RECT 65.665 3.629 66.165 3.825 ;
      RECT 65.685 3.623 65.735 3.872 ;
      RECT 65.81 2.1 65.82 2.362 ;
      RECT 65.8 2.157 65.81 2.365 ;
      RECT 65.775 2.162 65.8 2.371 ;
      RECT 65.75 2.166 65.775 2.383 ;
      RECT 65.74 2.169 65.75 2.393 ;
      RECT 65.735 2.17 65.74 2.398 ;
      RECT 65.73 2.171 65.735 2.403 ;
      RECT 65.725 2.172 65.73 2.405 ;
      RECT 65.7 2.175 65.725 2.408 ;
      RECT 65.67 2.181 65.7 2.411 ;
      RECT 65.605 2.192 65.67 2.414 ;
      RECT 65.56 2.2 65.605 2.418 ;
      RECT 65.545 2.2 65.56 2.426 ;
      RECT 65.54 2.201 65.545 2.433 ;
      RECT 65.535 2.203 65.54 2.436 ;
      RECT 65.53 2.207 65.535 2.439 ;
      RECT 65.52 2.215 65.53 2.443 ;
      RECT 65.515 2.228 65.52 2.448 ;
      RECT 65.51 2.236 65.515 2.45 ;
      RECT 65.505 2.242 65.51 2.45 ;
      RECT 65.5 2.246 65.505 2.453 ;
      RECT 65.495 2.248 65.5 2.456 ;
      RECT 65.49 2.251 65.495 2.459 ;
      RECT 65.48 2.256 65.49 2.463 ;
      RECT 65.475 2.262 65.48 2.468 ;
      RECT 65.465 2.268 65.475 2.472 ;
      RECT 65.45 2.275 65.465 2.478 ;
      RECT 65.421 2.289 65.45 2.488 ;
      RECT 65.335 2.324 65.421 2.52 ;
      RECT 65.315 2.357 65.335 2.549 ;
      RECT 65.295 2.37 65.315 2.56 ;
      RECT 65.275 2.382 65.295 2.571 ;
      RECT 65.225 2.404 65.275 2.591 ;
      RECT 65.21 2.422 65.225 2.608 ;
      RECT 65.205 2.428 65.21 2.611 ;
      RECT 65.2 2.432 65.205 2.614 ;
      RECT 65.195 2.436 65.2 2.618 ;
      RECT 65.19 2.438 65.195 2.621 ;
      RECT 65.18 2.445 65.19 2.624 ;
      RECT 65.175 2.45 65.18 2.628 ;
      RECT 65.17 2.452 65.175 2.631 ;
      RECT 65.165 2.456 65.17 2.634 ;
      RECT 65.16 2.458 65.165 2.638 ;
      RECT 65.145 2.463 65.16 2.643 ;
      RECT 65.14 2.468 65.145 2.646 ;
      RECT 65.135 2.476 65.14 2.649 ;
      RECT 65.13 2.478 65.135 2.652 ;
      RECT 65.125 2.48 65.13 2.655 ;
      RECT 65.115 2.482 65.125 2.661 ;
      RECT 65.08 2.496 65.115 2.673 ;
      RECT 65.07 2.511 65.08 2.683 ;
      RECT 64.995 2.54 65.07 2.707 ;
      RECT 64.99 2.565 64.995 2.73 ;
      RECT 64.975 2.569 64.99 2.736 ;
      RECT 64.965 2.577 64.975 2.741 ;
      RECT 64.935 2.59 64.965 2.745 ;
      RECT 64.925 2.605 64.935 2.75 ;
      RECT 64.915 2.61 64.925 2.753 ;
      RECT 64.91 2.612 64.915 2.755 ;
      RECT 64.895 2.615 64.91 2.758 ;
      RECT 64.89 2.617 64.895 2.761 ;
      RECT 64.87 2.622 64.89 2.765 ;
      RECT 64.84 2.627 64.87 2.773 ;
      RECT 64.815 2.634 64.84 2.781 ;
      RECT 64.81 2.639 64.815 2.786 ;
      RECT 64.78 2.642 64.81 2.79 ;
      RECT 64.74 2.645 64.78 2.8 ;
      RECT 64.705 2.642 64.74 2.812 ;
      RECT 64.695 2.638 64.705 2.819 ;
      RECT 64.67 2.634 64.695 2.825 ;
      RECT 64.665 2.63 64.67 2.83 ;
      RECT 64.625 2.627 64.665 2.83 ;
      RECT 64.61 2.612 64.625 2.831 ;
      RECT 64.587 2.6 64.61 2.831 ;
      RECT 64.501 2.6 64.587 2.832 ;
      RECT 64.415 2.6 64.501 2.834 ;
      RECT 64.395 2.6 64.415 2.831 ;
      RECT 64.39 2.605 64.395 2.826 ;
      RECT 64.385 2.61 64.39 2.824 ;
      RECT 64.375 2.62 64.385 2.822 ;
      RECT 64.37 2.626 64.375 2.815 ;
      RECT 64.365 2.628 64.37 2.8 ;
      RECT 64.36 2.632 64.365 2.79 ;
      RECT 65.82 2.1 66.07 2.36 ;
      RECT 63.545 3.635 63.805 3.895 ;
      RECT 65.84 3.125 65.845 3.335 ;
      RECT 65.845 3.13 65.855 3.33 ;
      RECT 65.795 3.125 65.84 3.35 ;
      RECT 65.785 3.125 65.795 3.37 ;
      RECT 65.766 3.125 65.785 3.375 ;
      RECT 65.68 3.125 65.766 3.372 ;
      RECT 65.65 3.127 65.68 3.37 ;
      RECT 65.595 3.137 65.65 3.368 ;
      RECT 65.53 3.151 65.595 3.366 ;
      RECT 65.525 3.159 65.53 3.365 ;
      RECT 65.51 3.162 65.525 3.363 ;
      RECT 65.445 3.172 65.51 3.359 ;
      RECT 65.397 3.186 65.445 3.36 ;
      RECT 65.311 3.203 65.397 3.374 ;
      RECT 65.225 3.224 65.311 3.391 ;
      RECT 65.205 3.237 65.225 3.401 ;
      RECT 65.16 3.245 65.205 3.408 ;
      RECT 65.125 3.253 65.16 3.416 ;
      RECT 65.091 3.261 65.125 3.424 ;
      RECT 65.005 3.275 65.091 3.436 ;
      RECT 64.97 3.292 65.005 3.448 ;
      RECT 64.961 3.301 64.97 3.452 ;
      RECT 64.875 3.319 64.961 3.469 ;
      RECT 64.816 3.346 64.875 3.496 ;
      RECT 64.73 3.373 64.816 3.524 ;
      RECT 64.71 3.395 64.73 3.544 ;
      RECT 64.65 3.41 64.71 3.56 ;
      RECT 64.64 3.422 64.65 3.573 ;
      RECT 64.635 3.427 64.64 3.576 ;
      RECT 64.625 3.43 64.635 3.579 ;
      RECT 64.62 3.432 64.625 3.582 ;
      RECT 64.59 3.44 64.62 3.589 ;
      RECT 64.575 3.447 64.59 3.597 ;
      RECT 64.565 3.452 64.575 3.601 ;
      RECT 64.56 3.455 64.565 3.604 ;
      RECT 64.55 3.457 64.56 3.607 ;
      RECT 64.515 3.467 64.55 3.616 ;
      RECT 64.44 3.49 64.515 3.638 ;
      RECT 64.42 3.508 64.44 3.656 ;
      RECT 64.39 3.515 64.42 3.666 ;
      RECT 64.37 3.523 64.39 3.676 ;
      RECT 64.36 3.529 64.37 3.683 ;
      RECT 64.341 3.534 64.36 3.689 ;
      RECT 64.255 3.554 64.341 3.709 ;
      RECT 64.24 3.574 64.255 3.728 ;
      RECT 64.195 3.586 64.24 3.739 ;
      RECT 64.13 3.607 64.195 3.762 ;
      RECT 64.09 3.627 64.13 3.783 ;
      RECT 64.08 3.637 64.09 3.793 ;
      RECT 64.03 3.649 64.08 3.804 ;
      RECT 64.01 3.665 64.03 3.816 ;
      RECT 63.98 3.675 64.01 3.822 ;
      RECT 63.97 3.68 63.98 3.824 ;
      RECT 63.901 3.681 63.97 3.83 ;
      RECT 63.815 3.683 63.901 3.84 ;
      RECT 63.805 3.684 63.815 3.845 ;
      RECT 65.075 3.71 65.265 3.92 ;
      RECT 65.065 3.715 65.275 3.913 ;
      RECT 65.05 3.715 65.275 3.878 ;
      RECT 64.97 3.6 65.23 3.86 ;
      RECT 63.885 3.13 64.07 3.425 ;
      RECT 63.875 3.13 64.07 3.423 ;
      RECT 63.86 3.13 64.075 3.418 ;
      RECT 63.86 3.13 64.08 3.415 ;
      RECT 63.855 3.13 64.08 3.413 ;
      RECT 63.85 3.385 64.08 3.403 ;
      RECT 63.855 3.13 64.115 3.39 ;
      RECT 63.815 2.165 64.075 2.425 ;
      RECT 63.625 2.09 63.711 2.423 ;
      RECT 63.6 2.094 63.755 2.419 ;
      RECT 63.711 2.086 63.755 2.419 ;
      RECT 63.711 2.087 63.76 2.418 ;
      RECT 63.625 2.092 63.775 2.417 ;
      RECT 63.6 2.1 63.815 2.416 ;
      RECT 63.595 2.095 63.775 2.411 ;
      RECT 63.585 2.11 63.815 2.318 ;
      RECT 63.585 2.162 64.015 2.318 ;
      RECT 63.585 2.155 63.995 2.318 ;
      RECT 63.585 2.142 63.965 2.318 ;
      RECT 63.585 2.13 63.905 2.318 ;
      RECT 63.585 2.115 63.88 2.318 ;
      RECT 62.785 2.745 62.92 3.04 ;
      RECT 63.045 2.768 63.05 2.955 ;
      RECT 63.765 2.665 63.91 2.9 ;
      RECT 63.925 2.665 63.93 2.89 ;
      RECT 63.96 2.676 63.965 2.87 ;
      RECT 63.955 2.668 63.96 2.875 ;
      RECT 63.935 2.665 63.955 2.88 ;
      RECT 63.93 2.665 63.935 2.888 ;
      RECT 63.92 2.665 63.925 2.893 ;
      RECT 63.91 2.665 63.92 2.898 ;
      RECT 63.74 2.667 63.765 2.9 ;
      RECT 63.69 2.674 63.74 2.9 ;
      RECT 63.685 2.679 63.69 2.9 ;
      RECT 63.646 2.684 63.685 2.901 ;
      RECT 63.56 2.696 63.646 2.902 ;
      RECT 63.551 2.706 63.56 2.902 ;
      RECT 63.465 2.715 63.551 2.904 ;
      RECT 63.441 2.725 63.465 2.906 ;
      RECT 63.355 2.736 63.441 2.907 ;
      RECT 63.325 2.747 63.355 2.909 ;
      RECT 63.295 2.752 63.325 2.911 ;
      RECT 63.27 2.758 63.295 2.914 ;
      RECT 63.255 2.763 63.27 2.915 ;
      RECT 63.21 2.769 63.255 2.915 ;
      RECT 63.205 2.774 63.21 2.916 ;
      RECT 63.185 2.774 63.205 2.918 ;
      RECT 63.165 2.772 63.185 2.923 ;
      RECT 63.13 2.771 63.165 2.93 ;
      RECT 63.1 2.77 63.13 2.94 ;
      RECT 63.05 2.769 63.1 2.95 ;
      RECT 62.96 2.766 63.045 3.04 ;
      RECT 62.935 2.76 62.96 3.04 ;
      RECT 62.92 2.75 62.935 3.04 ;
      RECT 62.735 2.745 62.785 2.96 ;
      RECT 62.725 2.75 62.735 2.95 ;
      RECT 62.965 3.225 63.225 3.485 ;
      RECT 62.965 3.225 63.255 3.378 ;
      RECT 62.965 3.225 63.29 3.363 ;
      RECT 63.22 3.145 63.41 3.355 ;
      RECT 63.21 3.15 63.42 3.348 ;
      RECT 63.175 3.22 63.42 3.348 ;
      RECT 63.205 3.162 63.225 3.485 ;
      RECT 63.19 3.21 63.42 3.348 ;
      RECT 63.195 3.182 63.225 3.485 ;
      RECT 62.275 2.25 62.345 3.355 ;
      RECT 63.01 2.355 63.27 2.615 ;
      RECT 62.59 2.401 62.605 2.61 ;
      RECT 62.926 2.414 63.01 2.565 ;
      RECT 62.84 2.411 62.926 2.565 ;
      RECT 62.801 2.409 62.84 2.565 ;
      RECT 62.715 2.407 62.801 2.565 ;
      RECT 62.655 2.405 62.715 2.576 ;
      RECT 62.62 2.403 62.655 2.594 ;
      RECT 62.605 2.401 62.62 2.605 ;
      RECT 62.575 2.401 62.59 2.618 ;
      RECT 62.565 2.401 62.575 2.623 ;
      RECT 62.54 2.4 62.565 2.628 ;
      RECT 62.525 2.395 62.54 2.634 ;
      RECT 62.52 2.388 62.525 2.639 ;
      RECT 62.495 2.379 62.52 2.645 ;
      RECT 62.45 2.358 62.495 2.658 ;
      RECT 62.44 2.342 62.45 2.668 ;
      RECT 62.425 2.335 62.44 2.678 ;
      RECT 62.415 2.328 62.425 2.695 ;
      RECT 62.41 2.325 62.415 2.725 ;
      RECT 62.405 2.323 62.41 2.755 ;
      RECT 62.4 2.321 62.405 2.792 ;
      RECT 62.385 2.317 62.4 2.859 ;
      RECT 62.385 3.15 62.395 3.35 ;
      RECT 62.38 2.313 62.385 2.985 ;
      RECT 62.38 3.137 62.385 3.355 ;
      RECT 62.375 2.311 62.38 3.07 ;
      RECT 62.375 3.127 62.38 3.355 ;
      RECT 62.36 2.282 62.375 3.355 ;
      RECT 62.345 2.255 62.36 3.355 ;
      RECT 62.27 2.25 62.275 2.605 ;
      RECT 62.27 2.66 62.275 3.355 ;
      RECT 62.255 2.25 62.27 2.583 ;
      RECT 62.265 2.682 62.27 3.355 ;
      RECT 62.255 2.722 62.265 3.355 ;
      RECT 62.22 2.25 62.255 2.525 ;
      RECT 62.25 2.757 62.255 3.355 ;
      RECT 62.235 2.812 62.25 3.355 ;
      RECT 62.23 2.877 62.235 3.355 ;
      RECT 62.215 2.925 62.23 3.355 ;
      RECT 62.19 2.25 62.22 2.48 ;
      RECT 62.21 2.98 62.215 3.355 ;
      RECT 62.195 3.04 62.21 3.355 ;
      RECT 62.19 3.088 62.195 3.353 ;
      RECT 62.185 2.25 62.19 2.473 ;
      RECT 62.185 3.12 62.19 3.348 ;
      RECT 62.16 2.25 62.185 2.465 ;
      RECT 62.15 2.255 62.16 2.455 ;
      RECT 62.365 3.53 62.385 3.77 ;
      RECT 61.595 3.46 61.6 3.67 ;
      RECT 62.875 3.533 62.885 3.728 ;
      RECT 62.87 3.523 62.875 3.731 ;
      RECT 62.79 3.52 62.87 3.754 ;
      RECT 62.786 3.52 62.79 3.776 ;
      RECT 62.7 3.52 62.786 3.786 ;
      RECT 62.685 3.52 62.7 3.794 ;
      RECT 62.656 3.521 62.685 3.792 ;
      RECT 62.57 3.526 62.656 3.788 ;
      RECT 62.557 3.53 62.57 3.784 ;
      RECT 62.471 3.53 62.557 3.78 ;
      RECT 62.385 3.53 62.471 3.774 ;
      RECT 62.301 3.53 62.365 3.768 ;
      RECT 62.215 3.53 62.301 3.763 ;
      RECT 62.195 3.53 62.215 3.759 ;
      RECT 62.135 3.525 62.195 3.756 ;
      RECT 62.107 3.519 62.135 3.753 ;
      RECT 62.021 3.514 62.107 3.749 ;
      RECT 61.935 3.508 62.021 3.743 ;
      RECT 61.86 3.49 61.935 3.738 ;
      RECT 61.825 3.467 61.86 3.734 ;
      RECT 61.815 3.457 61.825 3.733 ;
      RECT 61.76 3.455 61.815 3.732 ;
      RECT 61.685 3.455 61.76 3.728 ;
      RECT 61.675 3.455 61.685 3.723 ;
      RECT 61.66 3.455 61.675 3.715 ;
      RECT 61.61 3.457 61.66 3.693 ;
      RECT 61.6 3.46 61.61 3.673 ;
      RECT 61.59 3.465 61.595 3.668 ;
      RECT 61.585 3.47 61.59 3.663 ;
      RECT 61.71 2.635 61.97 2.895 ;
      RECT 61.71 2.65 61.99 2.86 ;
      RECT 61.71 2.655 62 2.855 ;
      RECT 59.695 2.115 59.955 2.375 ;
      RECT 59.685 2.145 59.955 2.355 ;
      RECT 61.605 2.06 61.865 2.32 ;
      RECT 61.6 2.135 61.605 2.321 ;
      RECT 61.575 2.14 61.6 2.323 ;
      RECT 61.56 2.147 61.575 2.326 ;
      RECT 61.5 2.165 61.56 2.331 ;
      RECT 61.47 2.185 61.5 2.338 ;
      RECT 61.445 2.193 61.47 2.343 ;
      RECT 61.42 2.201 61.445 2.345 ;
      RECT 61.402 2.205 61.42 2.344 ;
      RECT 61.316 2.203 61.402 2.344 ;
      RECT 61.23 2.201 61.316 2.344 ;
      RECT 61.144 2.199 61.23 2.343 ;
      RECT 61.058 2.197 61.144 2.343 ;
      RECT 60.972 2.195 61.058 2.343 ;
      RECT 60.886 2.193 60.972 2.343 ;
      RECT 60.8 2.191 60.886 2.342 ;
      RECT 60.782 2.19 60.8 2.342 ;
      RECT 60.696 2.189 60.782 2.342 ;
      RECT 60.61 2.187 60.696 2.342 ;
      RECT 60.524 2.186 60.61 2.341 ;
      RECT 60.438 2.185 60.524 2.341 ;
      RECT 60.352 2.183 60.438 2.341 ;
      RECT 60.266 2.182 60.352 2.341 ;
      RECT 60.18 2.18 60.266 2.34 ;
      RECT 60.156 2.178 60.18 2.34 ;
      RECT 60.07 2.171 60.156 2.34 ;
      RECT 60.041 2.163 60.07 2.34 ;
      RECT 59.955 2.155 60.041 2.34 ;
      RECT 59.675 2.152 59.685 2.35 ;
      RECT 61.18 3.115 61.185 3.465 ;
      RECT 60.95 3.205 61.09 3.465 ;
      RECT 61.425 2.89 61.47 3.1 ;
      RECT 61.48 2.901 61.49 3.095 ;
      RECT 61.47 2.893 61.48 3.1 ;
      RECT 61.405 2.89 61.425 3.105 ;
      RECT 61.375 2.89 61.405 3.128 ;
      RECT 61.365 2.89 61.375 3.153 ;
      RECT 61.36 2.89 61.365 3.163 ;
      RECT 61.305 2.89 61.36 3.203 ;
      RECT 61.3 2.89 61.305 3.243 ;
      RECT 61.295 2.892 61.3 3.248 ;
      RECT 61.28 2.902 61.295 3.259 ;
      RECT 61.235 2.96 61.28 3.295 ;
      RECT 61.225 3.015 61.235 3.329 ;
      RECT 61.21 3.042 61.225 3.345 ;
      RECT 61.2 3.069 61.21 3.465 ;
      RECT 61.185 3.092 61.2 3.465 ;
      RECT 61.175 3.132 61.18 3.465 ;
      RECT 61.17 3.142 61.175 3.465 ;
      RECT 61.165 3.157 61.17 3.465 ;
      RECT 61.155 3.162 61.165 3.465 ;
      RECT 61.09 3.185 61.155 3.465 ;
      RECT 60.59 2.68 60.78 2.89 ;
      RECT 59.165 2.605 59.425 2.865 ;
      RECT 59.515 2.6 59.61 2.81 ;
      RECT 59.49 2.615 59.5 2.81 ;
      RECT 60.78 2.687 60.79 2.885 ;
      RECT 60.58 2.687 60.59 2.885 ;
      RECT 60.565 2.702 60.58 2.875 ;
      RECT 60.56 2.71 60.565 2.868 ;
      RECT 60.55 2.713 60.56 2.865 ;
      RECT 60.515 2.712 60.55 2.863 ;
      RECT 60.486 2.708 60.515 2.86 ;
      RECT 60.4 2.703 60.486 2.857 ;
      RECT 60.34 2.697 60.4 2.853 ;
      RECT 60.311 2.693 60.34 2.85 ;
      RECT 60.225 2.685 60.311 2.847 ;
      RECT 60.216 2.679 60.225 2.845 ;
      RECT 60.13 2.674 60.216 2.843 ;
      RECT 60.107 2.669 60.13 2.84 ;
      RECT 60.021 2.663 60.107 2.837 ;
      RECT 59.935 2.654 60.021 2.832 ;
      RECT 59.925 2.649 59.935 2.83 ;
      RECT 59.906 2.648 59.925 2.829 ;
      RECT 59.82 2.643 59.906 2.825 ;
      RECT 59.8 2.638 59.82 2.821 ;
      RECT 59.74 2.633 59.8 2.818 ;
      RECT 59.715 2.623 59.74 2.816 ;
      RECT 59.71 2.616 59.715 2.815 ;
      RECT 59.7 2.607 59.71 2.814 ;
      RECT 59.696 2.6 59.7 2.814 ;
      RECT 59.61 2.6 59.696 2.812 ;
      RECT 59.5 2.607 59.515 2.81 ;
      RECT 59.485 2.617 59.49 2.81 ;
      RECT 59.465 2.62 59.485 2.807 ;
      RECT 59.435 2.62 59.465 2.803 ;
      RECT 59.425 2.62 59.435 2.803 ;
      RECT 60.34 3.115 60.6 3.375 ;
      RECT 60.27 3.125 60.6 3.335 ;
      RECT 60.26 3.132 60.6 3.33 ;
      RECT 59.68 3.12 59.94 3.38 ;
      RECT 59.68 3.16 60.045 3.37 ;
      RECT 59.68 3.162 60.05 3.369 ;
      RECT 59.68 3.17 60.055 3.366 ;
      RECT 58.605 2.245 58.705 3.77 ;
      RECT 58.795 3.385 58.845 3.645 ;
      RECT 58.79 2.258 58.795 2.445 ;
      RECT 58.785 3.366 58.795 3.645 ;
      RECT 58.785 2.255 58.79 2.453 ;
      RECT 58.77 2.249 58.785 2.46 ;
      RECT 58.78 3.354 58.785 3.728 ;
      RECT 58.77 3.342 58.78 3.765 ;
      RECT 58.76 2.245 58.77 2.467 ;
      RECT 58.76 3.327 58.77 3.77 ;
      RECT 58.755 2.245 58.76 2.475 ;
      RECT 58.735 3.297 58.76 3.77 ;
      RECT 58.715 2.245 58.755 2.523 ;
      RECT 58.725 3.257 58.735 3.77 ;
      RECT 58.715 3.212 58.725 3.77 ;
      RECT 58.71 2.245 58.715 2.593 ;
      RECT 58.71 3.17 58.715 3.77 ;
      RECT 58.705 2.245 58.71 3.07 ;
      RECT 58.705 3.152 58.71 3.77 ;
      RECT 58.595 2.248 58.605 3.77 ;
      RECT 58.58 2.255 58.595 3.766 ;
      RECT 58.575 2.265 58.58 3.761 ;
      RECT 58.57 2.465 58.575 3.653 ;
      RECT 58.565 2.55 58.57 3.205 ;
      RECT 57.44 7.77 57.73 8 ;
      RECT 57.5 6.29 57.67 8 ;
      RECT 57.45 6.655 57.8 7.005 ;
      RECT 57.44 6.29 57.73 6.52 ;
      RECT 57.035 2.395 57.14 2.965 ;
      RECT 57.035 2.73 57.36 2.96 ;
      RECT 57.035 2.76 57.53 2.93 ;
      RECT 57.035 2.395 57.225 2.96 ;
      RECT 56.45 2.36 56.74 2.59 ;
      RECT 56.45 2.395 57.225 2.565 ;
      RECT 56.51 0.88 56.68 2.59 ;
      RECT 56.45 0.88 56.74 1.11 ;
      RECT 56.45 7.77 56.74 8 ;
      RECT 56.51 6.29 56.68 8 ;
      RECT 56.45 6.29 56.74 6.52 ;
      RECT 56.45 6.325 57.305 6.485 ;
      RECT 57.135 5.92 57.305 6.485 ;
      RECT 56.45 6.32 56.845 6.485 ;
      RECT 57.07 5.92 57.36 6.15 ;
      RECT 57.07 5.95 57.53 6.12 ;
      RECT 56.08 2.73 56.37 2.96 ;
      RECT 56.08 2.76 56.54 2.93 ;
      RECT 56.145 1.655 56.31 2.96 ;
      RECT 54.66 1.625 54.95 1.855 ;
      RECT 54.66 1.655 56.31 1.825 ;
      RECT 54.72 0.885 54.89 1.855 ;
      RECT 54.66 0.885 54.95 1.115 ;
      RECT 54.66 7.765 54.95 7.995 ;
      RECT 54.72 7.025 54.89 7.995 ;
      RECT 54.72 7.12 56.31 7.29 ;
      RECT 56.14 5.92 56.31 7.29 ;
      RECT 54.66 7.025 54.95 7.255 ;
      RECT 56.08 5.92 56.37 6.15 ;
      RECT 56.08 5.95 56.54 6.12 ;
      RECT 52.695 3.43 53.045 3.78 ;
      RECT 52.785 2.025 52.955 3.78 ;
      RECT 55.09 1.965 55.44 2.315 ;
      RECT 52.785 2.025 54.405 2.2 ;
      RECT 52.785 2.025 55.44 2.195 ;
      RECT 55.115 6.655 55.44 6.98 ;
      RECT 50.545 6.615 50.895 6.965 ;
      RECT 55.09 6.655 55.44 6.885 ;
      RECT 50.33 6.655 50.895 6.885 ;
      RECT 50.16 6.685 55.44 6.855 ;
      RECT 54.315 2.365 54.635 2.685 ;
      RECT 54.285 2.365 54.635 2.595 ;
      RECT 54.115 2.395 54.635 2.565 ;
      RECT 54.315 6.225 54.635 6.545 ;
      RECT 54.285 6.285 54.635 6.515 ;
      RECT 54.115 6.315 54.635 6.485 ;
      RECT 50.095 3.665 50.135 3.925 ;
      RECT 50.135 3.645 50.14 3.655 ;
      RECT 51.465 2.89 51.475 3.111 ;
      RECT 51.395 2.885 51.465 3.236 ;
      RECT 51.385 2.885 51.395 3.363 ;
      RECT 51.36 2.885 51.385 3.41 ;
      RECT 51.335 2.885 51.36 3.488 ;
      RECT 51.315 2.885 51.335 3.558 ;
      RECT 51.29 2.885 51.315 3.598 ;
      RECT 51.28 2.885 51.29 3.618 ;
      RECT 51.27 2.887 51.28 3.626 ;
      RECT 51.265 2.892 51.27 3.083 ;
      RECT 51.265 3.092 51.27 3.627 ;
      RECT 51.26 3.137 51.265 3.628 ;
      RECT 51.25 3.202 51.26 3.629 ;
      RECT 51.24 3.297 51.25 3.631 ;
      RECT 51.235 3.35 51.24 3.633 ;
      RECT 51.23 3.37 51.235 3.634 ;
      RECT 51.175 3.395 51.23 3.64 ;
      RECT 51.135 3.43 51.175 3.649 ;
      RECT 51.125 3.447 51.135 3.654 ;
      RECT 51.116 3.453 51.125 3.656 ;
      RECT 51.03 3.491 51.116 3.667 ;
      RECT 51.025 3.53 51.03 3.677 ;
      RECT 50.95 3.537 51.025 3.687 ;
      RECT 50.93 3.547 50.95 3.698 ;
      RECT 50.9 3.554 50.93 3.706 ;
      RECT 50.875 3.561 50.9 3.713 ;
      RECT 50.851 3.567 50.875 3.718 ;
      RECT 50.765 3.58 50.851 3.73 ;
      RECT 50.687 3.587 50.765 3.748 ;
      RECT 50.601 3.582 50.687 3.766 ;
      RECT 50.515 3.577 50.601 3.786 ;
      RECT 50.435 3.571 50.515 3.803 ;
      RECT 50.37 3.567 50.435 3.832 ;
      RECT 50.365 3.281 50.37 3.305 ;
      RECT 50.355 3.557 50.37 3.86 ;
      RECT 50.36 3.275 50.365 3.345 ;
      RECT 50.355 3.269 50.36 3.415 ;
      RECT 50.35 3.263 50.355 3.493 ;
      RECT 50.35 3.54 50.355 3.925 ;
      RECT 50.342 3.26 50.35 3.925 ;
      RECT 50.256 3.258 50.342 3.925 ;
      RECT 50.17 3.256 50.256 3.925 ;
      RECT 50.16 3.257 50.17 3.925 ;
      RECT 50.155 3.262 50.16 3.925 ;
      RECT 50.145 3.275 50.155 3.925 ;
      RECT 50.14 3.297 50.145 3.925 ;
      RECT 50.135 3.657 50.14 3.925 ;
      RECT 50.765 3.125 50.77 3.345 ;
      RECT 51.27 2.16 51.305 2.42 ;
      RECT 51.255 2.16 51.27 2.428 ;
      RECT 51.226 2.16 51.255 2.45 ;
      RECT 51.14 2.16 51.226 2.51 ;
      RECT 51.12 2.16 51.14 2.575 ;
      RECT 51.06 2.16 51.12 2.74 ;
      RECT 51.055 2.16 51.06 2.888 ;
      RECT 51.05 2.16 51.055 2.9 ;
      RECT 51.045 2.16 51.05 2.926 ;
      RECT 51.015 2.346 51.045 3.006 ;
      RECT 51.01 2.394 51.015 3.095 ;
      RECT 51.005 2.408 51.01 3.11 ;
      RECT 51 2.427 51.005 3.14 ;
      RECT 50.995 2.442 51 3.156 ;
      RECT 50.99 2.457 50.995 3.178 ;
      RECT 50.985 2.477 50.99 3.2 ;
      RECT 50.975 2.497 50.985 3.233 ;
      RECT 50.96 2.539 50.975 3.295 ;
      RECT 50.955 2.57 50.96 3.335 ;
      RECT 50.95 2.582 50.955 3.34 ;
      RECT 50.945 2.594 50.95 3.345 ;
      RECT 50.94 2.607 50.945 3.345 ;
      RECT 50.935 2.625 50.94 3.345 ;
      RECT 50.93 2.645 50.935 3.345 ;
      RECT 50.925 2.657 50.93 3.345 ;
      RECT 50.92 2.67 50.925 3.345 ;
      RECT 50.9 2.705 50.92 3.345 ;
      RECT 50.85 2.807 50.9 3.345 ;
      RECT 50.845 2.892 50.85 3.345 ;
      RECT 50.84 2.9 50.845 3.345 ;
      RECT 50.835 2.917 50.84 3.345 ;
      RECT 50.83 2.932 50.835 3.345 ;
      RECT 50.795 2.997 50.83 3.345 ;
      RECT 50.78 3.062 50.795 3.345 ;
      RECT 50.775 3.092 50.78 3.345 ;
      RECT 50.77 3.117 50.775 3.345 ;
      RECT 50.755 3.127 50.765 3.345 ;
      RECT 50.74 3.14 50.755 3.338 ;
      RECT 50.485 2.73 50.555 2.94 ;
      RECT 50.275 2.707 50.28 2.9 ;
      RECT 47.73 2.635 47.99 2.895 ;
      RECT 50.565 2.917 50.57 2.92 ;
      RECT 50.555 2.735 50.565 2.935 ;
      RECT 50.456 2.728 50.485 2.94 ;
      RECT 50.37 2.72 50.456 2.94 ;
      RECT 50.355 2.714 50.37 2.938 ;
      RECT 50.335 2.713 50.355 2.925 ;
      RECT 50.33 2.712 50.335 2.908 ;
      RECT 50.28 2.709 50.33 2.903 ;
      RECT 50.25 2.706 50.275 2.898 ;
      RECT 50.23 2.704 50.25 2.893 ;
      RECT 50.215 2.702 50.23 2.89 ;
      RECT 50.185 2.7 50.215 2.888 ;
      RECT 50.12 2.696 50.185 2.88 ;
      RECT 50.09 2.691 50.12 2.875 ;
      RECT 50.07 2.689 50.09 2.873 ;
      RECT 50.04 2.686 50.07 2.868 ;
      RECT 49.98 2.682 50.04 2.86 ;
      RECT 49.975 2.679 49.98 2.855 ;
      RECT 49.905 2.677 49.975 2.85 ;
      RECT 49.876 2.673 49.905 2.843 ;
      RECT 49.79 2.668 49.876 2.835 ;
      RECT 49.756 2.663 49.79 2.827 ;
      RECT 49.67 2.655 49.756 2.819 ;
      RECT 49.631 2.648 49.67 2.811 ;
      RECT 49.545 2.643 49.631 2.803 ;
      RECT 49.48 2.637 49.545 2.793 ;
      RECT 49.46 2.632 49.48 2.788 ;
      RECT 49.451 2.629 49.46 2.787 ;
      RECT 49.365 2.625 49.451 2.781 ;
      RECT 49.325 2.621 49.365 2.773 ;
      RECT 49.305 2.617 49.325 2.771 ;
      RECT 49.245 2.617 49.305 2.768 ;
      RECT 49.225 2.62 49.245 2.766 ;
      RECT 49.204 2.62 49.225 2.766 ;
      RECT 49.118 2.622 49.204 2.77 ;
      RECT 49.032 2.624 49.118 2.776 ;
      RECT 48.946 2.626 49.032 2.783 ;
      RECT 48.86 2.629 48.946 2.789 ;
      RECT 48.826 2.63 48.86 2.794 ;
      RECT 48.74 2.633 48.826 2.799 ;
      RECT 48.711 2.64 48.74 2.804 ;
      RECT 48.625 2.64 48.711 2.809 ;
      RECT 48.592 2.64 48.625 2.814 ;
      RECT 48.506 2.642 48.592 2.819 ;
      RECT 48.42 2.644 48.506 2.826 ;
      RECT 48.356 2.646 48.42 2.832 ;
      RECT 48.27 2.648 48.356 2.838 ;
      RECT 48.267 2.65 48.27 2.841 ;
      RECT 48.181 2.651 48.267 2.845 ;
      RECT 48.095 2.654 48.181 2.852 ;
      RECT 48.076 2.656 48.095 2.856 ;
      RECT 47.99 2.658 48.076 2.861 ;
      RECT 47.72 2.67 47.73 2.865 ;
      RECT 49.9 7.765 50.19 7.995 ;
      RECT 49.96 7.025 50.13 7.995 ;
      RECT 49.85 7.055 50.225 7.425 ;
      RECT 49.9 7.025 50.19 7.425 ;
      RECT 49.955 2.25 50.14 2.46 ;
      RECT 49.95 2.251 50.145 2.458 ;
      RECT 49.945 2.256 50.155 2.453 ;
      RECT 49.94 2.232 49.945 2.45 ;
      RECT 49.91 2.229 49.94 2.443 ;
      RECT 49.905 2.225 49.91 2.434 ;
      RECT 49.87 2.256 50.155 2.429 ;
      RECT 49.645 2.165 49.905 2.425 ;
      RECT 49.945 2.234 49.95 2.453 ;
      RECT 49.95 2.235 49.955 2.458 ;
      RECT 49.645 2.247 50.025 2.425 ;
      RECT 49.645 2.245 50.01 2.425 ;
      RECT 49.645 2.24 50 2.425 ;
      RECT 49.6 3.155 49.65 3.44 ;
      RECT 49.545 3.125 49.55 3.44 ;
      RECT 49.515 3.105 49.52 3.44 ;
      RECT 49.665 3.155 49.725 3.415 ;
      RECT 49.66 3.155 49.665 3.423 ;
      RECT 49.65 3.155 49.66 3.435 ;
      RECT 49.565 3.145 49.6 3.44 ;
      RECT 49.56 3.132 49.565 3.44 ;
      RECT 49.55 3.127 49.56 3.44 ;
      RECT 49.53 3.117 49.545 3.44 ;
      RECT 49.52 3.11 49.53 3.44 ;
      RECT 49.51 3.102 49.515 3.44 ;
      RECT 49.48 3.092 49.51 3.44 ;
      RECT 49.465 3.08 49.48 3.44 ;
      RECT 49.45 3.07 49.465 3.435 ;
      RECT 49.43 3.06 49.45 3.41 ;
      RECT 49.42 3.052 49.43 3.387 ;
      RECT 49.39 3.035 49.42 3.377 ;
      RECT 49.385 3.012 49.39 3.368 ;
      RECT 49.38 2.999 49.385 3.366 ;
      RECT 49.365 2.975 49.38 3.36 ;
      RECT 49.36 2.951 49.365 3.354 ;
      RECT 49.35 2.94 49.36 3.349 ;
      RECT 49.345 2.93 49.35 3.345 ;
      RECT 49.34 2.922 49.345 3.342 ;
      RECT 49.33 2.917 49.34 3.338 ;
      RECT 49.325 2.912 49.33 3.334 ;
      RECT 49.24 2.91 49.325 3.309 ;
      RECT 49.21 2.91 49.24 3.275 ;
      RECT 49.195 2.91 49.21 3.258 ;
      RECT 49.14 2.91 49.195 3.203 ;
      RECT 49.135 2.915 49.14 3.152 ;
      RECT 49.125 2.92 49.135 3.142 ;
      RECT 49.12 2.93 49.125 3.128 ;
      RECT 49.07 3.67 49.33 3.93 ;
      RECT 48.99 3.685 49.33 3.906 ;
      RECT 48.97 3.685 49.33 3.901 ;
      RECT 48.946 3.685 49.33 3.899 ;
      RECT 48.86 3.685 49.33 3.894 ;
      RECT 48.71 3.625 48.97 3.89 ;
      RECT 48.665 3.685 49.33 3.885 ;
      RECT 48.66 3.692 49.33 3.88 ;
      RECT 48.675 3.68 48.99 3.89 ;
      RECT 48.565 2.115 48.825 2.375 ;
      RECT 48.565 2.172 48.83 2.368 ;
      RECT 48.565 2.202 48.835 2.3 ;
      RECT 48.625 2.633 48.74 2.635 ;
      RECT 48.711 2.63 48.74 2.635 ;
      RECT 47.735 3.634 47.76 3.874 ;
      RECT 47.72 3.637 47.81 3.868 ;
      RECT 47.715 3.642 47.896 3.863 ;
      RECT 47.71 3.65 47.96 3.861 ;
      RECT 47.71 3.65 47.97 3.86 ;
      RECT 47.705 3.657 47.98 3.853 ;
      RECT 47.705 3.657 48.066 3.842 ;
      RECT 47.7 3.692 48.066 3.838 ;
      RECT 47.7 3.692 48.075 3.827 ;
      RECT 47.98 3.565 48.24 3.825 ;
      RECT 47.69 3.742 48.24 3.823 ;
      RECT 47.96 3.61 47.98 3.858 ;
      RECT 47.896 3.613 47.96 3.862 ;
      RECT 47.81 3.618 47.896 3.867 ;
      RECT 47.74 3.629 48.24 3.825 ;
      RECT 47.76 3.623 47.81 3.872 ;
      RECT 47.885 2.1 47.895 2.362 ;
      RECT 47.875 2.157 47.885 2.365 ;
      RECT 47.85 2.162 47.875 2.371 ;
      RECT 47.825 2.166 47.85 2.383 ;
      RECT 47.815 2.169 47.825 2.393 ;
      RECT 47.81 2.17 47.815 2.398 ;
      RECT 47.805 2.171 47.81 2.403 ;
      RECT 47.8 2.172 47.805 2.405 ;
      RECT 47.775 2.175 47.8 2.408 ;
      RECT 47.745 2.181 47.775 2.411 ;
      RECT 47.68 2.192 47.745 2.414 ;
      RECT 47.635 2.2 47.68 2.418 ;
      RECT 47.62 2.2 47.635 2.426 ;
      RECT 47.615 2.201 47.62 2.433 ;
      RECT 47.61 2.203 47.615 2.436 ;
      RECT 47.605 2.207 47.61 2.439 ;
      RECT 47.595 2.215 47.605 2.443 ;
      RECT 47.59 2.228 47.595 2.448 ;
      RECT 47.585 2.236 47.59 2.45 ;
      RECT 47.58 2.242 47.585 2.45 ;
      RECT 47.575 2.246 47.58 2.453 ;
      RECT 47.57 2.248 47.575 2.456 ;
      RECT 47.565 2.251 47.57 2.459 ;
      RECT 47.555 2.256 47.565 2.463 ;
      RECT 47.55 2.262 47.555 2.468 ;
      RECT 47.54 2.268 47.55 2.472 ;
      RECT 47.525 2.275 47.54 2.478 ;
      RECT 47.496 2.289 47.525 2.488 ;
      RECT 47.41 2.324 47.496 2.52 ;
      RECT 47.39 2.357 47.41 2.549 ;
      RECT 47.37 2.37 47.39 2.56 ;
      RECT 47.35 2.382 47.37 2.571 ;
      RECT 47.3 2.404 47.35 2.591 ;
      RECT 47.285 2.422 47.3 2.608 ;
      RECT 47.28 2.428 47.285 2.611 ;
      RECT 47.275 2.432 47.28 2.614 ;
      RECT 47.27 2.436 47.275 2.618 ;
      RECT 47.265 2.438 47.27 2.621 ;
      RECT 47.255 2.445 47.265 2.624 ;
      RECT 47.25 2.45 47.255 2.628 ;
      RECT 47.245 2.452 47.25 2.631 ;
      RECT 47.24 2.456 47.245 2.634 ;
      RECT 47.235 2.458 47.24 2.638 ;
      RECT 47.22 2.463 47.235 2.643 ;
      RECT 47.215 2.468 47.22 2.646 ;
      RECT 47.21 2.476 47.215 2.649 ;
      RECT 47.205 2.478 47.21 2.652 ;
      RECT 47.2 2.48 47.205 2.655 ;
      RECT 47.19 2.482 47.2 2.661 ;
      RECT 47.155 2.496 47.19 2.673 ;
      RECT 47.145 2.511 47.155 2.683 ;
      RECT 47.07 2.54 47.145 2.707 ;
      RECT 47.065 2.565 47.07 2.73 ;
      RECT 47.05 2.569 47.065 2.736 ;
      RECT 47.04 2.577 47.05 2.741 ;
      RECT 47.01 2.59 47.04 2.745 ;
      RECT 47 2.605 47.01 2.75 ;
      RECT 46.99 2.61 47 2.753 ;
      RECT 46.985 2.612 46.99 2.755 ;
      RECT 46.97 2.615 46.985 2.758 ;
      RECT 46.965 2.617 46.97 2.761 ;
      RECT 46.945 2.622 46.965 2.765 ;
      RECT 46.915 2.627 46.945 2.773 ;
      RECT 46.89 2.634 46.915 2.781 ;
      RECT 46.885 2.639 46.89 2.786 ;
      RECT 46.855 2.642 46.885 2.79 ;
      RECT 46.815 2.645 46.855 2.8 ;
      RECT 46.78 2.642 46.815 2.812 ;
      RECT 46.77 2.638 46.78 2.819 ;
      RECT 46.745 2.634 46.77 2.825 ;
      RECT 46.74 2.63 46.745 2.83 ;
      RECT 46.7 2.627 46.74 2.83 ;
      RECT 46.685 2.612 46.7 2.831 ;
      RECT 46.662 2.6 46.685 2.831 ;
      RECT 46.576 2.6 46.662 2.832 ;
      RECT 46.49 2.6 46.576 2.834 ;
      RECT 46.47 2.6 46.49 2.831 ;
      RECT 46.465 2.605 46.47 2.826 ;
      RECT 46.46 2.61 46.465 2.824 ;
      RECT 46.45 2.62 46.46 2.822 ;
      RECT 46.445 2.626 46.45 2.815 ;
      RECT 46.44 2.628 46.445 2.8 ;
      RECT 46.435 2.632 46.44 2.79 ;
      RECT 47.895 2.1 48.145 2.36 ;
      RECT 45.62 3.635 45.88 3.895 ;
      RECT 47.915 3.125 47.92 3.335 ;
      RECT 47.92 3.13 47.93 3.33 ;
      RECT 47.87 3.125 47.915 3.35 ;
      RECT 47.86 3.125 47.87 3.37 ;
      RECT 47.841 3.125 47.86 3.375 ;
      RECT 47.755 3.125 47.841 3.372 ;
      RECT 47.725 3.127 47.755 3.37 ;
      RECT 47.67 3.137 47.725 3.368 ;
      RECT 47.605 3.151 47.67 3.366 ;
      RECT 47.6 3.159 47.605 3.365 ;
      RECT 47.585 3.162 47.6 3.363 ;
      RECT 47.52 3.172 47.585 3.359 ;
      RECT 47.472 3.186 47.52 3.36 ;
      RECT 47.386 3.203 47.472 3.374 ;
      RECT 47.3 3.224 47.386 3.391 ;
      RECT 47.28 3.237 47.3 3.401 ;
      RECT 47.235 3.245 47.28 3.408 ;
      RECT 47.2 3.253 47.235 3.416 ;
      RECT 47.166 3.261 47.2 3.424 ;
      RECT 47.08 3.275 47.166 3.436 ;
      RECT 47.045 3.292 47.08 3.448 ;
      RECT 47.036 3.301 47.045 3.452 ;
      RECT 46.95 3.319 47.036 3.469 ;
      RECT 46.891 3.346 46.95 3.496 ;
      RECT 46.805 3.373 46.891 3.524 ;
      RECT 46.785 3.395 46.805 3.544 ;
      RECT 46.725 3.41 46.785 3.56 ;
      RECT 46.715 3.422 46.725 3.573 ;
      RECT 46.71 3.427 46.715 3.576 ;
      RECT 46.7 3.43 46.71 3.579 ;
      RECT 46.695 3.432 46.7 3.582 ;
      RECT 46.665 3.44 46.695 3.589 ;
      RECT 46.65 3.447 46.665 3.597 ;
      RECT 46.64 3.452 46.65 3.601 ;
      RECT 46.635 3.455 46.64 3.604 ;
      RECT 46.625 3.457 46.635 3.607 ;
      RECT 46.59 3.467 46.625 3.616 ;
      RECT 46.515 3.49 46.59 3.638 ;
      RECT 46.495 3.508 46.515 3.656 ;
      RECT 46.465 3.515 46.495 3.666 ;
      RECT 46.445 3.523 46.465 3.676 ;
      RECT 46.435 3.529 46.445 3.683 ;
      RECT 46.416 3.534 46.435 3.689 ;
      RECT 46.33 3.554 46.416 3.709 ;
      RECT 46.315 3.574 46.33 3.728 ;
      RECT 46.27 3.586 46.315 3.739 ;
      RECT 46.205 3.607 46.27 3.762 ;
      RECT 46.165 3.627 46.205 3.783 ;
      RECT 46.155 3.637 46.165 3.793 ;
      RECT 46.105 3.649 46.155 3.804 ;
      RECT 46.085 3.665 46.105 3.816 ;
      RECT 46.055 3.675 46.085 3.822 ;
      RECT 46.045 3.68 46.055 3.824 ;
      RECT 45.976 3.681 46.045 3.83 ;
      RECT 45.89 3.683 45.976 3.84 ;
      RECT 45.88 3.684 45.89 3.845 ;
      RECT 47.15 3.71 47.34 3.92 ;
      RECT 47.14 3.715 47.35 3.913 ;
      RECT 47.125 3.715 47.35 3.878 ;
      RECT 47.045 3.6 47.305 3.86 ;
      RECT 45.96 3.13 46.145 3.425 ;
      RECT 45.95 3.13 46.145 3.423 ;
      RECT 45.935 3.13 46.15 3.418 ;
      RECT 45.935 3.13 46.155 3.415 ;
      RECT 45.93 3.13 46.155 3.413 ;
      RECT 45.925 3.385 46.155 3.403 ;
      RECT 45.93 3.13 46.19 3.39 ;
      RECT 45.89 2.165 46.15 2.425 ;
      RECT 45.7 2.09 45.786 2.423 ;
      RECT 45.675 2.094 45.83 2.419 ;
      RECT 45.786 2.086 45.83 2.419 ;
      RECT 45.786 2.087 45.835 2.418 ;
      RECT 45.7 2.092 45.85 2.417 ;
      RECT 45.675 2.1 45.89 2.416 ;
      RECT 45.67 2.095 45.85 2.411 ;
      RECT 45.66 2.11 45.89 2.318 ;
      RECT 45.66 2.162 46.09 2.318 ;
      RECT 45.66 2.155 46.07 2.318 ;
      RECT 45.66 2.142 46.04 2.318 ;
      RECT 45.66 2.13 45.98 2.318 ;
      RECT 45.66 2.115 45.955 2.318 ;
      RECT 44.86 2.745 44.995 3.04 ;
      RECT 45.12 2.768 45.125 2.955 ;
      RECT 45.84 2.665 45.985 2.9 ;
      RECT 46 2.665 46.005 2.89 ;
      RECT 46.035 2.676 46.04 2.87 ;
      RECT 46.03 2.668 46.035 2.875 ;
      RECT 46.01 2.665 46.03 2.88 ;
      RECT 46.005 2.665 46.01 2.888 ;
      RECT 45.995 2.665 46 2.893 ;
      RECT 45.985 2.665 45.995 2.898 ;
      RECT 45.815 2.667 45.84 2.9 ;
      RECT 45.765 2.674 45.815 2.9 ;
      RECT 45.76 2.679 45.765 2.9 ;
      RECT 45.721 2.684 45.76 2.901 ;
      RECT 45.635 2.696 45.721 2.902 ;
      RECT 45.626 2.706 45.635 2.902 ;
      RECT 45.54 2.715 45.626 2.904 ;
      RECT 45.516 2.725 45.54 2.906 ;
      RECT 45.43 2.736 45.516 2.907 ;
      RECT 45.4 2.747 45.43 2.909 ;
      RECT 45.37 2.752 45.4 2.911 ;
      RECT 45.345 2.758 45.37 2.914 ;
      RECT 45.33 2.763 45.345 2.915 ;
      RECT 45.285 2.769 45.33 2.915 ;
      RECT 45.28 2.774 45.285 2.916 ;
      RECT 45.26 2.774 45.28 2.918 ;
      RECT 45.24 2.772 45.26 2.923 ;
      RECT 45.205 2.771 45.24 2.93 ;
      RECT 45.175 2.77 45.205 2.94 ;
      RECT 45.125 2.769 45.175 2.95 ;
      RECT 45.035 2.766 45.12 3.04 ;
      RECT 45.01 2.76 45.035 3.04 ;
      RECT 44.995 2.75 45.01 3.04 ;
      RECT 44.81 2.745 44.86 2.96 ;
      RECT 44.8 2.75 44.81 2.95 ;
      RECT 45.04 3.225 45.3 3.485 ;
      RECT 45.04 3.225 45.33 3.378 ;
      RECT 45.04 3.225 45.365 3.363 ;
      RECT 45.295 3.145 45.485 3.355 ;
      RECT 45.285 3.15 45.495 3.348 ;
      RECT 45.25 3.22 45.495 3.348 ;
      RECT 45.28 3.162 45.3 3.485 ;
      RECT 45.265 3.21 45.495 3.348 ;
      RECT 45.27 3.182 45.3 3.485 ;
      RECT 44.35 2.25 44.42 3.355 ;
      RECT 45.085 2.355 45.345 2.615 ;
      RECT 44.665 2.401 44.68 2.61 ;
      RECT 45.001 2.414 45.085 2.565 ;
      RECT 44.915 2.411 45.001 2.565 ;
      RECT 44.876 2.409 44.915 2.565 ;
      RECT 44.79 2.407 44.876 2.565 ;
      RECT 44.73 2.405 44.79 2.576 ;
      RECT 44.695 2.403 44.73 2.594 ;
      RECT 44.68 2.401 44.695 2.605 ;
      RECT 44.65 2.401 44.665 2.618 ;
      RECT 44.64 2.401 44.65 2.623 ;
      RECT 44.615 2.4 44.64 2.628 ;
      RECT 44.6 2.395 44.615 2.634 ;
      RECT 44.595 2.388 44.6 2.639 ;
      RECT 44.57 2.379 44.595 2.645 ;
      RECT 44.525 2.358 44.57 2.658 ;
      RECT 44.515 2.342 44.525 2.668 ;
      RECT 44.5 2.335 44.515 2.678 ;
      RECT 44.49 2.328 44.5 2.695 ;
      RECT 44.485 2.325 44.49 2.725 ;
      RECT 44.48 2.323 44.485 2.755 ;
      RECT 44.475 2.321 44.48 2.792 ;
      RECT 44.46 2.317 44.475 2.859 ;
      RECT 44.46 3.15 44.47 3.35 ;
      RECT 44.455 2.313 44.46 2.985 ;
      RECT 44.455 3.137 44.46 3.355 ;
      RECT 44.45 2.311 44.455 3.07 ;
      RECT 44.45 3.127 44.455 3.355 ;
      RECT 44.435 2.282 44.45 3.355 ;
      RECT 44.42 2.255 44.435 3.355 ;
      RECT 44.345 2.25 44.35 2.605 ;
      RECT 44.345 2.66 44.35 3.355 ;
      RECT 44.33 2.25 44.345 2.583 ;
      RECT 44.34 2.682 44.345 3.355 ;
      RECT 44.33 2.722 44.34 3.355 ;
      RECT 44.295 2.25 44.33 2.525 ;
      RECT 44.325 2.757 44.33 3.355 ;
      RECT 44.31 2.812 44.325 3.355 ;
      RECT 44.305 2.877 44.31 3.355 ;
      RECT 44.29 2.925 44.305 3.355 ;
      RECT 44.265 2.25 44.295 2.48 ;
      RECT 44.285 2.98 44.29 3.355 ;
      RECT 44.27 3.04 44.285 3.355 ;
      RECT 44.265 3.088 44.27 3.353 ;
      RECT 44.26 2.25 44.265 2.473 ;
      RECT 44.26 3.12 44.265 3.348 ;
      RECT 44.235 2.25 44.26 2.465 ;
      RECT 44.225 2.255 44.235 2.455 ;
      RECT 44.44 3.53 44.46 3.77 ;
      RECT 43.67 3.46 43.675 3.67 ;
      RECT 44.95 3.533 44.96 3.728 ;
      RECT 44.945 3.523 44.95 3.731 ;
      RECT 44.865 3.52 44.945 3.754 ;
      RECT 44.861 3.52 44.865 3.776 ;
      RECT 44.775 3.52 44.861 3.786 ;
      RECT 44.76 3.52 44.775 3.794 ;
      RECT 44.731 3.521 44.76 3.792 ;
      RECT 44.645 3.526 44.731 3.788 ;
      RECT 44.632 3.53 44.645 3.784 ;
      RECT 44.546 3.53 44.632 3.78 ;
      RECT 44.46 3.53 44.546 3.774 ;
      RECT 44.376 3.53 44.44 3.768 ;
      RECT 44.29 3.53 44.376 3.763 ;
      RECT 44.27 3.53 44.29 3.759 ;
      RECT 44.21 3.525 44.27 3.756 ;
      RECT 44.182 3.519 44.21 3.753 ;
      RECT 44.096 3.514 44.182 3.749 ;
      RECT 44.01 3.508 44.096 3.743 ;
      RECT 43.935 3.49 44.01 3.738 ;
      RECT 43.9 3.467 43.935 3.734 ;
      RECT 43.89 3.457 43.9 3.733 ;
      RECT 43.835 3.455 43.89 3.732 ;
      RECT 43.76 3.455 43.835 3.728 ;
      RECT 43.75 3.455 43.76 3.723 ;
      RECT 43.735 3.455 43.75 3.715 ;
      RECT 43.685 3.457 43.735 3.693 ;
      RECT 43.675 3.46 43.685 3.673 ;
      RECT 43.665 3.465 43.67 3.668 ;
      RECT 43.66 3.47 43.665 3.663 ;
      RECT 43.785 2.635 44.045 2.895 ;
      RECT 43.785 2.65 44.065 2.86 ;
      RECT 43.785 2.655 44.075 2.855 ;
      RECT 41.77 2.115 42.03 2.375 ;
      RECT 41.76 2.145 42.03 2.355 ;
      RECT 43.68 2.06 43.94 2.32 ;
      RECT 43.675 2.135 43.68 2.321 ;
      RECT 43.65 2.14 43.675 2.323 ;
      RECT 43.635 2.147 43.65 2.326 ;
      RECT 43.575 2.165 43.635 2.331 ;
      RECT 43.545 2.185 43.575 2.338 ;
      RECT 43.52 2.193 43.545 2.343 ;
      RECT 43.495 2.201 43.52 2.345 ;
      RECT 43.477 2.205 43.495 2.344 ;
      RECT 43.391 2.203 43.477 2.344 ;
      RECT 43.305 2.201 43.391 2.344 ;
      RECT 43.219 2.199 43.305 2.343 ;
      RECT 43.133 2.197 43.219 2.343 ;
      RECT 43.047 2.195 43.133 2.343 ;
      RECT 42.961 2.193 43.047 2.343 ;
      RECT 42.875 2.191 42.961 2.342 ;
      RECT 42.857 2.19 42.875 2.342 ;
      RECT 42.771 2.189 42.857 2.342 ;
      RECT 42.685 2.187 42.771 2.342 ;
      RECT 42.599 2.186 42.685 2.341 ;
      RECT 42.513 2.185 42.599 2.341 ;
      RECT 42.427 2.183 42.513 2.341 ;
      RECT 42.341 2.182 42.427 2.341 ;
      RECT 42.255 2.18 42.341 2.34 ;
      RECT 42.231 2.178 42.255 2.34 ;
      RECT 42.145 2.171 42.231 2.34 ;
      RECT 42.116 2.163 42.145 2.34 ;
      RECT 42.03 2.155 42.116 2.34 ;
      RECT 41.75 2.152 41.76 2.35 ;
      RECT 43.255 3.115 43.26 3.465 ;
      RECT 43.025 3.205 43.165 3.465 ;
      RECT 43.5 2.89 43.545 3.1 ;
      RECT 43.555 2.901 43.565 3.095 ;
      RECT 43.545 2.893 43.555 3.1 ;
      RECT 43.48 2.89 43.5 3.105 ;
      RECT 43.45 2.89 43.48 3.128 ;
      RECT 43.44 2.89 43.45 3.153 ;
      RECT 43.435 2.89 43.44 3.163 ;
      RECT 43.38 2.89 43.435 3.203 ;
      RECT 43.375 2.89 43.38 3.243 ;
      RECT 43.37 2.892 43.375 3.248 ;
      RECT 43.355 2.902 43.37 3.259 ;
      RECT 43.31 2.96 43.355 3.295 ;
      RECT 43.3 3.015 43.31 3.329 ;
      RECT 43.285 3.042 43.3 3.345 ;
      RECT 43.275 3.069 43.285 3.465 ;
      RECT 43.26 3.092 43.275 3.465 ;
      RECT 43.25 3.132 43.255 3.465 ;
      RECT 43.245 3.142 43.25 3.465 ;
      RECT 43.24 3.157 43.245 3.465 ;
      RECT 43.23 3.162 43.24 3.465 ;
      RECT 43.165 3.185 43.23 3.465 ;
      RECT 42.665 2.68 42.855 2.89 ;
      RECT 41.24 2.605 41.5 2.865 ;
      RECT 41.59 2.6 41.685 2.81 ;
      RECT 41.565 2.615 41.575 2.81 ;
      RECT 42.855 2.687 42.865 2.885 ;
      RECT 42.655 2.687 42.665 2.885 ;
      RECT 42.64 2.702 42.655 2.875 ;
      RECT 42.635 2.71 42.64 2.868 ;
      RECT 42.625 2.713 42.635 2.865 ;
      RECT 42.59 2.712 42.625 2.863 ;
      RECT 42.561 2.708 42.59 2.86 ;
      RECT 42.475 2.703 42.561 2.857 ;
      RECT 42.415 2.697 42.475 2.853 ;
      RECT 42.386 2.693 42.415 2.85 ;
      RECT 42.3 2.685 42.386 2.847 ;
      RECT 42.291 2.679 42.3 2.845 ;
      RECT 42.205 2.674 42.291 2.843 ;
      RECT 42.182 2.669 42.205 2.84 ;
      RECT 42.096 2.663 42.182 2.837 ;
      RECT 42.01 2.654 42.096 2.832 ;
      RECT 42 2.649 42.01 2.83 ;
      RECT 41.981 2.648 42 2.829 ;
      RECT 41.895 2.643 41.981 2.825 ;
      RECT 41.875 2.638 41.895 2.821 ;
      RECT 41.815 2.633 41.875 2.818 ;
      RECT 41.79 2.623 41.815 2.816 ;
      RECT 41.785 2.616 41.79 2.815 ;
      RECT 41.775 2.607 41.785 2.814 ;
      RECT 41.771 2.6 41.775 2.814 ;
      RECT 41.685 2.6 41.771 2.812 ;
      RECT 41.575 2.607 41.59 2.81 ;
      RECT 41.56 2.617 41.565 2.81 ;
      RECT 41.54 2.62 41.56 2.807 ;
      RECT 41.51 2.62 41.54 2.803 ;
      RECT 41.5 2.62 41.51 2.803 ;
      RECT 42.415 3.115 42.675 3.375 ;
      RECT 42.345 3.125 42.675 3.335 ;
      RECT 42.335 3.132 42.675 3.33 ;
      RECT 41.755 3.12 42.015 3.38 ;
      RECT 41.755 3.16 42.12 3.37 ;
      RECT 41.755 3.162 42.125 3.369 ;
      RECT 41.755 3.17 42.13 3.366 ;
      RECT 40.68 2.245 40.78 3.77 ;
      RECT 40.87 3.385 40.92 3.645 ;
      RECT 40.865 2.258 40.87 2.445 ;
      RECT 40.86 3.366 40.87 3.645 ;
      RECT 40.86 2.255 40.865 2.453 ;
      RECT 40.845 2.249 40.86 2.46 ;
      RECT 40.855 3.354 40.86 3.728 ;
      RECT 40.845 3.342 40.855 3.765 ;
      RECT 40.835 2.245 40.845 2.467 ;
      RECT 40.835 3.327 40.845 3.77 ;
      RECT 40.83 2.245 40.835 2.475 ;
      RECT 40.81 3.297 40.835 3.77 ;
      RECT 40.79 2.245 40.83 2.523 ;
      RECT 40.8 3.257 40.81 3.77 ;
      RECT 40.79 3.212 40.8 3.77 ;
      RECT 40.785 2.245 40.79 2.593 ;
      RECT 40.785 3.17 40.79 3.77 ;
      RECT 40.78 2.245 40.785 3.07 ;
      RECT 40.78 3.152 40.785 3.77 ;
      RECT 40.67 2.248 40.68 3.77 ;
      RECT 40.655 2.255 40.67 3.766 ;
      RECT 40.65 2.265 40.655 3.761 ;
      RECT 40.645 2.465 40.65 3.653 ;
      RECT 40.64 2.55 40.645 3.205 ;
      RECT 39.515 7.77 39.805 8 ;
      RECT 39.575 6.29 39.745 8 ;
      RECT 39.565 6.66 39.92 7.015 ;
      RECT 39.515 6.29 39.805 6.52 ;
      RECT 39.11 2.395 39.215 2.965 ;
      RECT 39.11 2.73 39.435 2.96 ;
      RECT 39.11 2.76 39.605 2.93 ;
      RECT 39.11 2.395 39.3 2.96 ;
      RECT 38.525 2.36 38.815 2.59 ;
      RECT 38.525 2.395 39.3 2.565 ;
      RECT 38.585 0.88 38.755 2.59 ;
      RECT 38.525 0.88 38.815 1.11 ;
      RECT 38.525 7.77 38.815 8 ;
      RECT 38.585 6.29 38.755 8 ;
      RECT 38.525 6.29 38.815 6.52 ;
      RECT 38.525 6.325 39.38 6.485 ;
      RECT 39.21 5.92 39.38 6.485 ;
      RECT 38.525 6.32 38.92 6.485 ;
      RECT 39.145 5.92 39.435 6.15 ;
      RECT 39.145 5.95 39.605 6.12 ;
      RECT 38.155 2.73 38.445 2.96 ;
      RECT 38.155 2.76 38.615 2.93 ;
      RECT 38.22 1.655 38.385 2.96 ;
      RECT 36.735 1.625 37.025 1.855 ;
      RECT 36.735 1.655 38.385 1.825 ;
      RECT 36.795 0.885 36.965 1.855 ;
      RECT 36.735 0.885 37.025 1.115 ;
      RECT 36.735 7.765 37.025 7.995 ;
      RECT 36.795 7.025 36.965 7.995 ;
      RECT 36.795 7.12 38.385 7.29 ;
      RECT 38.215 5.92 38.385 7.29 ;
      RECT 36.735 7.025 37.025 7.255 ;
      RECT 38.155 5.92 38.445 6.15 ;
      RECT 38.155 5.95 38.615 6.12 ;
      RECT 34.77 3.43 35.12 3.78 ;
      RECT 34.86 2.025 35.03 3.78 ;
      RECT 37.165 1.965 37.515 2.315 ;
      RECT 34.86 2.025 36.48 2.2 ;
      RECT 34.86 2.025 37.515 2.195 ;
      RECT 37.19 6.655 37.515 6.98 ;
      RECT 32.615 6.61 32.965 6.96 ;
      RECT 37.165 6.655 37.515 6.885 ;
      RECT 32.405 6.655 32.965 6.885 ;
      RECT 32.235 6.685 37.515 6.855 ;
      RECT 36.39 2.365 36.71 2.685 ;
      RECT 36.36 2.365 36.71 2.595 ;
      RECT 36.19 2.395 36.71 2.565 ;
      RECT 36.39 6.225 36.71 6.545 ;
      RECT 36.36 6.285 36.71 6.515 ;
      RECT 36.19 6.315 36.71 6.485 ;
      RECT 32.17 3.665 32.21 3.925 ;
      RECT 32.21 3.645 32.215 3.655 ;
      RECT 33.54 2.89 33.55 3.111 ;
      RECT 33.47 2.885 33.54 3.236 ;
      RECT 33.46 2.885 33.47 3.363 ;
      RECT 33.435 2.885 33.46 3.41 ;
      RECT 33.41 2.885 33.435 3.488 ;
      RECT 33.39 2.885 33.41 3.558 ;
      RECT 33.365 2.885 33.39 3.598 ;
      RECT 33.355 2.885 33.365 3.618 ;
      RECT 33.345 2.887 33.355 3.626 ;
      RECT 33.34 2.892 33.345 3.083 ;
      RECT 33.34 3.092 33.345 3.627 ;
      RECT 33.335 3.137 33.34 3.628 ;
      RECT 33.325 3.202 33.335 3.629 ;
      RECT 33.315 3.297 33.325 3.631 ;
      RECT 33.31 3.35 33.315 3.633 ;
      RECT 33.305 3.37 33.31 3.634 ;
      RECT 33.25 3.395 33.305 3.64 ;
      RECT 33.21 3.43 33.25 3.649 ;
      RECT 33.2 3.447 33.21 3.654 ;
      RECT 33.191 3.453 33.2 3.656 ;
      RECT 33.105 3.491 33.191 3.667 ;
      RECT 33.1 3.53 33.105 3.677 ;
      RECT 33.025 3.537 33.1 3.687 ;
      RECT 33.005 3.547 33.025 3.698 ;
      RECT 32.975 3.554 33.005 3.706 ;
      RECT 32.95 3.561 32.975 3.713 ;
      RECT 32.926 3.567 32.95 3.718 ;
      RECT 32.84 3.58 32.926 3.73 ;
      RECT 32.762 3.587 32.84 3.748 ;
      RECT 32.676 3.582 32.762 3.766 ;
      RECT 32.59 3.577 32.676 3.786 ;
      RECT 32.51 3.571 32.59 3.803 ;
      RECT 32.445 3.567 32.51 3.832 ;
      RECT 32.44 3.281 32.445 3.305 ;
      RECT 32.43 3.557 32.445 3.86 ;
      RECT 32.435 3.275 32.44 3.345 ;
      RECT 32.43 3.269 32.435 3.415 ;
      RECT 32.425 3.263 32.43 3.493 ;
      RECT 32.425 3.54 32.43 3.925 ;
      RECT 32.417 3.26 32.425 3.925 ;
      RECT 32.331 3.258 32.417 3.925 ;
      RECT 32.245 3.256 32.331 3.925 ;
      RECT 32.235 3.257 32.245 3.925 ;
      RECT 32.23 3.262 32.235 3.925 ;
      RECT 32.22 3.275 32.23 3.925 ;
      RECT 32.215 3.297 32.22 3.925 ;
      RECT 32.21 3.657 32.215 3.925 ;
      RECT 32.84 3.125 32.845 3.345 ;
      RECT 33.345 2.16 33.38 2.42 ;
      RECT 33.33 2.16 33.345 2.428 ;
      RECT 33.301 2.16 33.33 2.45 ;
      RECT 33.215 2.16 33.301 2.51 ;
      RECT 33.195 2.16 33.215 2.575 ;
      RECT 33.135 2.16 33.195 2.74 ;
      RECT 33.13 2.16 33.135 2.888 ;
      RECT 33.125 2.16 33.13 2.9 ;
      RECT 33.12 2.16 33.125 2.926 ;
      RECT 33.09 2.346 33.12 3.006 ;
      RECT 33.085 2.394 33.09 3.095 ;
      RECT 33.08 2.408 33.085 3.11 ;
      RECT 33.075 2.427 33.08 3.14 ;
      RECT 33.07 2.442 33.075 3.156 ;
      RECT 33.065 2.457 33.07 3.178 ;
      RECT 33.06 2.477 33.065 3.2 ;
      RECT 33.05 2.497 33.06 3.233 ;
      RECT 33.035 2.539 33.05 3.295 ;
      RECT 33.03 2.57 33.035 3.335 ;
      RECT 33.025 2.582 33.03 3.34 ;
      RECT 33.02 2.594 33.025 3.345 ;
      RECT 33.015 2.607 33.02 3.345 ;
      RECT 33.01 2.625 33.015 3.345 ;
      RECT 33.005 2.645 33.01 3.345 ;
      RECT 33 2.657 33.005 3.345 ;
      RECT 32.995 2.67 33 3.345 ;
      RECT 32.975 2.705 32.995 3.345 ;
      RECT 32.925 2.807 32.975 3.345 ;
      RECT 32.92 2.892 32.925 3.345 ;
      RECT 32.915 2.9 32.92 3.345 ;
      RECT 32.91 2.917 32.915 3.345 ;
      RECT 32.905 2.932 32.91 3.345 ;
      RECT 32.87 2.997 32.905 3.345 ;
      RECT 32.855 3.062 32.87 3.345 ;
      RECT 32.85 3.092 32.855 3.345 ;
      RECT 32.845 3.117 32.85 3.345 ;
      RECT 32.83 3.127 32.84 3.345 ;
      RECT 32.815 3.14 32.83 3.338 ;
      RECT 32.56 2.73 32.63 2.94 ;
      RECT 32.35 2.707 32.355 2.9 ;
      RECT 29.805 2.635 30.065 2.895 ;
      RECT 32.64 2.917 32.645 2.92 ;
      RECT 32.63 2.735 32.64 2.935 ;
      RECT 32.531 2.728 32.56 2.94 ;
      RECT 32.445 2.72 32.531 2.94 ;
      RECT 32.43 2.714 32.445 2.938 ;
      RECT 32.41 2.713 32.43 2.925 ;
      RECT 32.405 2.712 32.41 2.908 ;
      RECT 32.355 2.709 32.405 2.903 ;
      RECT 32.325 2.706 32.35 2.898 ;
      RECT 32.305 2.704 32.325 2.893 ;
      RECT 32.29 2.702 32.305 2.89 ;
      RECT 32.26 2.7 32.29 2.888 ;
      RECT 32.195 2.696 32.26 2.88 ;
      RECT 32.165 2.691 32.195 2.875 ;
      RECT 32.145 2.689 32.165 2.873 ;
      RECT 32.115 2.686 32.145 2.868 ;
      RECT 32.055 2.682 32.115 2.86 ;
      RECT 32.05 2.679 32.055 2.855 ;
      RECT 31.98 2.677 32.05 2.85 ;
      RECT 31.951 2.673 31.98 2.843 ;
      RECT 31.865 2.668 31.951 2.835 ;
      RECT 31.831 2.663 31.865 2.827 ;
      RECT 31.745 2.655 31.831 2.819 ;
      RECT 31.706 2.648 31.745 2.811 ;
      RECT 31.62 2.643 31.706 2.803 ;
      RECT 31.555 2.637 31.62 2.793 ;
      RECT 31.535 2.632 31.555 2.788 ;
      RECT 31.526 2.629 31.535 2.787 ;
      RECT 31.44 2.625 31.526 2.781 ;
      RECT 31.4 2.621 31.44 2.773 ;
      RECT 31.38 2.617 31.4 2.771 ;
      RECT 31.32 2.617 31.38 2.768 ;
      RECT 31.3 2.62 31.32 2.766 ;
      RECT 31.279 2.62 31.3 2.766 ;
      RECT 31.193 2.622 31.279 2.77 ;
      RECT 31.107 2.624 31.193 2.776 ;
      RECT 31.021 2.626 31.107 2.783 ;
      RECT 30.935 2.629 31.021 2.789 ;
      RECT 30.901 2.63 30.935 2.794 ;
      RECT 30.815 2.633 30.901 2.799 ;
      RECT 30.786 2.64 30.815 2.804 ;
      RECT 30.7 2.64 30.786 2.809 ;
      RECT 30.667 2.64 30.7 2.814 ;
      RECT 30.581 2.642 30.667 2.819 ;
      RECT 30.495 2.644 30.581 2.826 ;
      RECT 30.431 2.646 30.495 2.832 ;
      RECT 30.345 2.648 30.431 2.838 ;
      RECT 30.342 2.65 30.345 2.841 ;
      RECT 30.256 2.651 30.342 2.845 ;
      RECT 30.17 2.654 30.256 2.852 ;
      RECT 30.151 2.656 30.17 2.856 ;
      RECT 30.065 2.658 30.151 2.861 ;
      RECT 29.795 2.67 29.805 2.865 ;
      RECT 31.975 7.765 32.265 7.995 ;
      RECT 32.035 7.025 32.205 7.995 ;
      RECT 31.925 7.055 32.3 7.425 ;
      RECT 31.975 7.025 32.265 7.425 ;
      RECT 32.03 2.25 32.215 2.46 ;
      RECT 32.025 2.251 32.22 2.458 ;
      RECT 32.02 2.256 32.23 2.453 ;
      RECT 32.015 2.232 32.02 2.45 ;
      RECT 31.985 2.229 32.015 2.443 ;
      RECT 31.98 2.225 31.985 2.434 ;
      RECT 31.945 2.256 32.23 2.429 ;
      RECT 31.72 2.165 31.98 2.425 ;
      RECT 32.02 2.234 32.025 2.453 ;
      RECT 32.025 2.235 32.03 2.458 ;
      RECT 31.72 2.247 32.1 2.425 ;
      RECT 31.72 2.245 32.085 2.425 ;
      RECT 31.72 2.24 32.075 2.425 ;
      RECT 31.675 3.155 31.725 3.44 ;
      RECT 31.62 3.125 31.625 3.44 ;
      RECT 31.59 3.105 31.595 3.44 ;
      RECT 31.74 3.155 31.8 3.415 ;
      RECT 31.735 3.155 31.74 3.423 ;
      RECT 31.725 3.155 31.735 3.435 ;
      RECT 31.64 3.145 31.675 3.44 ;
      RECT 31.635 3.132 31.64 3.44 ;
      RECT 31.625 3.127 31.635 3.44 ;
      RECT 31.605 3.117 31.62 3.44 ;
      RECT 31.595 3.11 31.605 3.44 ;
      RECT 31.585 3.102 31.59 3.44 ;
      RECT 31.555 3.092 31.585 3.44 ;
      RECT 31.54 3.08 31.555 3.44 ;
      RECT 31.525 3.07 31.54 3.435 ;
      RECT 31.505 3.06 31.525 3.41 ;
      RECT 31.495 3.052 31.505 3.387 ;
      RECT 31.465 3.035 31.495 3.377 ;
      RECT 31.46 3.012 31.465 3.368 ;
      RECT 31.455 2.999 31.46 3.366 ;
      RECT 31.44 2.975 31.455 3.36 ;
      RECT 31.435 2.951 31.44 3.354 ;
      RECT 31.425 2.94 31.435 3.349 ;
      RECT 31.42 2.93 31.425 3.345 ;
      RECT 31.415 2.922 31.42 3.342 ;
      RECT 31.405 2.917 31.415 3.338 ;
      RECT 31.4 2.912 31.405 3.334 ;
      RECT 31.315 2.91 31.4 3.309 ;
      RECT 31.285 2.91 31.315 3.275 ;
      RECT 31.27 2.91 31.285 3.258 ;
      RECT 31.215 2.91 31.27 3.203 ;
      RECT 31.21 2.915 31.215 3.152 ;
      RECT 31.2 2.92 31.21 3.142 ;
      RECT 31.195 2.93 31.2 3.128 ;
      RECT 31.145 3.67 31.405 3.93 ;
      RECT 31.065 3.685 31.405 3.906 ;
      RECT 31.045 3.685 31.405 3.901 ;
      RECT 31.021 3.685 31.405 3.899 ;
      RECT 30.935 3.685 31.405 3.894 ;
      RECT 30.785 3.625 31.045 3.89 ;
      RECT 30.74 3.685 31.405 3.885 ;
      RECT 30.735 3.692 31.405 3.88 ;
      RECT 30.75 3.68 31.065 3.89 ;
      RECT 30.64 2.115 30.9 2.375 ;
      RECT 30.64 2.172 30.905 2.368 ;
      RECT 30.64 2.202 30.91 2.3 ;
      RECT 30.7 2.633 30.815 2.635 ;
      RECT 30.786 2.63 30.815 2.635 ;
      RECT 29.81 3.634 29.835 3.874 ;
      RECT 29.795 3.637 29.885 3.868 ;
      RECT 29.79 3.642 29.971 3.863 ;
      RECT 29.785 3.65 30.035 3.861 ;
      RECT 29.785 3.65 30.045 3.86 ;
      RECT 29.78 3.657 30.055 3.853 ;
      RECT 29.78 3.657 30.141 3.842 ;
      RECT 29.775 3.692 30.141 3.838 ;
      RECT 29.775 3.692 30.15 3.827 ;
      RECT 30.055 3.565 30.315 3.825 ;
      RECT 29.765 3.742 30.315 3.823 ;
      RECT 30.035 3.61 30.055 3.858 ;
      RECT 29.971 3.613 30.035 3.862 ;
      RECT 29.885 3.618 29.971 3.867 ;
      RECT 29.815 3.629 30.315 3.825 ;
      RECT 29.835 3.623 29.885 3.872 ;
      RECT 29.96 2.1 29.97 2.362 ;
      RECT 29.95 2.157 29.96 2.365 ;
      RECT 29.925 2.162 29.95 2.371 ;
      RECT 29.9 2.166 29.925 2.383 ;
      RECT 29.89 2.169 29.9 2.393 ;
      RECT 29.885 2.17 29.89 2.398 ;
      RECT 29.88 2.171 29.885 2.403 ;
      RECT 29.875 2.172 29.88 2.405 ;
      RECT 29.85 2.175 29.875 2.408 ;
      RECT 29.82 2.181 29.85 2.411 ;
      RECT 29.755 2.192 29.82 2.414 ;
      RECT 29.71 2.2 29.755 2.418 ;
      RECT 29.695 2.2 29.71 2.426 ;
      RECT 29.69 2.201 29.695 2.433 ;
      RECT 29.685 2.203 29.69 2.436 ;
      RECT 29.68 2.207 29.685 2.439 ;
      RECT 29.67 2.215 29.68 2.443 ;
      RECT 29.665 2.228 29.67 2.448 ;
      RECT 29.66 2.236 29.665 2.45 ;
      RECT 29.655 2.242 29.66 2.45 ;
      RECT 29.65 2.246 29.655 2.453 ;
      RECT 29.645 2.248 29.65 2.456 ;
      RECT 29.64 2.251 29.645 2.459 ;
      RECT 29.63 2.256 29.64 2.463 ;
      RECT 29.625 2.262 29.63 2.468 ;
      RECT 29.615 2.268 29.625 2.472 ;
      RECT 29.6 2.275 29.615 2.478 ;
      RECT 29.571 2.289 29.6 2.488 ;
      RECT 29.485 2.324 29.571 2.52 ;
      RECT 29.465 2.357 29.485 2.549 ;
      RECT 29.445 2.37 29.465 2.56 ;
      RECT 29.425 2.382 29.445 2.571 ;
      RECT 29.375 2.404 29.425 2.591 ;
      RECT 29.36 2.422 29.375 2.608 ;
      RECT 29.355 2.428 29.36 2.611 ;
      RECT 29.35 2.432 29.355 2.614 ;
      RECT 29.345 2.436 29.35 2.618 ;
      RECT 29.34 2.438 29.345 2.621 ;
      RECT 29.33 2.445 29.34 2.624 ;
      RECT 29.325 2.45 29.33 2.628 ;
      RECT 29.32 2.452 29.325 2.631 ;
      RECT 29.315 2.456 29.32 2.634 ;
      RECT 29.31 2.458 29.315 2.638 ;
      RECT 29.295 2.463 29.31 2.643 ;
      RECT 29.29 2.468 29.295 2.646 ;
      RECT 29.285 2.476 29.29 2.649 ;
      RECT 29.28 2.478 29.285 2.652 ;
      RECT 29.275 2.48 29.28 2.655 ;
      RECT 29.265 2.482 29.275 2.661 ;
      RECT 29.23 2.496 29.265 2.673 ;
      RECT 29.22 2.511 29.23 2.683 ;
      RECT 29.145 2.54 29.22 2.707 ;
      RECT 29.14 2.565 29.145 2.73 ;
      RECT 29.125 2.569 29.14 2.736 ;
      RECT 29.115 2.577 29.125 2.741 ;
      RECT 29.085 2.59 29.115 2.745 ;
      RECT 29.075 2.605 29.085 2.75 ;
      RECT 29.065 2.61 29.075 2.753 ;
      RECT 29.06 2.612 29.065 2.755 ;
      RECT 29.045 2.615 29.06 2.758 ;
      RECT 29.04 2.617 29.045 2.761 ;
      RECT 29.02 2.622 29.04 2.765 ;
      RECT 28.99 2.627 29.02 2.773 ;
      RECT 28.965 2.634 28.99 2.781 ;
      RECT 28.96 2.639 28.965 2.786 ;
      RECT 28.93 2.642 28.96 2.79 ;
      RECT 28.89 2.645 28.93 2.8 ;
      RECT 28.855 2.642 28.89 2.812 ;
      RECT 28.845 2.638 28.855 2.819 ;
      RECT 28.82 2.634 28.845 2.825 ;
      RECT 28.815 2.63 28.82 2.83 ;
      RECT 28.775 2.627 28.815 2.83 ;
      RECT 28.76 2.612 28.775 2.831 ;
      RECT 28.737 2.6 28.76 2.831 ;
      RECT 28.651 2.6 28.737 2.832 ;
      RECT 28.565 2.6 28.651 2.834 ;
      RECT 28.545 2.6 28.565 2.831 ;
      RECT 28.54 2.605 28.545 2.826 ;
      RECT 28.535 2.61 28.54 2.824 ;
      RECT 28.525 2.62 28.535 2.822 ;
      RECT 28.52 2.626 28.525 2.815 ;
      RECT 28.515 2.628 28.52 2.8 ;
      RECT 28.51 2.632 28.515 2.79 ;
      RECT 29.97 2.1 30.22 2.36 ;
      RECT 27.695 3.635 27.955 3.895 ;
      RECT 29.99 3.125 29.995 3.335 ;
      RECT 29.995 3.13 30.005 3.33 ;
      RECT 29.945 3.125 29.99 3.35 ;
      RECT 29.935 3.125 29.945 3.37 ;
      RECT 29.916 3.125 29.935 3.375 ;
      RECT 29.83 3.125 29.916 3.372 ;
      RECT 29.8 3.127 29.83 3.37 ;
      RECT 29.745 3.137 29.8 3.368 ;
      RECT 29.68 3.151 29.745 3.366 ;
      RECT 29.675 3.159 29.68 3.365 ;
      RECT 29.66 3.162 29.675 3.363 ;
      RECT 29.595 3.172 29.66 3.359 ;
      RECT 29.547 3.186 29.595 3.36 ;
      RECT 29.461 3.203 29.547 3.374 ;
      RECT 29.375 3.224 29.461 3.391 ;
      RECT 29.355 3.237 29.375 3.401 ;
      RECT 29.31 3.245 29.355 3.408 ;
      RECT 29.275 3.253 29.31 3.416 ;
      RECT 29.241 3.261 29.275 3.424 ;
      RECT 29.155 3.275 29.241 3.436 ;
      RECT 29.12 3.292 29.155 3.448 ;
      RECT 29.111 3.301 29.12 3.452 ;
      RECT 29.025 3.319 29.111 3.469 ;
      RECT 28.966 3.346 29.025 3.496 ;
      RECT 28.88 3.373 28.966 3.524 ;
      RECT 28.86 3.395 28.88 3.544 ;
      RECT 28.8 3.41 28.86 3.56 ;
      RECT 28.79 3.422 28.8 3.573 ;
      RECT 28.785 3.427 28.79 3.576 ;
      RECT 28.775 3.43 28.785 3.579 ;
      RECT 28.77 3.432 28.775 3.582 ;
      RECT 28.74 3.44 28.77 3.589 ;
      RECT 28.725 3.447 28.74 3.597 ;
      RECT 28.715 3.452 28.725 3.601 ;
      RECT 28.71 3.455 28.715 3.604 ;
      RECT 28.7 3.457 28.71 3.607 ;
      RECT 28.665 3.467 28.7 3.616 ;
      RECT 28.59 3.49 28.665 3.638 ;
      RECT 28.57 3.508 28.59 3.656 ;
      RECT 28.54 3.515 28.57 3.666 ;
      RECT 28.52 3.523 28.54 3.676 ;
      RECT 28.51 3.529 28.52 3.683 ;
      RECT 28.491 3.534 28.51 3.689 ;
      RECT 28.405 3.554 28.491 3.709 ;
      RECT 28.39 3.574 28.405 3.728 ;
      RECT 28.345 3.586 28.39 3.739 ;
      RECT 28.28 3.607 28.345 3.762 ;
      RECT 28.24 3.627 28.28 3.783 ;
      RECT 28.23 3.637 28.24 3.793 ;
      RECT 28.18 3.649 28.23 3.804 ;
      RECT 28.16 3.665 28.18 3.816 ;
      RECT 28.13 3.675 28.16 3.822 ;
      RECT 28.12 3.68 28.13 3.824 ;
      RECT 28.051 3.681 28.12 3.83 ;
      RECT 27.965 3.683 28.051 3.84 ;
      RECT 27.955 3.684 27.965 3.845 ;
      RECT 29.225 3.71 29.415 3.92 ;
      RECT 29.215 3.715 29.425 3.913 ;
      RECT 29.2 3.715 29.425 3.878 ;
      RECT 29.12 3.6 29.38 3.86 ;
      RECT 28.035 3.13 28.22 3.425 ;
      RECT 28.025 3.13 28.22 3.423 ;
      RECT 28.01 3.13 28.225 3.418 ;
      RECT 28.01 3.13 28.23 3.415 ;
      RECT 28.005 3.13 28.23 3.413 ;
      RECT 28 3.385 28.23 3.403 ;
      RECT 28.005 3.13 28.265 3.39 ;
      RECT 27.965 2.165 28.225 2.425 ;
      RECT 27.775 2.09 27.861 2.423 ;
      RECT 27.75 2.094 27.905 2.419 ;
      RECT 27.861 2.086 27.905 2.419 ;
      RECT 27.861 2.087 27.91 2.418 ;
      RECT 27.775 2.092 27.925 2.417 ;
      RECT 27.75 2.1 27.965 2.416 ;
      RECT 27.745 2.095 27.925 2.411 ;
      RECT 27.735 2.11 27.965 2.318 ;
      RECT 27.735 2.162 28.165 2.318 ;
      RECT 27.735 2.155 28.145 2.318 ;
      RECT 27.735 2.142 28.115 2.318 ;
      RECT 27.735 2.13 28.055 2.318 ;
      RECT 27.735 2.115 28.03 2.318 ;
      RECT 26.935 2.745 27.07 3.04 ;
      RECT 27.195 2.768 27.2 2.955 ;
      RECT 27.915 2.665 28.06 2.9 ;
      RECT 28.075 2.665 28.08 2.89 ;
      RECT 28.11 2.676 28.115 2.87 ;
      RECT 28.105 2.668 28.11 2.875 ;
      RECT 28.085 2.665 28.105 2.88 ;
      RECT 28.08 2.665 28.085 2.888 ;
      RECT 28.07 2.665 28.075 2.893 ;
      RECT 28.06 2.665 28.07 2.898 ;
      RECT 27.89 2.667 27.915 2.9 ;
      RECT 27.84 2.674 27.89 2.9 ;
      RECT 27.835 2.679 27.84 2.9 ;
      RECT 27.796 2.684 27.835 2.901 ;
      RECT 27.71 2.696 27.796 2.902 ;
      RECT 27.701 2.706 27.71 2.902 ;
      RECT 27.615 2.715 27.701 2.904 ;
      RECT 27.591 2.725 27.615 2.906 ;
      RECT 27.505 2.736 27.591 2.907 ;
      RECT 27.475 2.747 27.505 2.909 ;
      RECT 27.445 2.752 27.475 2.911 ;
      RECT 27.42 2.758 27.445 2.914 ;
      RECT 27.405 2.763 27.42 2.915 ;
      RECT 27.36 2.769 27.405 2.915 ;
      RECT 27.355 2.774 27.36 2.916 ;
      RECT 27.335 2.774 27.355 2.918 ;
      RECT 27.315 2.772 27.335 2.923 ;
      RECT 27.28 2.771 27.315 2.93 ;
      RECT 27.25 2.77 27.28 2.94 ;
      RECT 27.2 2.769 27.25 2.95 ;
      RECT 27.11 2.766 27.195 3.04 ;
      RECT 27.085 2.76 27.11 3.04 ;
      RECT 27.07 2.75 27.085 3.04 ;
      RECT 26.885 2.745 26.935 2.96 ;
      RECT 26.875 2.75 26.885 2.95 ;
      RECT 27.115 3.225 27.375 3.485 ;
      RECT 27.115 3.225 27.405 3.378 ;
      RECT 27.115 3.225 27.44 3.363 ;
      RECT 27.37 3.145 27.56 3.355 ;
      RECT 27.36 3.15 27.57 3.348 ;
      RECT 27.325 3.22 27.57 3.348 ;
      RECT 27.355 3.162 27.375 3.485 ;
      RECT 27.34 3.21 27.57 3.348 ;
      RECT 27.345 3.182 27.375 3.485 ;
      RECT 26.425 2.25 26.495 3.355 ;
      RECT 27.16 2.355 27.42 2.615 ;
      RECT 26.74 2.401 26.755 2.61 ;
      RECT 27.076 2.414 27.16 2.565 ;
      RECT 26.99 2.411 27.076 2.565 ;
      RECT 26.951 2.409 26.99 2.565 ;
      RECT 26.865 2.407 26.951 2.565 ;
      RECT 26.805 2.405 26.865 2.576 ;
      RECT 26.77 2.403 26.805 2.594 ;
      RECT 26.755 2.401 26.77 2.605 ;
      RECT 26.725 2.401 26.74 2.618 ;
      RECT 26.715 2.401 26.725 2.623 ;
      RECT 26.69 2.4 26.715 2.628 ;
      RECT 26.675 2.395 26.69 2.634 ;
      RECT 26.67 2.388 26.675 2.639 ;
      RECT 26.645 2.379 26.67 2.645 ;
      RECT 26.6 2.358 26.645 2.658 ;
      RECT 26.59 2.342 26.6 2.668 ;
      RECT 26.575 2.335 26.59 2.678 ;
      RECT 26.565 2.328 26.575 2.695 ;
      RECT 26.56 2.325 26.565 2.725 ;
      RECT 26.555 2.323 26.56 2.755 ;
      RECT 26.55 2.321 26.555 2.792 ;
      RECT 26.535 2.317 26.55 2.859 ;
      RECT 26.535 3.15 26.545 3.35 ;
      RECT 26.53 2.313 26.535 2.985 ;
      RECT 26.53 3.137 26.535 3.355 ;
      RECT 26.525 2.311 26.53 3.07 ;
      RECT 26.525 3.127 26.53 3.355 ;
      RECT 26.51 2.282 26.525 3.355 ;
      RECT 26.495 2.255 26.51 3.355 ;
      RECT 26.42 2.25 26.425 2.605 ;
      RECT 26.42 2.66 26.425 3.355 ;
      RECT 26.405 2.25 26.42 2.583 ;
      RECT 26.415 2.682 26.42 3.355 ;
      RECT 26.405 2.722 26.415 3.355 ;
      RECT 26.37 2.25 26.405 2.525 ;
      RECT 26.4 2.757 26.405 3.355 ;
      RECT 26.385 2.812 26.4 3.355 ;
      RECT 26.38 2.877 26.385 3.355 ;
      RECT 26.365 2.925 26.38 3.355 ;
      RECT 26.34 2.25 26.37 2.48 ;
      RECT 26.36 2.98 26.365 3.355 ;
      RECT 26.345 3.04 26.36 3.355 ;
      RECT 26.34 3.088 26.345 3.353 ;
      RECT 26.335 2.25 26.34 2.473 ;
      RECT 26.335 3.12 26.34 3.348 ;
      RECT 26.31 2.25 26.335 2.465 ;
      RECT 26.3 2.255 26.31 2.455 ;
      RECT 26.515 3.53 26.535 3.77 ;
      RECT 25.745 3.46 25.75 3.67 ;
      RECT 27.025 3.533 27.035 3.728 ;
      RECT 27.02 3.523 27.025 3.731 ;
      RECT 26.94 3.52 27.02 3.754 ;
      RECT 26.936 3.52 26.94 3.776 ;
      RECT 26.85 3.52 26.936 3.786 ;
      RECT 26.835 3.52 26.85 3.794 ;
      RECT 26.806 3.521 26.835 3.792 ;
      RECT 26.72 3.526 26.806 3.788 ;
      RECT 26.707 3.53 26.72 3.784 ;
      RECT 26.621 3.53 26.707 3.78 ;
      RECT 26.535 3.53 26.621 3.774 ;
      RECT 26.451 3.53 26.515 3.768 ;
      RECT 26.365 3.53 26.451 3.763 ;
      RECT 26.345 3.53 26.365 3.759 ;
      RECT 26.285 3.525 26.345 3.756 ;
      RECT 26.257 3.519 26.285 3.753 ;
      RECT 26.171 3.514 26.257 3.749 ;
      RECT 26.085 3.508 26.171 3.743 ;
      RECT 26.01 3.49 26.085 3.738 ;
      RECT 25.975 3.467 26.01 3.734 ;
      RECT 25.965 3.457 25.975 3.733 ;
      RECT 25.91 3.455 25.965 3.732 ;
      RECT 25.835 3.455 25.91 3.728 ;
      RECT 25.825 3.455 25.835 3.723 ;
      RECT 25.81 3.455 25.825 3.715 ;
      RECT 25.76 3.457 25.81 3.693 ;
      RECT 25.75 3.46 25.76 3.673 ;
      RECT 25.74 3.465 25.745 3.668 ;
      RECT 25.735 3.47 25.74 3.663 ;
      RECT 25.86 2.635 26.12 2.895 ;
      RECT 25.86 2.65 26.14 2.86 ;
      RECT 25.86 2.655 26.15 2.855 ;
      RECT 23.845 2.115 24.105 2.375 ;
      RECT 23.835 2.145 24.105 2.355 ;
      RECT 25.755 2.06 26.015 2.32 ;
      RECT 25.75 2.135 25.755 2.321 ;
      RECT 25.725 2.14 25.75 2.323 ;
      RECT 25.71 2.147 25.725 2.326 ;
      RECT 25.65 2.165 25.71 2.331 ;
      RECT 25.62 2.185 25.65 2.338 ;
      RECT 25.595 2.193 25.62 2.343 ;
      RECT 25.57 2.201 25.595 2.345 ;
      RECT 25.552 2.205 25.57 2.344 ;
      RECT 25.466 2.203 25.552 2.344 ;
      RECT 25.38 2.201 25.466 2.344 ;
      RECT 25.294 2.199 25.38 2.343 ;
      RECT 25.208 2.197 25.294 2.343 ;
      RECT 25.122 2.195 25.208 2.343 ;
      RECT 25.036 2.193 25.122 2.343 ;
      RECT 24.95 2.191 25.036 2.342 ;
      RECT 24.932 2.19 24.95 2.342 ;
      RECT 24.846 2.189 24.932 2.342 ;
      RECT 24.76 2.187 24.846 2.342 ;
      RECT 24.674 2.186 24.76 2.341 ;
      RECT 24.588 2.185 24.674 2.341 ;
      RECT 24.502 2.183 24.588 2.341 ;
      RECT 24.416 2.182 24.502 2.341 ;
      RECT 24.33 2.18 24.416 2.34 ;
      RECT 24.306 2.178 24.33 2.34 ;
      RECT 24.22 2.171 24.306 2.34 ;
      RECT 24.191 2.163 24.22 2.34 ;
      RECT 24.105 2.155 24.191 2.34 ;
      RECT 23.825 2.152 23.835 2.35 ;
      RECT 25.33 3.115 25.335 3.465 ;
      RECT 25.1 3.205 25.24 3.465 ;
      RECT 25.575 2.89 25.62 3.1 ;
      RECT 25.63 2.901 25.64 3.095 ;
      RECT 25.62 2.893 25.63 3.1 ;
      RECT 25.555 2.89 25.575 3.105 ;
      RECT 25.525 2.89 25.555 3.128 ;
      RECT 25.515 2.89 25.525 3.153 ;
      RECT 25.51 2.89 25.515 3.163 ;
      RECT 25.455 2.89 25.51 3.203 ;
      RECT 25.45 2.89 25.455 3.243 ;
      RECT 25.445 2.892 25.45 3.248 ;
      RECT 25.43 2.902 25.445 3.259 ;
      RECT 25.385 2.96 25.43 3.295 ;
      RECT 25.375 3.015 25.385 3.329 ;
      RECT 25.36 3.042 25.375 3.345 ;
      RECT 25.35 3.069 25.36 3.465 ;
      RECT 25.335 3.092 25.35 3.465 ;
      RECT 25.325 3.132 25.33 3.465 ;
      RECT 25.32 3.142 25.325 3.465 ;
      RECT 25.315 3.157 25.32 3.465 ;
      RECT 25.305 3.162 25.315 3.465 ;
      RECT 25.24 3.185 25.305 3.465 ;
      RECT 24.74 2.68 24.93 2.89 ;
      RECT 23.315 2.605 23.575 2.865 ;
      RECT 23.665 2.6 23.76 2.81 ;
      RECT 23.64 2.615 23.65 2.81 ;
      RECT 24.93 2.687 24.94 2.885 ;
      RECT 24.73 2.687 24.74 2.885 ;
      RECT 24.715 2.702 24.73 2.875 ;
      RECT 24.71 2.71 24.715 2.868 ;
      RECT 24.7 2.713 24.71 2.865 ;
      RECT 24.665 2.712 24.7 2.863 ;
      RECT 24.636 2.708 24.665 2.86 ;
      RECT 24.55 2.703 24.636 2.857 ;
      RECT 24.49 2.697 24.55 2.853 ;
      RECT 24.461 2.693 24.49 2.85 ;
      RECT 24.375 2.685 24.461 2.847 ;
      RECT 24.366 2.679 24.375 2.845 ;
      RECT 24.28 2.674 24.366 2.843 ;
      RECT 24.257 2.669 24.28 2.84 ;
      RECT 24.171 2.663 24.257 2.837 ;
      RECT 24.085 2.654 24.171 2.832 ;
      RECT 24.075 2.649 24.085 2.83 ;
      RECT 24.056 2.648 24.075 2.829 ;
      RECT 23.97 2.643 24.056 2.825 ;
      RECT 23.95 2.638 23.97 2.821 ;
      RECT 23.89 2.633 23.95 2.818 ;
      RECT 23.865 2.623 23.89 2.816 ;
      RECT 23.86 2.616 23.865 2.815 ;
      RECT 23.85 2.607 23.86 2.814 ;
      RECT 23.846 2.6 23.85 2.814 ;
      RECT 23.76 2.6 23.846 2.812 ;
      RECT 23.65 2.607 23.665 2.81 ;
      RECT 23.635 2.617 23.64 2.81 ;
      RECT 23.615 2.62 23.635 2.807 ;
      RECT 23.585 2.62 23.615 2.803 ;
      RECT 23.575 2.62 23.585 2.803 ;
      RECT 24.49 3.115 24.75 3.375 ;
      RECT 24.42 3.125 24.75 3.335 ;
      RECT 24.41 3.132 24.75 3.33 ;
      RECT 23.83 3.12 24.09 3.38 ;
      RECT 23.83 3.16 24.195 3.37 ;
      RECT 23.83 3.162 24.2 3.369 ;
      RECT 23.83 3.17 24.205 3.366 ;
      RECT 22.755 2.245 22.855 3.77 ;
      RECT 22.945 3.385 22.995 3.645 ;
      RECT 22.94 2.258 22.945 2.445 ;
      RECT 22.935 3.366 22.945 3.645 ;
      RECT 22.935 2.255 22.94 2.453 ;
      RECT 22.92 2.249 22.935 2.46 ;
      RECT 22.93 3.354 22.935 3.728 ;
      RECT 22.92 3.342 22.93 3.765 ;
      RECT 22.91 2.245 22.92 2.467 ;
      RECT 22.91 3.327 22.92 3.77 ;
      RECT 22.905 2.245 22.91 2.475 ;
      RECT 22.885 3.297 22.91 3.77 ;
      RECT 22.865 2.245 22.905 2.523 ;
      RECT 22.875 3.257 22.885 3.77 ;
      RECT 22.865 3.212 22.875 3.77 ;
      RECT 22.86 2.245 22.865 2.593 ;
      RECT 22.86 3.17 22.865 3.77 ;
      RECT 22.855 2.245 22.86 3.07 ;
      RECT 22.855 3.152 22.86 3.77 ;
      RECT 22.745 2.248 22.755 3.77 ;
      RECT 22.73 2.255 22.745 3.766 ;
      RECT 22.725 2.265 22.73 3.761 ;
      RECT 22.72 2.465 22.725 3.653 ;
      RECT 22.715 2.55 22.72 3.205 ;
      RECT 21.59 7.77 21.88 8 ;
      RECT 21.65 6.29 21.82 8 ;
      RECT 21.645 6.655 21.995 7.005 ;
      RECT 21.59 6.29 21.88 6.52 ;
      RECT 21.185 2.395 21.29 2.965 ;
      RECT 21.185 2.73 21.51 2.96 ;
      RECT 21.185 2.76 21.68 2.93 ;
      RECT 21.185 2.395 21.375 2.96 ;
      RECT 20.6 2.36 20.89 2.59 ;
      RECT 20.6 2.395 21.375 2.565 ;
      RECT 20.66 0.88 20.83 2.59 ;
      RECT 20.6 0.88 20.89 1.11 ;
      RECT 20.6 7.77 20.89 8 ;
      RECT 20.66 6.29 20.83 8 ;
      RECT 20.6 6.29 20.89 6.52 ;
      RECT 20.6 6.325 21.455 6.485 ;
      RECT 21.285 5.92 21.455 6.485 ;
      RECT 20.6 6.32 20.995 6.485 ;
      RECT 21.22 5.92 21.51 6.15 ;
      RECT 21.22 5.95 21.68 6.12 ;
      RECT 20.23 2.73 20.52 2.96 ;
      RECT 20.23 2.76 20.69 2.93 ;
      RECT 20.295 1.655 20.46 2.96 ;
      RECT 18.81 1.625 19.1 1.855 ;
      RECT 18.81 1.655 20.46 1.825 ;
      RECT 18.87 0.885 19.04 1.855 ;
      RECT 18.81 0.885 19.1 1.115 ;
      RECT 18.81 7.765 19.1 7.995 ;
      RECT 18.87 7.025 19.04 7.995 ;
      RECT 18.87 7.12 20.46 7.29 ;
      RECT 20.29 5.92 20.46 7.29 ;
      RECT 18.81 7.025 19.1 7.255 ;
      RECT 20.23 5.92 20.52 6.15 ;
      RECT 20.23 5.95 20.69 6.12 ;
      RECT 16.845 3.43 17.195 3.78 ;
      RECT 16.935 2.025 17.105 3.78 ;
      RECT 19.24 1.965 19.59 2.315 ;
      RECT 16.935 2.025 18.555 2.2 ;
      RECT 16.935 2.025 19.59 2.195 ;
      RECT 19.265 6.655 19.59 6.98 ;
      RECT 14.66 6.605 15.01 6.955 ;
      RECT 19.24 6.655 19.59 6.885 ;
      RECT 14.48 6.655 15.01 6.885 ;
      RECT 14.31 6.685 19.59 6.855 ;
      RECT 18.465 2.365 18.785 2.685 ;
      RECT 18.435 2.365 18.785 2.595 ;
      RECT 18.265 2.395 18.785 2.565 ;
      RECT 18.465 6.225 18.785 6.545 ;
      RECT 18.435 6.285 18.785 6.515 ;
      RECT 18.265 6.315 18.785 6.485 ;
      RECT 14.245 3.665 14.285 3.925 ;
      RECT 14.285 3.645 14.29 3.655 ;
      RECT 15.615 2.89 15.625 3.111 ;
      RECT 15.545 2.885 15.615 3.236 ;
      RECT 15.535 2.885 15.545 3.363 ;
      RECT 15.51 2.885 15.535 3.41 ;
      RECT 15.485 2.885 15.51 3.488 ;
      RECT 15.465 2.885 15.485 3.558 ;
      RECT 15.44 2.885 15.465 3.598 ;
      RECT 15.43 2.885 15.44 3.618 ;
      RECT 15.42 2.887 15.43 3.626 ;
      RECT 15.415 2.892 15.42 3.083 ;
      RECT 15.415 3.092 15.42 3.627 ;
      RECT 15.41 3.137 15.415 3.628 ;
      RECT 15.4 3.202 15.41 3.629 ;
      RECT 15.39 3.297 15.4 3.631 ;
      RECT 15.385 3.35 15.39 3.633 ;
      RECT 15.38 3.37 15.385 3.634 ;
      RECT 15.325 3.395 15.38 3.64 ;
      RECT 15.285 3.43 15.325 3.649 ;
      RECT 15.275 3.447 15.285 3.654 ;
      RECT 15.266 3.453 15.275 3.656 ;
      RECT 15.18 3.491 15.266 3.667 ;
      RECT 15.175 3.53 15.18 3.677 ;
      RECT 15.1 3.537 15.175 3.687 ;
      RECT 15.08 3.547 15.1 3.698 ;
      RECT 15.05 3.554 15.08 3.706 ;
      RECT 15.025 3.561 15.05 3.713 ;
      RECT 15.001 3.567 15.025 3.718 ;
      RECT 14.915 3.58 15.001 3.73 ;
      RECT 14.837 3.587 14.915 3.748 ;
      RECT 14.751 3.582 14.837 3.766 ;
      RECT 14.665 3.577 14.751 3.786 ;
      RECT 14.585 3.571 14.665 3.803 ;
      RECT 14.52 3.567 14.585 3.832 ;
      RECT 14.515 3.281 14.52 3.305 ;
      RECT 14.505 3.557 14.52 3.86 ;
      RECT 14.51 3.275 14.515 3.345 ;
      RECT 14.505 3.269 14.51 3.415 ;
      RECT 14.5 3.263 14.505 3.493 ;
      RECT 14.5 3.54 14.505 3.925 ;
      RECT 14.492 3.26 14.5 3.925 ;
      RECT 14.406 3.258 14.492 3.925 ;
      RECT 14.32 3.256 14.406 3.925 ;
      RECT 14.31 3.257 14.32 3.925 ;
      RECT 14.305 3.262 14.31 3.925 ;
      RECT 14.295 3.275 14.305 3.925 ;
      RECT 14.29 3.297 14.295 3.925 ;
      RECT 14.285 3.657 14.29 3.925 ;
      RECT 14.915 3.125 14.92 3.345 ;
      RECT 15.42 2.16 15.455 2.42 ;
      RECT 15.405 2.16 15.42 2.428 ;
      RECT 15.376 2.16 15.405 2.45 ;
      RECT 15.29 2.16 15.376 2.51 ;
      RECT 15.27 2.16 15.29 2.575 ;
      RECT 15.21 2.16 15.27 2.74 ;
      RECT 15.205 2.16 15.21 2.888 ;
      RECT 15.2 2.16 15.205 2.9 ;
      RECT 15.195 2.16 15.2 2.926 ;
      RECT 15.165 2.346 15.195 3.006 ;
      RECT 15.16 2.394 15.165 3.095 ;
      RECT 15.155 2.408 15.16 3.11 ;
      RECT 15.15 2.427 15.155 3.14 ;
      RECT 15.145 2.442 15.15 3.156 ;
      RECT 15.14 2.457 15.145 3.178 ;
      RECT 15.135 2.477 15.14 3.2 ;
      RECT 15.125 2.497 15.135 3.233 ;
      RECT 15.11 2.539 15.125 3.295 ;
      RECT 15.105 2.57 15.11 3.335 ;
      RECT 15.1 2.582 15.105 3.34 ;
      RECT 15.095 2.594 15.1 3.345 ;
      RECT 15.09 2.607 15.095 3.345 ;
      RECT 15.085 2.625 15.09 3.345 ;
      RECT 15.08 2.645 15.085 3.345 ;
      RECT 15.075 2.657 15.08 3.345 ;
      RECT 15.07 2.67 15.075 3.345 ;
      RECT 15.05 2.705 15.07 3.345 ;
      RECT 15 2.807 15.05 3.345 ;
      RECT 14.995 2.892 15 3.345 ;
      RECT 14.99 2.9 14.995 3.345 ;
      RECT 14.985 2.917 14.99 3.345 ;
      RECT 14.98 2.932 14.985 3.345 ;
      RECT 14.945 2.997 14.98 3.345 ;
      RECT 14.93 3.062 14.945 3.345 ;
      RECT 14.925 3.092 14.93 3.345 ;
      RECT 14.92 3.117 14.925 3.345 ;
      RECT 14.905 3.127 14.915 3.345 ;
      RECT 14.89 3.14 14.905 3.338 ;
      RECT 14.635 2.73 14.705 2.94 ;
      RECT 14.425 2.707 14.43 2.9 ;
      RECT 11.88 2.635 12.14 2.895 ;
      RECT 14.715 2.917 14.72 2.92 ;
      RECT 14.705 2.735 14.715 2.935 ;
      RECT 14.606 2.728 14.635 2.94 ;
      RECT 14.52 2.72 14.606 2.94 ;
      RECT 14.505 2.714 14.52 2.938 ;
      RECT 14.485 2.713 14.505 2.925 ;
      RECT 14.48 2.712 14.485 2.908 ;
      RECT 14.43 2.709 14.48 2.903 ;
      RECT 14.4 2.706 14.425 2.898 ;
      RECT 14.38 2.704 14.4 2.893 ;
      RECT 14.365 2.702 14.38 2.89 ;
      RECT 14.335 2.7 14.365 2.888 ;
      RECT 14.27 2.696 14.335 2.88 ;
      RECT 14.24 2.691 14.27 2.875 ;
      RECT 14.22 2.689 14.24 2.873 ;
      RECT 14.19 2.686 14.22 2.868 ;
      RECT 14.13 2.682 14.19 2.86 ;
      RECT 14.125 2.679 14.13 2.855 ;
      RECT 14.055 2.677 14.125 2.85 ;
      RECT 14.026 2.673 14.055 2.843 ;
      RECT 13.94 2.668 14.026 2.835 ;
      RECT 13.906 2.663 13.94 2.827 ;
      RECT 13.82 2.655 13.906 2.819 ;
      RECT 13.781 2.648 13.82 2.811 ;
      RECT 13.695 2.643 13.781 2.803 ;
      RECT 13.63 2.637 13.695 2.793 ;
      RECT 13.61 2.632 13.63 2.788 ;
      RECT 13.601 2.629 13.61 2.787 ;
      RECT 13.515 2.625 13.601 2.781 ;
      RECT 13.475 2.621 13.515 2.773 ;
      RECT 13.455 2.617 13.475 2.771 ;
      RECT 13.395 2.617 13.455 2.768 ;
      RECT 13.375 2.62 13.395 2.766 ;
      RECT 13.354 2.62 13.375 2.766 ;
      RECT 13.268 2.622 13.354 2.77 ;
      RECT 13.182 2.624 13.268 2.776 ;
      RECT 13.096 2.626 13.182 2.783 ;
      RECT 13.01 2.629 13.096 2.789 ;
      RECT 12.976 2.63 13.01 2.794 ;
      RECT 12.89 2.633 12.976 2.799 ;
      RECT 12.861 2.64 12.89 2.804 ;
      RECT 12.775 2.64 12.861 2.809 ;
      RECT 12.742 2.64 12.775 2.814 ;
      RECT 12.656 2.642 12.742 2.819 ;
      RECT 12.57 2.644 12.656 2.826 ;
      RECT 12.506 2.646 12.57 2.832 ;
      RECT 12.42 2.648 12.506 2.838 ;
      RECT 12.417 2.65 12.42 2.841 ;
      RECT 12.331 2.651 12.417 2.845 ;
      RECT 12.245 2.654 12.331 2.852 ;
      RECT 12.226 2.656 12.245 2.856 ;
      RECT 12.14 2.658 12.226 2.861 ;
      RECT 11.87 2.67 11.88 2.865 ;
      RECT 14.05 7.765 14.34 7.995 ;
      RECT 14.11 7.025 14.28 7.995 ;
      RECT 14 7.055 14.375 7.425 ;
      RECT 14.05 7.025 14.34 7.425 ;
      RECT 14.105 2.25 14.29 2.46 ;
      RECT 14.1 2.251 14.295 2.458 ;
      RECT 14.095 2.256 14.305 2.453 ;
      RECT 14.09 2.232 14.095 2.45 ;
      RECT 14.06 2.229 14.09 2.443 ;
      RECT 14.055 2.225 14.06 2.434 ;
      RECT 14.02 2.256 14.305 2.429 ;
      RECT 13.795 2.165 14.055 2.425 ;
      RECT 14.095 2.234 14.1 2.453 ;
      RECT 14.1 2.235 14.105 2.458 ;
      RECT 13.795 2.247 14.175 2.425 ;
      RECT 13.795 2.245 14.16 2.425 ;
      RECT 13.795 2.24 14.15 2.425 ;
      RECT 13.75 3.155 13.8 3.44 ;
      RECT 13.695 3.125 13.7 3.44 ;
      RECT 13.665 3.105 13.67 3.44 ;
      RECT 13.815 3.155 13.875 3.415 ;
      RECT 13.81 3.155 13.815 3.423 ;
      RECT 13.8 3.155 13.81 3.435 ;
      RECT 13.715 3.145 13.75 3.44 ;
      RECT 13.71 3.132 13.715 3.44 ;
      RECT 13.7 3.127 13.71 3.44 ;
      RECT 13.68 3.117 13.695 3.44 ;
      RECT 13.67 3.11 13.68 3.44 ;
      RECT 13.66 3.102 13.665 3.44 ;
      RECT 13.63 3.092 13.66 3.44 ;
      RECT 13.615 3.08 13.63 3.44 ;
      RECT 13.6 3.07 13.615 3.435 ;
      RECT 13.58 3.06 13.6 3.41 ;
      RECT 13.57 3.052 13.58 3.387 ;
      RECT 13.54 3.035 13.57 3.377 ;
      RECT 13.535 3.012 13.54 3.368 ;
      RECT 13.53 2.999 13.535 3.366 ;
      RECT 13.515 2.975 13.53 3.36 ;
      RECT 13.51 2.951 13.515 3.354 ;
      RECT 13.5 2.94 13.51 3.349 ;
      RECT 13.495 2.93 13.5 3.345 ;
      RECT 13.49 2.922 13.495 3.342 ;
      RECT 13.48 2.917 13.49 3.338 ;
      RECT 13.475 2.912 13.48 3.334 ;
      RECT 13.39 2.91 13.475 3.309 ;
      RECT 13.36 2.91 13.39 3.275 ;
      RECT 13.345 2.91 13.36 3.258 ;
      RECT 13.29 2.91 13.345 3.203 ;
      RECT 13.285 2.915 13.29 3.152 ;
      RECT 13.275 2.92 13.285 3.142 ;
      RECT 13.27 2.93 13.275 3.128 ;
      RECT 13.22 3.67 13.48 3.93 ;
      RECT 13.14 3.685 13.48 3.906 ;
      RECT 13.12 3.685 13.48 3.901 ;
      RECT 13.096 3.685 13.48 3.899 ;
      RECT 13.01 3.685 13.48 3.894 ;
      RECT 12.86 3.625 13.12 3.89 ;
      RECT 12.815 3.685 13.48 3.885 ;
      RECT 12.81 3.692 13.48 3.88 ;
      RECT 12.825 3.68 13.14 3.89 ;
      RECT 12.715 2.115 12.975 2.375 ;
      RECT 12.715 2.172 12.98 2.368 ;
      RECT 12.715 2.202 12.985 2.3 ;
      RECT 12.775 2.633 12.89 2.635 ;
      RECT 12.861 2.63 12.89 2.635 ;
      RECT 11.885 3.634 11.91 3.874 ;
      RECT 11.87 3.637 11.96 3.868 ;
      RECT 11.865 3.642 12.046 3.863 ;
      RECT 11.86 3.65 12.11 3.861 ;
      RECT 11.86 3.65 12.12 3.86 ;
      RECT 11.855 3.657 12.13 3.853 ;
      RECT 11.855 3.657 12.216 3.842 ;
      RECT 11.85 3.692 12.216 3.838 ;
      RECT 11.85 3.692 12.225 3.827 ;
      RECT 12.13 3.565 12.39 3.825 ;
      RECT 11.84 3.742 12.39 3.823 ;
      RECT 12.11 3.61 12.13 3.858 ;
      RECT 12.046 3.613 12.11 3.862 ;
      RECT 11.96 3.618 12.046 3.867 ;
      RECT 11.89 3.629 12.39 3.825 ;
      RECT 11.91 3.623 11.96 3.872 ;
      RECT 12.035 2.1 12.045 2.362 ;
      RECT 12.025 2.157 12.035 2.365 ;
      RECT 12 2.162 12.025 2.371 ;
      RECT 11.975 2.166 12 2.383 ;
      RECT 11.965 2.169 11.975 2.393 ;
      RECT 11.96 2.17 11.965 2.398 ;
      RECT 11.955 2.171 11.96 2.403 ;
      RECT 11.95 2.172 11.955 2.405 ;
      RECT 11.925 2.175 11.95 2.408 ;
      RECT 11.895 2.181 11.925 2.411 ;
      RECT 11.83 2.192 11.895 2.414 ;
      RECT 11.785 2.2 11.83 2.418 ;
      RECT 11.77 2.2 11.785 2.426 ;
      RECT 11.765 2.201 11.77 2.433 ;
      RECT 11.76 2.203 11.765 2.436 ;
      RECT 11.755 2.207 11.76 2.439 ;
      RECT 11.745 2.215 11.755 2.443 ;
      RECT 11.74 2.228 11.745 2.448 ;
      RECT 11.735 2.236 11.74 2.45 ;
      RECT 11.73 2.242 11.735 2.45 ;
      RECT 11.725 2.246 11.73 2.453 ;
      RECT 11.72 2.248 11.725 2.456 ;
      RECT 11.715 2.251 11.72 2.459 ;
      RECT 11.705 2.256 11.715 2.463 ;
      RECT 11.7 2.262 11.705 2.468 ;
      RECT 11.69 2.268 11.7 2.472 ;
      RECT 11.675 2.275 11.69 2.478 ;
      RECT 11.646 2.289 11.675 2.488 ;
      RECT 11.56 2.324 11.646 2.52 ;
      RECT 11.54 2.357 11.56 2.549 ;
      RECT 11.52 2.37 11.54 2.56 ;
      RECT 11.5 2.382 11.52 2.571 ;
      RECT 11.45 2.404 11.5 2.591 ;
      RECT 11.435 2.422 11.45 2.608 ;
      RECT 11.43 2.428 11.435 2.611 ;
      RECT 11.425 2.432 11.43 2.614 ;
      RECT 11.42 2.436 11.425 2.618 ;
      RECT 11.415 2.438 11.42 2.621 ;
      RECT 11.405 2.445 11.415 2.624 ;
      RECT 11.4 2.45 11.405 2.628 ;
      RECT 11.395 2.452 11.4 2.631 ;
      RECT 11.39 2.456 11.395 2.634 ;
      RECT 11.385 2.458 11.39 2.638 ;
      RECT 11.37 2.463 11.385 2.643 ;
      RECT 11.365 2.468 11.37 2.646 ;
      RECT 11.36 2.476 11.365 2.649 ;
      RECT 11.355 2.478 11.36 2.652 ;
      RECT 11.35 2.48 11.355 2.655 ;
      RECT 11.34 2.482 11.35 2.661 ;
      RECT 11.305 2.496 11.34 2.673 ;
      RECT 11.295 2.511 11.305 2.683 ;
      RECT 11.22 2.54 11.295 2.707 ;
      RECT 11.215 2.565 11.22 2.73 ;
      RECT 11.2 2.569 11.215 2.736 ;
      RECT 11.19 2.577 11.2 2.741 ;
      RECT 11.16 2.59 11.19 2.745 ;
      RECT 11.15 2.605 11.16 2.75 ;
      RECT 11.14 2.61 11.15 2.753 ;
      RECT 11.135 2.612 11.14 2.755 ;
      RECT 11.12 2.615 11.135 2.758 ;
      RECT 11.115 2.617 11.12 2.761 ;
      RECT 11.095 2.622 11.115 2.765 ;
      RECT 11.065 2.627 11.095 2.773 ;
      RECT 11.04 2.634 11.065 2.781 ;
      RECT 11.035 2.639 11.04 2.786 ;
      RECT 11.005 2.642 11.035 2.79 ;
      RECT 10.965 2.645 11.005 2.8 ;
      RECT 10.93 2.642 10.965 2.812 ;
      RECT 10.92 2.638 10.93 2.819 ;
      RECT 10.895 2.634 10.92 2.825 ;
      RECT 10.89 2.63 10.895 2.83 ;
      RECT 10.85 2.627 10.89 2.83 ;
      RECT 10.835 2.612 10.85 2.831 ;
      RECT 10.812 2.6 10.835 2.831 ;
      RECT 10.726 2.6 10.812 2.832 ;
      RECT 10.64 2.6 10.726 2.834 ;
      RECT 10.62 2.6 10.64 2.831 ;
      RECT 10.615 2.605 10.62 2.826 ;
      RECT 10.61 2.61 10.615 2.824 ;
      RECT 10.6 2.62 10.61 2.822 ;
      RECT 10.595 2.626 10.6 2.815 ;
      RECT 10.59 2.628 10.595 2.8 ;
      RECT 10.585 2.632 10.59 2.79 ;
      RECT 12.045 2.1 12.295 2.36 ;
      RECT 9.77 3.635 10.03 3.895 ;
      RECT 12.065 3.125 12.07 3.335 ;
      RECT 12.07 3.13 12.08 3.33 ;
      RECT 12.02 3.125 12.065 3.35 ;
      RECT 12.01 3.125 12.02 3.37 ;
      RECT 11.991 3.125 12.01 3.375 ;
      RECT 11.905 3.125 11.991 3.372 ;
      RECT 11.875 3.127 11.905 3.37 ;
      RECT 11.82 3.137 11.875 3.368 ;
      RECT 11.755 3.151 11.82 3.366 ;
      RECT 11.75 3.159 11.755 3.365 ;
      RECT 11.735 3.162 11.75 3.363 ;
      RECT 11.67 3.172 11.735 3.359 ;
      RECT 11.622 3.186 11.67 3.36 ;
      RECT 11.536 3.203 11.622 3.374 ;
      RECT 11.45 3.224 11.536 3.391 ;
      RECT 11.43 3.237 11.45 3.401 ;
      RECT 11.385 3.245 11.43 3.408 ;
      RECT 11.35 3.253 11.385 3.416 ;
      RECT 11.316 3.261 11.35 3.424 ;
      RECT 11.23 3.275 11.316 3.436 ;
      RECT 11.195 3.292 11.23 3.448 ;
      RECT 11.186 3.301 11.195 3.452 ;
      RECT 11.1 3.319 11.186 3.469 ;
      RECT 11.041 3.346 11.1 3.496 ;
      RECT 10.955 3.373 11.041 3.524 ;
      RECT 10.935 3.395 10.955 3.544 ;
      RECT 10.875 3.41 10.935 3.56 ;
      RECT 10.865 3.422 10.875 3.573 ;
      RECT 10.86 3.427 10.865 3.576 ;
      RECT 10.85 3.43 10.86 3.579 ;
      RECT 10.845 3.432 10.85 3.582 ;
      RECT 10.815 3.44 10.845 3.589 ;
      RECT 10.8 3.447 10.815 3.597 ;
      RECT 10.79 3.452 10.8 3.601 ;
      RECT 10.785 3.455 10.79 3.604 ;
      RECT 10.775 3.457 10.785 3.607 ;
      RECT 10.74 3.467 10.775 3.616 ;
      RECT 10.665 3.49 10.74 3.638 ;
      RECT 10.645 3.508 10.665 3.656 ;
      RECT 10.615 3.515 10.645 3.666 ;
      RECT 10.595 3.523 10.615 3.676 ;
      RECT 10.585 3.529 10.595 3.683 ;
      RECT 10.566 3.534 10.585 3.689 ;
      RECT 10.48 3.554 10.566 3.709 ;
      RECT 10.465 3.574 10.48 3.728 ;
      RECT 10.42 3.586 10.465 3.739 ;
      RECT 10.355 3.607 10.42 3.762 ;
      RECT 10.315 3.627 10.355 3.783 ;
      RECT 10.305 3.637 10.315 3.793 ;
      RECT 10.255 3.649 10.305 3.804 ;
      RECT 10.235 3.665 10.255 3.816 ;
      RECT 10.205 3.675 10.235 3.822 ;
      RECT 10.195 3.68 10.205 3.824 ;
      RECT 10.126 3.681 10.195 3.83 ;
      RECT 10.04 3.683 10.126 3.84 ;
      RECT 10.03 3.684 10.04 3.845 ;
      RECT 11.3 3.71 11.49 3.92 ;
      RECT 11.29 3.715 11.5 3.913 ;
      RECT 11.275 3.715 11.5 3.878 ;
      RECT 11.195 3.6 11.455 3.86 ;
      RECT 10.11 3.13 10.295 3.425 ;
      RECT 10.1 3.13 10.295 3.423 ;
      RECT 10.085 3.13 10.3 3.418 ;
      RECT 10.085 3.13 10.305 3.415 ;
      RECT 10.08 3.13 10.305 3.413 ;
      RECT 10.075 3.385 10.305 3.403 ;
      RECT 10.08 3.13 10.34 3.39 ;
      RECT 10.04 2.165 10.3 2.425 ;
      RECT 9.85 2.09 9.936 2.423 ;
      RECT 9.825 2.094 9.98 2.419 ;
      RECT 9.936 2.086 9.98 2.419 ;
      RECT 9.936 2.087 9.985 2.418 ;
      RECT 9.85 2.092 10 2.417 ;
      RECT 9.825 2.1 10.04 2.416 ;
      RECT 9.82 2.095 10 2.411 ;
      RECT 9.81 2.11 10.04 2.318 ;
      RECT 9.81 2.162 10.24 2.318 ;
      RECT 9.81 2.155 10.22 2.318 ;
      RECT 9.81 2.142 10.19 2.318 ;
      RECT 9.81 2.13 10.13 2.318 ;
      RECT 9.81 2.115 10.105 2.318 ;
      RECT 9.01 2.745 9.145 3.04 ;
      RECT 9.27 2.768 9.275 2.955 ;
      RECT 9.99 2.665 10.135 2.9 ;
      RECT 10.15 2.665 10.155 2.89 ;
      RECT 10.185 2.676 10.19 2.87 ;
      RECT 10.18 2.668 10.185 2.875 ;
      RECT 10.16 2.665 10.18 2.88 ;
      RECT 10.155 2.665 10.16 2.888 ;
      RECT 10.145 2.665 10.15 2.893 ;
      RECT 10.135 2.665 10.145 2.898 ;
      RECT 9.965 2.667 9.99 2.9 ;
      RECT 9.915 2.674 9.965 2.9 ;
      RECT 9.91 2.679 9.915 2.9 ;
      RECT 9.871 2.684 9.91 2.901 ;
      RECT 9.785 2.696 9.871 2.902 ;
      RECT 9.776 2.706 9.785 2.902 ;
      RECT 9.69 2.715 9.776 2.904 ;
      RECT 9.666 2.725 9.69 2.906 ;
      RECT 9.58 2.736 9.666 2.907 ;
      RECT 9.55 2.747 9.58 2.909 ;
      RECT 9.52 2.752 9.55 2.911 ;
      RECT 9.495 2.758 9.52 2.914 ;
      RECT 9.48 2.763 9.495 2.915 ;
      RECT 9.435 2.769 9.48 2.915 ;
      RECT 9.43 2.774 9.435 2.916 ;
      RECT 9.41 2.774 9.43 2.918 ;
      RECT 9.39 2.772 9.41 2.923 ;
      RECT 9.355 2.771 9.39 2.93 ;
      RECT 9.325 2.77 9.355 2.94 ;
      RECT 9.275 2.769 9.325 2.95 ;
      RECT 9.185 2.766 9.27 3.04 ;
      RECT 9.16 2.76 9.185 3.04 ;
      RECT 9.145 2.75 9.16 3.04 ;
      RECT 8.96 2.745 9.01 2.96 ;
      RECT 8.95 2.75 8.96 2.95 ;
      RECT 9.19 3.225 9.45 3.485 ;
      RECT 9.19 3.225 9.48 3.378 ;
      RECT 9.19 3.225 9.515 3.363 ;
      RECT 9.445 3.145 9.635 3.355 ;
      RECT 9.435 3.15 9.645 3.348 ;
      RECT 9.4 3.22 9.645 3.348 ;
      RECT 9.43 3.162 9.45 3.485 ;
      RECT 9.415 3.21 9.645 3.348 ;
      RECT 9.42 3.182 9.45 3.485 ;
      RECT 8.5 2.25 8.57 3.355 ;
      RECT 9.235 2.355 9.495 2.615 ;
      RECT 8.815 2.401 8.83 2.61 ;
      RECT 9.151 2.414 9.235 2.565 ;
      RECT 9.065 2.411 9.151 2.565 ;
      RECT 9.026 2.409 9.065 2.565 ;
      RECT 8.94 2.407 9.026 2.565 ;
      RECT 8.88 2.405 8.94 2.576 ;
      RECT 8.845 2.403 8.88 2.594 ;
      RECT 8.83 2.401 8.845 2.605 ;
      RECT 8.8 2.401 8.815 2.618 ;
      RECT 8.79 2.401 8.8 2.623 ;
      RECT 8.765 2.4 8.79 2.628 ;
      RECT 8.75 2.395 8.765 2.634 ;
      RECT 8.745 2.388 8.75 2.639 ;
      RECT 8.72 2.379 8.745 2.645 ;
      RECT 8.675 2.358 8.72 2.658 ;
      RECT 8.665 2.342 8.675 2.668 ;
      RECT 8.65 2.335 8.665 2.678 ;
      RECT 8.64 2.328 8.65 2.695 ;
      RECT 8.635 2.325 8.64 2.725 ;
      RECT 8.63 2.323 8.635 2.755 ;
      RECT 8.625 2.321 8.63 2.792 ;
      RECT 8.61 2.317 8.625 2.859 ;
      RECT 8.61 3.15 8.62 3.35 ;
      RECT 8.605 2.313 8.61 2.985 ;
      RECT 8.605 3.137 8.61 3.355 ;
      RECT 8.6 2.311 8.605 3.07 ;
      RECT 8.6 3.127 8.605 3.355 ;
      RECT 8.585 2.282 8.6 3.355 ;
      RECT 8.57 2.255 8.585 3.355 ;
      RECT 8.495 2.25 8.5 2.605 ;
      RECT 8.495 2.66 8.5 3.355 ;
      RECT 8.48 2.25 8.495 2.583 ;
      RECT 8.49 2.682 8.495 3.355 ;
      RECT 8.48 2.722 8.49 3.355 ;
      RECT 8.445 2.25 8.48 2.525 ;
      RECT 8.475 2.757 8.48 3.355 ;
      RECT 8.46 2.812 8.475 3.355 ;
      RECT 8.455 2.877 8.46 3.355 ;
      RECT 8.44 2.925 8.455 3.355 ;
      RECT 8.415 2.25 8.445 2.48 ;
      RECT 8.435 2.98 8.44 3.355 ;
      RECT 8.42 3.04 8.435 3.355 ;
      RECT 8.415 3.088 8.42 3.353 ;
      RECT 8.41 2.25 8.415 2.473 ;
      RECT 8.41 3.12 8.415 3.348 ;
      RECT 8.385 2.25 8.41 2.465 ;
      RECT 8.375 2.255 8.385 2.455 ;
      RECT 8.59 3.53 8.61 3.77 ;
      RECT 7.82 3.46 7.825 3.67 ;
      RECT 9.1 3.533 9.11 3.728 ;
      RECT 9.095 3.523 9.1 3.731 ;
      RECT 9.015 3.52 9.095 3.754 ;
      RECT 9.011 3.52 9.015 3.776 ;
      RECT 8.925 3.52 9.011 3.786 ;
      RECT 8.91 3.52 8.925 3.794 ;
      RECT 8.881 3.521 8.91 3.792 ;
      RECT 8.795 3.526 8.881 3.788 ;
      RECT 8.782 3.53 8.795 3.784 ;
      RECT 8.696 3.53 8.782 3.78 ;
      RECT 8.61 3.53 8.696 3.774 ;
      RECT 8.526 3.53 8.59 3.768 ;
      RECT 8.44 3.53 8.526 3.763 ;
      RECT 8.42 3.53 8.44 3.759 ;
      RECT 8.36 3.525 8.42 3.756 ;
      RECT 8.332 3.519 8.36 3.753 ;
      RECT 8.246 3.514 8.332 3.749 ;
      RECT 8.16 3.508 8.246 3.743 ;
      RECT 8.085 3.49 8.16 3.738 ;
      RECT 8.05 3.467 8.085 3.734 ;
      RECT 8.04 3.457 8.05 3.733 ;
      RECT 7.985 3.455 8.04 3.732 ;
      RECT 7.91 3.455 7.985 3.728 ;
      RECT 7.9 3.455 7.91 3.723 ;
      RECT 7.885 3.455 7.9 3.715 ;
      RECT 7.835 3.457 7.885 3.693 ;
      RECT 7.825 3.46 7.835 3.673 ;
      RECT 7.815 3.465 7.82 3.668 ;
      RECT 7.81 3.47 7.815 3.663 ;
      RECT 7.935 2.635 8.195 2.895 ;
      RECT 7.935 2.65 8.215 2.86 ;
      RECT 7.935 2.655 8.225 2.855 ;
      RECT 5.92 2.115 6.18 2.375 ;
      RECT 5.91 2.145 6.18 2.355 ;
      RECT 7.83 2.06 8.09 2.32 ;
      RECT 7.825 2.135 7.83 2.321 ;
      RECT 7.8 2.14 7.825 2.323 ;
      RECT 7.785 2.147 7.8 2.326 ;
      RECT 7.725 2.165 7.785 2.331 ;
      RECT 7.695 2.185 7.725 2.338 ;
      RECT 7.67 2.193 7.695 2.343 ;
      RECT 7.645 2.201 7.67 2.345 ;
      RECT 7.627 2.205 7.645 2.344 ;
      RECT 7.541 2.203 7.627 2.344 ;
      RECT 7.455 2.201 7.541 2.344 ;
      RECT 7.369 2.199 7.455 2.343 ;
      RECT 7.283 2.197 7.369 2.343 ;
      RECT 7.197 2.195 7.283 2.343 ;
      RECT 7.111 2.193 7.197 2.343 ;
      RECT 7.025 2.191 7.111 2.342 ;
      RECT 7.007 2.19 7.025 2.342 ;
      RECT 6.921 2.189 7.007 2.342 ;
      RECT 6.835 2.187 6.921 2.342 ;
      RECT 6.749 2.186 6.835 2.341 ;
      RECT 6.663 2.185 6.749 2.341 ;
      RECT 6.577 2.183 6.663 2.341 ;
      RECT 6.491 2.182 6.577 2.341 ;
      RECT 6.405 2.18 6.491 2.34 ;
      RECT 6.381 2.178 6.405 2.34 ;
      RECT 6.295 2.171 6.381 2.34 ;
      RECT 6.266 2.163 6.295 2.34 ;
      RECT 6.18 2.155 6.266 2.34 ;
      RECT 5.9 2.152 5.91 2.35 ;
      RECT 7.405 3.115 7.41 3.465 ;
      RECT 7.175 3.205 7.315 3.465 ;
      RECT 7.65 2.89 7.695 3.1 ;
      RECT 7.705 2.901 7.715 3.095 ;
      RECT 7.695 2.893 7.705 3.1 ;
      RECT 7.63 2.89 7.65 3.105 ;
      RECT 7.6 2.89 7.63 3.128 ;
      RECT 7.59 2.89 7.6 3.153 ;
      RECT 7.585 2.89 7.59 3.163 ;
      RECT 7.53 2.89 7.585 3.203 ;
      RECT 7.525 2.89 7.53 3.243 ;
      RECT 7.52 2.892 7.525 3.248 ;
      RECT 7.505 2.902 7.52 3.259 ;
      RECT 7.46 2.96 7.505 3.295 ;
      RECT 7.45 3.015 7.46 3.329 ;
      RECT 7.435 3.042 7.45 3.345 ;
      RECT 7.425 3.069 7.435 3.465 ;
      RECT 7.41 3.092 7.425 3.465 ;
      RECT 7.4 3.132 7.405 3.465 ;
      RECT 7.395 3.142 7.4 3.465 ;
      RECT 7.39 3.157 7.395 3.465 ;
      RECT 7.38 3.162 7.39 3.465 ;
      RECT 7.315 3.185 7.38 3.465 ;
      RECT 6.815 2.68 7.005 2.89 ;
      RECT 5.39 2.605 5.65 2.865 ;
      RECT 5.74 2.6 5.835 2.81 ;
      RECT 5.715 2.615 5.725 2.81 ;
      RECT 7.005 2.687 7.015 2.885 ;
      RECT 6.805 2.687 6.815 2.885 ;
      RECT 6.79 2.702 6.805 2.875 ;
      RECT 6.785 2.71 6.79 2.868 ;
      RECT 6.775 2.713 6.785 2.865 ;
      RECT 6.74 2.712 6.775 2.863 ;
      RECT 6.711 2.708 6.74 2.86 ;
      RECT 6.625 2.703 6.711 2.857 ;
      RECT 6.565 2.697 6.625 2.853 ;
      RECT 6.536 2.693 6.565 2.85 ;
      RECT 6.45 2.685 6.536 2.847 ;
      RECT 6.441 2.679 6.45 2.845 ;
      RECT 6.355 2.674 6.441 2.843 ;
      RECT 6.332 2.669 6.355 2.84 ;
      RECT 6.246 2.663 6.332 2.837 ;
      RECT 6.16 2.654 6.246 2.832 ;
      RECT 6.15 2.649 6.16 2.83 ;
      RECT 6.131 2.648 6.15 2.829 ;
      RECT 6.045 2.643 6.131 2.825 ;
      RECT 6.025 2.638 6.045 2.821 ;
      RECT 5.965 2.633 6.025 2.818 ;
      RECT 5.94 2.623 5.965 2.816 ;
      RECT 5.935 2.616 5.94 2.815 ;
      RECT 5.925 2.607 5.935 2.814 ;
      RECT 5.921 2.6 5.925 2.814 ;
      RECT 5.835 2.6 5.921 2.812 ;
      RECT 5.725 2.607 5.74 2.81 ;
      RECT 5.71 2.617 5.715 2.81 ;
      RECT 5.69 2.62 5.71 2.807 ;
      RECT 5.66 2.62 5.69 2.803 ;
      RECT 5.65 2.62 5.66 2.803 ;
      RECT 6.565 3.115 6.825 3.375 ;
      RECT 6.495 3.125 6.825 3.335 ;
      RECT 6.485 3.132 6.825 3.33 ;
      RECT 5.905 3.12 6.165 3.38 ;
      RECT 5.905 3.16 6.27 3.37 ;
      RECT 5.905 3.162 6.275 3.369 ;
      RECT 5.905 3.17 6.28 3.366 ;
      RECT 4.83 2.245 4.93 3.77 ;
      RECT 5.02 3.385 5.07 3.645 ;
      RECT 5.015 2.258 5.02 2.445 ;
      RECT 5.01 3.366 5.02 3.645 ;
      RECT 5.01 2.255 5.015 2.453 ;
      RECT 4.995 2.249 5.01 2.46 ;
      RECT 5.005 3.354 5.01 3.728 ;
      RECT 4.995 3.342 5.005 3.765 ;
      RECT 4.985 2.245 4.995 2.467 ;
      RECT 4.985 3.327 4.995 3.77 ;
      RECT 4.98 2.245 4.985 2.475 ;
      RECT 4.96 3.297 4.985 3.77 ;
      RECT 4.94 2.245 4.98 2.523 ;
      RECT 4.95 3.257 4.96 3.77 ;
      RECT 4.94 3.212 4.95 3.77 ;
      RECT 4.935 2.245 4.94 2.593 ;
      RECT 4.935 3.17 4.94 3.77 ;
      RECT 4.93 2.245 4.935 3.07 ;
      RECT 4.93 3.152 4.935 3.77 ;
      RECT 4.82 2.248 4.83 3.77 ;
      RECT 4.805 2.255 4.82 3.766 ;
      RECT 4.8 2.265 4.805 3.761 ;
      RECT 4.795 2.465 4.8 3.653 ;
      RECT 4.79 2.55 4.795 3.205 ;
      RECT 3.02 7.765 3.31 7.995 ;
      RECT 3.08 7.025 3.25 7.995 ;
      RECT 2.99 7.025 3.34 7.315 ;
      RECT 2.615 6.285 2.965 6.575 ;
      RECT 2.475 6.315 2.965 6.485 ;
      RECT 88.52 1.14 88.895 1.51 ;
      RECT 82.5 2.225 82.76 2.485 ;
      RECT 70.595 1.14 70.97 1.51 ;
      RECT 64.575 2.225 64.835 2.485 ;
      RECT 52.67 1.14 53.045 1.51 ;
      RECT 46.65 2.225 46.91 2.485 ;
      RECT 34.745 1.14 35.12 1.51 ;
      RECT 28.725 2.225 28.985 2.485 ;
      RECT 16.82 1.14 17.195 1.51 ;
      RECT 10.8 2.225 11.06 2.485 ;
    LAYER mcon ;
      RECT 93.35 6.32 93.52 6.49 ;
      RECT 93.355 6.315 93.525 6.485 ;
      RECT 75.425 6.32 75.595 6.49 ;
      RECT 75.43 6.315 75.6 6.485 ;
      RECT 57.5 6.32 57.67 6.49 ;
      RECT 57.505 6.315 57.675 6.485 ;
      RECT 39.575 6.32 39.745 6.49 ;
      RECT 39.58 6.315 39.75 6.485 ;
      RECT 21.65 6.32 21.82 6.49 ;
      RECT 21.655 6.315 21.825 6.485 ;
      RECT 93.35 7.8 93.52 7.97 ;
      RECT 93 0.1 93.17 0.27 ;
      RECT 93 8.61 93.17 8.78 ;
      RECT 92.98 2.76 93.15 2.93 ;
      RECT 92.98 5.95 93.15 6.12 ;
      RECT 92.36 0.91 92.53 1.08 ;
      RECT 92.36 2.39 92.53 2.56 ;
      RECT 92.36 6.32 92.53 6.49 ;
      RECT 92.36 7.8 92.53 7.97 ;
      RECT 92.01 0.1 92.18 0.27 ;
      RECT 92.01 8.61 92.18 8.78 ;
      RECT 91.99 2.76 92.16 2.93 ;
      RECT 91.99 5.95 92.16 6.12 ;
      RECT 91.31 0.105 91.48 0.275 ;
      RECT 91.31 8.605 91.48 8.775 ;
      RECT 91 2.025 91.17 2.195 ;
      RECT 91 6.685 91.17 6.855 ;
      RECT 90.63 0.105 90.8 0.275 ;
      RECT 90.63 8.605 90.8 8.775 ;
      RECT 90.57 0.915 90.74 1.085 ;
      RECT 90.57 1.655 90.74 1.825 ;
      RECT 90.57 7.055 90.74 7.225 ;
      RECT 90.57 7.795 90.74 7.965 ;
      RECT 90.195 2.395 90.365 2.565 ;
      RECT 90.195 6.315 90.365 6.485 ;
      RECT 89.95 0.105 90.12 0.275 ;
      RECT 89.95 8.605 90.12 8.775 ;
      RECT 89.27 0.105 89.44 0.275 ;
      RECT 89.27 8.605 89.44 8.775 ;
      RECT 87.99 1.565 88.16 1.735 ;
      RECT 87.53 1.565 87.7 1.735 ;
      RECT 87.135 2.905 87.305 3.075 ;
      RECT 87.07 1.565 87.24 1.735 ;
      RECT 86.925 2.245 87.095 2.415 ;
      RECT 86.61 1.565 86.78 1.735 ;
      RECT 86.61 3.155 86.78 3.325 ;
      RECT 86.55 8.605 86.72 8.775 ;
      RECT 86.24 6.685 86.41 6.855 ;
      RECT 86.225 2.75 86.395 2.92 ;
      RECT 86.15 1.565 86.32 1.735 ;
      RECT 86.01 3.315 86.18 3.485 ;
      RECT 85.99 3.715 86.16 3.885 ;
      RECT 85.87 8.605 86.04 8.775 ;
      RECT 85.815 2.27 85.985 2.44 ;
      RECT 85.81 7.055 85.98 7.225 ;
      RECT 85.81 7.795 85.98 7.965 ;
      RECT 85.69 1.565 85.86 1.735 ;
      RECT 85.435 6.315 85.605 6.485 ;
      RECT 85.32 3.25 85.49 3.42 ;
      RECT 85.23 1.565 85.4 1.735 ;
      RECT 85.19 8.605 85.36 8.775 ;
      RECT 84.995 2.935 85.165 3.105 ;
      RECT 84.93 3.715 85.1 3.885 ;
      RECT 84.77 1.565 84.94 1.735 ;
      RECT 84.53 3.7 84.7 3.87 ;
      RECT 84.51 8.605 84.68 8.775 ;
      RECT 84.49 2.185 84.66 2.355 ;
      RECT 84.31 1.565 84.48 1.735 ;
      RECT 83.85 1.565 84.02 1.735 ;
      RECT 83.59 2.685 83.76 2.855 ;
      RECT 83.59 3.145 83.76 3.315 ;
      RECT 83.59 3.66 83.76 3.83 ;
      RECT 83.475 2.22 83.645 2.39 ;
      RECT 83.39 1.565 83.56 1.735 ;
      RECT 83.01 3.73 83.18 3.9 ;
      RECT 82.93 1.565 83.1 1.735 ;
      RECT 82.53 2.26 82.7 2.43 ;
      RECT 82.47 1.565 82.64 1.735 ;
      RECT 82.315 2.635 82.485 2.805 ;
      RECT 82.01 1.565 82.18 1.735 ;
      RECT 81.815 3.235 81.985 3.405 ;
      RECT 81.7 2.685 81.87 2.855 ;
      RECT 81.55 1.565 81.72 1.735 ;
      RECT 81.53 2.135 81.7 2.305 ;
      RECT 81.155 3.165 81.325 3.335 ;
      RECT 81.09 1.565 81.26 1.735 ;
      RECT 80.67 2.765 80.84 2.935 ;
      RECT 80.63 1.565 80.8 1.735 ;
      RECT 80.62 3.54 80.79 3.71 ;
      RECT 80.17 1.565 80.34 1.735 ;
      RECT 80.13 3.165 80.3 3.335 ;
      RECT 80.095 2.27 80.265 2.44 ;
      RECT 79.735 2.67 79.905 2.84 ;
      RECT 79.71 1.565 79.88 1.735 ;
      RECT 79.53 3.48 79.7 3.65 ;
      RECT 79.25 1.565 79.42 1.735 ;
      RECT 79.225 2.91 79.395 3.08 ;
      RECT 78.79 1.565 78.96 1.735 ;
      RECT 78.525 2.7 78.695 2.87 ;
      RECT 78.33 1.565 78.5 1.735 ;
      RECT 78.205 3.145 78.375 3.315 ;
      RECT 77.87 1.565 78.04 1.735 ;
      RECT 77.79 3.18 77.96 3.35 ;
      RECT 77.62 2.165 77.79 2.335 ;
      RECT 77.445 2.62 77.615 2.79 ;
      RECT 77.41 1.565 77.58 1.735 ;
      RECT 76.95 1.565 77.12 1.735 ;
      RECT 76.525 2.27 76.695 2.44 ;
      RECT 76.52 3.585 76.69 3.755 ;
      RECT 76.49 1.565 76.66 1.735 ;
      RECT 75.425 7.8 75.595 7.97 ;
      RECT 75.075 0.1 75.245 0.27 ;
      RECT 75.075 8.61 75.245 8.78 ;
      RECT 75.055 2.76 75.225 2.93 ;
      RECT 75.055 5.95 75.225 6.12 ;
      RECT 74.435 0.91 74.605 1.08 ;
      RECT 74.435 2.39 74.605 2.56 ;
      RECT 74.435 6.32 74.605 6.49 ;
      RECT 74.435 7.8 74.605 7.97 ;
      RECT 74.085 0.1 74.255 0.27 ;
      RECT 74.085 8.61 74.255 8.78 ;
      RECT 74.065 2.76 74.235 2.93 ;
      RECT 74.065 5.95 74.235 6.12 ;
      RECT 73.385 0.105 73.555 0.275 ;
      RECT 73.385 8.605 73.555 8.775 ;
      RECT 73.075 2.025 73.245 2.195 ;
      RECT 73.075 6.685 73.245 6.855 ;
      RECT 72.705 0.105 72.875 0.275 ;
      RECT 72.705 8.605 72.875 8.775 ;
      RECT 72.645 0.915 72.815 1.085 ;
      RECT 72.645 1.655 72.815 1.825 ;
      RECT 72.645 7.055 72.815 7.225 ;
      RECT 72.645 7.795 72.815 7.965 ;
      RECT 72.27 2.395 72.44 2.565 ;
      RECT 72.27 6.315 72.44 6.485 ;
      RECT 72.025 0.105 72.195 0.275 ;
      RECT 72.025 8.605 72.195 8.775 ;
      RECT 71.345 0.105 71.515 0.275 ;
      RECT 71.345 8.605 71.515 8.775 ;
      RECT 70.065 1.565 70.235 1.735 ;
      RECT 69.605 1.565 69.775 1.735 ;
      RECT 69.21 2.905 69.38 3.075 ;
      RECT 69.145 1.565 69.315 1.735 ;
      RECT 69 2.245 69.17 2.415 ;
      RECT 68.685 1.565 68.855 1.735 ;
      RECT 68.685 3.155 68.855 3.325 ;
      RECT 68.625 8.605 68.795 8.775 ;
      RECT 68.315 6.685 68.485 6.855 ;
      RECT 68.3 2.75 68.47 2.92 ;
      RECT 68.225 1.565 68.395 1.735 ;
      RECT 68.085 3.315 68.255 3.485 ;
      RECT 68.065 3.715 68.235 3.885 ;
      RECT 67.945 8.605 68.115 8.775 ;
      RECT 67.89 2.27 68.06 2.44 ;
      RECT 67.885 7.055 68.055 7.225 ;
      RECT 67.885 7.795 68.055 7.965 ;
      RECT 67.765 1.565 67.935 1.735 ;
      RECT 67.51 6.315 67.68 6.485 ;
      RECT 67.395 3.25 67.565 3.42 ;
      RECT 67.305 1.565 67.475 1.735 ;
      RECT 67.265 8.605 67.435 8.775 ;
      RECT 67.07 2.935 67.24 3.105 ;
      RECT 67.005 3.715 67.175 3.885 ;
      RECT 66.845 1.565 67.015 1.735 ;
      RECT 66.605 3.7 66.775 3.87 ;
      RECT 66.585 8.605 66.755 8.775 ;
      RECT 66.565 2.185 66.735 2.355 ;
      RECT 66.385 1.565 66.555 1.735 ;
      RECT 65.925 1.565 66.095 1.735 ;
      RECT 65.665 2.685 65.835 2.855 ;
      RECT 65.665 3.145 65.835 3.315 ;
      RECT 65.665 3.66 65.835 3.83 ;
      RECT 65.55 2.22 65.72 2.39 ;
      RECT 65.465 1.565 65.635 1.735 ;
      RECT 65.085 3.73 65.255 3.9 ;
      RECT 65.005 1.565 65.175 1.735 ;
      RECT 64.605 2.26 64.775 2.43 ;
      RECT 64.545 1.565 64.715 1.735 ;
      RECT 64.39 2.635 64.56 2.805 ;
      RECT 64.085 1.565 64.255 1.735 ;
      RECT 63.89 3.235 64.06 3.405 ;
      RECT 63.775 2.685 63.945 2.855 ;
      RECT 63.625 1.565 63.795 1.735 ;
      RECT 63.605 2.135 63.775 2.305 ;
      RECT 63.23 3.165 63.4 3.335 ;
      RECT 63.165 1.565 63.335 1.735 ;
      RECT 62.745 2.765 62.915 2.935 ;
      RECT 62.705 1.565 62.875 1.735 ;
      RECT 62.695 3.54 62.865 3.71 ;
      RECT 62.245 1.565 62.415 1.735 ;
      RECT 62.205 3.165 62.375 3.335 ;
      RECT 62.17 2.27 62.34 2.44 ;
      RECT 61.81 2.67 61.98 2.84 ;
      RECT 61.785 1.565 61.955 1.735 ;
      RECT 61.605 3.48 61.775 3.65 ;
      RECT 61.325 1.565 61.495 1.735 ;
      RECT 61.3 2.91 61.47 3.08 ;
      RECT 60.865 1.565 61.035 1.735 ;
      RECT 60.6 2.7 60.77 2.87 ;
      RECT 60.405 1.565 60.575 1.735 ;
      RECT 60.28 3.145 60.45 3.315 ;
      RECT 59.945 1.565 60.115 1.735 ;
      RECT 59.865 3.18 60.035 3.35 ;
      RECT 59.695 2.165 59.865 2.335 ;
      RECT 59.52 2.62 59.69 2.79 ;
      RECT 59.485 1.565 59.655 1.735 ;
      RECT 59.025 1.565 59.195 1.735 ;
      RECT 58.6 2.27 58.77 2.44 ;
      RECT 58.595 3.585 58.765 3.755 ;
      RECT 58.565 1.565 58.735 1.735 ;
      RECT 57.5 7.8 57.67 7.97 ;
      RECT 57.15 0.1 57.32 0.27 ;
      RECT 57.15 8.61 57.32 8.78 ;
      RECT 57.13 2.76 57.3 2.93 ;
      RECT 57.13 5.95 57.3 6.12 ;
      RECT 56.51 0.91 56.68 1.08 ;
      RECT 56.51 2.39 56.68 2.56 ;
      RECT 56.51 6.32 56.68 6.49 ;
      RECT 56.51 7.8 56.68 7.97 ;
      RECT 56.16 0.1 56.33 0.27 ;
      RECT 56.16 8.61 56.33 8.78 ;
      RECT 56.14 2.76 56.31 2.93 ;
      RECT 56.14 5.95 56.31 6.12 ;
      RECT 55.46 0.105 55.63 0.275 ;
      RECT 55.46 8.605 55.63 8.775 ;
      RECT 55.15 2.025 55.32 2.195 ;
      RECT 55.15 6.685 55.32 6.855 ;
      RECT 54.78 0.105 54.95 0.275 ;
      RECT 54.78 8.605 54.95 8.775 ;
      RECT 54.72 0.915 54.89 1.085 ;
      RECT 54.72 1.655 54.89 1.825 ;
      RECT 54.72 7.055 54.89 7.225 ;
      RECT 54.72 7.795 54.89 7.965 ;
      RECT 54.345 2.395 54.515 2.565 ;
      RECT 54.345 6.315 54.515 6.485 ;
      RECT 54.1 0.105 54.27 0.275 ;
      RECT 54.1 8.605 54.27 8.775 ;
      RECT 53.42 0.105 53.59 0.275 ;
      RECT 53.42 8.605 53.59 8.775 ;
      RECT 52.14 1.565 52.31 1.735 ;
      RECT 51.68 1.565 51.85 1.735 ;
      RECT 51.285 2.905 51.455 3.075 ;
      RECT 51.22 1.565 51.39 1.735 ;
      RECT 51.075 2.245 51.245 2.415 ;
      RECT 50.76 1.565 50.93 1.735 ;
      RECT 50.76 3.155 50.93 3.325 ;
      RECT 50.7 8.605 50.87 8.775 ;
      RECT 50.39 6.685 50.56 6.855 ;
      RECT 50.375 2.75 50.545 2.92 ;
      RECT 50.3 1.565 50.47 1.735 ;
      RECT 50.16 3.315 50.33 3.485 ;
      RECT 50.14 3.715 50.31 3.885 ;
      RECT 50.02 8.605 50.19 8.775 ;
      RECT 49.965 2.27 50.135 2.44 ;
      RECT 49.96 7.055 50.13 7.225 ;
      RECT 49.96 7.795 50.13 7.965 ;
      RECT 49.84 1.565 50.01 1.735 ;
      RECT 49.585 6.315 49.755 6.485 ;
      RECT 49.47 3.25 49.64 3.42 ;
      RECT 49.38 1.565 49.55 1.735 ;
      RECT 49.34 8.605 49.51 8.775 ;
      RECT 49.145 2.935 49.315 3.105 ;
      RECT 49.08 3.715 49.25 3.885 ;
      RECT 48.92 1.565 49.09 1.735 ;
      RECT 48.68 3.7 48.85 3.87 ;
      RECT 48.66 8.605 48.83 8.775 ;
      RECT 48.64 2.185 48.81 2.355 ;
      RECT 48.46 1.565 48.63 1.735 ;
      RECT 48 1.565 48.17 1.735 ;
      RECT 47.74 2.685 47.91 2.855 ;
      RECT 47.74 3.145 47.91 3.315 ;
      RECT 47.74 3.66 47.91 3.83 ;
      RECT 47.625 2.22 47.795 2.39 ;
      RECT 47.54 1.565 47.71 1.735 ;
      RECT 47.16 3.73 47.33 3.9 ;
      RECT 47.08 1.565 47.25 1.735 ;
      RECT 46.68 2.26 46.85 2.43 ;
      RECT 46.62 1.565 46.79 1.735 ;
      RECT 46.465 2.635 46.635 2.805 ;
      RECT 46.16 1.565 46.33 1.735 ;
      RECT 45.965 3.235 46.135 3.405 ;
      RECT 45.85 2.685 46.02 2.855 ;
      RECT 45.7 1.565 45.87 1.735 ;
      RECT 45.68 2.135 45.85 2.305 ;
      RECT 45.305 3.165 45.475 3.335 ;
      RECT 45.24 1.565 45.41 1.735 ;
      RECT 44.82 2.765 44.99 2.935 ;
      RECT 44.78 1.565 44.95 1.735 ;
      RECT 44.77 3.54 44.94 3.71 ;
      RECT 44.32 1.565 44.49 1.735 ;
      RECT 44.28 3.165 44.45 3.335 ;
      RECT 44.245 2.27 44.415 2.44 ;
      RECT 43.885 2.67 44.055 2.84 ;
      RECT 43.86 1.565 44.03 1.735 ;
      RECT 43.68 3.48 43.85 3.65 ;
      RECT 43.4 1.565 43.57 1.735 ;
      RECT 43.375 2.91 43.545 3.08 ;
      RECT 42.94 1.565 43.11 1.735 ;
      RECT 42.675 2.7 42.845 2.87 ;
      RECT 42.48 1.565 42.65 1.735 ;
      RECT 42.355 3.145 42.525 3.315 ;
      RECT 42.02 1.565 42.19 1.735 ;
      RECT 41.94 3.18 42.11 3.35 ;
      RECT 41.77 2.165 41.94 2.335 ;
      RECT 41.595 2.62 41.765 2.79 ;
      RECT 41.56 1.565 41.73 1.735 ;
      RECT 41.1 1.565 41.27 1.735 ;
      RECT 40.675 2.27 40.845 2.44 ;
      RECT 40.67 3.585 40.84 3.755 ;
      RECT 40.64 1.565 40.81 1.735 ;
      RECT 39.575 7.8 39.745 7.97 ;
      RECT 39.225 0.1 39.395 0.27 ;
      RECT 39.225 8.61 39.395 8.78 ;
      RECT 39.205 2.76 39.375 2.93 ;
      RECT 39.205 5.95 39.375 6.12 ;
      RECT 38.585 0.91 38.755 1.08 ;
      RECT 38.585 2.39 38.755 2.56 ;
      RECT 38.585 6.32 38.755 6.49 ;
      RECT 38.585 7.8 38.755 7.97 ;
      RECT 38.235 0.1 38.405 0.27 ;
      RECT 38.235 8.61 38.405 8.78 ;
      RECT 38.215 2.76 38.385 2.93 ;
      RECT 38.215 5.95 38.385 6.12 ;
      RECT 37.535 0.105 37.705 0.275 ;
      RECT 37.535 8.605 37.705 8.775 ;
      RECT 37.225 2.025 37.395 2.195 ;
      RECT 37.225 6.685 37.395 6.855 ;
      RECT 36.855 0.105 37.025 0.275 ;
      RECT 36.855 8.605 37.025 8.775 ;
      RECT 36.795 0.915 36.965 1.085 ;
      RECT 36.795 1.655 36.965 1.825 ;
      RECT 36.795 7.055 36.965 7.225 ;
      RECT 36.795 7.795 36.965 7.965 ;
      RECT 36.42 2.395 36.59 2.565 ;
      RECT 36.42 6.315 36.59 6.485 ;
      RECT 36.175 0.105 36.345 0.275 ;
      RECT 36.175 8.605 36.345 8.775 ;
      RECT 35.495 0.105 35.665 0.275 ;
      RECT 35.495 8.605 35.665 8.775 ;
      RECT 34.215 1.565 34.385 1.735 ;
      RECT 33.755 1.565 33.925 1.735 ;
      RECT 33.36 2.905 33.53 3.075 ;
      RECT 33.295 1.565 33.465 1.735 ;
      RECT 33.15 2.245 33.32 2.415 ;
      RECT 32.835 1.565 33.005 1.735 ;
      RECT 32.835 3.155 33.005 3.325 ;
      RECT 32.775 8.605 32.945 8.775 ;
      RECT 32.465 6.685 32.635 6.855 ;
      RECT 32.45 2.75 32.62 2.92 ;
      RECT 32.375 1.565 32.545 1.735 ;
      RECT 32.235 3.315 32.405 3.485 ;
      RECT 32.215 3.715 32.385 3.885 ;
      RECT 32.095 8.605 32.265 8.775 ;
      RECT 32.04 2.27 32.21 2.44 ;
      RECT 32.035 7.055 32.205 7.225 ;
      RECT 32.035 7.795 32.205 7.965 ;
      RECT 31.915 1.565 32.085 1.735 ;
      RECT 31.66 6.315 31.83 6.485 ;
      RECT 31.545 3.25 31.715 3.42 ;
      RECT 31.455 1.565 31.625 1.735 ;
      RECT 31.415 8.605 31.585 8.775 ;
      RECT 31.22 2.935 31.39 3.105 ;
      RECT 31.155 3.715 31.325 3.885 ;
      RECT 30.995 1.565 31.165 1.735 ;
      RECT 30.755 3.7 30.925 3.87 ;
      RECT 30.735 8.605 30.905 8.775 ;
      RECT 30.715 2.185 30.885 2.355 ;
      RECT 30.535 1.565 30.705 1.735 ;
      RECT 30.075 1.565 30.245 1.735 ;
      RECT 29.815 2.685 29.985 2.855 ;
      RECT 29.815 3.145 29.985 3.315 ;
      RECT 29.815 3.66 29.985 3.83 ;
      RECT 29.7 2.22 29.87 2.39 ;
      RECT 29.615 1.565 29.785 1.735 ;
      RECT 29.235 3.73 29.405 3.9 ;
      RECT 29.155 1.565 29.325 1.735 ;
      RECT 28.755 2.26 28.925 2.43 ;
      RECT 28.695 1.565 28.865 1.735 ;
      RECT 28.54 2.635 28.71 2.805 ;
      RECT 28.235 1.565 28.405 1.735 ;
      RECT 28.04 3.235 28.21 3.405 ;
      RECT 27.925 2.685 28.095 2.855 ;
      RECT 27.775 1.565 27.945 1.735 ;
      RECT 27.755 2.135 27.925 2.305 ;
      RECT 27.38 3.165 27.55 3.335 ;
      RECT 27.315 1.565 27.485 1.735 ;
      RECT 26.895 2.765 27.065 2.935 ;
      RECT 26.855 1.565 27.025 1.735 ;
      RECT 26.845 3.54 27.015 3.71 ;
      RECT 26.395 1.565 26.565 1.735 ;
      RECT 26.355 3.165 26.525 3.335 ;
      RECT 26.32 2.27 26.49 2.44 ;
      RECT 25.96 2.67 26.13 2.84 ;
      RECT 25.935 1.565 26.105 1.735 ;
      RECT 25.755 3.48 25.925 3.65 ;
      RECT 25.475 1.565 25.645 1.735 ;
      RECT 25.45 2.91 25.62 3.08 ;
      RECT 25.015 1.565 25.185 1.735 ;
      RECT 24.75 2.7 24.92 2.87 ;
      RECT 24.555 1.565 24.725 1.735 ;
      RECT 24.43 3.145 24.6 3.315 ;
      RECT 24.095 1.565 24.265 1.735 ;
      RECT 24.015 3.18 24.185 3.35 ;
      RECT 23.845 2.165 24.015 2.335 ;
      RECT 23.67 2.62 23.84 2.79 ;
      RECT 23.635 1.565 23.805 1.735 ;
      RECT 23.175 1.565 23.345 1.735 ;
      RECT 22.75 2.27 22.92 2.44 ;
      RECT 22.745 3.585 22.915 3.755 ;
      RECT 22.715 1.565 22.885 1.735 ;
      RECT 21.65 7.8 21.82 7.97 ;
      RECT 21.3 0.1 21.47 0.27 ;
      RECT 21.3 8.61 21.47 8.78 ;
      RECT 21.28 2.76 21.45 2.93 ;
      RECT 21.28 5.95 21.45 6.12 ;
      RECT 20.66 0.91 20.83 1.08 ;
      RECT 20.66 2.39 20.83 2.56 ;
      RECT 20.66 6.32 20.83 6.49 ;
      RECT 20.66 7.8 20.83 7.97 ;
      RECT 20.31 0.1 20.48 0.27 ;
      RECT 20.31 8.61 20.48 8.78 ;
      RECT 20.29 2.76 20.46 2.93 ;
      RECT 20.29 5.95 20.46 6.12 ;
      RECT 19.61 0.105 19.78 0.275 ;
      RECT 19.61 8.605 19.78 8.775 ;
      RECT 19.3 2.025 19.47 2.195 ;
      RECT 19.3 6.685 19.47 6.855 ;
      RECT 18.93 0.105 19.1 0.275 ;
      RECT 18.93 8.605 19.1 8.775 ;
      RECT 18.87 0.915 19.04 1.085 ;
      RECT 18.87 1.655 19.04 1.825 ;
      RECT 18.87 7.055 19.04 7.225 ;
      RECT 18.87 7.795 19.04 7.965 ;
      RECT 18.495 2.395 18.665 2.565 ;
      RECT 18.495 6.315 18.665 6.485 ;
      RECT 18.25 0.105 18.42 0.275 ;
      RECT 18.25 8.605 18.42 8.775 ;
      RECT 17.57 0.105 17.74 0.275 ;
      RECT 17.57 8.605 17.74 8.775 ;
      RECT 16.29 1.565 16.46 1.735 ;
      RECT 15.83 1.565 16 1.735 ;
      RECT 15.435 2.905 15.605 3.075 ;
      RECT 15.37 1.565 15.54 1.735 ;
      RECT 15.225 2.245 15.395 2.415 ;
      RECT 14.91 1.565 15.08 1.735 ;
      RECT 14.91 3.155 15.08 3.325 ;
      RECT 14.85 8.605 15.02 8.775 ;
      RECT 14.54 6.685 14.71 6.855 ;
      RECT 14.525 2.75 14.695 2.92 ;
      RECT 14.45 1.565 14.62 1.735 ;
      RECT 14.31 3.315 14.48 3.485 ;
      RECT 14.29 3.715 14.46 3.885 ;
      RECT 14.17 8.605 14.34 8.775 ;
      RECT 14.115 2.27 14.285 2.44 ;
      RECT 14.11 7.055 14.28 7.225 ;
      RECT 14.11 7.795 14.28 7.965 ;
      RECT 13.99 1.565 14.16 1.735 ;
      RECT 13.735 6.315 13.905 6.485 ;
      RECT 13.62 3.25 13.79 3.42 ;
      RECT 13.53 1.565 13.7 1.735 ;
      RECT 13.49 8.605 13.66 8.775 ;
      RECT 13.295 2.935 13.465 3.105 ;
      RECT 13.23 3.715 13.4 3.885 ;
      RECT 13.07 1.565 13.24 1.735 ;
      RECT 12.83 3.7 13 3.87 ;
      RECT 12.81 8.605 12.98 8.775 ;
      RECT 12.79 2.185 12.96 2.355 ;
      RECT 12.61 1.565 12.78 1.735 ;
      RECT 12.15 1.565 12.32 1.735 ;
      RECT 11.89 2.685 12.06 2.855 ;
      RECT 11.89 3.145 12.06 3.315 ;
      RECT 11.89 3.66 12.06 3.83 ;
      RECT 11.775 2.22 11.945 2.39 ;
      RECT 11.69 1.565 11.86 1.735 ;
      RECT 11.31 3.73 11.48 3.9 ;
      RECT 11.23 1.565 11.4 1.735 ;
      RECT 10.83 2.26 11 2.43 ;
      RECT 10.77 1.565 10.94 1.735 ;
      RECT 10.615 2.635 10.785 2.805 ;
      RECT 10.31 1.565 10.48 1.735 ;
      RECT 10.115 3.235 10.285 3.405 ;
      RECT 10 2.685 10.17 2.855 ;
      RECT 9.85 1.565 10.02 1.735 ;
      RECT 9.83 2.135 10 2.305 ;
      RECT 9.455 3.165 9.625 3.335 ;
      RECT 9.39 1.565 9.56 1.735 ;
      RECT 8.97 2.765 9.14 2.935 ;
      RECT 8.93 1.565 9.1 1.735 ;
      RECT 8.92 3.54 9.09 3.71 ;
      RECT 8.47 1.565 8.64 1.735 ;
      RECT 8.43 3.165 8.6 3.335 ;
      RECT 8.395 2.27 8.565 2.44 ;
      RECT 8.035 2.67 8.205 2.84 ;
      RECT 8.01 1.565 8.18 1.735 ;
      RECT 7.83 3.48 8 3.65 ;
      RECT 7.55 1.565 7.72 1.735 ;
      RECT 7.525 2.91 7.695 3.08 ;
      RECT 7.09 1.565 7.26 1.735 ;
      RECT 6.825 2.7 6.995 2.87 ;
      RECT 6.63 1.565 6.8 1.735 ;
      RECT 6.505 3.145 6.675 3.315 ;
      RECT 6.17 1.565 6.34 1.735 ;
      RECT 6.09 3.18 6.26 3.35 ;
      RECT 5.92 2.165 6.09 2.335 ;
      RECT 5.745 2.62 5.915 2.79 ;
      RECT 5.71 1.565 5.88 1.735 ;
      RECT 5.25 1.565 5.42 1.735 ;
      RECT 4.825 2.27 4.995 2.44 ;
      RECT 4.82 3.585 4.99 3.755 ;
      RECT 4.79 1.565 4.96 1.735 ;
      RECT 3.82 8.605 3.99 8.775 ;
      RECT 3.14 8.605 3.31 8.775 ;
      RECT 3.08 7.055 3.25 7.225 ;
      RECT 3.08 7.795 3.25 7.965 ;
      RECT 2.705 6.315 2.875 6.485 ;
      RECT 2.46 8.605 2.63 8.775 ;
      RECT 1.78 8.605 1.95 8.775 ;
    LAYER li1 ;
      RECT 87.395 0 87.565 2.235 ;
      RECT 86.435 0 86.605 2.235 ;
      RECT 85.475 0 85.645 2.235 ;
      RECT 84.955 0 85.125 2.235 ;
      RECT 83.995 0 84.165 2.235 ;
      RECT 82.995 0 83.165 2.235 ;
      RECT 82.035 0 82.205 2.235 ;
      RECT 80.555 0 80.725 2.235 ;
      RECT 78.635 0 78.805 2.235 ;
      RECT 77.155 0 77.325 2.235 ;
      RECT 69.47 0 69.64 2.235 ;
      RECT 68.51 0 68.68 2.235 ;
      RECT 67.55 0 67.72 2.235 ;
      RECT 67.03 0 67.2 2.235 ;
      RECT 66.07 0 66.24 2.235 ;
      RECT 65.07 0 65.24 2.235 ;
      RECT 64.11 0 64.28 2.235 ;
      RECT 62.63 0 62.8 2.235 ;
      RECT 60.71 0 60.88 2.235 ;
      RECT 59.23 0 59.4 2.235 ;
      RECT 51.545 0 51.715 2.235 ;
      RECT 50.585 0 50.755 2.235 ;
      RECT 49.625 0 49.795 2.235 ;
      RECT 49.105 0 49.275 2.235 ;
      RECT 48.145 0 48.315 2.235 ;
      RECT 47.145 0 47.315 2.235 ;
      RECT 46.185 0 46.355 2.235 ;
      RECT 44.705 0 44.875 2.235 ;
      RECT 42.785 0 42.955 2.235 ;
      RECT 41.305 0 41.475 2.235 ;
      RECT 33.62 0 33.79 2.235 ;
      RECT 32.66 0 32.83 2.235 ;
      RECT 31.7 0 31.87 2.235 ;
      RECT 31.18 0 31.35 2.235 ;
      RECT 30.22 0 30.39 2.235 ;
      RECT 29.22 0 29.39 2.235 ;
      RECT 28.26 0 28.43 2.235 ;
      RECT 26.78 0 26.95 2.235 ;
      RECT 24.86 0 25.03 2.235 ;
      RECT 23.38 0 23.55 2.235 ;
      RECT 15.695 0 15.865 2.235 ;
      RECT 14.735 0 14.905 2.235 ;
      RECT 13.775 0 13.945 2.235 ;
      RECT 13.255 0 13.425 2.235 ;
      RECT 12.295 0 12.465 2.235 ;
      RECT 11.295 0 11.465 2.235 ;
      RECT 10.335 0 10.505 2.235 ;
      RECT 8.855 0 9.025 2.235 ;
      RECT 6.935 0 7.105 2.235 ;
      RECT 5.455 0 5.625 2.235 ;
      RECT 76.345 0 88.305 1.735 ;
      RECT 58.42 0 70.38 1.735 ;
      RECT 40.495 0 52.455 1.735 ;
      RECT 22.57 0 34.53 1.735 ;
      RECT 4.645 0 16.605 1.735 ;
      RECT 76.34 0 88.305 1.68 ;
      RECT 58.415 0 70.38 1.68 ;
      RECT 40.49 0 52.455 1.68 ;
      RECT 22.565 0 34.53 1.68 ;
      RECT 4.64 0 16.605 1.68 ;
      RECT 89.19 0 89.36 0.935 ;
      RECT 71.265 0 71.435 0.935 ;
      RECT 53.34 0 53.51 0.935 ;
      RECT 35.415 0 35.585 0.935 ;
      RECT 17.49 0 17.66 0.935 ;
      RECT 92.92 0 93.09 0.93 ;
      RECT 91.93 0 92.1 0.93 ;
      RECT 74.995 0 75.165 0.93 ;
      RECT 74.005 0 74.175 0.93 ;
      RECT 57.07 0 57.24 0.93 ;
      RECT 56.08 0 56.25 0.93 ;
      RECT 39.145 0 39.315 0.93 ;
      RECT 38.155 0 38.325 0.93 ;
      RECT 21.22 0 21.39 0.93 ;
      RECT 20.23 0 20.4 0.93 ;
      RECT 93.715 0 93.895 0.305 ;
      RECT 75.79 0 91.765 0.305 ;
      RECT 57.865 0 73.84 0.305 ;
      RECT 39.94 0 55.915 0.305 ;
      RECT 22.015 0 37.99 0.305 ;
      RECT 1.48 0 20.065 0.305 ;
      RECT 1.48 0 93.895 0.3 ;
      RECT 1.46 8.58 93.895 8.88 ;
      RECT 93.715 8.575 93.895 8.88 ;
      RECT 92.92 7.95 93.09 8.88 ;
      RECT 91.93 7.95 92.1 8.88 ;
      RECT 75.79 8.575 91.765 8.88 ;
      RECT 74.995 7.95 75.165 8.88 ;
      RECT 74.005 7.95 74.175 8.88 ;
      RECT 57.865 8.575 73.84 8.88 ;
      RECT 57.07 7.95 57.24 8.88 ;
      RECT 56.08 7.95 56.25 8.88 ;
      RECT 39.94 8.575 55.915 8.88 ;
      RECT 39.145 7.95 39.315 8.88 ;
      RECT 38.155 7.95 38.325 8.88 ;
      RECT 22.015 8.575 37.99 8.88 ;
      RECT 21.22 7.95 21.39 8.88 ;
      RECT 20.23 7.95 20.4 8.88 ;
      RECT 1.46 8.575 20.065 8.88 ;
      RECT 89.19 7.945 89.36 8.88 ;
      RECT 84.43 7.945 84.6 8.88 ;
      RECT 71.265 7.945 71.435 8.88 ;
      RECT 66.505 7.945 66.675 8.88 ;
      RECT 53.34 7.945 53.51 8.88 ;
      RECT 48.58 7.945 48.75 8.88 ;
      RECT 35.415 7.945 35.585 8.88 ;
      RECT 30.655 7.945 30.825 8.88 ;
      RECT 17.49 7.945 17.66 8.88 ;
      RECT 12.73 7.945 12.9 8.88 ;
      RECT 1.7 7.945 1.87 8.88 ;
      RECT 93.35 5.02 93.52 6.49 ;
      RECT 93.35 6.315 93.525 6.485 ;
      RECT 92.98 1.74 93.15 2.93 ;
      RECT 92.98 1.74 93.45 1.91 ;
      RECT 92.98 6.97 93.45 7.14 ;
      RECT 92.98 5.95 93.15 7.14 ;
      RECT 91.99 1.74 92.16 2.93 ;
      RECT 91.99 1.74 92.46 1.91 ;
      RECT 91.99 6.97 92.46 7.14 ;
      RECT 91.99 5.95 92.16 7.14 ;
      RECT 90.14 2.635 90.31 3.865 ;
      RECT 90.195 0.855 90.365 2.805 ;
      RECT 90.14 0.575 90.31 1.025 ;
      RECT 90.14 7.855 90.31 8.305 ;
      RECT 90.195 6.075 90.365 8.025 ;
      RECT 90.14 5.015 90.31 6.245 ;
      RECT 89.62 0.575 89.79 3.865 ;
      RECT 89.62 2.075 90.025 2.405 ;
      RECT 89.62 1.235 90.025 1.565 ;
      RECT 89.62 5.015 89.79 8.305 ;
      RECT 89.62 7.315 90.025 7.645 ;
      RECT 89.62 6.475 90.025 6.805 ;
      RECT 87.72 3.392 87.735 3.443 ;
      RECT 87.715 3.372 87.72 3.49 ;
      RECT 87.7 3.362 87.715 3.558 ;
      RECT 87.675 3.342 87.7 3.613 ;
      RECT 87.635 3.327 87.675 3.633 ;
      RECT 87.59 3.321 87.635 3.661 ;
      RECT 87.52 3.311 87.59 3.678 ;
      RECT 87.5 3.303 87.52 3.678 ;
      RECT 87.44 3.297 87.5 3.67 ;
      RECT 87.381 3.288 87.44 3.658 ;
      RECT 87.295 3.277 87.381 3.641 ;
      RECT 87.273 3.268 87.295 3.629 ;
      RECT 87.187 3.261 87.273 3.616 ;
      RECT 87.101 3.248 87.187 3.597 ;
      RECT 87.015 3.236 87.101 3.577 ;
      RECT 86.985 3.225 87.015 3.564 ;
      RECT 86.935 3.211 86.985 3.556 ;
      RECT 86.915 3.2 86.935 3.548 ;
      RECT 86.866 3.189 86.915 3.54 ;
      RECT 86.78 3.168 86.866 3.525 ;
      RECT 86.735 3.155 86.78 3.51 ;
      RECT 86.69 3.155 86.735 3.49 ;
      RECT 86.635 3.155 86.69 3.425 ;
      RECT 86.61 3.155 86.635 3.348 ;
      RECT 87.135 2.892 87.305 3.075 ;
      RECT 87.135 2.892 87.32 3.033 ;
      RECT 87.135 2.892 87.325 2.975 ;
      RECT 87.195 2.66 87.33 2.951 ;
      RECT 87.195 2.664 87.335 2.934 ;
      RECT 87.14 2.827 87.335 2.934 ;
      RECT 87.165 2.672 87.305 3.075 ;
      RECT 87.165 2.676 87.345 2.875 ;
      RECT 87.15 2.762 87.345 2.875 ;
      RECT 87.16 2.692 87.305 3.075 ;
      RECT 87.16 2.695 87.355 2.788 ;
      RECT 87.155 2.712 87.355 2.788 ;
      RECT 86.925 1.932 87.095 2.415 ;
      RECT 86.92 1.927 87.07 2.405 ;
      RECT 86.92 1.934 87.1 2.399 ;
      RECT 86.91 1.928 87.07 2.378 ;
      RECT 86.91 1.944 87.115 2.337 ;
      RECT 86.88 1.929 87.07 2.3 ;
      RECT 86.88 1.959 87.125 2.24 ;
      RECT 86.875 1.931 87.07 2.238 ;
      RECT 86.855 1.94 87.1 2.195 ;
      RECT 86.83 1.956 87.115 2.107 ;
      RECT 86.83 1.975 87.14 2.098 ;
      RECT 86.825 2.012 87.14 2.05 ;
      RECT 86.83 1.992 87.145 2.018 ;
      RECT 86.925 1.926 87.035 2.415 ;
      RECT 87.011 1.925 87.035 2.415 ;
      RECT 86.245 2.71 86.25 2.921 ;
      RECT 86.845 2.71 86.85 2.895 ;
      RECT 86.91 2.75 86.915 2.863 ;
      RECT 86.905 2.742 86.91 2.869 ;
      RECT 86.9 2.732 86.905 2.877 ;
      RECT 86.895 2.722 86.9 2.886 ;
      RECT 86.89 2.712 86.895 2.89 ;
      RECT 86.85 2.71 86.89 2.893 ;
      RECT 86.822 2.709 86.845 2.897 ;
      RECT 86.736 2.706 86.822 2.904 ;
      RECT 86.65 2.702 86.736 2.915 ;
      RECT 86.63 2.7 86.65 2.921 ;
      RECT 86.612 2.699 86.63 2.924 ;
      RECT 86.526 2.697 86.612 2.931 ;
      RECT 86.44 2.692 86.526 2.944 ;
      RECT 86.421 2.689 86.44 2.949 ;
      RECT 86.335 2.687 86.421 2.94 ;
      RECT 86.325 2.687 86.335 2.933 ;
      RECT 86.25 2.7 86.325 2.927 ;
      RECT 86.235 2.711 86.245 2.921 ;
      RECT 86.225 2.713 86.235 2.92 ;
      RECT 86.215 2.717 86.225 2.916 ;
      RECT 86.21 2.72 86.215 2.91 ;
      RECT 86.2 2.722 86.21 2.904 ;
      RECT 86.195 2.725 86.2 2.898 ;
      RECT 86.175 3.311 86.18 3.515 ;
      RECT 86.16 3.298 86.175 3.608 ;
      RECT 86.145 3.279 86.16 3.885 ;
      RECT 86.11 3.245 86.145 3.885 ;
      RECT 86.106 3.215 86.11 3.885 ;
      RECT 86.02 3.097 86.106 3.885 ;
      RECT 86.01 2.972 86.02 3.885 ;
      RECT 85.995 2.94 86.01 3.885 ;
      RECT 85.99 2.915 85.995 3.885 ;
      RECT 85.985 2.905 85.99 3.841 ;
      RECT 85.97 2.877 85.985 3.746 ;
      RECT 85.955 2.843 85.97 3.645 ;
      RECT 85.95 2.821 85.955 3.598 ;
      RECT 85.945 2.81 85.95 3.568 ;
      RECT 85.94 2.8 85.945 3.534 ;
      RECT 85.93 2.787 85.94 3.502 ;
      RECT 85.905 2.763 85.93 3.428 ;
      RECT 85.9 2.743 85.905 3.353 ;
      RECT 85.895 2.737 85.9 3.328 ;
      RECT 85.89 2.732 85.895 3.293 ;
      RECT 85.885 2.727 85.89 3.268 ;
      RECT 85.88 2.725 85.885 3.248 ;
      RECT 85.875 2.725 85.88 3.233 ;
      RECT 85.87 2.725 85.875 3.193 ;
      RECT 85.86 2.725 85.87 3.165 ;
      RECT 85.85 2.725 85.86 3.11 ;
      RECT 85.835 2.725 85.85 3.048 ;
      RECT 85.83 2.724 85.835 2.993 ;
      RECT 85.815 2.723 85.83 2.973 ;
      RECT 85.755 2.721 85.815 2.947 ;
      RECT 85.72 2.722 85.755 2.927 ;
      RECT 85.715 2.724 85.72 2.917 ;
      RECT 85.705 2.743 85.715 2.907 ;
      RECT 85.7 2.77 85.705 2.838 ;
      RECT 85.815 2.195 85.985 2.44 ;
      RECT 85.85 1.966 85.985 2.44 ;
      RECT 85.85 1.968 85.995 2.435 ;
      RECT 85.85 1.97 86.02 2.423 ;
      RECT 85.85 1.973 86.045 2.405 ;
      RECT 85.85 1.978 86.095 2.378 ;
      RECT 85.85 1.983 86.115 2.343 ;
      RECT 85.83 1.985 86.125 2.318 ;
      RECT 85.82 2.08 86.125 2.318 ;
      RECT 85.85 1.965 85.96 2.44 ;
      RECT 85.86 1.962 85.955 2.44 ;
      RECT 85.38 3.227 85.57 3.585 ;
      RECT 85.38 3.239 85.605 3.584 ;
      RECT 85.38 3.267 85.625 3.582 ;
      RECT 85.38 3.292 85.63 3.581 ;
      RECT 85.38 3.35 85.645 3.58 ;
      RECT 85.365 3.223 85.525 3.565 ;
      RECT 85.345 3.232 85.57 3.518 ;
      RECT 85.32 3.243 85.605 3.455 ;
      RECT 85.32 3.327 85.64 3.455 ;
      RECT 85.32 3.302 85.635 3.455 ;
      RECT 85.38 3.218 85.525 3.585 ;
      RECT 85.466 3.217 85.525 3.585 ;
      RECT 85.466 3.216 85.51 3.585 ;
      RECT 85.38 7.855 85.55 8.305 ;
      RECT 85.435 6.075 85.605 8.025 ;
      RECT 85.38 5.015 85.55 6.245 ;
      RECT 84.86 5.015 85.03 8.305 ;
      RECT 84.86 7.315 85.265 7.645 ;
      RECT 84.86 6.475 85.265 6.805 ;
      RECT 85.165 2.732 85.17 3.11 ;
      RECT 85.16 2.7 85.165 3.11 ;
      RECT 85.155 2.672 85.16 3.11 ;
      RECT 85.15 2.652 85.155 3.11 ;
      RECT 85.095 2.635 85.15 3.11 ;
      RECT 85.055 2.62 85.095 3.11 ;
      RECT 85 2.607 85.055 3.11 ;
      RECT 84.965 2.598 85 3.11 ;
      RECT 84.961 2.596 84.965 3.109 ;
      RECT 84.875 2.592 84.961 3.092 ;
      RECT 84.79 2.584 84.875 3.055 ;
      RECT 84.78 2.58 84.79 3.028 ;
      RECT 84.77 2.58 84.78 3.01 ;
      RECT 84.76 2.582 84.77 2.993 ;
      RECT 84.755 2.587 84.76 2.979 ;
      RECT 84.75 2.591 84.755 2.966 ;
      RECT 84.74 2.596 84.75 2.95 ;
      RECT 84.725 2.61 84.74 2.925 ;
      RECT 84.72 2.616 84.725 2.905 ;
      RECT 84.715 2.618 84.72 2.898 ;
      RECT 84.71 2.622 84.715 2.773 ;
      RECT 84.89 3.422 85.135 3.885 ;
      RECT 84.81 3.395 85.13 3.881 ;
      RECT 84.74 3.43 85.135 3.874 ;
      RECT 84.53 3.685 85.135 3.87 ;
      RECT 84.71 3.453 85.135 3.87 ;
      RECT 84.55 3.645 85.135 3.87 ;
      RECT 84.7 3.465 85.135 3.87 ;
      RECT 84.585 3.582 85.135 3.87 ;
      RECT 84.64 3.507 85.135 3.87 ;
      RECT 84.89 3.372 85.13 3.885 ;
      RECT 84.92 3.365 85.13 3.885 ;
      RECT 84.91 3.367 85.13 3.885 ;
      RECT 84.92 3.362 85.05 3.885 ;
      RECT 84.475 1.925 84.561 2.364 ;
      RECT 84.47 1.925 84.561 2.362 ;
      RECT 84.47 1.925 84.63 2.361 ;
      RECT 84.47 1.925 84.66 2.358 ;
      RECT 84.455 1.932 84.66 2.349 ;
      RECT 84.455 1.932 84.665 2.345 ;
      RECT 84.45 1.942 84.665 2.338 ;
      RECT 84.445 1.947 84.665 2.313 ;
      RECT 84.445 1.947 84.68 2.295 ;
      RECT 84.47 1.925 84.7 2.21 ;
      RECT 84.44 1.952 84.7 2.208 ;
      RECT 84.45 1.945 84.705 2.146 ;
      RECT 84.44 2.067 84.71 2.129 ;
      RECT 84.425 1.962 84.705 2.08 ;
      RECT 84.42 1.972 84.705 1.98 ;
      RECT 84.5 2.743 84.505 2.82 ;
      RECT 84.49 2.737 84.5 3.01 ;
      RECT 84.48 2.729 84.49 3.031 ;
      RECT 84.47 2.72 84.48 3.053 ;
      RECT 84.465 2.715 84.47 3.07 ;
      RECT 84.425 2.715 84.465 3.11 ;
      RECT 84.405 2.715 84.425 3.165 ;
      RECT 84.4 2.715 84.405 3.193 ;
      RECT 84.39 2.715 84.4 3.208 ;
      RECT 84.355 2.715 84.39 3.25 ;
      RECT 84.35 2.715 84.355 3.293 ;
      RECT 84.34 2.715 84.35 3.308 ;
      RECT 84.325 2.715 84.34 3.328 ;
      RECT 84.31 2.715 84.325 3.355 ;
      RECT 84.305 2.716 84.31 3.373 ;
      RECT 84.285 2.717 84.305 3.38 ;
      RECT 84.23 2.718 84.285 3.4 ;
      RECT 84.22 2.719 84.23 3.414 ;
      RECT 84.215 2.722 84.22 3.413 ;
      RECT 84.175 2.795 84.215 3.411 ;
      RECT 84.16 2.875 84.175 3.409 ;
      RECT 84.135 2.93 84.16 3.407 ;
      RECT 84.12 2.995 84.135 3.406 ;
      RECT 84.075 3.027 84.12 3.403 ;
      RECT 83.99 3.05 84.075 3.398 ;
      RECT 83.965 3.07 83.99 3.393 ;
      RECT 83.895 3.075 83.965 3.389 ;
      RECT 83.875 3.077 83.895 3.386 ;
      RECT 83.79 3.088 83.875 3.38 ;
      RECT 83.785 3.099 83.79 3.375 ;
      RECT 83.775 3.101 83.785 3.375 ;
      RECT 83.74 3.105 83.775 3.373 ;
      RECT 83.69 3.115 83.74 3.36 ;
      RECT 83.67 3.123 83.69 3.345 ;
      RECT 83.59 3.135 83.67 3.328 ;
      RECT 83.755 2.685 83.925 2.895 ;
      RECT 83.871 2.681 83.925 2.895 ;
      RECT 83.676 2.685 83.925 2.886 ;
      RECT 83.676 2.685 83.93 2.875 ;
      RECT 83.59 2.685 83.93 2.866 ;
      RECT 83.59 2.693 83.94 2.81 ;
      RECT 83.59 2.705 83.945 2.723 ;
      RECT 83.59 2.712 83.95 2.715 ;
      RECT 83.785 2.683 83.925 2.895 ;
      RECT 83.54 3.628 83.785 3.96 ;
      RECT 83.535 3.62 83.54 3.957 ;
      RECT 83.505 3.64 83.785 3.938 ;
      RECT 83.485 3.672 83.785 3.911 ;
      RECT 83.535 3.625 83.712 3.957 ;
      RECT 83.535 3.622 83.626 3.957 ;
      RECT 83.475 1.97 83.645 2.39 ;
      RECT 83.47 1.97 83.645 2.388 ;
      RECT 83.47 1.97 83.67 2.378 ;
      RECT 83.47 1.97 83.69 2.353 ;
      RECT 83.465 1.97 83.69 2.348 ;
      RECT 83.465 1.97 83.7 2.338 ;
      RECT 83.465 1.97 83.705 2.333 ;
      RECT 83.465 1.975 83.71 2.328 ;
      RECT 83.465 2.007 83.725 2.318 ;
      RECT 83.465 2.077 83.75 2.301 ;
      RECT 83.445 2.077 83.75 2.293 ;
      RECT 83.445 2.137 83.76 2.27 ;
      RECT 83.445 2.177 83.77 2.215 ;
      RECT 83.43 1.97 83.705 2.195 ;
      RECT 83.42 1.985 83.71 2.093 ;
      RECT 83.01 3.375 83.18 3.9 ;
      RECT 83.005 3.375 83.18 3.893 ;
      RECT 82.995 3.375 83.185 3.858 ;
      RECT 82.99 3.385 83.185 3.83 ;
      RECT 82.985 3.405 83.185 3.813 ;
      RECT 82.995 3.38 83.19 3.803 ;
      RECT 82.98 3.425 83.19 3.795 ;
      RECT 82.975 3.445 83.19 3.78 ;
      RECT 82.97 3.475 83.19 3.77 ;
      RECT 82.96 3.52 83.19 3.745 ;
      RECT 82.99 3.39 83.195 3.728 ;
      RECT 82.955 3.572 83.195 3.723 ;
      RECT 82.99 3.4 83.2 3.693 ;
      RECT 82.95 3.605 83.2 3.69 ;
      RECT 82.945 3.63 83.2 3.67 ;
      RECT 82.985 3.417 83.21 3.61 ;
      RECT 82.98 3.439 83.22 3.503 ;
      RECT 82.93 2.686 82.945 2.955 ;
      RECT 82.885 2.67 82.93 3 ;
      RECT 82.88 2.658 82.885 3.05 ;
      RECT 82.87 2.654 82.88 3.083 ;
      RECT 82.865 2.651 82.87 3.111 ;
      RECT 82.85 2.653 82.865 3.153 ;
      RECT 82.845 2.657 82.85 3.193 ;
      RECT 82.825 2.662 82.845 3.245 ;
      RECT 82.821 2.667 82.825 3.302 ;
      RECT 82.735 2.686 82.821 3.339 ;
      RECT 82.725 2.707 82.735 3.375 ;
      RECT 82.72 2.715 82.725 3.376 ;
      RECT 82.715 2.757 82.72 3.377 ;
      RECT 82.7 2.845 82.715 3.378 ;
      RECT 82.69 2.995 82.7 3.38 ;
      RECT 82.685 3.04 82.69 3.382 ;
      RECT 82.65 3.082 82.685 3.385 ;
      RECT 82.645 3.1 82.65 3.388 ;
      RECT 82.568 3.106 82.645 3.394 ;
      RECT 82.482 3.12 82.568 3.407 ;
      RECT 82.396 3.134 82.482 3.421 ;
      RECT 82.31 3.148 82.396 3.434 ;
      RECT 82.25 3.16 82.31 3.446 ;
      RECT 82.225 3.167 82.25 3.453 ;
      RECT 82.211 3.17 82.225 3.458 ;
      RECT 82.125 3.178 82.211 3.474 ;
      RECT 82.12 3.185 82.125 3.489 ;
      RECT 82.096 3.185 82.12 3.496 ;
      RECT 82.01 3.188 82.096 3.524 ;
      RECT 81.925 3.192 82.01 3.568 ;
      RECT 81.86 3.196 81.925 3.605 ;
      RECT 81.835 3.199 81.86 3.621 ;
      RECT 81.76 3.212 81.835 3.625 ;
      RECT 81.735 3.23 81.76 3.629 ;
      RECT 81.725 3.237 81.735 3.631 ;
      RECT 81.71 3.24 81.725 3.632 ;
      RECT 81.65 3.252 81.71 3.636 ;
      RECT 81.64 3.266 81.65 3.64 ;
      RECT 81.585 3.276 81.64 3.628 ;
      RECT 81.56 3.297 81.585 3.611 ;
      RECT 81.54 3.317 81.56 3.602 ;
      RECT 81.535 3.33 81.54 3.597 ;
      RECT 81.52 3.342 81.535 3.593 ;
      RECT 82.755 1.997 82.76 2.02 ;
      RECT 82.75 1.988 82.755 2.06 ;
      RECT 82.745 1.986 82.75 2.103 ;
      RECT 82.74 1.977 82.745 2.138 ;
      RECT 82.735 1.967 82.74 2.21 ;
      RECT 82.73 1.957 82.735 2.275 ;
      RECT 82.725 1.954 82.73 2.315 ;
      RECT 82.7 1.948 82.725 2.405 ;
      RECT 82.665 1.936 82.7 2.43 ;
      RECT 82.655 1.927 82.665 2.43 ;
      RECT 82.52 1.925 82.53 2.413 ;
      RECT 82.51 1.925 82.52 2.38 ;
      RECT 82.505 1.925 82.51 2.355 ;
      RECT 82.5 1.925 82.505 2.343 ;
      RECT 82.495 1.925 82.5 2.325 ;
      RECT 82.485 1.925 82.495 2.29 ;
      RECT 82.48 1.927 82.485 2.268 ;
      RECT 82.475 1.933 82.48 2.253 ;
      RECT 82.47 1.939 82.475 2.238 ;
      RECT 82.455 1.951 82.47 2.211 ;
      RECT 82.45 1.962 82.455 2.179 ;
      RECT 82.445 1.972 82.45 2.163 ;
      RECT 82.435 1.98 82.445 2.132 ;
      RECT 82.43 1.99 82.435 2.106 ;
      RECT 82.425 2.047 82.43 2.089 ;
      RECT 82.53 1.925 82.655 2.43 ;
      RECT 82.245 2.612 82.505 2.91 ;
      RECT 82.24 2.619 82.505 2.908 ;
      RECT 82.245 2.614 82.52 2.903 ;
      RECT 82.235 2.627 82.52 2.9 ;
      RECT 82.235 2.632 82.525 2.893 ;
      RECT 82.23 2.64 82.525 2.89 ;
      RECT 82.23 2.657 82.53 2.688 ;
      RECT 82.245 2.609 82.476 2.91 ;
      RECT 82.3 2.608 82.476 2.91 ;
      RECT 82.3 2.605 82.39 2.91 ;
      RECT 82.3 2.602 82.386 2.91 ;
      RECT 81.99 2.875 81.995 2.888 ;
      RECT 81.985 2.842 81.99 2.893 ;
      RECT 81.98 2.797 81.985 2.9 ;
      RECT 81.975 2.752 81.98 2.908 ;
      RECT 81.97 2.72 81.975 2.916 ;
      RECT 81.965 2.68 81.97 2.917 ;
      RECT 81.95 2.66 81.965 2.919 ;
      RECT 81.875 2.642 81.95 2.931 ;
      RECT 81.865 2.635 81.875 2.942 ;
      RECT 81.86 2.635 81.865 2.944 ;
      RECT 81.83 2.641 81.86 2.948 ;
      RECT 81.79 2.654 81.83 2.948 ;
      RECT 81.765 2.665 81.79 2.934 ;
      RECT 81.75 2.671 81.765 2.917 ;
      RECT 81.74 2.673 81.75 2.908 ;
      RECT 81.735 2.674 81.74 2.903 ;
      RECT 81.73 2.675 81.735 2.898 ;
      RECT 81.725 2.676 81.73 2.895 ;
      RECT 81.7 2.681 81.725 2.885 ;
      RECT 81.69 2.697 81.7 2.872 ;
      RECT 81.685 2.717 81.69 2.867 ;
      RECT 81.695 2.11 81.7 2.306 ;
      RECT 81.68 2.074 81.695 2.308 ;
      RECT 81.67 2.056 81.68 2.313 ;
      RECT 81.66 2.042 81.67 2.317 ;
      RECT 81.615 2.026 81.66 2.327 ;
      RECT 81.61 2.016 81.615 2.336 ;
      RECT 81.565 2.005 81.61 2.342 ;
      RECT 81.56 1.993 81.565 2.349 ;
      RECT 81.545 1.988 81.56 2.353 ;
      RECT 81.53 1.98 81.545 2.358 ;
      RECT 81.52 1.973 81.53 2.363 ;
      RECT 81.51 1.97 81.52 2.368 ;
      RECT 81.5 1.97 81.51 2.369 ;
      RECT 81.495 1.967 81.5 2.368 ;
      RECT 81.46 1.962 81.485 2.367 ;
      RECT 81.436 1.958 81.46 2.366 ;
      RECT 81.35 1.949 81.436 2.363 ;
      RECT 81.335 1.941 81.35 2.36 ;
      RECT 81.313 1.94 81.335 2.359 ;
      RECT 81.227 1.94 81.313 2.357 ;
      RECT 81.141 1.94 81.227 2.355 ;
      RECT 81.055 1.94 81.141 2.352 ;
      RECT 81.045 1.94 81.055 2.343 ;
      RECT 81.015 1.94 81.045 2.303 ;
      RECT 81.005 1.95 81.015 2.258 ;
      RECT 81 1.99 81.005 2.243 ;
      RECT 80.995 2.005 81 2.23 ;
      RECT 80.965 2.085 80.995 2.192 ;
      RECT 81.485 1.965 81.495 2.368 ;
      RECT 81.31 2.73 81.325 3.335 ;
      RECT 81.315 2.725 81.325 3.335 ;
      RECT 81.48 2.725 81.485 2.908 ;
      RECT 81.47 2.725 81.48 2.938 ;
      RECT 81.455 2.725 81.47 2.998 ;
      RECT 81.45 2.725 81.455 3.043 ;
      RECT 81.445 2.725 81.45 3.073 ;
      RECT 81.44 2.725 81.445 3.093 ;
      RECT 81.43 2.725 81.44 3.128 ;
      RECT 81.415 2.725 81.43 3.16 ;
      RECT 81.37 2.725 81.415 3.188 ;
      RECT 81.365 2.725 81.37 3.218 ;
      RECT 81.36 2.725 81.365 3.23 ;
      RECT 81.355 2.725 81.36 3.238 ;
      RECT 81.345 2.725 81.355 3.253 ;
      RECT 81.34 2.725 81.345 3.275 ;
      RECT 81.33 2.725 81.34 3.298 ;
      RECT 81.325 2.725 81.33 3.318 ;
      RECT 81.29 2.74 81.31 3.335 ;
      RECT 81.265 2.757 81.29 3.335 ;
      RECT 81.26 2.767 81.265 3.335 ;
      RECT 81.23 2.782 81.26 3.335 ;
      RECT 81.155 2.824 81.23 3.335 ;
      RECT 81.15 2.855 81.155 3.318 ;
      RECT 81.145 2.859 81.15 3.3 ;
      RECT 81.14 2.863 81.145 3.263 ;
      RECT 81.135 3.047 81.14 3.23 ;
      RECT 80.62 3.236 80.706 3.801 ;
      RECT 80.575 3.238 80.74 3.795 ;
      RECT 80.706 3.235 80.74 3.795 ;
      RECT 80.62 3.237 80.825 3.789 ;
      RECT 80.575 3.247 80.835 3.785 ;
      RECT 80.55 3.239 80.825 3.781 ;
      RECT 80.545 3.242 80.825 3.776 ;
      RECT 80.52 3.257 80.835 3.77 ;
      RECT 80.52 3.282 80.875 3.765 ;
      RECT 80.48 3.29 80.875 3.74 ;
      RECT 80.48 3.317 80.89 3.738 ;
      RECT 80.48 3.347 80.9 3.725 ;
      RECT 80.475 3.492 80.9 3.713 ;
      RECT 80.48 3.421 80.92 3.71 ;
      RECT 80.48 3.478 80.925 3.518 ;
      RECT 80.67 2.757 80.84 2.935 ;
      RECT 80.62 2.696 80.67 2.92 ;
      RECT 80.355 2.676 80.62 2.905 ;
      RECT 80.315 2.74 80.79 2.905 ;
      RECT 80.315 2.73 80.745 2.905 ;
      RECT 80.315 2.727 80.735 2.905 ;
      RECT 80.315 2.715 80.725 2.905 ;
      RECT 80.315 2.7 80.67 2.905 ;
      RECT 80.355 2.672 80.556 2.905 ;
      RECT 80.365 2.65 80.556 2.905 ;
      RECT 80.39 2.635 80.47 2.905 ;
      RECT 80.145 3.165 80.265 3.61 ;
      RECT 80.13 3.165 80.265 3.609 ;
      RECT 80.085 3.187 80.265 3.604 ;
      RECT 80.045 3.236 80.265 3.598 ;
      RECT 80.045 3.236 80.27 3.573 ;
      RECT 80.045 3.236 80.29 3.463 ;
      RECT 80.04 3.266 80.29 3.46 ;
      RECT 80.13 3.165 80.3 3.355 ;
      RECT 79.79 1.95 79.795 2.395 ;
      RECT 79.6 1.95 79.62 2.36 ;
      RECT 79.57 1.95 79.575 2.335 ;
      RECT 80.25 2.257 80.265 2.445 ;
      RECT 80.245 2.242 80.25 2.451 ;
      RECT 80.225 2.215 80.245 2.454 ;
      RECT 80.175 2.182 80.225 2.463 ;
      RECT 80.145 2.162 80.175 2.467 ;
      RECT 80.126 2.15 80.145 2.463 ;
      RECT 80.04 2.122 80.126 2.453 ;
      RECT 80.03 2.097 80.04 2.443 ;
      RECT 79.96 2.065 80.03 2.435 ;
      RECT 79.935 2.025 79.96 2.427 ;
      RECT 79.915 2.007 79.935 2.421 ;
      RECT 79.905 1.997 79.915 2.418 ;
      RECT 79.895 1.99 79.905 2.416 ;
      RECT 79.875 1.977 79.895 2.413 ;
      RECT 79.865 1.967 79.875 2.41 ;
      RECT 79.855 1.96 79.865 2.408 ;
      RECT 79.805 1.952 79.855 2.402 ;
      RECT 79.795 1.95 79.805 2.396 ;
      RECT 79.765 1.95 79.79 2.393 ;
      RECT 79.736 1.95 79.765 2.388 ;
      RECT 79.65 1.95 79.736 2.378 ;
      RECT 79.62 1.95 79.65 2.365 ;
      RECT 79.575 1.95 79.6 2.348 ;
      RECT 79.56 1.95 79.57 2.33 ;
      RECT 79.54 1.957 79.56 2.315 ;
      RECT 79.535 1.972 79.54 2.303 ;
      RECT 79.53 1.977 79.535 2.243 ;
      RECT 79.525 1.982 79.53 2.085 ;
      RECT 79.52 1.985 79.525 2.003 ;
      RECT 79.785 2.67 79.871 2.991 ;
      RECT 79.785 2.67 79.905 2.984 ;
      RECT 79.735 2.67 79.905 2.98 ;
      RECT 79.735 2.672 79.991 2.978 ;
      RECT 79.735 2.674 80.015 2.972 ;
      RECT 79.735 2.681 80.025 2.971 ;
      RECT 79.735 2.69 80.03 2.968 ;
      RECT 79.735 2.696 80.035 2.963 ;
      RECT 79.735 2.74 80.04 2.96 ;
      RECT 79.735 2.832 80.045 2.957 ;
      RECT 79.26 3.275 79.295 3.595 ;
      RECT 79.845 3.46 79.85 3.642 ;
      RECT 79.8 3.342 79.845 3.661 ;
      RECT 79.785 3.319 79.8 3.684 ;
      RECT 79.775 3.309 79.785 3.694 ;
      RECT 79.755 3.304 79.775 3.707 ;
      RECT 79.73 3.302 79.755 3.728 ;
      RECT 79.711 3.301 79.73 3.74 ;
      RECT 79.625 3.298 79.711 3.74 ;
      RECT 79.555 3.293 79.625 3.728 ;
      RECT 79.48 3.289 79.555 3.703 ;
      RECT 79.415 3.285 79.48 3.67 ;
      RECT 79.345 3.282 79.415 3.63 ;
      RECT 79.315 3.278 79.345 3.605 ;
      RECT 79.295 3.276 79.315 3.598 ;
      RECT 79.211 3.274 79.26 3.596 ;
      RECT 79.125 3.271 79.211 3.597 ;
      RECT 79.05 3.27 79.125 3.599 ;
      RECT 78.965 3.27 79.05 3.625 ;
      RECT 78.888 3.271 78.965 3.65 ;
      RECT 78.802 3.272 78.888 3.65 ;
      RECT 78.716 3.272 78.802 3.65 ;
      RECT 78.63 3.273 78.716 3.65 ;
      RECT 78.61 3.274 78.63 3.642 ;
      RECT 78.595 3.28 78.61 3.627 ;
      RECT 78.56 3.3 78.595 3.607 ;
      RECT 78.55 3.32 78.56 3.589 ;
      RECT 79.52 2.625 79.525 2.895 ;
      RECT 79.515 2.616 79.52 2.9 ;
      RECT 79.505 2.606 79.515 2.912 ;
      RECT 79.5 2.595 79.505 2.923 ;
      RECT 79.48 2.589 79.5 2.941 ;
      RECT 79.435 2.586 79.48 2.99 ;
      RECT 79.42 2.585 79.435 3.035 ;
      RECT 79.415 2.585 79.42 3.048 ;
      RECT 79.405 2.585 79.415 3.06 ;
      RECT 79.4 2.586 79.405 3.075 ;
      RECT 79.38 2.594 79.4 3.08 ;
      RECT 79.35 2.61 79.38 3.08 ;
      RECT 79.34 2.622 79.345 3.08 ;
      RECT 79.305 2.637 79.34 3.08 ;
      RECT 79.275 2.657 79.305 3.08 ;
      RECT 79.265 2.682 79.275 3.08 ;
      RECT 79.26 2.71 79.265 3.08 ;
      RECT 79.255 2.74 79.26 3.08 ;
      RECT 79.25 2.757 79.255 3.08 ;
      RECT 79.24 2.785 79.25 3.08 ;
      RECT 79.23 2.82 79.24 3.08 ;
      RECT 79.225 2.855 79.23 3.08 ;
      RECT 79.345 2.62 79.35 3.08 ;
      RECT 78.86 2.722 79.045 2.895 ;
      RECT 78.82 2.64 79.005 2.893 ;
      RECT 78.781 2.645 79.005 2.889 ;
      RECT 78.695 2.654 79.005 2.884 ;
      RECT 78.611 2.67 79.01 2.879 ;
      RECT 78.525 2.69 79.035 2.873 ;
      RECT 78.525 2.71 79.04 2.873 ;
      RECT 78.611 2.68 79.035 2.879 ;
      RECT 78.695 2.655 79.01 2.884 ;
      RECT 78.86 2.637 79.005 2.895 ;
      RECT 78.86 2.632 78.96 2.895 ;
      RECT 78.946 2.626 78.96 2.895 ;
      RECT 78.335 1.95 78.34 2.349 ;
      RECT 78.08 1.95 78.115 2.347 ;
      RECT 77.675 1.985 77.68 2.341 ;
      RECT 78.42 1.988 78.425 2.243 ;
      RECT 78.415 1.986 78.42 2.249 ;
      RECT 78.41 1.985 78.415 2.256 ;
      RECT 78.385 1.978 78.41 2.28 ;
      RECT 78.38 1.971 78.385 2.304 ;
      RECT 78.375 1.967 78.38 2.313 ;
      RECT 78.365 1.962 78.375 2.326 ;
      RECT 78.36 1.959 78.365 2.335 ;
      RECT 78.355 1.957 78.36 2.34 ;
      RECT 78.34 1.953 78.355 2.35 ;
      RECT 78.325 1.947 78.335 2.349 ;
      RECT 78.287 1.945 78.325 2.349 ;
      RECT 78.201 1.947 78.287 2.349 ;
      RECT 78.115 1.949 78.201 2.348 ;
      RECT 78.044 1.95 78.08 2.347 ;
      RECT 77.958 1.952 78.044 2.347 ;
      RECT 77.872 1.954 77.958 2.346 ;
      RECT 77.786 1.956 77.872 2.346 ;
      RECT 77.7 1.959 77.786 2.345 ;
      RECT 77.69 1.965 77.7 2.344 ;
      RECT 77.68 1.977 77.69 2.342 ;
      RECT 77.62 2.012 77.675 2.338 ;
      RECT 77.615 2.042 77.62 2.1 ;
      RECT 78.36 3.122 78.375 3.315 ;
      RECT 78.355 3.09 78.36 3.315 ;
      RECT 78.345 3.065 78.355 3.315 ;
      RECT 78.34 3.037 78.345 3.315 ;
      RECT 78.31 2.96 78.34 3.315 ;
      RECT 78.285 2.842 78.31 3.315 ;
      RECT 78.28 2.78 78.285 3.315 ;
      RECT 78.27 2.767 78.28 3.315 ;
      RECT 78.25 2.757 78.27 3.315 ;
      RECT 78.235 2.74 78.25 3.315 ;
      RECT 78.205 2.728 78.235 3.315 ;
      RECT 78.2 2.727 78.205 3.26 ;
      RECT 78.195 2.727 78.2 3.218 ;
      RECT 78.18 2.726 78.195 3.17 ;
      RECT 78.165 2.726 78.18 3.108 ;
      RECT 78.145 2.726 78.165 3.068 ;
      RECT 78.14 2.726 78.145 3.053 ;
      RECT 78.115 2.725 78.14 3.048 ;
      RECT 78.045 2.724 78.115 3.035 ;
      RECT 78.03 2.723 78.045 3.02 ;
      RECT 78 2.722 78.03 3.003 ;
      RECT 77.995 2.722 78 2.988 ;
      RECT 77.945 2.721 77.995 2.968 ;
      RECT 77.88 2.72 77.945 2.923 ;
      RECT 77.875 2.72 77.88 2.895 ;
      RECT 77.96 3.257 77.965 3.514 ;
      RECT 77.94 3.176 77.96 3.531 ;
      RECT 77.92 3.17 77.94 3.56 ;
      RECT 77.86 3.157 77.92 3.58 ;
      RECT 77.815 3.141 77.86 3.581 ;
      RECT 77.731 3.129 77.815 3.569 ;
      RECT 77.645 3.116 77.731 3.553 ;
      RECT 77.635 3.109 77.645 3.545 ;
      RECT 77.59 3.106 77.635 3.485 ;
      RECT 77.57 3.102 77.59 3.4 ;
      RECT 77.555 3.1 77.57 3.353 ;
      RECT 77.525 3.097 77.555 3.323 ;
      RECT 77.49 3.093 77.525 3.3 ;
      RECT 77.447 3.088 77.49 3.288 ;
      RECT 77.361 3.079 77.447 3.297 ;
      RECT 77.275 3.068 77.361 3.309 ;
      RECT 77.21 3.059 77.275 3.318 ;
      RECT 77.19 3.05 77.21 3.323 ;
      RECT 77.185 3.043 77.19 3.325 ;
      RECT 77.145 3.028 77.185 3.322 ;
      RECT 77.125 3.007 77.145 3.317 ;
      RECT 77.11 2.995 77.125 3.31 ;
      RECT 77.105 2.987 77.11 3.303 ;
      RECT 77.09 2.967 77.105 3.296 ;
      RECT 77.085 2.83 77.09 3.29 ;
      RECT 77.005 2.719 77.085 3.262 ;
      RECT 76.996 2.712 77.005 3.228 ;
      RECT 76.91 2.706 76.996 3.153 ;
      RECT 76.885 2.697 76.91 3.065 ;
      RECT 76.855 2.692 76.885 3.04 ;
      RECT 76.79 2.701 76.855 3.025 ;
      RECT 76.77 2.717 76.79 3 ;
      RECT 76.76 2.723 76.77 2.948 ;
      RECT 76.74 2.745 76.76 2.83 ;
      RECT 77.395 2.71 77.565 2.895 ;
      RECT 77.395 2.71 77.6 2.893 ;
      RECT 77.445 2.62 77.615 2.884 ;
      RECT 77.395 2.777 77.62 2.877 ;
      RECT 77.41 2.655 77.615 2.884 ;
      RECT 76.61 3.388 76.675 3.831 ;
      RECT 76.55 3.413 76.675 3.829 ;
      RECT 76.55 3.413 76.73 3.823 ;
      RECT 76.535 3.438 76.73 3.822 ;
      RECT 76.675 3.375 76.75 3.819 ;
      RECT 76.61 3.4 76.83 3.813 ;
      RECT 76.535 3.439 76.875 3.807 ;
      RECT 76.52 3.466 76.875 3.798 ;
      RECT 76.535 3.459 76.895 3.79 ;
      RECT 76.52 3.468 76.9 3.773 ;
      RECT 76.515 3.485 76.9 3.6 ;
      RECT 76.52 2.207 76.555 2.445 ;
      RECT 76.52 2.207 76.585 2.444 ;
      RECT 76.52 2.207 76.7 2.44 ;
      RECT 76.52 2.207 76.755 2.418 ;
      RECT 76.53 2.15 76.81 2.318 ;
      RECT 76.635 1.99 76.665 2.441 ;
      RECT 76.665 1.985 76.845 2.198 ;
      RECT 76.535 2.126 76.845 2.198 ;
      RECT 76.585 2.022 76.635 2.442 ;
      RECT 76.555 2.078 76.845 2.198 ;
      RECT 75.425 5.02 75.595 6.49 ;
      RECT 75.425 6.315 75.6 6.485 ;
      RECT 75.055 1.74 75.225 2.93 ;
      RECT 75.055 1.74 75.525 1.91 ;
      RECT 75.055 6.97 75.525 7.14 ;
      RECT 75.055 5.95 75.225 7.14 ;
      RECT 74.065 1.74 74.235 2.93 ;
      RECT 74.065 1.74 74.535 1.91 ;
      RECT 74.065 6.97 74.535 7.14 ;
      RECT 74.065 5.95 74.235 7.14 ;
      RECT 72.215 2.635 72.385 3.865 ;
      RECT 72.27 0.855 72.44 2.805 ;
      RECT 72.215 0.575 72.385 1.025 ;
      RECT 72.215 7.855 72.385 8.305 ;
      RECT 72.27 6.075 72.44 8.025 ;
      RECT 72.215 5.015 72.385 6.245 ;
      RECT 71.695 0.575 71.865 3.865 ;
      RECT 71.695 2.075 72.1 2.405 ;
      RECT 71.695 1.235 72.1 1.565 ;
      RECT 71.695 5.015 71.865 8.305 ;
      RECT 71.695 7.315 72.1 7.645 ;
      RECT 71.695 6.475 72.1 6.805 ;
      RECT 69.795 3.392 69.81 3.443 ;
      RECT 69.79 3.372 69.795 3.49 ;
      RECT 69.775 3.362 69.79 3.558 ;
      RECT 69.75 3.342 69.775 3.613 ;
      RECT 69.71 3.327 69.75 3.633 ;
      RECT 69.665 3.321 69.71 3.661 ;
      RECT 69.595 3.311 69.665 3.678 ;
      RECT 69.575 3.303 69.595 3.678 ;
      RECT 69.515 3.297 69.575 3.67 ;
      RECT 69.456 3.288 69.515 3.658 ;
      RECT 69.37 3.277 69.456 3.641 ;
      RECT 69.348 3.268 69.37 3.629 ;
      RECT 69.262 3.261 69.348 3.616 ;
      RECT 69.176 3.248 69.262 3.597 ;
      RECT 69.09 3.236 69.176 3.577 ;
      RECT 69.06 3.225 69.09 3.564 ;
      RECT 69.01 3.211 69.06 3.556 ;
      RECT 68.99 3.2 69.01 3.548 ;
      RECT 68.941 3.189 68.99 3.54 ;
      RECT 68.855 3.168 68.941 3.525 ;
      RECT 68.81 3.155 68.855 3.51 ;
      RECT 68.765 3.155 68.81 3.49 ;
      RECT 68.71 3.155 68.765 3.425 ;
      RECT 68.685 3.155 68.71 3.348 ;
      RECT 69.21 2.892 69.38 3.075 ;
      RECT 69.21 2.892 69.395 3.033 ;
      RECT 69.21 2.892 69.4 2.975 ;
      RECT 69.27 2.66 69.405 2.951 ;
      RECT 69.27 2.664 69.41 2.934 ;
      RECT 69.215 2.827 69.41 2.934 ;
      RECT 69.24 2.672 69.38 3.075 ;
      RECT 69.24 2.676 69.42 2.875 ;
      RECT 69.225 2.762 69.42 2.875 ;
      RECT 69.235 2.692 69.38 3.075 ;
      RECT 69.235 2.695 69.43 2.788 ;
      RECT 69.23 2.712 69.43 2.788 ;
      RECT 69 1.932 69.17 2.415 ;
      RECT 68.995 1.927 69.145 2.405 ;
      RECT 68.995 1.934 69.175 2.399 ;
      RECT 68.985 1.928 69.145 2.378 ;
      RECT 68.985 1.944 69.19 2.337 ;
      RECT 68.955 1.929 69.145 2.3 ;
      RECT 68.955 1.959 69.2 2.24 ;
      RECT 68.95 1.931 69.145 2.238 ;
      RECT 68.93 1.94 69.175 2.195 ;
      RECT 68.905 1.956 69.19 2.107 ;
      RECT 68.905 1.975 69.215 2.098 ;
      RECT 68.9 2.012 69.215 2.05 ;
      RECT 68.905 1.992 69.22 2.018 ;
      RECT 69 1.926 69.11 2.415 ;
      RECT 69.086 1.925 69.11 2.415 ;
      RECT 68.32 2.71 68.325 2.921 ;
      RECT 68.92 2.71 68.925 2.895 ;
      RECT 68.985 2.75 68.99 2.863 ;
      RECT 68.98 2.742 68.985 2.869 ;
      RECT 68.975 2.732 68.98 2.877 ;
      RECT 68.97 2.722 68.975 2.886 ;
      RECT 68.965 2.712 68.97 2.89 ;
      RECT 68.925 2.71 68.965 2.893 ;
      RECT 68.897 2.709 68.92 2.897 ;
      RECT 68.811 2.706 68.897 2.904 ;
      RECT 68.725 2.702 68.811 2.915 ;
      RECT 68.705 2.7 68.725 2.921 ;
      RECT 68.687 2.699 68.705 2.924 ;
      RECT 68.601 2.697 68.687 2.931 ;
      RECT 68.515 2.692 68.601 2.944 ;
      RECT 68.496 2.689 68.515 2.949 ;
      RECT 68.41 2.687 68.496 2.94 ;
      RECT 68.4 2.687 68.41 2.933 ;
      RECT 68.325 2.7 68.4 2.927 ;
      RECT 68.31 2.711 68.32 2.921 ;
      RECT 68.3 2.713 68.31 2.92 ;
      RECT 68.29 2.717 68.3 2.916 ;
      RECT 68.285 2.72 68.29 2.91 ;
      RECT 68.275 2.722 68.285 2.904 ;
      RECT 68.27 2.725 68.275 2.898 ;
      RECT 68.25 3.311 68.255 3.515 ;
      RECT 68.235 3.298 68.25 3.608 ;
      RECT 68.22 3.279 68.235 3.885 ;
      RECT 68.185 3.245 68.22 3.885 ;
      RECT 68.181 3.215 68.185 3.885 ;
      RECT 68.095 3.097 68.181 3.885 ;
      RECT 68.085 2.972 68.095 3.885 ;
      RECT 68.07 2.94 68.085 3.885 ;
      RECT 68.065 2.915 68.07 3.885 ;
      RECT 68.06 2.905 68.065 3.841 ;
      RECT 68.045 2.877 68.06 3.746 ;
      RECT 68.03 2.843 68.045 3.645 ;
      RECT 68.025 2.821 68.03 3.598 ;
      RECT 68.02 2.81 68.025 3.568 ;
      RECT 68.015 2.8 68.02 3.534 ;
      RECT 68.005 2.787 68.015 3.502 ;
      RECT 67.98 2.763 68.005 3.428 ;
      RECT 67.975 2.743 67.98 3.353 ;
      RECT 67.97 2.737 67.975 3.328 ;
      RECT 67.965 2.732 67.97 3.293 ;
      RECT 67.96 2.727 67.965 3.268 ;
      RECT 67.955 2.725 67.96 3.248 ;
      RECT 67.95 2.725 67.955 3.233 ;
      RECT 67.945 2.725 67.95 3.193 ;
      RECT 67.935 2.725 67.945 3.165 ;
      RECT 67.925 2.725 67.935 3.11 ;
      RECT 67.91 2.725 67.925 3.048 ;
      RECT 67.905 2.724 67.91 2.993 ;
      RECT 67.89 2.723 67.905 2.973 ;
      RECT 67.83 2.721 67.89 2.947 ;
      RECT 67.795 2.722 67.83 2.927 ;
      RECT 67.79 2.724 67.795 2.917 ;
      RECT 67.78 2.743 67.79 2.907 ;
      RECT 67.775 2.77 67.78 2.838 ;
      RECT 67.89 2.195 68.06 2.44 ;
      RECT 67.925 1.966 68.06 2.44 ;
      RECT 67.925 1.968 68.07 2.435 ;
      RECT 67.925 1.97 68.095 2.423 ;
      RECT 67.925 1.973 68.12 2.405 ;
      RECT 67.925 1.978 68.17 2.378 ;
      RECT 67.925 1.983 68.19 2.343 ;
      RECT 67.905 1.985 68.2 2.318 ;
      RECT 67.895 2.08 68.2 2.318 ;
      RECT 67.925 1.965 68.035 2.44 ;
      RECT 67.935 1.962 68.03 2.44 ;
      RECT 67.455 3.227 67.645 3.585 ;
      RECT 67.455 3.239 67.68 3.584 ;
      RECT 67.455 3.267 67.7 3.582 ;
      RECT 67.455 3.292 67.705 3.581 ;
      RECT 67.455 3.35 67.72 3.58 ;
      RECT 67.44 3.223 67.6 3.565 ;
      RECT 67.42 3.232 67.645 3.518 ;
      RECT 67.395 3.243 67.68 3.455 ;
      RECT 67.395 3.327 67.715 3.455 ;
      RECT 67.395 3.302 67.71 3.455 ;
      RECT 67.455 3.218 67.6 3.585 ;
      RECT 67.541 3.217 67.6 3.585 ;
      RECT 67.541 3.216 67.585 3.585 ;
      RECT 67.455 7.855 67.625 8.305 ;
      RECT 67.51 6.075 67.68 8.025 ;
      RECT 67.455 5.015 67.625 6.245 ;
      RECT 66.935 5.015 67.105 8.305 ;
      RECT 66.935 7.315 67.34 7.645 ;
      RECT 66.935 6.475 67.34 6.805 ;
      RECT 67.24 2.732 67.245 3.11 ;
      RECT 67.235 2.7 67.24 3.11 ;
      RECT 67.23 2.672 67.235 3.11 ;
      RECT 67.225 2.652 67.23 3.11 ;
      RECT 67.17 2.635 67.225 3.11 ;
      RECT 67.13 2.62 67.17 3.11 ;
      RECT 67.075 2.607 67.13 3.11 ;
      RECT 67.04 2.598 67.075 3.11 ;
      RECT 67.036 2.596 67.04 3.109 ;
      RECT 66.95 2.592 67.036 3.092 ;
      RECT 66.865 2.584 66.95 3.055 ;
      RECT 66.855 2.58 66.865 3.028 ;
      RECT 66.845 2.58 66.855 3.01 ;
      RECT 66.835 2.582 66.845 2.993 ;
      RECT 66.83 2.587 66.835 2.979 ;
      RECT 66.825 2.591 66.83 2.966 ;
      RECT 66.815 2.596 66.825 2.95 ;
      RECT 66.8 2.61 66.815 2.925 ;
      RECT 66.795 2.616 66.8 2.905 ;
      RECT 66.79 2.618 66.795 2.898 ;
      RECT 66.785 2.622 66.79 2.773 ;
      RECT 66.965 3.422 67.21 3.885 ;
      RECT 66.885 3.395 67.205 3.881 ;
      RECT 66.815 3.43 67.21 3.874 ;
      RECT 66.605 3.685 67.21 3.87 ;
      RECT 66.785 3.453 67.21 3.87 ;
      RECT 66.625 3.645 67.21 3.87 ;
      RECT 66.775 3.465 67.21 3.87 ;
      RECT 66.66 3.582 67.21 3.87 ;
      RECT 66.715 3.507 67.21 3.87 ;
      RECT 66.965 3.372 67.205 3.885 ;
      RECT 66.995 3.365 67.205 3.885 ;
      RECT 66.985 3.367 67.205 3.885 ;
      RECT 66.995 3.362 67.125 3.885 ;
      RECT 66.55 1.925 66.636 2.364 ;
      RECT 66.545 1.925 66.636 2.362 ;
      RECT 66.545 1.925 66.705 2.361 ;
      RECT 66.545 1.925 66.735 2.358 ;
      RECT 66.53 1.932 66.735 2.349 ;
      RECT 66.53 1.932 66.74 2.345 ;
      RECT 66.525 1.942 66.74 2.338 ;
      RECT 66.52 1.947 66.74 2.313 ;
      RECT 66.52 1.947 66.755 2.295 ;
      RECT 66.545 1.925 66.775 2.21 ;
      RECT 66.515 1.952 66.775 2.208 ;
      RECT 66.525 1.945 66.78 2.146 ;
      RECT 66.515 2.067 66.785 2.129 ;
      RECT 66.5 1.962 66.78 2.08 ;
      RECT 66.495 1.972 66.78 1.98 ;
      RECT 66.575 2.743 66.58 2.82 ;
      RECT 66.565 2.737 66.575 3.01 ;
      RECT 66.555 2.729 66.565 3.031 ;
      RECT 66.545 2.72 66.555 3.053 ;
      RECT 66.54 2.715 66.545 3.07 ;
      RECT 66.5 2.715 66.54 3.11 ;
      RECT 66.48 2.715 66.5 3.165 ;
      RECT 66.475 2.715 66.48 3.193 ;
      RECT 66.465 2.715 66.475 3.208 ;
      RECT 66.43 2.715 66.465 3.25 ;
      RECT 66.425 2.715 66.43 3.293 ;
      RECT 66.415 2.715 66.425 3.308 ;
      RECT 66.4 2.715 66.415 3.328 ;
      RECT 66.385 2.715 66.4 3.355 ;
      RECT 66.38 2.716 66.385 3.373 ;
      RECT 66.36 2.717 66.38 3.38 ;
      RECT 66.305 2.718 66.36 3.4 ;
      RECT 66.295 2.719 66.305 3.414 ;
      RECT 66.29 2.722 66.295 3.413 ;
      RECT 66.25 2.795 66.29 3.411 ;
      RECT 66.235 2.875 66.25 3.409 ;
      RECT 66.21 2.93 66.235 3.407 ;
      RECT 66.195 2.995 66.21 3.406 ;
      RECT 66.15 3.027 66.195 3.403 ;
      RECT 66.065 3.05 66.15 3.398 ;
      RECT 66.04 3.07 66.065 3.393 ;
      RECT 65.97 3.075 66.04 3.389 ;
      RECT 65.95 3.077 65.97 3.386 ;
      RECT 65.865 3.088 65.95 3.38 ;
      RECT 65.86 3.099 65.865 3.375 ;
      RECT 65.85 3.101 65.86 3.375 ;
      RECT 65.815 3.105 65.85 3.373 ;
      RECT 65.765 3.115 65.815 3.36 ;
      RECT 65.745 3.123 65.765 3.345 ;
      RECT 65.665 3.135 65.745 3.328 ;
      RECT 65.83 2.685 66 2.895 ;
      RECT 65.946 2.681 66 2.895 ;
      RECT 65.751 2.685 66 2.886 ;
      RECT 65.751 2.685 66.005 2.875 ;
      RECT 65.665 2.685 66.005 2.866 ;
      RECT 65.665 2.693 66.015 2.81 ;
      RECT 65.665 2.705 66.02 2.723 ;
      RECT 65.665 2.712 66.025 2.715 ;
      RECT 65.86 2.683 66 2.895 ;
      RECT 65.615 3.628 65.86 3.96 ;
      RECT 65.61 3.62 65.615 3.957 ;
      RECT 65.58 3.64 65.86 3.938 ;
      RECT 65.56 3.672 65.86 3.911 ;
      RECT 65.61 3.625 65.787 3.957 ;
      RECT 65.61 3.622 65.701 3.957 ;
      RECT 65.55 1.97 65.72 2.39 ;
      RECT 65.545 1.97 65.72 2.388 ;
      RECT 65.545 1.97 65.745 2.378 ;
      RECT 65.545 1.97 65.765 2.353 ;
      RECT 65.54 1.97 65.765 2.348 ;
      RECT 65.54 1.97 65.775 2.338 ;
      RECT 65.54 1.97 65.78 2.333 ;
      RECT 65.54 1.975 65.785 2.328 ;
      RECT 65.54 2.007 65.8 2.318 ;
      RECT 65.54 2.077 65.825 2.301 ;
      RECT 65.52 2.077 65.825 2.293 ;
      RECT 65.52 2.137 65.835 2.27 ;
      RECT 65.52 2.177 65.845 2.215 ;
      RECT 65.505 1.97 65.78 2.195 ;
      RECT 65.495 1.985 65.785 2.093 ;
      RECT 65.085 3.375 65.255 3.9 ;
      RECT 65.08 3.375 65.255 3.893 ;
      RECT 65.07 3.375 65.26 3.858 ;
      RECT 65.065 3.385 65.26 3.83 ;
      RECT 65.06 3.405 65.26 3.813 ;
      RECT 65.07 3.38 65.265 3.803 ;
      RECT 65.055 3.425 65.265 3.795 ;
      RECT 65.05 3.445 65.265 3.78 ;
      RECT 65.045 3.475 65.265 3.77 ;
      RECT 65.035 3.52 65.265 3.745 ;
      RECT 65.065 3.39 65.27 3.728 ;
      RECT 65.03 3.572 65.27 3.723 ;
      RECT 65.065 3.4 65.275 3.693 ;
      RECT 65.025 3.605 65.275 3.69 ;
      RECT 65.02 3.63 65.275 3.67 ;
      RECT 65.06 3.417 65.285 3.61 ;
      RECT 65.055 3.439 65.295 3.503 ;
      RECT 65.005 2.686 65.02 2.955 ;
      RECT 64.96 2.67 65.005 3 ;
      RECT 64.955 2.658 64.96 3.05 ;
      RECT 64.945 2.654 64.955 3.083 ;
      RECT 64.94 2.651 64.945 3.111 ;
      RECT 64.925 2.653 64.94 3.153 ;
      RECT 64.92 2.657 64.925 3.193 ;
      RECT 64.9 2.662 64.92 3.245 ;
      RECT 64.896 2.667 64.9 3.302 ;
      RECT 64.81 2.686 64.896 3.339 ;
      RECT 64.8 2.707 64.81 3.375 ;
      RECT 64.795 2.715 64.8 3.376 ;
      RECT 64.79 2.757 64.795 3.377 ;
      RECT 64.775 2.845 64.79 3.378 ;
      RECT 64.765 2.995 64.775 3.38 ;
      RECT 64.76 3.04 64.765 3.382 ;
      RECT 64.725 3.082 64.76 3.385 ;
      RECT 64.72 3.1 64.725 3.388 ;
      RECT 64.643 3.106 64.72 3.394 ;
      RECT 64.557 3.12 64.643 3.407 ;
      RECT 64.471 3.134 64.557 3.421 ;
      RECT 64.385 3.148 64.471 3.434 ;
      RECT 64.325 3.16 64.385 3.446 ;
      RECT 64.3 3.167 64.325 3.453 ;
      RECT 64.286 3.17 64.3 3.458 ;
      RECT 64.2 3.178 64.286 3.474 ;
      RECT 64.195 3.185 64.2 3.489 ;
      RECT 64.171 3.185 64.195 3.496 ;
      RECT 64.085 3.188 64.171 3.524 ;
      RECT 64 3.192 64.085 3.568 ;
      RECT 63.935 3.196 64 3.605 ;
      RECT 63.91 3.199 63.935 3.621 ;
      RECT 63.835 3.212 63.91 3.625 ;
      RECT 63.81 3.23 63.835 3.629 ;
      RECT 63.8 3.237 63.81 3.631 ;
      RECT 63.785 3.24 63.8 3.632 ;
      RECT 63.725 3.252 63.785 3.636 ;
      RECT 63.715 3.266 63.725 3.64 ;
      RECT 63.66 3.276 63.715 3.628 ;
      RECT 63.635 3.297 63.66 3.611 ;
      RECT 63.615 3.317 63.635 3.602 ;
      RECT 63.61 3.33 63.615 3.597 ;
      RECT 63.595 3.342 63.61 3.593 ;
      RECT 64.83 1.997 64.835 2.02 ;
      RECT 64.825 1.988 64.83 2.06 ;
      RECT 64.82 1.986 64.825 2.103 ;
      RECT 64.815 1.977 64.82 2.138 ;
      RECT 64.81 1.967 64.815 2.21 ;
      RECT 64.805 1.957 64.81 2.275 ;
      RECT 64.8 1.954 64.805 2.315 ;
      RECT 64.775 1.948 64.8 2.405 ;
      RECT 64.74 1.936 64.775 2.43 ;
      RECT 64.73 1.927 64.74 2.43 ;
      RECT 64.595 1.925 64.605 2.413 ;
      RECT 64.585 1.925 64.595 2.38 ;
      RECT 64.58 1.925 64.585 2.355 ;
      RECT 64.575 1.925 64.58 2.343 ;
      RECT 64.57 1.925 64.575 2.325 ;
      RECT 64.56 1.925 64.57 2.29 ;
      RECT 64.555 1.927 64.56 2.268 ;
      RECT 64.55 1.933 64.555 2.253 ;
      RECT 64.545 1.939 64.55 2.238 ;
      RECT 64.53 1.951 64.545 2.211 ;
      RECT 64.525 1.962 64.53 2.179 ;
      RECT 64.52 1.972 64.525 2.163 ;
      RECT 64.51 1.98 64.52 2.132 ;
      RECT 64.505 1.99 64.51 2.106 ;
      RECT 64.5 2.047 64.505 2.089 ;
      RECT 64.605 1.925 64.73 2.43 ;
      RECT 64.32 2.612 64.58 2.91 ;
      RECT 64.315 2.619 64.58 2.908 ;
      RECT 64.32 2.614 64.595 2.903 ;
      RECT 64.31 2.627 64.595 2.9 ;
      RECT 64.31 2.632 64.6 2.893 ;
      RECT 64.305 2.64 64.6 2.89 ;
      RECT 64.305 2.657 64.605 2.688 ;
      RECT 64.32 2.609 64.551 2.91 ;
      RECT 64.375 2.608 64.551 2.91 ;
      RECT 64.375 2.605 64.465 2.91 ;
      RECT 64.375 2.602 64.461 2.91 ;
      RECT 64.065 2.875 64.07 2.888 ;
      RECT 64.06 2.842 64.065 2.893 ;
      RECT 64.055 2.797 64.06 2.9 ;
      RECT 64.05 2.752 64.055 2.908 ;
      RECT 64.045 2.72 64.05 2.916 ;
      RECT 64.04 2.68 64.045 2.917 ;
      RECT 64.025 2.66 64.04 2.919 ;
      RECT 63.95 2.642 64.025 2.931 ;
      RECT 63.94 2.635 63.95 2.942 ;
      RECT 63.935 2.635 63.94 2.944 ;
      RECT 63.905 2.641 63.935 2.948 ;
      RECT 63.865 2.654 63.905 2.948 ;
      RECT 63.84 2.665 63.865 2.934 ;
      RECT 63.825 2.671 63.84 2.917 ;
      RECT 63.815 2.673 63.825 2.908 ;
      RECT 63.81 2.674 63.815 2.903 ;
      RECT 63.805 2.675 63.81 2.898 ;
      RECT 63.8 2.676 63.805 2.895 ;
      RECT 63.775 2.681 63.8 2.885 ;
      RECT 63.765 2.697 63.775 2.872 ;
      RECT 63.76 2.717 63.765 2.867 ;
      RECT 63.77 2.11 63.775 2.306 ;
      RECT 63.755 2.074 63.77 2.308 ;
      RECT 63.745 2.056 63.755 2.313 ;
      RECT 63.735 2.042 63.745 2.317 ;
      RECT 63.69 2.026 63.735 2.327 ;
      RECT 63.685 2.016 63.69 2.336 ;
      RECT 63.64 2.005 63.685 2.342 ;
      RECT 63.635 1.993 63.64 2.349 ;
      RECT 63.62 1.988 63.635 2.353 ;
      RECT 63.605 1.98 63.62 2.358 ;
      RECT 63.595 1.973 63.605 2.363 ;
      RECT 63.585 1.97 63.595 2.368 ;
      RECT 63.575 1.97 63.585 2.369 ;
      RECT 63.57 1.967 63.575 2.368 ;
      RECT 63.535 1.962 63.56 2.367 ;
      RECT 63.511 1.958 63.535 2.366 ;
      RECT 63.425 1.949 63.511 2.363 ;
      RECT 63.41 1.941 63.425 2.36 ;
      RECT 63.388 1.94 63.41 2.359 ;
      RECT 63.302 1.94 63.388 2.357 ;
      RECT 63.216 1.94 63.302 2.355 ;
      RECT 63.13 1.94 63.216 2.352 ;
      RECT 63.12 1.94 63.13 2.343 ;
      RECT 63.09 1.94 63.12 2.303 ;
      RECT 63.08 1.95 63.09 2.258 ;
      RECT 63.075 1.99 63.08 2.243 ;
      RECT 63.07 2.005 63.075 2.23 ;
      RECT 63.04 2.085 63.07 2.192 ;
      RECT 63.56 1.965 63.57 2.368 ;
      RECT 63.385 2.73 63.4 3.335 ;
      RECT 63.39 2.725 63.4 3.335 ;
      RECT 63.555 2.725 63.56 2.908 ;
      RECT 63.545 2.725 63.555 2.938 ;
      RECT 63.53 2.725 63.545 2.998 ;
      RECT 63.525 2.725 63.53 3.043 ;
      RECT 63.52 2.725 63.525 3.073 ;
      RECT 63.515 2.725 63.52 3.093 ;
      RECT 63.505 2.725 63.515 3.128 ;
      RECT 63.49 2.725 63.505 3.16 ;
      RECT 63.445 2.725 63.49 3.188 ;
      RECT 63.44 2.725 63.445 3.218 ;
      RECT 63.435 2.725 63.44 3.23 ;
      RECT 63.43 2.725 63.435 3.238 ;
      RECT 63.42 2.725 63.43 3.253 ;
      RECT 63.415 2.725 63.42 3.275 ;
      RECT 63.405 2.725 63.415 3.298 ;
      RECT 63.4 2.725 63.405 3.318 ;
      RECT 63.365 2.74 63.385 3.335 ;
      RECT 63.34 2.757 63.365 3.335 ;
      RECT 63.335 2.767 63.34 3.335 ;
      RECT 63.305 2.782 63.335 3.335 ;
      RECT 63.23 2.824 63.305 3.335 ;
      RECT 63.225 2.855 63.23 3.318 ;
      RECT 63.22 2.859 63.225 3.3 ;
      RECT 63.215 2.863 63.22 3.263 ;
      RECT 63.21 3.047 63.215 3.23 ;
      RECT 62.695 3.236 62.781 3.801 ;
      RECT 62.65 3.238 62.815 3.795 ;
      RECT 62.781 3.235 62.815 3.795 ;
      RECT 62.695 3.237 62.9 3.789 ;
      RECT 62.65 3.247 62.91 3.785 ;
      RECT 62.625 3.239 62.9 3.781 ;
      RECT 62.62 3.242 62.9 3.776 ;
      RECT 62.595 3.257 62.91 3.77 ;
      RECT 62.595 3.282 62.95 3.765 ;
      RECT 62.555 3.29 62.95 3.74 ;
      RECT 62.555 3.317 62.965 3.738 ;
      RECT 62.555 3.347 62.975 3.725 ;
      RECT 62.55 3.492 62.975 3.713 ;
      RECT 62.555 3.421 62.995 3.71 ;
      RECT 62.555 3.478 63 3.518 ;
      RECT 62.745 2.757 62.915 2.935 ;
      RECT 62.695 2.696 62.745 2.92 ;
      RECT 62.43 2.676 62.695 2.905 ;
      RECT 62.39 2.74 62.865 2.905 ;
      RECT 62.39 2.73 62.82 2.905 ;
      RECT 62.39 2.727 62.81 2.905 ;
      RECT 62.39 2.715 62.8 2.905 ;
      RECT 62.39 2.7 62.745 2.905 ;
      RECT 62.43 2.672 62.631 2.905 ;
      RECT 62.44 2.65 62.631 2.905 ;
      RECT 62.465 2.635 62.545 2.905 ;
      RECT 62.22 3.165 62.34 3.61 ;
      RECT 62.205 3.165 62.34 3.609 ;
      RECT 62.16 3.187 62.34 3.604 ;
      RECT 62.12 3.236 62.34 3.598 ;
      RECT 62.12 3.236 62.345 3.573 ;
      RECT 62.12 3.236 62.365 3.463 ;
      RECT 62.115 3.266 62.365 3.46 ;
      RECT 62.205 3.165 62.375 3.355 ;
      RECT 61.865 1.95 61.87 2.395 ;
      RECT 61.675 1.95 61.695 2.36 ;
      RECT 61.645 1.95 61.65 2.335 ;
      RECT 62.325 2.257 62.34 2.445 ;
      RECT 62.32 2.242 62.325 2.451 ;
      RECT 62.3 2.215 62.32 2.454 ;
      RECT 62.25 2.182 62.3 2.463 ;
      RECT 62.22 2.162 62.25 2.467 ;
      RECT 62.201 2.15 62.22 2.463 ;
      RECT 62.115 2.122 62.201 2.453 ;
      RECT 62.105 2.097 62.115 2.443 ;
      RECT 62.035 2.065 62.105 2.435 ;
      RECT 62.01 2.025 62.035 2.427 ;
      RECT 61.99 2.007 62.01 2.421 ;
      RECT 61.98 1.997 61.99 2.418 ;
      RECT 61.97 1.99 61.98 2.416 ;
      RECT 61.95 1.977 61.97 2.413 ;
      RECT 61.94 1.967 61.95 2.41 ;
      RECT 61.93 1.96 61.94 2.408 ;
      RECT 61.88 1.952 61.93 2.402 ;
      RECT 61.87 1.95 61.88 2.396 ;
      RECT 61.84 1.95 61.865 2.393 ;
      RECT 61.811 1.95 61.84 2.388 ;
      RECT 61.725 1.95 61.811 2.378 ;
      RECT 61.695 1.95 61.725 2.365 ;
      RECT 61.65 1.95 61.675 2.348 ;
      RECT 61.635 1.95 61.645 2.33 ;
      RECT 61.615 1.957 61.635 2.315 ;
      RECT 61.61 1.972 61.615 2.303 ;
      RECT 61.605 1.977 61.61 2.243 ;
      RECT 61.6 1.982 61.605 2.085 ;
      RECT 61.595 1.985 61.6 2.003 ;
      RECT 61.86 2.67 61.946 2.991 ;
      RECT 61.86 2.67 61.98 2.984 ;
      RECT 61.81 2.67 61.98 2.98 ;
      RECT 61.81 2.672 62.066 2.978 ;
      RECT 61.81 2.674 62.09 2.972 ;
      RECT 61.81 2.681 62.1 2.971 ;
      RECT 61.81 2.69 62.105 2.968 ;
      RECT 61.81 2.696 62.11 2.963 ;
      RECT 61.81 2.74 62.115 2.96 ;
      RECT 61.81 2.832 62.12 2.957 ;
      RECT 61.335 3.275 61.37 3.595 ;
      RECT 61.92 3.46 61.925 3.642 ;
      RECT 61.875 3.342 61.92 3.661 ;
      RECT 61.86 3.319 61.875 3.684 ;
      RECT 61.85 3.309 61.86 3.694 ;
      RECT 61.83 3.304 61.85 3.707 ;
      RECT 61.805 3.302 61.83 3.728 ;
      RECT 61.786 3.301 61.805 3.74 ;
      RECT 61.7 3.298 61.786 3.74 ;
      RECT 61.63 3.293 61.7 3.728 ;
      RECT 61.555 3.289 61.63 3.703 ;
      RECT 61.49 3.285 61.555 3.67 ;
      RECT 61.42 3.282 61.49 3.63 ;
      RECT 61.39 3.278 61.42 3.605 ;
      RECT 61.37 3.276 61.39 3.598 ;
      RECT 61.286 3.274 61.335 3.596 ;
      RECT 61.2 3.271 61.286 3.597 ;
      RECT 61.125 3.27 61.2 3.599 ;
      RECT 61.04 3.27 61.125 3.625 ;
      RECT 60.963 3.271 61.04 3.65 ;
      RECT 60.877 3.272 60.963 3.65 ;
      RECT 60.791 3.272 60.877 3.65 ;
      RECT 60.705 3.273 60.791 3.65 ;
      RECT 60.685 3.274 60.705 3.642 ;
      RECT 60.67 3.28 60.685 3.627 ;
      RECT 60.635 3.3 60.67 3.607 ;
      RECT 60.625 3.32 60.635 3.589 ;
      RECT 61.595 2.625 61.6 2.895 ;
      RECT 61.59 2.616 61.595 2.9 ;
      RECT 61.58 2.606 61.59 2.912 ;
      RECT 61.575 2.595 61.58 2.923 ;
      RECT 61.555 2.589 61.575 2.941 ;
      RECT 61.51 2.586 61.555 2.99 ;
      RECT 61.495 2.585 61.51 3.035 ;
      RECT 61.49 2.585 61.495 3.048 ;
      RECT 61.48 2.585 61.49 3.06 ;
      RECT 61.475 2.586 61.48 3.075 ;
      RECT 61.455 2.594 61.475 3.08 ;
      RECT 61.425 2.61 61.455 3.08 ;
      RECT 61.415 2.622 61.42 3.08 ;
      RECT 61.38 2.637 61.415 3.08 ;
      RECT 61.35 2.657 61.38 3.08 ;
      RECT 61.34 2.682 61.35 3.08 ;
      RECT 61.335 2.71 61.34 3.08 ;
      RECT 61.33 2.74 61.335 3.08 ;
      RECT 61.325 2.757 61.33 3.08 ;
      RECT 61.315 2.785 61.325 3.08 ;
      RECT 61.305 2.82 61.315 3.08 ;
      RECT 61.3 2.855 61.305 3.08 ;
      RECT 61.42 2.62 61.425 3.08 ;
      RECT 60.935 2.722 61.12 2.895 ;
      RECT 60.895 2.64 61.08 2.893 ;
      RECT 60.856 2.645 61.08 2.889 ;
      RECT 60.77 2.654 61.08 2.884 ;
      RECT 60.686 2.67 61.085 2.879 ;
      RECT 60.6 2.69 61.11 2.873 ;
      RECT 60.6 2.71 61.115 2.873 ;
      RECT 60.686 2.68 61.11 2.879 ;
      RECT 60.77 2.655 61.085 2.884 ;
      RECT 60.935 2.637 61.08 2.895 ;
      RECT 60.935 2.632 61.035 2.895 ;
      RECT 61.021 2.626 61.035 2.895 ;
      RECT 60.41 1.95 60.415 2.349 ;
      RECT 60.155 1.95 60.19 2.347 ;
      RECT 59.75 1.985 59.755 2.341 ;
      RECT 60.495 1.988 60.5 2.243 ;
      RECT 60.49 1.986 60.495 2.249 ;
      RECT 60.485 1.985 60.49 2.256 ;
      RECT 60.46 1.978 60.485 2.28 ;
      RECT 60.455 1.971 60.46 2.304 ;
      RECT 60.45 1.967 60.455 2.313 ;
      RECT 60.44 1.962 60.45 2.326 ;
      RECT 60.435 1.959 60.44 2.335 ;
      RECT 60.43 1.957 60.435 2.34 ;
      RECT 60.415 1.953 60.43 2.35 ;
      RECT 60.4 1.947 60.41 2.349 ;
      RECT 60.362 1.945 60.4 2.349 ;
      RECT 60.276 1.947 60.362 2.349 ;
      RECT 60.19 1.949 60.276 2.348 ;
      RECT 60.119 1.95 60.155 2.347 ;
      RECT 60.033 1.952 60.119 2.347 ;
      RECT 59.947 1.954 60.033 2.346 ;
      RECT 59.861 1.956 59.947 2.346 ;
      RECT 59.775 1.959 59.861 2.345 ;
      RECT 59.765 1.965 59.775 2.344 ;
      RECT 59.755 1.977 59.765 2.342 ;
      RECT 59.695 2.012 59.75 2.338 ;
      RECT 59.69 2.042 59.695 2.1 ;
      RECT 60.435 3.122 60.45 3.315 ;
      RECT 60.43 3.09 60.435 3.315 ;
      RECT 60.42 3.065 60.43 3.315 ;
      RECT 60.415 3.037 60.42 3.315 ;
      RECT 60.385 2.96 60.415 3.315 ;
      RECT 60.36 2.842 60.385 3.315 ;
      RECT 60.355 2.78 60.36 3.315 ;
      RECT 60.345 2.767 60.355 3.315 ;
      RECT 60.325 2.757 60.345 3.315 ;
      RECT 60.31 2.74 60.325 3.315 ;
      RECT 60.28 2.728 60.31 3.315 ;
      RECT 60.275 2.727 60.28 3.26 ;
      RECT 60.27 2.727 60.275 3.218 ;
      RECT 60.255 2.726 60.27 3.17 ;
      RECT 60.24 2.726 60.255 3.108 ;
      RECT 60.22 2.726 60.24 3.068 ;
      RECT 60.215 2.726 60.22 3.053 ;
      RECT 60.19 2.725 60.215 3.048 ;
      RECT 60.12 2.724 60.19 3.035 ;
      RECT 60.105 2.723 60.12 3.02 ;
      RECT 60.075 2.722 60.105 3.003 ;
      RECT 60.07 2.722 60.075 2.988 ;
      RECT 60.02 2.721 60.07 2.968 ;
      RECT 59.955 2.72 60.02 2.923 ;
      RECT 59.95 2.72 59.955 2.895 ;
      RECT 60.035 3.257 60.04 3.514 ;
      RECT 60.015 3.176 60.035 3.531 ;
      RECT 59.995 3.17 60.015 3.56 ;
      RECT 59.935 3.157 59.995 3.58 ;
      RECT 59.89 3.141 59.935 3.581 ;
      RECT 59.806 3.129 59.89 3.569 ;
      RECT 59.72 3.116 59.806 3.553 ;
      RECT 59.71 3.109 59.72 3.545 ;
      RECT 59.665 3.106 59.71 3.485 ;
      RECT 59.645 3.102 59.665 3.4 ;
      RECT 59.63 3.1 59.645 3.353 ;
      RECT 59.6 3.097 59.63 3.323 ;
      RECT 59.565 3.093 59.6 3.3 ;
      RECT 59.522 3.088 59.565 3.288 ;
      RECT 59.436 3.079 59.522 3.297 ;
      RECT 59.35 3.068 59.436 3.309 ;
      RECT 59.285 3.059 59.35 3.318 ;
      RECT 59.265 3.05 59.285 3.323 ;
      RECT 59.26 3.043 59.265 3.325 ;
      RECT 59.22 3.028 59.26 3.322 ;
      RECT 59.2 3.007 59.22 3.317 ;
      RECT 59.185 2.995 59.2 3.31 ;
      RECT 59.18 2.987 59.185 3.303 ;
      RECT 59.165 2.967 59.18 3.296 ;
      RECT 59.16 2.83 59.165 3.29 ;
      RECT 59.08 2.719 59.16 3.262 ;
      RECT 59.071 2.712 59.08 3.228 ;
      RECT 58.985 2.706 59.071 3.153 ;
      RECT 58.96 2.697 58.985 3.065 ;
      RECT 58.93 2.692 58.96 3.04 ;
      RECT 58.865 2.701 58.93 3.025 ;
      RECT 58.845 2.717 58.865 3 ;
      RECT 58.835 2.723 58.845 2.948 ;
      RECT 58.815 2.745 58.835 2.83 ;
      RECT 59.47 2.71 59.64 2.895 ;
      RECT 59.47 2.71 59.675 2.893 ;
      RECT 59.52 2.62 59.69 2.884 ;
      RECT 59.47 2.777 59.695 2.877 ;
      RECT 59.485 2.655 59.69 2.884 ;
      RECT 58.685 3.388 58.75 3.831 ;
      RECT 58.625 3.413 58.75 3.829 ;
      RECT 58.625 3.413 58.805 3.823 ;
      RECT 58.61 3.438 58.805 3.822 ;
      RECT 58.75 3.375 58.825 3.819 ;
      RECT 58.685 3.4 58.905 3.813 ;
      RECT 58.61 3.439 58.95 3.807 ;
      RECT 58.595 3.466 58.95 3.798 ;
      RECT 58.61 3.459 58.97 3.79 ;
      RECT 58.595 3.468 58.975 3.773 ;
      RECT 58.59 3.485 58.975 3.6 ;
      RECT 58.595 2.207 58.63 2.445 ;
      RECT 58.595 2.207 58.66 2.444 ;
      RECT 58.595 2.207 58.775 2.44 ;
      RECT 58.595 2.207 58.83 2.418 ;
      RECT 58.605 2.15 58.885 2.318 ;
      RECT 58.71 1.99 58.74 2.441 ;
      RECT 58.74 1.985 58.92 2.198 ;
      RECT 58.61 2.126 58.92 2.198 ;
      RECT 58.66 2.022 58.71 2.442 ;
      RECT 58.63 2.078 58.92 2.198 ;
      RECT 57.5 5.02 57.67 6.49 ;
      RECT 57.5 6.315 57.675 6.485 ;
      RECT 57.13 1.74 57.3 2.93 ;
      RECT 57.13 1.74 57.6 1.91 ;
      RECT 57.13 6.97 57.6 7.14 ;
      RECT 57.13 5.95 57.3 7.14 ;
      RECT 56.14 1.74 56.31 2.93 ;
      RECT 56.14 1.74 56.61 1.91 ;
      RECT 56.14 6.97 56.61 7.14 ;
      RECT 56.14 5.95 56.31 7.14 ;
      RECT 54.29 2.635 54.46 3.865 ;
      RECT 54.345 0.855 54.515 2.805 ;
      RECT 54.29 0.575 54.46 1.025 ;
      RECT 54.29 7.855 54.46 8.305 ;
      RECT 54.345 6.075 54.515 8.025 ;
      RECT 54.29 5.015 54.46 6.245 ;
      RECT 53.77 0.575 53.94 3.865 ;
      RECT 53.77 2.075 54.175 2.405 ;
      RECT 53.77 1.235 54.175 1.565 ;
      RECT 53.77 5.015 53.94 8.305 ;
      RECT 53.77 7.315 54.175 7.645 ;
      RECT 53.77 6.475 54.175 6.805 ;
      RECT 51.87 3.392 51.885 3.443 ;
      RECT 51.865 3.372 51.87 3.49 ;
      RECT 51.85 3.362 51.865 3.558 ;
      RECT 51.825 3.342 51.85 3.613 ;
      RECT 51.785 3.327 51.825 3.633 ;
      RECT 51.74 3.321 51.785 3.661 ;
      RECT 51.67 3.311 51.74 3.678 ;
      RECT 51.65 3.303 51.67 3.678 ;
      RECT 51.59 3.297 51.65 3.67 ;
      RECT 51.531 3.288 51.59 3.658 ;
      RECT 51.445 3.277 51.531 3.641 ;
      RECT 51.423 3.268 51.445 3.629 ;
      RECT 51.337 3.261 51.423 3.616 ;
      RECT 51.251 3.248 51.337 3.597 ;
      RECT 51.165 3.236 51.251 3.577 ;
      RECT 51.135 3.225 51.165 3.564 ;
      RECT 51.085 3.211 51.135 3.556 ;
      RECT 51.065 3.2 51.085 3.548 ;
      RECT 51.016 3.189 51.065 3.54 ;
      RECT 50.93 3.168 51.016 3.525 ;
      RECT 50.885 3.155 50.93 3.51 ;
      RECT 50.84 3.155 50.885 3.49 ;
      RECT 50.785 3.155 50.84 3.425 ;
      RECT 50.76 3.155 50.785 3.348 ;
      RECT 51.285 2.892 51.455 3.075 ;
      RECT 51.285 2.892 51.47 3.033 ;
      RECT 51.285 2.892 51.475 2.975 ;
      RECT 51.345 2.66 51.48 2.951 ;
      RECT 51.345 2.664 51.485 2.934 ;
      RECT 51.29 2.827 51.485 2.934 ;
      RECT 51.315 2.672 51.455 3.075 ;
      RECT 51.315 2.676 51.495 2.875 ;
      RECT 51.3 2.762 51.495 2.875 ;
      RECT 51.31 2.692 51.455 3.075 ;
      RECT 51.31 2.695 51.505 2.788 ;
      RECT 51.305 2.712 51.505 2.788 ;
      RECT 51.075 1.932 51.245 2.415 ;
      RECT 51.07 1.927 51.22 2.405 ;
      RECT 51.07 1.934 51.25 2.399 ;
      RECT 51.06 1.928 51.22 2.378 ;
      RECT 51.06 1.944 51.265 2.337 ;
      RECT 51.03 1.929 51.22 2.3 ;
      RECT 51.03 1.959 51.275 2.24 ;
      RECT 51.025 1.931 51.22 2.238 ;
      RECT 51.005 1.94 51.25 2.195 ;
      RECT 50.98 1.956 51.265 2.107 ;
      RECT 50.98 1.975 51.29 2.098 ;
      RECT 50.975 2.012 51.29 2.05 ;
      RECT 50.98 1.992 51.295 2.018 ;
      RECT 51.075 1.926 51.185 2.415 ;
      RECT 51.161 1.925 51.185 2.415 ;
      RECT 50.395 2.71 50.4 2.921 ;
      RECT 50.995 2.71 51 2.895 ;
      RECT 51.06 2.75 51.065 2.863 ;
      RECT 51.055 2.742 51.06 2.869 ;
      RECT 51.05 2.732 51.055 2.877 ;
      RECT 51.045 2.722 51.05 2.886 ;
      RECT 51.04 2.712 51.045 2.89 ;
      RECT 51 2.71 51.04 2.893 ;
      RECT 50.972 2.709 50.995 2.897 ;
      RECT 50.886 2.706 50.972 2.904 ;
      RECT 50.8 2.702 50.886 2.915 ;
      RECT 50.78 2.7 50.8 2.921 ;
      RECT 50.762 2.699 50.78 2.924 ;
      RECT 50.676 2.697 50.762 2.931 ;
      RECT 50.59 2.692 50.676 2.944 ;
      RECT 50.571 2.689 50.59 2.949 ;
      RECT 50.485 2.687 50.571 2.94 ;
      RECT 50.475 2.687 50.485 2.933 ;
      RECT 50.4 2.7 50.475 2.927 ;
      RECT 50.385 2.711 50.395 2.921 ;
      RECT 50.375 2.713 50.385 2.92 ;
      RECT 50.365 2.717 50.375 2.916 ;
      RECT 50.36 2.72 50.365 2.91 ;
      RECT 50.35 2.722 50.36 2.904 ;
      RECT 50.345 2.725 50.35 2.898 ;
      RECT 50.325 3.311 50.33 3.515 ;
      RECT 50.31 3.298 50.325 3.608 ;
      RECT 50.295 3.279 50.31 3.885 ;
      RECT 50.26 3.245 50.295 3.885 ;
      RECT 50.256 3.215 50.26 3.885 ;
      RECT 50.17 3.097 50.256 3.885 ;
      RECT 50.16 2.972 50.17 3.885 ;
      RECT 50.145 2.94 50.16 3.885 ;
      RECT 50.14 2.915 50.145 3.885 ;
      RECT 50.135 2.905 50.14 3.841 ;
      RECT 50.12 2.877 50.135 3.746 ;
      RECT 50.105 2.843 50.12 3.645 ;
      RECT 50.1 2.821 50.105 3.598 ;
      RECT 50.095 2.81 50.1 3.568 ;
      RECT 50.09 2.8 50.095 3.534 ;
      RECT 50.08 2.787 50.09 3.502 ;
      RECT 50.055 2.763 50.08 3.428 ;
      RECT 50.05 2.743 50.055 3.353 ;
      RECT 50.045 2.737 50.05 3.328 ;
      RECT 50.04 2.732 50.045 3.293 ;
      RECT 50.035 2.727 50.04 3.268 ;
      RECT 50.03 2.725 50.035 3.248 ;
      RECT 50.025 2.725 50.03 3.233 ;
      RECT 50.02 2.725 50.025 3.193 ;
      RECT 50.01 2.725 50.02 3.165 ;
      RECT 50 2.725 50.01 3.11 ;
      RECT 49.985 2.725 50 3.048 ;
      RECT 49.98 2.724 49.985 2.993 ;
      RECT 49.965 2.723 49.98 2.973 ;
      RECT 49.905 2.721 49.965 2.947 ;
      RECT 49.87 2.722 49.905 2.927 ;
      RECT 49.865 2.724 49.87 2.917 ;
      RECT 49.855 2.743 49.865 2.907 ;
      RECT 49.85 2.77 49.855 2.838 ;
      RECT 49.965 2.195 50.135 2.44 ;
      RECT 50 1.966 50.135 2.44 ;
      RECT 50 1.968 50.145 2.435 ;
      RECT 50 1.97 50.17 2.423 ;
      RECT 50 1.973 50.195 2.405 ;
      RECT 50 1.978 50.245 2.378 ;
      RECT 50 1.983 50.265 2.343 ;
      RECT 49.98 1.985 50.275 2.318 ;
      RECT 49.97 2.08 50.275 2.318 ;
      RECT 50 1.965 50.11 2.44 ;
      RECT 50.01 1.962 50.105 2.44 ;
      RECT 49.53 3.227 49.72 3.585 ;
      RECT 49.53 3.239 49.755 3.584 ;
      RECT 49.53 3.267 49.775 3.582 ;
      RECT 49.53 3.292 49.78 3.581 ;
      RECT 49.53 3.35 49.795 3.58 ;
      RECT 49.515 3.223 49.675 3.565 ;
      RECT 49.495 3.232 49.72 3.518 ;
      RECT 49.47 3.243 49.755 3.455 ;
      RECT 49.47 3.327 49.79 3.455 ;
      RECT 49.47 3.302 49.785 3.455 ;
      RECT 49.53 3.218 49.675 3.585 ;
      RECT 49.616 3.217 49.675 3.585 ;
      RECT 49.616 3.216 49.66 3.585 ;
      RECT 49.53 7.855 49.7 8.305 ;
      RECT 49.585 6.075 49.755 8.025 ;
      RECT 49.53 5.015 49.7 6.245 ;
      RECT 49.01 5.015 49.18 8.305 ;
      RECT 49.01 7.315 49.415 7.645 ;
      RECT 49.01 6.475 49.415 6.805 ;
      RECT 49.315 2.732 49.32 3.11 ;
      RECT 49.31 2.7 49.315 3.11 ;
      RECT 49.305 2.672 49.31 3.11 ;
      RECT 49.3 2.652 49.305 3.11 ;
      RECT 49.245 2.635 49.3 3.11 ;
      RECT 49.205 2.62 49.245 3.11 ;
      RECT 49.15 2.607 49.205 3.11 ;
      RECT 49.115 2.598 49.15 3.11 ;
      RECT 49.111 2.596 49.115 3.109 ;
      RECT 49.025 2.592 49.111 3.092 ;
      RECT 48.94 2.584 49.025 3.055 ;
      RECT 48.93 2.58 48.94 3.028 ;
      RECT 48.92 2.58 48.93 3.01 ;
      RECT 48.91 2.582 48.92 2.993 ;
      RECT 48.905 2.587 48.91 2.979 ;
      RECT 48.9 2.591 48.905 2.966 ;
      RECT 48.89 2.596 48.9 2.95 ;
      RECT 48.875 2.61 48.89 2.925 ;
      RECT 48.87 2.616 48.875 2.905 ;
      RECT 48.865 2.618 48.87 2.898 ;
      RECT 48.86 2.622 48.865 2.773 ;
      RECT 49.04 3.422 49.285 3.885 ;
      RECT 48.96 3.395 49.28 3.881 ;
      RECT 48.89 3.43 49.285 3.874 ;
      RECT 48.68 3.685 49.285 3.87 ;
      RECT 48.86 3.453 49.285 3.87 ;
      RECT 48.7 3.645 49.285 3.87 ;
      RECT 48.85 3.465 49.285 3.87 ;
      RECT 48.735 3.582 49.285 3.87 ;
      RECT 48.79 3.507 49.285 3.87 ;
      RECT 49.04 3.372 49.28 3.885 ;
      RECT 49.07 3.365 49.28 3.885 ;
      RECT 49.06 3.367 49.28 3.885 ;
      RECT 49.07 3.362 49.2 3.885 ;
      RECT 48.625 1.925 48.711 2.364 ;
      RECT 48.62 1.925 48.711 2.362 ;
      RECT 48.62 1.925 48.78 2.361 ;
      RECT 48.62 1.925 48.81 2.358 ;
      RECT 48.605 1.932 48.81 2.349 ;
      RECT 48.605 1.932 48.815 2.345 ;
      RECT 48.6 1.942 48.815 2.338 ;
      RECT 48.595 1.947 48.815 2.313 ;
      RECT 48.595 1.947 48.83 2.295 ;
      RECT 48.62 1.925 48.85 2.21 ;
      RECT 48.59 1.952 48.85 2.208 ;
      RECT 48.6 1.945 48.855 2.146 ;
      RECT 48.59 2.067 48.86 2.129 ;
      RECT 48.575 1.962 48.855 2.08 ;
      RECT 48.57 1.972 48.855 1.98 ;
      RECT 48.65 2.743 48.655 2.82 ;
      RECT 48.64 2.737 48.65 3.01 ;
      RECT 48.63 2.729 48.64 3.031 ;
      RECT 48.62 2.72 48.63 3.053 ;
      RECT 48.615 2.715 48.62 3.07 ;
      RECT 48.575 2.715 48.615 3.11 ;
      RECT 48.555 2.715 48.575 3.165 ;
      RECT 48.55 2.715 48.555 3.193 ;
      RECT 48.54 2.715 48.55 3.208 ;
      RECT 48.505 2.715 48.54 3.25 ;
      RECT 48.5 2.715 48.505 3.293 ;
      RECT 48.49 2.715 48.5 3.308 ;
      RECT 48.475 2.715 48.49 3.328 ;
      RECT 48.46 2.715 48.475 3.355 ;
      RECT 48.455 2.716 48.46 3.373 ;
      RECT 48.435 2.717 48.455 3.38 ;
      RECT 48.38 2.718 48.435 3.4 ;
      RECT 48.37 2.719 48.38 3.414 ;
      RECT 48.365 2.722 48.37 3.413 ;
      RECT 48.325 2.795 48.365 3.411 ;
      RECT 48.31 2.875 48.325 3.409 ;
      RECT 48.285 2.93 48.31 3.407 ;
      RECT 48.27 2.995 48.285 3.406 ;
      RECT 48.225 3.027 48.27 3.403 ;
      RECT 48.14 3.05 48.225 3.398 ;
      RECT 48.115 3.07 48.14 3.393 ;
      RECT 48.045 3.075 48.115 3.389 ;
      RECT 48.025 3.077 48.045 3.386 ;
      RECT 47.94 3.088 48.025 3.38 ;
      RECT 47.935 3.099 47.94 3.375 ;
      RECT 47.925 3.101 47.935 3.375 ;
      RECT 47.89 3.105 47.925 3.373 ;
      RECT 47.84 3.115 47.89 3.36 ;
      RECT 47.82 3.123 47.84 3.345 ;
      RECT 47.74 3.135 47.82 3.328 ;
      RECT 47.905 2.685 48.075 2.895 ;
      RECT 48.021 2.681 48.075 2.895 ;
      RECT 47.826 2.685 48.075 2.886 ;
      RECT 47.826 2.685 48.08 2.875 ;
      RECT 47.74 2.685 48.08 2.866 ;
      RECT 47.74 2.693 48.09 2.81 ;
      RECT 47.74 2.705 48.095 2.723 ;
      RECT 47.74 2.712 48.1 2.715 ;
      RECT 47.935 2.683 48.075 2.895 ;
      RECT 47.69 3.628 47.935 3.96 ;
      RECT 47.685 3.62 47.69 3.957 ;
      RECT 47.655 3.64 47.935 3.938 ;
      RECT 47.635 3.672 47.935 3.911 ;
      RECT 47.685 3.625 47.862 3.957 ;
      RECT 47.685 3.622 47.776 3.957 ;
      RECT 47.625 1.97 47.795 2.39 ;
      RECT 47.62 1.97 47.795 2.388 ;
      RECT 47.62 1.97 47.82 2.378 ;
      RECT 47.62 1.97 47.84 2.353 ;
      RECT 47.615 1.97 47.84 2.348 ;
      RECT 47.615 1.97 47.85 2.338 ;
      RECT 47.615 1.97 47.855 2.333 ;
      RECT 47.615 1.975 47.86 2.328 ;
      RECT 47.615 2.007 47.875 2.318 ;
      RECT 47.615 2.077 47.9 2.301 ;
      RECT 47.595 2.077 47.9 2.293 ;
      RECT 47.595 2.137 47.91 2.27 ;
      RECT 47.595 2.177 47.92 2.215 ;
      RECT 47.58 1.97 47.855 2.195 ;
      RECT 47.57 1.985 47.86 2.093 ;
      RECT 47.16 3.375 47.33 3.9 ;
      RECT 47.155 3.375 47.33 3.893 ;
      RECT 47.145 3.375 47.335 3.858 ;
      RECT 47.14 3.385 47.335 3.83 ;
      RECT 47.135 3.405 47.335 3.813 ;
      RECT 47.145 3.38 47.34 3.803 ;
      RECT 47.13 3.425 47.34 3.795 ;
      RECT 47.125 3.445 47.34 3.78 ;
      RECT 47.12 3.475 47.34 3.77 ;
      RECT 47.11 3.52 47.34 3.745 ;
      RECT 47.14 3.39 47.345 3.728 ;
      RECT 47.105 3.572 47.345 3.723 ;
      RECT 47.14 3.4 47.35 3.693 ;
      RECT 47.1 3.605 47.35 3.69 ;
      RECT 47.095 3.63 47.35 3.67 ;
      RECT 47.135 3.417 47.36 3.61 ;
      RECT 47.13 3.439 47.37 3.503 ;
      RECT 47.08 2.686 47.095 2.955 ;
      RECT 47.035 2.67 47.08 3 ;
      RECT 47.03 2.658 47.035 3.05 ;
      RECT 47.02 2.654 47.03 3.083 ;
      RECT 47.015 2.651 47.02 3.111 ;
      RECT 47 2.653 47.015 3.153 ;
      RECT 46.995 2.657 47 3.193 ;
      RECT 46.975 2.662 46.995 3.245 ;
      RECT 46.971 2.667 46.975 3.302 ;
      RECT 46.885 2.686 46.971 3.339 ;
      RECT 46.875 2.707 46.885 3.375 ;
      RECT 46.87 2.715 46.875 3.376 ;
      RECT 46.865 2.757 46.87 3.377 ;
      RECT 46.85 2.845 46.865 3.378 ;
      RECT 46.84 2.995 46.85 3.38 ;
      RECT 46.835 3.04 46.84 3.382 ;
      RECT 46.8 3.082 46.835 3.385 ;
      RECT 46.795 3.1 46.8 3.388 ;
      RECT 46.718 3.106 46.795 3.394 ;
      RECT 46.632 3.12 46.718 3.407 ;
      RECT 46.546 3.134 46.632 3.421 ;
      RECT 46.46 3.148 46.546 3.434 ;
      RECT 46.4 3.16 46.46 3.446 ;
      RECT 46.375 3.167 46.4 3.453 ;
      RECT 46.361 3.17 46.375 3.458 ;
      RECT 46.275 3.178 46.361 3.474 ;
      RECT 46.27 3.185 46.275 3.489 ;
      RECT 46.246 3.185 46.27 3.496 ;
      RECT 46.16 3.188 46.246 3.524 ;
      RECT 46.075 3.192 46.16 3.568 ;
      RECT 46.01 3.196 46.075 3.605 ;
      RECT 45.985 3.199 46.01 3.621 ;
      RECT 45.91 3.212 45.985 3.625 ;
      RECT 45.885 3.23 45.91 3.629 ;
      RECT 45.875 3.237 45.885 3.631 ;
      RECT 45.86 3.24 45.875 3.632 ;
      RECT 45.8 3.252 45.86 3.636 ;
      RECT 45.79 3.266 45.8 3.64 ;
      RECT 45.735 3.276 45.79 3.628 ;
      RECT 45.71 3.297 45.735 3.611 ;
      RECT 45.69 3.317 45.71 3.602 ;
      RECT 45.685 3.33 45.69 3.597 ;
      RECT 45.67 3.342 45.685 3.593 ;
      RECT 46.905 1.997 46.91 2.02 ;
      RECT 46.9 1.988 46.905 2.06 ;
      RECT 46.895 1.986 46.9 2.103 ;
      RECT 46.89 1.977 46.895 2.138 ;
      RECT 46.885 1.967 46.89 2.21 ;
      RECT 46.88 1.957 46.885 2.275 ;
      RECT 46.875 1.954 46.88 2.315 ;
      RECT 46.85 1.948 46.875 2.405 ;
      RECT 46.815 1.936 46.85 2.43 ;
      RECT 46.805 1.927 46.815 2.43 ;
      RECT 46.67 1.925 46.68 2.413 ;
      RECT 46.66 1.925 46.67 2.38 ;
      RECT 46.655 1.925 46.66 2.355 ;
      RECT 46.65 1.925 46.655 2.343 ;
      RECT 46.645 1.925 46.65 2.325 ;
      RECT 46.635 1.925 46.645 2.29 ;
      RECT 46.63 1.927 46.635 2.268 ;
      RECT 46.625 1.933 46.63 2.253 ;
      RECT 46.62 1.939 46.625 2.238 ;
      RECT 46.605 1.951 46.62 2.211 ;
      RECT 46.6 1.962 46.605 2.179 ;
      RECT 46.595 1.972 46.6 2.163 ;
      RECT 46.585 1.98 46.595 2.132 ;
      RECT 46.58 1.99 46.585 2.106 ;
      RECT 46.575 2.047 46.58 2.089 ;
      RECT 46.68 1.925 46.805 2.43 ;
      RECT 46.395 2.612 46.655 2.91 ;
      RECT 46.39 2.619 46.655 2.908 ;
      RECT 46.395 2.614 46.67 2.903 ;
      RECT 46.385 2.627 46.67 2.9 ;
      RECT 46.385 2.632 46.675 2.893 ;
      RECT 46.38 2.64 46.675 2.89 ;
      RECT 46.38 2.657 46.68 2.688 ;
      RECT 46.395 2.609 46.626 2.91 ;
      RECT 46.45 2.608 46.626 2.91 ;
      RECT 46.45 2.605 46.54 2.91 ;
      RECT 46.45 2.602 46.536 2.91 ;
      RECT 46.14 2.875 46.145 2.888 ;
      RECT 46.135 2.842 46.14 2.893 ;
      RECT 46.13 2.797 46.135 2.9 ;
      RECT 46.125 2.752 46.13 2.908 ;
      RECT 46.12 2.72 46.125 2.916 ;
      RECT 46.115 2.68 46.12 2.917 ;
      RECT 46.1 2.66 46.115 2.919 ;
      RECT 46.025 2.642 46.1 2.931 ;
      RECT 46.015 2.635 46.025 2.942 ;
      RECT 46.01 2.635 46.015 2.944 ;
      RECT 45.98 2.641 46.01 2.948 ;
      RECT 45.94 2.654 45.98 2.948 ;
      RECT 45.915 2.665 45.94 2.934 ;
      RECT 45.9 2.671 45.915 2.917 ;
      RECT 45.89 2.673 45.9 2.908 ;
      RECT 45.885 2.674 45.89 2.903 ;
      RECT 45.88 2.675 45.885 2.898 ;
      RECT 45.875 2.676 45.88 2.895 ;
      RECT 45.85 2.681 45.875 2.885 ;
      RECT 45.84 2.697 45.85 2.872 ;
      RECT 45.835 2.717 45.84 2.867 ;
      RECT 45.845 2.11 45.85 2.306 ;
      RECT 45.83 2.074 45.845 2.308 ;
      RECT 45.82 2.056 45.83 2.313 ;
      RECT 45.81 2.042 45.82 2.317 ;
      RECT 45.765 2.026 45.81 2.327 ;
      RECT 45.76 2.016 45.765 2.336 ;
      RECT 45.715 2.005 45.76 2.342 ;
      RECT 45.71 1.993 45.715 2.349 ;
      RECT 45.695 1.988 45.71 2.353 ;
      RECT 45.68 1.98 45.695 2.358 ;
      RECT 45.67 1.973 45.68 2.363 ;
      RECT 45.66 1.97 45.67 2.368 ;
      RECT 45.65 1.97 45.66 2.369 ;
      RECT 45.645 1.967 45.65 2.368 ;
      RECT 45.61 1.962 45.635 2.367 ;
      RECT 45.586 1.958 45.61 2.366 ;
      RECT 45.5 1.949 45.586 2.363 ;
      RECT 45.485 1.941 45.5 2.36 ;
      RECT 45.463 1.94 45.485 2.359 ;
      RECT 45.377 1.94 45.463 2.357 ;
      RECT 45.291 1.94 45.377 2.355 ;
      RECT 45.205 1.94 45.291 2.352 ;
      RECT 45.195 1.94 45.205 2.343 ;
      RECT 45.165 1.94 45.195 2.303 ;
      RECT 45.155 1.95 45.165 2.258 ;
      RECT 45.15 1.99 45.155 2.243 ;
      RECT 45.145 2.005 45.15 2.23 ;
      RECT 45.115 2.085 45.145 2.192 ;
      RECT 45.635 1.965 45.645 2.368 ;
      RECT 45.46 2.73 45.475 3.335 ;
      RECT 45.465 2.725 45.475 3.335 ;
      RECT 45.63 2.725 45.635 2.908 ;
      RECT 45.62 2.725 45.63 2.938 ;
      RECT 45.605 2.725 45.62 2.998 ;
      RECT 45.6 2.725 45.605 3.043 ;
      RECT 45.595 2.725 45.6 3.073 ;
      RECT 45.59 2.725 45.595 3.093 ;
      RECT 45.58 2.725 45.59 3.128 ;
      RECT 45.565 2.725 45.58 3.16 ;
      RECT 45.52 2.725 45.565 3.188 ;
      RECT 45.515 2.725 45.52 3.218 ;
      RECT 45.51 2.725 45.515 3.23 ;
      RECT 45.505 2.725 45.51 3.238 ;
      RECT 45.495 2.725 45.505 3.253 ;
      RECT 45.49 2.725 45.495 3.275 ;
      RECT 45.48 2.725 45.49 3.298 ;
      RECT 45.475 2.725 45.48 3.318 ;
      RECT 45.44 2.74 45.46 3.335 ;
      RECT 45.415 2.757 45.44 3.335 ;
      RECT 45.41 2.767 45.415 3.335 ;
      RECT 45.38 2.782 45.41 3.335 ;
      RECT 45.305 2.824 45.38 3.335 ;
      RECT 45.3 2.855 45.305 3.318 ;
      RECT 45.295 2.859 45.3 3.3 ;
      RECT 45.29 2.863 45.295 3.263 ;
      RECT 45.285 3.047 45.29 3.23 ;
      RECT 44.77 3.236 44.856 3.801 ;
      RECT 44.725 3.238 44.89 3.795 ;
      RECT 44.856 3.235 44.89 3.795 ;
      RECT 44.77 3.237 44.975 3.789 ;
      RECT 44.725 3.247 44.985 3.785 ;
      RECT 44.7 3.239 44.975 3.781 ;
      RECT 44.695 3.242 44.975 3.776 ;
      RECT 44.67 3.257 44.985 3.77 ;
      RECT 44.67 3.282 45.025 3.765 ;
      RECT 44.63 3.29 45.025 3.74 ;
      RECT 44.63 3.317 45.04 3.738 ;
      RECT 44.63 3.347 45.05 3.725 ;
      RECT 44.625 3.492 45.05 3.713 ;
      RECT 44.63 3.421 45.07 3.71 ;
      RECT 44.63 3.478 45.075 3.518 ;
      RECT 44.82 2.757 44.99 2.935 ;
      RECT 44.77 2.696 44.82 2.92 ;
      RECT 44.505 2.676 44.77 2.905 ;
      RECT 44.465 2.74 44.94 2.905 ;
      RECT 44.465 2.73 44.895 2.905 ;
      RECT 44.465 2.727 44.885 2.905 ;
      RECT 44.465 2.715 44.875 2.905 ;
      RECT 44.465 2.7 44.82 2.905 ;
      RECT 44.505 2.672 44.706 2.905 ;
      RECT 44.515 2.65 44.706 2.905 ;
      RECT 44.54 2.635 44.62 2.905 ;
      RECT 44.295 3.165 44.415 3.61 ;
      RECT 44.28 3.165 44.415 3.609 ;
      RECT 44.235 3.187 44.415 3.604 ;
      RECT 44.195 3.236 44.415 3.598 ;
      RECT 44.195 3.236 44.42 3.573 ;
      RECT 44.195 3.236 44.44 3.463 ;
      RECT 44.19 3.266 44.44 3.46 ;
      RECT 44.28 3.165 44.45 3.355 ;
      RECT 43.94 1.95 43.945 2.395 ;
      RECT 43.75 1.95 43.77 2.36 ;
      RECT 43.72 1.95 43.725 2.335 ;
      RECT 44.4 2.257 44.415 2.445 ;
      RECT 44.395 2.242 44.4 2.451 ;
      RECT 44.375 2.215 44.395 2.454 ;
      RECT 44.325 2.182 44.375 2.463 ;
      RECT 44.295 2.162 44.325 2.467 ;
      RECT 44.276 2.15 44.295 2.463 ;
      RECT 44.19 2.122 44.276 2.453 ;
      RECT 44.18 2.097 44.19 2.443 ;
      RECT 44.11 2.065 44.18 2.435 ;
      RECT 44.085 2.025 44.11 2.427 ;
      RECT 44.065 2.007 44.085 2.421 ;
      RECT 44.055 1.997 44.065 2.418 ;
      RECT 44.045 1.99 44.055 2.416 ;
      RECT 44.025 1.977 44.045 2.413 ;
      RECT 44.015 1.967 44.025 2.41 ;
      RECT 44.005 1.96 44.015 2.408 ;
      RECT 43.955 1.952 44.005 2.402 ;
      RECT 43.945 1.95 43.955 2.396 ;
      RECT 43.915 1.95 43.94 2.393 ;
      RECT 43.886 1.95 43.915 2.388 ;
      RECT 43.8 1.95 43.886 2.378 ;
      RECT 43.77 1.95 43.8 2.365 ;
      RECT 43.725 1.95 43.75 2.348 ;
      RECT 43.71 1.95 43.72 2.33 ;
      RECT 43.69 1.957 43.71 2.315 ;
      RECT 43.685 1.972 43.69 2.303 ;
      RECT 43.68 1.977 43.685 2.243 ;
      RECT 43.675 1.982 43.68 2.085 ;
      RECT 43.67 1.985 43.675 2.003 ;
      RECT 43.935 2.67 44.021 2.991 ;
      RECT 43.935 2.67 44.055 2.984 ;
      RECT 43.885 2.67 44.055 2.98 ;
      RECT 43.885 2.672 44.141 2.978 ;
      RECT 43.885 2.674 44.165 2.972 ;
      RECT 43.885 2.681 44.175 2.971 ;
      RECT 43.885 2.69 44.18 2.968 ;
      RECT 43.885 2.696 44.185 2.963 ;
      RECT 43.885 2.74 44.19 2.96 ;
      RECT 43.885 2.832 44.195 2.957 ;
      RECT 43.41 3.275 43.445 3.595 ;
      RECT 43.995 3.46 44 3.642 ;
      RECT 43.95 3.342 43.995 3.661 ;
      RECT 43.935 3.319 43.95 3.684 ;
      RECT 43.925 3.309 43.935 3.694 ;
      RECT 43.905 3.304 43.925 3.707 ;
      RECT 43.88 3.302 43.905 3.728 ;
      RECT 43.861 3.301 43.88 3.74 ;
      RECT 43.775 3.298 43.861 3.74 ;
      RECT 43.705 3.293 43.775 3.728 ;
      RECT 43.63 3.289 43.705 3.703 ;
      RECT 43.565 3.285 43.63 3.67 ;
      RECT 43.495 3.282 43.565 3.63 ;
      RECT 43.465 3.278 43.495 3.605 ;
      RECT 43.445 3.276 43.465 3.598 ;
      RECT 43.361 3.274 43.41 3.596 ;
      RECT 43.275 3.271 43.361 3.597 ;
      RECT 43.2 3.27 43.275 3.599 ;
      RECT 43.115 3.27 43.2 3.625 ;
      RECT 43.038 3.271 43.115 3.65 ;
      RECT 42.952 3.272 43.038 3.65 ;
      RECT 42.866 3.272 42.952 3.65 ;
      RECT 42.78 3.273 42.866 3.65 ;
      RECT 42.76 3.274 42.78 3.642 ;
      RECT 42.745 3.28 42.76 3.627 ;
      RECT 42.71 3.3 42.745 3.607 ;
      RECT 42.7 3.32 42.71 3.589 ;
      RECT 43.67 2.625 43.675 2.895 ;
      RECT 43.665 2.616 43.67 2.9 ;
      RECT 43.655 2.606 43.665 2.912 ;
      RECT 43.65 2.595 43.655 2.923 ;
      RECT 43.63 2.589 43.65 2.941 ;
      RECT 43.585 2.586 43.63 2.99 ;
      RECT 43.57 2.585 43.585 3.035 ;
      RECT 43.565 2.585 43.57 3.048 ;
      RECT 43.555 2.585 43.565 3.06 ;
      RECT 43.55 2.586 43.555 3.075 ;
      RECT 43.53 2.594 43.55 3.08 ;
      RECT 43.5 2.61 43.53 3.08 ;
      RECT 43.49 2.622 43.495 3.08 ;
      RECT 43.455 2.637 43.49 3.08 ;
      RECT 43.425 2.657 43.455 3.08 ;
      RECT 43.415 2.682 43.425 3.08 ;
      RECT 43.41 2.71 43.415 3.08 ;
      RECT 43.405 2.74 43.41 3.08 ;
      RECT 43.4 2.757 43.405 3.08 ;
      RECT 43.39 2.785 43.4 3.08 ;
      RECT 43.38 2.82 43.39 3.08 ;
      RECT 43.375 2.855 43.38 3.08 ;
      RECT 43.495 2.62 43.5 3.08 ;
      RECT 43.01 2.722 43.195 2.895 ;
      RECT 42.97 2.64 43.155 2.893 ;
      RECT 42.931 2.645 43.155 2.889 ;
      RECT 42.845 2.654 43.155 2.884 ;
      RECT 42.761 2.67 43.16 2.879 ;
      RECT 42.675 2.69 43.185 2.873 ;
      RECT 42.675 2.71 43.19 2.873 ;
      RECT 42.761 2.68 43.185 2.879 ;
      RECT 42.845 2.655 43.16 2.884 ;
      RECT 43.01 2.637 43.155 2.895 ;
      RECT 43.01 2.632 43.11 2.895 ;
      RECT 43.096 2.626 43.11 2.895 ;
      RECT 42.485 1.95 42.49 2.349 ;
      RECT 42.23 1.95 42.265 2.347 ;
      RECT 41.825 1.985 41.83 2.341 ;
      RECT 42.57 1.988 42.575 2.243 ;
      RECT 42.565 1.986 42.57 2.249 ;
      RECT 42.56 1.985 42.565 2.256 ;
      RECT 42.535 1.978 42.56 2.28 ;
      RECT 42.53 1.971 42.535 2.304 ;
      RECT 42.525 1.967 42.53 2.313 ;
      RECT 42.515 1.962 42.525 2.326 ;
      RECT 42.51 1.959 42.515 2.335 ;
      RECT 42.505 1.957 42.51 2.34 ;
      RECT 42.49 1.953 42.505 2.35 ;
      RECT 42.475 1.947 42.485 2.349 ;
      RECT 42.437 1.945 42.475 2.349 ;
      RECT 42.351 1.947 42.437 2.349 ;
      RECT 42.265 1.949 42.351 2.348 ;
      RECT 42.194 1.95 42.23 2.347 ;
      RECT 42.108 1.952 42.194 2.347 ;
      RECT 42.022 1.954 42.108 2.346 ;
      RECT 41.936 1.956 42.022 2.346 ;
      RECT 41.85 1.959 41.936 2.345 ;
      RECT 41.84 1.965 41.85 2.344 ;
      RECT 41.83 1.977 41.84 2.342 ;
      RECT 41.77 2.012 41.825 2.338 ;
      RECT 41.765 2.042 41.77 2.1 ;
      RECT 42.51 3.122 42.525 3.315 ;
      RECT 42.505 3.09 42.51 3.315 ;
      RECT 42.495 3.065 42.505 3.315 ;
      RECT 42.49 3.037 42.495 3.315 ;
      RECT 42.46 2.96 42.49 3.315 ;
      RECT 42.435 2.842 42.46 3.315 ;
      RECT 42.43 2.78 42.435 3.315 ;
      RECT 42.42 2.767 42.43 3.315 ;
      RECT 42.4 2.757 42.42 3.315 ;
      RECT 42.385 2.74 42.4 3.315 ;
      RECT 42.355 2.728 42.385 3.315 ;
      RECT 42.35 2.727 42.355 3.26 ;
      RECT 42.345 2.727 42.35 3.218 ;
      RECT 42.33 2.726 42.345 3.17 ;
      RECT 42.315 2.726 42.33 3.108 ;
      RECT 42.295 2.726 42.315 3.068 ;
      RECT 42.29 2.726 42.295 3.053 ;
      RECT 42.265 2.725 42.29 3.048 ;
      RECT 42.195 2.724 42.265 3.035 ;
      RECT 42.18 2.723 42.195 3.02 ;
      RECT 42.15 2.722 42.18 3.003 ;
      RECT 42.145 2.722 42.15 2.988 ;
      RECT 42.095 2.721 42.145 2.968 ;
      RECT 42.03 2.72 42.095 2.923 ;
      RECT 42.025 2.72 42.03 2.895 ;
      RECT 42.11 3.257 42.115 3.514 ;
      RECT 42.09 3.176 42.11 3.531 ;
      RECT 42.07 3.17 42.09 3.56 ;
      RECT 42.01 3.157 42.07 3.58 ;
      RECT 41.965 3.141 42.01 3.581 ;
      RECT 41.881 3.129 41.965 3.569 ;
      RECT 41.795 3.116 41.881 3.553 ;
      RECT 41.785 3.109 41.795 3.545 ;
      RECT 41.74 3.106 41.785 3.485 ;
      RECT 41.72 3.102 41.74 3.4 ;
      RECT 41.705 3.1 41.72 3.353 ;
      RECT 41.675 3.097 41.705 3.323 ;
      RECT 41.64 3.093 41.675 3.3 ;
      RECT 41.597 3.088 41.64 3.288 ;
      RECT 41.511 3.079 41.597 3.297 ;
      RECT 41.425 3.068 41.511 3.309 ;
      RECT 41.36 3.059 41.425 3.318 ;
      RECT 41.34 3.05 41.36 3.323 ;
      RECT 41.335 3.043 41.34 3.325 ;
      RECT 41.295 3.028 41.335 3.322 ;
      RECT 41.275 3.007 41.295 3.317 ;
      RECT 41.26 2.995 41.275 3.31 ;
      RECT 41.255 2.987 41.26 3.303 ;
      RECT 41.24 2.967 41.255 3.296 ;
      RECT 41.235 2.83 41.24 3.29 ;
      RECT 41.155 2.719 41.235 3.262 ;
      RECT 41.146 2.712 41.155 3.228 ;
      RECT 41.06 2.706 41.146 3.153 ;
      RECT 41.035 2.697 41.06 3.065 ;
      RECT 41.005 2.692 41.035 3.04 ;
      RECT 40.94 2.701 41.005 3.025 ;
      RECT 40.92 2.717 40.94 3 ;
      RECT 40.91 2.723 40.92 2.948 ;
      RECT 40.89 2.745 40.91 2.83 ;
      RECT 41.545 2.71 41.715 2.895 ;
      RECT 41.545 2.71 41.75 2.893 ;
      RECT 41.595 2.62 41.765 2.884 ;
      RECT 41.545 2.777 41.77 2.877 ;
      RECT 41.56 2.655 41.765 2.884 ;
      RECT 40.76 3.388 40.825 3.831 ;
      RECT 40.7 3.413 40.825 3.829 ;
      RECT 40.7 3.413 40.88 3.823 ;
      RECT 40.685 3.438 40.88 3.822 ;
      RECT 40.825 3.375 40.9 3.819 ;
      RECT 40.76 3.4 40.98 3.813 ;
      RECT 40.685 3.439 41.025 3.807 ;
      RECT 40.67 3.466 41.025 3.798 ;
      RECT 40.685 3.459 41.045 3.79 ;
      RECT 40.67 3.468 41.05 3.773 ;
      RECT 40.665 3.485 41.05 3.6 ;
      RECT 40.67 2.207 40.705 2.445 ;
      RECT 40.67 2.207 40.735 2.444 ;
      RECT 40.67 2.207 40.85 2.44 ;
      RECT 40.67 2.207 40.905 2.418 ;
      RECT 40.68 2.15 40.96 2.318 ;
      RECT 40.785 1.99 40.815 2.441 ;
      RECT 40.815 1.985 40.995 2.198 ;
      RECT 40.685 2.126 40.995 2.198 ;
      RECT 40.735 2.022 40.785 2.442 ;
      RECT 40.705 2.078 40.995 2.198 ;
      RECT 39.575 5.02 39.745 6.49 ;
      RECT 39.575 6.315 39.75 6.485 ;
      RECT 39.205 1.74 39.375 2.93 ;
      RECT 39.205 1.74 39.675 1.91 ;
      RECT 39.205 6.97 39.675 7.14 ;
      RECT 39.205 5.95 39.375 7.14 ;
      RECT 38.215 1.74 38.385 2.93 ;
      RECT 38.215 1.74 38.685 1.91 ;
      RECT 38.215 6.97 38.685 7.14 ;
      RECT 38.215 5.95 38.385 7.14 ;
      RECT 36.365 2.635 36.535 3.865 ;
      RECT 36.42 0.855 36.59 2.805 ;
      RECT 36.365 0.575 36.535 1.025 ;
      RECT 36.365 7.855 36.535 8.305 ;
      RECT 36.42 6.075 36.59 8.025 ;
      RECT 36.365 5.015 36.535 6.245 ;
      RECT 35.845 0.575 36.015 3.865 ;
      RECT 35.845 2.075 36.25 2.405 ;
      RECT 35.845 1.235 36.25 1.565 ;
      RECT 35.845 5.015 36.015 8.305 ;
      RECT 35.845 7.315 36.25 7.645 ;
      RECT 35.845 6.475 36.25 6.805 ;
      RECT 33.945 3.392 33.96 3.443 ;
      RECT 33.94 3.372 33.945 3.49 ;
      RECT 33.925 3.362 33.94 3.558 ;
      RECT 33.9 3.342 33.925 3.613 ;
      RECT 33.86 3.327 33.9 3.633 ;
      RECT 33.815 3.321 33.86 3.661 ;
      RECT 33.745 3.311 33.815 3.678 ;
      RECT 33.725 3.303 33.745 3.678 ;
      RECT 33.665 3.297 33.725 3.67 ;
      RECT 33.606 3.288 33.665 3.658 ;
      RECT 33.52 3.277 33.606 3.641 ;
      RECT 33.498 3.268 33.52 3.629 ;
      RECT 33.412 3.261 33.498 3.616 ;
      RECT 33.326 3.248 33.412 3.597 ;
      RECT 33.24 3.236 33.326 3.577 ;
      RECT 33.21 3.225 33.24 3.564 ;
      RECT 33.16 3.211 33.21 3.556 ;
      RECT 33.14 3.2 33.16 3.548 ;
      RECT 33.091 3.189 33.14 3.54 ;
      RECT 33.005 3.168 33.091 3.525 ;
      RECT 32.96 3.155 33.005 3.51 ;
      RECT 32.915 3.155 32.96 3.49 ;
      RECT 32.86 3.155 32.915 3.425 ;
      RECT 32.835 3.155 32.86 3.348 ;
      RECT 33.36 2.892 33.53 3.075 ;
      RECT 33.36 2.892 33.545 3.033 ;
      RECT 33.36 2.892 33.55 2.975 ;
      RECT 33.42 2.66 33.555 2.951 ;
      RECT 33.42 2.664 33.56 2.934 ;
      RECT 33.365 2.827 33.56 2.934 ;
      RECT 33.39 2.672 33.53 3.075 ;
      RECT 33.39 2.676 33.57 2.875 ;
      RECT 33.375 2.762 33.57 2.875 ;
      RECT 33.385 2.692 33.53 3.075 ;
      RECT 33.385 2.695 33.58 2.788 ;
      RECT 33.38 2.712 33.58 2.788 ;
      RECT 33.15 1.932 33.32 2.415 ;
      RECT 33.145 1.927 33.295 2.405 ;
      RECT 33.145 1.934 33.325 2.399 ;
      RECT 33.135 1.928 33.295 2.378 ;
      RECT 33.135 1.944 33.34 2.337 ;
      RECT 33.105 1.929 33.295 2.3 ;
      RECT 33.105 1.959 33.35 2.24 ;
      RECT 33.1 1.931 33.295 2.238 ;
      RECT 33.08 1.94 33.325 2.195 ;
      RECT 33.055 1.956 33.34 2.107 ;
      RECT 33.055 1.975 33.365 2.098 ;
      RECT 33.05 2.012 33.365 2.05 ;
      RECT 33.055 1.992 33.37 2.018 ;
      RECT 33.15 1.926 33.26 2.415 ;
      RECT 33.236 1.925 33.26 2.415 ;
      RECT 32.47 2.71 32.475 2.921 ;
      RECT 33.07 2.71 33.075 2.895 ;
      RECT 33.135 2.75 33.14 2.863 ;
      RECT 33.13 2.742 33.135 2.869 ;
      RECT 33.125 2.732 33.13 2.877 ;
      RECT 33.12 2.722 33.125 2.886 ;
      RECT 33.115 2.712 33.12 2.89 ;
      RECT 33.075 2.71 33.115 2.893 ;
      RECT 33.047 2.709 33.07 2.897 ;
      RECT 32.961 2.706 33.047 2.904 ;
      RECT 32.875 2.702 32.961 2.915 ;
      RECT 32.855 2.7 32.875 2.921 ;
      RECT 32.837 2.699 32.855 2.924 ;
      RECT 32.751 2.697 32.837 2.931 ;
      RECT 32.665 2.692 32.751 2.944 ;
      RECT 32.646 2.689 32.665 2.949 ;
      RECT 32.56 2.687 32.646 2.94 ;
      RECT 32.55 2.687 32.56 2.933 ;
      RECT 32.475 2.7 32.55 2.927 ;
      RECT 32.46 2.711 32.47 2.921 ;
      RECT 32.45 2.713 32.46 2.92 ;
      RECT 32.44 2.717 32.45 2.916 ;
      RECT 32.435 2.72 32.44 2.91 ;
      RECT 32.425 2.722 32.435 2.904 ;
      RECT 32.42 2.725 32.425 2.898 ;
      RECT 32.4 3.311 32.405 3.515 ;
      RECT 32.385 3.298 32.4 3.608 ;
      RECT 32.37 3.279 32.385 3.885 ;
      RECT 32.335 3.245 32.37 3.885 ;
      RECT 32.331 3.215 32.335 3.885 ;
      RECT 32.245 3.097 32.331 3.885 ;
      RECT 32.235 2.972 32.245 3.885 ;
      RECT 32.22 2.94 32.235 3.885 ;
      RECT 32.215 2.915 32.22 3.885 ;
      RECT 32.21 2.905 32.215 3.841 ;
      RECT 32.195 2.877 32.21 3.746 ;
      RECT 32.18 2.843 32.195 3.645 ;
      RECT 32.175 2.821 32.18 3.598 ;
      RECT 32.17 2.81 32.175 3.568 ;
      RECT 32.165 2.8 32.17 3.534 ;
      RECT 32.155 2.787 32.165 3.502 ;
      RECT 32.13 2.763 32.155 3.428 ;
      RECT 32.125 2.743 32.13 3.353 ;
      RECT 32.12 2.737 32.125 3.328 ;
      RECT 32.115 2.732 32.12 3.293 ;
      RECT 32.11 2.727 32.115 3.268 ;
      RECT 32.105 2.725 32.11 3.248 ;
      RECT 32.1 2.725 32.105 3.233 ;
      RECT 32.095 2.725 32.1 3.193 ;
      RECT 32.085 2.725 32.095 3.165 ;
      RECT 32.075 2.725 32.085 3.11 ;
      RECT 32.06 2.725 32.075 3.048 ;
      RECT 32.055 2.724 32.06 2.993 ;
      RECT 32.04 2.723 32.055 2.973 ;
      RECT 31.98 2.721 32.04 2.947 ;
      RECT 31.945 2.722 31.98 2.927 ;
      RECT 31.94 2.724 31.945 2.917 ;
      RECT 31.93 2.743 31.94 2.907 ;
      RECT 31.925 2.77 31.93 2.838 ;
      RECT 32.04 2.195 32.21 2.44 ;
      RECT 32.075 1.966 32.21 2.44 ;
      RECT 32.075 1.968 32.22 2.435 ;
      RECT 32.075 1.97 32.245 2.423 ;
      RECT 32.075 1.973 32.27 2.405 ;
      RECT 32.075 1.978 32.32 2.378 ;
      RECT 32.075 1.983 32.34 2.343 ;
      RECT 32.055 1.985 32.35 2.318 ;
      RECT 32.045 2.08 32.35 2.318 ;
      RECT 32.075 1.965 32.185 2.44 ;
      RECT 32.085 1.962 32.18 2.44 ;
      RECT 31.605 3.227 31.795 3.585 ;
      RECT 31.605 3.239 31.83 3.584 ;
      RECT 31.605 3.267 31.85 3.582 ;
      RECT 31.605 3.292 31.855 3.581 ;
      RECT 31.605 3.35 31.87 3.58 ;
      RECT 31.59 3.223 31.75 3.565 ;
      RECT 31.57 3.232 31.795 3.518 ;
      RECT 31.545 3.243 31.83 3.455 ;
      RECT 31.545 3.327 31.865 3.455 ;
      RECT 31.545 3.302 31.86 3.455 ;
      RECT 31.605 3.218 31.75 3.585 ;
      RECT 31.691 3.217 31.75 3.585 ;
      RECT 31.691 3.216 31.735 3.585 ;
      RECT 31.605 7.855 31.775 8.305 ;
      RECT 31.66 6.075 31.83 8.025 ;
      RECT 31.605 5.015 31.775 6.245 ;
      RECT 31.085 5.015 31.255 8.305 ;
      RECT 31.085 7.315 31.49 7.645 ;
      RECT 31.085 6.475 31.49 6.805 ;
      RECT 31.39 2.732 31.395 3.11 ;
      RECT 31.385 2.7 31.39 3.11 ;
      RECT 31.38 2.672 31.385 3.11 ;
      RECT 31.375 2.652 31.38 3.11 ;
      RECT 31.32 2.635 31.375 3.11 ;
      RECT 31.28 2.62 31.32 3.11 ;
      RECT 31.225 2.607 31.28 3.11 ;
      RECT 31.19 2.598 31.225 3.11 ;
      RECT 31.186 2.596 31.19 3.109 ;
      RECT 31.1 2.592 31.186 3.092 ;
      RECT 31.015 2.584 31.1 3.055 ;
      RECT 31.005 2.58 31.015 3.028 ;
      RECT 30.995 2.58 31.005 3.01 ;
      RECT 30.985 2.582 30.995 2.993 ;
      RECT 30.98 2.587 30.985 2.979 ;
      RECT 30.975 2.591 30.98 2.966 ;
      RECT 30.965 2.596 30.975 2.95 ;
      RECT 30.95 2.61 30.965 2.925 ;
      RECT 30.945 2.616 30.95 2.905 ;
      RECT 30.94 2.618 30.945 2.898 ;
      RECT 30.935 2.622 30.94 2.773 ;
      RECT 31.115 3.422 31.36 3.885 ;
      RECT 31.035 3.395 31.355 3.881 ;
      RECT 30.965 3.43 31.36 3.874 ;
      RECT 30.755 3.685 31.36 3.87 ;
      RECT 30.935 3.453 31.36 3.87 ;
      RECT 30.775 3.645 31.36 3.87 ;
      RECT 30.925 3.465 31.36 3.87 ;
      RECT 30.81 3.582 31.36 3.87 ;
      RECT 30.865 3.507 31.36 3.87 ;
      RECT 31.115 3.372 31.355 3.885 ;
      RECT 31.145 3.365 31.355 3.885 ;
      RECT 31.135 3.367 31.355 3.885 ;
      RECT 31.145 3.362 31.275 3.885 ;
      RECT 30.7 1.925 30.786 2.364 ;
      RECT 30.695 1.925 30.786 2.362 ;
      RECT 30.695 1.925 30.855 2.361 ;
      RECT 30.695 1.925 30.885 2.358 ;
      RECT 30.68 1.932 30.885 2.349 ;
      RECT 30.68 1.932 30.89 2.345 ;
      RECT 30.675 1.942 30.89 2.338 ;
      RECT 30.67 1.947 30.89 2.313 ;
      RECT 30.67 1.947 30.905 2.295 ;
      RECT 30.695 1.925 30.925 2.21 ;
      RECT 30.665 1.952 30.925 2.208 ;
      RECT 30.675 1.945 30.93 2.146 ;
      RECT 30.665 2.067 30.935 2.129 ;
      RECT 30.65 1.962 30.93 2.08 ;
      RECT 30.645 1.972 30.93 1.98 ;
      RECT 30.725 2.743 30.73 2.82 ;
      RECT 30.715 2.737 30.725 3.01 ;
      RECT 30.705 2.729 30.715 3.031 ;
      RECT 30.695 2.72 30.705 3.053 ;
      RECT 30.69 2.715 30.695 3.07 ;
      RECT 30.65 2.715 30.69 3.11 ;
      RECT 30.63 2.715 30.65 3.165 ;
      RECT 30.625 2.715 30.63 3.193 ;
      RECT 30.615 2.715 30.625 3.208 ;
      RECT 30.58 2.715 30.615 3.25 ;
      RECT 30.575 2.715 30.58 3.293 ;
      RECT 30.565 2.715 30.575 3.308 ;
      RECT 30.55 2.715 30.565 3.328 ;
      RECT 30.535 2.715 30.55 3.355 ;
      RECT 30.53 2.716 30.535 3.373 ;
      RECT 30.51 2.717 30.53 3.38 ;
      RECT 30.455 2.718 30.51 3.4 ;
      RECT 30.445 2.719 30.455 3.414 ;
      RECT 30.44 2.722 30.445 3.413 ;
      RECT 30.4 2.795 30.44 3.411 ;
      RECT 30.385 2.875 30.4 3.409 ;
      RECT 30.36 2.93 30.385 3.407 ;
      RECT 30.345 2.995 30.36 3.406 ;
      RECT 30.3 3.027 30.345 3.403 ;
      RECT 30.215 3.05 30.3 3.398 ;
      RECT 30.19 3.07 30.215 3.393 ;
      RECT 30.12 3.075 30.19 3.389 ;
      RECT 30.1 3.077 30.12 3.386 ;
      RECT 30.015 3.088 30.1 3.38 ;
      RECT 30.01 3.099 30.015 3.375 ;
      RECT 30 3.101 30.01 3.375 ;
      RECT 29.965 3.105 30 3.373 ;
      RECT 29.915 3.115 29.965 3.36 ;
      RECT 29.895 3.123 29.915 3.345 ;
      RECT 29.815 3.135 29.895 3.328 ;
      RECT 29.98 2.685 30.15 2.895 ;
      RECT 30.096 2.681 30.15 2.895 ;
      RECT 29.901 2.685 30.15 2.886 ;
      RECT 29.901 2.685 30.155 2.875 ;
      RECT 29.815 2.685 30.155 2.866 ;
      RECT 29.815 2.693 30.165 2.81 ;
      RECT 29.815 2.705 30.17 2.723 ;
      RECT 29.815 2.712 30.175 2.715 ;
      RECT 30.01 2.683 30.15 2.895 ;
      RECT 29.765 3.628 30.01 3.96 ;
      RECT 29.76 3.62 29.765 3.957 ;
      RECT 29.73 3.64 30.01 3.938 ;
      RECT 29.71 3.672 30.01 3.911 ;
      RECT 29.76 3.625 29.937 3.957 ;
      RECT 29.76 3.622 29.851 3.957 ;
      RECT 29.7 1.97 29.87 2.39 ;
      RECT 29.695 1.97 29.87 2.388 ;
      RECT 29.695 1.97 29.895 2.378 ;
      RECT 29.695 1.97 29.915 2.353 ;
      RECT 29.69 1.97 29.915 2.348 ;
      RECT 29.69 1.97 29.925 2.338 ;
      RECT 29.69 1.97 29.93 2.333 ;
      RECT 29.69 1.975 29.935 2.328 ;
      RECT 29.69 2.007 29.95 2.318 ;
      RECT 29.69 2.077 29.975 2.301 ;
      RECT 29.67 2.077 29.975 2.293 ;
      RECT 29.67 2.137 29.985 2.27 ;
      RECT 29.67 2.177 29.995 2.215 ;
      RECT 29.655 1.97 29.93 2.195 ;
      RECT 29.645 1.985 29.935 2.093 ;
      RECT 29.235 3.375 29.405 3.9 ;
      RECT 29.23 3.375 29.405 3.893 ;
      RECT 29.22 3.375 29.41 3.858 ;
      RECT 29.215 3.385 29.41 3.83 ;
      RECT 29.21 3.405 29.41 3.813 ;
      RECT 29.22 3.38 29.415 3.803 ;
      RECT 29.205 3.425 29.415 3.795 ;
      RECT 29.2 3.445 29.415 3.78 ;
      RECT 29.195 3.475 29.415 3.77 ;
      RECT 29.185 3.52 29.415 3.745 ;
      RECT 29.215 3.39 29.42 3.728 ;
      RECT 29.18 3.572 29.42 3.723 ;
      RECT 29.215 3.4 29.425 3.693 ;
      RECT 29.175 3.605 29.425 3.69 ;
      RECT 29.17 3.63 29.425 3.67 ;
      RECT 29.21 3.417 29.435 3.61 ;
      RECT 29.205 3.439 29.445 3.503 ;
      RECT 29.155 2.686 29.17 2.955 ;
      RECT 29.11 2.67 29.155 3 ;
      RECT 29.105 2.658 29.11 3.05 ;
      RECT 29.095 2.654 29.105 3.083 ;
      RECT 29.09 2.651 29.095 3.111 ;
      RECT 29.075 2.653 29.09 3.153 ;
      RECT 29.07 2.657 29.075 3.193 ;
      RECT 29.05 2.662 29.07 3.245 ;
      RECT 29.046 2.667 29.05 3.302 ;
      RECT 28.96 2.686 29.046 3.339 ;
      RECT 28.95 2.707 28.96 3.375 ;
      RECT 28.945 2.715 28.95 3.376 ;
      RECT 28.94 2.757 28.945 3.377 ;
      RECT 28.925 2.845 28.94 3.378 ;
      RECT 28.915 2.995 28.925 3.38 ;
      RECT 28.91 3.04 28.915 3.382 ;
      RECT 28.875 3.082 28.91 3.385 ;
      RECT 28.87 3.1 28.875 3.388 ;
      RECT 28.793 3.106 28.87 3.394 ;
      RECT 28.707 3.12 28.793 3.407 ;
      RECT 28.621 3.134 28.707 3.421 ;
      RECT 28.535 3.148 28.621 3.434 ;
      RECT 28.475 3.16 28.535 3.446 ;
      RECT 28.45 3.167 28.475 3.453 ;
      RECT 28.436 3.17 28.45 3.458 ;
      RECT 28.35 3.178 28.436 3.474 ;
      RECT 28.345 3.185 28.35 3.489 ;
      RECT 28.321 3.185 28.345 3.496 ;
      RECT 28.235 3.188 28.321 3.524 ;
      RECT 28.15 3.192 28.235 3.568 ;
      RECT 28.085 3.196 28.15 3.605 ;
      RECT 28.06 3.199 28.085 3.621 ;
      RECT 27.985 3.212 28.06 3.625 ;
      RECT 27.96 3.23 27.985 3.629 ;
      RECT 27.95 3.237 27.96 3.631 ;
      RECT 27.935 3.24 27.95 3.632 ;
      RECT 27.875 3.252 27.935 3.636 ;
      RECT 27.865 3.266 27.875 3.64 ;
      RECT 27.81 3.276 27.865 3.628 ;
      RECT 27.785 3.297 27.81 3.611 ;
      RECT 27.765 3.317 27.785 3.602 ;
      RECT 27.76 3.33 27.765 3.597 ;
      RECT 27.745 3.342 27.76 3.593 ;
      RECT 28.98 1.997 28.985 2.02 ;
      RECT 28.975 1.988 28.98 2.06 ;
      RECT 28.97 1.986 28.975 2.103 ;
      RECT 28.965 1.977 28.97 2.138 ;
      RECT 28.96 1.967 28.965 2.21 ;
      RECT 28.955 1.957 28.96 2.275 ;
      RECT 28.95 1.954 28.955 2.315 ;
      RECT 28.925 1.948 28.95 2.405 ;
      RECT 28.89 1.936 28.925 2.43 ;
      RECT 28.88 1.927 28.89 2.43 ;
      RECT 28.745 1.925 28.755 2.413 ;
      RECT 28.735 1.925 28.745 2.38 ;
      RECT 28.73 1.925 28.735 2.355 ;
      RECT 28.725 1.925 28.73 2.343 ;
      RECT 28.72 1.925 28.725 2.325 ;
      RECT 28.71 1.925 28.72 2.29 ;
      RECT 28.705 1.927 28.71 2.268 ;
      RECT 28.7 1.933 28.705 2.253 ;
      RECT 28.695 1.939 28.7 2.238 ;
      RECT 28.68 1.951 28.695 2.211 ;
      RECT 28.675 1.962 28.68 2.179 ;
      RECT 28.67 1.972 28.675 2.163 ;
      RECT 28.66 1.98 28.67 2.132 ;
      RECT 28.655 1.99 28.66 2.106 ;
      RECT 28.65 2.047 28.655 2.089 ;
      RECT 28.755 1.925 28.88 2.43 ;
      RECT 28.47 2.612 28.73 2.91 ;
      RECT 28.465 2.619 28.73 2.908 ;
      RECT 28.47 2.614 28.745 2.903 ;
      RECT 28.46 2.627 28.745 2.9 ;
      RECT 28.46 2.632 28.75 2.893 ;
      RECT 28.455 2.64 28.75 2.89 ;
      RECT 28.455 2.657 28.755 2.688 ;
      RECT 28.47 2.609 28.701 2.91 ;
      RECT 28.525 2.608 28.701 2.91 ;
      RECT 28.525 2.605 28.615 2.91 ;
      RECT 28.525 2.602 28.611 2.91 ;
      RECT 28.215 2.875 28.22 2.888 ;
      RECT 28.21 2.842 28.215 2.893 ;
      RECT 28.205 2.797 28.21 2.9 ;
      RECT 28.2 2.752 28.205 2.908 ;
      RECT 28.195 2.72 28.2 2.916 ;
      RECT 28.19 2.68 28.195 2.917 ;
      RECT 28.175 2.66 28.19 2.919 ;
      RECT 28.1 2.642 28.175 2.931 ;
      RECT 28.09 2.635 28.1 2.942 ;
      RECT 28.085 2.635 28.09 2.944 ;
      RECT 28.055 2.641 28.085 2.948 ;
      RECT 28.015 2.654 28.055 2.948 ;
      RECT 27.99 2.665 28.015 2.934 ;
      RECT 27.975 2.671 27.99 2.917 ;
      RECT 27.965 2.673 27.975 2.908 ;
      RECT 27.96 2.674 27.965 2.903 ;
      RECT 27.955 2.675 27.96 2.898 ;
      RECT 27.95 2.676 27.955 2.895 ;
      RECT 27.925 2.681 27.95 2.885 ;
      RECT 27.915 2.697 27.925 2.872 ;
      RECT 27.91 2.717 27.915 2.867 ;
      RECT 27.92 2.11 27.925 2.306 ;
      RECT 27.905 2.074 27.92 2.308 ;
      RECT 27.895 2.056 27.905 2.313 ;
      RECT 27.885 2.042 27.895 2.317 ;
      RECT 27.84 2.026 27.885 2.327 ;
      RECT 27.835 2.016 27.84 2.336 ;
      RECT 27.79 2.005 27.835 2.342 ;
      RECT 27.785 1.993 27.79 2.349 ;
      RECT 27.77 1.988 27.785 2.353 ;
      RECT 27.755 1.98 27.77 2.358 ;
      RECT 27.745 1.973 27.755 2.363 ;
      RECT 27.735 1.97 27.745 2.368 ;
      RECT 27.725 1.97 27.735 2.369 ;
      RECT 27.72 1.967 27.725 2.368 ;
      RECT 27.685 1.962 27.71 2.367 ;
      RECT 27.661 1.958 27.685 2.366 ;
      RECT 27.575 1.949 27.661 2.363 ;
      RECT 27.56 1.941 27.575 2.36 ;
      RECT 27.538 1.94 27.56 2.359 ;
      RECT 27.452 1.94 27.538 2.357 ;
      RECT 27.366 1.94 27.452 2.355 ;
      RECT 27.28 1.94 27.366 2.352 ;
      RECT 27.27 1.94 27.28 2.343 ;
      RECT 27.24 1.94 27.27 2.303 ;
      RECT 27.23 1.95 27.24 2.258 ;
      RECT 27.225 1.99 27.23 2.243 ;
      RECT 27.22 2.005 27.225 2.23 ;
      RECT 27.19 2.085 27.22 2.192 ;
      RECT 27.71 1.965 27.72 2.368 ;
      RECT 27.535 2.73 27.55 3.335 ;
      RECT 27.54 2.725 27.55 3.335 ;
      RECT 27.705 2.725 27.71 2.908 ;
      RECT 27.695 2.725 27.705 2.938 ;
      RECT 27.68 2.725 27.695 2.998 ;
      RECT 27.675 2.725 27.68 3.043 ;
      RECT 27.67 2.725 27.675 3.073 ;
      RECT 27.665 2.725 27.67 3.093 ;
      RECT 27.655 2.725 27.665 3.128 ;
      RECT 27.64 2.725 27.655 3.16 ;
      RECT 27.595 2.725 27.64 3.188 ;
      RECT 27.59 2.725 27.595 3.218 ;
      RECT 27.585 2.725 27.59 3.23 ;
      RECT 27.58 2.725 27.585 3.238 ;
      RECT 27.57 2.725 27.58 3.253 ;
      RECT 27.565 2.725 27.57 3.275 ;
      RECT 27.555 2.725 27.565 3.298 ;
      RECT 27.55 2.725 27.555 3.318 ;
      RECT 27.515 2.74 27.535 3.335 ;
      RECT 27.49 2.757 27.515 3.335 ;
      RECT 27.485 2.767 27.49 3.335 ;
      RECT 27.455 2.782 27.485 3.335 ;
      RECT 27.38 2.824 27.455 3.335 ;
      RECT 27.375 2.855 27.38 3.318 ;
      RECT 27.37 2.859 27.375 3.3 ;
      RECT 27.365 2.863 27.37 3.263 ;
      RECT 27.36 3.047 27.365 3.23 ;
      RECT 26.845 3.236 26.931 3.801 ;
      RECT 26.8 3.238 26.965 3.795 ;
      RECT 26.931 3.235 26.965 3.795 ;
      RECT 26.845 3.237 27.05 3.789 ;
      RECT 26.8 3.247 27.06 3.785 ;
      RECT 26.775 3.239 27.05 3.781 ;
      RECT 26.77 3.242 27.05 3.776 ;
      RECT 26.745 3.257 27.06 3.77 ;
      RECT 26.745 3.282 27.1 3.765 ;
      RECT 26.705 3.29 27.1 3.74 ;
      RECT 26.705 3.317 27.115 3.738 ;
      RECT 26.705 3.347 27.125 3.725 ;
      RECT 26.7 3.492 27.125 3.713 ;
      RECT 26.705 3.421 27.145 3.71 ;
      RECT 26.705 3.478 27.15 3.518 ;
      RECT 26.895 2.757 27.065 2.935 ;
      RECT 26.845 2.696 26.895 2.92 ;
      RECT 26.58 2.676 26.845 2.905 ;
      RECT 26.54 2.74 27.015 2.905 ;
      RECT 26.54 2.73 26.97 2.905 ;
      RECT 26.54 2.727 26.96 2.905 ;
      RECT 26.54 2.715 26.95 2.905 ;
      RECT 26.54 2.7 26.895 2.905 ;
      RECT 26.58 2.672 26.781 2.905 ;
      RECT 26.59 2.65 26.781 2.905 ;
      RECT 26.615 2.635 26.695 2.905 ;
      RECT 26.37 3.165 26.49 3.61 ;
      RECT 26.355 3.165 26.49 3.609 ;
      RECT 26.31 3.187 26.49 3.604 ;
      RECT 26.27 3.236 26.49 3.598 ;
      RECT 26.27 3.236 26.495 3.573 ;
      RECT 26.27 3.236 26.515 3.463 ;
      RECT 26.265 3.266 26.515 3.46 ;
      RECT 26.355 3.165 26.525 3.355 ;
      RECT 26.015 1.95 26.02 2.395 ;
      RECT 25.825 1.95 25.845 2.36 ;
      RECT 25.795 1.95 25.8 2.335 ;
      RECT 26.475 2.257 26.49 2.445 ;
      RECT 26.47 2.242 26.475 2.451 ;
      RECT 26.45 2.215 26.47 2.454 ;
      RECT 26.4 2.182 26.45 2.463 ;
      RECT 26.37 2.162 26.4 2.467 ;
      RECT 26.351 2.15 26.37 2.463 ;
      RECT 26.265 2.122 26.351 2.453 ;
      RECT 26.255 2.097 26.265 2.443 ;
      RECT 26.185 2.065 26.255 2.435 ;
      RECT 26.16 2.025 26.185 2.427 ;
      RECT 26.14 2.007 26.16 2.421 ;
      RECT 26.13 1.997 26.14 2.418 ;
      RECT 26.12 1.99 26.13 2.416 ;
      RECT 26.1 1.977 26.12 2.413 ;
      RECT 26.09 1.967 26.1 2.41 ;
      RECT 26.08 1.96 26.09 2.408 ;
      RECT 26.03 1.952 26.08 2.402 ;
      RECT 26.02 1.95 26.03 2.396 ;
      RECT 25.99 1.95 26.015 2.393 ;
      RECT 25.961 1.95 25.99 2.388 ;
      RECT 25.875 1.95 25.961 2.378 ;
      RECT 25.845 1.95 25.875 2.365 ;
      RECT 25.8 1.95 25.825 2.348 ;
      RECT 25.785 1.95 25.795 2.33 ;
      RECT 25.765 1.957 25.785 2.315 ;
      RECT 25.76 1.972 25.765 2.303 ;
      RECT 25.755 1.977 25.76 2.243 ;
      RECT 25.75 1.982 25.755 2.085 ;
      RECT 25.745 1.985 25.75 2.003 ;
      RECT 26.01 2.67 26.096 2.991 ;
      RECT 26.01 2.67 26.13 2.984 ;
      RECT 25.96 2.67 26.13 2.98 ;
      RECT 25.96 2.672 26.216 2.978 ;
      RECT 25.96 2.674 26.24 2.972 ;
      RECT 25.96 2.681 26.25 2.971 ;
      RECT 25.96 2.69 26.255 2.968 ;
      RECT 25.96 2.696 26.26 2.963 ;
      RECT 25.96 2.74 26.265 2.96 ;
      RECT 25.96 2.832 26.27 2.957 ;
      RECT 25.485 3.275 25.52 3.595 ;
      RECT 26.07 3.46 26.075 3.642 ;
      RECT 26.025 3.342 26.07 3.661 ;
      RECT 26.01 3.319 26.025 3.684 ;
      RECT 26 3.309 26.01 3.694 ;
      RECT 25.98 3.304 26 3.707 ;
      RECT 25.955 3.302 25.98 3.728 ;
      RECT 25.936 3.301 25.955 3.74 ;
      RECT 25.85 3.298 25.936 3.74 ;
      RECT 25.78 3.293 25.85 3.728 ;
      RECT 25.705 3.289 25.78 3.703 ;
      RECT 25.64 3.285 25.705 3.67 ;
      RECT 25.57 3.282 25.64 3.63 ;
      RECT 25.54 3.278 25.57 3.605 ;
      RECT 25.52 3.276 25.54 3.598 ;
      RECT 25.436 3.274 25.485 3.596 ;
      RECT 25.35 3.271 25.436 3.597 ;
      RECT 25.275 3.27 25.35 3.599 ;
      RECT 25.19 3.27 25.275 3.625 ;
      RECT 25.113 3.271 25.19 3.65 ;
      RECT 25.027 3.272 25.113 3.65 ;
      RECT 24.941 3.272 25.027 3.65 ;
      RECT 24.855 3.273 24.941 3.65 ;
      RECT 24.835 3.274 24.855 3.642 ;
      RECT 24.82 3.28 24.835 3.627 ;
      RECT 24.785 3.3 24.82 3.607 ;
      RECT 24.775 3.32 24.785 3.589 ;
      RECT 25.745 2.625 25.75 2.895 ;
      RECT 25.74 2.616 25.745 2.9 ;
      RECT 25.73 2.606 25.74 2.912 ;
      RECT 25.725 2.595 25.73 2.923 ;
      RECT 25.705 2.589 25.725 2.941 ;
      RECT 25.66 2.586 25.705 2.99 ;
      RECT 25.645 2.585 25.66 3.035 ;
      RECT 25.64 2.585 25.645 3.048 ;
      RECT 25.63 2.585 25.64 3.06 ;
      RECT 25.625 2.586 25.63 3.075 ;
      RECT 25.605 2.594 25.625 3.08 ;
      RECT 25.575 2.61 25.605 3.08 ;
      RECT 25.565 2.622 25.57 3.08 ;
      RECT 25.53 2.637 25.565 3.08 ;
      RECT 25.5 2.657 25.53 3.08 ;
      RECT 25.49 2.682 25.5 3.08 ;
      RECT 25.485 2.71 25.49 3.08 ;
      RECT 25.48 2.74 25.485 3.08 ;
      RECT 25.475 2.757 25.48 3.08 ;
      RECT 25.465 2.785 25.475 3.08 ;
      RECT 25.455 2.82 25.465 3.08 ;
      RECT 25.45 2.855 25.455 3.08 ;
      RECT 25.57 2.62 25.575 3.08 ;
      RECT 25.085 2.722 25.27 2.895 ;
      RECT 25.045 2.64 25.23 2.893 ;
      RECT 25.006 2.645 25.23 2.889 ;
      RECT 24.92 2.654 25.23 2.884 ;
      RECT 24.836 2.67 25.235 2.879 ;
      RECT 24.75 2.69 25.26 2.873 ;
      RECT 24.75 2.71 25.265 2.873 ;
      RECT 24.836 2.68 25.26 2.879 ;
      RECT 24.92 2.655 25.235 2.884 ;
      RECT 25.085 2.637 25.23 2.895 ;
      RECT 25.085 2.632 25.185 2.895 ;
      RECT 25.171 2.626 25.185 2.895 ;
      RECT 24.56 1.95 24.565 2.349 ;
      RECT 24.305 1.95 24.34 2.347 ;
      RECT 23.9 1.985 23.905 2.341 ;
      RECT 24.645 1.988 24.65 2.243 ;
      RECT 24.64 1.986 24.645 2.249 ;
      RECT 24.635 1.985 24.64 2.256 ;
      RECT 24.61 1.978 24.635 2.28 ;
      RECT 24.605 1.971 24.61 2.304 ;
      RECT 24.6 1.967 24.605 2.313 ;
      RECT 24.59 1.962 24.6 2.326 ;
      RECT 24.585 1.959 24.59 2.335 ;
      RECT 24.58 1.957 24.585 2.34 ;
      RECT 24.565 1.953 24.58 2.35 ;
      RECT 24.55 1.947 24.56 2.349 ;
      RECT 24.512 1.945 24.55 2.349 ;
      RECT 24.426 1.947 24.512 2.349 ;
      RECT 24.34 1.949 24.426 2.348 ;
      RECT 24.269 1.95 24.305 2.347 ;
      RECT 24.183 1.952 24.269 2.347 ;
      RECT 24.097 1.954 24.183 2.346 ;
      RECT 24.011 1.956 24.097 2.346 ;
      RECT 23.925 1.959 24.011 2.345 ;
      RECT 23.915 1.965 23.925 2.344 ;
      RECT 23.905 1.977 23.915 2.342 ;
      RECT 23.845 2.012 23.9 2.338 ;
      RECT 23.84 2.042 23.845 2.1 ;
      RECT 24.585 3.122 24.6 3.315 ;
      RECT 24.58 3.09 24.585 3.315 ;
      RECT 24.57 3.065 24.58 3.315 ;
      RECT 24.565 3.037 24.57 3.315 ;
      RECT 24.535 2.96 24.565 3.315 ;
      RECT 24.51 2.842 24.535 3.315 ;
      RECT 24.505 2.78 24.51 3.315 ;
      RECT 24.495 2.767 24.505 3.315 ;
      RECT 24.475 2.757 24.495 3.315 ;
      RECT 24.46 2.74 24.475 3.315 ;
      RECT 24.43 2.728 24.46 3.315 ;
      RECT 24.425 2.727 24.43 3.26 ;
      RECT 24.42 2.727 24.425 3.218 ;
      RECT 24.405 2.726 24.42 3.17 ;
      RECT 24.39 2.726 24.405 3.108 ;
      RECT 24.37 2.726 24.39 3.068 ;
      RECT 24.365 2.726 24.37 3.053 ;
      RECT 24.34 2.725 24.365 3.048 ;
      RECT 24.27 2.724 24.34 3.035 ;
      RECT 24.255 2.723 24.27 3.02 ;
      RECT 24.225 2.722 24.255 3.003 ;
      RECT 24.22 2.722 24.225 2.988 ;
      RECT 24.17 2.721 24.22 2.968 ;
      RECT 24.105 2.72 24.17 2.923 ;
      RECT 24.1 2.72 24.105 2.895 ;
      RECT 24.185 3.257 24.19 3.514 ;
      RECT 24.165 3.176 24.185 3.531 ;
      RECT 24.145 3.17 24.165 3.56 ;
      RECT 24.085 3.157 24.145 3.58 ;
      RECT 24.04 3.141 24.085 3.581 ;
      RECT 23.956 3.129 24.04 3.569 ;
      RECT 23.87 3.116 23.956 3.553 ;
      RECT 23.86 3.109 23.87 3.545 ;
      RECT 23.815 3.106 23.86 3.485 ;
      RECT 23.795 3.102 23.815 3.4 ;
      RECT 23.78 3.1 23.795 3.353 ;
      RECT 23.75 3.097 23.78 3.323 ;
      RECT 23.715 3.093 23.75 3.3 ;
      RECT 23.672 3.088 23.715 3.288 ;
      RECT 23.586 3.079 23.672 3.297 ;
      RECT 23.5 3.068 23.586 3.309 ;
      RECT 23.435 3.059 23.5 3.318 ;
      RECT 23.415 3.05 23.435 3.323 ;
      RECT 23.41 3.043 23.415 3.325 ;
      RECT 23.37 3.028 23.41 3.322 ;
      RECT 23.35 3.007 23.37 3.317 ;
      RECT 23.335 2.995 23.35 3.31 ;
      RECT 23.33 2.987 23.335 3.303 ;
      RECT 23.315 2.967 23.33 3.296 ;
      RECT 23.31 2.83 23.315 3.29 ;
      RECT 23.23 2.719 23.31 3.262 ;
      RECT 23.221 2.712 23.23 3.228 ;
      RECT 23.135 2.706 23.221 3.153 ;
      RECT 23.11 2.697 23.135 3.065 ;
      RECT 23.08 2.692 23.11 3.04 ;
      RECT 23.015 2.701 23.08 3.025 ;
      RECT 22.995 2.717 23.015 3 ;
      RECT 22.985 2.723 22.995 2.948 ;
      RECT 22.965 2.745 22.985 2.83 ;
      RECT 23.62 2.71 23.79 2.895 ;
      RECT 23.62 2.71 23.825 2.893 ;
      RECT 23.67 2.62 23.84 2.884 ;
      RECT 23.62 2.777 23.845 2.877 ;
      RECT 23.635 2.655 23.84 2.884 ;
      RECT 22.835 3.388 22.9 3.831 ;
      RECT 22.775 3.413 22.9 3.829 ;
      RECT 22.775 3.413 22.955 3.823 ;
      RECT 22.76 3.438 22.955 3.822 ;
      RECT 22.9 3.375 22.975 3.819 ;
      RECT 22.835 3.4 23.055 3.813 ;
      RECT 22.76 3.439 23.1 3.807 ;
      RECT 22.745 3.466 23.1 3.798 ;
      RECT 22.76 3.459 23.12 3.79 ;
      RECT 22.745 3.468 23.125 3.773 ;
      RECT 22.74 3.485 23.125 3.6 ;
      RECT 22.745 2.207 22.78 2.445 ;
      RECT 22.745 2.207 22.81 2.444 ;
      RECT 22.745 2.207 22.925 2.44 ;
      RECT 22.745 2.207 22.98 2.418 ;
      RECT 22.755 2.15 23.035 2.318 ;
      RECT 22.86 1.99 22.89 2.441 ;
      RECT 22.89 1.985 23.07 2.198 ;
      RECT 22.76 2.126 23.07 2.198 ;
      RECT 22.81 2.022 22.86 2.442 ;
      RECT 22.78 2.078 23.07 2.198 ;
      RECT 21.65 5.02 21.82 6.49 ;
      RECT 21.65 6.315 21.825 6.485 ;
      RECT 21.28 1.74 21.45 2.93 ;
      RECT 21.28 1.74 21.75 1.91 ;
      RECT 21.28 6.97 21.75 7.14 ;
      RECT 21.28 5.95 21.45 7.14 ;
      RECT 20.29 1.74 20.46 2.93 ;
      RECT 20.29 1.74 20.76 1.91 ;
      RECT 20.29 6.97 20.76 7.14 ;
      RECT 20.29 5.95 20.46 7.14 ;
      RECT 18.44 2.635 18.61 3.865 ;
      RECT 18.495 0.855 18.665 2.805 ;
      RECT 18.44 0.575 18.61 1.025 ;
      RECT 18.44 7.855 18.61 8.305 ;
      RECT 18.495 6.075 18.665 8.025 ;
      RECT 18.44 5.015 18.61 6.245 ;
      RECT 17.92 0.575 18.09 3.865 ;
      RECT 17.92 2.075 18.325 2.405 ;
      RECT 17.92 1.235 18.325 1.565 ;
      RECT 17.92 5.015 18.09 8.305 ;
      RECT 17.92 7.315 18.325 7.645 ;
      RECT 17.92 6.475 18.325 6.805 ;
      RECT 16.02 3.392 16.035 3.443 ;
      RECT 16.015 3.372 16.02 3.49 ;
      RECT 16 3.362 16.015 3.558 ;
      RECT 15.975 3.342 16 3.613 ;
      RECT 15.935 3.327 15.975 3.633 ;
      RECT 15.89 3.321 15.935 3.661 ;
      RECT 15.82 3.311 15.89 3.678 ;
      RECT 15.8 3.303 15.82 3.678 ;
      RECT 15.74 3.297 15.8 3.67 ;
      RECT 15.681 3.288 15.74 3.658 ;
      RECT 15.595 3.277 15.681 3.641 ;
      RECT 15.573 3.268 15.595 3.629 ;
      RECT 15.487 3.261 15.573 3.616 ;
      RECT 15.401 3.248 15.487 3.597 ;
      RECT 15.315 3.236 15.401 3.577 ;
      RECT 15.285 3.225 15.315 3.564 ;
      RECT 15.235 3.211 15.285 3.556 ;
      RECT 15.215 3.2 15.235 3.548 ;
      RECT 15.166 3.189 15.215 3.54 ;
      RECT 15.08 3.168 15.166 3.525 ;
      RECT 15.035 3.155 15.08 3.51 ;
      RECT 14.99 3.155 15.035 3.49 ;
      RECT 14.935 3.155 14.99 3.425 ;
      RECT 14.91 3.155 14.935 3.348 ;
      RECT 15.435 2.892 15.605 3.075 ;
      RECT 15.435 2.892 15.62 3.033 ;
      RECT 15.435 2.892 15.625 2.975 ;
      RECT 15.495 2.66 15.63 2.951 ;
      RECT 15.495 2.664 15.635 2.934 ;
      RECT 15.44 2.827 15.635 2.934 ;
      RECT 15.465 2.672 15.605 3.075 ;
      RECT 15.465 2.676 15.645 2.875 ;
      RECT 15.45 2.762 15.645 2.875 ;
      RECT 15.46 2.692 15.605 3.075 ;
      RECT 15.46 2.695 15.655 2.788 ;
      RECT 15.455 2.712 15.655 2.788 ;
      RECT 15.225 1.932 15.395 2.415 ;
      RECT 15.22 1.927 15.37 2.405 ;
      RECT 15.22 1.934 15.4 2.399 ;
      RECT 15.21 1.928 15.37 2.378 ;
      RECT 15.21 1.944 15.415 2.337 ;
      RECT 15.18 1.929 15.37 2.3 ;
      RECT 15.18 1.959 15.425 2.24 ;
      RECT 15.175 1.931 15.37 2.238 ;
      RECT 15.155 1.94 15.4 2.195 ;
      RECT 15.13 1.956 15.415 2.107 ;
      RECT 15.13 1.975 15.44 2.098 ;
      RECT 15.125 2.012 15.44 2.05 ;
      RECT 15.13 1.992 15.445 2.018 ;
      RECT 15.225 1.926 15.335 2.415 ;
      RECT 15.311 1.925 15.335 2.415 ;
      RECT 14.545 2.71 14.55 2.921 ;
      RECT 15.145 2.71 15.15 2.895 ;
      RECT 15.21 2.75 15.215 2.863 ;
      RECT 15.205 2.742 15.21 2.869 ;
      RECT 15.2 2.732 15.205 2.877 ;
      RECT 15.195 2.722 15.2 2.886 ;
      RECT 15.19 2.712 15.195 2.89 ;
      RECT 15.15 2.71 15.19 2.893 ;
      RECT 15.122 2.709 15.145 2.897 ;
      RECT 15.036 2.706 15.122 2.904 ;
      RECT 14.95 2.702 15.036 2.915 ;
      RECT 14.93 2.7 14.95 2.921 ;
      RECT 14.912 2.699 14.93 2.924 ;
      RECT 14.826 2.697 14.912 2.931 ;
      RECT 14.74 2.692 14.826 2.944 ;
      RECT 14.721 2.689 14.74 2.949 ;
      RECT 14.635 2.687 14.721 2.94 ;
      RECT 14.625 2.687 14.635 2.933 ;
      RECT 14.55 2.7 14.625 2.927 ;
      RECT 14.535 2.711 14.545 2.921 ;
      RECT 14.525 2.713 14.535 2.92 ;
      RECT 14.515 2.717 14.525 2.916 ;
      RECT 14.51 2.72 14.515 2.91 ;
      RECT 14.5 2.722 14.51 2.904 ;
      RECT 14.495 2.725 14.5 2.898 ;
      RECT 14.475 3.311 14.48 3.515 ;
      RECT 14.46 3.298 14.475 3.608 ;
      RECT 14.445 3.279 14.46 3.885 ;
      RECT 14.41 3.245 14.445 3.885 ;
      RECT 14.406 3.215 14.41 3.885 ;
      RECT 14.32 3.097 14.406 3.885 ;
      RECT 14.31 2.972 14.32 3.885 ;
      RECT 14.295 2.94 14.31 3.885 ;
      RECT 14.29 2.915 14.295 3.885 ;
      RECT 14.285 2.905 14.29 3.841 ;
      RECT 14.27 2.877 14.285 3.746 ;
      RECT 14.255 2.843 14.27 3.645 ;
      RECT 14.25 2.821 14.255 3.598 ;
      RECT 14.245 2.81 14.25 3.568 ;
      RECT 14.24 2.8 14.245 3.534 ;
      RECT 14.23 2.787 14.24 3.502 ;
      RECT 14.205 2.763 14.23 3.428 ;
      RECT 14.2 2.743 14.205 3.353 ;
      RECT 14.195 2.737 14.2 3.328 ;
      RECT 14.19 2.732 14.195 3.293 ;
      RECT 14.185 2.727 14.19 3.268 ;
      RECT 14.18 2.725 14.185 3.248 ;
      RECT 14.175 2.725 14.18 3.233 ;
      RECT 14.17 2.725 14.175 3.193 ;
      RECT 14.16 2.725 14.17 3.165 ;
      RECT 14.15 2.725 14.16 3.11 ;
      RECT 14.135 2.725 14.15 3.048 ;
      RECT 14.13 2.724 14.135 2.993 ;
      RECT 14.115 2.723 14.13 2.973 ;
      RECT 14.055 2.721 14.115 2.947 ;
      RECT 14.02 2.722 14.055 2.927 ;
      RECT 14.015 2.724 14.02 2.917 ;
      RECT 14.005 2.743 14.015 2.907 ;
      RECT 14 2.77 14.005 2.838 ;
      RECT 14.115 2.195 14.285 2.44 ;
      RECT 14.15 1.966 14.285 2.44 ;
      RECT 14.15 1.968 14.295 2.435 ;
      RECT 14.15 1.97 14.32 2.423 ;
      RECT 14.15 1.973 14.345 2.405 ;
      RECT 14.15 1.978 14.395 2.378 ;
      RECT 14.15 1.983 14.415 2.343 ;
      RECT 14.13 1.985 14.425 2.318 ;
      RECT 14.12 2.08 14.425 2.318 ;
      RECT 14.15 1.965 14.26 2.44 ;
      RECT 14.16 1.962 14.255 2.44 ;
      RECT 13.68 3.227 13.87 3.585 ;
      RECT 13.68 3.239 13.905 3.584 ;
      RECT 13.68 3.267 13.925 3.582 ;
      RECT 13.68 3.292 13.93 3.581 ;
      RECT 13.68 3.35 13.945 3.58 ;
      RECT 13.665 3.223 13.825 3.565 ;
      RECT 13.645 3.232 13.87 3.518 ;
      RECT 13.62 3.243 13.905 3.455 ;
      RECT 13.62 3.327 13.94 3.455 ;
      RECT 13.62 3.302 13.935 3.455 ;
      RECT 13.68 3.218 13.825 3.585 ;
      RECT 13.766 3.217 13.825 3.585 ;
      RECT 13.766 3.216 13.81 3.585 ;
      RECT 13.68 7.855 13.85 8.305 ;
      RECT 13.735 6.075 13.905 8.025 ;
      RECT 13.68 5.015 13.85 6.245 ;
      RECT 13.16 5.015 13.33 8.305 ;
      RECT 13.16 7.315 13.565 7.645 ;
      RECT 13.16 6.475 13.565 6.805 ;
      RECT 13.465 2.732 13.47 3.11 ;
      RECT 13.46 2.7 13.465 3.11 ;
      RECT 13.455 2.672 13.46 3.11 ;
      RECT 13.45 2.652 13.455 3.11 ;
      RECT 13.395 2.635 13.45 3.11 ;
      RECT 13.355 2.62 13.395 3.11 ;
      RECT 13.3 2.607 13.355 3.11 ;
      RECT 13.265 2.598 13.3 3.11 ;
      RECT 13.261 2.596 13.265 3.109 ;
      RECT 13.175 2.592 13.261 3.092 ;
      RECT 13.09 2.584 13.175 3.055 ;
      RECT 13.08 2.58 13.09 3.028 ;
      RECT 13.07 2.58 13.08 3.01 ;
      RECT 13.06 2.582 13.07 2.993 ;
      RECT 13.055 2.587 13.06 2.979 ;
      RECT 13.05 2.591 13.055 2.966 ;
      RECT 13.04 2.596 13.05 2.95 ;
      RECT 13.025 2.61 13.04 2.925 ;
      RECT 13.02 2.616 13.025 2.905 ;
      RECT 13.015 2.618 13.02 2.898 ;
      RECT 13.01 2.622 13.015 2.773 ;
      RECT 13.19 3.422 13.435 3.885 ;
      RECT 13.11 3.395 13.43 3.881 ;
      RECT 13.04 3.43 13.435 3.874 ;
      RECT 12.83 3.685 13.435 3.87 ;
      RECT 13.01 3.453 13.435 3.87 ;
      RECT 12.85 3.645 13.435 3.87 ;
      RECT 13 3.465 13.435 3.87 ;
      RECT 12.885 3.582 13.435 3.87 ;
      RECT 12.94 3.507 13.435 3.87 ;
      RECT 13.19 3.372 13.43 3.885 ;
      RECT 13.22 3.365 13.43 3.885 ;
      RECT 13.21 3.367 13.43 3.885 ;
      RECT 13.22 3.362 13.35 3.885 ;
      RECT 12.775 1.925 12.861 2.364 ;
      RECT 12.77 1.925 12.861 2.362 ;
      RECT 12.77 1.925 12.93 2.361 ;
      RECT 12.77 1.925 12.96 2.358 ;
      RECT 12.755 1.932 12.96 2.349 ;
      RECT 12.755 1.932 12.965 2.345 ;
      RECT 12.75 1.942 12.965 2.338 ;
      RECT 12.745 1.947 12.965 2.313 ;
      RECT 12.745 1.947 12.98 2.295 ;
      RECT 12.77 1.925 13 2.21 ;
      RECT 12.74 1.952 13 2.208 ;
      RECT 12.75 1.945 13.005 2.146 ;
      RECT 12.74 2.067 13.01 2.129 ;
      RECT 12.725 1.962 13.005 2.08 ;
      RECT 12.72 1.972 13.005 1.98 ;
      RECT 12.8 2.743 12.805 2.82 ;
      RECT 12.79 2.737 12.8 3.01 ;
      RECT 12.78 2.729 12.79 3.031 ;
      RECT 12.77 2.72 12.78 3.053 ;
      RECT 12.765 2.715 12.77 3.07 ;
      RECT 12.725 2.715 12.765 3.11 ;
      RECT 12.705 2.715 12.725 3.165 ;
      RECT 12.7 2.715 12.705 3.193 ;
      RECT 12.69 2.715 12.7 3.208 ;
      RECT 12.655 2.715 12.69 3.25 ;
      RECT 12.65 2.715 12.655 3.293 ;
      RECT 12.64 2.715 12.65 3.308 ;
      RECT 12.625 2.715 12.64 3.328 ;
      RECT 12.61 2.715 12.625 3.355 ;
      RECT 12.605 2.716 12.61 3.373 ;
      RECT 12.585 2.717 12.605 3.38 ;
      RECT 12.53 2.718 12.585 3.4 ;
      RECT 12.52 2.719 12.53 3.414 ;
      RECT 12.515 2.722 12.52 3.413 ;
      RECT 12.475 2.795 12.515 3.411 ;
      RECT 12.46 2.875 12.475 3.409 ;
      RECT 12.435 2.93 12.46 3.407 ;
      RECT 12.42 2.995 12.435 3.406 ;
      RECT 12.375 3.027 12.42 3.403 ;
      RECT 12.29 3.05 12.375 3.398 ;
      RECT 12.265 3.07 12.29 3.393 ;
      RECT 12.195 3.075 12.265 3.389 ;
      RECT 12.175 3.077 12.195 3.386 ;
      RECT 12.09 3.088 12.175 3.38 ;
      RECT 12.085 3.099 12.09 3.375 ;
      RECT 12.075 3.101 12.085 3.375 ;
      RECT 12.04 3.105 12.075 3.373 ;
      RECT 11.99 3.115 12.04 3.36 ;
      RECT 11.97 3.123 11.99 3.345 ;
      RECT 11.89 3.135 11.97 3.328 ;
      RECT 12.055 2.685 12.225 2.895 ;
      RECT 12.171 2.681 12.225 2.895 ;
      RECT 11.976 2.685 12.225 2.886 ;
      RECT 11.976 2.685 12.23 2.875 ;
      RECT 11.89 2.685 12.23 2.866 ;
      RECT 11.89 2.693 12.24 2.81 ;
      RECT 11.89 2.705 12.245 2.723 ;
      RECT 11.89 2.712 12.25 2.715 ;
      RECT 12.085 2.683 12.225 2.895 ;
      RECT 11.84 3.628 12.085 3.96 ;
      RECT 11.835 3.62 11.84 3.957 ;
      RECT 11.805 3.64 12.085 3.938 ;
      RECT 11.785 3.672 12.085 3.911 ;
      RECT 11.835 3.625 12.012 3.957 ;
      RECT 11.835 3.622 11.926 3.957 ;
      RECT 11.775 1.97 11.945 2.39 ;
      RECT 11.77 1.97 11.945 2.388 ;
      RECT 11.77 1.97 11.97 2.378 ;
      RECT 11.77 1.97 11.99 2.353 ;
      RECT 11.765 1.97 11.99 2.348 ;
      RECT 11.765 1.97 12 2.338 ;
      RECT 11.765 1.97 12.005 2.333 ;
      RECT 11.765 1.975 12.01 2.328 ;
      RECT 11.765 2.007 12.025 2.318 ;
      RECT 11.765 2.077 12.05 2.301 ;
      RECT 11.745 2.077 12.05 2.293 ;
      RECT 11.745 2.137 12.06 2.27 ;
      RECT 11.745 2.177 12.07 2.215 ;
      RECT 11.73 1.97 12.005 2.195 ;
      RECT 11.72 1.985 12.01 2.093 ;
      RECT 11.31 3.375 11.48 3.9 ;
      RECT 11.305 3.375 11.48 3.893 ;
      RECT 11.295 3.375 11.485 3.858 ;
      RECT 11.29 3.385 11.485 3.83 ;
      RECT 11.285 3.405 11.485 3.813 ;
      RECT 11.295 3.38 11.49 3.803 ;
      RECT 11.28 3.425 11.49 3.795 ;
      RECT 11.275 3.445 11.49 3.78 ;
      RECT 11.27 3.475 11.49 3.77 ;
      RECT 11.26 3.52 11.49 3.745 ;
      RECT 11.29 3.39 11.495 3.728 ;
      RECT 11.255 3.572 11.495 3.723 ;
      RECT 11.29 3.4 11.5 3.693 ;
      RECT 11.25 3.605 11.5 3.69 ;
      RECT 11.245 3.63 11.5 3.67 ;
      RECT 11.285 3.417 11.51 3.61 ;
      RECT 11.28 3.439 11.52 3.503 ;
      RECT 11.23 2.686 11.245 2.955 ;
      RECT 11.185 2.67 11.23 3 ;
      RECT 11.18 2.658 11.185 3.05 ;
      RECT 11.17 2.654 11.18 3.083 ;
      RECT 11.165 2.651 11.17 3.111 ;
      RECT 11.15 2.653 11.165 3.153 ;
      RECT 11.145 2.657 11.15 3.193 ;
      RECT 11.125 2.662 11.145 3.245 ;
      RECT 11.121 2.667 11.125 3.302 ;
      RECT 11.035 2.686 11.121 3.339 ;
      RECT 11.025 2.707 11.035 3.375 ;
      RECT 11.02 2.715 11.025 3.376 ;
      RECT 11.015 2.757 11.02 3.377 ;
      RECT 11 2.845 11.015 3.378 ;
      RECT 10.99 2.995 11 3.38 ;
      RECT 10.985 3.04 10.99 3.382 ;
      RECT 10.95 3.082 10.985 3.385 ;
      RECT 10.945 3.1 10.95 3.388 ;
      RECT 10.868 3.106 10.945 3.394 ;
      RECT 10.782 3.12 10.868 3.407 ;
      RECT 10.696 3.134 10.782 3.421 ;
      RECT 10.61 3.148 10.696 3.434 ;
      RECT 10.55 3.16 10.61 3.446 ;
      RECT 10.525 3.167 10.55 3.453 ;
      RECT 10.511 3.17 10.525 3.458 ;
      RECT 10.425 3.178 10.511 3.474 ;
      RECT 10.42 3.185 10.425 3.489 ;
      RECT 10.396 3.185 10.42 3.496 ;
      RECT 10.31 3.188 10.396 3.524 ;
      RECT 10.225 3.192 10.31 3.568 ;
      RECT 10.16 3.196 10.225 3.605 ;
      RECT 10.135 3.199 10.16 3.621 ;
      RECT 10.06 3.212 10.135 3.625 ;
      RECT 10.035 3.23 10.06 3.629 ;
      RECT 10.025 3.237 10.035 3.631 ;
      RECT 10.01 3.24 10.025 3.632 ;
      RECT 9.95 3.252 10.01 3.636 ;
      RECT 9.94 3.266 9.95 3.64 ;
      RECT 9.885 3.276 9.94 3.628 ;
      RECT 9.86 3.297 9.885 3.611 ;
      RECT 9.84 3.317 9.86 3.602 ;
      RECT 9.835 3.33 9.84 3.597 ;
      RECT 9.82 3.342 9.835 3.593 ;
      RECT 11.055 1.997 11.06 2.02 ;
      RECT 11.05 1.988 11.055 2.06 ;
      RECT 11.045 1.986 11.05 2.103 ;
      RECT 11.04 1.977 11.045 2.138 ;
      RECT 11.035 1.967 11.04 2.21 ;
      RECT 11.03 1.957 11.035 2.275 ;
      RECT 11.025 1.954 11.03 2.315 ;
      RECT 11 1.948 11.025 2.405 ;
      RECT 10.965 1.936 11 2.43 ;
      RECT 10.955 1.927 10.965 2.43 ;
      RECT 10.82 1.925 10.83 2.413 ;
      RECT 10.81 1.925 10.82 2.38 ;
      RECT 10.805 1.925 10.81 2.355 ;
      RECT 10.8 1.925 10.805 2.343 ;
      RECT 10.795 1.925 10.8 2.325 ;
      RECT 10.785 1.925 10.795 2.29 ;
      RECT 10.78 1.927 10.785 2.268 ;
      RECT 10.775 1.933 10.78 2.253 ;
      RECT 10.77 1.939 10.775 2.238 ;
      RECT 10.755 1.951 10.77 2.211 ;
      RECT 10.75 1.962 10.755 2.179 ;
      RECT 10.745 1.972 10.75 2.163 ;
      RECT 10.735 1.98 10.745 2.132 ;
      RECT 10.73 1.99 10.735 2.106 ;
      RECT 10.725 2.047 10.73 2.089 ;
      RECT 10.83 1.925 10.955 2.43 ;
      RECT 10.545 2.612 10.805 2.91 ;
      RECT 10.54 2.619 10.805 2.908 ;
      RECT 10.545 2.614 10.82 2.903 ;
      RECT 10.535 2.627 10.82 2.9 ;
      RECT 10.535 2.632 10.825 2.893 ;
      RECT 10.53 2.64 10.825 2.89 ;
      RECT 10.53 2.657 10.83 2.688 ;
      RECT 10.545 2.609 10.776 2.91 ;
      RECT 10.6 2.608 10.776 2.91 ;
      RECT 10.6 2.605 10.69 2.91 ;
      RECT 10.6 2.602 10.686 2.91 ;
      RECT 10.29 2.875 10.295 2.888 ;
      RECT 10.285 2.842 10.29 2.893 ;
      RECT 10.28 2.797 10.285 2.9 ;
      RECT 10.275 2.752 10.28 2.908 ;
      RECT 10.27 2.72 10.275 2.916 ;
      RECT 10.265 2.68 10.27 2.917 ;
      RECT 10.25 2.66 10.265 2.919 ;
      RECT 10.175 2.642 10.25 2.931 ;
      RECT 10.165 2.635 10.175 2.942 ;
      RECT 10.16 2.635 10.165 2.944 ;
      RECT 10.13 2.641 10.16 2.948 ;
      RECT 10.09 2.654 10.13 2.948 ;
      RECT 10.065 2.665 10.09 2.934 ;
      RECT 10.05 2.671 10.065 2.917 ;
      RECT 10.04 2.673 10.05 2.908 ;
      RECT 10.035 2.674 10.04 2.903 ;
      RECT 10.03 2.675 10.035 2.898 ;
      RECT 10.025 2.676 10.03 2.895 ;
      RECT 10 2.681 10.025 2.885 ;
      RECT 9.99 2.697 10 2.872 ;
      RECT 9.985 2.717 9.99 2.867 ;
      RECT 9.995 2.11 10 2.306 ;
      RECT 9.98 2.074 9.995 2.308 ;
      RECT 9.97 2.056 9.98 2.313 ;
      RECT 9.96 2.042 9.97 2.317 ;
      RECT 9.915 2.026 9.96 2.327 ;
      RECT 9.91 2.016 9.915 2.336 ;
      RECT 9.865 2.005 9.91 2.342 ;
      RECT 9.86 1.993 9.865 2.349 ;
      RECT 9.845 1.988 9.86 2.353 ;
      RECT 9.83 1.98 9.845 2.358 ;
      RECT 9.82 1.973 9.83 2.363 ;
      RECT 9.81 1.97 9.82 2.368 ;
      RECT 9.8 1.97 9.81 2.369 ;
      RECT 9.795 1.967 9.8 2.368 ;
      RECT 9.76 1.962 9.785 2.367 ;
      RECT 9.736 1.958 9.76 2.366 ;
      RECT 9.65 1.949 9.736 2.363 ;
      RECT 9.635 1.941 9.65 2.36 ;
      RECT 9.613 1.94 9.635 2.359 ;
      RECT 9.527 1.94 9.613 2.357 ;
      RECT 9.441 1.94 9.527 2.355 ;
      RECT 9.355 1.94 9.441 2.352 ;
      RECT 9.345 1.94 9.355 2.343 ;
      RECT 9.315 1.94 9.345 2.303 ;
      RECT 9.305 1.95 9.315 2.258 ;
      RECT 9.3 1.99 9.305 2.243 ;
      RECT 9.295 2.005 9.3 2.23 ;
      RECT 9.265 2.085 9.295 2.192 ;
      RECT 9.785 1.965 9.795 2.368 ;
      RECT 9.61 2.73 9.625 3.335 ;
      RECT 9.615 2.725 9.625 3.335 ;
      RECT 9.78 2.725 9.785 2.908 ;
      RECT 9.77 2.725 9.78 2.938 ;
      RECT 9.755 2.725 9.77 2.998 ;
      RECT 9.75 2.725 9.755 3.043 ;
      RECT 9.745 2.725 9.75 3.073 ;
      RECT 9.74 2.725 9.745 3.093 ;
      RECT 9.73 2.725 9.74 3.128 ;
      RECT 9.715 2.725 9.73 3.16 ;
      RECT 9.67 2.725 9.715 3.188 ;
      RECT 9.665 2.725 9.67 3.218 ;
      RECT 9.66 2.725 9.665 3.23 ;
      RECT 9.655 2.725 9.66 3.238 ;
      RECT 9.645 2.725 9.655 3.253 ;
      RECT 9.64 2.725 9.645 3.275 ;
      RECT 9.63 2.725 9.64 3.298 ;
      RECT 9.625 2.725 9.63 3.318 ;
      RECT 9.59 2.74 9.61 3.335 ;
      RECT 9.565 2.757 9.59 3.335 ;
      RECT 9.56 2.767 9.565 3.335 ;
      RECT 9.53 2.782 9.56 3.335 ;
      RECT 9.455 2.824 9.53 3.335 ;
      RECT 9.45 2.855 9.455 3.318 ;
      RECT 9.445 2.859 9.45 3.3 ;
      RECT 9.44 2.863 9.445 3.263 ;
      RECT 9.435 3.047 9.44 3.23 ;
      RECT 8.92 3.236 9.006 3.801 ;
      RECT 8.875 3.238 9.04 3.795 ;
      RECT 9.006 3.235 9.04 3.795 ;
      RECT 8.92 3.237 9.125 3.789 ;
      RECT 8.875 3.247 9.135 3.785 ;
      RECT 8.85 3.239 9.125 3.781 ;
      RECT 8.845 3.242 9.125 3.776 ;
      RECT 8.82 3.257 9.135 3.77 ;
      RECT 8.82 3.282 9.175 3.765 ;
      RECT 8.78 3.29 9.175 3.74 ;
      RECT 8.78 3.317 9.19 3.738 ;
      RECT 8.78 3.347 9.2 3.725 ;
      RECT 8.775 3.492 9.2 3.713 ;
      RECT 8.78 3.421 9.22 3.71 ;
      RECT 8.78 3.478 9.225 3.518 ;
      RECT 8.97 2.757 9.14 2.935 ;
      RECT 8.92 2.696 8.97 2.92 ;
      RECT 8.655 2.676 8.92 2.905 ;
      RECT 8.615 2.74 9.09 2.905 ;
      RECT 8.615 2.73 9.045 2.905 ;
      RECT 8.615 2.727 9.035 2.905 ;
      RECT 8.615 2.715 9.025 2.905 ;
      RECT 8.615 2.7 8.97 2.905 ;
      RECT 8.655 2.672 8.856 2.905 ;
      RECT 8.665 2.65 8.856 2.905 ;
      RECT 8.69 2.635 8.77 2.905 ;
      RECT 8.445 3.165 8.565 3.61 ;
      RECT 8.43 3.165 8.565 3.609 ;
      RECT 8.385 3.187 8.565 3.604 ;
      RECT 8.345 3.236 8.565 3.598 ;
      RECT 8.345 3.236 8.57 3.573 ;
      RECT 8.345 3.236 8.59 3.463 ;
      RECT 8.34 3.266 8.59 3.46 ;
      RECT 8.43 3.165 8.6 3.355 ;
      RECT 8.09 1.95 8.095 2.395 ;
      RECT 7.9 1.95 7.92 2.36 ;
      RECT 7.87 1.95 7.875 2.335 ;
      RECT 8.55 2.257 8.565 2.445 ;
      RECT 8.545 2.242 8.55 2.451 ;
      RECT 8.525 2.215 8.545 2.454 ;
      RECT 8.475 2.182 8.525 2.463 ;
      RECT 8.445 2.162 8.475 2.467 ;
      RECT 8.426 2.15 8.445 2.463 ;
      RECT 8.34 2.122 8.426 2.453 ;
      RECT 8.33 2.097 8.34 2.443 ;
      RECT 8.26 2.065 8.33 2.435 ;
      RECT 8.235 2.025 8.26 2.427 ;
      RECT 8.215 2.007 8.235 2.421 ;
      RECT 8.205 1.997 8.215 2.418 ;
      RECT 8.195 1.99 8.205 2.416 ;
      RECT 8.175 1.977 8.195 2.413 ;
      RECT 8.165 1.967 8.175 2.41 ;
      RECT 8.155 1.96 8.165 2.408 ;
      RECT 8.105 1.952 8.155 2.402 ;
      RECT 8.095 1.95 8.105 2.396 ;
      RECT 8.065 1.95 8.09 2.393 ;
      RECT 8.036 1.95 8.065 2.388 ;
      RECT 7.95 1.95 8.036 2.378 ;
      RECT 7.92 1.95 7.95 2.365 ;
      RECT 7.875 1.95 7.9 2.348 ;
      RECT 7.86 1.95 7.87 2.33 ;
      RECT 7.84 1.957 7.86 2.315 ;
      RECT 7.835 1.972 7.84 2.303 ;
      RECT 7.83 1.977 7.835 2.243 ;
      RECT 7.825 1.982 7.83 2.085 ;
      RECT 7.82 1.985 7.825 2.003 ;
      RECT 8.085 2.67 8.171 2.991 ;
      RECT 8.085 2.67 8.205 2.984 ;
      RECT 8.035 2.67 8.205 2.98 ;
      RECT 8.035 2.672 8.291 2.978 ;
      RECT 8.035 2.674 8.315 2.972 ;
      RECT 8.035 2.681 8.325 2.971 ;
      RECT 8.035 2.69 8.33 2.968 ;
      RECT 8.035 2.696 8.335 2.963 ;
      RECT 8.035 2.74 8.34 2.96 ;
      RECT 8.035 2.832 8.345 2.957 ;
      RECT 7.56 3.275 7.595 3.595 ;
      RECT 8.145 3.46 8.15 3.642 ;
      RECT 8.1 3.342 8.145 3.661 ;
      RECT 8.085 3.319 8.1 3.684 ;
      RECT 8.075 3.309 8.085 3.694 ;
      RECT 8.055 3.304 8.075 3.707 ;
      RECT 8.03 3.302 8.055 3.728 ;
      RECT 8.011 3.301 8.03 3.74 ;
      RECT 7.925 3.298 8.011 3.74 ;
      RECT 7.855 3.293 7.925 3.728 ;
      RECT 7.78 3.289 7.855 3.703 ;
      RECT 7.715 3.285 7.78 3.67 ;
      RECT 7.645 3.282 7.715 3.63 ;
      RECT 7.615 3.278 7.645 3.605 ;
      RECT 7.595 3.276 7.615 3.598 ;
      RECT 7.511 3.274 7.56 3.596 ;
      RECT 7.425 3.271 7.511 3.597 ;
      RECT 7.35 3.27 7.425 3.599 ;
      RECT 7.265 3.27 7.35 3.625 ;
      RECT 7.188 3.271 7.265 3.65 ;
      RECT 7.102 3.272 7.188 3.65 ;
      RECT 7.016 3.272 7.102 3.65 ;
      RECT 6.93 3.273 7.016 3.65 ;
      RECT 6.91 3.274 6.93 3.642 ;
      RECT 6.895 3.28 6.91 3.627 ;
      RECT 6.86 3.3 6.895 3.607 ;
      RECT 6.85 3.32 6.86 3.589 ;
      RECT 7.82 2.625 7.825 2.895 ;
      RECT 7.815 2.616 7.82 2.9 ;
      RECT 7.805 2.606 7.815 2.912 ;
      RECT 7.8 2.595 7.805 2.923 ;
      RECT 7.78 2.589 7.8 2.941 ;
      RECT 7.735 2.586 7.78 2.99 ;
      RECT 7.72 2.585 7.735 3.035 ;
      RECT 7.715 2.585 7.72 3.048 ;
      RECT 7.705 2.585 7.715 3.06 ;
      RECT 7.7 2.586 7.705 3.075 ;
      RECT 7.68 2.594 7.7 3.08 ;
      RECT 7.65 2.61 7.68 3.08 ;
      RECT 7.64 2.622 7.645 3.08 ;
      RECT 7.605 2.637 7.64 3.08 ;
      RECT 7.575 2.657 7.605 3.08 ;
      RECT 7.565 2.682 7.575 3.08 ;
      RECT 7.56 2.71 7.565 3.08 ;
      RECT 7.555 2.74 7.56 3.08 ;
      RECT 7.55 2.757 7.555 3.08 ;
      RECT 7.54 2.785 7.55 3.08 ;
      RECT 7.53 2.82 7.54 3.08 ;
      RECT 7.525 2.855 7.53 3.08 ;
      RECT 7.645 2.62 7.65 3.08 ;
      RECT 7.16 2.722 7.345 2.895 ;
      RECT 7.12 2.64 7.305 2.893 ;
      RECT 7.081 2.645 7.305 2.889 ;
      RECT 6.995 2.654 7.305 2.884 ;
      RECT 6.911 2.67 7.31 2.879 ;
      RECT 6.825 2.69 7.335 2.873 ;
      RECT 6.825 2.71 7.34 2.873 ;
      RECT 6.911 2.68 7.335 2.879 ;
      RECT 6.995 2.655 7.31 2.884 ;
      RECT 7.16 2.637 7.305 2.895 ;
      RECT 7.16 2.632 7.26 2.895 ;
      RECT 7.246 2.626 7.26 2.895 ;
      RECT 6.635 1.95 6.64 2.349 ;
      RECT 6.38 1.95 6.415 2.347 ;
      RECT 5.975 1.985 5.98 2.341 ;
      RECT 6.72 1.988 6.725 2.243 ;
      RECT 6.715 1.986 6.72 2.249 ;
      RECT 6.71 1.985 6.715 2.256 ;
      RECT 6.685 1.978 6.71 2.28 ;
      RECT 6.68 1.971 6.685 2.304 ;
      RECT 6.675 1.967 6.68 2.313 ;
      RECT 6.665 1.962 6.675 2.326 ;
      RECT 6.66 1.959 6.665 2.335 ;
      RECT 6.655 1.957 6.66 2.34 ;
      RECT 6.64 1.953 6.655 2.35 ;
      RECT 6.625 1.947 6.635 2.349 ;
      RECT 6.587 1.945 6.625 2.349 ;
      RECT 6.501 1.947 6.587 2.349 ;
      RECT 6.415 1.949 6.501 2.348 ;
      RECT 6.344 1.95 6.38 2.347 ;
      RECT 6.258 1.952 6.344 2.347 ;
      RECT 6.172 1.954 6.258 2.346 ;
      RECT 6.086 1.956 6.172 2.346 ;
      RECT 6 1.959 6.086 2.345 ;
      RECT 5.99 1.965 6 2.344 ;
      RECT 5.98 1.977 5.99 2.342 ;
      RECT 5.92 2.012 5.975 2.338 ;
      RECT 5.915 2.042 5.92 2.1 ;
      RECT 6.66 3.122 6.675 3.315 ;
      RECT 6.655 3.09 6.66 3.315 ;
      RECT 6.645 3.065 6.655 3.315 ;
      RECT 6.64 3.037 6.645 3.315 ;
      RECT 6.61 2.96 6.64 3.315 ;
      RECT 6.585 2.842 6.61 3.315 ;
      RECT 6.58 2.78 6.585 3.315 ;
      RECT 6.57 2.767 6.58 3.315 ;
      RECT 6.55 2.757 6.57 3.315 ;
      RECT 6.535 2.74 6.55 3.315 ;
      RECT 6.505 2.728 6.535 3.315 ;
      RECT 6.5 2.727 6.505 3.26 ;
      RECT 6.495 2.727 6.5 3.218 ;
      RECT 6.48 2.726 6.495 3.17 ;
      RECT 6.465 2.726 6.48 3.108 ;
      RECT 6.445 2.726 6.465 3.068 ;
      RECT 6.44 2.726 6.445 3.053 ;
      RECT 6.415 2.725 6.44 3.048 ;
      RECT 6.345 2.724 6.415 3.035 ;
      RECT 6.33 2.723 6.345 3.02 ;
      RECT 6.3 2.722 6.33 3.003 ;
      RECT 6.295 2.722 6.3 2.988 ;
      RECT 6.245 2.721 6.295 2.968 ;
      RECT 6.18 2.72 6.245 2.923 ;
      RECT 6.175 2.72 6.18 2.895 ;
      RECT 6.26 3.257 6.265 3.514 ;
      RECT 6.24 3.176 6.26 3.531 ;
      RECT 6.22 3.17 6.24 3.56 ;
      RECT 6.16 3.157 6.22 3.58 ;
      RECT 6.115 3.141 6.16 3.581 ;
      RECT 6.031 3.129 6.115 3.569 ;
      RECT 5.945 3.116 6.031 3.553 ;
      RECT 5.935 3.109 5.945 3.545 ;
      RECT 5.89 3.106 5.935 3.485 ;
      RECT 5.87 3.102 5.89 3.4 ;
      RECT 5.855 3.1 5.87 3.353 ;
      RECT 5.825 3.097 5.855 3.323 ;
      RECT 5.79 3.093 5.825 3.3 ;
      RECT 5.747 3.088 5.79 3.288 ;
      RECT 5.661 3.079 5.747 3.297 ;
      RECT 5.575 3.068 5.661 3.309 ;
      RECT 5.51 3.059 5.575 3.318 ;
      RECT 5.49 3.05 5.51 3.323 ;
      RECT 5.485 3.043 5.49 3.325 ;
      RECT 5.445 3.028 5.485 3.322 ;
      RECT 5.425 3.007 5.445 3.317 ;
      RECT 5.41 2.995 5.425 3.31 ;
      RECT 5.405 2.987 5.41 3.303 ;
      RECT 5.39 2.967 5.405 3.296 ;
      RECT 5.385 2.83 5.39 3.29 ;
      RECT 5.305 2.719 5.385 3.262 ;
      RECT 5.296 2.712 5.305 3.228 ;
      RECT 5.21 2.706 5.296 3.153 ;
      RECT 5.185 2.697 5.21 3.065 ;
      RECT 5.155 2.692 5.185 3.04 ;
      RECT 5.09 2.701 5.155 3.025 ;
      RECT 5.07 2.717 5.09 3 ;
      RECT 5.06 2.723 5.07 2.948 ;
      RECT 5.04 2.745 5.06 2.83 ;
      RECT 5.695 2.71 5.865 2.895 ;
      RECT 5.695 2.71 5.9 2.893 ;
      RECT 5.745 2.62 5.915 2.884 ;
      RECT 5.695 2.777 5.92 2.877 ;
      RECT 5.71 2.655 5.915 2.884 ;
      RECT 4.91 3.388 4.975 3.831 ;
      RECT 4.85 3.413 4.975 3.829 ;
      RECT 4.85 3.413 5.03 3.823 ;
      RECT 4.835 3.438 5.03 3.822 ;
      RECT 4.975 3.375 5.05 3.819 ;
      RECT 4.91 3.4 5.13 3.813 ;
      RECT 4.835 3.439 5.175 3.807 ;
      RECT 4.82 3.466 5.175 3.798 ;
      RECT 4.835 3.459 5.195 3.79 ;
      RECT 4.82 3.468 5.2 3.773 ;
      RECT 4.815 3.485 5.2 3.6 ;
      RECT 4.82 2.207 4.855 2.445 ;
      RECT 4.82 2.207 4.885 2.444 ;
      RECT 4.82 2.207 5 2.44 ;
      RECT 4.82 2.207 5.055 2.418 ;
      RECT 4.83 2.15 5.11 2.318 ;
      RECT 4.935 1.99 4.965 2.441 ;
      RECT 4.965 1.985 5.145 2.198 ;
      RECT 4.835 2.126 5.145 2.198 ;
      RECT 4.885 2.022 4.935 2.442 ;
      RECT 4.855 2.078 5.145 2.198 ;
      RECT 2.65 7.855 2.82 8.305 ;
      RECT 2.705 6.075 2.875 8.025 ;
      RECT 2.65 5.015 2.82 6.245 ;
      RECT 2.13 5.015 2.3 8.305 ;
      RECT 2.13 7.315 2.535 7.645 ;
      RECT 2.13 6.475 2.535 6.805 ;
      RECT 93.35 7.8 93.52 8.31 ;
      RECT 92.36 0.57 92.53 1.08 ;
      RECT 92.36 2.39 92.53 3.86 ;
      RECT 92.36 5.02 92.53 6.49 ;
      RECT 92.36 7.8 92.53 8.31 ;
      RECT 91 0.575 91.17 3.865 ;
      RECT 91 5.015 91.17 8.305 ;
      RECT 90.57 0.575 90.74 1.085 ;
      RECT 90.57 1.655 90.74 3.865 ;
      RECT 90.57 5.015 90.74 7.225 ;
      RECT 90.57 7.795 90.74 8.305 ;
      RECT 86.24 5.015 86.41 8.305 ;
      RECT 85.81 5.015 85.98 7.225 ;
      RECT 85.81 7.795 85.98 8.305 ;
      RECT 75.425 7.8 75.595 8.31 ;
      RECT 74.435 0.57 74.605 1.08 ;
      RECT 74.435 2.39 74.605 3.86 ;
      RECT 74.435 5.02 74.605 6.49 ;
      RECT 74.435 7.8 74.605 8.31 ;
      RECT 73.075 0.575 73.245 3.865 ;
      RECT 73.075 5.015 73.245 8.305 ;
      RECT 72.645 0.575 72.815 1.085 ;
      RECT 72.645 1.655 72.815 3.865 ;
      RECT 72.645 5.015 72.815 7.225 ;
      RECT 72.645 7.795 72.815 8.305 ;
      RECT 68.315 5.015 68.485 8.305 ;
      RECT 67.885 5.015 68.055 7.225 ;
      RECT 67.885 7.795 68.055 8.305 ;
      RECT 57.5 7.8 57.67 8.31 ;
      RECT 56.51 0.57 56.68 1.08 ;
      RECT 56.51 2.39 56.68 3.86 ;
      RECT 56.51 5.02 56.68 6.49 ;
      RECT 56.51 7.8 56.68 8.31 ;
      RECT 55.15 0.575 55.32 3.865 ;
      RECT 55.15 5.015 55.32 8.305 ;
      RECT 54.72 0.575 54.89 1.085 ;
      RECT 54.72 1.655 54.89 3.865 ;
      RECT 54.72 5.015 54.89 7.225 ;
      RECT 54.72 7.795 54.89 8.305 ;
      RECT 50.39 5.015 50.56 8.305 ;
      RECT 49.96 5.015 50.13 7.225 ;
      RECT 49.96 7.795 50.13 8.305 ;
      RECT 39.575 7.8 39.745 8.31 ;
      RECT 38.585 0.57 38.755 1.08 ;
      RECT 38.585 2.39 38.755 3.86 ;
      RECT 38.585 5.02 38.755 6.49 ;
      RECT 38.585 7.8 38.755 8.31 ;
      RECT 37.225 0.575 37.395 3.865 ;
      RECT 37.225 5.015 37.395 8.305 ;
      RECT 36.795 0.575 36.965 1.085 ;
      RECT 36.795 1.655 36.965 3.865 ;
      RECT 36.795 5.015 36.965 7.225 ;
      RECT 36.795 7.795 36.965 8.305 ;
      RECT 32.465 5.015 32.635 8.305 ;
      RECT 32.035 5.015 32.205 7.225 ;
      RECT 32.035 7.795 32.205 8.305 ;
      RECT 21.65 7.8 21.82 8.31 ;
      RECT 20.66 0.57 20.83 1.08 ;
      RECT 20.66 2.39 20.83 3.86 ;
      RECT 20.66 5.02 20.83 6.49 ;
      RECT 20.66 7.8 20.83 8.31 ;
      RECT 19.3 0.575 19.47 3.865 ;
      RECT 19.3 5.015 19.47 8.305 ;
      RECT 18.87 0.575 19.04 1.085 ;
      RECT 18.87 1.655 19.04 3.865 ;
      RECT 18.87 5.015 19.04 7.225 ;
      RECT 18.87 7.795 19.04 8.305 ;
      RECT 14.54 5.015 14.71 8.305 ;
      RECT 14.11 5.015 14.28 7.225 ;
      RECT 14.11 7.795 14.28 8.305 ;
      RECT 3.08 5.015 3.25 7.225 ;
      RECT 3.08 7.795 3.25 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2at_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2at_8_b0r2
  CLASS BLOCK ;
  ORIGIN 0 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2at_8_b0r2 ;
  SIZE 92.575 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 20.335 0.915 20.505 1.085 ;
        RECT 20.33 0.91 20.5 1.08 ;
        RECT 20.33 2.39 20.5 2.56 ;
      LAYER li1 ;
        RECT 20.335 0.915 20.505 1.085 ;
        RECT 20.33 0.57 20.5 1.08 ;
        RECT 20.33 2.39 20.5 3.86 ;
      LAYER met1 ;
        RECT 20.27 2.36 20.56 2.59 ;
        RECT 20.27 0.88 20.56 1.11 ;
        RECT 20.33 0.88 20.5 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 38.26 0.915 38.43 1.085 ;
        RECT 38.255 0.91 38.425 1.08 ;
        RECT 38.255 2.39 38.425 2.56 ;
      LAYER li1 ;
        RECT 38.26 0.915 38.43 1.085 ;
        RECT 38.255 0.57 38.425 1.08 ;
        RECT 38.255 2.39 38.425 3.86 ;
      LAYER met1 ;
        RECT 38.195 2.36 38.485 2.59 ;
        RECT 38.195 0.88 38.485 1.11 ;
        RECT 38.255 0.88 38.425 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 56.185 0.915 56.355 1.085 ;
        RECT 56.18 0.91 56.35 1.08 ;
        RECT 56.18 2.39 56.35 2.56 ;
      LAYER li1 ;
        RECT 56.185 0.915 56.355 1.085 ;
        RECT 56.18 0.57 56.35 1.08 ;
        RECT 56.18 2.39 56.35 3.86 ;
      LAYER met1 ;
        RECT 56.12 2.36 56.41 2.59 ;
        RECT 56.12 0.88 56.41 1.11 ;
        RECT 56.18 0.88 56.35 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 74.11 0.915 74.28 1.085 ;
        RECT 74.105 0.91 74.275 1.08 ;
        RECT 74.105 2.39 74.275 2.56 ;
      LAYER li1 ;
        RECT 74.11 0.915 74.28 1.085 ;
        RECT 74.105 0.57 74.275 1.08 ;
        RECT 74.105 2.39 74.275 3.86 ;
      LAYER met1 ;
        RECT 74.045 2.36 74.335 2.59 ;
        RECT 74.045 0.88 74.335 1.11 ;
        RECT 74.105 0.88 74.275 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 92.035 0.915 92.205 1.085 ;
        RECT 92.03 0.91 92.2 1.08 ;
        RECT 92.03 2.39 92.2 2.56 ;
      LAYER li1 ;
        RECT 92.035 0.915 92.205 1.085 ;
        RECT 92.03 0.57 92.2 1.08 ;
        RECT 92.03 2.39 92.2 3.86 ;
      LAYER met1 ;
        RECT 91.97 2.36 92.26 2.59 ;
        RECT 91.97 0.88 92.26 1.11 ;
        RECT 92.03 0.88 92.2 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 16.18 1.66 16.35 2.935 ;
        RECT 16.18 5.945 16.35 7.22 ;
        RECT 11.42 5.945 11.59 7.22 ;
      LAYER met2 ;
        RECT 16.1 2.705 16.45 3.055 ;
        RECT 16.09 5.84 16.44 6.19 ;
        RECT 16.165 2.705 16.34 6.19 ;
      LAYER met1 ;
        RECT 16.1 2.765 16.58 2.935 ;
        RECT 16.1 2.705 16.45 3.055 ;
        RECT 11.36 5.945 16.58 6.115 ;
        RECT 16.09 5.84 16.44 6.19 ;
        RECT 11.36 5.915 11.65 6.145 ;
      LAYER via1 ;
        RECT 16.19 5.94 16.34 6.09 ;
        RECT 16.2 2.805 16.35 2.955 ;
      LAYER mcon ;
        RECT 11.42 5.945 11.59 6.115 ;
        RECT 16.18 5.945 16.35 6.115 ;
        RECT 16.18 2.765 16.35 2.935 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 34.105 1.66 34.275 2.935 ;
        RECT 34.105 5.945 34.275 7.22 ;
        RECT 29.345 5.945 29.515 7.22 ;
      LAYER met2 ;
        RECT 34.025 2.705 34.375 3.055 ;
        RECT 34.015 5.84 34.365 6.19 ;
        RECT 34.09 2.705 34.265 6.19 ;
      LAYER met1 ;
        RECT 34.025 2.765 34.505 2.935 ;
        RECT 34.025 2.705 34.375 3.055 ;
        RECT 29.285 5.945 34.505 6.115 ;
        RECT 34.015 5.84 34.365 6.19 ;
        RECT 29.285 5.915 29.575 6.145 ;
      LAYER via1 ;
        RECT 34.115 5.94 34.265 6.09 ;
        RECT 34.125 2.805 34.275 2.955 ;
      LAYER mcon ;
        RECT 29.345 5.945 29.515 6.115 ;
        RECT 34.105 5.945 34.275 6.115 ;
        RECT 34.105 2.765 34.275 2.935 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 52.03 1.66 52.2 2.935 ;
        RECT 52.03 5.945 52.2 7.22 ;
        RECT 47.27 5.945 47.44 7.22 ;
      LAYER met2 ;
        RECT 51.95 2.705 52.3 3.055 ;
        RECT 51.94 5.84 52.29 6.19 ;
        RECT 52.015 2.705 52.19 6.19 ;
      LAYER met1 ;
        RECT 51.95 2.765 52.43 2.935 ;
        RECT 51.95 2.705 52.3 3.055 ;
        RECT 47.21 5.945 52.43 6.115 ;
        RECT 51.94 5.84 52.29 6.19 ;
        RECT 47.21 5.915 47.5 6.145 ;
      LAYER via1 ;
        RECT 52.04 5.94 52.19 6.09 ;
        RECT 52.05 2.805 52.2 2.955 ;
      LAYER mcon ;
        RECT 47.27 5.945 47.44 6.115 ;
        RECT 52.03 5.945 52.2 6.115 ;
        RECT 52.03 2.765 52.2 2.935 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 69.955 1.66 70.125 2.935 ;
        RECT 69.955 5.945 70.125 7.22 ;
        RECT 65.195 5.945 65.365 7.22 ;
      LAYER met2 ;
        RECT 69.875 2.705 70.225 3.055 ;
        RECT 69.865 5.84 70.215 6.19 ;
        RECT 69.94 2.705 70.115 6.19 ;
      LAYER met1 ;
        RECT 69.875 2.765 70.355 2.935 ;
        RECT 69.875 2.705 70.225 3.055 ;
        RECT 65.135 5.945 70.355 6.115 ;
        RECT 69.865 5.84 70.215 6.19 ;
        RECT 65.135 5.915 65.425 6.145 ;
      LAYER via1 ;
        RECT 69.965 5.94 70.115 6.09 ;
        RECT 69.975 2.805 70.125 2.955 ;
      LAYER mcon ;
        RECT 65.195 5.945 65.365 6.115 ;
        RECT 69.955 5.945 70.125 6.115 ;
        RECT 69.955 2.765 70.125 2.935 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 87.88 1.66 88.05 2.935 ;
        RECT 87.88 5.945 88.05 7.22 ;
        RECT 83.12 5.945 83.29 7.22 ;
      LAYER met2 ;
        RECT 87.8 2.705 88.15 3.055 ;
        RECT 87.79 5.84 88.14 6.19 ;
        RECT 87.865 2.705 88.04 6.19 ;
      LAYER met1 ;
        RECT 87.8 2.765 88.28 2.935 ;
        RECT 87.8 2.705 88.15 3.055 ;
        RECT 83.06 5.945 88.28 6.115 ;
        RECT 87.79 5.84 88.14 6.19 ;
        RECT 83.06 5.915 83.35 6.145 ;
      LAYER via1 ;
        RECT 87.89 5.94 88.04 6.09 ;
        RECT 87.9 2.805 88.05 2.955 ;
      LAYER mcon ;
        RECT 83.12 5.945 83.29 6.115 ;
        RECT 87.88 5.945 88.05 6.115 ;
        RECT 87.88 2.765 88.05 2.935 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 0.39 5.945 0.56 7.22 ;
      LAYER met1 ;
        RECT 0.33 5.945 0.79 6.115 ;
        RECT 0.33 5.915 0.62 6.145 ;
      LAYER mcon ;
        RECT 0.39 5.945 0.56 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0 4.285 92.575 4.745 ;
        RECT 86.615 4.135 92.575 4.745 ;
        RECT 90.44 4.13 92.42 4.75 ;
        RECT 91.6 3.4 91.77 5.48 ;
        RECT 90.61 3.4 90.78 5.48 ;
        RECT 87.87 3.405 88.04 5.475 ;
        RECT 85.115 3.785 85.285 4.745 ;
        RECT 83.11 4.285 83.28 5.475 ;
        RECT 82.675 3.785 82.845 4.745 ;
        RECT 80.715 3.785 80.885 4.745 ;
        RECT 79.755 3.785 79.925 4.745 ;
        RECT 77.795 3.785 77.965 4.745 ;
        RECT 76.795 3.785 76.965 4.745 ;
        RECT 75.835 3.785 76.005 4.745 ;
        RECT 68.69 4.135 74.65 4.745 ;
        RECT 72.515 4.13 74.495 4.75 ;
        RECT 73.675 3.4 73.845 5.48 ;
        RECT 72.685 3.4 72.855 5.48 ;
        RECT 69.945 3.405 70.115 5.475 ;
        RECT 67.19 3.785 67.36 4.745 ;
        RECT 65.185 4.285 65.355 5.475 ;
        RECT 64.75 3.785 64.92 4.745 ;
        RECT 62.79 3.785 62.96 4.745 ;
        RECT 61.83 3.785 62 4.745 ;
        RECT 59.87 3.785 60.04 4.745 ;
        RECT 58.87 3.785 59.04 4.745 ;
        RECT 57.91 3.785 58.08 4.745 ;
        RECT 50.765 4.135 56.725 4.745 ;
        RECT 54.59 4.13 56.57 4.75 ;
        RECT 55.75 3.4 55.92 5.48 ;
        RECT 54.76 3.4 54.93 5.48 ;
        RECT 52.02 3.405 52.19 5.475 ;
        RECT 49.265 3.785 49.435 4.745 ;
        RECT 47.26 4.285 47.43 5.475 ;
        RECT 46.825 3.785 46.995 4.745 ;
        RECT 44.865 3.785 45.035 4.745 ;
        RECT 43.905 3.785 44.075 4.745 ;
        RECT 41.945 3.785 42.115 4.745 ;
        RECT 40.945 3.785 41.115 4.745 ;
        RECT 39.985 3.785 40.155 4.745 ;
        RECT 32.84 4.135 38.8 4.745 ;
        RECT 36.665 4.13 38.645 4.75 ;
        RECT 37.825 3.4 37.995 5.48 ;
        RECT 36.835 3.4 37.005 5.48 ;
        RECT 34.095 3.405 34.265 5.475 ;
        RECT 31.34 3.785 31.51 4.745 ;
        RECT 29.335 4.285 29.505 5.475 ;
        RECT 28.9 3.785 29.07 4.745 ;
        RECT 26.94 3.785 27.11 4.745 ;
        RECT 25.98 3.785 26.15 4.745 ;
        RECT 24.02 3.785 24.19 4.745 ;
        RECT 23.02 3.785 23.19 4.745 ;
        RECT 22.06 3.785 22.23 4.745 ;
        RECT 14.915 4.135 20.875 4.745 ;
        RECT 18.74 4.13 20.72 4.75 ;
        RECT 19.9 3.4 20.07 5.48 ;
        RECT 18.91 3.4 19.08 5.48 ;
        RECT 16.17 3.405 16.34 5.475 ;
        RECT 13.415 3.785 13.585 4.745 ;
        RECT 11.41 4.285 11.58 5.475 ;
        RECT 10.975 3.785 11.145 4.745 ;
        RECT 9.015 3.785 9.185 4.745 ;
        RECT 8.055 3.785 8.225 4.745 ;
        RECT 6.095 3.785 6.265 4.745 ;
        RECT 5.095 3.785 5.265 4.745 ;
        RECT 4.135 3.785 4.305 4.745 ;
        RECT 2.19 4.285 2.36 8.305 ;
        RECT 0.38 4.285 0.55 5.475 ;
      LAYER met1 ;
        RECT 0 4.285 92.575 4.745 ;
        RECT 75.025 4.135 92.575 4.745 ;
        RECT 90.44 4.13 92.42 4.75 ;
        RECT 75.025 4.13 86.985 4.745 ;
        RECT 57.1 4.135 74.65 4.745 ;
        RECT 72.515 4.13 74.495 4.75 ;
        RECT 57.1 4.13 69.06 4.745 ;
        RECT 39.175 4.135 56.725 4.745 ;
        RECT 54.59 4.13 56.57 4.75 ;
        RECT 39.175 4.13 51.135 4.745 ;
        RECT 21.25 4.135 38.8 4.745 ;
        RECT 36.665 4.13 38.645 4.75 ;
        RECT 21.25 4.13 33.21 4.745 ;
        RECT 3.325 4.135 20.875 4.745 ;
        RECT 18.74 4.13 20.72 4.75 ;
        RECT 3.325 4.13 15.285 4.745 ;
        RECT 2.13 6.655 2.42 6.885 ;
        RECT 1.96 6.685 2.42 6.855 ;
      LAYER mcon ;
        RECT 2.19 6.685 2.36 6.855 ;
        RECT 2.5 4.545 2.67 4.715 ;
        RECT 3.47 4.285 3.64 4.455 ;
        RECT 3.93 4.285 4.1 4.455 ;
        RECT 4.39 4.285 4.56 4.455 ;
        RECT 4.85 4.285 5.02 4.455 ;
        RECT 5.31 4.285 5.48 4.455 ;
        RECT 5.77 4.285 5.94 4.455 ;
        RECT 6.23 4.285 6.4 4.455 ;
        RECT 6.69 4.285 6.86 4.455 ;
        RECT 7.15 4.285 7.32 4.455 ;
        RECT 7.61 4.285 7.78 4.455 ;
        RECT 8.07 4.285 8.24 4.455 ;
        RECT 8.53 4.285 8.7 4.455 ;
        RECT 8.99 4.285 9.16 4.455 ;
        RECT 9.45 4.285 9.62 4.455 ;
        RECT 9.91 4.285 10.08 4.455 ;
        RECT 10.37 4.285 10.54 4.455 ;
        RECT 10.83 4.285 11 4.455 ;
        RECT 11.29 4.285 11.46 4.455 ;
        RECT 11.75 4.285 11.92 4.455 ;
        RECT 12.21 4.285 12.38 4.455 ;
        RECT 12.67 4.285 12.84 4.455 ;
        RECT 13.13 4.285 13.3 4.455 ;
        RECT 13.53 4.545 13.7 4.715 ;
        RECT 13.59 4.285 13.76 4.455 ;
        RECT 14.05 4.285 14.22 4.455 ;
        RECT 14.51 4.285 14.68 4.455 ;
        RECT 14.97 4.285 15.14 4.455 ;
        RECT 18.29 4.545 18.46 4.715 ;
        RECT 18.29 4.165 18.46 4.335 ;
        RECT 18.99 4.55 19.16 4.72 ;
        RECT 18.99 4.16 19.16 4.33 ;
        RECT 19.98 4.55 20.15 4.72 ;
        RECT 19.98 4.16 20.15 4.33 ;
        RECT 21.395 4.285 21.565 4.455 ;
        RECT 21.855 4.285 22.025 4.455 ;
        RECT 22.315 4.285 22.485 4.455 ;
        RECT 22.775 4.285 22.945 4.455 ;
        RECT 23.235 4.285 23.405 4.455 ;
        RECT 23.695 4.285 23.865 4.455 ;
        RECT 24.155 4.285 24.325 4.455 ;
        RECT 24.615 4.285 24.785 4.455 ;
        RECT 25.075 4.285 25.245 4.455 ;
        RECT 25.535 4.285 25.705 4.455 ;
        RECT 25.995 4.285 26.165 4.455 ;
        RECT 26.455 4.285 26.625 4.455 ;
        RECT 26.915 4.285 27.085 4.455 ;
        RECT 27.375 4.285 27.545 4.455 ;
        RECT 27.835 4.285 28.005 4.455 ;
        RECT 28.295 4.285 28.465 4.455 ;
        RECT 28.755 4.285 28.925 4.455 ;
        RECT 29.215 4.285 29.385 4.455 ;
        RECT 29.675 4.285 29.845 4.455 ;
        RECT 30.135 4.285 30.305 4.455 ;
        RECT 30.595 4.285 30.765 4.455 ;
        RECT 31.055 4.285 31.225 4.455 ;
        RECT 31.455 4.545 31.625 4.715 ;
        RECT 31.515 4.285 31.685 4.455 ;
        RECT 31.975 4.285 32.145 4.455 ;
        RECT 32.435 4.285 32.605 4.455 ;
        RECT 32.895 4.285 33.065 4.455 ;
        RECT 36.215 4.545 36.385 4.715 ;
        RECT 36.215 4.165 36.385 4.335 ;
        RECT 36.915 4.55 37.085 4.72 ;
        RECT 36.915 4.16 37.085 4.33 ;
        RECT 37.905 4.55 38.075 4.72 ;
        RECT 37.905 4.16 38.075 4.33 ;
        RECT 39.32 4.285 39.49 4.455 ;
        RECT 39.78 4.285 39.95 4.455 ;
        RECT 40.24 4.285 40.41 4.455 ;
        RECT 40.7 4.285 40.87 4.455 ;
        RECT 41.16 4.285 41.33 4.455 ;
        RECT 41.62 4.285 41.79 4.455 ;
        RECT 42.08 4.285 42.25 4.455 ;
        RECT 42.54 4.285 42.71 4.455 ;
        RECT 43 4.285 43.17 4.455 ;
        RECT 43.46 4.285 43.63 4.455 ;
        RECT 43.92 4.285 44.09 4.455 ;
        RECT 44.38 4.285 44.55 4.455 ;
        RECT 44.84 4.285 45.01 4.455 ;
        RECT 45.3 4.285 45.47 4.455 ;
        RECT 45.76 4.285 45.93 4.455 ;
        RECT 46.22 4.285 46.39 4.455 ;
        RECT 46.68 4.285 46.85 4.455 ;
        RECT 47.14 4.285 47.31 4.455 ;
        RECT 47.6 4.285 47.77 4.455 ;
        RECT 48.06 4.285 48.23 4.455 ;
        RECT 48.52 4.285 48.69 4.455 ;
        RECT 48.98 4.285 49.15 4.455 ;
        RECT 49.38 4.545 49.55 4.715 ;
        RECT 49.44 4.285 49.61 4.455 ;
        RECT 49.9 4.285 50.07 4.455 ;
        RECT 50.36 4.285 50.53 4.455 ;
        RECT 50.82 4.285 50.99 4.455 ;
        RECT 54.14 4.545 54.31 4.715 ;
        RECT 54.14 4.165 54.31 4.335 ;
        RECT 54.84 4.55 55.01 4.72 ;
        RECT 54.84 4.16 55.01 4.33 ;
        RECT 55.83 4.55 56 4.72 ;
        RECT 55.83 4.16 56 4.33 ;
        RECT 57.245 4.285 57.415 4.455 ;
        RECT 57.705 4.285 57.875 4.455 ;
        RECT 58.165 4.285 58.335 4.455 ;
        RECT 58.625 4.285 58.795 4.455 ;
        RECT 59.085 4.285 59.255 4.455 ;
        RECT 59.545 4.285 59.715 4.455 ;
        RECT 60.005 4.285 60.175 4.455 ;
        RECT 60.465 4.285 60.635 4.455 ;
        RECT 60.925 4.285 61.095 4.455 ;
        RECT 61.385 4.285 61.555 4.455 ;
        RECT 61.845 4.285 62.015 4.455 ;
        RECT 62.305 4.285 62.475 4.455 ;
        RECT 62.765 4.285 62.935 4.455 ;
        RECT 63.225 4.285 63.395 4.455 ;
        RECT 63.685 4.285 63.855 4.455 ;
        RECT 64.145 4.285 64.315 4.455 ;
        RECT 64.605 4.285 64.775 4.455 ;
        RECT 65.065 4.285 65.235 4.455 ;
        RECT 65.525 4.285 65.695 4.455 ;
        RECT 65.985 4.285 66.155 4.455 ;
        RECT 66.445 4.285 66.615 4.455 ;
        RECT 66.905 4.285 67.075 4.455 ;
        RECT 67.305 4.545 67.475 4.715 ;
        RECT 67.365 4.285 67.535 4.455 ;
        RECT 67.825 4.285 67.995 4.455 ;
        RECT 68.285 4.285 68.455 4.455 ;
        RECT 68.745 4.285 68.915 4.455 ;
        RECT 72.065 4.545 72.235 4.715 ;
        RECT 72.065 4.165 72.235 4.335 ;
        RECT 72.765 4.55 72.935 4.72 ;
        RECT 72.765 4.16 72.935 4.33 ;
        RECT 73.755 4.55 73.925 4.72 ;
        RECT 73.755 4.16 73.925 4.33 ;
        RECT 75.17 4.285 75.34 4.455 ;
        RECT 75.63 4.285 75.8 4.455 ;
        RECT 76.09 4.285 76.26 4.455 ;
        RECT 76.55 4.285 76.72 4.455 ;
        RECT 77.01 4.285 77.18 4.455 ;
        RECT 77.47 4.285 77.64 4.455 ;
        RECT 77.93 4.285 78.1 4.455 ;
        RECT 78.39 4.285 78.56 4.455 ;
        RECT 78.85 4.285 79.02 4.455 ;
        RECT 79.31 4.285 79.48 4.455 ;
        RECT 79.77 4.285 79.94 4.455 ;
        RECT 80.23 4.285 80.4 4.455 ;
        RECT 80.69 4.285 80.86 4.455 ;
        RECT 81.15 4.285 81.32 4.455 ;
        RECT 81.61 4.285 81.78 4.455 ;
        RECT 82.07 4.285 82.24 4.455 ;
        RECT 82.53 4.285 82.7 4.455 ;
        RECT 82.99 4.285 83.16 4.455 ;
        RECT 83.45 4.285 83.62 4.455 ;
        RECT 83.91 4.285 84.08 4.455 ;
        RECT 84.37 4.285 84.54 4.455 ;
        RECT 84.83 4.285 85 4.455 ;
        RECT 85.23 4.545 85.4 4.715 ;
        RECT 85.29 4.285 85.46 4.455 ;
        RECT 85.75 4.285 85.92 4.455 ;
        RECT 86.21 4.285 86.38 4.455 ;
        RECT 86.67 4.285 86.84 4.455 ;
        RECT 89.99 4.545 90.16 4.715 ;
        RECT 89.99 4.165 90.16 4.335 ;
        RECT 90.69 4.55 90.86 4.72 ;
        RECT 90.69 4.16 90.86 4.33 ;
        RECT 91.68 4.55 91.85 4.72 ;
        RECT 91.68 4.16 91.85 4.33 ;
    END
  END vccd1
  OBS
    LAYER met3 ;
      RECT 84.38 7.055 84.755 7.425 ;
      RECT 84.415 4.925 84.725 7.425 ;
      RECT 84.415 4.925 87.51 5.235 ;
      RECT 87.2 1.125 87.51 5.235 ;
      RECT 87.2 1.14 87.575 1.51 ;
      RECT 84.33 3.685 84.885 4.015 ;
      RECT 84.33 2.02 84.63 4.015 ;
      RECT 80.395 3.125 80.95 3.455 ;
      RECT 80.65 2.02 80.95 3.455 ;
      RECT 81.445 1.885 81.595 2.535 ;
      RECT 80.65 2.02 84.63 2.32 ;
      RECT 79.165 0.96 79.465 3.91 ;
      RECT 79.155 2.565 79.885 2.895 ;
      RECT 79.12 0.96 79.495 1.33 ;
      RECT 77.715 3.125 78.445 3.455 ;
      RECT 77.73 0.96 78.03 3.455 ;
      RECT 75.605 2.565 76.335 2.895 ;
      RECT 75.76 0.93 76.06 2.895 ;
      RECT 77.685 0.96 78.06 1.33 ;
      RECT 75.715 0.93 76.09 1.3 ;
      RECT 75.715 0.97 78.06 1.27 ;
      RECT 66.455 7.055 66.83 7.425 ;
      RECT 66.49 4.925 66.8 7.425 ;
      RECT 66.49 4.925 69.585 5.235 ;
      RECT 69.275 1.125 69.585 5.235 ;
      RECT 69.275 1.14 69.65 1.51 ;
      RECT 66.405 3.685 66.96 4.015 ;
      RECT 66.405 2.02 66.705 4.015 ;
      RECT 62.47 3.125 63.025 3.455 ;
      RECT 62.725 2.02 63.025 3.455 ;
      RECT 63.52 1.885 63.67 2.535 ;
      RECT 62.725 2.02 66.705 2.32 ;
      RECT 61.24 0.96 61.54 3.91 ;
      RECT 61.23 2.565 61.96 2.895 ;
      RECT 61.195 0.96 61.57 1.33 ;
      RECT 59.79 3.125 60.52 3.455 ;
      RECT 59.805 0.96 60.105 3.455 ;
      RECT 57.68 2.565 58.41 2.895 ;
      RECT 57.835 0.93 58.135 2.895 ;
      RECT 59.76 0.96 60.135 1.33 ;
      RECT 57.79 0.93 58.165 1.3 ;
      RECT 57.79 0.97 60.135 1.27 ;
      RECT 48.53 7.055 48.905 7.425 ;
      RECT 48.565 4.925 48.875 7.425 ;
      RECT 48.565 4.925 51.66 5.235 ;
      RECT 51.35 1.125 51.66 5.235 ;
      RECT 51.35 1.14 51.725 1.51 ;
      RECT 48.48 3.685 49.035 4.015 ;
      RECT 48.48 2.02 48.78 4.015 ;
      RECT 44.545 3.125 45.1 3.455 ;
      RECT 44.8 2.02 45.1 3.455 ;
      RECT 45.595 1.885 45.745 2.535 ;
      RECT 44.8 2.02 48.78 2.32 ;
      RECT 43.315 0.96 43.615 3.91 ;
      RECT 43.305 2.565 44.035 2.895 ;
      RECT 43.27 0.96 43.645 1.33 ;
      RECT 41.865 3.125 42.595 3.455 ;
      RECT 41.88 0.96 42.18 3.455 ;
      RECT 39.755 2.565 40.485 2.895 ;
      RECT 39.91 0.93 40.21 2.895 ;
      RECT 41.835 0.96 42.21 1.33 ;
      RECT 39.865 0.93 40.24 1.3 ;
      RECT 39.865 0.97 42.21 1.27 ;
      RECT 30.605 7.055 30.98 7.425 ;
      RECT 30.64 4.925 30.95 7.425 ;
      RECT 30.64 4.925 33.735 5.235 ;
      RECT 33.425 1.125 33.735 5.235 ;
      RECT 33.425 1.14 33.8 1.51 ;
      RECT 30.555 3.685 31.11 4.015 ;
      RECT 30.555 2.02 30.855 4.015 ;
      RECT 26.62 3.125 27.175 3.455 ;
      RECT 26.875 2.02 27.175 3.455 ;
      RECT 27.67 1.885 27.82 2.535 ;
      RECT 26.875 2.02 30.855 2.32 ;
      RECT 25.39 0.96 25.69 3.91 ;
      RECT 25.38 2.565 26.11 2.895 ;
      RECT 25.345 0.96 25.72 1.33 ;
      RECT 23.94 3.125 24.67 3.455 ;
      RECT 23.955 0.96 24.255 3.455 ;
      RECT 21.83 2.565 22.56 2.895 ;
      RECT 21.985 0.93 22.285 2.895 ;
      RECT 23.91 0.96 24.285 1.33 ;
      RECT 21.94 0.93 22.315 1.3 ;
      RECT 21.94 0.97 24.285 1.27 ;
      RECT 12.68 7.055 13.055 7.425 ;
      RECT 12.715 4.925 13.025 7.425 ;
      RECT 12.715 4.925 15.81 5.235 ;
      RECT 15.5 1.125 15.81 5.235 ;
      RECT 15.5 1.14 15.875 1.51 ;
      RECT 12.63 3.685 13.185 4.015 ;
      RECT 12.63 2.02 12.93 4.015 ;
      RECT 8.695 3.125 9.25 3.455 ;
      RECT 8.95 2.02 9.25 3.455 ;
      RECT 9.745 1.885 9.895 2.535 ;
      RECT 8.95 2.02 12.93 2.32 ;
      RECT 7.465 0.96 7.765 3.91 ;
      RECT 7.455 2.565 8.185 2.895 ;
      RECT 7.42 0.96 7.795 1.33 ;
      RECT 6.015 3.125 6.745 3.455 ;
      RECT 6.03 0.96 6.33 3.455 ;
      RECT 3.905 2.565 4.635 2.895 ;
      RECT 4.06 0.93 4.36 2.895 ;
      RECT 5.985 0.96 6.36 1.33 ;
      RECT 4.015 0.93 4.39 1.3 ;
      RECT 4.015 0.97 6.36 1.27 ;
      RECT 85.515 2.005 86.245 2.335 ;
      RECT 83.295 3.685 84.025 4.015 ;
      RECT 81.595 3.685 82.325 4.015 ;
      RECT 76.64 2.565 77.37 2.895 ;
      RECT 75.275 3.685 76.005 4.015 ;
      RECT 67.59 2.005 68.32 2.335 ;
      RECT 65.37 3.685 66.1 4.015 ;
      RECT 63.67 3.685 64.4 4.015 ;
      RECT 58.715 2.565 59.445 2.895 ;
      RECT 57.35 3.685 58.08 4.015 ;
      RECT 49.665 2.005 50.395 2.335 ;
      RECT 47.445 3.685 48.175 4.015 ;
      RECT 45.745 3.685 46.475 4.015 ;
      RECT 40.79 2.565 41.52 2.895 ;
      RECT 39.425 3.685 40.155 4.015 ;
      RECT 31.74 2.005 32.47 2.335 ;
      RECT 29.52 3.685 30.25 4.015 ;
      RECT 27.82 3.685 28.55 4.015 ;
      RECT 22.865 2.565 23.595 2.895 ;
      RECT 21.5 3.685 22.23 4.015 ;
      RECT 13.815 2.005 14.545 2.335 ;
      RECT 11.595 3.685 12.325 4.015 ;
      RECT 9.895 3.685 10.625 4.015 ;
      RECT 4.94 2.565 5.67 2.895 ;
      RECT 3.575 3.685 4.305 4.015 ;
    LAYER via2 ;
      RECT 87.29 1.225 87.49 1.425 ;
      RECT 85.58 2.07 85.78 2.27 ;
      RECT 84.62 3.75 84.82 3.95 ;
      RECT 84.47 7.14 84.67 7.34 ;
      RECT 83.62 3.75 83.82 3.95 ;
      RECT 81.66 3.75 81.86 3.95 ;
      RECT 80.46 3.19 80.66 3.39 ;
      RECT 79.22 2.63 79.42 2.83 ;
      RECT 79.21 1.045 79.41 1.245 ;
      RECT 77.78 3.19 77.98 3.39 ;
      RECT 77.775 1.04 77.975 1.24 ;
      RECT 77.04 2.63 77.24 2.83 ;
      RECT 75.82 2.63 76.02 2.83 ;
      RECT 75.805 1.015 76.005 1.215 ;
      RECT 75.34 3.75 75.54 3.95 ;
      RECT 69.365 1.225 69.565 1.425 ;
      RECT 67.655 2.07 67.855 2.27 ;
      RECT 66.695 3.75 66.895 3.95 ;
      RECT 66.545 7.14 66.745 7.34 ;
      RECT 65.695 3.75 65.895 3.95 ;
      RECT 63.735 3.75 63.935 3.95 ;
      RECT 62.535 3.19 62.735 3.39 ;
      RECT 61.295 2.63 61.495 2.83 ;
      RECT 61.285 1.045 61.485 1.245 ;
      RECT 59.855 3.19 60.055 3.39 ;
      RECT 59.85 1.04 60.05 1.24 ;
      RECT 59.115 2.63 59.315 2.83 ;
      RECT 57.895 2.63 58.095 2.83 ;
      RECT 57.88 1.015 58.08 1.215 ;
      RECT 57.415 3.75 57.615 3.95 ;
      RECT 51.44 1.225 51.64 1.425 ;
      RECT 49.73 2.07 49.93 2.27 ;
      RECT 48.77 3.75 48.97 3.95 ;
      RECT 48.62 7.14 48.82 7.34 ;
      RECT 47.77 3.75 47.97 3.95 ;
      RECT 45.81 3.75 46.01 3.95 ;
      RECT 44.61 3.19 44.81 3.39 ;
      RECT 43.37 2.63 43.57 2.83 ;
      RECT 43.36 1.045 43.56 1.245 ;
      RECT 41.93 3.19 42.13 3.39 ;
      RECT 41.925 1.04 42.125 1.24 ;
      RECT 41.19 2.63 41.39 2.83 ;
      RECT 39.97 2.63 40.17 2.83 ;
      RECT 39.955 1.015 40.155 1.215 ;
      RECT 39.49 3.75 39.69 3.95 ;
      RECT 33.515 1.225 33.715 1.425 ;
      RECT 31.805 2.07 32.005 2.27 ;
      RECT 30.845 3.75 31.045 3.95 ;
      RECT 30.695 7.14 30.895 7.34 ;
      RECT 29.845 3.75 30.045 3.95 ;
      RECT 27.885 3.75 28.085 3.95 ;
      RECT 26.685 3.19 26.885 3.39 ;
      RECT 25.445 2.63 25.645 2.83 ;
      RECT 25.435 1.045 25.635 1.245 ;
      RECT 24.005 3.19 24.205 3.39 ;
      RECT 24 1.04 24.2 1.24 ;
      RECT 23.265 2.63 23.465 2.83 ;
      RECT 22.045 2.63 22.245 2.83 ;
      RECT 22.03 1.015 22.23 1.215 ;
      RECT 21.565 3.75 21.765 3.95 ;
      RECT 15.59 1.225 15.79 1.425 ;
      RECT 13.88 2.07 14.08 2.27 ;
      RECT 12.92 3.75 13.12 3.95 ;
      RECT 12.77 7.14 12.97 7.34 ;
      RECT 11.92 3.75 12.12 3.95 ;
      RECT 9.96 3.75 10.16 3.95 ;
      RECT 8.76 3.19 8.96 3.39 ;
      RECT 7.52 2.63 7.72 2.83 ;
      RECT 7.51 1.045 7.71 1.245 ;
      RECT 6.08 3.19 6.28 3.39 ;
      RECT 6.075 1.04 6.275 1.24 ;
      RECT 5.34 2.63 5.54 2.83 ;
      RECT 4.12 2.63 4.32 2.83 ;
      RECT 4.105 1.015 4.305 1.215 ;
      RECT 3.64 3.75 3.84 3.95 ;
    LAYER met2 ;
      RECT 1.385 8.4 92.2 8.57 ;
      RECT 92.03 7.275 92.2 8.57 ;
      RECT 1.385 6.255 1.555 8.57 ;
      RECT 92 7.275 92.35 7.625 ;
      RECT 1.325 6.255 1.615 6.605 ;
      RECT 88.845 6.225 89.165 6.545 ;
      RECT 88.875 5.695 89.045 6.545 ;
      RECT 88.875 5.695 89.05 6.045 ;
      RECT 88.875 5.695 89.85 5.87 ;
      RECT 89.675 1.965 89.85 5.87 ;
      RECT 89.62 1.965 89.97 2.315 ;
      RECT 89.645 6.655 89.97 6.98 ;
      RECT 88.53 6.745 89.97 6.915 ;
      RECT 88.53 2.395 88.69 6.915 ;
      RECT 88.845 2.365 89.165 2.685 ;
      RECT 88.53 2.395 89.165 2.565 ;
      RECT 87.2 1.14 87.575 1.51 ;
      RECT 79.12 0.96 79.495 1.33 ;
      RECT 77.685 0.96 78.06 1.33 ;
      RECT 77.685 1.08 87.505 1.25 ;
      RECT 81.805 4.36 87.485 4.53 ;
      RECT 87.315 3.425 87.485 4.53 ;
      RECT 81.615 3.6 81.64 4.53 ;
      RECT 81.87 3.71 81.9 3.99 ;
      RECT 81.575 3.6 81.64 3.86 ;
      RECT 87.225 3.43 87.575 3.78 ;
      RECT 81.405 2.225 81.44 2.485 ;
      RECT 81.18 2.225 81.24 2.485 ;
      RECT 81.86 3.69 81.87 3.99 ;
      RECT 81.855 3.65 81.86 3.99 ;
      RECT 81.84 3.605 81.855 3.99 ;
      RECT 81.835 3.57 81.84 3.99 ;
      RECT 81.83 3.55 81.835 3.99 ;
      RECT 81.805 3.487 81.83 3.99 ;
      RECT 81.8 3.425 81.805 4.53 ;
      RECT 81.78 3.375 81.8 4.53 ;
      RECT 81.77 3.305 81.78 4.53 ;
      RECT 81.725 3.245 81.77 4.53 ;
      RECT 81.64 3.206 81.725 4.53 ;
      RECT 81.635 3.197 81.64 3.57 ;
      RECT 81.625 3.196 81.635 3.553 ;
      RECT 81.6 3.177 81.625 3.523 ;
      RECT 81.595 3.152 81.6 3.502 ;
      RECT 81.585 3.13 81.595 3.493 ;
      RECT 81.58 3.101 81.585 3.483 ;
      RECT 81.54 3.027 81.58 3.455 ;
      RECT 81.52 2.928 81.54 3.42 ;
      RECT 81.505 2.864 81.52 3.403 ;
      RECT 81.475 2.788 81.505 3.375 ;
      RECT 81.455 2.703 81.475 3.348 ;
      RECT 81.415 2.599 81.455 3.255 ;
      RECT 81.41 2.52 81.415 3.163 ;
      RECT 81.405 2.503 81.41 3.14 ;
      RECT 81.4 2.225 81.405 3.12 ;
      RECT 81.37 2.225 81.4 3.058 ;
      RECT 81.365 2.225 81.37 2.99 ;
      RECT 81.355 2.225 81.365 2.955 ;
      RECT 81.345 2.225 81.355 2.92 ;
      RECT 81.28 2.225 81.345 2.775 ;
      RECT 81.275 2.225 81.28 2.645 ;
      RECT 81.245 2.225 81.275 2.578 ;
      RECT 81.24 2.225 81.245 2.503 ;
      RECT 85.575 2.16 85.835 2.42 ;
      RECT 85.57 2.16 85.835 2.368 ;
      RECT 85.565 2.16 85.835 2.338 ;
      RECT 85.54 2.03 85.82 2.31 ;
      RECT 74.055 6.655 74.405 7.005 ;
      RECT 85.3 6.61 85.65 6.96 ;
      RECT 74.055 6.685 85.65 6.885 ;
      RECT 84.58 3.71 84.86 3.99 ;
      RECT 84.62 3.665 84.885 3.925 ;
      RECT 84.61 3.7 84.885 3.925 ;
      RECT 84.615 3.685 84.86 3.99 ;
      RECT 84.62 3.662 84.83 3.99 ;
      RECT 84.62 3.66 84.815 3.99 ;
      RECT 84.66 3.65 84.815 3.99 ;
      RECT 84.63 3.655 84.815 3.99 ;
      RECT 84.66 3.647 84.76 3.99 ;
      RECT 84.685 3.64 84.76 3.99 ;
      RECT 84.665 3.642 84.76 3.99 ;
      RECT 83.995 3.155 84.255 3.415 ;
      RECT 84.045 3.147 84.235 3.415 ;
      RECT 84.05 3.067 84.235 3.415 ;
      RECT 84.17 2.455 84.235 3.415 ;
      RECT 84.075 2.852 84.235 3.415 ;
      RECT 84.15 2.54 84.235 3.415 ;
      RECT 84.185 2.165 84.321 2.893 ;
      RECT 84.13 2.662 84.321 2.893 ;
      RECT 84.145 2.602 84.235 3.415 ;
      RECT 84.185 2.165 84.345 2.558 ;
      RECT 84.185 2.165 84.355 2.455 ;
      RECT 84.175 2.165 84.435 2.425 ;
      RECT 83.58 3.71 83.86 3.99 ;
      RECT 83.6 3.67 83.86 3.99 ;
      RECT 83.24 3.625 83.345 3.885 ;
      RECT 83.095 2.115 83.185 2.375 ;
      RECT 83.635 3.18 83.64 3.22 ;
      RECT 83.63 3.17 83.635 3.305 ;
      RECT 83.625 3.16 83.63 3.398 ;
      RECT 83.615 3.14 83.625 3.454 ;
      RECT 83.535 3.068 83.615 3.534 ;
      RECT 83.57 3.712 83.58 3.937 ;
      RECT 83.565 3.709 83.57 3.932 ;
      RECT 83.55 3.706 83.565 3.925 ;
      RECT 83.515 3.7 83.55 3.907 ;
      RECT 83.53 3.003 83.535 3.608 ;
      RECT 83.51 2.954 83.53 3.623 ;
      RECT 83.5 3.687 83.515 3.89 ;
      RECT 83.505 2.896 83.51 3.638 ;
      RECT 83.5 2.874 83.505 3.648 ;
      RECT 83.465 2.784 83.5 3.885 ;
      RECT 83.45 2.662 83.465 3.885 ;
      RECT 83.445 2.615 83.45 3.885 ;
      RECT 83.42 2.54 83.445 3.885 ;
      RECT 83.405 2.455 83.42 3.885 ;
      RECT 83.4 2.402 83.405 3.885 ;
      RECT 83.395 2.382 83.4 3.885 ;
      RECT 83.39 2.357 83.395 3.119 ;
      RECT 83.375 3.317 83.395 3.885 ;
      RECT 83.385 2.335 83.39 3.096 ;
      RECT 83.375 2.287 83.385 3.061 ;
      RECT 83.37 2.25 83.375 3.027 ;
      RECT 83.37 3.397 83.375 3.885 ;
      RECT 83.355 2.227 83.37 2.982 ;
      RECT 83.35 3.495 83.37 3.885 ;
      RECT 83.3 2.115 83.355 2.824 ;
      RECT 83.345 3.617 83.35 3.885 ;
      RECT 83.285 2.115 83.3 2.663 ;
      RECT 83.28 2.115 83.285 2.615 ;
      RECT 83.275 2.115 83.28 2.603 ;
      RECT 83.23 2.115 83.275 2.54 ;
      RECT 83.205 2.115 83.23 2.458 ;
      RECT 83.19 2.115 83.205 2.41 ;
      RECT 83.185 2.115 83.19 2.38 ;
      RECT 82.51 3.565 82.555 3.825 ;
      RECT 82.415 2.1 82.56 2.36 ;
      RECT 82.92 2.722 82.93 2.813 ;
      RECT 82.905 2.66 82.92 2.869 ;
      RECT 82.9 2.607 82.905 2.915 ;
      RECT 82.85 2.554 82.9 3.041 ;
      RECT 82.845 2.509 82.85 3.188 ;
      RECT 82.835 2.497 82.845 3.23 ;
      RECT 82.8 2.461 82.835 3.335 ;
      RECT 82.795 2.429 82.8 3.441 ;
      RECT 82.78 2.411 82.795 3.486 ;
      RECT 82.775 2.394 82.78 2.72 ;
      RECT 82.77 2.775 82.78 3.543 ;
      RECT 82.765 2.38 82.775 2.693 ;
      RECT 82.76 2.83 82.77 3.825 ;
      RECT 82.755 2.366 82.765 2.678 ;
      RECT 82.755 2.88 82.76 3.825 ;
      RECT 82.74 2.343 82.755 2.658 ;
      RECT 82.72 3.002 82.755 3.825 ;
      RECT 82.735 2.325 82.74 2.64 ;
      RECT 82.73 2.317 82.735 2.63 ;
      RECT 82.7 2.285 82.73 2.594 ;
      RECT 82.71 3.13 82.72 3.825 ;
      RECT 82.705 3.157 82.71 3.825 ;
      RECT 82.7 3.207 82.705 3.825 ;
      RECT 82.69 2.251 82.7 2.559 ;
      RECT 82.65 3.275 82.7 3.825 ;
      RECT 82.675 2.228 82.69 2.535 ;
      RECT 82.65 2.1 82.675 2.498 ;
      RECT 82.645 2.1 82.65 2.47 ;
      RECT 82.615 3.375 82.65 3.825 ;
      RECT 82.64 2.1 82.645 2.463 ;
      RECT 82.635 2.1 82.64 2.453 ;
      RECT 82.62 2.1 82.635 2.438 ;
      RECT 82.605 2.1 82.62 2.41 ;
      RECT 82.57 3.48 82.615 3.825 ;
      RECT 82.59 2.1 82.605 2.383 ;
      RECT 82.56 2.1 82.59 2.368 ;
      RECT 82.555 3.552 82.57 3.825 ;
      RECT 82.48 2.635 82.52 2.895 ;
      RECT 82.255 2.582 82.26 2.84 ;
      RECT 78.21 2.06 78.47 2.32 ;
      RECT 78.21 2.085 78.485 2.3 ;
      RECT 80.6 1.91 80.605 2.055 ;
      RECT 82.47 2.63 82.48 2.895 ;
      RECT 82.45 2.622 82.47 2.895 ;
      RECT 82.432 2.618 82.45 2.895 ;
      RECT 82.346 2.607 82.432 2.895 ;
      RECT 82.26 2.59 82.346 2.895 ;
      RECT 82.205 2.577 82.255 2.825 ;
      RECT 82.171 2.569 82.205 2.8 ;
      RECT 82.085 2.558 82.171 2.765 ;
      RECT 82.05 2.535 82.085 2.73 ;
      RECT 82.04 2.497 82.05 2.716 ;
      RECT 82.035 2.47 82.04 2.712 ;
      RECT 82.03 2.457 82.035 2.709 ;
      RECT 82.02 2.437 82.03 2.705 ;
      RECT 82.015 2.412 82.02 2.701 ;
      RECT 81.99 2.367 82.015 2.695 ;
      RECT 81.98 2.308 81.99 2.687 ;
      RECT 81.97 2.276 81.98 2.678 ;
      RECT 81.95 2.228 81.97 2.658 ;
      RECT 81.945 2.188 81.95 2.628 ;
      RECT 81.93 2.162 81.945 2.602 ;
      RECT 81.925 2.14 81.93 2.578 ;
      RECT 81.91 2.112 81.925 2.554 ;
      RECT 81.895 2.085 81.91 2.518 ;
      RECT 81.88 2.062 81.895 2.48 ;
      RECT 81.875 2.052 81.88 2.455 ;
      RECT 81.865 2.045 81.875 2.438 ;
      RECT 81.85 2.032 81.865 2.408 ;
      RECT 81.845 2.022 81.85 2.383 ;
      RECT 81.84 2.017 81.845 2.37 ;
      RECT 81.83 2.01 81.84 2.35 ;
      RECT 81.825 2.003 81.83 2.335 ;
      RECT 81.8 1.996 81.825 2.293 ;
      RECT 81.785 1.986 81.8 2.243 ;
      RECT 81.775 1.981 81.785 2.213 ;
      RECT 81.765 1.977 81.775 2.188 ;
      RECT 81.75 1.974 81.765 2.178 ;
      RECT 81.7 1.971 81.75 2.163 ;
      RECT 81.68 1.969 81.7 2.148 ;
      RECT 81.631 1.967 81.68 2.143 ;
      RECT 81.545 1.963 81.631 2.138 ;
      RECT 81.506 1.96 81.545 2.134 ;
      RECT 81.42 1.956 81.506 2.129 ;
      RECT 81.37 1.953 81.42 2.123 ;
      RECT 81.321 1.95 81.37 2.118 ;
      RECT 81.235 1.947 81.321 2.113 ;
      RECT 81.231 1.945 81.235 2.11 ;
      RECT 81.145 1.942 81.231 2.105 ;
      RECT 81.096 1.938 81.145 2.098 ;
      RECT 81.01 1.935 81.096 2.093 ;
      RECT 80.986 1.932 81.01 2.089 ;
      RECT 80.9 1.93 80.986 2.084 ;
      RECT 80.835 1.926 80.9 2.077 ;
      RECT 80.832 1.925 80.835 2.074 ;
      RECT 80.746 1.922 80.832 2.071 ;
      RECT 80.66 1.916 80.746 2.064 ;
      RECT 80.63 1.912 80.66 2.06 ;
      RECT 80.605 1.91 80.63 2.058 ;
      RECT 80.55 1.907 80.6 2.055 ;
      RECT 80.47 1.906 80.55 2.055 ;
      RECT 80.415 1.908 80.47 2.058 ;
      RECT 80.4 1.909 80.415 2.062 ;
      RECT 80.345 1.917 80.4 2.072 ;
      RECT 80.315 1.925 80.345 2.085 ;
      RECT 80.296 1.926 80.315 2.091 ;
      RECT 80.21 1.929 80.296 2.096 ;
      RECT 80.14 1.934 80.21 2.105 ;
      RECT 80.121 1.937 80.14 2.111 ;
      RECT 80.035 1.941 80.121 2.116 ;
      RECT 79.995 1.945 80.035 2.123 ;
      RECT 79.986 1.947 79.995 2.126 ;
      RECT 79.9 1.951 79.986 2.131 ;
      RECT 79.897 1.954 79.9 2.135 ;
      RECT 79.811 1.957 79.897 2.139 ;
      RECT 79.725 1.963 79.811 2.147 ;
      RECT 79.701 1.967 79.725 2.151 ;
      RECT 79.615 1.971 79.701 2.156 ;
      RECT 79.57 1.976 79.615 2.163 ;
      RECT 79.49 1.981 79.57 2.17 ;
      RECT 79.41 1.987 79.49 2.185 ;
      RECT 79.385 1.991 79.41 2.198 ;
      RECT 79.32 1.994 79.385 2.21 ;
      RECT 79.265 1.999 79.32 2.225 ;
      RECT 79.235 2.002 79.265 2.243 ;
      RECT 79.225 2.004 79.235 2.256 ;
      RECT 79.165 2.019 79.225 2.266 ;
      RECT 79.15 2.036 79.165 2.275 ;
      RECT 79.145 2.045 79.15 2.275 ;
      RECT 79.135 2.055 79.145 2.275 ;
      RECT 79.125 2.072 79.135 2.275 ;
      RECT 79.105 2.082 79.125 2.276 ;
      RECT 79.06 2.092 79.105 2.277 ;
      RECT 79.025 2.101 79.06 2.279 ;
      RECT 78.96 2.106 79.025 2.281 ;
      RECT 78.88 2.107 78.96 2.284 ;
      RECT 78.876 2.105 78.88 2.285 ;
      RECT 78.79 2.102 78.876 2.287 ;
      RECT 78.743 2.099 78.79 2.289 ;
      RECT 78.657 2.095 78.743 2.292 ;
      RECT 78.571 2.091 78.657 2.295 ;
      RECT 78.485 2.087 78.571 2.299 ;
      RECT 80.42 3.15 80.7 3.43 ;
      RECT 80.46 3.13 80.72 3.39 ;
      RECT 80.45 3.14 80.72 3.39 ;
      RECT 80.46 3.067 80.675 3.43 ;
      RECT 80.515 2.99 80.67 3.43 ;
      RECT 80.52 2.775 80.67 3.43 ;
      RECT 80.51 2.577 80.66 2.828 ;
      RECT 80.5 2.577 80.66 2.695 ;
      RECT 80.495 2.455 80.655 2.598 ;
      RECT 80.48 2.455 80.655 2.503 ;
      RECT 80.475 2.165 80.65 2.48 ;
      RECT 80.46 2.165 80.65 2.45 ;
      RECT 80.42 2.165 80.68 2.425 ;
      RECT 80.33 3.635 80.41 3.895 ;
      RECT 79.735 2.355 79.74 2.62 ;
      RECT 79.615 2.355 79.74 2.615 ;
      RECT 80.29 3.6 80.33 3.895 ;
      RECT 80.245 3.522 80.29 3.895 ;
      RECT 80.225 3.45 80.245 3.895 ;
      RECT 80.215 3.402 80.225 3.895 ;
      RECT 80.18 3.335 80.215 3.895 ;
      RECT 80.15 3.235 80.18 3.895 ;
      RECT 80.13 3.16 80.15 3.695 ;
      RECT 80.12 3.11 80.13 3.65 ;
      RECT 80.115 3.087 80.12 3.623 ;
      RECT 80.11 3.072 80.115 3.61 ;
      RECT 80.105 3.057 80.11 3.588 ;
      RECT 80.1 3.042 80.105 3.57 ;
      RECT 80.075 2.997 80.1 3.525 ;
      RECT 80.065 2.945 80.075 3.468 ;
      RECT 80.055 2.915 80.065 3.435 ;
      RECT 80.045 2.88 80.055 3.403 ;
      RECT 80.01 2.812 80.045 3.335 ;
      RECT 80.005 2.751 80.01 3.27 ;
      RECT 79.995 2.739 80.005 3.25 ;
      RECT 79.99 2.727 79.995 3.23 ;
      RECT 79.985 2.719 79.99 3.218 ;
      RECT 79.98 2.711 79.985 3.198 ;
      RECT 79.97 2.699 79.98 3.17 ;
      RECT 79.96 2.683 79.97 3.14 ;
      RECT 79.935 2.655 79.96 3.078 ;
      RECT 79.925 2.626 79.935 3.023 ;
      RECT 79.91 2.605 79.925 2.983 ;
      RECT 79.905 2.589 79.91 2.955 ;
      RECT 79.9 2.577 79.905 2.945 ;
      RECT 79.895 2.572 79.9 2.918 ;
      RECT 79.89 2.565 79.895 2.905 ;
      RECT 79.875 2.548 79.89 2.878 ;
      RECT 79.865 2.355 79.875 2.838 ;
      RECT 79.855 2.355 79.865 2.805 ;
      RECT 79.845 2.355 79.855 2.78 ;
      RECT 79.775 2.355 79.845 2.715 ;
      RECT 79.765 2.355 79.775 2.663 ;
      RECT 79.75 2.355 79.765 2.645 ;
      RECT 79.74 2.355 79.75 2.63 ;
      RECT 79.57 3.225 79.83 3.485 ;
      RECT 78.105 3.26 78.11 3.467 ;
      RECT 77.74 3.15 77.815 3.465 ;
      RECT 77.555 3.205 77.71 3.465 ;
      RECT 77.74 3.15 77.845 3.43 ;
      RECT 79.555 3.322 79.57 3.483 ;
      RECT 79.53 3.33 79.555 3.488 ;
      RECT 79.505 3.337 79.53 3.493 ;
      RECT 79.442 3.348 79.505 3.502 ;
      RECT 79.356 3.367 79.442 3.519 ;
      RECT 79.27 3.389 79.356 3.538 ;
      RECT 79.255 3.402 79.27 3.549 ;
      RECT 79.215 3.41 79.255 3.556 ;
      RECT 79.195 3.415 79.215 3.563 ;
      RECT 79.157 3.416 79.195 3.566 ;
      RECT 79.071 3.419 79.157 3.567 ;
      RECT 78.985 3.423 79.071 3.568 ;
      RECT 78.936 3.425 78.985 3.57 ;
      RECT 78.85 3.425 78.936 3.572 ;
      RECT 78.81 3.42 78.85 3.574 ;
      RECT 78.8 3.414 78.81 3.575 ;
      RECT 78.76 3.409 78.8 3.572 ;
      RECT 78.75 3.402 78.76 3.568 ;
      RECT 78.735 3.398 78.75 3.566 ;
      RECT 78.718 3.394 78.735 3.564 ;
      RECT 78.632 3.384 78.718 3.556 ;
      RECT 78.546 3.366 78.632 3.542 ;
      RECT 78.46 3.349 78.546 3.528 ;
      RECT 78.435 3.337 78.46 3.519 ;
      RECT 78.365 3.327 78.435 3.512 ;
      RECT 78.32 3.315 78.365 3.503 ;
      RECT 78.26 3.302 78.32 3.495 ;
      RECT 78.255 3.294 78.26 3.49 ;
      RECT 78.22 3.289 78.255 3.488 ;
      RECT 78.165 3.28 78.22 3.481 ;
      RECT 78.125 3.269 78.165 3.473 ;
      RECT 78.11 3.262 78.125 3.469 ;
      RECT 78.09 3.255 78.105 3.466 ;
      RECT 78.075 3.245 78.09 3.464 ;
      RECT 78.06 3.232 78.075 3.461 ;
      RECT 78.035 3.215 78.06 3.457 ;
      RECT 78.02 3.197 78.035 3.454 ;
      RECT 77.995 3.15 78.02 3.452 ;
      RECT 77.971 3.15 77.995 3.449 ;
      RECT 77.885 3.15 77.971 3.441 ;
      RECT 77.845 3.15 77.885 3.433 ;
      RECT 77.71 3.197 77.74 3.465 ;
      RECT 79.39 2.78 79.65 3.04 ;
      RECT 79.35 2.78 79.65 2.918 ;
      RECT 79.315 2.78 79.65 2.903 ;
      RECT 79.26 2.78 79.65 2.883 ;
      RECT 79.18 2.59 79.46 2.87 ;
      RECT 79.18 2.772 79.53 2.87 ;
      RECT 79.18 2.715 79.515 2.87 ;
      RECT 79.18 2.662 79.465 2.87 ;
      RECT 77.01 2.59 77.205 3.375 ;
      RECT 77.09 1.205 77.205 3.375 ;
      RECT 76.945 3.115 77.005 3.375 ;
      RECT 78.315 2.635 78.575 2.895 ;
      RECT 77 2.59 77.205 2.87 ;
      RECT 78.31 2.645 78.575 2.83 ;
      RECT 78.025 2.62 78.035 2.77 ;
      RECT 77.26 1.205 77.34 1.55 ;
      RECT 76.995 1.205 77.205 1.55 ;
      RECT 78.3 2.645 78.31 2.829 ;
      RECT 78.29 2.644 78.3 2.826 ;
      RECT 78.281 2.643 78.29 2.824 ;
      RECT 78.195 2.639 78.281 2.814 ;
      RECT 78.121 2.631 78.195 2.796 ;
      RECT 78.035 2.624 78.121 2.779 ;
      RECT 77.975 2.62 78.025 2.769 ;
      RECT 77.94 2.619 77.975 2.766 ;
      RECT 77.885 2.619 77.94 2.768 ;
      RECT 77.85 2.619 77.885 2.772 ;
      RECT 77.764 2.618 77.85 2.779 ;
      RECT 77.678 2.617 77.764 2.789 ;
      RECT 77.592 2.616 77.678 2.8 ;
      RECT 77.506 2.616 77.592 2.81 ;
      RECT 77.42 2.615 77.506 2.82 ;
      RECT 77.385 2.615 77.42 2.86 ;
      RECT 77.38 2.615 77.385 2.903 ;
      RECT 77.355 2.615 77.38 2.92 ;
      RECT 77.28 2.615 77.355 2.935 ;
      RECT 77.26 2.59 77.28 2.948 ;
      RECT 77.255 1.205 77.26 2.958 ;
      RECT 77.23 1.205 77.255 3 ;
      RECT 77.205 1.205 77.23 3.078 ;
      RECT 77.005 2.997 77.01 3.375 ;
      RECT 76.34 2.949 76.355 3.405 ;
      RECT 76.335 3.021 76.441 3.403 ;
      RECT 76.355 2.115 76.49 3.401 ;
      RECT 76.34 2.965 76.495 3.4 ;
      RECT 76.34 3.015 76.5 3.398 ;
      RECT 76.325 3.08 76.5 3.397 ;
      RECT 76.335 3.072 76.505 3.394 ;
      RECT 76.315 3.12 76.505 3.389 ;
      RECT 76.315 3.12 76.52 3.386 ;
      RECT 76.31 3.12 76.52 3.383 ;
      RECT 76.285 3.12 76.545 3.38 ;
      RECT 76.355 2.115 76.515 2.768 ;
      RECT 76.35 2.115 76.515 2.74 ;
      RECT 76.345 2.115 76.515 2.568 ;
      RECT 76.345 2.115 76.535 2.508 ;
      RECT 76.3 2.115 76.56 2.375 ;
      RECT 75.78 2.59 76.06 2.87 ;
      RECT 75.77 2.605 76.06 2.865 ;
      RECT 75.725 2.667 76.06 2.863 ;
      RECT 75.8 2.582 75.965 2.87 ;
      RECT 75.8 2.567 75.921 2.87 ;
      RECT 75.835 2.56 75.921 2.87 ;
      RECT 75.3 3.71 75.58 3.99 ;
      RECT 75.26 3.672 75.555 3.783 ;
      RECT 75.245 3.622 75.535 3.678 ;
      RECT 75.19 3.385 75.45 3.645 ;
      RECT 75.19 3.587 75.53 3.645 ;
      RECT 75.19 3.527 75.525 3.645 ;
      RECT 75.19 3.477 75.505 3.645 ;
      RECT 75.19 3.457 75.5 3.645 ;
      RECT 75.19 3.435 75.495 3.645 ;
      RECT 75.19 3.42 75.465 3.645 ;
      RECT 70.92 6.225 71.24 6.545 ;
      RECT 70.95 5.695 71.12 6.545 ;
      RECT 70.95 5.695 71.125 6.045 ;
      RECT 70.95 5.695 71.925 5.87 ;
      RECT 71.75 1.965 71.925 5.87 ;
      RECT 71.695 1.965 72.045 2.315 ;
      RECT 71.72 6.655 72.045 6.98 ;
      RECT 70.605 6.745 72.045 6.915 ;
      RECT 70.605 2.395 70.765 6.915 ;
      RECT 70.92 2.365 71.24 2.685 ;
      RECT 70.605 2.395 71.24 2.565 ;
      RECT 69.275 1.14 69.65 1.51 ;
      RECT 61.195 0.96 61.57 1.33 ;
      RECT 59.76 0.96 60.135 1.33 ;
      RECT 59.76 1.08 69.58 1.25 ;
      RECT 63.88 4.36 69.56 4.53 ;
      RECT 69.39 3.425 69.56 4.53 ;
      RECT 63.69 3.6 63.715 4.53 ;
      RECT 63.945 3.71 63.975 3.99 ;
      RECT 63.65 3.6 63.715 3.86 ;
      RECT 69.3 3.43 69.65 3.78 ;
      RECT 63.48 2.225 63.515 2.485 ;
      RECT 63.255 2.225 63.315 2.485 ;
      RECT 63.935 3.69 63.945 3.99 ;
      RECT 63.93 3.65 63.935 3.99 ;
      RECT 63.915 3.605 63.93 3.99 ;
      RECT 63.91 3.57 63.915 3.99 ;
      RECT 63.905 3.55 63.91 3.99 ;
      RECT 63.88 3.487 63.905 3.99 ;
      RECT 63.875 3.425 63.88 4.53 ;
      RECT 63.855 3.375 63.875 4.53 ;
      RECT 63.845 3.305 63.855 4.53 ;
      RECT 63.8 3.245 63.845 4.53 ;
      RECT 63.715 3.206 63.8 4.53 ;
      RECT 63.71 3.197 63.715 3.57 ;
      RECT 63.7 3.196 63.71 3.553 ;
      RECT 63.675 3.177 63.7 3.523 ;
      RECT 63.67 3.152 63.675 3.502 ;
      RECT 63.66 3.13 63.67 3.493 ;
      RECT 63.655 3.101 63.66 3.483 ;
      RECT 63.615 3.027 63.655 3.455 ;
      RECT 63.595 2.928 63.615 3.42 ;
      RECT 63.58 2.864 63.595 3.403 ;
      RECT 63.55 2.788 63.58 3.375 ;
      RECT 63.53 2.703 63.55 3.348 ;
      RECT 63.49 2.599 63.53 3.255 ;
      RECT 63.485 2.52 63.49 3.163 ;
      RECT 63.48 2.503 63.485 3.14 ;
      RECT 63.475 2.225 63.48 3.12 ;
      RECT 63.445 2.225 63.475 3.058 ;
      RECT 63.44 2.225 63.445 2.99 ;
      RECT 63.43 2.225 63.44 2.955 ;
      RECT 63.42 2.225 63.43 2.92 ;
      RECT 63.355 2.225 63.42 2.775 ;
      RECT 63.35 2.225 63.355 2.645 ;
      RECT 63.32 2.225 63.35 2.578 ;
      RECT 63.315 2.225 63.32 2.503 ;
      RECT 67.65 2.16 67.91 2.42 ;
      RECT 67.645 2.16 67.91 2.368 ;
      RECT 67.64 2.16 67.91 2.338 ;
      RECT 67.615 2.03 67.895 2.31 ;
      RECT 56.13 6.655 56.48 7.005 ;
      RECT 67.095 6.61 67.445 6.96 ;
      RECT 56.13 6.685 67.445 6.885 ;
      RECT 66.655 3.71 66.935 3.99 ;
      RECT 66.695 3.665 66.96 3.925 ;
      RECT 66.685 3.7 66.96 3.925 ;
      RECT 66.69 3.685 66.935 3.99 ;
      RECT 66.695 3.662 66.905 3.99 ;
      RECT 66.695 3.66 66.89 3.99 ;
      RECT 66.735 3.65 66.89 3.99 ;
      RECT 66.705 3.655 66.89 3.99 ;
      RECT 66.735 3.647 66.835 3.99 ;
      RECT 66.76 3.64 66.835 3.99 ;
      RECT 66.74 3.642 66.835 3.99 ;
      RECT 66.07 3.155 66.33 3.415 ;
      RECT 66.12 3.147 66.31 3.415 ;
      RECT 66.125 3.067 66.31 3.415 ;
      RECT 66.245 2.455 66.31 3.415 ;
      RECT 66.15 2.852 66.31 3.415 ;
      RECT 66.225 2.54 66.31 3.415 ;
      RECT 66.26 2.165 66.396 2.893 ;
      RECT 66.205 2.662 66.396 2.893 ;
      RECT 66.22 2.602 66.31 3.415 ;
      RECT 66.26 2.165 66.42 2.558 ;
      RECT 66.26 2.165 66.43 2.455 ;
      RECT 66.25 2.165 66.51 2.425 ;
      RECT 65.655 3.71 65.935 3.99 ;
      RECT 65.675 3.67 65.935 3.99 ;
      RECT 65.315 3.625 65.42 3.885 ;
      RECT 65.17 2.115 65.26 2.375 ;
      RECT 65.71 3.18 65.715 3.22 ;
      RECT 65.705 3.17 65.71 3.305 ;
      RECT 65.7 3.16 65.705 3.398 ;
      RECT 65.69 3.14 65.7 3.454 ;
      RECT 65.61 3.068 65.69 3.534 ;
      RECT 65.645 3.712 65.655 3.937 ;
      RECT 65.64 3.709 65.645 3.932 ;
      RECT 65.625 3.706 65.64 3.925 ;
      RECT 65.59 3.7 65.625 3.907 ;
      RECT 65.605 3.003 65.61 3.608 ;
      RECT 65.585 2.954 65.605 3.623 ;
      RECT 65.575 3.687 65.59 3.89 ;
      RECT 65.58 2.896 65.585 3.638 ;
      RECT 65.575 2.874 65.58 3.648 ;
      RECT 65.54 2.784 65.575 3.885 ;
      RECT 65.525 2.662 65.54 3.885 ;
      RECT 65.52 2.615 65.525 3.885 ;
      RECT 65.495 2.54 65.52 3.885 ;
      RECT 65.48 2.455 65.495 3.885 ;
      RECT 65.475 2.402 65.48 3.885 ;
      RECT 65.47 2.382 65.475 3.885 ;
      RECT 65.465 2.357 65.47 3.119 ;
      RECT 65.45 3.317 65.47 3.885 ;
      RECT 65.46 2.335 65.465 3.096 ;
      RECT 65.45 2.287 65.46 3.061 ;
      RECT 65.445 2.25 65.45 3.027 ;
      RECT 65.445 3.397 65.45 3.885 ;
      RECT 65.43 2.227 65.445 2.982 ;
      RECT 65.425 3.495 65.445 3.885 ;
      RECT 65.375 2.115 65.43 2.824 ;
      RECT 65.42 3.617 65.425 3.885 ;
      RECT 65.36 2.115 65.375 2.663 ;
      RECT 65.355 2.115 65.36 2.615 ;
      RECT 65.35 2.115 65.355 2.603 ;
      RECT 65.305 2.115 65.35 2.54 ;
      RECT 65.28 2.115 65.305 2.458 ;
      RECT 65.265 2.115 65.28 2.41 ;
      RECT 65.26 2.115 65.265 2.38 ;
      RECT 64.585 3.565 64.63 3.825 ;
      RECT 64.49 2.1 64.635 2.36 ;
      RECT 64.995 2.722 65.005 2.813 ;
      RECT 64.98 2.66 64.995 2.869 ;
      RECT 64.975 2.607 64.98 2.915 ;
      RECT 64.925 2.554 64.975 3.041 ;
      RECT 64.92 2.509 64.925 3.188 ;
      RECT 64.91 2.497 64.92 3.23 ;
      RECT 64.875 2.461 64.91 3.335 ;
      RECT 64.87 2.429 64.875 3.441 ;
      RECT 64.855 2.411 64.87 3.486 ;
      RECT 64.85 2.394 64.855 2.72 ;
      RECT 64.845 2.775 64.855 3.543 ;
      RECT 64.84 2.38 64.85 2.693 ;
      RECT 64.835 2.83 64.845 3.825 ;
      RECT 64.83 2.366 64.84 2.678 ;
      RECT 64.83 2.88 64.835 3.825 ;
      RECT 64.815 2.343 64.83 2.658 ;
      RECT 64.795 3.002 64.83 3.825 ;
      RECT 64.81 2.325 64.815 2.64 ;
      RECT 64.805 2.317 64.81 2.63 ;
      RECT 64.775 2.285 64.805 2.594 ;
      RECT 64.785 3.13 64.795 3.825 ;
      RECT 64.78 3.157 64.785 3.825 ;
      RECT 64.775 3.207 64.78 3.825 ;
      RECT 64.765 2.251 64.775 2.559 ;
      RECT 64.725 3.275 64.775 3.825 ;
      RECT 64.75 2.228 64.765 2.535 ;
      RECT 64.725 2.1 64.75 2.498 ;
      RECT 64.72 2.1 64.725 2.47 ;
      RECT 64.69 3.375 64.725 3.825 ;
      RECT 64.715 2.1 64.72 2.463 ;
      RECT 64.71 2.1 64.715 2.453 ;
      RECT 64.695 2.1 64.71 2.438 ;
      RECT 64.68 2.1 64.695 2.41 ;
      RECT 64.645 3.48 64.69 3.825 ;
      RECT 64.665 2.1 64.68 2.383 ;
      RECT 64.635 2.1 64.665 2.368 ;
      RECT 64.63 3.552 64.645 3.825 ;
      RECT 64.555 2.635 64.595 2.895 ;
      RECT 64.33 2.582 64.335 2.84 ;
      RECT 60.285 2.06 60.545 2.32 ;
      RECT 60.285 2.085 60.56 2.3 ;
      RECT 62.675 1.91 62.68 2.055 ;
      RECT 64.545 2.63 64.555 2.895 ;
      RECT 64.525 2.622 64.545 2.895 ;
      RECT 64.507 2.618 64.525 2.895 ;
      RECT 64.421 2.607 64.507 2.895 ;
      RECT 64.335 2.59 64.421 2.895 ;
      RECT 64.28 2.577 64.33 2.825 ;
      RECT 64.246 2.569 64.28 2.8 ;
      RECT 64.16 2.558 64.246 2.765 ;
      RECT 64.125 2.535 64.16 2.73 ;
      RECT 64.115 2.497 64.125 2.716 ;
      RECT 64.11 2.47 64.115 2.712 ;
      RECT 64.105 2.457 64.11 2.709 ;
      RECT 64.095 2.437 64.105 2.705 ;
      RECT 64.09 2.412 64.095 2.701 ;
      RECT 64.065 2.367 64.09 2.695 ;
      RECT 64.055 2.308 64.065 2.687 ;
      RECT 64.045 2.276 64.055 2.678 ;
      RECT 64.025 2.228 64.045 2.658 ;
      RECT 64.02 2.188 64.025 2.628 ;
      RECT 64.005 2.162 64.02 2.602 ;
      RECT 64 2.14 64.005 2.578 ;
      RECT 63.985 2.112 64 2.554 ;
      RECT 63.97 2.085 63.985 2.518 ;
      RECT 63.955 2.062 63.97 2.48 ;
      RECT 63.95 2.052 63.955 2.455 ;
      RECT 63.94 2.045 63.95 2.438 ;
      RECT 63.925 2.032 63.94 2.408 ;
      RECT 63.92 2.022 63.925 2.383 ;
      RECT 63.915 2.017 63.92 2.37 ;
      RECT 63.905 2.01 63.915 2.35 ;
      RECT 63.9 2.003 63.905 2.335 ;
      RECT 63.875 1.996 63.9 2.293 ;
      RECT 63.86 1.986 63.875 2.243 ;
      RECT 63.85 1.981 63.86 2.213 ;
      RECT 63.84 1.977 63.85 2.188 ;
      RECT 63.825 1.974 63.84 2.178 ;
      RECT 63.775 1.971 63.825 2.163 ;
      RECT 63.755 1.969 63.775 2.148 ;
      RECT 63.706 1.967 63.755 2.143 ;
      RECT 63.62 1.963 63.706 2.138 ;
      RECT 63.581 1.96 63.62 2.134 ;
      RECT 63.495 1.956 63.581 2.129 ;
      RECT 63.445 1.953 63.495 2.123 ;
      RECT 63.396 1.95 63.445 2.118 ;
      RECT 63.31 1.947 63.396 2.113 ;
      RECT 63.306 1.945 63.31 2.11 ;
      RECT 63.22 1.942 63.306 2.105 ;
      RECT 63.171 1.938 63.22 2.098 ;
      RECT 63.085 1.935 63.171 2.093 ;
      RECT 63.061 1.932 63.085 2.089 ;
      RECT 62.975 1.93 63.061 2.084 ;
      RECT 62.91 1.926 62.975 2.077 ;
      RECT 62.907 1.925 62.91 2.074 ;
      RECT 62.821 1.922 62.907 2.071 ;
      RECT 62.735 1.916 62.821 2.064 ;
      RECT 62.705 1.912 62.735 2.06 ;
      RECT 62.68 1.91 62.705 2.058 ;
      RECT 62.625 1.907 62.675 2.055 ;
      RECT 62.545 1.906 62.625 2.055 ;
      RECT 62.49 1.908 62.545 2.058 ;
      RECT 62.475 1.909 62.49 2.062 ;
      RECT 62.42 1.917 62.475 2.072 ;
      RECT 62.39 1.925 62.42 2.085 ;
      RECT 62.371 1.926 62.39 2.091 ;
      RECT 62.285 1.929 62.371 2.096 ;
      RECT 62.215 1.934 62.285 2.105 ;
      RECT 62.196 1.937 62.215 2.111 ;
      RECT 62.11 1.941 62.196 2.116 ;
      RECT 62.07 1.945 62.11 2.123 ;
      RECT 62.061 1.947 62.07 2.126 ;
      RECT 61.975 1.951 62.061 2.131 ;
      RECT 61.972 1.954 61.975 2.135 ;
      RECT 61.886 1.957 61.972 2.139 ;
      RECT 61.8 1.963 61.886 2.147 ;
      RECT 61.776 1.967 61.8 2.151 ;
      RECT 61.69 1.971 61.776 2.156 ;
      RECT 61.645 1.976 61.69 2.163 ;
      RECT 61.565 1.981 61.645 2.17 ;
      RECT 61.485 1.987 61.565 2.185 ;
      RECT 61.46 1.991 61.485 2.198 ;
      RECT 61.395 1.994 61.46 2.21 ;
      RECT 61.34 1.999 61.395 2.225 ;
      RECT 61.31 2.002 61.34 2.243 ;
      RECT 61.3 2.004 61.31 2.256 ;
      RECT 61.24 2.019 61.3 2.266 ;
      RECT 61.225 2.036 61.24 2.275 ;
      RECT 61.22 2.045 61.225 2.275 ;
      RECT 61.21 2.055 61.22 2.275 ;
      RECT 61.2 2.072 61.21 2.275 ;
      RECT 61.18 2.082 61.2 2.276 ;
      RECT 61.135 2.092 61.18 2.277 ;
      RECT 61.1 2.101 61.135 2.279 ;
      RECT 61.035 2.106 61.1 2.281 ;
      RECT 60.955 2.107 61.035 2.284 ;
      RECT 60.951 2.105 60.955 2.285 ;
      RECT 60.865 2.102 60.951 2.287 ;
      RECT 60.818 2.099 60.865 2.289 ;
      RECT 60.732 2.095 60.818 2.292 ;
      RECT 60.646 2.091 60.732 2.295 ;
      RECT 60.56 2.087 60.646 2.299 ;
      RECT 62.495 3.15 62.775 3.43 ;
      RECT 62.535 3.13 62.795 3.39 ;
      RECT 62.525 3.14 62.795 3.39 ;
      RECT 62.535 3.067 62.75 3.43 ;
      RECT 62.59 2.99 62.745 3.43 ;
      RECT 62.595 2.775 62.745 3.43 ;
      RECT 62.585 2.577 62.735 2.828 ;
      RECT 62.575 2.577 62.735 2.695 ;
      RECT 62.57 2.455 62.73 2.598 ;
      RECT 62.555 2.455 62.73 2.503 ;
      RECT 62.55 2.165 62.725 2.48 ;
      RECT 62.535 2.165 62.725 2.45 ;
      RECT 62.495 2.165 62.755 2.425 ;
      RECT 62.405 3.635 62.485 3.895 ;
      RECT 61.81 2.355 61.815 2.62 ;
      RECT 61.69 2.355 61.815 2.615 ;
      RECT 62.365 3.6 62.405 3.895 ;
      RECT 62.32 3.522 62.365 3.895 ;
      RECT 62.3 3.45 62.32 3.895 ;
      RECT 62.29 3.402 62.3 3.895 ;
      RECT 62.255 3.335 62.29 3.895 ;
      RECT 62.225 3.235 62.255 3.895 ;
      RECT 62.205 3.16 62.225 3.695 ;
      RECT 62.195 3.11 62.205 3.65 ;
      RECT 62.19 3.087 62.195 3.623 ;
      RECT 62.185 3.072 62.19 3.61 ;
      RECT 62.18 3.057 62.185 3.588 ;
      RECT 62.175 3.042 62.18 3.57 ;
      RECT 62.15 2.997 62.175 3.525 ;
      RECT 62.14 2.945 62.15 3.468 ;
      RECT 62.13 2.915 62.14 3.435 ;
      RECT 62.12 2.88 62.13 3.403 ;
      RECT 62.085 2.812 62.12 3.335 ;
      RECT 62.08 2.751 62.085 3.27 ;
      RECT 62.07 2.739 62.08 3.25 ;
      RECT 62.065 2.727 62.07 3.23 ;
      RECT 62.06 2.719 62.065 3.218 ;
      RECT 62.055 2.711 62.06 3.198 ;
      RECT 62.045 2.699 62.055 3.17 ;
      RECT 62.035 2.683 62.045 3.14 ;
      RECT 62.01 2.655 62.035 3.078 ;
      RECT 62 2.626 62.01 3.023 ;
      RECT 61.985 2.605 62 2.983 ;
      RECT 61.98 2.589 61.985 2.955 ;
      RECT 61.975 2.577 61.98 2.945 ;
      RECT 61.97 2.572 61.975 2.918 ;
      RECT 61.965 2.565 61.97 2.905 ;
      RECT 61.95 2.548 61.965 2.878 ;
      RECT 61.94 2.355 61.95 2.838 ;
      RECT 61.93 2.355 61.94 2.805 ;
      RECT 61.92 2.355 61.93 2.78 ;
      RECT 61.85 2.355 61.92 2.715 ;
      RECT 61.84 2.355 61.85 2.663 ;
      RECT 61.825 2.355 61.84 2.645 ;
      RECT 61.815 2.355 61.825 2.63 ;
      RECT 61.645 3.225 61.905 3.485 ;
      RECT 60.18 3.26 60.185 3.467 ;
      RECT 59.815 3.15 59.89 3.465 ;
      RECT 59.63 3.205 59.785 3.465 ;
      RECT 59.815 3.15 59.92 3.43 ;
      RECT 61.63 3.322 61.645 3.483 ;
      RECT 61.605 3.33 61.63 3.488 ;
      RECT 61.58 3.337 61.605 3.493 ;
      RECT 61.517 3.348 61.58 3.502 ;
      RECT 61.431 3.367 61.517 3.519 ;
      RECT 61.345 3.389 61.431 3.538 ;
      RECT 61.33 3.402 61.345 3.549 ;
      RECT 61.29 3.41 61.33 3.556 ;
      RECT 61.27 3.415 61.29 3.563 ;
      RECT 61.232 3.416 61.27 3.566 ;
      RECT 61.146 3.419 61.232 3.567 ;
      RECT 61.06 3.423 61.146 3.568 ;
      RECT 61.011 3.425 61.06 3.57 ;
      RECT 60.925 3.425 61.011 3.572 ;
      RECT 60.885 3.42 60.925 3.574 ;
      RECT 60.875 3.414 60.885 3.575 ;
      RECT 60.835 3.409 60.875 3.572 ;
      RECT 60.825 3.402 60.835 3.568 ;
      RECT 60.81 3.398 60.825 3.566 ;
      RECT 60.793 3.394 60.81 3.564 ;
      RECT 60.707 3.384 60.793 3.556 ;
      RECT 60.621 3.366 60.707 3.542 ;
      RECT 60.535 3.349 60.621 3.528 ;
      RECT 60.51 3.337 60.535 3.519 ;
      RECT 60.44 3.327 60.51 3.512 ;
      RECT 60.395 3.315 60.44 3.503 ;
      RECT 60.335 3.302 60.395 3.495 ;
      RECT 60.33 3.294 60.335 3.49 ;
      RECT 60.295 3.289 60.33 3.488 ;
      RECT 60.24 3.28 60.295 3.481 ;
      RECT 60.2 3.269 60.24 3.473 ;
      RECT 60.185 3.262 60.2 3.469 ;
      RECT 60.165 3.255 60.18 3.466 ;
      RECT 60.15 3.245 60.165 3.464 ;
      RECT 60.135 3.232 60.15 3.461 ;
      RECT 60.11 3.215 60.135 3.457 ;
      RECT 60.095 3.197 60.11 3.454 ;
      RECT 60.07 3.15 60.095 3.452 ;
      RECT 60.046 3.15 60.07 3.449 ;
      RECT 59.96 3.15 60.046 3.441 ;
      RECT 59.92 3.15 59.96 3.433 ;
      RECT 59.785 3.197 59.815 3.465 ;
      RECT 61.465 2.78 61.725 3.04 ;
      RECT 61.425 2.78 61.725 2.918 ;
      RECT 61.39 2.78 61.725 2.903 ;
      RECT 61.335 2.78 61.725 2.883 ;
      RECT 61.255 2.59 61.535 2.87 ;
      RECT 61.255 2.772 61.605 2.87 ;
      RECT 61.255 2.715 61.59 2.87 ;
      RECT 61.255 2.662 61.54 2.87 ;
      RECT 59.085 2.59 59.28 3.375 ;
      RECT 59.165 1.205 59.28 3.375 ;
      RECT 59.02 3.115 59.08 3.375 ;
      RECT 60.39 2.635 60.65 2.895 ;
      RECT 59.075 2.59 59.28 2.87 ;
      RECT 60.385 2.645 60.65 2.83 ;
      RECT 60.1 2.62 60.11 2.77 ;
      RECT 59.335 1.205 59.415 1.55 ;
      RECT 59.07 1.205 59.28 1.55 ;
      RECT 60.375 2.645 60.385 2.829 ;
      RECT 60.365 2.644 60.375 2.826 ;
      RECT 60.356 2.643 60.365 2.824 ;
      RECT 60.27 2.639 60.356 2.814 ;
      RECT 60.196 2.631 60.27 2.796 ;
      RECT 60.11 2.624 60.196 2.779 ;
      RECT 60.05 2.62 60.1 2.769 ;
      RECT 60.015 2.619 60.05 2.766 ;
      RECT 59.96 2.619 60.015 2.768 ;
      RECT 59.925 2.619 59.96 2.772 ;
      RECT 59.839 2.618 59.925 2.779 ;
      RECT 59.753 2.617 59.839 2.789 ;
      RECT 59.667 2.616 59.753 2.8 ;
      RECT 59.581 2.616 59.667 2.81 ;
      RECT 59.495 2.615 59.581 2.82 ;
      RECT 59.46 2.615 59.495 2.86 ;
      RECT 59.455 2.615 59.46 2.903 ;
      RECT 59.43 2.615 59.455 2.92 ;
      RECT 59.355 2.615 59.43 2.935 ;
      RECT 59.335 2.59 59.355 2.948 ;
      RECT 59.33 1.205 59.335 2.958 ;
      RECT 59.305 1.205 59.33 3 ;
      RECT 59.28 1.205 59.305 3.078 ;
      RECT 59.08 2.997 59.085 3.375 ;
      RECT 58.415 2.949 58.43 3.405 ;
      RECT 58.41 3.021 58.516 3.403 ;
      RECT 58.43 2.115 58.565 3.401 ;
      RECT 58.415 2.965 58.57 3.4 ;
      RECT 58.415 3.015 58.575 3.398 ;
      RECT 58.4 3.08 58.575 3.397 ;
      RECT 58.41 3.072 58.58 3.394 ;
      RECT 58.39 3.12 58.58 3.389 ;
      RECT 58.39 3.12 58.595 3.386 ;
      RECT 58.385 3.12 58.595 3.383 ;
      RECT 58.36 3.12 58.62 3.38 ;
      RECT 58.43 2.115 58.59 2.768 ;
      RECT 58.425 2.115 58.59 2.74 ;
      RECT 58.42 2.115 58.59 2.568 ;
      RECT 58.42 2.115 58.61 2.508 ;
      RECT 58.375 2.115 58.635 2.375 ;
      RECT 57.855 2.59 58.135 2.87 ;
      RECT 57.845 2.605 58.135 2.865 ;
      RECT 57.8 2.667 58.135 2.863 ;
      RECT 57.875 2.582 58.04 2.87 ;
      RECT 57.875 2.567 57.996 2.87 ;
      RECT 57.91 2.56 57.996 2.87 ;
      RECT 57.375 3.71 57.655 3.99 ;
      RECT 57.335 3.672 57.63 3.783 ;
      RECT 57.32 3.622 57.61 3.678 ;
      RECT 57.265 3.385 57.525 3.645 ;
      RECT 57.265 3.587 57.605 3.645 ;
      RECT 57.265 3.527 57.6 3.645 ;
      RECT 57.265 3.477 57.58 3.645 ;
      RECT 57.265 3.457 57.575 3.645 ;
      RECT 57.265 3.435 57.57 3.645 ;
      RECT 57.265 3.42 57.54 3.645 ;
      RECT 52.995 6.225 53.315 6.545 ;
      RECT 53.025 5.695 53.195 6.545 ;
      RECT 53.025 5.695 53.2 6.045 ;
      RECT 53.025 5.695 54 5.87 ;
      RECT 53.825 1.965 54 5.87 ;
      RECT 53.77 1.965 54.12 2.315 ;
      RECT 53.795 6.655 54.12 6.98 ;
      RECT 52.68 6.745 54.12 6.915 ;
      RECT 52.68 2.395 52.84 6.915 ;
      RECT 52.995 2.365 53.315 2.685 ;
      RECT 52.68 2.395 53.315 2.565 ;
      RECT 51.35 1.14 51.725 1.51 ;
      RECT 43.27 0.96 43.645 1.33 ;
      RECT 41.835 0.96 42.21 1.33 ;
      RECT 41.835 1.08 51.655 1.25 ;
      RECT 45.955 4.36 51.635 4.53 ;
      RECT 51.465 3.425 51.635 4.53 ;
      RECT 45.765 3.6 45.79 4.53 ;
      RECT 46.02 3.71 46.05 3.99 ;
      RECT 45.725 3.6 45.79 3.86 ;
      RECT 51.375 3.43 51.725 3.78 ;
      RECT 45.555 2.225 45.59 2.485 ;
      RECT 45.33 2.225 45.39 2.485 ;
      RECT 46.01 3.69 46.02 3.99 ;
      RECT 46.005 3.65 46.01 3.99 ;
      RECT 45.99 3.605 46.005 3.99 ;
      RECT 45.985 3.57 45.99 3.99 ;
      RECT 45.98 3.55 45.985 3.99 ;
      RECT 45.955 3.487 45.98 3.99 ;
      RECT 45.95 3.425 45.955 4.53 ;
      RECT 45.93 3.375 45.95 4.53 ;
      RECT 45.92 3.305 45.93 4.53 ;
      RECT 45.875 3.245 45.92 4.53 ;
      RECT 45.79 3.206 45.875 4.53 ;
      RECT 45.785 3.197 45.79 3.57 ;
      RECT 45.775 3.196 45.785 3.553 ;
      RECT 45.75 3.177 45.775 3.523 ;
      RECT 45.745 3.152 45.75 3.502 ;
      RECT 45.735 3.13 45.745 3.493 ;
      RECT 45.73 3.101 45.735 3.483 ;
      RECT 45.69 3.027 45.73 3.455 ;
      RECT 45.67 2.928 45.69 3.42 ;
      RECT 45.655 2.864 45.67 3.403 ;
      RECT 45.625 2.788 45.655 3.375 ;
      RECT 45.605 2.703 45.625 3.348 ;
      RECT 45.565 2.599 45.605 3.255 ;
      RECT 45.56 2.52 45.565 3.163 ;
      RECT 45.555 2.503 45.56 3.14 ;
      RECT 45.55 2.225 45.555 3.12 ;
      RECT 45.52 2.225 45.55 3.058 ;
      RECT 45.515 2.225 45.52 2.99 ;
      RECT 45.505 2.225 45.515 2.955 ;
      RECT 45.495 2.225 45.505 2.92 ;
      RECT 45.43 2.225 45.495 2.775 ;
      RECT 45.425 2.225 45.43 2.645 ;
      RECT 45.395 2.225 45.425 2.578 ;
      RECT 45.39 2.225 45.395 2.503 ;
      RECT 49.725 2.16 49.985 2.42 ;
      RECT 49.72 2.16 49.985 2.368 ;
      RECT 49.715 2.16 49.985 2.338 ;
      RECT 49.69 2.03 49.97 2.31 ;
      RECT 38.25 6.66 38.6 7.01 ;
      RECT 49.225 6.615 49.575 6.965 ;
      RECT 38.25 6.69 49.575 6.89 ;
      RECT 48.73 3.71 49.01 3.99 ;
      RECT 48.77 3.665 49.035 3.925 ;
      RECT 48.76 3.7 49.035 3.925 ;
      RECT 48.765 3.685 49.01 3.99 ;
      RECT 48.77 3.662 48.98 3.99 ;
      RECT 48.77 3.66 48.965 3.99 ;
      RECT 48.81 3.65 48.965 3.99 ;
      RECT 48.78 3.655 48.965 3.99 ;
      RECT 48.81 3.647 48.91 3.99 ;
      RECT 48.835 3.64 48.91 3.99 ;
      RECT 48.815 3.642 48.91 3.99 ;
      RECT 48.145 3.155 48.405 3.415 ;
      RECT 48.195 3.147 48.385 3.415 ;
      RECT 48.2 3.067 48.385 3.415 ;
      RECT 48.32 2.455 48.385 3.415 ;
      RECT 48.225 2.852 48.385 3.415 ;
      RECT 48.3 2.54 48.385 3.415 ;
      RECT 48.335 2.165 48.471 2.893 ;
      RECT 48.28 2.662 48.471 2.893 ;
      RECT 48.295 2.602 48.385 3.415 ;
      RECT 48.335 2.165 48.495 2.558 ;
      RECT 48.335 2.165 48.505 2.455 ;
      RECT 48.325 2.165 48.585 2.425 ;
      RECT 47.73 3.71 48.01 3.99 ;
      RECT 47.75 3.67 48.01 3.99 ;
      RECT 47.39 3.625 47.495 3.885 ;
      RECT 47.245 2.115 47.335 2.375 ;
      RECT 47.785 3.18 47.79 3.22 ;
      RECT 47.78 3.17 47.785 3.305 ;
      RECT 47.775 3.16 47.78 3.398 ;
      RECT 47.765 3.14 47.775 3.454 ;
      RECT 47.685 3.068 47.765 3.534 ;
      RECT 47.72 3.712 47.73 3.937 ;
      RECT 47.715 3.709 47.72 3.932 ;
      RECT 47.7 3.706 47.715 3.925 ;
      RECT 47.665 3.7 47.7 3.907 ;
      RECT 47.68 3.003 47.685 3.608 ;
      RECT 47.66 2.954 47.68 3.623 ;
      RECT 47.65 3.687 47.665 3.89 ;
      RECT 47.655 2.896 47.66 3.638 ;
      RECT 47.65 2.874 47.655 3.648 ;
      RECT 47.615 2.784 47.65 3.885 ;
      RECT 47.6 2.662 47.615 3.885 ;
      RECT 47.595 2.615 47.6 3.885 ;
      RECT 47.57 2.54 47.595 3.885 ;
      RECT 47.555 2.455 47.57 3.885 ;
      RECT 47.55 2.402 47.555 3.885 ;
      RECT 47.545 2.382 47.55 3.885 ;
      RECT 47.54 2.357 47.545 3.119 ;
      RECT 47.525 3.317 47.545 3.885 ;
      RECT 47.535 2.335 47.54 3.096 ;
      RECT 47.525 2.287 47.535 3.061 ;
      RECT 47.52 2.25 47.525 3.027 ;
      RECT 47.52 3.397 47.525 3.885 ;
      RECT 47.505 2.227 47.52 2.982 ;
      RECT 47.5 3.495 47.52 3.885 ;
      RECT 47.45 2.115 47.505 2.824 ;
      RECT 47.495 3.617 47.5 3.885 ;
      RECT 47.435 2.115 47.45 2.663 ;
      RECT 47.43 2.115 47.435 2.615 ;
      RECT 47.425 2.115 47.43 2.603 ;
      RECT 47.38 2.115 47.425 2.54 ;
      RECT 47.355 2.115 47.38 2.458 ;
      RECT 47.34 2.115 47.355 2.41 ;
      RECT 47.335 2.115 47.34 2.38 ;
      RECT 46.66 3.565 46.705 3.825 ;
      RECT 46.565 2.1 46.71 2.36 ;
      RECT 47.07 2.722 47.08 2.813 ;
      RECT 47.055 2.66 47.07 2.869 ;
      RECT 47.05 2.607 47.055 2.915 ;
      RECT 47 2.554 47.05 3.041 ;
      RECT 46.995 2.509 47 3.188 ;
      RECT 46.985 2.497 46.995 3.23 ;
      RECT 46.95 2.461 46.985 3.335 ;
      RECT 46.945 2.429 46.95 3.441 ;
      RECT 46.93 2.411 46.945 3.486 ;
      RECT 46.925 2.394 46.93 2.72 ;
      RECT 46.92 2.775 46.93 3.543 ;
      RECT 46.915 2.38 46.925 2.693 ;
      RECT 46.91 2.83 46.92 3.825 ;
      RECT 46.905 2.366 46.915 2.678 ;
      RECT 46.905 2.88 46.91 3.825 ;
      RECT 46.89 2.343 46.905 2.658 ;
      RECT 46.87 3.002 46.905 3.825 ;
      RECT 46.885 2.325 46.89 2.64 ;
      RECT 46.88 2.317 46.885 2.63 ;
      RECT 46.85 2.285 46.88 2.594 ;
      RECT 46.86 3.13 46.87 3.825 ;
      RECT 46.855 3.157 46.86 3.825 ;
      RECT 46.85 3.207 46.855 3.825 ;
      RECT 46.84 2.251 46.85 2.559 ;
      RECT 46.8 3.275 46.85 3.825 ;
      RECT 46.825 2.228 46.84 2.535 ;
      RECT 46.8 2.1 46.825 2.498 ;
      RECT 46.795 2.1 46.8 2.47 ;
      RECT 46.765 3.375 46.8 3.825 ;
      RECT 46.79 2.1 46.795 2.463 ;
      RECT 46.785 2.1 46.79 2.453 ;
      RECT 46.77 2.1 46.785 2.438 ;
      RECT 46.755 2.1 46.77 2.41 ;
      RECT 46.72 3.48 46.765 3.825 ;
      RECT 46.74 2.1 46.755 2.383 ;
      RECT 46.71 2.1 46.74 2.368 ;
      RECT 46.705 3.552 46.72 3.825 ;
      RECT 46.63 2.635 46.67 2.895 ;
      RECT 46.405 2.582 46.41 2.84 ;
      RECT 42.36 2.06 42.62 2.32 ;
      RECT 42.36 2.085 42.635 2.3 ;
      RECT 44.75 1.91 44.755 2.055 ;
      RECT 46.62 2.63 46.63 2.895 ;
      RECT 46.6 2.622 46.62 2.895 ;
      RECT 46.582 2.618 46.6 2.895 ;
      RECT 46.496 2.607 46.582 2.895 ;
      RECT 46.41 2.59 46.496 2.895 ;
      RECT 46.355 2.577 46.405 2.825 ;
      RECT 46.321 2.569 46.355 2.8 ;
      RECT 46.235 2.558 46.321 2.765 ;
      RECT 46.2 2.535 46.235 2.73 ;
      RECT 46.19 2.497 46.2 2.716 ;
      RECT 46.185 2.47 46.19 2.712 ;
      RECT 46.18 2.457 46.185 2.709 ;
      RECT 46.17 2.437 46.18 2.705 ;
      RECT 46.165 2.412 46.17 2.701 ;
      RECT 46.14 2.367 46.165 2.695 ;
      RECT 46.13 2.308 46.14 2.687 ;
      RECT 46.12 2.276 46.13 2.678 ;
      RECT 46.1 2.228 46.12 2.658 ;
      RECT 46.095 2.188 46.1 2.628 ;
      RECT 46.08 2.162 46.095 2.602 ;
      RECT 46.075 2.14 46.08 2.578 ;
      RECT 46.06 2.112 46.075 2.554 ;
      RECT 46.045 2.085 46.06 2.518 ;
      RECT 46.03 2.062 46.045 2.48 ;
      RECT 46.025 2.052 46.03 2.455 ;
      RECT 46.015 2.045 46.025 2.438 ;
      RECT 46 2.032 46.015 2.408 ;
      RECT 45.995 2.022 46 2.383 ;
      RECT 45.99 2.017 45.995 2.37 ;
      RECT 45.98 2.01 45.99 2.35 ;
      RECT 45.975 2.003 45.98 2.335 ;
      RECT 45.95 1.996 45.975 2.293 ;
      RECT 45.935 1.986 45.95 2.243 ;
      RECT 45.925 1.981 45.935 2.213 ;
      RECT 45.915 1.977 45.925 2.188 ;
      RECT 45.9 1.974 45.915 2.178 ;
      RECT 45.85 1.971 45.9 2.163 ;
      RECT 45.83 1.969 45.85 2.148 ;
      RECT 45.781 1.967 45.83 2.143 ;
      RECT 45.695 1.963 45.781 2.138 ;
      RECT 45.656 1.96 45.695 2.134 ;
      RECT 45.57 1.956 45.656 2.129 ;
      RECT 45.52 1.953 45.57 2.123 ;
      RECT 45.471 1.95 45.52 2.118 ;
      RECT 45.385 1.947 45.471 2.113 ;
      RECT 45.381 1.945 45.385 2.11 ;
      RECT 45.295 1.942 45.381 2.105 ;
      RECT 45.246 1.938 45.295 2.098 ;
      RECT 45.16 1.935 45.246 2.093 ;
      RECT 45.136 1.932 45.16 2.089 ;
      RECT 45.05 1.93 45.136 2.084 ;
      RECT 44.985 1.926 45.05 2.077 ;
      RECT 44.982 1.925 44.985 2.074 ;
      RECT 44.896 1.922 44.982 2.071 ;
      RECT 44.81 1.916 44.896 2.064 ;
      RECT 44.78 1.912 44.81 2.06 ;
      RECT 44.755 1.91 44.78 2.058 ;
      RECT 44.7 1.907 44.75 2.055 ;
      RECT 44.62 1.906 44.7 2.055 ;
      RECT 44.565 1.908 44.62 2.058 ;
      RECT 44.55 1.909 44.565 2.062 ;
      RECT 44.495 1.917 44.55 2.072 ;
      RECT 44.465 1.925 44.495 2.085 ;
      RECT 44.446 1.926 44.465 2.091 ;
      RECT 44.36 1.929 44.446 2.096 ;
      RECT 44.29 1.934 44.36 2.105 ;
      RECT 44.271 1.937 44.29 2.111 ;
      RECT 44.185 1.941 44.271 2.116 ;
      RECT 44.145 1.945 44.185 2.123 ;
      RECT 44.136 1.947 44.145 2.126 ;
      RECT 44.05 1.951 44.136 2.131 ;
      RECT 44.047 1.954 44.05 2.135 ;
      RECT 43.961 1.957 44.047 2.139 ;
      RECT 43.875 1.963 43.961 2.147 ;
      RECT 43.851 1.967 43.875 2.151 ;
      RECT 43.765 1.971 43.851 2.156 ;
      RECT 43.72 1.976 43.765 2.163 ;
      RECT 43.64 1.981 43.72 2.17 ;
      RECT 43.56 1.987 43.64 2.185 ;
      RECT 43.535 1.991 43.56 2.198 ;
      RECT 43.47 1.994 43.535 2.21 ;
      RECT 43.415 1.999 43.47 2.225 ;
      RECT 43.385 2.002 43.415 2.243 ;
      RECT 43.375 2.004 43.385 2.256 ;
      RECT 43.315 2.019 43.375 2.266 ;
      RECT 43.3 2.036 43.315 2.275 ;
      RECT 43.295 2.045 43.3 2.275 ;
      RECT 43.285 2.055 43.295 2.275 ;
      RECT 43.275 2.072 43.285 2.275 ;
      RECT 43.255 2.082 43.275 2.276 ;
      RECT 43.21 2.092 43.255 2.277 ;
      RECT 43.175 2.101 43.21 2.279 ;
      RECT 43.11 2.106 43.175 2.281 ;
      RECT 43.03 2.107 43.11 2.284 ;
      RECT 43.026 2.105 43.03 2.285 ;
      RECT 42.94 2.102 43.026 2.287 ;
      RECT 42.893 2.099 42.94 2.289 ;
      RECT 42.807 2.095 42.893 2.292 ;
      RECT 42.721 2.091 42.807 2.295 ;
      RECT 42.635 2.087 42.721 2.299 ;
      RECT 44.57 3.15 44.85 3.43 ;
      RECT 44.61 3.13 44.87 3.39 ;
      RECT 44.6 3.14 44.87 3.39 ;
      RECT 44.61 3.067 44.825 3.43 ;
      RECT 44.665 2.99 44.82 3.43 ;
      RECT 44.67 2.775 44.82 3.43 ;
      RECT 44.66 2.577 44.81 2.828 ;
      RECT 44.65 2.577 44.81 2.695 ;
      RECT 44.645 2.455 44.805 2.598 ;
      RECT 44.63 2.455 44.805 2.503 ;
      RECT 44.625 2.165 44.8 2.48 ;
      RECT 44.61 2.165 44.8 2.45 ;
      RECT 44.57 2.165 44.83 2.425 ;
      RECT 44.48 3.635 44.56 3.895 ;
      RECT 43.885 2.355 43.89 2.62 ;
      RECT 43.765 2.355 43.89 2.615 ;
      RECT 44.44 3.6 44.48 3.895 ;
      RECT 44.395 3.522 44.44 3.895 ;
      RECT 44.375 3.45 44.395 3.895 ;
      RECT 44.365 3.402 44.375 3.895 ;
      RECT 44.33 3.335 44.365 3.895 ;
      RECT 44.3 3.235 44.33 3.895 ;
      RECT 44.28 3.16 44.3 3.695 ;
      RECT 44.27 3.11 44.28 3.65 ;
      RECT 44.265 3.087 44.27 3.623 ;
      RECT 44.26 3.072 44.265 3.61 ;
      RECT 44.255 3.057 44.26 3.588 ;
      RECT 44.25 3.042 44.255 3.57 ;
      RECT 44.225 2.997 44.25 3.525 ;
      RECT 44.215 2.945 44.225 3.468 ;
      RECT 44.205 2.915 44.215 3.435 ;
      RECT 44.195 2.88 44.205 3.403 ;
      RECT 44.16 2.812 44.195 3.335 ;
      RECT 44.155 2.751 44.16 3.27 ;
      RECT 44.145 2.739 44.155 3.25 ;
      RECT 44.14 2.727 44.145 3.23 ;
      RECT 44.135 2.719 44.14 3.218 ;
      RECT 44.13 2.711 44.135 3.198 ;
      RECT 44.12 2.699 44.13 3.17 ;
      RECT 44.11 2.683 44.12 3.14 ;
      RECT 44.085 2.655 44.11 3.078 ;
      RECT 44.075 2.626 44.085 3.023 ;
      RECT 44.06 2.605 44.075 2.983 ;
      RECT 44.055 2.589 44.06 2.955 ;
      RECT 44.05 2.577 44.055 2.945 ;
      RECT 44.045 2.572 44.05 2.918 ;
      RECT 44.04 2.565 44.045 2.905 ;
      RECT 44.025 2.548 44.04 2.878 ;
      RECT 44.015 2.355 44.025 2.838 ;
      RECT 44.005 2.355 44.015 2.805 ;
      RECT 43.995 2.355 44.005 2.78 ;
      RECT 43.925 2.355 43.995 2.715 ;
      RECT 43.915 2.355 43.925 2.663 ;
      RECT 43.9 2.355 43.915 2.645 ;
      RECT 43.89 2.355 43.9 2.63 ;
      RECT 43.72 3.225 43.98 3.485 ;
      RECT 42.255 3.26 42.26 3.467 ;
      RECT 41.89 3.15 41.965 3.465 ;
      RECT 41.705 3.205 41.86 3.465 ;
      RECT 41.89 3.15 41.995 3.43 ;
      RECT 43.705 3.322 43.72 3.483 ;
      RECT 43.68 3.33 43.705 3.488 ;
      RECT 43.655 3.337 43.68 3.493 ;
      RECT 43.592 3.348 43.655 3.502 ;
      RECT 43.506 3.367 43.592 3.519 ;
      RECT 43.42 3.389 43.506 3.538 ;
      RECT 43.405 3.402 43.42 3.549 ;
      RECT 43.365 3.41 43.405 3.556 ;
      RECT 43.345 3.415 43.365 3.563 ;
      RECT 43.307 3.416 43.345 3.566 ;
      RECT 43.221 3.419 43.307 3.567 ;
      RECT 43.135 3.423 43.221 3.568 ;
      RECT 43.086 3.425 43.135 3.57 ;
      RECT 43 3.425 43.086 3.572 ;
      RECT 42.96 3.42 43 3.574 ;
      RECT 42.95 3.414 42.96 3.575 ;
      RECT 42.91 3.409 42.95 3.572 ;
      RECT 42.9 3.402 42.91 3.568 ;
      RECT 42.885 3.398 42.9 3.566 ;
      RECT 42.868 3.394 42.885 3.564 ;
      RECT 42.782 3.384 42.868 3.556 ;
      RECT 42.696 3.366 42.782 3.542 ;
      RECT 42.61 3.349 42.696 3.528 ;
      RECT 42.585 3.337 42.61 3.519 ;
      RECT 42.515 3.327 42.585 3.512 ;
      RECT 42.47 3.315 42.515 3.503 ;
      RECT 42.41 3.302 42.47 3.495 ;
      RECT 42.405 3.294 42.41 3.49 ;
      RECT 42.37 3.289 42.405 3.488 ;
      RECT 42.315 3.28 42.37 3.481 ;
      RECT 42.275 3.269 42.315 3.473 ;
      RECT 42.26 3.262 42.275 3.469 ;
      RECT 42.24 3.255 42.255 3.466 ;
      RECT 42.225 3.245 42.24 3.464 ;
      RECT 42.21 3.232 42.225 3.461 ;
      RECT 42.185 3.215 42.21 3.457 ;
      RECT 42.17 3.197 42.185 3.454 ;
      RECT 42.145 3.15 42.17 3.452 ;
      RECT 42.121 3.15 42.145 3.449 ;
      RECT 42.035 3.15 42.121 3.441 ;
      RECT 41.995 3.15 42.035 3.433 ;
      RECT 41.86 3.197 41.89 3.465 ;
      RECT 43.54 2.78 43.8 3.04 ;
      RECT 43.5 2.78 43.8 2.918 ;
      RECT 43.465 2.78 43.8 2.903 ;
      RECT 43.41 2.78 43.8 2.883 ;
      RECT 43.33 2.59 43.61 2.87 ;
      RECT 43.33 2.772 43.68 2.87 ;
      RECT 43.33 2.715 43.665 2.87 ;
      RECT 43.33 2.662 43.615 2.87 ;
      RECT 41.16 2.59 41.355 3.375 ;
      RECT 41.24 1.205 41.355 3.375 ;
      RECT 41.095 3.115 41.155 3.375 ;
      RECT 42.465 2.635 42.725 2.895 ;
      RECT 41.15 2.59 41.355 2.87 ;
      RECT 42.46 2.645 42.725 2.83 ;
      RECT 42.175 2.62 42.185 2.77 ;
      RECT 41.41 1.205 41.49 1.55 ;
      RECT 41.145 1.205 41.355 1.55 ;
      RECT 42.45 2.645 42.46 2.829 ;
      RECT 42.44 2.644 42.45 2.826 ;
      RECT 42.431 2.643 42.44 2.824 ;
      RECT 42.345 2.639 42.431 2.814 ;
      RECT 42.271 2.631 42.345 2.796 ;
      RECT 42.185 2.624 42.271 2.779 ;
      RECT 42.125 2.62 42.175 2.769 ;
      RECT 42.09 2.619 42.125 2.766 ;
      RECT 42.035 2.619 42.09 2.768 ;
      RECT 42 2.619 42.035 2.772 ;
      RECT 41.914 2.618 42 2.779 ;
      RECT 41.828 2.617 41.914 2.789 ;
      RECT 41.742 2.616 41.828 2.8 ;
      RECT 41.656 2.616 41.742 2.81 ;
      RECT 41.57 2.615 41.656 2.82 ;
      RECT 41.535 2.615 41.57 2.86 ;
      RECT 41.53 2.615 41.535 2.903 ;
      RECT 41.505 2.615 41.53 2.92 ;
      RECT 41.43 2.615 41.505 2.935 ;
      RECT 41.41 2.59 41.43 2.948 ;
      RECT 41.405 1.205 41.41 2.958 ;
      RECT 41.38 1.205 41.405 3 ;
      RECT 41.355 1.205 41.38 3.078 ;
      RECT 41.155 2.997 41.16 3.375 ;
      RECT 40.49 2.949 40.505 3.405 ;
      RECT 40.485 3.021 40.591 3.403 ;
      RECT 40.505 2.115 40.64 3.401 ;
      RECT 40.49 2.965 40.645 3.4 ;
      RECT 40.49 3.015 40.65 3.398 ;
      RECT 40.475 3.08 40.65 3.397 ;
      RECT 40.485 3.072 40.655 3.394 ;
      RECT 40.465 3.12 40.655 3.389 ;
      RECT 40.465 3.12 40.67 3.386 ;
      RECT 40.46 3.12 40.67 3.383 ;
      RECT 40.435 3.12 40.695 3.38 ;
      RECT 40.505 2.115 40.665 2.768 ;
      RECT 40.5 2.115 40.665 2.74 ;
      RECT 40.495 2.115 40.665 2.568 ;
      RECT 40.495 2.115 40.685 2.508 ;
      RECT 40.45 2.115 40.71 2.375 ;
      RECT 39.93 2.59 40.21 2.87 ;
      RECT 39.92 2.605 40.21 2.865 ;
      RECT 39.875 2.667 40.21 2.863 ;
      RECT 39.95 2.582 40.115 2.87 ;
      RECT 39.95 2.567 40.071 2.87 ;
      RECT 39.985 2.56 40.071 2.87 ;
      RECT 39.45 3.71 39.73 3.99 ;
      RECT 39.41 3.672 39.705 3.783 ;
      RECT 39.395 3.622 39.685 3.678 ;
      RECT 39.34 3.385 39.6 3.645 ;
      RECT 39.34 3.587 39.68 3.645 ;
      RECT 39.34 3.527 39.675 3.645 ;
      RECT 39.34 3.477 39.655 3.645 ;
      RECT 39.34 3.457 39.65 3.645 ;
      RECT 39.34 3.435 39.645 3.645 ;
      RECT 39.34 3.42 39.615 3.645 ;
      RECT 35.07 6.225 35.39 6.545 ;
      RECT 35.1 5.695 35.27 6.545 ;
      RECT 35.1 5.695 35.275 6.045 ;
      RECT 35.1 5.695 36.075 5.87 ;
      RECT 35.9 1.965 36.075 5.87 ;
      RECT 35.845 1.965 36.195 2.315 ;
      RECT 35.87 6.655 36.195 6.98 ;
      RECT 34.755 6.745 36.195 6.915 ;
      RECT 34.755 2.395 34.915 6.915 ;
      RECT 35.07 2.365 35.39 2.685 ;
      RECT 34.755 2.395 35.39 2.565 ;
      RECT 33.425 1.14 33.8 1.51 ;
      RECT 25.345 0.96 25.72 1.33 ;
      RECT 23.91 0.96 24.285 1.33 ;
      RECT 23.91 1.08 33.73 1.25 ;
      RECT 28.03 4.36 33.71 4.53 ;
      RECT 33.54 3.425 33.71 4.53 ;
      RECT 27.84 3.6 27.865 4.53 ;
      RECT 28.095 3.71 28.125 3.99 ;
      RECT 27.8 3.6 27.865 3.86 ;
      RECT 33.45 3.43 33.8 3.78 ;
      RECT 27.63 2.225 27.665 2.485 ;
      RECT 27.405 2.225 27.465 2.485 ;
      RECT 28.085 3.69 28.095 3.99 ;
      RECT 28.08 3.65 28.085 3.99 ;
      RECT 28.065 3.605 28.08 3.99 ;
      RECT 28.06 3.57 28.065 3.99 ;
      RECT 28.055 3.55 28.06 3.99 ;
      RECT 28.03 3.487 28.055 3.99 ;
      RECT 28.025 3.425 28.03 4.53 ;
      RECT 28.005 3.375 28.025 4.53 ;
      RECT 27.995 3.305 28.005 4.53 ;
      RECT 27.95 3.245 27.995 4.53 ;
      RECT 27.865 3.206 27.95 4.53 ;
      RECT 27.86 3.197 27.865 3.57 ;
      RECT 27.85 3.196 27.86 3.553 ;
      RECT 27.825 3.177 27.85 3.523 ;
      RECT 27.82 3.152 27.825 3.502 ;
      RECT 27.81 3.13 27.82 3.493 ;
      RECT 27.805 3.101 27.81 3.483 ;
      RECT 27.765 3.027 27.805 3.455 ;
      RECT 27.745 2.928 27.765 3.42 ;
      RECT 27.73 2.864 27.745 3.403 ;
      RECT 27.7 2.788 27.73 3.375 ;
      RECT 27.68 2.703 27.7 3.348 ;
      RECT 27.64 2.599 27.68 3.255 ;
      RECT 27.635 2.52 27.64 3.163 ;
      RECT 27.63 2.503 27.635 3.14 ;
      RECT 27.625 2.225 27.63 3.12 ;
      RECT 27.595 2.225 27.625 3.058 ;
      RECT 27.59 2.225 27.595 2.99 ;
      RECT 27.58 2.225 27.59 2.955 ;
      RECT 27.57 2.225 27.58 2.92 ;
      RECT 27.505 2.225 27.57 2.775 ;
      RECT 27.5 2.225 27.505 2.645 ;
      RECT 27.47 2.225 27.5 2.578 ;
      RECT 27.465 2.225 27.47 2.503 ;
      RECT 31.8 2.16 32.06 2.42 ;
      RECT 31.795 2.16 32.06 2.368 ;
      RECT 31.79 2.16 32.06 2.338 ;
      RECT 31.765 2.03 32.045 2.31 ;
      RECT 20.325 6.655 20.675 7.005 ;
      RECT 31.295 6.61 31.645 6.96 ;
      RECT 20.325 6.685 31.645 6.885 ;
      RECT 30.805 3.71 31.085 3.99 ;
      RECT 30.845 3.665 31.11 3.925 ;
      RECT 30.835 3.7 31.11 3.925 ;
      RECT 30.84 3.685 31.085 3.99 ;
      RECT 30.845 3.662 31.055 3.99 ;
      RECT 30.845 3.66 31.04 3.99 ;
      RECT 30.885 3.65 31.04 3.99 ;
      RECT 30.855 3.655 31.04 3.99 ;
      RECT 30.885 3.647 30.985 3.99 ;
      RECT 30.91 3.64 30.985 3.99 ;
      RECT 30.89 3.642 30.985 3.99 ;
      RECT 30.22 3.155 30.48 3.415 ;
      RECT 30.27 3.147 30.46 3.415 ;
      RECT 30.275 3.067 30.46 3.415 ;
      RECT 30.395 2.455 30.46 3.415 ;
      RECT 30.3 2.852 30.46 3.415 ;
      RECT 30.375 2.54 30.46 3.415 ;
      RECT 30.41 2.165 30.546 2.893 ;
      RECT 30.355 2.662 30.546 2.893 ;
      RECT 30.37 2.602 30.46 3.415 ;
      RECT 30.41 2.165 30.57 2.558 ;
      RECT 30.41 2.165 30.58 2.455 ;
      RECT 30.4 2.165 30.66 2.425 ;
      RECT 29.805 3.71 30.085 3.99 ;
      RECT 29.825 3.67 30.085 3.99 ;
      RECT 29.465 3.625 29.57 3.885 ;
      RECT 29.32 2.115 29.41 2.375 ;
      RECT 29.86 3.18 29.865 3.22 ;
      RECT 29.855 3.17 29.86 3.305 ;
      RECT 29.85 3.16 29.855 3.398 ;
      RECT 29.84 3.14 29.85 3.454 ;
      RECT 29.76 3.068 29.84 3.534 ;
      RECT 29.795 3.712 29.805 3.937 ;
      RECT 29.79 3.709 29.795 3.932 ;
      RECT 29.775 3.706 29.79 3.925 ;
      RECT 29.74 3.7 29.775 3.907 ;
      RECT 29.755 3.003 29.76 3.608 ;
      RECT 29.735 2.954 29.755 3.623 ;
      RECT 29.725 3.687 29.74 3.89 ;
      RECT 29.73 2.896 29.735 3.638 ;
      RECT 29.725 2.874 29.73 3.648 ;
      RECT 29.69 2.784 29.725 3.885 ;
      RECT 29.675 2.662 29.69 3.885 ;
      RECT 29.67 2.615 29.675 3.885 ;
      RECT 29.645 2.54 29.67 3.885 ;
      RECT 29.63 2.455 29.645 3.885 ;
      RECT 29.625 2.402 29.63 3.885 ;
      RECT 29.62 2.382 29.625 3.885 ;
      RECT 29.615 2.357 29.62 3.119 ;
      RECT 29.6 3.317 29.62 3.885 ;
      RECT 29.61 2.335 29.615 3.096 ;
      RECT 29.6 2.287 29.61 3.061 ;
      RECT 29.595 2.25 29.6 3.027 ;
      RECT 29.595 3.397 29.6 3.885 ;
      RECT 29.58 2.227 29.595 2.982 ;
      RECT 29.575 3.495 29.595 3.885 ;
      RECT 29.525 2.115 29.58 2.824 ;
      RECT 29.57 3.617 29.575 3.885 ;
      RECT 29.51 2.115 29.525 2.663 ;
      RECT 29.505 2.115 29.51 2.615 ;
      RECT 29.5 2.115 29.505 2.603 ;
      RECT 29.455 2.115 29.5 2.54 ;
      RECT 29.43 2.115 29.455 2.458 ;
      RECT 29.415 2.115 29.43 2.41 ;
      RECT 29.41 2.115 29.415 2.38 ;
      RECT 28.735 3.565 28.78 3.825 ;
      RECT 28.64 2.1 28.785 2.36 ;
      RECT 29.145 2.722 29.155 2.813 ;
      RECT 29.13 2.66 29.145 2.869 ;
      RECT 29.125 2.607 29.13 2.915 ;
      RECT 29.075 2.554 29.125 3.041 ;
      RECT 29.07 2.509 29.075 3.188 ;
      RECT 29.06 2.497 29.07 3.23 ;
      RECT 29.025 2.461 29.06 3.335 ;
      RECT 29.02 2.429 29.025 3.441 ;
      RECT 29.005 2.411 29.02 3.486 ;
      RECT 29 2.394 29.005 2.72 ;
      RECT 28.995 2.775 29.005 3.543 ;
      RECT 28.99 2.38 29 2.693 ;
      RECT 28.985 2.83 28.995 3.825 ;
      RECT 28.98 2.366 28.99 2.678 ;
      RECT 28.98 2.88 28.985 3.825 ;
      RECT 28.965 2.343 28.98 2.658 ;
      RECT 28.945 3.002 28.98 3.825 ;
      RECT 28.96 2.325 28.965 2.64 ;
      RECT 28.955 2.317 28.96 2.63 ;
      RECT 28.925 2.285 28.955 2.594 ;
      RECT 28.935 3.13 28.945 3.825 ;
      RECT 28.93 3.157 28.935 3.825 ;
      RECT 28.925 3.207 28.93 3.825 ;
      RECT 28.915 2.251 28.925 2.559 ;
      RECT 28.875 3.275 28.925 3.825 ;
      RECT 28.9 2.228 28.915 2.535 ;
      RECT 28.875 2.1 28.9 2.498 ;
      RECT 28.87 2.1 28.875 2.47 ;
      RECT 28.84 3.375 28.875 3.825 ;
      RECT 28.865 2.1 28.87 2.463 ;
      RECT 28.86 2.1 28.865 2.453 ;
      RECT 28.845 2.1 28.86 2.438 ;
      RECT 28.83 2.1 28.845 2.41 ;
      RECT 28.795 3.48 28.84 3.825 ;
      RECT 28.815 2.1 28.83 2.383 ;
      RECT 28.785 2.1 28.815 2.368 ;
      RECT 28.78 3.552 28.795 3.825 ;
      RECT 28.705 2.635 28.745 2.895 ;
      RECT 28.48 2.582 28.485 2.84 ;
      RECT 24.435 2.06 24.695 2.32 ;
      RECT 24.435 2.085 24.71 2.3 ;
      RECT 26.825 1.91 26.83 2.055 ;
      RECT 28.695 2.63 28.705 2.895 ;
      RECT 28.675 2.622 28.695 2.895 ;
      RECT 28.657 2.618 28.675 2.895 ;
      RECT 28.571 2.607 28.657 2.895 ;
      RECT 28.485 2.59 28.571 2.895 ;
      RECT 28.43 2.577 28.48 2.825 ;
      RECT 28.396 2.569 28.43 2.8 ;
      RECT 28.31 2.558 28.396 2.765 ;
      RECT 28.275 2.535 28.31 2.73 ;
      RECT 28.265 2.497 28.275 2.716 ;
      RECT 28.26 2.47 28.265 2.712 ;
      RECT 28.255 2.457 28.26 2.709 ;
      RECT 28.245 2.437 28.255 2.705 ;
      RECT 28.24 2.412 28.245 2.701 ;
      RECT 28.215 2.367 28.24 2.695 ;
      RECT 28.205 2.308 28.215 2.687 ;
      RECT 28.195 2.276 28.205 2.678 ;
      RECT 28.175 2.228 28.195 2.658 ;
      RECT 28.17 2.188 28.175 2.628 ;
      RECT 28.155 2.162 28.17 2.602 ;
      RECT 28.15 2.14 28.155 2.578 ;
      RECT 28.135 2.112 28.15 2.554 ;
      RECT 28.12 2.085 28.135 2.518 ;
      RECT 28.105 2.062 28.12 2.48 ;
      RECT 28.1 2.052 28.105 2.455 ;
      RECT 28.09 2.045 28.1 2.438 ;
      RECT 28.075 2.032 28.09 2.408 ;
      RECT 28.07 2.022 28.075 2.383 ;
      RECT 28.065 2.017 28.07 2.37 ;
      RECT 28.055 2.01 28.065 2.35 ;
      RECT 28.05 2.003 28.055 2.335 ;
      RECT 28.025 1.996 28.05 2.293 ;
      RECT 28.01 1.986 28.025 2.243 ;
      RECT 28 1.981 28.01 2.213 ;
      RECT 27.99 1.977 28 2.188 ;
      RECT 27.975 1.974 27.99 2.178 ;
      RECT 27.925 1.971 27.975 2.163 ;
      RECT 27.905 1.969 27.925 2.148 ;
      RECT 27.856 1.967 27.905 2.143 ;
      RECT 27.77 1.963 27.856 2.138 ;
      RECT 27.731 1.96 27.77 2.134 ;
      RECT 27.645 1.956 27.731 2.129 ;
      RECT 27.595 1.953 27.645 2.123 ;
      RECT 27.546 1.95 27.595 2.118 ;
      RECT 27.46 1.947 27.546 2.113 ;
      RECT 27.456 1.945 27.46 2.11 ;
      RECT 27.37 1.942 27.456 2.105 ;
      RECT 27.321 1.938 27.37 2.098 ;
      RECT 27.235 1.935 27.321 2.093 ;
      RECT 27.211 1.932 27.235 2.089 ;
      RECT 27.125 1.93 27.211 2.084 ;
      RECT 27.06 1.926 27.125 2.077 ;
      RECT 27.057 1.925 27.06 2.074 ;
      RECT 26.971 1.922 27.057 2.071 ;
      RECT 26.885 1.916 26.971 2.064 ;
      RECT 26.855 1.912 26.885 2.06 ;
      RECT 26.83 1.91 26.855 2.058 ;
      RECT 26.775 1.907 26.825 2.055 ;
      RECT 26.695 1.906 26.775 2.055 ;
      RECT 26.64 1.908 26.695 2.058 ;
      RECT 26.625 1.909 26.64 2.062 ;
      RECT 26.57 1.917 26.625 2.072 ;
      RECT 26.54 1.925 26.57 2.085 ;
      RECT 26.521 1.926 26.54 2.091 ;
      RECT 26.435 1.929 26.521 2.096 ;
      RECT 26.365 1.934 26.435 2.105 ;
      RECT 26.346 1.937 26.365 2.111 ;
      RECT 26.26 1.941 26.346 2.116 ;
      RECT 26.22 1.945 26.26 2.123 ;
      RECT 26.211 1.947 26.22 2.126 ;
      RECT 26.125 1.951 26.211 2.131 ;
      RECT 26.122 1.954 26.125 2.135 ;
      RECT 26.036 1.957 26.122 2.139 ;
      RECT 25.95 1.963 26.036 2.147 ;
      RECT 25.926 1.967 25.95 2.151 ;
      RECT 25.84 1.971 25.926 2.156 ;
      RECT 25.795 1.976 25.84 2.163 ;
      RECT 25.715 1.981 25.795 2.17 ;
      RECT 25.635 1.987 25.715 2.185 ;
      RECT 25.61 1.991 25.635 2.198 ;
      RECT 25.545 1.994 25.61 2.21 ;
      RECT 25.49 1.999 25.545 2.225 ;
      RECT 25.46 2.002 25.49 2.243 ;
      RECT 25.45 2.004 25.46 2.256 ;
      RECT 25.39 2.019 25.45 2.266 ;
      RECT 25.375 2.036 25.39 2.275 ;
      RECT 25.37 2.045 25.375 2.275 ;
      RECT 25.36 2.055 25.37 2.275 ;
      RECT 25.35 2.072 25.36 2.275 ;
      RECT 25.33 2.082 25.35 2.276 ;
      RECT 25.285 2.092 25.33 2.277 ;
      RECT 25.25 2.101 25.285 2.279 ;
      RECT 25.185 2.106 25.25 2.281 ;
      RECT 25.105 2.107 25.185 2.284 ;
      RECT 25.101 2.105 25.105 2.285 ;
      RECT 25.015 2.102 25.101 2.287 ;
      RECT 24.968 2.099 25.015 2.289 ;
      RECT 24.882 2.095 24.968 2.292 ;
      RECT 24.796 2.091 24.882 2.295 ;
      RECT 24.71 2.087 24.796 2.299 ;
      RECT 26.645 3.15 26.925 3.43 ;
      RECT 26.685 3.13 26.945 3.39 ;
      RECT 26.675 3.14 26.945 3.39 ;
      RECT 26.685 3.067 26.9 3.43 ;
      RECT 26.74 2.99 26.895 3.43 ;
      RECT 26.745 2.775 26.895 3.43 ;
      RECT 26.735 2.577 26.885 2.828 ;
      RECT 26.725 2.577 26.885 2.695 ;
      RECT 26.72 2.455 26.88 2.598 ;
      RECT 26.705 2.455 26.88 2.503 ;
      RECT 26.7 2.165 26.875 2.48 ;
      RECT 26.685 2.165 26.875 2.45 ;
      RECT 26.645 2.165 26.905 2.425 ;
      RECT 26.555 3.635 26.635 3.895 ;
      RECT 25.96 2.355 25.965 2.62 ;
      RECT 25.84 2.355 25.965 2.615 ;
      RECT 26.515 3.6 26.555 3.895 ;
      RECT 26.47 3.522 26.515 3.895 ;
      RECT 26.45 3.45 26.47 3.895 ;
      RECT 26.44 3.402 26.45 3.895 ;
      RECT 26.405 3.335 26.44 3.895 ;
      RECT 26.375 3.235 26.405 3.895 ;
      RECT 26.355 3.16 26.375 3.695 ;
      RECT 26.345 3.11 26.355 3.65 ;
      RECT 26.34 3.087 26.345 3.623 ;
      RECT 26.335 3.072 26.34 3.61 ;
      RECT 26.33 3.057 26.335 3.588 ;
      RECT 26.325 3.042 26.33 3.57 ;
      RECT 26.3 2.997 26.325 3.525 ;
      RECT 26.29 2.945 26.3 3.468 ;
      RECT 26.28 2.915 26.29 3.435 ;
      RECT 26.27 2.88 26.28 3.403 ;
      RECT 26.235 2.812 26.27 3.335 ;
      RECT 26.23 2.751 26.235 3.27 ;
      RECT 26.22 2.739 26.23 3.25 ;
      RECT 26.215 2.727 26.22 3.23 ;
      RECT 26.21 2.719 26.215 3.218 ;
      RECT 26.205 2.711 26.21 3.198 ;
      RECT 26.195 2.699 26.205 3.17 ;
      RECT 26.185 2.683 26.195 3.14 ;
      RECT 26.16 2.655 26.185 3.078 ;
      RECT 26.15 2.626 26.16 3.023 ;
      RECT 26.135 2.605 26.15 2.983 ;
      RECT 26.13 2.589 26.135 2.955 ;
      RECT 26.125 2.577 26.13 2.945 ;
      RECT 26.12 2.572 26.125 2.918 ;
      RECT 26.115 2.565 26.12 2.905 ;
      RECT 26.1 2.548 26.115 2.878 ;
      RECT 26.09 2.355 26.1 2.838 ;
      RECT 26.08 2.355 26.09 2.805 ;
      RECT 26.07 2.355 26.08 2.78 ;
      RECT 26 2.355 26.07 2.715 ;
      RECT 25.99 2.355 26 2.663 ;
      RECT 25.975 2.355 25.99 2.645 ;
      RECT 25.965 2.355 25.975 2.63 ;
      RECT 25.795 3.225 26.055 3.485 ;
      RECT 24.33 3.26 24.335 3.467 ;
      RECT 23.965 3.15 24.04 3.465 ;
      RECT 23.78 3.205 23.935 3.465 ;
      RECT 23.965 3.15 24.07 3.43 ;
      RECT 25.78 3.322 25.795 3.483 ;
      RECT 25.755 3.33 25.78 3.488 ;
      RECT 25.73 3.337 25.755 3.493 ;
      RECT 25.667 3.348 25.73 3.502 ;
      RECT 25.581 3.367 25.667 3.519 ;
      RECT 25.495 3.389 25.581 3.538 ;
      RECT 25.48 3.402 25.495 3.549 ;
      RECT 25.44 3.41 25.48 3.556 ;
      RECT 25.42 3.415 25.44 3.563 ;
      RECT 25.382 3.416 25.42 3.566 ;
      RECT 25.296 3.419 25.382 3.567 ;
      RECT 25.21 3.423 25.296 3.568 ;
      RECT 25.161 3.425 25.21 3.57 ;
      RECT 25.075 3.425 25.161 3.572 ;
      RECT 25.035 3.42 25.075 3.574 ;
      RECT 25.025 3.414 25.035 3.575 ;
      RECT 24.985 3.409 25.025 3.572 ;
      RECT 24.975 3.402 24.985 3.568 ;
      RECT 24.96 3.398 24.975 3.566 ;
      RECT 24.943 3.394 24.96 3.564 ;
      RECT 24.857 3.384 24.943 3.556 ;
      RECT 24.771 3.366 24.857 3.542 ;
      RECT 24.685 3.349 24.771 3.528 ;
      RECT 24.66 3.337 24.685 3.519 ;
      RECT 24.59 3.327 24.66 3.512 ;
      RECT 24.545 3.315 24.59 3.503 ;
      RECT 24.485 3.302 24.545 3.495 ;
      RECT 24.48 3.294 24.485 3.49 ;
      RECT 24.445 3.289 24.48 3.488 ;
      RECT 24.39 3.28 24.445 3.481 ;
      RECT 24.35 3.269 24.39 3.473 ;
      RECT 24.335 3.262 24.35 3.469 ;
      RECT 24.315 3.255 24.33 3.466 ;
      RECT 24.3 3.245 24.315 3.464 ;
      RECT 24.285 3.232 24.3 3.461 ;
      RECT 24.26 3.215 24.285 3.457 ;
      RECT 24.245 3.197 24.26 3.454 ;
      RECT 24.22 3.15 24.245 3.452 ;
      RECT 24.196 3.15 24.22 3.449 ;
      RECT 24.11 3.15 24.196 3.441 ;
      RECT 24.07 3.15 24.11 3.433 ;
      RECT 23.935 3.197 23.965 3.465 ;
      RECT 25.615 2.78 25.875 3.04 ;
      RECT 25.575 2.78 25.875 2.918 ;
      RECT 25.54 2.78 25.875 2.903 ;
      RECT 25.485 2.78 25.875 2.883 ;
      RECT 25.405 2.59 25.685 2.87 ;
      RECT 25.405 2.772 25.755 2.87 ;
      RECT 25.405 2.715 25.74 2.87 ;
      RECT 25.405 2.662 25.69 2.87 ;
      RECT 23.235 2.59 23.43 3.375 ;
      RECT 23.315 1.205 23.43 3.375 ;
      RECT 23.17 3.115 23.23 3.375 ;
      RECT 24.54 2.635 24.8 2.895 ;
      RECT 23.225 2.59 23.43 2.87 ;
      RECT 24.535 2.645 24.8 2.83 ;
      RECT 24.25 2.62 24.26 2.77 ;
      RECT 23.485 1.205 23.565 1.55 ;
      RECT 23.22 1.205 23.43 1.55 ;
      RECT 24.525 2.645 24.535 2.829 ;
      RECT 24.515 2.644 24.525 2.826 ;
      RECT 24.506 2.643 24.515 2.824 ;
      RECT 24.42 2.639 24.506 2.814 ;
      RECT 24.346 2.631 24.42 2.796 ;
      RECT 24.26 2.624 24.346 2.779 ;
      RECT 24.2 2.62 24.25 2.769 ;
      RECT 24.165 2.619 24.2 2.766 ;
      RECT 24.11 2.619 24.165 2.768 ;
      RECT 24.075 2.619 24.11 2.772 ;
      RECT 23.989 2.618 24.075 2.779 ;
      RECT 23.903 2.617 23.989 2.789 ;
      RECT 23.817 2.616 23.903 2.8 ;
      RECT 23.731 2.616 23.817 2.81 ;
      RECT 23.645 2.615 23.731 2.82 ;
      RECT 23.61 2.615 23.645 2.86 ;
      RECT 23.605 2.615 23.61 2.903 ;
      RECT 23.58 2.615 23.605 2.92 ;
      RECT 23.505 2.615 23.58 2.935 ;
      RECT 23.485 2.59 23.505 2.948 ;
      RECT 23.48 1.205 23.485 2.958 ;
      RECT 23.455 1.205 23.48 3 ;
      RECT 23.43 1.205 23.455 3.078 ;
      RECT 23.23 2.997 23.235 3.375 ;
      RECT 22.565 2.949 22.58 3.405 ;
      RECT 22.56 3.021 22.666 3.403 ;
      RECT 22.58 2.115 22.715 3.401 ;
      RECT 22.565 2.965 22.72 3.4 ;
      RECT 22.565 3.015 22.725 3.398 ;
      RECT 22.55 3.08 22.725 3.397 ;
      RECT 22.56 3.072 22.73 3.394 ;
      RECT 22.54 3.12 22.73 3.389 ;
      RECT 22.54 3.12 22.745 3.386 ;
      RECT 22.535 3.12 22.745 3.383 ;
      RECT 22.51 3.12 22.77 3.38 ;
      RECT 22.58 2.115 22.74 2.768 ;
      RECT 22.575 2.115 22.74 2.74 ;
      RECT 22.57 2.115 22.74 2.568 ;
      RECT 22.57 2.115 22.76 2.508 ;
      RECT 22.525 2.115 22.785 2.375 ;
      RECT 22.005 2.59 22.285 2.87 ;
      RECT 21.995 2.605 22.285 2.865 ;
      RECT 21.95 2.667 22.285 2.863 ;
      RECT 22.025 2.582 22.19 2.87 ;
      RECT 22.025 2.567 22.146 2.87 ;
      RECT 22.06 2.56 22.146 2.87 ;
      RECT 21.525 3.71 21.805 3.99 ;
      RECT 21.485 3.672 21.78 3.783 ;
      RECT 21.47 3.622 21.76 3.678 ;
      RECT 21.415 3.385 21.675 3.645 ;
      RECT 21.415 3.587 21.755 3.645 ;
      RECT 21.415 3.527 21.75 3.645 ;
      RECT 21.415 3.477 21.73 3.645 ;
      RECT 21.415 3.457 21.725 3.645 ;
      RECT 21.415 3.435 21.72 3.645 ;
      RECT 21.415 3.42 21.69 3.645 ;
      RECT 17.145 6.225 17.465 6.545 ;
      RECT 17.175 5.695 17.345 6.545 ;
      RECT 17.175 5.695 17.35 6.045 ;
      RECT 17.175 5.695 18.15 5.87 ;
      RECT 17.975 1.965 18.15 5.87 ;
      RECT 17.92 1.965 18.27 2.315 ;
      RECT 17.945 6.655 18.27 6.98 ;
      RECT 16.83 6.745 18.27 6.915 ;
      RECT 16.83 2.395 16.99 6.915 ;
      RECT 17.145 2.365 17.465 2.685 ;
      RECT 16.83 2.395 17.465 2.565 ;
      RECT 15.5 1.14 15.875 1.51 ;
      RECT 7.42 0.96 7.795 1.33 ;
      RECT 5.985 0.96 6.36 1.33 ;
      RECT 5.985 1.08 15.805 1.25 ;
      RECT 10.105 4.36 15.785 4.53 ;
      RECT 15.615 3.425 15.785 4.53 ;
      RECT 9.915 3.6 9.94 4.53 ;
      RECT 10.17 3.71 10.2 3.99 ;
      RECT 9.875 3.6 9.94 3.86 ;
      RECT 15.525 3.43 15.875 3.78 ;
      RECT 9.705 2.225 9.74 2.485 ;
      RECT 9.48 2.225 9.54 2.485 ;
      RECT 10.16 3.69 10.17 3.99 ;
      RECT 10.155 3.65 10.16 3.99 ;
      RECT 10.14 3.605 10.155 3.99 ;
      RECT 10.135 3.57 10.14 3.99 ;
      RECT 10.13 3.55 10.135 3.99 ;
      RECT 10.105 3.487 10.13 3.99 ;
      RECT 10.1 3.425 10.105 4.53 ;
      RECT 10.08 3.375 10.1 4.53 ;
      RECT 10.07 3.305 10.08 4.53 ;
      RECT 10.025 3.245 10.07 4.53 ;
      RECT 9.94 3.206 10.025 4.53 ;
      RECT 9.935 3.197 9.94 3.57 ;
      RECT 9.925 3.196 9.935 3.553 ;
      RECT 9.9 3.177 9.925 3.523 ;
      RECT 9.895 3.152 9.9 3.502 ;
      RECT 9.885 3.13 9.895 3.493 ;
      RECT 9.88 3.101 9.885 3.483 ;
      RECT 9.84 3.027 9.88 3.455 ;
      RECT 9.82 2.928 9.84 3.42 ;
      RECT 9.805 2.864 9.82 3.403 ;
      RECT 9.775 2.788 9.805 3.375 ;
      RECT 9.755 2.703 9.775 3.348 ;
      RECT 9.715 2.599 9.755 3.255 ;
      RECT 9.71 2.52 9.715 3.163 ;
      RECT 9.705 2.503 9.71 3.14 ;
      RECT 9.7 2.225 9.705 3.12 ;
      RECT 9.67 2.225 9.7 3.058 ;
      RECT 9.665 2.225 9.67 2.99 ;
      RECT 9.655 2.225 9.665 2.955 ;
      RECT 9.645 2.225 9.655 2.92 ;
      RECT 9.58 2.225 9.645 2.775 ;
      RECT 9.575 2.225 9.58 2.645 ;
      RECT 9.545 2.225 9.575 2.578 ;
      RECT 9.54 2.225 9.545 2.503 ;
      RECT 13.875 2.16 14.135 2.42 ;
      RECT 13.87 2.16 14.135 2.368 ;
      RECT 13.865 2.16 14.135 2.338 ;
      RECT 13.84 2.03 14.12 2.31 ;
      RECT 1.7 6.995 1.99 7.345 ;
      RECT 1.7 7.055 3.01 7.225 ;
      RECT 2.84 6.685 3.01 7.225 ;
      RECT 13.34 6.605 13.69 6.955 ;
      RECT 2.84 6.685 13.69 6.855 ;
      RECT 12.88 3.71 13.16 3.99 ;
      RECT 12.92 3.665 13.185 3.925 ;
      RECT 12.91 3.7 13.185 3.925 ;
      RECT 12.915 3.685 13.16 3.99 ;
      RECT 12.92 3.662 13.13 3.99 ;
      RECT 12.92 3.66 13.115 3.99 ;
      RECT 12.96 3.65 13.115 3.99 ;
      RECT 12.93 3.655 13.115 3.99 ;
      RECT 12.96 3.647 13.06 3.99 ;
      RECT 12.985 3.64 13.06 3.99 ;
      RECT 12.965 3.642 13.06 3.99 ;
      RECT 12.295 3.155 12.555 3.415 ;
      RECT 12.345 3.147 12.535 3.415 ;
      RECT 12.35 3.067 12.535 3.415 ;
      RECT 12.47 2.455 12.535 3.415 ;
      RECT 12.375 2.852 12.535 3.415 ;
      RECT 12.45 2.54 12.535 3.415 ;
      RECT 12.485 2.165 12.621 2.893 ;
      RECT 12.43 2.662 12.621 2.893 ;
      RECT 12.445 2.602 12.535 3.415 ;
      RECT 12.485 2.165 12.645 2.558 ;
      RECT 12.485 2.165 12.655 2.455 ;
      RECT 12.475 2.165 12.735 2.425 ;
      RECT 11.88 3.71 12.16 3.99 ;
      RECT 11.9 3.67 12.16 3.99 ;
      RECT 11.54 3.625 11.645 3.885 ;
      RECT 11.395 2.115 11.485 2.375 ;
      RECT 11.935 3.18 11.94 3.22 ;
      RECT 11.93 3.17 11.935 3.305 ;
      RECT 11.925 3.16 11.93 3.398 ;
      RECT 11.915 3.14 11.925 3.454 ;
      RECT 11.835 3.068 11.915 3.534 ;
      RECT 11.87 3.712 11.88 3.937 ;
      RECT 11.865 3.709 11.87 3.932 ;
      RECT 11.85 3.706 11.865 3.925 ;
      RECT 11.815 3.7 11.85 3.907 ;
      RECT 11.83 3.003 11.835 3.608 ;
      RECT 11.81 2.954 11.83 3.623 ;
      RECT 11.8 3.687 11.815 3.89 ;
      RECT 11.805 2.896 11.81 3.638 ;
      RECT 11.8 2.874 11.805 3.648 ;
      RECT 11.765 2.784 11.8 3.885 ;
      RECT 11.75 2.662 11.765 3.885 ;
      RECT 11.745 2.615 11.75 3.885 ;
      RECT 11.72 2.54 11.745 3.885 ;
      RECT 11.705 2.455 11.72 3.885 ;
      RECT 11.7 2.402 11.705 3.885 ;
      RECT 11.695 2.382 11.7 3.885 ;
      RECT 11.69 2.357 11.695 3.119 ;
      RECT 11.675 3.317 11.695 3.885 ;
      RECT 11.685 2.335 11.69 3.096 ;
      RECT 11.675 2.287 11.685 3.061 ;
      RECT 11.67 2.25 11.675 3.027 ;
      RECT 11.67 3.397 11.675 3.885 ;
      RECT 11.655 2.227 11.67 2.982 ;
      RECT 11.65 3.495 11.67 3.885 ;
      RECT 11.6 2.115 11.655 2.824 ;
      RECT 11.645 3.617 11.65 3.885 ;
      RECT 11.585 2.115 11.6 2.663 ;
      RECT 11.58 2.115 11.585 2.615 ;
      RECT 11.575 2.115 11.58 2.603 ;
      RECT 11.53 2.115 11.575 2.54 ;
      RECT 11.505 2.115 11.53 2.458 ;
      RECT 11.49 2.115 11.505 2.41 ;
      RECT 11.485 2.115 11.49 2.38 ;
      RECT 10.81 3.565 10.855 3.825 ;
      RECT 10.715 2.1 10.86 2.36 ;
      RECT 11.22 2.722 11.23 2.813 ;
      RECT 11.205 2.66 11.22 2.869 ;
      RECT 11.2 2.607 11.205 2.915 ;
      RECT 11.15 2.554 11.2 3.041 ;
      RECT 11.145 2.509 11.15 3.188 ;
      RECT 11.135 2.497 11.145 3.23 ;
      RECT 11.1 2.461 11.135 3.335 ;
      RECT 11.095 2.429 11.1 3.441 ;
      RECT 11.08 2.411 11.095 3.486 ;
      RECT 11.075 2.394 11.08 2.72 ;
      RECT 11.07 2.775 11.08 3.543 ;
      RECT 11.065 2.38 11.075 2.693 ;
      RECT 11.06 2.83 11.07 3.825 ;
      RECT 11.055 2.366 11.065 2.678 ;
      RECT 11.055 2.88 11.06 3.825 ;
      RECT 11.04 2.343 11.055 2.658 ;
      RECT 11.02 3.002 11.055 3.825 ;
      RECT 11.035 2.325 11.04 2.64 ;
      RECT 11.03 2.317 11.035 2.63 ;
      RECT 11 2.285 11.03 2.594 ;
      RECT 11.01 3.13 11.02 3.825 ;
      RECT 11.005 3.157 11.01 3.825 ;
      RECT 11 3.207 11.005 3.825 ;
      RECT 10.99 2.251 11 2.559 ;
      RECT 10.95 3.275 11 3.825 ;
      RECT 10.975 2.228 10.99 2.535 ;
      RECT 10.95 2.1 10.975 2.498 ;
      RECT 10.945 2.1 10.95 2.47 ;
      RECT 10.915 3.375 10.95 3.825 ;
      RECT 10.94 2.1 10.945 2.463 ;
      RECT 10.935 2.1 10.94 2.453 ;
      RECT 10.92 2.1 10.935 2.438 ;
      RECT 10.905 2.1 10.92 2.41 ;
      RECT 10.87 3.48 10.915 3.825 ;
      RECT 10.89 2.1 10.905 2.383 ;
      RECT 10.86 2.1 10.89 2.368 ;
      RECT 10.855 3.552 10.87 3.825 ;
      RECT 10.78 2.635 10.82 2.895 ;
      RECT 10.555 2.582 10.56 2.84 ;
      RECT 6.51 2.06 6.77 2.32 ;
      RECT 6.51 2.085 6.785 2.3 ;
      RECT 8.9 1.91 8.905 2.055 ;
      RECT 10.77 2.63 10.78 2.895 ;
      RECT 10.75 2.622 10.77 2.895 ;
      RECT 10.732 2.618 10.75 2.895 ;
      RECT 10.646 2.607 10.732 2.895 ;
      RECT 10.56 2.59 10.646 2.895 ;
      RECT 10.505 2.577 10.555 2.825 ;
      RECT 10.471 2.569 10.505 2.8 ;
      RECT 10.385 2.558 10.471 2.765 ;
      RECT 10.35 2.535 10.385 2.73 ;
      RECT 10.34 2.497 10.35 2.716 ;
      RECT 10.335 2.47 10.34 2.712 ;
      RECT 10.33 2.457 10.335 2.709 ;
      RECT 10.32 2.437 10.33 2.705 ;
      RECT 10.315 2.412 10.32 2.701 ;
      RECT 10.29 2.367 10.315 2.695 ;
      RECT 10.28 2.308 10.29 2.687 ;
      RECT 10.27 2.276 10.28 2.678 ;
      RECT 10.25 2.228 10.27 2.658 ;
      RECT 10.245 2.188 10.25 2.628 ;
      RECT 10.23 2.162 10.245 2.602 ;
      RECT 10.225 2.14 10.23 2.578 ;
      RECT 10.21 2.112 10.225 2.554 ;
      RECT 10.195 2.085 10.21 2.518 ;
      RECT 10.18 2.062 10.195 2.48 ;
      RECT 10.175 2.052 10.18 2.455 ;
      RECT 10.165 2.045 10.175 2.438 ;
      RECT 10.15 2.032 10.165 2.408 ;
      RECT 10.145 2.022 10.15 2.383 ;
      RECT 10.14 2.017 10.145 2.37 ;
      RECT 10.13 2.01 10.14 2.35 ;
      RECT 10.125 2.003 10.13 2.335 ;
      RECT 10.1 1.996 10.125 2.293 ;
      RECT 10.085 1.986 10.1 2.243 ;
      RECT 10.075 1.981 10.085 2.213 ;
      RECT 10.065 1.977 10.075 2.188 ;
      RECT 10.05 1.974 10.065 2.178 ;
      RECT 10 1.971 10.05 2.163 ;
      RECT 9.98 1.969 10 2.148 ;
      RECT 9.931 1.967 9.98 2.143 ;
      RECT 9.845 1.963 9.931 2.138 ;
      RECT 9.806 1.96 9.845 2.134 ;
      RECT 9.72 1.956 9.806 2.129 ;
      RECT 9.67 1.953 9.72 2.123 ;
      RECT 9.621 1.95 9.67 2.118 ;
      RECT 9.535 1.947 9.621 2.113 ;
      RECT 9.531 1.945 9.535 2.11 ;
      RECT 9.445 1.942 9.531 2.105 ;
      RECT 9.396 1.938 9.445 2.098 ;
      RECT 9.31 1.935 9.396 2.093 ;
      RECT 9.286 1.932 9.31 2.089 ;
      RECT 9.2 1.93 9.286 2.084 ;
      RECT 9.135 1.926 9.2 2.077 ;
      RECT 9.132 1.925 9.135 2.074 ;
      RECT 9.046 1.922 9.132 2.071 ;
      RECT 8.96 1.916 9.046 2.064 ;
      RECT 8.93 1.912 8.96 2.06 ;
      RECT 8.905 1.91 8.93 2.058 ;
      RECT 8.85 1.907 8.9 2.055 ;
      RECT 8.77 1.906 8.85 2.055 ;
      RECT 8.715 1.908 8.77 2.058 ;
      RECT 8.7 1.909 8.715 2.062 ;
      RECT 8.645 1.917 8.7 2.072 ;
      RECT 8.615 1.925 8.645 2.085 ;
      RECT 8.596 1.926 8.615 2.091 ;
      RECT 8.51 1.929 8.596 2.096 ;
      RECT 8.44 1.934 8.51 2.105 ;
      RECT 8.421 1.937 8.44 2.111 ;
      RECT 8.335 1.941 8.421 2.116 ;
      RECT 8.295 1.945 8.335 2.123 ;
      RECT 8.286 1.947 8.295 2.126 ;
      RECT 8.2 1.951 8.286 2.131 ;
      RECT 8.197 1.954 8.2 2.135 ;
      RECT 8.111 1.957 8.197 2.139 ;
      RECT 8.025 1.963 8.111 2.147 ;
      RECT 8.001 1.967 8.025 2.151 ;
      RECT 7.915 1.971 8.001 2.156 ;
      RECT 7.87 1.976 7.915 2.163 ;
      RECT 7.79 1.981 7.87 2.17 ;
      RECT 7.71 1.987 7.79 2.185 ;
      RECT 7.685 1.991 7.71 2.198 ;
      RECT 7.62 1.994 7.685 2.21 ;
      RECT 7.565 1.999 7.62 2.225 ;
      RECT 7.535 2.002 7.565 2.243 ;
      RECT 7.525 2.004 7.535 2.256 ;
      RECT 7.465 2.019 7.525 2.266 ;
      RECT 7.45 2.036 7.465 2.275 ;
      RECT 7.445 2.045 7.45 2.275 ;
      RECT 7.435 2.055 7.445 2.275 ;
      RECT 7.425 2.072 7.435 2.275 ;
      RECT 7.405 2.082 7.425 2.276 ;
      RECT 7.36 2.092 7.405 2.277 ;
      RECT 7.325 2.101 7.36 2.279 ;
      RECT 7.26 2.106 7.325 2.281 ;
      RECT 7.18 2.107 7.26 2.284 ;
      RECT 7.176 2.105 7.18 2.285 ;
      RECT 7.09 2.102 7.176 2.287 ;
      RECT 7.043 2.099 7.09 2.289 ;
      RECT 6.957 2.095 7.043 2.292 ;
      RECT 6.871 2.091 6.957 2.295 ;
      RECT 6.785 2.087 6.871 2.299 ;
      RECT 8.72 3.15 9 3.43 ;
      RECT 8.76 3.13 9.02 3.39 ;
      RECT 8.75 3.14 9.02 3.39 ;
      RECT 8.76 3.067 8.975 3.43 ;
      RECT 8.815 2.99 8.97 3.43 ;
      RECT 8.82 2.775 8.97 3.43 ;
      RECT 8.81 2.577 8.96 2.828 ;
      RECT 8.8 2.577 8.96 2.695 ;
      RECT 8.795 2.455 8.955 2.598 ;
      RECT 8.78 2.455 8.955 2.503 ;
      RECT 8.775 2.165 8.95 2.48 ;
      RECT 8.76 2.165 8.95 2.45 ;
      RECT 8.72 2.165 8.98 2.425 ;
      RECT 8.63 3.635 8.71 3.895 ;
      RECT 8.035 2.355 8.04 2.62 ;
      RECT 7.915 2.355 8.04 2.615 ;
      RECT 8.59 3.6 8.63 3.895 ;
      RECT 8.545 3.522 8.59 3.895 ;
      RECT 8.525 3.45 8.545 3.895 ;
      RECT 8.515 3.402 8.525 3.895 ;
      RECT 8.48 3.335 8.515 3.895 ;
      RECT 8.45 3.235 8.48 3.895 ;
      RECT 8.43 3.16 8.45 3.695 ;
      RECT 8.42 3.11 8.43 3.65 ;
      RECT 8.415 3.087 8.42 3.623 ;
      RECT 8.41 3.072 8.415 3.61 ;
      RECT 8.405 3.057 8.41 3.588 ;
      RECT 8.4 3.042 8.405 3.57 ;
      RECT 8.375 2.997 8.4 3.525 ;
      RECT 8.365 2.945 8.375 3.468 ;
      RECT 8.355 2.915 8.365 3.435 ;
      RECT 8.345 2.88 8.355 3.403 ;
      RECT 8.31 2.812 8.345 3.335 ;
      RECT 8.305 2.751 8.31 3.27 ;
      RECT 8.295 2.739 8.305 3.25 ;
      RECT 8.29 2.727 8.295 3.23 ;
      RECT 8.285 2.719 8.29 3.218 ;
      RECT 8.28 2.711 8.285 3.198 ;
      RECT 8.27 2.699 8.28 3.17 ;
      RECT 8.26 2.683 8.27 3.14 ;
      RECT 8.235 2.655 8.26 3.078 ;
      RECT 8.225 2.626 8.235 3.023 ;
      RECT 8.21 2.605 8.225 2.983 ;
      RECT 8.205 2.589 8.21 2.955 ;
      RECT 8.2 2.577 8.205 2.945 ;
      RECT 8.195 2.572 8.2 2.918 ;
      RECT 8.19 2.565 8.195 2.905 ;
      RECT 8.175 2.548 8.19 2.878 ;
      RECT 8.165 2.355 8.175 2.838 ;
      RECT 8.155 2.355 8.165 2.805 ;
      RECT 8.145 2.355 8.155 2.78 ;
      RECT 8.075 2.355 8.145 2.715 ;
      RECT 8.065 2.355 8.075 2.663 ;
      RECT 8.05 2.355 8.065 2.645 ;
      RECT 8.04 2.355 8.05 2.63 ;
      RECT 7.87 3.225 8.13 3.485 ;
      RECT 6.405 3.26 6.41 3.467 ;
      RECT 6.04 3.15 6.115 3.465 ;
      RECT 5.855 3.205 6.01 3.465 ;
      RECT 6.04 3.15 6.145 3.43 ;
      RECT 7.855 3.322 7.87 3.483 ;
      RECT 7.83 3.33 7.855 3.488 ;
      RECT 7.805 3.337 7.83 3.493 ;
      RECT 7.742 3.348 7.805 3.502 ;
      RECT 7.656 3.367 7.742 3.519 ;
      RECT 7.57 3.389 7.656 3.538 ;
      RECT 7.555 3.402 7.57 3.549 ;
      RECT 7.515 3.41 7.555 3.556 ;
      RECT 7.495 3.415 7.515 3.563 ;
      RECT 7.457 3.416 7.495 3.566 ;
      RECT 7.371 3.419 7.457 3.567 ;
      RECT 7.285 3.423 7.371 3.568 ;
      RECT 7.236 3.425 7.285 3.57 ;
      RECT 7.15 3.425 7.236 3.572 ;
      RECT 7.11 3.42 7.15 3.574 ;
      RECT 7.1 3.414 7.11 3.575 ;
      RECT 7.06 3.409 7.1 3.572 ;
      RECT 7.05 3.402 7.06 3.568 ;
      RECT 7.035 3.398 7.05 3.566 ;
      RECT 7.018 3.394 7.035 3.564 ;
      RECT 6.932 3.384 7.018 3.556 ;
      RECT 6.846 3.366 6.932 3.542 ;
      RECT 6.76 3.349 6.846 3.528 ;
      RECT 6.735 3.337 6.76 3.519 ;
      RECT 6.665 3.327 6.735 3.512 ;
      RECT 6.62 3.315 6.665 3.503 ;
      RECT 6.56 3.302 6.62 3.495 ;
      RECT 6.555 3.294 6.56 3.49 ;
      RECT 6.52 3.289 6.555 3.488 ;
      RECT 6.465 3.28 6.52 3.481 ;
      RECT 6.425 3.269 6.465 3.473 ;
      RECT 6.41 3.262 6.425 3.469 ;
      RECT 6.39 3.255 6.405 3.466 ;
      RECT 6.375 3.245 6.39 3.464 ;
      RECT 6.36 3.232 6.375 3.461 ;
      RECT 6.335 3.215 6.36 3.457 ;
      RECT 6.32 3.197 6.335 3.454 ;
      RECT 6.295 3.15 6.32 3.452 ;
      RECT 6.271 3.15 6.295 3.449 ;
      RECT 6.185 3.15 6.271 3.441 ;
      RECT 6.145 3.15 6.185 3.433 ;
      RECT 6.01 3.197 6.04 3.465 ;
      RECT 7.69 2.78 7.95 3.04 ;
      RECT 7.65 2.78 7.95 2.918 ;
      RECT 7.615 2.78 7.95 2.903 ;
      RECT 7.56 2.78 7.95 2.883 ;
      RECT 7.48 2.59 7.76 2.87 ;
      RECT 7.48 2.772 7.83 2.87 ;
      RECT 7.48 2.715 7.815 2.87 ;
      RECT 7.48 2.662 7.765 2.87 ;
      RECT 5.31 2.59 5.505 3.375 ;
      RECT 5.39 1.205 5.505 3.375 ;
      RECT 5.245 3.115 5.305 3.375 ;
      RECT 6.615 2.635 6.875 2.895 ;
      RECT 5.3 2.59 5.505 2.87 ;
      RECT 6.61 2.645 6.875 2.83 ;
      RECT 6.325 2.62 6.335 2.77 ;
      RECT 5.56 1.205 5.64 1.55 ;
      RECT 5.295 1.205 5.505 1.55 ;
      RECT 6.6 2.645 6.61 2.829 ;
      RECT 6.59 2.644 6.6 2.826 ;
      RECT 6.581 2.643 6.59 2.824 ;
      RECT 6.495 2.639 6.581 2.814 ;
      RECT 6.421 2.631 6.495 2.796 ;
      RECT 6.335 2.624 6.421 2.779 ;
      RECT 6.275 2.62 6.325 2.769 ;
      RECT 6.24 2.619 6.275 2.766 ;
      RECT 6.185 2.619 6.24 2.768 ;
      RECT 6.15 2.619 6.185 2.772 ;
      RECT 6.064 2.618 6.15 2.779 ;
      RECT 5.978 2.617 6.064 2.789 ;
      RECT 5.892 2.616 5.978 2.8 ;
      RECT 5.806 2.616 5.892 2.81 ;
      RECT 5.72 2.615 5.806 2.82 ;
      RECT 5.685 2.615 5.72 2.86 ;
      RECT 5.68 2.615 5.685 2.903 ;
      RECT 5.655 2.615 5.68 2.92 ;
      RECT 5.58 2.615 5.655 2.935 ;
      RECT 5.56 2.59 5.58 2.948 ;
      RECT 5.555 1.205 5.56 2.958 ;
      RECT 5.53 1.205 5.555 3 ;
      RECT 5.505 1.205 5.53 3.078 ;
      RECT 5.305 2.997 5.31 3.375 ;
      RECT 4.64 2.949 4.655 3.405 ;
      RECT 4.635 3.021 4.741 3.403 ;
      RECT 4.655 2.115 4.79 3.401 ;
      RECT 4.64 2.965 4.795 3.4 ;
      RECT 4.64 3.015 4.8 3.398 ;
      RECT 4.625 3.08 4.8 3.397 ;
      RECT 4.635 3.072 4.805 3.394 ;
      RECT 4.615 3.12 4.805 3.389 ;
      RECT 4.615 3.12 4.82 3.386 ;
      RECT 4.61 3.12 4.82 3.383 ;
      RECT 4.585 3.12 4.845 3.38 ;
      RECT 4.655 2.115 4.815 2.768 ;
      RECT 4.65 2.115 4.815 2.74 ;
      RECT 4.645 2.115 4.815 2.568 ;
      RECT 4.645 2.115 4.835 2.508 ;
      RECT 4.6 2.115 4.86 2.375 ;
      RECT 4.08 2.59 4.36 2.87 ;
      RECT 4.07 2.605 4.36 2.865 ;
      RECT 4.025 2.667 4.36 2.863 ;
      RECT 4.1 2.582 4.265 2.87 ;
      RECT 4.1 2.567 4.221 2.87 ;
      RECT 4.135 2.56 4.221 2.87 ;
      RECT 3.6 3.71 3.88 3.99 ;
      RECT 3.56 3.672 3.855 3.783 ;
      RECT 3.545 3.622 3.835 3.678 ;
      RECT 3.49 3.385 3.75 3.645 ;
      RECT 3.49 3.587 3.83 3.645 ;
      RECT 3.49 3.527 3.825 3.645 ;
      RECT 3.49 3.477 3.805 3.645 ;
      RECT 3.49 3.457 3.8 3.645 ;
      RECT 3.49 3.435 3.795 3.645 ;
      RECT 3.49 3.42 3.765 3.645 ;
      RECT 84.38 7.055 84.755 7.425 ;
      RECT 75.715 0.93 76.09 1.3 ;
      RECT 66.455 7.055 66.83 7.425 ;
      RECT 57.79 0.93 58.165 1.3 ;
      RECT 48.53 7.055 48.905 7.425 ;
      RECT 39.865 0.93 40.24 1.3 ;
      RECT 30.605 7.055 30.98 7.425 ;
      RECT 21.94 0.93 22.315 1.3 ;
      RECT 12.68 7.055 13.055 7.425 ;
      RECT 4.015 0.93 4.39 1.3 ;
    LAYER via1 ;
      RECT 92.1 7.375 92.25 7.525 ;
      RECT 89.735 6.74 89.885 6.89 ;
      RECT 89.72 2.065 89.87 2.215 ;
      RECT 88.93 2.45 89.08 2.6 ;
      RECT 88.93 6.325 89.08 6.475 ;
      RECT 87.325 3.53 87.475 3.68 ;
      RECT 87.315 1.25 87.465 1.4 ;
      RECT 85.63 2.215 85.78 2.365 ;
      RECT 85.4 6.71 85.55 6.86 ;
      RECT 84.68 3.72 84.83 3.87 ;
      RECT 84.495 7.165 84.645 7.315 ;
      RECT 84.23 2.22 84.38 2.37 ;
      RECT 84.05 3.21 84.2 3.36 ;
      RECT 83.655 3.725 83.805 3.875 ;
      RECT 83.295 3.68 83.445 3.83 ;
      RECT 83.15 2.17 83.3 2.32 ;
      RECT 82.565 3.62 82.715 3.77 ;
      RECT 82.47 2.155 82.62 2.305 ;
      RECT 82.315 2.69 82.465 2.84 ;
      RECT 81.63 3.655 81.78 3.805 ;
      RECT 81.235 2.28 81.385 2.43 ;
      RECT 80.515 3.185 80.665 3.335 ;
      RECT 80.475 2.22 80.625 2.37 ;
      RECT 80.205 3.69 80.355 3.84 ;
      RECT 79.67 2.41 79.82 2.56 ;
      RECT 79.625 3.28 79.775 3.43 ;
      RECT 79.445 2.835 79.595 2.985 ;
      RECT 78.37 2.69 78.52 2.84 ;
      RECT 78.265 2.115 78.415 2.265 ;
      RECT 77.61 3.26 77.76 3.41 ;
      RECT 77.09 1.3 77.24 1.45 ;
      RECT 77 3.17 77.15 3.32 ;
      RECT 76.355 2.17 76.505 2.32 ;
      RECT 76.34 3.175 76.49 3.325 ;
      RECT 75.825 2.66 75.975 2.81 ;
      RECT 75.245 3.44 75.395 3.59 ;
      RECT 74.155 6.755 74.305 6.905 ;
      RECT 71.81 6.74 71.96 6.89 ;
      RECT 71.795 2.065 71.945 2.215 ;
      RECT 71.005 2.45 71.155 2.6 ;
      RECT 71.005 6.325 71.155 6.475 ;
      RECT 69.4 3.53 69.55 3.68 ;
      RECT 69.39 1.25 69.54 1.4 ;
      RECT 67.705 2.215 67.855 2.365 ;
      RECT 67.195 6.71 67.345 6.86 ;
      RECT 66.755 3.72 66.905 3.87 ;
      RECT 66.57 7.165 66.72 7.315 ;
      RECT 66.305 2.22 66.455 2.37 ;
      RECT 66.125 3.21 66.275 3.36 ;
      RECT 65.73 3.725 65.88 3.875 ;
      RECT 65.37 3.68 65.52 3.83 ;
      RECT 65.225 2.17 65.375 2.32 ;
      RECT 64.64 3.62 64.79 3.77 ;
      RECT 64.545 2.155 64.695 2.305 ;
      RECT 64.39 2.69 64.54 2.84 ;
      RECT 63.705 3.655 63.855 3.805 ;
      RECT 63.31 2.28 63.46 2.43 ;
      RECT 62.59 3.185 62.74 3.335 ;
      RECT 62.55 2.22 62.7 2.37 ;
      RECT 62.28 3.69 62.43 3.84 ;
      RECT 61.745 2.41 61.895 2.56 ;
      RECT 61.7 3.28 61.85 3.43 ;
      RECT 61.52 2.835 61.67 2.985 ;
      RECT 60.445 2.69 60.595 2.84 ;
      RECT 60.34 2.115 60.49 2.265 ;
      RECT 59.685 3.26 59.835 3.41 ;
      RECT 59.165 1.3 59.315 1.45 ;
      RECT 59.075 3.17 59.225 3.32 ;
      RECT 58.43 2.17 58.58 2.32 ;
      RECT 58.415 3.175 58.565 3.325 ;
      RECT 57.9 2.66 58.05 2.81 ;
      RECT 57.32 3.44 57.47 3.59 ;
      RECT 56.23 6.755 56.38 6.905 ;
      RECT 53.885 6.74 54.035 6.89 ;
      RECT 53.87 2.065 54.02 2.215 ;
      RECT 53.08 2.45 53.23 2.6 ;
      RECT 53.08 6.325 53.23 6.475 ;
      RECT 51.475 3.53 51.625 3.68 ;
      RECT 51.465 1.25 51.615 1.4 ;
      RECT 49.78 2.215 49.93 2.365 ;
      RECT 49.325 6.715 49.475 6.865 ;
      RECT 48.83 3.72 48.98 3.87 ;
      RECT 48.645 7.165 48.795 7.315 ;
      RECT 48.38 2.22 48.53 2.37 ;
      RECT 48.2 3.21 48.35 3.36 ;
      RECT 47.805 3.725 47.955 3.875 ;
      RECT 47.445 3.68 47.595 3.83 ;
      RECT 47.3 2.17 47.45 2.32 ;
      RECT 46.715 3.62 46.865 3.77 ;
      RECT 46.62 2.155 46.77 2.305 ;
      RECT 46.465 2.69 46.615 2.84 ;
      RECT 45.78 3.655 45.93 3.805 ;
      RECT 45.385 2.28 45.535 2.43 ;
      RECT 44.665 3.185 44.815 3.335 ;
      RECT 44.625 2.22 44.775 2.37 ;
      RECT 44.355 3.69 44.505 3.84 ;
      RECT 43.82 2.41 43.97 2.56 ;
      RECT 43.775 3.28 43.925 3.43 ;
      RECT 43.595 2.835 43.745 2.985 ;
      RECT 42.52 2.69 42.67 2.84 ;
      RECT 42.415 2.115 42.565 2.265 ;
      RECT 41.76 3.26 41.91 3.41 ;
      RECT 41.24 1.3 41.39 1.45 ;
      RECT 41.15 3.17 41.3 3.32 ;
      RECT 40.505 2.17 40.655 2.32 ;
      RECT 40.49 3.175 40.64 3.325 ;
      RECT 39.975 2.66 40.125 2.81 ;
      RECT 39.395 3.44 39.545 3.59 ;
      RECT 38.35 6.76 38.5 6.91 ;
      RECT 35.96 6.74 36.11 6.89 ;
      RECT 35.945 2.065 36.095 2.215 ;
      RECT 35.155 2.45 35.305 2.6 ;
      RECT 35.155 6.325 35.305 6.475 ;
      RECT 33.55 3.53 33.7 3.68 ;
      RECT 33.54 1.25 33.69 1.4 ;
      RECT 31.855 2.215 32.005 2.365 ;
      RECT 31.395 6.71 31.545 6.86 ;
      RECT 30.905 3.72 31.055 3.87 ;
      RECT 30.72 7.165 30.87 7.315 ;
      RECT 30.455 2.22 30.605 2.37 ;
      RECT 30.275 3.21 30.425 3.36 ;
      RECT 29.88 3.725 30.03 3.875 ;
      RECT 29.52 3.68 29.67 3.83 ;
      RECT 29.375 2.17 29.525 2.32 ;
      RECT 28.79 3.62 28.94 3.77 ;
      RECT 28.695 2.155 28.845 2.305 ;
      RECT 28.54 2.69 28.69 2.84 ;
      RECT 27.855 3.655 28.005 3.805 ;
      RECT 27.46 2.28 27.61 2.43 ;
      RECT 26.74 3.185 26.89 3.335 ;
      RECT 26.7 2.22 26.85 2.37 ;
      RECT 26.43 3.69 26.58 3.84 ;
      RECT 25.895 2.41 26.045 2.56 ;
      RECT 25.85 3.28 26 3.43 ;
      RECT 25.67 2.835 25.82 2.985 ;
      RECT 24.595 2.69 24.745 2.84 ;
      RECT 24.49 2.115 24.64 2.265 ;
      RECT 23.835 3.26 23.985 3.41 ;
      RECT 23.315 1.3 23.465 1.45 ;
      RECT 23.225 3.17 23.375 3.32 ;
      RECT 22.58 2.17 22.73 2.32 ;
      RECT 22.565 3.175 22.715 3.325 ;
      RECT 22.05 2.66 22.2 2.81 ;
      RECT 21.47 3.44 21.62 3.59 ;
      RECT 20.425 6.755 20.575 6.905 ;
      RECT 18.035 6.74 18.185 6.89 ;
      RECT 18.02 2.065 18.17 2.215 ;
      RECT 17.23 2.45 17.38 2.6 ;
      RECT 17.23 6.325 17.38 6.475 ;
      RECT 15.625 3.53 15.775 3.68 ;
      RECT 15.615 1.25 15.765 1.4 ;
      RECT 13.93 2.215 14.08 2.365 ;
      RECT 13.44 6.705 13.59 6.855 ;
      RECT 12.98 3.72 13.13 3.87 ;
      RECT 12.795 7.165 12.945 7.315 ;
      RECT 12.53 2.22 12.68 2.37 ;
      RECT 12.35 3.21 12.5 3.36 ;
      RECT 11.955 3.725 12.105 3.875 ;
      RECT 11.595 3.68 11.745 3.83 ;
      RECT 11.45 2.17 11.6 2.32 ;
      RECT 10.865 3.62 11.015 3.77 ;
      RECT 10.77 2.155 10.92 2.305 ;
      RECT 10.615 2.69 10.765 2.84 ;
      RECT 9.93 3.655 10.08 3.805 ;
      RECT 9.535 2.28 9.685 2.43 ;
      RECT 8.815 3.185 8.965 3.335 ;
      RECT 8.775 2.22 8.925 2.37 ;
      RECT 8.505 3.69 8.655 3.84 ;
      RECT 7.97 2.41 8.12 2.56 ;
      RECT 7.925 3.28 8.075 3.43 ;
      RECT 7.745 2.835 7.895 2.985 ;
      RECT 6.67 2.69 6.82 2.84 ;
      RECT 6.565 2.115 6.715 2.265 ;
      RECT 5.91 3.26 6.06 3.41 ;
      RECT 5.39 1.3 5.54 1.45 ;
      RECT 5.3 3.17 5.45 3.32 ;
      RECT 4.655 2.17 4.805 2.32 ;
      RECT 4.64 3.175 4.79 3.325 ;
      RECT 4.125 2.66 4.275 2.81 ;
      RECT 3.545 3.44 3.695 3.59 ;
      RECT 1.77 7.095 1.92 7.245 ;
      RECT 1.395 6.355 1.545 6.505 ;
    LAYER met1 ;
      RECT 75.025 1.285 86.985 1.89 ;
      RECT 79.45 0 86.985 1.89 ;
      RECT 57.1 1.285 69.06 1.89 ;
      RECT 61.525 0 69.06 1.89 ;
      RECT 39.175 1.285 51.135 1.89 ;
      RECT 43.6 0 51.135 1.89 ;
      RECT 21.25 1.285 33.21 1.89 ;
      RECT 25.675 0 33.21 1.89 ;
      RECT 3.325 1.285 15.285 1.89 ;
      RECT 7.75 0 15.285 1.89 ;
      RECT 75.02 0 75.765 1.68 ;
      RECT 57.095 0 57.84 1.68 ;
      RECT 39.17 0 39.915 1.68 ;
      RECT 21.245 0 21.99 1.68 ;
      RECT 3.32 0 4.065 1.68 ;
      RECT 78.015 0 79.17 1.89 ;
      RECT 75.02 1.255 77.735 1.68 ;
      RECT 76.045 0 77.735 1.89 ;
      RECT 60.09 0 61.245 1.89 ;
      RECT 57.095 1.255 59.81 1.68 ;
      RECT 58.12 0 59.81 1.89 ;
      RECT 42.165 0 43.32 1.89 ;
      RECT 39.17 1.255 41.885 1.68 ;
      RECT 40.195 0 41.885 1.89 ;
      RECT 24.24 0 25.395 1.89 ;
      RECT 21.245 1.255 23.96 1.68 ;
      RECT 22.27 0 23.96 1.89 ;
      RECT 6.315 0 7.47 1.89 ;
      RECT 3.32 1.255 6.035 1.68 ;
      RECT 4.345 0 6.035 1.89 ;
      RECT 76.045 0 86.985 1.005 ;
      RECT 58.12 0 69.06 1.005 ;
      RECT 40.195 0 51.135 1.005 ;
      RECT 22.27 0 33.21 1.005 ;
      RECT 4.345 0 15.285 1.005 ;
      RECT 75.02 0 86.985 0.975 ;
      RECT 57.095 0 69.06 0.975 ;
      RECT 39.17 0 51.135 0.975 ;
      RECT 21.245 0 33.21 0.975 ;
      RECT 3.32 0 15.285 0.975 ;
      RECT 92.395 0 92.575 0.305 ;
      RECT 74.47 0 90.445 0.305 ;
      RECT 56.545 0 72.52 0.305 ;
      RECT 38.62 0 54.595 0.305 ;
      RECT 20.695 0 36.67 0.305 ;
      RECT 0 0 18.745 0.305 ;
      RECT 0 0 92.575 0.3 ;
      RECT 0 8.58 92.575 8.88 ;
      RECT 92.395 8.575 92.575 8.88 ;
      RECT 74.47 8.575 90.445 8.88 ;
      RECT 56.545 8.575 72.52 8.88 ;
      RECT 38.62 8.575 54.595 8.88 ;
      RECT 20.695 8.575 36.67 8.88 ;
      RECT 0 8.575 18.745 8.88 ;
      RECT 83.72 6.315 83.89 8.88 ;
      RECT 65.795 6.315 65.965 8.88 ;
      RECT 47.87 6.315 48.04 8.88 ;
      RECT 29.945 6.315 30.115 8.88 ;
      RECT 12.02 6.315 12.19 8.88 ;
      RECT 84.055 6.285 84.345 6.515 ;
      RECT 66.13 6.285 66.42 6.515 ;
      RECT 48.205 6.285 48.495 6.515 ;
      RECT 30.28 6.285 30.57 6.515 ;
      RECT 12.355 6.285 12.645 6.515 ;
      RECT 83.72 6.315 84.345 6.485 ;
      RECT 65.795 6.315 66.42 6.485 ;
      RECT 47.87 6.315 48.495 6.485 ;
      RECT 29.945 6.315 30.57 6.485 ;
      RECT 12.02 6.315 12.645 6.485 ;
      RECT 91.97 7.77 92.26 8 ;
      RECT 92.03 6.29 92.2 8 ;
      RECT 92 7.275 92.35 7.625 ;
      RECT 91.97 6.29 92.26 6.52 ;
      RECT 91.565 2.395 91.67 2.965 ;
      RECT 91.565 2.73 91.89 2.96 ;
      RECT 91.565 2.76 92.06 2.93 ;
      RECT 91.565 2.395 91.755 2.96 ;
      RECT 90.98 2.36 91.27 2.59 ;
      RECT 90.98 2.395 91.755 2.565 ;
      RECT 91.04 0.88 91.21 2.59 ;
      RECT 90.98 0.88 91.27 1.11 ;
      RECT 90.98 7.77 91.27 8 ;
      RECT 91.04 6.29 91.21 8 ;
      RECT 90.98 6.29 91.27 6.52 ;
      RECT 90.98 6.325 91.835 6.485 ;
      RECT 91.665 5.92 91.835 6.485 ;
      RECT 90.98 6.32 91.375 6.485 ;
      RECT 91.6 5.92 91.89 6.15 ;
      RECT 91.6 5.95 92.06 6.12 ;
      RECT 90.61 2.73 90.9 2.96 ;
      RECT 90.61 2.76 91.07 2.93 ;
      RECT 90.675 1.655 90.84 2.96 ;
      RECT 89.19 1.625 89.48 1.855 ;
      RECT 89.19 1.655 90.84 1.825 ;
      RECT 89.25 0.885 89.42 1.855 ;
      RECT 89.19 0.885 89.48 1.115 ;
      RECT 89.19 7.765 89.48 7.995 ;
      RECT 89.25 7.025 89.42 7.995 ;
      RECT 89.25 7.12 90.84 7.29 ;
      RECT 90.67 5.92 90.84 7.29 ;
      RECT 89.19 7.025 89.48 7.255 ;
      RECT 90.61 5.92 90.9 6.15 ;
      RECT 90.61 5.95 91.07 6.12 ;
      RECT 87.225 3.43 87.575 3.78 ;
      RECT 87.315 2.025 87.485 3.78 ;
      RECT 89.62 1.965 89.97 2.315 ;
      RECT 87.315 2.025 88.935 2.2 ;
      RECT 87.315 2.025 89.97 2.195 ;
      RECT 89.645 6.655 89.97 6.98 ;
      RECT 85.3 6.61 85.65 6.96 ;
      RECT 89.62 6.655 89.97 6.885 ;
      RECT 84.86 6.655 85.15 6.885 ;
      RECT 84.69 6.685 89.97 6.855 ;
      RECT 88.845 2.365 89.165 2.685 ;
      RECT 88.815 2.365 89.165 2.595 ;
      RECT 88.645 2.395 89.165 2.565 ;
      RECT 88.845 6.225 89.165 6.545 ;
      RECT 88.815 6.285 89.165 6.515 ;
      RECT 88.645 6.315 89.165 6.485 ;
      RECT 84.625 3.665 84.665 3.925 ;
      RECT 84.665 3.645 84.67 3.655 ;
      RECT 85.995 2.89 86.005 3.111 ;
      RECT 85.925 2.885 85.995 3.236 ;
      RECT 85.915 2.885 85.925 3.363 ;
      RECT 85.89 2.885 85.915 3.41 ;
      RECT 85.865 2.885 85.89 3.488 ;
      RECT 85.845 2.885 85.865 3.558 ;
      RECT 85.82 2.885 85.845 3.598 ;
      RECT 85.81 2.885 85.82 3.618 ;
      RECT 85.8 2.887 85.81 3.626 ;
      RECT 85.795 2.892 85.8 3.083 ;
      RECT 85.795 3.092 85.8 3.627 ;
      RECT 85.79 3.137 85.795 3.628 ;
      RECT 85.78 3.202 85.79 3.629 ;
      RECT 85.77 3.297 85.78 3.631 ;
      RECT 85.765 3.35 85.77 3.633 ;
      RECT 85.76 3.37 85.765 3.634 ;
      RECT 85.705 3.395 85.76 3.64 ;
      RECT 85.665 3.43 85.705 3.649 ;
      RECT 85.655 3.447 85.665 3.654 ;
      RECT 85.646 3.453 85.655 3.656 ;
      RECT 85.56 3.491 85.646 3.667 ;
      RECT 85.555 3.53 85.56 3.677 ;
      RECT 85.48 3.537 85.555 3.687 ;
      RECT 85.46 3.547 85.48 3.698 ;
      RECT 85.43 3.554 85.46 3.706 ;
      RECT 85.405 3.561 85.43 3.713 ;
      RECT 85.381 3.567 85.405 3.718 ;
      RECT 85.295 3.58 85.381 3.73 ;
      RECT 85.217 3.587 85.295 3.748 ;
      RECT 85.131 3.582 85.217 3.766 ;
      RECT 85.045 3.577 85.131 3.786 ;
      RECT 84.965 3.571 85.045 3.803 ;
      RECT 84.9 3.567 84.965 3.832 ;
      RECT 84.895 3.281 84.9 3.305 ;
      RECT 84.885 3.557 84.9 3.86 ;
      RECT 84.89 3.275 84.895 3.345 ;
      RECT 84.885 3.269 84.89 3.415 ;
      RECT 84.88 3.263 84.885 3.493 ;
      RECT 84.88 3.54 84.885 3.925 ;
      RECT 84.872 3.26 84.88 3.925 ;
      RECT 84.786 3.258 84.872 3.925 ;
      RECT 84.7 3.256 84.786 3.925 ;
      RECT 84.69 3.257 84.7 3.925 ;
      RECT 84.685 3.262 84.69 3.925 ;
      RECT 84.675 3.275 84.685 3.925 ;
      RECT 84.67 3.297 84.675 3.925 ;
      RECT 84.665 3.657 84.67 3.925 ;
      RECT 85.295 3.125 85.3 3.345 ;
      RECT 85.8 2.16 85.835 2.42 ;
      RECT 85.785 2.16 85.8 2.428 ;
      RECT 85.756 2.16 85.785 2.45 ;
      RECT 85.67 2.16 85.756 2.51 ;
      RECT 85.65 2.16 85.67 2.575 ;
      RECT 85.59 2.16 85.65 2.74 ;
      RECT 85.585 2.16 85.59 2.888 ;
      RECT 85.58 2.16 85.585 2.9 ;
      RECT 85.575 2.16 85.58 2.926 ;
      RECT 85.545 2.346 85.575 3.006 ;
      RECT 85.54 2.394 85.545 3.095 ;
      RECT 85.535 2.408 85.54 3.11 ;
      RECT 85.53 2.427 85.535 3.14 ;
      RECT 85.525 2.442 85.53 3.156 ;
      RECT 85.52 2.457 85.525 3.178 ;
      RECT 85.515 2.477 85.52 3.2 ;
      RECT 85.505 2.497 85.515 3.233 ;
      RECT 85.49 2.539 85.505 3.295 ;
      RECT 85.485 2.57 85.49 3.335 ;
      RECT 85.48 2.582 85.485 3.34 ;
      RECT 85.475 2.594 85.48 3.345 ;
      RECT 85.47 2.607 85.475 3.345 ;
      RECT 85.465 2.625 85.47 3.345 ;
      RECT 85.46 2.645 85.465 3.345 ;
      RECT 85.455 2.657 85.46 3.345 ;
      RECT 85.45 2.67 85.455 3.345 ;
      RECT 85.43 2.705 85.45 3.345 ;
      RECT 85.38 2.807 85.43 3.345 ;
      RECT 85.375 2.892 85.38 3.345 ;
      RECT 85.37 2.9 85.375 3.345 ;
      RECT 85.365 2.917 85.37 3.345 ;
      RECT 85.36 2.932 85.365 3.345 ;
      RECT 85.325 2.997 85.36 3.345 ;
      RECT 85.31 3.062 85.325 3.345 ;
      RECT 85.305 3.092 85.31 3.345 ;
      RECT 85.3 3.117 85.305 3.345 ;
      RECT 85.285 3.127 85.295 3.345 ;
      RECT 85.27 3.14 85.285 3.338 ;
      RECT 85.015 2.73 85.085 2.94 ;
      RECT 84.805 2.707 84.81 2.9 ;
      RECT 82.26 2.635 82.52 2.895 ;
      RECT 85.095 2.917 85.1 2.92 ;
      RECT 85.085 2.735 85.095 2.935 ;
      RECT 84.986 2.728 85.015 2.94 ;
      RECT 84.9 2.72 84.986 2.94 ;
      RECT 84.885 2.714 84.9 2.938 ;
      RECT 84.865 2.713 84.885 2.925 ;
      RECT 84.86 2.712 84.865 2.908 ;
      RECT 84.81 2.709 84.86 2.903 ;
      RECT 84.78 2.706 84.805 2.898 ;
      RECT 84.76 2.704 84.78 2.893 ;
      RECT 84.745 2.702 84.76 2.89 ;
      RECT 84.715 2.7 84.745 2.888 ;
      RECT 84.65 2.696 84.715 2.88 ;
      RECT 84.62 2.691 84.65 2.875 ;
      RECT 84.6 2.689 84.62 2.873 ;
      RECT 84.57 2.686 84.6 2.868 ;
      RECT 84.51 2.682 84.57 2.86 ;
      RECT 84.505 2.679 84.51 2.855 ;
      RECT 84.435 2.677 84.505 2.85 ;
      RECT 84.406 2.673 84.435 2.843 ;
      RECT 84.32 2.668 84.406 2.835 ;
      RECT 84.286 2.663 84.32 2.827 ;
      RECT 84.2 2.655 84.286 2.819 ;
      RECT 84.161 2.648 84.2 2.811 ;
      RECT 84.075 2.643 84.161 2.803 ;
      RECT 84.01 2.637 84.075 2.793 ;
      RECT 83.99 2.632 84.01 2.788 ;
      RECT 83.981 2.629 83.99 2.787 ;
      RECT 83.895 2.625 83.981 2.781 ;
      RECT 83.855 2.621 83.895 2.773 ;
      RECT 83.835 2.617 83.855 2.771 ;
      RECT 83.775 2.617 83.835 2.768 ;
      RECT 83.755 2.62 83.775 2.766 ;
      RECT 83.734 2.62 83.755 2.766 ;
      RECT 83.648 2.622 83.734 2.77 ;
      RECT 83.562 2.624 83.648 2.776 ;
      RECT 83.476 2.626 83.562 2.783 ;
      RECT 83.39 2.629 83.476 2.789 ;
      RECT 83.356 2.63 83.39 2.794 ;
      RECT 83.27 2.633 83.356 2.799 ;
      RECT 83.241 2.64 83.27 2.804 ;
      RECT 83.155 2.64 83.241 2.809 ;
      RECT 83.122 2.64 83.155 2.814 ;
      RECT 83.036 2.642 83.122 2.819 ;
      RECT 82.95 2.644 83.036 2.826 ;
      RECT 82.886 2.646 82.95 2.832 ;
      RECT 82.8 2.648 82.886 2.838 ;
      RECT 82.797 2.65 82.8 2.841 ;
      RECT 82.711 2.651 82.797 2.845 ;
      RECT 82.625 2.654 82.711 2.852 ;
      RECT 82.606 2.656 82.625 2.856 ;
      RECT 82.52 2.658 82.606 2.861 ;
      RECT 82.25 2.67 82.26 2.865 ;
      RECT 84.43 7.765 84.72 7.995 ;
      RECT 84.49 7.025 84.66 7.995 ;
      RECT 84.38 7.055 84.755 7.425 ;
      RECT 84.43 7.025 84.72 7.425 ;
      RECT 84.485 2.25 84.67 2.46 ;
      RECT 84.48 2.251 84.675 2.458 ;
      RECT 84.475 2.256 84.685 2.453 ;
      RECT 84.47 2.232 84.475 2.45 ;
      RECT 84.44 2.229 84.47 2.443 ;
      RECT 84.435 2.225 84.44 2.434 ;
      RECT 84.4 2.256 84.685 2.429 ;
      RECT 84.175 2.165 84.435 2.425 ;
      RECT 84.475 2.234 84.48 2.453 ;
      RECT 84.48 2.235 84.485 2.458 ;
      RECT 84.175 2.247 84.555 2.425 ;
      RECT 84.175 2.245 84.54 2.425 ;
      RECT 84.175 2.24 84.53 2.425 ;
      RECT 84.13 3.155 84.18 3.44 ;
      RECT 84.075 3.125 84.08 3.44 ;
      RECT 84.045 3.105 84.05 3.44 ;
      RECT 84.195 3.155 84.255 3.415 ;
      RECT 84.19 3.155 84.195 3.423 ;
      RECT 84.18 3.155 84.19 3.435 ;
      RECT 84.095 3.145 84.13 3.44 ;
      RECT 84.09 3.132 84.095 3.44 ;
      RECT 84.08 3.127 84.09 3.44 ;
      RECT 84.06 3.117 84.075 3.44 ;
      RECT 84.05 3.11 84.06 3.44 ;
      RECT 84.04 3.102 84.045 3.44 ;
      RECT 84.01 3.092 84.04 3.44 ;
      RECT 83.995 3.08 84.01 3.44 ;
      RECT 83.98 3.07 83.995 3.435 ;
      RECT 83.96 3.06 83.98 3.41 ;
      RECT 83.95 3.052 83.96 3.387 ;
      RECT 83.92 3.035 83.95 3.377 ;
      RECT 83.915 3.012 83.92 3.368 ;
      RECT 83.91 2.999 83.915 3.366 ;
      RECT 83.895 2.975 83.91 3.36 ;
      RECT 83.89 2.951 83.895 3.354 ;
      RECT 83.88 2.94 83.89 3.349 ;
      RECT 83.875 2.93 83.88 3.345 ;
      RECT 83.87 2.922 83.875 3.342 ;
      RECT 83.86 2.917 83.87 3.338 ;
      RECT 83.855 2.912 83.86 3.334 ;
      RECT 83.77 2.91 83.855 3.309 ;
      RECT 83.74 2.91 83.77 3.275 ;
      RECT 83.725 2.91 83.74 3.258 ;
      RECT 83.67 2.91 83.725 3.203 ;
      RECT 83.665 2.915 83.67 3.152 ;
      RECT 83.655 2.92 83.665 3.142 ;
      RECT 83.65 2.93 83.655 3.128 ;
      RECT 83.6 3.67 83.86 3.93 ;
      RECT 83.52 3.685 83.86 3.906 ;
      RECT 83.5 3.685 83.86 3.901 ;
      RECT 83.476 3.685 83.86 3.899 ;
      RECT 83.39 3.685 83.86 3.894 ;
      RECT 83.24 3.625 83.5 3.89 ;
      RECT 83.195 3.685 83.86 3.885 ;
      RECT 83.19 3.692 83.86 3.88 ;
      RECT 83.205 3.68 83.52 3.89 ;
      RECT 83.095 2.115 83.355 2.375 ;
      RECT 83.095 2.172 83.36 2.368 ;
      RECT 83.095 2.202 83.365 2.3 ;
      RECT 83.155 2.633 83.27 2.635 ;
      RECT 83.241 2.63 83.27 2.635 ;
      RECT 82.265 3.634 82.29 3.874 ;
      RECT 82.25 3.637 82.34 3.868 ;
      RECT 82.245 3.642 82.426 3.863 ;
      RECT 82.24 3.65 82.49 3.861 ;
      RECT 82.24 3.65 82.5 3.86 ;
      RECT 82.235 3.657 82.51 3.853 ;
      RECT 82.235 3.657 82.596 3.842 ;
      RECT 82.23 3.692 82.596 3.838 ;
      RECT 82.23 3.692 82.605 3.827 ;
      RECT 82.51 3.565 82.77 3.825 ;
      RECT 82.22 3.742 82.77 3.823 ;
      RECT 82.49 3.61 82.51 3.858 ;
      RECT 82.426 3.613 82.49 3.862 ;
      RECT 82.34 3.618 82.426 3.867 ;
      RECT 82.27 3.629 82.77 3.825 ;
      RECT 82.29 3.623 82.34 3.872 ;
      RECT 82.415 2.1 82.425 2.362 ;
      RECT 82.405 2.157 82.415 2.365 ;
      RECT 82.38 2.162 82.405 2.371 ;
      RECT 82.355 2.166 82.38 2.383 ;
      RECT 82.345 2.169 82.355 2.393 ;
      RECT 82.34 2.17 82.345 2.398 ;
      RECT 82.335 2.171 82.34 2.403 ;
      RECT 82.33 2.172 82.335 2.405 ;
      RECT 82.305 2.175 82.33 2.408 ;
      RECT 82.275 2.181 82.305 2.411 ;
      RECT 82.21 2.192 82.275 2.414 ;
      RECT 82.165 2.2 82.21 2.418 ;
      RECT 82.15 2.2 82.165 2.426 ;
      RECT 82.145 2.201 82.15 2.433 ;
      RECT 82.14 2.203 82.145 2.436 ;
      RECT 82.135 2.207 82.14 2.439 ;
      RECT 82.125 2.215 82.135 2.443 ;
      RECT 82.12 2.228 82.125 2.448 ;
      RECT 82.115 2.236 82.12 2.45 ;
      RECT 82.11 2.242 82.115 2.45 ;
      RECT 82.105 2.246 82.11 2.453 ;
      RECT 82.1 2.248 82.105 2.456 ;
      RECT 82.095 2.251 82.1 2.459 ;
      RECT 82.085 2.256 82.095 2.463 ;
      RECT 82.08 2.262 82.085 2.468 ;
      RECT 82.07 2.268 82.08 2.472 ;
      RECT 82.055 2.275 82.07 2.478 ;
      RECT 82.026 2.289 82.055 2.488 ;
      RECT 81.94 2.324 82.026 2.52 ;
      RECT 81.92 2.357 81.94 2.549 ;
      RECT 81.9 2.37 81.92 2.56 ;
      RECT 81.88 2.382 81.9 2.571 ;
      RECT 81.83 2.404 81.88 2.591 ;
      RECT 81.815 2.422 81.83 2.608 ;
      RECT 81.81 2.428 81.815 2.611 ;
      RECT 81.805 2.432 81.81 2.614 ;
      RECT 81.8 2.436 81.805 2.618 ;
      RECT 81.795 2.438 81.8 2.621 ;
      RECT 81.785 2.445 81.795 2.624 ;
      RECT 81.78 2.45 81.785 2.628 ;
      RECT 81.775 2.452 81.78 2.631 ;
      RECT 81.77 2.456 81.775 2.634 ;
      RECT 81.765 2.458 81.77 2.638 ;
      RECT 81.75 2.463 81.765 2.643 ;
      RECT 81.745 2.468 81.75 2.646 ;
      RECT 81.74 2.476 81.745 2.649 ;
      RECT 81.735 2.478 81.74 2.652 ;
      RECT 81.73 2.48 81.735 2.655 ;
      RECT 81.72 2.482 81.73 2.661 ;
      RECT 81.685 2.496 81.72 2.673 ;
      RECT 81.675 2.511 81.685 2.683 ;
      RECT 81.6 2.54 81.675 2.707 ;
      RECT 81.595 2.565 81.6 2.73 ;
      RECT 81.58 2.569 81.595 2.736 ;
      RECT 81.57 2.577 81.58 2.741 ;
      RECT 81.54 2.59 81.57 2.745 ;
      RECT 81.53 2.605 81.54 2.75 ;
      RECT 81.52 2.61 81.53 2.753 ;
      RECT 81.515 2.612 81.52 2.755 ;
      RECT 81.5 2.615 81.515 2.758 ;
      RECT 81.495 2.617 81.5 2.761 ;
      RECT 81.475 2.622 81.495 2.765 ;
      RECT 81.445 2.627 81.475 2.773 ;
      RECT 81.42 2.634 81.445 2.781 ;
      RECT 81.415 2.639 81.42 2.786 ;
      RECT 81.385 2.642 81.415 2.79 ;
      RECT 81.345 2.645 81.385 2.8 ;
      RECT 81.31 2.642 81.345 2.812 ;
      RECT 81.3 2.638 81.31 2.819 ;
      RECT 81.275 2.634 81.3 2.825 ;
      RECT 81.27 2.63 81.275 2.83 ;
      RECT 81.23 2.627 81.27 2.83 ;
      RECT 81.215 2.612 81.23 2.831 ;
      RECT 81.192 2.6 81.215 2.831 ;
      RECT 81.106 2.6 81.192 2.832 ;
      RECT 81.02 2.6 81.106 2.834 ;
      RECT 81 2.6 81.02 2.831 ;
      RECT 80.995 2.605 81 2.826 ;
      RECT 80.99 2.61 80.995 2.824 ;
      RECT 80.98 2.62 80.99 2.822 ;
      RECT 80.975 2.626 80.98 2.815 ;
      RECT 80.97 2.628 80.975 2.8 ;
      RECT 80.965 2.632 80.97 2.79 ;
      RECT 82.425 2.1 82.675 2.36 ;
      RECT 80.15 3.635 80.41 3.895 ;
      RECT 82.445 3.125 82.45 3.335 ;
      RECT 82.45 3.13 82.46 3.33 ;
      RECT 82.4 3.125 82.445 3.35 ;
      RECT 82.39 3.125 82.4 3.37 ;
      RECT 82.371 3.125 82.39 3.375 ;
      RECT 82.285 3.125 82.371 3.372 ;
      RECT 82.255 3.127 82.285 3.37 ;
      RECT 82.2 3.137 82.255 3.368 ;
      RECT 82.135 3.151 82.2 3.366 ;
      RECT 82.13 3.159 82.135 3.365 ;
      RECT 82.115 3.162 82.13 3.363 ;
      RECT 82.05 3.172 82.115 3.359 ;
      RECT 82.002 3.186 82.05 3.36 ;
      RECT 81.916 3.203 82.002 3.374 ;
      RECT 81.83 3.224 81.916 3.391 ;
      RECT 81.81 3.237 81.83 3.401 ;
      RECT 81.765 3.245 81.81 3.408 ;
      RECT 81.73 3.253 81.765 3.416 ;
      RECT 81.696 3.261 81.73 3.424 ;
      RECT 81.61 3.275 81.696 3.436 ;
      RECT 81.575 3.292 81.61 3.448 ;
      RECT 81.566 3.301 81.575 3.452 ;
      RECT 81.48 3.319 81.566 3.469 ;
      RECT 81.421 3.346 81.48 3.496 ;
      RECT 81.335 3.373 81.421 3.524 ;
      RECT 81.315 3.395 81.335 3.544 ;
      RECT 81.255 3.41 81.315 3.56 ;
      RECT 81.245 3.422 81.255 3.573 ;
      RECT 81.24 3.427 81.245 3.576 ;
      RECT 81.23 3.43 81.24 3.579 ;
      RECT 81.225 3.432 81.23 3.582 ;
      RECT 81.195 3.44 81.225 3.589 ;
      RECT 81.18 3.447 81.195 3.597 ;
      RECT 81.17 3.452 81.18 3.601 ;
      RECT 81.165 3.455 81.17 3.604 ;
      RECT 81.155 3.457 81.165 3.607 ;
      RECT 81.12 3.467 81.155 3.616 ;
      RECT 81.045 3.49 81.12 3.638 ;
      RECT 81.025 3.508 81.045 3.656 ;
      RECT 80.995 3.515 81.025 3.666 ;
      RECT 80.975 3.523 80.995 3.676 ;
      RECT 80.965 3.529 80.975 3.683 ;
      RECT 80.946 3.534 80.965 3.689 ;
      RECT 80.86 3.554 80.946 3.709 ;
      RECT 80.845 3.574 80.86 3.728 ;
      RECT 80.8 3.586 80.845 3.739 ;
      RECT 80.735 3.607 80.8 3.762 ;
      RECT 80.695 3.627 80.735 3.783 ;
      RECT 80.685 3.637 80.695 3.793 ;
      RECT 80.635 3.649 80.685 3.804 ;
      RECT 80.615 3.665 80.635 3.816 ;
      RECT 80.585 3.675 80.615 3.822 ;
      RECT 80.575 3.68 80.585 3.824 ;
      RECT 80.506 3.681 80.575 3.83 ;
      RECT 80.42 3.683 80.506 3.84 ;
      RECT 80.41 3.684 80.42 3.845 ;
      RECT 81.68 3.71 81.87 3.92 ;
      RECT 81.67 3.715 81.88 3.913 ;
      RECT 81.655 3.715 81.88 3.878 ;
      RECT 81.575 3.6 81.835 3.86 ;
      RECT 80.49 3.13 80.675 3.425 ;
      RECT 80.48 3.13 80.675 3.423 ;
      RECT 80.465 3.13 80.68 3.418 ;
      RECT 80.465 3.13 80.685 3.415 ;
      RECT 80.46 3.13 80.685 3.413 ;
      RECT 80.455 3.385 80.685 3.403 ;
      RECT 80.46 3.13 80.72 3.39 ;
      RECT 80.42 2.165 80.68 2.425 ;
      RECT 80.23 2.09 80.316 2.423 ;
      RECT 80.205 2.094 80.36 2.419 ;
      RECT 80.316 2.086 80.36 2.419 ;
      RECT 80.316 2.087 80.365 2.418 ;
      RECT 80.23 2.092 80.38 2.417 ;
      RECT 80.205 2.1 80.42 2.416 ;
      RECT 80.2 2.095 80.38 2.411 ;
      RECT 80.19 2.11 80.42 2.318 ;
      RECT 80.19 2.162 80.62 2.318 ;
      RECT 80.19 2.155 80.6 2.318 ;
      RECT 80.19 2.142 80.57 2.318 ;
      RECT 80.19 2.13 80.51 2.318 ;
      RECT 80.19 2.115 80.485 2.318 ;
      RECT 79.39 2.745 79.525 3.04 ;
      RECT 79.65 2.768 79.655 2.955 ;
      RECT 80.37 2.665 80.515 2.9 ;
      RECT 80.53 2.665 80.535 2.89 ;
      RECT 80.565 2.676 80.57 2.87 ;
      RECT 80.56 2.668 80.565 2.875 ;
      RECT 80.54 2.665 80.56 2.88 ;
      RECT 80.535 2.665 80.54 2.888 ;
      RECT 80.525 2.665 80.53 2.893 ;
      RECT 80.515 2.665 80.525 2.898 ;
      RECT 80.345 2.667 80.37 2.9 ;
      RECT 80.295 2.674 80.345 2.9 ;
      RECT 80.29 2.679 80.295 2.9 ;
      RECT 80.251 2.684 80.29 2.901 ;
      RECT 80.165 2.696 80.251 2.902 ;
      RECT 80.156 2.706 80.165 2.902 ;
      RECT 80.07 2.715 80.156 2.904 ;
      RECT 80.046 2.725 80.07 2.906 ;
      RECT 79.96 2.736 80.046 2.907 ;
      RECT 79.93 2.747 79.96 2.909 ;
      RECT 79.9 2.752 79.93 2.911 ;
      RECT 79.875 2.758 79.9 2.914 ;
      RECT 79.86 2.763 79.875 2.915 ;
      RECT 79.815 2.769 79.86 2.915 ;
      RECT 79.81 2.774 79.815 2.916 ;
      RECT 79.79 2.774 79.81 2.918 ;
      RECT 79.77 2.772 79.79 2.923 ;
      RECT 79.735 2.771 79.77 2.93 ;
      RECT 79.705 2.77 79.735 2.94 ;
      RECT 79.655 2.769 79.705 2.95 ;
      RECT 79.565 2.766 79.65 3.04 ;
      RECT 79.54 2.76 79.565 3.04 ;
      RECT 79.525 2.75 79.54 3.04 ;
      RECT 79.34 2.745 79.39 2.96 ;
      RECT 79.33 2.75 79.34 2.95 ;
      RECT 79.57 3.225 79.83 3.485 ;
      RECT 79.57 3.225 79.86 3.378 ;
      RECT 79.57 3.225 79.895 3.363 ;
      RECT 79.825 3.145 80.015 3.355 ;
      RECT 79.815 3.15 80.025 3.348 ;
      RECT 79.78 3.22 80.025 3.348 ;
      RECT 79.81 3.162 79.83 3.485 ;
      RECT 79.795 3.21 80.025 3.348 ;
      RECT 79.8 3.182 79.83 3.485 ;
      RECT 78.88 2.25 78.95 3.355 ;
      RECT 79.615 2.355 79.875 2.615 ;
      RECT 79.195 2.401 79.21 2.61 ;
      RECT 79.531 2.414 79.615 2.565 ;
      RECT 79.445 2.411 79.531 2.565 ;
      RECT 79.406 2.409 79.445 2.565 ;
      RECT 79.32 2.407 79.406 2.565 ;
      RECT 79.26 2.405 79.32 2.576 ;
      RECT 79.225 2.403 79.26 2.594 ;
      RECT 79.21 2.401 79.225 2.605 ;
      RECT 79.18 2.401 79.195 2.618 ;
      RECT 79.17 2.401 79.18 2.623 ;
      RECT 79.145 2.4 79.17 2.628 ;
      RECT 79.13 2.395 79.145 2.634 ;
      RECT 79.125 2.388 79.13 2.639 ;
      RECT 79.1 2.379 79.125 2.645 ;
      RECT 79.055 2.358 79.1 2.658 ;
      RECT 79.045 2.342 79.055 2.668 ;
      RECT 79.03 2.335 79.045 2.678 ;
      RECT 79.02 2.328 79.03 2.695 ;
      RECT 79.015 2.325 79.02 2.725 ;
      RECT 79.01 2.323 79.015 2.755 ;
      RECT 79.005 2.321 79.01 2.792 ;
      RECT 78.99 2.317 79.005 2.859 ;
      RECT 78.99 3.15 79 3.35 ;
      RECT 78.985 2.313 78.99 2.985 ;
      RECT 78.985 3.137 78.99 3.355 ;
      RECT 78.98 2.311 78.985 3.07 ;
      RECT 78.98 3.127 78.985 3.355 ;
      RECT 78.965 2.282 78.98 3.355 ;
      RECT 78.95 2.255 78.965 3.355 ;
      RECT 78.875 2.25 78.88 2.605 ;
      RECT 78.875 2.66 78.88 3.355 ;
      RECT 78.86 2.25 78.875 2.583 ;
      RECT 78.87 2.682 78.875 3.355 ;
      RECT 78.86 2.722 78.87 3.355 ;
      RECT 78.825 2.25 78.86 2.525 ;
      RECT 78.855 2.757 78.86 3.355 ;
      RECT 78.84 2.812 78.855 3.355 ;
      RECT 78.835 2.877 78.84 3.355 ;
      RECT 78.82 2.925 78.835 3.355 ;
      RECT 78.795 2.25 78.825 2.48 ;
      RECT 78.815 2.98 78.82 3.355 ;
      RECT 78.8 3.04 78.815 3.355 ;
      RECT 78.795 3.088 78.8 3.353 ;
      RECT 78.79 2.25 78.795 2.473 ;
      RECT 78.79 3.12 78.795 3.348 ;
      RECT 78.765 2.25 78.79 2.465 ;
      RECT 78.755 2.255 78.765 2.455 ;
      RECT 78.97 3.53 78.99 3.77 ;
      RECT 78.2 3.46 78.205 3.67 ;
      RECT 79.48 3.533 79.49 3.728 ;
      RECT 79.475 3.523 79.48 3.731 ;
      RECT 79.395 3.52 79.475 3.754 ;
      RECT 79.391 3.52 79.395 3.776 ;
      RECT 79.305 3.52 79.391 3.786 ;
      RECT 79.29 3.52 79.305 3.794 ;
      RECT 79.261 3.521 79.29 3.792 ;
      RECT 79.175 3.526 79.261 3.788 ;
      RECT 79.162 3.53 79.175 3.784 ;
      RECT 79.076 3.53 79.162 3.78 ;
      RECT 78.99 3.53 79.076 3.774 ;
      RECT 78.906 3.53 78.97 3.768 ;
      RECT 78.82 3.53 78.906 3.763 ;
      RECT 78.8 3.53 78.82 3.759 ;
      RECT 78.74 3.525 78.8 3.756 ;
      RECT 78.712 3.519 78.74 3.753 ;
      RECT 78.626 3.514 78.712 3.749 ;
      RECT 78.54 3.508 78.626 3.743 ;
      RECT 78.465 3.49 78.54 3.738 ;
      RECT 78.43 3.467 78.465 3.734 ;
      RECT 78.42 3.457 78.43 3.733 ;
      RECT 78.365 3.455 78.42 3.732 ;
      RECT 78.29 3.455 78.365 3.728 ;
      RECT 78.28 3.455 78.29 3.723 ;
      RECT 78.265 3.455 78.28 3.715 ;
      RECT 78.215 3.457 78.265 3.693 ;
      RECT 78.205 3.46 78.215 3.673 ;
      RECT 78.195 3.465 78.2 3.668 ;
      RECT 78.19 3.47 78.195 3.663 ;
      RECT 78.315 2.635 78.575 2.895 ;
      RECT 78.315 2.65 78.595 2.86 ;
      RECT 78.315 2.655 78.605 2.855 ;
      RECT 76.3 2.115 76.56 2.375 ;
      RECT 76.29 2.145 76.56 2.355 ;
      RECT 78.21 2.06 78.47 2.32 ;
      RECT 78.205 2.135 78.21 2.321 ;
      RECT 78.18 2.14 78.205 2.323 ;
      RECT 78.165 2.147 78.18 2.326 ;
      RECT 78.105 2.165 78.165 2.331 ;
      RECT 78.075 2.185 78.105 2.338 ;
      RECT 78.05 2.193 78.075 2.343 ;
      RECT 78.025 2.201 78.05 2.345 ;
      RECT 78.007 2.205 78.025 2.344 ;
      RECT 77.921 2.203 78.007 2.344 ;
      RECT 77.835 2.201 77.921 2.344 ;
      RECT 77.749 2.199 77.835 2.343 ;
      RECT 77.663 2.197 77.749 2.343 ;
      RECT 77.577 2.195 77.663 2.343 ;
      RECT 77.491 2.193 77.577 2.343 ;
      RECT 77.405 2.191 77.491 2.342 ;
      RECT 77.387 2.19 77.405 2.342 ;
      RECT 77.301 2.189 77.387 2.342 ;
      RECT 77.215 2.187 77.301 2.342 ;
      RECT 77.129 2.186 77.215 2.341 ;
      RECT 77.043 2.185 77.129 2.341 ;
      RECT 76.957 2.183 77.043 2.341 ;
      RECT 76.871 2.182 76.957 2.341 ;
      RECT 76.785 2.18 76.871 2.34 ;
      RECT 76.761 2.178 76.785 2.34 ;
      RECT 76.675 2.171 76.761 2.34 ;
      RECT 76.646 2.163 76.675 2.34 ;
      RECT 76.56 2.155 76.646 2.34 ;
      RECT 76.28 2.152 76.29 2.35 ;
      RECT 77.785 3.115 77.79 3.465 ;
      RECT 77.555 3.205 77.695 3.465 ;
      RECT 78.03 2.89 78.075 3.1 ;
      RECT 78.085 2.901 78.095 3.095 ;
      RECT 78.075 2.893 78.085 3.1 ;
      RECT 78.01 2.89 78.03 3.105 ;
      RECT 77.98 2.89 78.01 3.128 ;
      RECT 77.97 2.89 77.98 3.153 ;
      RECT 77.965 2.89 77.97 3.163 ;
      RECT 77.91 2.89 77.965 3.203 ;
      RECT 77.905 2.89 77.91 3.243 ;
      RECT 77.9 2.892 77.905 3.248 ;
      RECT 77.885 2.902 77.9 3.259 ;
      RECT 77.84 2.96 77.885 3.295 ;
      RECT 77.83 3.015 77.84 3.329 ;
      RECT 77.815 3.042 77.83 3.345 ;
      RECT 77.805 3.069 77.815 3.465 ;
      RECT 77.79 3.092 77.805 3.465 ;
      RECT 77.78 3.132 77.785 3.465 ;
      RECT 77.775 3.142 77.78 3.465 ;
      RECT 77.77 3.157 77.775 3.465 ;
      RECT 77.76 3.162 77.77 3.465 ;
      RECT 77.695 3.185 77.76 3.465 ;
      RECT 77.195 2.68 77.385 2.89 ;
      RECT 75.77 2.605 76.03 2.865 ;
      RECT 76.12 2.6 76.215 2.81 ;
      RECT 76.095 2.615 76.105 2.81 ;
      RECT 77.385 2.687 77.395 2.885 ;
      RECT 77.185 2.687 77.195 2.885 ;
      RECT 77.17 2.702 77.185 2.875 ;
      RECT 77.165 2.71 77.17 2.868 ;
      RECT 77.155 2.713 77.165 2.865 ;
      RECT 77.12 2.712 77.155 2.863 ;
      RECT 77.091 2.708 77.12 2.86 ;
      RECT 77.005 2.703 77.091 2.857 ;
      RECT 76.945 2.697 77.005 2.853 ;
      RECT 76.916 2.693 76.945 2.85 ;
      RECT 76.83 2.685 76.916 2.847 ;
      RECT 76.821 2.679 76.83 2.845 ;
      RECT 76.735 2.674 76.821 2.843 ;
      RECT 76.712 2.669 76.735 2.84 ;
      RECT 76.626 2.663 76.712 2.837 ;
      RECT 76.54 2.654 76.626 2.832 ;
      RECT 76.53 2.649 76.54 2.83 ;
      RECT 76.511 2.648 76.53 2.829 ;
      RECT 76.425 2.643 76.511 2.825 ;
      RECT 76.405 2.638 76.425 2.821 ;
      RECT 76.345 2.633 76.405 2.818 ;
      RECT 76.32 2.623 76.345 2.816 ;
      RECT 76.315 2.616 76.32 2.815 ;
      RECT 76.305 2.607 76.315 2.814 ;
      RECT 76.301 2.6 76.305 2.814 ;
      RECT 76.215 2.6 76.301 2.812 ;
      RECT 76.105 2.607 76.12 2.81 ;
      RECT 76.09 2.617 76.095 2.81 ;
      RECT 76.07 2.62 76.09 2.807 ;
      RECT 76.04 2.62 76.07 2.803 ;
      RECT 76.03 2.62 76.04 2.803 ;
      RECT 76.945 3.115 77.205 3.375 ;
      RECT 76.875 3.125 77.205 3.335 ;
      RECT 76.865 3.132 77.205 3.33 ;
      RECT 76.285 3.12 76.545 3.38 ;
      RECT 76.285 3.16 76.65 3.37 ;
      RECT 76.285 3.162 76.655 3.369 ;
      RECT 76.285 3.17 76.66 3.366 ;
      RECT 75.21 2.245 75.31 3.77 ;
      RECT 75.4 3.385 75.45 3.645 ;
      RECT 75.395 2.258 75.4 2.445 ;
      RECT 75.39 3.366 75.4 3.645 ;
      RECT 75.39 2.255 75.395 2.453 ;
      RECT 75.375 2.249 75.39 2.46 ;
      RECT 75.385 3.354 75.39 3.728 ;
      RECT 75.375 3.342 75.385 3.765 ;
      RECT 75.365 2.245 75.375 2.467 ;
      RECT 75.365 3.327 75.375 3.77 ;
      RECT 75.36 2.245 75.365 2.475 ;
      RECT 75.34 3.297 75.365 3.77 ;
      RECT 75.32 2.245 75.36 2.523 ;
      RECT 75.33 3.257 75.34 3.77 ;
      RECT 75.32 3.212 75.33 3.77 ;
      RECT 75.315 2.245 75.32 2.593 ;
      RECT 75.315 3.17 75.32 3.77 ;
      RECT 75.31 2.245 75.315 3.07 ;
      RECT 75.31 3.152 75.315 3.77 ;
      RECT 75.2 2.248 75.21 3.77 ;
      RECT 75.185 2.255 75.2 3.766 ;
      RECT 75.18 2.265 75.185 3.761 ;
      RECT 75.175 2.465 75.18 3.653 ;
      RECT 75.17 2.55 75.175 3.205 ;
      RECT 74.045 7.77 74.335 8 ;
      RECT 74.105 6.29 74.275 8 ;
      RECT 74.055 6.655 74.405 7.005 ;
      RECT 74.045 6.29 74.335 6.52 ;
      RECT 73.64 2.395 73.745 2.965 ;
      RECT 73.64 2.73 73.965 2.96 ;
      RECT 73.64 2.76 74.135 2.93 ;
      RECT 73.64 2.395 73.83 2.96 ;
      RECT 73.055 2.36 73.345 2.59 ;
      RECT 73.055 2.395 73.83 2.565 ;
      RECT 73.115 0.88 73.285 2.59 ;
      RECT 73.055 0.88 73.345 1.11 ;
      RECT 73.055 7.77 73.345 8 ;
      RECT 73.115 6.29 73.285 8 ;
      RECT 73.055 6.29 73.345 6.52 ;
      RECT 73.055 6.325 73.91 6.485 ;
      RECT 73.74 5.92 73.91 6.485 ;
      RECT 73.055 6.32 73.45 6.485 ;
      RECT 73.675 5.92 73.965 6.15 ;
      RECT 73.675 5.95 74.135 6.12 ;
      RECT 72.685 2.73 72.975 2.96 ;
      RECT 72.685 2.76 73.145 2.93 ;
      RECT 72.75 1.655 72.915 2.96 ;
      RECT 71.265 1.625 71.555 1.855 ;
      RECT 71.265 1.655 72.915 1.825 ;
      RECT 71.325 0.885 71.495 1.855 ;
      RECT 71.265 0.885 71.555 1.115 ;
      RECT 71.265 7.765 71.555 7.995 ;
      RECT 71.325 7.025 71.495 7.995 ;
      RECT 71.325 7.12 72.915 7.29 ;
      RECT 72.745 5.92 72.915 7.29 ;
      RECT 71.265 7.025 71.555 7.255 ;
      RECT 72.685 5.92 72.975 6.15 ;
      RECT 72.685 5.95 73.145 6.12 ;
      RECT 69.3 3.43 69.65 3.78 ;
      RECT 69.39 2.025 69.56 3.78 ;
      RECT 71.695 1.965 72.045 2.315 ;
      RECT 69.39 2.025 71.01 2.2 ;
      RECT 69.39 2.025 72.045 2.195 ;
      RECT 71.72 6.655 72.045 6.98 ;
      RECT 67.095 6.61 67.445 6.96 ;
      RECT 71.695 6.655 72.045 6.885 ;
      RECT 66.935 6.655 67.445 6.885 ;
      RECT 66.765 6.685 72.045 6.855 ;
      RECT 70.92 2.365 71.24 2.685 ;
      RECT 70.89 2.365 71.24 2.595 ;
      RECT 70.72 2.395 71.24 2.565 ;
      RECT 70.92 6.225 71.24 6.545 ;
      RECT 70.89 6.285 71.24 6.515 ;
      RECT 70.72 6.315 71.24 6.485 ;
      RECT 66.7 3.665 66.74 3.925 ;
      RECT 66.74 3.645 66.745 3.655 ;
      RECT 68.07 2.89 68.08 3.111 ;
      RECT 68 2.885 68.07 3.236 ;
      RECT 67.99 2.885 68 3.363 ;
      RECT 67.965 2.885 67.99 3.41 ;
      RECT 67.94 2.885 67.965 3.488 ;
      RECT 67.92 2.885 67.94 3.558 ;
      RECT 67.895 2.885 67.92 3.598 ;
      RECT 67.885 2.885 67.895 3.618 ;
      RECT 67.875 2.887 67.885 3.626 ;
      RECT 67.87 2.892 67.875 3.083 ;
      RECT 67.87 3.092 67.875 3.627 ;
      RECT 67.865 3.137 67.87 3.628 ;
      RECT 67.855 3.202 67.865 3.629 ;
      RECT 67.845 3.297 67.855 3.631 ;
      RECT 67.84 3.35 67.845 3.633 ;
      RECT 67.835 3.37 67.84 3.634 ;
      RECT 67.78 3.395 67.835 3.64 ;
      RECT 67.74 3.43 67.78 3.649 ;
      RECT 67.73 3.447 67.74 3.654 ;
      RECT 67.721 3.453 67.73 3.656 ;
      RECT 67.635 3.491 67.721 3.667 ;
      RECT 67.63 3.53 67.635 3.677 ;
      RECT 67.555 3.537 67.63 3.687 ;
      RECT 67.535 3.547 67.555 3.698 ;
      RECT 67.505 3.554 67.535 3.706 ;
      RECT 67.48 3.561 67.505 3.713 ;
      RECT 67.456 3.567 67.48 3.718 ;
      RECT 67.37 3.58 67.456 3.73 ;
      RECT 67.292 3.587 67.37 3.748 ;
      RECT 67.206 3.582 67.292 3.766 ;
      RECT 67.12 3.577 67.206 3.786 ;
      RECT 67.04 3.571 67.12 3.803 ;
      RECT 66.975 3.567 67.04 3.832 ;
      RECT 66.97 3.281 66.975 3.305 ;
      RECT 66.96 3.557 66.975 3.86 ;
      RECT 66.965 3.275 66.97 3.345 ;
      RECT 66.96 3.269 66.965 3.415 ;
      RECT 66.955 3.263 66.96 3.493 ;
      RECT 66.955 3.54 66.96 3.925 ;
      RECT 66.947 3.26 66.955 3.925 ;
      RECT 66.861 3.258 66.947 3.925 ;
      RECT 66.775 3.256 66.861 3.925 ;
      RECT 66.765 3.257 66.775 3.925 ;
      RECT 66.76 3.262 66.765 3.925 ;
      RECT 66.75 3.275 66.76 3.925 ;
      RECT 66.745 3.297 66.75 3.925 ;
      RECT 66.74 3.657 66.745 3.925 ;
      RECT 67.37 3.125 67.375 3.345 ;
      RECT 67.875 2.16 67.91 2.42 ;
      RECT 67.86 2.16 67.875 2.428 ;
      RECT 67.831 2.16 67.86 2.45 ;
      RECT 67.745 2.16 67.831 2.51 ;
      RECT 67.725 2.16 67.745 2.575 ;
      RECT 67.665 2.16 67.725 2.74 ;
      RECT 67.66 2.16 67.665 2.888 ;
      RECT 67.655 2.16 67.66 2.9 ;
      RECT 67.65 2.16 67.655 2.926 ;
      RECT 67.62 2.346 67.65 3.006 ;
      RECT 67.615 2.394 67.62 3.095 ;
      RECT 67.61 2.408 67.615 3.11 ;
      RECT 67.605 2.427 67.61 3.14 ;
      RECT 67.6 2.442 67.605 3.156 ;
      RECT 67.595 2.457 67.6 3.178 ;
      RECT 67.59 2.477 67.595 3.2 ;
      RECT 67.58 2.497 67.59 3.233 ;
      RECT 67.565 2.539 67.58 3.295 ;
      RECT 67.56 2.57 67.565 3.335 ;
      RECT 67.555 2.582 67.56 3.34 ;
      RECT 67.55 2.594 67.555 3.345 ;
      RECT 67.545 2.607 67.55 3.345 ;
      RECT 67.54 2.625 67.545 3.345 ;
      RECT 67.535 2.645 67.54 3.345 ;
      RECT 67.53 2.657 67.535 3.345 ;
      RECT 67.525 2.67 67.53 3.345 ;
      RECT 67.505 2.705 67.525 3.345 ;
      RECT 67.455 2.807 67.505 3.345 ;
      RECT 67.45 2.892 67.455 3.345 ;
      RECT 67.445 2.9 67.45 3.345 ;
      RECT 67.44 2.917 67.445 3.345 ;
      RECT 67.435 2.932 67.44 3.345 ;
      RECT 67.4 2.997 67.435 3.345 ;
      RECT 67.385 3.062 67.4 3.345 ;
      RECT 67.38 3.092 67.385 3.345 ;
      RECT 67.375 3.117 67.38 3.345 ;
      RECT 67.36 3.127 67.37 3.345 ;
      RECT 67.345 3.14 67.36 3.338 ;
      RECT 67.09 2.73 67.16 2.94 ;
      RECT 66.88 2.707 66.885 2.9 ;
      RECT 64.335 2.635 64.595 2.895 ;
      RECT 67.17 2.917 67.175 2.92 ;
      RECT 67.16 2.735 67.17 2.935 ;
      RECT 67.061 2.728 67.09 2.94 ;
      RECT 66.975 2.72 67.061 2.94 ;
      RECT 66.96 2.714 66.975 2.938 ;
      RECT 66.94 2.713 66.96 2.925 ;
      RECT 66.935 2.712 66.94 2.908 ;
      RECT 66.885 2.709 66.935 2.903 ;
      RECT 66.855 2.706 66.88 2.898 ;
      RECT 66.835 2.704 66.855 2.893 ;
      RECT 66.82 2.702 66.835 2.89 ;
      RECT 66.79 2.7 66.82 2.888 ;
      RECT 66.725 2.696 66.79 2.88 ;
      RECT 66.695 2.691 66.725 2.875 ;
      RECT 66.675 2.689 66.695 2.873 ;
      RECT 66.645 2.686 66.675 2.868 ;
      RECT 66.585 2.682 66.645 2.86 ;
      RECT 66.58 2.679 66.585 2.855 ;
      RECT 66.51 2.677 66.58 2.85 ;
      RECT 66.481 2.673 66.51 2.843 ;
      RECT 66.395 2.668 66.481 2.835 ;
      RECT 66.361 2.663 66.395 2.827 ;
      RECT 66.275 2.655 66.361 2.819 ;
      RECT 66.236 2.648 66.275 2.811 ;
      RECT 66.15 2.643 66.236 2.803 ;
      RECT 66.085 2.637 66.15 2.793 ;
      RECT 66.065 2.632 66.085 2.788 ;
      RECT 66.056 2.629 66.065 2.787 ;
      RECT 65.97 2.625 66.056 2.781 ;
      RECT 65.93 2.621 65.97 2.773 ;
      RECT 65.91 2.617 65.93 2.771 ;
      RECT 65.85 2.617 65.91 2.768 ;
      RECT 65.83 2.62 65.85 2.766 ;
      RECT 65.809 2.62 65.83 2.766 ;
      RECT 65.723 2.622 65.809 2.77 ;
      RECT 65.637 2.624 65.723 2.776 ;
      RECT 65.551 2.626 65.637 2.783 ;
      RECT 65.465 2.629 65.551 2.789 ;
      RECT 65.431 2.63 65.465 2.794 ;
      RECT 65.345 2.633 65.431 2.799 ;
      RECT 65.316 2.64 65.345 2.804 ;
      RECT 65.23 2.64 65.316 2.809 ;
      RECT 65.197 2.64 65.23 2.814 ;
      RECT 65.111 2.642 65.197 2.819 ;
      RECT 65.025 2.644 65.111 2.826 ;
      RECT 64.961 2.646 65.025 2.832 ;
      RECT 64.875 2.648 64.961 2.838 ;
      RECT 64.872 2.65 64.875 2.841 ;
      RECT 64.786 2.651 64.872 2.845 ;
      RECT 64.7 2.654 64.786 2.852 ;
      RECT 64.681 2.656 64.7 2.856 ;
      RECT 64.595 2.658 64.681 2.861 ;
      RECT 64.325 2.67 64.335 2.865 ;
      RECT 66.505 7.765 66.795 7.995 ;
      RECT 66.565 7.025 66.735 7.995 ;
      RECT 66.455 7.055 66.83 7.425 ;
      RECT 66.505 7.025 66.795 7.425 ;
      RECT 66.56 2.25 66.745 2.46 ;
      RECT 66.555 2.251 66.75 2.458 ;
      RECT 66.55 2.256 66.76 2.453 ;
      RECT 66.545 2.232 66.55 2.45 ;
      RECT 66.515 2.229 66.545 2.443 ;
      RECT 66.51 2.225 66.515 2.434 ;
      RECT 66.475 2.256 66.76 2.429 ;
      RECT 66.25 2.165 66.51 2.425 ;
      RECT 66.55 2.234 66.555 2.453 ;
      RECT 66.555 2.235 66.56 2.458 ;
      RECT 66.25 2.247 66.63 2.425 ;
      RECT 66.25 2.245 66.615 2.425 ;
      RECT 66.25 2.24 66.605 2.425 ;
      RECT 66.205 3.155 66.255 3.44 ;
      RECT 66.15 3.125 66.155 3.44 ;
      RECT 66.12 3.105 66.125 3.44 ;
      RECT 66.27 3.155 66.33 3.415 ;
      RECT 66.265 3.155 66.27 3.423 ;
      RECT 66.255 3.155 66.265 3.435 ;
      RECT 66.17 3.145 66.205 3.44 ;
      RECT 66.165 3.132 66.17 3.44 ;
      RECT 66.155 3.127 66.165 3.44 ;
      RECT 66.135 3.117 66.15 3.44 ;
      RECT 66.125 3.11 66.135 3.44 ;
      RECT 66.115 3.102 66.12 3.44 ;
      RECT 66.085 3.092 66.115 3.44 ;
      RECT 66.07 3.08 66.085 3.44 ;
      RECT 66.055 3.07 66.07 3.435 ;
      RECT 66.035 3.06 66.055 3.41 ;
      RECT 66.025 3.052 66.035 3.387 ;
      RECT 65.995 3.035 66.025 3.377 ;
      RECT 65.99 3.012 65.995 3.368 ;
      RECT 65.985 2.999 65.99 3.366 ;
      RECT 65.97 2.975 65.985 3.36 ;
      RECT 65.965 2.951 65.97 3.354 ;
      RECT 65.955 2.94 65.965 3.349 ;
      RECT 65.95 2.93 65.955 3.345 ;
      RECT 65.945 2.922 65.95 3.342 ;
      RECT 65.935 2.917 65.945 3.338 ;
      RECT 65.93 2.912 65.935 3.334 ;
      RECT 65.845 2.91 65.93 3.309 ;
      RECT 65.815 2.91 65.845 3.275 ;
      RECT 65.8 2.91 65.815 3.258 ;
      RECT 65.745 2.91 65.8 3.203 ;
      RECT 65.74 2.915 65.745 3.152 ;
      RECT 65.73 2.92 65.74 3.142 ;
      RECT 65.725 2.93 65.73 3.128 ;
      RECT 65.675 3.67 65.935 3.93 ;
      RECT 65.595 3.685 65.935 3.906 ;
      RECT 65.575 3.685 65.935 3.901 ;
      RECT 65.551 3.685 65.935 3.899 ;
      RECT 65.465 3.685 65.935 3.894 ;
      RECT 65.315 3.625 65.575 3.89 ;
      RECT 65.27 3.685 65.935 3.885 ;
      RECT 65.265 3.692 65.935 3.88 ;
      RECT 65.28 3.68 65.595 3.89 ;
      RECT 65.17 2.115 65.43 2.375 ;
      RECT 65.17 2.172 65.435 2.368 ;
      RECT 65.17 2.202 65.44 2.3 ;
      RECT 65.23 2.633 65.345 2.635 ;
      RECT 65.316 2.63 65.345 2.635 ;
      RECT 64.34 3.634 64.365 3.874 ;
      RECT 64.325 3.637 64.415 3.868 ;
      RECT 64.32 3.642 64.501 3.863 ;
      RECT 64.315 3.65 64.565 3.861 ;
      RECT 64.315 3.65 64.575 3.86 ;
      RECT 64.31 3.657 64.585 3.853 ;
      RECT 64.31 3.657 64.671 3.842 ;
      RECT 64.305 3.692 64.671 3.838 ;
      RECT 64.305 3.692 64.68 3.827 ;
      RECT 64.585 3.565 64.845 3.825 ;
      RECT 64.295 3.742 64.845 3.823 ;
      RECT 64.565 3.61 64.585 3.858 ;
      RECT 64.501 3.613 64.565 3.862 ;
      RECT 64.415 3.618 64.501 3.867 ;
      RECT 64.345 3.629 64.845 3.825 ;
      RECT 64.365 3.623 64.415 3.872 ;
      RECT 64.49 2.1 64.5 2.362 ;
      RECT 64.48 2.157 64.49 2.365 ;
      RECT 64.455 2.162 64.48 2.371 ;
      RECT 64.43 2.166 64.455 2.383 ;
      RECT 64.42 2.169 64.43 2.393 ;
      RECT 64.415 2.17 64.42 2.398 ;
      RECT 64.41 2.171 64.415 2.403 ;
      RECT 64.405 2.172 64.41 2.405 ;
      RECT 64.38 2.175 64.405 2.408 ;
      RECT 64.35 2.181 64.38 2.411 ;
      RECT 64.285 2.192 64.35 2.414 ;
      RECT 64.24 2.2 64.285 2.418 ;
      RECT 64.225 2.2 64.24 2.426 ;
      RECT 64.22 2.201 64.225 2.433 ;
      RECT 64.215 2.203 64.22 2.436 ;
      RECT 64.21 2.207 64.215 2.439 ;
      RECT 64.2 2.215 64.21 2.443 ;
      RECT 64.195 2.228 64.2 2.448 ;
      RECT 64.19 2.236 64.195 2.45 ;
      RECT 64.185 2.242 64.19 2.45 ;
      RECT 64.18 2.246 64.185 2.453 ;
      RECT 64.175 2.248 64.18 2.456 ;
      RECT 64.17 2.251 64.175 2.459 ;
      RECT 64.16 2.256 64.17 2.463 ;
      RECT 64.155 2.262 64.16 2.468 ;
      RECT 64.145 2.268 64.155 2.472 ;
      RECT 64.13 2.275 64.145 2.478 ;
      RECT 64.101 2.289 64.13 2.488 ;
      RECT 64.015 2.324 64.101 2.52 ;
      RECT 63.995 2.357 64.015 2.549 ;
      RECT 63.975 2.37 63.995 2.56 ;
      RECT 63.955 2.382 63.975 2.571 ;
      RECT 63.905 2.404 63.955 2.591 ;
      RECT 63.89 2.422 63.905 2.608 ;
      RECT 63.885 2.428 63.89 2.611 ;
      RECT 63.88 2.432 63.885 2.614 ;
      RECT 63.875 2.436 63.88 2.618 ;
      RECT 63.87 2.438 63.875 2.621 ;
      RECT 63.86 2.445 63.87 2.624 ;
      RECT 63.855 2.45 63.86 2.628 ;
      RECT 63.85 2.452 63.855 2.631 ;
      RECT 63.845 2.456 63.85 2.634 ;
      RECT 63.84 2.458 63.845 2.638 ;
      RECT 63.825 2.463 63.84 2.643 ;
      RECT 63.82 2.468 63.825 2.646 ;
      RECT 63.815 2.476 63.82 2.649 ;
      RECT 63.81 2.478 63.815 2.652 ;
      RECT 63.805 2.48 63.81 2.655 ;
      RECT 63.795 2.482 63.805 2.661 ;
      RECT 63.76 2.496 63.795 2.673 ;
      RECT 63.75 2.511 63.76 2.683 ;
      RECT 63.675 2.54 63.75 2.707 ;
      RECT 63.67 2.565 63.675 2.73 ;
      RECT 63.655 2.569 63.67 2.736 ;
      RECT 63.645 2.577 63.655 2.741 ;
      RECT 63.615 2.59 63.645 2.745 ;
      RECT 63.605 2.605 63.615 2.75 ;
      RECT 63.595 2.61 63.605 2.753 ;
      RECT 63.59 2.612 63.595 2.755 ;
      RECT 63.575 2.615 63.59 2.758 ;
      RECT 63.57 2.617 63.575 2.761 ;
      RECT 63.55 2.622 63.57 2.765 ;
      RECT 63.52 2.627 63.55 2.773 ;
      RECT 63.495 2.634 63.52 2.781 ;
      RECT 63.49 2.639 63.495 2.786 ;
      RECT 63.46 2.642 63.49 2.79 ;
      RECT 63.42 2.645 63.46 2.8 ;
      RECT 63.385 2.642 63.42 2.812 ;
      RECT 63.375 2.638 63.385 2.819 ;
      RECT 63.35 2.634 63.375 2.825 ;
      RECT 63.345 2.63 63.35 2.83 ;
      RECT 63.305 2.627 63.345 2.83 ;
      RECT 63.29 2.612 63.305 2.831 ;
      RECT 63.267 2.6 63.29 2.831 ;
      RECT 63.181 2.6 63.267 2.832 ;
      RECT 63.095 2.6 63.181 2.834 ;
      RECT 63.075 2.6 63.095 2.831 ;
      RECT 63.07 2.605 63.075 2.826 ;
      RECT 63.065 2.61 63.07 2.824 ;
      RECT 63.055 2.62 63.065 2.822 ;
      RECT 63.05 2.626 63.055 2.815 ;
      RECT 63.045 2.628 63.05 2.8 ;
      RECT 63.04 2.632 63.045 2.79 ;
      RECT 64.5 2.1 64.75 2.36 ;
      RECT 62.225 3.635 62.485 3.895 ;
      RECT 64.52 3.125 64.525 3.335 ;
      RECT 64.525 3.13 64.535 3.33 ;
      RECT 64.475 3.125 64.52 3.35 ;
      RECT 64.465 3.125 64.475 3.37 ;
      RECT 64.446 3.125 64.465 3.375 ;
      RECT 64.36 3.125 64.446 3.372 ;
      RECT 64.33 3.127 64.36 3.37 ;
      RECT 64.275 3.137 64.33 3.368 ;
      RECT 64.21 3.151 64.275 3.366 ;
      RECT 64.205 3.159 64.21 3.365 ;
      RECT 64.19 3.162 64.205 3.363 ;
      RECT 64.125 3.172 64.19 3.359 ;
      RECT 64.077 3.186 64.125 3.36 ;
      RECT 63.991 3.203 64.077 3.374 ;
      RECT 63.905 3.224 63.991 3.391 ;
      RECT 63.885 3.237 63.905 3.401 ;
      RECT 63.84 3.245 63.885 3.408 ;
      RECT 63.805 3.253 63.84 3.416 ;
      RECT 63.771 3.261 63.805 3.424 ;
      RECT 63.685 3.275 63.771 3.436 ;
      RECT 63.65 3.292 63.685 3.448 ;
      RECT 63.641 3.301 63.65 3.452 ;
      RECT 63.555 3.319 63.641 3.469 ;
      RECT 63.496 3.346 63.555 3.496 ;
      RECT 63.41 3.373 63.496 3.524 ;
      RECT 63.39 3.395 63.41 3.544 ;
      RECT 63.33 3.41 63.39 3.56 ;
      RECT 63.32 3.422 63.33 3.573 ;
      RECT 63.315 3.427 63.32 3.576 ;
      RECT 63.305 3.43 63.315 3.579 ;
      RECT 63.3 3.432 63.305 3.582 ;
      RECT 63.27 3.44 63.3 3.589 ;
      RECT 63.255 3.447 63.27 3.597 ;
      RECT 63.245 3.452 63.255 3.601 ;
      RECT 63.24 3.455 63.245 3.604 ;
      RECT 63.23 3.457 63.24 3.607 ;
      RECT 63.195 3.467 63.23 3.616 ;
      RECT 63.12 3.49 63.195 3.638 ;
      RECT 63.1 3.508 63.12 3.656 ;
      RECT 63.07 3.515 63.1 3.666 ;
      RECT 63.05 3.523 63.07 3.676 ;
      RECT 63.04 3.529 63.05 3.683 ;
      RECT 63.021 3.534 63.04 3.689 ;
      RECT 62.935 3.554 63.021 3.709 ;
      RECT 62.92 3.574 62.935 3.728 ;
      RECT 62.875 3.586 62.92 3.739 ;
      RECT 62.81 3.607 62.875 3.762 ;
      RECT 62.77 3.627 62.81 3.783 ;
      RECT 62.76 3.637 62.77 3.793 ;
      RECT 62.71 3.649 62.76 3.804 ;
      RECT 62.69 3.665 62.71 3.816 ;
      RECT 62.66 3.675 62.69 3.822 ;
      RECT 62.65 3.68 62.66 3.824 ;
      RECT 62.581 3.681 62.65 3.83 ;
      RECT 62.495 3.683 62.581 3.84 ;
      RECT 62.485 3.684 62.495 3.845 ;
      RECT 63.755 3.71 63.945 3.92 ;
      RECT 63.745 3.715 63.955 3.913 ;
      RECT 63.73 3.715 63.955 3.878 ;
      RECT 63.65 3.6 63.91 3.86 ;
      RECT 62.565 3.13 62.75 3.425 ;
      RECT 62.555 3.13 62.75 3.423 ;
      RECT 62.54 3.13 62.755 3.418 ;
      RECT 62.54 3.13 62.76 3.415 ;
      RECT 62.535 3.13 62.76 3.413 ;
      RECT 62.53 3.385 62.76 3.403 ;
      RECT 62.535 3.13 62.795 3.39 ;
      RECT 62.495 2.165 62.755 2.425 ;
      RECT 62.305 2.09 62.391 2.423 ;
      RECT 62.28 2.094 62.435 2.419 ;
      RECT 62.391 2.086 62.435 2.419 ;
      RECT 62.391 2.087 62.44 2.418 ;
      RECT 62.305 2.092 62.455 2.417 ;
      RECT 62.28 2.1 62.495 2.416 ;
      RECT 62.275 2.095 62.455 2.411 ;
      RECT 62.265 2.11 62.495 2.318 ;
      RECT 62.265 2.162 62.695 2.318 ;
      RECT 62.265 2.155 62.675 2.318 ;
      RECT 62.265 2.142 62.645 2.318 ;
      RECT 62.265 2.13 62.585 2.318 ;
      RECT 62.265 2.115 62.56 2.318 ;
      RECT 61.465 2.745 61.6 3.04 ;
      RECT 61.725 2.768 61.73 2.955 ;
      RECT 62.445 2.665 62.59 2.9 ;
      RECT 62.605 2.665 62.61 2.89 ;
      RECT 62.64 2.676 62.645 2.87 ;
      RECT 62.635 2.668 62.64 2.875 ;
      RECT 62.615 2.665 62.635 2.88 ;
      RECT 62.61 2.665 62.615 2.888 ;
      RECT 62.6 2.665 62.605 2.893 ;
      RECT 62.59 2.665 62.6 2.898 ;
      RECT 62.42 2.667 62.445 2.9 ;
      RECT 62.37 2.674 62.42 2.9 ;
      RECT 62.365 2.679 62.37 2.9 ;
      RECT 62.326 2.684 62.365 2.901 ;
      RECT 62.24 2.696 62.326 2.902 ;
      RECT 62.231 2.706 62.24 2.902 ;
      RECT 62.145 2.715 62.231 2.904 ;
      RECT 62.121 2.725 62.145 2.906 ;
      RECT 62.035 2.736 62.121 2.907 ;
      RECT 62.005 2.747 62.035 2.909 ;
      RECT 61.975 2.752 62.005 2.911 ;
      RECT 61.95 2.758 61.975 2.914 ;
      RECT 61.935 2.763 61.95 2.915 ;
      RECT 61.89 2.769 61.935 2.915 ;
      RECT 61.885 2.774 61.89 2.916 ;
      RECT 61.865 2.774 61.885 2.918 ;
      RECT 61.845 2.772 61.865 2.923 ;
      RECT 61.81 2.771 61.845 2.93 ;
      RECT 61.78 2.77 61.81 2.94 ;
      RECT 61.73 2.769 61.78 2.95 ;
      RECT 61.64 2.766 61.725 3.04 ;
      RECT 61.615 2.76 61.64 3.04 ;
      RECT 61.6 2.75 61.615 3.04 ;
      RECT 61.415 2.745 61.465 2.96 ;
      RECT 61.405 2.75 61.415 2.95 ;
      RECT 61.645 3.225 61.905 3.485 ;
      RECT 61.645 3.225 61.935 3.378 ;
      RECT 61.645 3.225 61.97 3.363 ;
      RECT 61.9 3.145 62.09 3.355 ;
      RECT 61.89 3.15 62.1 3.348 ;
      RECT 61.855 3.22 62.1 3.348 ;
      RECT 61.885 3.162 61.905 3.485 ;
      RECT 61.87 3.21 62.1 3.348 ;
      RECT 61.875 3.182 61.905 3.485 ;
      RECT 60.955 2.25 61.025 3.355 ;
      RECT 61.69 2.355 61.95 2.615 ;
      RECT 61.27 2.401 61.285 2.61 ;
      RECT 61.606 2.414 61.69 2.565 ;
      RECT 61.52 2.411 61.606 2.565 ;
      RECT 61.481 2.409 61.52 2.565 ;
      RECT 61.395 2.407 61.481 2.565 ;
      RECT 61.335 2.405 61.395 2.576 ;
      RECT 61.3 2.403 61.335 2.594 ;
      RECT 61.285 2.401 61.3 2.605 ;
      RECT 61.255 2.401 61.27 2.618 ;
      RECT 61.245 2.401 61.255 2.623 ;
      RECT 61.22 2.4 61.245 2.628 ;
      RECT 61.205 2.395 61.22 2.634 ;
      RECT 61.2 2.388 61.205 2.639 ;
      RECT 61.175 2.379 61.2 2.645 ;
      RECT 61.13 2.358 61.175 2.658 ;
      RECT 61.12 2.342 61.13 2.668 ;
      RECT 61.105 2.335 61.12 2.678 ;
      RECT 61.095 2.328 61.105 2.695 ;
      RECT 61.09 2.325 61.095 2.725 ;
      RECT 61.085 2.323 61.09 2.755 ;
      RECT 61.08 2.321 61.085 2.792 ;
      RECT 61.065 2.317 61.08 2.859 ;
      RECT 61.065 3.15 61.075 3.35 ;
      RECT 61.06 2.313 61.065 2.985 ;
      RECT 61.06 3.137 61.065 3.355 ;
      RECT 61.055 2.311 61.06 3.07 ;
      RECT 61.055 3.127 61.06 3.355 ;
      RECT 61.04 2.282 61.055 3.355 ;
      RECT 61.025 2.255 61.04 3.355 ;
      RECT 60.95 2.25 60.955 2.605 ;
      RECT 60.95 2.66 60.955 3.355 ;
      RECT 60.935 2.25 60.95 2.583 ;
      RECT 60.945 2.682 60.95 3.355 ;
      RECT 60.935 2.722 60.945 3.355 ;
      RECT 60.9 2.25 60.935 2.525 ;
      RECT 60.93 2.757 60.935 3.355 ;
      RECT 60.915 2.812 60.93 3.355 ;
      RECT 60.91 2.877 60.915 3.355 ;
      RECT 60.895 2.925 60.91 3.355 ;
      RECT 60.87 2.25 60.9 2.48 ;
      RECT 60.89 2.98 60.895 3.355 ;
      RECT 60.875 3.04 60.89 3.355 ;
      RECT 60.87 3.088 60.875 3.353 ;
      RECT 60.865 2.25 60.87 2.473 ;
      RECT 60.865 3.12 60.87 3.348 ;
      RECT 60.84 2.25 60.865 2.465 ;
      RECT 60.83 2.255 60.84 2.455 ;
      RECT 61.045 3.53 61.065 3.77 ;
      RECT 60.275 3.46 60.28 3.67 ;
      RECT 61.555 3.533 61.565 3.728 ;
      RECT 61.55 3.523 61.555 3.731 ;
      RECT 61.47 3.52 61.55 3.754 ;
      RECT 61.466 3.52 61.47 3.776 ;
      RECT 61.38 3.52 61.466 3.786 ;
      RECT 61.365 3.52 61.38 3.794 ;
      RECT 61.336 3.521 61.365 3.792 ;
      RECT 61.25 3.526 61.336 3.788 ;
      RECT 61.237 3.53 61.25 3.784 ;
      RECT 61.151 3.53 61.237 3.78 ;
      RECT 61.065 3.53 61.151 3.774 ;
      RECT 60.981 3.53 61.045 3.768 ;
      RECT 60.895 3.53 60.981 3.763 ;
      RECT 60.875 3.53 60.895 3.759 ;
      RECT 60.815 3.525 60.875 3.756 ;
      RECT 60.787 3.519 60.815 3.753 ;
      RECT 60.701 3.514 60.787 3.749 ;
      RECT 60.615 3.508 60.701 3.743 ;
      RECT 60.54 3.49 60.615 3.738 ;
      RECT 60.505 3.467 60.54 3.734 ;
      RECT 60.495 3.457 60.505 3.733 ;
      RECT 60.44 3.455 60.495 3.732 ;
      RECT 60.365 3.455 60.44 3.728 ;
      RECT 60.355 3.455 60.365 3.723 ;
      RECT 60.34 3.455 60.355 3.715 ;
      RECT 60.29 3.457 60.34 3.693 ;
      RECT 60.28 3.46 60.29 3.673 ;
      RECT 60.27 3.465 60.275 3.668 ;
      RECT 60.265 3.47 60.27 3.663 ;
      RECT 60.39 2.635 60.65 2.895 ;
      RECT 60.39 2.65 60.67 2.86 ;
      RECT 60.39 2.655 60.68 2.855 ;
      RECT 58.375 2.115 58.635 2.375 ;
      RECT 58.365 2.145 58.635 2.355 ;
      RECT 60.285 2.06 60.545 2.32 ;
      RECT 60.28 2.135 60.285 2.321 ;
      RECT 60.255 2.14 60.28 2.323 ;
      RECT 60.24 2.147 60.255 2.326 ;
      RECT 60.18 2.165 60.24 2.331 ;
      RECT 60.15 2.185 60.18 2.338 ;
      RECT 60.125 2.193 60.15 2.343 ;
      RECT 60.1 2.201 60.125 2.345 ;
      RECT 60.082 2.205 60.1 2.344 ;
      RECT 59.996 2.203 60.082 2.344 ;
      RECT 59.91 2.201 59.996 2.344 ;
      RECT 59.824 2.199 59.91 2.343 ;
      RECT 59.738 2.197 59.824 2.343 ;
      RECT 59.652 2.195 59.738 2.343 ;
      RECT 59.566 2.193 59.652 2.343 ;
      RECT 59.48 2.191 59.566 2.342 ;
      RECT 59.462 2.19 59.48 2.342 ;
      RECT 59.376 2.189 59.462 2.342 ;
      RECT 59.29 2.187 59.376 2.342 ;
      RECT 59.204 2.186 59.29 2.341 ;
      RECT 59.118 2.185 59.204 2.341 ;
      RECT 59.032 2.183 59.118 2.341 ;
      RECT 58.946 2.182 59.032 2.341 ;
      RECT 58.86 2.18 58.946 2.34 ;
      RECT 58.836 2.178 58.86 2.34 ;
      RECT 58.75 2.171 58.836 2.34 ;
      RECT 58.721 2.163 58.75 2.34 ;
      RECT 58.635 2.155 58.721 2.34 ;
      RECT 58.355 2.152 58.365 2.35 ;
      RECT 59.86 3.115 59.865 3.465 ;
      RECT 59.63 3.205 59.77 3.465 ;
      RECT 60.105 2.89 60.15 3.1 ;
      RECT 60.16 2.901 60.17 3.095 ;
      RECT 60.15 2.893 60.16 3.1 ;
      RECT 60.085 2.89 60.105 3.105 ;
      RECT 60.055 2.89 60.085 3.128 ;
      RECT 60.045 2.89 60.055 3.153 ;
      RECT 60.04 2.89 60.045 3.163 ;
      RECT 59.985 2.89 60.04 3.203 ;
      RECT 59.98 2.89 59.985 3.243 ;
      RECT 59.975 2.892 59.98 3.248 ;
      RECT 59.96 2.902 59.975 3.259 ;
      RECT 59.915 2.96 59.96 3.295 ;
      RECT 59.905 3.015 59.915 3.329 ;
      RECT 59.89 3.042 59.905 3.345 ;
      RECT 59.88 3.069 59.89 3.465 ;
      RECT 59.865 3.092 59.88 3.465 ;
      RECT 59.855 3.132 59.86 3.465 ;
      RECT 59.85 3.142 59.855 3.465 ;
      RECT 59.845 3.157 59.85 3.465 ;
      RECT 59.835 3.162 59.845 3.465 ;
      RECT 59.77 3.185 59.835 3.465 ;
      RECT 59.27 2.68 59.46 2.89 ;
      RECT 57.845 2.605 58.105 2.865 ;
      RECT 58.195 2.6 58.29 2.81 ;
      RECT 58.17 2.615 58.18 2.81 ;
      RECT 59.46 2.687 59.47 2.885 ;
      RECT 59.26 2.687 59.27 2.885 ;
      RECT 59.245 2.702 59.26 2.875 ;
      RECT 59.24 2.71 59.245 2.868 ;
      RECT 59.23 2.713 59.24 2.865 ;
      RECT 59.195 2.712 59.23 2.863 ;
      RECT 59.166 2.708 59.195 2.86 ;
      RECT 59.08 2.703 59.166 2.857 ;
      RECT 59.02 2.697 59.08 2.853 ;
      RECT 58.991 2.693 59.02 2.85 ;
      RECT 58.905 2.685 58.991 2.847 ;
      RECT 58.896 2.679 58.905 2.845 ;
      RECT 58.81 2.674 58.896 2.843 ;
      RECT 58.787 2.669 58.81 2.84 ;
      RECT 58.701 2.663 58.787 2.837 ;
      RECT 58.615 2.654 58.701 2.832 ;
      RECT 58.605 2.649 58.615 2.83 ;
      RECT 58.586 2.648 58.605 2.829 ;
      RECT 58.5 2.643 58.586 2.825 ;
      RECT 58.48 2.638 58.5 2.821 ;
      RECT 58.42 2.633 58.48 2.818 ;
      RECT 58.395 2.623 58.42 2.816 ;
      RECT 58.39 2.616 58.395 2.815 ;
      RECT 58.38 2.607 58.39 2.814 ;
      RECT 58.376 2.6 58.38 2.814 ;
      RECT 58.29 2.6 58.376 2.812 ;
      RECT 58.18 2.607 58.195 2.81 ;
      RECT 58.165 2.617 58.17 2.81 ;
      RECT 58.145 2.62 58.165 2.807 ;
      RECT 58.115 2.62 58.145 2.803 ;
      RECT 58.105 2.62 58.115 2.803 ;
      RECT 59.02 3.115 59.28 3.375 ;
      RECT 58.95 3.125 59.28 3.335 ;
      RECT 58.94 3.132 59.28 3.33 ;
      RECT 58.36 3.12 58.62 3.38 ;
      RECT 58.36 3.16 58.725 3.37 ;
      RECT 58.36 3.162 58.73 3.369 ;
      RECT 58.36 3.17 58.735 3.366 ;
      RECT 57.285 2.245 57.385 3.77 ;
      RECT 57.475 3.385 57.525 3.645 ;
      RECT 57.47 2.258 57.475 2.445 ;
      RECT 57.465 3.366 57.475 3.645 ;
      RECT 57.465 2.255 57.47 2.453 ;
      RECT 57.45 2.249 57.465 2.46 ;
      RECT 57.46 3.354 57.465 3.728 ;
      RECT 57.45 3.342 57.46 3.765 ;
      RECT 57.44 2.245 57.45 2.467 ;
      RECT 57.44 3.327 57.45 3.77 ;
      RECT 57.435 2.245 57.44 2.475 ;
      RECT 57.415 3.297 57.44 3.77 ;
      RECT 57.395 2.245 57.435 2.523 ;
      RECT 57.405 3.257 57.415 3.77 ;
      RECT 57.395 3.212 57.405 3.77 ;
      RECT 57.39 2.245 57.395 2.593 ;
      RECT 57.39 3.17 57.395 3.77 ;
      RECT 57.385 2.245 57.39 3.07 ;
      RECT 57.385 3.152 57.39 3.77 ;
      RECT 57.275 2.248 57.285 3.77 ;
      RECT 57.26 2.255 57.275 3.766 ;
      RECT 57.255 2.265 57.26 3.761 ;
      RECT 57.25 2.465 57.255 3.653 ;
      RECT 57.245 2.55 57.25 3.205 ;
      RECT 56.12 7.77 56.41 8 ;
      RECT 56.18 6.29 56.35 8 ;
      RECT 56.13 6.655 56.48 7.005 ;
      RECT 56.12 6.29 56.41 6.52 ;
      RECT 55.715 2.395 55.82 2.965 ;
      RECT 55.715 2.73 56.04 2.96 ;
      RECT 55.715 2.76 56.21 2.93 ;
      RECT 55.715 2.395 55.905 2.96 ;
      RECT 55.13 2.36 55.42 2.59 ;
      RECT 55.13 2.395 55.905 2.565 ;
      RECT 55.19 0.88 55.36 2.59 ;
      RECT 55.13 0.88 55.42 1.11 ;
      RECT 55.13 7.77 55.42 8 ;
      RECT 55.19 6.29 55.36 8 ;
      RECT 55.13 6.29 55.42 6.52 ;
      RECT 55.13 6.325 55.985 6.485 ;
      RECT 55.815 5.92 55.985 6.485 ;
      RECT 55.13 6.32 55.525 6.485 ;
      RECT 55.75 5.92 56.04 6.15 ;
      RECT 55.75 5.95 56.21 6.12 ;
      RECT 54.76 2.73 55.05 2.96 ;
      RECT 54.76 2.76 55.22 2.93 ;
      RECT 54.825 1.655 54.99 2.96 ;
      RECT 53.34 1.625 53.63 1.855 ;
      RECT 53.34 1.655 54.99 1.825 ;
      RECT 53.4 0.885 53.57 1.855 ;
      RECT 53.34 0.885 53.63 1.115 ;
      RECT 53.34 7.765 53.63 7.995 ;
      RECT 53.4 7.025 53.57 7.995 ;
      RECT 53.4 7.12 54.99 7.29 ;
      RECT 54.82 5.92 54.99 7.29 ;
      RECT 53.34 7.025 53.63 7.255 ;
      RECT 54.76 5.92 55.05 6.15 ;
      RECT 54.76 5.95 55.22 6.12 ;
      RECT 51.375 3.43 51.725 3.78 ;
      RECT 51.465 2.025 51.635 3.78 ;
      RECT 53.77 1.965 54.12 2.315 ;
      RECT 51.465 2.025 53.085 2.2 ;
      RECT 51.465 2.025 54.12 2.195 ;
      RECT 53.795 6.655 54.12 6.98 ;
      RECT 49.225 6.615 49.575 6.965 ;
      RECT 53.77 6.655 54.12 6.885 ;
      RECT 49.01 6.655 49.575 6.885 ;
      RECT 48.84 6.685 54.12 6.855 ;
      RECT 52.995 2.365 53.315 2.685 ;
      RECT 52.965 2.365 53.315 2.595 ;
      RECT 52.795 2.395 53.315 2.565 ;
      RECT 52.995 6.225 53.315 6.545 ;
      RECT 52.965 6.285 53.315 6.515 ;
      RECT 52.795 6.315 53.315 6.485 ;
      RECT 48.775 3.665 48.815 3.925 ;
      RECT 48.815 3.645 48.82 3.655 ;
      RECT 50.145 2.89 50.155 3.111 ;
      RECT 50.075 2.885 50.145 3.236 ;
      RECT 50.065 2.885 50.075 3.363 ;
      RECT 50.04 2.885 50.065 3.41 ;
      RECT 50.015 2.885 50.04 3.488 ;
      RECT 49.995 2.885 50.015 3.558 ;
      RECT 49.97 2.885 49.995 3.598 ;
      RECT 49.96 2.885 49.97 3.618 ;
      RECT 49.95 2.887 49.96 3.626 ;
      RECT 49.945 2.892 49.95 3.083 ;
      RECT 49.945 3.092 49.95 3.627 ;
      RECT 49.94 3.137 49.945 3.628 ;
      RECT 49.93 3.202 49.94 3.629 ;
      RECT 49.92 3.297 49.93 3.631 ;
      RECT 49.915 3.35 49.92 3.633 ;
      RECT 49.91 3.37 49.915 3.634 ;
      RECT 49.855 3.395 49.91 3.64 ;
      RECT 49.815 3.43 49.855 3.649 ;
      RECT 49.805 3.447 49.815 3.654 ;
      RECT 49.796 3.453 49.805 3.656 ;
      RECT 49.71 3.491 49.796 3.667 ;
      RECT 49.705 3.53 49.71 3.677 ;
      RECT 49.63 3.537 49.705 3.687 ;
      RECT 49.61 3.547 49.63 3.698 ;
      RECT 49.58 3.554 49.61 3.706 ;
      RECT 49.555 3.561 49.58 3.713 ;
      RECT 49.531 3.567 49.555 3.718 ;
      RECT 49.445 3.58 49.531 3.73 ;
      RECT 49.367 3.587 49.445 3.748 ;
      RECT 49.281 3.582 49.367 3.766 ;
      RECT 49.195 3.577 49.281 3.786 ;
      RECT 49.115 3.571 49.195 3.803 ;
      RECT 49.05 3.567 49.115 3.832 ;
      RECT 49.045 3.281 49.05 3.305 ;
      RECT 49.035 3.557 49.05 3.86 ;
      RECT 49.04 3.275 49.045 3.345 ;
      RECT 49.035 3.269 49.04 3.415 ;
      RECT 49.03 3.263 49.035 3.493 ;
      RECT 49.03 3.54 49.035 3.925 ;
      RECT 49.022 3.26 49.03 3.925 ;
      RECT 48.936 3.258 49.022 3.925 ;
      RECT 48.85 3.256 48.936 3.925 ;
      RECT 48.84 3.257 48.85 3.925 ;
      RECT 48.835 3.262 48.84 3.925 ;
      RECT 48.825 3.275 48.835 3.925 ;
      RECT 48.82 3.297 48.825 3.925 ;
      RECT 48.815 3.657 48.82 3.925 ;
      RECT 49.445 3.125 49.45 3.345 ;
      RECT 49.95 2.16 49.985 2.42 ;
      RECT 49.935 2.16 49.95 2.428 ;
      RECT 49.906 2.16 49.935 2.45 ;
      RECT 49.82 2.16 49.906 2.51 ;
      RECT 49.8 2.16 49.82 2.575 ;
      RECT 49.74 2.16 49.8 2.74 ;
      RECT 49.735 2.16 49.74 2.888 ;
      RECT 49.73 2.16 49.735 2.9 ;
      RECT 49.725 2.16 49.73 2.926 ;
      RECT 49.695 2.346 49.725 3.006 ;
      RECT 49.69 2.394 49.695 3.095 ;
      RECT 49.685 2.408 49.69 3.11 ;
      RECT 49.68 2.427 49.685 3.14 ;
      RECT 49.675 2.442 49.68 3.156 ;
      RECT 49.67 2.457 49.675 3.178 ;
      RECT 49.665 2.477 49.67 3.2 ;
      RECT 49.655 2.497 49.665 3.233 ;
      RECT 49.64 2.539 49.655 3.295 ;
      RECT 49.635 2.57 49.64 3.335 ;
      RECT 49.63 2.582 49.635 3.34 ;
      RECT 49.625 2.594 49.63 3.345 ;
      RECT 49.62 2.607 49.625 3.345 ;
      RECT 49.615 2.625 49.62 3.345 ;
      RECT 49.61 2.645 49.615 3.345 ;
      RECT 49.605 2.657 49.61 3.345 ;
      RECT 49.6 2.67 49.605 3.345 ;
      RECT 49.58 2.705 49.6 3.345 ;
      RECT 49.53 2.807 49.58 3.345 ;
      RECT 49.525 2.892 49.53 3.345 ;
      RECT 49.52 2.9 49.525 3.345 ;
      RECT 49.515 2.917 49.52 3.345 ;
      RECT 49.51 2.932 49.515 3.345 ;
      RECT 49.475 2.997 49.51 3.345 ;
      RECT 49.46 3.062 49.475 3.345 ;
      RECT 49.455 3.092 49.46 3.345 ;
      RECT 49.45 3.117 49.455 3.345 ;
      RECT 49.435 3.127 49.445 3.345 ;
      RECT 49.42 3.14 49.435 3.338 ;
      RECT 49.165 2.73 49.235 2.94 ;
      RECT 48.955 2.707 48.96 2.9 ;
      RECT 46.41 2.635 46.67 2.895 ;
      RECT 49.245 2.917 49.25 2.92 ;
      RECT 49.235 2.735 49.245 2.935 ;
      RECT 49.136 2.728 49.165 2.94 ;
      RECT 49.05 2.72 49.136 2.94 ;
      RECT 49.035 2.714 49.05 2.938 ;
      RECT 49.015 2.713 49.035 2.925 ;
      RECT 49.01 2.712 49.015 2.908 ;
      RECT 48.96 2.709 49.01 2.903 ;
      RECT 48.93 2.706 48.955 2.898 ;
      RECT 48.91 2.704 48.93 2.893 ;
      RECT 48.895 2.702 48.91 2.89 ;
      RECT 48.865 2.7 48.895 2.888 ;
      RECT 48.8 2.696 48.865 2.88 ;
      RECT 48.77 2.691 48.8 2.875 ;
      RECT 48.75 2.689 48.77 2.873 ;
      RECT 48.72 2.686 48.75 2.868 ;
      RECT 48.66 2.682 48.72 2.86 ;
      RECT 48.655 2.679 48.66 2.855 ;
      RECT 48.585 2.677 48.655 2.85 ;
      RECT 48.556 2.673 48.585 2.843 ;
      RECT 48.47 2.668 48.556 2.835 ;
      RECT 48.436 2.663 48.47 2.827 ;
      RECT 48.35 2.655 48.436 2.819 ;
      RECT 48.311 2.648 48.35 2.811 ;
      RECT 48.225 2.643 48.311 2.803 ;
      RECT 48.16 2.637 48.225 2.793 ;
      RECT 48.14 2.632 48.16 2.788 ;
      RECT 48.131 2.629 48.14 2.787 ;
      RECT 48.045 2.625 48.131 2.781 ;
      RECT 48.005 2.621 48.045 2.773 ;
      RECT 47.985 2.617 48.005 2.771 ;
      RECT 47.925 2.617 47.985 2.768 ;
      RECT 47.905 2.62 47.925 2.766 ;
      RECT 47.884 2.62 47.905 2.766 ;
      RECT 47.798 2.622 47.884 2.77 ;
      RECT 47.712 2.624 47.798 2.776 ;
      RECT 47.626 2.626 47.712 2.783 ;
      RECT 47.54 2.629 47.626 2.789 ;
      RECT 47.506 2.63 47.54 2.794 ;
      RECT 47.42 2.633 47.506 2.799 ;
      RECT 47.391 2.64 47.42 2.804 ;
      RECT 47.305 2.64 47.391 2.809 ;
      RECT 47.272 2.64 47.305 2.814 ;
      RECT 47.186 2.642 47.272 2.819 ;
      RECT 47.1 2.644 47.186 2.826 ;
      RECT 47.036 2.646 47.1 2.832 ;
      RECT 46.95 2.648 47.036 2.838 ;
      RECT 46.947 2.65 46.95 2.841 ;
      RECT 46.861 2.651 46.947 2.845 ;
      RECT 46.775 2.654 46.861 2.852 ;
      RECT 46.756 2.656 46.775 2.856 ;
      RECT 46.67 2.658 46.756 2.861 ;
      RECT 46.4 2.67 46.41 2.865 ;
      RECT 48.58 7.765 48.87 7.995 ;
      RECT 48.64 7.025 48.81 7.995 ;
      RECT 48.53 7.055 48.905 7.425 ;
      RECT 48.58 7.025 48.87 7.425 ;
      RECT 48.635 2.25 48.82 2.46 ;
      RECT 48.63 2.251 48.825 2.458 ;
      RECT 48.625 2.256 48.835 2.453 ;
      RECT 48.62 2.232 48.625 2.45 ;
      RECT 48.59 2.229 48.62 2.443 ;
      RECT 48.585 2.225 48.59 2.434 ;
      RECT 48.55 2.256 48.835 2.429 ;
      RECT 48.325 2.165 48.585 2.425 ;
      RECT 48.625 2.234 48.63 2.453 ;
      RECT 48.63 2.235 48.635 2.458 ;
      RECT 48.325 2.247 48.705 2.425 ;
      RECT 48.325 2.245 48.69 2.425 ;
      RECT 48.325 2.24 48.68 2.425 ;
      RECT 48.28 3.155 48.33 3.44 ;
      RECT 48.225 3.125 48.23 3.44 ;
      RECT 48.195 3.105 48.2 3.44 ;
      RECT 48.345 3.155 48.405 3.415 ;
      RECT 48.34 3.155 48.345 3.423 ;
      RECT 48.33 3.155 48.34 3.435 ;
      RECT 48.245 3.145 48.28 3.44 ;
      RECT 48.24 3.132 48.245 3.44 ;
      RECT 48.23 3.127 48.24 3.44 ;
      RECT 48.21 3.117 48.225 3.44 ;
      RECT 48.2 3.11 48.21 3.44 ;
      RECT 48.19 3.102 48.195 3.44 ;
      RECT 48.16 3.092 48.19 3.44 ;
      RECT 48.145 3.08 48.16 3.44 ;
      RECT 48.13 3.07 48.145 3.435 ;
      RECT 48.11 3.06 48.13 3.41 ;
      RECT 48.1 3.052 48.11 3.387 ;
      RECT 48.07 3.035 48.1 3.377 ;
      RECT 48.065 3.012 48.07 3.368 ;
      RECT 48.06 2.999 48.065 3.366 ;
      RECT 48.045 2.975 48.06 3.36 ;
      RECT 48.04 2.951 48.045 3.354 ;
      RECT 48.03 2.94 48.04 3.349 ;
      RECT 48.025 2.93 48.03 3.345 ;
      RECT 48.02 2.922 48.025 3.342 ;
      RECT 48.01 2.917 48.02 3.338 ;
      RECT 48.005 2.912 48.01 3.334 ;
      RECT 47.92 2.91 48.005 3.309 ;
      RECT 47.89 2.91 47.92 3.275 ;
      RECT 47.875 2.91 47.89 3.258 ;
      RECT 47.82 2.91 47.875 3.203 ;
      RECT 47.815 2.915 47.82 3.152 ;
      RECT 47.805 2.92 47.815 3.142 ;
      RECT 47.8 2.93 47.805 3.128 ;
      RECT 47.75 3.67 48.01 3.93 ;
      RECT 47.67 3.685 48.01 3.906 ;
      RECT 47.65 3.685 48.01 3.901 ;
      RECT 47.626 3.685 48.01 3.899 ;
      RECT 47.54 3.685 48.01 3.894 ;
      RECT 47.39 3.625 47.65 3.89 ;
      RECT 47.345 3.685 48.01 3.885 ;
      RECT 47.34 3.692 48.01 3.88 ;
      RECT 47.355 3.68 47.67 3.89 ;
      RECT 47.245 2.115 47.505 2.375 ;
      RECT 47.245 2.172 47.51 2.368 ;
      RECT 47.245 2.202 47.515 2.3 ;
      RECT 47.305 2.633 47.42 2.635 ;
      RECT 47.391 2.63 47.42 2.635 ;
      RECT 46.415 3.634 46.44 3.874 ;
      RECT 46.4 3.637 46.49 3.868 ;
      RECT 46.395 3.642 46.576 3.863 ;
      RECT 46.39 3.65 46.64 3.861 ;
      RECT 46.39 3.65 46.65 3.86 ;
      RECT 46.385 3.657 46.66 3.853 ;
      RECT 46.385 3.657 46.746 3.842 ;
      RECT 46.38 3.692 46.746 3.838 ;
      RECT 46.38 3.692 46.755 3.827 ;
      RECT 46.66 3.565 46.92 3.825 ;
      RECT 46.37 3.742 46.92 3.823 ;
      RECT 46.64 3.61 46.66 3.858 ;
      RECT 46.576 3.613 46.64 3.862 ;
      RECT 46.49 3.618 46.576 3.867 ;
      RECT 46.42 3.629 46.92 3.825 ;
      RECT 46.44 3.623 46.49 3.872 ;
      RECT 46.565 2.1 46.575 2.362 ;
      RECT 46.555 2.157 46.565 2.365 ;
      RECT 46.53 2.162 46.555 2.371 ;
      RECT 46.505 2.166 46.53 2.383 ;
      RECT 46.495 2.169 46.505 2.393 ;
      RECT 46.49 2.17 46.495 2.398 ;
      RECT 46.485 2.171 46.49 2.403 ;
      RECT 46.48 2.172 46.485 2.405 ;
      RECT 46.455 2.175 46.48 2.408 ;
      RECT 46.425 2.181 46.455 2.411 ;
      RECT 46.36 2.192 46.425 2.414 ;
      RECT 46.315 2.2 46.36 2.418 ;
      RECT 46.3 2.2 46.315 2.426 ;
      RECT 46.295 2.201 46.3 2.433 ;
      RECT 46.29 2.203 46.295 2.436 ;
      RECT 46.285 2.207 46.29 2.439 ;
      RECT 46.275 2.215 46.285 2.443 ;
      RECT 46.27 2.228 46.275 2.448 ;
      RECT 46.265 2.236 46.27 2.45 ;
      RECT 46.26 2.242 46.265 2.45 ;
      RECT 46.255 2.246 46.26 2.453 ;
      RECT 46.25 2.248 46.255 2.456 ;
      RECT 46.245 2.251 46.25 2.459 ;
      RECT 46.235 2.256 46.245 2.463 ;
      RECT 46.23 2.262 46.235 2.468 ;
      RECT 46.22 2.268 46.23 2.472 ;
      RECT 46.205 2.275 46.22 2.478 ;
      RECT 46.176 2.289 46.205 2.488 ;
      RECT 46.09 2.324 46.176 2.52 ;
      RECT 46.07 2.357 46.09 2.549 ;
      RECT 46.05 2.37 46.07 2.56 ;
      RECT 46.03 2.382 46.05 2.571 ;
      RECT 45.98 2.404 46.03 2.591 ;
      RECT 45.965 2.422 45.98 2.608 ;
      RECT 45.96 2.428 45.965 2.611 ;
      RECT 45.955 2.432 45.96 2.614 ;
      RECT 45.95 2.436 45.955 2.618 ;
      RECT 45.945 2.438 45.95 2.621 ;
      RECT 45.935 2.445 45.945 2.624 ;
      RECT 45.93 2.45 45.935 2.628 ;
      RECT 45.925 2.452 45.93 2.631 ;
      RECT 45.92 2.456 45.925 2.634 ;
      RECT 45.915 2.458 45.92 2.638 ;
      RECT 45.9 2.463 45.915 2.643 ;
      RECT 45.895 2.468 45.9 2.646 ;
      RECT 45.89 2.476 45.895 2.649 ;
      RECT 45.885 2.478 45.89 2.652 ;
      RECT 45.88 2.48 45.885 2.655 ;
      RECT 45.87 2.482 45.88 2.661 ;
      RECT 45.835 2.496 45.87 2.673 ;
      RECT 45.825 2.511 45.835 2.683 ;
      RECT 45.75 2.54 45.825 2.707 ;
      RECT 45.745 2.565 45.75 2.73 ;
      RECT 45.73 2.569 45.745 2.736 ;
      RECT 45.72 2.577 45.73 2.741 ;
      RECT 45.69 2.59 45.72 2.745 ;
      RECT 45.68 2.605 45.69 2.75 ;
      RECT 45.67 2.61 45.68 2.753 ;
      RECT 45.665 2.612 45.67 2.755 ;
      RECT 45.65 2.615 45.665 2.758 ;
      RECT 45.645 2.617 45.65 2.761 ;
      RECT 45.625 2.622 45.645 2.765 ;
      RECT 45.595 2.627 45.625 2.773 ;
      RECT 45.57 2.634 45.595 2.781 ;
      RECT 45.565 2.639 45.57 2.786 ;
      RECT 45.535 2.642 45.565 2.79 ;
      RECT 45.495 2.645 45.535 2.8 ;
      RECT 45.46 2.642 45.495 2.812 ;
      RECT 45.45 2.638 45.46 2.819 ;
      RECT 45.425 2.634 45.45 2.825 ;
      RECT 45.42 2.63 45.425 2.83 ;
      RECT 45.38 2.627 45.42 2.83 ;
      RECT 45.365 2.612 45.38 2.831 ;
      RECT 45.342 2.6 45.365 2.831 ;
      RECT 45.256 2.6 45.342 2.832 ;
      RECT 45.17 2.6 45.256 2.834 ;
      RECT 45.15 2.6 45.17 2.831 ;
      RECT 45.145 2.605 45.15 2.826 ;
      RECT 45.14 2.61 45.145 2.824 ;
      RECT 45.13 2.62 45.14 2.822 ;
      RECT 45.125 2.626 45.13 2.815 ;
      RECT 45.12 2.628 45.125 2.8 ;
      RECT 45.115 2.632 45.12 2.79 ;
      RECT 46.575 2.1 46.825 2.36 ;
      RECT 44.3 3.635 44.56 3.895 ;
      RECT 46.595 3.125 46.6 3.335 ;
      RECT 46.6 3.13 46.61 3.33 ;
      RECT 46.55 3.125 46.595 3.35 ;
      RECT 46.54 3.125 46.55 3.37 ;
      RECT 46.521 3.125 46.54 3.375 ;
      RECT 46.435 3.125 46.521 3.372 ;
      RECT 46.405 3.127 46.435 3.37 ;
      RECT 46.35 3.137 46.405 3.368 ;
      RECT 46.285 3.151 46.35 3.366 ;
      RECT 46.28 3.159 46.285 3.365 ;
      RECT 46.265 3.162 46.28 3.363 ;
      RECT 46.2 3.172 46.265 3.359 ;
      RECT 46.152 3.186 46.2 3.36 ;
      RECT 46.066 3.203 46.152 3.374 ;
      RECT 45.98 3.224 46.066 3.391 ;
      RECT 45.96 3.237 45.98 3.401 ;
      RECT 45.915 3.245 45.96 3.408 ;
      RECT 45.88 3.253 45.915 3.416 ;
      RECT 45.846 3.261 45.88 3.424 ;
      RECT 45.76 3.275 45.846 3.436 ;
      RECT 45.725 3.292 45.76 3.448 ;
      RECT 45.716 3.301 45.725 3.452 ;
      RECT 45.63 3.319 45.716 3.469 ;
      RECT 45.571 3.346 45.63 3.496 ;
      RECT 45.485 3.373 45.571 3.524 ;
      RECT 45.465 3.395 45.485 3.544 ;
      RECT 45.405 3.41 45.465 3.56 ;
      RECT 45.395 3.422 45.405 3.573 ;
      RECT 45.39 3.427 45.395 3.576 ;
      RECT 45.38 3.43 45.39 3.579 ;
      RECT 45.375 3.432 45.38 3.582 ;
      RECT 45.345 3.44 45.375 3.589 ;
      RECT 45.33 3.447 45.345 3.597 ;
      RECT 45.32 3.452 45.33 3.601 ;
      RECT 45.315 3.455 45.32 3.604 ;
      RECT 45.305 3.457 45.315 3.607 ;
      RECT 45.27 3.467 45.305 3.616 ;
      RECT 45.195 3.49 45.27 3.638 ;
      RECT 45.175 3.508 45.195 3.656 ;
      RECT 45.145 3.515 45.175 3.666 ;
      RECT 45.125 3.523 45.145 3.676 ;
      RECT 45.115 3.529 45.125 3.683 ;
      RECT 45.096 3.534 45.115 3.689 ;
      RECT 45.01 3.554 45.096 3.709 ;
      RECT 44.995 3.574 45.01 3.728 ;
      RECT 44.95 3.586 44.995 3.739 ;
      RECT 44.885 3.607 44.95 3.762 ;
      RECT 44.845 3.627 44.885 3.783 ;
      RECT 44.835 3.637 44.845 3.793 ;
      RECT 44.785 3.649 44.835 3.804 ;
      RECT 44.765 3.665 44.785 3.816 ;
      RECT 44.735 3.675 44.765 3.822 ;
      RECT 44.725 3.68 44.735 3.824 ;
      RECT 44.656 3.681 44.725 3.83 ;
      RECT 44.57 3.683 44.656 3.84 ;
      RECT 44.56 3.684 44.57 3.845 ;
      RECT 45.83 3.71 46.02 3.92 ;
      RECT 45.82 3.715 46.03 3.913 ;
      RECT 45.805 3.715 46.03 3.878 ;
      RECT 45.725 3.6 45.985 3.86 ;
      RECT 44.64 3.13 44.825 3.425 ;
      RECT 44.63 3.13 44.825 3.423 ;
      RECT 44.615 3.13 44.83 3.418 ;
      RECT 44.615 3.13 44.835 3.415 ;
      RECT 44.61 3.13 44.835 3.413 ;
      RECT 44.605 3.385 44.835 3.403 ;
      RECT 44.61 3.13 44.87 3.39 ;
      RECT 44.57 2.165 44.83 2.425 ;
      RECT 44.38 2.09 44.466 2.423 ;
      RECT 44.355 2.094 44.51 2.419 ;
      RECT 44.466 2.086 44.51 2.419 ;
      RECT 44.466 2.087 44.515 2.418 ;
      RECT 44.38 2.092 44.53 2.417 ;
      RECT 44.355 2.1 44.57 2.416 ;
      RECT 44.35 2.095 44.53 2.411 ;
      RECT 44.34 2.11 44.57 2.318 ;
      RECT 44.34 2.162 44.77 2.318 ;
      RECT 44.34 2.155 44.75 2.318 ;
      RECT 44.34 2.142 44.72 2.318 ;
      RECT 44.34 2.13 44.66 2.318 ;
      RECT 44.34 2.115 44.635 2.318 ;
      RECT 43.54 2.745 43.675 3.04 ;
      RECT 43.8 2.768 43.805 2.955 ;
      RECT 44.52 2.665 44.665 2.9 ;
      RECT 44.68 2.665 44.685 2.89 ;
      RECT 44.715 2.676 44.72 2.87 ;
      RECT 44.71 2.668 44.715 2.875 ;
      RECT 44.69 2.665 44.71 2.88 ;
      RECT 44.685 2.665 44.69 2.888 ;
      RECT 44.675 2.665 44.68 2.893 ;
      RECT 44.665 2.665 44.675 2.898 ;
      RECT 44.495 2.667 44.52 2.9 ;
      RECT 44.445 2.674 44.495 2.9 ;
      RECT 44.44 2.679 44.445 2.9 ;
      RECT 44.401 2.684 44.44 2.901 ;
      RECT 44.315 2.696 44.401 2.902 ;
      RECT 44.306 2.706 44.315 2.902 ;
      RECT 44.22 2.715 44.306 2.904 ;
      RECT 44.196 2.725 44.22 2.906 ;
      RECT 44.11 2.736 44.196 2.907 ;
      RECT 44.08 2.747 44.11 2.909 ;
      RECT 44.05 2.752 44.08 2.911 ;
      RECT 44.025 2.758 44.05 2.914 ;
      RECT 44.01 2.763 44.025 2.915 ;
      RECT 43.965 2.769 44.01 2.915 ;
      RECT 43.96 2.774 43.965 2.916 ;
      RECT 43.94 2.774 43.96 2.918 ;
      RECT 43.92 2.772 43.94 2.923 ;
      RECT 43.885 2.771 43.92 2.93 ;
      RECT 43.855 2.77 43.885 2.94 ;
      RECT 43.805 2.769 43.855 2.95 ;
      RECT 43.715 2.766 43.8 3.04 ;
      RECT 43.69 2.76 43.715 3.04 ;
      RECT 43.675 2.75 43.69 3.04 ;
      RECT 43.49 2.745 43.54 2.96 ;
      RECT 43.48 2.75 43.49 2.95 ;
      RECT 43.72 3.225 43.98 3.485 ;
      RECT 43.72 3.225 44.01 3.378 ;
      RECT 43.72 3.225 44.045 3.363 ;
      RECT 43.975 3.145 44.165 3.355 ;
      RECT 43.965 3.15 44.175 3.348 ;
      RECT 43.93 3.22 44.175 3.348 ;
      RECT 43.96 3.162 43.98 3.485 ;
      RECT 43.945 3.21 44.175 3.348 ;
      RECT 43.95 3.182 43.98 3.485 ;
      RECT 43.03 2.25 43.1 3.355 ;
      RECT 43.765 2.355 44.025 2.615 ;
      RECT 43.345 2.401 43.36 2.61 ;
      RECT 43.681 2.414 43.765 2.565 ;
      RECT 43.595 2.411 43.681 2.565 ;
      RECT 43.556 2.409 43.595 2.565 ;
      RECT 43.47 2.407 43.556 2.565 ;
      RECT 43.41 2.405 43.47 2.576 ;
      RECT 43.375 2.403 43.41 2.594 ;
      RECT 43.36 2.401 43.375 2.605 ;
      RECT 43.33 2.401 43.345 2.618 ;
      RECT 43.32 2.401 43.33 2.623 ;
      RECT 43.295 2.4 43.32 2.628 ;
      RECT 43.28 2.395 43.295 2.634 ;
      RECT 43.275 2.388 43.28 2.639 ;
      RECT 43.25 2.379 43.275 2.645 ;
      RECT 43.205 2.358 43.25 2.658 ;
      RECT 43.195 2.342 43.205 2.668 ;
      RECT 43.18 2.335 43.195 2.678 ;
      RECT 43.17 2.328 43.18 2.695 ;
      RECT 43.165 2.325 43.17 2.725 ;
      RECT 43.16 2.323 43.165 2.755 ;
      RECT 43.155 2.321 43.16 2.792 ;
      RECT 43.14 2.317 43.155 2.859 ;
      RECT 43.14 3.15 43.15 3.35 ;
      RECT 43.135 2.313 43.14 2.985 ;
      RECT 43.135 3.137 43.14 3.355 ;
      RECT 43.13 2.311 43.135 3.07 ;
      RECT 43.13 3.127 43.135 3.355 ;
      RECT 43.115 2.282 43.13 3.355 ;
      RECT 43.1 2.255 43.115 3.355 ;
      RECT 43.025 2.25 43.03 2.605 ;
      RECT 43.025 2.66 43.03 3.355 ;
      RECT 43.01 2.25 43.025 2.583 ;
      RECT 43.02 2.682 43.025 3.355 ;
      RECT 43.01 2.722 43.02 3.355 ;
      RECT 42.975 2.25 43.01 2.525 ;
      RECT 43.005 2.757 43.01 3.355 ;
      RECT 42.99 2.812 43.005 3.355 ;
      RECT 42.985 2.877 42.99 3.355 ;
      RECT 42.97 2.925 42.985 3.355 ;
      RECT 42.945 2.25 42.975 2.48 ;
      RECT 42.965 2.98 42.97 3.355 ;
      RECT 42.95 3.04 42.965 3.355 ;
      RECT 42.945 3.088 42.95 3.353 ;
      RECT 42.94 2.25 42.945 2.473 ;
      RECT 42.94 3.12 42.945 3.348 ;
      RECT 42.915 2.25 42.94 2.465 ;
      RECT 42.905 2.255 42.915 2.455 ;
      RECT 43.12 3.53 43.14 3.77 ;
      RECT 42.35 3.46 42.355 3.67 ;
      RECT 43.63 3.533 43.64 3.728 ;
      RECT 43.625 3.523 43.63 3.731 ;
      RECT 43.545 3.52 43.625 3.754 ;
      RECT 43.541 3.52 43.545 3.776 ;
      RECT 43.455 3.52 43.541 3.786 ;
      RECT 43.44 3.52 43.455 3.794 ;
      RECT 43.411 3.521 43.44 3.792 ;
      RECT 43.325 3.526 43.411 3.788 ;
      RECT 43.312 3.53 43.325 3.784 ;
      RECT 43.226 3.53 43.312 3.78 ;
      RECT 43.14 3.53 43.226 3.774 ;
      RECT 43.056 3.53 43.12 3.768 ;
      RECT 42.97 3.53 43.056 3.763 ;
      RECT 42.95 3.53 42.97 3.759 ;
      RECT 42.89 3.525 42.95 3.756 ;
      RECT 42.862 3.519 42.89 3.753 ;
      RECT 42.776 3.514 42.862 3.749 ;
      RECT 42.69 3.508 42.776 3.743 ;
      RECT 42.615 3.49 42.69 3.738 ;
      RECT 42.58 3.467 42.615 3.734 ;
      RECT 42.57 3.457 42.58 3.733 ;
      RECT 42.515 3.455 42.57 3.732 ;
      RECT 42.44 3.455 42.515 3.728 ;
      RECT 42.43 3.455 42.44 3.723 ;
      RECT 42.415 3.455 42.43 3.715 ;
      RECT 42.365 3.457 42.415 3.693 ;
      RECT 42.355 3.46 42.365 3.673 ;
      RECT 42.345 3.465 42.35 3.668 ;
      RECT 42.34 3.47 42.345 3.663 ;
      RECT 42.465 2.635 42.725 2.895 ;
      RECT 42.465 2.65 42.745 2.86 ;
      RECT 42.465 2.655 42.755 2.855 ;
      RECT 40.45 2.115 40.71 2.375 ;
      RECT 40.44 2.145 40.71 2.355 ;
      RECT 42.36 2.06 42.62 2.32 ;
      RECT 42.355 2.135 42.36 2.321 ;
      RECT 42.33 2.14 42.355 2.323 ;
      RECT 42.315 2.147 42.33 2.326 ;
      RECT 42.255 2.165 42.315 2.331 ;
      RECT 42.225 2.185 42.255 2.338 ;
      RECT 42.2 2.193 42.225 2.343 ;
      RECT 42.175 2.201 42.2 2.345 ;
      RECT 42.157 2.205 42.175 2.344 ;
      RECT 42.071 2.203 42.157 2.344 ;
      RECT 41.985 2.201 42.071 2.344 ;
      RECT 41.899 2.199 41.985 2.343 ;
      RECT 41.813 2.197 41.899 2.343 ;
      RECT 41.727 2.195 41.813 2.343 ;
      RECT 41.641 2.193 41.727 2.343 ;
      RECT 41.555 2.191 41.641 2.342 ;
      RECT 41.537 2.19 41.555 2.342 ;
      RECT 41.451 2.189 41.537 2.342 ;
      RECT 41.365 2.187 41.451 2.342 ;
      RECT 41.279 2.186 41.365 2.341 ;
      RECT 41.193 2.185 41.279 2.341 ;
      RECT 41.107 2.183 41.193 2.341 ;
      RECT 41.021 2.182 41.107 2.341 ;
      RECT 40.935 2.18 41.021 2.34 ;
      RECT 40.911 2.178 40.935 2.34 ;
      RECT 40.825 2.171 40.911 2.34 ;
      RECT 40.796 2.163 40.825 2.34 ;
      RECT 40.71 2.155 40.796 2.34 ;
      RECT 40.43 2.152 40.44 2.35 ;
      RECT 41.935 3.115 41.94 3.465 ;
      RECT 41.705 3.205 41.845 3.465 ;
      RECT 42.18 2.89 42.225 3.1 ;
      RECT 42.235 2.901 42.245 3.095 ;
      RECT 42.225 2.893 42.235 3.1 ;
      RECT 42.16 2.89 42.18 3.105 ;
      RECT 42.13 2.89 42.16 3.128 ;
      RECT 42.12 2.89 42.13 3.153 ;
      RECT 42.115 2.89 42.12 3.163 ;
      RECT 42.06 2.89 42.115 3.203 ;
      RECT 42.055 2.89 42.06 3.243 ;
      RECT 42.05 2.892 42.055 3.248 ;
      RECT 42.035 2.902 42.05 3.259 ;
      RECT 41.99 2.96 42.035 3.295 ;
      RECT 41.98 3.015 41.99 3.329 ;
      RECT 41.965 3.042 41.98 3.345 ;
      RECT 41.955 3.069 41.965 3.465 ;
      RECT 41.94 3.092 41.955 3.465 ;
      RECT 41.93 3.132 41.935 3.465 ;
      RECT 41.925 3.142 41.93 3.465 ;
      RECT 41.92 3.157 41.925 3.465 ;
      RECT 41.91 3.162 41.92 3.465 ;
      RECT 41.845 3.185 41.91 3.465 ;
      RECT 41.345 2.68 41.535 2.89 ;
      RECT 39.92 2.605 40.18 2.865 ;
      RECT 40.27 2.6 40.365 2.81 ;
      RECT 40.245 2.615 40.255 2.81 ;
      RECT 41.535 2.687 41.545 2.885 ;
      RECT 41.335 2.687 41.345 2.885 ;
      RECT 41.32 2.702 41.335 2.875 ;
      RECT 41.315 2.71 41.32 2.868 ;
      RECT 41.305 2.713 41.315 2.865 ;
      RECT 41.27 2.712 41.305 2.863 ;
      RECT 41.241 2.708 41.27 2.86 ;
      RECT 41.155 2.703 41.241 2.857 ;
      RECT 41.095 2.697 41.155 2.853 ;
      RECT 41.066 2.693 41.095 2.85 ;
      RECT 40.98 2.685 41.066 2.847 ;
      RECT 40.971 2.679 40.98 2.845 ;
      RECT 40.885 2.674 40.971 2.843 ;
      RECT 40.862 2.669 40.885 2.84 ;
      RECT 40.776 2.663 40.862 2.837 ;
      RECT 40.69 2.654 40.776 2.832 ;
      RECT 40.68 2.649 40.69 2.83 ;
      RECT 40.661 2.648 40.68 2.829 ;
      RECT 40.575 2.643 40.661 2.825 ;
      RECT 40.555 2.638 40.575 2.821 ;
      RECT 40.495 2.633 40.555 2.818 ;
      RECT 40.47 2.623 40.495 2.816 ;
      RECT 40.465 2.616 40.47 2.815 ;
      RECT 40.455 2.607 40.465 2.814 ;
      RECT 40.451 2.6 40.455 2.814 ;
      RECT 40.365 2.6 40.451 2.812 ;
      RECT 40.255 2.607 40.27 2.81 ;
      RECT 40.24 2.617 40.245 2.81 ;
      RECT 40.22 2.62 40.24 2.807 ;
      RECT 40.19 2.62 40.22 2.803 ;
      RECT 40.18 2.62 40.19 2.803 ;
      RECT 41.095 3.115 41.355 3.375 ;
      RECT 41.025 3.125 41.355 3.335 ;
      RECT 41.015 3.132 41.355 3.33 ;
      RECT 40.435 3.12 40.695 3.38 ;
      RECT 40.435 3.16 40.8 3.37 ;
      RECT 40.435 3.162 40.805 3.369 ;
      RECT 40.435 3.17 40.81 3.366 ;
      RECT 39.36 2.245 39.46 3.77 ;
      RECT 39.55 3.385 39.6 3.645 ;
      RECT 39.545 2.258 39.55 2.445 ;
      RECT 39.54 3.366 39.55 3.645 ;
      RECT 39.54 2.255 39.545 2.453 ;
      RECT 39.525 2.249 39.54 2.46 ;
      RECT 39.535 3.354 39.54 3.728 ;
      RECT 39.525 3.342 39.535 3.765 ;
      RECT 39.515 2.245 39.525 2.467 ;
      RECT 39.515 3.327 39.525 3.77 ;
      RECT 39.51 2.245 39.515 2.475 ;
      RECT 39.49 3.297 39.515 3.77 ;
      RECT 39.47 2.245 39.51 2.523 ;
      RECT 39.48 3.257 39.49 3.77 ;
      RECT 39.47 3.212 39.48 3.77 ;
      RECT 39.465 2.245 39.47 2.593 ;
      RECT 39.465 3.17 39.47 3.77 ;
      RECT 39.46 2.245 39.465 3.07 ;
      RECT 39.46 3.152 39.465 3.77 ;
      RECT 39.35 2.248 39.36 3.77 ;
      RECT 39.335 2.255 39.35 3.766 ;
      RECT 39.33 2.265 39.335 3.761 ;
      RECT 39.325 2.465 39.33 3.653 ;
      RECT 39.32 2.55 39.325 3.205 ;
      RECT 38.195 7.77 38.485 8 ;
      RECT 38.255 6.29 38.425 8 ;
      RECT 38.245 6.66 38.6 7.015 ;
      RECT 38.195 6.29 38.485 6.52 ;
      RECT 37.79 2.395 37.895 2.965 ;
      RECT 37.79 2.73 38.115 2.96 ;
      RECT 37.79 2.76 38.285 2.93 ;
      RECT 37.79 2.395 37.98 2.96 ;
      RECT 37.205 2.36 37.495 2.59 ;
      RECT 37.205 2.395 37.98 2.565 ;
      RECT 37.265 0.88 37.435 2.59 ;
      RECT 37.205 0.88 37.495 1.11 ;
      RECT 37.205 7.77 37.495 8 ;
      RECT 37.265 6.29 37.435 8 ;
      RECT 37.205 6.29 37.495 6.52 ;
      RECT 37.205 6.325 38.06 6.485 ;
      RECT 37.89 5.92 38.06 6.485 ;
      RECT 37.205 6.32 37.6 6.485 ;
      RECT 37.825 5.92 38.115 6.15 ;
      RECT 37.825 5.95 38.285 6.12 ;
      RECT 36.835 2.73 37.125 2.96 ;
      RECT 36.835 2.76 37.295 2.93 ;
      RECT 36.9 1.655 37.065 2.96 ;
      RECT 35.415 1.625 35.705 1.855 ;
      RECT 35.415 1.655 37.065 1.825 ;
      RECT 35.475 0.885 35.645 1.855 ;
      RECT 35.415 0.885 35.705 1.115 ;
      RECT 35.415 7.765 35.705 7.995 ;
      RECT 35.475 7.025 35.645 7.995 ;
      RECT 35.475 7.12 37.065 7.29 ;
      RECT 36.895 5.92 37.065 7.29 ;
      RECT 35.415 7.025 35.705 7.255 ;
      RECT 36.835 5.92 37.125 6.15 ;
      RECT 36.835 5.95 37.295 6.12 ;
      RECT 33.45 3.43 33.8 3.78 ;
      RECT 33.54 2.025 33.71 3.78 ;
      RECT 35.845 1.965 36.195 2.315 ;
      RECT 33.54 2.025 35.16 2.2 ;
      RECT 33.54 2.025 36.195 2.195 ;
      RECT 35.87 6.655 36.195 6.98 ;
      RECT 31.295 6.61 31.645 6.96 ;
      RECT 35.845 6.655 36.195 6.885 ;
      RECT 31.085 6.655 31.645 6.885 ;
      RECT 30.915 6.685 36.195 6.855 ;
      RECT 35.07 2.365 35.39 2.685 ;
      RECT 35.04 2.365 35.39 2.595 ;
      RECT 34.87 2.395 35.39 2.565 ;
      RECT 35.07 6.225 35.39 6.545 ;
      RECT 35.04 6.285 35.39 6.515 ;
      RECT 34.87 6.315 35.39 6.485 ;
      RECT 30.85 3.665 30.89 3.925 ;
      RECT 30.89 3.645 30.895 3.655 ;
      RECT 32.22 2.89 32.23 3.111 ;
      RECT 32.15 2.885 32.22 3.236 ;
      RECT 32.14 2.885 32.15 3.363 ;
      RECT 32.115 2.885 32.14 3.41 ;
      RECT 32.09 2.885 32.115 3.488 ;
      RECT 32.07 2.885 32.09 3.558 ;
      RECT 32.045 2.885 32.07 3.598 ;
      RECT 32.035 2.885 32.045 3.618 ;
      RECT 32.025 2.887 32.035 3.626 ;
      RECT 32.02 2.892 32.025 3.083 ;
      RECT 32.02 3.092 32.025 3.627 ;
      RECT 32.015 3.137 32.02 3.628 ;
      RECT 32.005 3.202 32.015 3.629 ;
      RECT 31.995 3.297 32.005 3.631 ;
      RECT 31.99 3.35 31.995 3.633 ;
      RECT 31.985 3.37 31.99 3.634 ;
      RECT 31.93 3.395 31.985 3.64 ;
      RECT 31.89 3.43 31.93 3.649 ;
      RECT 31.88 3.447 31.89 3.654 ;
      RECT 31.871 3.453 31.88 3.656 ;
      RECT 31.785 3.491 31.871 3.667 ;
      RECT 31.78 3.53 31.785 3.677 ;
      RECT 31.705 3.537 31.78 3.687 ;
      RECT 31.685 3.547 31.705 3.698 ;
      RECT 31.655 3.554 31.685 3.706 ;
      RECT 31.63 3.561 31.655 3.713 ;
      RECT 31.606 3.567 31.63 3.718 ;
      RECT 31.52 3.58 31.606 3.73 ;
      RECT 31.442 3.587 31.52 3.748 ;
      RECT 31.356 3.582 31.442 3.766 ;
      RECT 31.27 3.577 31.356 3.786 ;
      RECT 31.19 3.571 31.27 3.803 ;
      RECT 31.125 3.567 31.19 3.832 ;
      RECT 31.12 3.281 31.125 3.305 ;
      RECT 31.11 3.557 31.125 3.86 ;
      RECT 31.115 3.275 31.12 3.345 ;
      RECT 31.11 3.269 31.115 3.415 ;
      RECT 31.105 3.263 31.11 3.493 ;
      RECT 31.105 3.54 31.11 3.925 ;
      RECT 31.097 3.26 31.105 3.925 ;
      RECT 31.011 3.258 31.097 3.925 ;
      RECT 30.925 3.256 31.011 3.925 ;
      RECT 30.915 3.257 30.925 3.925 ;
      RECT 30.91 3.262 30.915 3.925 ;
      RECT 30.9 3.275 30.91 3.925 ;
      RECT 30.895 3.297 30.9 3.925 ;
      RECT 30.89 3.657 30.895 3.925 ;
      RECT 31.52 3.125 31.525 3.345 ;
      RECT 32.025 2.16 32.06 2.42 ;
      RECT 32.01 2.16 32.025 2.428 ;
      RECT 31.981 2.16 32.01 2.45 ;
      RECT 31.895 2.16 31.981 2.51 ;
      RECT 31.875 2.16 31.895 2.575 ;
      RECT 31.815 2.16 31.875 2.74 ;
      RECT 31.81 2.16 31.815 2.888 ;
      RECT 31.805 2.16 31.81 2.9 ;
      RECT 31.8 2.16 31.805 2.926 ;
      RECT 31.77 2.346 31.8 3.006 ;
      RECT 31.765 2.394 31.77 3.095 ;
      RECT 31.76 2.408 31.765 3.11 ;
      RECT 31.755 2.427 31.76 3.14 ;
      RECT 31.75 2.442 31.755 3.156 ;
      RECT 31.745 2.457 31.75 3.178 ;
      RECT 31.74 2.477 31.745 3.2 ;
      RECT 31.73 2.497 31.74 3.233 ;
      RECT 31.715 2.539 31.73 3.295 ;
      RECT 31.71 2.57 31.715 3.335 ;
      RECT 31.705 2.582 31.71 3.34 ;
      RECT 31.7 2.594 31.705 3.345 ;
      RECT 31.695 2.607 31.7 3.345 ;
      RECT 31.69 2.625 31.695 3.345 ;
      RECT 31.685 2.645 31.69 3.345 ;
      RECT 31.68 2.657 31.685 3.345 ;
      RECT 31.675 2.67 31.68 3.345 ;
      RECT 31.655 2.705 31.675 3.345 ;
      RECT 31.605 2.807 31.655 3.345 ;
      RECT 31.6 2.892 31.605 3.345 ;
      RECT 31.595 2.9 31.6 3.345 ;
      RECT 31.59 2.917 31.595 3.345 ;
      RECT 31.585 2.932 31.59 3.345 ;
      RECT 31.55 2.997 31.585 3.345 ;
      RECT 31.535 3.062 31.55 3.345 ;
      RECT 31.53 3.092 31.535 3.345 ;
      RECT 31.525 3.117 31.53 3.345 ;
      RECT 31.51 3.127 31.52 3.345 ;
      RECT 31.495 3.14 31.51 3.338 ;
      RECT 31.24 2.73 31.31 2.94 ;
      RECT 31.03 2.707 31.035 2.9 ;
      RECT 28.485 2.635 28.745 2.895 ;
      RECT 31.32 2.917 31.325 2.92 ;
      RECT 31.31 2.735 31.32 2.935 ;
      RECT 31.211 2.728 31.24 2.94 ;
      RECT 31.125 2.72 31.211 2.94 ;
      RECT 31.11 2.714 31.125 2.938 ;
      RECT 31.09 2.713 31.11 2.925 ;
      RECT 31.085 2.712 31.09 2.908 ;
      RECT 31.035 2.709 31.085 2.903 ;
      RECT 31.005 2.706 31.03 2.898 ;
      RECT 30.985 2.704 31.005 2.893 ;
      RECT 30.97 2.702 30.985 2.89 ;
      RECT 30.94 2.7 30.97 2.888 ;
      RECT 30.875 2.696 30.94 2.88 ;
      RECT 30.845 2.691 30.875 2.875 ;
      RECT 30.825 2.689 30.845 2.873 ;
      RECT 30.795 2.686 30.825 2.868 ;
      RECT 30.735 2.682 30.795 2.86 ;
      RECT 30.73 2.679 30.735 2.855 ;
      RECT 30.66 2.677 30.73 2.85 ;
      RECT 30.631 2.673 30.66 2.843 ;
      RECT 30.545 2.668 30.631 2.835 ;
      RECT 30.511 2.663 30.545 2.827 ;
      RECT 30.425 2.655 30.511 2.819 ;
      RECT 30.386 2.648 30.425 2.811 ;
      RECT 30.3 2.643 30.386 2.803 ;
      RECT 30.235 2.637 30.3 2.793 ;
      RECT 30.215 2.632 30.235 2.788 ;
      RECT 30.206 2.629 30.215 2.787 ;
      RECT 30.12 2.625 30.206 2.781 ;
      RECT 30.08 2.621 30.12 2.773 ;
      RECT 30.06 2.617 30.08 2.771 ;
      RECT 30 2.617 30.06 2.768 ;
      RECT 29.98 2.62 30 2.766 ;
      RECT 29.959 2.62 29.98 2.766 ;
      RECT 29.873 2.622 29.959 2.77 ;
      RECT 29.787 2.624 29.873 2.776 ;
      RECT 29.701 2.626 29.787 2.783 ;
      RECT 29.615 2.629 29.701 2.789 ;
      RECT 29.581 2.63 29.615 2.794 ;
      RECT 29.495 2.633 29.581 2.799 ;
      RECT 29.466 2.64 29.495 2.804 ;
      RECT 29.38 2.64 29.466 2.809 ;
      RECT 29.347 2.64 29.38 2.814 ;
      RECT 29.261 2.642 29.347 2.819 ;
      RECT 29.175 2.644 29.261 2.826 ;
      RECT 29.111 2.646 29.175 2.832 ;
      RECT 29.025 2.648 29.111 2.838 ;
      RECT 29.022 2.65 29.025 2.841 ;
      RECT 28.936 2.651 29.022 2.845 ;
      RECT 28.85 2.654 28.936 2.852 ;
      RECT 28.831 2.656 28.85 2.856 ;
      RECT 28.745 2.658 28.831 2.861 ;
      RECT 28.475 2.67 28.485 2.865 ;
      RECT 30.655 7.765 30.945 7.995 ;
      RECT 30.715 7.025 30.885 7.995 ;
      RECT 30.605 7.055 30.98 7.425 ;
      RECT 30.655 7.025 30.945 7.425 ;
      RECT 30.71 2.25 30.895 2.46 ;
      RECT 30.705 2.251 30.9 2.458 ;
      RECT 30.7 2.256 30.91 2.453 ;
      RECT 30.695 2.232 30.7 2.45 ;
      RECT 30.665 2.229 30.695 2.443 ;
      RECT 30.66 2.225 30.665 2.434 ;
      RECT 30.625 2.256 30.91 2.429 ;
      RECT 30.4 2.165 30.66 2.425 ;
      RECT 30.7 2.234 30.705 2.453 ;
      RECT 30.705 2.235 30.71 2.458 ;
      RECT 30.4 2.247 30.78 2.425 ;
      RECT 30.4 2.245 30.765 2.425 ;
      RECT 30.4 2.24 30.755 2.425 ;
      RECT 30.355 3.155 30.405 3.44 ;
      RECT 30.3 3.125 30.305 3.44 ;
      RECT 30.27 3.105 30.275 3.44 ;
      RECT 30.42 3.155 30.48 3.415 ;
      RECT 30.415 3.155 30.42 3.423 ;
      RECT 30.405 3.155 30.415 3.435 ;
      RECT 30.32 3.145 30.355 3.44 ;
      RECT 30.315 3.132 30.32 3.44 ;
      RECT 30.305 3.127 30.315 3.44 ;
      RECT 30.285 3.117 30.3 3.44 ;
      RECT 30.275 3.11 30.285 3.44 ;
      RECT 30.265 3.102 30.27 3.44 ;
      RECT 30.235 3.092 30.265 3.44 ;
      RECT 30.22 3.08 30.235 3.44 ;
      RECT 30.205 3.07 30.22 3.435 ;
      RECT 30.185 3.06 30.205 3.41 ;
      RECT 30.175 3.052 30.185 3.387 ;
      RECT 30.145 3.035 30.175 3.377 ;
      RECT 30.14 3.012 30.145 3.368 ;
      RECT 30.135 2.999 30.14 3.366 ;
      RECT 30.12 2.975 30.135 3.36 ;
      RECT 30.115 2.951 30.12 3.354 ;
      RECT 30.105 2.94 30.115 3.349 ;
      RECT 30.1 2.93 30.105 3.345 ;
      RECT 30.095 2.922 30.1 3.342 ;
      RECT 30.085 2.917 30.095 3.338 ;
      RECT 30.08 2.912 30.085 3.334 ;
      RECT 29.995 2.91 30.08 3.309 ;
      RECT 29.965 2.91 29.995 3.275 ;
      RECT 29.95 2.91 29.965 3.258 ;
      RECT 29.895 2.91 29.95 3.203 ;
      RECT 29.89 2.915 29.895 3.152 ;
      RECT 29.88 2.92 29.89 3.142 ;
      RECT 29.875 2.93 29.88 3.128 ;
      RECT 29.825 3.67 30.085 3.93 ;
      RECT 29.745 3.685 30.085 3.906 ;
      RECT 29.725 3.685 30.085 3.901 ;
      RECT 29.701 3.685 30.085 3.899 ;
      RECT 29.615 3.685 30.085 3.894 ;
      RECT 29.465 3.625 29.725 3.89 ;
      RECT 29.42 3.685 30.085 3.885 ;
      RECT 29.415 3.692 30.085 3.88 ;
      RECT 29.43 3.68 29.745 3.89 ;
      RECT 29.32 2.115 29.58 2.375 ;
      RECT 29.32 2.172 29.585 2.368 ;
      RECT 29.32 2.202 29.59 2.3 ;
      RECT 29.38 2.633 29.495 2.635 ;
      RECT 29.466 2.63 29.495 2.635 ;
      RECT 28.49 3.634 28.515 3.874 ;
      RECT 28.475 3.637 28.565 3.868 ;
      RECT 28.47 3.642 28.651 3.863 ;
      RECT 28.465 3.65 28.715 3.861 ;
      RECT 28.465 3.65 28.725 3.86 ;
      RECT 28.46 3.657 28.735 3.853 ;
      RECT 28.46 3.657 28.821 3.842 ;
      RECT 28.455 3.692 28.821 3.838 ;
      RECT 28.455 3.692 28.83 3.827 ;
      RECT 28.735 3.565 28.995 3.825 ;
      RECT 28.445 3.742 28.995 3.823 ;
      RECT 28.715 3.61 28.735 3.858 ;
      RECT 28.651 3.613 28.715 3.862 ;
      RECT 28.565 3.618 28.651 3.867 ;
      RECT 28.495 3.629 28.995 3.825 ;
      RECT 28.515 3.623 28.565 3.872 ;
      RECT 28.64 2.1 28.65 2.362 ;
      RECT 28.63 2.157 28.64 2.365 ;
      RECT 28.605 2.162 28.63 2.371 ;
      RECT 28.58 2.166 28.605 2.383 ;
      RECT 28.57 2.169 28.58 2.393 ;
      RECT 28.565 2.17 28.57 2.398 ;
      RECT 28.56 2.171 28.565 2.403 ;
      RECT 28.555 2.172 28.56 2.405 ;
      RECT 28.53 2.175 28.555 2.408 ;
      RECT 28.5 2.181 28.53 2.411 ;
      RECT 28.435 2.192 28.5 2.414 ;
      RECT 28.39 2.2 28.435 2.418 ;
      RECT 28.375 2.2 28.39 2.426 ;
      RECT 28.37 2.201 28.375 2.433 ;
      RECT 28.365 2.203 28.37 2.436 ;
      RECT 28.36 2.207 28.365 2.439 ;
      RECT 28.35 2.215 28.36 2.443 ;
      RECT 28.345 2.228 28.35 2.448 ;
      RECT 28.34 2.236 28.345 2.45 ;
      RECT 28.335 2.242 28.34 2.45 ;
      RECT 28.33 2.246 28.335 2.453 ;
      RECT 28.325 2.248 28.33 2.456 ;
      RECT 28.32 2.251 28.325 2.459 ;
      RECT 28.31 2.256 28.32 2.463 ;
      RECT 28.305 2.262 28.31 2.468 ;
      RECT 28.295 2.268 28.305 2.472 ;
      RECT 28.28 2.275 28.295 2.478 ;
      RECT 28.251 2.289 28.28 2.488 ;
      RECT 28.165 2.324 28.251 2.52 ;
      RECT 28.145 2.357 28.165 2.549 ;
      RECT 28.125 2.37 28.145 2.56 ;
      RECT 28.105 2.382 28.125 2.571 ;
      RECT 28.055 2.404 28.105 2.591 ;
      RECT 28.04 2.422 28.055 2.608 ;
      RECT 28.035 2.428 28.04 2.611 ;
      RECT 28.03 2.432 28.035 2.614 ;
      RECT 28.025 2.436 28.03 2.618 ;
      RECT 28.02 2.438 28.025 2.621 ;
      RECT 28.01 2.445 28.02 2.624 ;
      RECT 28.005 2.45 28.01 2.628 ;
      RECT 28 2.452 28.005 2.631 ;
      RECT 27.995 2.456 28 2.634 ;
      RECT 27.99 2.458 27.995 2.638 ;
      RECT 27.975 2.463 27.99 2.643 ;
      RECT 27.97 2.468 27.975 2.646 ;
      RECT 27.965 2.476 27.97 2.649 ;
      RECT 27.96 2.478 27.965 2.652 ;
      RECT 27.955 2.48 27.96 2.655 ;
      RECT 27.945 2.482 27.955 2.661 ;
      RECT 27.91 2.496 27.945 2.673 ;
      RECT 27.9 2.511 27.91 2.683 ;
      RECT 27.825 2.54 27.9 2.707 ;
      RECT 27.82 2.565 27.825 2.73 ;
      RECT 27.805 2.569 27.82 2.736 ;
      RECT 27.795 2.577 27.805 2.741 ;
      RECT 27.765 2.59 27.795 2.745 ;
      RECT 27.755 2.605 27.765 2.75 ;
      RECT 27.745 2.61 27.755 2.753 ;
      RECT 27.74 2.612 27.745 2.755 ;
      RECT 27.725 2.615 27.74 2.758 ;
      RECT 27.72 2.617 27.725 2.761 ;
      RECT 27.7 2.622 27.72 2.765 ;
      RECT 27.67 2.627 27.7 2.773 ;
      RECT 27.645 2.634 27.67 2.781 ;
      RECT 27.64 2.639 27.645 2.786 ;
      RECT 27.61 2.642 27.64 2.79 ;
      RECT 27.57 2.645 27.61 2.8 ;
      RECT 27.535 2.642 27.57 2.812 ;
      RECT 27.525 2.638 27.535 2.819 ;
      RECT 27.5 2.634 27.525 2.825 ;
      RECT 27.495 2.63 27.5 2.83 ;
      RECT 27.455 2.627 27.495 2.83 ;
      RECT 27.44 2.612 27.455 2.831 ;
      RECT 27.417 2.6 27.44 2.831 ;
      RECT 27.331 2.6 27.417 2.832 ;
      RECT 27.245 2.6 27.331 2.834 ;
      RECT 27.225 2.6 27.245 2.831 ;
      RECT 27.22 2.605 27.225 2.826 ;
      RECT 27.215 2.61 27.22 2.824 ;
      RECT 27.205 2.62 27.215 2.822 ;
      RECT 27.2 2.626 27.205 2.815 ;
      RECT 27.195 2.628 27.2 2.8 ;
      RECT 27.19 2.632 27.195 2.79 ;
      RECT 28.65 2.1 28.9 2.36 ;
      RECT 26.375 3.635 26.635 3.895 ;
      RECT 28.67 3.125 28.675 3.335 ;
      RECT 28.675 3.13 28.685 3.33 ;
      RECT 28.625 3.125 28.67 3.35 ;
      RECT 28.615 3.125 28.625 3.37 ;
      RECT 28.596 3.125 28.615 3.375 ;
      RECT 28.51 3.125 28.596 3.372 ;
      RECT 28.48 3.127 28.51 3.37 ;
      RECT 28.425 3.137 28.48 3.368 ;
      RECT 28.36 3.151 28.425 3.366 ;
      RECT 28.355 3.159 28.36 3.365 ;
      RECT 28.34 3.162 28.355 3.363 ;
      RECT 28.275 3.172 28.34 3.359 ;
      RECT 28.227 3.186 28.275 3.36 ;
      RECT 28.141 3.203 28.227 3.374 ;
      RECT 28.055 3.224 28.141 3.391 ;
      RECT 28.035 3.237 28.055 3.401 ;
      RECT 27.99 3.245 28.035 3.408 ;
      RECT 27.955 3.253 27.99 3.416 ;
      RECT 27.921 3.261 27.955 3.424 ;
      RECT 27.835 3.275 27.921 3.436 ;
      RECT 27.8 3.292 27.835 3.448 ;
      RECT 27.791 3.301 27.8 3.452 ;
      RECT 27.705 3.319 27.791 3.469 ;
      RECT 27.646 3.346 27.705 3.496 ;
      RECT 27.56 3.373 27.646 3.524 ;
      RECT 27.54 3.395 27.56 3.544 ;
      RECT 27.48 3.41 27.54 3.56 ;
      RECT 27.47 3.422 27.48 3.573 ;
      RECT 27.465 3.427 27.47 3.576 ;
      RECT 27.455 3.43 27.465 3.579 ;
      RECT 27.45 3.432 27.455 3.582 ;
      RECT 27.42 3.44 27.45 3.589 ;
      RECT 27.405 3.447 27.42 3.597 ;
      RECT 27.395 3.452 27.405 3.601 ;
      RECT 27.39 3.455 27.395 3.604 ;
      RECT 27.38 3.457 27.39 3.607 ;
      RECT 27.345 3.467 27.38 3.616 ;
      RECT 27.27 3.49 27.345 3.638 ;
      RECT 27.25 3.508 27.27 3.656 ;
      RECT 27.22 3.515 27.25 3.666 ;
      RECT 27.2 3.523 27.22 3.676 ;
      RECT 27.19 3.529 27.2 3.683 ;
      RECT 27.171 3.534 27.19 3.689 ;
      RECT 27.085 3.554 27.171 3.709 ;
      RECT 27.07 3.574 27.085 3.728 ;
      RECT 27.025 3.586 27.07 3.739 ;
      RECT 26.96 3.607 27.025 3.762 ;
      RECT 26.92 3.627 26.96 3.783 ;
      RECT 26.91 3.637 26.92 3.793 ;
      RECT 26.86 3.649 26.91 3.804 ;
      RECT 26.84 3.665 26.86 3.816 ;
      RECT 26.81 3.675 26.84 3.822 ;
      RECT 26.8 3.68 26.81 3.824 ;
      RECT 26.731 3.681 26.8 3.83 ;
      RECT 26.645 3.683 26.731 3.84 ;
      RECT 26.635 3.684 26.645 3.845 ;
      RECT 27.905 3.71 28.095 3.92 ;
      RECT 27.895 3.715 28.105 3.913 ;
      RECT 27.88 3.715 28.105 3.878 ;
      RECT 27.8 3.6 28.06 3.86 ;
      RECT 26.715 3.13 26.9 3.425 ;
      RECT 26.705 3.13 26.9 3.423 ;
      RECT 26.69 3.13 26.905 3.418 ;
      RECT 26.69 3.13 26.91 3.415 ;
      RECT 26.685 3.13 26.91 3.413 ;
      RECT 26.68 3.385 26.91 3.403 ;
      RECT 26.685 3.13 26.945 3.39 ;
      RECT 26.645 2.165 26.905 2.425 ;
      RECT 26.455 2.09 26.541 2.423 ;
      RECT 26.43 2.094 26.585 2.419 ;
      RECT 26.541 2.086 26.585 2.419 ;
      RECT 26.541 2.087 26.59 2.418 ;
      RECT 26.455 2.092 26.605 2.417 ;
      RECT 26.43 2.1 26.645 2.416 ;
      RECT 26.425 2.095 26.605 2.411 ;
      RECT 26.415 2.11 26.645 2.318 ;
      RECT 26.415 2.162 26.845 2.318 ;
      RECT 26.415 2.155 26.825 2.318 ;
      RECT 26.415 2.142 26.795 2.318 ;
      RECT 26.415 2.13 26.735 2.318 ;
      RECT 26.415 2.115 26.71 2.318 ;
      RECT 25.615 2.745 25.75 3.04 ;
      RECT 25.875 2.768 25.88 2.955 ;
      RECT 26.595 2.665 26.74 2.9 ;
      RECT 26.755 2.665 26.76 2.89 ;
      RECT 26.79 2.676 26.795 2.87 ;
      RECT 26.785 2.668 26.79 2.875 ;
      RECT 26.765 2.665 26.785 2.88 ;
      RECT 26.76 2.665 26.765 2.888 ;
      RECT 26.75 2.665 26.755 2.893 ;
      RECT 26.74 2.665 26.75 2.898 ;
      RECT 26.57 2.667 26.595 2.9 ;
      RECT 26.52 2.674 26.57 2.9 ;
      RECT 26.515 2.679 26.52 2.9 ;
      RECT 26.476 2.684 26.515 2.901 ;
      RECT 26.39 2.696 26.476 2.902 ;
      RECT 26.381 2.706 26.39 2.902 ;
      RECT 26.295 2.715 26.381 2.904 ;
      RECT 26.271 2.725 26.295 2.906 ;
      RECT 26.185 2.736 26.271 2.907 ;
      RECT 26.155 2.747 26.185 2.909 ;
      RECT 26.125 2.752 26.155 2.911 ;
      RECT 26.1 2.758 26.125 2.914 ;
      RECT 26.085 2.763 26.1 2.915 ;
      RECT 26.04 2.769 26.085 2.915 ;
      RECT 26.035 2.774 26.04 2.916 ;
      RECT 26.015 2.774 26.035 2.918 ;
      RECT 25.995 2.772 26.015 2.923 ;
      RECT 25.96 2.771 25.995 2.93 ;
      RECT 25.93 2.77 25.96 2.94 ;
      RECT 25.88 2.769 25.93 2.95 ;
      RECT 25.79 2.766 25.875 3.04 ;
      RECT 25.765 2.76 25.79 3.04 ;
      RECT 25.75 2.75 25.765 3.04 ;
      RECT 25.565 2.745 25.615 2.96 ;
      RECT 25.555 2.75 25.565 2.95 ;
      RECT 25.795 3.225 26.055 3.485 ;
      RECT 25.795 3.225 26.085 3.378 ;
      RECT 25.795 3.225 26.12 3.363 ;
      RECT 26.05 3.145 26.24 3.355 ;
      RECT 26.04 3.15 26.25 3.348 ;
      RECT 26.005 3.22 26.25 3.348 ;
      RECT 26.035 3.162 26.055 3.485 ;
      RECT 26.02 3.21 26.25 3.348 ;
      RECT 26.025 3.182 26.055 3.485 ;
      RECT 25.105 2.25 25.175 3.355 ;
      RECT 25.84 2.355 26.1 2.615 ;
      RECT 25.42 2.401 25.435 2.61 ;
      RECT 25.756 2.414 25.84 2.565 ;
      RECT 25.67 2.411 25.756 2.565 ;
      RECT 25.631 2.409 25.67 2.565 ;
      RECT 25.545 2.407 25.631 2.565 ;
      RECT 25.485 2.405 25.545 2.576 ;
      RECT 25.45 2.403 25.485 2.594 ;
      RECT 25.435 2.401 25.45 2.605 ;
      RECT 25.405 2.401 25.42 2.618 ;
      RECT 25.395 2.401 25.405 2.623 ;
      RECT 25.37 2.4 25.395 2.628 ;
      RECT 25.355 2.395 25.37 2.634 ;
      RECT 25.35 2.388 25.355 2.639 ;
      RECT 25.325 2.379 25.35 2.645 ;
      RECT 25.28 2.358 25.325 2.658 ;
      RECT 25.27 2.342 25.28 2.668 ;
      RECT 25.255 2.335 25.27 2.678 ;
      RECT 25.245 2.328 25.255 2.695 ;
      RECT 25.24 2.325 25.245 2.725 ;
      RECT 25.235 2.323 25.24 2.755 ;
      RECT 25.23 2.321 25.235 2.792 ;
      RECT 25.215 2.317 25.23 2.859 ;
      RECT 25.215 3.15 25.225 3.35 ;
      RECT 25.21 2.313 25.215 2.985 ;
      RECT 25.21 3.137 25.215 3.355 ;
      RECT 25.205 2.311 25.21 3.07 ;
      RECT 25.205 3.127 25.21 3.355 ;
      RECT 25.19 2.282 25.205 3.355 ;
      RECT 25.175 2.255 25.19 3.355 ;
      RECT 25.1 2.25 25.105 2.605 ;
      RECT 25.1 2.66 25.105 3.355 ;
      RECT 25.085 2.25 25.1 2.583 ;
      RECT 25.095 2.682 25.1 3.355 ;
      RECT 25.085 2.722 25.095 3.355 ;
      RECT 25.05 2.25 25.085 2.525 ;
      RECT 25.08 2.757 25.085 3.355 ;
      RECT 25.065 2.812 25.08 3.355 ;
      RECT 25.06 2.877 25.065 3.355 ;
      RECT 25.045 2.925 25.06 3.355 ;
      RECT 25.02 2.25 25.05 2.48 ;
      RECT 25.04 2.98 25.045 3.355 ;
      RECT 25.025 3.04 25.04 3.355 ;
      RECT 25.02 3.088 25.025 3.353 ;
      RECT 25.015 2.25 25.02 2.473 ;
      RECT 25.015 3.12 25.02 3.348 ;
      RECT 24.99 2.25 25.015 2.465 ;
      RECT 24.98 2.255 24.99 2.455 ;
      RECT 25.195 3.53 25.215 3.77 ;
      RECT 24.425 3.46 24.43 3.67 ;
      RECT 25.705 3.533 25.715 3.728 ;
      RECT 25.7 3.523 25.705 3.731 ;
      RECT 25.62 3.52 25.7 3.754 ;
      RECT 25.616 3.52 25.62 3.776 ;
      RECT 25.53 3.52 25.616 3.786 ;
      RECT 25.515 3.52 25.53 3.794 ;
      RECT 25.486 3.521 25.515 3.792 ;
      RECT 25.4 3.526 25.486 3.788 ;
      RECT 25.387 3.53 25.4 3.784 ;
      RECT 25.301 3.53 25.387 3.78 ;
      RECT 25.215 3.53 25.301 3.774 ;
      RECT 25.131 3.53 25.195 3.768 ;
      RECT 25.045 3.53 25.131 3.763 ;
      RECT 25.025 3.53 25.045 3.759 ;
      RECT 24.965 3.525 25.025 3.756 ;
      RECT 24.937 3.519 24.965 3.753 ;
      RECT 24.851 3.514 24.937 3.749 ;
      RECT 24.765 3.508 24.851 3.743 ;
      RECT 24.69 3.49 24.765 3.738 ;
      RECT 24.655 3.467 24.69 3.734 ;
      RECT 24.645 3.457 24.655 3.733 ;
      RECT 24.59 3.455 24.645 3.732 ;
      RECT 24.515 3.455 24.59 3.728 ;
      RECT 24.505 3.455 24.515 3.723 ;
      RECT 24.49 3.455 24.505 3.715 ;
      RECT 24.44 3.457 24.49 3.693 ;
      RECT 24.43 3.46 24.44 3.673 ;
      RECT 24.42 3.465 24.425 3.668 ;
      RECT 24.415 3.47 24.42 3.663 ;
      RECT 24.54 2.635 24.8 2.895 ;
      RECT 24.54 2.65 24.82 2.86 ;
      RECT 24.54 2.655 24.83 2.855 ;
      RECT 22.525 2.115 22.785 2.375 ;
      RECT 22.515 2.145 22.785 2.355 ;
      RECT 24.435 2.06 24.695 2.32 ;
      RECT 24.43 2.135 24.435 2.321 ;
      RECT 24.405 2.14 24.43 2.323 ;
      RECT 24.39 2.147 24.405 2.326 ;
      RECT 24.33 2.165 24.39 2.331 ;
      RECT 24.3 2.185 24.33 2.338 ;
      RECT 24.275 2.193 24.3 2.343 ;
      RECT 24.25 2.201 24.275 2.345 ;
      RECT 24.232 2.205 24.25 2.344 ;
      RECT 24.146 2.203 24.232 2.344 ;
      RECT 24.06 2.201 24.146 2.344 ;
      RECT 23.974 2.199 24.06 2.343 ;
      RECT 23.888 2.197 23.974 2.343 ;
      RECT 23.802 2.195 23.888 2.343 ;
      RECT 23.716 2.193 23.802 2.343 ;
      RECT 23.63 2.191 23.716 2.342 ;
      RECT 23.612 2.19 23.63 2.342 ;
      RECT 23.526 2.189 23.612 2.342 ;
      RECT 23.44 2.187 23.526 2.342 ;
      RECT 23.354 2.186 23.44 2.341 ;
      RECT 23.268 2.185 23.354 2.341 ;
      RECT 23.182 2.183 23.268 2.341 ;
      RECT 23.096 2.182 23.182 2.341 ;
      RECT 23.01 2.18 23.096 2.34 ;
      RECT 22.986 2.178 23.01 2.34 ;
      RECT 22.9 2.171 22.986 2.34 ;
      RECT 22.871 2.163 22.9 2.34 ;
      RECT 22.785 2.155 22.871 2.34 ;
      RECT 22.505 2.152 22.515 2.35 ;
      RECT 24.01 3.115 24.015 3.465 ;
      RECT 23.78 3.205 23.92 3.465 ;
      RECT 24.255 2.89 24.3 3.1 ;
      RECT 24.31 2.901 24.32 3.095 ;
      RECT 24.3 2.893 24.31 3.1 ;
      RECT 24.235 2.89 24.255 3.105 ;
      RECT 24.205 2.89 24.235 3.128 ;
      RECT 24.195 2.89 24.205 3.153 ;
      RECT 24.19 2.89 24.195 3.163 ;
      RECT 24.135 2.89 24.19 3.203 ;
      RECT 24.13 2.89 24.135 3.243 ;
      RECT 24.125 2.892 24.13 3.248 ;
      RECT 24.11 2.902 24.125 3.259 ;
      RECT 24.065 2.96 24.11 3.295 ;
      RECT 24.055 3.015 24.065 3.329 ;
      RECT 24.04 3.042 24.055 3.345 ;
      RECT 24.03 3.069 24.04 3.465 ;
      RECT 24.015 3.092 24.03 3.465 ;
      RECT 24.005 3.132 24.01 3.465 ;
      RECT 24 3.142 24.005 3.465 ;
      RECT 23.995 3.157 24 3.465 ;
      RECT 23.985 3.162 23.995 3.465 ;
      RECT 23.92 3.185 23.985 3.465 ;
      RECT 23.42 2.68 23.61 2.89 ;
      RECT 21.995 2.605 22.255 2.865 ;
      RECT 22.345 2.6 22.44 2.81 ;
      RECT 22.32 2.615 22.33 2.81 ;
      RECT 23.61 2.687 23.62 2.885 ;
      RECT 23.41 2.687 23.42 2.885 ;
      RECT 23.395 2.702 23.41 2.875 ;
      RECT 23.39 2.71 23.395 2.868 ;
      RECT 23.38 2.713 23.39 2.865 ;
      RECT 23.345 2.712 23.38 2.863 ;
      RECT 23.316 2.708 23.345 2.86 ;
      RECT 23.23 2.703 23.316 2.857 ;
      RECT 23.17 2.697 23.23 2.853 ;
      RECT 23.141 2.693 23.17 2.85 ;
      RECT 23.055 2.685 23.141 2.847 ;
      RECT 23.046 2.679 23.055 2.845 ;
      RECT 22.96 2.674 23.046 2.843 ;
      RECT 22.937 2.669 22.96 2.84 ;
      RECT 22.851 2.663 22.937 2.837 ;
      RECT 22.765 2.654 22.851 2.832 ;
      RECT 22.755 2.649 22.765 2.83 ;
      RECT 22.736 2.648 22.755 2.829 ;
      RECT 22.65 2.643 22.736 2.825 ;
      RECT 22.63 2.638 22.65 2.821 ;
      RECT 22.57 2.633 22.63 2.818 ;
      RECT 22.545 2.623 22.57 2.816 ;
      RECT 22.54 2.616 22.545 2.815 ;
      RECT 22.53 2.607 22.54 2.814 ;
      RECT 22.526 2.6 22.53 2.814 ;
      RECT 22.44 2.6 22.526 2.812 ;
      RECT 22.33 2.607 22.345 2.81 ;
      RECT 22.315 2.617 22.32 2.81 ;
      RECT 22.295 2.62 22.315 2.807 ;
      RECT 22.265 2.62 22.295 2.803 ;
      RECT 22.255 2.62 22.265 2.803 ;
      RECT 23.17 3.115 23.43 3.375 ;
      RECT 23.1 3.125 23.43 3.335 ;
      RECT 23.09 3.132 23.43 3.33 ;
      RECT 22.51 3.12 22.77 3.38 ;
      RECT 22.51 3.16 22.875 3.37 ;
      RECT 22.51 3.162 22.88 3.369 ;
      RECT 22.51 3.17 22.885 3.366 ;
      RECT 21.435 2.245 21.535 3.77 ;
      RECT 21.625 3.385 21.675 3.645 ;
      RECT 21.62 2.258 21.625 2.445 ;
      RECT 21.615 3.366 21.625 3.645 ;
      RECT 21.615 2.255 21.62 2.453 ;
      RECT 21.6 2.249 21.615 2.46 ;
      RECT 21.61 3.354 21.615 3.728 ;
      RECT 21.6 3.342 21.61 3.765 ;
      RECT 21.59 2.245 21.6 2.467 ;
      RECT 21.59 3.327 21.6 3.77 ;
      RECT 21.585 2.245 21.59 2.475 ;
      RECT 21.565 3.297 21.59 3.77 ;
      RECT 21.545 2.245 21.585 2.523 ;
      RECT 21.555 3.257 21.565 3.77 ;
      RECT 21.545 3.212 21.555 3.77 ;
      RECT 21.54 2.245 21.545 2.593 ;
      RECT 21.54 3.17 21.545 3.77 ;
      RECT 21.535 2.245 21.54 3.07 ;
      RECT 21.535 3.152 21.54 3.77 ;
      RECT 21.425 2.248 21.435 3.77 ;
      RECT 21.41 2.255 21.425 3.766 ;
      RECT 21.405 2.265 21.41 3.761 ;
      RECT 21.4 2.465 21.405 3.653 ;
      RECT 21.395 2.55 21.4 3.205 ;
      RECT 20.27 7.77 20.56 8 ;
      RECT 20.33 6.29 20.5 8 ;
      RECT 20.325 6.655 20.675 7.005 ;
      RECT 20.27 6.29 20.56 6.52 ;
      RECT 19.865 2.395 19.97 2.965 ;
      RECT 19.865 2.73 20.19 2.96 ;
      RECT 19.865 2.76 20.36 2.93 ;
      RECT 19.865 2.395 20.055 2.96 ;
      RECT 19.28 2.36 19.57 2.59 ;
      RECT 19.28 2.395 20.055 2.565 ;
      RECT 19.34 0.88 19.51 2.59 ;
      RECT 19.28 0.88 19.57 1.11 ;
      RECT 19.28 7.77 19.57 8 ;
      RECT 19.34 6.29 19.51 8 ;
      RECT 19.28 6.29 19.57 6.52 ;
      RECT 19.28 6.325 20.135 6.485 ;
      RECT 19.965 5.92 20.135 6.485 ;
      RECT 19.28 6.32 19.675 6.485 ;
      RECT 19.9 5.92 20.19 6.15 ;
      RECT 19.9 5.95 20.36 6.12 ;
      RECT 18.91 2.73 19.2 2.96 ;
      RECT 18.91 2.76 19.37 2.93 ;
      RECT 18.975 1.655 19.14 2.96 ;
      RECT 17.49 1.625 17.78 1.855 ;
      RECT 17.49 1.655 19.14 1.825 ;
      RECT 17.55 0.885 17.72 1.855 ;
      RECT 17.49 0.885 17.78 1.115 ;
      RECT 17.49 7.765 17.78 7.995 ;
      RECT 17.55 7.025 17.72 7.995 ;
      RECT 17.55 7.12 19.14 7.29 ;
      RECT 18.97 5.92 19.14 7.29 ;
      RECT 17.49 7.025 17.78 7.255 ;
      RECT 18.91 5.92 19.2 6.15 ;
      RECT 18.91 5.95 19.37 6.12 ;
      RECT 15.525 3.43 15.875 3.78 ;
      RECT 15.615 2.025 15.785 3.78 ;
      RECT 17.92 1.965 18.27 2.315 ;
      RECT 15.615 2.025 17.235 2.2 ;
      RECT 15.615 2.025 18.27 2.195 ;
      RECT 17.945 6.655 18.27 6.98 ;
      RECT 13.34 6.605 13.69 6.955 ;
      RECT 17.92 6.655 18.27 6.885 ;
      RECT 13.16 6.655 13.69 6.885 ;
      RECT 12.99 6.685 18.27 6.855 ;
      RECT 17.145 2.365 17.465 2.685 ;
      RECT 17.115 2.365 17.465 2.595 ;
      RECT 16.945 2.395 17.465 2.565 ;
      RECT 17.145 6.225 17.465 6.545 ;
      RECT 17.115 6.285 17.465 6.515 ;
      RECT 16.945 6.315 17.465 6.485 ;
      RECT 12.925 3.665 12.965 3.925 ;
      RECT 12.965 3.645 12.97 3.655 ;
      RECT 14.295 2.89 14.305 3.111 ;
      RECT 14.225 2.885 14.295 3.236 ;
      RECT 14.215 2.885 14.225 3.363 ;
      RECT 14.19 2.885 14.215 3.41 ;
      RECT 14.165 2.885 14.19 3.488 ;
      RECT 14.145 2.885 14.165 3.558 ;
      RECT 14.12 2.885 14.145 3.598 ;
      RECT 14.11 2.885 14.12 3.618 ;
      RECT 14.1 2.887 14.11 3.626 ;
      RECT 14.095 2.892 14.1 3.083 ;
      RECT 14.095 3.092 14.1 3.627 ;
      RECT 14.09 3.137 14.095 3.628 ;
      RECT 14.08 3.202 14.09 3.629 ;
      RECT 14.07 3.297 14.08 3.631 ;
      RECT 14.065 3.35 14.07 3.633 ;
      RECT 14.06 3.37 14.065 3.634 ;
      RECT 14.005 3.395 14.06 3.64 ;
      RECT 13.965 3.43 14.005 3.649 ;
      RECT 13.955 3.447 13.965 3.654 ;
      RECT 13.946 3.453 13.955 3.656 ;
      RECT 13.86 3.491 13.946 3.667 ;
      RECT 13.855 3.53 13.86 3.677 ;
      RECT 13.78 3.537 13.855 3.687 ;
      RECT 13.76 3.547 13.78 3.698 ;
      RECT 13.73 3.554 13.76 3.706 ;
      RECT 13.705 3.561 13.73 3.713 ;
      RECT 13.681 3.567 13.705 3.718 ;
      RECT 13.595 3.58 13.681 3.73 ;
      RECT 13.517 3.587 13.595 3.748 ;
      RECT 13.431 3.582 13.517 3.766 ;
      RECT 13.345 3.577 13.431 3.786 ;
      RECT 13.265 3.571 13.345 3.803 ;
      RECT 13.2 3.567 13.265 3.832 ;
      RECT 13.195 3.281 13.2 3.305 ;
      RECT 13.185 3.557 13.2 3.86 ;
      RECT 13.19 3.275 13.195 3.345 ;
      RECT 13.185 3.269 13.19 3.415 ;
      RECT 13.18 3.263 13.185 3.493 ;
      RECT 13.18 3.54 13.185 3.925 ;
      RECT 13.172 3.26 13.18 3.925 ;
      RECT 13.086 3.258 13.172 3.925 ;
      RECT 13 3.256 13.086 3.925 ;
      RECT 12.99 3.257 13 3.925 ;
      RECT 12.985 3.262 12.99 3.925 ;
      RECT 12.975 3.275 12.985 3.925 ;
      RECT 12.97 3.297 12.975 3.925 ;
      RECT 12.965 3.657 12.97 3.925 ;
      RECT 13.595 3.125 13.6 3.345 ;
      RECT 14.1 2.16 14.135 2.42 ;
      RECT 14.085 2.16 14.1 2.428 ;
      RECT 14.056 2.16 14.085 2.45 ;
      RECT 13.97 2.16 14.056 2.51 ;
      RECT 13.95 2.16 13.97 2.575 ;
      RECT 13.89 2.16 13.95 2.74 ;
      RECT 13.885 2.16 13.89 2.888 ;
      RECT 13.88 2.16 13.885 2.9 ;
      RECT 13.875 2.16 13.88 2.926 ;
      RECT 13.845 2.346 13.875 3.006 ;
      RECT 13.84 2.394 13.845 3.095 ;
      RECT 13.835 2.408 13.84 3.11 ;
      RECT 13.83 2.427 13.835 3.14 ;
      RECT 13.825 2.442 13.83 3.156 ;
      RECT 13.82 2.457 13.825 3.178 ;
      RECT 13.815 2.477 13.82 3.2 ;
      RECT 13.805 2.497 13.815 3.233 ;
      RECT 13.79 2.539 13.805 3.295 ;
      RECT 13.785 2.57 13.79 3.335 ;
      RECT 13.78 2.582 13.785 3.34 ;
      RECT 13.775 2.594 13.78 3.345 ;
      RECT 13.77 2.607 13.775 3.345 ;
      RECT 13.765 2.625 13.77 3.345 ;
      RECT 13.76 2.645 13.765 3.345 ;
      RECT 13.755 2.657 13.76 3.345 ;
      RECT 13.75 2.67 13.755 3.345 ;
      RECT 13.73 2.705 13.75 3.345 ;
      RECT 13.68 2.807 13.73 3.345 ;
      RECT 13.675 2.892 13.68 3.345 ;
      RECT 13.67 2.9 13.675 3.345 ;
      RECT 13.665 2.917 13.67 3.345 ;
      RECT 13.66 2.932 13.665 3.345 ;
      RECT 13.625 2.997 13.66 3.345 ;
      RECT 13.61 3.062 13.625 3.345 ;
      RECT 13.605 3.092 13.61 3.345 ;
      RECT 13.6 3.117 13.605 3.345 ;
      RECT 13.585 3.127 13.595 3.345 ;
      RECT 13.57 3.14 13.585 3.338 ;
      RECT 13.315 2.73 13.385 2.94 ;
      RECT 13.105 2.707 13.11 2.9 ;
      RECT 10.56 2.635 10.82 2.895 ;
      RECT 13.395 2.917 13.4 2.92 ;
      RECT 13.385 2.735 13.395 2.935 ;
      RECT 13.286 2.728 13.315 2.94 ;
      RECT 13.2 2.72 13.286 2.94 ;
      RECT 13.185 2.714 13.2 2.938 ;
      RECT 13.165 2.713 13.185 2.925 ;
      RECT 13.16 2.712 13.165 2.908 ;
      RECT 13.11 2.709 13.16 2.903 ;
      RECT 13.08 2.706 13.105 2.898 ;
      RECT 13.06 2.704 13.08 2.893 ;
      RECT 13.045 2.702 13.06 2.89 ;
      RECT 13.015 2.7 13.045 2.888 ;
      RECT 12.95 2.696 13.015 2.88 ;
      RECT 12.92 2.691 12.95 2.875 ;
      RECT 12.9 2.689 12.92 2.873 ;
      RECT 12.87 2.686 12.9 2.868 ;
      RECT 12.81 2.682 12.87 2.86 ;
      RECT 12.805 2.679 12.81 2.855 ;
      RECT 12.735 2.677 12.805 2.85 ;
      RECT 12.706 2.673 12.735 2.843 ;
      RECT 12.62 2.668 12.706 2.835 ;
      RECT 12.586 2.663 12.62 2.827 ;
      RECT 12.5 2.655 12.586 2.819 ;
      RECT 12.461 2.648 12.5 2.811 ;
      RECT 12.375 2.643 12.461 2.803 ;
      RECT 12.31 2.637 12.375 2.793 ;
      RECT 12.29 2.632 12.31 2.788 ;
      RECT 12.281 2.629 12.29 2.787 ;
      RECT 12.195 2.625 12.281 2.781 ;
      RECT 12.155 2.621 12.195 2.773 ;
      RECT 12.135 2.617 12.155 2.771 ;
      RECT 12.075 2.617 12.135 2.768 ;
      RECT 12.055 2.62 12.075 2.766 ;
      RECT 12.034 2.62 12.055 2.766 ;
      RECT 11.948 2.622 12.034 2.77 ;
      RECT 11.862 2.624 11.948 2.776 ;
      RECT 11.776 2.626 11.862 2.783 ;
      RECT 11.69 2.629 11.776 2.789 ;
      RECT 11.656 2.63 11.69 2.794 ;
      RECT 11.57 2.633 11.656 2.799 ;
      RECT 11.541 2.64 11.57 2.804 ;
      RECT 11.455 2.64 11.541 2.809 ;
      RECT 11.422 2.64 11.455 2.814 ;
      RECT 11.336 2.642 11.422 2.819 ;
      RECT 11.25 2.644 11.336 2.826 ;
      RECT 11.186 2.646 11.25 2.832 ;
      RECT 11.1 2.648 11.186 2.838 ;
      RECT 11.097 2.65 11.1 2.841 ;
      RECT 11.011 2.651 11.097 2.845 ;
      RECT 10.925 2.654 11.011 2.852 ;
      RECT 10.906 2.656 10.925 2.856 ;
      RECT 10.82 2.658 10.906 2.861 ;
      RECT 10.55 2.67 10.56 2.865 ;
      RECT 12.73 7.765 13.02 7.995 ;
      RECT 12.79 7.025 12.96 7.995 ;
      RECT 12.68 7.055 13.055 7.425 ;
      RECT 12.73 7.025 13.02 7.425 ;
      RECT 12.785 2.25 12.97 2.46 ;
      RECT 12.78 2.251 12.975 2.458 ;
      RECT 12.775 2.256 12.985 2.453 ;
      RECT 12.77 2.232 12.775 2.45 ;
      RECT 12.74 2.229 12.77 2.443 ;
      RECT 12.735 2.225 12.74 2.434 ;
      RECT 12.7 2.256 12.985 2.429 ;
      RECT 12.475 2.165 12.735 2.425 ;
      RECT 12.775 2.234 12.78 2.453 ;
      RECT 12.78 2.235 12.785 2.458 ;
      RECT 12.475 2.247 12.855 2.425 ;
      RECT 12.475 2.245 12.84 2.425 ;
      RECT 12.475 2.24 12.83 2.425 ;
      RECT 12.43 3.155 12.48 3.44 ;
      RECT 12.375 3.125 12.38 3.44 ;
      RECT 12.345 3.105 12.35 3.44 ;
      RECT 12.495 3.155 12.555 3.415 ;
      RECT 12.49 3.155 12.495 3.423 ;
      RECT 12.48 3.155 12.49 3.435 ;
      RECT 12.395 3.145 12.43 3.44 ;
      RECT 12.39 3.132 12.395 3.44 ;
      RECT 12.38 3.127 12.39 3.44 ;
      RECT 12.36 3.117 12.375 3.44 ;
      RECT 12.35 3.11 12.36 3.44 ;
      RECT 12.34 3.102 12.345 3.44 ;
      RECT 12.31 3.092 12.34 3.44 ;
      RECT 12.295 3.08 12.31 3.44 ;
      RECT 12.28 3.07 12.295 3.435 ;
      RECT 12.26 3.06 12.28 3.41 ;
      RECT 12.25 3.052 12.26 3.387 ;
      RECT 12.22 3.035 12.25 3.377 ;
      RECT 12.215 3.012 12.22 3.368 ;
      RECT 12.21 2.999 12.215 3.366 ;
      RECT 12.195 2.975 12.21 3.36 ;
      RECT 12.19 2.951 12.195 3.354 ;
      RECT 12.18 2.94 12.19 3.349 ;
      RECT 12.175 2.93 12.18 3.345 ;
      RECT 12.17 2.922 12.175 3.342 ;
      RECT 12.16 2.917 12.17 3.338 ;
      RECT 12.155 2.912 12.16 3.334 ;
      RECT 12.07 2.91 12.155 3.309 ;
      RECT 12.04 2.91 12.07 3.275 ;
      RECT 12.025 2.91 12.04 3.258 ;
      RECT 11.97 2.91 12.025 3.203 ;
      RECT 11.965 2.915 11.97 3.152 ;
      RECT 11.955 2.92 11.965 3.142 ;
      RECT 11.95 2.93 11.955 3.128 ;
      RECT 11.9 3.67 12.16 3.93 ;
      RECT 11.82 3.685 12.16 3.906 ;
      RECT 11.8 3.685 12.16 3.901 ;
      RECT 11.776 3.685 12.16 3.899 ;
      RECT 11.69 3.685 12.16 3.894 ;
      RECT 11.54 3.625 11.8 3.89 ;
      RECT 11.495 3.685 12.16 3.885 ;
      RECT 11.49 3.692 12.16 3.88 ;
      RECT 11.505 3.68 11.82 3.89 ;
      RECT 11.395 2.115 11.655 2.375 ;
      RECT 11.395 2.172 11.66 2.368 ;
      RECT 11.395 2.202 11.665 2.3 ;
      RECT 11.455 2.633 11.57 2.635 ;
      RECT 11.541 2.63 11.57 2.635 ;
      RECT 10.565 3.634 10.59 3.874 ;
      RECT 10.55 3.637 10.64 3.868 ;
      RECT 10.545 3.642 10.726 3.863 ;
      RECT 10.54 3.65 10.79 3.861 ;
      RECT 10.54 3.65 10.8 3.86 ;
      RECT 10.535 3.657 10.81 3.853 ;
      RECT 10.535 3.657 10.896 3.842 ;
      RECT 10.53 3.692 10.896 3.838 ;
      RECT 10.53 3.692 10.905 3.827 ;
      RECT 10.81 3.565 11.07 3.825 ;
      RECT 10.52 3.742 11.07 3.823 ;
      RECT 10.79 3.61 10.81 3.858 ;
      RECT 10.726 3.613 10.79 3.862 ;
      RECT 10.64 3.618 10.726 3.867 ;
      RECT 10.57 3.629 11.07 3.825 ;
      RECT 10.59 3.623 10.64 3.872 ;
      RECT 10.715 2.1 10.725 2.362 ;
      RECT 10.705 2.157 10.715 2.365 ;
      RECT 10.68 2.162 10.705 2.371 ;
      RECT 10.655 2.166 10.68 2.383 ;
      RECT 10.645 2.169 10.655 2.393 ;
      RECT 10.64 2.17 10.645 2.398 ;
      RECT 10.635 2.171 10.64 2.403 ;
      RECT 10.63 2.172 10.635 2.405 ;
      RECT 10.605 2.175 10.63 2.408 ;
      RECT 10.575 2.181 10.605 2.411 ;
      RECT 10.51 2.192 10.575 2.414 ;
      RECT 10.465 2.2 10.51 2.418 ;
      RECT 10.45 2.2 10.465 2.426 ;
      RECT 10.445 2.201 10.45 2.433 ;
      RECT 10.44 2.203 10.445 2.436 ;
      RECT 10.435 2.207 10.44 2.439 ;
      RECT 10.425 2.215 10.435 2.443 ;
      RECT 10.42 2.228 10.425 2.448 ;
      RECT 10.415 2.236 10.42 2.45 ;
      RECT 10.41 2.242 10.415 2.45 ;
      RECT 10.405 2.246 10.41 2.453 ;
      RECT 10.4 2.248 10.405 2.456 ;
      RECT 10.395 2.251 10.4 2.459 ;
      RECT 10.385 2.256 10.395 2.463 ;
      RECT 10.38 2.262 10.385 2.468 ;
      RECT 10.37 2.268 10.38 2.472 ;
      RECT 10.355 2.275 10.37 2.478 ;
      RECT 10.326 2.289 10.355 2.488 ;
      RECT 10.24 2.324 10.326 2.52 ;
      RECT 10.22 2.357 10.24 2.549 ;
      RECT 10.2 2.37 10.22 2.56 ;
      RECT 10.18 2.382 10.2 2.571 ;
      RECT 10.13 2.404 10.18 2.591 ;
      RECT 10.115 2.422 10.13 2.608 ;
      RECT 10.11 2.428 10.115 2.611 ;
      RECT 10.105 2.432 10.11 2.614 ;
      RECT 10.1 2.436 10.105 2.618 ;
      RECT 10.095 2.438 10.1 2.621 ;
      RECT 10.085 2.445 10.095 2.624 ;
      RECT 10.08 2.45 10.085 2.628 ;
      RECT 10.075 2.452 10.08 2.631 ;
      RECT 10.07 2.456 10.075 2.634 ;
      RECT 10.065 2.458 10.07 2.638 ;
      RECT 10.05 2.463 10.065 2.643 ;
      RECT 10.045 2.468 10.05 2.646 ;
      RECT 10.04 2.476 10.045 2.649 ;
      RECT 10.035 2.478 10.04 2.652 ;
      RECT 10.03 2.48 10.035 2.655 ;
      RECT 10.02 2.482 10.03 2.661 ;
      RECT 9.985 2.496 10.02 2.673 ;
      RECT 9.975 2.511 9.985 2.683 ;
      RECT 9.9 2.54 9.975 2.707 ;
      RECT 9.895 2.565 9.9 2.73 ;
      RECT 9.88 2.569 9.895 2.736 ;
      RECT 9.87 2.577 9.88 2.741 ;
      RECT 9.84 2.59 9.87 2.745 ;
      RECT 9.83 2.605 9.84 2.75 ;
      RECT 9.82 2.61 9.83 2.753 ;
      RECT 9.815 2.612 9.82 2.755 ;
      RECT 9.8 2.615 9.815 2.758 ;
      RECT 9.795 2.617 9.8 2.761 ;
      RECT 9.775 2.622 9.795 2.765 ;
      RECT 9.745 2.627 9.775 2.773 ;
      RECT 9.72 2.634 9.745 2.781 ;
      RECT 9.715 2.639 9.72 2.786 ;
      RECT 9.685 2.642 9.715 2.79 ;
      RECT 9.645 2.645 9.685 2.8 ;
      RECT 9.61 2.642 9.645 2.812 ;
      RECT 9.6 2.638 9.61 2.819 ;
      RECT 9.575 2.634 9.6 2.825 ;
      RECT 9.57 2.63 9.575 2.83 ;
      RECT 9.53 2.627 9.57 2.83 ;
      RECT 9.515 2.612 9.53 2.831 ;
      RECT 9.492 2.6 9.515 2.831 ;
      RECT 9.406 2.6 9.492 2.832 ;
      RECT 9.32 2.6 9.406 2.834 ;
      RECT 9.3 2.6 9.32 2.831 ;
      RECT 9.295 2.605 9.3 2.826 ;
      RECT 9.29 2.61 9.295 2.824 ;
      RECT 9.28 2.62 9.29 2.822 ;
      RECT 9.275 2.626 9.28 2.815 ;
      RECT 9.27 2.628 9.275 2.8 ;
      RECT 9.265 2.632 9.27 2.79 ;
      RECT 10.725 2.1 10.975 2.36 ;
      RECT 8.45 3.635 8.71 3.895 ;
      RECT 10.745 3.125 10.75 3.335 ;
      RECT 10.75 3.13 10.76 3.33 ;
      RECT 10.7 3.125 10.745 3.35 ;
      RECT 10.69 3.125 10.7 3.37 ;
      RECT 10.671 3.125 10.69 3.375 ;
      RECT 10.585 3.125 10.671 3.372 ;
      RECT 10.555 3.127 10.585 3.37 ;
      RECT 10.5 3.137 10.555 3.368 ;
      RECT 10.435 3.151 10.5 3.366 ;
      RECT 10.43 3.159 10.435 3.365 ;
      RECT 10.415 3.162 10.43 3.363 ;
      RECT 10.35 3.172 10.415 3.359 ;
      RECT 10.302 3.186 10.35 3.36 ;
      RECT 10.216 3.203 10.302 3.374 ;
      RECT 10.13 3.224 10.216 3.391 ;
      RECT 10.11 3.237 10.13 3.401 ;
      RECT 10.065 3.245 10.11 3.408 ;
      RECT 10.03 3.253 10.065 3.416 ;
      RECT 9.996 3.261 10.03 3.424 ;
      RECT 9.91 3.275 9.996 3.436 ;
      RECT 9.875 3.292 9.91 3.448 ;
      RECT 9.866 3.301 9.875 3.452 ;
      RECT 9.78 3.319 9.866 3.469 ;
      RECT 9.721 3.346 9.78 3.496 ;
      RECT 9.635 3.373 9.721 3.524 ;
      RECT 9.615 3.395 9.635 3.544 ;
      RECT 9.555 3.41 9.615 3.56 ;
      RECT 9.545 3.422 9.555 3.573 ;
      RECT 9.54 3.427 9.545 3.576 ;
      RECT 9.53 3.43 9.54 3.579 ;
      RECT 9.525 3.432 9.53 3.582 ;
      RECT 9.495 3.44 9.525 3.589 ;
      RECT 9.48 3.447 9.495 3.597 ;
      RECT 9.47 3.452 9.48 3.601 ;
      RECT 9.465 3.455 9.47 3.604 ;
      RECT 9.455 3.457 9.465 3.607 ;
      RECT 9.42 3.467 9.455 3.616 ;
      RECT 9.345 3.49 9.42 3.638 ;
      RECT 9.325 3.508 9.345 3.656 ;
      RECT 9.295 3.515 9.325 3.666 ;
      RECT 9.275 3.523 9.295 3.676 ;
      RECT 9.265 3.529 9.275 3.683 ;
      RECT 9.246 3.534 9.265 3.689 ;
      RECT 9.16 3.554 9.246 3.709 ;
      RECT 9.145 3.574 9.16 3.728 ;
      RECT 9.1 3.586 9.145 3.739 ;
      RECT 9.035 3.607 9.1 3.762 ;
      RECT 8.995 3.627 9.035 3.783 ;
      RECT 8.985 3.637 8.995 3.793 ;
      RECT 8.935 3.649 8.985 3.804 ;
      RECT 8.915 3.665 8.935 3.816 ;
      RECT 8.885 3.675 8.915 3.822 ;
      RECT 8.875 3.68 8.885 3.824 ;
      RECT 8.806 3.681 8.875 3.83 ;
      RECT 8.72 3.683 8.806 3.84 ;
      RECT 8.71 3.684 8.72 3.845 ;
      RECT 9.98 3.71 10.17 3.92 ;
      RECT 9.97 3.715 10.18 3.913 ;
      RECT 9.955 3.715 10.18 3.878 ;
      RECT 9.875 3.6 10.135 3.86 ;
      RECT 8.79 3.13 8.975 3.425 ;
      RECT 8.78 3.13 8.975 3.423 ;
      RECT 8.765 3.13 8.98 3.418 ;
      RECT 8.765 3.13 8.985 3.415 ;
      RECT 8.76 3.13 8.985 3.413 ;
      RECT 8.755 3.385 8.985 3.403 ;
      RECT 8.76 3.13 9.02 3.39 ;
      RECT 8.72 2.165 8.98 2.425 ;
      RECT 8.53 2.09 8.616 2.423 ;
      RECT 8.505 2.094 8.66 2.419 ;
      RECT 8.616 2.086 8.66 2.419 ;
      RECT 8.616 2.087 8.665 2.418 ;
      RECT 8.53 2.092 8.68 2.417 ;
      RECT 8.505 2.1 8.72 2.416 ;
      RECT 8.5 2.095 8.68 2.411 ;
      RECT 8.49 2.11 8.72 2.318 ;
      RECT 8.49 2.162 8.92 2.318 ;
      RECT 8.49 2.155 8.9 2.318 ;
      RECT 8.49 2.142 8.87 2.318 ;
      RECT 8.49 2.13 8.81 2.318 ;
      RECT 8.49 2.115 8.785 2.318 ;
      RECT 7.69 2.745 7.825 3.04 ;
      RECT 7.95 2.768 7.955 2.955 ;
      RECT 8.67 2.665 8.815 2.9 ;
      RECT 8.83 2.665 8.835 2.89 ;
      RECT 8.865 2.676 8.87 2.87 ;
      RECT 8.86 2.668 8.865 2.875 ;
      RECT 8.84 2.665 8.86 2.88 ;
      RECT 8.835 2.665 8.84 2.888 ;
      RECT 8.825 2.665 8.83 2.893 ;
      RECT 8.815 2.665 8.825 2.898 ;
      RECT 8.645 2.667 8.67 2.9 ;
      RECT 8.595 2.674 8.645 2.9 ;
      RECT 8.59 2.679 8.595 2.9 ;
      RECT 8.551 2.684 8.59 2.901 ;
      RECT 8.465 2.696 8.551 2.902 ;
      RECT 8.456 2.706 8.465 2.902 ;
      RECT 8.37 2.715 8.456 2.904 ;
      RECT 8.346 2.725 8.37 2.906 ;
      RECT 8.26 2.736 8.346 2.907 ;
      RECT 8.23 2.747 8.26 2.909 ;
      RECT 8.2 2.752 8.23 2.911 ;
      RECT 8.175 2.758 8.2 2.914 ;
      RECT 8.16 2.763 8.175 2.915 ;
      RECT 8.115 2.769 8.16 2.915 ;
      RECT 8.11 2.774 8.115 2.916 ;
      RECT 8.09 2.774 8.11 2.918 ;
      RECT 8.07 2.772 8.09 2.923 ;
      RECT 8.035 2.771 8.07 2.93 ;
      RECT 8.005 2.77 8.035 2.94 ;
      RECT 7.955 2.769 8.005 2.95 ;
      RECT 7.865 2.766 7.95 3.04 ;
      RECT 7.84 2.76 7.865 3.04 ;
      RECT 7.825 2.75 7.84 3.04 ;
      RECT 7.64 2.745 7.69 2.96 ;
      RECT 7.63 2.75 7.64 2.95 ;
      RECT 7.87 3.225 8.13 3.485 ;
      RECT 7.87 3.225 8.16 3.378 ;
      RECT 7.87 3.225 8.195 3.363 ;
      RECT 8.125 3.145 8.315 3.355 ;
      RECT 8.115 3.15 8.325 3.348 ;
      RECT 8.08 3.22 8.325 3.348 ;
      RECT 8.11 3.162 8.13 3.485 ;
      RECT 8.095 3.21 8.325 3.348 ;
      RECT 8.1 3.182 8.13 3.485 ;
      RECT 7.18 2.25 7.25 3.355 ;
      RECT 7.915 2.355 8.175 2.615 ;
      RECT 7.495 2.401 7.51 2.61 ;
      RECT 7.831 2.414 7.915 2.565 ;
      RECT 7.745 2.411 7.831 2.565 ;
      RECT 7.706 2.409 7.745 2.565 ;
      RECT 7.62 2.407 7.706 2.565 ;
      RECT 7.56 2.405 7.62 2.576 ;
      RECT 7.525 2.403 7.56 2.594 ;
      RECT 7.51 2.401 7.525 2.605 ;
      RECT 7.48 2.401 7.495 2.618 ;
      RECT 7.47 2.401 7.48 2.623 ;
      RECT 7.445 2.4 7.47 2.628 ;
      RECT 7.43 2.395 7.445 2.634 ;
      RECT 7.425 2.388 7.43 2.639 ;
      RECT 7.4 2.379 7.425 2.645 ;
      RECT 7.355 2.358 7.4 2.658 ;
      RECT 7.345 2.342 7.355 2.668 ;
      RECT 7.33 2.335 7.345 2.678 ;
      RECT 7.32 2.328 7.33 2.695 ;
      RECT 7.315 2.325 7.32 2.725 ;
      RECT 7.31 2.323 7.315 2.755 ;
      RECT 7.305 2.321 7.31 2.792 ;
      RECT 7.29 2.317 7.305 2.859 ;
      RECT 7.29 3.15 7.3 3.35 ;
      RECT 7.285 2.313 7.29 2.985 ;
      RECT 7.285 3.137 7.29 3.355 ;
      RECT 7.28 2.311 7.285 3.07 ;
      RECT 7.28 3.127 7.285 3.355 ;
      RECT 7.265 2.282 7.28 3.355 ;
      RECT 7.25 2.255 7.265 3.355 ;
      RECT 7.175 2.25 7.18 2.605 ;
      RECT 7.175 2.66 7.18 3.355 ;
      RECT 7.16 2.25 7.175 2.583 ;
      RECT 7.17 2.682 7.175 3.355 ;
      RECT 7.16 2.722 7.17 3.355 ;
      RECT 7.125 2.25 7.16 2.525 ;
      RECT 7.155 2.757 7.16 3.355 ;
      RECT 7.14 2.812 7.155 3.355 ;
      RECT 7.135 2.877 7.14 3.355 ;
      RECT 7.12 2.925 7.135 3.355 ;
      RECT 7.095 2.25 7.125 2.48 ;
      RECT 7.115 2.98 7.12 3.355 ;
      RECT 7.1 3.04 7.115 3.355 ;
      RECT 7.095 3.088 7.1 3.353 ;
      RECT 7.09 2.25 7.095 2.473 ;
      RECT 7.09 3.12 7.095 3.348 ;
      RECT 7.065 2.25 7.09 2.465 ;
      RECT 7.055 2.255 7.065 2.455 ;
      RECT 7.27 3.53 7.29 3.77 ;
      RECT 6.5 3.46 6.505 3.67 ;
      RECT 7.78 3.533 7.79 3.728 ;
      RECT 7.775 3.523 7.78 3.731 ;
      RECT 7.695 3.52 7.775 3.754 ;
      RECT 7.691 3.52 7.695 3.776 ;
      RECT 7.605 3.52 7.691 3.786 ;
      RECT 7.59 3.52 7.605 3.794 ;
      RECT 7.561 3.521 7.59 3.792 ;
      RECT 7.475 3.526 7.561 3.788 ;
      RECT 7.462 3.53 7.475 3.784 ;
      RECT 7.376 3.53 7.462 3.78 ;
      RECT 7.29 3.53 7.376 3.774 ;
      RECT 7.206 3.53 7.27 3.768 ;
      RECT 7.12 3.53 7.206 3.763 ;
      RECT 7.1 3.53 7.12 3.759 ;
      RECT 7.04 3.525 7.1 3.756 ;
      RECT 7.012 3.519 7.04 3.753 ;
      RECT 6.926 3.514 7.012 3.749 ;
      RECT 6.84 3.508 6.926 3.743 ;
      RECT 6.765 3.49 6.84 3.738 ;
      RECT 6.73 3.467 6.765 3.734 ;
      RECT 6.72 3.457 6.73 3.733 ;
      RECT 6.665 3.455 6.72 3.732 ;
      RECT 6.59 3.455 6.665 3.728 ;
      RECT 6.58 3.455 6.59 3.723 ;
      RECT 6.565 3.455 6.58 3.715 ;
      RECT 6.515 3.457 6.565 3.693 ;
      RECT 6.505 3.46 6.515 3.673 ;
      RECT 6.495 3.465 6.5 3.668 ;
      RECT 6.49 3.47 6.495 3.663 ;
      RECT 6.615 2.635 6.875 2.895 ;
      RECT 6.615 2.65 6.895 2.86 ;
      RECT 6.615 2.655 6.905 2.855 ;
      RECT 4.6 2.115 4.86 2.375 ;
      RECT 4.59 2.145 4.86 2.355 ;
      RECT 6.51 2.06 6.77 2.32 ;
      RECT 6.505 2.135 6.51 2.321 ;
      RECT 6.48 2.14 6.505 2.323 ;
      RECT 6.465 2.147 6.48 2.326 ;
      RECT 6.405 2.165 6.465 2.331 ;
      RECT 6.375 2.185 6.405 2.338 ;
      RECT 6.35 2.193 6.375 2.343 ;
      RECT 6.325 2.201 6.35 2.345 ;
      RECT 6.307 2.205 6.325 2.344 ;
      RECT 6.221 2.203 6.307 2.344 ;
      RECT 6.135 2.201 6.221 2.344 ;
      RECT 6.049 2.199 6.135 2.343 ;
      RECT 5.963 2.197 6.049 2.343 ;
      RECT 5.877 2.195 5.963 2.343 ;
      RECT 5.791 2.193 5.877 2.343 ;
      RECT 5.705 2.191 5.791 2.342 ;
      RECT 5.687 2.19 5.705 2.342 ;
      RECT 5.601 2.189 5.687 2.342 ;
      RECT 5.515 2.187 5.601 2.342 ;
      RECT 5.429 2.186 5.515 2.341 ;
      RECT 5.343 2.185 5.429 2.341 ;
      RECT 5.257 2.183 5.343 2.341 ;
      RECT 5.171 2.182 5.257 2.341 ;
      RECT 5.085 2.18 5.171 2.34 ;
      RECT 5.061 2.178 5.085 2.34 ;
      RECT 4.975 2.171 5.061 2.34 ;
      RECT 4.946 2.163 4.975 2.34 ;
      RECT 4.86 2.155 4.946 2.34 ;
      RECT 4.58 2.152 4.59 2.35 ;
      RECT 6.085 3.115 6.09 3.465 ;
      RECT 5.855 3.205 5.995 3.465 ;
      RECT 6.33 2.89 6.375 3.1 ;
      RECT 6.385 2.901 6.395 3.095 ;
      RECT 6.375 2.893 6.385 3.1 ;
      RECT 6.31 2.89 6.33 3.105 ;
      RECT 6.28 2.89 6.31 3.128 ;
      RECT 6.27 2.89 6.28 3.153 ;
      RECT 6.265 2.89 6.27 3.163 ;
      RECT 6.21 2.89 6.265 3.203 ;
      RECT 6.205 2.89 6.21 3.243 ;
      RECT 6.2 2.892 6.205 3.248 ;
      RECT 6.185 2.902 6.2 3.259 ;
      RECT 6.14 2.96 6.185 3.295 ;
      RECT 6.13 3.015 6.14 3.329 ;
      RECT 6.115 3.042 6.13 3.345 ;
      RECT 6.105 3.069 6.115 3.465 ;
      RECT 6.09 3.092 6.105 3.465 ;
      RECT 6.08 3.132 6.085 3.465 ;
      RECT 6.075 3.142 6.08 3.465 ;
      RECT 6.07 3.157 6.075 3.465 ;
      RECT 6.06 3.162 6.07 3.465 ;
      RECT 5.995 3.185 6.06 3.465 ;
      RECT 5.495 2.68 5.685 2.89 ;
      RECT 4.07 2.605 4.33 2.865 ;
      RECT 4.42 2.6 4.515 2.81 ;
      RECT 4.395 2.615 4.405 2.81 ;
      RECT 5.685 2.687 5.695 2.885 ;
      RECT 5.485 2.687 5.495 2.885 ;
      RECT 5.47 2.702 5.485 2.875 ;
      RECT 5.465 2.71 5.47 2.868 ;
      RECT 5.455 2.713 5.465 2.865 ;
      RECT 5.42 2.712 5.455 2.863 ;
      RECT 5.391 2.708 5.42 2.86 ;
      RECT 5.305 2.703 5.391 2.857 ;
      RECT 5.245 2.697 5.305 2.853 ;
      RECT 5.216 2.693 5.245 2.85 ;
      RECT 5.13 2.685 5.216 2.847 ;
      RECT 5.121 2.679 5.13 2.845 ;
      RECT 5.035 2.674 5.121 2.843 ;
      RECT 5.012 2.669 5.035 2.84 ;
      RECT 4.926 2.663 5.012 2.837 ;
      RECT 4.84 2.654 4.926 2.832 ;
      RECT 4.83 2.649 4.84 2.83 ;
      RECT 4.811 2.648 4.83 2.829 ;
      RECT 4.725 2.643 4.811 2.825 ;
      RECT 4.705 2.638 4.725 2.821 ;
      RECT 4.645 2.633 4.705 2.818 ;
      RECT 4.62 2.623 4.645 2.816 ;
      RECT 4.615 2.616 4.62 2.815 ;
      RECT 4.605 2.607 4.615 2.814 ;
      RECT 4.601 2.6 4.605 2.814 ;
      RECT 4.515 2.6 4.601 2.812 ;
      RECT 4.405 2.607 4.42 2.81 ;
      RECT 4.39 2.617 4.395 2.81 ;
      RECT 4.37 2.62 4.39 2.807 ;
      RECT 4.34 2.62 4.37 2.803 ;
      RECT 4.33 2.62 4.34 2.803 ;
      RECT 5.245 3.115 5.505 3.375 ;
      RECT 5.175 3.125 5.505 3.335 ;
      RECT 5.165 3.132 5.505 3.33 ;
      RECT 4.585 3.12 4.845 3.38 ;
      RECT 4.585 3.16 4.95 3.37 ;
      RECT 4.585 3.162 4.955 3.369 ;
      RECT 4.585 3.17 4.96 3.366 ;
      RECT 3.51 2.245 3.61 3.77 ;
      RECT 3.7 3.385 3.75 3.645 ;
      RECT 3.695 2.258 3.7 2.445 ;
      RECT 3.69 3.366 3.7 3.645 ;
      RECT 3.69 2.255 3.695 2.453 ;
      RECT 3.675 2.249 3.69 2.46 ;
      RECT 3.685 3.354 3.69 3.728 ;
      RECT 3.675 3.342 3.685 3.765 ;
      RECT 3.665 2.245 3.675 2.467 ;
      RECT 3.665 3.327 3.675 3.77 ;
      RECT 3.66 2.245 3.665 2.475 ;
      RECT 3.64 3.297 3.665 3.77 ;
      RECT 3.62 2.245 3.66 2.523 ;
      RECT 3.63 3.257 3.64 3.77 ;
      RECT 3.62 3.212 3.63 3.77 ;
      RECT 3.615 2.245 3.62 2.593 ;
      RECT 3.615 3.17 3.62 3.77 ;
      RECT 3.61 2.245 3.615 3.07 ;
      RECT 3.61 3.152 3.615 3.77 ;
      RECT 3.5 2.248 3.51 3.77 ;
      RECT 3.485 2.255 3.5 3.766 ;
      RECT 3.48 2.265 3.485 3.761 ;
      RECT 3.475 2.465 3.48 3.653 ;
      RECT 3.47 2.55 3.475 3.205 ;
      RECT 1.7 7.765 1.99 7.995 ;
      RECT 1.76 7.025 1.93 7.995 ;
      RECT 1.67 7.025 2.02 7.315 ;
      RECT 1.295 6.285 1.645 6.575 ;
      RECT 1.155 6.315 1.645 6.485 ;
      RECT 87.2 1.14 87.575 1.51 ;
      RECT 81.18 2.225 81.44 2.485 ;
      RECT 69.275 1.14 69.65 1.51 ;
      RECT 63.255 2.225 63.515 2.485 ;
      RECT 51.35 1.14 51.725 1.51 ;
      RECT 45.33 2.225 45.59 2.485 ;
      RECT 33.425 1.14 33.8 1.51 ;
      RECT 27.405 2.225 27.665 2.485 ;
      RECT 15.5 1.14 15.875 1.51 ;
      RECT 9.48 2.225 9.74 2.485 ;
    LAYER mcon ;
      RECT 92.03 6.32 92.2 6.49 ;
      RECT 92.035 6.315 92.205 6.485 ;
      RECT 74.105 6.32 74.275 6.49 ;
      RECT 74.11 6.315 74.28 6.485 ;
      RECT 56.18 6.32 56.35 6.49 ;
      RECT 56.185 6.315 56.355 6.485 ;
      RECT 38.255 6.32 38.425 6.49 ;
      RECT 38.26 6.315 38.43 6.485 ;
      RECT 20.33 6.32 20.5 6.49 ;
      RECT 20.335 6.315 20.505 6.485 ;
      RECT 92.03 7.8 92.2 7.97 ;
      RECT 91.68 0.1 91.85 0.27 ;
      RECT 91.68 8.61 91.85 8.78 ;
      RECT 91.66 2.76 91.83 2.93 ;
      RECT 91.66 5.95 91.83 6.12 ;
      RECT 91.04 0.91 91.21 1.08 ;
      RECT 91.04 2.39 91.21 2.56 ;
      RECT 91.04 6.32 91.21 6.49 ;
      RECT 91.04 7.8 91.21 7.97 ;
      RECT 90.69 0.1 90.86 0.27 ;
      RECT 90.69 8.61 90.86 8.78 ;
      RECT 90.67 2.76 90.84 2.93 ;
      RECT 90.67 5.95 90.84 6.12 ;
      RECT 89.99 0.105 90.16 0.275 ;
      RECT 89.99 8.605 90.16 8.775 ;
      RECT 89.68 2.025 89.85 2.195 ;
      RECT 89.68 6.685 89.85 6.855 ;
      RECT 89.31 0.105 89.48 0.275 ;
      RECT 89.31 8.605 89.48 8.775 ;
      RECT 89.25 0.915 89.42 1.085 ;
      RECT 89.25 1.655 89.42 1.825 ;
      RECT 89.25 7.055 89.42 7.225 ;
      RECT 89.25 7.795 89.42 7.965 ;
      RECT 88.875 2.395 89.045 2.565 ;
      RECT 88.875 6.315 89.045 6.485 ;
      RECT 88.63 0.105 88.8 0.275 ;
      RECT 88.63 8.605 88.8 8.775 ;
      RECT 87.95 0.105 88.12 0.275 ;
      RECT 87.95 8.605 88.12 8.775 ;
      RECT 86.67 1.565 86.84 1.735 ;
      RECT 86.21 1.565 86.38 1.735 ;
      RECT 85.815 2.905 85.985 3.075 ;
      RECT 85.75 1.565 85.92 1.735 ;
      RECT 85.605 2.245 85.775 2.415 ;
      RECT 85.29 1.565 85.46 1.735 ;
      RECT 85.29 3.155 85.46 3.325 ;
      RECT 85.23 8.605 85.4 8.775 ;
      RECT 84.92 6.685 85.09 6.855 ;
      RECT 84.905 2.75 85.075 2.92 ;
      RECT 84.83 1.565 85 1.735 ;
      RECT 84.69 3.315 84.86 3.485 ;
      RECT 84.67 3.715 84.84 3.885 ;
      RECT 84.55 8.605 84.72 8.775 ;
      RECT 84.495 2.27 84.665 2.44 ;
      RECT 84.49 7.055 84.66 7.225 ;
      RECT 84.49 7.795 84.66 7.965 ;
      RECT 84.37 1.565 84.54 1.735 ;
      RECT 84.115 6.315 84.285 6.485 ;
      RECT 84 3.25 84.17 3.42 ;
      RECT 83.91 1.565 84.08 1.735 ;
      RECT 83.87 8.605 84.04 8.775 ;
      RECT 83.675 2.935 83.845 3.105 ;
      RECT 83.61 3.715 83.78 3.885 ;
      RECT 83.45 1.565 83.62 1.735 ;
      RECT 83.21 3.7 83.38 3.87 ;
      RECT 83.19 8.605 83.36 8.775 ;
      RECT 83.17 2.185 83.34 2.355 ;
      RECT 82.99 1.565 83.16 1.735 ;
      RECT 82.53 1.565 82.7 1.735 ;
      RECT 82.27 2.685 82.44 2.855 ;
      RECT 82.27 3.145 82.44 3.315 ;
      RECT 82.27 3.66 82.44 3.83 ;
      RECT 82.155 2.22 82.325 2.39 ;
      RECT 82.07 1.565 82.24 1.735 ;
      RECT 81.69 3.73 81.86 3.9 ;
      RECT 81.61 1.565 81.78 1.735 ;
      RECT 81.21 2.26 81.38 2.43 ;
      RECT 81.15 1.565 81.32 1.735 ;
      RECT 80.995 2.635 81.165 2.805 ;
      RECT 80.69 1.565 80.86 1.735 ;
      RECT 80.495 3.235 80.665 3.405 ;
      RECT 80.38 2.685 80.55 2.855 ;
      RECT 80.23 1.565 80.4 1.735 ;
      RECT 80.21 2.135 80.38 2.305 ;
      RECT 79.835 3.165 80.005 3.335 ;
      RECT 79.77 1.565 79.94 1.735 ;
      RECT 79.35 2.765 79.52 2.935 ;
      RECT 79.31 1.565 79.48 1.735 ;
      RECT 79.3 3.54 79.47 3.71 ;
      RECT 78.85 1.565 79.02 1.735 ;
      RECT 78.81 3.165 78.98 3.335 ;
      RECT 78.775 2.27 78.945 2.44 ;
      RECT 78.415 2.67 78.585 2.84 ;
      RECT 78.39 1.565 78.56 1.735 ;
      RECT 78.21 3.48 78.38 3.65 ;
      RECT 77.93 1.565 78.1 1.735 ;
      RECT 77.905 2.91 78.075 3.08 ;
      RECT 77.47 1.565 77.64 1.735 ;
      RECT 77.205 2.7 77.375 2.87 ;
      RECT 77.01 1.565 77.18 1.735 ;
      RECT 76.885 3.145 77.055 3.315 ;
      RECT 76.55 1.565 76.72 1.735 ;
      RECT 76.47 3.18 76.64 3.35 ;
      RECT 76.3 2.165 76.47 2.335 ;
      RECT 76.125 2.62 76.295 2.79 ;
      RECT 76.09 1.565 76.26 1.735 ;
      RECT 75.63 1.565 75.8 1.735 ;
      RECT 75.205 2.27 75.375 2.44 ;
      RECT 75.2 3.585 75.37 3.755 ;
      RECT 75.17 1.565 75.34 1.735 ;
      RECT 74.105 7.8 74.275 7.97 ;
      RECT 73.755 0.1 73.925 0.27 ;
      RECT 73.755 8.61 73.925 8.78 ;
      RECT 73.735 2.76 73.905 2.93 ;
      RECT 73.735 5.95 73.905 6.12 ;
      RECT 73.115 0.91 73.285 1.08 ;
      RECT 73.115 2.39 73.285 2.56 ;
      RECT 73.115 6.32 73.285 6.49 ;
      RECT 73.115 7.8 73.285 7.97 ;
      RECT 72.765 0.1 72.935 0.27 ;
      RECT 72.765 8.61 72.935 8.78 ;
      RECT 72.745 2.76 72.915 2.93 ;
      RECT 72.745 5.95 72.915 6.12 ;
      RECT 72.065 0.105 72.235 0.275 ;
      RECT 72.065 8.605 72.235 8.775 ;
      RECT 71.755 2.025 71.925 2.195 ;
      RECT 71.755 6.685 71.925 6.855 ;
      RECT 71.385 0.105 71.555 0.275 ;
      RECT 71.385 8.605 71.555 8.775 ;
      RECT 71.325 0.915 71.495 1.085 ;
      RECT 71.325 1.655 71.495 1.825 ;
      RECT 71.325 7.055 71.495 7.225 ;
      RECT 71.325 7.795 71.495 7.965 ;
      RECT 70.95 2.395 71.12 2.565 ;
      RECT 70.95 6.315 71.12 6.485 ;
      RECT 70.705 0.105 70.875 0.275 ;
      RECT 70.705 8.605 70.875 8.775 ;
      RECT 70.025 0.105 70.195 0.275 ;
      RECT 70.025 8.605 70.195 8.775 ;
      RECT 68.745 1.565 68.915 1.735 ;
      RECT 68.285 1.565 68.455 1.735 ;
      RECT 67.89 2.905 68.06 3.075 ;
      RECT 67.825 1.565 67.995 1.735 ;
      RECT 67.68 2.245 67.85 2.415 ;
      RECT 67.365 1.565 67.535 1.735 ;
      RECT 67.365 3.155 67.535 3.325 ;
      RECT 67.305 8.605 67.475 8.775 ;
      RECT 66.995 6.685 67.165 6.855 ;
      RECT 66.98 2.75 67.15 2.92 ;
      RECT 66.905 1.565 67.075 1.735 ;
      RECT 66.765 3.315 66.935 3.485 ;
      RECT 66.745 3.715 66.915 3.885 ;
      RECT 66.625 8.605 66.795 8.775 ;
      RECT 66.57 2.27 66.74 2.44 ;
      RECT 66.565 7.055 66.735 7.225 ;
      RECT 66.565 7.795 66.735 7.965 ;
      RECT 66.445 1.565 66.615 1.735 ;
      RECT 66.19 6.315 66.36 6.485 ;
      RECT 66.075 3.25 66.245 3.42 ;
      RECT 65.985 1.565 66.155 1.735 ;
      RECT 65.945 8.605 66.115 8.775 ;
      RECT 65.75 2.935 65.92 3.105 ;
      RECT 65.685 3.715 65.855 3.885 ;
      RECT 65.525 1.565 65.695 1.735 ;
      RECT 65.285 3.7 65.455 3.87 ;
      RECT 65.265 8.605 65.435 8.775 ;
      RECT 65.245 2.185 65.415 2.355 ;
      RECT 65.065 1.565 65.235 1.735 ;
      RECT 64.605 1.565 64.775 1.735 ;
      RECT 64.345 2.685 64.515 2.855 ;
      RECT 64.345 3.145 64.515 3.315 ;
      RECT 64.345 3.66 64.515 3.83 ;
      RECT 64.23 2.22 64.4 2.39 ;
      RECT 64.145 1.565 64.315 1.735 ;
      RECT 63.765 3.73 63.935 3.9 ;
      RECT 63.685 1.565 63.855 1.735 ;
      RECT 63.285 2.26 63.455 2.43 ;
      RECT 63.225 1.565 63.395 1.735 ;
      RECT 63.07 2.635 63.24 2.805 ;
      RECT 62.765 1.565 62.935 1.735 ;
      RECT 62.57 3.235 62.74 3.405 ;
      RECT 62.455 2.685 62.625 2.855 ;
      RECT 62.305 1.565 62.475 1.735 ;
      RECT 62.285 2.135 62.455 2.305 ;
      RECT 61.91 3.165 62.08 3.335 ;
      RECT 61.845 1.565 62.015 1.735 ;
      RECT 61.425 2.765 61.595 2.935 ;
      RECT 61.385 1.565 61.555 1.735 ;
      RECT 61.375 3.54 61.545 3.71 ;
      RECT 60.925 1.565 61.095 1.735 ;
      RECT 60.885 3.165 61.055 3.335 ;
      RECT 60.85 2.27 61.02 2.44 ;
      RECT 60.49 2.67 60.66 2.84 ;
      RECT 60.465 1.565 60.635 1.735 ;
      RECT 60.285 3.48 60.455 3.65 ;
      RECT 60.005 1.565 60.175 1.735 ;
      RECT 59.98 2.91 60.15 3.08 ;
      RECT 59.545 1.565 59.715 1.735 ;
      RECT 59.28 2.7 59.45 2.87 ;
      RECT 59.085 1.565 59.255 1.735 ;
      RECT 58.96 3.145 59.13 3.315 ;
      RECT 58.625 1.565 58.795 1.735 ;
      RECT 58.545 3.18 58.715 3.35 ;
      RECT 58.375 2.165 58.545 2.335 ;
      RECT 58.2 2.62 58.37 2.79 ;
      RECT 58.165 1.565 58.335 1.735 ;
      RECT 57.705 1.565 57.875 1.735 ;
      RECT 57.28 2.27 57.45 2.44 ;
      RECT 57.275 3.585 57.445 3.755 ;
      RECT 57.245 1.565 57.415 1.735 ;
      RECT 56.18 7.8 56.35 7.97 ;
      RECT 55.83 0.1 56 0.27 ;
      RECT 55.83 8.61 56 8.78 ;
      RECT 55.81 2.76 55.98 2.93 ;
      RECT 55.81 5.95 55.98 6.12 ;
      RECT 55.19 0.91 55.36 1.08 ;
      RECT 55.19 2.39 55.36 2.56 ;
      RECT 55.19 6.32 55.36 6.49 ;
      RECT 55.19 7.8 55.36 7.97 ;
      RECT 54.84 0.1 55.01 0.27 ;
      RECT 54.84 8.61 55.01 8.78 ;
      RECT 54.82 2.76 54.99 2.93 ;
      RECT 54.82 5.95 54.99 6.12 ;
      RECT 54.14 0.105 54.31 0.275 ;
      RECT 54.14 8.605 54.31 8.775 ;
      RECT 53.83 2.025 54 2.195 ;
      RECT 53.83 6.685 54 6.855 ;
      RECT 53.46 0.105 53.63 0.275 ;
      RECT 53.46 8.605 53.63 8.775 ;
      RECT 53.4 0.915 53.57 1.085 ;
      RECT 53.4 1.655 53.57 1.825 ;
      RECT 53.4 7.055 53.57 7.225 ;
      RECT 53.4 7.795 53.57 7.965 ;
      RECT 53.025 2.395 53.195 2.565 ;
      RECT 53.025 6.315 53.195 6.485 ;
      RECT 52.78 0.105 52.95 0.275 ;
      RECT 52.78 8.605 52.95 8.775 ;
      RECT 52.1 0.105 52.27 0.275 ;
      RECT 52.1 8.605 52.27 8.775 ;
      RECT 50.82 1.565 50.99 1.735 ;
      RECT 50.36 1.565 50.53 1.735 ;
      RECT 49.965 2.905 50.135 3.075 ;
      RECT 49.9 1.565 50.07 1.735 ;
      RECT 49.755 2.245 49.925 2.415 ;
      RECT 49.44 1.565 49.61 1.735 ;
      RECT 49.44 3.155 49.61 3.325 ;
      RECT 49.38 8.605 49.55 8.775 ;
      RECT 49.07 6.685 49.24 6.855 ;
      RECT 49.055 2.75 49.225 2.92 ;
      RECT 48.98 1.565 49.15 1.735 ;
      RECT 48.84 3.315 49.01 3.485 ;
      RECT 48.82 3.715 48.99 3.885 ;
      RECT 48.7 8.605 48.87 8.775 ;
      RECT 48.645 2.27 48.815 2.44 ;
      RECT 48.64 7.055 48.81 7.225 ;
      RECT 48.64 7.795 48.81 7.965 ;
      RECT 48.52 1.565 48.69 1.735 ;
      RECT 48.265 6.315 48.435 6.485 ;
      RECT 48.15 3.25 48.32 3.42 ;
      RECT 48.06 1.565 48.23 1.735 ;
      RECT 48.02 8.605 48.19 8.775 ;
      RECT 47.825 2.935 47.995 3.105 ;
      RECT 47.76 3.715 47.93 3.885 ;
      RECT 47.6 1.565 47.77 1.735 ;
      RECT 47.36 3.7 47.53 3.87 ;
      RECT 47.34 8.605 47.51 8.775 ;
      RECT 47.32 2.185 47.49 2.355 ;
      RECT 47.14 1.565 47.31 1.735 ;
      RECT 46.68 1.565 46.85 1.735 ;
      RECT 46.42 2.685 46.59 2.855 ;
      RECT 46.42 3.145 46.59 3.315 ;
      RECT 46.42 3.66 46.59 3.83 ;
      RECT 46.305 2.22 46.475 2.39 ;
      RECT 46.22 1.565 46.39 1.735 ;
      RECT 45.84 3.73 46.01 3.9 ;
      RECT 45.76 1.565 45.93 1.735 ;
      RECT 45.36 2.26 45.53 2.43 ;
      RECT 45.3 1.565 45.47 1.735 ;
      RECT 45.145 2.635 45.315 2.805 ;
      RECT 44.84 1.565 45.01 1.735 ;
      RECT 44.645 3.235 44.815 3.405 ;
      RECT 44.53 2.685 44.7 2.855 ;
      RECT 44.38 1.565 44.55 1.735 ;
      RECT 44.36 2.135 44.53 2.305 ;
      RECT 43.985 3.165 44.155 3.335 ;
      RECT 43.92 1.565 44.09 1.735 ;
      RECT 43.5 2.765 43.67 2.935 ;
      RECT 43.46 1.565 43.63 1.735 ;
      RECT 43.45 3.54 43.62 3.71 ;
      RECT 43 1.565 43.17 1.735 ;
      RECT 42.96 3.165 43.13 3.335 ;
      RECT 42.925 2.27 43.095 2.44 ;
      RECT 42.565 2.67 42.735 2.84 ;
      RECT 42.54 1.565 42.71 1.735 ;
      RECT 42.36 3.48 42.53 3.65 ;
      RECT 42.08 1.565 42.25 1.735 ;
      RECT 42.055 2.91 42.225 3.08 ;
      RECT 41.62 1.565 41.79 1.735 ;
      RECT 41.355 2.7 41.525 2.87 ;
      RECT 41.16 1.565 41.33 1.735 ;
      RECT 41.035 3.145 41.205 3.315 ;
      RECT 40.7 1.565 40.87 1.735 ;
      RECT 40.62 3.18 40.79 3.35 ;
      RECT 40.45 2.165 40.62 2.335 ;
      RECT 40.275 2.62 40.445 2.79 ;
      RECT 40.24 1.565 40.41 1.735 ;
      RECT 39.78 1.565 39.95 1.735 ;
      RECT 39.355 2.27 39.525 2.44 ;
      RECT 39.35 3.585 39.52 3.755 ;
      RECT 39.32 1.565 39.49 1.735 ;
      RECT 38.255 7.8 38.425 7.97 ;
      RECT 37.905 0.1 38.075 0.27 ;
      RECT 37.905 8.61 38.075 8.78 ;
      RECT 37.885 2.76 38.055 2.93 ;
      RECT 37.885 5.95 38.055 6.12 ;
      RECT 37.265 0.91 37.435 1.08 ;
      RECT 37.265 2.39 37.435 2.56 ;
      RECT 37.265 6.32 37.435 6.49 ;
      RECT 37.265 7.8 37.435 7.97 ;
      RECT 36.915 0.1 37.085 0.27 ;
      RECT 36.915 8.61 37.085 8.78 ;
      RECT 36.895 2.76 37.065 2.93 ;
      RECT 36.895 5.95 37.065 6.12 ;
      RECT 36.215 0.105 36.385 0.275 ;
      RECT 36.215 8.605 36.385 8.775 ;
      RECT 35.905 2.025 36.075 2.195 ;
      RECT 35.905 6.685 36.075 6.855 ;
      RECT 35.535 0.105 35.705 0.275 ;
      RECT 35.535 8.605 35.705 8.775 ;
      RECT 35.475 0.915 35.645 1.085 ;
      RECT 35.475 1.655 35.645 1.825 ;
      RECT 35.475 7.055 35.645 7.225 ;
      RECT 35.475 7.795 35.645 7.965 ;
      RECT 35.1 2.395 35.27 2.565 ;
      RECT 35.1 6.315 35.27 6.485 ;
      RECT 34.855 0.105 35.025 0.275 ;
      RECT 34.855 8.605 35.025 8.775 ;
      RECT 34.175 0.105 34.345 0.275 ;
      RECT 34.175 8.605 34.345 8.775 ;
      RECT 32.895 1.565 33.065 1.735 ;
      RECT 32.435 1.565 32.605 1.735 ;
      RECT 32.04 2.905 32.21 3.075 ;
      RECT 31.975 1.565 32.145 1.735 ;
      RECT 31.83 2.245 32 2.415 ;
      RECT 31.515 1.565 31.685 1.735 ;
      RECT 31.515 3.155 31.685 3.325 ;
      RECT 31.455 8.605 31.625 8.775 ;
      RECT 31.145 6.685 31.315 6.855 ;
      RECT 31.13 2.75 31.3 2.92 ;
      RECT 31.055 1.565 31.225 1.735 ;
      RECT 30.915 3.315 31.085 3.485 ;
      RECT 30.895 3.715 31.065 3.885 ;
      RECT 30.775 8.605 30.945 8.775 ;
      RECT 30.72 2.27 30.89 2.44 ;
      RECT 30.715 7.055 30.885 7.225 ;
      RECT 30.715 7.795 30.885 7.965 ;
      RECT 30.595 1.565 30.765 1.735 ;
      RECT 30.34 6.315 30.51 6.485 ;
      RECT 30.225 3.25 30.395 3.42 ;
      RECT 30.135 1.565 30.305 1.735 ;
      RECT 30.095 8.605 30.265 8.775 ;
      RECT 29.9 2.935 30.07 3.105 ;
      RECT 29.835 3.715 30.005 3.885 ;
      RECT 29.675 1.565 29.845 1.735 ;
      RECT 29.435 3.7 29.605 3.87 ;
      RECT 29.415 8.605 29.585 8.775 ;
      RECT 29.395 2.185 29.565 2.355 ;
      RECT 29.215 1.565 29.385 1.735 ;
      RECT 28.755 1.565 28.925 1.735 ;
      RECT 28.495 2.685 28.665 2.855 ;
      RECT 28.495 3.145 28.665 3.315 ;
      RECT 28.495 3.66 28.665 3.83 ;
      RECT 28.38 2.22 28.55 2.39 ;
      RECT 28.295 1.565 28.465 1.735 ;
      RECT 27.915 3.73 28.085 3.9 ;
      RECT 27.835 1.565 28.005 1.735 ;
      RECT 27.435 2.26 27.605 2.43 ;
      RECT 27.375 1.565 27.545 1.735 ;
      RECT 27.22 2.635 27.39 2.805 ;
      RECT 26.915 1.565 27.085 1.735 ;
      RECT 26.72 3.235 26.89 3.405 ;
      RECT 26.605 2.685 26.775 2.855 ;
      RECT 26.455 1.565 26.625 1.735 ;
      RECT 26.435 2.135 26.605 2.305 ;
      RECT 26.06 3.165 26.23 3.335 ;
      RECT 25.995 1.565 26.165 1.735 ;
      RECT 25.575 2.765 25.745 2.935 ;
      RECT 25.535 1.565 25.705 1.735 ;
      RECT 25.525 3.54 25.695 3.71 ;
      RECT 25.075 1.565 25.245 1.735 ;
      RECT 25.035 3.165 25.205 3.335 ;
      RECT 25 2.27 25.17 2.44 ;
      RECT 24.64 2.67 24.81 2.84 ;
      RECT 24.615 1.565 24.785 1.735 ;
      RECT 24.435 3.48 24.605 3.65 ;
      RECT 24.155 1.565 24.325 1.735 ;
      RECT 24.13 2.91 24.3 3.08 ;
      RECT 23.695 1.565 23.865 1.735 ;
      RECT 23.43 2.7 23.6 2.87 ;
      RECT 23.235 1.565 23.405 1.735 ;
      RECT 23.11 3.145 23.28 3.315 ;
      RECT 22.775 1.565 22.945 1.735 ;
      RECT 22.695 3.18 22.865 3.35 ;
      RECT 22.525 2.165 22.695 2.335 ;
      RECT 22.35 2.62 22.52 2.79 ;
      RECT 22.315 1.565 22.485 1.735 ;
      RECT 21.855 1.565 22.025 1.735 ;
      RECT 21.43 2.27 21.6 2.44 ;
      RECT 21.425 3.585 21.595 3.755 ;
      RECT 21.395 1.565 21.565 1.735 ;
      RECT 20.33 7.8 20.5 7.97 ;
      RECT 19.98 0.1 20.15 0.27 ;
      RECT 19.98 8.61 20.15 8.78 ;
      RECT 19.96 2.76 20.13 2.93 ;
      RECT 19.96 5.95 20.13 6.12 ;
      RECT 19.34 0.91 19.51 1.08 ;
      RECT 19.34 2.39 19.51 2.56 ;
      RECT 19.34 6.32 19.51 6.49 ;
      RECT 19.34 7.8 19.51 7.97 ;
      RECT 18.99 0.1 19.16 0.27 ;
      RECT 18.99 8.61 19.16 8.78 ;
      RECT 18.97 2.76 19.14 2.93 ;
      RECT 18.97 5.95 19.14 6.12 ;
      RECT 18.29 0.105 18.46 0.275 ;
      RECT 18.29 8.605 18.46 8.775 ;
      RECT 17.98 2.025 18.15 2.195 ;
      RECT 17.98 6.685 18.15 6.855 ;
      RECT 17.61 0.105 17.78 0.275 ;
      RECT 17.61 8.605 17.78 8.775 ;
      RECT 17.55 0.915 17.72 1.085 ;
      RECT 17.55 1.655 17.72 1.825 ;
      RECT 17.55 7.055 17.72 7.225 ;
      RECT 17.55 7.795 17.72 7.965 ;
      RECT 17.175 2.395 17.345 2.565 ;
      RECT 17.175 6.315 17.345 6.485 ;
      RECT 16.93 0.105 17.1 0.275 ;
      RECT 16.93 8.605 17.1 8.775 ;
      RECT 16.25 0.105 16.42 0.275 ;
      RECT 16.25 8.605 16.42 8.775 ;
      RECT 14.97 1.565 15.14 1.735 ;
      RECT 14.51 1.565 14.68 1.735 ;
      RECT 14.115 2.905 14.285 3.075 ;
      RECT 14.05 1.565 14.22 1.735 ;
      RECT 13.905 2.245 14.075 2.415 ;
      RECT 13.59 1.565 13.76 1.735 ;
      RECT 13.59 3.155 13.76 3.325 ;
      RECT 13.53 8.605 13.7 8.775 ;
      RECT 13.22 6.685 13.39 6.855 ;
      RECT 13.205 2.75 13.375 2.92 ;
      RECT 13.13 1.565 13.3 1.735 ;
      RECT 12.99 3.315 13.16 3.485 ;
      RECT 12.97 3.715 13.14 3.885 ;
      RECT 12.85 8.605 13.02 8.775 ;
      RECT 12.795 2.27 12.965 2.44 ;
      RECT 12.79 7.055 12.96 7.225 ;
      RECT 12.79 7.795 12.96 7.965 ;
      RECT 12.67 1.565 12.84 1.735 ;
      RECT 12.415 6.315 12.585 6.485 ;
      RECT 12.3 3.25 12.47 3.42 ;
      RECT 12.21 1.565 12.38 1.735 ;
      RECT 12.17 8.605 12.34 8.775 ;
      RECT 11.975 2.935 12.145 3.105 ;
      RECT 11.91 3.715 12.08 3.885 ;
      RECT 11.75 1.565 11.92 1.735 ;
      RECT 11.51 3.7 11.68 3.87 ;
      RECT 11.49 8.605 11.66 8.775 ;
      RECT 11.47 2.185 11.64 2.355 ;
      RECT 11.29 1.565 11.46 1.735 ;
      RECT 10.83 1.565 11 1.735 ;
      RECT 10.57 2.685 10.74 2.855 ;
      RECT 10.57 3.145 10.74 3.315 ;
      RECT 10.57 3.66 10.74 3.83 ;
      RECT 10.455 2.22 10.625 2.39 ;
      RECT 10.37 1.565 10.54 1.735 ;
      RECT 9.99 3.73 10.16 3.9 ;
      RECT 9.91 1.565 10.08 1.735 ;
      RECT 9.51 2.26 9.68 2.43 ;
      RECT 9.45 1.565 9.62 1.735 ;
      RECT 9.295 2.635 9.465 2.805 ;
      RECT 8.99 1.565 9.16 1.735 ;
      RECT 8.795 3.235 8.965 3.405 ;
      RECT 8.68 2.685 8.85 2.855 ;
      RECT 8.53 1.565 8.7 1.735 ;
      RECT 8.51 2.135 8.68 2.305 ;
      RECT 8.135 3.165 8.305 3.335 ;
      RECT 8.07 1.565 8.24 1.735 ;
      RECT 7.65 2.765 7.82 2.935 ;
      RECT 7.61 1.565 7.78 1.735 ;
      RECT 7.6 3.54 7.77 3.71 ;
      RECT 7.15 1.565 7.32 1.735 ;
      RECT 7.11 3.165 7.28 3.335 ;
      RECT 7.075 2.27 7.245 2.44 ;
      RECT 6.715 2.67 6.885 2.84 ;
      RECT 6.69 1.565 6.86 1.735 ;
      RECT 6.51 3.48 6.68 3.65 ;
      RECT 6.23 1.565 6.4 1.735 ;
      RECT 6.205 2.91 6.375 3.08 ;
      RECT 5.77 1.565 5.94 1.735 ;
      RECT 5.505 2.7 5.675 2.87 ;
      RECT 5.31 1.565 5.48 1.735 ;
      RECT 5.185 3.145 5.355 3.315 ;
      RECT 4.85 1.565 5.02 1.735 ;
      RECT 4.77 3.18 4.94 3.35 ;
      RECT 4.6 2.165 4.77 2.335 ;
      RECT 4.425 2.62 4.595 2.79 ;
      RECT 4.39 1.565 4.56 1.735 ;
      RECT 3.93 1.565 4.1 1.735 ;
      RECT 3.505 2.27 3.675 2.44 ;
      RECT 3.5 3.585 3.67 3.755 ;
      RECT 3.47 1.565 3.64 1.735 ;
      RECT 2.5 8.605 2.67 8.775 ;
      RECT 1.82 8.605 1.99 8.775 ;
      RECT 1.76 7.055 1.93 7.225 ;
      RECT 1.76 7.795 1.93 7.965 ;
      RECT 1.385 6.315 1.555 6.485 ;
      RECT 1.14 8.605 1.31 8.775 ;
      RECT 0.46 8.605 0.63 8.775 ;
    LAYER li1 ;
      RECT 86.075 0 86.245 2.235 ;
      RECT 85.115 0 85.285 2.235 ;
      RECT 84.155 0 84.325 2.235 ;
      RECT 83.635 0 83.805 2.235 ;
      RECT 82.675 0 82.845 2.235 ;
      RECT 81.675 0 81.845 2.235 ;
      RECT 80.715 0 80.885 2.235 ;
      RECT 79.235 0 79.405 2.235 ;
      RECT 77.315 0 77.485 2.235 ;
      RECT 75.835 0 76.005 2.235 ;
      RECT 68.15 0 68.32 2.235 ;
      RECT 67.19 0 67.36 2.235 ;
      RECT 66.23 0 66.4 2.235 ;
      RECT 65.71 0 65.88 2.235 ;
      RECT 64.75 0 64.92 2.235 ;
      RECT 63.75 0 63.92 2.235 ;
      RECT 62.79 0 62.96 2.235 ;
      RECT 61.31 0 61.48 2.235 ;
      RECT 59.39 0 59.56 2.235 ;
      RECT 57.91 0 58.08 2.235 ;
      RECT 50.225 0 50.395 2.235 ;
      RECT 49.265 0 49.435 2.235 ;
      RECT 48.305 0 48.475 2.235 ;
      RECT 47.785 0 47.955 2.235 ;
      RECT 46.825 0 46.995 2.235 ;
      RECT 45.825 0 45.995 2.235 ;
      RECT 44.865 0 45.035 2.235 ;
      RECT 43.385 0 43.555 2.235 ;
      RECT 41.465 0 41.635 2.235 ;
      RECT 39.985 0 40.155 2.235 ;
      RECT 32.3 0 32.47 2.235 ;
      RECT 31.34 0 31.51 2.235 ;
      RECT 30.38 0 30.55 2.235 ;
      RECT 29.86 0 30.03 2.235 ;
      RECT 28.9 0 29.07 2.235 ;
      RECT 27.9 0 28.07 2.235 ;
      RECT 26.94 0 27.11 2.235 ;
      RECT 25.46 0 25.63 2.235 ;
      RECT 23.54 0 23.71 2.235 ;
      RECT 22.06 0 22.23 2.235 ;
      RECT 14.375 0 14.545 2.235 ;
      RECT 13.415 0 13.585 2.235 ;
      RECT 12.455 0 12.625 2.235 ;
      RECT 11.935 0 12.105 2.235 ;
      RECT 10.975 0 11.145 2.235 ;
      RECT 9.975 0 10.145 2.235 ;
      RECT 9.015 0 9.185 2.235 ;
      RECT 7.535 0 7.705 2.235 ;
      RECT 5.615 0 5.785 2.235 ;
      RECT 4.135 0 4.305 2.235 ;
      RECT 75.025 0 86.985 1.735 ;
      RECT 57.1 0 69.06 1.735 ;
      RECT 39.175 0 51.135 1.735 ;
      RECT 21.25 0 33.21 1.735 ;
      RECT 3.325 0 15.285 1.735 ;
      RECT 75.02 0 86.985 1.68 ;
      RECT 57.095 0 69.06 1.68 ;
      RECT 39.17 0 51.135 1.68 ;
      RECT 21.245 0 33.21 1.68 ;
      RECT 3.32 0 15.285 1.68 ;
      RECT 87.87 0 88.04 0.935 ;
      RECT 69.945 0 70.115 0.935 ;
      RECT 52.02 0 52.19 0.935 ;
      RECT 34.095 0 34.265 0.935 ;
      RECT 16.17 0 16.34 0.935 ;
      RECT 91.6 0 91.77 0.93 ;
      RECT 90.61 0 90.78 0.93 ;
      RECT 73.675 0 73.845 0.93 ;
      RECT 72.685 0 72.855 0.93 ;
      RECT 55.75 0 55.92 0.93 ;
      RECT 54.76 0 54.93 0.93 ;
      RECT 37.825 0 37.995 0.93 ;
      RECT 36.835 0 37.005 0.93 ;
      RECT 19.9 0 20.07 0.93 ;
      RECT 18.91 0 19.08 0.93 ;
      RECT 92.395 0 92.575 0.305 ;
      RECT 74.47 0 90.445 0.305 ;
      RECT 56.545 0 72.52 0.305 ;
      RECT 38.62 0 54.595 0.305 ;
      RECT 20.695 0 36.67 0.305 ;
      RECT 0 0 18.745 0.305 ;
      RECT 0 0 92.575 0.3 ;
      RECT 0 8.58 92.575 8.88 ;
      RECT 92.395 8.575 92.575 8.88 ;
      RECT 91.6 7.95 91.77 8.88 ;
      RECT 90.61 7.95 90.78 8.88 ;
      RECT 74.47 8.575 90.445 8.88 ;
      RECT 73.675 7.95 73.845 8.88 ;
      RECT 72.685 7.95 72.855 8.88 ;
      RECT 56.545 8.575 72.52 8.88 ;
      RECT 55.75 7.95 55.92 8.88 ;
      RECT 54.76 7.95 54.93 8.88 ;
      RECT 38.62 8.575 54.595 8.88 ;
      RECT 37.825 7.95 37.995 8.88 ;
      RECT 36.835 7.95 37.005 8.88 ;
      RECT 20.695 8.575 36.67 8.88 ;
      RECT 19.9 7.95 20.07 8.88 ;
      RECT 18.91 7.95 19.08 8.88 ;
      RECT 0 8.575 18.745 8.88 ;
      RECT 87.87 7.945 88.04 8.88 ;
      RECT 83.11 7.945 83.28 8.88 ;
      RECT 69.945 7.945 70.115 8.88 ;
      RECT 65.185 7.945 65.355 8.88 ;
      RECT 52.02 7.945 52.19 8.88 ;
      RECT 47.26 7.945 47.43 8.88 ;
      RECT 34.095 7.945 34.265 8.88 ;
      RECT 29.335 7.945 29.505 8.88 ;
      RECT 16.17 7.945 16.34 8.88 ;
      RECT 11.41 7.945 11.58 8.88 ;
      RECT 0.38 7.945 0.55 8.88 ;
      RECT 92.03 5.02 92.2 6.49 ;
      RECT 92.03 6.315 92.205 6.485 ;
      RECT 91.66 1.74 91.83 2.93 ;
      RECT 91.66 1.74 92.13 1.91 ;
      RECT 91.66 6.97 92.13 7.14 ;
      RECT 91.66 5.95 91.83 7.14 ;
      RECT 90.67 1.74 90.84 2.93 ;
      RECT 90.67 1.74 91.14 1.91 ;
      RECT 90.67 6.97 91.14 7.14 ;
      RECT 90.67 5.95 90.84 7.14 ;
      RECT 88.82 2.635 88.99 3.865 ;
      RECT 88.875 0.855 89.045 2.805 ;
      RECT 88.82 0.575 88.99 1.025 ;
      RECT 88.82 7.855 88.99 8.305 ;
      RECT 88.875 6.075 89.045 8.025 ;
      RECT 88.82 5.015 88.99 6.245 ;
      RECT 88.3 0.575 88.47 3.865 ;
      RECT 88.3 2.075 88.705 2.405 ;
      RECT 88.3 1.235 88.705 1.565 ;
      RECT 88.3 5.015 88.47 8.305 ;
      RECT 88.3 7.315 88.705 7.645 ;
      RECT 88.3 6.475 88.705 6.805 ;
      RECT 86.4 3.392 86.415 3.443 ;
      RECT 86.395 3.372 86.4 3.49 ;
      RECT 86.38 3.362 86.395 3.558 ;
      RECT 86.355 3.342 86.38 3.613 ;
      RECT 86.315 3.327 86.355 3.633 ;
      RECT 86.27 3.321 86.315 3.661 ;
      RECT 86.2 3.311 86.27 3.678 ;
      RECT 86.18 3.303 86.2 3.678 ;
      RECT 86.12 3.297 86.18 3.67 ;
      RECT 86.061 3.288 86.12 3.658 ;
      RECT 85.975 3.277 86.061 3.641 ;
      RECT 85.953 3.268 85.975 3.629 ;
      RECT 85.867 3.261 85.953 3.616 ;
      RECT 85.781 3.248 85.867 3.597 ;
      RECT 85.695 3.236 85.781 3.577 ;
      RECT 85.665 3.225 85.695 3.564 ;
      RECT 85.615 3.211 85.665 3.556 ;
      RECT 85.595 3.2 85.615 3.548 ;
      RECT 85.546 3.189 85.595 3.54 ;
      RECT 85.46 3.168 85.546 3.525 ;
      RECT 85.415 3.155 85.46 3.51 ;
      RECT 85.37 3.155 85.415 3.49 ;
      RECT 85.315 3.155 85.37 3.425 ;
      RECT 85.29 3.155 85.315 3.348 ;
      RECT 85.815 2.892 85.985 3.075 ;
      RECT 85.815 2.892 86 3.033 ;
      RECT 85.815 2.892 86.005 2.975 ;
      RECT 85.875 2.66 86.01 2.951 ;
      RECT 85.875 2.664 86.015 2.934 ;
      RECT 85.82 2.827 86.015 2.934 ;
      RECT 85.845 2.672 85.985 3.075 ;
      RECT 85.845 2.676 86.025 2.875 ;
      RECT 85.83 2.762 86.025 2.875 ;
      RECT 85.84 2.692 85.985 3.075 ;
      RECT 85.84 2.695 86.035 2.788 ;
      RECT 85.835 2.712 86.035 2.788 ;
      RECT 85.605 1.932 85.775 2.415 ;
      RECT 85.6 1.927 85.75 2.405 ;
      RECT 85.6 1.934 85.78 2.399 ;
      RECT 85.59 1.928 85.75 2.378 ;
      RECT 85.59 1.944 85.795 2.337 ;
      RECT 85.56 1.929 85.75 2.3 ;
      RECT 85.56 1.959 85.805 2.24 ;
      RECT 85.555 1.931 85.75 2.238 ;
      RECT 85.535 1.94 85.78 2.195 ;
      RECT 85.51 1.956 85.795 2.107 ;
      RECT 85.51 1.975 85.82 2.098 ;
      RECT 85.505 2.012 85.82 2.05 ;
      RECT 85.51 1.992 85.825 2.018 ;
      RECT 85.605 1.926 85.715 2.415 ;
      RECT 85.691 1.925 85.715 2.415 ;
      RECT 84.925 2.71 84.93 2.921 ;
      RECT 85.525 2.71 85.53 2.895 ;
      RECT 85.59 2.75 85.595 2.863 ;
      RECT 85.585 2.742 85.59 2.869 ;
      RECT 85.58 2.732 85.585 2.877 ;
      RECT 85.575 2.722 85.58 2.886 ;
      RECT 85.57 2.712 85.575 2.89 ;
      RECT 85.53 2.71 85.57 2.893 ;
      RECT 85.502 2.709 85.525 2.897 ;
      RECT 85.416 2.706 85.502 2.904 ;
      RECT 85.33 2.702 85.416 2.915 ;
      RECT 85.31 2.7 85.33 2.921 ;
      RECT 85.292 2.699 85.31 2.924 ;
      RECT 85.206 2.697 85.292 2.931 ;
      RECT 85.12 2.692 85.206 2.944 ;
      RECT 85.101 2.689 85.12 2.949 ;
      RECT 85.015 2.687 85.101 2.94 ;
      RECT 85.005 2.687 85.015 2.933 ;
      RECT 84.93 2.7 85.005 2.927 ;
      RECT 84.915 2.711 84.925 2.921 ;
      RECT 84.905 2.713 84.915 2.92 ;
      RECT 84.895 2.717 84.905 2.916 ;
      RECT 84.89 2.72 84.895 2.91 ;
      RECT 84.88 2.722 84.89 2.904 ;
      RECT 84.875 2.725 84.88 2.898 ;
      RECT 84.855 3.311 84.86 3.515 ;
      RECT 84.84 3.298 84.855 3.608 ;
      RECT 84.825 3.279 84.84 3.885 ;
      RECT 84.79 3.245 84.825 3.885 ;
      RECT 84.786 3.215 84.79 3.885 ;
      RECT 84.7 3.097 84.786 3.885 ;
      RECT 84.69 2.972 84.7 3.885 ;
      RECT 84.675 2.94 84.69 3.885 ;
      RECT 84.67 2.915 84.675 3.885 ;
      RECT 84.665 2.905 84.67 3.841 ;
      RECT 84.65 2.877 84.665 3.746 ;
      RECT 84.635 2.843 84.65 3.645 ;
      RECT 84.63 2.821 84.635 3.598 ;
      RECT 84.625 2.81 84.63 3.568 ;
      RECT 84.62 2.8 84.625 3.534 ;
      RECT 84.61 2.787 84.62 3.502 ;
      RECT 84.585 2.763 84.61 3.428 ;
      RECT 84.58 2.743 84.585 3.353 ;
      RECT 84.575 2.737 84.58 3.328 ;
      RECT 84.57 2.732 84.575 3.293 ;
      RECT 84.565 2.727 84.57 3.268 ;
      RECT 84.56 2.725 84.565 3.248 ;
      RECT 84.555 2.725 84.56 3.233 ;
      RECT 84.55 2.725 84.555 3.193 ;
      RECT 84.54 2.725 84.55 3.165 ;
      RECT 84.53 2.725 84.54 3.11 ;
      RECT 84.515 2.725 84.53 3.048 ;
      RECT 84.51 2.724 84.515 2.993 ;
      RECT 84.495 2.723 84.51 2.973 ;
      RECT 84.435 2.721 84.495 2.947 ;
      RECT 84.4 2.722 84.435 2.927 ;
      RECT 84.395 2.724 84.4 2.917 ;
      RECT 84.385 2.743 84.395 2.907 ;
      RECT 84.38 2.77 84.385 2.838 ;
      RECT 84.495 2.195 84.665 2.44 ;
      RECT 84.53 1.966 84.665 2.44 ;
      RECT 84.53 1.968 84.675 2.435 ;
      RECT 84.53 1.97 84.7 2.423 ;
      RECT 84.53 1.973 84.725 2.405 ;
      RECT 84.53 1.978 84.775 2.378 ;
      RECT 84.53 1.983 84.795 2.343 ;
      RECT 84.51 1.985 84.805 2.318 ;
      RECT 84.5 2.08 84.805 2.318 ;
      RECT 84.53 1.965 84.64 2.44 ;
      RECT 84.54 1.962 84.635 2.44 ;
      RECT 84.06 3.227 84.25 3.585 ;
      RECT 84.06 3.239 84.285 3.584 ;
      RECT 84.06 3.267 84.305 3.582 ;
      RECT 84.06 3.292 84.31 3.581 ;
      RECT 84.06 3.35 84.325 3.58 ;
      RECT 84.045 3.223 84.205 3.565 ;
      RECT 84.025 3.232 84.25 3.518 ;
      RECT 84 3.243 84.285 3.455 ;
      RECT 84 3.327 84.32 3.455 ;
      RECT 84 3.302 84.315 3.455 ;
      RECT 84.06 3.218 84.205 3.585 ;
      RECT 84.146 3.217 84.205 3.585 ;
      RECT 84.146 3.216 84.19 3.585 ;
      RECT 84.06 7.855 84.23 8.305 ;
      RECT 84.115 6.075 84.285 8.025 ;
      RECT 84.06 5.015 84.23 6.245 ;
      RECT 83.54 5.015 83.71 8.305 ;
      RECT 83.54 7.315 83.945 7.645 ;
      RECT 83.54 6.475 83.945 6.805 ;
      RECT 83.845 2.732 83.85 3.11 ;
      RECT 83.84 2.7 83.845 3.11 ;
      RECT 83.835 2.672 83.84 3.11 ;
      RECT 83.83 2.652 83.835 3.11 ;
      RECT 83.775 2.635 83.83 3.11 ;
      RECT 83.735 2.62 83.775 3.11 ;
      RECT 83.68 2.607 83.735 3.11 ;
      RECT 83.645 2.598 83.68 3.11 ;
      RECT 83.641 2.596 83.645 3.109 ;
      RECT 83.555 2.592 83.641 3.092 ;
      RECT 83.47 2.584 83.555 3.055 ;
      RECT 83.46 2.58 83.47 3.028 ;
      RECT 83.45 2.58 83.46 3.01 ;
      RECT 83.44 2.582 83.45 2.993 ;
      RECT 83.435 2.587 83.44 2.979 ;
      RECT 83.43 2.591 83.435 2.966 ;
      RECT 83.42 2.596 83.43 2.95 ;
      RECT 83.405 2.61 83.42 2.925 ;
      RECT 83.4 2.616 83.405 2.905 ;
      RECT 83.395 2.618 83.4 2.898 ;
      RECT 83.39 2.622 83.395 2.773 ;
      RECT 83.57 3.422 83.815 3.885 ;
      RECT 83.49 3.395 83.81 3.881 ;
      RECT 83.42 3.43 83.815 3.874 ;
      RECT 83.21 3.685 83.815 3.87 ;
      RECT 83.39 3.453 83.815 3.87 ;
      RECT 83.23 3.645 83.815 3.87 ;
      RECT 83.38 3.465 83.815 3.87 ;
      RECT 83.265 3.582 83.815 3.87 ;
      RECT 83.32 3.507 83.815 3.87 ;
      RECT 83.57 3.372 83.81 3.885 ;
      RECT 83.6 3.365 83.81 3.885 ;
      RECT 83.59 3.367 83.81 3.885 ;
      RECT 83.6 3.362 83.73 3.885 ;
      RECT 83.155 1.925 83.241 2.364 ;
      RECT 83.15 1.925 83.241 2.362 ;
      RECT 83.15 1.925 83.31 2.361 ;
      RECT 83.15 1.925 83.34 2.358 ;
      RECT 83.135 1.932 83.34 2.349 ;
      RECT 83.135 1.932 83.345 2.345 ;
      RECT 83.13 1.942 83.345 2.338 ;
      RECT 83.125 1.947 83.345 2.313 ;
      RECT 83.125 1.947 83.36 2.295 ;
      RECT 83.15 1.925 83.38 2.21 ;
      RECT 83.12 1.952 83.38 2.208 ;
      RECT 83.13 1.945 83.385 2.146 ;
      RECT 83.12 2.067 83.39 2.129 ;
      RECT 83.105 1.962 83.385 2.08 ;
      RECT 83.1 1.972 83.385 1.98 ;
      RECT 83.18 2.743 83.185 2.82 ;
      RECT 83.17 2.737 83.18 3.01 ;
      RECT 83.16 2.729 83.17 3.031 ;
      RECT 83.15 2.72 83.16 3.053 ;
      RECT 83.145 2.715 83.15 3.07 ;
      RECT 83.105 2.715 83.145 3.11 ;
      RECT 83.085 2.715 83.105 3.165 ;
      RECT 83.08 2.715 83.085 3.193 ;
      RECT 83.07 2.715 83.08 3.208 ;
      RECT 83.035 2.715 83.07 3.25 ;
      RECT 83.03 2.715 83.035 3.293 ;
      RECT 83.02 2.715 83.03 3.308 ;
      RECT 83.005 2.715 83.02 3.328 ;
      RECT 82.99 2.715 83.005 3.355 ;
      RECT 82.985 2.716 82.99 3.373 ;
      RECT 82.965 2.717 82.985 3.38 ;
      RECT 82.91 2.718 82.965 3.4 ;
      RECT 82.9 2.719 82.91 3.414 ;
      RECT 82.895 2.722 82.9 3.413 ;
      RECT 82.855 2.795 82.895 3.411 ;
      RECT 82.84 2.875 82.855 3.409 ;
      RECT 82.815 2.93 82.84 3.407 ;
      RECT 82.8 2.995 82.815 3.406 ;
      RECT 82.755 3.027 82.8 3.403 ;
      RECT 82.67 3.05 82.755 3.398 ;
      RECT 82.645 3.07 82.67 3.393 ;
      RECT 82.575 3.075 82.645 3.389 ;
      RECT 82.555 3.077 82.575 3.386 ;
      RECT 82.47 3.088 82.555 3.38 ;
      RECT 82.465 3.099 82.47 3.375 ;
      RECT 82.455 3.101 82.465 3.375 ;
      RECT 82.42 3.105 82.455 3.373 ;
      RECT 82.37 3.115 82.42 3.36 ;
      RECT 82.35 3.123 82.37 3.345 ;
      RECT 82.27 3.135 82.35 3.328 ;
      RECT 82.435 2.685 82.605 2.895 ;
      RECT 82.551 2.681 82.605 2.895 ;
      RECT 82.356 2.685 82.605 2.886 ;
      RECT 82.356 2.685 82.61 2.875 ;
      RECT 82.27 2.685 82.61 2.866 ;
      RECT 82.27 2.693 82.62 2.81 ;
      RECT 82.27 2.705 82.625 2.723 ;
      RECT 82.27 2.712 82.63 2.715 ;
      RECT 82.465 2.683 82.605 2.895 ;
      RECT 82.22 3.628 82.465 3.96 ;
      RECT 82.215 3.62 82.22 3.957 ;
      RECT 82.185 3.64 82.465 3.938 ;
      RECT 82.165 3.672 82.465 3.911 ;
      RECT 82.215 3.625 82.392 3.957 ;
      RECT 82.215 3.622 82.306 3.957 ;
      RECT 82.155 1.97 82.325 2.39 ;
      RECT 82.15 1.97 82.325 2.388 ;
      RECT 82.15 1.97 82.35 2.378 ;
      RECT 82.15 1.97 82.37 2.353 ;
      RECT 82.145 1.97 82.37 2.348 ;
      RECT 82.145 1.97 82.38 2.338 ;
      RECT 82.145 1.97 82.385 2.333 ;
      RECT 82.145 1.975 82.39 2.328 ;
      RECT 82.145 2.007 82.405 2.318 ;
      RECT 82.145 2.077 82.43 2.301 ;
      RECT 82.125 2.077 82.43 2.293 ;
      RECT 82.125 2.137 82.44 2.27 ;
      RECT 82.125 2.177 82.45 2.215 ;
      RECT 82.11 1.97 82.385 2.195 ;
      RECT 82.1 1.985 82.39 2.093 ;
      RECT 81.69 3.375 81.86 3.9 ;
      RECT 81.685 3.375 81.86 3.893 ;
      RECT 81.675 3.375 81.865 3.858 ;
      RECT 81.67 3.385 81.865 3.83 ;
      RECT 81.665 3.405 81.865 3.813 ;
      RECT 81.675 3.38 81.87 3.803 ;
      RECT 81.66 3.425 81.87 3.795 ;
      RECT 81.655 3.445 81.87 3.78 ;
      RECT 81.65 3.475 81.87 3.77 ;
      RECT 81.64 3.52 81.87 3.745 ;
      RECT 81.67 3.39 81.875 3.728 ;
      RECT 81.635 3.572 81.875 3.723 ;
      RECT 81.67 3.4 81.88 3.693 ;
      RECT 81.63 3.605 81.88 3.69 ;
      RECT 81.625 3.63 81.88 3.67 ;
      RECT 81.665 3.417 81.89 3.61 ;
      RECT 81.66 3.439 81.9 3.503 ;
      RECT 81.61 2.686 81.625 2.955 ;
      RECT 81.565 2.67 81.61 3 ;
      RECT 81.56 2.658 81.565 3.05 ;
      RECT 81.55 2.654 81.56 3.083 ;
      RECT 81.545 2.651 81.55 3.111 ;
      RECT 81.53 2.653 81.545 3.153 ;
      RECT 81.525 2.657 81.53 3.193 ;
      RECT 81.505 2.662 81.525 3.245 ;
      RECT 81.501 2.667 81.505 3.302 ;
      RECT 81.415 2.686 81.501 3.339 ;
      RECT 81.405 2.707 81.415 3.375 ;
      RECT 81.4 2.715 81.405 3.376 ;
      RECT 81.395 2.757 81.4 3.377 ;
      RECT 81.38 2.845 81.395 3.378 ;
      RECT 81.37 2.995 81.38 3.38 ;
      RECT 81.365 3.04 81.37 3.382 ;
      RECT 81.33 3.082 81.365 3.385 ;
      RECT 81.325 3.1 81.33 3.388 ;
      RECT 81.248 3.106 81.325 3.394 ;
      RECT 81.162 3.12 81.248 3.407 ;
      RECT 81.076 3.134 81.162 3.421 ;
      RECT 80.99 3.148 81.076 3.434 ;
      RECT 80.93 3.16 80.99 3.446 ;
      RECT 80.905 3.167 80.93 3.453 ;
      RECT 80.891 3.17 80.905 3.458 ;
      RECT 80.805 3.178 80.891 3.474 ;
      RECT 80.8 3.185 80.805 3.489 ;
      RECT 80.776 3.185 80.8 3.496 ;
      RECT 80.69 3.188 80.776 3.524 ;
      RECT 80.605 3.192 80.69 3.568 ;
      RECT 80.54 3.196 80.605 3.605 ;
      RECT 80.515 3.199 80.54 3.621 ;
      RECT 80.44 3.212 80.515 3.625 ;
      RECT 80.415 3.23 80.44 3.629 ;
      RECT 80.405 3.237 80.415 3.631 ;
      RECT 80.39 3.24 80.405 3.632 ;
      RECT 80.33 3.252 80.39 3.636 ;
      RECT 80.32 3.266 80.33 3.64 ;
      RECT 80.265 3.276 80.32 3.628 ;
      RECT 80.24 3.297 80.265 3.611 ;
      RECT 80.22 3.317 80.24 3.602 ;
      RECT 80.215 3.33 80.22 3.597 ;
      RECT 80.2 3.342 80.215 3.593 ;
      RECT 81.435 1.997 81.44 2.02 ;
      RECT 81.43 1.988 81.435 2.06 ;
      RECT 81.425 1.986 81.43 2.103 ;
      RECT 81.42 1.977 81.425 2.138 ;
      RECT 81.415 1.967 81.42 2.21 ;
      RECT 81.41 1.957 81.415 2.275 ;
      RECT 81.405 1.954 81.41 2.315 ;
      RECT 81.38 1.948 81.405 2.405 ;
      RECT 81.345 1.936 81.38 2.43 ;
      RECT 81.335 1.927 81.345 2.43 ;
      RECT 81.2 1.925 81.21 2.413 ;
      RECT 81.19 1.925 81.2 2.38 ;
      RECT 81.185 1.925 81.19 2.355 ;
      RECT 81.18 1.925 81.185 2.343 ;
      RECT 81.175 1.925 81.18 2.325 ;
      RECT 81.165 1.925 81.175 2.29 ;
      RECT 81.16 1.927 81.165 2.268 ;
      RECT 81.155 1.933 81.16 2.253 ;
      RECT 81.15 1.939 81.155 2.238 ;
      RECT 81.135 1.951 81.15 2.211 ;
      RECT 81.13 1.962 81.135 2.179 ;
      RECT 81.125 1.972 81.13 2.163 ;
      RECT 81.115 1.98 81.125 2.132 ;
      RECT 81.11 1.99 81.115 2.106 ;
      RECT 81.105 2.047 81.11 2.089 ;
      RECT 81.21 1.925 81.335 2.43 ;
      RECT 80.925 2.612 81.185 2.91 ;
      RECT 80.92 2.619 81.185 2.908 ;
      RECT 80.925 2.614 81.2 2.903 ;
      RECT 80.915 2.627 81.2 2.9 ;
      RECT 80.915 2.632 81.205 2.893 ;
      RECT 80.91 2.64 81.205 2.89 ;
      RECT 80.91 2.657 81.21 2.688 ;
      RECT 80.925 2.609 81.156 2.91 ;
      RECT 80.98 2.608 81.156 2.91 ;
      RECT 80.98 2.605 81.07 2.91 ;
      RECT 80.98 2.602 81.066 2.91 ;
      RECT 80.67 2.875 80.675 2.888 ;
      RECT 80.665 2.842 80.67 2.893 ;
      RECT 80.66 2.797 80.665 2.9 ;
      RECT 80.655 2.752 80.66 2.908 ;
      RECT 80.65 2.72 80.655 2.916 ;
      RECT 80.645 2.68 80.65 2.917 ;
      RECT 80.63 2.66 80.645 2.919 ;
      RECT 80.555 2.642 80.63 2.931 ;
      RECT 80.545 2.635 80.555 2.942 ;
      RECT 80.54 2.635 80.545 2.944 ;
      RECT 80.51 2.641 80.54 2.948 ;
      RECT 80.47 2.654 80.51 2.948 ;
      RECT 80.445 2.665 80.47 2.934 ;
      RECT 80.43 2.671 80.445 2.917 ;
      RECT 80.42 2.673 80.43 2.908 ;
      RECT 80.415 2.674 80.42 2.903 ;
      RECT 80.41 2.675 80.415 2.898 ;
      RECT 80.405 2.676 80.41 2.895 ;
      RECT 80.38 2.681 80.405 2.885 ;
      RECT 80.37 2.697 80.38 2.872 ;
      RECT 80.365 2.717 80.37 2.867 ;
      RECT 80.375 2.11 80.38 2.306 ;
      RECT 80.36 2.074 80.375 2.308 ;
      RECT 80.35 2.056 80.36 2.313 ;
      RECT 80.34 2.042 80.35 2.317 ;
      RECT 80.295 2.026 80.34 2.327 ;
      RECT 80.29 2.016 80.295 2.336 ;
      RECT 80.245 2.005 80.29 2.342 ;
      RECT 80.24 1.993 80.245 2.349 ;
      RECT 80.225 1.988 80.24 2.353 ;
      RECT 80.21 1.98 80.225 2.358 ;
      RECT 80.2 1.973 80.21 2.363 ;
      RECT 80.19 1.97 80.2 2.368 ;
      RECT 80.18 1.97 80.19 2.369 ;
      RECT 80.175 1.967 80.18 2.368 ;
      RECT 80.14 1.962 80.165 2.367 ;
      RECT 80.116 1.958 80.14 2.366 ;
      RECT 80.03 1.949 80.116 2.363 ;
      RECT 80.015 1.941 80.03 2.36 ;
      RECT 79.993 1.94 80.015 2.359 ;
      RECT 79.907 1.94 79.993 2.357 ;
      RECT 79.821 1.94 79.907 2.355 ;
      RECT 79.735 1.94 79.821 2.352 ;
      RECT 79.725 1.94 79.735 2.343 ;
      RECT 79.695 1.94 79.725 2.303 ;
      RECT 79.685 1.95 79.695 2.258 ;
      RECT 79.68 1.99 79.685 2.243 ;
      RECT 79.675 2.005 79.68 2.23 ;
      RECT 79.645 2.085 79.675 2.192 ;
      RECT 80.165 1.965 80.175 2.368 ;
      RECT 79.99 2.73 80.005 3.335 ;
      RECT 79.995 2.725 80.005 3.335 ;
      RECT 80.16 2.725 80.165 2.908 ;
      RECT 80.15 2.725 80.16 2.938 ;
      RECT 80.135 2.725 80.15 2.998 ;
      RECT 80.13 2.725 80.135 3.043 ;
      RECT 80.125 2.725 80.13 3.073 ;
      RECT 80.12 2.725 80.125 3.093 ;
      RECT 80.11 2.725 80.12 3.128 ;
      RECT 80.095 2.725 80.11 3.16 ;
      RECT 80.05 2.725 80.095 3.188 ;
      RECT 80.045 2.725 80.05 3.218 ;
      RECT 80.04 2.725 80.045 3.23 ;
      RECT 80.035 2.725 80.04 3.238 ;
      RECT 80.025 2.725 80.035 3.253 ;
      RECT 80.02 2.725 80.025 3.275 ;
      RECT 80.01 2.725 80.02 3.298 ;
      RECT 80.005 2.725 80.01 3.318 ;
      RECT 79.97 2.74 79.99 3.335 ;
      RECT 79.945 2.757 79.97 3.335 ;
      RECT 79.94 2.767 79.945 3.335 ;
      RECT 79.91 2.782 79.94 3.335 ;
      RECT 79.835 2.824 79.91 3.335 ;
      RECT 79.83 2.855 79.835 3.318 ;
      RECT 79.825 2.859 79.83 3.3 ;
      RECT 79.82 2.863 79.825 3.263 ;
      RECT 79.815 3.047 79.82 3.23 ;
      RECT 79.3 3.236 79.386 3.801 ;
      RECT 79.255 3.238 79.42 3.795 ;
      RECT 79.386 3.235 79.42 3.795 ;
      RECT 79.3 3.237 79.505 3.789 ;
      RECT 79.255 3.247 79.515 3.785 ;
      RECT 79.23 3.239 79.505 3.781 ;
      RECT 79.225 3.242 79.505 3.776 ;
      RECT 79.2 3.257 79.515 3.77 ;
      RECT 79.2 3.282 79.555 3.765 ;
      RECT 79.16 3.29 79.555 3.74 ;
      RECT 79.16 3.317 79.57 3.738 ;
      RECT 79.16 3.347 79.58 3.725 ;
      RECT 79.155 3.492 79.58 3.713 ;
      RECT 79.16 3.421 79.6 3.71 ;
      RECT 79.16 3.478 79.605 3.518 ;
      RECT 79.35 2.757 79.52 2.935 ;
      RECT 79.3 2.696 79.35 2.92 ;
      RECT 79.035 2.676 79.3 2.905 ;
      RECT 78.995 2.74 79.47 2.905 ;
      RECT 78.995 2.73 79.425 2.905 ;
      RECT 78.995 2.727 79.415 2.905 ;
      RECT 78.995 2.715 79.405 2.905 ;
      RECT 78.995 2.7 79.35 2.905 ;
      RECT 79.035 2.672 79.236 2.905 ;
      RECT 79.045 2.65 79.236 2.905 ;
      RECT 79.07 2.635 79.15 2.905 ;
      RECT 78.825 3.165 78.945 3.61 ;
      RECT 78.81 3.165 78.945 3.609 ;
      RECT 78.765 3.187 78.945 3.604 ;
      RECT 78.725 3.236 78.945 3.598 ;
      RECT 78.725 3.236 78.95 3.573 ;
      RECT 78.725 3.236 78.97 3.463 ;
      RECT 78.72 3.266 78.97 3.46 ;
      RECT 78.81 3.165 78.98 3.355 ;
      RECT 78.47 1.95 78.475 2.395 ;
      RECT 78.28 1.95 78.3 2.36 ;
      RECT 78.25 1.95 78.255 2.335 ;
      RECT 78.93 2.257 78.945 2.445 ;
      RECT 78.925 2.242 78.93 2.451 ;
      RECT 78.905 2.215 78.925 2.454 ;
      RECT 78.855 2.182 78.905 2.463 ;
      RECT 78.825 2.162 78.855 2.467 ;
      RECT 78.806 2.15 78.825 2.463 ;
      RECT 78.72 2.122 78.806 2.453 ;
      RECT 78.71 2.097 78.72 2.443 ;
      RECT 78.64 2.065 78.71 2.435 ;
      RECT 78.615 2.025 78.64 2.427 ;
      RECT 78.595 2.007 78.615 2.421 ;
      RECT 78.585 1.997 78.595 2.418 ;
      RECT 78.575 1.99 78.585 2.416 ;
      RECT 78.555 1.977 78.575 2.413 ;
      RECT 78.545 1.967 78.555 2.41 ;
      RECT 78.535 1.96 78.545 2.408 ;
      RECT 78.485 1.952 78.535 2.402 ;
      RECT 78.475 1.95 78.485 2.396 ;
      RECT 78.445 1.95 78.47 2.393 ;
      RECT 78.416 1.95 78.445 2.388 ;
      RECT 78.33 1.95 78.416 2.378 ;
      RECT 78.3 1.95 78.33 2.365 ;
      RECT 78.255 1.95 78.28 2.348 ;
      RECT 78.24 1.95 78.25 2.33 ;
      RECT 78.22 1.957 78.24 2.315 ;
      RECT 78.215 1.972 78.22 2.303 ;
      RECT 78.21 1.977 78.215 2.243 ;
      RECT 78.205 1.982 78.21 2.085 ;
      RECT 78.2 1.985 78.205 2.003 ;
      RECT 78.465 2.67 78.551 2.991 ;
      RECT 78.465 2.67 78.585 2.984 ;
      RECT 78.415 2.67 78.585 2.98 ;
      RECT 78.415 2.672 78.671 2.978 ;
      RECT 78.415 2.674 78.695 2.972 ;
      RECT 78.415 2.681 78.705 2.971 ;
      RECT 78.415 2.69 78.71 2.968 ;
      RECT 78.415 2.696 78.715 2.963 ;
      RECT 78.415 2.74 78.72 2.96 ;
      RECT 78.415 2.832 78.725 2.957 ;
      RECT 77.94 3.275 77.975 3.595 ;
      RECT 78.525 3.46 78.53 3.642 ;
      RECT 78.48 3.342 78.525 3.661 ;
      RECT 78.465 3.319 78.48 3.684 ;
      RECT 78.455 3.309 78.465 3.694 ;
      RECT 78.435 3.304 78.455 3.707 ;
      RECT 78.41 3.302 78.435 3.728 ;
      RECT 78.391 3.301 78.41 3.74 ;
      RECT 78.305 3.298 78.391 3.74 ;
      RECT 78.235 3.293 78.305 3.728 ;
      RECT 78.16 3.289 78.235 3.703 ;
      RECT 78.095 3.285 78.16 3.67 ;
      RECT 78.025 3.282 78.095 3.63 ;
      RECT 77.995 3.278 78.025 3.605 ;
      RECT 77.975 3.276 77.995 3.598 ;
      RECT 77.891 3.274 77.94 3.596 ;
      RECT 77.805 3.271 77.891 3.597 ;
      RECT 77.73 3.27 77.805 3.599 ;
      RECT 77.645 3.27 77.73 3.625 ;
      RECT 77.568 3.271 77.645 3.65 ;
      RECT 77.482 3.272 77.568 3.65 ;
      RECT 77.396 3.272 77.482 3.65 ;
      RECT 77.31 3.273 77.396 3.65 ;
      RECT 77.29 3.274 77.31 3.642 ;
      RECT 77.275 3.28 77.29 3.627 ;
      RECT 77.24 3.3 77.275 3.607 ;
      RECT 77.23 3.32 77.24 3.589 ;
      RECT 78.2 2.625 78.205 2.895 ;
      RECT 78.195 2.616 78.2 2.9 ;
      RECT 78.185 2.606 78.195 2.912 ;
      RECT 78.18 2.595 78.185 2.923 ;
      RECT 78.16 2.589 78.18 2.941 ;
      RECT 78.115 2.586 78.16 2.99 ;
      RECT 78.1 2.585 78.115 3.035 ;
      RECT 78.095 2.585 78.1 3.048 ;
      RECT 78.085 2.585 78.095 3.06 ;
      RECT 78.08 2.586 78.085 3.075 ;
      RECT 78.06 2.594 78.08 3.08 ;
      RECT 78.03 2.61 78.06 3.08 ;
      RECT 78.02 2.622 78.025 3.08 ;
      RECT 77.985 2.637 78.02 3.08 ;
      RECT 77.955 2.657 77.985 3.08 ;
      RECT 77.945 2.682 77.955 3.08 ;
      RECT 77.94 2.71 77.945 3.08 ;
      RECT 77.935 2.74 77.94 3.08 ;
      RECT 77.93 2.757 77.935 3.08 ;
      RECT 77.92 2.785 77.93 3.08 ;
      RECT 77.91 2.82 77.92 3.08 ;
      RECT 77.905 2.855 77.91 3.08 ;
      RECT 78.025 2.62 78.03 3.08 ;
      RECT 77.54 2.722 77.725 2.895 ;
      RECT 77.5 2.64 77.685 2.893 ;
      RECT 77.461 2.645 77.685 2.889 ;
      RECT 77.375 2.654 77.685 2.884 ;
      RECT 77.291 2.67 77.69 2.879 ;
      RECT 77.205 2.69 77.715 2.873 ;
      RECT 77.205 2.71 77.72 2.873 ;
      RECT 77.291 2.68 77.715 2.879 ;
      RECT 77.375 2.655 77.69 2.884 ;
      RECT 77.54 2.637 77.685 2.895 ;
      RECT 77.54 2.632 77.64 2.895 ;
      RECT 77.626 2.626 77.64 2.895 ;
      RECT 77.015 1.95 77.02 2.349 ;
      RECT 76.76 1.95 76.795 2.347 ;
      RECT 76.355 1.985 76.36 2.341 ;
      RECT 77.1 1.988 77.105 2.243 ;
      RECT 77.095 1.986 77.1 2.249 ;
      RECT 77.09 1.985 77.095 2.256 ;
      RECT 77.065 1.978 77.09 2.28 ;
      RECT 77.06 1.971 77.065 2.304 ;
      RECT 77.055 1.967 77.06 2.313 ;
      RECT 77.045 1.962 77.055 2.326 ;
      RECT 77.04 1.959 77.045 2.335 ;
      RECT 77.035 1.957 77.04 2.34 ;
      RECT 77.02 1.953 77.035 2.35 ;
      RECT 77.005 1.947 77.015 2.349 ;
      RECT 76.967 1.945 77.005 2.349 ;
      RECT 76.881 1.947 76.967 2.349 ;
      RECT 76.795 1.949 76.881 2.348 ;
      RECT 76.724 1.95 76.76 2.347 ;
      RECT 76.638 1.952 76.724 2.347 ;
      RECT 76.552 1.954 76.638 2.346 ;
      RECT 76.466 1.956 76.552 2.346 ;
      RECT 76.38 1.959 76.466 2.345 ;
      RECT 76.37 1.965 76.38 2.344 ;
      RECT 76.36 1.977 76.37 2.342 ;
      RECT 76.3 2.012 76.355 2.338 ;
      RECT 76.295 2.042 76.3 2.1 ;
      RECT 77.04 3.122 77.055 3.315 ;
      RECT 77.035 3.09 77.04 3.315 ;
      RECT 77.025 3.065 77.035 3.315 ;
      RECT 77.02 3.037 77.025 3.315 ;
      RECT 76.99 2.96 77.02 3.315 ;
      RECT 76.965 2.842 76.99 3.315 ;
      RECT 76.96 2.78 76.965 3.315 ;
      RECT 76.95 2.767 76.96 3.315 ;
      RECT 76.93 2.757 76.95 3.315 ;
      RECT 76.915 2.74 76.93 3.315 ;
      RECT 76.885 2.728 76.915 3.315 ;
      RECT 76.88 2.727 76.885 3.26 ;
      RECT 76.875 2.727 76.88 3.218 ;
      RECT 76.86 2.726 76.875 3.17 ;
      RECT 76.845 2.726 76.86 3.108 ;
      RECT 76.825 2.726 76.845 3.068 ;
      RECT 76.82 2.726 76.825 3.053 ;
      RECT 76.795 2.725 76.82 3.048 ;
      RECT 76.725 2.724 76.795 3.035 ;
      RECT 76.71 2.723 76.725 3.02 ;
      RECT 76.68 2.722 76.71 3.003 ;
      RECT 76.675 2.722 76.68 2.988 ;
      RECT 76.625 2.721 76.675 2.968 ;
      RECT 76.56 2.72 76.625 2.923 ;
      RECT 76.555 2.72 76.56 2.895 ;
      RECT 76.64 3.257 76.645 3.514 ;
      RECT 76.62 3.176 76.64 3.531 ;
      RECT 76.6 3.17 76.62 3.56 ;
      RECT 76.54 3.157 76.6 3.58 ;
      RECT 76.495 3.141 76.54 3.581 ;
      RECT 76.411 3.129 76.495 3.569 ;
      RECT 76.325 3.116 76.411 3.553 ;
      RECT 76.315 3.109 76.325 3.545 ;
      RECT 76.27 3.106 76.315 3.485 ;
      RECT 76.25 3.102 76.27 3.4 ;
      RECT 76.235 3.1 76.25 3.353 ;
      RECT 76.205 3.097 76.235 3.323 ;
      RECT 76.17 3.093 76.205 3.3 ;
      RECT 76.127 3.088 76.17 3.288 ;
      RECT 76.041 3.079 76.127 3.297 ;
      RECT 75.955 3.068 76.041 3.309 ;
      RECT 75.89 3.059 75.955 3.318 ;
      RECT 75.87 3.05 75.89 3.323 ;
      RECT 75.865 3.043 75.87 3.325 ;
      RECT 75.825 3.028 75.865 3.322 ;
      RECT 75.805 3.007 75.825 3.317 ;
      RECT 75.79 2.995 75.805 3.31 ;
      RECT 75.785 2.987 75.79 3.303 ;
      RECT 75.77 2.967 75.785 3.296 ;
      RECT 75.765 2.83 75.77 3.29 ;
      RECT 75.685 2.719 75.765 3.262 ;
      RECT 75.676 2.712 75.685 3.228 ;
      RECT 75.59 2.706 75.676 3.153 ;
      RECT 75.565 2.697 75.59 3.065 ;
      RECT 75.535 2.692 75.565 3.04 ;
      RECT 75.47 2.701 75.535 3.025 ;
      RECT 75.45 2.717 75.47 3 ;
      RECT 75.44 2.723 75.45 2.948 ;
      RECT 75.42 2.745 75.44 2.83 ;
      RECT 76.075 2.71 76.245 2.895 ;
      RECT 76.075 2.71 76.28 2.893 ;
      RECT 76.125 2.62 76.295 2.884 ;
      RECT 76.075 2.777 76.3 2.877 ;
      RECT 76.09 2.655 76.295 2.884 ;
      RECT 75.29 3.388 75.355 3.831 ;
      RECT 75.23 3.413 75.355 3.829 ;
      RECT 75.23 3.413 75.41 3.823 ;
      RECT 75.215 3.438 75.41 3.822 ;
      RECT 75.355 3.375 75.43 3.819 ;
      RECT 75.29 3.4 75.51 3.813 ;
      RECT 75.215 3.439 75.555 3.807 ;
      RECT 75.2 3.466 75.555 3.798 ;
      RECT 75.215 3.459 75.575 3.79 ;
      RECT 75.2 3.468 75.58 3.773 ;
      RECT 75.195 3.485 75.58 3.6 ;
      RECT 75.2 2.207 75.235 2.445 ;
      RECT 75.2 2.207 75.265 2.444 ;
      RECT 75.2 2.207 75.38 2.44 ;
      RECT 75.2 2.207 75.435 2.418 ;
      RECT 75.21 2.15 75.49 2.318 ;
      RECT 75.315 1.99 75.345 2.441 ;
      RECT 75.345 1.985 75.525 2.198 ;
      RECT 75.215 2.126 75.525 2.198 ;
      RECT 75.265 2.022 75.315 2.442 ;
      RECT 75.235 2.078 75.525 2.198 ;
      RECT 74.105 5.02 74.275 6.49 ;
      RECT 74.105 6.315 74.28 6.485 ;
      RECT 73.735 1.74 73.905 2.93 ;
      RECT 73.735 1.74 74.205 1.91 ;
      RECT 73.735 6.97 74.205 7.14 ;
      RECT 73.735 5.95 73.905 7.14 ;
      RECT 72.745 1.74 72.915 2.93 ;
      RECT 72.745 1.74 73.215 1.91 ;
      RECT 72.745 6.97 73.215 7.14 ;
      RECT 72.745 5.95 72.915 7.14 ;
      RECT 70.895 2.635 71.065 3.865 ;
      RECT 70.95 0.855 71.12 2.805 ;
      RECT 70.895 0.575 71.065 1.025 ;
      RECT 70.895 7.855 71.065 8.305 ;
      RECT 70.95 6.075 71.12 8.025 ;
      RECT 70.895 5.015 71.065 6.245 ;
      RECT 70.375 0.575 70.545 3.865 ;
      RECT 70.375 2.075 70.78 2.405 ;
      RECT 70.375 1.235 70.78 1.565 ;
      RECT 70.375 5.015 70.545 8.305 ;
      RECT 70.375 7.315 70.78 7.645 ;
      RECT 70.375 6.475 70.78 6.805 ;
      RECT 68.475 3.392 68.49 3.443 ;
      RECT 68.47 3.372 68.475 3.49 ;
      RECT 68.455 3.362 68.47 3.558 ;
      RECT 68.43 3.342 68.455 3.613 ;
      RECT 68.39 3.327 68.43 3.633 ;
      RECT 68.345 3.321 68.39 3.661 ;
      RECT 68.275 3.311 68.345 3.678 ;
      RECT 68.255 3.303 68.275 3.678 ;
      RECT 68.195 3.297 68.255 3.67 ;
      RECT 68.136 3.288 68.195 3.658 ;
      RECT 68.05 3.277 68.136 3.641 ;
      RECT 68.028 3.268 68.05 3.629 ;
      RECT 67.942 3.261 68.028 3.616 ;
      RECT 67.856 3.248 67.942 3.597 ;
      RECT 67.77 3.236 67.856 3.577 ;
      RECT 67.74 3.225 67.77 3.564 ;
      RECT 67.69 3.211 67.74 3.556 ;
      RECT 67.67 3.2 67.69 3.548 ;
      RECT 67.621 3.189 67.67 3.54 ;
      RECT 67.535 3.168 67.621 3.525 ;
      RECT 67.49 3.155 67.535 3.51 ;
      RECT 67.445 3.155 67.49 3.49 ;
      RECT 67.39 3.155 67.445 3.425 ;
      RECT 67.365 3.155 67.39 3.348 ;
      RECT 67.89 2.892 68.06 3.075 ;
      RECT 67.89 2.892 68.075 3.033 ;
      RECT 67.89 2.892 68.08 2.975 ;
      RECT 67.95 2.66 68.085 2.951 ;
      RECT 67.95 2.664 68.09 2.934 ;
      RECT 67.895 2.827 68.09 2.934 ;
      RECT 67.92 2.672 68.06 3.075 ;
      RECT 67.92 2.676 68.1 2.875 ;
      RECT 67.905 2.762 68.1 2.875 ;
      RECT 67.915 2.692 68.06 3.075 ;
      RECT 67.915 2.695 68.11 2.788 ;
      RECT 67.91 2.712 68.11 2.788 ;
      RECT 67.68 1.932 67.85 2.415 ;
      RECT 67.675 1.927 67.825 2.405 ;
      RECT 67.675 1.934 67.855 2.399 ;
      RECT 67.665 1.928 67.825 2.378 ;
      RECT 67.665 1.944 67.87 2.337 ;
      RECT 67.635 1.929 67.825 2.3 ;
      RECT 67.635 1.959 67.88 2.24 ;
      RECT 67.63 1.931 67.825 2.238 ;
      RECT 67.61 1.94 67.855 2.195 ;
      RECT 67.585 1.956 67.87 2.107 ;
      RECT 67.585 1.975 67.895 2.098 ;
      RECT 67.58 2.012 67.895 2.05 ;
      RECT 67.585 1.992 67.9 2.018 ;
      RECT 67.68 1.926 67.79 2.415 ;
      RECT 67.766 1.925 67.79 2.415 ;
      RECT 67 2.71 67.005 2.921 ;
      RECT 67.6 2.71 67.605 2.895 ;
      RECT 67.665 2.75 67.67 2.863 ;
      RECT 67.66 2.742 67.665 2.869 ;
      RECT 67.655 2.732 67.66 2.877 ;
      RECT 67.65 2.722 67.655 2.886 ;
      RECT 67.645 2.712 67.65 2.89 ;
      RECT 67.605 2.71 67.645 2.893 ;
      RECT 67.577 2.709 67.6 2.897 ;
      RECT 67.491 2.706 67.577 2.904 ;
      RECT 67.405 2.702 67.491 2.915 ;
      RECT 67.385 2.7 67.405 2.921 ;
      RECT 67.367 2.699 67.385 2.924 ;
      RECT 67.281 2.697 67.367 2.931 ;
      RECT 67.195 2.692 67.281 2.944 ;
      RECT 67.176 2.689 67.195 2.949 ;
      RECT 67.09 2.687 67.176 2.94 ;
      RECT 67.08 2.687 67.09 2.933 ;
      RECT 67.005 2.7 67.08 2.927 ;
      RECT 66.99 2.711 67 2.921 ;
      RECT 66.98 2.713 66.99 2.92 ;
      RECT 66.97 2.717 66.98 2.916 ;
      RECT 66.965 2.72 66.97 2.91 ;
      RECT 66.955 2.722 66.965 2.904 ;
      RECT 66.95 2.725 66.955 2.898 ;
      RECT 66.93 3.311 66.935 3.515 ;
      RECT 66.915 3.298 66.93 3.608 ;
      RECT 66.9 3.279 66.915 3.885 ;
      RECT 66.865 3.245 66.9 3.885 ;
      RECT 66.861 3.215 66.865 3.885 ;
      RECT 66.775 3.097 66.861 3.885 ;
      RECT 66.765 2.972 66.775 3.885 ;
      RECT 66.75 2.94 66.765 3.885 ;
      RECT 66.745 2.915 66.75 3.885 ;
      RECT 66.74 2.905 66.745 3.841 ;
      RECT 66.725 2.877 66.74 3.746 ;
      RECT 66.71 2.843 66.725 3.645 ;
      RECT 66.705 2.821 66.71 3.598 ;
      RECT 66.7 2.81 66.705 3.568 ;
      RECT 66.695 2.8 66.7 3.534 ;
      RECT 66.685 2.787 66.695 3.502 ;
      RECT 66.66 2.763 66.685 3.428 ;
      RECT 66.655 2.743 66.66 3.353 ;
      RECT 66.65 2.737 66.655 3.328 ;
      RECT 66.645 2.732 66.65 3.293 ;
      RECT 66.64 2.727 66.645 3.268 ;
      RECT 66.635 2.725 66.64 3.248 ;
      RECT 66.63 2.725 66.635 3.233 ;
      RECT 66.625 2.725 66.63 3.193 ;
      RECT 66.615 2.725 66.625 3.165 ;
      RECT 66.605 2.725 66.615 3.11 ;
      RECT 66.59 2.725 66.605 3.048 ;
      RECT 66.585 2.724 66.59 2.993 ;
      RECT 66.57 2.723 66.585 2.973 ;
      RECT 66.51 2.721 66.57 2.947 ;
      RECT 66.475 2.722 66.51 2.927 ;
      RECT 66.47 2.724 66.475 2.917 ;
      RECT 66.46 2.743 66.47 2.907 ;
      RECT 66.455 2.77 66.46 2.838 ;
      RECT 66.57 2.195 66.74 2.44 ;
      RECT 66.605 1.966 66.74 2.44 ;
      RECT 66.605 1.968 66.75 2.435 ;
      RECT 66.605 1.97 66.775 2.423 ;
      RECT 66.605 1.973 66.8 2.405 ;
      RECT 66.605 1.978 66.85 2.378 ;
      RECT 66.605 1.983 66.87 2.343 ;
      RECT 66.585 1.985 66.88 2.318 ;
      RECT 66.575 2.08 66.88 2.318 ;
      RECT 66.605 1.965 66.715 2.44 ;
      RECT 66.615 1.962 66.71 2.44 ;
      RECT 66.135 3.227 66.325 3.585 ;
      RECT 66.135 3.239 66.36 3.584 ;
      RECT 66.135 3.267 66.38 3.582 ;
      RECT 66.135 3.292 66.385 3.581 ;
      RECT 66.135 3.35 66.4 3.58 ;
      RECT 66.12 3.223 66.28 3.565 ;
      RECT 66.1 3.232 66.325 3.518 ;
      RECT 66.075 3.243 66.36 3.455 ;
      RECT 66.075 3.327 66.395 3.455 ;
      RECT 66.075 3.302 66.39 3.455 ;
      RECT 66.135 3.218 66.28 3.585 ;
      RECT 66.221 3.217 66.28 3.585 ;
      RECT 66.221 3.216 66.265 3.585 ;
      RECT 66.135 7.855 66.305 8.305 ;
      RECT 66.19 6.075 66.36 8.025 ;
      RECT 66.135 5.015 66.305 6.245 ;
      RECT 65.615 5.015 65.785 8.305 ;
      RECT 65.615 7.315 66.02 7.645 ;
      RECT 65.615 6.475 66.02 6.805 ;
      RECT 65.92 2.732 65.925 3.11 ;
      RECT 65.915 2.7 65.92 3.11 ;
      RECT 65.91 2.672 65.915 3.11 ;
      RECT 65.905 2.652 65.91 3.11 ;
      RECT 65.85 2.635 65.905 3.11 ;
      RECT 65.81 2.62 65.85 3.11 ;
      RECT 65.755 2.607 65.81 3.11 ;
      RECT 65.72 2.598 65.755 3.11 ;
      RECT 65.716 2.596 65.72 3.109 ;
      RECT 65.63 2.592 65.716 3.092 ;
      RECT 65.545 2.584 65.63 3.055 ;
      RECT 65.535 2.58 65.545 3.028 ;
      RECT 65.525 2.58 65.535 3.01 ;
      RECT 65.515 2.582 65.525 2.993 ;
      RECT 65.51 2.587 65.515 2.979 ;
      RECT 65.505 2.591 65.51 2.966 ;
      RECT 65.495 2.596 65.505 2.95 ;
      RECT 65.48 2.61 65.495 2.925 ;
      RECT 65.475 2.616 65.48 2.905 ;
      RECT 65.47 2.618 65.475 2.898 ;
      RECT 65.465 2.622 65.47 2.773 ;
      RECT 65.645 3.422 65.89 3.885 ;
      RECT 65.565 3.395 65.885 3.881 ;
      RECT 65.495 3.43 65.89 3.874 ;
      RECT 65.285 3.685 65.89 3.87 ;
      RECT 65.465 3.453 65.89 3.87 ;
      RECT 65.305 3.645 65.89 3.87 ;
      RECT 65.455 3.465 65.89 3.87 ;
      RECT 65.34 3.582 65.89 3.87 ;
      RECT 65.395 3.507 65.89 3.87 ;
      RECT 65.645 3.372 65.885 3.885 ;
      RECT 65.675 3.365 65.885 3.885 ;
      RECT 65.665 3.367 65.885 3.885 ;
      RECT 65.675 3.362 65.805 3.885 ;
      RECT 65.23 1.925 65.316 2.364 ;
      RECT 65.225 1.925 65.316 2.362 ;
      RECT 65.225 1.925 65.385 2.361 ;
      RECT 65.225 1.925 65.415 2.358 ;
      RECT 65.21 1.932 65.415 2.349 ;
      RECT 65.21 1.932 65.42 2.345 ;
      RECT 65.205 1.942 65.42 2.338 ;
      RECT 65.2 1.947 65.42 2.313 ;
      RECT 65.2 1.947 65.435 2.295 ;
      RECT 65.225 1.925 65.455 2.21 ;
      RECT 65.195 1.952 65.455 2.208 ;
      RECT 65.205 1.945 65.46 2.146 ;
      RECT 65.195 2.067 65.465 2.129 ;
      RECT 65.18 1.962 65.46 2.08 ;
      RECT 65.175 1.972 65.46 1.98 ;
      RECT 65.255 2.743 65.26 2.82 ;
      RECT 65.245 2.737 65.255 3.01 ;
      RECT 65.235 2.729 65.245 3.031 ;
      RECT 65.225 2.72 65.235 3.053 ;
      RECT 65.22 2.715 65.225 3.07 ;
      RECT 65.18 2.715 65.22 3.11 ;
      RECT 65.16 2.715 65.18 3.165 ;
      RECT 65.155 2.715 65.16 3.193 ;
      RECT 65.145 2.715 65.155 3.208 ;
      RECT 65.11 2.715 65.145 3.25 ;
      RECT 65.105 2.715 65.11 3.293 ;
      RECT 65.095 2.715 65.105 3.308 ;
      RECT 65.08 2.715 65.095 3.328 ;
      RECT 65.065 2.715 65.08 3.355 ;
      RECT 65.06 2.716 65.065 3.373 ;
      RECT 65.04 2.717 65.06 3.38 ;
      RECT 64.985 2.718 65.04 3.4 ;
      RECT 64.975 2.719 64.985 3.414 ;
      RECT 64.97 2.722 64.975 3.413 ;
      RECT 64.93 2.795 64.97 3.411 ;
      RECT 64.915 2.875 64.93 3.409 ;
      RECT 64.89 2.93 64.915 3.407 ;
      RECT 64.875 2.995 64.89 3.406 ;
      RECT 64.83 3.027 64.875 3.403 ;
      RECT 64.745 3.05 64.83 3.398 ;
      RECT 64.72 3.07 64.745 3.393 ;
      RECT 64.65 3.075 64.72 3.389 ;
      RECT 64.63 3.077 64.65 3.386 ;
      RECT 64.545 3.088 64.63 3.38 ;
      RECT 64.54 3.099 64.545 3.375 ;
      RECT 64.53 3.101 64.54 3.375 ;
      RECT 64.495 3.105 64.53 3.373 ;
      RECT 64.445 3.115 64.495 3.36 ;
      RECT 64.425 3.123 64.445 3.345 ;
      RECT 64.345 3.135 64.425 3.328 ;
      RECT 64.51 2.685 64.68 2.895 ;
      RECT 64.626 2.681 64.68 2.895 ;
      RECT 64.431 2.685 64.68 2.886 ;
      RECT 64.431 2.685 64.685 2.875 ;
      RECT 64.345 2.685 64.685 2.866 ;
      RECT 64.345 2.693 64.695 2.81 ;
      RECT 64.345 2.705 64.7 2.723 ;
      RECT 64.345 2.712 64.705 2.715 ;
      RECT 64.54 2.683 64.68 2.895 ;
      RECT 64.295 3.628 64.54 3.96 ;
      RECT 64.29 3.62 64.295 3.957 ;
      RECT 64.26 3.64 64.54 3.938 ;
      RECT 64.24 3.672 64.54 3.911 ;
      RECT 64.29 3.625 64.467 3.957 ;
      RECT 64.29 3.622 64.381 3.957 ;
      RECT 64.23 1.97 64.4 2.39 ;
      RECT 64.225 1.97 64.4 2.388 ;
      RECT 64.225 1.97 64.425 2.378 ;
      RECT 64.225 1.97 64.445 2.353 ;
      RECT 64.22 1.97 64.445 2.348 ;
      RECT 64.22 1.97 64.455 2.338 ;
      RECT 64.22 1.97 64.46 2.333 ;
      RECT 64.22 1.975 64.465 2.328 ;
      RECT 64.22 2.007 64.48 2.318 ;
      RECT 64.22 2.077 64.505 2.301 ;
      RECT 64.2 2.077 64.505 2.293 ;
      RECT 64.2 2.137 64.515 2.27 ;
      RECT 64.2 2.177 64.525 2.215 ;
      RECT 64.185 1.97 64.46 2.195 ;
      RECT 64.175 1.985 64.465 2.093 ;
      RECT 63.765 3.375 63.935 3.9 ;
      RECT 63.76 3.375 63.935 3.893 ;
      RECT 63.75 3.375 63.94 3.858 ;
      RECT 63.745 3.385 63.94 3.83 ;
      RECT 63.74 3.405 63.94 3.813 ;
      RECT 63.75 3.38 63.945 3.803 ;
      RECT 63.735 3.425 63.945 3.795 ;
      RECT 63.73 3.445 63.945 3.78 ;
      RECT 63.725 3.475 63.945 3.77 ;
      RECT 63.715 3.52 63.945 3.745 ;
      RECT 63.745 3.39 63.95 3.728 ;
      RECT 63.71 3.572 63.95 3.723 ;
      RECT 63.745 3.4 63.955 3.693 ;
      RECT 63.705 3.605 63.955 3.69 ;
      RECT 63.7 3.63 63.955 3.67 ;
      RECT 63.74 3.417 63.965 3.61 ;
      RECT 63.735 3.439 63.975 3.503 ;
      RECT 63.685 2.686 63.7 2.955 ;
      RECT 63.64 2.67 63.685 3 ;
      RECT 63.635 2.658 63.64 3.05 ;
      RECT 63.625 2.654 63.635 3.083 ;
      RECT 63.62 2.651 63.625 3.111 ;
      RECT 63.605 2.653 63.62 3.153 ;
      RECT 63.6 2.657 63.605 3.193 ;
      RECT 63.58 2.662 63.6 3.245 ;
      RECT 63.576 2.667 63.58 3.302 ;
      RECT 63.49 2.686 63.576 3.339 ;
      RECT 63.48 2.707 63.49 3.375 ;
      RECT 63.475 2.715 63.48 3.376 ;
      RECT 63.47 2.757 63.475 3.377 ;
      RECT 63.455 2.845 63.47 3.378 ;
      RECT 63.445 2.995 63.455 3.38 ;
      RECT 63.44 3.04 63.445 3.382 ;
      RECT 63.405 3.082 63.44 3.385 ;
      RECT 63.4 3.1 63.405 3.388 ;
      RECT 63.323 3.106 63.4 3.394 ;
      RECT 63.237 3.12 63.323 3.407 ;
      RECT 63.151 3.134 63.237 3.421 ;
      RECT 63.065 3.148 63.151 3.434 ;
      RECT 63.005 3.16 63.065 3.446 ;
      RECT 62.98 3.167 63.005 3.453 ;
      RECT 62.966 3.17 62.98 3.458 ;
      RECT 62.88 3.178 62.966 3.474 ;
      RECT 62.875 3.185 62.88 3.489 ;
      RECT 62.851 3.185 62.875 3.496 ;
      RECT 62.765 3.188 62.851 3.524 ;
      RECT 62.68 3.192 62.765 3.568 ;
      RECT 62.615 3.196 62.68 3.605 ;
      RECT 62.59 3.199 62.615 3.621 ;
      RECT 62.515 3.212 62.59 3.625 ;
      RECT 62.49 3.23 62.515 3.629 ;
      RECT 62.48 3.237 62.49 3.631 ;
      RECT 62.465 3.24 62.48 3.632 ;
      RECT 62.405 3.252 62.465 3.636 ;
      RECT 62.395 3.266 62.405 3.64 ;
      RECT 62.34 3.276 62.395 3.628 ;
      RECT 62.315 3.297 62.34 3.611 ;
      RECT 62.295 3.317 62.315 3.602 ;
      RECT 62.29 3.33 62.295 3.597 ;
      RECT 62.275 3.342 62.29 3.593 ;
      RECT 63.51 1.997 63.515 2.02 ;
      RECT 63.505 1.988 63.51 2.06 ;
      RECT 63.5 1.986 63.505 2.103 ;
      RECT 63.495 1.977 63.5 2.138 ;
      RECT 63.49 1.967 63.495 2.21 ;
      RECT 63.485 1.957 63.49 2.275 ;
      RECT 63.48 1.954 63.485 2.315 ;
      RECT 63.455 1.948 63.48 2.405 ;
      RECT 63.42 1.936 63.455 2.43 ;
      RECT 63.41 1.927 63.42 2.43 ;
      RECT 63.275 1.925 63.285 2.413 ;
      RECT 63.265 1.925 63.275 2.38 ;
      RECT 63.26 1.925 63.265 2.355 ;
      RECT 63.255 1.925 63.26 2.343 ;
      RECT 63.25 1.925 63.255 2.325 ;
      RECT 63.24 1.925 63.25 2.29 ;
      RECT 63.235 1.927 63.24 2.268 ;
      RECT 63.23 1.933 63.235 2.253 ;
      RECT 63.225 1.939 63.23 2.238 ;
      RECT 63.21 1.951 63.225 2.211 ;
      RECT 63.205 1.962 63.21 2.179 ;
      RECT 63.2 1.972 63.205 2.163 ;
      RECT 63.19 1.98 63.2 2.132 ;
      RECT 63.185 1.99 63.19 2.106 ;
      RECT 63.18 2.047 63.185 2.089 ;
      RECT 63.285 1.925 63.41 2.43 ;
      RECT 63 2.612 63.26 2.91 ;
      RECT 62.995 2.619 63.26 2.908 ;
      RECT 63 2.614 63.275 2.903 ;
      RECT 62.99 2.627 63.275 2.9 ;
      RECT 62.99 2.632 63.28 2.893 ;
      RECT 62.985 2.64 63.28 2.89 ;
      RECT 62.985 2.657 63.285 2.688 ;
      RECT 63 2.609 63.231 2.91 ;
      RECT 63.055 2.608 63.231 2.91 ;
      RECT 63.055 2.605 63.145 2.91 ;
      RECT 63.055 2.602 63.141 2.91 ;
      RECT 62.745 2.875 62.75 2.888 ;
      RECT 62.74 2.842 62.745 2.893 ;
      RECT 62.735 2.797 62.74 2.9 ;
      RECT 62.73 2.752 62.735 2.908 ;
      RECT 62.725 2.72 62.73 2.916 ;
      RECT 62.72 2.68 62.725 2.917 ;
      RECT 62.705 2.66 62.72 2.919 ;
      RECT 62.63 2.642 62.705 2.931 ;
      RECT 62.62 2.635 62.63 2.942 ;
      RECT 62.615 2.635 62.62 2.944 ;
      RECT 62.585 2.641 62.615 2.948 ;
      RECT 62.545 2.654 62.585 2.948 ;
      RECT 62.52 2.665 62.545 2.934 ;
      RECT 62.505 2.671 62.52 2.917 ;
      RECT 62.495 2.673 62.505 2.908 ;
      RECT 62.49 2.674 62.495 2.903 ;
      RECT 62.485 2.675 62.49 2.898 ;
      RECT 62.48 2.676 62.485 2.895 ;
      RECT 62.455 2.681 62.48 2.885 ;
      RECT 62.445 2.697 62.455 2.872 ;
      RECT 62.44 2.717 62.445 2.867 ;
      RECT 62.45 2.11 62.455 2.306 ;
      RECT 62.435 2.074 62.45 2.308 ;
      RECT 62.425 2.056 62.435 2.313 ;
      RECT 62.415 2.042 62.425 2.317 ;
      RECT 62.37 2.026 62.415 2.327 ;
      RECT 62.365 2.016 62.37 2.336 ;
      RECT 62.32 2.005 62.365 2.342 ;
      RECT 62.315 1.993 62.32 2.349 ;
      RECT 62.3 1.988 62.315 2.353 ;
      RECT 62.285 1.98 62.3 2.358 ;
      RECT 62.275 1.973 62.285 2.363 ;
      RECT 62.265 1.97 62.275 2.368 ;
      RECT 62.255 1.97 62.265 2.369 ;
      RECT 62.25 1.967 62.255 2.368 ;
      RECT 62.215 1.962 62.24 2.367 ;
      RECT 62.191 1.958 62.215 2.366 ;
      RECT 62.105 1.949 62.191 2.363 ;
      RECT 62.09 1.941 62.105 2.36 ;
      RECT 62.068 1.94 62.09 2.359 ;
      RECT 61.982 1.94 62.068 2.357 ;
      RECT 61.896 1.94 61.982 2.355 ;
      RECT 61.81 1.94 61.896 2.352 ;
      RECT 61.8 1.94 61.81 2.343 ;
      RECT 61.77 1.94 61.8 2.303 ;
      RECT 61.76 1.95 61.77 2.258 ;
      RECT 61.755 1.99 61.76 2.243 ;
      RECT 61.75 2.005 61.755 2.23 ;
      RECT 61.72 2.085 61.75 2.192 ;
      RECT 62.24 1.965 62.25 2.368 ;
      RECT 62.065 2.73 62.08 3.335 ;
      RECT 62.07 2.725 62.08 3.335 ;
      RECT 62.235 2.725 62.24 2.908 ;
      RECT 62.225 2.725 62.235 2.938 ;
      RECT 62.21 2.725 62.225 2.998 ;
      RECT 62.205 2.725 62.21 3.043 ;
      RECT 62.2 2.725 62.205 3.073 ;
      RECT 62.195 2.725 62.2 3.093 ;
      RECT 62.185 2.725 62.195 3.128 ;
      RECT 62.17 2.725 62.185 3.16 ;
      RECT 62.125 2.725 62.17 3.188 ;
      RECT 62.12 2.725 62.125 3.218 ;
      RECT 62.115 2.725 62.12 3.23 ;
      RECT 62.11 2.725 62.115 3.238 ;
      RECT 62.1 2.725 62.11 3.253 ;
      RECT 62.095 2.725 62.1 3.275 ;
      RECT 62.085 2.725 62.095 3.298 ;
      RECT 62.08 2.725 62.085 3.318 ;
      RECT 62.045 2.74 62.065 3.335 ;
      RECT 62.02 2.757 62.045 3.335 ;
      RECT 62.015 2.767 62.02 3.335 ;
      RECT 61.985 2.782 62.015 3.335 ;
      RECT 61.91 2.824 61.985 3.335 ;
      RECT 61.905 2.855 61.91 3.318 ;
      RECT 61.9 2.859 61.905 3.3 ;
      RECT 61.895 2.863 61.9 3.263 ;
      RECT 61.89 3.047 61.895 3.23 ;
      RECT 61.375 3.236 61.461 3.801 ;
      RECT 61.33 3.238 61.495 3.795 ;
      RECT 61.461 3.235 61.495 3.795 ;
      RECT 61.375 3.237 61.58 3.789 ;
      RECT 61.33 3.247 61.59 3.785 ;
      RECT 61.305 3.239 61.58 3.781 ;
      RECT 61.3 3.242 61.58 3.776 ;
      RECT 61.275 3.257 61.59 3.77 ;
      RECT 61.275 3.282 61.63 3.765 ;
      RECT 61.235 3.29 61.63 3.74 ;
      RECT 61.235 3.317 61.645 3.738 ;
      RECT 61.235 3.347 61.655 3.725 ;
      RECT 61.23 3.492 61.655 3.713 ;
      RECT 61.235 3.421 61.675 3.71 ;
      RECT 61.235 3.478 61.68 3.518 ;
      RECT 61.425 2.757 61.595 2.935 ;
      RECT 61.375 2.696 61.425 2.92 ;
      RECT 61.11 2.676 61.375 2.905 ;
      RECT 61.07 2.74 61.545 2.905 ;
      RECT 61.07 2.73 61.5 2.905 ;
      RECT 61.07 2.727 61.49 2.905 ;
      RECT 61.07 2.715 61.48 2.905 ;
      RECT 61.07 2.7 61.425 2.905 ;
      RECT 61.11 2.672 61.311 2.905 ;
      RECT 61.12 2.65 61.311 2.905 ;
      RECT 61.145 2.635 61.225 2.905 ;
      RECT 60.9 3.165 61.02 3.61 ;
      RECT 60.885 3.165 61.02 3.609 ;
      RECT 60.84 3.187 61.02 3.604 ;
      RECT 60.8 3.236 61.02 3.598 ;
      RECT 60.8 3.236 61.025 3.573 ;
      RECT 60.8 3.236 61.045 3.463 ;
      RECT 60.795 3.266 61.045 3.46 ;
      RECT 60.885 3.165 61.055 3.355 ;
      RECT 60.545 1.95 60.55 2.395 ;
      RECT 60.355 1.95 60.375 2.36 ;
      RECT 60.325 1.95 60.33 2.335 ;
      RECT 61.005 2.257 61.02 2.445 ;
      RECT 61 2.242 61.005 2.451 ;
      RECT 60.98 2.215 61 2.454 ;
      RECT 60.93 2.182 60.98 2.463 ;
      RECT 60.9 2.162 60.93 2.467 ;
      RECT 60.881 2.15 60.9 2.463 ;
      RECT 60.795 2.122 60.881 2.453 ;
      RECT 60.785 2.097 60.795 2.443 ;
      RECT 60.715 2.065 60.785 2.435 ;
      RECT 60.69 2.025 60.715 2.427 ;
      RECT 60.67 2.007 60.69 2.421 ;
      RECT 60.66 1.997 60.67 2.418 ;
      RECT 60.65 1.99 60.66 2.416 ;
      RECT 60.63 1.977 60.65 2.413 ;
      RECT 60.62 1.967 60.63 2.41 ;
      RECT 60.61 1.96 60.62 2.408 ;
      RECT 60.56 1.952 60.61 2.402 ;
      RECT 60.55 1.95 60.56 2.396 ;
      RECT 60.52 1.95 60.545 2.393 ;
      RECT 60.491 1.95 60.52 2.388 ;
      RECT 60.405 1.95 60.491 2.378 ;
      RECT 60.375 1.95 60.405 2.365 ;
      RECT 60.33 1.95 60.355 2.348 ;
      RECT 60.315 1.95 60.325 2.33 ;
      RECT 60.295 1.957 60.315 2.315 ;
      RECT 60.29 1.972 60.295 2.303 ;
      RECT 60.285 1.977 60.29 2.243 ;
      RECT 60.28 1.982 60.285 2.085 ;
      RECT 60.275 1.985 60.28 2.003 ;
      RECT 60.54 2.67 60.626 2.991 ;
      RECT 60.54 2.67 60.66 2.984 ;
      RECT 60.49 2.67 60.66 2.98 ;
      RECT 60.49 2.672 60.746 2.978 ;
      RECT 60.49 2.674 60.77 2.972 ;
      RECT 60.49 2.681 60.78 2.971 ;
      RECT 60.49 2.69 60.785 2.968 ;
      RECT 60.49 2.696 60.79 2.963 ;
      RECT 60.49 2.74 60.795 2.96 ;
      RECT 60.49 2.832 60.8 2.957 ;
      RECT 60.015 3.275 60.05 3.595 ;
      RECT 60.6 3.46 60.605 3.642 ;
      RECT 60.555 3.342 60.6 3.661 ;
      RECT 60.54 3.319 60.555 3.684 ;
      RECT 60.53 3.309 60.54 3.694 ;
      RECT 60.51 3.304 60.53 3.707 ;
      RECT 60.485 3.302 60.51 3.728 ;
      RECT 60.466 3.301 60.485 3.74 ;
      RECT 60.38 3.298 60.466 3.74 ;
      RECT 60.31 3.293 60.38 3.728 ;
      RECT 60.235 3.289 60.31 3.703 ;
      RECT 60.17 3.285 60.235 3.67 ;
      RECT 60.1 3.282 60.17 3.63 ;
      RECT 60.07 3.278 60.1 3.605 ;
      RECT 60.05 3.276 60.07 3.598 ;
      RECT 59.966 3.274 60.015 3.596 ;
      RECT 59.88 3.271 59.966 3.597 ;
      RECT 59.805 3.27 59.88 3.599 ;
      RECT 59.72 3.27 59.805 3.625 ;
      RECT 59.643 3.271 59.72 3.65 ;
      RECT 59.557 3.272 59.643 3.65 ;
      RECT 59.471 3.272 59.557 3.65 ;
      RECT 59.385 3.273 59.471 3.65 ;
      RECT 59.365 3.274 59.385 3.642 ;
      RECT 59.35 3.28 59.365 3.627 ;
      RECT 59.315 3.3 59.35 3.607 ;
      RECT 59.305 3.32 59.315 3.589 ;
      RECT 60.275 2.625 60.28 2.895 ;
      RECT 60.27 2.616 60.275 2.9 ;
      RECT 60.26 2.606 60.27 2.912 ;
      RECT 60.255 2.595 60.26 2.923 ;
      RECT 60.235 2.589 60.255 2.941 ;
      RECT 60.19 2.586 60.235 2.99 ;
      RECT 60.175 2.585 60.19 3.035 ;
      RECT 60.17 2.585 60.175 3.048 ;
      RECT 60.16 2.585 60.17 3.06 ;
      RECT 60.155 2.586 60.16 3.075 ;
      RECT 60.135 2.594 60.155 3.08 ;
      RECT 60.105 2.61 60.135 3.08 ;
      RECT 60.095 2.622 60.1 3.08 ;
      RECT 60.06 2.637 60.095 3.08 ;
      RECT 60.03 2.657 60.06 3.08 ;
      RECT 60.02 2.682 60.03 3.08 ;
      RECT 60.015 2.71 60.02 3.08 ;
      RECT 60.01 2.74 60.015 3.08 ;
      RECT 60.005 2.757 60.01 3.08 ;
      RECT 59.995 2.785 60.005 3.08 ;
      RECT 59.985 2.82 59.995 3.08 ;
      RECT 59.98 2.855 59.985 3.08 ;
      RECT 60.1 2.62 60.105 3.08 ;
      RECT 59.615 2.722 59.8 2.895 ;
      RECT 59.575 2.64 59.76 2.893 ;
      RECT 59.536 2.645 59.76 2.889 ;
      RECT 59.45 2.654 59.76 2.884 ;
      RECT 59.366 2.67 59.765 2.879 ;
      RECT 59.28 2.69 59.79 2.873 ;
      RECT 59.28 2.71 59.795 2.873 ;
      RECT 59.366 2.68 59.79 2.879 ;
      RECT 59.45 2.655 59.765 2.884 ;
      RECT 59.615 2.637 59.76 2.895 ;
      RECT 59.615 2.632 59.715 2.895 ;
      RECT 59.701 2.626 59.715 2.895 ;
      RECT 59.09 1.95 59.095 2.349 ;
      RECT 58.835 1.95 58.87 2.347 ;
      RECT 58.43 1.985 58.435 2.341 ;
      RECT 59.175 1.988 59.18 2.243 ;
      RECT 59.17 1.986 59.175 2.249 ;
      RECT 59.165 1.985 59.17 2.256 ;
      RECT 59.14 1.978 59.165 2.28 ;
      RECT 59.135 1.971 59.14 2.304 ;
      RECT 59.13 1.967 59.135 2.313 ;
      RECT 59.12 1.962 59.13 2.326 ;
      RECT 59.115 1.959 59.12 2.335 ;
      RECT 59.11 1.957 59.115 2.34 ;
      RECT 59.095 1.953 59.11 2.35 ;
      RECT 59.08 1.947 59.09 2.349 ;
      RECT 59.042 1.945 59.08 2.349 ;
      RECT 58.956 1.947 59.042 2.349 ;
      RECT 58.87 1.949 58.956 2.348 ;
      RECT 58.799 1.95 58.835 2.347 ;
      RECT 58.713 1.952 58.799 2.347 ;
      RECT 58.627 1.954 58.713 2.346 ;
      RECT 58.541 1.956 58.627 2.346 ;
      RECT 58.455 1.959 58.541 2.345 ;
      RECT 58.445 1.965 58.455 2.344 ;
      RECT 58.435 1.977 58.445 2.342 ;
      RECT 58.375 2.012 58.43 2.338 ;
      RECT 58.37 2.042 58.375 2.1 ;
      RECT 59.115 3.122 59.13 3.315 ;
      RECT 59.11 3.09 59.115 3.315 ;
      RECT 59.1 3.065 59.11 3.315 ;
      RECT 59.095 3.037 59.1 3.315 ;
      RECT 59.065 2.96 59.095 3.315 ;
      RECT 59.04 2.842 59.065 3.315 ;
      RECT 59.035 2.78 59.04 3.315 ;
      RECT 59.025 2.767 59.035 3.315 ;
      RECT 59.005 2.757 59.025 3.315 ;
      RECT 58.99 2.74 59.005 3.315 ;
      RECT 58.96 2.728 58.99 3.315 ;
      RECT 58.955 2.727 58.96 3.26 ;
      RECT 58.95 2.727 58.955 3.218 ;
      RECT 58.935 2.726 58.95 3.17 ;
      RECT 58.92 2.726 58.935 3.108 ;
      RECT 58.9 2.726 58.92 3.068 ;
      RECT 58.895 2.726 58.9 3.053 ;
      RECT 58.87 2.725 58.895 3.048 ;
      RECT 58.8 2.724 58.87 3.035 ;
      RECT 58.785 2.723 58.8 3.02 ;
      RECT 58.755 2.722 58.785 3.003 ;
      RECT 58.75 2.722 58.755 2.988 ;
      RECT 58.7 2.721 58.75 2.968 ;
      RECT 58.635 2.72 58.7 2.923 ;
      RECT 58.63 2.72 58.635 2.895 ;
      RECT 58.715 3.257 58.72 3.514 ;
      RECT 58.695 3.176 58.715 3.531 ;
      RECT 58.675 3.17 58.695 3.56 ;
      RECT 58.615 3.157 58.675 3.58 ;
      RECT 58.57 3.141 58.615 3.581 ;
      RECT 58.486 3.129 58.57 3.569 ;
      RECT 58.4 3.116 58.486 3.553 ;
      RECT 58.39 3.109 58.4 3.545 ;
      RECT 58.345 3.106 58.39 3.485 ;
      RECT 58.325 3.102 58.345 3.4 ;
      RECT 58.31 3.1 58.325 3.353 ;
      RECT 58.28 3.097 58.31 3.323 ;
      RECT 58.245 3.093 58.28 3.3 ;
      RECT 58.202 3.088 58.245 3.288 ;
      RECT 58.116 3.079 58.202 3.297 ;
      RECT 58.03 3.068 58.116 3.309 ;
      RECT 57.965 3.059 58.03 3.318 ;
      RECT 57.945 3.05 57.965 3.323 ;
      RECT 57.94 3.043 57.945 3.325 ;
      RECT 57.9 3.028 57.94 3.322 ;
      RECT 57.88 3.007 57.9 3.317 ;
      RECT 57.865 2.995 57.88 3.31 ;
      RECT 57.86 2.987 57.865 3.303 ;
      RECT 57.845 2.967 57.86 3.296 ;
      RECT 57.84 2.83 57.845 3.29 ;
      RECT 57.76 2.719 57.84 3.262 ;
      RECT 57.751 2.712 57.76 3.228 ;
      RECT 57.665 2.706 57.751 3.153 ;
      RECT 57.64 2.697 57.665 3.065 ;
      RECT 57.61 2.692 57.64 3.04 ;
      RECT 57.545 2.701 57.61 3.025 ;
      RECT 57.525 2.717 57.545 3 ;
      RECT 57.515 2.723 57.525 2.948 ;
      RECT 57.495 2.745 57.515 2.83 ;
      RECT 58.15 2.71 58.32 2.895 ;
      RECT 58.15 2.71 58.355 2.893 ;
      RECT 58.2 2.62 58.37 2.884 ;
      RECT 58.15 2.777 58.375 2.877 ;
      RECT 58.165 2.655 58.37 2.884 ;
      RECT 57.365 3.388 57.43 3.831 ;
      RECT 57.305 3.413 57.43 3.829 ;
      RECT 57.305 3.413 57.485 3.823 ;
      RECT 57.29 3.438 57.485 3.822 ;
      RECT 57.43 3.375 57.505 3.819 ;
      RECT 57.365 3.4 57.585 3.813 ;
      RECT 57.29 3.439 57.63 3.807 ;
      RECT 57.275 3.466 57.63 3.798 ;
      RECT 57.29 3.459 57.65 3.79 ;
      RECT 57.275 3.468 57.655 3.773 ;
      RECT 57.27 3.485 57.655 3.6 ;
      RECT 57.275 2.207 57.31 2.445 ;
      RECT 57.275 2.207 57.34 2.444 ;
      RECT 57.275 2.207 57.455 2.44 ;
      RECT 57.275 2.207 57.51 2.418 ;
      RECT 57.285 2.15 57.565 2.318 ;
      RECT 57.39 1.99 57.42 2.441 ;
      RECT 57.42 1.985 57.6 2.198 ;
      RECT 57.29 2.126 57.6 2.198 ;
      RECT 57.34 2.022 57.39 2.442 ;
      RECT 57.31 2.078 57.6 2.198 ;
      RECT 56.18 5.02 56.35 6.49 ;
      RECT 56.18 6.315 56.355 6.485 ;
      RECT 55.81 1.74 55.98 2.93 ;
      RECT 55.81 1.74 56.28 1.91 ;
      RECT 55.81 6.97 56.28 7.14 ;
      RECT 55.81 5.95 55.98 7.14 ;
      RECT 54.82 1.74 54.99 2.93 ;
      RECT 54.82 1.74 55.29 1.91 ;
      RECT 54.82 6.97 55.29 7.14 ;
      RECT 54.82 5.95 54.99 7.14 ;
      RECT 52.97 2.635 53.14 3.865 ;
      RECT 53.025 0.855 53.195 2.805 ;
      RECT 52.97 0.575 53.14 1.025 ;
      RECT 52.97 7.855 53.14 8.305 ;
      RECT 53.025 6.075 53.195 8.025 ;
      RECT 52.97 5.015 53.14 6.245 ;
      RECT 52.45 0.575 52.62 3.865 ;
      RECT 52.45 2.075 52.855 2.405 ;
      RECT 52.45 1.235 52.855 1.565 ;
      RECT 52.45 5.015 52.62 8.305 ;
      RECT 52.45 7.315 52.855 7.645 ;
      RECT 52.45 6.475 52.855 6.805 ;
      RECT 50.55 3.392 50.565 3.443 ;
      RECT 50.545 3.372 50.55 3.49 ;
      RECT 50.53 3.362 50.545 3.558 ;
      RECT 50.505 3.342 50.53 3.613 ;
      RECT 50.465 3.327 50.505 3.633 ;
      RECT 50.42 3.321 50.465 3.661 ;
      RECT 50.35 3.311 50.42 3.678 ;
      RECT 50.33 3.303 50.35 3.678 ;
      RECT 50.27 3.297 50.33 3.67 ;
      RECT 50.211 3.288 50.27 3.658 ;
      RECT 50.125 3.277 50.211 3.641 ;
      RECT 50.103 3.268 50.125 3.629 ;
      RECT 50.017 3.261 50.103 3.616 ;
      RECT 49.931 3.248 50.017 3.597 ;
      RECT 49.845 3.236 49.931 3.577 ;
      RECT 49.815 3.225 49.845 3.564 ;
      RECT 49.765 3.211 49.815 3.556 ;
      RECT 49.745 3.2 49.765 3.548 ;
      RECT 49.696 3.189 49.745 3.54 ;
      RECT 49.61 3.168 49.696 3.525 ;
      RECT 49.565 3.155 49.61 3.51 ;
      RECT 49.52 3.155 49.565 3.49 ;
      RECT 49.465 3.155 49.52 3.425 ;
      RECT 49.44 3.155 49.465 3.348 ;
      RECT 49.965 2.892 50.135 3.075 ;
      RECT 49.965 2.892 50.15 3.033 ;
      RECT 49.965 2.892 50.155 2.975 ;
      RECT 50.025 2.66 50.16 2.951 ;
      RECT 50.025 2.664 50.165 2.934 ;
      RECT 49.97 2.827 50.165 2.934 ;
      RECT 49.995 2.672 50.135 3.075 ;
      RECT 49.995 2.676 50.175 2.875 ;
      RECT 49.98 2.762 50.175 2.875 ;
      RECT 49.99 2.692 50.135 3.075 ;
      RECT 49.99 2.695 50.185 2.788 ;
      RECT 49.985 2.712 50.185 2.788 ;
      RECT 49.755 1.932 49.925 2.415 ;
      RECT 49.75 1.927 49.9 2.405 ;
      RECT 49.75 1.934 49.93 2.399 ;
      RECT 49.74 1.928 49.9 2.378 ;
      RECT 49.74 1.944 49.945 2.337 ;
      RECT 49.71 1.929 49.9 2.3 ;
      RECT 49.71 1.959 49.955 2.24 ;
      RECT 49.705 1.931 49.9 2.238 ;
      RECT 49.685 1.94 49.93 2.195 ;
      RECT 49.66 1.956 49.945 2.107 ;
      RECT 49.66 1.975 49.97 2.098 ;
      RECT 49.655 2.012 49.97 2.05 ;
      RECT 49.66 1.992 49.975 2.018 ;
      RECT 49.755 1.926 49.865 2.415 ;
      RECT 49.841 1.925 49.865 2.415 ;
      RECT 49.075 2.71 49.08 2.921 ;
      RECT 49.675 2.71 49.68 2.895 ;
      RECT 49.74 2.75 49.745 2.863 ;
      RECT 49.735 2.742 49.74 2.869 ;
      RECT 49.73 2.732 49.735 2.877 ;
      RECT 49.725 2.722 49.73 2.886 ;
      RECT 49.72 2.712 49.725 2.89 ;
      RECT 49.68 2.71 49.72 2.893 ;
      RECT 49.652 2.709 49.675 2.897 ;
      RECT 49.566 2.706 49.652 2.904 ;
      RECT 49.48 2.702 49.566 2.915 ;
      RECT 49.46 2.7 49.48 2.921 ;
      RECT 49.442 2.699 49.46 2.924 ;
      RECT 49.356 2.697 49.442 2.931 ;
      RECT 49.27 2.692 49.356 2.944 ;
      RECT 49.251 2.689 49.27 2.949 ;
      RECT 49.165 2.687 49.251 2.94 ;
      RECT 49.155 2.687 49.165 2.933 ;
      RECT 49.08 2.7 49.155 2.927 ;
      RECT 49.065 2.711 49.075 2.921 ;
      RECT 49.055 2.713 49.065 2.92 ;
      RECT 49.045 2.717 49.055 2.916 ;
      RECT 49.04 2.72 49.045 2.91 ;
      RECT 49.03 2.722 49.04 2.904 ;
      RECT 49.025 2.725 49.03 2.898 ;
      RECT 49.005 3.311 49.01 3.515 ;
      RECT 48.99 3.298 49.005 3.608 ;
      RECT 48.975 3.279 48.99 3.885 ;
      RECT 48.94 3.245 48.975 3.885 ;
      RECT 48.936 3.215 48.94 3.885 ;
      RECT 48.85 3.097 48.936 3.885 ;
      RECT 48.84 2.972 48.85 3.885 ;
      RECT 48.825 2.94 48.84 3.885 ;
      RECT 48.82 2.915 48.825 3.885 ;
      RECT 48.815 2.905 48.82 3.841 ;
      RECT 48.8 2.877 48.815 3.746 ;
      RECT 48.785 2.843 48.8 3.645 ;
      RECT 48.78 2.821 48.785 3.598 ;
      RECT 48.775 2.81 48.78 3.568 ;
      RECT 48.77 2.8 48.775 3.534 ;
      RECT 48.76 2.787 48.77 3.502 ;
      RECT 48.735 2.763 48.76 3.428 ;
      RECT 48.73 2.743 48.735 3.353 ;
      RECT 48.725 2.737 48.73 3.328 ;
      RECT 48.72 2.732 48.725 3.293 ;
      RECT 48.715 2.727 48.72 3.268 ;
      RECT 48.71 2.725 48.715 3.248 ;
      RECT 48.705 2.725 48.71 3.233 ;
      RECT 48.7 2.725 48.705 3.193 ;
      RECT 48.69 2.725 48.7 3.165 ;
      RECT 48.68 2.725 48.69 3.11 ;
      RECT 48.665 2.725 48.68 3.048 ;
      RECT 48.66 2.724 48.665 2.993 ;
      RECT 48.645 2.723 48.66 2.973 ;
      RECT 48.585 2.721 48.645 2.947 ;
      RECT 48.55 2.722 48.585 2.927 ;
      RECT 48.545 2.724 48.55 2.917 ;
      RECT 48.535 2.743 48.545 2.907 ;
      RECT 48.53 2.77 48.535 2.838 ;
      RECT 48.645 2.195 48.815 2.44 ;
      RECT 48.68 1.966 48.815 2.44 ;
      RECT 48.68 1.968 48.825 2.435 ;
      RECT 48.68 1.97 48.85 2.423 ;
      RECT 48.68 1.973 48.875 2.405 ;
      RECT 48.68 1.978 48.925 2.378 ;
      RECT 48.68 1.983 48.945 2.343 ;
      RECT 48.66 1.985 48.955 2.318 ;
      RECT 48.65 2.08 48.955 2.318 ;
      RECT 48.68 1.965 48.79 2.44 ;
      RECT 48.69 1.962 48.785 2.44 ;
      RECT 48.21 3.227 48.4 3.585 ;
      RECT 48.21 3.239 48.435 3.584 ;
      RECT 48.21 3.267 48.455 3.582 ;
      RECT 48.21 3.292 48.46 3.581 ;
      RECT 48.21 3.35 48.475 3.58 ;
      RECT 48.195 3.223 48.355 3.565 ;
      RECT 48.175 3.232 48.4 3.518 ;
      RECT 48.15 3.243 48.435 3.455 ;
      RECT 48.15 3.327 48.47 3.455 ;
      RECT 48.15 3.302 48.465 3.455 ;
      RECT 48.21 3.218 48.355 3.585 ;
      RECT 48.296 3.217 48.355 3.585 ;
      RECT 48.296 3.216 48.34 3.585 ;
      RECT 48.21 7.855 48.38 8.305 ;
      RECT 48.265 6.075 48.435 8.025 ;
      RECT 48.21 5.015 48.38 6.245 ;
      RECT 47.69 5.015 47.86 8.305 ;
      RECT 47.69 7.315 48.095 7.645 ;
      RECT 47.69 6.475 48.095 6.805 ;
      RECT 47.995 2.732 48 3.11 ;
      RECT 47.99 2.7 47.995 3.11 ;
      RECT 47.985 2.672 47.99 3.11 ;
      RECT 47.98 2.652 47.985 3.11 ;
      RECT 47.925 2.635 47.98 3.11 ;
      RECT 47.885 2.62 47.925 3.11 ;
      RECT 47.83 2.607 47.885 3.11 ;
      RECT 47.795 2.598 47.83 3.11 ;
      RECT 47.791 2.596 47.795 3.109 ;
      RECT 47.705 2.592 47.791 3.092 ;
      RECT 47.62 2.584 47.705 3.055 ;
      RECT 47.61 2.58 47.62 3.028 ;
      RECT 47.6 2.58 47.61 3.01 ;
      RECT 47.59 2.582 47.6 2.993 ;
      RECT 47.585 2.587 47.59 2.979 ;
      RECT 47.58 2.591 47.585 2.966 ;
      RECT 47.57 2.596 47.58 2.95 ;
      RECT 47.555 2.61 47.57 2.925 ;
      RECT 47.55 2.616 47.555 2.905 ;
      RECT 47.545 2.618 47.55 2.898 ;
      RECT 47.54 2.622 47.545 2.773 ;
      RECT 47.72 3.422 47.965 3.885 ;
      RECT 47.64 3.395 47.96 3.881 ;
      RECT 47.57 3.43 47.965 3.874 ;
      RECT 47.36 3.685 47.965 3.87 ;
      RECT 47.54 3.453 47.965 3.87 ;
      RECT 47.38 3.645 47.965 3.87 ;
      RECT 47.53 3.465 47.965 3.87 ;
      RECT 47.415 3.582 47.965 3.87 ;
      RECT 47.47 3.507 47.965 3.87 ;
      RECT 47.72 3.372 47.96 3.885 ;
      RECT 47.75 3.365 47.96 3.885 ;
      RECT 47.74 3.367 47.96 3.885 ;
      RECT 47.75 3.362 47.88 3.885 ;
      RECT 47.305 1.925 47.391 2.364 ;
      RECT 47.3 1.925 47.391 2.362 ;
      RECT 47.3 1.925 47.46 2.361 ;
      RECT 47.3 1.925 47.49 2.358 ;
      RECT 47.285 1.932 47.49 2.349 ;
      RECT 47.285 1.932 47.495 2.345 ;
      RECT 47.28 1.942 47.495 2.338 ;
      RECT 47.275 1.947 47.495 2.313 ;
      RECT 47.275 1.947 47.51 2.295 ;
      RECT 47.3 1.925 47.53 2.21 ;
      RECT 47.27 1.952 47.53 2.208 ;
      RECT 47.28 1.945 47.535 2.146 ;
      RECT 47.27 2.067 47.54 2.129 ;
      RECT 47.255 1.962 47.535 2.08 ;
      RECT 47.25 1.972 47.535 1.98 ;
      RECT 47.33 2.743 47.335 2.82 ;
      RECT 47.32 2.737 47.33 3.01 ;
      RECT 47.31 2.729 47.32 3.031 ;
      RECT 47.3 2.72 47.31 3.053 ;
      RECT 47.295 2.715 47.3 3.07 ;
      RECT 47.255 2.715 47.295 3.11 ;
      RECT 47.235 2.715 47.255 3.165 ;
      RECT 47.23 2.715 47.235 3.193 ;
      RECT 47.22 2.715 47.23 3.208 ;
      RECT 47.185 2.715 47.22 3.25 ;
      RECT 47.18 2.715 47.185 3.293 ;
      RECT 47.17 2.715 47.18 3.308 ;
      RECT 47.155 2.715 47.17 3.328 ;
      RECT 47.14 2.715 47.155 3.355 ;
      RECT 47.135 2.716 47.14 3.373 ;
      RECT 47.115 2.717 47.135 3.38 ;
      RECT 47.06 2.718 47.115 3.4 ;
      RECT 47.05 2.719 47.06 3.414 ;
      RECT 47.045 2.722 47.05 3.413 ;
      RECT 47.005 2.795 47.045 3.411 ;
      RECT 46.99 2.875 47.005 3.409 ;
      RECT 46.965 2.93 46.99 3.407 ;
      RECT 46.95 2.995 46.965 3.406 ;
      RECT 46.905 3.027 46.95 3.403 ;
      RECT 46.82 3.05 46.905 3.398 ;
      RECT 46.795 3.07 46.82 3.393 ;
      RECT 46.725 3.075 46.795 3.389 ;
      RECT 46.705 3.077 46.725 3.386 ;
      RECT 46.62 3.088 46.705 3.38 ;
      RECT 46.615 3.099 46.62 3.375 ;
      RECT 46.605 3.101 46.615 3.375 ;
      RECT 46.57 3.105 46.605 3.373 ;
      RECT 46.52 3.115 46.57 3.36 ;
      RECT 46.5 3.123 46.52 3.345 ;
      RECT 46.42 3.135 46.5 3.328 ;
      RECT 46.585 2.685 46.755 2.895 ;
      RECT 46.701 2.681 46.755 2.895 ;
      RECT 46.506 2.685 46.755 2.886 ;
      RECT 46.506 2.685 46.76 2.875 ;
      RECT 46.42 2.685 46.76 2.866 ;
      RECT 46.42 2.693 46.77 2.81 ;
      RECT 46.42 2.705 46.775 2.723 ;
      RECT 46.42 2.712 46.78 2.715 ;
      RECT 46.615 2.683 46.755 2.895 ;
      RECT 46.37 3.628 46.615 3.96 ;
      RECT 46.365 3.62 46.37 3.957 ;
      RECT 46.335 3.64 46.615 3.938 ;
      RECT 46.315 3.672 46.615 3.911 ;
      RECT 46.365 3.625 46.542 3.957 ;
      RECT 46.365 3.622 46.456 3.957 ;
      RECT 46.305 1.97 46.475 2.39 ;
      RECT 46.3 1.97 46.475 2.388 ;
      RECT 46.3 1.97 46.5 2.378 ;
      RECT 46.3 1.97 46.52 2.353 ;
      RECT 46.295 1.97 46.52 2.348 ;
      RECT 46.295 1.97 46.53 2.338 ;
      RECT 46.295 1.97 46.535 2.333 ;
      RECT 46.295 1.975 46.54 2.328 ;
      RECT 46.295 2.007 46.555 2.318 ;
      RECT 46.295 2.077 46.58 2.301 ;
      RECT 46.275 2.077 46.58 2.293 ;
      RECT 46.275 2.137 46.59 2.27 ;
      RECT 46.275 2.177 46.6 2.215 ;
      RECT 46.26 1.97 46.535 2.195 ;
      RECT 46.25 1.985 46.54 2.093 ;
      RECT 45.84 3.375 46.01 3.9 ;
      RECT 45.835 3.375 46.01 3.893 ;
      RECT 45.825 3.375 46.015 3.858 ;
      RECT 45.82 3.385 46.015 3.83 ;
      RECT 45.815 3.405 46.015 3.813 ;
      RECT 45.825 3.38 46.02 3.803 ;
      RECT 45.81 3.425 46.02 3.795 ;
      RECT 45.805 3.445 46.02 3.78 ;
      RECT 45.8 3.475 46.02 3.77 ;
      RECT 45.79 3.52 46.02 3.745 ;
      RECT 45.82 3.39 46.025 3.728 ;
      RECT 45.785 3.572 46.025 3.723 ;
      RECT 45.82 3.4 46.03 3.693 ;
      RECT 45.78 3.605 46.03 3.69 ;
      RECT 45.775 3.63 46.03 3.67 ;
      RECT 45.815 3.417 46.04 3.61 ;
      RECT 45.81 3.439 46.05 3.503 ;
      RECT 45.76 2.686 45.775 2.955 ;
      RECT 45.715 2.67 45.76 3 ;
      RECT 45.71 2.658 45.715 3.05 ;
      RECT 45.7 2.654 45.71 3.083 ;
      RECT 45.695 2.651 45.7 3.111 ;
      RECT 45.68 2.653 45.695 3.153 ;
      RECT 45.675 2.657 45.68 3.193 ;
      RECT 45.655 2.662 45.675 3.245 ;
      RECT 45.651 2.667 45.655 3.302 ;
      RECT 45.565 2.686 45.651 3.339 ;
      RECT 45.555 2.707 45.565 3.375 ;
      RECT 45.55 2.715 45.555 3.376 ;
      RECT 45.545 2.757 45.55 3.377 ;
      RECT 45.53 2.845 45.545 3.378 ;
      RECT 45.52 2.995 45.53 3.38 ;
      RECT 45.515 3.04 45.52 3.382 ;
      RECT 45.48 3.082 45.515 3.385 ;
      RECT 45.475 3.1 45.48 3.388 ;
      RECT 45.398 3.106 45.475 3.394 ;
      RECT 45.312 3.12 45.398 3.407 ;
      RECT 45.226 3.134 45.312 3.421 ;
      RECT 45.14 3.148 45.226 3.434 ;
      RECT 45.08 3.16 45.14 3.446 ;
      RECT 45.055 3.167 45.08 3.453 ;
      RECT 45.041 3.17 45.055 3.458 ;
      RECT 44.955 3.178 45.041 3.474 ;
      RECT 44.95 3.185 44.955 3.489 ;
      RECT 44.926 3.185 44.95 3.496 ;
      RECT 44.84 3.188 44.926 3.524 ;
      RECT 44.755 3.192 44.84 3.568 ;
      RECT 44.69 3.196 44.755 3.605 ;
      RECT 44.665 3.199 44.69 3.621 ;
      RECT 44.59 3.212 44.665 3.625 ;
      RECT 44.565 3.23 44.59 3.629 ;
      RECT 44.555 3.237 44.565 3.631 ;
      RECT 44.54 3.24 44.555 3.632 ;
      RECT 44.48 3.252 44.54 3.636 ;
      RECT 44.47 3.266 44.48 3.64 ;
      RECT 44.415 3.276 44.47 3.628 ;
      RECT 44.39 3.297 44.415 3.611 ;
      RECT 44.37 3.317 44.39 3.602 ;
      RECT 44.365 3.33 44.37 3.597 ;
      RECT 44.35 3.342 44.365 3.593 ;
      RECT 45.585 1.997 45.59 2.02 ;
      RECT 45.58 1.988 45.585 2.06 ;
      RECT 45.575 1.986 45.58 2.103 ;
      RECT 45.57 1.977 45.575 2.138 ;
      RECT 45.565 1.967 45.57 2.21 ;
      RECT 45.56 1.957 45.565 2.275 ;
      RECT 45.555 1.954 45.56 2.315 ;
      RECT 45.53 1.948 45.555 2.405 ;
      RECT 45.495 1.936 45.53 2.43 ;
      RECT 45.485 1.927 45.495 2.43 ;
      RECT 45.35 1.925 45.36 2.413 ;
      RECT 45.34 1.925 45.35 2.38 ;
      RECT 45.335 1.925 45.34 2.355 ;
      RECT 45.33 1.925 45.335 2.343 ;
      RECT 45.325 1.925 45.33 2.325 ;
      RECT 45.315 1.925 45.325 2.29 ;
      RECT 45.31 1.927 45.315 2.268 ;
      RECT 45.305 1.933 45.31 2.253 ;
      RECT 45.3 1.939 45.305 2.238 ;
      RECT 45.285 1.951 45.3 2.211 ;
      RECT 45.28 1.962 45.285 2.179 ;
      RECT 45.275 1.972 45.28 2.163 ;
      RECT 45.265 1.98 45.275 2.132 ;
      RECT 45.26 1.99 45.265 2.106 ;
      RECT 45.255 2.047 45.26 2.089 ;
      RECT 45.36 1.925 45.485 2.43 ;
      RECT 45.075 2.612 45.335 2.91 ;
      RECT 45.07 2.619 45.335 2.908 ;
      RECT 45.075 2.614 45.35 2.903 ;
      RECT 45.065 2.627 45.35 2.9 ;
      RECT 45.065 2.632 45.355 2.893 ;
      RECT 45.06 2.64 45.355 2.89 ;
      RECT 45.06 2.657 45.36 2.688 ;
      RECT 45.075 2.609 45.306 2.91 ;
      RECT 45.13 2.608 45.306 2.91 ;
      RECT 45.13 2.605 45.22 2.91 ;
      RECT 45.13 2.602 45.216 2.91 ;
      RECT 44.82 2.875 44.825 2.888 ;
      RECT 44.815 2.842 44.82 2.893 ;
      RECT 44.81 2.797 44.815 2.9 ;
      RECT 44.805 2.752 44.81 2.908 ;
      RECT 44.8 2.72 44.805 2.916 ;
      RECT 44.795 2.68 44.8 2.917 ;
      RECT 44.78 2.66 44.795 2.919 ;
      RECT 44.705 2.642 44.78 2.931 ;
      RECT 44.695 2.635 44.705 2.942 ;
      RECT 44.69 2.635 44.695 2.944 ;
      RECT 44.66 2.641 44.69 2.948 ;
      RECT 44.62 2.654 44.66 2.948 ;
      RECT 44.595 2.665 44.62 2.934 ;
      RECT 44.58 2.671 44.595 2.917 ;
      RECT 44.57 2.673 44.58 2.908 ;
      RECT 44.565 2.674 44.57 2.903 ;
      RECT 44.56 2.675 44.565 2.898 ;
      RECT 44.555 2.676 44.56 2.895 ;
      RECT 44.53 2.681 44.555 2.885 ;
      RECT 44.52 2.697 44.53 2.872 ;
      RECT 44.515 2.717 44.52 2.867 ;
      RECT 44.525 2.11 44.53 2.306 ;
      RECT 44.51 2.074 44.525 2.308 ;
      RECT 44.5 2.056 44.51 2.313 ;
      RECT 44.49 2.042 44.5 2.317 ;
      RECT 44.445 2.026 44.49 2.327 ;
      RECT 44.44 2.016 44.445 2.336 ;
      RECT 44.395 2.005 44.44 2.342 ;
      RECT 44.39 1.993 44.395 2.349 ;
      RECT 44.375 1.988 44.39 2.353 ;
      RECT 44.36 1.98 44.375 2.358 ;
      RECT 44.35 1.973 44.36 2.363 ;
      RECT 44.34 1.97 44.35 2.368 ;
      RECT 44.33 1.97 44.34 2.369 ;
      RECT 44.325 1.967 44.33 2.368 ;
      RECT 44.29 1.962 44.315 2.367 ;
      RECT 44.266 1.958 44.29 2.366 ;
      RECT 44.18 1.949 44.266 2.363 ;
      RECT 44.165 1.941 44.18 2.36 ;
      RECT 44.143 1.94 44.165 2.359 ;
      RECT 44.057 1.94 44.143 2.357 ;
      RECT 43.971 1.94 44.057 2.355 ;
      RECT 43.885 1.94 43.971 2.352 ;
      RECT 43.875 1.94 43.885 2.343 ;
      RECT 43.845 1.94 43.875 2.303 ;
      RECT 43.835 1.95 43.845 2.258 ;
      RECT 43.83 1.99 43.835 2.243 ;
      RECT 43.825 2.005 43.83 2.23 ;
      RECT 43.795 2.085 43.825 2.192 ;
      RECT 44.315 1.965 44.325 2.368 ;
      RECT 44.14 2.73 44.155 3.335 ;
      RECT 44.145 2.725 44.155 3.335 ;
      RECT 44.31 2.725 44.315 2.908 ;
      RECT 44.3 2.725 44.31 2.938 ;
      RECT 44.285 2.725 44.3 2.998 ;
      RECT 44.28 2.725 44.285 3.043 ;
      RECT 44.275 2.725 44.28 3.073 ;
      RECT 44.27 2.725 44.275 3.093 ;
      RECT 44.26 2.725 44.27 3.128 ;
      RECT 44.245 2.725 44.26 3.16 ;
      RECT 44.2 2.725 44.245 3.188 ;
      RECT 44.195 2.725 44.2 3.218 ;
      RECT 44.19 2.725 44.195 3.23 ;
      RECT 44.185 2.725 44.19 3.238 ;
      RECT 44.175 2.725 44.185 3.253 ;
      RECT 44.17 2.725 44.175 3.275 ;
      RECT 44.16 2.725 44.17 3.298 ;
      RECT 44.155 2.725 44.16 3.318 ;
      RECT 44.12 2.74 44.14 3.335 ;
      RECT 44.095 2.757 44.12 3.335 ;
      RECT 44.09 2.767 44.095 3.335 ;
      RECT 44.06 2.782 44.09 3.335 ;
      RECT 43.985 2.824 44.06 3.335 ;
      RECT 43.98 2.855 43.985 3.318 ;
      RECT 43.975 2.859 43.98 3.3 ;
      RECT 43.97 2.863 43.975 3.263 ;
      RECT 43.965 3.047 43.97 3.23 ;
      RECT 43.45 3.236 43.536 3.801 ;
      RECT 43.405 3.238 43.57 3.795 ;
      RECT 43.536 3.235 43.57 3.795 ;
      RECT 43.45 3.237 43.655 3.789 ;
      RECT 43.405 3.247 43.665 3.785 ;
      RECT 43.38 3.239 43.655 3.781 ;
      RECT 43.375 3.242 43.655 3.776 ;
      RECT 43.35 3.257 43.665 3.77 ;
      RECT 43.35 3.282 43.705 3.765 ;
      RECT 43.31 3.29 43.705 3.74 ;
      RECT 43.31 3.317 43.72 3.738 ;
      RECT 43.31 3.347 43.73 3.725 ;
      RECT 43.305 3.492 43.73 3.713 ;
      RECT 43.31 3.421 43.75 3.71 ;
      RECT 43.31 3.478 43.755 3.518 ;
      RECT 43.5 2.757 43.67 2.935 ;
      RECT 43.45 2.696 43.5 2.92 ;
      RECT 43.185 2.676 43.45 2.905 ;
      RECT 43.145 2.74 43.62 2.905 ;
      RECT 43.145 2.73 43.575 2.905 ;
      RECT 43.145 2.727 43.565 2.905 ;
      RECT 43.145 2.715 43.555 2.905 ;
      RECT 43.145 2.7 43.5 2.905 ;
      RECT 43.185 2.672 43.386 2.905 ;
      RECT 43.195 2.65 43.386 2.905 ;
      RECT 43.22 2.635 43.3 2.905 ;
      RECT 42.975 3.165 43.095 3.61 ;
      RECT 42.96 3.165 43.095 3.609 ;
      RECT 42.915 3.187 43.095 3.604 ;
      RECT 42.875 3.236 43.095 3.598 ;
      RECT 42.875 3.236 43.1 3.573 ;
      RECT 42.875 3.236 43.12 3.463 ;
      RECT 42.87 3.266 43.12 3.46 ;
      RECT 42.96 3.165 43.13 3.355 ;
      RECT 42.62 1.95 42.625 2.395 ;
      RECT 42.43 1.95 42.45 2.36 ;
      RECT 42.4 1.95 42.405 2.335 ;
      RECT 43.08 2.257 43.095 2.445 ;
      RECT 43.075 2.242 43.08 2.451 ;
      RECT 43.055 2.215 43.075 2.454 ;
      RECT 43.005 2.182 43.055 2.463 ;
      RECT 42.975 2.162 43.005 2.467 ;
      RECT 42.956 2.15 42.975 2.463 ;
      RECT 42.87 2.122 42.956 2.453 ;
      RECT 42.86 2.097 42.87 2.443 ;
      RECT 42.79 2.065 42.86 2.435 ;
      RECT 42.765 2.025 42.79 2.427 ;
      RECT 42.745 2.007 42.765 2.421 ;
      RECT 42.735 1.997 42.745 2.418 ;
      RECT 42.725 1.99 42.735 2.416 ;
      RECT 42.705 1.977 42.725 2.413 ;
      RECT 42.695 1.967 42.705 2.41 ;
      RECT 42.685 1.96 42.695 2.408 ;
      RECT 42.635 1.952 42.685 2.402 ;
      RECT 42.625 1.95 42.635 2.396 ;
      RECT 42.595 1.95 42.62 2.393 ;
      RECT 42.566 1.95 42.595 2.388 ;
      RECT 42.48 1.95 42.566 2.378 ;
      RECT 42.45 1.95 42.48 2.365 ;
      RECT 42.405 1.95 42.43 2.348 ;
      RECT 42.39 1.95 42.4 2.33 ;
      RECT 42.37 1.957 42.39 2.315 ;
      RECT 42.365 1.972 42.37 2.303 ;
      RECT 42.36 1.977 42.365 2.243 ;
      RECT 42.355 1.982 42.36 2.085 ;
      RECT 42.35 1.985 42.355 2.003 ;
      RECT 42.615 2.67 42.701 2.991 ;
      RECT 42.615 2.67 42.735 2.984 ;
      RECT 42.565 2.67 42.735 2.98 ;
      RECT 42.565 2.672 42.821 2.978 ;
      RECT 42.565 2.674 42.845 2.972 ;
      RECT 42.565 2.681 42.855 2.971 ;
      RECT 42.565 2.69 42.86 2.968 ;
      RECT 42.565 2.696 42.865 2.963 ;
      RECT 42.565 2.74 42.87 2.96 ;
      RECT 42.565 2.832 42.875 2.957 ;
      RECT 42.09 3.275 42.125 3.595 ;
      RECT 42.675 3.46 42.68 3.642 ;
      RECT 42.63 3.342 42.675 3.661 ;
      RECT 42.615 3.319 42.63 3.684 ;
      RECT 42.605 3.309 42.615 3.694 ;
      RECT 42.585 3.304 42.605 3.707 ;
      RECT 42.56 3.302 42.585 3.728 ;
      RECT 42.541 3.301 42.56 3.74 ;
      RECT 42.455 3.298 42.541 3.74 ;
      RECT 42.385 3.293 42.455 3.728 ;
      RECT 42.31 3.289 42.385 3.703 ;
      RECT 42.245 3.285 42.31 3.67 ;
      RECT 42.175 3.282 42.245 3.63 ;
      RECT 42.145 3.278 42.175 3.605 ;
      RECT 42.125 3.276 42.145 3.598 ;
      RECT 42.041 3.274 42.09 3.596 ;
      RECT 41.955 3.271 42.041 3.597 ;
      RECT 41.88 3.27 41.955 3.599 ;
      RECT 41.795 3.27 41.88 3.625 ;
      RECT 41.718 3.271 41.795 3.65 ;
      RECT 41.632 3.272 41.718 3.65 ;
      RECT 41.546 3.272 41.632 3.65 ;
      RECT 41.46 3.273 41.546 3.65 ;
      RECT 41.44 3.274 41.46 3.642 ;
      RECT 41.425 3.28 41.44 3.627 ;
      RECT 41.39 3.3 41.425 3.607 ;
      RECT 41.38 3.32 41.39 3.589 ;
      RECT 42.35 2.625 42.355 2.895 ;
      RECT 42.345 2.616 42.35 2.9 ;
      RECT 42.335 2.606 42.345 2.912 ;
      RECT 42.33 2.595 42.335 2.923 ;
      RECT 42.31 2.589 42.33 2.941 ;
      RECT 42.265 2.586 42.31 2.99 ;
      RECT 42.25 2.585 42.265 3.035 ;
      RECT 42.245 2.585 42.25 3.048 ;
      RECT 42.235 2.585 42.245 3.06 ;
      RECT 42.23 2.586 42.235 3.075 ;
      RECT 42.21 2.594 42.23 3.08 ;
      RECT 42.18 2.61 42.21 3.08 ;
      RECT 42.17 2.622 42.175 3.08 ;
      RECT 42.135 2.637 42.17 3.08 ;
      RECT 42.105 2.657 42.135 3.08 ;
      RECT 42.095 2.682 42.105 3.08 ;
      RECT 42.09 2.71 42.095 3.08 ;
      RECT 42.085 2.74 42.09 3.08 ;
      RECT 42.08 2.757 42.085 3.08 ;
      RECT 42.07 2.785 42.08 3.08 ;
      RECT 42.06 2.82 42.07 3.08 ;
      RECT 42.055 2.855 42.06 3.08 ;
      RECT 42.175 2.62 42.18 3.08 ;
      RECT 41.69 2.722 41.875 2.895 ;
      RECT 41.65 2.64 41.835 2.893 ;
      RECT 41.611 2.645 41.835 2.889 ;
      RECT 41.525 2.654 41.835 2.884 ;
      RECT 41.441 2.67 41.84 2.879 ;
      RECT 41.355 2.69 41.865 2.873 ;
      RECT 41.355 2.71 41.87 2.873 ;
      RECT 41.441 2.68 41.865 2.879 ;
      RECT 41.525 2.655 41.84 2.884 ;
      RECT 41.69 2.637 41.835 2.895 ;
      RECT 41.69 2.632 41.79 2.895 ;
      RECT 41.776 2.626 41.79 2.895 ;
      RECT 41.165 1.95 41.17 2.349 ;
      RECT 40.91 1.95 40.945 2.347 ;
      RECT 40.505 1.985 40.51 2.341 ;
      RECT 41.25 1.988 41.255 2.243 ;
      RECT 41.245 1.986 41.25 2.249 ;
      RECT 41.24 1.985 41.245 2.256 ;
      RECT 41.215 1.978 41.24 2.28 ;
      RECT 41.21 1.971 41.215 2.304 ;
      RECT 41.205 1.967 41.21 2.313 ;
      RECT 41.195 1.962 41.205 2.326 ;
      RECT 41.19 1.959 41.195 2.335 ;
      RECT 41.185 1.957 41.19 2.34 ;
      RECT 41.17 1.953 41.185 2.35 ;
      RECT 41.155 1.947 41.165 2.349 ;
      RECT 41.117 1.945 41.155 2.349 ;
      RECT 41.031 1.947 41.117 2.349 ;
      RECT 40.945 1.949 41.031 2.348 ;
      RECT 40.874 1.95 40.91 2.347 ;
      RECT 40.788 1.952 40.874 2.347 ;
      RECT 40.702 1.954 40.788 2.346 ;
      RECT 40.616 1.956 40.702 2.346 ;
      RECT 40.53 1.959 40.616 2.345 ;
      RECT 40.52 1.965 40.53 2.344 ;
      RECT 40.51 1.977 40.52 2.342 ;
      RECT 40.45 2.012 40.505 2.338 ;
      RECT 40.445 2.042 40.45 2.1 ;
      RECT 41.19 3.122 41.205 3.315 ;
      RECT 41.185 3.09 41.19 3.315 ;
      RECT 41.175 3.065 41.185 3.315 ;
      RECT 41.17 3.037 41.175 3.315 ;
      RECT 41.14 2.96 41.17 3.315 ;
      RECT 41.115 2.842 41.14 3.315 ;
      RECT 41.11 2.78 41.115 3.315 ;
      RECT 41.1 2.767 41.11 3.315 ;
      RECT 41.08 2.757 41.1 3.315 ;
      RECT 41.065 2.74 41.08 3.315 ;
      RECT 41.035 2.728 41.065 3.315 ;
      RECT 41.03 2.727 41.035 3.26 ;
      RECT 41.025 2.727 41.03 3.218 ;
      RECT 41.01 2.726 41.025 3.17 ;
      RECT 40.995 2.726 41.01 3.108 ;
      RECT 40.975 2.726 40.995 3.068 ;
      RECT 40.97 2.726 40.975 3.053 ;
      RECT 40.945 2.725 40.97 3.048 ;
      RECT 40.875 2.724 40.945 3.035 ;
      RECT 40.86 2.723 40.875 3.02 ;
      RECT 40.83 2.722 40.86 3.003 ;
      RECT 40.825 2.722 40.83 2.988 ;
      RECT 40.775 2.721 40.825 2.968 ;
      RECT 40.71 2.72 40.775 2.923 ;
      RECT 40.705 2.72 40.71 2.895 ;
      RECT 40.79 3.257 40.795 3.514 ;
      RECT 40.77 3.176 40.79 3.531 ;
      RECT 40.75 3.17 40.77 3.56 ;
      RECT 40.69 3.157 40.75 3.58 ;
      RECT 40.645 3.141 40.69 3.581 ;
      RECT 40.561 3.129 40.645 3.569 ;
      RECT 40.475 3.116 40.561 3.553 ;
      RECT 40.465 3.109 40.475 3.545 ;
      RECT 40.42 3.106 40.465 3.485 ;
      RECT 40.4 3.102 40.42 3.4 ;
      RECT 40.385 3.1 40.4 3.353 ;
      RECT 40.355 3.097 40.385 3.323 ;
      RECT 40.32 3.093 40.355 3.3 ;
      RECT 40.277 3.088 40.32 3.288 ;
      RECT 40.191 3.079 40.277 3.297 ;
      RECT 40.105 3.068 40.191 3.309 ;
      RECT 40.04 3.059 40.105 3.318 ;
      RECT 40.02 3.05 40.04 3.323 ;
      RECT 40.015 3.043 40.02 3.325 ;
      RECT 39.975 3.028 40.015 3.322 ;
      RECT 39.955 3.007 39.975 3.317 ;
      RECT 39.94 2.995 39.955 3.31 ;
      RECT 39.935 2.987 39.94 3.303 ;
      RECT 39.92 2.967 39.935 3.296 ;
      RECT 39.915 2.83 39.92 3.29 ;
      RECT 39.835 2.719 39.915 3.262 ;
      RECT 39.826 2.712 39.835 3.228 ;
      RECT 39.74 2.706 39.826 3.153 ;
      RECT 39.715 2.697 39.74 3.065 ;
      RECT 39.685 2.692 39.715 3.04 ;
      RECT 39.62 2.701 39.685 3.025 ;
      RECT 39.6 2.717 39.62 3 ;
      RECT 39.59 2.723 39.6 2.948 ;
      RECT 39.57 2.745 39.59 2.83 ;
      RECT 40.225 2.71 40.395 2.895 ;
      RECT 40.225 2.71 40.43 2.893 ;
      RECT 40.275 2.62 40.445 2.884 ;
      RECT 40.225 2.777 40.45 2.877 ;
      RECT 40.24 2.655 40.445 2.884 ;
      RECT 39.44 3.388 39.505 3.831 ;
      RECT 39.38 3.413 39.505 3.829 ;
      RECT 39.38 3.413 39.56 3.823 ;
      RECT 39.365 3.438 39.56 3.822 ;
      RECT 39.505 3.375 39.58 3.819 ;
      RECT 39.44 3.4 39.66 3.813 ;
      RECT 39.365 3.439 39.705 3.807 ;
      RECT 39.35 3.466 39.705 3.798 ;
      RECT 39.365 3.459 39.725 3.79 ;
      RECT 39.35 3.468 39.73 3.773 ;
      RECT 39.345 3.485 39.73 3.6 ;
      RECT 39.35 2.207 39.385 2.445 ;
      RECT 39.35 2.207 39.415 2.444 ;
      RECT 39.35 2.207 39.53 2.44 ;
      RECT 39.35 2.207 39.585 2.418 ;
      RECT 39.36 2.15 39.64 2.318 ;
      RECT 39.465 1.99 39.495 2.441 ;
      RECT 39.495 1.985 39.675 2.198 ;
      RECT 39.365 2.126 39.675 2.198 ;
      RECT 39.415 2.022 39.465 2.442 ;
      RECT 39.385 2.078 39.675 2.198 ;
      RECT 38.255 5.02 38.425 6.49 ;
      RECT 38.255 6.315 38.43 6.485 ;
      RECT 37.885 1.74 38.055 2.93 ;
      RECT 37.885 1.74 38.355 1.91 ;
      RECT 37.885 6.97 38.355 7.14 ;
      RECT 37.885 5.95 38.055 7.14 ;
      RECT 36.895 1.74 37.065 2.93 ;
      RECT 36.895 1.74 37.365 1.91 ;
      RECT 36.895 6.97 37.365 7.14 ;
      RECT 36.895 5.95 37.065 7.14 ;
      RECT 35.045 2.635 35.215 3.865 ;
      RECT 35.1 0.855 35.27 2.805 ;
      RECT 35.045 0.575 35.215 1.025 ;
      RECT 35.045 7.855 35.215 8.305 ;
      RECT 35.1 6.075 35.27 8.025 ;
      RECT 35.045 5.015 35.215 6.245 ;
      RECT 34.525 0.575 34.695 3.865 ;
      RECT 34.525 2.075 34.93 2.405 ;
      RECT 34.525 1.235 34.93 1.565 ;
      RECT 34.525 5.015 34.695 8.305 ;
      RECT 34.525 7.315 34.93 7.645 ;
      RECT 34.525 6.475 34.93 6.805 ;
      RECT 32.625 3.392 32.64 3.443 ;
      RECT 32.62 3.372 32.625 3.49 ;
      RECT 32.605 3.362 32.62 3.558 ;
      RECT 32.58 3.342 32.605 3.613 ;
      RECT 32.54 3.327 32.58 3.633 ;
      RECT 32.495 3.321 32.54 3.661 ;
      RECT 32.425 3.311 32.495 3.678 ;
      RECT 32.405 3.303 32.425 3.678 ;
      RECT 32.345 3.297 32.405 3.67 ;
      RECT 32.286 3.288 32.345 3.658 ;
      RECT 32.2 3.277 32.286 3.641 ;
      RECT 32.178 3.268 32.2 3.629 ;
      RECT 32.092 3.261 32.178 3.616 ;
      RECT 32.006 3.248 32.092 3.597 ;
      RECT 31.92 3.236 32.006 3.577 ;
      RECT 31.89 3.225 31.92 3.564 ;
      RECT 31.84 3.211 31.89 3.556 ;
      RECT 31.82 3.2 31.84 3.548 ;
      RECT 31.771 3.189 31.82 3.54 ;
      RECT 31.685 3.168 31.771 3.525 ;
      RECT 31.64 3.155 31.685 3.51 ;
      RECT 31.595 3.155 31.64 3.49 ;
      RECT 31.54 3.155 31.595 3.425 ;
      RECT 31.515 3.155 31.54 3.348 ;
      RECT 32.04 2.892 32.21 3.075 ;
      RECT 32.04 2.892 32.225 3.033 ;
      RECT 32.04 2.892 32.23 2.975 ;
      RECT 32.1 2.66 32.235 2.951 ;
      RECT 32.1 2.664 32.24 2.934 ;
      RECT 32.045 2.827 32.24 2.934 ;
      RECT 32.07 2.672 32.21 3.075 ;
      RECT 32.07 2.676 32.25 2.875 ;
      RECT 32.055 2.762 32.25 2.875 ;
      RECT 32.065 2.692 32.21 3.075 ;
      RECT 32.065 2.695 32.26 2.788 ;
      RECT 32.06 2.712 32.26 2.788 ;
      RECT 31.83 1.932 32 2.415 ;
      RECT 31.825 1.927 31.975 2.405 ;
      RECT 31.825 1.934 32.005 2.399 ;
      RECT 31.815 1.928 31.975 2.378 ;
      RECT 31.815 1.944 32.02 2.337 ;
      RECT 31.785 1.929 31.975 2.3 ;
      RECT 31.785 1.959 32.03 2.24 ;
      RECT 31.78 1.931 31.975 2.238 ;
      RECT 31.76 1.94 32.005 2.195 ;
      RECT 31.735 1.956 32.02 2.107 ;
      RECT 31.735 1.975 32.045 2.098 ;
      RECT 31.73 2.012 32.045 2.05 ;
      RECT 31.735 1.992 32.05 2.018 ;
      RECT 31.83 1.926 31.94 2.415 ;
      RECT 31.916 1.925 31.94 2.415 ;
      RECT 31.15 2.71 31.155 2.921 ;
      RECT 31.75 2.71 31.755 2.895 ;
      RECT 31.815 2.75 31.82 2.863 ;
      RECT 31.81 2.742 31.815 2.869 ;
      RECT 31.805 2.732 31.81 2.877 ;
      RECT 31.8 2.722 31.805 2.886 ;
      RECT 31.795 2.712 31.8 2.89 ;
      RECT 31.755 2.71 31.795 2.893 ;
      RECT 31.727 2.709 31.75 2.897 ;
      RECT 31.641 2.706 31.727 2.904 ;
      RECT 31.555 2.702 31.641 2.915 ;
      RECT 31.535 2.7 31.555 2.921 ;
      RECT 31.517 2.699 31.535 2.924 ;
      RECT 31.431 2.697 31.517 2.931 ;
      RECT 31.345 2.692 31.431 2.944 ;
      RECT 31.326 2.689 31.345 2.949 ;
      RECT 31.24 2.687 31.326 2.94 ;
      RECT 31.23 2.687 31.24 2.933 ;
      RECT 31.155 2.7 31.23 2.927 ;
      RECT 31.14 2.711 31.15 2.921 ;
      RECT 31.13 2.713 31.14 2.92 ;
      RECT 31.12 2.717 31.13 2.916 ;
      RECT 31.115 2.72 31.12 2.91 ;
      RECT 31.105 2.722 31.115 2.904 ;
      RECT 31.1 2.725 31.105 2.898 ;
      RECT 31.08 3.311 31.085 3.515 ;
      RECT 31.065 3.298 31.08 3.608 ;
      RECT 31.05 3.279 31.065 3.885 ;
      RECT 31.015 3.245 31.05 3.885 ;
      RECT 31.011 3.215 31.015 3.885 ;
      RECT 30.925 3.097 31.011 3.885 ;
      RECT 30.915 2.972 30.925 3.885 ;
      RECT 30.9 2.94 30.915 3.885 ;
      RECT 30.895 2.915 30.9 3.885 ;
      RECT 30.89 2.905 30.895 3.841 ;
      RECT 30.875 2.877 30.89 3.746 ;
      RECT 30.86 2.843 30.875 3.645 ;
      RECT 30.855 2.821 30.86 3.598 ;
      RECT 30.85 2.81 30.855 3.568 ;
      RECT 30.845 2.8 30.85 3.534 ;
      RECT 30.835 2.787 30.845 3.502 ;
      RECT 30.81 2.763 30.835 3.428 ;
      RECT 30.805 2.743 30.81 3.353 ;
      RECT 30.8 2.737 30.805 3.328 ;
      RECT 30.795 2.732 30.8 3.293 ;
      RECT 30.79 2.727 30.795 3.268 ;
      RECT 30.785 2.725 30.79 3.248 ;
      RECT 30.78 2.725 30.785 3.233 ;
      RECT 30.775 2.725 30.78 3.193 ;
      RECT 30.765 2.725 30.775 3.165 ;
      RECT 30.755 2.725 30.765 3.11 ;
      RECT 30.74 2.725 30.755 3.048 ;
      RECT 30.735 2.724 30.74 2.993 ;
      RECT 30.72 2.723 30.735 2.973 ;
      RECT 30.66 2.721 30.72 2.947 ;
      RECT 30.625 2.722 30.66 2.927 ;
      RECT 30.62 2.724 30.625 2.917 ;
      RECT 30.61 2.743 30.62 2.907 ;
      RECT 30.605 2.77 30.61 2.838 ;
      RECT 30.72 2.195 30.89 2.44 ;
      RECT 30.755 1.966 30.89 2.44 ;
      RECT 30.755 1.968 30.9 2.435 ;
      RECT 30.755 1.97 30.925 2.423 ;
      RECT 30.755 1.973 30.95 2.405 ;
      RECT 30.755 1.978 31 2.378 ;
      RECT 30.755 1.983 31.02 2.343 ;
      RECT 30.735 1.985 31.03 2.318 ;
      RECT 30.725 2.08 31.03 2.318 ;
      RECT 30.755 1.965 30.865 2.44 ;
      RECT 30.765 1.962 30.86 2.44 ;
      RECT 30.285 3.227 30.475 3.585 ;
      RECT 30.285 3.239 30.51 3.584 ;
      RECT 30.285 3.267 30.53 3.582 ;
      RECT 30.285 3.292 30.535 3.581 ;
      RECT 30.285 3.35 30.55 3.58 ;
      RECT 30.27 3.223 30.43 3.565 ;
      RECT 30.25 3.232 30.475 3.518 ;
      RECT 30.225 3.243 30.51 3.455 ;
      RECT 30.225 3.327 30.545 3.455 ;
      RECT 30.225 3.302 30.54 3.455 ;
      RECT 30.285 3.218 30.43 3.585 ;
      RECT 30.371 3.217 30.43 3.585 ;
      RECT 30.371 3.216 30.415 3.585 ;
      RECT 30.285 7.855 30.455 8.305 ;
      RECT 30.34 6.075 30.51 8.025 ;
      RECT 30.285 5.015 30.455 6.245 ;
      RECT 29.765 5.015 29.935 8.305 ;
      RECT 29.765 7.315 30.17 7.645 ;
      RECT 29.765 6.475 30.17 6.805 ;
      RECT 30.07 2.732 30.075 3.11 ;
      RECT 30.065 2.7 30.07 3.11 ;
      RECT 30.06 2.672 30.065 3.11 ;
      RECT 30.055 2.652 30.06 3.11 ;
      RECT 30 2.635 30.055 3.11 ;
      RECT 29.96 2.62 30 3.11 ;
      RECT 29.905 2.607 29.96 3.11 ;
      RECT 29.87 2.598 29.905 3.11 ;
      RECT 29.866 2.596 29.87 3.109 ;
      RECT 29.78 2.592 29.866 3.092 ;
      RECT 29.695 2.584 29.78 3.055 ;
      RECT 29.685 2.58 29.695 3.028 ;
      RECT 29.675 2.58 29.685 3.01 ;
      RECT 29.665 2.582 29.675 2.993 ;
      RECT 29.66 2.587 29.665 2.979 ;
      RECT 29.655 2.591 29.66 2.966 ;
      RECT 29.645 2.596 29.655 2.95 ;
      RECT 29.63 2.61 29.645 2.925 ;
      RECT 29.625 2.616 29.63 2.905 ;
      RECT 29.62 2.618 29.625 2.898 ;
      RECT 29.615 2.622 29.62 2.773 ;
      RECT 29.795 3.422 30.04 3.885 ;
      RECT 29.715 3.395 30.035 3.881 ;
      RECT 29.645 3.43 30.04 3.874 ;
      RECT 29.435 3.685 30.04 3.87 ;
      RECT 29.615 3.453 30.04 3.87 ;
      RECT 29.455 3.645 30.04 3.87 ;
      RECT 29.605 3.465 30.04 3.87 ;
      RECT 29.49 3.582 30.04 3.87 ;
      RECT 29.545 3.507 30.04 3.87 ;
      RECT 29.795 3.372 30.035 3.885 ;
      RECT 29.825 3.365 30.035 3.885 ;
      RECT 29.815 3.367 30.035 3.885 ;
      RECT 29.825 3.362 29.955 3.885 ;
      RECT 29.38 1.925 29.466 2.364 ;
      RECT 29.375 1.925 29.466 2.362 ;
      RECT 29.375 1.925 29.535 2.361 ;
      RECT 29.375 1.925 29.565 2.358 ;
      RECT 29.36 1.932 29.565 2.349 ;
      RECT 29.36 1.932 29.57 2.345 ;
      RECT 29.355 1.942 29.57 2.338 ;
      RECT 29.35 1.947 29.57 2.313 ;
      RECT 29.35 1.947 29.585 2.295 ;
      RECT 29.375 1.925 29.605 2.21 ;
      RECT 29.345 1.952 29.605 2.208 ;
      RECT 29.355 1.945 29.61 2.146 ;
      RECT 29.345 2.067 29.615 2.129 ;
      RECT 29.33 1.962 29.61 2.08 ;
      RECT 29.325 1.972 29.61 1.98 ;
      RECT 29.405 2.743 29.41 2.82 ;
      RECT 29.395 2.737 29.405 3.01 ;
      RECT 29.385 2.729 29.395 3.031 ;
      RECT 29.375 2.72 29.385 3.053 ;
      RECT 29.37 2.715 29.375 3.07 ;
      RECT 29.33 2.715 29.37 3.11 ;
      RECT 29.31 2.715 29.33 3.165 ;
      RECT 29.305 2.715 29.31 3.193 ;
      RECT 29.295 2.715 29.305 3.208 ;
      RECT 29.26 2.715 29.295 3.25 ;
      RECT 29.255 2.715 29.26 3.293 ;
      RECT 29.245 2.715 29.255 3.308 ;
      RECT 29.23 2.715 29.245 3.328 ;
      RECT 29.215 2.715 29.23 3.355 ;
      RECT 29.21 2.716 29.215 3.373 ;
      RECT 29.19 2.717 29.21 3.38 ;
      RECT 29.135 2.718 29.19 3.4 ;
      RECT 29.125 2.719 29.135 3.414 ;
      RECT 29.12 2.722 29.125 3.413 ;
      RECT 29.08 2.795 29.12 3.411 ;
      RECT 29.065 2.875 29.08 3.409 ;
      RECT 29.04 2.93 29.065 3.407 ;
      RECT 29.025 2.995 29.04 3.406 ;
      RECT 28.98 3.027 29.025 3.403 ;
      RECT 28.895 3.05 28.98 3.398 ;
      RECT 28.87 3.07 28.895 3.393 ;
      RECT 28.8 3.075 28.87 3.389 ;
      RECT 28.78 3.077 28.8 3.386 ;
      RECT 28.695 3.088 28.78 3.38 ;
      RECT 28.69 3.099 28.695 3.375 ;
      RECT 28.68 3.101 28.69 3.375 ;
      RECT 28.645 3.105 28.68 3.373 ;
      RECT 28.595 3.115 28.645 3.36 ;
      RECT 28.575 3.123 28.595 3.345 ;
      RECT 28.495 3.135 28.575 3.328 ;
      RECT 28.66 2.685 28.83 2.895 ;
      RECT 28.776 2.681 28.83 2.895 ;
      RECT 28.581 2.685 28.83 2.886 ;
      RECT 28.581 2.685 28.835 2.875 ;
      RECT 28.495 2.685 28.835 2.866 ;
      RECT 28.495 2.693 28.845 2.81 ;
      RECT 28.495 2.705 28.85 2.723 ;
      RECT 28.495 2.712 28.855 2.715 ;
      RECT 28.69 2.683 28.83 2.895 ;
      RECT 28.445 3.628 28.69 3.96 ;
      RECT 28.44 3.62 28.445 3.957 ;
      RECT 28.41 3.64 28.69 3.938 ;
      RECT 28.39 3.672 28.69 3.911 ;
      RECT 28.44 3.625 28.617 3.957 ;
      RECT 28.44 3.622 28.531 3.957 ;
      RECT 28.38 1.97 28.55 2.39 ;
      RECT 28.375 1.97 28.55 2.388 ;
      RECT 28.375 1.97 28.575 2.378 ;
      RECT 28.375 1.97 28.595 2.353 ;
      RECT 28.37 1.97 28.595 2.348 ;
      RECT 28.37 1.97 28.605 2.338 ;
      RECT 28.37 1.97 28.61 2.333 ;
      RECT 28.37 1.975 28.615 2.328 ;
      RECT 28.37 2.007 28.63 2.318 ;
      RECT 28.37 2.077 28.655 2.301 ;
      RECT 28.35 2.077 28.655 2.293 ;
      RECT 28.35 2.137 28.665 2.27 ;
      RECT 28.35 2.177 28.675 2.215 ;
      RECT 28.335 1.97 28.61 2.195 ;
      RECT 28.325 1.985 28.615 2.093 ;
      RECT 27.915 3.375 28.085 3.9 ;
      RECT 27.91 3.375 28.085 3.893 ;
      RECT 27.9 3.375 28.09 3.858 ;
      RECT 27.895 3.385 28.09 3.83 ;
      RECT 27.89 3.405 28.09 3.813 ;
      RECT 27.9 3.38 28.095 3.803 ;
      RECT 27.885 3.425 28.095 3.795 ;
      RECT 27.88 3.445 28.095 3.78 ;
      RECT 27.875 3.475 28.095 3.77 ;
      RECT 27.865 3.52 28.095 3.745 ;
      RECT 27.895 3.39 28.1 3.728 ;
      RECT 27.86 3.572 28.1 3.723 ;
      RECT 27.895 3.4 28.105 3.693 ;
      RECT 27.855 3.605 28.105 3.69 ;
      RECT 27.85 3.63 28.105 3.67 ;
      RECT 27.89 3.417 28.115 3.61 ;
      RECT 27.885 3.439 28.125 3.503 ;
      RECT 27.835 2.686 27.85 2.955 ;
      RECT 27.79 2.67 27.835 3 ;
      RECT 27.785 2.658 27.79 3.05 ;
      RECT 27.775 2.654 27.785 3.083 ;
      RECT 27.77 2.651 27.775 3.111 ;
      RECT 27.755 2.653 27.77 3.153 ;
      RECT 27.75 2.657 27.755 3.193 ;
      RECT 27.73 2.662 27.75 3.245 ;
      RECT 27.726 2.667 27.73 3.302 ;
      RECT 27.64 2.686 27.726 3.339 ;
      RECT 27.63 2.707 27.64 3.375 ;
      RECT 27.625 2.715 27.63 3.376 ;
      RECT 27.62 2.757 27.625 3.377 ;
      RECT 27.605 2.845 27.62 3.378 ;
      RECT 27.595 2.995 27.605 3.38 ;
      RECT 27.59 3.04 27.595 3.382 ;
      RECT 27.555 3.082 27.59 3.385 ;
      RECT 27.55 3.1 27.555 3.388 ;
      RECT 27.473 3.106 27.55 3.394 ;
      RECT 27.387 3.12 27.473 3.407 ;
      RECT 27.301 3.134 27.387 3.421 ;
      RECT 27.215 3.148 27.301 3.434 ;
      RECT 27.155 3.16 27.215 3.446 ;
      RECT 27.13 3.167 27.155 3.453 ;
      RECT 27.116 3.17 27.13 3.458 ;
      RECT 27.03 3.178 27.116 3.474 ;
      RECT 27.025 3.185 27.03 3.489 ;
      RECT 27.001 3.185 27.025 3.496 ;
      RECT 26.915 3.188 27.001 3.524 ;
      RECT 26.83 3.192 26.915 3.568 ;
      RECT 26.765 3.196 26.83 3.605 ;
      RECT 26.74 3.199 26.765 3.621 ;
      RECT 26.665 3.212 26.74 3.625 ;
      RECT 26.64 3.23 26.665 3.629 ;
      RECT 26.63 3.237 26.64 3.631 ;
      RECT 26.615 3.24 26.63 3.632 ;
      RECT 26.555 3.252 26.615 3.636 ;
      RECT 26.545 3.266 26.555 3.64 ;
      RECT 26.49 3.276 26.545 3.628 ;
      RECT 26.465 3.297 26.49 3.611 ;
      RECT 26.445 3.317 26.465 3.602 ;
      RECT 26.44 3.33 26.445 3.597 ;
      RECT 26.425 3.342 26.44 3.593 ;
      RECT 27.66 1.997 27.665 2.02 ;
      RECT 27.655 1.988 27.66 2.06 ;
      RECT 27.65 1.986 27.655 2.103 ;
      RECT 27.645 1.977 27.65 2.138 ;
      RECT 27.64 1.967 27.645 2.21 ;
      RECT 27.635 1.957 27.64 2.275 ;
      RECT 27.63 1.954 27.635 2.315 ;
      RECT 27.605 1.948 27.63 2.405 ;
      RECT 27.57 1.936 27.605 2.43 ;
      RECT 27.56 1.927 27.57 2.43 ;
      RECT 27.425 1.925 27.435 2.413 ;
      RECT 27.415 1.925 27.425 2.38 ;
      RECT 27.41 1.925 27.415 2.355 ;
      RECT 27.405 1.925 27.41 2.343 ;
      RECT 27.4 1.925 27.405 2.325 ;
      RECT 27.39 1.925 27.4 2.29 ;
      RECT 27.385 1.927 27.39 2.268 ;
      RECT 27.38 1.933 27.385 2.253 ;
      RECT 27.375 1.939 27.38 2.238 ;
      RECT 27.36 1.951 27.375 2.211 ;
      RECT 27.355 1.962 27.36 2.179 ;
      RECT 27.35 1.972 27.355 2.163 ;
      RECT 27.34 1.98 27.35 2.132 ;
      RECT 27.335 1.99 27.34 2.106 ;
      RECT 27.33 2.047 27.335 2.089 ;
      RECT 27.435 1.925 27.56 2.43 ;
      RECT 27.15 2.612 27.41 2.91 ;
      RECT 27.145 2.619 27.41 2.908 ;
      RECT 27.15 2.614 27.425 2.903 ;
      RECT 27.14 2.627 27.425 2.9 ;
      RECT 27.14 2.632 27.43 2.893 ;
      RECT 27.135 2.64 27.43 2.89 ;
      RECT 27.135 2.657 27.435 2.688 ;
      RECT 27.15 2.609 27.381 2.91 ;
      RECT 27.205 2.608 27.381 2.91 ;
      RECT 27.205 2.605 27.295 2.91 ;
      RECT 27.205 2.602 27.291 2.91 ;
      RECT 26.895 2.875 26.9 2.888 ;
      RECT 26.89 2.842 26.895 2.893 ;
      RECT 26.885 2.797 26.89 2.9 ;
      RECT 26.88 2.752 26.885 2.908 ;
      RECT 26.875 2.72 26.88 2.916 ;
      RECT 26.87 2.68 26.875 2.917 ;
      RECT 26.855 2.66 26.87 2.919 ;
      RECT 26.78 2.642 26.855 2.931 ;
      RECT 26.77 2.635 26.78 2.942 ;
      RECT 26.765 2.635 26.77 2.944 ;
      RECT 26.735 2.641 26.765 2.948 ;
      RECT 26.695 2.654 26.735 2.948 ;
      RECT 26.67 2.665 26.695 2.934 ;
      RECT 26.655 2.671 26.67 2.917 ;
      RECT 26.645 2.673 26.655 2.908 ;
      RECT 26.64 2.674 26.645 2.903 ;
      RECT 26.635 2.675 26.64 2.898 ;
      RECT 26.63 2.676 26.635 2.895 ;
      RECT 26.605 2.681 26.63 2.885 ;
      RECT 26.595 2.697 26.605 2.872 ;
      RECT 26.59 2.717 26.595 2.867 ;
      RECT 26.6 2.11 26.605 2.306 ;
      RECT 26.585 2.074 26.6 2.308 ;
      RECT 26.575 2.056 26.585 2.313 ;
      RECT 26.565 2.042 26.575 2.317 ;
      RECT 26.52 2.026 26.565 2.327 ;
      RECT 26.515 2.016 26.52 2.336 ;
      RECT 26.47 2.005 26.515 2.342 ;
      RECT 26.465 1.993 26.47 2.349 ;
      RECT 26.45 1.988 26.465 2.353 ;
      RECT 26.435 1.98 26.45 2.358 ;
      RECT 26.425 1.973 26.435 2.363 ;
      RECT 26.415 1.97 26.425 2.368 ;
      RECT 26.405 1.97 26.415 2.369 ;
      RECT 26.4 1.967 26.405 2.368 ;
      RECT 26.365 1.962 26.39 2.367 ;
      RECT 26.341 1.958 26.365 2.366 ;
      RECT 26.255 1.949 26.341 2.363 ;
      RECT 26.24 1.941 26.255 2.36 ;
      RECT 26.218 1.94 26.24 2.359 ;
      RECT 26.132 1.94 26.218 2.357 ;
      RECT 26.046 1.94 26.132 2.355 ;
      RECT 25.96 1.94 26.046 2.352 ;
      RECT 25.95 1.94 25.96 2.343 ;
      RECT 25.92 1.94 25.95 2.303 ;
      RECT 25.91 1.95 25.92 2.258 ;
      RECT 25.905 1.99 25.91 2.243 ;
      RECT 25.9 2.005 25.905 2.23 ;
      RECT 25.87 2.085 25.9 2.192 ;
      RECT 26.39 1.965 26.4 2.368 ;
      RECT 26.215 2.73 26.23 3.335 ;
      RECT 26.22 2.725 26.23 3.335 ;
      RECT 26.385 2.725 26.39 2.908 ;
      RECT 26.375 2.725 26.385 2.938 ;
      RECT 26.36 2.725 26.375 2.998 ;
      RECT 26.355 2.725 26.36 3.043 ;
      RECT 26.35 2.725 26.355 3.073 ;
      RECT 26.345 2.725 26.35 3.093 ;
      RECT 26.335 2.725 26.345 3.128 ;
      RECT 26.32 2.725 26.335 3.16 ;
      RECT 26.275 2.725 26.32 3.188 ;
      RECT 26.27 2.725 26.275 3.218 ;
      RECT 26.265 2.725 26.27 3.23 ;
      RECT 26.26 2.725 26.265 3.238 ;
      RECT 26.25 2.725 26.26 3.253 ;
      RECT 26.245 2.725 26.25 3.275 ;
      RECT 26.235 2.725 26.245 3.298 ;
      RECT 26.23 2.725 26.235 3.318 ;
      RECT 26.195 2.74 26.215 3.335 ;
      RECT 26.17 2.757 26.195 3.335 ;
      RECT 26.165 2.767 26.17 3.335 ;
      RECT 26.135 2.782 26.165 3.335 ;
      RECT 26.06 2.824 26.135 3.335 ;
      RECT 26.055 2.855 26.06 3.318 ;
      RECT 26.05 2.859 26.055 3.3 ;
      RECT 26.045 2.863 26.05 3.263 ;
      RECT 26.04 3.047 26.045 3.23 ;
      RECT 25.525 3.236 25.611 3.801 ;
      RECT 25.48 3.238 25.645 3.795 ;
      RECT 25.611 3.235 25.645 3.795 ;
      RECT 25.525 3.237 25.73 3.789 ;
      RECT 25.48 3.247 25.74 3.785 ;
      RECT 25.455 3.239 25.73 3.781 ;
      RECT 25.45 3.242 25.73 3.776 ;
      RECT 25.425 3.257 25.74 3.77 ;
      RECT 25.425 3.282 25.78 3.765 ;
      RECT 25.385 3.29 25.78 3.74 ;
      RECT 25.385 3.317 25.795 3.738 ;
      RECT 25.385 3.347 25.805 3.725 ;
      RECT 25.38 3.492 25.805 3.713 ;
      RECT 25.385 3.421 25.825 3.71 ;
      RECT 25.385 3.478 25.83 3.518 ;
      RECT 25.575 2.757 25.745 2.935 ;
      RECT 25.525 2.696 25.575 2.92 ;
      RECT 25.26 2.676 25.525 2.905 ;
      RECT 25.22 2.74 25.695 2.905 ;
      RECT 25.22 2.73 25.65 2.905 ;
      RECT 25.22 2.727 25.64 2.905 ;
      RECT 25.22 2.715 25.63 2.905 ;
      RECT 25.22 2.7 25.575 2.905 ;
      RECT 25.26 2.672 25.461 2.905 ;
      RECT 25.27 2.65 25.461 2.905 ;
      RECT 25.295 2.635 25.375 2.905 ;
      RECT 25.05 3.165 25.17 3.61 ;
      RECT 25.035 3.165 25.17 3.609 ;
      RECT 24.99 3.187 25.17 3.604 ;
      RECT 24.95 3.236 25.17 3.598 ;
      RECT 24.95 3.236 25.175 3.573 ;
      RECT 24.95 3.236 25.195 3.463 ;
      RECT 24.945 3.266 25.195 3.46 ;
      RECT 25.035 3.165 25.205 3.355 ;
      RECT 24.695 1.95 24.7 2.395 ;
      RECT 24.505 1.95 24.525 2.36 ;
      RECT 24.475 1.95 24.48 2.335 ;
      RECT 25.155 2.257 25.17 2.445 ;
      RECT 25.15 2.242 25.155 2.451 ;
      RECT 25.13 2.215 25.15 2.454 ;
      RECT 25.08 2.182 25.13 2.463 ;
      RECT 25.05 2.162 25.08 2.467 ;
      RECT 25.031 2.15 25.05 2.463 ;
      RECT 24.945 2.122 25.031 2.453 ;
      RECT 24.935 2.097 24.945 2.443 ;
      RECT 24.865 2.065 24.935 2.435 ;
      RECT 24.84 2.025 24.865 2.427 ;
      RECT 24.82 2.007 24.84 2.421 ;
      RECT 24.81 1.997 24.82 2.418 ;
      RECT 24.8 1.99 24.81 2.416 ;
      RECT 24.78 1.977 24.8 2.413 ;
      RECT 24.77 1.967 24.78 2.41 ;
      RECT 24.76 1.96 24.77 2.408 ;
      RECT 24.71 1.952 24.76 2.402 ;
      RECT 24.7 1.95 24.71 2.396 ;
      RECT 24.67 1.95 24.695 2.393 ;
      RECT 24.641 1.95 24.67 2.388 ;
      RECT 24.555 1.95 24.641 2.378 ;
      RECT 24.525 1.95 24.555 2.365 ;
      RECT 24.48 1.95 24.505 2.348 ;
      RECT 24.465 1.95 24.475 2.33 ;
      RECT 24.445 1.957 24.465 2.315 ;
      RECT 24.44 1.972 24.445 2.303 ;
      RECT 24.435 1.977 24.44 2.243 ;
      RECT 24.43 1.982 24.435 2.085 ;
      RECT 24.425 1.985 24.43 2.003 ;
      RECT 24.69 2.67 24.776 2.991 ;
      RECT 24.69 2.67 24.81 2.984 ;
      RECT 24.64 2.67 24.81 2.98 ;
      RECT 24.64 2.672 24.896 2.978 ;
      RECT 24.64 2.674 24.92 2.972 ;
      RECT 24.64 2.681 24.93 2.971 ;
      RECT 24.64 2.69 24.935 2.968 ;
      RECT 24.64 2.696 24.94 2.963 ;
      RECT 24.64 2.74 24.945 2.96 ;
      RECT 24.64 2.832 24.95 2.957 ;
      RECT 24.165 3.275 24.2 3.595 ;
      RECT 24.75 3.46 24.755 3.642 ;
      RECT 24.705 3.342 24.75 3.661 ;
      RECT 24.69 3.319 24.705 3.684 ;
      RECT 24.68 3.309 24.69 3.694 ;
      RECT 24.66 3.304 24.68 3.707 ;
      RECT 24.635 3.302 24.66 3.728 ;
      RECT 24.616 3.301 24.635 3.74 ;
      RECT 24.53 3.298 24.616 3.74 ;
      RECT 24.46 3.293 24.53 3.728 ;
      RECT 24.385 3.289 24.46 3.703 ;
      RECT 24.32 3.285 24.385 3.67 ;
      RECT 24.25 3.282 24.32 3.63 ;
      RECT 24.22 3.278 24.25 3.605 ;
      RECT 24.2 3.276 24.22 3.598 ;
      RECT 24.116 3.274 24.165 3.596 ;
      RECT 24.03 3.271 24.116 3.597 ;
      RECT 23.955 3.27 24.03 3.599 ;
      RECT 23.87 3.27 23.955 3.625 ;
      RECT 23.793 3.271 23.87 3.65 ;
      RECT 23.707 3.272 23.793 3.65 ;
      RECT 23.621 3.272 23.707 3.65 ;
      RECT 23.535 3.273 23.621 3.65 ;
      RECT 23.515 3.274 23.535 3.642 ;
      RECT 23.5 3.28 23.515 3.627 ;
      RECT 23.465 3.3 23.5 3.607 ;
      RECT 23.455 3.32 23.465 3.589 ;
      RECT 24.425 2.625 24.43 2.895 ;
      RECT 24.42 2.616 24.425 2.9 ;
      RECT 24.41 2.606 24.42 2.912 ;
      RECT 24.405 2.595 24.41 2.923 ;
      RECT 24.385 2.589 24.405 2.941 ;
      RECT 24.34 2.586 24.385 2.99 ;
      RECT 24.325 2.585 24.34 3.035 ;
      RECT 24.32 2.585 24.325 3.048 ;
      RECT 24.31 2.585 24.32 3.06 ;
      RECT 24.305 2.586 24.31 3.075 ;
      RECT 24.285 2.594 24.305 3.08 ;
      RECT 24.255 2.61 24.285 3.08 ;
      RECT 24.245 2.622 24.25 3.08 ;
      RECT 24.21 2.637 24.245 3.08 ;
      RECT 24.18 2.657 24.21 3.08 ;
      RECT 24.17 2.682 24.18 3.08 ;
      RECT 24.165 2.71 24.17 3.08 ;
      RECT 24.16 2.74 24.165 3.08 ;
      RECT 24.155 2.757 24.16 3.08 ;
      RECT 24.145 2.785 24.155 3.08 ;
      RECT 24.135 2.82 24.145 3.08 ;
      RECT 24.13 2.855 24.135 3.08 ;
      RECT 24.25 2.62 24.255 3.08 ;
      RECT 23.765 2.722 23.95 2.895 ;
      RECT 23.725 2.64 23.91 2.893 ;
      RECT 23.686 2.645 23.91 2.889 ;
      RECT 23.6 2.654 23.91 2.884 ;
      RECT 23.516 2.67 23.915 2.879 ;
      RECT 23.43 2.69 23.94 2.873 ;
      RECT 23.43 2.71 23.945 2.873 ;
      RECT 23.516 2.68 23.94 2.879 ;
      RECT 23.6 2.655 23.915 2.884 ;
      RECT 23.765 2.637 23.91 2.895 ;
      RECT 23.765 2.632 23.865 2.895 ;
      RECT 23.851 2.626 23.865 2.895 ;
      RECT 23.24 1.95 23.245 2.349 ;
      RECT 22.985 1.95 23.02 2.347 ;
      RECT 22.58 1.985 22.585 2.341 ;
      RECT 23.325 1.988 23.33 2.243 ;
      RECT 23.32 1.986 23.325 2.249 ;
      RECT 23.315 1.985 23.32 2.256 ;
      RECT 23.29 1.978 23.315 2.28 ;
      RECT 23.285 1.971 23.29 2.304 ;
      RECT 23.28 1.967 23.285 2.313 ;
      RECT 23.27 1.962 23.28 2.326 ;
      RECT 23.265 1.959 23.27 2.335 ;
      RECT 23.26 1.957 23.265 2.34 ;
      RECT 23.245 1.953 23.26 2.35 ;
      RECT 23.23 1.947 23.24 2.349 ;
      RECT 23.192 1.945 23.23 2.349 ;
      RECT 23.106 1.947 23.192 2.349 ;
      RECT 23.02 1.949 23.106 2.348 ;
      RECT 22.949 1.95 22.985 2.347 ;
      RECT 22.863 1.952 22.949 2.347 ;
      RECT 22.777 1.954 22.863 2.346 ;
      RECT 22.691 1.956 22.777 2.346 ;
      RECT 22.605 1.959 22.691 2.345 ;
      RECT 22.595 1.965 22.605 2.344 ;
      RECT 22.585 1.977 22.595 2.342 ;
      RECT 22.525 2.012 22.58 2.338 ;
      RECT 22.52 2.042 22.525 2.1 ;
      RECT 23.265 3.122 23.28 3.315 ;
      RECT 23.26 3.09 23.265 3.315 ;
      RECT 23.25 3.065 23.26 3.315 ;
      RECT 23.245 3.037 23.25 3.315 ;
      RECT 23.215 2.96 23.245 3.315 ;
      RECT 23.19 2.842 23.215 3.315 ;
      RECT 23.185 2.78 23.19 3.315 ;
      RECT 23.175 2.767 23.185 3.315 ;
      RECT 23.155 2.757 23.175 3.315 ;
      RECT 23.14 2.74 23.155 3.315 ;
      RECT 23.11 2.728 23.14 3.315 ;
      RECT 23.105 2.727 23.11 3.26 ;
      RECT 23.1 2.727 23.105 3.218 ;
      RECT 23.085 2.726 23.1 3.17 ;
      RECT 23.07 2.726 23.085 3.108 ;
      RECT 23.05 2.726 23.07 3.068 ;
      RECT 23.045 2.726 23.05 3.053 ;
      RECT 23.02 2.725 23.045 3.048 ;
      RECT 22.95 2.724 23.02 3.035 ;
      RECT 22.935 2.723 22.95 3.02 ;
      RECT 22.905 2.722 22.935 3.003 ;
      RECT 22.9 2.722 22.905 2.988 ;
      RECT 22.85 2.721 22.9 2.968 ;
      RECT 22.785 2.72 22.85 2.923 ;
      RECT 22.78 2.72 22.785 2.895 ;
      RECT 22.865 3.257 22.87 3.514 ;
      RECT 22.845 3.176 22.865 3.531 ;
      RECT 22.825 3.17 22.845 3.56 ;
      RECT 22.765 3.157 22.825 3.58 ;
      RECT 22.72 3.141 22.765 3.581 ;
      RECT 22.636 3.129 22.72 3.569 ;
      RECT 22.55 3.116 22.636 3.553 ;
      RECT 22.54 3.109 22.55 3.545 ;
      RECT 22.495 3.106 22.54 3.485 ;
      RECT 22.475 3.102 22.495 3.4 ;
      RECT 22.46 3.1 22.475 3.353 ;
      RECT 22.43 3.097 22.46 3.323 ;
      RECT 22.395 3.093 22.43 3.3 ;
      RECT 22.352 3.088 22.395 3.288 ;
      RECT 22.266 3.079 22.352 3.297 ;
      RECT 22.18 3.068 22.266 3.309 ;
      RECT 22.115 3.059 22.18 3.318 ;
      RECT 22.095 3.05 22.115 3.323 ;
      RECT 22.09 3.043 22.095 3.325 ;
      RECT 22.05 3.028 22.09 3.322 ;
      RECT 22.03 3.007 22.05 3.317 ;
      RECT 22.015 2.995 22.03 3.31 ;
      RECT 22.01 2.987 22.015 3.303 ;
      RECT 21.995 2.967 22.01 3.296 ;
      RECT 21.99 2.83 21.995 3.29 ;
      RECT 21.91 2.719 21.99 3.262 ;
      RECT 21.901 2.712 21.91 3.228 ;
      RECT 21.815 2.706 21.901 3.153 ;
      RECT 21.79 2.697 21.815 3.065 ;
      RECT 21.76 2.692 21.79 3.04 ;
      RECT 21.695 2.701 21.76 3.025 ;
      RECT 21.675 2.717 21.695 3 ;
      RECT 21.665 2.723 21.675 2.948 ;
      RECT 21.645 2.745 21.665 2.83 ;
      RECT 22.3 2.71 22.47 2.895 ;
      RECT 22.3 2.71 22.505 2.893 ;
      RECT 22.35 2.62 22.52 2.884 ;
      RECT 22.3 2.777 22.525 2.877 ;
      RECT 22.315 2.655 22.52 2.884 ;
      RECT 21.515 3.388 21.58 3.831 ;
      RECT 21.455 3.413 21.58 3.829 ;
      RECT 21.455 3.413 21.635 3.823 ;
      RECT 21.44 3.438 21.635 3.822 ;
      RECT 21.58 3.375 21.655 3.819 ;
      RECT 21.515 3.4 21.735 3.813 ;
      RECT 21.44 3.439 21.78 3.807 ;
      RECT 21.425 3.466 21.78 3.798 ;
      RECT 21.44 3.459 21.8 3.79 ;
      RECT 21.425 3.468 21.805 3.773 ;
      RECT 21.42 3.485 21.805 3.6 ;
      RECT 21.425 2.207 21.46 2.445 ;
      RECT 21.425 2.207 21.49 2.444 ;
      RECT 21.425 2.207 21.605 2.44 ;
      RECT 21.425 2.207 21.66 2.418 ;
      RECT 21.435 2.15 21.715 2.318 ;
      RECT 21.54 1.99 21.57 2.441 ;
      RECT 21.57 1.985 21.75 2.198 ;
      RECT 21.44 2.126 21.75 2.198 ;
      RECT 21.49 2.022 21.54 2.442 ;
      RECT 21.46 2.078 21.75 2.198 ;
      RECT 20.33 5.02 20.5 6.49 ;
      RECT 20.33 6.315 20.505 6.485 ;
      RECT 19.96 1.74 20.13 2.93 ;
      RECT 19.96 1.74 20.43 1.91 ;
      RECT 19.96 6.97 20.43 7.14 ;
      RECT 19.96 5.95 20.13 7.14 ;
      RECT 18.97 1.74 19.14 2.93 ;
      RECT 18.97 1.74 19.44 1.91 ;
      RECT 18.97 6.97 19.44 7.14 ;
      RECT 18.97 5.95 19.14 7.14 ;
      RECT 17.12 2.635 17.29 3.865 ;
      RECT 17.175 0.855 17.345 2.805 ;
      RECT 17.12 0.575 17.29 1.025 ;
      RECT 17.12 7.855 17.29 8.305 ;
      RECT 17.175 6.075 17.345 8.025 ;
      RECT 17.12 5.015 17.29 6.245 ;
      RECT 16.6 0.575 16.77 3.865 ;
      RECT 16.6 2.075 17.005 2.405 ;
      RECT 16.6 1.235 17.005 1.565 ;
      RECT 16.6 5.015 16.77 8.305 ;
      RECT 16.6 7.315 17.005 7.645 ;
      RECT 16.6 6.475 17.005 6.805 ;
      RECT 14.7 3.392 14.715 3.443 ;
      RECT 14.695 3.372 14.7 3.49 ;
      RECT 14.68 3.362 14.695 3.558 ;
      RECT 14.655 3.342 14.68 3.613 ;
      RECT 14.615 3.327 14.655 3.633 ;
      RECT 14.57 3.321 14.615 3.661 ;
      RECT 14.5 3.311 14.57 3.678 ;
      RECT 14.48 3.303 14.5 3.678 ;
      RECT 14.42 3.297 14.48 3.67 ;
      RECT 14.361 3.288 14.42 3.658 ;
      RECT 14.275 3.277 14.361 3.641 ;
      RECT 14.253 3.268 14.275 3.629 ;
      RECT 14.167 3.261 14.253 3.616 ;
      RECT 14.081 3.248 14.167 3.597 ;
      RECT 13.995 3.236 14.081 3.577 ;
      RECT 13.965 3.225 13.995 3.564 ;
      RECT 13.915 3.211 13.965 3.556 ;
      RECT 13.895 3.2 13.915 3.548 ;
      RECT 13.846 3.189 13.895 3.54 ;
      RECT 13.76 3.168 13.846 3.525 ;
      RECT 13.715 3.155 13.76 3.51 ;
      RECT 13.67 3.155 13.715 3.49 ;
      RECT 13.615 3.155 13.67 3.425 ;
      RECT 13.59 3.155 13.615 3.348 ;
      RECT 14.115 2.892 14.285 3.075 ;
      RECT 14.115 2.892 14.3 3.033 ;
      RECT 14.115 2.892 14.305 2.975 ;
      RECT 14.175 2.66 14.31 2.951 ;
      RECT 14.175 2.664 14.315 2.934 ;
      RECT 14.12 2.827 14.315 2.934 ;
      RECT 14.145 2.672 14.285 3.075 ;
      RECT 14.145 2.676 14.325 2.875 ;
      RECT 14.13 2.762 14.325 2.875 ;
      RECT 14.14 2.692 14.285 3.075 ;
      RECT 14.14 2.695 14.335 2.788 ;
      RECT 14.135 2.712 14.335 2.788 ;
      RECT 13.905 1.932 14.075 2.415 ;
      RECT 13.9 1.927 14.05 2.405 ;
      RECT 13.9 1.934 14.08 2.399 ;
      RECT 13.89 1.928 14.05 2.378 ;
      RECT 13.89 1.944 14.095 2.337 ;
      RECT 13.86 1.929 14.05 2.3 ;
      RECT 13.86 1.959 14.105 2.24 ;
      RECT 13.855 1.931 14.05 2.238 ;
      RECT 13.835 1.94 14.08 2.195 ;
      RECT 13.81 1.956 14.095 2.107 ;
      RECT 13.81 1.975 14.12 2.098 ;
      RECT 13.805 2.012 14.12 2.05 ;
      RECT 13.81 1.992 14.125 2.018 ;
      RECT 13.905 1.926 14.015 2.415 ;
      RECT 13.991 1.925 14.015 2.415 ;
      RECT 13.225 2.71 13.23 2.921 ;
      RECT 13.825 2.71 13.83 2.895 ;
      RECT 13.89 2.75 13.895 2.863 ;
      RECT 13.885 2.742 13.89 2.869 ;
      RECT 13.88 2.732 13.885 2.877 ;
      RECT 13.875 2.722 13.88 2.886 ;
      RECT 13.87 2.712 13.875 2.89 ;
      RECT 13.83 2.71 13.87 2.893 ;
      RECT 13.802 2.709 13.825 2.897 ;
      RECT 13.716 2.706 13.802 2.904 ;
      RECT 13.63 2.702 13.716 2.915 ;
      RECT 13.61 2.7 13.63 2.921 ;
      RECT 13.592 2.699 13.61 2.924 ;
      RECT 13.506 2.697 13.592 2.931 ;
      RECT 13.42 2.692 13.506 2.944 ;
      RECT 13.401 2.689 13.42 2.949 ;
      RECT 13.315 2.687 13.401 2.94 ;
      RECT 13.305 2.687 13.315 2.933 ;
      RECT 13.23 2.7 13.305 2.927 ;
      RECT 13.215 2.711 13.225 2.921 ;
      RECT 13.205 2.713 13.215 2.92 ;
      RECT 13.195 2.717 13.205 2.916 ;
      RECT 13.19 2.72 13.195 2.91 ;
      RECT 13.18 2.722 13.19 2.904 ;
      RECT 13.175 2.725 13.18 2.898 ;
      RECT 13.155 3.311 13.16 3.515 ;
      RECT 13.14 3.298 13.155 3.608 ;
      RECT 13.125 3.279 13.14 3.885 ;
      RECT 13.09 3.245 13.125 3.885 ;
      RECT 13.086 3.215 13.09 3.885 ;
      RECT 13 3.097 13.086 3.885 ;
      RECT 12.99 2.972 13 3.885 ;
      RECT 12.975 2.94 12.99 3.885 ;
      RECT 12.97 2.915 12.975 3.885 ;
      RECT 12.965 2.905 12.97 3.841 ;
      RECT 12.95 2.877 12.965 3.746 ;
      RECT 12.935 2.843 12.95 3.645 ;
      RECT 12.93 2.821 12.935 3.598 ;
      RECT 12.925 2.81 12.93 3.568 ;
      RECT 12.92 2.8 12.925 3.534 ;
      RECT 12.91 2.787 12.92 3.502 ;
      RECT 12.885 2.763 12.91 3.428 ;
      RECT 12.88 2.743 12.885 3.353 ;
      RECT 12.875 2.737 12.88 3.328 ;
      RECT 12.87 2.732 12.875 3.293 ;
      RECT 12.865 2.727 12.87 3.268 ;
      RECT 12.86 2.725 12.865 3.248 ;
      RECT 12.855 2.725 12.86 3.233 ;
      RECT 12.85 2.725 12.855 3.193 ;
      RECT 12.84 2.725 12.85 3.165 ;
      RECT 12.83 2.725 12.84 3.11 ;
      RECT 12.815 2.725 12.83 3.048 ;
      RECT 12.81 2.724 12.815 2.993 ;
      RECT 12.795 2.723 12.81 2.973 ;
      RECT 12.735 2.721 12.795 2.947 ;
      RECT 12.7 2.722 12.735 2.927 ;
      RECT 12.695 2.724 12.7 2.917 ;
      RECT 12.685 2.743 12.695 2.907 ;
      RECT 12.68 2.77 12.685 2.838 ;
      RECT 12.795 2.195 12.965 2.44 ;
      RECT 12.83 1.966 12.965 2.44 ;
      RECT 12.83 1.968 12.975 2.435 ;
      RECT 12.83 1.97 13 2.423 ;
      RECT 12.83 1.973 13.025 2.405 ;
      RECT 12.83 1.978 13.075 2.378 ;
      RECT 12.83 1.983 13.095 2.343 ;
      RECT 12.81 1.985 13.105 2.318 ;
      RECT 12.8 2.08 13.105 2.318 ;
      RECT 12.83 1.965 12.94 2.44 ;
      RECT 12.84 1.962 12.935 2.44 ;
      RECT 12.36 3.227 12.55 3.585 ;
      RECT 12.36 3.239 12.585 3.584 ;
      RECT 12.36 3.267 12.605 3.582 ;
      RECT 12.36 3.292 12.61 3.581 ;
      RECT 12.36 3.35 12.625 3.58 ;
      RECT 12.345 3.223 12.505 3.565 ;
      RECT 12.325 3.232 12.55 3.518 ;
      RECT 12.3 3.243 12.585 3.455 ;
      RECT 12.3 3.327 12.62 3.455 ;
      RECT 12.3 3.302 12.615 3.455 ;
      RECT 12.36 3.218 12.505 3.585 ;
      RECT 12.446 3.217 12.505 3.585 ;
      RECT 12.446 3.216 12.49 3.585 ;
      RECT 12.36 7.855 12.53 8.305 ;
      RECT 12.415 6.075 12.585 8.025 ;
      RECT 12.36 5.015 12.53 6.245 ;
      RECT 11.84 5.015 12.01 8.305 ;
      RECT 11.84 7.315 12.245 7.645 ;
      RECT 11.84 6.475 12.245 6.805 ;
      RECT 12.145 2.732 12.15 3.11 ;
      RECT 12.14 2.7 12.145 3.11 ;
      RECT 12.135 2.672 12.14 3.11 ;
      RECT 12.13 2.652 12.135 3.11 ;
      RECT 12.075 2.635 12.13 3.11 ;
      RECT 12.035 2.62 12.075 3.11 ;
      RECT 11.98 2.607 12.035 3.11 ;
      RECT 11.945 2.598 11.98 3.11 ;
      RECT 11.941 2.596 11.945 3.109 ;
      RECT 11.855 2.592 11.941 3.092 ;
      RECT 11.77 2.584 11.855 3.055 ;
      RECT 11.76 2.58 11.77 3.028 ;
      RECT 11.75 2.58 11.76 3.01 ;
      RECT 11.74 2.582 11.75 2.993 ;
      RECT 11.735 2.587 11.74 2.979 ;
      RECT 11.73 2.591 11.735 2.966 ;
      RECT 11.72 2.596 11.73 2.95 ;
      RECT 11.705 2.61 11.72 2.925 ;
      RECT 11.7 2.616 11.705 2.905 ;
      RECT 11.695 2.618 11.7 2.898 ;
      RECT 11.69 2.622 11.695 2.773 ;
      RECT 11.87 3.422 12.115 3.885 ;
      RECT 11.79 3.395 12.11 3.881 ;
      RECT 11.72 3.43 12.115 3.874 ;
      RECT 11.51 3.685 12.115 3.87 ;
      RECT 11.69 3.453 12.115 3.87 ;
      RECT 11.53 3.645 12.115 3.87 ;
      RECT 11.68 3.465 12.115 3.87 ;
      RECT 11.565 3.582 12.115 3.87 ;
      RECT 11.62 3.507 12.115 3.87 ;
      RECT 11.87 3.372 12.11 3.885 ;
      RECT 11.9 3.365 12.11 3.885 ;
      RECT 11.89 3.367 12.11 3.885 ;
      RECT 11.9 3.362 12.03 3.885 ;
      RECT 11.455 1.925 11.541 2.364 ;
      RECT 11.45 1.925 11.541 2.362 ;
      RECT 11.45 1.925 11.61 2.361 ;
      RECT 11.45 1.925 11.64 2.358 ;
      RECT 11.435 1.932 11.64 2.349 ;
      RECT 11.435 1.932 11.645 2.345 ;
      RECT 11.43 1.942 11.645 2.338 ;
      RECT 11.425 1.947 11.645 2.313 ;
      RECT 11.425 1.947 11.66 2.295 ;
      RECT 11.45 1.925 11.68 2.21 ;
      RECT 11.42 1.952 11.68 2.208 ;
      RECT 11.43 1.945 11.685 2.146 ;
      RECT 11.42 2.067 11.69 2.129 ;
      RECT 11.405 1.962 11.685 2.08 ;
      RECT 11.4 1.972 11.685 1.98 ;
      RECT 11.48 2.743 11.485 2.82 ;
      RECT 11.47 2.737 11.48 3.01 ;
      RECT 11.46 2.729 11.47 3.031 ;
      RECT 11.45 2.72 11.46 3.053 ;
      RECT 11.445 2.715 11.45 3.07 ;
      RECT 11.405 2.715 11.445 3.11 ;
      RECT 11.385 2.715 11.405 3.165 ;
      RECT 11.38 2.715 11.385 3.193 ;
      RECT 11.37 2.715 11.38 3.208 ;
      RECT 11.335 2.715 11.37 3.25 ;
      RECT 11.33 2.715 11.335 3.293 ;
      RECT 11.32 2.715 11.33 3.308 ;
      RECT 11.305 2.715 11.32 3.328 ;
      RECT 11.29 2.715 11.305 3.355 ;
      RECT 11.285 2.716 11.29 3.373 ;
      RECT 11.265 2.717 11.285 3.38 ;
      RECT 11.21 2.718 11.265 3.4 ;
      RECT 11.2 2.719 11.21 3.414 ;
      RECT 11.195 2.722 11.2 3.413 ;
      RECT 11.155 2.795 11.195 3.411 ;
      RECT 11.14 2.875 11.155 3.409 ;
      RECT 11.115 2.93 11.14 3.407 ;
      RECT 11.1 2.995 11.115 3.406 ;
      RECT 11.055 3.027 11.1 3.403 ;
      RECT 10.97 3.05 11.055 3.398 ;
      RECT 10.945 3.07 10.97 3.393 ;
      RECT 10.875 3.075 10.945 3.389 ;
      RECT 10.855 3.077 10.875 3.386 ;
      RECT 10.77 3.088 10.855 3.38 ;
      RECT 10.765 3.099 10.77 3.375 ;
      RECT 10.755 3.101 10.765 3.375 ;
      RECT 10.72 3.105 10.755 3.373 ;
      RECT 10.67 3.115 10.72 3.36 ;
      RECT 10.65 3.123 10.67 3.345 ;
      RECT 10.57 3.135 10.65 3.328 ;
      RECT 10.735 2.685 10.905 2.895 ;
      RECT 10.851 2.681 10.905 2.895 ;
      RECT 10.656 2.685 10.905 2.886 ;
      RECT 10.656 2.685 10.91 2.875 ;
      RECT 10.57 2.685 10.91 2.866 ;
      RECT 10.57 2.693 10.92 2.81 ;
      RECT 10.57 2.705 10.925 2.723 ;
      RECT 10.57 2.712 10.93 2.715 ;
      RECT 10.765 2.683 10.905 2.895 ;
      RECT 10.52 3.628 10.765 3.96 ;
      RECT 10.515 3.62 10.52 3.957 ;
      RECT 10.485 3.64 10.765 3.938 ;
      RECT 10.465 3.672 10.765 3.911 ;
      RECT 10.515 3.625 10.692 3.957 ;
      RECT 10.515 3.622 10.606 3.957 ;
      RECT 10.455 1.97 10.625 2.39 ;
      RECT 10.45 1.97 10.625 2.388 ;
      RECT 10.45 1.97 10.65 2.378 ;
      RECT 10.45 1.97 10.67 2.353 ;
      RECT 10.445 1.97 10.67 2.348 ;
      RECT 10.445 1.97 10.68 2.338 ;
      RECT 10.445 1.97 10.685 2.333 ;
      RECT 10.445 1.975 10.69 2.328 ;
      RECT 10.445 2.007 10.705 2.318 ;
      RECT 10.445 2.077 10.73 2.301 ;
      RECT 10.425 2.077 10.73 2.293 ;
      RECT 10.425 2.137 10.74 2.27 ;
      RECT 10.425 2.177 10.75 2.215 ;
      RECT 10.41 1.97 10.685 2.195 ;
      RECT 10.4 1.985 10.69 2.093 ;
      RECT 9.99 3.375 10.16 3.9 ;
      RECT 9.985 3.375 10.16 3.893 ;
      RECT 9.975 3.375 10.165 3.858 ;
      RECT 9.97 3.385 10.165 3.83 ;
      RECT 9.965 3.405 10.165 3.813 ;
      RECT 9.975 3.38 10.17 3.803 ;
      RECT 9.96 3.425 10.17 3.795 ;
      RECT 9.955 3.445 10.17 3.78 ;
      RECT 9.95 3.475 10.17 3.77 ;
      RECT 9.94 3.52 10.17 3.745 ;
      RECT 9.97 3.39 10.175 3.728 ;
      RECT 9.935 3.572 10.175 3.723 ;
      RECT 9.97 3.4 10.18 3.693 ;
      RECT 9.93 3.605 10.18 3.69 ;
      RECT 9.925 3.63 10.18 3.67 ;
      RECT 9.965 3.417 10.19 3.61 ;
      RECT 9.96 3.439 10.2 3.503 ;
      RECT 9.91 2.686 9.925 2.955 ;
      RECT 9.865 2.67 9.91 3 ;
      RECT 9.86 2.658 9.865 3.05 ;
      RECT 9.85 2.654 9.86 3.083 ;
      RECT 9.845 2.651 9.85 3.111 ;
      RECT 9.83 2.653 9.845 3.153 ;
      RECT 9.825 2.657 9.83 3.193 ;
      RECT 9.805 2.662 9.825 3.245 ;
      RECT 9.801 2.667 9.805 3.302 ;
      RECT 9.715 2.686 9.801 3.339 ;
      RECT 9.705 2.707 9.715 3.375 ;
      RECT 9.7 2.715 9.705 3.376 ;
      RECT 9.695 2.757 9.7 3.377 ;
      RECT 9.68 2.845 9.695 3.378 ;
      RECT 9.67 2.995 9.68 3.38 ;
      RECT 9.665 3.04 9.67 3.382 ;
      RECT 9.63 3.082 9.665 3.385 ;
      RECT 9.625 3.1 9.63 3.388 ;
      RECT 9.548 3.106 9.625 3.394 ;
      RECT 9.462 3.12 9.548 3.407 ;
      RECT 9.376 3.134 9.462 3.421 ;
      RECT 9.29 3.148 9.376 3.434 ;
      RECT 9.23 3.16 9.29 3.446 ;
      RECT 9.205 3.167 9.23 3.453 ;
      RECT 9.191 3.17 9.205 3.458 ;
      RECT 9.105 3.178 9.191 3.474 ;
      RECT 9.1 3.185 9.105 3.489 ;
      RECT 9.076 3.185 9.1 3.496 ;
      RECT 8.99 3.188 9.076 3.524 ;
      RECT 8.905 3.192 8.99 3.568 ;
      RECT 8.84 3.196 8.905 3.605 ;
      RECT 8.815 3.199 8.84 3.621 ;
      RECT 8.74 3.212 8.815 3.625 ;
      RECT 8.715 3.23 8.74 3.629 ;
      RECT 8.705 3.237 8.715 3.631 ;
      RECT 8.69 3.24 8.705 3.632 ;
      RECT 8.63 3.252 8.69 3.636 ;
      RECT 8.62 3.266 8.63 3.64 ;
      RECT 8.565 3.276 8.62 3.628 ;
      RECT 8.54 3.297 8.565 3.611 ;
      RECT 8.52 3.317 8.54 3.602 ;
      RECT 8.515 3.33 8.52 3.597 ;
      RECT 8.5 3.342 8.515 3.593 ;
      RECT 9.735 1.997 9.74 2.02 ;
      RECT 9.73 1.988 9.735 2.06 ;
      RECT 9.725 1.986 9.73 2.103 ;
      RECT 9.72 1.977 9.725 2.138 ;
      RECT 9.715 1.967 9.72 2.21 ;
      RECT 9.71 1.957 9.715 2.275 ;
      RECT 9.705 1.954 9.71 2.315 ;
      RECT 9.68 1.948 9.705 2.405 ;
      RECT 9.645 1.936 9.68 2.43 ;
      RECT 9.635 1.927 9.645 2.43 ;
      RECT 9.5 1.925 9.51 2.413 ;
      RECT 9.49 1.925 9.5 2.38 ;
      RECT 9.485 1.925 9.49 2.355 ;
      RECT 9.48 1.925 9.485 2.343 ;
      RECT 9.475 1.925 9.48 2.325 ;
      RECT 9.465 1.925 9.475 2.29 ;
      RECT 9.46 1.927 9.465 2.268 ;
      RECT 9.455 1.933 9.46 2.253 ;
      RECT 9.45 1.939 9.455 2.238 ;
      RECT 9.435 1.951 9.45 2.211 ;
      RECT 9.43 1.962 9.435 2.179 ;
      RECT 9.425 1.972 9.43 2.163 ;
      RECT 9.415 1.98 9.425 2.132 ;
      RECT 9.41 1.99 9.415 2.106 ;
      RECT 9.405 2.047 9.41 2.089 ;
      RECT 9.51 1.925 9.635 2.43 ;
      RECT 9.225 2.612 9.485 2.91 ;
      RECT 9.22 2.619 9.485 2.908 ;
      RECT 9.225 2.614 9.5 2.903 ;
      RECT 9.215 2.627 9.5 2.9 ;
      RECT 9.215 2.632 9.505 2.893 ;
      RECT 9.21 2.64 9.505 2.89 ;
      RECT 9.21 2.657 9.51 2.688 ;
      RECT 9.225 2.609 9.456 2.91 ;
      RECT 9.28 2.608 9.456 2.91 ;
      RECT 9.28 2.605 9.37 2.91 ;
      RECT 9.28 2.602 9.366 2.91 ;
      RECT 8.97 2.875 8.975 2.888 ;
      RECT 8.965 2.842 8.97 2.893 ;
      RECT 8.96 2.797 8.965 2.9 ;
      RECT 8.955 2.752 8.96 2.908 ;
      RECT 8.95 2.72 8.955 2.916 ;
      RECT 8.945 2.68 8.95 2.917 ;
      RECT 8.93 2.66 8.945 2.919 ;
      RECT 8.855 2.642 8.93 2.931 ;
      RECT 8.845 2.635 8.855 2.942 ;
      RECT 8.84 2.635 8.845 2.944 ;
      RECT 8.81 2.641 8.84 2.948 ;
      RECT 8.77 2.654 8.81 2.948 ;
      RECT 8.745 2.665 8.77 2.934 ;
      RECT 8.73 2.671 8.745 2.917 ;
      RECT 8.72 2.673 8.73 2.908 ;
      RECT 8.715 2.674 8.72 2.903 ;
      RECT 8.71 2.675 8.715 2.898 ;
      RECT 8.705 2.676 8.71 2.895 ;
      RECT 8.68 2.681 8.705 2.885 ;
      RECT 8.67 2.697 8.68 2.872 ;
      RECT 8.665 2.717 8.67 2.867 ;
      RECT 8.675 2.11 8.68 2.306 ;
      RECT 8.66 2.074 8.675 2.308 ;
      RECT 8.65 2.056 8.66 2.313 ;
      RECT 8.64 2.042 8.65 2.317 ;
      RECT 8.595 2.026 8.64 2.327 ;
      RECT 8.59 2.016 8.595 2.336 ;
      RECT 8.545 2.005 8.59 2.342 ;
      RECT 8.54 1.993 8.545 2.349 ;
      RECT 8.525 1.988 8.54 2.353 ;
      RECT 8.51 1.98 8.525 2.358 ;
      RECT 8.5 1.973 8.51 2.363 ;
      RECT 8.49 1.97 8.5 2.368 ;
      RECT 8.48 1.97 8.49 2.369 ;
      RECT 8.475 1.967 8.48 2.368 ;
      RECT 8.44 1.962 8.465 2.367 ;
      RECT 8.416 1.958 8.44 2.366 ;
      RECT 8.33 1.949 8.416 2.363 ;
      RECT 8.315 1.941 8.33 2.36 ;
      RECT 8.293 1.94 8.315 2.359 ;
      RECT 8.207 1.94 8.293 2.357 ;
      RECT 8.121 1.94 8.207 2.355 ;
      RECT 8.035 1.94 8.121 2.352 ;
      RECT 8.025 1.94 8.035 2.343 ;
      RECT 7.995 1.94 8.025 2.303 ;
      RECT 7.985 1.95 7.995 2.258 ;
      RECT 7.98 1.99 7.985 2.243 ;
      RECT 7.975 2.005 7.98 2.23 ;
      RECT 7.945 2.085 7.975 2.192 ;
      RECT 8.465 1.965 8.475 2.368 ;
      RECT 8.29 2.73 8.305 3.335 ;
      RECT 8.295 2.725 8.305 3.335 ;
      RECT 8.46 2.725 8.465 2.908 ;
      RECT 8.45 2.725 8.46 2.938 ;
      RECT 8.435 2.725 8.45 2.998 ;
      RECT 8.43 2.725 8.435 3.043 ;
      RECT 8.425 2.725 8.43 3.073 ;
      RECT 8.42 2.725 8.425 3.093 ;
      RECT 8.41 2.725 8.42 3.128 ;
      RECT 8.395 2.725 8.41 3.16 ;
      RECT 8.35 2.725 8.395 3.188 ;
      RECT 8.345 2.725 8.35 3.218 ;
      RECT 8.34 2.725 8.345 3.23 ;
      RECT 8.335 2.725 8.34 3.238 ;
      RECT 8.325 2.725 8.335 3.253 ;
      RECT 8.32 2.725 8.325 3.275 ;
      RECT 8.31 2.725 8.32 3.298 ;
      RECT 8.305 2.725 8.31 3.318 ;
      RECT 8.27 2.74 8.29 3.335 ;
      RECT 8.245 2.757 8.27 3.335 ;
      RECT 8.24 2.767 8.245 3.335 ;
      RECT 8.21 2.782 8.24 3.335 ;
      RECT 8.135 2.824 8.21 3.335 ;
      RECT 8.13 2.855 8.135 3.318 ;
      RECT 8.125 2.859 8.13 3.3 ;
      RECT 8.12 2.863 8.125 3.263 ;
      RECT 8.115 3.047 8.12 3.23 ;
      RECT 7.6 3.236 7.686 3.801 ;
      RECT 7.555 3.238 7.72 3.795 ;
      RECT 7.686 3.235 7.72 3.795 ;
      RECT 7.6 3.237 7.805 3.789 ;
      RECT 7.555 3.247 7.815 3.785 ;
      RECT 7.53 3.239 7.805 3.781 ;
      RECT 7.525 3.242 7.805 3.776 ;
      RECT 7.5 3.257 7.815 3.77 ;
      RECT 7.5 3.282 7.855 3.765 ;
      RECT 7.46 3.29 7.855 3.74 ;
      RECT 7.46 3.317 7.87 3.738 ;
      RECT 7.46 3.347 7.88 3.725 ;
      RECT 7.455 3.492 7.88 3.713 ;
      RECT 7.46 3.421 7.9 3.71 ;
      RECT 7.46 3.478 7.905 3.518 ;
      RECT 7.65 2.757 7.82 2.935 ;
      RECT 7.6 2.696 7.65 2.92 ;
      RECT 7.335 2.676 7.6 2.905 ;
      RECT 7.295 2.74 7.77 2.905 ;
      RECT 7.295 2.73 7.725 2.905 ;
      RECT 7.295 2.727 7.715 2.905 ;
      RECT 7.295 2.715 7.705 2.905 ;
      RECT 7.295 2.7 7.65 2.905 ;
      RECT 7.335 2.672 7.536 2.905 ;
      RECT 7.345 2.65 7.536 2.905 ;
      RECT 7.37 2.635 7.45 2.905 ;
      RECT 7.125 3.165 7.245 3.61 ;
      RECT 7.11 3.165 7.245 3.609 ;
      RECT 7.065 3.187 7.245 3.604 ;
      RECT 7.025 3.236 7.245 3.598 ;
      RECT 7.025 3.236 7.25 3.573 ;
      RECT 7.025 3.236 7.27 3.463 ;
      RECT 7.02 3.266 7.27 3.46 ;
      RECT 7.11 3.165 7.28 3.355 ;
      RECT 6.77 1.95 6.775 2.395 ;
      RECT 6.58 1.95 6.6 2.36 ;
      RECT 6.55 1.95 6.555 2.335 ;
      RECT 7.23 2.257 7.245 2.445 ;
      RECT 7.225 2.242 7.23 2.451 ;
      RECT 7.205 2.215 7.225 2.454 ;
      RECT 7.155 2.182 7.205 2.463 ;
      RECT 7.125 2.162 7.155 2.467 ;
      RECT 7.106 2.15 7.125 2.463 ;
      RECT 7.02 2.122 7.106 2.453 ;
      RECT 7.01 2.097 7.02 2.443 ;
      RECT 6.94 2.065 7.01 2.435 ;
      RECT 6.915 2.025 6.94 2.427 ;
      RECT 6.895 2.007 6.915 2.421 ;
      RECT 6.885 1.997 6.895 2.418 ;
      RECT 6.875 1.99 6.885 2.416 ;
      RECT 6.855 1.977 6.875 2.413 ;
      RECT 6.845 1.967 6.855 2.41 ;
      RECT 6.835 1.96 6.845 2.408 ;
      RECT 6.785 1.952 6.835 2.402 ;
      RECT 6.775 1.95 6.785 2.396 ;
      RECT 6.745 1.95 6.77 2.393 ;
      RECT 6.716 1.95 6.745 2.388 ;
      RECT 6.63 1.95 6.716 2.378 ;
      RECT 6.6 1.95 6.63 2.365 ;
      RECT 6.555 1.95 6.58 2.348 ;
      RECT 6.54 1.95 6.55 2.33 ;
      RECT 6.52 1.957 6.54 2.315 ;
      RECT 6.515 1.972 6.52 2.303 ;
      RECT 6.51 1.977 6.515 2.243 ;
      RECT 6.505 1.982 6.51 2.085 ;
      RECT 6.5 1.985 6.505 2.003 ;
      RECT 6.765 2.67 6.851 2.991 ;
      RECT 6.765 2.67 6.885 2.984 ;
      RECT 6.715 2.67 6.885 2.98 ;
      RECT 6.715 2.672 6.971 2.978 ;
      RECT 6.715 2.674 6.995 2.972 ;
      RECT 6.715 2.681 7.005 2.971 ;
      RECT 6.715 2.69 7.01 2.968 ;
      RECT 6.715 2.696 7.015 2.963 ;
      RECT 6.715 2.74 7.02 2.96 ;
      RECT 6.715 2.832 7.025 2.957 ;
      RECT 6.24 3.275 6.275 3.595 ;
      RECT 6.825 3.46 6.83 3.642 ;
      RECT 6.78 3.342 6.825 3.661 ;
      RECT 6.765 3.319 6.78 3.684 ;
      RECT 6.755 3.309 6.765 3.694 ;
      RECT 6.735 3.304 6.755 3.707 ;
      RECT 6.71 3.302 6.735 3.728 ;
      RECT 6.691 3.301 6.71 3.74 ;
      RECT 6.605 3.298 6.691 3.74 ;
      RECT 6.535 3.293 6.605 3.728 ;
      RECT 6.46 3.289 6.535 3.703 ;
      RECT 6.395 3.285 6.46 3.67 ;
      RECT 6.325 3.282 6.395 3.63 ;
      RECT 6.295 3.278 6.325 3.605 ;
      RECT 6.275 3.276 6.295 3.598 ;
      RECT 6.191 3.274 6.24 3.596 ;
      RECT 6.105 3.271 6.191 3.597 ;
      RECT 6.03 3.27 6.105 3.599 ;
      RECT 5.945 3.27 6.03 3.625 ;
      RECT 5.868 3.271 5.945 3.65 ;
      RECT 5.782 3.272 5.868 3.65 ;
      RECT 5.696 3.272 5.782 3.65 ;
      RECT 5.61 3.273 5.696 3.65 ;
      RECT 5.59 3.274 5.61 3.642 ;
      RECT 5.575 3.28 5.59 3.627 ;
      RECT 5.54 3.3 5.575 3.607 ;
      RECT 5.53 3.32 5.54 3.589 ;
      RECT 6.5 2.625 6.505 2.895 ;
      RECT 6.495 2.616 6.5 2.9 ;
      RECT 6.485 2.606 6.495 2.912 ;
      RECT 6.48 2.595 6.485 2.923 ;
      RECT 6.46 2.589 6.48 2.941 ;
      RECT 6.415 2.586 6.46 2.99 ;
      RECT 6.4 2.585 6.415 3.035 ;
      RECT 6.395 2.585 6.4 3.048 ;
      RECT 6.385 2.585 6.395 3.06 ;
      RECT 6.38 2.586 6.385 3.075 ;
      RECT 6.36 2.594 6.38 3.08 ;
      RECT 6.33 2.61 6.36 3.08 ;
      RECT 6.32 2.622 6.325 3.08 ;
      RECT 6.285 2.637 6.32 3.08 ;
      RECT 6.255 2.657 6.285 3.08 ;
      RECT 6.245 2.682 6.255 3.08 ;
      RECT 6.24 2.71 6.245 3.08 ;
      RECT 6.235 2.74 6.24 3.08 ;
      RECT 6.23 2.757 6.235 3.08 ;
      RECT 6.22 2.785 6.23 3.08 ;
      RECT 6.21 2.82 6.22 3.08 ;
      RECT 6.205 2.855 6.21 3.08 ;
      RECT 6.325 2.62 6.33 3.08 ;
      RECT 5.84 2.722 6.025 2.895 ;
      RECT 5.8 2.64 5.985 2.893 ;
      RECT 5.761 2.645 5.985 2.889 ;
      RECT 5.675 2.654 5.985 2.884 ;
      RECT 5.591 2.67 5.99 2.879 ;
      RECT 5.505 2.69 6.015 2.873 ;
      RECT 5.505 2.71 6.02 2.873 ;
      RECT 5.591 2.68 6.015 2.879 ;
      RECT 5.675 2.655 5.99 2.884 ;
      RECT 5.84 2.637 5.985 2.895 ;
      RECT 5.84 2.632 5.94 2.895 ;
      RECT 5.926 2.626 5.94 2.895 ;
      RECT 5.315 1.95 5.32 2.349 ;
      RECT 5.06 1.95 5.095 2.347 ;
      RECT 4.655 1.985 4.66 2.341 ;
      RECT 5.4 1.988 5.405 2.243 ;
      RECT 5.395 1.986 5.4 2.249 ;
      RECT 5.39 1.985 5.395 2.256 ;
      RECT 5.365 1.978 5.39 2.28 ;
      RECT 5.36 1.971 5.365 2.304 ;
      RECT 5.355 1.967 5.36 2.313 ;
      RECT 5.345 1.962 5.355 2.326 ;
      RECT 5.34 1.959 5.345 2.335 ;
      RECT 5.335 1.957 5.34 2.34 ;
      RECT 5.32 1.953 5.335 2.35 ;
      RECT 5.305 1.947 5.315 2.349 ;
      RECT 5.267 1.945 5.305 2.349 ;
      RECT 5.181 1.947 5.267 2.349 ;
      RECT 5.095 1.949 5.181 2.348 ;
      RECT 5.024 1.95 5.06 2.347 ;
      RECT 4.938 1.952 5.024 2.347 ;
      RECT 4.852 1.954 4.938 2.346 ;
      RECT 4.766 1.956 4.852 2.346 ;
      RECT 4.68 1.959 4.766 2.345 ;
      RECT 4.67 1.965 4.68 2.344 ;
      RECT 4.66 1.977 4.67 2.342 ;
      RECT 4.6 2.012 4.655 2.338 ;
      RECT 4.595 2.042 4.6 2.1 ;
      RECT 5.34 3.122 5.355 3.315 ;
      RECT 5.335 3.09 5.34 3.315 ;
      RECT 5.325 3.065 5.335 3.315 ;
      RECT 5.32 3.037 5.325 3.315 ;
      RECT 5.29 2.96 5.32 3.315 ;
      RECT 5.265 2.842 5.29 3.315 ;
      RECT 5.26 2.78 5.265 3.315 ;
      RECT 5.25 2.767 5.26 3.315 ;
      RECT 5.23 2.757 5.25 3.315 ;
      RECT 5.215 2.74 5.23 3.315 ;
      RECT 5.185 2.728 5.215 3.315 ;
      RECT 5.18 2.727 5.185 3.26 ;
      RECT 5.175 2.727 5.18 3.218 ;
      RECT 5.16 2.726 5.175 3.17 ;
      RECT 5.145 2.726 5.16 3.108 ;
      RECT 5.125 2.726 5.145 3.068 ;
      RECT 5.12 2.726 5.125 3.053 ;
      RECT 5.095 2.725 5.12 3.048 ;
      RECT 5.025 2.724 5.095 3.035 ;
      RECT 5.01 2.723 5.025 3.02 ;
      RECT 4.98 2.722 5.01 3.003 ;
      RECT 4.975 2.722 4.98 2.988 ;
      RECT 4.925 2.721 4.975 2.968 ;
      RECT 4.86 2.72 4.925 2.923 ;
      RECT 4.855 2.72 4.86 2.895 ;
      RECT 4.94 3.257 4.945 3.514 ;
      RECT 4.92 3.176 4.94 3.531 ;
      RECT 4.9 3.17 4.92 3.56 ;
      RECT 4.84 3.157 4.9 3.58 ;
      RECT 4.795 3.141 4.84 3.581 ;
      RECT 4.711 3.129 4.795 3.569 ;
      RECT 4.625 3.116 4.711 3.553 ;
      RECT 4.615 3.109 4.625 3.545 ;
      RECT 4.57 3.106 4.615 3.485 ;
      RECT 4.55 3.102 4.57 3.4 ;
      RECT 4.535 3.1 4.55 3.353 ;
      RECT 4.505 3.097 4.535 3.323 ;
      RECT 4.47 3.093 4.505 3.3 ;
      RECT 4.427 3.088 4.47 3.288 ;
      RECT 4.341 3.079 4.427 3.297 ;
      RECT 4.255 3.068 4.341 3.309 ;
      RECT 4.19 3.059 4.255 3.318 ;
      RECT 4.17 3.05 4.19 3.323 ;
      RECT 4.165 3.043 4.17 3.325 ;
      RECT 4.125 3.028 4.165 3.322 ;
      RECT 4.105 3.007 4.125 3.317 ;
      RECT 4.09 2.995 4.105 3.31 ;
      RECT 4.085 2.987 4.09 3.303 ;
      RECT 4.07 2.967 4.085 3.296 ;
      RECT 4.065 2.83 4.07 3.29 ;
      RECT 3.985 2.719 4.065 3.262 ;
      RECT 3.976 2.712 3.985 3.228 ;
      RECT 3.89 2.706 3.976 3.153 ;
      RECT 3.865 2.697 3.89 3.065 ;
      RECT 3.835 2.692 3.865 3.04 ;
      RECT 3.77 2.701 3.835 3.025 ;
      RECT 3.75 2.717 3.77 3 ;
      RECT 3.74 2.723 3.75 2.948 ;
      RECT 3.72 2.745 3.74 2.83 ;
      RECT 4.375 2.71 4.545 2.895 ;
      RECT 4.375 2.71 4.58 2.893 ;
      RECT 4.425 2.62 4.595 2.884 ;
      RECT 4.375 2.777 4.6 2.877 ;
      RECT 4.39 2.655 4.595 2.884 ;
      RECT 3.59 3.388 3.655 3.831 ;
      RECT 3.53 3.413 3.655 3.829 ;
      RECT 3.53 3.413 3.71 3.823 ;
      RECT 3.515 3.438 3.71 3.822 ;
      RECT 3.655 3.375 3.73 3.819 ;
      RECT 3.59 3.4 3.81 3.813 ;
      RECT 3.515 3.439 3.855 3.807 ;
      RECT 3.5 3.466 3.855 3.798 ;
      RECT 3.515 3.459 3.875 3.79 ;
      RECT 3.5 3.468 3.88 3.773 ;
      RECT 3.495 3.485 3.88 3.6 ;
      RECT 3.5 2.207 3.535 2.445 ;
      RECT 3.5 2.207 3.565 2.444 ;
      RECT 3.5 2.207 3.68 2.44 ;
      RECT 3.5 2.207 3.735 2.418 ;
      RECT 3.51 2.15 3.79 2.318 ;
      RECT 3.615 1.99 3.645 2.441 ;
      RECT 3.645 1.985 3.825 2.198 ;
      RECT 3.515 2.126 3.825 2.198 ;
      RECT 3.565 2.022 3.615 2.442 ;
      RECT 3.535 2.078 3.825 2.198 ;
      RECT 1.33 7.855 1.5 8.305 ;
      RECT 1.385 6.075 1.555 8.025 ;
      RECT 1.33 5.015 1.5 6.245 ;
      RECT 0.81 5.015 0.98 8.305 ;
      RECT 0.81 7.315 1.215 7.645 ;
      RECT 0.81 6.475 1.215 6.805 ;
      RECT 92.03 7.8 92.2 8.31 ;
      RECT 91.04 0.57 91.21 1.08 ;
      RECT 91.04 2.39 91.21 3.86 ;
      RECT 91.04 5.02 91.21 6.49 ;
      RECT 91.04 7.8 91.21 8.31 ;
      RECT 89.68 0.575 89.85 3.865 ;
      RECT 89.68 5.015 89.85 8.305 ;
      RECT 89.25 0.575 89.42 1.085 ;
      RECT 89.25 1.655 89.42 3.865 ;
      RECT 89.25 5.015 89.42 7.225 ;
      RECT 89.25 7.795 89.42 8.305 ;
      RECT 84.92 5.015 85.09 8.305 ;
      RECT 84.49 5.015 84.66 7.225 ;
      RECT 84.49 7.795 84.66 8.305 ;
      RECT 74.105 7.8 74.275 8.31 ;
      RECT 73.115 0.57 73.285 1.08 ;
      RECT 73.115 2.39 73.285 3.86 ;
      RECT 73.115 5.02 73.285 6.49 ;
      RECT 73.115 7.8 73.285 8.31 ;
      RECT 71.755 0.575 71.925 3.865 ;
      RECT 71.755 5.015 71.925 8.305 ;
      RECT 71.325 0.575 71.495 1.085 ;
      RECT 71.325 1.655 71.495 3.865 ;
      RECT 71.325 5.015 71.495 7.225 ;
      RECT 71.325 7.795 71.495 8.305 ;
      RECT 66.995 5.015 67.165 8.305 ;
      RECT 66.565 5.015 66.735 7.225 ;
      RECT 66.565 7.795 66.735 8.305 ;
      RECT 56.18 7.8 56.35 8.31 ;
      RECT 55.19 0.57 55.36 1.08 ;
      RECT 55.19 2.39 55.36 3.86 ;
      RECT 55.19 5.02 55.36 6.49 ;
      RECT 55.19 7.8 55.36 8.31 ;
      RECT 53.83 0.575 54 3.865 ;
      RECT 53.83 5.015 54 8.305 ;
      RECT 53.4 0.575 53.57 1.085 ;
      RECT 53.4 1.655 53.57 3.865 ;
      RECT 53.4 5.015 53.57 7.225 ;
      RECT 53.4 7.795 53.57 8.305 ;
      RECT 49.07 5.015 49.24 8.305 ;
      RECT 48.64 5.015 48.81 7.225 ;
      RECT 48.64 7.795 48.81 8.305 ;
      RECT 38.255 7.8 38.425 8.31 ;
      RECT 37.265 0.57 37.435 1.08 ;
      RECT 37.265 2.39 37.435 3.86 ;
      RECT 37.265 5.02 37.435 6.49 ;
      RECT 37.265 7.8 37.435 8.31 ;
      RECT 35.905 0.575 36.075 3.865 ;
      RECT 35.905 5.015 36.075 8.305 ;
      RECT 35.475 0.575 35.645 1.085 ;
      RECT 35.475 1.655 35.645 3.865 ;
      RECT 35.475 5.015 35.645 7.225 ;
      RECT 35.475 7.795 35.645 8.305 ;
      RECT 31.145 5.015 31.315 8.305 ;
      RECT 30.715 5.015 30.885 7.225 ;
      RECT 30.715 7.795 30.885 8.305 ;
      RECT 20.33 7.8 20.5 8.31 ;
      RECT 19.34 0.57 19.51 1.08 ;
      RECT 19.34 2.39 19.51 3.86 ;
      RECT 19.34 5.02 19.51 6.49 ;
      RECT 19.34 7.8 19.51 8.31 ;
      RECT 17.98 0.575 18.15 3.865 ;
      RECT 17.98 5.015 18.15 8.305 ;
      RECT 17.55 0.575 17.72 1.085 ;
      RECT 17.55 1.655 17.72 3.865 ;
      RECT 17.55 5.015 17.72 7.225 ;
      RECT 17.55 7.795 17.72 8.305 ;
      RECT 13.22 5.015 13.39 8.305 ;
      RECT 12.79 5.015 12.96 7.225 ;
      RECT 12.79 7.795 12.96 8.305 ;
      RECT 1.76 5.015 1.93 7.225 ;
      RECT 1.76 7.795 1.93 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2at_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2ca_8_b0r1
  CLASS BLOCK ;
  ORIGIN 0.025 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ca_8_b0r1 ;
  SIZE 85.755 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 18.825 0.915 18.995 1.085 ;
        RECT 18.82 0.91 18.99 1.08 ;
        RECT 18.825 2.395 18.995 2.565 ;
        RECT 18.82 2.39 18.99 2.56 ;
      LAYER li1 ;
        RECT 18.825 0.915 18.995 1.085 ;
        RECT 18.82 0.57 18.99 1.08 ;
        RECT 18.82 2.395 18.995 2.565 ;
        RECT 18.82 2.39 18.99 3.86 ;
      LAYER met1 ;
        RECT 18.76 2.36 19.05 2.59 ;
        RECT 18.76 0.88 19.05 1.11 ;
        RECT 18.82 0.88 18.99 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 35.41 0.915 35.58 1.085 ;
        RECT 35.405 0.91 35.575 1.08 ;
        RECT 35.41 2.395 35.58 2.565 ;
        RECT 35.405 2.39 35.575 2.56 ;
      LAYER li1 ;
        RECT 35.41 0.915 35.58 1.085 ;
        RECT 35.405 0.57 35.575 1.08 ;
        RECT 35.405 2.395 35.58 2.565 ;
        RECT 35.405 2.39 35.575 3.86 ;
      LAYER met1 ;
        RECT 35.345 2.36 35.635 2.59 ;
        RECT 35.345 0.88 35.635 1.11 ;
        RECT 35.405 0.88 35.575 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 51.995 0.915 52.165 1.085 ;
        RECT 51.99 0.91 52.16 1.08 ;
        RECT 51.995 2.395 52.165 2.565 ;
        RECT 51.99 2.39 52.16 2.56 ;
      LAYER li1 ;
        RECT 51.995 0.915 52.165 1.085 ;
        RECT 51.99 0.57 52.16 1.08 ;
        RECT 51.99 2.395 52.165 2.565 ;
        RECT 51.99 2.39 52.16 3.86 ;
      LAYER met1 ;
        RECT 51.93 2.36 52.22 2.59 ;
        RECT 51.93 0.88 52.22 1.11 ;
        RECT 51.99 0.88 52.16 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 68.58 0.915 68.75 1.085 ;
        RECT 68.575 0.91 68.745 1.08 ;
        RECT 68.58 2.395 68.75 2.565 ;
        RECT 68.575 2.39 68.745 2.56 ;
      LAYER li1 ;
        RECT 68.58 0.915 68.75 1.085 ;
        RECT 68.575 0.57 68.745 1.08 ;
        RECT 68.575 2.395 68.75 2.565 ;
        RECT 68.575 2.39 68.745 3.86 ;
      LAYER met1 ;
        RECT 68.515 2.36 68.805 2.59 ;
        RECT 68.515 0.88 68.805 1.11 ;
        RECT 68.575 0.88 68.745 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 85.16 0.915 85.33 1.085 ;
        RECT 85.155 0.91 85.325 1.08 ;
        RECT 85.16 2.395 85.33 2.565 ;
        RECT 85.155 2.39 85.325 2.56 ;
      LAYER li1 ;
        RECT 85.16 0.915 85.33 1.085 ;
        RECT 85.155 0.57 85.325 1.08 ;
        RECT 85.155 2.395 85.33 2.565 ;
        RECT 85.155 2.39 85.325 3.86 ;
      LAYER met1 ;
        RECT 85.095 2.36 85.385 2.59 ;
        RECT 85.095 0.88 85.385 1.11 ;
        RECT 85.155 0.88 85.325 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 14.67 1.66 14.84 2.935 ;
        RECT 14.67 5.945 14.84 7.22 ;
        RECT 3.445 5.945 3.615 7.22 ;
      LAYER met2 ;
        RECT 14.595 5.865 14.92 6.19 ;
        RECT 14.59 3.635 14.915 3.96 ;
        RECT 5.75 7.885 14.835 8.055 ;
        RECT 14.66 3.635 14.835 8.055 ;
        RECT 5.695 5.86 5.975 6.2 ;
        RECT 5.75 5.86 5.92 8.055 ;
      LAYER met1 ;
        RECT 14.61 2.765 15.07 2.935 ;
        RECT 14.59 3.635 14.915 3.96 ;
        RECT 14.61 2.735 14.9 2.965 ;
        RECT 14.665 2.735 14.845 3.96 ;
        RECT 14.595 5.945 15.07 6.115 ;
        RECT 14.595 5.865 14.92 6.19 ;
        RECT 5.665 5.89 6.005 6.17 ;
        RECT 3.385 5.945 6.005 6.115 ;
        RECT 3.385 5.915 3.675 6.145 ;
      LAYER via1 ;
        RECT 5.76 5.955 5.91 6.105 ;
        RECT 14.68 3.72 14.83 3.87 ;
        RECT 14.685 5.95 14.835 6.1 ;
      LAYER mcon ;
        RECT 3.445 5.945 3.615 6.115 ;
        RECT 14.67 5.945 14.84 6.115 ;
        RECT 14.67 2.765 14.84 2.935 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 31.255 1.66 31.425 2.935 ;
        RECT 31.255 5.945 31.425 7.22 ;
        RECT 20.03 5.945 20.2 7.22 ;
      LAYER met2 ;
        RECT 31.18 5.865 31.505 6.19 ;
        RECT 31.175 3.635 31.5 3.96 ;
        RECT 22.335 7.885 31.42 8.055 ;
        RECT 31.245 3.635 31.42 8.055 ;
        RECT 22.28 5.86 22.56 6.2 ;
        RECT 22.335 5.86 22.505 8.055 ;
      LAYER met1 ;
        RECT 31.195 2.765 31.655 2.935 ;
        RECT 31.175 3.635 31.5 3.96 ;
        RECT 31.195 2.735 31.485 2.965 ;
        RECT 31.25 2.735 31.43 3.96 ;
        RECT 31.18 5.945 31.655 6.115 ;
        RECT 31.18 5.865 31.505 6.19 ;
        RECT 22.25 5.89 22.59 6.17 ;
        RECT 19.97 5.945 22.59 6.115 ;
        RECT 19.97 5.915 20.26 6.145 ;
      LAYER via1 ;
        RECT 22.345 5.955 22.495 6.105 ;
        RECT 31.265 3.72 31.415 3.87 ;
        RECT 31.27 5.95 31.42 6.1 ;
      LAYER mcon ;
        RECT 20.03 5.945 20.2 6.115 ;
        RECT 31.255 5.945 31.425 6.115 ;
        RECT 31.255 2.765 31.425 2.935 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 47.84 1.66 48.01 2.935 ;
        RECT 47.84 5.945 48.01 7.22 ;
        RECT 36.615 5.945 36.785 7.22 ;
      LAYER met2 ;
        RECT 47.765 5.865 48.09 6.19 ;
        RECT 47.76 3.635 48.085 3.96 ;
        RECT 38.92 7.885 48.005 8.055 ;
        RECT 47.83 3.635 48.005 8.055 ;
        RECT 38.865 5.86 39.145 6.2 ;
        RECT 38.92 5.86 39.09 8.055 ;
      LAYER met1 ;
        RECT 47.78 2.765 48.24 2.935 ;
        RECT 47.76 3.635 48.085 3.96 ;
        RECT 47.78 2.735 48.07 2.965 ;
        RECT 47.835 2.735 48.015 3.96 ;
        RECT 47.765 5.945 48.24 6.115 ;
        RECT 47.765 5.865 48.09 6.19 ;
        RECT 38.835 5.89 39.175 6.17 ;
        RECT 36.555 5.945 39.175 6.115 ;
        RECT 36.555 5.915 36.845 6.145 ;
      LAYER via1 ;
        RECT 38.93 5.955 39.08 6.105 ;
        RECT 47.85 3.72 48 3.87 ;
        RECT 47.855 5.95 48.005 6.1 ;
      LAYER mcon ;
        RECT 36.615 5.945 36.785 6.115 ;
        RECT 47.84 5.945 48.01 6.115 ;
        RECT 47.84 2.765 48.01 2.935 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 64.425 1.66 64.595 2.935 ;
        RECT 64.425 5.945 64.595 7.22 ;
        RECT 53.2 5.945 53.37 7.22 ;
      LAYER met2 ;
        RECT 64.35 5.865 64.675 6.19 ;
        RECT 64.345 3.635 64.67 3.96 ;
        RECT 55.505 7.885 64.59 8.055 ;
        RECT 64.415 3.635 64.59 8.055 ;
        RECT 55.45 5.86 55.73 6.2 ;
        RECT 55.505 5.86 55.675 8.055 ;
      LAYER met1 ;
        RECT 64.365 2.765 64.825 2.935 ;
        RECT 64.345 3.635 64.67 3.96 ;
        RECT 64.365 2.735 64.655 2.965 ;
        RECT 64.42 2.735 64.6 3.96 ;
        RECT 64.35 5.945 64.825 6.115 ;
        RECT 64.35 5.865 64.675 6.19 ;
        RECT 55.42 5.89 55.76 6.17 ;
        RECT 53.14 5.945 55.76 6.115 ;
        RECT 53.14 5.915 53.43 6.145 ;
      LAYER via1 ;
        RECT 55.515 5.955 55.665 6.105 ;
        RECT 64.435 3.72 64.585 3.87 ;
        RECT 64.44 5.95 64.59 6.1 ;
      LAYER mcon ;
        RECT 53.2 5.945 53.37 6.115 ;
        RECT 64.425 5.945 64.595 6.115 ;
        RECT 64.425 2.765 64.595 2.935 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 81.005 1.66 81.175 2.935 ;
        RECT 81.005 5.945 81.175 7.22 ;
        RECT 69.78 5.945 69.95 7.22 ;
      LAYER met2 ;
        RECT 80.93 5.865 81.255 6.19 ;
        RECT 80.925 3.635 81.25 3.96 ;
        RECT 72.085 7.885 81.17 8.055 ;
        RECT 80.995 3.635 81.17 8.055 ;
        RECT 72.03 5.86 72.31 6.2 ;
        RECT 72.085 5.86 72.255 8.055 ;
      LAYER met1 ;
        RECT 80.945 2.765 81.405 2.935 ;
        RECT 80.925 3.635 81.25 3.96 ;
        RECT 80.945 2.735 81.235 2.965 ;
        RECT 81 2.735 81.18 3.96 ;
        RECT 80.93 5.945 81.405 6.115 ;
        RECT 80.93 5.865 81.255 6.19 ;
        RECT 72 5.89 72.34 6.17 ;
        RECT 69.72 5.945 72.34 6.115 ;
        RECT 69.72 5.915 70.01 6.145 ;
      LAYER via1 ;
        RECT 72.095 5.955 72.245 6.105 ;
        RECT 81.015 3.72 81.165 3.87 ;
        RECT 81.02 5.95 81.17 6.1 ;
      LAYER mcon ;
        RECT 69.78 5.945 69.95 6.115 ;
        RECT 81.005 5.945 81.175 6.115 ;
        RECT 81.005 2.765 81.175 2.935 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 0.215 5.945 0.385 7.22 ;
      LAYER met1 ;
        RECT 0.155 5.945 0.615 6.115 ;
        RECT 0.155 5.915 0.445 6.145 ;
      LAYER mcon ;
        RECT 0.215 5.945 0.385 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 79.76 4.135 85.7 4.745 ;
        RECT 83.565 4.13 85.545 4.75 ;
        RECT 84.725 3.4 84.895 5.48 ;
        RECT 83.735 3.4 83.905 5.48 ;
        RECT 80.995 3.405 81.165 5.475 ;
        RECT 79.63 4.135 85.7 4.67 ;
        RECT 79.305 3.205 79.635 4.515 ;
        RECT -0.025 4.345 85.7 4.515 ;
        RECT 77.565 3.8 77.82 4.515 ;
        RECT 77 4.345 77.375 4.895 ;
        RECT 76.565 3.42 76.895 3.665 ;
        RECT 76.565 3.42 76.75 3.79 ;
        RECT 76.135 3.69 76.74 4.515 ;
        RECT 76.185 3.69 76.45 5.295 ;
        RECT 75.265 3.8 75.48 4.515 ;
        RECT 75.025 4.345 75.305 5.185 ;
        RECT 74.255 3.475 74.585 3.665 ;
        RECT 73.835 3.84 74.45 4.515 ;
        RECT 74.255 3.475 74.45 4.515 ;
        RECT 74.025 3.84 74.355 5.235 ;
        RECT 72.915 3.835 73.175 4.515 ;
        RECT 69.115 4.13 72.69 4.74 ;
        RECT 69.595 4.13 72.345 4.745 ;
        RECT 69.77 4.13 69.94 5.475 ;
        RECT 63.18 4.135 69.12 4.745 ;
        RECT 66.985 4.13 68.965 4.75 ;
        RECT 68.145 3.4 68.315 5.48 ;
        RECT 67.155 3.4 67.325 5.48 ;
        RECT 64.415 3.405 64.585 5.475 ;
        RECT 63.05 4.135 72.69 4.67 ;
        RECT 62.725 3.205 63.055 4.515 ;
        RECT 60.985 3.8 61.24 4.515 ;
        RECT 60.42 4.345 60.795 4.895 ;
        RECT 59.985 3.42 60.315 3.665 ;
        RECT 59.985 3.42 60.17 3.79 ;
        RECT 59.555 3.69 60.16 4.515 ;
        RECT 59.605 3.69 59.87 5.295 ;
        RECT 58.685 3.8 58.9 4.515 ;
        RECT 58.445 4.345 58.725 5.185 ;
        RECT 57.675 3.475 58.005 3.665 ;
        RECT 57.255 3.84 57.87 4.515 ;
        RECT 57.675 3.475 57.87 4.515 ;
        RECT 57.445 3.84 57.775 5.235 ;
        RECT 56.335 3.835 56.595 4.515 ;
        RECT 52.535 4.13 56.11 4.74 ;
        RECT 53.015 4.13 55.765 4.745 ;
        RECT 53.19 4.13 53.36 5.475 ;
        RECT 46.595 4.135 52.535 4.745 ;
        RECT 50.4 4.13 52.38 4.75 ;
        RECT 51.56 3.4 51.73 5.48 ;
        RECT 50.57 3.4 50.74 5.48 ;
        RECT 47.83 3.405 48 5.475 ;
        RECT 46.465 4.135 56.11 4.67 ;
        RECT 46.14 3.205 46.47 4.515 ;
        RECT 44.4 3.8 44.655 4.515 ;
        RECT 43.835 4.345 44.21 4.895 ;
        RECT 43.4 3.42 43.73 3.665 ;
        RECT 43.4 3.42 43.585 3.79 ;
        RECT 42.97 3.69 43.575 4.515 ;
        RECT 43.02 3.69 43.285 5.295 ;
        RECT 42.1 3.8 42.315 4.515 ;
        RECT 41.86 4.345 42.14 5.185 ;
        RECT 41.09 3.475 41.42 3.665 ;
        RECT 40.67 3.84 41.285 4.515 ;
        RECT 41.09 3.475 41.285 4.515 ;
        RECT 40.86 3.84 41.19 5.235 ;
        RECT 39.75 3.835 40.01 4.515 ;
        RECT 35.95 4.13 39.525 4.74 ;
        RECT 36.43 4.13 39.18 4.745 ;
        RECT 36.605 4.13 36.775 5.475 ;
        RECT 30.01 4.135 35.95 4.745 ;
        RECT 33.815 4.13 35.795 4.75 ;
        RECT 34.975 3.4 35.145 5.48 ;
        RECT 33.985 3.4 34.155 5.48 ;
        RECT 31.245 3.405 31.415 5.475 ;
        RECT 29.88 4.135 39.525 4.67 ;
        RECT 29.555 3.205 29.885 4.515 ;
        RECT 27.815 3.8 28.07 4.515 ;
        RECT 27.25 4.345 27.625 4.895 ;
        RECT 26.815 3.42 27.145 3.665 ;
        RECT 26.815 3.42 27 3.79 ;
        RECT 26.385 3.69 26.99 4.515 ;
        RECT 26.435 3.69 26.7 5.295 ;
        RECT 25.515 3.8 25.73 4.515 ;
        RECT 25.275 4.345 25.555 5.185 ;
        RECT 24.505 3.475 24.835 3.665 ;
        RECT 24.085 3.84 24.7 4.515 ;
        RECT 24.505 3.475 24.7 4.515 ;
        RECT 24.275 3.84 24.605 5.235 ;
        RECT 23.165 3.835 23.425 4.515 ;
        RECT 19.365 4.13 22.94 4.74 ;
        RECT 19.845 4.13 22.595 4.745 ;
        RECT 20.02 4.13 20.19 5.475 ;
        RECT 13.425 4.135 19.365 4.745 ;
        RECT 17.23 4.13 19.21 4.75 ;
        RECT 18.39 3.4 18.56 5.48 ;
        RECT 17.4 3.4 17.57 5.48 ;
        RECT 14.66 3.405 14.83 5.475 ;
        RECT 13.295 4.135 22.94 4.67 ;
        RECT 12.97 3.205 13.3 4.515 ;
        RECT 11.23 3.8 11.485 4.515 ;
        RECT 10.665 4.345 11.04 4.895 ;
        RECT 10.23 3.42 10.56 3.665 ;
        RECT 10.23 3.42 10.415 3.79 ;
        RECT 9.8 3.69 10.405 4.515 ;
        RECT 9.85 3.69 10.115 5.295 ;
        RECT 8.93 3.8 9.145 4.515 ;
        RECT 8.69 4.345 8.97 5.185 ;
        RECT 7.92 3.475 8.25 3.665 ;
        RECT 7.5 3.84 8.115 4.515 ;
        RECT 7.92 3.475 8.115 4.515 ;
        RECT 7.69 3.84 8.02 5.235 ;
        RECT 6.58 3.835 6.84 4.515 ;
        RECT -0.025 4.13 6.355 4.74 ;
        RECT 3.26 4.13 6.01 4.745 ;
        RECT 3.435 4.13 3.605 5.475 ;
        RECT -0.025 4.13 2.78 4.745 ;
        RECT 2.015 4.13 2.185 8.305 ;
        RECT 0.205 4.13 0.375 5.475 ;
      LAYER met1 ;
        RECT 79.76 4.15 85.7 4.745 ;
        RECT 80.22 4.135 85.7 4.745 ;
        RECT 83.565 4.13 85.545 4.75 ;
        RECT -0.025 4.19 85.7 4.67 ;
        RECT 79.63 4.15 85.7 4.67 ;
        RECT 69.115 4.13 72.69 4.74 ;
        RECT 69.595 4.13 72.345 4.745 ;
        RECT 63.18 4.15 69.12 4.745 ;
        RECT 63.64 4.135 72.69 4.74 ;
        RECT 66.985 4.13 68.965 4.75 ;
        RECT 63.05 4.15 72.69 4.67 ;
        RECT 52.535 4.13 56.11 4.74 ;
        RECT 53.015 4.13 55.765 4.745 ;
        RECT 46.595 4.15 52.535 4.745 ;
        RECT 47.055 4.135 56.11 4.74 ;
        RECT 50.4 4.13 52.38 4.75 ;
        RECT 46.465 4.15 56.11 4.67 ;
        RECT 35.95 4.13 39.525 4.74 ;
        RECT 36.43 4.13 39.18 4.745 ;
        RECT 30.01 4.15 35.95 4.745 ;
        RECT 30.47 4.135 39.525 4.74 ;
        RECT 33.815 4.13 35.795 4.75 ;
        RECT 29.88 4.15 39.525 4.67 ;
        RECT 19.365 4.13 22.94 4.74 ;
        RECT 19.845 4.13 22.595 4.745 ;
        RECT 13.425 4.15 19.365 4.745 ;
        RECT 13.885 4.135 22.94 4.74 ;
        RECT 17.23 4.13 19.21 4.75 ;
        RECT 13.295 4.15 22.94 4.67 ;
        RECT -0.025 4.13 6.355 4.74 ;
        RECT 3.26 4.13 6.01 4.745 ;
        RECT -0.025 4.13 2.78 4.745 ;
        RECT 1.955 6.655 2.245 6.885 ;
        RECT 1.785 6.685 2.245 6.855 ;
      LAYER mcon ;
        RECT 2.015 6.685 2.185 6.855 ;
        RECT 2.325 4.545 2.495 4.715 ;
        RECT 5.555 4.545 5.725 4.715 ;
        RECT 6.64 4.345 6.81 4.515 ;
        RECT 7.1 4.345 7.27 4.515 ;
        RECT 7.56 4.345 7.73 4.515 ;
        RECT 8.02 4.345 8.19 4.515 ;
        RECT 8.48 4.345 8.65 4.515 ;
        RECT 8.94 4.345 9.11 4.515 ;
        RECT 9.4 4.345 9.57 4.515 ;
        RECT 9.86 4.345 10.03 4.515 ;
        RECT 10.32 4.345 10.49 4.515 ;
        RECT 10.78 4.345 10.95 4.515 ;
        RECT 11.24 4.345 11.41 4.515 ;
        RECT 11.7 4.345 11.87 4.515 ;
        RECT 12.16 4.345 12.33 4.515 ;
        RECT 12.62 4.345 12.79 4.515 ;
        RECT 13.08 4.345 13.25 4.515 ;
        RECT 16.78 4.545 16.95 4.715 ;
        RECT 16.78 4.165 16.95 4.335 ;
        RECT 17.48 4.55 17.65 4.72 ;
        RECT 17.48 4.16 17.65 4.33 ;
        RECT 18.47 4.55 18.64 4.72 ;
        RECT 18.47 4.16 18.64 4.33 ;
        RECT 22.14 4.545 22.31 4.715 ;
        RECT 23.225 4.345 23.395 4.515 ;
        RECT 23.685 4.345 23.855 4.515 ;
        RECT 24.145 4.345 24.315 4.515 ;
        RECT 24.605 4.345 24.775 4.515 ;
        RECT 25.065 4.345 25.235 4.515 ;
        RECT 25.525 4.345 25.695 4.515 ;
        RECT 25.985 4.345 26.155 4.515 ;
        RECT 26.445 4.345 26.615 4.515 ;
        RECT 26.905 4.345 27.075 4.515 ;
        RECT 27.365 4.345 27.535 4.515 ;
        RECT 27.825 4.345 27.995 4.515 ;
        RECT 28.285 4.345 28.455 4.515 ;
        RECT 28.745 4.345 28.915 4.515 ;
        RECT 29.205 4.345 29.375 4.515 ;
        RECT 29.665 4.345 29.835 4.515 ;
        RECT 33.365 4.545 33.535 4.715 ;
        RECT 33.365 4.165 33.535 4.335 ;
        RECT 34.065 4.55 34.235 4.72 ;
        RECT 34.065 4.16 34.235 4.33 ;
        RECT 35.055 4.55 35.225 4.72 ;
        RECT 35.055 4.16 35.225 4.33 ;
        RECT 38.725 4.545 38.895 4.715 ;
        RECT 39.81 4.345 39.98 4.515 ;
        RECT 40.27 4.345 40.44 4.515 ;
        RECT 40.73 4.345 40.9 4.515 ;
        RECT 41.19 4.345 41.36 4.515 ;
        RECT 41.65 4.345 41.82 4.515 ;
        RECT 42.11 4.345 42.28 4.515 ;
        RECT 42.57 4.345 42.74 4.515 ;
        RECT 43.03 4.345 43.2 4.515 ;
        RECT 43.49 4.345 43.66 4.515 ;
        RECT 43.95 4.345 44.12 4.515 ;
        RECT 44.41 4.345 44.58 4.515 ;
        RECT 44.87 4.345 45.04 4.515 ;
        RECT 45.33 4.345 45.5 4.515 ;
        RECT 45.79 4.345 45.96 4.515 ;
        RECT 46.25 4.345 46.42 4.515 ;
        RECT 49.95 4.545 50.12 4.715 ;
        RECT 49.95 4.165 50.12 4.335 ;
        RECT 50.65 4.55 50.82 4.72 ;
        RECT 50.65 4.16 50.82 4.33 ;
        RECT 51.64 4.55 51.81 4.72 ;
        RECT 51.64 4.16 51.81 4.33 ;
        RECT 55.31 4.545 55.48 4.715 ;
        RECT 56.395 4.345 56.565 4.515 ;
        RECT 56.855 4.345 57.025 4.515 ;
        RECT 57.315 4.345 57.485 4.515 ;
        RECT 57.775 4.345 57.945 4.515 ;
        RECT 58.235 4.345 58.405 4.515 ;
        RECT 58.695 4.345 58.865 4.515 ;
        RECT 59.155 4.345 59.325 4.515 ;
        RECT 59.615 4.345 59.785 4.515 ;
        RECT 60.075 4.345 60.245 4.515 ;
        RECT 60.535 4.345 60.705 4.515 ;
        RECT 60.995 4.345 61.165 4.515 ;
        RECT 61.455 4.345 61.625 4.515 ;
        RECT 61.915 4.345 62.085 4.515 ;
        RECT 62.375 4.345 62.545 4.515 ;
        RECT 62.835 4.345 63.005 4.515 ;
        RECT 66.535 4.545 66.705 4.715 ;
        RECT 66.535 4.165 66.705 4.335 ;
        RECT 67.235 4.55 67.405 4.72 ;
        RECT 67.235 4.16 67.405 4.33 ;
        RECT 68.225 4.55 68.395 4.72 ;
        RECT 68.225 4.16 68.395 4.33 ;
        RECT 71.89 4.545 72.06 4.715 ;
        RECT 72.975 4.345 73.145 4.515 ;
        RECT 73.435 4.345 73.605 4.515 ;
        RECT 73.895 4.345 74.065 4.515 ;
        RECT 74.355 4.345 74.525 4.515 ;
        RECT 74.815 4.345 74.985 4.515 ;
        RECT 75.275 4.345 75.445 4.515 ;
        RECT 75.735 4.345 75.905 4.515 ;
        RECT 76.195 4.345 76.365 4.515 ;
        RECT 76.655 4.345 76.825 4.515 ;
        RECT 77.115 4.345 77.285 4.515 ;
        RECT 77.575 4.345 77.745 4.515 ;
        RECT 78.035 4.345 78.205 4.515 ;
        RECT 78.495 4.345 78.665 4.515 ;
        RECT 78.955 4.345 79.125 4.515 ;
        RECT 79.415 4.345 79.585 4.515 ;
        RECT 83.115 4.545 83.285 4.715 ;
        RECT 83.115 4.165 83.285 4.335 ;
        RECT 83.815 4.55 83.985 4.72 ;
        RECT 83.815 4.16 83.985 4.33 ;
        RECT 84.805 4.55 84.975 4.72 ;
        RECT 84.805 4.16 84.975 4.33 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 75.205 6.475 75.535 6.805 ;
        RECT 75.175 6.49 75.475 6.905 ;
        RECT 74.735 6.49 75.535 6.79 ;
        RECT 58.625 6.475 58.955 6.805 ;
        RECT 58.595 6.49 58.895 6.905 ;
        RECT 58.155 6.49 58.955 6.79 ;
        RECT 42.04 6.475 42.37 6.805 ;
        RECT 42.01 6.49 42.31 6.905 ;
        RECT 41.57 6.49 42.37 6.79 ;
        RECT 25.455 6.475 25.785 6.805 ;
        RECT 25.425 6.49 25.725 6.905 ;
        RECT 24.985 6.49 25.785 6.79 ;
        RECT 8.87 6.475 9.2 6.805 ;
        RECT 8.84 6.49 9.14 6.905 ;
        RECT 8.4 6.49 9.2 6.79 ;
      LAYER li1 ;
        RECT -0.025 8.57 85.73 8.88 ;
        RECT 84.725 7.95 84.895 8.88 ;
        RECT 83.735 7.95 83.905 8.88 ;
        RECT 80.995 7.945 81.165 8.88 ;
        RECT 72.535 7.18 79.735 8.88 ;
        RECT 72.83 7.065 79.73 8.88 ;
        RECT 78.265 6.555 78.715 8.88 ;
        RECT 76.175 6.665 76.505 8.88 ;
        RECT 74.105 6.605 74.355 8.88 ;
        RECT 69.77 7.945 69.94 8.88 ;
        RECT 68.145 7.95 68.315 8.88 ;
        RECT 67.155 7.95 67.325 8.88 ;
        RECT 64.415 7.945 64.585 8.88 ;
        RECT 55.955 7.18 63.155 8.88 ;
        RECT 56.25 7.065 63.15 8.88 ;
        RECT 61.685 6.555 62.135 8.88 ;
        RECT 59.595 6.665 59.925 8.88 ;
        RECT 57.525 6.605 57.775 8.88 ;
        RECT 53.19 7.945 53.36 8.88 ;
        RECT 51.56 7.95 51.73 8.88 ;
        RECT 50.57 7.95 50.74 8.88 ;
        RECT 47.83 7.945 48 8.88 ;
        RECT 39.37 7.18 46.57 8.88 ;
        RECT 39.665 7.065 46.565 8.88 ;
        RECT 45.1 6.555 45.55 8.88 ;
        RECT 43.01 6.665 43.34 8.88 ;
        RECT 40.94 6.605 41.19 8.88 ;
        RECT 36.605 7.945 36.775 8.88 ;
        RECT 34.975 7.95 35.145 8.88 ;
        RECT 33.985 7.95 34.155 8.88 ;
        RECT 31.245 7.945 31.415 8.88 ;
        RECT 22.785 7.18 29.985 8.88 ;
        RECT 23.08 7.065 29.98 8.88 ;
        RECT 28.515 6.555 28.965 8.88 ;
        RECT 26.425 6.665 26.755 8.88 ;
        RECT 24.355 6.605 24.605 8.88 ;
        RECT 20.02 7.945 20.19 8.88 ;
        RECT 18.39 7.95 18.56 8.88 ;
        RECT 17.4 7.95 17.57 8.88 ;
        RECT 14.66 7.945 14.83 8.88 ;
        RECT 6.2 7.18 13.4 8.88 ;
        RECT 6.495 7.065 13.395 8.88 ;
        RECT 11.93 6.555 12.38 8.88 ;
        RECT 9.84 6.665 10.17 8.88 ;
        RECT 7.77 6.605 8.02 8.88 ;
        RECT 3.435 7.945 3.605 8.88 ;
        RECT 0.205 7.945 0.375 8.88 ;
        RECT -0.025 0 85.705 0.31 ;
        RECT 84.725 0 84.895 0.93 ;
        RECT 83.735 0 83.905 0.93 ;
        RECT 80.995 0 81.165 0.935 ;
        RECT 72.83 0 79.92 1.795 ;
        RECT 79.365 0 79.635 2.605 ;
        RECT 78.455 0 78.695 2.605 ;
        RECT 77.585 0 77.835 2.335 ;
        RECT 75.205 0 75.535 2.255 ;
        RECT 72.915 0 73.175 2.615 ;
        RECT 72.575 0 79.92 1.655 ;
        RECT 68.145 0 68.315 0.93 ;
        RECT 67.155 0 67.325 0.93 ;
        RECT 64.415 0 64.585 0.935 ;
        RECT 56.25 0 63.34 1.795 ;
        RECT 62.785 0 63.055 2.605 ;
        RECT 61.875 0 62.115 2.605 ;
        RECT 61.005 0 61.255 2.335 ;
        RECT 58.625 0 58.955 2.255 ;
        RECT 56.335 0 56.595 2.615 ;
        RECT 55.995 0 63.34 1.655 ;
        RECT 51.56 0 51.73 0.93 ;
        RECT 50.57 0 50.74 0.93 ;
        RECT 47.83 0 48 0.935 ;
        RECT 39.665 0 46.755 1.795 ;
        RECT 46.2 0 46.47 2.605 ;
        RECT 45.29 0 45.53 2.605 ;
        RECT 44.42 0 44.67 2.335 ;
        RECT 42.04 0 42.37 2.255 ;
        RECT 39.75 0 40.01 2.615 ;
        RECT 39.41 0 46.755 1.655 ;
        RECT 34.975 0 35.145 0.93 ;
        RECT 33.985 0 34.155 0.93 ;
        RECT 31.245 0 31.415 0.935 ;
        RECT 23.08 0 30.17 1.795 ;
        RECT 29.615 0 29.885 2.605 ;
        RECT 28.705 0 28.945 2.605 ;
        RECT 27.835 0 28.085 2.335 ;
        RECT 25.455 0 25.785 2.255 ;
        RECT 23.165 0 23.425 2.615 ;
        RECT 22.825 0 30.17 1.655 ;
        RECT 18.39 0 18.56 0.93 ;
        RECT 17.4 0 17.57 0.93 ;
        RECT 14.66 0 14.83 0.935 ;
        RECT 6.495 0 13.585 1.795 ;
        RECT 13.03 0 13.3 2.605 ;
        RECT 12.12 0 12.36 2.605 ;
        RECT 11.25 0 11.5 2.335 ;
        RECT 8.87 0 9.2 2.255 ;
        RECT 6.58 0 6.84 2.615 ;
        RECT 6.24 0 13.585 1.655 ;
        RECT 76.475 5.825 76.8 6.155 ;
        RECT 74.255 5.825 74.595 6.075 ;
        RECT 70.775 6.075 70.945 8.025 ;
        RECT 70.72 7.855 70.89 8.305 ;
        RECT 70.72 5.015 70.89 6.245 ;
        RECT 59.895 5.825 60.22 6.155 ;
        RECT 57.675 5.825 58.015 6.075 ;
        RECT 54.195 6.075 54.365 8.025 ;
        RECT 54.14 7.855 54.31 8.305 ;
        RECT 54.14 5.015 54.31 6.245 ;
        RECT 43.31 5.825 43.635 6.155 ;
        RECT 41.09 5.825 41.43 6.075 ;
        RECT 37.61 6.075 37.78 8.025 ;
        RECT 37.555 7.855 37.725 8.305 ;
        RECT 37.555 5.015 37.725 6.245 ;
        RECT 26.725 5.825 27.05 6.155 ;
        RECT 24.505 5.825 24.845 6.075 ;
        RECT 21.025 6.075 21.195 8.025 ;
        RECT 20.97 7.855 21.14 8.305 ;
        RECT 20.97 5.015 21.14 6.245 ;
        RECT 10.14 5.825 10.465 6.155 ;
        RECT 7.92 5.825 8.26 6.075 ;
        RECT 4.44 6.075 4.61 8.025 ;
        RECT 4.385 7.855 4.555 8.305 ;
        RECT 4.385 5.015 4.555 6.245 ;
      LAYER met2 ;
        RECT 75.23 6.455 75.51 6.825 ;
        RECT 58.65 6.455 58.93 6.825 ;
        RECT 42.065 6.455 42.345 6.825 ;
        RECT 25.48 6.455 25.76 6.825 ;
        RECT 8.895 6.455 9.175 6.825 ;
      LAYER met1 ;
        RECT -0.025 8.57 85.73 8.88 ;
        RECT 72.535 7.18 79.735 8.88 ;
        RECT 72.83 6.91 79.73 8.88 ;
        RECT 76.425 5.845 76.715 6.075 ;
        RECT 74.29 6.57 76.64 6.71 ;
        RECT 76.5 5.845 76.64 6.71 ;
        RECT 75.22 6.51 75.54 6.77 ;
        RECT 75.255 6.51 75.51 8.88 ;
        RECT 74.215 5.845 74.505 6.075 ;
        RECT 74.29 5.845 74.43 6.71 ;
        RECT 70.715 6.285 71.005 6.515 ;
        RECT 70.555 6.315 70.725 8.88 ;
        RECT 70.545 6.315 71.005 6.485 ;
        RECT 55.955 7.18 63.155 8.88 ;
        RECT 56.25 6.91 63.15 8.88 ;
        RECT 59.845 5.845 60.135 6.075 ;
        RECT 57.71 6.57 60.06 6.71 ;
        RECT 59.92 5.845 60.06 6.71 ;
        RECT 58.64 6.51 58.96 6.77 ;
        RECT 58.675 6.51 58.93 8.88 ;
        RECT 57.635 5.845 57.925 6.075 ;
        RECT 57.71 5.845 57.85 6.71 ;
        RECT 54.135 6.285 54.425 6.515 ;
        RECT 53.975 6.315 54.145 8.88 ;
        RECT 53.965 6.315 54.425 6.485 ;
        RECT 39.37 7.18 46.57 8.88 ;
        RECT 39.665 6.91 46.565 8.88 ;
        RECT 43.26 5.845 43.55 6.075 ;
        RECT 41.125 6.57 43.475 6.71 ;
        RECT 43.335 5.845 43.475 6.71 ;
        RECT 42.055 6.51 42.375 6.77 ;
        RECT 42.09 6.51 42.345 8.88 ;
        RECT 41.05 5.845 41.34 6.075 ;
        RECT 41.125 5.845 41.265 6.71 ;
        RECT 37.55 6.285 37.84 6.515 ;
        RECT 37.39 6.315 37.56 8.88 ;
        RECT 37.38 6.315 37.84 6.485 ;
        RECT 22.785 7.18 29.985 8.88 ;
        RECT 23.08 6.91 29.98 8.88 ;
        RECT 26.675 5.845 26.965 6.075 ;
        RECT 24.54 6.57 26.89 6.71 ;
        RECT 26.75 5.845 26.89 6.71 ;
        RECT 25.47 6.51 25.79 6.77 ;
        RECT 25.505 6.51 25.76 8.88 ;
        RECT 24.465 5.845 24.755 6.075 ;
        RECT 24.54 5.845 24.68 6.71 ;
        RECT 20.965 6.285 21.255 6.515 ;
        RECT 20.805 6.315 20.975 8.88 ;
        RECT 20.795 6.315 21.255 6.485 ;
        RECT 6.2 7.18 13.4 8.88 ;
        RECT 6.495 6.91 13.395 8.88 ;
        RECT 10.09 5.845 10.38 6.075 ;
        RECT 7.955 6.57 10.305 6.71 ;
        RECT 10.165 5.845 10.305 6.71 ;
        RECT 8.885 6.51 9.205 6.77 ;
        RECT 8.92 6.51 9.175 8.88 ;
        RECT 7.88 5.845 8.17 6.075 ;
        RECT 7.955 5.845 8.095 6.71 ;
        RECT 4.38 6.285 4.67 6.515 ;
        RECT 4.22 6.315 4.39 8.88 ;
        RECT 4.21 6.315 4.67 6.485 ;
        RECT -0.025 0 85.705 0.31 ;
        RECT 72.83 0 79.92 1.795 ;
        RECT 72.83 0 79.73 1.95 ;
        RECT 72.575 0 79.92 1.655 ;
        RECT 56.25 0 63.34 1.795 ;
        RECT 56.25 0 63.15 1.95 ;
        RECT 55.995 0 63.34 1.655 ;
        RECT 39.665 0 46.755 1.795 ;
        RECT 39.665 0 46.565 1.95 ;
        RECT 39.41 0 46.755 1.655 ;
        RECT 23.08 0 30.17 1.795 ;
        RECT 23.08 0 29.98 1.95 ;
        RECT 22.825 0 30.17 1.655 ;
        RECT 6.495 0 13.585 1.795 ;
        RECT 6.495 0 13.395 1.95 ;
        RECT 6.24 0 13.585 1.655 ;
      LAYER via2 ;
        RECT 8.935 6.54 9.135 6.74 ;
        RECT 25.52 6.54 25.72 6.74 ;
        RECT 42.105 6.54 42.305 6.74 ;
        RECT 58.69 6.54 58.89 6.74 ;
        RECT 75.27 6.54 75.47 6.74 ;
      LAYER via1 ;
        RECT 8.97 6.565 9.12 6.715 ;
        RECT 25.555 6.565 25.705 6.715 ;
        RECT 42.14 6.565 42.29 6.715 ;
        RECT 58.725 6.565 58.875 6.715 ;
        RECT 75.305 6.565 75.455 6.715 ;
      LAYER mcon ;
        RECT 0.285 8.605 0.455 8.775 ;
        RECT 0.965 8.605 1.135 8.775 ;
        RECT 1.645 8.605 1.815 8.775 ;
        RECT 2.325 8.605 2.495 8.775 ;
        RECT 3.515 8.605 3.685 8.775 ;
        RECT 4.195 8.605 4.365 8.775 ;
        RECT 4.44 6.315 4.61 6.485 ;
        RECT 4.875 8.605 5.045 8.775 ;
        RECT 5.555 8.605 5.725 8.775 ;
        RECT 6.64 7.065 6.81 7.235 ;
        RECT 6.64 1.625 6.81 1.795 ;
        RECT 7.1 7.065 7.27 7.235 ;
        RECT 7.1 1.625 7.27 1.795 ;
        RECT 7.56 7.065 7.73 7.235 ;
        RECT 7.56 1.625 7.73 1.795 ;
        RECT 7.94 5.875 8.11 6.045 ;
        RECT 8.02 7.065 8.19 7.235 ;
        RECT 8.02 1.625 8.19 1.795 ;
        RECT 8.48 7.065 8.65 7.235 ;
        RECT 8.48 1.625 8.65 1.795 ;
        RECT 8.94 7.065 9.11 7.235 ;
        RECT 8.94 1.625 9.11 1.795 ;
        RECT 9.4 7.065 9.57 7.235 ;
        RECT 9.4 1.625 9.57 1.795 ;
        RECT 9.86 7.065 10.03 7.235 ;
        RECT 9.86 1.625 10.03 1.795 ;
        RECT 10.15 5.875 10.32 6.045 ;
        RECT 10.32 7.065 10.49 7.235 ;
        RECT 10.32 1.625 10.49 1.795 ;
        RECT 10.78 7.065 10.95 7.235 ;
        RECT 10.78 1.625 10.95 1.795 ;
        RECT 11.24 7.065 11.41 7.235 ;
        RECT 11.24 1.625 11.41 1.795 ;
        RECT 11.7 7.065 11.87 7.235 ;
        RECT 11.7 1.625 11.87 1.795 ;
        RECT 12.16 7.065 12.33 7.235 ;
        RECT 12.16 1.625 12.33 1.795 ;
        RECT 12.62 7.065 12.79 7.235 ;
        RECT 12.62 1.625 12.79 1.795 ;
        RECT 13.08 7.065 13.25 7.235 ;
        RECT 13.08 1.625 13.25 1.795 ;
        RECT 14.74 8.605 14.91 8.775 ;
        RECT 14.74 0.105 14.91 0.275 ;
        RECT 15.42 8.605 15.59 8.775 ;
        RECT 15.42 0.105 15.59 0.275 ;
        RECT 16.1 8.605 16.27 8.775 ;
        RECT 16.1 0.105 16.27 0.275 ;
        RECT 16.78 8.605 16.95 8.775 ;
        RECT 16.78 0.105 16.95 0.275 ;
        RECT 17.48 8.61 17.65 8.78 ;
        RECT 17.48 0.1 17.65 0.27 ;
        RECT 18.47 8.61 18.64 8.78 ;
        RECT 18.47 0.1 18.64 0.27 ;
        RECT 20.1 8.605 20.27 8.775 ;
        RECT 20.78 8.605 20.95 8.775 ;
        RECT 21.025 6.315 21.195 6.485 ;
        RECT 21.46 8.605 21.63 8.775 ;
        RECT 22.14 8.605 22.31 8.775 ;
        RECT 23.225 7.065 23.395 7.235 ;
        RECT 23.225 1.625 23.395 1.795 ;
        RECT 23.685 7.065 23.855 7.235 ;
        RECT 23.685 1.625 23.855 1.795 ;
        RECT 24.145 7.065 24.315 7.235 ;
        RECT 24.145 1.625 24.315 1.795 ;
        RECT 24.525 5.875 24.695 6.045 ;
        RECT 24.605 7.065 24.775 7.235 ;
        RECT 24.605 1.625 24.775 1.795 ;
        RECT 25.065 7.065 25.235 7.235 ;
        RECT 25.065 1.625 25.235 1.795 ;
        RECT 25.525 7.065 25.695 7.235 ;
        RECT 25.525 1.625 25.695 1.795 ;
        RECT 25.985 7.065 26.155 7.235 ;
        RECT 25.985 1.625 26.155 1.795 ;
        RECT 26.445 7.065 26.615 7.235 ;
        RECT 26.445 1.625 26.615 1.795 ;
        RECT 26.735 5.875 26.905 6.045 ;
        RECT 26.905 7.065 27.075 7.235 ;
        RECT 26.905 1.625 27.075 1.795 ;
        RECT 27.365 7.065 27.535 7.235 ;
        RECT 27.365 1.625 27.535 1.795 ;
        RECT 27.825 7.065 27.995 7.235 ;
        RECT 27.825 1.625 27.995 1.795 ;
        RECT 28.285 7.065 28.455 7.235 ;
        RECT 28.285 1.625 28.455 1.795 ;
        RECT 28.745 7.065 28.915 7.235 ;
        RECT 28.745 1.625 28.915 1.795 ;
        RECT 29.205 7.065 29.375 7.235 ;
        RECT 29.205 1.625 29.375 1.795 ;
        RECT 29.665 7.065 29.835 7.235 ;
        RECT 29.665 1.625 29.835 1.795 ;
        RECT 31.325 8.605 31.495 8.775 ;
        RECT 31.325 0.105 31.495 0.275 ;
        RECT 32.005 8.605 32.175 8.775 ;
        RECT 32.005 0.105 32.175 0.275 ;
        RECT 32.685 8.605 32.855 8.775 ;
        RECT 32.685 0.105 32.855 0.275 ;
        RECT 33.365 8.605 33.535 8.775 ;
        RECT 33.365 0.105 33.535 0.275 ;
        RECT 34.065 8.61 34.235 8.78 ;
        RECT 34.065 0.1 34.235 0.27 ;
        RECT 35.055 8.61 35.225 8.78 ;
        RECT 35.055 0.1 35.225 0.27 ;
        RECT 36.685 8.605 36.855 8.775 ;
        RECT 37.365 8.605 37.535 8.775 ;
        RECT 37.61 6.315 37.78 6.485 ;
        RECT 38.045 8.605 38.215 8.775 ;
        RECT 38.725 8.605 38.895 8.775 ;
        RECT 39.81 7.065 39.98 7.235 ;
        RECT 39.81 1.625 39.98 1.795 ;
        RECT 40.27 7.065 40.44 7.235 ;
        RECT 40.27 1.625 40.44 1.795 ;
        RECT 40.73 7.065 40.9 7.235 ;
        RECT 40.73 1.625 40.9 1.795 ;
        RECT 41.11 5.875 41.28 6.045 ;
        RECT 41.19 7.065 41.36 7.235 ;
        RECT 41.19 1.625 41.36 1.795 ;
        RECT 41.65 7.065 41.82 7.235 ;
        RECT 41.65 1.625 41.82 1.795 ;
        RECT 42.11 7.065 42.28 7.235 ;
        RECT 42.11 1.625 42.28 1.795 ;
        RECT 42.57 7.065 42.74 7.235 ;
        RECT 42.57 1.625 42.74 1.795 ;
        RECT 43.03 7.065 43.2 7.235 ;
        RECT 43.03 1.625 43.2 1.795 ;
        RECT 43.32 5.875 43.49 6.045 ;
        RECT 43.49 7.065 43.66 7.235 ;
        RECT 43.49 1.625 43.66 1.795 ;
        RECT 43.95 7.065 44.12 7.235 ;
        RECT 43.95 1.625 44.12 1.795 ;
        RECT 44.41 7.065 44.58 7.235 ;
        RECT 44.41 1.625 44.58 1.795 ;
        RECT 44.87 7.065 45.04 7.235 ;
        RECT 44.87 1.625 45.04 1.795 ;
        RECT 45.33 7.065 45.5 7.235 ;
        RECT 45.33 1.625 45.5 1.795 ;
        RECT 45.79 7.065 45.96 7.235 ;
        RECT 45.79 1.625 45.96 1.795 ;
        RECT 46.25 7.065 46.42 7.235 ;
        RECT 46.25 1.625 46.42 1.795 ;
        RECT 47.91 8.605 48.08 8.775 ;
        RECT 47.91 0.105 48.08 0.275 ;
        RECT 48.59 8.605 48.76 8.775 ;
        RECT 48.59 0.105 48.76 0.275 ;
        RECT 49.27 8.605 49.44 8.775 ;
        RECT 49.27 0.105 49.44 0.275 ;
        RECT 49.95 8.605 50.12 8.775 ;
        RECT 49.95 0.105 50.12 0.275 ;
        RECT 50.65 8.61 50.82 8.78 ;
        RECT 50.65 0.1 50.82 0.27 ;
        RECT 51.64 8.61 51.81 8.78 ;
        RECT 51.64 0.1 51.81 0.27 ;
        RECT 53.27 8.605 53.44 8.775 ;
        RECT 53.95 8.605 54.12 8.775 ;
        RECT 54.195 6.315 54.365 6.485 ;
        RECT 54.63 8.605 54.8 8.775 ;
        RECT 55.31 8.605 55.48 8.775 ;
        RECT 56.395 7.065 56.565 7.235 ;
        RECT 56.395 1.625 56.565 1.795 ;
        RECT 56.855 7.065 57.025 7.235 ;
        RECT 56.855 1.625 57.025 1.795 ;
        RECT 57.315 7.065 57.485 7.235 ;
        RECT 57.315 1.625 57.485 1.795 ;
        RECT 57.695 5.875 57.865 6.045 ;
        RECT 57.775 7.065 57.945 7.235 ;
        RECT 57.775 1.625 57.945 1.795 ;
        RECT 58.235 7.065 58.405 7.235 ;
        RECT 58.235 1.625 58.405 1.795 ;
        RECT 58.695 7.065 58.865 7.235 ;
        RECT 58.695 1.625 58.865 1.795 ;
        RECT 59.155 7.065 59.325 7.235 ;
        RECT 59.155 1.625 59.325 1.795 ;
        RECT 59.615 7.065 59.785 7.235 ;
        RECT 59.615 1.625 59.785 1.795 ;
        RECT 59.905 5.875 60.075 6.045 ;
        RECT 60.075 7.065 60.245 7.235 ;
        RECT 60.075 1.625 60.245 1.795 ;
        RECT 60.535 7.065 60.705 7.235 ;
        RECT 60.535 1.625 60.705 1.795 ;
        RECT 60.995 7.065 61.165 7.235 ;
        RECT 60.995 1.625 61.165 1.795 ;
        RECT 61.455 7.065 61.625 7.235 ;
        RECT 61.455 1.625 61.625 1.795 ;
        RECT 61.915 7.065 62.085 7.235 ;
        RECT 61.915 1.625 62.085 1.795 ;
        RECT 62.375 7.065 62.545 7.235 ;
        RECT 62.375 1.625 62.545 1.795 ;
        RECT 62.835 7.065 63.005 7.235 ;
        RECT 62.835 1.625 63.005 1.795 ;
        RECT 64.495 8.605 64.665 8.775 ;
        RECT 64.495 0.105 64.665 0.275 ;
        RECT 65.175 8.605 65.345 8.775 ;
        RECT 65.175 0.105 65.345 0.275 ;
        RECT 65.855 8.605 66.025 8.775 ;
        RECT 65.855 0.105 66.025 0.275 ;
        RECT 66.535 8.605 66.705 8.775 ;
        RECT 66.535 0.105 66.705 0.275 ;
        RECT 67.235 8.61 67.405 8.78 ;
        RECT 67.235 0.1 67.405 0.27 ;
        RECT 68.225 8.61 68.395 8.78 ;
        RECT 68.225 0.1 68.395 0.27 ;
        RECT 69.85 8.605 70.02 8.775 ;
        RECT 70.53 8.605 70.7 8.775 ;
        RECT 70.775 6.315 70.945 6.485 ;
        RECT 71.21 8.605 71.38 8.775 ;
        RECT 71.89 8.605 72.06 8.775 ;
        RECT 72.975 7.065 73.145 7.235 ;
        RECT 72.975 1.625 73.145 1.795 ;
        RECT 73.435 7.065 73.605 7.235 ;
        RECT 73.435 1.625 73.605 1.795 ;
        RECT 73.895 7.065 74.065 7.235 ;
        RECT 73.895 1.625 74.065 1.795 ;
        RECT 74.275 5.875 74.445 6.045 ;
        RECT 74.355 7.065 74.525 7.235 ;
        RECT 74.355 1.625 74.525 1.795 ;
        RECT 74.815 7.065 74.985 7.235 ;
        RECT 74.815 1.625 74.985 1.795 ;
        RECT 75.275 7.065 75.445 7.235 ;
        RECT 75.275 1.625 75.445 1.795 ;
        RECT 75.735 7.065 75.905 7.235 ;
        RECT 75.735 1.625 75.905 1.795 ;
        RECT 76.195 7.065 76.365 7.235 ;
        RECT 76.195 1.625 76.365 1.795 ;
        RECT 76.485 5.875 76.655 6.045 ;
        RECT 76.655 7.065 76.825 7.235 ;
        RECT 76.655 1.625 76.825 1.795 ;
        RECT 77.115 7.065 77.285 7.235 ;
        RECT 77.115 1.625 77.285 1.795 ;
        RECT 77.575 7.065 77.745 7.235 ;
        RECT 77.575 1.625 77.745 1.795 ;
        RECT 78.035 7.065 78.205 7.235 ;
        RECT 78.035 1.625 78.205 1.795 ;
        RECT 78.495 7.065 78.665 7.235 ;
        RECT 78.495 1.625 78.665 1.795 ;
        RECT 78.955 7.065 79.125 7.235 ;
        RECT 78.955 1.625 79.125 1.795 ;
        RECT 79.415 7.065 79.585 7.235 ;
        RECT 79.415 1.625 79.585 1.795 ;
        RECT 81.075 8.605 81.245 8.775 ;
        RECT 81.075 0.105 81.245 0.275 ;
        RECT 81.755 8.605 81.925 8.775 ;
        RECT 81.755 0.105 81.925 0.275 ;
        RECT 82.435 8.605 82.605 8.775 ;
        RECT 82.435 0.105 82.605 0.275 ;
        RECT 83.115 8.605 83.285 8.775 ;
        RECT 83.115 0.105 83.285 0.275 ;
        RECT 83.815 8.61 83.985 8.78 ;
        RECT 83.815 0.1 83.985 0.27 ;
        RECT 84.805 8.61 84.975 8.78 ;
        RECT 84.805 0.1 84.975 0.27 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 77.605 2.735 77.935 3.065 ;
      RECT 77.605 2.75 78.405 3.05 ;
      RECT 77.605 2.73 77.925 3.065 ;
      RECT 71.925 7.97 76.205 8.27 ;
      RECT 75.9 5.795 76.2 8.27 ;
      RECT 71.925 7.03 72.225 8.27 ;
      RECT 71.05 6.995 71.42 7.365 ;
      RECT 71.05 7.03 72.225 7.33 ;
      RECT 76.925 5.795 77.255 6.125 ;
      RECT 75.275 5.795 76.21 6.125 ;
      RECT 75.275 5.81 77.725 6.11 ;
      RECT 75.275 5.795 77.255 6.11 ;
      RECT 76.93 5.79 77.23 6.125 ;
      RECT 75.275 3.765 75.605 6.125 ;
      RECT 75.275 3.765 77.57 4.095 ;
      RECT 75.275 3.765 77.935 4.085 ;
      RECT 77.605 3.755 77.935 4.085 ;
      RECT 75.275 3.77 78.405 4.07 ;
      RECT 77.61 3.705 77.91 4.085 ;
      RECT 76.905 3.075 77.235 3.405 ;
      RECT 76.435 3.09 77.235 3.39 ;
      RECT 76.93 3.06 77.23 3.405 ;
      RECT 76.245 4.775 76.575 5.105 ;
      RECT 76.245 4.79 77.045 5.09 ;
      RECT 75.565 2.39 75.895 2.72 ;
      RECT 75.095 2.41 75.455 2.71 ;
      RECT 75.455 2.405 75.895 2.705 ;
      RECT 61.025 2.735 61.355 3.065 ;
      RECT 61.025 2.75 61.825 3.05 ;
      RECT 61.025 2.73 61.345 3.065 ;
      RECT 55.345 7.97 59.625 8.27 ;
      RECT 59.32 5.795 59.62 8.27 ;
      RECT 55.345 7.03 55.645 8.27 ;
      RECT 54.47 6.995 54.84 7.365 ;
      RECT 54.47 7.03 55.645 7.33 ;
      RECT 60.345 5.795 60.675 6.125 ;
      RECT 58.695 5.795 59.63 6.125 ;
      RECT 58.695 5.81 61.145 6.11 ;
      RECT 58.695 5.795 60.675 6.11 ;
      RECT 60.35 5.79 60.65 6.125 ;
      RECT 58.695 3.765 59.025 6.125 ;
      RECT 58.695 3.765 60.99 4.095 ;
      RECT 58.695 3.765 61.355 4.085 ;
      RECT 61.025 3.755 61.355 4.085 ;
      RECT 58.695 3.77 61.825 4.07 ;
      RECT 61.03 3.705 61.33 4.085 ;
      RECT 60.325 3.075 60.655 3.405 ;
      RECT 59.855 3.09 60.655 3.39 ;
      RECT 60.35 3.06 60.65 3.405 ;
      RECT 59.665 4.775 59.995 5.105 ;
      RECT 59.665 4.79 60.465 5.09 ;
      RECT 58.985 2.39 59.315 2.72 ;
      RECT 58.515 2.41 58.875 2.71 ;
      RECT 58.875 2.405 59.315 2.705 ;
      RECT 44.44 2.735 44.77 3.065 ;
      RECT 44.44 2.75 45.24 3.05 ;
      RECT 44.44 2.73 44.76 3.065 ;
      RECT 38.76 7.97 43.04 8.27 ;
      RECT 42.735 5.795 43.035 8.27 ;
      RECT 38.76 7.03 39.06 8.27 ;
      RECT 37.885 6.995 38.255 7.365 ;
      RECT 37.885 7.03 39.06 7.33 ;
      RECT 43.76 5.795 44.09 6.125 ;
      RECT 42.11 5.795 43.045 6.125 ;
      RECT 42.11 5.81 44.56 6.11 ;
      RECT 42.11 5.795 44.09 6.11 ;
      RECT 43.765 5.79 44.065 6.125 ;
      RECT 42.11 3.765 42.44 6.125 ;
      RECT 42.11 3.765 44.405 4.095 ;
      RECT 42.11 3.765 44.77 4.085 ;
      RECT 44.44 3.755 44.77 4.085 ;
      RECT 42.11 3.77 45.24 4.07 ;
      RECT 44.445 3.705 44.745 4.085 ;
      RECT 43.74 3.075 44.07 3.405 ;
      RECT 43.27 3.09 44.07 3.39 ;
      RECT 43.765 3.06 44.065 3.405 ;
      RECT 43.08 4.775 43.41 5.105 ;
      RECT 43.08 4.79 43.88 5.09 ;
      RECT 42.4 2.39 42.73 2.72 ;
      RECT 41.93 2.41 42.29 2.71 ;
      RECT 42.29 2.405 42.73 2.705 ;
      RECT 27.855 2.735 28.185 3.065 ;
      RECT 27.855 2.75 28.655 3.05 ;
      RECT 27.855 2.73 28.175 3.065 ;
      RECT 22.175 7.97 26.455 8.27 ;
      RECT 26.15 5.795 26.45 8.27 ;
      RECT 22.175 7.03 22.475 8.27 ;
      RECT 21.3 6.995 21.67 7.365 ;
      RECT 21.3 7.03 22.475 7.33 ;
      RECT 27.175 5.795 27.505 6.125 ;
      RECT 25.525 5.795 26.46 6.125 ;
      RECT 25.525 5.81 27.975 6.11 ;
      RECT 25.525 5.795 27.505 6.11 ;
      RECT 27.18 5.79 27.48 6.125 ;
      RECT 25.525 3.765 25.855 6.125 ;
      RECT 25.525 3.765 27.82 4.095 ;
      RECT 25.525 3.765 28.185 4.085 ;
      RECT 27.855 3.755 28.185 4.085 ;
      RECT 25.525 3.77 28.655 4.07 ;
      RECT 27.86 3.705 28.16 4.085 ;
      RECT 27.155 3.075 27.485 3.405 ;
      RECT 26.685 3.09 27.485 3.39 ;
      RECT 27.18 3.06 27.48 3.405 ;
      RECT 26.495 4.775 26.825 5.105 ;
      RECT 26.495 4.79 27.295 5.09 ;
      RECT 25.815 2.39 26.145 2.72 ;
      RECT 25.345 2.41 25.705 2.71 ;
      RECT 25.705 2.405 26.145 2.705 ;
      RECT 11.27 2.735 11.6 3.065 ;
      RECT 11.27 2.75 12.07 3.05 ;
      RECT 11.27 2.73 11.59 3.065 ;
      RECT 5.59 7.97 9.87 8.27 ;
      RECT 9.565 5.795 9.865 8.27 ;
      RECT 5.59 7.03 5.89 8.27 ;
      RECT 4.715 6.995 5.085 7.365 ;
      RECT 4.715 7.03 5.89 7.33 ;
      RECT 10.59 5.795 10.92 6.125 ;
      RECT 8.94 5.795 9.875 6.125 ;
      RECT 8.94 5.81 11.39 6.11 ;
      RECT 8.94 5.795 10.92 6.11 ;
      RECT 10.595 5.79 10.895 6.125 ;
      RECT 8.94 3.765 9.27 6.125 ;
      RECT 8.94 3.765 11.235 4.095 ;
      RECT 8.94 3.765 11.6 4.085 ;
      RECT 11.27 3.755 11.6 4.085 ;
      RECT 8.94 3.77 12.07 4.07 ;
      RECT 11.275 3.705 11.575 4.085 ;
      RECT 10.57 3.075 10.9 3.405 ;
      RECT 10.1 3.09 10.9 3.39 ;
      RECT 10.595 3.06 10.895 3.405 ;
      RECT 9.91 4.775 10.24 5.105 ;
      RECT 9.91 4.79 10.71 5.09 ;
      RECT 9.23 2.39 9.56 2.72 ;
      RECT 8.76 2.41 9.12 2.71 ;
      RECT 9.12 2.405 9.56 2.705 ;
    LAYER via2 ;
      RECT 77.67 2.8 77.87 3 ;
      RECT 77.67 3.82 77.87 4.02 ;
      RECT 76.99 5.86 77.19 6.06 ;
      RECT 76.97 3.14 77.17 3.34 ;
      RECT 76.31 4.84 76.51 5.04 ;
      RECT 75.945 5.86 76.145 6.06 ;
      RECT 75.63 2.455 75.83 2.655 ;
      RECT 71.135 7.08 71.335 7.28 ;
      RECT 61.09 2.8 61.29 3 ;
      RECT 61.09 3.82 61.29 4.02 ;
      RECT 60.41 5.86 60.61 6.06 ;
      RECT 60.39 3.14 60.59 3.34 ;
      RECT 59.73 4.84 59.93 5.04 ;
      RECT 59.365 5.86 59.565 6.06 ;
      RECT 59.05 2.455 59.25 2.655 ;
      RECT 54.555 7.08 54.755 7.28 ;
      RECT 44.505 2.8 44.705 3 ;
      RECT 44.505 3.82 44.705 4.02 ;
      RECT 43.825 5.86 44.025 6.06 ;
      RECT 43.805 3.14 44.005 3.34 ;
      RECT 43.145 4.84 43.345 5.04 ;
      RECT 42.78 5.86 42.98 6.06 ;
      RECT 42.465 2.455 42.665 2.655 ;
      RECT 37.97 7.08 38.17 7.28 ;
      RECT 27.92 2.8 28.12 3 ;
      RECT 27.92 3.82 28.12 4.02 ;
      RECT 27.24 5.86 27.44 6.06 ;
      RECT 27.22 3.14 27.42 3.34 ;
      RECT 26.56 4.84 26.76 5.04 ;
      RECT 26.195 5.86 26.395 6.06 ;
      RECT 25.88 2.455 26.08 2.655 ;
      RECT 21.385 7.08 21.585 7.28 ;
      RECT 11.335 2.8 11.535 3 ;
      RECT 11.335 3.82 11.535 4.02 ;
      RECT 10.655 5.86 10.855 6.06 ;
      RECT 10.635 3.14 10.835 3.34 ;
      RECT 9.975 4.84 10.175 5.04 ;
      RECT 9.61 5.86 9.81 6.06 ;
      RECT 9.295 2.455 9.495 2.655 ;
      RECT 4.8 7.08 5 7.28 ;
    LAYER met2 ;
      RECT 1.205 8.6 85.33 8.77 ;
      RECT 85.16 7.3 85.33 8.77 ;
      RECT 1.205 6.255 1.375 8.77 ;
      RECT 85.125 7.3 85.45 7.625 ;
      RECT 1.15 6.255 1.43 6.595 ;
      RECT 81.97 6.28 82.29 6.605 ;
      RECT 82 5.695 82.17 6.605 ;
      RECT 82 5.695 82.175 6.045 ;
      RECT 82 5.695 82.975 5.87 ;
      RECT 82.8 1.965 82.975 5.87 ;
      RECT 82.745 1.965 83.095 2.315 ;
      RECT 71.635 8.29 81.815 8.46 ;
      RECT 81.655 2.395 81.815 8.46 ;
      RECT 71.635 6.6 71.805 8.46 ;
      RECT 82.77 6.655 83.095 6.98 ;
      RECT 68.58 6.655 68.905 6.98 ;
      RECT 71.58 6.6 71.86 6.94 ;
      RECT 81.655 6.745 83.095 6.915 ;
      RECT 68.58 6.685 71.86 6.855 ;
      RECT 81.97 2.365 82.29 2.685 ;
      RECT 81.655 2.395 82.29 2.565 ;
      RECT 79.715 3.185 80.04 3.51 ;
      RECT 79.715 3.215 80.545 3.4 ;
      RECT 80.375 1.995 80.545 3.4 ;
      RECT 80.3 1.995 80.625 2.32 ;
      RECT 79.33 4.78 79.59 5.1 ;
      RECT 79.39 2.74 79.53 5.1 ;
      RECT 79.33 2.74 79.59 3.06 ;
      RECT 78.31 5.8 78.57 6.12 ;
      RECT 77.69 5.89 78.57 6.03 ;
      RECT 77.69 3.735 77.83 6.03 ;
      RECT 77.63 3.735 77.91 4.105 ;
      RECT 76.95 5.775 77.23 6.145 ;
      RECT 77.01 3.85 77.15 6.145 ;
      RECT 77.01 3.85 77.49 3.99 ;
      RECT 77.35 2.06 77.49 3.99 ;
      RECT 77.29 2.06 77.55 2.38 ;
      RECT 76.27 4.755 76.55 5.125 ;
      RECT 76.33 2.4 76.47 5.125 ;
      RECT 76.27 2.4 76.53 2.72 ;
      RECT 75.905 5.775 76.185 6.145 ;
      RECT 75.905 5.8 76.19 6.12 ;
      RECT 65.39 6.28 65.71 6.605 ;
      RECT 65.42 5.695 65.59 6.605 ;
      RECT 65.42 5.695 65.595 6.045 ;
      RECT 65.42 5.695 66.395 5.87 ;
      RECT 66.22 1.965 66.395 5.87 ;
      RECT 66.165 1.965 66.515 2.315 ;
      RECT 55.055 8.29 65.235 8.46 ;
      RECT 65.075 2.395 65.235 8.46 ;
      RECT 55.055 6.6 55.225 8.46 ;
      RECT 66.19 6.655 66.515 6.98 ;
      RECT 51.995 6.655 52.32 6.98 ;
      RECT 55 6.6 55.28 6.94 ;
      RECT 65.075 6.745 66.515 6.915 ;
      RECT 51.995 6.685 55.28 6.855 ;
      RECT 65.39 2.365 65.71 2.685 ;
      RECT 65.075 2.395 65.71 2.565 ;
      RECT 63.135 3.185 63.46 3.51 ;
      RECT 63.135 3.215 63.965 3.4 ;
      RECT 63.795 1.995 63.965 3.4 ;
      RECT 63.72 1.995 64.045 2.32 ;
      RECT 62.75 4.78 63.01 5.1 ;
      RECT 62.81 2.74 62.95 5.1 ;
      RECT 62.75 2.74 63.01 3.06 ;
      RECT 61.73 5.8 61.99 6.12 ;
      RECT 61.11 5.89 61.99 6.03 ;
      RECT 61.11 3.735 61.25 6.03 ;
      RECT 61.05 3.735 61.33 4.105 ;
      RECT 60.37 5.775 60.65 6.145 ;
      RECT 60.43 3.85 60.57 6.145 ;
      RECT 60.43 3.85 60.91 3.99 ;
      RECT 60.77 2.06 60.91 3.99 ;
      RECT 60.71 2.06 60.97 2.38 ;
      RECT 59.69 4.755 59.97 5.125 ;
      RECT 59.75 2.4 59.89 5.125 ;
      RECT 59.69 2.4 59.95 2.72 ;
      RECT 59.325 5.775 59.605 6.145 ;
      RECT 59.325 5.8 59.61 6.12 ;
      RECT 48.805 6.28 49.125 6.605 ;
      RECT 48.835 5.695 49.005 6.605 ;
      RECT 48.835 5.695 49.01 6.045 ;
      RECT 48.835 5.695 49.81 5.87 ;
      RECT 49.635 1.965 49.81 5.87 ;
      RECT 49.58 1.965 49.93 2.315 ;
      RECT 38.47 8.29 48.65 8.46 ;
      RECT 48.49 2.395 48.65 8.46 ;
      RECT 38.47 6.6 38.64 8.46 ;
      RECT 49.605 6.655 49.93 6.98 ;
      RECT 35.41 6.655 35.735 6.98 ;
      RECT 38.415 6.6 38.695 6.94 ;
      RECT 48.49 6.745 49.93 6.915 ;
      RECT 35.41 6.685 38.695 6.855 ;
      RECT 48.805 2.365 49.125 2.685 ;
      RECT 48.49 2.395 49.125 2.565 ;
      RECT 46.55 3.185 46.875 3.51 ;
      RECT 46.55 3.215 47.38 3.4 ;
      RECT 47.21 1.995 47.38 3.4 ;
      RECT 47.135 1.995 47.46 2.32 ;
      RECT 46.165 4.78 46.425 5.1 ;
      RECT 46.225 2.74 46.365 5.1 ;
      RECT 46.165 2.74 46.425 3.06 ;
      RECT 45.145 5.8 45.405 6.12 ;
      RECT 44.525 5.89 45.405 6.03 ;
      RECT 44.525 3.735 44.665 6.03 ;
      RECT 44.465 3.735 44.745 4.105 ;
      RECT 43.785 5.775 44.065 6.145 ;
      RECT 43.845 3.85 43.985 6.145 ;
      RECT 43.845 3.85 44.325 3.99 ;
      RECT 44.185 2.06 44.325 3.99 ;
      RECT 44.125 2.06 44.385 2.38 ;
      RECT 43.105 4.755 43.385 5.125 ;
      RECT 43.165 2.4 43.305 5.125 ;
      RECT 43.105 2.4 43.365 2.72 ;
      RECT 42.74 5.775 43.02 6.145 ;
      RECT 42.74 5.8 43.025 6.12 ;
      RECT 32.22 6.28 32.54 6.605 ;
      RECT 32.25 5.695 32.42 6.605 ;
      RECT 32.25 5.695 32.425 6.045 ;
      RECT 32.25 5.695 33.225 5.87 ;
      RECT 33.05 1.965 33.225 5.87 ;
      RECT 32.995 1.965 33.345 2.315 ;
      RECT 21.885 8.29 32.065 8.46 ;
      RECT 31.905 2.395 32.065 8.46 ;
      RECT 21.885 6.6 22.055 8.46 ;
      RECT 33.02 6.655 33.345 6.98 ;
      RECT 18.825 6.655 19.15 6.98 ;
      RECT 21.83 6.6 22.11 6.94 ;
      RECT 31.905 6.745 33.345 6.915 ;
      RECT 18.825 6.685 22.11 6.855 ;
      RECT 32.22 2.365 32.54 2.685 ;
      RECT 31.905 2.395 32.54 2.565 ;
      RECT 29.965 3.185 30.29 3.51 ;
      RECT 29.965 3.215 30.795 3.4 ;
      RECT 30.625 1.995 30.795 3.4 ;
      RECT 30.55 1.995 30.875 2.32 ;
      RECT 29.58 4.78 29.84 5.1 ;
      RECT 29.64 2.74 29.78 5.1 ;
      RECT 29.58 2.74 29.84 3.06 ;
      RECT 28.56 5.8 28.82 6.12 ;
      RECT 27.94 5.89 28.82 6.03 ;
      RECT 27.94 3.735 28.08 6.03 ;
      RECT 27.88 3.735 28.16 4.105 ;
      RECT 27.2 5.775 27.48 6.145 ;
      RECT 27.26 3.85 27.4 6.145 ;
      RECT 27.26 3.85 27.74 3.99 ;
      RECT 27.6 2.06 27.74 3.99 ;
      RECT 27.54 2.06 27.8 2.38 ;
      RECT 26.52 4.755 26.8 5.125 ;
      RECT 26.58 2.4 26.72 5.125 ;
      RECT 26.52 2.4 26.78 2.72 ;
      RECT 26.155 5.775 26.435 6.145 ;
      RECT 26.155 5.8 26.44 6.12 ;
      RECT 15.635 6.28 15.955 6.605 ;
      RECT 15.665 5.695 15.835 6.605 ;
      RECT 15.665 5.695 15.84 6.045 ;
      RECT 15.665 5.695 16.64 5.87 ;
      RECT 16.465 1.965 16.64 5.87 ;
      RECT 16.41 1.965 16.76 2.315 ;
      RECT 5.3 8.29 15.48 8.46 ;
      RECT 15.32 2.395 15.48 8.46 ;
      RECT 5.3 6.6 5.47 8.46 ;
      RECT 1.525 6.995 1.805 7.335 ;
      RECT 1.525 7.06 2.69 7.23 ;
      RECT 2.52 6.685 2.69 7.23 ;
      RECT 16.435 6.655 16.76 6.98 ;
      RECT 5.245 6.6 5.525 6.94 ;
      RECT 15.32 6.745 16.76 6.915 ;
      RECT 2.52 6.685 5.525 6.855 ;
      RECT 15.635 2.365 15.955 2.685 ;
      RECT 15.32 2.395 15.955 2.565 ;
      RECT 13.38 3.185 13.705 3.51 ;
      RECT 13.38 3.215 14.21 3.4 ;
      RECT 14.04 1.995 14.21 3.4 ;
      RECT 13.965 1.995 14.29 2.32 ;
      RECT 12.995 4.78 13.255 5.1 ;
      RECT 13.055 2.74 13.195 5.1 ;
      RECT 12.995 2.74 13.255 3.06 ;
      RECT 11.975 5.8 12.235 6.12 ;
      RECT 11.355 5.89 12.235 6.03 ;
      RECT 11.355 3.735 11.495 6.03 ;
      RECT 11.295 3.735 11.575 4.105 ;
      RECT 10.615 5.775 10.895 6.145 ;
      RECT 10.675 3.85 10.815 6.145 ;
      RECT 10.675 3.85 11.155 3.99 ;
      RECT 11.015 2.06 11.155 3.99 ;
      RECT 10.955 2.06 11.215 2.38 ;
      RECT 9.935 4.755 10.215 5.125 ;
      RECT 9.995 2.4 10.135 5.125 ;
      RECT 9.935 2.4 10.195 2.72 ;
      RECT 9.57 5.775 9.85 6.145 ;
      RECT 9.57 5.8 9.855 6.12 ;
      RECT 77.63 2.715 77.91 3.085 ;
      RECT 76.93 3.055 77.21 3.425 ;
      RECT 75.59 2.37 75.87 2.74 ;
      RECT 71.05 6.995 71.425 7.365 ;
      RECT 61.05 2.715 61.33 3.085 ;
      RECT 60.35 3.055 60.63 3.425 ;
      RECT 59.01 2.37 59.29 2.74 ;
      RECT 54.47 6.995 54.84 7.365 ;
      RECT 44.465 2.715 44.745 3.085 ;
      RECT 43.765 3.055 44.045 3.425 ;
      RECT 42.425 2.37 42.705 2.74 ;
      RECT 37.885 6.995 38.255 7.365 ;
      RECT 27.88 2.715 28.16 3.085 ;
      RECT 27.18 3.055 27.46 3.425 ;
      RECT 25.84 2.37 26.12 2.74 ;
      RECT 21.3 6.995 21.67 7.365 ;
      RECT 11.295 2.715 11.575 3.085 ;
      RECT 10.595 3.055 10.875 3.425 ;
      RECT 9.255 2.37 9.535 2.74 ;
      RECT 4.715 6.995 5.085 7.365 ;
    LAYER via1 ;
      RECT 85.215 7.385 85.365 7.535 ;
      RECT 82.86 6.74 83.01 6.89 ;
      RECT 82.845 2.065 82.995 2.215 ;
      RECT 82.055 2.45 82.205 2.6 ;
      RECT 82.055 6.37 82.205 6.52 ;
      RECT 80.39 2.08 80.54 2.23 ;
      RECT 79.805 3.27 79.955 3.42 ;
      RECT 79.385 2.825 79.535 2.975 ;
      RECT 79.385 4.865 79.535 5.015 ;
      RECT 78.365 5.885 78.515 6.035 ;
      RECT 77.685 2.825 77.835 2.975 ;
      RECT 77.685 3.845 77.835 3.995 ;
      RECT 77.345 2.145 77.495 2.295 ;
      RECT 77.005 3.165 77.155 3.315 ;
      RECT 77.005 5.885 77.155 6.035 ;
      RECT 76.325 2.485 76.475 2.635 ;
      RECT 76.325 4.865 76.475 5.015 ;
      RECT 75.985 5.885 76.135 6.035 ;
      RECT 75.645 2.48 75.795 2.63 ;
      RECT 71.645 6.695 71.795 6.845 ;
      RECT 71.16 7.105 71.31 7.255 ;
      RECT 68.67 6.74 68.82 6.89 ;
      RECT 66.28 6.74 66.43 6.89 ;
      RECT 66.265 2.065 66.415 2.215 ;
      RECT 65.475 2.45 65.625 2.6 ;
      RECT 65.475 6.37 65.625 6.52 ;
      RECT 63.81 2.08 63.96 2.23 ;
      RECT 63.225 3.27 63.375 3.42 ;
      RECT 62.805 2.825 62.955 2.975 ;
      RECT 62.805 4.865 62.955 5.015 ;
      RECT 61.785 5.885 61.935 6.035 ;
      RECT 61.105 2.825 61.255 2.975 ;
      RECT 61.105 3.845 61.255 3.995 ;
      RECT 60.765 2.145 60.915 2.295 ;
      RECT 60.425 3.165 60.575 3.315 ;
      RECT 60.425 5.885 60.575 6.035 ;
      RECT 59.745 2.485 59.895 2.635 ;
      RECT 59.745 4.865 59.895 5.015 ;
      RECT 59.405 5.885 59.555 6.035 ;
      RECT 59.065 2.48 59.215 2.63 ;
      RECT 55.065 6.695 55.215 6.845 ;
      RECT 54.58 7.105 54.73 7.255 ;
      RECT 52.085 6.74 52.235 6.89 ;
      RECT 49.695 6.74 49.845 6.89 ;
      RECT 49.68 2.065 49.83 2.215 ;
      RECT 48.89 2.45 49.04 2.6 ;
      RECT 48.89 6.37 49.04 6.52 ;
      RECT 47.225 2.08 47.375 2.23 ;
      RECT 46.64 3.27 46.79 3.42 ;
      RECT 46.22 2.825 46.37 2.975 ;
      RECT 46.22 4.865 46.37 5.015 ;
      RECT 45.2 5.885 45.35 6.035 ;
      RECT 44.52 2.825 44.67 2.975 ;
      RECT 44.52 3.845 44.67 3.995 ;
      RECT 44.18 2.145 44.33 2.295 ;
      RECT 43.84 3.165 43.99 3.315 ;
      RECT 43.84 5.885 43.99 6.035 ;
      RECT 43.16 2.485 43.31 2.635 ;
      RECT 43.16 4.865 43.31 5.015 ;
      RECT 42.82 5.885 42.97 6.035 ;
      RECT 42.48 2.48 42.63 2.63 ;
      RECT 38.48 6.695 38.63 6.845 ;
      RECT 37.995 7.105 38.145 7.255 ;
      RECT 35.5 6.74 35.65 6.89 ;
      RECT 33.11 6.74 33.26 6.89 ;
      RECT 33.095 2.065 33.245 2.215 ;
      RECT 32.305 2.45 32.455 2.6 ;
      RECT 32.305 6.37 32.455 6.52 ;
      RECT 30.64 2.08 30.79 2.23 ;
      RECT 30.055 3.27 30.205 3.42 ;
      RECT 29.635 2.825 29.785 2.975 ;
      RECT 29.635 4.865 29.785 5.015 ;
      RECT 28.615 5.885 28.765 6.035 ;
      RECT 27.935 2.825 28.085 2.975 ;
      RECT 27.935 3.845 28.085 3.995 ;
      RECT 27.595 2.145 27.745 2.295 ;
      RECT 27.255 3.165 27.405 3.315 ;
      RECT 27.255 5.885 27.405 6.035 ;
      RECT 26.575 2.485 26.725 2.635 ;
      RECT 26.575 4.865 26.725 5.015 ;
      RECT 26.235 5.885 26.385 6.035 ;
      RECT 25.895 2.48 26.045 2.63 ;
      RECT 21.895 6.695 22.045 6.845 ;
      RECT 21.41 7.105 21.56 7.255 ;
      RECT 18.915 6.74 19.065 6.89 ;
      RECT 16.525 6.74 16.675 6.89 ;
      RECT 16.51 2.065 16.66 2.215 ;
      RECT 15.72 2.45 15.87 2.6 ;
      RECT 15.72 6.37 15.87 6.52 ;
      RECT 14.055 2.08 14.205 2.23 ;
      RECT 13.47 3.27 13.62 3.42 ;
      RECT 13.05 2.825 13.2 2.975 ;
      RECT 13.05 4.865 13.2 5.015 ;
      RECT 12.03 5.885 12.18 6.035 ;
      RECT 11.35 2.825 11.5 2.975 ;
      RECT 11.35 3.845 11.5 3.995 ;
      RECT 11.01 2.145 11.16 2.295 ;
      RECT 10.67 3.165 10.82 3.315 ;
      RECT 10.67 5.885 10.82 6.035 ;
      RECT 9.99 2.485 10.14 2.635 ;
      RECT 9.99 4.865 10.14 5.015 ;
      RECT 9.65 5.885 9.8 6.035 ;
      RECT 9.31 2.48 9.46 2.63 ;
      RECT 5.31 6.695 5.46 6.845 ;
      RECT 4.825 7.105 4.975 7.255 ;
      RECT 1.59 7.09 1.74 7.24 ;
      RECT 1.215 6.35 1.365 6.5 ;
    LAYER met1 ;
      RECT 85.095 7.77 85.385 8 ;
      RECT 85.155 6.29 85.325 8 ;
      RECT 85.125 7.3 85.45 7.625 ;
      RECT 85.095 6.29 85.385 6.52 ;
      RECT 84.69 2.395 84.795 2.965 ;
      RECT 84.69 2.73 85.015 2.96 ;
      RECT 84.69 2.76 85.185 2.93 ;
      RECT 84.69 2.395 84.88 2.96 ;
      RECT 84.105 2.36 84.395 2.59 ;
      RECT 84.105 2.395 84.88 2.565 ;
      RECT 84.165 0.88 84.335 2.59 ;
      RECT 84.105 0.88 84.395 1.11 ;
      RECT 84.105 7.77 84.395 8 ;
      RECT 84.165 6.29 84.335 8 ;
      RECT 84.105 6.29 84.395 6.52 ;
      RECT 84.105 6.325 84.96 6.485 ;
      RECT 84.79 5.92 84.96 6.485 ;
      RECT 84.105 6.32 84.5 6.485 ;
      RECT 84.725 5.92 85.015 6.15 ;
      RECT 84.725 5.95 85.185 6.12 ;
      RECT 83.735 2.73 84.025 2.96 ;
      RECT 83.735 2.76 84.195 2.93 ;
      RECT 83.8 1.655 83.965 2.96 ;
      RECT 82.315 1.625 82.605 1.855 ;
      RECT 82.315 1.655 83.965 1.825 ;
      RECT 82.375 0.885 82.545 1.855 ;
      RECT 82.315 0.885 82.605 1.115 ;
      RECT 82.315 7.765 82.605 7.995 ;
      RECT 82.375 7.025 82.545 7.995 ;
      RECT 82.375 7.12 83.965 7.29 ;
      RECT 83.795 5.92 83.965 7.29 ;
      RECT 82.315 7.025 82.605 7.255 ;
      RECT 83.735 5.92 84.025 6.15 ;
      RECT 83.735 5.95 84.195 6.12 ;
      RECT 80.3 1.995 80.625 2.32 ;
      RECT 82.745 1.965 83.095 2.315 ;
      RECT 80.3 2.025 83.095 2.195 ;
      RECT 82.77 6.655 83.095 6.98 ;
      RECT 82.745 6.655 83.095 6.885 ;
      RECT 82.575 6.685 83.095 6.855 ;
      RECT 81.97 2.365 82.29 2.685 ;
      RECT 81.94 2.365 82.29 2.595 ;
      RECT 81.655 2.395 82.29 2.565 ;
      RECT 81.97 6.28 82.29 6.605 ;
      RECT 81.94 6.285 82.29 6.515 ;
      RECT 81.77 6.315 82.29 6.485 ;
      RECT 79.715 3.185 80.04 3.51 ;
      RECT 76.92 3.11 77.24 3.37 ;
      RECT 78.895 3.125 79.185 3.355 ;
      RECT 79.615 3.185 80.04 3.325 ;
      RECT 76.92 3.17 79.755 3.31 ;
      RECT 79.3 2.77 79.62 3.03 ;
      RECT 79.025 2.83 79.62 2.97 ;
      RECT 78.28 5.83 78.6 6.09 ;
      RECT 78.28 5.89 78.875 6.03 ;
      RECT 77.6 2.77 77.92 3.03 ;
      RECT 72.86 2.785 73.15 3.015 ;
      RECT 72.86 2.83 77.92 2.97 ;
      RECT 77.69 2.49 77.83 3.03 ;
      RECT 77.69 2.49 78.17 2.63 ;
      RECT 78.03 2.105 78.17 2.63 ;
      RECT 77.955 2.105 78.245 2.335 ;
      RECT 77.6 3.79 77.92 4.05 ;
      RECT 76.935 3.805 77.225 4.035 ;
      RECT 74.725 3.805 75.015 4.035 ;
      RECT 74.725 3.85 77.92 3.99 ;
      RECT 75.9 5.83 76.22 6.09 ;
      RECT 77.615 5.845 77.905 6.075 ;
      RECT 75.235 5.845 75.525 6.075 ;
      RECT 75.235 5.89 76.22 6.03 ;
      RECT 77.69 5.55 77.83 6.075 ;
      RECT 75.99 5.55 76.13 6.09 ;
      RECT 75.99 5.55 77.83 5.69 ;
      RECT 74.895 2.445 75.185 2.675 ;
      RECT 74.97 2.15 75.11 2.675 ;
      RECT 77.26 2.09 77.58 2.35 ;
      RECT 77.16 2.105 77.58 2.335 ;
      RECT 74.97 2.15 77.58 2.29 ;
      RECT 76.24 2.43 76.56 2.69 ;
      RECT 76.24 2.49 76.835 2.63 ;
      RECT 76.24 4.81 76.56 5.07 ;
      RECT 73.535 4.825 73.825 5.055 ;
      RECT 73.535 4.87 76.56 5.01 ;
      RECT 75.565 2.39 75.895 2.72 ;
      RECT 75.56 2.425 75.895 2.685 ;
      RECT 75.91 2.445 76.025 2.675 ;
      RECT 75.56 2.44 75.91 2.67 ;
      RECT 75.56 2.49 76.04 2.63 ;
      RECT 75.445 2.49 75.455 2.63 ;
      RECT 75.455 2.485 76.025 2.625 ;
      RECT 71.55 6.63 71.89 6.91 ;
      RECT 71.52 6.655 71.89 6.885 ;
      RECT 71.35 6.685 71.89 6.855 ;
      RECT 71.09 7.765 71.38 7.995 ;
      RECT 71.15 6.995 71.32 7.995 ;
      RECT 71.05 6.995 71.42 7.365 ;
      RECT 68.515 7.77 68.805 8 ;
      RECT 68.575 6.29 68.745 8 ;
      RECT 68.575 6.655 68.905 6.98 ;
      RECT 68.515 6.29 68.805 6.52 ;
      RECT 68.11 2.395 68.215 2.965 ;
      RECT 68.11 2.73 68.435 2.96 ;
      RECT 68.11 2.76 68.605 2.93 ;
      RECT 68.11 2.395 68.3 2.96 ;
      RECT 67.525 2.36 67.815 2.59 ;
      RECT 67.525 2.395 68.3 2.565 ;
      RECT 67.585 0.88 67.755 2.59 ;
      RECT 67.525 0.88 67.815 1.11 ;
      RECT 67.525 7.77 67.815 8 ;
      RECT 67.585 6.29 67.755 8 ;
      RECT 67.525 6.29 67.815 6.52 ;
      RECT 67.525 6.325 68.38 6.485 ;
      RECT 68.21 5.92 68.38 6.485 ;
      RECT 67.525 6.32 67.92 6.485 ;
      RECT 68.145 5.92 68.435 6.15 ;
      RECT 68.145 5.95 68.605 6.12 ;
      RECT 67.155 2.73 67.445 2.96 ;
      RECT 67.155 2.76 67.615 2.93 ;
      RECT 67.22 1.655 67.385 2.96 ;
      RECT 65.735 1.625 66.025 1.855 ;
      RECT 65.735 1.655 67.385 1.825 ;
      RECT 65.795 0.885 65.965 1.855 ;
      RECT 65.735 0.885 66.025 1.115 ;
      RECT 65.735 7.765 66.025 7.995 ;
      RECT 65.795 7.025 65.965 7.995 ;
      RECT 65.795 7.12 67.385 7.29 ;
      RECT 67.215 5.92 67.385 7.29 ;
      RECT 65.735 7.025 66.025 7.255 ;
      RECT 67.155 5.92 67.445 6.15 ;
      RECT 67.155 5.95 67.615 6.12 ;
      RECT 63.72 1.995 64.045 2.32 ;
      RECT 66.165 1.965 66.515 2.315 ;
      RECT 63.72 2.025 66.515 2.195 ;
      RECT 66.19 6.655 66.515 6.98 ;
      RECT 66.165 6.655 66.515 6.885 ;
      RECT 65.995 6.685 66.515 6.855 ;
      RECT 65.39 2.365 65.71 2.685 ;
      RECT 65.36 2.365 65.71 2.595 ;
      RECT 65.075 2.395 65.71 2.565 ;
      RECT 65.39 6.28 65.71 6.605 ;
      RECT 65.36 6.285 65.71 6.515 ;
      RECT 65.19 6.315 65.71 6.485 ;
      RECT 63.135 3.185 63.46 3.51 ;
      RECT 60.34 3.11 60.66 3.37 ;
      RECT 62.315 3.125 62.605 3.355 ;
      RECT 63.035 3.185 63.46 3.325 ;
      RECT 60.34 3.17 63.175 3.31 ;
      RECT 62.72 2.77 63.04 3.03 ;
      RECT 62.445 2.83 63.04 2.97 ;
      RECT 61.7 5.83 62.02 6.09 ;
      RECT 61.7 5.89 62.295 6.03 ;
      RECT 61.02 2.77 61.34 3.03 ;
      RECT 56.28 2.785 56.57 3.015 ;
      RECT 56.28 2.83 61.34 2.97 ;
      RECT 61.11 2.49 61.25 3.03 ;
      RECT 61.11 2.49 61.59 2.63 ;
      RECT 61.45 2.105 61.59 2.63 ;
      RECT 61.375 2.105 61.665 2.335 ;
      RECT 61.02 3.79 61.34 4.05 ;
      RECT 60.355 3.805 60.645 4.035 ;
      RECT 58.145 3.805 58.435 4.035 ;
      RECT 58.145 3.85 61.34 3.99 ;
      RECT 59.32 5.83 59.64 6.09 ;
      RECT 61.035 5.845 61.325 6.075 ;
      RECT 58.655 5.845 58.945 6.075 ;
      RECT 58.655 5.89 59.64 6.03 ;
      RECT 61.11 5.55 61.25 6.075 ;
      RECT 59.41 5.55 59.55 6.09 ;
      RECT 59.41 5.55 61.25 5.69 ;
      RECT 58.315 2.445 58.605 2.675 ;
      RECT 58.39 2.15 58.53 2.675 ;
      RECT 60.68 2.09 61 2.35 ;
      RECT 60.58 2.105 61 2.335 ;
      RECT 58.39 2.15 61 2.29 ;
      RECT 59.66 2.43 59.98 2.69 ;
      RECT 59.66 2.49 60.255 2.63 ;
      RECT 59.66 4.81 59.98 5.07 ;
      RECT 56.955 4.825 57.245 5.055 ;
      RECT 56.955 4.87 59.98 5.01 ;
      RECT 58.985 2.39 59.315 2.72 ;
      RECT 58.98 2.425 59.315 2.685 ;
      RECT 59.33 2.445 59.445 2.675 ;
      RECT 58.98 2.44 59.33 2.67 ;
      RECT 58.98 2.49 59.46 2.63 ;
      RECT 58.865 2.49 58.875 2.63 ;
      RECT 58.875 2.485 59.445 2.625 ;
      RECT 54.97 6.63 55.31 6.91 ;
      RECT 54.94 6.655 55.31 6.885 ;
      RECT 54.77 6.685 55.31 6.855 ;
      RECT 54.51 7.765 54.8 7.995 ;
      RECT 54.57 6.995 54.74 7.995 ;
      RECT 54.47 6.995 54.84 7.365 ;
      RECT 51.93 7.77 52.22 8 ;
      RECT 51.99 6.29 52.16 8 ;
      RECT 51.99 6.655 52.32 6.98 ;
      RECT 51.93 6.29 52.22 6.52 ;
      RECT 51.525 2.395 51.63 2.965 ;
      RECT 51.525 2.73 51.85 2.96 ;
      RECT 51.525 2.76 52.02 2.93 ;
      RECT 51.525 2.395 51.715 2.96 ;
      RECT 50.94 2.36 51.23 2.59 ;
      RECT 50.94 2.395 51.715 2.565 ;
      RECT 51 0.88 51.17 2.59 ;
      RECT 50.94 0.88 51.23 1.11 ;
      RECT 50.94 7.77 51.23 8 ;
      RECT 51 6.29 51.17 8 ;
      RECT 50.94 6.29 51.23 6.52 ;
      RECT 50.94 6.325 51.795 6.485 ;
      RECT 51.625 5.92 51.795 6.485 ;
      RECT 50.94 6.32 51.335 6.485 ;
      RECT 51.56 5.92 51.85 6.15 ;
      RECT 51.56 5.95 52.02 6.12 ;
      RECT 50.57 2.73 50.86 2.96 ;
      RECT 50.57 2.76 51.03 2.93 ;
      RECT 50.635 1.655 50.8 2.96 ;
      RECT 49.15 1.625 49.44 1.855 ;
      RECT 49.15 1.655 50.8 1.825 ;
      RECT 49.21 0.885 49.38 1.855 ;
      RECT 49.15 0.885 49.44 1.115 ;
      RECT 49.15 7.765 49.44 7.995 ;
      RECT 49.21 7.025 49.38 7.995 ;
      RECT 49.21 7.12 50.8 7.29 ;
      RECT 50.63 5.92 50.8 7.29 ;
      RECT 49.15 7.025 49.44 7.255 ;
      RECT 50.57 5.92 50.86 6.15 ;
      RECT 50.57 5.95 51.03 6.12 ;
      RECT 47.135 1.995 47.46 2.32 ;
      RECT 49.58 1.965 49.93 2.315 ;
      RECT 47.135 2.025 49.93 2.195 ;
      RECT 49.605 6.655 49.93 6.98 ;
      RECT 49.58 6.655 49.93 6.885 ;
      RECT 49.41 6.685 49.93 6.855 ;
      RECT 48.805 2.365 49.125 2.685 ;
      RECT 48.775 2.365 49.125 2.595 ;
      RECT 48.49 2.395 49.125 2.565 ;
      RECT 48.805 6.28 49.125 6.605 ;
      RECT 48.775 6.285 49.125 6.515 ;
      RECT 48.605 6.315 49.125 6.485 ;
      RECT 46.55 3.185 46.875 3.51 ;
      RECT 43.755 3.11 44.075 3.37 ;
      RECT 45.73 3.125 46.02 3.355 ;
      RECT 46.45 3.185 46.875 3.325 ;
      RECT 43.755 3.17 46.59 3.31 ;
      RECT 46.135 2.77 46.455 3.03 ;
      RECT 45.86 2.83 46.455 2.97 ;
      RECT 45.115 5.83 45.435 6.09 ;
      RECT 45.115 5.89 45.71 6.03 ;
      RECT 44.435 2.77 44.755 3.03 ;
      RECT 39.695 2.785 39.985 3.015 ;
      RECT 39.695 2.83 44.755 2.97 ;
      RECT 44.525 2.49 44.665 3.03 ;
      RECT 44.525 2.49 45.005 2.63 ;
      RECT 44.865 2.105 45.005 2.63 ;
      RECT 44.79 2.105 45.08 2.335 ;
      RECT 44.435 3.79 44.755 4.05 ;
      RECT 43.77 3.805 44.06 4.035 ;
      RECT 41.56 3.805 41.85 4.035 ;
      RECT 41.56 3.85 44.755 3.99 ;
      RECT 42.735 5.83 43.055 6.09 ;
      RECT 44.45 5.845 44.74 6.075 ;
      RECT 42.07 5.845 42.36 6.075 ;
      RECT 42.07 5.89 43.055 6.03 ;
      RECT 44.525 5.55 44.665 6.075 ;
      RECT 42.825 5.55 42.965 6.09 ;
      RECT 42.825 5.55 44.665 5.69 ;
      RECT 41.73 2.445 42.02 2.675 ;
      RECT 41.805 2.15 41.945 2.675 ;
      RECT 44.095 2.09 44.415 2.35 ;
      RECT 43.995 2.105 44.415 2.335 ;
      RECT 41.805 2.15 44.415 2.29 ;
      RECT 43.075 2.43 43.395 2.69 ;
      RECT 43.075 2.49 43.67 2.63 ;
      RECT 43.075 4.81 43.395 5.07 ;
      RECT 40.37 4.825 40.66 5.055 ;
      RECT 40.37 4.87 43.395 5.01 ;
      RECT 42.4 2.39 42.73 2.72 ;
      RECT 42.395 2.425 42.73 2.685 ;
      RECT 42.745 2.445 42.86 2.675 ;
      RECT 42.395 2.44 42.745 2.67 ;
      RECT 42.395 2.49 42.875 2.63 ;
      RECT 42.28 2.49 42.29 2.63 ;
      RECT 42.29 2.485 42.86 2.625 ;
      RECT 38.385 6.63 38.725 6.91 ;
      RECT 38.355 6.655 38.725 6.885 ;
      RECT 38.185 6.685 38.725 6.855 ;
      RECT 37.925 7.765 38.215 7.995 ;
      RECT 37.985 6.995 38.155 7.995 ;
      RECT 37.885 6.995 38.255 7.365 ;
      RECT 35.345 7.77 35.635 8 ;
      RECT 35.405 6.29 35.575 8 ;
      RECT 35.405 6.655 35.735 6.98 ;
      RECT 35.345 6.29 35.635 6.52 ;
      RECT 34.94 2.395 35.045 2.965 ;
      RECT 34.94 2.73 35.265 2.96 ;
      RECT 34.94 2.76 35.435 2.93 ;
      RECT 34.94 2.395 35.13 2.96 ;
      RECT 34.355 2.36 34.645 2.59 ;
      RECT 34.355 2.395 35.13 2.565 ;
      RECT 34.415 0.88 34.585 2.59 ;
      RECT 34.355 0.88 34.645 1.11 ;
      RECT 34.355 7.77 34.645 8 ;
      RECT 34.415 6.29 34.585 8 ;
      RECT 34.355 6.29 34.645 6.52 ;
      RECT 34.355 6.325 35.21 6.485 ;
      RECT 35.04 5.92 35.21 6.485 ;
      RECT 34.355 6.32 34.75 6.485 ;
      RECT 34.975 5.92 35.265 6.15 ;
      RECT 34.975 5.95 35.435 6.12 ;
      RECT 33.985 2.73 34.275 2.96 ;
      RECT 33.985 2.76 34.445 2.93 ;
      RECT 34.05 1.655 34.215 2.96 ;
      RECT 32.565 1.625 32.855 1.855 ;
      RECT 32.565 1.655 34.215 1.825 ;
      RECT 32.625 0.885 32.795 1.855 ;
      RECT 32.565 0.885 32.855 1.115 ;
      RECT 32.565 7.765 32.855 7.995 ;
      RECT 32.625 7.025 32.795 7.995 ;
      RECT 32.625 7.12 34.215 7.29 ;
      RECT 34.045 5.92 34.215 7.29 ;
      RECT 32.565 7.025 32.855 7.255 ;
      RECT 33.985 5.92 34.275 6.15 ;
      RECT 33.985 5.95 34.445 6.12 ;
      RECT 30.55 1.995 30.875 2.32 ;
      RECT 32.995 1.965 33.345 2.315 ;
      RECT 30.55 2.025 33.345 2.195 ;
      RECT 33.02 6.655 33.345 6.98 ;
      RECT 32.995 6.655 33.345 6.885 ;
      RECT 32.825 6.685 33.345 6.855 ;
      RECT 32.22 2.365 32.54 2.685 ;
      RECT 32.19 2.365 32.54 2.595 ;
      RECT 31.905 2.395 32.54 2.565 ;
      RECT 32.22 6.28 32.54 6.605 ;
      RECT 32.19 6.285 32.54 6.515 ;
      RECT 32.02 6.315 32.54 6.485 ;
      RECT 29.965 3.185 30.29 3.51 ;
      RECT 27.17 3.11 27.49 3.37 ;
      RECT 29.145 3.125 29.435 3.355 ;
      RECT 29.865 3.185 30.29 3.325 ;
      RECT 27.17 3.17 30.005 3.31 ;
      RECT 29.55 2.77 29.87 3.03 ;
      RECT 29.275 2.83 29.87 2.97 ;
      RECT 28.53 5.83 28.85 6.09 ;
      RECT 28.53 5.89 29.125 6.03 ;
      RECT 27.85 2.77 28.17 3.03 ;
      RECT 23.11 2.785 23.4 3.015 ;
      RECT 23.11 2.83 28.17 2.97 ;
      RECT 27.94 2.49 28.08 3.03 ;
      RECT 27.94 2.49 28.42 2.63 ;
      RECT 28.28 2.105 28.42 2.63 ;
      RECT 28.205 2.105 28.495 2.335 ;
      RECT 27.85 3.79 28.17 4.05 ;
      RECT 27.185 3.805 27.475 4.035 ;
      RECT 24.975 3.805 25.265 4.035 ;
      RECT 24.975 3.85 28.17 3.99 ;
      RECT 26.15 5.83 26.47 6.09 ;
      RECT 27.865 5.845 28.155 6.075 ;
      RECT 25.485 5.845 25.775 6.075 ;
      RECT 25.485 5.89 26.47 6.03 ;
      RECT 27.94 5.55 28.08 6.075 ;
      RECT 26.24 5.55 26.38 6.09 ;
      RECT 26.24 5.55 28.08 5.69 ;
      RECT 25.145 2.445 25.435 2.675 ;
      RECT 25.22 2.15 25.36 2.675 ;
      RECT 27.51 2.09 27.83 2.35 ;
      RECT 27.41 2.105 27.83 2.335 ;
      RECT 25.22 2.15 27.83 2.29 ;
      RECT 26.49 2.43 26.81 2.69 ;
      RECT 26.49 2.49 27.085 2.63 ;
      RECT 26.49 4.81 26.81 5.07 ;
      RECT 23.785 4.825 24.075 5.055 ;
      RECT 23.785 4.87 26.81 5.01 ;
      RECT 25.815 2.39 26.145 2.72 ;
      RECT 25.81 2.425 26.145 2.685 ;
      RECT 26.16 2.445 26.275 2.675 ;
      RECT 25.81 2.44 26.16 2.67 ;
      RECT 25.81 2.49 26.29 2.63 ;
      RECT 25.695 2.49 25.705 2.63 ;
      RECT 25.705 2.485 26.275 2.625 ;
      RECT 21.8 6.63 22.14 6.91 ;
      RECT 21.77 6.655 22.14 6.885 ;
      RECT 21.6 6.685 22.14 6.855 ;
      RECT 21.34 7.765 21.63 7.995 ;
      RECT 21.4 6.995 21.57 7.995 ;
      RECT 21.3 6.995 21.67 7.365 ;
      RECT 18.76 7.77 19.05 8 ;
      RECT 18.82 6.29 18.99 8 ;
      RECT 18.82 6.655 19.15 6.98 ;
      RECT 18.76 6.29 19.05 6.52 ;
      RECT 18.355 2.395 18.46 2.965 ;
      RECT 18.355 2.73 18.68 2.96 ;
      RECT 18.355 2.76 18.85 2.93 ;
      RECT 18.355 2.395 18.545 2.96 ;
      RECT 17.77 2.36 18.06 2.59 ;
      RECT 17.77 2.395 18.545 2.565 ;
      RECT 17.83 0.88 18 2.59 ;
      RECT 17.77 0.88 18.06 1.11 ;
      RECT 17.77 7.77 18.06 8 ;
      RECT 17.83 6.29 18 8 ;
      RECT 17.77 6.29 18.06 6.52 ;
      RECT 17.77 6.325 18.625 6.485 ;
      RECT 18.455 5.92 18.625 6.485 ;
      RECT 17.77 6.32 18.165 6.485 ;
      RECT 18.39 5.92 18.68 6.15 ;
      RECT 18.39 5.95 18.85 6.12 ;
      RECT 17.4 2.73 17.69 2.96 ;
      RECT 17.4 2.76 17.86 2.93 ;
      RECT 17.465 1.655 17.63 2.96 ;
      RECT 15.98 1.625 16.27 1.855 ;
      RECT 15.98 1.655 17.63 1.825 ;
      RECT 16.04 0.885 16.21 1.855 ;
      RECT 15.98 0.885 16.27 1.115 ;
      RECT 15.98 7.765 16.27 7.995 ;
      RECT 16.04 7.025 16.21 7.995 ;
      RECT 16.04 7.12 17.63 7.29 ;
      RECT 17.46 5.92 17.63 7.29 ;
      RECT 15.98 7.025 16.27 7.255 ;
      RECT 17.4 5.92 17.69 6.15 ;
      RECT 17.4 5.95 17.86 6.12 ;
      RECT 13.965 1.995 14.29 2.32 ;
      RECT 16.41 1.965 16.76 2.315 ;
      RECT 13.965 2.025 16.76 2.195 ;
      RECT 16.435 6.655 16.76 6.98 ;
      RECT 16.41 6.655 16.76 6.885 ;
      RECT 16.24 6.685 16.76 6.855 ;
      RECT 15.635 2.365 15.955 2.685 ;
      RECT 15.605 2.365 15.955 2.595 ;
      RECT 15.32 2.395 15.955 2.565 ;
      RECT 15.635 6.28 15.955 6.605 ;
      RECT 15.605 6.285 15.955 6.515 ;
      RECT 15.435 6.315 15.955 6.485 ;
      RECT 13.38 3.185 13.705 3.51 ;
      RECT 10.585 3.11 10.905 3.37 ;
      RECT 12.56 3.125 12.85 3.355 ;
      RECT 13.28 3.185 13.705 3.325 ;
      RECT 10.585 3.17 13.42 3.31 ;
      RECT 12.965 2.77 13.285 3.03 ;
      RECT 12.69 2.83 13.285 2.97 ;
      RECT 11.945 5.83 12.265 6.09 ;
      RECT 11.945 5.89 12.54 6.03 ;
      RECT 11.265 2.77 11.585 3.03 ;
      RECT 6.525 2.785 6.815 3.015 ;
      RECT 6.525 2.83 11.585 2.97 ;
      RECT 11.355 2.49 11.495 3.03 ;
      RECT 11.355 2.49 11.835 2.63 ;
      RECT 11.695 2.105 11.835 2.63 ;
      RECT 11.62 2.105 11.91 2.335 ;
      RECT 11.265 3.79 11.585 4.05 ;
      RECT 10.6 3.805 10.89 4.035 ;
      RECT 8.39 3.805 8.68 4.035 ;
      RECT 8.39 3.85 11.585 3.99 ;
      RECT 9.565 5.83 9.885 6.09 ;
      RECT 11.28 5.845 11.57 6.075 ;
      RECT 8.9 5.845 9.19 6.075 ;
      RECT 8.9 5.89 9.885 6.03 ;
      RECT 11.355 5.55 11.495 6.075 ;
      RECT 9.655 5.55 9.795 6.09 ;
      RECT 9.655 5.55 11.495 5.69 ;
      RECT 8.56 2.445 8.85 2.675 ;
      RECT 8.635 2.15 8.775 2.675 ;
      RECT 10.925 2.09 11.245 2.35 ;
      RECT 10.825 2.105 11.245 2.335 ;
      RECT 8.635 2.15 11.245 2.29 ;
      RECT 9.905 2.43 10.225 2.69 ;
      RECT 9.905 2.49 10.5 2.63 ;
      RECT 9.905 4.81 10.225 5.07 ;
      RECT 7.2 4.825 7.49 5.055 ;
      RECT 7.2 4.87 10.225 5.01 ;
      RECT 9.23 2.39 9.56 2.72 ;
      RECT 9.225 2.425 9.56 2.685 ;
      RECT 9.575 2.445 9.69 2.675 ;
      RECT 9.225 2.44 9.575 2.67 ;
      RECT 9.225 2.49 9.705 2.63 ;
      RECT 9.11 2.49 9.12 2.63 ;
      RECT 9.12 2.485 9.69 2.625 ;
      RECT 5.215 6.63 5.555 6.91 ;
      RECT 5.185 6.655 5.555 6.885 ;
      RECT 5.015 6.685 5.555 6.855 ;
      RECT 4.755 7.765 5.045 7.995 ;
      RECT 4.815 6.995 4.985 7.995 ;
      RECT 4.715 6.995 5.085 7.365 ;
      RECT 1.525 7.765 1.815 7.995 ;
      RECT 1.585 7.025 1.755 7.995 ;
      RECT 1.495 7.025 1.835 7.305 ;
      RECT 1.12 6.285 1.46 6.565 ;
      RECT 0.98 6.315 1.46 6.485 ;
      RECT 78.975 4.81 79.62 5.07 ;
      RECT 76.92 5.83 77.24 6.09 ;
      RECT 62.395 4.81 63.04 5.07 ;
      RECT 60.34 5.83 60.66 6.09 ;
      RECT 45.81 4.81 46.455 5.07 ;
      RECT 43.755 5.83 44.075 6.09 ;
      RECT 29.225 4.81 29.87 5.07 ;
      RECT 27.17 5.83 27.49 6.09 ;
      RECT 12.64 4.81 13.285 5.07 ;
      RECT 10.585 5.83 10.905 6.09 ;
    LAYER mcon ;
      RECT 85.155 6.32 85.325 6.49 ;
      RECT 85.16 6.315 85.33 6.485 ;
      RECT 68.575 6.32 68.745 6.49 ;
      RECT 68.58 6.315 68.75 6.485 ;
      RECT 51.99 6.32 52.16 6.49 ;
      RECT 51.995 6.315 52.165 6.485 ;
      RECT 35.405 6.32 35.575 6.49 ;
      RECT 35.41 6.315 35.58 6.485 ;
      RECT 18.82 6.32 18.99 6.49 ;
      RECT 18.825 6.315 18.995 6.485 ;
      RECT 85.155 7.8 85.325 7.97 ;
      RECT 84.785 2.76 84.955 2.93 ;
      RECT 84.785 5.95 84.955 6.12 ;
      RECT 84.165 0.91 84.335 1.08 ;
      RECT 84.165 2.39 84.335 2.56 ;
      RECT 84.165 6.32 84.335 6.49 ;
      RECT 84.165 7.8 84.335 7.97 ;
      RECT 83.795 2.76 83.965 2.93 ;
      RECT 83.795 5.95 83.965 6.12 ;
      RECT 82.805 2.025 82.975 2.195 ;
      RECT 82.805 6.685 82.975 6.855 ;
      RECT 82.375 0.915 82.545 1.085 ;
      RECT 82.375 1.655 82.545 1.825 ;
      RECT 82.375 7.055 82.545 7.225 ;
      RECT 82.375 7.795 82.545 7.965 ;
      RECT 82 2.395 82.17 2.565 ;
      RECT 82 6.315 82.17 6.485 ;
      RECT 79.375 2.815 79.545 2.985 ;
      RECT 79.035 4.855 79.205 5.025 ;
      RECT 78.955 3.155 79.125 3.325 ;
      RECT 78.355 5.875 78.525 6.045 ;
      RECT 78.015 2.135 78.185 2.305 ;
      RECT 77.675 5.875 77.845 6.045 ;
      RECT 77.22 2.135 77.39 2.305 ;
      RECT 76.995 3.835 77.165 4.005 ;
      RECT 76.995 5.875 77.165 6.045 ;
      RECT 76.315 2.475 76.485 2.645 ;
      RECT 75.295 5.875 75.465 6.045 ;
      RECT 74.955 2.475 75.125 2.645 ;
      RECT 74.785 3.835 74.955 4.005 ;
      RECT 73.595 4.855 73.765 5.025 ;
      RECT 72.92 2.815 73.09 2.985 ;
      RECT 71.58 6.685 71.75 6.855 ;
      RECT 71.15 7.055 71.32 7.225 ;
      RECT 71.15 7.795 71.32 7.965 ;
      RECT 68.575 7.8 68.745 7.97 ;
      RECT 68.205 2.76 68.375 2.93 ;
      RECT 68.205 5.95 68.375 6.12 ;
      RECT 67.585 0.91 67.755 1.08 ;
      RECT 67.585 2.39 67.755 2.56 ;
      RECT 67.585 6.32 67.755 6.49 ;
      RECT 67.585 7.8 67.755 7.97 ;
      RECT 67.215 2.76 67.385 2.93 ;
      RECT 67.215 5.95 67.385 6.12 ;
      RECT 66.225 2.025 66.395 2.195 ;
      RECT 66.225 6.685 66.395 6.855 ;
      RECT 65.795 0.915 65.965 1.085 ;
      RECT 65.795 1.655 65.965 1.825 ;
      RECT 65.795 7.055 65.965 7.225 ;
      RECT 65.795 7.795 65.965 7.965 ;
      RECT 65.42 2.395 65.59 2.565 ;
      RECT 65.42 6.315 65.59 6.485 ;
      RECT 62.795 2.815 62.965 2.985 ;
      RECT 62.455 4.855 62.625 5.025 ;
      RECT 62.375 3.155 62.545 3.325 ;
      RECT 61.775 5.875 61.945 6.045 ;
      RECT 61.435 2.135 61.605 2.305 ;
      RECT 61.095 5.875 61.265 6.045 ;
      RECT 60.64 2.135 60.81 2.305 ;
      RECT 60.415 3.835 60.585 4.005 ;
      RECT 60.415 5.875 60.585 6.045 ;
      RECT 59.735 2.475 59.905 2.645 ;
      RECT 58.715 5.875 58.885 6.045 ;
      RECT 58.375 2.475 58.545 2.645 ;
      RECT 58.205 3.835 58.375 4.005 ;
      RECT 57.015 4.855 57.185 5.025 ;
      RECT 56.34 2.815 56.51 2.985 ;
      RECT 55 6.685 55.17 6.855 ;
      RECT 54.57 7.055 54.74 7.225 ;
      RECT 54.57 7.795 54.74 7.965 ;
      RECT 51.99 7.8 52.16 7.97 ;
      RECT 51.62 2.76 51.79 2.93 ;
      RECT 51.62 5.95 51.79 6.12 ;
      RECT 51 0.91 51.17 1.08 ;
      RECT 51 2.39 51.17 2.56 ;
      RECT 51 6.32 51.17 6.49 ;
      RECT 51 7.8 51.17 7.97 ;
      RECT 50.63 2.76 50.8 2.93 ;
      RECT 50.63 5.95 50.8 6.12 ;
      RECT 49.64 2.025 49.81 2.195 ;
      RECT 49.64 6.685 49.81 6.855 ;
      RECT 49.21 0.915 49.38 1.085 ;
      RECT 49.21 1.655 49.38 1.825 ;
      RECT 49.21 7.055 49.38 7.225 ;
      RECT 49.21 7.795 49.38 7.965 ;
      RECT 48.835 2.395 49.005 2.565 ;
      RECT 48.835 6.315 49.005 6.485 ;
      RECT 46.21 2.815 46.38 2.985 ;
      RECT 45.87 4.855 46.04 5.025 ;
      RECT 45.79 3.155 45.96 3.325 ;
      RECT 45.19 5.875 45.36 6.045 ;
      RECT 44.85 2.135 45.02 2.305 ;
      RECT 44.51 5.875 44.68 6.045 ;
      RECT 44.055 2.135 44.225 2.305 ;
      RECT 43.83 3.835 44 4.005 ;
      RECT 43.83 5.875 44 6.045 ;
      RECT 43.15 2.475 43.32 2.645 ;
      RECT 42.13 5.875 42.3 6.045 ;
      RECT 41.79 2.475 41.96 2.645 ;
      RECT 41.62 3.835 41.79 4.005 ;
      RECT 40.43 4.855 40.6 5.025 ;
      RECT 39.755 2.815 39.925 2.985 ;
      RECT 38.415 6.685 38.585 6.855 ;
      RECT 37.985 7.055 38.155 7.225 ;
      RECT 37.985 7.795 38.155 7.965 ;
      RECT 35.405 7.8 35.575 7.97 ;
      RECT 35.035 2.76 35.205 2.93 ;
      RECT 35.035 5.95 35.205 6.12 ;
      RECT 34.415 0.91 34.585 1.08 ;
      RECT 34.415 2.39 34.585 2.56 ;
      RECT 34.415 6.32 34.585 6.49 ;
      RECT 34.415 7.8 34.585 7.97 ;
      RECT 34.045 2.76 34.215 2.93 ;
      RECT 34.045 5.95 34.215 6.12 ;
      RECT 33.055 2.025 33.225 2.195 ;
      RECT 33.055 6.685 33.225 6.855 ;
      RECT 32.625 0.915 32.795 1.085 ;
      RECT 32.625 1.655 32.795 1.825 ;
      RECT 32.625 7.055 32.795 7.225 ;
      RECT 32.625 7.795 32.795 7.965 ;
      RECT 32.25 2.395 32.42 2.565 ;
      RECT 32.25 6.315 32.42 6.485 ;
      RECT 29.625 2.815 29.795 2.985 ;
      RECT 29.285 4.855 29.455 5.025 ;
      RECT 29.205 3.155 29.375 3.325 ;
      RECT 28.605 5.875 28.775 6.045 ;
      RECT 28.265 2.135 28.435 2.305 ;
      RECT 27.925 5.875 28.095 6.045 ;
      RECT 27.47 2.135 27.64 2.305 ;
      RECT 27.245 3.835 27.415 4.005 ;
      RECT 27.245 5.875 27.415 6.045 ;
      RECT 26.565 2.475 26.735 2.645 ;
      RECT 25.545 5.875 25.715 6.045 ;
      RECT 25.205 2.475 25.375 2.645 ;
      RECT 25.035 3.835 25.205 4.005 ;
      RECT 23.845 4.855 24.015 5.025 ;
      RECT 23.17 2.815 23.34 2.985 ;
      RECT 21.83 6.685 22 6.855 ;
      RECT 21.4 7.055 21.57 7.225 ;
      RECT 21.4 7.795 21.57 7.965 ;
      RECT 18.82 7.8 18.99 7.97 ;
      RECT 18.45 2.76 18.62 2.93 ;
      RECT 18.45 5.95 18.62 6.12 ;
      RECT 17.83 0.91 18 1.08 ;
      RECT 17.83 2.39 18 2.56 ;
      RECT 17.83 6.32 18 6.49 ;
      RECT 17.83 7.8 18 7.97 ;
      RECT 17.46 2.76 17.63 2.93 ;
      RECT 17.46 5.95 17.63 6.12 ;
      RECT 16.47 2.025 16.64 2.195 ;
      RECT 16.47 6.685 16.64 6.855 ;
      RECT 16.04 0.915 16.21 1.085 ;
      RECT 16.04 1.655 16.21 1.825 ;
      RECT 16.04 7.055 16.21 7.225 ;
      RECT 16.04 7.795 16.21 7.965 ;
      RECT 15.665 2.395 15.835 2.565 ;
      RECT 15.665 6.315 15.835 6.485 ;
      RECT 13.04 2.815 13.21 2.985 ;
      RECT 12.7 4.855 12.87 5.025 ;
      RECT 12.62 3.155 12.79 3.325 ;
      RECT 12.02 5.875 12.19 6.045 ;
      RECT 11.68 2.135 11.85 2.305 ;
      RECT 11.34 5.875 11.51 6.045 ;
      RECT 10.885 2.135 11.055 2.305 ;
      RECT 10.66 3.835 10.83 4.005 ;
      RECT 10.66 5.875 10.83 6.045 ;
      RECT 9.98 2.475 10.15 2.645 ;
      RECT 8.96 5.875 9.13 6.045 ;
      RECT 8.62 2.475 8.79 2.645 ;
      RECT 8.45 3.835 8.62 4.005 ;
      RECT 7.26 4.855 7.43 5.025 ;
      RECT 6.585 2.815 6.755 2.985 ;
      RECT 5.245 6.685 5.415 6.855 ;
      RECT 4.815 7.055 4.985 7.225 ;
      RECT 4.815 7.795 4.985 7.965 ;
      RECT 1.585 7.055 1.755 7.225 ;
      RECT 1.585 7.795 1.755 7.965 ;
      RECT 1.21 6.315 1.38 6.485 ;
    LAYER li1 ;
      RECT 85.155 5.02 85.325 6.49 ;
      RECT 85.155 6.315 85.33 6.485 ;
      RECT 84.785 1.74 84.955 2.93 ;
      RECT 84.785 1.74 85.255 1.91 ;
      RECT 84.785 6.97 85.255 7.14 ;
      RECT 84.785 5.95 84.955 7.14 ;
      RECT 83.795 1.74 83.965 2.93 ;
      RECT 83.795 1.74 84.265 1.91 ;
      RECT 83.795 6.97 84.265 7.14 ;
      RECT 83.795 5.95 83.965 7.14 ;
      RECT 81.945 2.635 82.115 3.865 ;
      RECT 82 0.855 82.17 2.805 ;
      RECT 81.945 0.575 82.115 1.025 ;
      RECT 81.945 7.855 82.115 8.305 ;
      RECT 82 6.075 82.17 8.025 ;
      RECT 81.945 5.015 82.115 6.245 ;
      RECT 81.425 0.575 81.595 3.865 ;
      RECT 81.425 2.075 81.83 2.405 ;
      RECT 81.425 1.235 81.83 1.565 ;
      RECT 81.425 5.015 81.595 8.305 ;
      RECT 81.425 7.315 81.83 7.645 ;
      RECT 81.425 6.475 81.83 6.805 ;
      RECT 76.685 6.645 77.99 6.895 ;
      RECT 76.685 6.325 76.865 6.895 ;
      RECT 76.135 6.325 76.865 6.495 ;
      RECT 76.135 5.485 76.305 6.495 ;
      RECT 76.97 5.525 78.715 5.705 ;
      RECT 78.385 4.685 78.715 5.705 ;
      RECT 76.135 5.485 77.195 5.655 ;
      RECT 78.385 4.855 79.205 5.025 ;
      RECT 77.545 4.685 77.875 4.895 ;
      RECT 77.545 4.685 78.715 4.855 ;
      RECT 78.445 3.205 78.775 4.16 ;
      RECT 78.445 3.205 79.125 3.375 ;
      RECT 78.955 1.965 79.125 3.375 ;
      RECT 78.865 1.965 79.195 2.605 ;
      RECT 77.99 3.475 78.265 4.175 ;
      RECT 78.095 1.965 78.265 4.175 ;
      RECT 78.435 2.785 78.785 3.035 ;
      RECT 78.095 2.815 78.785 2.985 ;
      RECT 78.005 1.965 78.265 2.445 ;
      RECT 77.335 5.115 78.215 5.355 ;
      RECT 77.985 5.025 78.215 5.355 ;
      RECT 76.685 5.115 78.215 5.315 ;
      RECT 77.6 5.065 78.215 5.355 ;
      RECT 76.685 4.985 76.855 5.315 ;
      RECT 77.57 5.875 77.82 6.475 ;
      RECT 77.57 5.875 78.045 6.075 ;
      RECT 77.065 3.095 77.82 3.595 ;
      RECT 76.135 2.9 76.395 3.52 ;
      RECT 77.05 3.04 77.065 3.345 ;
      RECT 77.035 3.025 77.055 3.31 ;
      RECT 77.695 2.7 77.925 3.3 ;
      RECT 77.01 2.97 77.03 3.285 ;
      RECT 76.99 3.095 77.925 3.27 ;
      RECT 76.965 3.095 77.925 3.26 ;
      RECT 76.895 3.095 77.925 3.25 ;
      RECT 76.875 3.095 77.925 3.22 ;
      RECT 76.855 2.005 77.025 3.19 ;
      RECT 76.825 3.095 77.925 3.16 ;
      RECT 76.79 3.095 77.925 3.135 ;
      RECT 76.76 3.09 77.15 3.1 ;
      RECT 76.76 3.08 77.125 3.1 ;
      RECT 76.76 3.075 77.11 3.1 ;
      RECT 76.76 3.065 77.095 3.1 ;
      RECT 76.135 2.9 77.025 3.07 ;
      RECT 76.135 3.055 77.085 3.07 ;
      RECT 76.135 3.05 77.075 3.07 ;
      RECT 77.03 2.995 77.04 3.3 ;
      RECT 76.135 3.03 77.06 3.07 ;
      RECT 76.135 3.01 77.045 3.07 ;
      RECT 76.135 2.005 77.025 2.175 ;
      RECT 77.195 2.5 77.525 2.925 ;
      RECT 77.195 2.015 77.415 2.925 ;
      RECT 77.11 5.875 77.32 6.475 ;
      RECT 76.97 5.875 77.32 6.075 ;
      RECT 75.69 3.475 75.965 4.175 ;
      RECT 75.91 1.965 75.965 4.175 ;
      RECT 75.795 2.77 75.965 4.175 ;
      RECT 75.795 1.965 75.965 2.765 ;
      RECT 75.705 1.965 75.965 2.44 ;
      RECT 73.835 3.135 74.085 3.67 ;
      RECT 74.805 3.135 75.52 3.6 ;
      RECT 73.835 3.135 75.625 3.305 ;
      RECT 75.395 2.77 75.625 3.305 ;
      RECT 74.39 2.015 74.645 3.305 ;
      RECT 75.395 2.705 75.455 3.6 ;
      RECT 75.455 2.7 75.625 2.765 ;
      RECT 73.855 2.015 74.645 2.28 ;
      RECT 74.815 5.825 75.49 6.075 ;
      RECT 75.225 5.465 75.49 6.075 ;
      RECT 74.975 6.245 75.305 6.795 ;
      RECT 73.915 6.245 75.305 6.435 ;
      RECT 73.915 5.405 74.085 6.435 ;
      RECT 73.795 5.825 74.085 6.155 ;
      RECT 73.915 5.405 74.855 5.575 ;
      RECT 74.555 4.855 74.855 5.575 ;
      RECT 74.815 2.435 75.225 2.955 ;
      RECT 74.815 2.015 75.015 2.955 ;
      RECT 73.425 2.195 73.595 4.175 ;
      RECT 73.425 2.705 74.22 2.955 ;
      RECT 73.425 2.195 73.675 2.955 ;
      RECT 73.345 2.195 73.675 2.615 ;
      RECT 73.375 6.605 73.935 6.895 ;
      RECT 73.375 4.685 73.625 6.895 ;
      RECT 73.375 4.685 73.835 5.235 ;
      RECT 70.2 5.015 70.37 8.305 ;
      RECT 70.2 7.315 70.605 7.645 ;
      RECT 70.2 6.475 70.605 6.805 ;
      RECT 68.575 5.02 68.745 6.49 ;
      RECT 68.575 6.315 68.75 6.485 ;
      RECT 68.205 1.74 68.375 2.93 ;
      RECT 68.205 1.74 68.675 1.91 ;
      RECT 68.205 6.97 68.675 7.14 ;
      RECT 68.205 5.95 68.375 7.14 ;
      RECT 67.215 1.74 67.385 2.93 ;
      RECT 67.215 1.74 67.685 1.91 ;
      RECT 67.215 6.97 67.685 7.14 ;
      RECT 67.215 5.95 67.385 7.14 ;
      RECT 65.365 2.635 65.535 3.865 ;
      RECT 65.42 0.855 65.59 2.805 ;
      RECT 65.365 0.575 65.535 1.025 ;
      RECT 65.365 7.855 65.535 8.305 ;
      RECT 65.42 6.075 65.59 8.025 ;
      RECT 65.365 5.015 65.535 6.245 ;
      RECT 64.845 0.575 65.015 3.865 ;
      RECT 64.845 2.075 65.25 2.405 ;
      RECT 64.845 1.235 65.25 1.565 ;
      RECT 64.845 5.015 65.015 8.305 ;
      RECT 64.845 7.315 65.25 7.645 ;
      RECT 64.845 6.475 65.25 6.805 ;
      RECT 60.105 6.645 61.41 6.895 ;
      RECT 60.105 6.325 60.285 6.895 ;
      RECT 59.555 6.325 60.285 6.495 ;
      RECT 59.555 5.485 59.725 6.495 ;
      RECT 60.39 5.525 62.135 5.705 ;
      RECT 61.805 4.685 62.135 5.705 ;
      RECT 59.555 5.485 60.615 5.655 ;
      RECT 61.805 4.855 62.625 5.025 ;
      RECT 60.965 4.685 61.295 4.895 ;
      RECT 60.965 4.685 62.135 4.855 ;
      RECT 61.865 3.205 62.195 4.16 ;
      RECT 61.865 3.205 62.545 3.375 ;
      RECT 62.375 1.965 62.545 3.375 ;
      RECT 62.285 1.965 62.615 2.605 ;
      RECT 61.41 3.475 61.685 4.175 ;
      RECT 61.515 1.965 61.685 4.175 ;
      RECT 61.855 2.785 62.205 3.035 ;
      RECT 61.515 2.815 62.205 2.985 ;
      RECT 61.425 1.965 61.685 2.445 ;
      RECT 60.755 5.115 61.635 5.355 ;
      RECT 61.405 5.025 61.635 5.355 ;
      RECT 60.105 5.115 61.635 5.315 ;
      RECT 61.02 5.065 61.635 5.355 ;
      RECT 60.105 4.985 60.275 5.315 ;
      RECT 60.99 5.875 61.24 6.475 ;
      RECT 60.99 5.875 61.465 6.075 ;
      RECT 60.485 3.095 61.24 3.595 ;
      RECT 59.555 2.9 59.815 3.52 ;
      RECT 60.47 3.04 60.485 3.345 ;
      RECT 60.455 3.025 60.475 3.31 ;
      RECT 61.115 2.7 61.345 3.3 ;
      RECT 60.43 2.97 60.45 3.285 ;
      RECT 60.41 3.095 61.345 3.27 ;
      RECT 60.385 3.095 61.345 3.26 ;
      RECT 60.315 3.095 61.345 3.25 ;
      RECT 60.295 3.095 61.345 3.22 ;
      RECT 60.275 2.005 60.445 3.19 ;
      RECT 60.245 3.095 61.345 3.16 ;
      RECT 60.21 3.095 61.345 3.135 ;
      RECT 60.18 3.09 60.57 3.1 ;
      RECT 60.18 3.08 60.545 3.1 ;
      RECT 60.18 3.075 60.53 3.1 ;
      RECT 60.18 3.065 60.515 3.1 ;
      RECT 59.555 2.9 60.445 3.07 ;
      RECT 59.555 3.055 60.505 3.07 ;
      RECT 59.555 3.05 60.495 3.07 ;
      RECT 60.45 2.995 60.46 3.3 ;
      RECT 59.555 3.03 60.48 3.07 ;
      RECT 59.555 3.01 60.465 3.07 ;
      RECT 59.555 2.005 60.445 2.175 ;
      RECT 60.615 2.5 60.945 2.925 ;
      RECT 60.615 2.015 60.835 2.925 ;
      RECT 60.53 5.875 60.74 6.475 ;
      RECT 60.39 5.875 60.74 6.075 ;
      RECT 59.11 3.475 59.385 4.175 ;
      RECT 59.33 1.965 59.385 4.175 ;
      RECT 59.215 2.77 59.385 4.175 ;
      RECT 59.215 1.965 59.385 2.765 ;
      RECT 59.125 1.965 59.385 2.44 ;
      RECT 57.255 3.135 57.505 3.67 ;
      RECT 58.225 3.135 58.94 3.6 ;
      RECT 57.255 3.135 59.045 3.305 ;
      RECT 58.815 2.77 59.045 3.305 ;
      RECT 57.81 2.015 58.065 3.305 ;
      RECT 58.815 2.705 58.875 3.6 ;
      RECT 58.875 2.7 59.045 2.765 ;
      RECT 57.275 2.015 58.065 2.28 ;
      RECT 58.235 5.825 58.91 6.075 ;
      RECT 58.645 5.465 58.91 6.075 ;
      RECT 58.395 6.245 58.725 6.795 ;
      RECT 57.335 6.245 58.725 6.435 ;
      RECT 57.335 5.405 57.505 6.435 ;
      RECT 57.215 5.825 57.505 6.155 ;
      RECT 57.335 5.405 58.275 5.575 ;
      RECT 57.975 4.855 58.275 5.575 ;
      RECT 58.235 2.435 58.645 2.955 ;
      RECT 58.235 2.015 58.435 2.955 ;
      RECT 56.845 2.195 57.015 4.175 ;
      RECT 56.845 2.705 57.64 2.955 ;
      RECT 56.845 2.195 57.095 2.955 ;
      RECT 56.765 2.195 57.095 2.615 ;
      RECT 56.795 6.605 57.355 6.895 ;
      RECT 56.795 4.685 57.045 6.895 ;
      RECT 56.795 4.685 57.255 5.235 ;
      RECT 53.62 5.015 53.79 8.305 ;
      RECT 53.62 7.315 54.025 7.645 ;
      RECT 53.62 6.475 54.025 6.805 ;
      RECT 51.99 5.02 52.16 6.49 ;
      RECT 51.99 6.315 52.165 6.485 ;
      RECT 51.62 1.74 51.79 2.93 ;
      RECT 51.62 1.74 52.09 1.91 ;
      RECT 51.62 6.97 52.09 7.14 ;
      RECT 51.62 5.95 51.79 7.14 ;
      RECT 50.63 1.74 50.8 2.93 ;
      RECT 50.63 1.74 51.1 1.91 ;
      RECT 50.63 6.97 51.1 7.14 ;
      RECT 50.63 5.95 50.8 7.14 ;
      RECT 48.78 2.635 48.95 3.865 ;
      RECT 48.835 0.855 49.005 2.805 ;
      RECT 48.78 0.575 48.95 1.025 ;
      RECT 48.78 7.855 48.95 8.305 ;
      RECT 48.835 6.075 49.005 8.025 ;
      RECT 48.78 5.015 48.95 6.245 ;
      RECT 48.26 0.575 48.43 3.865 ;
      RECT 48.26 2.075 48.665 2.405 ;
      RECT 48.26 1.235 48.665 1.565 ;
      RECT 48.26 5.015 48.43 8.305 ;
      RECT 48.26 7.315 48.665 7.645 ;
      RECT 48.26 6.475 48.665 6.805 ;
      RECT 43.52 6.645 44.825 6.895 ;
      RECT 43.52 6.325 43.7 6.895 ;
      RECT 42.97 6.325 43.7 6.495 ;
      RECT 42.97 5.485 43.14 6.495 ;
      RECT 43.805 5.525 45.55 5.705 ;
      RECT 45.22 4.685 45.55 5.705 ;
      RECT 42.97 5.485 44.03 5.655 ;
      RECT 45.22 4.855 46.04 5.025 ;
      RECT 44.38 4.685 44.71 4.895 ;
      RECT 44.38 4.685 45.55 4.855 ;
      RECT 45.28 3.205 45.61 4.16 ;
      RECT 45.28 3.205 45.96 3.375 ;
      RECT 45.79 1.965 45.96 3.375 ;
      RECT 45.7 1.965 46.03 2.605 ;
      RECT 44.825 3.475 45.1 4.175 ;
      RECT 44.93 1.965 45.1 4.175 ;
      RECT 45.27 2.785 45.62 3.035 ;
      RECT 44.93 2.815 45.62 2.985 ;
      RECT 44.84 1.965 45.1 2.445 ;
      RECT 44.17 5.115 45.05 5.355 ;
      RECT 44.82 5.025 45.05 5.355 ;
      RECT 43.52 5.115 45.05 5.315 ;
      RECT 44.435 5.065 45.05 5.355 ;
      RECT 43.52 4.985 43.69 5.315 ;
      RECT 44.405 5.875 44.655 6.475 ;
      RECT 44.405 5.875 44.88 6.075 ;
      RECT 43.9 3.095 44.655 3.595 ;
      RECT 42.97 2.9 43.23 3.52 ;
      RECT 43.885 3.04 43.9 3.345 ;
      RECT 43.87 3.025 43.89 3.31 ;
      RECT 44.53 2.7 44.76 3.3 ;
      RECT 43.845 2.97 43.865 3.285 ;
      RECT 43.825 3.095 44.76 3.27 ;
      RECT 43.8 3.095 44.76 3.26 ;
      RECT 43.73 3.095 44.76 3.25 ;
      RECT 43.71 3.095 44.76 3.22 ;
      RECT 43.69 2.005 43.86 3.19 ;
      RECT 43.66 3.095 44.76 3.16 ;
      RECT 43.625 3.095 44.76 3.135 ;
      RECT 43.595 3.09 43.985 3.1 ;
      RECT 43.595 3.08 43.96 3.1 ;
      RECT 43.595 3.075 43.945 3.1 ;
      RECT 43.595 3.065 43.93 3.1 ;
      RECT 42.97 2.9 43.86 3.07 ;
      RECT 42.97 3.055 43.92 3.07 ;
      RECT 42.97 3.05 43.91 3.07 ;
      RECT 43.865 2.995 43.875 3.3 ;
      RECT 42.97 3.03 43.895 3.07 ;
      RECT 42.97 3.01 43.88 3.07 ;
      RECT 42.97 2.005 43.86 2.175 ;
      RECT 44.03 2.5 44.36 2.925 ;
      RECT 44.03 2.015 44.25 2.925 ;
      RECT 43.945 5.875 44.155 6.475 ;
      RECT 43.805 5.875 44.155 6.075 ;
      RECT 42.525 3.475 42.8 4.175 ;
      RECT 42.745 1.965 42.8 4.175 ;
      RECT 42.63 2.77 42.8 4.175 ;
      RECT 42.63 1.965 42.8 2.765 ;
      RECT 42.54 1.965 42.8 2.44 ;
      RECT 40.67 3.135 40.92 3.67 ;
      RECT 41.64 3.135 42.355 3.6 ;
      RECT 40.67 3.135 42.46 3.305 ;
      RECT 42.23 2.77 42.46 3.305 ;
      RECT 41.225 2.015 41.48 3.305 ;
      RECT 42.23 2.705 42.29 3.6 ;
      RECT 42.29 2.7 42.46 2.765 ;
      RECT 40.69 2.015 41.48 2.28 ;
      RECT 41.65 5.825 42.325 6.075 ;
      RECT 42.06 5.465 42.325 6.075 ;
      RECT 41.81 6.245 42.14 6.795 ;
      RECT 40.75 6.245 42.14 6.435 ;
      RECT 40.75 5.405 40.92 6.435 ;
      RECT 40.63 5.825 40.92 6.155 ;
      RECT 40.75 5.405 41.69 5.575 ;
      RECT 41.39 4.855 41.69 5.575 ;
      RECT 41.65 2.435 42.06 2.955 ;
      RECT 41.65 2.015 41.85 2.955 ;
      RECT 40.26 2.195 40.43 4.175 ;
      RECT 40.26 2.705 41.055 2.955 ;
      RECT 40.26 2.195 40.51 2.955 ;
      RECT 40.18 2.195 40.51 2.615 ;
      RECT 40.21 6.605 40.77 6.895 ;
      RECT 40.21 4.685 40.46 6.895 ;
      RECT 40.21 4.685 40.67 5.235 ;
      RECT 37.035 5.015 37.205 8.305 ;
      RECT 37.035 7.315 37.44 7.645 ;
      RECT 37.035 6.475 37.44 6.805 ;
      RECT 35.405 5.02 35.575 6.49 ;
      RECT 35.405 6.315 35.58 6.485 ;
      RECT 35.035 1.74 35.205 2.93 ;
      RECT 35.035 1.74 35.505 1.91 ;
      RECT 35.035 6.97 35.505 7.14 ;
      RECT 35.035 5.95 35.205 7.14 ;
      RECT 34.045 1.74 34.215 2.93 ;
      RECT 34.045 1.74 34.515 1.91 ;
      RECT 34.045 6.97 34.515 7.14 ;
      RECT 34.045 5.95 34.215 7.14 ;
      RECT 32.195 2.635 32.365 3.865 ;
      RECT 32.25 0.855 32.42 2.805 ;
      RECT 32.195 0.575 32.365 1.025 ;
      RECT 32.195 7.855 32.365 8.305 ;
      RECT 32.25 6.075 32.42 8.025 ;
      RECT 32.195 5.015 32.365 6.245 ;
      RECT 31.675 0.575 31.845 3.865 ;
      RECT 31.675 2.075 32.08 2.405 ;
      RECT 31.675 1.235 32.08 1.565 ;
      RECT 31.675 5.015 31.845 8.305 ;
      RECT 31.675 7.315 32.08 7.645 ;
      RECT 31.675 6.475 32.08 6.805 ;
      RECT 26.935 6.645 28.24 6.895 ;
      RECT 26.935 6.325 27.115 6.895 ;
      RECT 26.385 6.325 27.115 6.495 ;
      RECT 26.385 5.485 26.555 6.495 ;
      RECT 27.22 5.525 28.965 5.705 ;
      RECT 28.635 4.685 28.965 5.705 ;
      RECT 26.385 5.485 27.445 5.655 ;
      RECT 28.635 4.855 29.455 5.025 ;
      RECT 27.795 4.685 28.125 4.895 ;
      RECT 27.795 4.685 28.965 4.855 ;
      RECT 28.695 3.205 29.025 4.16 ;
      RECT 28.695 3.205 29.375 3.375 ;
      RECT 29.205 1.965 29.375 3.375 ;
      RECT 29.115 1.965 29.445 2.605 ;
      RECT 28.24 3.475 28.515 4.175 ;
      RECT 28.345 1.965 28.515 4.175 ;
      RECT 28.685 2.785 29.035 3.035 ;
      RECT 28.345 2.815 29.035 2.985 ;
      RECT 28.255 1.965 28.515 2.445 ;
      RECT 27.585 5.115 28.465 5.355 ;
      RECT 28.235 5.025 28.465 5.355 ;
      RECT 26.935 5.115 28.465 5.315 ;
      RECT 27.85 5.065 28.465 5.355 ;
      RECT 26.935 4.985 27.105 5.315 ;
      RECT 27.82 5.875 28.07 6.475 ;
      RECT 27.82 5.875 28.295 6.075 ;
      RECT 27.315 3.095 28.07 3.595 ;
      RECT 26.385 2.9 26.645 3.52 ;
      RECT 27.3 3.04 27.315 3.345 ;
      RECT 27.285 3.025 27.305 3.31 ;
      RECT 27.945 2.7 28.175 3.3 ;
      RECT 27.26 2.97 27.28 3.285 ;
      RECT 27.24 3.095 28.175 3.27 ;
      RECT 27.215 3.095 28.175 3.26 ;
      RECT 27.145 3.095 28.175 3.25 ;
      RECT 27.125 3.095 28.175 3.22 ;
      RECT 27.105 2.005 27.275 3.19 ;
      RECT 27.075 3.095 28.175 3.16 ;
      RECT 27.04 3.095 28.175 3.135 ;
      RECT 27.01 3.09 27.4 3.1 ;
      RECT 27.01 3.08 27.375 3.1 ;
      RECT 27.01 3.075 27.36 3.1 ;
      RECT 27.01 3.065 27.345 3.1 ;
      RECT 26.385 2.9 27.275 3.07 ;
      RECT 26.385 3.055 27.335 3.07 ;
      RECT 26.385 3.05 27.325 3.07 ;
      RECT 27.28 2.995 27.29 3.3 ;
      RECT 26.385 3.03 27.31 3.07 ;
      RECT 26.385 3.01 27.295 3.07 ;
      RECT 26.385 2.005 27.275 2.175 ;
      RECT 27.445 2.5 27.775 2.925 ;
      RECT 27.445 2.015 27.665 2.925 ;
      RECT 27.36 5.875 27.57 6.475 ;
      RECT 27.22 5.875 27.57 6.075 ;
      RECT 25.94 3.475 26.215 4.175 ;
      RECT 26.16 1.965 26.215 4.175 ;
      RECT 26.045 2.77 26.215 4.175 ;
      RECT 26.045 1.965 26.215 2.765 ;
      RECT 25.955 1.965 26.215 2.44 ;
      RECT 24.085 3.135 24.335 3.67 ;
      RECT 25.055 3.135 25.77 3.6 ;
      RECT 24.085 3.135 25.875 3.305 ;
      RECT 25.645 2.77 25.875 3.305 ;
      RECT 24.64 2.015 24.895 3.305 ;
      RECT 25.645 2.705 25.705 3.6 ;
      RECT 25.705 2.7 25.875 2.765 ;
      RECT 24.105 2.015 24.895 2.28 ;
      RECT 25.065 5.825 25.74 6.075 ;
      RECT 25.475 5.465 25.74 6.075 ;
      RECT 25.225 6.245 25.555 6.795 ;
      RECT 24.165 6.245 25.555 6.435 ;
      RECT 24.165 5.405 24.335 6.435 ;
      RECT 24.045 5.825 24.335 6.155 ;
      RECT 24.165 5.405 25.105 5.575 ;
      RECT 24.805 4.855 25.105 5.575 ;
      RECT 25.065 2.435 25.475 2.955 ;
      RECT 25.065 2.015 25.265 2.955 ;
      RECT 23.675 2.195 23.845 4.175 ;
      RECT 23.675 2.705 24.47 2.955 ;
      RECT 23.675 2.195 23.925 2.955 ;
      RECT 23.595 2.195 23.925 2.615 ;
      RECT 23.625 6.605 24.185 6.895 ;
      RECT 23.625 4.685 23.875 6.895 ;
      RECT 23.625 4.685 24.085 5.235 ;
      RECT 20.45 5.015 20.62 8.305 ;
      RECT 20.45 7.315 20.855 7.645 ;
      RECT 20.45 6.475 20.855 6.805 ;
      RECT 18.82 5.02 18.99 6.49 ;
      RECT 18.82 6.315 18.995 6.485 ;
      RECT 18.45 1.74 18.62 2.93 ;
      RECT 18.45 1.74 18.92 1.91 ;
      RECT 18.45 6.97 18.92 7.14 ;
      RECT 18.45 5.95 18.62 7.14 ;
      RECT 17.46 1.74 17.63 2.93 ;
      RECT 17.46 1.74 17.93 1.91 ;
      RECT 17.46 6.97 17.93 7.14 ;
      RECT 17.46 5.95 17.63 7.14 ;
      RECT 15.61 2.635 15.78 3.865 ;
      RECT 15.665 0.855 15.835 2.805 ;
      RECT 15.61 0.575 15.78 1.025 ;
      RECT 15.61 7.855 15.78 8.305 ;
      RECT 15.665 6.075 15.835 8.025 ;
      RECT 15.61 5.015 15.78 6.245 ;
      RECT 15.09 0.575 15.26 3.865 ;
      RECT 15.09 2.075 15.495 2.405 ;
      RECT 15.09 1.235 15.495 1.565 ;
      RECT 15.09 5.015 15.26 8.305 ;
      RECT 15.09 7.315 15.495 7.645 ;
      RECT 15.09 6.475 15.495 6.805 ;
      RECT 10.35 6.645 11.655 6.895 ;
      RECT 10.35 6.325 10.53 6.895 ;
      RECT 9.8 6.325 10.53 6.495 ;
      RECT 9.8 5.485 9.97 6.495 ;
      RECT 10.635 5.525 12.38 5.705 ;
      RECT 12.05 4.685 12.38 5.705 ;
      RECT 9.8 5.485 10.86 5.655 ;
      RECT 12.05 4.855 12.87 5.025 ;
      RECT 11.21 4.685 11.54 4.895 ;
      RECT 11.21 4.685 12.38 4.855 ;
      RECT 12.11 3.205 12.44 4.16 ;
      RECT 12.11 3.205 12.79 3.375 ;
      RECT 12.62 1.965 12.79 3.375 ;
      RECT 12.53 1.965 12.86 2.605 ;
      RECT 11.655 3.475 11.93 4.175 ;
      RECT 11.76 1.965 11.93 4.175 ;
      RECT 12.1 2.785 12.45 3.035 ;
      RECT 11.76 2.815 12.45 2.985 ;
      RECT 11.67 1.965 11.93 2.445 ;
      RECT 11 5.115 11.88 5.355 ;
      RECT 11.65 5.025 11.88 5.355 ;
      RECT 10.35 5.115 11.88 5.315 ;
      RECT 11.265 5.065 11.88 5.355 ;
      RECT 10.35 4.985 10.52 5.315 ;
      RECT 11.235 5.875 11.485 6.475 ;
      RECT 11.235 5.875 11.71 6.075 ;
      RECT 10.73 3.095 11.485 3.595 ;
      RECT 9.8 2.9 10.06 3.52 ;
      RECT 10.715 3.04 10.73 3.345 ;
      RECT 10.7 3.025 10.72 3.31 ;
      RECT 11.36 2.7 11.59 3.3 ;
      RECT 10.675 2.97 10.695 3.285 ;
      RECT 10.655 3.095 11.59 3.27 ;
      RECT 10.63 3.095 11.59 3.26 ;
      RECT 10.56 3.095 11.59 3.25 ;
      RECT 10.54 3.095 11.59 3.22 ;
      RECT 10.52 2.005 10.69 3.19 ;
      RECT 10.49 3.095 11.59 3.16 ;
      RECT 10.455 3.095 11.59 3.135 ;
      RECT 10.425 3.09 10.815 3.1 ;
      RECT 10.425 3.08 10.79 3.1 ;
      RECT 10.425 3.075 10.775 3.1 ;
      RECT 10.425 3.065 10.76 3.1 ;
      RECT 9.8 2.9 10.69 3.07 ;
      RECT 9.8 3.055 10.75 3.07 ;
      RECT 9.8 3.05 10.74 3.07 ;
      RECT 10.695 2.995 10.705 3.3 ;
      RECT 9.8 3.03 10.725 3.07 ;
      RECT 9.8 3.01 10.71 3.07 ;
      RECT 9.8 2.005 10.69 2.175 ;
      RECT 10.86 2.5 11.19 2.925 ;
      RECT 10.86 2.015 11.08 2.925 ;
      RECT 10.775 5.875 10.985 6.475 ;
      RECT 10.635 5.875 10.985 6.075 ;
      RECT 9.355 3.475 9.63 4.175 ;
      RECT 9.575 1.965 9.63 4.175 ;
      RECT 9.46 2.77 9.63 4.175 ;
      RECT 9.46 1.965 9.63 2.765 ;
      RECT 9.37 1.965 9.63 2.44 ;
      RECT 7.5 3.135 7.75 3.67 ;
      RECT 8.47 3.135 9.185 3.6 ;
      RECT 7.5 3.135 9.29 3.305 ;
      RECT 9.06 2.77 9.29 3.305 ;
      RECT 8.055 2.015 8.31 3.305 ;
      RECT 9.06 2.705 9.12 3.6 ;
      RECT 9.12 2.7 9.29 2.765 ;
      RECT 7.52 2.015 8.31 2.28 ;
      RECT 8.48 5.825 9.155 6.075 ;
      RECT 8.89 5.465 9.155 6.075 ;
      RECT 8.64 6.245 8.97 6.795 ;
      RECT 7.58 6.245 8.97 6.435 ;
      RECT 7.58 5.405 7.75 6.435 ;
      RECT 7.46 5.825 7.75 6.155 ;
      RECT 7.58 5.405 8.52 5.575 ;
      RECT 8.22 4.855 8.52 5.575 ;
      RECT 8.48 2.435 8.89 2.955 ;
      RECT 8.48 2.015 8.68 2.955 ;
      RECT 7.09 2.195 7.26 4.175 ;
      RECT 7.09 2.705 7.885 2.955 ;
      RECT 7.09 2.195 7.34 2.955 ;
      RECT 7.01 2.195 7.34 2.615 ;
      RECT 7.04 6.605 7.6 6.895 ;
      RECT 7.04 4.685 7.29 6.895 ;
      RECT 7.04 4.685 7.5 5.235 ;
      RECT 3.865 5.015 4.035 8.305 ;
      RECT 3.865 7.315 4.27 7.645 ;
      RECT 3.865 6.475 4.27 6.805 ;
      RECT 1.155 7.855 1.325 8.305 ;
      RECT 1.21 6.075 1.38 8.025 ;
      RECT 1.155 5.015 1.325 6.245 ;
      RECT 0.635 5.015 0.805 8.305 ;
      RECT 0.635 7.315 1.04 7.645 ;
      RECT 0.635 6.475 1.04 6.805 ;
      RECT 85.155 7.8 85.325 8.31 ;
      RECT 84.165 0.57 84.335 1.08 ;
      RECT 84.165 2.39 84.335 3.86 ;
      RECT 84.165 5.02 84.335 6.49 ;
      RECT 84.165 7.8 84.335 8.31 ;
      RECT 82.805 0.575 82.975 3.865 ;
      RECT 82.805 5.015 82.975 8.305 ;
      RECT 82.375 0.575 82.545 1.085 ;
      RECT 82.375 1.655 82.545 3.865 ;
      RECT 82.375 5.015 82.545 7.225 ;
      RECT 82.375 7.795 82.545 8.305 ;
      RECT 79.295 2.785 79.645 3.035 ;
      RECT 78.235 5.875 78.685 6.385 ;
      RECT 76.915 3.835 77.395 4.175 ;
      RECT 76.135 2.345 76.685 2.73 ;
      RECT 74.62 3.835 75.095 4.175 ;
      RECT 72.915 2.785 73.255 3.665 ;
      RECT 71.58 5.015 71.75 8.305 ;
      RECT 71.15 5.015 71.32 7.225 ;
      RECT 71.15 7.795 71.32 8.305 ;
      RECT 68.575 7.8 68.745 8.31 ;
      RECT 67.585 0.57 67.755 1.08 ;
      RECT 67.585 2.39 67.755 3.86 ;
      RECT 67.585 5.02 67.755 6.49 ;
      RECT 67.585 7.8 67.755 8.31 ;
      RECT 66.225 0.575 66.395 3.865 ;
      RECT 66.225 5.015 66.395 8.305 ;
      RECT 65.795 0.575 65.965 1.085 ;
      RECT 65.795 1.655 65.965 3.865 ;
      RECT 65.795 5.015 65.965 7.225 ;
      RECT 65.795 7.795 65.965 8.305 ;
      RECT 62.715 2.785 63.065 3.035 ;
      RECT 61.655 5.875 62.105 6.385 ;
      RECT 60.335 3.835 60.815 4.175 ;
      RECT 59.555 2.345 60.105 2.73 ;
      RECT 58.04 3.835 58.515 4.175 ;
      RECT 56.335 2.785 56.675 3.665 ;
      RECT 55 5.015 55.17 8.305 ;
      RECT 54.57 5.015 54.74 7.225 ;
      RECT 54.57 7.795 54.74 8.305 ;
      RECT 51.99 7.8 52.16 8.31 ;
      RECT 51 0.57 51.17 1.08 ;
      RECT 51 2.39 51.17 3.86 ;
      RECT 51 5.02 51.17 6.49 ;
      RECT 51 7.8 51.17 8.31 ;
      RECT 49.64 0.575 49.81 3.865 ;
      RECT 49.64 5.015 49.81 8.305 ;
      RECT 49.21 0.575 49.38 1.085 ;
      RECT 49.21 1.655 49.38 3.865 ;
      RECT 49.21 5.015 49.38 7.225 ;
      RECT 49.21 7.795 49.38 8.305 ;
      RECT 46.13 2.785 46.48 3.035 ;
      RECT 45.07 5.875 45.52 6.385 ;
      RECT 43.75 3.835 44.23 4.175 ;
      RECT 42.97 2.345 43.52 2.73 ;
      RECT 41.455 3.835 41.93 4.175 ;
      RECT 39.75 2.785 40.09 3.665 ;
      RECT 38.415 5.015 38.585 8.305 ;
      RECT 37.985 5.015 38.155 7.225 ;
      RECT 37.985 7.795 38.155 8.305 ;
      RECT 35.405 7.8 35.575 8.31 ;
      RECT 34.415 0.57 34.585 1.08 ;
      RECT 34.415 2.39 34.585 3.86 ;
      RECT 34.415 5.02 34.585 6.49 ;
      RECT 34.415 7.8 34.585 8.31 ;
      RECT 33.055 0.575 33.225 3.865 ;
      RECT 33.055 5.015 33.225 8.305 ;
      RECT 32.625 0.575 32.795 1.085 ;
      RECT 32.625 1.655 32.795 3.865 ;
      RECT 32.625 5.015 32.795 7.225 ;
      RECT 32.625 7.795 32.795 8.305 ;
      RECT 29.545 2.785 29.895 3.035 ;
      RECT 28.485 5.875 28.935 6.385 ;
      RECT 27.165 3.835 27.645 4.175 ;
      RECT 26.385 2.345 26.935 2.73 ;
      RECT 24.87 3.835 25.345 4.175 ;
      RECT 23.165 2.785 23.505 3.665 ;
      RECT 21.83 5.015 22 8.305 ;
      RECT 21.4 5.015 21.57 7.225 ;
      RECT 21.4 7.795 21.57 8.305 ;
      RECT 18.82 7.8 18.99 8.31 ;
      RECT 17.83 0.57 18 1.08 ;
      RECT 17.83 2.39 18 3.86 ;
      RECT 17.83 5.02 18 6.49 ;
      RECT 17.83 7.8 18 8.31 ;
      RECT 16.47 0.575 16.64 3.865 ;
      RECT 16.47 5.015 16.64 8.305 ;
      RECT 16.04 0.575 16.21 1.085 ;
      RECT 16.04 1.655 16.21 3.865 ;
      RECT 16.04 5.015 16.21 7.225 ;
      RECT 16.04 7.795 16.21 8.305 ;
      RECT 12.96 2.785 13.31 3.035 ;
      RECT 11.9 5.875 12.35 6.385 ;
      RECT 10.58 3.835 11.06 4.175 ;
      RECT 9.8 2.345 10.35 2.73 ;
      RECT 8.285 3.835 8.76 4.175 ;
      RECT 6.58 2.785 6.92 3.665 ;
      RECT 5.245 5.015 5.415 8.305 ;
      RECT 4.815 5.015 4.985 7.225 ;
      RECT 4.815 7.795 4.985 8.305 ;
      RECT 1.585 5.015 1.755 7.225 ;
      RECT 1.585 7.795 1.755 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2ca_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2ca_8_b0r2
  CLASS BLOCK ;
  ORIGIN 2.955 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ca_8_b0r2 ;
  SIZE 85.88 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 16.05 0.915 16.22 1.085 ;
        RECT 16.045 0.91 16.215 1.08 ;
        RECT 16.05 2.395 16.22 2.565 ;
        RECT 16.045 2.39 16.215 2.56 ;
      LAYER li1 ;
        RECT 16.05 0.915 16.22 1.085 ;
        RECT 16.045 0.57 16.215 1.08 ;
        RECT 16.045 2.395 16.22 2.565 ;
        RECT 16.045 2.39 16.215 3.86 ;
      LAYER met1 ;
        RECT 15.985 2.36 16.275 2.59 ;
        RECT 15.985 0.88 16.275 1.11 ;
        RECT 16.045 0.88 16.215 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 32.635 0.915 32.805 1.085 ;
        RECT 32.63 0.91 32.8 1.08 ;
        RECT 32.635 2.395 32.805 2.565 ;
        RECT 32.63 2.39 32.8 2.56 ;
      LAYER li1 ;
        RECT 32.635 0.915 32.805 1.085 ;
        RECT 32.63 0.57 32.8 1.08 ;
        RECT 32.63 2.395 32.805 2.565 ;
        RECT 32.63 2.39 32.8 3.86 ;
      LAYER met1 ;
        RECT 32.57 2.36 32.86 2.59 ;
        RECT 32.57 0.88 32.86 1.11 ;
        RECT 32.63 0.88 32.8 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 49.22 0.915 49.39 1.085 ;
        RECT 49.215 0.91 49.385 1.08 ;
        RECT 49.22 2.395 49.39 2.565 ;
        RECT 49.215 2.39 49.385 2.56 ;
      LAYER li1 ;
        RECT 49.22 0.915 49.39 1.085 ;
        RECT 49.215 0.57 49.385 1.08 ;
        RECT 49.215 2.395 49.39 2.565 ;
        RECT 49.215 2.39 49.385 3.86 ;
      LAYER met1 ;
        RECT 49.155 2.36 49.445 2.59 ;
        RECT 49.155 0.88 49.445 1.11 ;
        RECT 49.215 0.88 49.385 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 65.805 0.915 65.975 1.085 ;
        RECT 65.8 0.91 65.97 1.08 ;
        RECT 65.805 2.395 65.975 2.565 ;
        RECT 65.8 2.39 65.97 2.56 ;
      LAYER li1 ;
        RECT 65.805 0.915 65.975 1.085 ;
        RECT 65.8 0.57 65.97 1.08 ;
        RECT 65.8 2.395 65.975 2.565 ;
        RECT 65.8 2.39 65.97 3.86 ;
      LAYER met1 ;
        RECT 65.74 2.36 66.03 2.59 ;
        RECT 65.74 0.88 66.03 1.11 ;
        RECT 65.8 0.88 65.97 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 82.385 0.915 82.555 1.085 ;
        RECT 82.38 0.91 82.55 1.08 ;
        RECT 82.385 2.395 82.555 2.565 ;
        RECT 82.38 2.39 82.55 2.56 ;
      LAYER li1 ;
        RECT 82.385 0.915 82.555 1.085 ;
        RECT 82.38 0.57 82.55 1.08 ;
        RECT 82.38 2.395 82.555 2.565 ;
        RECT 82.38 2.39 82.55 3.86 ;
      LAYER met1 ;
        RECT 82.32 2.36 82.61 2.59 ;
        RECT 82.32 0.88 82.61 1.11 ;
        RECT 82.38 0.88 82.55 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 11.895 1.66 12.065 2.935 ;
        RECT 11.895 5.945 12.065 7.22 ;
        RECT 0.67 5.945 0.84 7.22 ;
      LAYER met2 ;
        RECT 11.82 5.865 12.145 6.19 ;
        RECT 11.815 3.635 12.14 3.96 ;
        RECT 2.975 7.885 12.06 8.055 ;
        RECT 11.885 3.635 12.06 8.055 ;
        RECT 2.92 5.86 3.2 6.2 ;
        RECT 2.975 5.86 3.145 8.055 ;
      LAYER met1 ;
        RECT 11.835 2.765 12.295 2.935 ;
        RECT 11.815 3.635 12.14 3.96 ;
        RECT 11.835 2.735 12.125 2.965 ;
        RECT 11.89 2.735 12.07 3.96 ;
        RECT 11.82 5.945 12.295 6.115 ;
        RECT 11.82 5.865 12.145 6.19 ;
        RECT 2.89 5.89 3.23 6.17 ;
        RECT 0.61 5.945 3.23 6.115 ;
        RECT 0.61 5.915 0.9 6.145 ;
      LAYER via1 ;
        RECT 2.985 5.955 3.135 6.105 ;
        RECT 11.905 3.72 12.055 3.87 ;
        RECT 11.91 5.95 12.06 6.1 ;
      LAYER mcon ;
        RECT 0.67 5.945 0.84 6.115 ;
        RECT 11.895 5.945 12.065 6.115 ;
        RECT 11.895 2.765 12.065 2.935 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 28.48 1.66 28.65 2.935 ;
        RECT 28.48 5.945 28.65 7.22 ;
        RECT 17.255 5.945 17.425 7.22 ;
      LAYER met2 ;
        RECT 28.405 5.865 28.73 6.19 ;
        RECT 28.4 3.635 28.725 3.96 ;
        RECT 19.56 7.885 28.645 8.055 ;
        RECT 28.47 3.635 28.645 8.055 ;
        RECT 19.505 5.86 19.785 6.2 ;
        RECT 19.56 5.86 19.73 8.055 ;
      LAYER met1 ;
        RECT 28.42 2.765 28.88 2.935 ;
        RECT 28.4 3.635 28.725 3.96 ;
        RECT 28.42 2.735 28.71 2.965 ;
        RECT 28.475 2.735 28.655 3.96 ;
        RECT 28.405 5.945 28.88 6.115 ;
        RECT 28.405 5.865 28.73 6.19 ;
        RECT 19.475 5.89 19.815 6.17 ;
        RECT 17.195 5.945 19.815 6.115 ;
        RECT 17.195 5.915 17.485 6.145 ;
      LAYER via1 ;
        RECT 19.57 5.955 19.72 6.105 ;
        RECT 28.49 3.72 28.64 3.87 ;
        RECT 28.495 5.95 28.645 6.1 ;
      LAYER mcon ;
        RECT 17.255 5.945 17.425 6.115 ;
        RECT 28.48 5.945 28.65 6.115 ;
        RECT 28.48 2.765 28.65 2.935 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 45.065 1.66 45.235 2.935 ;
        RECT 45.065 5.945 45.235 7.22 ;
        RECT 33.84 5.945 34.01 7.22 ;
      LAYER met2 ;
        RECT 44.99 5.865 45.315 6.19 ;
        RECT 44.985 3.635 45.31 3.96 ;
        RECT 36.145 7.885 45.23 8.055 ;
        RECT 45.055 3.635 45.23 8.055 ;
        RECT 36.09 5.86 36.37 6.2 ;
        RECT 36.145 5.86 36.315 8.055 ;
      LAYER met1 ;
        RECT 45.005 2.765 45.465 2.935 ;
        RECT 44.985 3.635 45.31 3.96 ;
        RECT 45.005 2.735 45.295 2.965 ;
        RECT 45.06 2.735 45.24 3.96 ;
        RECT 44.99 5.945 45.465 6.115 ;
        RECT 44.99 5.865 45.315 6.19 ;
        RECT 36.06 5.89 36.4 6.17 ;
        RECT 33.78 5.945 36.4 6.115 ;
        RECT 33.78 5.915 34.07 6.145 ;
      LAYER via1 ;
        RECT 36.155 5.955 36.305 6.105 ;
        RECT 45.075 3.72 45.225 3.87 ;
        RECT 45.08 5.95 45.23 6.1 ;
      LAYER mcon ;
        RECT 33.84 5.945 34.01 6.115 ;
        RECT 45.065 5.945 45.235 6.115 ;
        RECT 45.065 2.765 45.235 2.935 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 61.65 1.66 61.82 2.935 ;
        RECT 61.65 5.945 61.82 7.22 ;
        RECT 50.425 5.945 50.595 7.22 ;
      LAYER met2 ;
        RECT 61.575 5.865 61.9 6.19 ;
        RECT 61.57 3.635 61.895 3.96 ;
        RECT 52.73 7.885 61.815 8.055 ;
        RECT 61.64 3.635 61.815 8.055 ;
        RECT 52.675 5.86 52.955 6.2 ;
        RECT 52.73 5.86 52.9 8.055 ;
      LAYER met1 ;
        RECT 61.59 2.765 62.05 2.935 ;
        RECT 61.57 3.635 61.895 3.96 ;
        RECT 61.59 2.735 61.88 2.965 ;
        RECT 61.645 2.735 61.825 3.96 ;
        RECT 61.575 5.945 62.05 6.115 ;
        RECT 61.575 5.865 61.9 6.19 ;
        RECT 52.645 5.89 52.985 6.17 ;
        RECT 50.365 5.945 52.985 6.115 ;
        RECT 50.365 5.915 50.655 6.145 ;
      LAYER via1 ;
        RECT 52.74 5.955 52.89 6.105 ;
        RECT 61.66 3.72 61.81 3.87 ;
        RECT 61.665 5.95 61.815 6.1 ;
      LAYER mcon ;
        RECT 50.425 5.945 50.595 6.115 ;
        RECT 61.65 5.945 61.82 6.115 ;
        RECT 61.65 2.765 61.82 2.935 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 78.23 1.66 78.4 2.935 ;
        RECT 78.23 5.945 78.4 7.22 ;
        RECT 67.005 5.945 67.175 7.22 ;
      LAYER met2 ;
        RECT 78.155 5.865 78.48 6.19 ;
        RECT 78.15 3.635 78.475 3.96 ;
        RECT 69.31 7.885 78.395 8.055 ;
        RECT 78.22 3.635 78.395 8.055 ;
        RECT 69.255 5.86 69.535 6.2 ;
        RECT 69.31 5.86 69.48 8.055 ;
      LAYER met1 ;
        RECT 78.17 2.765 78.63 2.935 ;
        RECT 78.15 3.635 78.475 3.96 ;
        RECT 78.17 2.735 78.46 2.965 ;
        RECT 78.225 2.735 78.405 3.96 ;
        RECT 78.155 5.945 78.63 6.115 ;
        RECT 78.155 5.865 78.48 6.19 ;
        RECT 69.225 5.89 69.565 6.17 ;
        RECT 66.945 5.945 69.565 6.115 ;
        RECT 66.945 5.915 67.235 6.145 ;
      LAYER via1 ;
        RECT 69.32 5.955 69.47 6.105 ;
        RECT 78.24 3.72 78.39 3.87 ;
        RECT 78.245 5.95 78.395 6.1 ;
      LAYER mcon ;
        RECT 67.005 5.945 67.175 6.115 ;
        RECT 78.23 5.945 78.4 6.115 ;
        RECT 78.23 2.765 78.4 2.935 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT -2.56 5.945 -2.39 7.22 ;
      LAYER met1 ;
        RECT -2.62 5.945 -2.16 6.115 ;
        RECT -2.62 5.915 -2.33 6.145 ;
      LAYER mcon ;
        RECT -2.56 5.945 -2.39 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 76.985 4.135 82.925 4.745 ;
        RECT 80.79 4.13 82.77 4.75 ;
        RECT 81.95 3.4 82.12 5.48 ;
        RECT 80.96 3.4 81.13 5.48 ;
        RECT 78.22 3.405 78.39 5.475 ;
        RECT 76.855 4.135 82.925 4.67 ;
        RECT 76.53 3.205 76.86 4.515 ;
        RECT -2.955 4.345 82.925 4.515 ;
        RECT 74.79 3.8 75.045 4.515 ;
        RECT 74.225 4.345 74.6 4.895 ;
        RECT 73.79 3.42 74.12 3.665 ;
        RECT 73.79 3.42 73.975 3.79 ;
        RECT 73.36 3.69 73.965 4.515 ;
        RECT 73.41 3.69 73.675 5.295 ;
        RECT 72.49 3.8 72.705 4.515 ;
        RECT 72.25 4.345 72.53 5.185 ;
        RECT 71.48 3.475 71.81 3.665 ;
        RECT 71.06 3.84 71.675 4.515 ;
        RECT 71.48 3.475 71.675 4.515 ;
        RECT 71.25 3.84 71.58 5.235 ;
        RECT 70.14 3.835 70.4 4.515 ;
        RECT 66.34 4.13 69.915 4.74 ;
        RECT 66.82 4.13 69.57 4.745 ;
        RECT 66.995 4.13 67.165 5.475 ;
        RECT 60.405 4.135 66.345 4.745 ;
        RECT 64.21 4.13 66.19 4.75 ;
        RECT 65.37 3.4 65.54 5.48 ;
        RECT 64.38 3.4 64.55 5.48 ;
        RECT 61.64 3.405 61.81 5.475 ;
        RECT 60.275 4.135 69.915 4.67 ;
        RECT 59.95 3.205 60.28 4.515 ;
        RECT 58.21 3.8 58.465 4.515 ;
        RECT 57.645 4.345 58.02 4.895 ;
        RECT 57.21 3.42 57.54 3.665 ;
        RECT 57.21 3.42 57.395 3.79 ;
        RECT 56.78 3.69 57.385 4.515 ;
        RECT 56.83 3.69 57.095 5.295 ;
        RECT 55.91 3.8 56.125 4.515 ;
        RECT 55.67 4.345 55.95 5.185 ;
        RECT 54.9 3.475 55.23 3.665 ;
        RECT 54.48 3.84 55.095 4.515 ;
        RECT 54.9 3.475 55.095 4.515 ;
        RECT 54.67 3.84 55 5.235 ;
        RECT 53.56 3.835 53.82 4.515 ;
        RECT 49.76 4.13 53.335 4.74 ;
        RECT 50.24 4.13 52.99 4.745 ;
        RECT 50.415 4.13 50.585 5.475 ;
        RECT 43.82 4.135 49.76 4.745 ;
        RECT 47.625 4.13 49.605 4.75 ;
        RECT 48.785 3.4 48.955 5.48 ;
        RECT 47.795 3.4 47.965 5.48 ;
        RECT 45.055 3.405 45.225 5.475 ;
        RECT 43.69 4.135 53.335 4.67 ;
        RECT 43.365 3.205 43.695 4.515 ;
        RECT 41.625 3.8 41.88 4.515 ;
        RECT 41.06 4.345 41.435 4.895 ;
        RECT 40.625 3.42 40.955 3.665 ;
        RECT 40.625 3.42 40.81 3.79 ;
        RECT 40.195 3.69 40.8 4.515 ;
        RECT 40.245 3.69 40.51 5.295 ;
        RECT 39.325 3.8 39.54 4.515 ;
        RECT 39.085 4.345 39.365 5.185 ;
        RECT 38.315 3.475 38.645 3.665 ;
        RECT 37.895 3.84 38.51 4.515 ;
        RECT 38.315 3.475 38.51 4.515 ;
        RECT 38.085 3.84 38.415 5.235 ;
        RECT 36.975 3.835 37.235 4.515 ;
        RECT 33.175 4.13 36.75 4.74 ;
        RECT 33.655 4.13 36.405 4.745 ;
        RECT 33.83 4.13 34 5.475 ;
        RECT 27.235 4.135 33.175 4.745 ;
        RECT 31.04 4.13 33.02 4.75 ;
        RECT 32.2 3.4 32.37 5.48 ;
        RECT 31.21 3.4 31.38 5.48 ;
        RECT 28.47 3.405 28.64 5.475 ;
        RECT 27.105 4.135 36.75 4.67 ;
        RECT 26.78 3.205 27.11 4.515 ;
        RECT 25.04 3.8 25.295 4.515 ;
        RECT 24.475 4.345 24.85 4.895 ;
        RECT 24.04 3.42 24.37 3.665 ;
        RECT 24.04 3.42 24.225 3.79 ;
        RECT 23.61 3.69 24.215 4.515 ;
        RECT 23.66 3.69 23.925 5.295 ;
        RECT 22.74 3.8 22.955 4.515 ;
        RECT 22.5 4.345 22.78 5.185 ;
        RECT 21.73 3.475 22.06 3.665 ;
        RECT 21.31 3.84 21.925 4.515 ;
        RECT 21.73 3.475 21.925 4.515 ;
        RECT 21.5 3.84 21.83 5.235 ;
        RECT 20.39 3.835 20.65 4.515 ;
        RECT 16.59 4.13 20.165 4.74 ;
        RECT 17.07 4.13 19.82 4.745 ;
        RECT 17.245 4.13 17.415 5.475 ;
        RECT 10.65 4.135 16.59 4.745 ;
        RECT 14.455 4.13 16.435 4.75 ;
        RECT 15.615 3.4 15.785 5.48 ;
        RECT 14.625 3.4 14.795 5.48 ;
        RECT 11.885 3.405 12.055 5.475 ;
        RECT 10.52 4.135 20.165 4.67 ;
        RECT 10.195 3.205 10.525 4.515 ;
        RECT 8.455 3.8 8.71 4.515 ;
        RECT 7.89 4.345 8.265 4.895 ;
        RECT 7.455 3.42 7.785 3.665 ;
        RECT 7.455 3.42 7.64 3.79 ;
        RECT 7.025 3.69 7.63 4.515 ;
        RECT 7.075 3.69 7.34 5.295 ;
        RECT 6.155 3.8 6.37 4.515 ;
        RECT 5.915 4.345 6.195 5.185 ;
        RECT 5.145 3.475 5.475 3.665 ;
        RECT 4.725 3.84 5.34 4.515 ;
        RECT 5.145 3.475 5.34 4.515 ;
        RECT 4.915 3.84 5.245 5.235 ;
        RECT 3.805 3.835 4.065 4.515 ;
        RECT -2.955 4.13 3.58 4.74 ;
        RECT 0.485 4.13 3.235 4.745 ;
        RECT 0.66 4.13 0.83 5.475 ;
        RECT -2.955 4.13 0.005 4.745 ;
        RECT -0.76 4.13 -0.59 8.305 ;
        RECT -2.57 4.13 -2.4 5.475 ;
      LAYER met1 ;
        RECT 76.985 4.15 82.925 4.745 ;
        RECT 77.445 4.135 82.925 4.745 ;
        RECT 80.79 4.13 82.77 4.75 ;
        RECT -2.955 4.19 82.925 4.67 ;
        RECT 76.855 4.15 82.925 4.67 ;
        RECT 66.34 4.13 69.915 4.74 ;
        RECT 66.82 4.13 69.57 4.745 ;
        RECT 60.405 4.15 66.345 4.745 ;
        RECT 60.865 4.135 69.915 4.74 ;
        RECT 64.21 4.13 66.19 4.75 ;
        RECT 60.275 4.15 69.915 4.67 ;
        RECT 49.76 4.13 53.335 4.74 ;
        RECT 50.24 4.13 52.99 4.745 ;
        RECT 43.82 4.15 49.76 4.745 ;
        RECT 44.28 4.135 53.335 4.74 ;
        RECT 47.625 4.13 49.605 4.75 ;
        RECT 43.69 4.15 53.335 4.67 ;
        RECT 33.175 4.13 36.75 4.74 ;
        RECT 33.655 4.13 36.405 4.745 ;
        RECT 27.235 4.15 33.175 4.745 ;
        RECT 27.695 4.135 36.75 4.74 ;
        RECT 31.04 4.13 33.02 4.75 ;
        RECT 27.105 4.15 36.75 4.67 ;
        RECT 16.59 4.13 20.165 4.74 ;
        RECT 17.07 4.13 19.82 4.745 ;
        RECT 10.65 4.15 16.59 4.745 ;
        RECT 11.11 4.135 20.165 4.74 ;
        RECT 14.455 4.13 16.435 4.75 ;
        RECT 10.52 4.15 20.165 4.67 ;
        RECT -2.955 4.13 3.58 4.74 ;
        RECT 0.485 4.13 3.235 4.745 ;
        RECT -2.955 4.13 0.005 4.745 ;
        RECT -0.82 6.655 -0.53 6.885 ;
        RECT -0.99 6.685 -0.53 6.855 ;
      LAYER mcon ;
        RECT -0.76 6.685 -0.59 6.855 ;
        RECT -0.45 4.545 -0.28 4.715 ;
        RECT 2.78 4.545 2.95 4.715 ;
        RECT 3.865 4.345 4.035 4.515 ;
        RECT 4.325 4.345 4.495 4.515 ;
        RECT 4.785 4.345 4.955 4.515 ;
        RECT 5.245 4.345 5.415 4.515 ;
        RECT 5.705 4.345 5.875 4.515 ;
        RECT 6.165 4.345 6.335 4.515 ;
        RECT 6.625 4.345 6.795 4.515 ;
        RECT 7.085 4.345 7.255 4.515 ;
        RECT 7.545 4.345 7.715 4.515 ;
        RECT 8.005 4.345 8.175 4.515 ;
        RECT 8.465 4.345 8.635 4.515 ;
        RECT 8.925 4.345 9.095 4.515 ;
        RECT 9.385 4.345 9.555 4.515 ;
        RECT 9.845 4.345 10.015 4.515 ;
        RECT 10.305 4.345 10.475 4.515 ;
        RECT 14.005 4.545 14.175 4.715 ;
        RECT 14.005 4.165 14.175 4.335 ;
        RECT 14.705 4.55 14.875 4.72 ;
        RECT 14.705 4.16 14.875 4.33 ;
        RECT 15.695 4.55 15.865 4.72 ;
        RECT 15.695 4.16 15.865 4.33 ;
        RECT 19.365 4.545 19.535 4.715 ;
        RECT 20.45 4.345 20.62 4.515 ;
        RECT 20.91 4.345 21.08 4.515 ;
        RECT 21.37 4.345 21.54 4.515 ;
        RECT 21.83 4.345 22 4.515 ;
        RECT 22.29 4.345 22.46 4.515 ;
        RECT 22.75 4.345 22.92 4.515 ;
        RECT 23.21 4.345 23.38 4.515 ;
        RECT 23.67 4.345 23.84 4.515 ;
        RECT 24.13 4.345 24.3 4.515 ;
        RECT 24.59 4.345 24.76 4.515 ;
        RECT 25.05 4.345 25.22 4.515 ;
        RECT 25.51 4.345 25.68 4.515 ;
        RECT 25.97 4.345 26.14 4.515 ;
        RECT 26.43 4.345 26.6 4.515 ;
        RECT 26.89 4.345 27.06 4.515 ;
        RECT 30.59 4.545 30.76 4.715 ;
        RECT 30.59 4.165 30.76 4.335 ;
        RECT 31.29 4.55 31.46 4.72 ;
        RECT 31.29 4.16 31.46 4.33 ;
        RECT 32.28 4.55 32.45 4.72 ;
        RECT 32.28 4.16 32.45 4.33 ;
        RECT 35.95 4.545 36.12 4.715 ;
        RECT 37.035 4.345 37.205 4.515 ;
        RECT 37.495 4.345 37.665 4.515 ;
        RECT 37.955 4.345 38.125 4.515 ;
        RECT 38.415 4.345 38.585 4.515 ;
        RECT 38.875 4.345 39.045 4.515 ;
        RECT 39.335 4.345 39.505 4.515 ;
        RECT 39.795 4.345 39.965 4.515 ;
        RECT 40.255 4.345 40.425 4.515 ;
        RECT 40.715 4.345 40.885 4.515 ;
        RECT 41.175 4.345 41.345 4.515 ;
        RECT 41.635 4.345 41.805 4.515 ;
        RECT 42.095 4.345 42.265 4.515 ;
        RECT 42.555 4.345 42.725 4.515 ;
        RECT 43.015 4.345 43.185 4.515 ;
        RECT 43.475 4.345 43.645 4.515 ;
        RECT 47.175 4.545 47.345 4.715 ;
        RECT 47.175 4.165 47.345 4.335 ;
        RECT 47.875 4.55 48.045 4.72 ;
        RECT 47.875 4.16 48.045 4.33 ;
        RECT 48.865 4.55 49.035 4.72 ;
        RECT 48.865 4.16 49.035 4.33 ;
        RECT 52.535 4.545 52.705 4.715 ;
        RECT 53.62 4.345 53.79 4.515 ;
        RECT 54.08 4.345 54.25 4.515 ;
        RECT 54.54 4.345 54.71 4.515 ;
        RECT 55 4.345 55.17 4.515 ;
        RECT 55.46 4.345 55.63 4.515 ;
        RECT 55.92 4.345 56.09 4.515 ;
        RECT 56.38 4.345 56.55 4.515 ;
        RECT 56.84 4.345 57.01 4.515 ;
        RECT 57.3 4.345 57.47 4.515 ;
        RECT 57.76 4.345 57.93 4.515 ;
        RECT 58.22 4.345 58.39 4.515 ;
        RECT 58.68 4.345 58.85 4.515 ;
        RECT 59.14 4.345 59.31 4.515 ;
        RECT 59.6 4.345 59.77 4.515 ;
        RECT 60.06 4.345 60.23 4.515 ;
        RECT 63.76 4.545 63.93 4.715 ;
        RECT 63.76 4.165 63.93 4.335 ;
        RECT 64.46 4.55 64.63 4.72 ;
        RECT 64.46 4.16 64.63 4.33 ;
        RECT 65.45 4.55 65.62 4.72 ;
        RECT 65.45 4.16 65.62 4.33 ;
        RECT 69.115 4.545 69.285 4.715 ;
        RECT 70.2 4.345 70.37 4.515 ;
        RECT 70.66 4.345 70.83 4.515 ;
        RECT 71.12 4.345 71.29 4.515 ;
        RECT 71.58 4.345 71.75 4.515 ;
        RECT 72.04 4.345 72.21 4.515 ;
        RECT 72.5 4.345 72.67 4.515 ;
        RECT 72.96 4.345 73.13 4.515 ;
        RECT 73.42 4.345 73.59 4.515 ;
        RECT 73.88 4.345 74.05 4.515 ;
        RECT 74.34 4.345 74.51 4.515 ;
        RECT 74.8 4.345 74.97 4.515 ;
        RECT 75.26 4.345 75.43 4.515 ;
        RECT 75.72 4.345 75.89 4.515 ;
        RECT 76.18 4.345 76.35 4.515 ;
        RECT 76.64 4.345 76.81 4.515 ;
        RECT 80.34 4.545 80.51 4.715 ;
        RECT 80.34 4.165 80.51 4.335 ;
        RECT 81.04 4.55 81.21 4.72 ;
        RECT 81.04 4.16 81.21 4.33 ;
        RECT 82.03 4.55 82.2 4.72 ;
        RECT 82.03 4.16 82.2 4.33 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 72.43 6.475 72.76 6.805 ;
        RECT 72.4 6.49 72.7 6.905 ;
        RECT 71.96 6.49 72.76 6.79 ;
        RECT 55.85 6.475 56.18 6.805 ;
        RECT 55.82 6.49 56.12 6.905 ;
        RECT 55.38 6.49 56.18 6.79 ;
        RECT 39.265 6.475 39.595 6.805 ;
        RECT 39.235 6.49 39.535 6.905 ;
        RECT 38.795 6.49 39.595 6.79 ;
        RECT 22.68 6.475 23.01 6.805 ;
        RECT 22.65 6.49 22.95 6.905 ;
        RECT 22.21 6.49 23.01 6.79 ;
        RECT 6.095 6.475 6.425 6.805 ;
        RECT 6.065 6.49 6.365 6.905 ;
        RECT 5.625 6.49 6.425 6.79 ;
      LAYER li1 ;
        RECT 82.745 0 82.925 0.305 ;
        RECT -2.955 0 82.925 0.3 ;
        RECT 81.95 0 82.12 0.93 ;
        RECT 80.96 0 81.13 0.93 ;
        RECT 66.165 0 80.795 0.305 ;
        RECT 78.22 0 78.39 0.935 ;
        RECT 70.055 0 77.145 1.795 ;
        RECT 76.59 0 76.86 2.605 ;
        RECT 75.68 0 75.92 2.605 ;
        RECT 74.81 0 75.06 2.335 ;
        RECT 72.43 0 72.76 2.255 ;
        RECT 70.14 0 70.4 2.615 ;
        RECT 69.8 0 77.145 1.655 ;
        RECT 65.37 0 65.54 0.93 ;
        RECT 64.38 0 64.55 0.93 ;
        RECT 49.58 0 64.215 0.305 ;
        RECT 61.64 0 61.81 0.935 ;
        RECT 53.475 0 60.565 1.795 ;
        RECT 60.01 0 60.28 2.605 ;
        RECT 59.1 0 59.34 2.605 ;
        RECT 58.23 0 58.48 2.335 ;
        RECT 55.85 0 56.18 2.255 ;
        RECT 53.56 0 53.82 2.615 ;
        RECT 53.22 0 60.565 1.655 ;
        RECT 48.785 0 48.955 0.93 ;
        RECT 47.795 0 47.965 0.93 ;
        RECT 32.995 0 47.63 0.305 ;
        RECT 45.055 0 45.225 0.935 ;
        RECT 36.89 0 43.98 1.795 ;
        RECT 43.425 0 43.695 2.605 ;
        RECT 42.515 0 42.755 2.605 ;
        RECT 41.645 0 41.895 2.335 ;
        RECT 39.265 0 39.595 2.255 ;
        RECT 36.975 0 37.235 2.615 ;
        RECT 36.635 0 43.98 1.655 ;
        RECT 32.2 0 32.37 0.93 ;
        RECT 31.21 0 31.38 0.93 ;
        RECT 16.41 0 31.045 0.305 ;
        RECT 28.47 0 28.64 0.935 ;
        RECT 20.305 0 27.395 1.795 ;
        RECT 26.84 0 27.11 2.605 ;
        RECT 25.93 0 26.17 2.605 ;
        RECT 25.06 0 25.31 2.335 ;
        RECT 22.68 0 23.01 2.255 ;
        RECT 20.39 0 20.65 2.615 ;
        RECT 20.05 0 27.395 1.655 ;
        RECT 15.615 0 15.785 0.93 ;
        RECT 14.625 0 14.795 0.93 ;
        RECT -2.955 0 14.46 0.305 ;
        RECT 11.885 0 12.055 0.935 ;
        RECT 3.72 0 10.81 1.795 ;
        RECT 10.255 0 10.525 2.605 ;
        RECT 9.345 0 9.585 2.605 ;
        RECT 8.475 0 8.725 2.335 ;
        RECT 6.095 0 6.425 2.255 ;
        RECT 3.805 0 4.065 2.615 ;
        RECT 3.465 0 10.81 1.655 ;
        RECT -2.955 8.58 82.925 8.88 ;
        RECT 82.745 8.575 82.925 8.88 ;
        RECT 81.95 7.95 82.12 8.88 ;
        RECT 80.96 7.95 81.13 8.88 ;
        RECT 66.165 8.575 80.795 8.88 ;
        RECT 78.22 7.945 78.39 8.88 ;
        RECT 69.76 7.18 76.96 8.88 ;
        RECT 70.055 7.065 76.955 8.88 ;
        RECT 75.49 6.555 75.94 8.88 ;
        RECT 73.4 6.665 73.73 8.88 ;
        RECT 71.33 6.605 71.58 8.88 ;
        RECT 66.995 7.945 67.165 8.88 ;
        RECT 65.37 7.95 65.54 8.88 ;
        RECT 64.38 7.95 64.55 8.88 ;
        RECT 49.58 8.575 64.215 8.88 ;
        RECT 61.64 7.945 61.81 8.88 ;
        RECT 53.18 7.18 60.38 8.88 ;
        RECT 53.475 7.065 60.375 8.88 ;
        RECT 58.91 6.555 59.36 8.88 ;
        RECT 56.82 6.665 57.15 8.88 ;
        RECT 54.75 6.605 55 8.88 ;
        RECT 50.415 7.945 50.585 8.88 ;
        RECT 48.785 7.95 48.955 8.88 ;
        RECT 47.795 7.95 47.965 8.88 ;
        RECT 32.995 8.575 47.63 8.88 ;
        RECT 45.055 7.945 45.225 8.88 ;
        RECT 36.595 7.18 43.795 8.88 ;
        RECT 36.89 7.065 43.79 8.88 ;
        RECT 42.325 6.555 42.775 8.88 ;
        RECT 40.235 6.665 40.565 8.88 ;
        RECT 38.165 6.605 38.415 8.88 ;
        RECT 33.83 7.945 34 8.88 ;
        RECT 32.2 7.95 32.37 8.88 ;
        RECT 31.21 7.95 31.38 8.88 ;
        RECT 16.41 8.575 31.045 8.88 ;
        RECT 28.47 7.945 28.64 8.88 ;
        RECT 20.01 7.18 27.21 8.88 ;
        RECT 20.305 7.065 27.205 8.88 ;
        RECT 25.74 6.555 26.19 8.88 ;
        RECT 23.65 6.665 23.98 8.88 ;
        RECT 21.58 6.605 21.83 8.88 ;
        RECT 17.245 7.945 17.415 8.88 ;
        RECT 15.615 7.95 15.785 8.88 ;
        RECT 14.625 7.95 14.795 8.88 ;
        RECT -2.955 8.575 14.46 8.88 ;
        RECT 11.885 7.945 12.055 8.88 ;
        RECT 3.425 7.18 10.625 8.88 ;
        RECT 3.72 7.065 10.62 8.88 ;
        RECT 9.155 6.555 9.605 8.88 ;
        RECT 7.065 6.665 7.395 8.88 ;
        RECT 4.995 6.605 5.245 8.88 ;
        RECT 0.66 7.945 0.83 8.88 ;
        RECT -2.57 7.945 -2.4 8.88 ;
        RECT 73.7 5.825 74.025 6.155 ;
        RECT 71.48 5.825 71.82 6.075 ;
        RECT 68 6.075 68.17 8.025 ;
        RECT 67.945 7.855 68.115 8.305 ;
        RECT 67.945 5.015 68.115 6.245 ;
        RECT 57.12 5.825 57.445 6.155 ;
        RECT 54.9 5.825 55.24 6.075 ;
        RECT 51.42 6.075 51.59 8.025 ;
        RECT 51.365 7.855 51.535 8.305 ;
        RECT 51.365 5.015 51.535 6.245 ;
        RECT 40.535 5.825 40.86 6.155 ;
        RECT 38.315 5.825 38.655 6.075 ;
        RECT 34.835 6.075 35.005 8.025 ;
        RECT 34.78 7.855 34.95 8.305 ;
        RECT 34.78 5.015 34.95 6.245 ;
        RECT 23.95 5.825 24.275 6.155 ;
        RECT 21.73 5.825 22.07 6.075 ;
        RECT 18.25 6.075 18.42 8.025 ;
        RECT 18.195 7.855 18.365 8.305 ;
        RECT 18.195 5.015 18.365 6.245 ;
        RECT 7.365 5.825 7.69 6.155 ;
        RECT 5.145 5.825 5.485 6.075 ;
        RECT 1.665 6.075 1.835 8.025 ;
        RECT 1.61 7.855 1.78 8.305 ;
        RECT 1.61 5.015 1.78 6.245 ;
      LAYER met2 ;
        RECT 72.455 6.455 72.735 6.825 ;
        RECT 55.875 6.455 56.155 6.825 ;
        RECT 39.29 6.455 39.57 6.825 ;
        RECT 22.705 6.455 22.985 6.825 ;
        RECT 6.12 6.455 6.4 6.825 ;
      LAYER met1 ;
        RECT 82.745 0 82.925 0.305 ;
        RECT -2.955 0 82.925 0.3 ;
        RECT 66.165 0 80.795 0.305 ;
        RECT 70.055 0 77.145 1.795 ;
        RECT 70.055 0 76.955 1.95 ;
        RECT 69.8 0 77.145 1.655 ;
        RECT 49.58 0 64.215 0.305 ;
        RECT 53.475 0 60.565 1.795 ;
        RECT 53.475 0 60.375 1.95 ;
        RECT 53.22 0 60.565 1.655 ;
        RECT 32.995 0 47.63 0.305 ;
        RECT 36.89 0 43.98 1.795 ;
        RECT 36.89 0 43.79 1.95 ;
        RECT 36.635 0 43.98 1.655 ;
        RECT 16.41 0 31.045 0.305 ;
        RECT 20.305 0 27.395 1.795 ;
        RECT 20.305 0 27.205 1.95 ;
        RECT 20.05 0 27.395 1.655 ;
        RECT -2.955 0 14.46 0.305 ;
        RECT 3.72 0 10.81 1.795 ;
        RECT 3.72 0 10.62 1.95 ;
        RECT 3.465 0 10.81 1.655 ;
        RECT -2.955 8.58 82.925 8.88 ;
        RECT 82.745 8.575 82.925 8.88 ;
        RECT 66.165 8.575 80.795 8.88 ;
        RECT 69.76 7.18 76.96 8.88 ;
        RECT 70.055 6.91 76.955 8.88 ;
        RECT 73.65 5.845 73.94 6.075 ;
        RECT 71.515 6.57 73.865 6.71 ;
        RECT 73.725 5.845 73.865 6.71 ;
        RECT 72.445 6.51 72.765 6.77 ;
        RECT 72.48 6.51 72.735 8.88 ;
        RECT 71.44 5.845 71.73 6.075 ;
        RECT 71.515 5.845 71.655 6.71 ;
        RECT 67.94 6.285 68.23 6.515 ;
        RECT 67.78 6.315 67.95 8.88 ;
        RECT 67.77 6.315 68.23 6.485 ;
        RECT 49.58 8.575 64.215 8.88 ;
        RECT 53.18 7.18 60.38 8.88 ;
        RECT 53.475 6.91 60.375 8.88 ;
        RECT 57.07 5.845 57.36 6.075 ;
        RECT 54.935 6.57 57.285 6.71 ;
        RECT 57.145 5.845 57.285 6.71 ;
        RECT 55.865 6.51 56.185 6.77 ;
        RECT 55.9 6.51 56.155 8.88 ;
        RECT 54.86 5.845 55.15 6.075 ;
        RECT 54.935 5.845 55.075 6.71 ;
        RECT 51.36 6.285 51.65 6.515 ;
        RECT 51.2 6.315 51.37 8.88 ;
        RECT 51.19 6.315 51.65 6.485 ;
        RECT 32.995 8.575 47.63 8.88 ;
        RECT 36.595 7.18 43.795 8.88 ;
        RECT 36.89 6.91 43.79 8.88 ;
        RECT 40.485 5.845 40.775 6.075 ;
        RECT 38.35 6.57 40.7 6.71 ;
        RECT 40.56 5.845 40.7 6.71 ;
        RECT 39.28 6.51 39.6 6.77 ;
        RECT 39.315 6.51 39.57 8.88 ;
        RECT 38.275 5.845 38.565 6.075 ;
        RECT 38.35 5.845 38.49 6.71 ;
        RECT 34.775 6.285 35.065 6.515 ;
        RECT 34.615 6.315 34.785 8.88 ;
        RECT 34.605 6.315 35.065 6.485 ;
        RECT 16.41 8.575 31.045 8.88 ;
        RECT 20.01 7.18 27.21 8.88 ;
        RECT 20.305 6.91 27.205 8.88 ;
        RECT 23.9 5.845 24.19 6.075 ;
        RECT 21.765 6.57 24.115 6.71 ;
        RECT 23.975 5.845 24.115 6.71 ;
        RECT 22.695 6.51 23.015 6.77 ;
        RECT 22.73 6.51 22.985 8.88 ;
        RECT 21.69 5.845 21.98 6.075 ;
        RECT 21.765 5.845 21.905 6.71 ;
        RECT 18.19 6.285 18.48 6.515 ;
        RECT 18.03 6.315 18.2 8.88 ;
        RECT 18.02 6.315 18.48 6.485 ;
        RECT -2.955 8.575 14.46 8.88 ;
        RECT 3.425 7.18 10.625 8.88 ;
        RECT 3.72 6.91 10.62 8.88 ;
        RECT 7.315 5.845 7.605 6.075 ;
        RECT 5.18 6.57 7.53 6.71 ;
        RECT 7.39 5.845 7.53 6.71 ;
        RECT 6.11 6.51 6.43 6.77 ;
        RECT 6.145 6.51 6.4 8.88 ;
        RECT 5.105 5.845 5.395 6.075 ;
        RECT 5.18 5.845 5.32 6.71 ;
        RECT 1.605 6.285 1.895 6.515 ;
        RECT 1.445 6.315 1.615 8.88 ;
        RECT 1.435 6.315 1.895 6.485 ;
      LAYER via2 ;
        RECT 6.16 6.54 6.36 6.74 ;
        RECT 22.745 6.54 22.945 6.74 ;
        RECT 39.33 6.54 39.53 6.74 ;
        RECT 55.915 6.54 56.115 6.74 ;
        RECT 72.495 6.54 72.695 6.74 ;
      LAYER via1 ;
        RECT 6.195 6.565 6.345 6.715 ;
        RECT 22.78 6.565 22.93 6.715 ;
        RECT 39.365 6.565 39.515 6.715 ;
        RECT 55.95 6.565 56.1 6.715 ;
        RECT 72.53 6.565 72.68 6.715 ;
      LAYER mcon ;
        RECT -2.49 8.605 -2.32 8.775 ;
        RECT -1.81 8.605 -1.64 8.775 ;
        RECT -1.13 8.605 -0.96 8.775 ;
        RECT -0.45 8.605 -0.28 8.775 ;
        RECT 0.74 8.605 0.91 8.775 ;
        RECT 1.42 8.605 1.59 8.775 ;
        RECT 1.665 6.315 1.835 6.485 ;
        RECT 2.1 8.605 2.27 8.775 ;
        RECT 2.78 8.605 2.95 8.775 ;
        RECT 3.865 7.065 4.035 7.235 ;
        RECT 3.865 1.625 4.035 1.795 ;
        RECT 4.325 7.065 4.495 7.235 ;
        RECT 4.325 1.625 4.495 1.795 ;
        RECT 4.785 7.065 4.955 7.235 ;
        RECT 4.785 1.625 4.955 1.795 ;
        RECT 5.165 5.875 5.335 6.045 ;
        RECT 5.245 7.065 5.415 7.235 ;
        RECT 5.245 1.625 5.415 1.795 ;
        RECT 5.705 7.065 5.875 7.235 ;
        RECT 5.705 1.625 5.875 1.795 ;
        RECT 6.165 7.065 6.335 7.235 ;
        RECT 6.165 1.625 6.335 1.795 ;
        RECT 6.625 7.065 6.795 7.235 ;
        RECT 6.625 1.625 6.795 1.795 ;
        RECT 7.085 7.065 7.255 7.235 ;
        RECT 7.085 1.625 7.255 1.795 ;
        RECT 7.375 5.875 7.545 6.045 ;
        RECT 7.545 7.065 7.715 7.235 ;
        RECT 7.545 1.625 7.715 1.795 ;
        RECT 8.005 7.065 8.175 7.235 ;
        RECT 8.005 1.625 8.175 1.795 ;
        RECT 8.465 7.065 8.635 7.235 ;
        RECT 8.465 1.625 8.635 1.795 ;
        RECT 8.925 7.065 9.095 7.235 ;
        RECT 8.925 1.625 9.095 1.795 ;
        RECT 9.385 7.065 9.555 7.235 ;
        RECT 9.385 1.625 9.555 1.795 ;
        RECT 9.845 7.065 10.015 7.235 ;
        RECT 9.845 1.625 10.015 1.795 ;
        RECT 10.305 7.065 10.475 7.235 ;
        RECT 10.305 1.625 10.475 1.795 ;
        RECT 11.965 8.605 12.135 8.775 ;
        RECT 11.965 0.105 12.135 0.275 ;
        RECT 12.645 8.605 12.815 8.775 ;
        RECT 12.645 0.105 12.815 0.275 ;
        RECT 13.325 8.605 13.495 8.775 ;
        RECT 13.325 0.105 13.495 0.275 ;
        RECT 14.005 8.605 14.175 8.775 ;
        RECT 14.005 0.105 14.175 0.275 ;
        RECT 14.705 8.61 14.875 8.78 ;
        RECT 14.705 0.1 14.875 0.27 ;
        RECT 15.695 8.61 15.865 8.78 ;
        RECT 15.695 0.1 15.865 0.27 ;
        RECT 17.325 8.605 17.495 8.775 ;
        RECT 18.005 8.605 18.175 8.775 ;
        RECT 18.25 6.315 18.42 6.485 ;
        RECT 18.685 8.605 18.855 8.775 ;
        RECT 19.365 8.605 19.535 8.775 ;
        RECT 20.45 7.065 20.62 7.235 ;
        RECT 20.45 1.625 20.62 1.795 ;
        RECT 20.91 7.065 21.08 7.235 ;
        RECT 20.91 1.625 21.08 1.795 ;
        RECT 21.37 7.065 21.54 7.235 ;
        RECT 21.37 1.625 21.54 1.795 ;
        RECT 21.75 5.875 21.92 6.045 ;
        RECT 21.83 7.065 22 7.235 ;
        RECT 21.83 1.625 22 1.795 ;
        RECT 22.29 7.065 22.46 7.235 ;
        RECT 22.29 1.625 22.46 1.795 ;
        RECT 22.75 7.065 22.92 7.235 ;
        RECT 22.75 1.625 22.92 1.795 ;
        RECT 23.21 7.065 23.38 7.235 ;
        RECT 23.21 1.625 23.38 1.795 ;
        RECT 23.67 7.065 23.84 7.235 ;
        RECT 23.67 1.625 23.84 1.795 ;
        RECT 23.96 5.875 24.13 6.045 ;
        RECT 24.13 7.065 24.3 7.235 ;
        RECT 24.13 1.625 24.3 1.795 ;
        RECT 24.59 7.065 24.76 7.235 ;
        RECT 24.59 1.625 24.76 1.795 ;
        RECT 25.05 7.065 25.22 7.235 ;
        RECT 25.05 1.625 25.22 1.795 ;
        RECT 25.51 7.065 25.68 7.235 ;
        RECT 25.51 1.625 25.68 1.795 ;
        RECT 25.97 7.065 26.14 7.235 ;
        RECT 25.97 1.625 26.14 1.795 ;
        RECT 26.43 7.065 26.6 7.235 ;
        RECT 26.43 1.625 26.6 1.795 ;
        RECT 26.89 7.065 27.06 7.235 ;
        RECT 26.89 1.625 27.06 1.795 ;
        RECT 28.55 8.605 28.72 8.775 ;
        RECT 28.55 0.105 28.72 0.275 ;
        RECT 29.23 8.605 29.4 8.775 ;
        RECT 29.23 0.105 29.4 0.275 ;
        RECT 29.91 8.605 30.08 8.775 ;
        RECT 29.91 0.105 30.08 0.275 ;
        RECT 30.59 8.605 30.76 8.775 ;
        RECT 30.59 0.105 30.76 0.275 ;
        RECT 31.29 8.61 31.46 8.78 ;
        RECT 31.29 0.1 31.46 0.27 ;
        RECT 32.28 8.61 32.45 8.78 ;
        RECT 32.28 0.1 32.45 0.27 ;
        RECT 33.91 8.605 34.08 8.775 ;
        RECT 34.59 8.605 34.76 8.775 ;
        RECT 34.835 6.315 35.005 6.485 ;
        RECT 35.27 8.605 35.44 8.775 ;
        RECT 35.95 8.605 36.12 8.775 ;
        RECT 37.035 7.065 37.205 7.235 ;
        RECT 37.035 1.625 37.205 1.795 ;
        RECT 37.495 7.065 37.665 7.235 ;
        RECT 37.495 1.625 37.665 1.795 ;
        RECT 37.955 7.065 38.125 7.235 ;
        RECT 37.955 1.625 38.125 1.795 ;
        RECT 38.335 5.875 38.505 6.045 ;
        RECT 38.415 7.065 38.585 7.235 ;
        RECT 38.415 1.625 38.585 1.795 ;
        RECT 38.875 7.065 39.045 7.235 ;
        RECT 38.875 1.625 39.045 1.795 ;
        RECT 39.335 7.065 39.505 7.235 ;
        RECT 39.335 1.625 39.505 1.795 ;
        RECT 39.795 7.065 39.965 7.235 ;
        RECT 39.795 1.625 39.965 1.795 ;
        RECT 40.255 7.065 40.425 7.235 ;
        RECT 40.255 1.625 40.425 1.795 ;
        RECT 40.545 5.875 40.715 6.045 ;
        RECT 40.715 7.065 40.885 7.235 ;
        RECT 40.715 1.625 40.885 1.795 ;
        RECT 41.175 7.065 41.345 7.235 ;
        RECT 41.175 1.625 41.345 1.795 ;
        RECT 41.635 7.065 41.805 7.235 ;
        RECT 41.635 1.625 41.805 1.795 ;
        RECT 42.095 7.065 42.265 7.235 ;
        RECT 42.095 1.625 42.265 1.795 ;
        RECT 42.555 7.065 42.725 7.235 ;
        RECT 42.555 1.625 42.725 1.795 ;
        RECT 43.015 7.065 43.185 7.235 ;
        RECT 43.015 1.625 43.185 1.795 ;
        RECT 43.475 7.065 43.645 7.235 ;
        RECT 43.475 1.625 43.645 1.795 ;
        RECT 45.135 8.605 45.305 8.775 ;
        RECT 45.135 0.105 45.305 0.275 ;
        RECT 45.815 8.605 45.985 8.775 ;
        RECT 45.815 0.105 45.985 0.275 ;
        RECT 46.495 8.605 46.665 8.775 ;
        RECT 46.495 0.105 46.665 0.275 ;
        RECT 47.175 8.605 47.345 8.775 ;
        RECT 47.175 0.105 47.345 0.275 ;
        RECT 47.875 8.61 48.045 8.78 ;
        RECT 47.875 0.1 48.045 0.27 ;
        RECT 48.865 8.61 49.035 8.78 ;
        RECT 48.865 0.1 49.035 0.27 ;
        RECT 50.495 8.605 50.665 8.775 ;
        RECT 51.175 8.605 51.345 8.775 ;
        RECT 51.42 6.315 51.59 6.485 ;
        RECT 51.855 8.605 52.025 8.775 ;
        RECT 52.535 8.605 52.705 8.775 ;
        RECT 53.62 7.065 53.79 7.235 ;
        RECT 53.62 1.625 53.79 1.795 ;
        RECT 54.08 7.065 54.25 7.235 ;
        RECT 54.08 1.625 54.25 1.795 ;
        RECT 54.54 7.065 54.71 7.235 ;
        RECT 54.54 1.625 54.71 1.795 ;
        RECT 54.92 5.875 55.09 6.045 ;
        RECT 55 7.065 55.17 7.235 ;
        RECT 55 1.625 55.17 1.795 ;
        RECT 55.46 7.065 55.63 7.235 ;
        RECT 55.46 1.625 55.63 1.795 ;
        RECT 55.92 7.065 56.09 7.235 ;
        RECT 55.92 1.625 56.09 1.795 ;
        RECT 56.38 7.065 56.55 7.235 ;
        RECT 56.38 1.625 56.55 1.795 ;
        RECT 56.84 7.065 57.01 7.235 ;
        RECT 56.84 1.625 57.01 1.795 ;
        RECT 57.13 5.875 57.3 6.045 ;
        RECT 57.3 7.065 57.47 7.235 ;
        RECT 57.3 1.625 57.47 1.795 ;
        RECT 57.76 7.065 57.93 7.235 ;
        RECT 57.76 1.625 57.93 1.795 ;
        RECT 58.22 7.065 58.39 7.235 ;
        RECT 58.22 1.625 58.39 1.795 ;
        RECT 58.68 7.065 58.85 7.235 ;
        RECT 58.68 1.625 58.85 1.795 ;
        RECT 59.14 7.065 59.31 7.235 ;
        RECT 59.14 1.625 59.31 1.795 ;
        RECT 59.6 7.065 59.77 7.235 ;
        RECT 59.6 1.625 59.77 1.795 ;
        RECT 60.06 7.065 60.23 7.235 ;
        RECT 60.06 1.625 60.23 1.795 ;
        RECT 61.72 8.605 61.89 8.775 ;
        RECT 61.72 0.105 61.89 0.275 ;
        RECT 62.4 8.605 62.57 8.775 ;
        RECT 62.4 0.105 62.57 0.275 ;
        RECT 63.08 8.605 63.25 8.775 ;
        RECT 63.08 0.105 63.25 0.275 ;
        RECT 63.76 8.605 63.93 8.775 ;
        RECT 63.76 0.105 63.93 0.275 ;
        RECT 64.46 8.61 64.63 8.78 ;
        RECT 64.46 0.1 64.63 0.27 ;
        RECT 65.45 8.61 65.62 8.78 ;
        RECT 65.45 0.1 65.62 0.27 ;
        RECT 67.075 8.605 67.245 8.775 ;
        RECT 67.755 8.605 67.925 8.775 ;
        RECT 68 6.315 68.17 6.485 ;
        RECT 68.435 8.605 68.605 8.775 ;
        RECT 69.115 8.605 69.285 8.775 ;
        RECT 70.2 7.065 70.37 7.235 ;
        RECT 70.2 1.625 70.37 1.795 ;
        RECT 70.66 7.065 70.83 7.235 ;
        RECT 70.66 1.625 70.83 1.795 ;
        RECT 71.12 7.065 71.29 7.235 ;
        RECT 71.12 1.625 71.29 1.795 ;
        RECT 71.5 5.875 71.67 6.045 ;
        RECT 71.58 7.065 71.75 7.235 ;
        RECT 71.58 1.625 71.75 1.795 ;
        RECT 72.04 7.065 72.21 7.235 ;
        RECT 72.04 1.625 72.21 1.795 ;
        RECT 72.5 7.065 72.67 7.235 ;
        RECT 72.5 1.625 72.67 1.795 ;
        RECT 72.96 7.065 73.13 7.235 ;
        RECT 72.96 1.625 73.13 1.795 ;
        RECT 73.42 7.065 73.59 7.235 ;
        RECT 73.42 1.625 73.59 1.795 ;
        RECT 73.71 5.875 73.88 6.045 ;
        RECT 73.88 7.065 74.05 7.235 ;
        RECT 73.88 1.625 74.05 1.795 ;
        RECT 74.34 7.065 74.51 7.235 ;
        RECT 74.34 1.625 74.51 1.795 ;
        RECT 74.8 7.065 74.97 7.235 ;
        RECT 74.8 1.625 74.97 1.795 ;
        RECT 75.26 7.065 75.43 7.235 ;
        RECT 75.26 1.625 75.43 1.795 ;
        RECT 75.72 7.065 75.89 7.235 ;
        RECT 75.72 1.625 75.89 1.795 ;
        RECT 76.18 7.065 76.35 7.235 ;
        RECT 76.18 1.625 76.35 1.795 ;
        RECT 76.64 7.065 76.81 7.235 ;
        RECT 76.64 1.625 76.81 1.795 ;
        RECT 78.3 8.605 78.47 8.775 ;
        RECT 78.3 0.105 78.47 0.275 ;
        RECT 78.98 8.605 79.15 8.775 ;
        RECT 78.98 0.105 79.15 0.275 ;
        RECT 79.66 8.605 79.83 8.775 ;
        RECT 79.66 0.105 79.83 0.275 ;
        RECT 80.34 8.605 80.51 8.775 ;
        RECT 80.34 0.105 80.51 0.275 ;
        RECT 81.04 8.61 81.21 8.78 ;
        RECT 81.04 0.1 81.21 0.27 ;
        RECT 82.03 8.61 82.2 8.78 ;
        RECT 82.03 0.1 82.2 0.27 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 74.83 2.735 75.16 3.065 ;
      RECT 74.83 2.75 75.63 3.05 ;
      RECT 74.83 2.73 75.15 3.065 ;
      RECT 69.15 7.97 73.43 8.27 ;
      RECT 73.125 5.795 73.425 8.27 ;
      RECT 69.15 7.03 69.45 8.27 ;
      RECT 68.275 6.995 68.645 7.365 ;
      RECT 68.275 7.03 69.45 7.33 ;
      RECT 74.15 5.795 74.48 6.125 ;
      RECT 72.5 5.795 73.435 6.125 ;
      RECT 72.5 5.81 74.95 6.11 ;
      RECT 72.5 5.795 74.48 6.11 ;
      RECT 74.155 5.79 74.455 6.125 ;
      RECT 72.5 3.765 72.83 6.125 ;
      RECT 72.5 3.765 74.795 4.095 ;
      RECT 72.5 3.765 75.16 4.085 ;
      RECT 74.83 3.755 75.16 4.085 ;
      RECT 72.5 3.77 75.63 4.07 ;
      RECT 74.835 3.705 75.135 4.085 ;
      RECT 74.13 3.075 74.46 3.405 ;
      RECT 73.66 3.09 74.46 3.39 ;
      RECT 74.155 3.06 74.455 3.405 ;
      RECT 73.47 4.775 73.8 5.105 ;
      RECT 73.47 4.79 74.27 5.09 ;
      RECT 72.79 2.39 73.12 2.72 ;
      RECT 72.32 2.41 72.68 2.71 ;
      RECT 72.68 2.405 73.12 2.705 ;
      RECT 58.25 2.735 58.58 3.065 ;
      RECT 58.25 2.75 59.05 3.05 ;
      RECT 58.25 2.73 58.57 3.065 ;
      RECT 52.57 7.97 56.85 8.27 ;
      RECT 56.545 5.795 56.845 8.27 ;
      RECT 52.57 7.03 52.87 8.27 ;
      RECT 51.695 6.995 52.065 7.365 ;
      RECT 51.695 7.03 52.87 7.33 ;
      RECT 57.57 5.795 57.9 6.125 ;
      RECT 55.92 5.795 56.855 6.125 ;
      RECT 55.92 5.81 58.37 6.11 ;
      RECT 55.92 5.795 57.9 6.11 ;
      RECT 57.575 5.79 57.875 6.125 ;
      RECT 55.92 3.765 56.25 6.125 ;
      RECT 55.92 3.765 58.215 4.095 ;
      RECT 55.92 3.765 58.58 4.085 ;
      RECT 58.25 3.755 58.58 4.085 ;
      RECT 55.92 3.77 59.05 4.07 ;
      RECT 58.255 3.705 58.555 4.085 ;
      RECT 57.55 3.075 57.88 3.405 ;
      RECT 57.08 3.09 57.88 3.39 ;
      RECT 57.575 3.06 57.875 3.405 ;
      RECT 56.89 4.775 57.22 5.105 ;
      RECT 56.89 4.79 57.69 5.09 ;
      RECT 56.21 2.39 56.54 2.72 ;
      RECT 55.74 2.41 56.1 2.71 ;
      RECT 56.1 2.405 56.54 2.705 ;
      RECT 41.665 2.735 41.995 3.065 ;
      RECT 41.665 2.75 42.465 3.05 ;
      RECT 41.665 2.73 41.985 3.065 ;
      RECT 35.985 7.97 40.265 8.27 ;
      RECT 39.96 5.795 40.26 8.27 ;
      RECT 35.985 7.03 36.285 8.27 ;
      RECT 35.11 6.995 35.48 7.365 ;
      RECT 35.11 7.03 36.285 7.33 ;
      RECT 40.985 5.795 41.315 6.125 ;
      RECT 39.335 5.795 40.27 6.125 ;
      RECT 39.335 5.81 41.785 6.11 ;
      RECT 39.335 5.795 41.315 6.11 ;
      RECT 40.99 5.79 41.29 6.125 ;
      RECT 39.335 3.765 39.665 6.125 ;
      RECT 39.335 3.765 41.63 4.095 ;
      RECT 39.335 3.765 41.995 4.085 ;
      RECT 41.665 3.755 41.995 4.085 ;
      RECT 39.335 3.77 42.465 4.07 ;
      RECT 41.67 3.705 41.97 4.085 ;
      RECT 40.965 3.075 41.295 3.405 ;
      RECT 40.495 3.09 41.295 3.39 ;
      RECT 40.99 3.06 41.29 3.405 ;
      RECT 40.305 4.775 40.635 5.105 ;
      RECT 40.305 4.79 41.105 5.09 ;
      RECT 39.625 2.39 39.955 2.72 ;
      RECT 39.155 2.41 39.515 2.71 ;
      RECT 39.515 2.405 39.955 2.705 ;
      RECT 25.08 2.735 25.41 3.065 ;
      RECT 25.08 2.75 25.88 3.05 ;
      RECT 25.08 2.73 25.4 3.065 ;
      RECT 19.4 7.97 23.68 8.27 ;
      RECT 23.375 5.795 23.675 8.27 ;
      RECT 19.4 7.03 19.7 8.27 ;
      RECT 18.525 6.995 18.895 7.365 ;
      RECT 18.525 7.03 19.7 7.33 ;
      RECT 24.4 5.795 24.73 6.125 ;
      RECT 22.75 5.795 23.685 6.125 ;
      RECT 22.75 5.81 25.2 6.11 ;
      RECT 22.75 5.795 24.73 6.11 ;
      RECT 24.405 5.79 24.705 6.125 ;
      RECT 22.75 3.765 23.08 6.125 ;
      RECT 22.75 3.765 25.045 4.095 ;
      RECT 22.75 3.765 25.41 4.085 ;
      RECT 25.08 3.755 25.41 4.085 ;
      RECT 22.75 3.77 25.88 4.07 ;
      RECT 25.085 3.705 25.385 4.085 ;
      RECT 24.38 3.075 24.71 3.405 ;
      RECT 23.91 3.09 24.71 3.39 ;
      RECT 24.405 3.06 24.705 3.405 ;
      RECT 23.72 4.775 24.05 5.105 ;
      RECT 23.72 4.79 24.52 5.09 ;
      RECT 23.04 2.39 23.37 2.72 ;
      RECT 22.57 2.41 22.93 2.71 ;
      RECT 22.93 2.405 23.37 2.705 ;
      RECT 8.495 2.735 8.825 3.065 ;
      RECT 8.495 2.75 9.295 3.05 ;
      RECT 8.495 2.73 8.815 3.065 ;
      RECT 2.815 7.97 7.095 8.27 ;
      RECT 6.79 5.795 7.09 8.27 ;
      RECT 2.815 7.03 3.115 8.27 ;
      RECT 1.94 6.995 2.31 7.365 ;
      RECT 1.94 7.03 3.115 7.33 ;
      RECT 7.815 5.795 8.145 6.125 ;
      RECT 6.165 5.795 7.1 6.125 ;
      RECT 6.165 5.81 8.615 6.11 ;
      RECT 6.165 5.795 8.145 6.11 ;
      RECT 7.82 5.79 8.12 6.125 ;
      RECT 6.165 3.765 6.495 6.125 ;
      RECT 6.165 3.765 8.46 4.095 ;
      RECT 6.165 3.765 8.825 4.085 ;
      RECT 8.495 3.755 8.825 4.085 ;
      RECT 6.165 3.77 9.295 4.07 ;
      RECT 8.5 3.705 8.8 4.085 ;
      RECT 7.795 3.075 8.125 3.405 ;
      RECT 7.325 3.09 8.125 3.39 ;
      RECT 7.82 3.06 8.12 3.405 ;
      RECT 7.135 4.775 7.465 5.105 ;
      RECT 7.135 4.79 7.935 5.09 ;
      RECT 6.455 2.39 6.785 2.72 ;
      RECT 5.985 2.41 6.345 2.71 ;
      RECT 6.345 2.405 6.785 2.705 ;
    LAYER via2 ;
      RECT 74.895 2.8 75.095 3 ;
      RECT 74.895 3.82 75.095 4.02 ;
      RECT 74.215 5.86 74.415 6.06 ;
      RECT 74.195 3.14 74.395 3.34 ;
      RECT 73.535 4.84 73.735 5.04 ;
      RECT 73.17 5.86 73.37 6.06 ;
      RECT 72.855 2.455 73.055 2.655 ;
      RECT 68.36 7.08 68.56 7.28 ;
      RECT 58.315 2.8 58.515 3 ;
      RECT 58.315 3.82 58.515 4.02 ;
      RECT 57.635 5.86 57.835 6.06 ;
      RECT 57.615 3.14 57.815 3.34 ;
      RECT 56.955 4.84 57.155 5.04 ;
      RECT 56.59 5.86 56.79 6.06 ;
      RECT 56.275 2.455 56.475 2.655 ;
      RECT 51.78 7.08 51.98 7.28 ;
      RECT 41.73 2.8 41.93 3 ;
      RECT 41.73 3.82 41.93 4.02 ;
      RECT 41.05 5.86 41.25 6.06 ;
      RECT 41.03 3.14 41.23 3.34 ;
      RECT 40.37 4.84 40.57 5.04 ;
      RECT 40.005 5.86 40.205 6.06 ;
      RECT 39.69 2.455 39.89 2.655 ;
      RECT 35.195 7.08 35.395 7.28 ;
      RECT 25.145 2.8 25.345 3 ;
      RECT 25.145 3.82 25.345 4.02 ;
      RECT 24.465 5.86 24.665 6.06 ;
      RECT 24.445 3.14 24.645 3.34 ;
      RECT 23.785 4.84 23.985 5.04 ;
      RECT 23.42 5.86 23.62 6.06 ;
      RECT 23.105 2.455 23.305 2.655 ;
      RECT 18.61 7.08 18.81 7.28 ;
      RECT 8.56 2.8 8.76 3 ;
      RECT 8.56 3.82 8.76 4.02 ;
      RECT 7.88 5.86 8.08 6.06 ;
      RECT 7.86 3.14 8.06 3.34 ;
      RECT 7.2 4.84 7.4 5.04 ;
      RECT 6.835 5.86 7.035 6.06 ;
      RECT 6.52 2.455 6.72 2.655 ;
      RECT 2.025 7.08 2.225 7.28 ;
    LAYER met2 ;
      RECT -1.585 8.6 82.555 8.77 ;
      RECT 82.385 7.3 82.555 8.77 ;
      RECT -1.585 6.255 -1.415 8.77 ;
      RECT 82.35 7.3 82.675 7.625 ;
      RECT -1.625 6.255 -1.345 6.595 ;
      RECT 79.195 6.28 79.515 6.605 ;
      RECT 79.225 5.695 79.395 6.605 ;
      RECT 79.225 5.695 79.4 6.045 ;
      RECT 79.225 5.695 80.2 5.87 ;
      RECT 80.025 1.965 80.2 5.87 ;
      RECT 79.97 1.965 80.32 2.315 ;
      RECT 68.86 8.29 79.04 8.46 ;
      RECT 78.88 2.395 79.04 8.46 ;
      RECT 68.86 6.6 69.03 8.46 ;
      RECT 79.995 6.655 80.32 6.98 ;
      RECT 65.805 6.655 66.13 6.98 ;
      RECT 68.805 6.6 69.085 6.94 ;
      RECT 78.88 6.745 80.32 6.915 ;
      RECT 65.805 6.685 69.085 6.855 ;
      RECT 79.195 2.365 79.515 2.685 ;
      RECT 78.88 2.395 79.515 2.565 ;
      RECT 72.815 2.37 73.095 2.74 ;
      RECT 72.86 1.605 73.03 2.74 ;
      RECT 77.525 1.995 77.85 2.32 ;
      RECT 77.6 1.605 77.77 2.32 ;
      RECT 72.86 1.605 77.77 1.775 ;
      RECT 76.555 4.78 76.815 5.1 ;
      RECT 76.615 2.74 76.755 5.1 ;
      RECT 76.555 2.74 76.815 3.06 ;
      RECT 75.535 5.8 75.795 6.12 ;
      RECT 74.915 5.89 75.795 6.03 ;
      RECT 74.915 3.735 75.055 6.03 ;
      RECT 74.855 3.735 75.135 4.105 ;
      RECT 74.175 5.775 74.455 6.145 ;
      RECT 74.235 3.85 74.375 6.145 ;
      RECT 74.235 3.85 74.715 3.99 ;
      RECT 74.575 2.06 74.715 3.99 ;
      RECT 74.515 2.06 74.775 2.38 ;
      RECT 73.495 4.755 73.775 5.125 ;
      RECT 73.555 2.4 73.695 5.125 ;
      RECT 73.495 2.4 73.755 2.72 ;
      RECT 73.13 5.775 73.41 6.145 ;
      RECT 73.13 5.8 73.415 6.12 ;
      RECT 68.275 6.995 68.645 7.365 ;
      RECT 68.275 6.995 68.65 7.005 ;
      RECT 62.615 6.28 62.935 6.605 ;
      RECT 62.645 5.695 62.815 6.605 ;
      RECT 62.645 5.695 62.82 6.045 ;
      RECT 62.645 5.695 63.62 5.87 ;
      RECT 63.445 1.965 63.62 5.87 ;
      RECT 63.39 1.965 63.74 2.315 ;
      RECT 52.28 8.29 62.46 8.46 ;
      RECT 62.3 2.395 62.46 8.46 ;
      RECT 52.28 6.6 52.45 8.46 ;
      RECT 63.415 6.655 63.74 6.98 ;
      RECT 49.22 6.655 49.545 6.98 ;
      RECT 52.225 6.6 52.505 6.94 ;
      RECT 62.3 6.745 63.74 6.915 ;
      RECT 49.22 6.685 52.505 6.855 ;
      RECT 62.615 2.365 62.935 2.685 ;
      RECT 62.3 2.395 62.935 2.565 ;
      RECT 56.235 2.37 56.515 2.74 ;
      RECT 56.28 1.605 56.45 2.74 ;
      RECT 60.945 1.995 61.27 2.32 ;
      RECT 61.02 1.605 61.19 2.32 ;
      RECT 56.28 1.605 61.19 1.775 ;
      RECT 59.975 4.78 60.235 5.1 ;
      RECT 60.035 2.74 60.175 5.1 ;
      RECT 59.975 2.74 60.235 3.06 ;
      RECT 58.955 5.8 59.215 6.12 ;
      RECT 58.335 5.89 59.215 6.03 ;
      RECT 58.335 3.735 58.475 6.03 ;
      RECT 58.275 3.735 58.555 4.105 ;
      RECT 57.595 5.775 57.875 6.145 ;
      RECT 57.655 3.85 57.795 6.145 ;
      RECT 57.655 3.85 58.135 3.99 ;
      RECT 57.995 2.06 58.135 3.99 ;
      RECT 57.935 2.06 58.195 2.38 ;
      RECT 56.915 4.755 57.195 5.125 ;
      RECT 56.975 2.4 57.115 5.125 ;
      RECT 56.915 2.4 57.175 2.72 ;
      RECT 56.55 5.775 56.83 6.145 ;
      RECT 56.55 5.8 56.835 6.12 ;
      RECT 46.03 6.28 46.35 6.605 ;
      RECT 46.06 5.695 46.23 6.605 ;
      RECT 46.06 5.695 46.235 6.045 ;
      RECT 46.06 5.695 47.035 5.87 ;
      RECT 46.86 1.965 47.035 5.87 ;
      RECT 46.805 1.965 47.155 2.315 ;
      RECT 35.695 8.29 45.875 8.46 ;
      RECT 45.715 2.395 45.875 8.46 ;
      RECT 35.695 6.6 35.865 8.46 ;
      RECT 46.83 6.655 47.155 6.98 ;
      RECT 32.635 6.655 32.96 6.98 ;
      RECT 35.64 6.6 35.92 6.94 ;
      RECT 45.715 6.745 47.155 6.915 ;
      RECT 32.635 6.685 35.92 6.855 ;
      RECT 46.03 2.365 46.35 2.685 ;
      RECT 45.715 2.395 46.35 2.565 ;
      RECT 39.65 2.37 39.93 2.74 ;
      RECT 39.695 1.605 39.865 2.74 ;
      RECT 44.36 1.995 44.685 2.32 ;
      RECT 44.435 1.605 44.605 2.32 ;
      RECT 39.695 1.605 44.605 1.775 ;
      RECT 43.39 4.78 43.65 5.1 ;
      RECT 43.45 2.74 43.59 5.1 ;
      RECT 43.39 2.74 43.65 3.06 ;
      RECT 42.37 5.8 42.63 6.12 ;
      RECT 41.75 5.89 42.63 6.03 ;
      RECT 41.75 3.735 41.89 6.03 ;
      RECT 41.69 3.735 41.97 4.105 ;
      RECT 41.01 5.775 41.29 6.145 ;
      RECT 41.07 3.85 41.21 6.145 ;
      RECT 41.07 3.85 41.55 3.99 ;
      RECT 41.41 2.06 41.55 3.99 ;
      RECT 41.35 2.06 41.61 2.38 ;
      RECT 40.33 4.755 40.61 5.125 ;
      RECT 40.39 2.4 40.53 5.125 ;
      RECT 40.33 2.4 40.59 2.72 ;
      RECT 39.965 5.775 40.245 6.145 ;
      RECT 39.965 5.8 40.25 6.12 ;
      RECT 29.445 6.28 29.765 6.605 ;
      RECT 29.475 5.695 29.645 6.605 ;
      RECT 29.475 5.695 29.65 6.045 ;
      RECT 29.475 5.695 30.45 5.87 ;
      RECT 30.275 1.965 30.45 5.87 ;
      RECT 30.22 1.965 30.57 2.315 ;
      RECT 19.11 8.29 29.29 8.46 ;
      RECT 29.13 2.395 29.29 8.46 ;
      RECT 19.11 6.6 19.28 8.46 ;
      RECT 30.245 6.655 30.57 6.98 ;
      RECT 16.05 6.655 16.375 6.98 ;
      RECT 19.055 6.6 19.335 6.94 ;
      RECT 29.13 6.745 30.57 6.915 ;
      RECT 16.05 6.685 19.335 6.855 ;
      RECT 29.445 2.365 29.765 2.685 ;
      RECT 29.13 2.395 29.765 2.565 ;
      RECT 23.065 2.37 23.345 2.74 ;
      RECT 23.11 1.605 23.28 2.74 ;
      RECT 27.775 1.995 28.1 2.32 ;
      RECT 27.85 1.605 28.02 2.32 ;
      RECT 23.11 1.605 28.02 1.775 ;
      RECT 26.805 4.78 27.065 5.1 ;
      RECT 26.865 2.74 27.005 5.1 ;
      RECT 26.805 2.74 27.065 3.06 ;
      RECT 25.785 5.8 26.045 6.12 ;
      RECT 25.165 5.89 26.045 6.03 ;
      RECT 25.165 3.735 25.305 6.03 ;
      RECT 25.105 3.735 25.385 4.105 ;
      RECT 24.425 5.775 24.705 6.145 ;
      RECT 24.485 3.85 24.625 6.145 ;
      RECT 24.485 3.85 24.965 3.99 ;
      RECT 24.825 2.06 24.965 3.99 ;
      RECT 24.765 2.06 25.025 2.38 ;
      RECT 23.745 4.755 24.025 5.125 ;
      RECT 23.805 2.4 23.945 5.125 ;
      RECT 23.745 2.4 24.005 2.72 ;
      RECT 23.38 5.775 23.66 6.145 ;
      RECT 23.38 5.8 23.665 6.12 ;
      RECT 12.86 6.28 13.18 6.605 ;
      RECT 12.89 5.695 13.06 6.605 ;
      RECT 12.89 5.695 13.065 6.045 ;
      RECT 12.89 5.695 13.865 5.87 ;
      RECT 13.69 1.965 13.865 5.87 ;
      RECT 13.635 1.965 13.985 2.315 ;
      RECT 2.525 8.29 12.705 8.46 ;
      RECT 12.545 2.395 12.705 8.46 ;
      RECT 2.525 6.6 2.695 8.46 ;
      RECT -1.24 6.995 -0.96 7.335 ;
      RECT -1.24 7.06 -0.05 7.23 ;
      RECT -0.22 6.685 -0.05 7.23 ;
      RECT 13.66 6.655 13.985 6.98 ;
      RECT 2.47 6.6 2.75 6.94 ;
      RECT 12.545 6.745 13.985 6.915 ;
      RECT -0.22 6.685 2.75 6.855 ;
      RECT 12.86 2.365 13.18 2.685 ;
      RECT 12.545 2.395 13.18 2.565 ;
      RECT 6.48 2.37 6.76 2.74 ;
      RECT 6.525 1.605 6.695 2.74 ;
      RECT 11.19 1.995 11.515 2.32 ;
      RECT 11.265 1.605 11.435 2.32 ;
      RECT 6.525 1.605 11.435 1.775 ;
      RECT 10.22 4.78 10.48 5.1 ;
      RECT 10.28 2.74 10.42 5.1 ;
      RECT 10.22 2.74 10.48 3.06 ;
      RECT 9.2 5.8 9.46 6.12 ;
      RECT 8.58 5.89 9.46 6.03 ;
      RECT 8.58 3.735 8.72 6.03 ;
      RECT 8.52 3.735 8.8 4.105 ;
      RECT 7.84 5.775 8.12 6.145 ;
      RECT 7.9 3.85 8.04 6.145 ;
      RECT 7.9 3.85 8.38 3.99 ;
      RECT 8.24 2.06 8.38 3.99 ;
      RECT 8.18 2.06 8.44 2.38 ;
      RECT 7.16 4.755 7.44 5.125 ;
      RECT 7.22 2.4 7.36 5.125 ;
      RECT 7.16 2.4 7.42 2.72 ;
      RECT 6.795 5.775 7.075 6.145 ;
      RECT 6.795 5.8 7.08 6.12 ;
      RECT 74.855 2.715 75.135 3.085 ;
      RECT 74.155 3.055 74.435 3.425 ;
      RECT 58.275 2.715 58.555 3.085 ;
      RECT 57.575 3.055 57.855 3.425 ;
      RECT 51.695 6.995 52.065 7.365 ;
      RECT 41.69 2.715 41.97 3.085 ;
      RECT 40.99 3.055 41.27 3.425 ;
      RECT 35.11 6.995 35.48 7.365 ;
      RECT 25.105 2.715 25.385 3.085 ;
      RECT 24.405 3.055 24.685 3.425 ;
      RECT 18.525 6.995 18.895 7.365 ;
      RECT 8.52 2.715 8.8 3.085 ;
      RECT 7.82 3.055 8.1 3.425 ;
      RECT 1.94 6.995 2.31 7.365 ;
    LAYER via1 ;
      RECT 82.44 7.385 82.59 7.535 ;
      RECT 80.085 6.74 80.235 6.89 ;
      RECT 80.07 2.065 80.22 2.215 ;
      RECT 79.28 2.45 79.43 2.6 ;
      RECT 79.28 6.37 79.43 6.52 ;
      RECT 77.615 2.08 77.765 2.23 ;
      RECT 76.61 2.825 76.76 2.975 ;
      RECT 76.61 4.865 76.76 5.015 ;
      RECT 75.59 5.885 75.74 6.035 ;
      RECT 74.91 2.825 75.06 2.975 ;
      RECT 74.91 3.845 75.06 3.995 ;
      RECT 74.57 2.145 74.72 2.295 ;
      RECT 74.23 3.165 74.38 3.315 ;
      RECT 74.23 5.885 74.38 6.035 ;
      RECT 73.55 2.485 73.7 2.635 ;
      RECT 73.55 4.865 73.7 5.015 ;
      RECT 73.21 5.885 73.36 6.035 ;
      RECT 72.87 2.48 73.02 2.63 ;
      RECT 68.87 6.695 69.02 6.845 ;
      RECT 68.385 7.105 68.535 7.255 ;
      RECT 65.895 6.74 66.045 6.89 ;
      RECT 63.505 6.74 63.655 6.89 ;
      RECT 63.49 2.065 63.64 2.215 ;
      RECT 62.7 2.45 62.85 2.6 ;
      RECT 62.7 6.37 62.85 6.52 ;
      RECT 61.035 2.08 61.185 2.23 ;
      RECT 60.03 2.825 60.18 2.975 ;
      RECT 60.03 4.865 60.18 5.015 ;
      RECT 59.01 5.885 59.16 6.035 ;
      RECT 58.33 2.825 58.48 2.975 ;
      RECT 58.33 3.845 58.48 3.995 ;
      RECT 57.99 2.145 58.14 2.295 ;
      RECT 57.65 3.165 57.8 3.315 ;
      RECT 57.65 5.885 57.8 6.035 ;
      RECT 56.97 2.485 57.12 2.635 ;
      RECT 56.97 4.865 57.12 5.015 ;
      RECT 56.63 5.885 56.78 6.035 ;
      RECT 56.29 2.48 56.44 2.63 ;
      RECT 52.29 6.695 52.44 6.845 ;
      RECT 51.805 7.105 51.955 7.255 ;
      RECT 49.31 6.74 49.46 6.89 ;
      RECT 46.92 6.74 47.07 6.89 ;
      RECT 46.905 2.065 47.055 2.215 ;
      RECT 46.115 2.45 46.265 2.6 ;
      RECT 46.115 6.37 46.265 6.52 ;
      RECT 44.45 2.08 44.6 2.23 ;
      RECT 43.445 2.825 43.595 2.975 ;
      RECT 43.445 4.865 43.595 5.015 ;
      RECT 42.425 5.885 42.575 6.035 ;
      RECT 41.745 2.825 41.895 2.975 ;
      RECT 41.745 3.845 41.895 3.995 ;
      RECT 41.405 2.145 41.555 2.295 ;
      RECT 41.065 3.165 41.215 3.315 ;
      RECT 41.065 5.885 41.215 6.035 ;
      RECT 40.385 2.485 40.535 2.635 ;
      RECT 40.385 4.865 40.535 5.015 ;
      RECT 40.045 5.885 40.195 6.035 ;
      RECT 39.705 2.48 39.855 2.63 ;
      RECT 35.705 6.695 35.855 6.845 ;
      RECT 35.22 7.105 35.37 7.255 ;
      RECT 32.725 6.74 32.875 6.89 ;
      RECT 30.335 6.74 30.485 6.89 ;
      RECT 30.32 2.065 30.47 2.215 ;
      RECT 29.53 2.45 29.68 2.6 ;
      RECT 29.53 6.37 29.68 6.52 ;
      RECT 27.865 2.08 28.015 2.23 ;
      RECT 26.86 2.825 27.01 2.975 ;
      RECT 26.86 4.865 27.01 5.015 ;
      RECT 25.84 5.885 25.99 6.035 ;
      RECT 25.16 2.825 25.31 2.975 ;
      RECT 25.16 3.845 25.31 3.995 ;
      RECT 24.82 2.145 24.97 2.295 ;
      RECT 24.48 3.165 24.63 3.315 ;
      RECT 24.48 5.885 24.63 6.035 ;
      RECT 23.8 2.485 23.95 2.635 ;
      RECT 23.8 4.865 23.95 5.015 ;
      RECT 23.46 5.885 23.61 6.035 ;
      RECT 23.12 2.48 23.27 2.63 ;
      RECT 19.12 6.695 19.27 6.845 ;
      RECT 18.635 7.105 18.785 7.255 ;
      RECT 16.14 6.74 16.29 6.89 ;
      RECT 13.75 6.74 13.9 6.89 ;
      RECT 13.735 2.065 13.885 2.215 ;
      RECT 12.945 2.45 13.095 2.6 ;
      RECT 12.945 6.37 13.095 6.52 ;
      RECT 11.28 2.08 11.43 2.23 ;
      RECT 10.275 2.825 10.425 2.975 ;
      RECT 10.275 4.865 10.425 5.015 ;
      RECT 9.255 5.885 9.405 6.035 ;
      RECT 8.575 2.825 8.725 2.975 ;
      RECT 8.575 3.845 8.725 3.995 ;
      RECT 8.235 2.145 8.385 2.295 ;
      RECT 7.895 3.165 8.045 3.315 ;
      RECT 7.895 5.885 8.045 6.035 ;
      RECT 7.215 2.485 7.365 2.635 ;
      RECT 7.215 4.865 7.365 5.015 ;
      RECT 6.875 5.885 7.025 6.035 ;
      RECT 6.535 2.48 6.685 2.63 ;
      RECT 2.535 6.695 2.685 6.845 ;
      RECT 2.05 7.105 2.2 7.255 ;
      RECT -1.175 7.09 -1.025 7.24 ;
      RECT -1.56 6.35 -1.41 6.5 ;
    LAYER met1 ;
      RECT 82.32 7.77 82.61 8 ;
      RECT 82.38 6.29 82.55 8 ;
      RECT 82.35 7.3 82.675 7.625 ;
      RECT 82.32 6.29 82.61 6.52 ;
      RECT 81.915 2.395 82.02 2.965 ;
      RECT 81.915 2.73 82.24 2.96 ;
      RECT 81.915 2.76 82.41 2.93 ;
      RECT 81.915 2.395 82.105 2.96 ;
      RECT 81.33 2.36 81.62 2.59 ;
      RECT 81.33 2.395 82.105 2.565 ;
      RECT 81.39 0.88 81.56 2.59 ;
      RECT 81.33 0.88 81.62 1.11 ;
      RECT 81.33 7.77 81.62 8 ;
      RECT 81.39 6.29 81.56 8 ;
      RECT 81.33 6.29 81.62 6.52 ;
      RECT 81.33 6.325 82.185 6.485 ;
      RECT 82.015 5.92 82.185 6.485 ;
      RECT 81.33 6.32 81.725 6.485 ;
      RECT 81.95 5.92 82.24 6.15 ;
      RECT 81.95 5.95 82.41 6.12 ;
      RECT 80.96 2.73 81.25 2.96 ;
      RECT 80.96 2.76 81.42 2.93 ;
      RECT 81.025 1.655 81.19 2.96 ;
      RECT 79.54 1.625 79.83 1.855 ;
      RECT 79.54 1.655 81.19 1.825 ;
      RECT 79.6 0.885 79.77 1.855 ;
      RECT 79.54 0.885 79.83 1.115 ;
      RECT 79.54 7.765 79.83 7.995 ;
      RECT 79.6 7.025 79.77 7.995 ;
      RECT 79.6 7.12 81.19 7.29 ;
      RECT 81.02 5.92 81.19 7.29 ;
      RECT 79.54 7.025 79.83 7.255 ;
      RECT 80.96 5.92 81.25 6.15 ;
      RECT 80.96 5.95 81.42 6.12 ;
      RECT 77.525 1.995 77.85 2.32 ;
      RECT 79.97 1.965 80.32 2.315 ;
      RECT 77.525 2.025 80.32 2.195 ;
      RECT 79.995 6.655 80.32 6.98 ;
      RECT 79.97 6.655 80.32 6.885 ;
      RECT 79.8 6.685 80.32 6.855 ;
      RECT 79.195 2.365 79.515 2.685 ;
      RECT 79.165 2.365 79.515 2.595 ;
      RECT 78.88 2.395 79.515 2.565 ;
      RECT 79.195 6.28 79.515 6.605 ;
      RECT 79.165 6.285 79.515 6.515 ;
      RECT 78.995 6.315 79.515 6.485 ;
      RECT 76.525 2.77 76.845 3.03 ;
      RECT 76.25 2.83 76.845 2.97 ;
      RECT 74.145 3.11 74.465 3.37 ;
      RECT 76.12 3.125 76.41 3.355 ;
      RECT 74.145 3.17 76.41 3.31 ;
      RECT 75.505 5.83 75.825 6.09 ;
      RECT 75.505 5.89 76.1 6.03 ;
      RECT 74.825 2.77 75.145 3.03 ;
      RECT 70.085 2.785 70.375 3.015 ;
      RECT 70.085 2.83 75.145 2.97 ;
      RECT 74.915 2.49 75.055 3.03 ;
      RECT 74.915 2.49 75.395 2.63 ;
      RECT 75.255 2.105 75.395 2.63 ;
      RECT 75.18 2.105 75.47 2.335 ;
      RECT 74.825 3.79 75.145 4.05 ;
      RECT 74.16 3.805 74.45 4.035 ;
      RECT 71.95 3.805 72.24 4.035 ;
      RECT 71.95 3.85 75.145 3.99 ;
      RECT 73.125 5.83 73.445 6.09 ;
      RECT 74.84 5.845 75.13 6.075 ;
      RECT 72.46 5.845 72.75 6.075 ;
      RECT 72.46 5.89 73.445 6.03 ;
      RECT 74.915 5.55 75.055 6.075 ;
      RECT 73.215 5.55 73.355 6.09 ;
      RECT 73.215 5.55 75.055 5.69 ;
      RECT 72.12 2.445 72.41 2.675 ;
      RECT 72.195 2.15 72.335 2.675 ;
      RECT 74.485 2.09 74.805 2.35 ;
      RECT 74.385 2.105 74.805 2.335 ;
      RECT 72.195 2.15 74.805 2.29 ;
      RECT 73.465 2.43 73.785 2.69 ;
      RECT 73.465 2.49 74.06 2.63 ;
      RECT 73.465 4.81 73.785 5.07 ;
      RECT 70.76 4.825 71.05 5.055 ;
      RECT 70.76 4.87 73.785 5.01 ;
      RECT 72.79 2.39 73.12 2.72 ;
      RECT 72.785 2.425 73.12 2.685 ;
      RECT 73.135 2.445 73.25 2.675 ;
      RECT 72.785 2.44 73.135 2.67 ;
      RECT 72.785 2.49 73.265 2.63 ;
      RECT 72.67 2.49 72.68 2.63 ;
      RECT 72.68 2.485 73.25 2.625 ;
      RECT 68.775 6.63 69.115 6.91 ;
      RECT 68.745 6.655 69.115 6.885 ;
      RECT 68.575 6.685 69.115 6.855 ;
      RECT 68.315 7.765 68.605 7.995 ;
      RECT 68.375 6.995 68.545 7.995 ;
      RECT 68.275 6.995 68.645 7.365 ;
      RECT 65.74 7.77 66.03 8 ;
      RECT 65.8 6.29 65.97 8 ;
      RECT 65.8 6.655 66.13 6.98 ;
      RECT 65.74 6.29 66.03 6.52 ;
      RECT 65.335 2.395 65.44 2.965 ;
      RECT 65.335 2.73 65.66 2.96 ;
      RECT 65.335 2.76 65.83 2.93 ;
      RECT 65.335 2.395 65.525 2.96 ;
      RECT 64.75 2.36 65.04 2.59 ;
      RECT 64.75 2.395 65.525 2.565 ;
      RECT 64.81 0.88 64.98 2.59 ;
      RECT 64.75 0.88 65.04 1.11 ;
      RECT 64.75 7.77 65.04 8 ;
      RECT 64.81 6.29 64.98 8 ;
      RECT 64.75 6.29 65.04 6.52 ;
      RECT 64.75 6.325 65.605 6.485 ;
      RECT 65.435 5.92 65.605 6.485 ;
      RECT 64.75 6.32 65.145 6.485 ;
      RECT 65.37 5.92 65.66 6.15 ;
      RECT 65.37 5.95 65.83 6.12 ;
      RECT 64.38 2.73 64.67 2.96 ;
      RECT 64.38 2.76 64.84 2.93 ;
      RECT 64.445 1.655 64.61 2.96 ;
      RECT 62.96 1.625 63.25 1.855 ;
      RECT 62.96 1.655 64.61 1.825 ;
      RECT 63.02 0.885 63.19 1.855 ;
      RECT 62.96 0.885 63.25 1.115 ;
      RECT 62.96 7.765 63.25 7.995 ;
      RECT 63.02 7.025 63.19 7.995 ;
      RECT 63.02 7.12 64.61 7.29 ;
      RECT 64.44 5.92 64.61 7.29 ;
      RECT 62.96 7.025 63.25 7.255 ;
      RECT 64.38 5.92 64.67 6.15 ;
      RECT 64.38 5.95 64.84 6.12 ;
      RECT 60.945 1.995 61.27 2.32 ;
      RECT 63.39 1.965 63.74 2.315 ;
      RECT 60.945 2.025 63.74 2.195 ;
      RECT 63.415 6.655 63.74 6.98 ;
      RECT 63.39 6.655 63.74 6.885 ;
      RECT 63.22 6.685 63.74 6.855 ;
      RECT 62.615 2.365 62.935 2.685 ;
      RECT 62.585 2.365 62.935 2.595 ;
      RECT 62.3 2.395 62.935 2.565 ;
      RECT 62.615 6.28 62.935 6.605 ;
      RECT 62.585 6.285 62.935 6.515 ;
      RECT 62.415 6.315 62.935 6.485 ;
      RECT 59.945 2.77 60.265 3.03 ;
      RECT 59.67 2.83 60.265 2.97 ;
      RECT 57.565 3.11 57.885 3.37 ;
      RECT 59.54 3.125 59.83 3.355 ;
      RECT 57.565 3.17 59.83 3.31 ;
      RECT 58.925 5.83 59.245 6.09 ;
      RECT 58.925 5.89 59.52 6.03 ;
      RECT 58.245 2.77 58.565 3.03 ;
      RECT 53.505 2.785 53.795 3.015 ;
      RECT 53.505 2.83 58.565 2.97 ;
      RECT 58.335 2.49 58.475 3.03 ;
      RECT 58.335 2.49 58.815 2.63 ;
      RECT 58.675 2.105 58.815 2.63 ;
      RECT 58.6 2.105 58.89 2.335 ;
      RECT 58.245 3.79 58.565 4.05 ;
      RECT 57.58 3.805 57.87 4.035 ;
      RECT 55.37 3.805 55.66 4.035 ;
      RECT 55.37 3.85 58.565 3.99 ;
      RECT 56.545 5.83 56.865 6.09 ;
      RECT 58.26 5.845 58.55 6.075 ;
      RECT 55.88 5.845 56.17 6.075 ;
      RECT 55.88 5.89 56.865 6.03 ;
      RECT 58.335 5.55 58.475 6.075 ;
      RECT 56.635 5.55 56.775 6.09 ;
      RECT 56.635 5.55 58.475 5.69 ;
      RECT 55.54 2.445 55.83 2.675 ;
      RECT 55.615 2.15 55.755 2.675 ;
      RECT 57.905 2.09 58.225 2.35 ;
      RECT 57.805 2.105 58.225 2.335 ;
      RECT 55.615 2.15 58.225 2.29 ;
      RECT 56.885 2.43 57.205 2.69 ;
      RECT 56.885 2.49 57.48 2.63 ;
      RECT 56.885 4.81 57.205 5.07 ;
      RECT 54.18 4.825 54.47 5.055 ;
      RECT 54.18 4.87 57.205 5.01 ;
      RECT 56.21 2.39 56.54 2.72 ;
      RECT 56.205 2.425 56.54 2.685 ;
      RECT 56.555 2.445 56.67 2.675 ;
      RECT 56.205 2.44 56.555 2.67 ;
      RECT 56.205 2.49 56.685 2.63 ;
      RECT 56.09 2.49 56.1 2.63 ;
      RECT 56.1 2.485 56.67 2.625 ;
      RECT 52.195 6.63 52.535 6.91 ;
      RECT 52.165 6.655 52.535 6.885 ;
      RECT 51.995 6.685 52.535 6.855 ;
      RECT 51.735 7.765 52.025 7.995 ;
      RECT 51.795 6.995 51.965 7.995 ;
      RECT 51.695 6.995 52.065 7.365 ;
      RECT 49.155 7.77 49.445 8 ;
      RECT 49.215 6.29 49.385 8 ;
      RECT 49.215 6.655 49.545 6.98 ;
      RECT 49.155 6.29 49.445 6.52 ;
      RECT 48.75 2.395 48.855 2.965 ;
      RECT 48.75 2.73 49.075 2.96 ;
      RECT 48.75 2.76 49.245 2.93 ;
      RECT 48.75 2.395 48.94 2.96 ;
      RECT 48.165 2.36 48.455 2.59 ;
      RECT 48.165 2.395 48.94 2.565 ;
      RECT 48.225 0.88 48.395 2.59 ;
      RECT 48.165 0.88 48.455 1.11 ;
      RECT 48.165 7.77 48.455 8 ;
      RECT 48.225 6.29 48.395 8 ;
      RECT 48.165 6.29 48.455 6.52 ;
      RECT 48.165 6.325 49.02 6.485 ;
      RECT 48.85 5.92 49.02 6.485 ;
      RECT 48.165 6.32 48.56 6.485 ;
      RECT 48.785 5.92 49.075 6.15 ;
      RECT 48.785 5.95 49.245 6.12 ;
      RECT 47.795 2.73 48.085 2.96 ;
      RECT 47.795 2.76 48.255 2.93 ;
      RECT 47.86 1.655 48.025 2.96 ;
      RECT 46.375 1.625 46.665 1.855 ;
      RECT 46.375 1.655 48.025 1.825 ;
      RECT 46.435 0.885 46.605 1.855 ;
      RECT 46.375 0.885 46.665 1.115 ;
      RECT 46.375 7.765 46.665 7.995 ;
      RECT 46.435 7.025 46.605 7.995 ;
      RECT 46.435 7.12 48.025 7.29 ;
      RECT 47.855 5.92 48.025 7.29 ;
      RECT 46.375 7.025 46.665 7.255 ;
      RECT 47.795 5.92 48.085 6.15 ;
      RECT 47.795 5.95 48.255 6.12 ;
      RECT 44.36 1.995 44.685 2.32 ;
      RECT 46.805 1.965 47.155 2.315 ;
      RECT 44.36 2.025 47.155 2.195 ;
      RECT 46.83 6.655 47.155 6.98 ;
      RECT 46.805 6.655 47.155 6.885 ;
      RECT 46.635 6.685 47.155 6.855 ;
      RECT 46.03 2.365 46.35 2.685 ;
      RECT 46 2.365 46.35 2.595 ;
      RECT 45.715 2.395 46.35 2.565 ;
      RECT 46.03 6.28 46.35 6.605 ;
      RECT 46 6.285 46.35 6.515 ;
      RECT 45.83 6.315 46.35 6.485 ;
      RECT 43.36 2.77 43.68 3.03 ;
      RECT 43.085 2.83 43.68 2.97 ;
      RECT 40.98 3.11 41.3 3.37 ;
      RECT 42.955 3.125 43.245 3.355 ;
      RECT 40.98 3.17 43.245 3.31 ;
      RECT 42.34 5.83 42.66 6.09 ;
      RECT 42.34 5.89 42.935 6.03 ;
      RECT 41.66 2.77 41.98 3.03 ;
      RECT 36.92 2.785 37.21 3.015 ;
      RECT 36.92 2.83 41.98 2.97 ;
      RECT 41.75 2.49 41.89 3.03 ;
      RECT 41.75 2.49 42.23 2.63 ;
      RECT 42.09 2.105 42.23 2.63 ;
      RECT 42.015 2.105 42.305 2.335 ;
      RECT 41.66 3.79 41.98 4.05 ;
      RECT 40.995 3.805 41.285 4.035 ;
      RECT 38.785 3.805 39.075 4.035 ;
      RECT 38.785 3.85 41.98 3.99 ;
      RECT 39.96 5.83 40.28 6.09 ;
      RECT 41.675 5.845 41.965 6.075 ;
      RECT 39.295 5.845 39.585 6.075 ;
      RECT 39.295 5.89 40.28 6.03 ;
      RECT 41.75 5.55 41.89 6.075 ;
      RECT 40.05 5.55 40.19 6.09 ;
      RECT 40.05 5.55 41.89 5.69 ;
      RECT 38.955 2.445 39.245 2.675 ;
      RECT 39.03 2.15 39.17 2.675 ;
      RECT 41.32 2.09 41.64 2.35 ;
      RECT 41.22 2.105 41.64 2.335 ;
      RECT 39.03 2.15 41.64 2.29 ;
      RECT 40.3 2.43 40.62 2.69 ;
      RECT 40.3 2.49 40.895 2.63 ;
      RECT 40.3 4.81 40.62 5.07 ;
      RECT 37.595 4.825 37.885 5.055 ;
      RECT 37.595 4.87 40.62 5.01 ;
      RECT 39.625 2.39 39.955 2.72 ;
      RECT 39.62 2.425 39.955 2.685 ;
      RECT 39.97 2.445 40.085 2.675 ;
      RECT 39.62 2.44 39.97 2.67 ;
      RECT 39.62 2.49 40.1 2.63 ;
      RECT 39.505 2.49 39.515 2.63 ;
      RECT 39.515 2.485 40.085 2.625 ;
      RECT 35.61 6.63 35.95 6.91 ;
      RECT 35.58 6.655 35.95 6.885 ;
      RECT 35.41 6.685 35.95 6.855 ;
      RECT 35.15 7.765 35.44 7.995 ;
      RECT 35.21 6.995 35.38 7.995 ;
      RECT 35.11 6.995 35.48 7.365 ;
      RECT 32.57 7.77 32.86 8 ;
      RECT 32.63 6.29 32.8 8 ;
      RECT 32.63 6.655 32.96 6.98 ;
      RECT 32.57 6.29 32.86 6.52 ;
      RECT 32.165 2.395 32.27 2.965 ;
      RECT 32.165 2.73 32.49 2.96 ;
      RECT 32.165 2.76 32.66 2.93 ;
      RECT 32.165 2.395 32.355 2.96 ;
      RECT 31.58 2.36 31.87 2.59 ;
      RECT 31.58 2.395 32.355 2.565 ;
      RECT 31.64 0.88 31.81 2.59 ;
      RECT 31.58 0.88 31.87 1.11 ;
      RECT 31.58 7.77 31.87 8 ;
      RECT 31.64 6.29 31.81 8 ;
      RECT 31.58 6.29 31.87 6.52 ;
      RECT 31.58 6.325 32.435 6.485 ;
      RECT 32.265 5.92 32.435 6.485 ;
      RECT 31.58 6.32 31.975 6.485 ;
      RECT 32.2 5.92 32.49 6.15 ;
      RECT 32.2 5.95 32.66 6.12 ;
      RECT 31.21 2.73 31.5 2.96 ;
      RECT 31.21 2.76 31.67 2.93 ;
      RECT 31.275 1.655 31.44 2.96 ;
      RECT 29.79 1.625 30.08 1.855 ;
      RECT 29.79 1.655 31.44 1.825 ;
      RECT 29.85 0.885 30.02 1.855 ;
      RECT 29.79 0.885 30.08 1.115 ;
      RECT 29.79 7.765 30.08 7.995 ;
      RECT 29.85 7.025 30.02 7.995 ;
      RECT 29.85 7.12 31.44 7.29 ;
      RECT 31.27 5.92 31.44 7.29 ;
      RECT 29.79 7.025 30.08 7.255 ;
      RECT 31.21 5.92 31.5 6.15 ;
      RECT 31.21 5.95 31.67 6.12 ;
      RECT 27.775 1.995 28.1 2.32 ;
      RECT 30.22 1.965 30.57 2.315 ;
      RECT 27.775 2.025 30.57 2.195 ;
      RECT 30.245 6.655 30.57 6.98 ;
      RECT 30.22 6.655 30.57 6.885 ;
      RECT 30.05 6.685 30.57 6.855 ;
      RECT 29.445 2.365 29.765 2.685 ;
      RECT 29.415 2.365 29.765 2.595 ;
      RECT 29.13 2.395 29.765 2.565 ;
      RECT 29.445 6.28 29.765 6.605 ;
      RECT 29.415 6.285 29.765 6.515 ;
      RECT 29.245 6.315 29.765 6.485 ;
      RECT 26.775 2.77 27.095 3.03 ;
      RECT 26.5 2.83 27.095 2.97 ;
      RECT 24.395 3.11 24.715 3.37 ;
      RECT 26.37 3.125 26.66 3.355 ;
      RECT 24.395 3.17 26.66 3.31 ;
      RECT 25.755 5.83 26.075 6.09 ;
      RECT 25.755 5.89 26.35 6.03 ;
      RECT 25.075 2.77 25.395 3.03 ;
      RECT 20.335 2.785 20.625 3.015 ;
      RECT 20.335 2.83 25.395 2.97 ;
      RECT 25.165 2.49 25.305 3.03 ;
      RECT 25.165 2.49 25.645 2.63 ;
      RECT 25.505 2.105 25.645 2.63 ;
      RECT 25.43 2.105 25.72 2.335 ;
      RECT 25.075 3.79 25.395 4.05 ;
      RECT 24.41 3.805 24.7 4.035 ;
      RECT 22.2 3.805 22.49 4.035 ;
      RECT 22.2 3.85 25.395 3.99 ;
      RECT 23.375 5.83 23.695 6.09 ;
      RECT 25.09 5.845 25.38 6.075 ;
      RECT 22.71 5.845 23 6.075 ;
      RECT 22.71 5.89 23.695 6.03 ;
      RECT 25.165 5.55 25.305 6.075 ;
      RECT 23.465 5.55 23.605 6.09 ;
      RECT 23.465 5.55 25.305 5.69 ;
      RECT 22.37 2.445 22.66 2.675 ;
      RECT 22.445 2.15 22.585 2.675 ;
      RECT 24.735 2.09 25.055 2.35 ;
      RECT 24.635 2.105 25.055 2.335 ;
      RECT 22.445 2.15 25.055 2.29 ;
      RECT 23.715 2.43 24.035 2.69 ;
      RECT 23.715 2.49 24.31 2.63 ;
      RECT 23.715 4.81 24.035 5.07 ;
      RECT 21.01 4.825 21.3 5.055 ;
      RECT 21.01 4.87 24.035 5.01 ;
      RECT 23.04 2.39 23.37 2.72 ;
      RECT 23.035 2.425 23.37 2.685 ;
      RECT 23.385 2.445 23.5 2.675 ;
      RECT 23.035 2.44 23.385 2.67 ;
      RECT 23.035 2.49 23.515 2.63 ;
      RECT 22.92 2.49 22.93 2.63 ;
      RECT 22.93 2.485 23.5 2.625 ;
      RECT 19.025 6.63 19.365 6.91 ;
      RECT 18.995 6.655 19.365 6.885 ;
      RECT 18.825 6.685 19.365 6.855 ;
      RECT 18.565 7.765 18.855 7.995 ;
      RECT 18.625 6.995 18.795 7.995 ;
      RECT 18.525 6.995 18.895 7.365 ;
      RECT 15.985 7.77 16.275 8 ;
      RECT 16.045 6.29 16.215 8 ;
      RECT 16.045 6.655 16.375 6.98 ;
      RECT 15.985 6.29 16.275 6.52 ;
      RECT 15.58 2.395 15.685 2.965 ;
      RECT 15.58 2.73 15.905 2.96 ;
      RECT 15.58 2.76 16.075 2.93 ;
      RECT 15.58 2.395 15.77 2.96 ;
      RECT 14.995 2.36 15.285 2.59 ;
      RECT 14.995 2.395 15.77 2.565 ;
      RECT 15.055 0.88 15.225 2.59 ;
      RECT 14.995 0.88 15.285 1.11 ;
      RECT 14.995 7.77 15.285 8 ;
      RECT 15.055 6.29 15.225 8 ;
      RECT 14.995 6.29 15.285 6.52 ;
      RECT 14.995 6.325 15.85 6.485 ;
      RECT 15.68 5.92 15.85 6.485 ;
      RECT 14.995 6.32 15.39 6.485 ;
      RECT 15.615 5.92 15.905 6.15 ;
      RECT 15.615 5.95 16.075 6.12 ;
      RECT 14.625 2.73 14.915 2.96 ;
      RECT 14.625 2.76 15.085 2.93 ;
      RECT 14.69 1.655 14.855 2.96 ;
      RECT 13.205 1.625 13.495 1.855 ;
      RECT 13.205 1.655 14.855 1.825 ;
      RECT 13.265 0.885 13.435 1.855 ;
      RECT 13.205 0.885 13.495 1.115 ;
      RECT 13.205 7.765 13.495 7.995 ;
      RECT 13.265 7.025 13.435 7.995 ;
      RECT 13.265 7.12 14.855 7.29 ;
      RECT 14.685 5.92 14.855 7.29 ;
      RECT 13.205 7.025 13.495 7.255 ;
      RECT 14.625 5.92 14.915 6.15 ;
      RECT 14.625 5.95 15.085 6.12 ;
      RECT 11.19 1.995 11.515 2.32 ;
      RECT 13.635 1.965 13.985 2.315 ;
      RECT 11.19 2.025 13.985 2.195 ;
      RECT 13.66 6.655 13.985 6.98 ;
      RECT 13.635 6.655 13.985 6.885 ;
      RECT 13.465 6.685 13.985 6.855 ;
      RECT 12.86 2.365 13.18 2.685 ;
      RECT 12.83 2.365 13.18 2.595 ;
      RECT 12.545 2.395 13.18 2.565 ;
      RECT 12.86 6.28 13.18 6.605 ;
      RECT 12.83 6.285 13.18 6.515 ;
      RECT 12.66 6.315 13.18 6.485 ;
      RECT 10.19 2.77 10.51 3.03 ;
      RECT 9.915 2.83 10.51 2.97 ;
      RECT 7.81 3.11 8.13 3.37 ;
      RECT 9.785 3.125 10.075 3.355 ;
      RECT 7.81 3.17 10.075 3.31 ;
      RECT 9.17 5.83 9.49 6.09 ;
      RECT 9.17 5.89 9.765 6.03 ;
      RECT 8.49 2.77 8.81 3.03 ;
      RECT 3.75 2.785 4.04 3.015 ;
      RECT 3.75 2.83 8.81 2.97 ;
      RECT 8.58 2.49 8.72 3.03 ;
      RECT 8.58 2.49 9.06 2.63 ;
      RECT 8.92 2.105 9.06 2.63 ;
      RECT 8.845 2.105 9.135 2.335 ;
      RECT 8.49 3.79 8.81 4.05 ;
      RECT 7.825 3.805 8.115 4.035 ;
      RECT 5.615 3.805 5.905 4.035 ;
      RECT 5.615 3.85 8.81 3.99 ;
      RECT 6.79 5.83 7.11 6.09 ;
      RECT 8.505 5.845 8.795 6.075 ;
      RECT 6.125 5.845 6.415 6.075 ;
      RECT 6.125 5.89 7.11 6.03 ;
      RECT 8.58 5.55 8.72 6.075 ;
      RECT 6.88 5.55 7.02 6.09 ;
      RECT 6.88 5.55 8.72 5.69 ;
      RECT 5.785 2.445 6.075 2.675 ;
      RECT 5.86 2.15 6 2.675 ;
      RECT 8.15 2.09 8.47 2.35 ;
      RECT 8.05 2.105 8.47 2.335 ;
      RECT 5.86 2.15 8.47 2.29 ;
      RECT 7.13 2.43 7.45 2.69 ;
      RECT 7.13 2.49 7.725 2.63 ;
      RECT 7.13 4.81 7.45 5.07 ;
      RECT 4.425 4.825 4.715 5.055 ;
      RECT 4.425 4.87 7.45 5.01 ;
      RECT 6.455 2.39 6.785 2.72 ;
      RECT 6.45 2.425 6.785 2.685 ;
      RECT 6.8 2.445 6.915 2.675 ;
      RECT 6.45 2.44 6.8 2.67 ;
      RECT 6.45 2.49 6.93 2.63 ;
      RECT 6.335 2.49 6.345 2.63 ;
      RECT 6.345 2.485 6.915 2.625 ;
      RECT 2.44 6.63 2.78 6.91 ;
      RECT 2.41 6.655 2.78 6.885 ;
      RECT 2.24 6.685 2.78 6.855 ;
      RECT 1.98 7.765 2.27 7.995 ;
      RECT 2.04 6.995 2.21 7.995 ;
      RECT 1.94 6.995 2.31 7.365 ;
      RECT -1.25 7.765 -0.96 7.995 ;
      RECT -1.19 7.025 -1.02 7.995 ;
      RECT -1.27 7.025 -0.93 7.305 ;
      RECT -1.655 6.285 -1.315 6.565 ;
      RECT -1.795 6.315 -1.315 6.485 ;
      RECT 76.2 4.81 76.845 5.07 ;
      RECT 74.145 5.83 74.465 6.09 ;
      RECT 59.62 4.81 60.265 5.07 ;
      RECT 57.565 5.83 57.885 6.09 ;
      RECT 43.035 4.81 43.68 5.07 ;
      RECT 40.98 5.83 41.3 6.09 ;
      RECT 26.45 4.81 27.095 5.07 ;
      RECT 24.395 5.83 24.715 6.09 ;
      RECT 9.865 4.81 10.51 5.07 ;
      RECT 7.81 5.83 8.13 6.09 ;
    LAYER mcon ;
      RECT 82.38 6.32 82.55 6.49 ;
      RECT 82.385 6.315 82.555 6.485 ;
      RECT 65.8 6.32 65.97 6.49 ;
      RECT 65.805 6.315 65.975 6.485 ;
      RECT 49.215 6.32 49.385 6.49 ;
      RECT 49.22 6.315 49.39 6.485 ;
      RECT 32.63 6.32 32.8 6.49 ;
      RECT 32.635 6.315 32.805 6.485 ;
      RECT 16.045 6.32 16.215 6.49 ;
      RECT 16.05 6.315 16.22 6.485 ;
      RECT 82.38 7.8 82.55 7.97 ;
      RECT 82.01 2.76 82.18 2.93 ;
      RECT 82.01 5.95 82.18 6.12 ;
      RECT 81.39 0.91 81.56 1.08 ;
      RECT 81.39 2.39 81.56 2.56 ;
      RECT 81.39 6.32 81.56 6.49 ;
      RECT 81.39 7.8 81.56 7.97 ;
      RECT 81.02 2.76 81.19 2.93 ;
      RECT 81.02 5.95 81.19 6.12 ;
      RECT 80.03 2.025 80.2 2.195 ;
      RECT 80.03 6.685 80.2 6.855 ;
      RECT 79.6 0.915 79.77 1.085 ;
      RECT 79.6 1.655 79.77 1.825 ;
      RECT 79.6 7.055 79.77 7.225 ;
      RECT 79.6 7.795 79.77 7.965 ;
      RECT 79.225 2.395 79.395 2.565 ;
      RECT 79.225 6.315 79.395 6.485 ;
      RECT 76.6 2.815 76.77 2.985 ;
      RECT 76.26 4.855 76.43 5.025 ;
      RECT 76.18 3.155 76.35 3.325 ;
      RECT 75.58 5.875 75.75 6.045 ;
      RECT 75.24 2.135 75.41 2.305 ;
      RECT 74.9 5.875 75.07 6.045 ;
      RECT 74.445 2.135 74.615 2.305 ;
      RECT 74.22 3.835 74.39 4.005 ;
      RECT 74.22 5.875 74.39 6.045 ;
      RECT 73.54 2.475 73.71 2.645 ;
      RECT 72.52 5.875 72.69 6.045 ;
      RECT 72.18 2.475 72.35 2.645 ;
      RECT 72.01 3.835 72.18 4.005 ;
      RECT 70.82 4.855 70.99 5.025 ;
      RECT 70.145 2.815 70.315 2.985 ;
      RECT 68.805 6.685 68.975 6.855 ;
      RECT 68.375 7.055 68.545 7.225 ;
      RECT 68.375 7.795 68.545 7.965 ;
      RECT 65.8 7.8 65.97 7.97 ;
      RECT 65.43 2.76 65.6 2.93 ;
      RECT 65.43 5.95 65.6 6.12 ;
      RECT 64.81 0.91 64.98 1.08 ;
      RECT 64.81 2.39 64.98 2.56 ;
      RECT 64.81 6.32 64.98 6.49 ;
      RECT 64.81 7.8 64.98 7.97 ;
      RECT 64.44 2.76 64.61 2.93 ;
      RECT 64.44 5.95 64.61 6.12 ;
      RECT 63.45 2.025 63.62 2.195 ;
      RECT 63.45 6.685 63.62 6.855 ;
      RECT 63.02 0.915 63.19 1.085 ;
      RECT 63.02 1.655 63.19 1.825 ;
      RECT 63.02 7.055 63.19 7.225 ;
      RECT 63.02 7.795 63.19 7.965 ;
      RECT 62.645 2.395 62.815 2.565 ;
      RECT 62.645 6.315 62.815 6.485 ;
      RECT 60.02 2.815 60.19 2.985 ;
      RECT 59.68 4.855 59.85 5.025 ;
      RECT 59.6 3.155 59.77 3.325 ;
      RECT 59 5.875 59.17 6.045 ;
      RECT 58.66 2.135 58.83 2.305 ;
      RECT 58.32 5.875 58.49 6.045 ;
      RECT 57.865 2.135 58.035 2.305 ;
      RECT 57.64 3.835 57.81 4.005 ;
      RECT 57.64 5.875 57.81 6.045 ;
      RECT 56.96 2.475 57.13 2.645 ;
      RECT 55.94 5.875 56.11 6.045 ;
      RECT 55.6 2.475 55.77 2.645 ;
      RECT 55.43 3.835 55.6 4.005 ;
      RECT 54.24 4.855 54.41 5.025 ;
      RECT 53.565 2.815 53.735 2.985 ;
      RECT 52.225 6.685 52.395 6.855 ;
      RECT 51.795 7.055 51.965 7.225 ;
      RECT 51.795 7.795 51.965 7.965 ;
      RECT 49.215 7.8 49.385 7.97 ;
      RECT 48.845 2.76 49.015 2.93 ;
      RECT 48.845 5.95 49.015 6.12 ;
      RECT 48.225 0.91 48.395 1.08 ;
      RECT 48.225 2.39 48.395 2.56 ;
      RECT 48.225 6.32 48.395 6.49 ;
      RECT 48.225 7.8 48.395 7.97 ;
      RECT 47.855 2.76 48.025 2.93 ;
      RECT 47.855 5.95 48.025 6.12 ;
      RECT 46.865 2.025 47.035 2.195 ;
      RECT 46.865 6.685 47.035 6.855 ;
      RECT 46.435 0.915 46.605 1.085 ;
      RECT 46.435 1.655 46.605 1.825 ;
      RECT 46.435 7.055 46.605 7.225 ;
      RECT 46.435 7.795 46.605 7.965 ;
      RECT 46.06 2.395 46.23 2.565 ;
      RECT 46.06 6.315 46.23 6.485 ;
      RECT 43.435 2.815 43.605 2.985 ;
      RECT 43.095 4.855 43.265 5.025 ;
      RECT 43.015 3.155 43.185 3.325 ;
      RECT 42.415 5.875 42.585 6.045 ;
      RECT 42.075 2.135 42.245 2.305 ;
      RECT 41.735 5.875 41.905 6.045 ;
      RECT 41.28 2.135 41.45 2.305 ;
      RECT 41.055 3.835 41.225 4.005 ;
      RECT 41.055 5.875 41.225 6.045 ;
      RECT 40.375 2.475 40.545 2.645 ;
      RECT 39.355 5.875 39.525 6.045 ;
      RECT 39.015 2.475 39.185 2.645 ;
      RECT 38.845 3.835 39.015 4.005 ;
      RECT 37.655 4.855 37.825 5.025 ;
      RECT 36.98 2.815 37.15 2.985 ;
      RECT 35.64 6.685 35.81 6.855 ;
      RECT 35.21 7.055 35.38 7.225 ;
      RECT 35.21 7.795 35.38 7.965 ;
      RECT 32.63 7.8 32.8 7.97 ;
      RECT 32.26 2.76 32.43 2.93 ;
      RECT 32.26 5.95 32.43 6.12 ;
      RECT 31.64 0.91 31.81 1.08 ;
      RECT 31.64 2.39 31.81 2.56 ;
      RECT 31.64 6.32 31.81 6.49 ;
      RECT 31.64 7.8 31.81 7.97 ;
      RECT 31.27 2.76 31.44 2.93 ;
      RECT 31.27 5.95 31.44 6.12 ;
      RECT 30.28 2.025 30.45 2.195 ;
      RECT 30.28 6.685 30.45 6.855 ;
      RECT 29.85 0.915 30.02 1.085 ;
      RECT 29.85 1.655 30.02 1.825 ;
      RECT 29.85 7.055 30.02 7.225 ;
      RECT 29.85 7.795 30.02 7.965 ;
      RECT 29.475 2.395 29.645 2.565 ;
      RECT 29.475 6.315 29.645 6.485 ;
      RECT 26.85 2.815 27.02 2.985 ;
      RECT 26.51 4.855 26.68 5.025 ;
      RECT 26.43 3.155 26.6 3.325 ;
      RECT 25.83 5.875 26 6.045 ;
      RECT 25.49 2.135 25.66 2.305 ;
      RECT 25.15 5.875 25.32 6.045 ;
      RECT 24.695 2.135 24.865 2.305 ;
      RECT 24.47 3.835 24.64 4.005 ;
      RECT 24.47 5.875 24.64 6.045 ;
      RECT 23.79 2.475 23.96 2.645 ;
      RECT 22.77 5.875 22.94 6.045 ;
      RECT 22.43 2.475 22.6 2.645 ;
      RECT 22.26 3.835 22.43 4.005 ;
      RECT 21.07 4.855 21.24 5.025 ;
      RECT 20.395 2.815 20.565 2.985 ;
      RECT 19.055 6.685 19.225 6.855 ;
      RECT 18.625 7.055 18.795 7.225 ;
      RECT 18.625 7.795 18.795 7.965 ;
      RECT 16.045 7.8 16.215 7.97 ;
      RECT 15.675 2.76 15.845 2.93 ;
      RECT 15.675 5.95 15.845 6.12 ;
      RECT 15.055 0.91 15.225 1.08 ;
      RECT 15.055 2.39 15.225 2.56 ;
      RECT 15.055 6.32 15.225 6.49 ;
      RECT 15.055 7.8 15.225 7.97 ;
      RECT 14.685 2.76 14.855 2.93 ;
      RECT 14.685 5.95 14.855 6.12 ;
      RECT 13.695 2.025 13.865 2.195 ;
      RECT 13.695 6.685 13.865 6.855 ;
      RECT 13.265 0.915 13.435 1.085 ;
      RECT 13.265 1.655 13.435 1.825 ;
      RECT 13.265 7.055 13.435 7.225 ;
      RECT 13.265 7.795 13.435 7.965 ;
      RECT 12.89 2.395 13.06 2.565 ;
      RECT 12.89 6.315 13.06 6.485 ;
      RECT 10.265 2.815 10.435 2.985 ;
      RECT 9.925 4.855 10.095 5.025 ;
      RECT 9.845 3.155 10.015 3.325 ;
      RECT 9.245 5.875 9.415 6.045 ;
      RECT 8.905 2.135 9.075 2.305 ;
      RECT 8.565 5.875 8.735 6.045 ;
      RECT 8.11 2.135 8.28 2.305 ;
      RECT 7.885 3.835 8.055 4.005 ;
      RECT 7.885 5.875 8.055 6.045 ;
      RECT 7.205 2.475 7.375 2.645 ;
      RECT 6.185 5.875 6.355 6.045 ;
      RECT 5.845 2.475 6.015 2.645 ;
      RECT 5.675 3.835 5.845 4.005 ;
      RECT 4.485 4.855 4.655 5.025 ;
      RECT 3.81 2.815 3.98 2.985 ;
      RECT 2.47 6.685 2.64 6.855 ;
      RECT 2.04 7.055 2.21 7.225 ;
      RECT 2.04 7.795 2.21 7.965 ;
      RECT -1.19 7.055 -1.02 7.225 ;
      RECT -1.19 7.795 -1.02 7.965 ;
      RECT -1.565 6.315 -1.395 6.485 ;
    LAYER li1 ;
      RECT 82.38 5.02 82.55 6.49 ;
      RECT 82.38 6.315 82.555 6.485 ;
      RECT 82.01 1.74 82.18 2.93 ;
      RECT 82.01 1.74 82.48 1.91 ;
      RECT 82.01 6.97 82.48 7.14 ;
      RECT 82.01 5.95 82.18 7.14 ;
      RECT 81.02 1.74 81.19 2.93 ;
      RECT 81.02 1.74 81.49 1.91 ;
      RECT 81.02 6.97 81.49 7.14 ;
      RECT 81.02 5.95 81.19 7.14 ;
      RECT 79.17 2.635 79.34 3.865 ;
      RECT 79.225 0.855 79.395 2.805 ;
      RECT 79.17 0.575 79.34 1.025 ;
      RECT 79.17 7.855 79.34 8.305 ;
      RECT 79.225 6.075 79.395 8.025 ;
      RECT 79.17 5.015 79.34 6.245 ;
      RECT 78.65 0.575 78.82 3.865 ;
      RECT 78.65 2.075 79.055 2.405 ;
      RECT 78.65 1.235 79.055 1.565 ;
      RECT 78.65 5.015 78.82 8.305 ;
      RECT 78.65 7.315 79.055 7.645 ;
      RECT 78.65 6.475 79.055 6.805 ;
      RECT 73.91 6.645 75.215 6.895 ;
      RECT 73.91 6.325 74.09 6.895 ;
      RECT 73.36 6.325 74.09 6.495 ;
      RECT 73.36 5.485 73.53 6.495 ;
      RECT 74.195 5.525 75.94 5.705 ;
      RECT 75.61 4.685 75.94 5.705 ;
      RECT 73.36 5.485 74.42 5.655 ;
      RECT 75.61 4.855 76.43 5.025 ;
      RECT 74.77 4.685 75.1 4.895 ;
      RECT 74.77 4.685 75.94 4.855 ;
      RECT 75.67 3.205 76 4.16 ;
      RECT 75.67 3.205 76.35 3.375 ;
      RECT 76.18 1.965 76.35 3.375 ;
      RECT 76.09 1.965 76.42 2.605 ;
      RECT 75.215 3.475 75.49 4.175 ;
      RECT 75.32 1.965 75.49 4.175 ;
      RECT 75.66 2.785 76.01 3.035 ;
      RECT 75.32 2.815 76.01 2.985 ;
      RECT 75.23 1.965 75.49 2.445 ;
      RECT 74.56 5.115 75.44 5.355 ;
      RECT 75.21 5.025 75.44 5.355 ;
      RECT 73.91 5.115 75.44 5.315 ;
      RECT 74.825 5.065 75.44 5.355 ;
      RECT 73.91 4.985 74.08 5.315 ;
      RECT 74.795 5.875 75.045 6.475 ;
      RECT 74.795 5.875 75.27 6.075 ;
      RECT 74.29 3.095 75.045 3.595 ;
      RECT 73.36 2.9 73.62 3.52 ;
      RECT 74.275 3.04 74.29 3.345 ;
      RECT 74.26 3.025 74.28 3.31 ;
      RECT 74.92 2.7 75.15 3.3 ;
      RECT 74.235 2.97 74.255 3.285 ;
      RECT 74.215 3.095 75.15 3.27 ;
      RECT 74.19 3.095 75.15 3.26 ;
      RECT 74.12 3.095 75.15 3.25 ;
      RECT 74.1 3.095 75.15 3.22 ;
      RECT 74.08 2.005 74.25 3.19 ;
      RECT 74.05 3.095 75.15 3.16 ;
      RECT 74.015 3.095 75.15 3.135 ;
      RECT 73.985 3.09 74.375 3.1 ;
      RECT 73.985 3.08 74.35 3.1 ;
      RECT 73.985 3.075 74.335 3.1 ;
      RECT 73.985 3.065 74.32 3.1 ;
      RECT 73.36 2.9 74.25 3.07 ;
      RECT 73.36 3.055 74.31 3.07 ;
      RECT 73.36 3.05 74.3 3.07 ;
      RECT 74.255 2.995 74.265 3.3 ;
      RECT 73.36 3.03 74.285 3.07 ;
      RECT 73.36 3.01 74.27 3.07 ;
      RECT 73.36 2.005 74.25 2.175 ;
      RECT 74.42 2.5 74.75 2.925 ;
      RECT 74.42 2.015 74.64 2.925 ;
      RECT 74.335 5.875 74.545 6.475 ;
      RECT 74.195 5.875 74.545 6.075 ;
      RECT 72.915 3.475 73.19 4.175 ;
      RECT 73.135 1.965 73.19 4.175 ;
      RECT 73.02 2.77 73.19 4.175 ;
      RECT 73.02 1.965 73.19 2.765 ;
      RECT 72.93 1.965 73.19 2.44 ;
      RECT 71.06 3.135 71.31 3.67 ;
      RECT 72.03 3.135 72.745 3.6 ;
      RECT 71.06 3.135 72.85 3.305 ;
      RECT 72.62 2.77 72.85 3.305 ;
      RECT 71.615 2.015 71.87 3.305 ;
      RECT 72.62 2.705 72.68 3.6 ;
      RECT 72.68 2.7 72.85 2.765 ;
      RECT 71.08 2.015 71.87 2.28 ;
      RECT 72.04 5.825 72.715 6.075 ;
      RECT 72.45 5.465 72.715 6.075 ;
      RECT 72.2 6.245 72.53 6.795 ;
      RECT 71.14 6.245 72.53 6.435 ;
      RECT 71.14 5.405 71.31 6.435 ;
      RECT 71.02 5.825 71.31 6.155 ;
      RECT 71.14 5.405 72.08 5.575 ;
      RECT 71.78 4.855 72.08 5.575 ;
      RECT 72.04 2.435 72.45 2.955 ;
      RECT 72.04 2.015 72.24 2.955 ;
      RECT 70.65 2.195 70.82 4.175 ;
      RECT 70.65 2.705 71.445 2.955 ;
      RECT 70.65 2.195 70.9 2.955 ;
      RECT 70.57 2.195 70.9 2.615 ;
      RECT 70.6 6.605 71.16 6.895 ;
      RECT 70.6 4.685 70.85 6.895 ;
      RECT 70.6 4.685 71.06 5.235 ;
      RECT 67.425 5.015 67.595 8.305 ;
      RECT 67.425 7.315 67.83 7.645 ;
      RECT 67.425 6.475 67.83 6.805 ;
      RECT 65.8 5.02 65.97 6.49 ;
      RECT 65.8 6.315 65.975 6.485 ;
      RECT 65.43 1.74 65.6 2.93 ;
      RECT 65.43 1.74 65.9 1.91 ;
      RECT 65.43 6.97 65.9 7.14 ;
      RECT 65.43 5.95 65.6 7.14 ;
      RECT 64.44 1.74 64.61 2.93 ;
      RECT 64.44 1.74 64.91 1.91 ;
      RECT 64.44 6.97 64.91 7.14 ;
      RECT 64.44 5.95 64.61 7.14 ;
      RECT 62.59 2.635 62.76 3.865 ;
      RECT 62.645 0.855 62.815 2.805 ;
      RECT 62.59 0.575 62.76 1.025 ;
      RECT 62.59 7.855 62.76 8.305 ;
      RECT 62.645 6.075 62.815 8.025 ;
      RECT 62.59 5.015 62.76 6.245 ;
      RECT 62.07 0.575 62.24 3.865 ;
      RECT 62.07 2.075 62.475 2.405 ;
      RECT 62.07 1.235 62.475 1.565 ;
      RECT 62.07 5.015 62.24 8.305 ;
      RECT 62.07 7.315 62.475 7.645 ;
      RECT 62.07 6.475 62.475 6.805 ;
      RECT 57.33 6.645 58.635 6.895 ;
      RECT 57.33 6.325 57.51 6.895 ;
      RECT 56.78 6.325 57.51 6.495 ;
      RECT 56.78 5.485 56.95 6.495 ;
      RECT 57.615 5.525 59.36 5.705 ;
      RECT 59.03 4.685 59.36 5.705 ;
      RECT 56.78 5.485 57.84 5.655 ;
      RECT 59.03 4.855 59.85 5.025 ;
      RECT 58.19 4.685 58.52 4.895 ;
      RECT 58.19 4.685 59.36 4.855 ;
      RECT 59.09 3.205 59.42 4.16 ;
      RECT 59.09 3.205 59.77 3.375 ;
      RECT 59.6 1.965 59.77 3.375 ;
      RECT 59.51 1.965 59.84 2.605 ;
      RECT 58.635 3.475 58.91 4.175 ;
      RECT 58.74 1.965 58.91 4.175 ;
      RECT 59.08 2.785 59.43 3.035 ;
      RECT 58.74 2.815 59.43 2.985 ;
      RECT 58.65 1.965 58.91 2.445 ;
      RECT 57.98 5.115 58.86 5.355 ;
      RECT 58.63 5.025 58.86 5.355 ;
      RECT 57.33 5.115 58.86 5.315 ;
      RECT 58.245 5.065 58.86 5.355 ;
      RECT 57.33 4.985 57.5 5.315 ;
      RECT 58.215 5.875 58.465 6.475 ;
      RECT 58.215 5.875 58.69 6.075 ;
      RECT 57.71 3.095 58.465 3.595 ;
      RECT 56.78 2.9 57.04 3.52 ;
      RECT 57.695 3.04 57.71 3.345 ;
      RECT 57.68 3.025 57.7 3.31 ;
      RECT 58.34 2.7 58.57 3.3 ;
      RECT 57.655 2.97 57.675 3.285 ;
      RECT 57.635 3.095 58.57 3.27 ;
      RECT 57.61 3.095 58.57 3.26 ;
      RECT 57.54 3.095 58.57 3.25 ;
      RECT 57.52 3.095 58.57 3.22 ;
      RECT 57.5 2.005 57.67 3.19 ;
      RECT 57.47 3.095 58.57 3.16 ;
      RECT 57.435 3.095 58.57 3.135 ;
      RECT 57.405 3.09 57.795 3.1 ;
      RECT 57.405 3.08 57.77 3.1 ;
      RECT 57.405 3.075 57.755 3.1 ;
      RECT 57.405 3.065 57.74 3.1 ;
      RECT 56.78 2.9 57.67 3.07 ;
      RECT 56.78 3.055 57.73 3.07 ;
      RECT 56.78 3.05 57.72 3.07 ;
      RECT 57.675 2.995 57.685 3.3 ;
      RECT 56.78 3.03 57.705 3.07 ;
      RECT 56.78 3.01 57.69 3.07 ;
      RECT 56.78 2.005 57.67 2.175 ;
      RECT 57.84 2.5 58.17 2.925 ;
      RECT 57.84 2.015 58.06 2.925 ;
      RECT 57.755 5.875 57.965 6.475 ;
      RECT 57.615 5.875 57.965 6.075 ;
      RECT 56.335 3.475 56.61 4.175 ;
      RECT 56.555 1.965 56.61 4.175 ;
      RECT 56.44 2.77 56.61 4.175 ;
      RECT 56.44 1.965 56.61 2.765 ;
      RECT 56.35 1.965 56.61 2.44 ;
      RECT 54.48 3.135 54.73 3.67 ;
      RECT 55.45 3.135 56.165 3.6 ;
      RECT 54.48 3.135 56.27 3.305 ;
      RECT 56.04 2.77 56.27 3.305 ;
      RECT 55.035 2.015 55.29 3.305 ;
      RECT 56.04 2.705 56.1 3.6 ;
      RECT 56.1 2.7 56.27 2.765 ;
      RECT 54.5 2.015 55.29 2.28 ;
      RECT 55.46 5.825 56.135 6.075 ;
      RECT 55.87 5.465 56.135 6.075 ;
      RECT 55.62 6.245 55.95 6.795 ;
      RECT 54.56 6.245 55.95 6.435 ;
      RECT 54.56 5.405 54.73 6.435 ;
      RECT 54.44 5.825 54.73 6.155 ;
      RECT 54.56 5.405 55.5 5.575 ;
      RECT 55.2 4.855 55.5 5.575 ;
      RECT 55.46 2.435 55.87 2.955 ;
      RECT 55.46 2.015 55.66 2.955 ;
      RECT 54.07 2.195 54.24 4.175 ;
      RECT 54.07 2.705 54.865 2.955 ;
      RECT 54.07 2.195 54.32 2.955 ;
      RECT 53.99 2.195 54.32 2.615 ;
      RECT 54.02 6.605 54.58 6.895 ;
      RECT 54.02 4.685 54.27 6.895 ;
      RECT 54.02 4.685 54.48 5.235 ;
      RECT 50.845 5.015 51.015 8.305 ;
      RECT 50.845 7.315 51.25 7.645 ;
      RECT 50.845 6.475 51.25 6.805 ;
      RECT 49.215 5.02 49.385 6.49 ;
      RECT 49.215 6.315 49.39 6.485 ;
      RECT 48.845 1.74 49.015 2.93 ;
      RECT 48.845 1.74 49.315 1.91 ;
      RECT 48.845 6.97 49.315 7.14 ;
      RECT 48.845 5.95 49.015 7.14 ;
      RECT 47.855 1.74 48.025 2.93 ;
      RECT 47.855 1.74 48.325 1.91 ;
      RECT 47.855 6.97 48.325 7.14 ;
      RECT 47.855 5.95 48.025 7.14 ;
      RECT 46.005 2.635 46.175 3.865 ;
      RECT 46.06 0.855 46.23 2.805 ;
      RECT 46.005 0.575 46.175 1.025 ;
      RECT 46.005 7.855 46.175 8.305 ;
      RECT 46.06 6.075 46.23 8.025 ;
      RECT 46.005 5.015 46.175 6.245 ;
      RECT 45.485 0.575 45.655 3.865 ;
      RECT 45.485 2.075 45.89 2.405 ;
      RECT 45.485 1.235 45.89 1.565 ;
      RECT 45.485 5.015 45.655 8.305 ;
      RECT 45.485 7.315 45.89 7.645 ;
      RECT 45.485 6.475 45.89 6.805 ;
      RECT 40.745 6.645 42.05 6.895 ;
      RECT 40.745 6.325 40.925 6.895 ;
      RECT 40.195 6.325 40.925 6.495 ;
      RECT 40.195 5.485 40.365 6.495 ;
      RECT 41.03 5.525 42.775 5.705 ;
      RECT 42.445 4.685 42.775 5.705 ;
      RECT 40.195 5.485 41.255 5.655 ;
      RECT 42.445 4.855 43.265 5.025 ;
      RECT 41.605 4.685 41.935 4.895 ;
      RECT 41.605 4.685 42.775 4.855 ;
      RECT 42.505 3.205 42.835 4.16 ;
      RECT 42.505 3.205 43.185 3.375 ;
      RECT 43.015 1.965 43.185 3.375 ;
      RECT 42.925 1.965 43.255 2.605 ;
      RECT 42.05 3.475 42.325 4.175 ;
      RECT 42.155 1.965 42.325 4.175 ;
      RECT 42.495 2.785 42.845 3.035 ;
      RECT 42.155 2.815 42.845 2.985 ;
      RECT 42.065 1.965 42.325 2.445 ;
      RECT 41.395 5.115 42.275 5.355 ;
      RECT 42.045 5.025 42.275 5.355 ;
      RECT 40.745 5.115 42.275 5.315 ;
      RECT 41.66 5.065 42.275 5.355 ;
      RECT 40.745 4.985 40.915 5.315 ;
      RECT 41.63 5.875 41.88 6.475 ;
      RECT 41.63 5.875 42.105 6.075 ;
      RECT 41.125 3.095 41.88 3.595 ;
      RECT 40.195 2.9 40.455 3.52 ;
      RECT 41.11 3.04 41.125 3.345 ;
      RECT 41.095 3.025 41.115 3.31 ;
      RECT 41.755 2.7 41.985 3.3 ;
      RECT 41.07 2.97 41.09 3.285 ;
      RECT 41.05 3.095 41.985 3.27 ;
      RECT 41.025 3.095 41.985 3.26 ;
      RECT 40.955 3.095 41.985 3.25 ;
      RECT 40.935 3.095 41.985 3.22 ;
      RECT 40.915 2.005 41.085 3.19 ;
      RECT 40.885 3.095 41.985 3.16 ;
      RECT 40.85 3.095 41.985 3.135 ;
      RECT 40.82 3.09 41.21 3.1 ;
      RECT 40.82 3.08 41.185 3.1 ;
      RECT 40.82 3.075 41.17 3.1 ;
      RECT 40.82 3.065 41.155 3.1 ;
      RECT 40.195 2.9 41.085 3.07 ;
      RECT 40.195 3.055 41.145 3.07 ;
      RECT 40.195 3.05 41.135 3.07 ;
      RECT 41.09 2.995 41.1 3.3 ;
      RECT 40.195 3.03 41.12 3.07 ;
      RECT 40.195 3.01 41.105 3.07 ;
      RECT 40.195 2.005 41.085 2.175 ;
      RECT 41.255 2.5 41.585 2.925 ;
      RECT 41.255 2.015 41.475 2.925 ;
      RECT 41.17 5.875 41.38 6.475 ;
      RECT 41.03 5.875 41.38 6.075 ;
      RECT 39.75 3.475 40.025 4.175 ;
      RECT 39.97 1.965 40.025 4.175 ;
      RECT 39.855 2.77 40.025 4.175 ;
      RECT 39.855 1.965 40.025 2.765 ;
      RECT 39.765 1.965 40.025 2.44 ;
      RECT 37.895 3.135 38.145 3.67 ;
      RECT 38.865 3.135 39.58 3.6 ;
      RECT 37.895 3.135 39.685 3.305 ;
      RECT 39.455 2.77 39.685 3.305 ;
      RECT 38.45 2.015 38.705 3.305 ;
      RECT 39.455 2.705 39.515 3.6 ;
      RECT 39.515 2.7 39.685 2.765 ;
      RECT 37.915 2.015 38.705 2.28 ;
      RECT 38.875 5.825 39.55 6.075 ;
      RECT 39.285 5.465 39.55 6.075 ;
      RECT 39.035 6.245 39.365 6.795 ;
      RECT 37.975 6.245 39.365 6.435 ;
      RECT 37.975 5.405 38.145 6.435 ;
      RECT 37.855 5.825 38.145 6.155 ;
      RECT 37.975 5.405 38.915 5.575 ;
      RECT 38.615 4.855 38.915 5.575 ;
      RECT 38.875 2.435 39.285 2.955 ;
      RECT 38.875 2.015 39.075 2.955 ;
      RECT 37.485 2.195 37.655 4.175 ;
      RECT 37.485 2.705 38.28 2.955 ;
      RECT 37.485 2.195 37.735 2.955 ;
      RECT 37.405 2.195 37.735 2.615 ;
      RECT 37.435 6.605 37.995 6.895 ;
      RECT 37.435 4.685 37.685 6.895 ;
      RECT 37.435 4.685 37.895 5.235 ;
      RECT 34.26 5.015 34.43 8.305 ;
      RECT 34.26 7.315 34.665 7.645 ;
      RECT 34.26 6.475 34.665 6.805 ;
      RECT 32.63 5.02 32.8 6.49 ;
      RECT 32.63 6.315 32.805 6.485 ;
      RECT 32.26 1.74 32.43 2.93 ;
      RECT 32.26 1.74 32.73 1.91 ;
      RECT 32.26 6.97 32.73 7.14 ;
      RECT 32.26 5.95 32.43 7.14 ;
      RECT 31.27 1.74 31.44 2.93 ;
      RECT 31.27 1.74 31.74 1.91 ;
      RECT 31.27 6.97 31.74 7.14 ;
      RECT 31.27 5.95 31.44 7.14 ;
      RECT 29.42 2.635 29.59 3.865 ;
      RECT 29.475 0.855 29.645 2.805 ;
      RECT 29.42 0.575 29.59 1.025 ;
      RECT 29.42 7.855 29.59 8.305 ;
      RECT 29.475 6.075 29.645 8.025 ;
      RECT 29.42 5.015 29.59 6.245 ;
      RECT 28.9 0.575 29.07 3.865 ;
      RECT 28.9 2.075 29.305 2.405 ;
      RECT 28.9 1.235 29.305 1.565 ;
      RECT 28.9 5.015 29.07 8.305 ;
      RECT 28.9 7.315 29.305 7.645 ;
      RECT 28.9 6.475 29.305 6.805 ;
      RECT 24.16 6.645 25.465 6.895 ;
      RECT 24.16 6.325 24.34 6.895 ;
      RECT 23.61 6.325 24.34 6.495 ;
      RECT 23.61 5.485 23.78 6.495 ;
      RECT 24.445 5.525 26.19 5.705 ;
      RECT 25.86 4.685 26.19 5.705 ;
      RECT 23.61 5.485 24.67 5.655 ;
      RECT 25.86 4.855 26.68 5.025 ;
      RECT 25.02 4.685 25.35 4.895 ;
      RECT 25.02 4.685 26.19 4.855 ;
      RECT 25.92 3.205 26.25 4.16 ;
      RECT 25.92 3.205 26.6 3.375 ;
      RECT 26.43 1.965 26.6 3.375 ;
      RECT 26.34 1.965 26.67 2.605 ;
      RECT 25.465 3.475 25.74 4.175 ;
      RECT 25.57 1.965 25.74 4.175 ;
      RECT 25.91 2.785 26.26 3.035 ;
      RECT 25.57 2.815 26.26 2.985 ;
      RECT 25.48 1.965 25.74 2.445 ;
      RECT 24.81 5.115 25.69 5.355 ;
      RECT 25.46 5.025 25.69 5.355 ;
      RECT 24.16 5.115 25.69 5.315 ;
      RECT 25.075 5.065 25.69 5.355 ;
      RECT 24.16 4.985 24.33 5.315 ;
      RECT 25.045 5.875 25.295 6.475 ;
      RECT 25.045 5.875 25.52 6.075 ;
      RECT 24.54 3.095 25.295 3.595 ;
      RECT 23.61 2.9 23.87 3.52 ;
      RECT 24.525 3.04 24.54 3.345 ;
      RECT 24.51 3.025 24.53 3.31 ;
      RECT 25.17 2.7 25.4 3.3 ;
      RECT 24.485 2.97 24.505 3.285 ;
      RECT 24.465 3.095 25.4 3.27 ;
      RECT 24.44 3.095 25.4 3.26 ;
      RECT 24.37 3.095 25.4 3.25 ;
      RECT 24.35 3.095 25.4 3.22 ;
      RECT 24.33 2.005 24.5 3.19 ;
      RECT 24.3 3.095 25.4 3.16 ;
      RECT 24.265 3.095 25.4 3.135 ;
      RECT 24.235 3.09 24.625 3.1 ;
      RECT 24.235 3.08 24.6 3.1 ;
      RECT 24.235 3.075 24.585 3.1 ;
      RECT 24.235 3.065 24.57 3.1 ;
      RECT 23.61 2.9 24.5 3.07 ;
      RECT 23.61 3.055 24.56 3.07 ;
      RECT 23.61 3.05 24.55 3.07 ;
      RECT 24.505 2.995 24.515 3.3 ;
      RECT 23.61 3.03 24.535 3.07 ;
      RECT 23.61 3.01 24.52 3.07 ;
      RECT 23.61 2.005 24.5 2.175 ;
      RECT 24.67 2.5 25 2.925 ;
      RECT 24.67 2.015 24.89 2.925 ;
      RECT 24.585 5.875 24.795 6.475 ;
      RECT 24.445 5.875 24.795 6.075 ;
      RECT 23.165 3.475 23.44 4.175 ;
      RECT 23.385 1.965 23.44 4.175 ;
      RECT 23.27 2.77 23.44 4.175 ;
      RECT 23.27 1.965 23.44 2.765 ;
      RECT 23.18 1.965 23.44 2.44 ;
      RECT 21.31 3.135 21.56 3.67 ;
      RECT 22.28 3.135 22.995 3.6 ;
      RECT 21.31 3.135 23.1 3.305 ;
      RECT 22.87 2.77 23.1 3.305 ;
      RECT 21.865 2.015 22.12 3.305 ;
      RECT 22.87 2.705 22.93 3.6 ;
      RECT 22.93 2.7 23.1 2.765 ;
      RECT 21.33 2.015 22.12 2.28 ;
      RECT 22.29 5.825 22.965 6.075 ;
      RECT 22.7 5.465 22.965 6.075 ;
      RECT 22.45 6.245 22.78 6.795 ;
      RECT 21.39 6.245 22.78 6.435 ;
      RECT 21.39 5.405 21.56 6.435 ;
      RECT 21.27 5.825 21.56 6.155 ;
      RECT 21.39 5.405 22.33 5.575 ;
      RECT 22.03 4.855 22.33 5.575 ;
      RECT 22.29 2.435 22.7 2.955 ;
      RECT 22.29 2.015 22.49 2.955 ;
      RECT 20.9 2.195 21.07 4.175 ;
      RECT 20.9 2.705 21.695 2.955 ;
      RECT 20.9 2.195 21.15 2.955 ;
      RECT 20.82 2.195 21.15 2.615 ;
      RECT 20.85 6.605 21.41 6.895 ;
      RECT 20.85 4.685 21.1 6.895 ;
      RECT 20.85 4.685 21.31 5.235 ;
      RECT 17.675 5.015 17.845 8.305 ;
      RECT 17.675 7.315 18.08 7.645 ;
      RECT 17.675 6.475 18.08 6.805 ;
      RECT 16.045 5.02 16.215 6.49 ;
      RECT 16.045 6.315 16.22 6.485 ;
      RECT 15.675 1.74 15.845 2.93 ;
      RECT 15.675 1.74 16.145 1.91 ;
      RECT 15.675 6.97 16.145 7.14 ;
      RECT 15.675 5.95 15.845 7.14 ;
      RECT 14.685 1.74 14.855 2.93 ;
      RECT 14.685 1.74 15.155 1.91 ;
      RECT 14.685 6.97 15.155 7.14 ;
      RECT 14.685 5.95 14.855 7.14 ;
      RECT 12.835 2.635 13.005 3.865 ;
      RECT 12.89 0.855 13.06 2.805 ;
      RECT 12.835 0.575 13.005 1.025 ;
      RECT 12.835 7.855 13.005 8.305 ;
      RECT 12.89 6.075 13.06 8.025 ;
      RECT 12.835 5.015 13.005 6.245 ;
      RECT 12.315 0.575 12.485 3.865 ;
      RECT 12.315 2.075 12.72 2.405 ;
      RECT 12.315 1.235 12.72 1.565 ;
      RECT 12.315 5.015 12.485 8.305 ;
      RECT 12.315 7.315 12.72 7.645 ;
      RECT 12.315 6.475 12.72 6.805 ;
      RECT 7.575 6.645 8.88 6.895 ;
      RECT 7.575 6.325 7.755 6.895 ;
      RECT 7.025 6.325 7.755 6.495 ;
      RECT 7.025 5.485 7.195 6.495 ;
      RECT 7.86 5.525 9.605 5.705 ;
      RECT 9.275 4.685 9.605 5.705 ;
      RECT 7.025 5.485 8.085 5.655 ;
      RECT 9.275 4.855 10.095 5.025 ;
      RECT 8.435 4.685 8.765 4.895 ;
      RECT 8.435 4.685 9.605 4.855 ;
      RECT 9.335 3.205 9.665 4.16 ;
      RECT 9.335 3.205 10.015 3.375 ;
      RECT 9.845 1.965 10.015 3.375 ;
      RECT 9.755 1.965 10.085 2.605 ;
      RECT 8.88 3.475 9.155 4.175 ;
      RECT 8.985 1.965 9.155 4.175 ;
      RECT 9.325 2.785 9.675 3.035 ;
      RECT 8.985 2.815 9.675 2.985 ;
      RECT 8.895 1.965 9.155 2.445 ;
      RECT 8.225 5.115 9.105 5.355 ;
      RECT 8.875 5.025 9.105 5.355 ;
      RECT 7.575 5.115 9.105 5.315 ;
      RECT 8.49 5.065 9.105 5.355 ;
      RECT 7.575 4.985 7.745 5.315 ;
      RECT 8.46 5.875 8.71 6.475 ;
      RECT 8.46 5.875 8.935 6.075 ;
      RECT 7.955 3.095 8.71 3.595 ;
      RECT 7.025 2.9 7.285 3.52 ;
      RECT 7.94 3.04 7.955 3.345 ;
      RECT 7.925 3.025 7.945 3.31 ;
      RECT 8.585 2.7 8.815 3.3 ;
      RECT 7.9 2.97 7.92 3.285 ;
      RECT 7.88 3.095 8.815 3.27 ;
      RECT 7.855 3.095 8.815 3.26 ;
      RECT 7.785 3.095 8.815 3.25 ;
      RECT 7.765 3.095 8.815 3.22 ;
      RECT 7.745 2.005 7.915 3.19 ;
      RECT 7.715 3.095 8.815 3.16 ;
      RECT 7.68 3.095 8.815 3.135 ;
      RECT 7.65 3.09 8.04 3.1 ;
      RECT 7.65 3.08 8.015 3.1 ;
      RECT 7.65 3.075 8 3.1 ;
      RECT 7.65 3.065 7.985 3.1 ;
      RECT 7.025 2.9 7.915 3.07 ;
      RECT 7.025 3.055 7.975 3.07 ;
      RECT 7.025 3.05 7.965 3.07 ;
      RECT 7.92 2.995 7.93 3.3 ;
      RECT 7.025 3.03 7.95 3.07 ;
      RECT 7.025 3.01 7.935 3.07 ;
      RECT 7.025 2.005 7.915 2.175 ;
      RECT 8.085 2.5 8.415 2.925 ;
      RECT 8.085 2.015 8.305 2.925 ;
      RECT 8 5.875 8.21 6.475 ;
      RECT 7.86 5.875 8.21 6.075 ;
      RECT 6.58 3.475 6.855 4.175 ;
      RECT 6.8 1.965 6.855 4.175 ;
      RECT 6.685 2.77 6.855 4.175 ;
      RECT 6.685 1.965 6.855 2.765 ;
      RECT 6.595 1.965 6.855 2.44 ;
      RECT 4.725 3.135 4.975 3.67 ;
      RECT 5.695 3.135 6.41 3.6 ;
      RECT 4.725 3.135 6.515 3.305 ;
      RECT 6.285 2.77 6.515 3.305 ;
      RECT 5.28 2.015 5.535 3.305 ;
      RECT 6.285 2.705 6.345 3.6 ;
      RECT 6.345 2.7 6.515 2.765 ;
      RECT 4.745 2.015 5.535 2.28 ;
      RECT 5.705 5.825 6.38 6.075 ;
      RECT 6.115 5.465 6.38 6.075 ;
      RECT 5.865 6.245 6.195 6.795 ;
      RECT 4.805 6.245 6.195 6.435 ;
      RECT 4.805 5.405 4.975 6.435 ;
      RECT 4.685 5.825 4.975 6.155 ;
      RECT 4.805 5.405 5.745 5.575 ;
      RECT 5.445 4.855 5.745 5.575 ;
      RECT 5.705 2.435 6.115 2.955 ;
      RECT 5.705 2.015 5.905 2.955 ;
      RECT 4.315 2.195 4.485 4.175 ;
      RECT 4.315 2.705 5.11 2.955 ;
      RECT 4.315 2.195 4.565 2.955 ;
      RECT 4.235 2.195 4.565 2.615 ;
      RECT 4.265 6.605 4.825 6.895 ;
      RECT 4.265 4.685 4.515 6.895 ;
      RECT 4.265 4.685 4.725 5.235 ;
      RECT 1.09 5.015 1.26 8.305 ;
      RECT 1.09 7.315 1.495 7.645 ;
      RECT 1.09 6.475 1.495 6.805 ;
      RECT -1.62 7.855 -1.45 8.305 ;
      RECT -1.565 6.075 -1.395 8.025 ;
      RECT -1.62 5.015 -1.45 6.245 ;
      RECT -2.14 5.015 -1.97 8.305 ;
      RECT -2.14 7.315 -1.735 7.645 ;
      RECT -2.14 6.475 -1.735 6.805 ;
      RECT 82.38 7.8 82.55 8.31 ;
      RECT 81.39 0.57 81.56 1.08 ;
      RECT 81.39 2.39 81.56 3.86 ;
      RECT 81.39 5.02 81.56 6.49 ;
      RECT 81.39 7.8 81.56 8.31 ;
      RECT 80.03 0.575 80.2 3.865 ;
      RECT 80.03 5.015 80.2 8.305 ;
      RECT 79.6 0.575 79.77 1.085 ;
      RECT 79.6 1.655 79.77 3.865 ;
      RECT 79.6 5.015 79.77 7.225 ;
      RECT 79.6 7.795 79.77 8.305 ;
      RECT 76.52 2.785 76.87 3.035 ;
      RECT 75.46 5.875 75.91 6.385 ;
      RECT 74.14 3.835 74.62 4.175 ;
      RECT 73.36 2.345 73.91 2.73 ;
      RECT 71.845 3.835 72.32 4.175 ;
      RECT 70.14 2.785 70.48 3.665 ;
      RECT 68.805 5.015 68.975 8.305 ;
      RECT 68.375 5.015 68.545 7.225 ;
      RECT 68.375 7.795 68.545 8.305 ;
      RECT 65.8 7.8 65.97 8.31 ;
      RECT 64.81 0.57 64.98 1.08 ;
      RECT 64.81 2.39 64.98 3.86 ;
      RECT 64.81 5.02 64.98 6.49 ;
      RECT 64.81 7.8 64.98 8.31 ;
      RECT 63.45 0.575 63.62 3.865 ;
      RECT 63.45 5.015 63.62 8.305 ;
      RECT 63.02 0.575 63.19 1.085 ;
      RECT 63.02 1.655 63.19 3.865 ;
      RECT 63.02 5.015 63.19 7.225 ;
      RECT 63.02 7.795 63.19 8.305 ;
      RECT 59.94 2.785 60.29 3.035 ;
      RECT 58.88 5.875 59.33 6.385 ;
      RECT 57.56 3.835 58.04 4.175 ;
      RECT 56.78 2.345 57.33 2.73 ;
      RECT 55.265 3.835 55.74 4.175 ;
      RECT 53.56 2.785 53.9 3.665 ;
      RECT 52.225 5.015 52.395 8.305 ;
      RECT 51.795 5.015 51.965 7.225 ;
      RECT 51.795 7.795 51.965 8.305 ;
      RECT 49.215 7.8 49.385 8.31 ;
      RECT 48.225 0.57 48.395 1.08 ;
      RECT 48.225 2.39 48.395 3.86 ;
      RECT 48.225 5.02 48.395 6.49 ;
      RECT 48.225 7.8 48.395 8.31 ;
      RECT 46.865 0.575 47.035 3.865 ;
      RECT 46.865 5.015 47.035 8.305 ;
      RECT 46.435 0.575 46.605 1.085 ;
      RECT 46.435 1.655 46.605 3.865 ;
      RECT 46.435 5.015 46.605 7.225 ;
      RECT 46.435 7.795 46.605 8.305 ;
      RECT 43.355 2.785 43.705 3.035 ;
      RECT 42.295 5.875 42.745 6.385 ;
      RECT 40.975 3.835 41.455 4.175 ;
      RECT 40.195 2.345 40.745 2.73 ;
      RECT 38.68 3.835 39.155 4.175 ;
      RECT 36.975 2.785 37.315 3.665 ;
      RECT 35.64 5.015 35.81 8.305 ;
      RECT 35.21 5.015 35.38 7.225 ;
      RECT 35.21 7.795 35.38 8.305 ;
      RECT 32.63 7.8 32.8 8.31 ;
      RECT 31.64 0.57 31.81 1.08 ;
      RECT 31.64 2.39 31.81 3.86 ;
      RECT 31.64 5.02 31.81 6.49 ;
      RECT 31.64 7.8 31.81 8.31 ;
      RECT 30.28 0.575 30.45 3.865 ;
      RECT 30.28 5.015 30.45 8.305 ;
      RECT 29.85 0.575 30.02 1.085 ;
      RECT 29.85 1.655 30.02 3.865 ;
      RECT 29.85 5.015 30.02 7.225 ;
      RECT 29.85 7.795 30.02 8.305 ;
      RECT 26.77 2.785 27.12 3.035 ;
      RECT 25.71 5.875 26.16 6.385 ;
      RECT 24.39 3.835 24.87 4.175 ;
      RECT 23.61 2.345 24.16 2.73 ;
      RECT 22.095 3.835 22.57 4.175 ;
      RECT 20.39 2.785 20.73 3.665 ;
      RECT 19.055 5.015 19.225 8.305 ;
      RECT 18.625 5.015 18.795 7.225 ;
      RECT 18.625 7.795 18.795 8.305 ;
      RECT 16.045 7.8 16.215 8.31 ;
      RECT 15.055 0.57 15.225 1.08 ;
      RECT 15.055 2.39 15.225 3.86 ;
      RECT 15.055 5.02 15.225 6.49 ;
      RECT 15.055 7.8 15.225 8.31 ;
      RECT 13.695 0.575 13.865 3.865 ;
      RECT 13.695 5.015 13.865 8.305 ;
      RECT 13.265 0.575 13.435 1.085 ;
      RECT 13.265 1.655 13.435 3.865 ;
      RECT 13.265 5.015 13.435 7.225 ;
      RECT 13.265 7.795 13.435 8.305 ;
      RECT 10.185 2.785 10.535 3.035 ;
      RECT 9.125 5.875 9.575 6.385 ;
      RECT 7.805 3.835 8.285 4.175 ;
      RECT 7.025 2.345 7.575 2.73 ;
      RECT 5.51 3.835 5.985 4.175 ;
      RECT 3.805 2.785 4.145 3.665 ;
      RECT 2.47 5.015 2.64 8.305 ;
      RECT 2.04 5.015 2.21 7.225 ;
      RECT 2.04 7.795 2.21 8.305 ;
      RECT -1.19 5.015 -1.02 7.225 ;
      RECT -1.19 7.795 -1.02 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2ca_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2ct_8_b0r1
  CLASS BLOCK ;
  ORIGIN 3.44 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ct_8_b0r1 ;
  SIZE 88.91 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 16.05 0.915 16.22 1.085 ;
        RECT 16.045 0.91 16.215 1.08 ;
        RECT 16.045 2.39 16.215 2.56 ;
      LAYER li1 ;
        RECT 16.05 0.915 16.22 1.085 ;
        RECT 16.045 0.57 16.215 1.08 ;
        RECT 16.045 2.39 16.215 3.86 ;
      LAYER met1 ;
        RECT 15.985 2.36 16.275 2.59 ;
        RECT 15.985 0.88 16.275 1.11 ;
        RECT 16.045 0.88 16.215 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 33.27 0.915 33.44 1.085 ;
        RECT 33.265 0.91 33.435 1.08 ;
        RECT 33.265 2.39 33.435 2.56 ;
      LAYER li1 ;
        RECT 33.27 0.915 33.44 1.085 ;
        RECT 33.265 0.57 33.435 1.08 ;
        RECT 33.265 2.39 33.435 3.86 ;
      LAYER met1 ;
        RECT 33.205 2.36 33.495 2.59 ;
        RECT 33.205 0.88 33.495 1.11 ;
        RECT 33.265 0.88 33.435 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 50.49 0.915 50.66 1.085 ;
        RECT 50.485 0.91 50.655 1.08 ;
        RECT 50.485 2.39 50.655 2.56 ;
      LAYER li1 ;
        RECT 50.49 0.915 50.66 1.085 ;
        RECT 50.485 0.57 50.655 1.08 ;
        RECT 50.485 2.39 50.655 3.86 ;
      LAYER met1 ;
        RECT 50.425 2.36 50.715 2.59 ;
        RECT 50.425 0.88 50.715 1.11 ;
        RECT 50.485 0.88 50.655 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 67.71 0.915 67.88 1.085 ;
        RECT 67.705 0.91 67.875 1.08 ;
        RECT 67.705 2.39 67.875 2.56 ;
      LAYER li1 ;
        RECT 67.71 0.915 67.88 1.085 ;
        RECT 67.705 0.57 67.875 1.08 ;
        RECT 67.705 2.39 67.875 3.86 ;
      LAYER met1 ;
        RECT 67.645 2.36 67.935 2.59 ;
        RECT 67.645 0.88 67.935 1.11 ;
        RECT 67.705 0.88 67.875 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 84.93 0.915 85.1 1.085 ;
        RECT 84.925 0.91 85.095 1.08 ;
        RECT 84.925 2.39 85.095 2.56 ;
      LAYER li1 ;
        RECT 84.93 0.915 85.1 1.085 ;
        RECT 84.925 0.57 85.095 1.08 ;
        RECT 84.925 2.39 85.095 3.86 ;
      LAYER met1 ;
        RECT 84.865 2.36 85.155 2.59 ;
        RECT 84.865 0.88 85.155 1.11 ;
        RECT 84.925 0.88 85.095 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 11.895 1.66 12.065 2.935 ;
        RECT 11.895 5.94 12.065 7.22 ;
        RECT 11.885 5.94 12.065 6.18 ;
        RECT 0.21 5.945 0.38 7.22 ;
      LAYER met2 ;
        RECT 11.815 5.855 12.14 6.18 ;
        RECT 11.815 3.495 12.14 3.82 ;
        RECT 2.515 7.55 12.065 7.72 ;
        RECT 11.895 5.855 12.065 7.72 ;
        RECT 11.885 3.495 12.055 6.18 ;
        RECT 2.46 5.86 2.74 6.2 ;
        RECT 2.515 5.86 2.685 7.72 ;
      LAYER met1 ;
        RECT 11.835 2.765 12.295 2.935 ;
        RECT 11.815 3.495 12.14 3.82 ;
        RECT 11.835 2.735 12.125 2.965 ;
        RECT 11.895 2.735 12.065 3.82 ;
        RECT 11.815 5.945 12.295 6.115 ;
        RECT 11.815 5.855 12.14 6.18 ;
        RECT 2.43 5.89 2.77 6.17 ;
        RECT 0.15 5.945 2.77 6.115 ;
        RECT 0.15 5.915 0.44 6.145 ;
      LAYER via1 ;
        RECT 2.525 5.955 2.675 6.105 ;
        RECT 11.905 5.94 12.055 6.09 ;
        RECT 11.905 3.58 12.055 3.73 ;
      LAYER mcon ;
        RECT 0.21 5.945 0.38 6.115 ;
        RECT 11.895 5.945 12.065 6.115 ;
        RECT 11.895 2.765 12.065 2.935 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 29.115 1.66 29.285 2.935 ;
        RECT 29.115 5.94 29.285 7.22 ;
        RECT 29.105 5.94 29.285 6.18 ;
        RECT 17.43 5.945 17.6 7.22 ;
      LAYER met2 ;
        RECT 29.035 5.855 29.36 6.18 ;
        RECT 29.035 3.495 29.36 3.82 ;
        RECT 19.735 7.55 29.285 7.72 ;
        RECT 29.115 5.855 29.285 7.72 ;
        RECT 29.105 3.495 29.275 6.18 ;
        RECT 19.68 5.86 19.96 6.2 ;
        RECT 19.735 5.86 19.905 7.72 ;
      LAYER met1 ;
        RECT 29.055 2.765 29.515 2.935 ;
        RECT 29.035 3.495 29.36 3.82 ;
        RECT 29.055 2.735 29.345 2.965 ;
        RECT 29.115 2.735 29.285 3.82 ;
        RECT 29.035 5.945 29.515 6.115 ;
        RECT 29.035 5.855 29.36 6.18 ;
        RECT 19.65 5.89 19.99 6.17 ;
        RECT 17.37 5.945 19.99 6.115 ;
        RECT 17.37 5.915 17.66 6.145 ;
      LAYER via1 ;
        RECT 19.745 5.955 19.895 6.105 ;
        RECT 29.125 5.94 29.275 6.09 ;
        RECT 29.125 3.58 29.275 3.73 ;
      LAYER mcon ;
        RECT 17.43 5.945 17.6 6.115 ;
        RECT 29.115 5.945 29.285 6.115 ;
        RECT 29.115 2.765 29.285 2.935 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 46.335 1.66 46.505 2.935 ;
        RECT 46.335 5.94 46.505 7.22 ;
        RECT 46.325 5.94 46.505 6.18 ;
        RECT 34.65 5.945 34.82 7.22 ;
      LAYER met2 ;
        RECT 46.255 5.855 46.58 6.18 ;
        RECT 46.255 3.495 46.58 3.82 ;
        RECT 36.955 7.55 46.505 7.72 ;
        RECT 46.335 5.855 46.505 7.72 ;
        RECT 46.325 3.495 46.495 6.18 ;
        RECT 36.9 5.86 37.18 6.2 ;
        RECT 36.955 5.86 37.125 7.72 ;
      LAYER met1 ;
        RECT 46.275 2.765 46.735 2.935 ;
        RECT 46.255 3.495 46.58 3.82 ;
        RECT 46.275 2.735 46.565 2.965 ;
        RECT 46.335 2.735 46.505 3.82 ;
        RECT 46.255 5.945 46.735 6.115 ;
        RECT 46.255 5.855 46.58 6.18 ;
        RECT 36.87 5.89 37.21 6.17 ;
        RECT 34.59 5.945 37.21 6.115 ;
        RECT 34.59 5.915 34.88 6.145 ;
      LAYER via1 ;
        RECT 36.965 5.955 37.115 6.105 ;
        RECT 46.345 5.94 46.495 6.09 ;
        RECT 46.345 3.58 46.495 3.73 ;
      LAYER mcon ;
        RECT 34.65 5.945 34.82 6.115 ;
        RECT 46.335 5.945 46.505 6.115 ;
        RECT 46.335 2.765 46.505 2.935 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 63.555 1.66 63.725 2.935 ;
        RECT 63.555 5.94 63.725 7.22 ;
        RECT 63.545 5.94 63.725 6.18 ;
        RECT 51.87 5.945 52.04 7.22 ;
      LAYER met2 ;
        RECT 63.475 5.855 63.8 6.18 ;
        RECT 63.475 3.495 63.8 3.82 ;
        RECT 54.175 7.55 63.725 7.72 ;
        RECT 63.555 5.855 63.725 7.72 ;
        RECT 63.545 3.495 63.715 6.18 ;
        RECT 54.12 5.86 54.4 6.2 ;
        RECT 54.175 5.86 54.345 7.72 ;
      LAYER met1 ;
        RECT 63.495 2.765 63.955 2.935 ;
        RECT 63.475 3.495 63.8 3.82 ;
        RECT 63.495 2.735 63.785 2.965 ;
        RECT 63.555 2.735 63.725 3.82 ;
        RECT 63.475 5.945 63.955 6.115 ;
        RECT 63.475 5.855 63.8 6.18 ;
        RECT 54.09 5.89 54.43 6.17 ;
        RECT 51.81 5.945 54.43 6.115 ;
        RECT 51.81 5.915 52.1 6.145 ;
      LAYER via1 ;
        RECT 54.185 5.955 54.335 6.105 ;
        RECT 63.565 5.94 63.715 6.09 ;
        RECT 63.565 3.58 63.715 3.73 ;
      LAYER mcon ;
        RECT 51.87 5.945 52.04 6.115 ;
        RECT 63.555 5.945 63.725 6.115 ;
        RECT 63.555 2.765 63.725 2.935 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 80.775 1.66 80.945 2.935 ;
        RECT 80.775 5.94 80.945 7.22 ;
        RECT 80.765 5.94 80.945 6.18 ;
        RECT 69.09 5.945 69.26 7.22 ;
      LAYER met2 ;
        RECT 80.695 5.855 81.02 6.18 ;
        RECT 80.695 3.495 81.02 3.82 ;
        RECT 71.395 7.55 80.945 7.72 ;
        RECT 80.775 5.855 80.945 7.72 ;
        RECT 80.765 3.495 80.935 6.18 ;
        RECT 71.34 5.86 71.62 6.2 ;
        RECT 71.395 5.86 71.565 7.72 ;
      LAYER met1 ;
        RECT 80.715 2.765 81.175 2.935 ;
        RECT 80.695 3.495 81.02 3.82 ;
        RECT 80.715 2.735 81.005 2.965 ;
        RECT 80.775 2.735 80.945 3.82 ;
        RECT 80.695 5.945 81.175 6.115 ;
        RECT 80.695 5.855 81.02 6.18 ;
        RECT 71.31 5.89 71.65 6.17 ;
        RECT 69.03 5.945 71.65 6.115 ;
        RECT 69.03 5.915 69.32 6.145 ;
      LAYER via1 ;
        RECT 71.405 5.955 71.555 6.105 ;
        RECT 80.785 5.94 80.935 6.09 ;
        RECT 80.785 3.58 80.935 3.73 ;
      LAYER mcon ;
        RECT 69.09 5.945 69.26 6.115 ;
        RECT 80.775 5.945 80.945 6.115 ;
        RECT 80.775 2.765 80.945 2.935 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT -3.2 5.945 -3.03 7.22 ;
      LAYER met1 ;
        RECT -3.26 5.945 -2.8 6.115 ;
        RECT -3.26 5.915 -2.97 6.145 ;
      LAYER mcon ;
        RECT -3.2 5.945 -3.03 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 79.485 4.135 85.47 4.745 ;
        RECT 83.335 4.13 85.315 4.75 ;
        RECT 84.495 3.4 84.665 5.48 ;
        RECT 83.505 3.4 83.675 5.48 ;
        RECT 80.765 3.405 80.935 5.475 ;
        RECT -3.44 4.345 85.47 4.515 ;
        RECT 79.48 4.135 85.47 4.515 ;
        RECT 78.57 4.345 78.85 5.655 ;
        RECT 78.17 3.495 78.34 4.515 ;
        RECT 77.64 4.345 77.9 5.655 ;
        RECT 77.33 3.835 77.5 4.515 ;
        RECT 77.19 4.345 77.47 5.655 ;
        RECT 76.26 4.345 76.52 5.655 ;
        RECT 75.83 4.345 76.09 5.655 ;
        RECT 75.75 3.205 76.08 4.515 ;
        RECT 74.88 4.345 75.16 5.655 ;
        RECT 73.51 3.205 73.84 4.515 ;
        RECT 73.53 3.205 73.79 5.655 ;
        RECT 73.06 3.205 73.29 4.515 ;
        RECT 72.58 4.345 72.86 5.655 ;
        RECT 62.265 4.345 72.41 4.74 ;
        RECT 62.26 4.135 72.39 4.515 ;
        RECT 72.18 3.205 72.39 4.74 ;
        RECT 68.245 4.13 72.39 4.74 ;
        RECT 68.905 4.13 71.655 4.745 ;
        RECT 69.08 4.13 69.25 5.475 ;
        RECT 62.265 4.135 68.25 4.745 ;
        RECT 66.115 4.13 68.095 4.75 ;
        RECT 67.275 3.4 67.445 5.48 ;
        RECT 66.285 3.4 66.455 5.48 ;
        RECT 63.545 3.405 63.715 5.475 ;
        RECT 61.35 4.345 61.63 5.655 ;
        RECT 60.95 3.495 61.12 4.515 ;
        RECT 60.42 4.345 60.68 5.655 ;
        RECT 60.11 3.835 60.28 4.515 ;
        RECT 59.97 4.345 60.25 5.655 ;
        RECT 59.04 4.345 59.3 5.655 ;
        RECT 58.61 4.345 58.87 5.655 ;
        RECT 58.53 3.205 58.86 4.515 ;
        RECT 57.66 4.345 57.94 5.655 ;
        RECT 56.29 3.205 56.62 4.515 ;
        RECT 56.31 3.205 56.57 5.655 ;
        RECT 55.84 3.205 56.07 4.515 ;
        RECT 55.36 4.345 55.64 5.655 ;
        RECT 45.045 4.345 55.19 4.74 ;
        RECT 45.04 4.135 55.17 4.515 ;
        RECT 54.96 3.205 55.17 4.74 ;
        RECT 51.025 4.13 55.17 4.74 ;
        RECT 51.685 4.13 54.435 4.745 ;
        RECT 51.86 4.13 52.03 5.475 ;
        RECT 45.045 4.135 51.03 4.745 ;
        RECT 48.895 4.13 50.875 4.75 ;
        RECT 50.055 3.4 50.225 5.48 ;
        RECT 49.065 3.4 49.235 5.48 ;
        RECT 46.325 3.405 46.495 5.475 ;
        RECT 44.13 4.345 44.41 5.655 ;
        RECT 43.73 3.495 43.9 4.515 ;
        RECT 43.2 4.345 43.46 5.655 ;
        RECT 42.89 3.835 43.06 4.515 ;
        RECT 42.75 4.345 43.03 5.655 ;
        RECT 41.82 4.345 42.08 5.655 ;
        RECT 41.39 4.345 41.65 5.655 ;
        RECT 41.31 3.205 41.64 4.515 ;
        RECT 40.44 4.345 40.72 5.655 ;
        RECT 39.07 3.205 39.4 4.515 ;
        RECT 39.09 3.205 39.35 5.655 ;
        RECT 38.62 3.205 38.85 4.515 ;
        RECT 38.14 4.345 38.42 5.655 ;
        RECT 27.825 4.345 37.97 4.74 ;
        RECT 27.82 4.135 37.95 4.515 ;
        RECT 37.74 3.205 37.95 4.74 ;
        RECT 33.805 4.13 37.95 4.74 ;
        RECT 34.465 4.13 37.215 4.745 ;
        RECT 34.64 4.13 34.81 5.475 ;
        RECT 27.825 4.135 33.81 4.745 ;
        RECT 31.675 4.13 33.655 4.75 ;
        RECT 32.835 3.4 33.005 5.48 ;
        RECT 31.845 3.4 32.015 5.48 ;
        RECT 29.105 3.405 29.275 5.475 ;
        RECT 26.91 4.345 27.19 5.655 ;
        RECT 26.51 3.495 26.68 4.515 ;
        RECT 25.98 4.345 26.24 5.655 ;
        RECT 25.67 3.835 25.84 4.515 ;
        RECT 25.53 4.345 25.81 5.655 ;
        RECT 24.6 4.345 24.86 5.655 ;
        RECT 24.17 4.345 24.43 5.655 ;
        RECT 24.09 3.205 24.42 4.515 ;
        RECT 23.22 4.345 23.5 5.655 ;
        RECT 21.85 3.205 22.18 4.515 ;
        RECT 21.87 3.205 22.13 5.655 ;
        RECT 21.4 3.205 21.63 4.515 ;
        RECT 20.92 4.345 21.2 5.655 ;
        RECT 10.605 4.345 20.75 4.74 ;
        RECT 10.6 4.135 20.73 4.515 ;
        RECT 20.52 3.205 20.73 4.74 ;
        RECT 16.585 4.13 20.73 4.74 ;
        RECT 17.245 4.13 19.995 4.745 ;
        RECT 17.42 4.13 17.59 5.475 ;
        RECT 10.605 4.135 16.59 4.745 ;
        RECT 14.455 4.13 16.435 4.75 ;
        RECT 15.615 3.4 15.785 5.48 ;
        RECT 14.625 3.4 14.795 5.48 ;
        RECT 11.885 3.405 12.055 5.475 ;
        RECT 9.69 4.345 9.97 5.655 ;
        RECT 9.29 3.495 9.46 4.515 ;
        RECT 8.76 4.345 9.02 5.655 ;
        RECT 8.45 3.835 8.62 4.515 ;
        RECT 8.31 4.345 8.59 5.655 ;
        RECT 7.38 4.345 7.64 5.655 ;
        RECT 6.95 4.345 7.21 5.655 ;
        RECT 6.87 3.205 7.2 4.515 ;
        RECT 6 4.345 6.28 5.655 ;
        RECT 4.63 3.205 4.96 4.515 ;
        RECT 4.65 3.205 4.91 5.655 ;
        RECT 4.18 3.205 4.41 4.515 ;
        RECT 3.7 4.345 3.98 5.655 ;
        RECT -3.44 4.345 3.53 4.74 ;
        RECT -3.44 4.13 3.51 4.74 ;
        RECT 3.3 3.205 3.51 4.74 ;
        RECT 0.025 4.13 2.775 4.745 ;
        RECT 0.2 4.13 0.37 5.475 ;
        RECT -3.385 4.13 -0.635 4.745 ;
        RECT -1.4 4.13 -1.23 8.305 ;
        RECT -3.21 4.13 -3.04 5.475 ;
      LAYER met1 ;
        RECT 79.485 4.135 85.47 4.745 ;
        RECT 83.335 4.13 85.315 4.75 ;
        RECT -3.44 4.19 85.47 4.67 ;
        RECT 79.48 4.135 85.47 4.67 ;
        RECT 62.265 4.19 72.41 4.74 ;
        RECT 62.26 4.135 72.39 4.67 ;
        RECT 68.245 4.13 72.39 4.74 ;
        RECT 68.905 4.13 71.655 4.745 ;
        RECT 62.265 4.135 68.25 4.745 ;
        RECT 66.115 4.13 68.095 4.75 ;
        RECT 45.045 4.19 55.19 4.74 ;
        RECT 45.04 4.135 55.17 4.67 ;
        RECT 51.025 4.13 55.17 4.74 ;
        RECT 51.685 4.13 54.435 4.745 ;
        RECT 45.045 4.135 51.03 4.745 ;
        RECT 48.895 4.13 50.875 4.75 ;
        RECT 27.825 4.19 37.97 4.74 ;
        RECT 27.82 4.135 37.95 4.67 ;
        RECT 33.805 4.13 37.95 4.74 ;
        RECT 34.465 4.13 37.215 4.745 ;
        RECT 27.825 4.135 33.81 4.745 ;
        RECT 31.675 4.13 33.655 4.75 ;
        RECT 10.605 4.19 20.75 4.74 ;
        RECT 10.6 4.135 20.73 4.67 ;
        RECT 16.585 4.13 20.73 4.74 ;
        RECT 17.245 4.13 19.995 4.745 ;
        RECT 10.605 4.135 16.59 4.745 ;
        RECT 14.455 4.13 16.435 4.75 ;
        RECT -3.44 4.19 3.53 4.74 ;
        RECT -3.44 4.13 3.51 4.74 ;
        RECT 0.025 4.13 2.775 4.745 ;
        RECT -3.385 4.13 -0.635 4.745 ;
        RECT -1.46 6.655 -1.17 6.885 ;
        RECT -1.63 6.685 -1.17 6.855 ;
      LAYER mcon ;
        RECT -1.4 6.685 -1.23 6.855 ;
        RECT -1.09 4.545 -0.92 4.715 ;
        RECT 2.32 4.545 2.49 4.715 ;
        RECT 3.3 4.345 3.47 4.515 ;
        RECT 3.76 4.345 3.93 4.515 ;
        RECT 4.22 4.345 4.39 4.515 ;
        RECT 4.68 4.345 4.85 4.515 ;
        RECT 5.14 4.345 5.31 4.515 ;
        RECT 5.6 4.345 5.77 4.515 ;
        RECT 6.06 4.345 6.23 4.515 ;
        RECT 6.52 4.345 6.69 4.515 ;
        RECT 6.98 4.345 7.15 4.515 ;
        RECT 7.44 4.345 7.61 4.515 ;
        RECT 7.9 4.345 8.07 4.515 ;
        RECT 8.36 4.345 8.53 4.515 ;
        RECT 8.82 4.345 8.99 4.515 ;
        RECT 9.28 4.345 9.45 4.515 ;
        RECT 9.74 4.345 9.91 4.515 ;
        RECT 10.2 4.345 10.37 4.515 ;
        RECT 14.005 4.545 14.175 4.715 ;
        RECT 14.005 4.165 14.175 4.335 ;
        RECT 14.705 4.55 14.875 4.72 ;
        RECT 14.705 4.16 14.875 4.33 ;
        RECT 15.695 4.55 15.865 4.72 ;
        RECT 15.695 4.16 15.865 4.33 ;
        RECT 19.54 4.545 19.71 4.715 ;
        RECT 20.52 4.345 20.69 4.515 ;
        RECT 20.98 4.345 21.15 4.515 ;
        RECT 21.44 4.345 21.61 4.515 ;
        RECT 21.9 4.345 22.07 4.515 ;
        RECT 22.36 4.345 22.53 4.515 ;
        RECT 22.82 4.345 22.99 4.515 ;
        RECT 23.28 4.345 23.45 4.515 ;
        RECT 23.74 4.345 23.91 4.515 ;
        RECT 24.2 4.345 24.37 4.515 ;
        RECT 24.66 4.345 24.83 4.515 ;
        RECT 25.12 4.345 25.29 4.515 ;
        RECT 25.58 4.345 25.75 4.515 ;
        RECT 26.04 4.345 26.21 4.515 ;
        RECT 26.5 4.345 26.67 4.515 ;
        RECT 26.96 4.345 27.13 4.515 ;
        RECT 27.42 4.345 27.59 4.515 ;
        RECT 31.225 4.545 31.395 4.715 ;
        RECT 31.225 4.165 31.395 4.335 ;
        RECT 31.925 4.55 32.095 4.72 ;
        RECT 31.925 4.16 32.095 4.33 ;
        RECT 32.915 4.55 33.085 4.72 ;
        RECT 32.915 4.16 33.085 4.33 ;
        RECT 36.76 4.545 36.93 4.715 ;
        RECT 37.74 4.345 37.91 4.515 ;
        RECT 38.2 4.345 38.37 4.515 ;
        RECT 38.66 4.345 38.83 4.515 ;
        RECT 39.12 4.345 39.29 4.515 ;
        RECT 39.58 4.345 39.75 4.515 ;
        RECT 40.04 4.345 40.21 4.515 ;
        RECT 40.5 4.345 40.67 4.515 ;
        RECT 40.96 4.345 41.13 4.515 ;
        RECT 41.42 4.345 41.59 4.515 ;
        RECT 41.88 4.345 42.05 4.515 ;
        RECT 42.34 4.345 42.51 4.515 ;
        RECT 42.8 4.345 42.97 4.515 ;
        RECT 43.26 4.345 43.43 4.515 ;
        RECT 43.72 4.345 43.89 4.515 ;
        RECT 44.18 4.345 44.35 4.515 ;
        RECT 44.64 4.345 44.81 4.515 ;
        RECT 48.445 4.545 48.615 4.715 ;
        RECT 48.445 4.165 48.615 4.335 ;
        RECT 49.145 4.55 49.315 4.72 ;
        RECT 49.145 4.16 49.315 4.33 ;
        RECT 50.135 4.55 50.305 4.72 ;
        RECT 50.135 4.16 50.305 4.33 ;
        RECT 53.98 4.545 54.15 4.715 ;
        RECT 54.96 4.345 55.13 4.515 ;
        RECT 55.42 4.345 55.59 4.515 ;
        RECT 55.88 4.345 56.05 4.515 ;
        RECT 56.34 4.345 56.51 4.515 ;
        RECT 56.8 4.345 56.97 4.515 ;
        RECT 57.26 4.345 57.43 4.515 ;
        RECT 57.72 4.345 57.89 4.515 ;
        RECT 58.18 4.345 58.35 4.515 ;
        RECT 58.64 4.345 58.81 4.515 ;
        RECT 59.1 4.345 59.27 4.515 ;
        RECT 59.56 4.345 59.73 4.515 ;
        RECT 60.02 4.345 60.19 4.515 ;
        RECT 60.48 4.345 60.65 4.515 ;
        RECT 60.94 4.345 61.11 4.515 ;
        RECT 61.4 4.345 61.57 4.515 ;
        RECT 61.86 4.345 62.03 4.515 ;
        RECT 65.665 4.545 65.835 4.715 ;
        RECT 65.665 4.165 65.835 4.335 ;
        RECT 66.365 4.55 66.535 4.72 ;
        RECT 66.365 4.16 66.535 4.33 ;
        RECT 67.355 4.55 67.525 4.72 ;
        RECT 67.355 4.16 67.525 4.33 ;
        RECT 71.2 4.545 71.37 4.715 ;
        RECT 72.18 4.345 72.35 4.515 ;
        RECT 72.64 4.345 72.81 4.515 ;
        RECT 73.1 4.345 73.27 4.515 ;
        RECT 73.56 4.345 73.73 4.515 ;
        RECT 74.02 4.345 74.19 4.515 ;
        RECT 74.48 4.345 74.65 4.515 ;
        RECT 74.94 4.345 75.11 4.515 ;
        RECT 75.4 4.345 75.57 4.515 ;
        RECT 75.86 4.345 76.03 4.515 ;
        RECT 76.32 4.345 76.49 4.515 ;
        RECT 76.78 4.345 76.95 4.515 ;
        RECT 77.24 4.345 77.41 4.515 ;
        RECT 77.7 4.345 77.87 4.515 ;
        RECT 78.16 4.345 78.33 4.515 ;
        RECT 78.62 4.345 78.79 4.515 ;
        RECT 79.08 4.345 79.25 4.515 ;
        RECT 82.885 4.545 83.055 4.715 ;
        RECT 82.885 4.165 83.055 4.335 ;
        RECT 83.585 4.55 83.755 4.72 ;
        RECT 83.585 4.16 83.755 4.33 ;
        RECT 84.575 4.55 84.745 4.72 ;
        RECT 84.575 4.16 84.745 4.33 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 74.42 5.79 74.75 6.12 ;
        RECT 73.95 5.805 74.75 6.105 ;
        RECT 57.2 5.79 57.53 6.12 ;
        RECT 56.73 5.805 57.53 6.105 ;
        RECT 39.98 5.79 40.31 6.12 ;
        RECT 39.51 5.805 40.31 6.105 ;
        RECT 22.76 5.79 23.09 6.12 ;
        RECT 22.29 5.805 23.09 6.105 ;
        RECT 5.54 5.79 5.87 6.12 ;
        RECT 5.07 5.805 5.87 6.105 ;
      LAYER li1 ;
        RECT 85.29 0 85.47 0.305 ;
        RECT -3.44 0 85.47 0.3 ;
        RECT 84.495 0 84.665 0.93 ;
        RECT 83.505 0 83.675 0.93 ;
        RECT 68.07 0 83.34 0.305 ;
        RECT 80.765 0 80.935 0.935 ;
        RECT 72.035 0 79.69 1.795 ;
        RECT 78.93 0 79.26 2.185 ;
        RECT 78.09 0 78.42 2.185 ;
        RECT 76.26 0 76.55 2.63 ;
        RECT 75.81 0 76.08 2.605 ;
        RECT 74.9 0 75.14 2.605 ;
        RECT 74.45 0 74.69 2.605 ;
        RECT 73.51 0 73.78 2.605 ;
        RECT 73.06 0 73.29 2.615 ;
        RECT 72.18 0 72.39 2.615 ;
        RECT 72.03 0 79.69 1.635 ;
        RECT 67.275 0 67.445 0.93 ;
        RECT 66.285 0 66.455 0.93 ;
        RECT 50.85 0 66.12 0.305 ;
        RECT 63.545 0 63.715 0.935 ;
        RECT 54.815 0 62.47 1.795 ;
        RECT 61.71 0 62.04 2.185 ;
        RECT 60.87 0 61.2 2.185 ;
        RECT 59.04 0 59.33 2.63 ;
        RECT 58.59 0 58.86 2.605 ;
        RECT 57.68 0 57.92 2.605 ;
        RECT 57.23 0 57.47 2.605 ;
        RECT 56.29 0 56.56 2.605 ;
        RECT 55.84 0 56.07 2.615 ;
        RECT 54.96 0 55.17 2.615 ;
        RECT 54.81 0 62.47 1.635 ;
        RECT 50.055 0 50.225 0.93 ;
        RECT 49.065 0 49.235 0.93 ;
        RECT 33.63 0 48.9 0.305 ;
        RECT 46.325 0 46.495 0.935 ;
        RECT 37.595 0 45.25 1.795 ;
        RECT 44.49 0 44.82 2.185 ;
        RECT 43.65 0 43.98 2.185 ;
        RECT 41.82 0 42.11 2.63 ;
        RECT 41.37 0 41.64 2.605 ;
        RECT 40.46 0 40.7 2.605 ;
        RECT 40.01 0 40.25 2.605 ;
        RECT 39.07 0 39.34 2.605 ;
        RECT 38.62 0 38.85 2.615 ;
        RECT 37.74 0 37.95 2.615 ;
        RECT 37.59 0 45.25 1.635 ;
        RECT 32.835 0 33.005 0.93 ;
        RECT 31.845 0 32.015 0.93 ;
        RECT 16.41 0 31.68 0.305 ;
        RECT 29.105 0 29.275 0.935 ;
        RECT 20.375 0 28.03 1.795 ;
        RECT 27.27 0 27.6 2.185 ;
        RECT 26.43 0 26.76 2.185 ;
        RECT 24.6 0 24.89 2.63 ;
        RECT 24.15 0 24.42 2.605 ;
        RECT 23.24 0 23.48 2.605 ;
        RECT 22.79 0 23.03 2.605 ;
        RECT 21.85 0 22.12 2.605 ;
        RECT 21.4 0 21.63 2.615 ;
        RECT 20.52 0 20.73 2.615 ;
        RECT 20.37 0 28.03 1.635 ;
        RECT 15.615 0 15.785 0.93 ;
        RECT 14.625 0 14.795 0.93 ;
        RECT -3.44 0 14.46 0.305 ;
        RECT 11.885 0 12.055 0.935 ;
        RECT 3.155 0 10.81 1.795 ;
        RECT 10.05 0 10.38 2.185 ;
        RECT 9.21 0 9.54 2.185 ;
        RECT 7.38 0 7.67 2.63 ;
        RECT 6.93 0 7.2 2.605 ;
        RECT 6.02 0 6.26 2.605 ;
        RECT 5.57 0 5.81 2.605 ;
        RECT 4.63 0 4.9 2.605 ;
        RECT 4.18 0 4.41 2.615 ;
        RECT 3.3 0 3.51 2.615 ;
        RECT 3.15 0 10.81 1.635 ;
        RECT -3.44 8.58 85.47 8.88 ;
        RECT 85.29 8.575 85.47 8.88 ;
        RECT 84.495 7.95 84.665 8.88 ;
        RECT 83.505 7.95 83.675 8.88 ;
        RECT 68.07 8.575 83.34 8.88 ;
        RECT 80.765 7.945 80.935 8.88 ;
        RECT 72.305 7.18 79.505 8.88 ;
        RECT 72.035 7.065 79.395 7.235 ;
        RECT 78.54 6.265 78.85 8.88 ;
        RECT 77.16 6.265 77.47 8.88 ;
        RECT 74.89 5.825 75.225 6.095 ;
        RECT 74.88 6.265 75.19 8.88 ;
        RECT 74.5 5.875 75.225 6.045 ;
        RECT 74.51 5.875 74.68 8.88 ;
        RECT 72.58 6.265 72.89 8.88 ;
        RECT 69.08 7.945 69.25 8.88 ;
        RECT 67.275 7.95 67.445 8.88 ;
        RECT 66.285 7.95 66.455 8.88 ;
        RECT 50.85 8.575 66.12 8.88 ;
        RECT 63.545 7.945 63.715 8.88 ;
        RECT 55.085 7.18 62.285 8.88 ;
        RECT 54.815 7.065 62.175 7.235 ;
        RECT 61.32 6.265 61.63 8.88 ;
        RECT 59.94 6.265 60.25 8.88 ;
        RECT 57.67 5.825 58.005 6.095 ;
        RECT 57.66 6.265 57.97 8.88 ;
        RECT 57.28 5.875 58.005 6.045 ;
        RECT 57.29 5.875 57.46 8.88 ;
        RECT 55.36 6.265 55.67 8.88 ;
        RECT 51.86 7.945 52.03 8.88 ;
        RECT 50.055 7.95 50.225 8.88 ;
        RECT 49.065 7.95 49.235 8.88 ;
        RECT 33.63 8.575 48.9 8.88 ;
        RECT 46.325 7.945 46.495 8.88 ;
        RECT 37.865 7.18 45.065 8.88 ;
        RECT 37.595 7.065 44.955 7.235 ;
        RECT 44.1 6.265 44.41 8.88 ;
        RECT 42.72 6.265 43.03 8.88 ;
        RECT 40.45 5.825 40.785 6.095 ;
        RECT 40.44 6.265 40.75 8.88 ;
        RECT 40.06 5.875 40.785 6.045 ;
        RECT 40.07 5.875 40.24 8.88 ;
        RECT 38.14 6.265 38.45 8.88 ;
        RECT 34.64 7.945 34.81 8.88 ;
        RECT 32.835 7.95 33.005 8.88 ;
        RECT 31.845 7.95 32.015 8.88 ;
        RECT 16.41 8.575 31.68 8.88 ;
        RECT 29.105 7.945 29.275 8.88 ;
        RECT 20.645 7.18 27.845 8.88 ;
        RECT 20.375 7.065 27.735 7.235 ;
        RECT 26.88 6.265 27.19 8.88 ;
        RECT 25.5 6.265 25.81 8.88 ;
        RECT 23.23 5.825 23.565 6.095 ;
        RECT 23.22 6.265 23.53 8.88 ;
        RECT 22.84 5.875 23.565 6.045 ;
        RECT 22.85 5.875 23.02 8.88 ;
        RECT 20.92 6.265 21.23 8.88 ;
        RECT 17.42 7.945 17.59 8.88 ;
        RECT 15.615 7.95 15.785 8.88 ;
        RECT 14.625 7.95 14.795 8.88 ;
        RECT -3.44 8.575 14.46 8.88 ;
        RECT 11.885 7.945 12.055 8.88 ;
        RECT 3.425 7.18 10.625 8.88 ;
        RECT 3.155 7.065 10.515 7.235 ;
        RECT 9.66 6.265 9.97 8.88 ;
        RECT 8.28 6.265 8.59 8.88 ;
        RECT 6.01 5.825 6.345 6.095 ;
        RECT 6 6.265 6.31 8.88 ;
        RECT 5.62 5.875 6.345 6.045 ;
        RECT 5.63 5.875 5.8 8.88 ;
        RECT 3.7 6.265 4.01 8.88 ;
        RECT 0.2 7.945 0.37 8.88 ;
        RECT -3.21 7.945 -3.04 8.88 ;
        RECT 72.59 5.825 72.925 6.095 ;
        RECT 72.12 5.875 72.925 6.045 ;
        RECT 70.085 6.075 70.255 8.025 ;
        RECT 70.03 7.855 70.2 8.305 ;
        RECT 70.03 5.015 70.2 6.245 ;
        RECT 55.37 5.825 55.705 6.095 ;
        RECT 54.9 5.875 55.705 6.045 ;
        RECT 52.865 6.075 53.035 8.025 ;
        RECT 52.81 7.855 52.98 8.305 ;
        RECT 52.81 5.015 52.98 6.245 ;
        RECT 38.15 5.825 38.485 6.095 ;
        RECT 37.68 5.875 38.485 6.045 ;
        RECT 35.645 6.075 35.815 8.025 ;
        RECT 35.59 7.855 35.76 8.305 ;
        RECT 35.59 5.015 35.76 6.245 ;
        RECT 20.93 5.825 21.265 6.095 ;
        RECT 20.46 5.875 21.265 6.045 ;
        RECT 18.425 6.075 18.595 8.025 ;
        RECT 18.37 7.855 18.54 8.305 ;
        RECT 18.37 5.015 18.54 6.245 ;
        RECT 3.71 5.825 4.045 6.095 ;
        RECT 3.24 5.875 4.045 6.045 ;
        RECT 1.205 6.075 1.375 8.025 ;
        RECT 1.15 7.855 1.32 8.305 ;
        RECT 1.15 5.015 1.32 6.245 ;
      LAYER met2 ;
        RECT 74.445 5.77 74.725 6.14 ;
        RECT 57.225 5.77 57.505 6.14 ;
        RECT 40.005 5.77 40.285 6.14 ;
        RECT 22.785 5.77 23.065 6.14 ;
        RECT 5.565 5.77 5.845 6.14 ;
      LAYER met1 ;
        RECT 85.29 0 85.47 0.305 ;
        RECT -3.44 0 85.47 0.3 ;
        RECT 68.07 0 83.34 0.305 ;
        RECT 72.035 0 79.69 1.795 ;
        RECT 72.035 0 79.395 1.95 ;
        RECT 72.03 0 79.69 1.635 ;
        RECT 50.85 0 66.12 0.305 ;
        RECT 54.815 0 62.47 1.795 ;
        RECT 54.815 0 62.175 1.95 ;
        RECT 54.81 0 62.47 1.635 ;
        RECT 33.63 0 48.9 0.305 ;
        RECT 37.595 0 45.25 1.795 ;
        RECT 37.595 0 44.955 1.95 ;
        RECT 37.59 0 45.25 1.635 ;
        RECT 16.41 0 31.68 0.305 ;
        RECT 20.375 0 28.03 1.795 ;
        RECT 20.375 0 27.735 1.95 ;
        RECT 20.37 0 28.03 1.635 ;
        RECT -3.44 0 14.46 0.305 ;
        RECT 3.155 0 10.81 1.795 ;
        RECT 3.155 0 10.515 1.95 ;
        RECT 3.15 0 10.81 1.635 ;
        RECT -3.44 8.58 85.47 8.88 ;
        RECT 85.29 8.575 85.47 8.88 ;
        RECT 68.07 8.575 83.34 8.88 ;
        RECT 72.305 7.18 79.505 8.88 ;
        RECT 72.035 6.91 79.395 7.39 ;
        RECT 70.025 6.285 70.315 6.515 ;
        RECT 69.625 6.315 70.315 6.485 ;
        RECT 69.625 6.315 69.795 8.88 ;
        RECT 50.85 8.575 66.12 8.88 ;
        RECT 55.085 7.18 62.285 8.88 ;
        RECT 54.815 6.91 62.175 7.39 ;
        RECT 52.805 6.285 53.095 6.515 ;
        RECT 52.405 6.315 53.095 6.485 ;
        RECT 52.405 6.315 52.575 8.88 ;
        RECT 33.63 8.575 48.9 8.88 ;
        RECT 37.865 7.18 45.065 8.88 ;
        RECT 37.595 6.91 44.955 7.39 ;
        RECT 35.585 6.285 35.875 6.515 ;
        RECT 35.185 6.315 35.875 6.485 ;
        RECT 35.185 6.315 35.355 8.88 ;
        RECT 16.41 8.575 31.68 8.88 ;
        RECT 20.645 7.18 27.845 8.88 ;
        RECT 20.375 6.91 27.735 7.39 ;
        RECT 18.365 6.285 18.655 6.515 ;
        RECT 17.965 6.315 18.655 6.485 ;
        RECT 17.965 6.315 18.135 8.88 ;
        RECT -3.44 8.575 14.46 8.88 ;
        RECT 3.425 7.18 10.625 8.88 ;
        RECT 3.155 6.91 10.515 7.39 ;
        RECT 1.145 6.285 1.435 6.515 ;
        RECT 0.745 6.315 1.435 6.485 ;
        RECT 0.745 6.315 0.915 8.88 ;
        RECT 74.425 5.83 74.745 6.09 ;
        RECT 72.06 5.89 74.745 6.03 ;
        RECT 72.06 5.845 72.35 6.075 ;
        RECT 57.205 5.83 57.525 6.09 ;
        RECT 54.84 5.89 57.525 6.03 ;
        RECT 54.84 5.845 55.13 6.075 ;
        RECT 39.985 5.83 40.305 6.09 ;
        RECT 37.62 5.89 40.305 6.03 ;
        RECT 37.62 5.845 37.91 6.075 ;
        RECT 22.765 5.83 23.085 6.09 ;
        RECT 20.4 5.89 23.085 6.03 ;
        RECT 20.4 5.845 20.69 6.075 ;
        RECT 5.545 5.83 5.865 6.09 ;
        RECT 3.18 5.89 5.865 6.03 ;
        RECT 3.18 5.845 3.47 6.075 ;
      LAYER via2 ;
        RECT 5.605 5.855 5.805 6.055 ;
        RECT 22.825 5.855 23.025 6.055 ;
        RECT 40.045 5.855 40.245 6.055 ;
        RECT 57.265 5.855 57.465 6.055 ;
        RECT 74.485 5.855 74.685 6.055 ;
      LAYER via1 ;
        RECT 5.63 5.885 5.78 6.035 ;
        RECT 22.85 5.885 23 6.035 ;
        RECT 40.07 5.885 40.22 6.035 ;
        RECT 57.29 5.885 57.44 6.035 ;
        RECT 74.51 5.885 74.66 6.035 ;
      LAYER mcon ;
        RECT -3.13 8.605 -2.96 8.775 ;
        RECT -2.45 8.605 -2.28 8.775 ;
        RECT -1.77 8.605 -1.6 8.775 ;
        RECT -1.09 8.605 -0.92 8.775 ;
        RECT 0.28 8.605 0.45 8.775 ;
        RECT 0.96 8.605 1.13 8.775 ;
        RECT 1.205 6.315 1.375 6.485 ;
        RECT 1.64 8.605 1.81 8.775 ;
        RECT 2.32 8.605 2.49 8.775 ;
        RECT 3.24 5.875 3.41 6.045 ;
        RECT 3.3 7.065 3.47 7.235 ;
        RECT 3.3 1.625 3.47 1.795 ;
        RECT 3.76 7.065 3.93 7.235 ;
        RECT 3.76 1.625 3.93 1.795 ;
        RECT 4.22 7.065 4.39 7.235 ;
        RECT 4.22 1.625 4.39 1.795 ;
        RECT 4.68 7.065 4.85 7.235 ;
        RECT 4.68 1.625 4.85 1.795 ;
        RECT 5.14 7.065 5.31 7.235 ;
        RECT 5.14 1.625 5.31 1.795 ;
        RECT 5.6 7.065 5.77 7.235 ;
        RECT 5.6 1.625 5.77 1.795 ;
        RECT 5.62 5.875 5.79 6.045 ;
        RECT 6.06 7.065 6.23 7.235 ;
        RECT 6.06 1.625 6.23 1.795 ;
        RECT 6.52 7.065 6.69 7.235 ;
        RECT 6.52 1.625 6.69 1.795 ;
        RECT 6.98 7.065 7.15 7.235 ;
        RECT 6.98 1.625 7.15 1.795 ;
        RECT 7.44 7.065 7.61 7.235 ;
        RECT 7.44 1.625 7.61 1.795 ;
        RECT 7.9 7.065 8.07 7.235 ;
        RECT 7.9 1.625 8.07 1.795 ;
        RECT 8.36 7.065 8.53 7.235 ;
        RECT 8.36 1.625 8.53 1.795 ;
        RECT 8.82 7.065 8.99 7.235 ;
        RECT 8.82 1.625 8.99 1.795 ;
        RECT 9.28 7.065 9.45 7.235 ;
        RECT 9.28 1.625 9.45 1.795 ;
        RECT 9.74 7.065 9.91 7.235 ;
        RECT 9.74 1.625 9.91 1.795 ;
        RECT 10.2 7.065 10.37 7.235 ;
        RECT 10.2 1.625 10.37 1.795 ;
        RECT 11.965 8.605 12.135 8.775 ;
        RECT 11.965 0.105 12.135 0.275 ;
        RECT 12.645 8.605 12.815 8.775 ;
        RECT 12.645 0.105 12.815 0.275 ;
        RECT 13.325 8.605 13.495 8.775 ;
        RECT 13.325 0.105 13.495 0.275 ;
        RECT 14.005 8.605 14.175 8.775 ;
        RECT 14.005 0.105 14.175 0.275 ;
        RECT 14.705 8.61 14.875 8.78 ;
        RECT 14.705 0.1 14.875 0.27 ;
        RECT 15.695 8.61 15.865 8.78 ;
        RECT 15.695 0.1 15.865 0.27 ;
        RECT 17.5 8.605 17.67 8.775 ;
        RECT 18.18 8.605 18.35 8.775 ;
        RECT 18.425 6.315 18.595 6.485 ;
        RECT 18.86 8.605 19.03 8.775 ;
        RECT 19.54 8.605 19.71 8.775 ;
        RECT 20.46 5.875 20.63 6.045 ;
        RECT 20.52 7.065 20.69 7.235 ;
        RECT 20.52 1.625 20.69 1.795 ;
        RECT 20.98 7.065 21.15 7.235 ;
        RECT 20.98 1.625 21.15 1.795 ;
        RECT 21.44 7.065 21.61 7.235 ;
        RECT 21.44 1.625 21.61 1.795 ;
        RECT 21.9 7.065 22.07 7.235 ;
        RECT 21.9 1.625 22.07 1.795 ;
        RECT 22.36 7.065 22.53 7.235 ;
        RECT 22.36 1.625 22.53 1.795 ;
        RECT 22.82 7.065 22.99 7.235 ;
        RECT 22.82 1.625 22.99 1.795 ;
        RECT 22.84 5.875 23.01 6.045 ;
        RECT 23.28 7.065 23.45 7.235 ;
        RECT 23.28 1.625 23.45 1.795 ;
        RECT 23.74 7.065 23.91 7.235 ;
        RECT 23.74 1.625 23.91 1.795 ;
        RECT 24.2 7.065 24.37 7.235 ;
        RECT 24.2 1.625 24.37 1.795 ;
        RECT 24.66 7.065 24.83 7.235 ;
        RECT 24.66 1.625 24.83 1.795 ;
        RECT 25.12 7.065 25.29 7.235 ;
        RECT 25.12 1.625 25.29 1.795 ;
        RECT 25.58 7.065 25.75 7.235 ;
        RECT 25.58 1.625 25.75 1.795 ;
        RECT 26.04 7.065 26.21 7.235 ;
        RECT 26.04 1.625 26.21 1.795 ;
        RECT 26.5 7.065 26.67 7.235 ;
        RECT 26.5 1.625 26.67 1.795 ;
        RECT 26.96 7.065 27.13 7.235 ;
        RECT 26.96 1.625 27.13 1.795 ;
        RECT 27.42 7.065 27.59 7.235 ;
        RECT 27.42 1.625 27.59 1.795 ;
        RECT 29.185 8.605 29.355 8.775 ;
        RECT 29.185 0.105 29.355 0.275 ;
        RECT 29.865 8.605 30.035 8.775 ;
        RECT 29.865 0.105 30.035 0.275 ;
        RECT 30.545 8.605 30.715 8.775 ;
        RECT 30.545 0.105 30.715 0.275 ;
        RECT 31.225 8.605 31.395 8.775 ;
        RECT 31.225 0.105 31.395 0.275 ;
        RECT 31.925 8.61 32.095 8.78 ;
        RECT 31.925 0.1 32.095 0.27 ;
        RECT 32.915 8.61 33.085 8.78 ;
        RECT 32.915 0.1 33.085 0.27 ;
        RECT 34.72 8.605 34.89 8.775 ;
        RECT 35.4 8.605 35.57 8.775 ;
        RECT 35.645 6.315 35.815 6.485 ;
        RECT 36.08 8.605 36.25 8.775 ;
        RECT 36.76 8.605 36.93 8.775 ;
        RECT 37.68 5.875 37.85 6.045 ;
        RECT 37.74 7.065 37.91 7.235 ;
        RECT 37.74 1.625 37.91 1.795 ;
        RECT 38.2 7.065 38.37 7.235 ;
        RECT 38.2 1.625 38.37 1.795 ;
        RECT 38.66 7.065 38.83 7.235 ;
        RECT 38.66 1.625 38.83 1.795 ;
        RECT 39.12 7.065 39.29 7.235 ;
        RECT 39.12 1.625 39.29 1.795 ;
        RECT 39.58 7.065 39.75 7.235 ;
        RECT 39.58 1.625 39.75 1.795 ;
        RECT 40.04 7.065 40.21 7.235 ;
        RECT 40.04 1.625 40.21 1.795 ;
        RECT 40.06 5.875 40.23 6.045 ;
        RECT 40.5 7.065 40.67 7.235 ;
        RECT 40.5 1.625 40.67 1.795 ;
        RECT 40.96 7.065 41.13 7.235 ;
        RECT 40.96 1.625 41.13 1.795 ;
        RECT 41.42 7.065 41.59 7.235 ;
        RECT 41.42 1.625 41.59 1.795 ;
        RECT 41.88 7.065 42.05 7.235 ;
        RECT 41.88 1.625 42.05 1.795 ;
        RECT 42.34 7.065 42.51 7.235 ;
        RECT 42.34 1.625 42.51 1.795 ;
        RECT 42.8 7.065 42.97 7.235 ;
        RECT 42.8 1.625 42.97 1.795 ;
        RECT 43.26 7.065 43.43 7.235 ;
        RECT 43.26 1.625 43.43 1.795 ;
        RECT 43.72 7.065 43.89 7.235 ;
        RECT 43.72 1.625 43.89 1.795 ;
        RECT 44.18 7.065 44.35 7.235 ;
        RECT 44.18 1.625 44.35 1.795 ;
        RECT 44.64 7.065 44.81 7.235 ;
        RECT 44.64 1.625 44.81 1.795 ;
        RECT 46.405 8.605 46.575 8.775 ;
        RECT 46.405 0.105 46.575 0.275 ;
        RECT 47.085 8.605 47.255 8.775 ;
        RECT 47.085 0.105 47.255 0.275 ;
        RECT 47.765 8.605 47.935 8.775 ;
        RECT 47.765 0.105 47.935 0.275 ;
        RECT 48.445 8.605 48.615 8.775 ;
        RECT 48.445 0.105 48.615 0.275 ;
        RECT 49.145 8.61 49.315 8.78 ;
        RECT 49.145 0.1 49.315 0.27 ;
        RECT 50.135 8.61 50.305 8.78 ;
        RECT 50.135 0.1 50.305 0.27 ;
        RECT 51.94 8.605 52.11 8.775 ;
        RECT 52.62 8.605 52.79 8.775 ;
        RECT 52.865 6.315 53.035 6.485 ;
        RECT 53.3 8.605 53.47 8.775 ;
        RECT 53.98 8.605 54.15 8.775 ;
        RECT 54.9 5.875 55.07 6.045 ;
        RECT 54.96 7.065 55.13 7.235 ;
        RECT 54.96 1.625 55.13 1.795 ;
        RECT 55.42 7.065 55.59 7.235 ;
        RECT 55.42 1.625 55.59 1.795 ;
        RECT 55.88 7.065 56.05 7.235 ;
        RECT 55.88 1.625 56.05 1.795 ;
        RECT 56.34 7.065 56.51 7.235 ;
        RECT 56.34 1.625 56.51 1.795 ;
        RECT 56.8 7.065 56.97 7.235 ;
        RECT 56.8 1.625 56.97 1.795 ;
        RECT 57.26 7.065 57.43 7.235 ;
        RECT 57.26 1.625 57.43 1.795 ;
        RECT 57.28 5.875 57.45 6.045 ;
        RECT 57.72 7.065 57.89 7.235 ;
        RECT 57.72 1.625 57.89 1.795 ;
        RECT 58.18 7.065 58.35 7.235 ;
        RECT 58.18 1.625 58.35 1.795 ;
        RECT 58.64 7.065 58.81 7.235 ;
        RECT 58.64 1.625 58.81 1.795 ;
        RECT 59.1 7.065 59.27 7.235 ;
        RECT 59.1 1.625 59.27 1.795 ;
        RECT 59.56 7.065 59.73 7.235 ;
        RECT 59.56 1.625 59.73 1.795 ;
        RECT 60.02 7.065 60.19 7.235 ;
        RECT 60.02 1.625 60.19 1.795 ;
        RECT 60.48 7.065 60.65 7.235 ;
        RECT 60.48 1.625 60.65 1.795 ;
        RECT 60.94 7.065 61.11 7.235 ;
        RECT 60.94 1.625 61.11 1.795 ;
        RECT 61.4 7.065 61.57 7.235 ;
        RECT 61.4 1.625 61.57 1.795 ;
        RECT 61.86 7.065 62.03 7.235 ;
        RECT 61.86 1.625 62.03 1.795 ;
        RECT 63.625 8.605 63.795 8.775 ;
        RECT 63.625 0.105 63.795 0.275 ;
        RECT 64.305 8.605 64.475 8.775 ;
        RECT 64.305 0.105 64.475 0.275 ;
        RECT 64.985 8.605 65.155 8.775 ;
        RECT 64.985 0.105 65.155 0.275 ;
        RECT 65.665 8.605 65.835 8.775 ;
        RECT 65.665 0.105 65.835 0.275 ;
        RECT 66.365 8.61 66.535 8.78 ;
        RECT 66.365 0.1 66.535 0.27 ;
        RECT 67.355 8.61 67.525 8.78 ;
        RECT 67.355 0.1 67.525 0.27 ;
        RECT 69.16 8.605 69.33 8.775 ;
        RECT 69.84 8.605 70.01 8.775 ;
        RECT 70.085 6.315 70.255 6.485 ;
        RECT 70.52 8.605 70.69 8.775 ;
        RECT 71.2 8.605 71.37 8.775 ;
        RECT 72.12 5.875 72.29 6.045 ;
        RECT 72.18 7.065 72.35 7.235 ;
        RECT 72.18 1.625 72.35 1.795 ;
        RECT 72.64 7.065 72.81 7.235 ;
        RECT 72.64 1.625 72.81 1.795 ;
        RECT 73.1 7.065 73.27 7.235 ;
        RECT 73.1 1.625 73.27 1.795 ;
        RECT 73.56 7.065 73.73 7.235 ;
        RECT 73.56 1.625 73.73 1.795 ;
        RECT 74.02 7.065 74.19 7.235 ;
        RECT 74.02 1.625 74.19 1.795 ;
        RECT 74.48 7.065 74.65 7.235 ;
        RECT 74.48 1.625 74.65 1.795 ;
        RECT 74.5 5.875 74.67 6.045 ;
        RECT 74.94 7.065 75.11 7.235 ;
        RECT 74.94 1.625 75.11 1.795 ;
        RECT 75.4 7.065 75.57 7.235 ;
        RECT 75.4 1.625 75.57 1.795 ;
        RECT 75.86 7.065 76.03 7.235 ;
        RECT 75.86 1.625 76.03 1.795 ;
        RECT 76.32 7.065 76.49 7.235 ;
        RECT 76.32 1.625 76.49 1.795 ;
        RECT 76.78 7.065 76.95 7.235 ;
        RECT 76.78 1.625 76.95 1.795 ;
        RECT 77.24 7.065 77.41 7.235 ;
        RECT 77.24 1.625 77.41 1.795 ;
        RECT 77.7 7.065 77.87 7.235 ;
        RECT 77.7 1.625 77.87 1.795 ;
        RECT 78.16 7.065 78.33 7.235 ;
        RECT 78.16 1.625 78.33 1.795 ;
        RECT 78.62 7.065 78.79 7.235 ;
        RECT 78.62 1.625 78.79 1.795 ;
        RECT 79.08 7.065 79.25 7.235 ;
        RECT 79.08 1.625 79.25 1.795 ;
        RECT 80.845 8.605 81.015 8.775 ;
        RECT 80.845 0.105 81.015 0.275 ;
        RECT 81.525 8.605 81.695 8.775 ;
        RECT 81.525 0.105 81.695 0.275 ;
        RECT 82.205 8.605 82.375 8.775 ;
        RECT 82.205 0.105 82.375 0.275 ;
        RECT 82.885 8.605 83.055 8.775 ;
        RECT 82.885 0.105 83.055 0.275 ;
        RECT 83.585 8.61 83.755 8.78 ;
        RECT 83.585 0.1 83.755 0.27 ;
        RECT 84.575 8.61 84.745 8.78 ;
        RECT 84.575 0.1 84.745 0.27 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 71.5 7.435 77.515 7.735 ;
      RECT 77.215 5.805 77.515 7.735 ;
      RECT 76.16 5.785 76.46 7.735 ;
      RECT 75.13 6.48 75.43 7.735 ;
      RECT 71.5 7.035 71.8 7.735 ;
      RECT 70.365 7 70.735 7.37 ;
      RECT 70.365 7.035 71.8 7.335 ;
      RECT 75.1 6.48 75.43 6.81 ;
      RECT 74.63 6.495 75.43 6.795 ;
      RECT 75.01 6.455 75.31 6.795 ;
      RECT 77.14 5.805 77.515 6.17 ;
      RECT 77.205 5.765 77.505 6.17 ;
      RECT 76.12 5.785 76.46 6.135 ;
      RECT 76.135 5.745 76.435 6.135 ;
      RECT 76.11 5.79 76.46 6.12 ;
      RECT 77.14 5.805 77.95 6.105 ;
      RECT 75.64 5.805 76.46 6.105 ;
      RECT 77.15 5.79 77.505 6.17 ;
      RECT 76.8 3.755 77.13 4.085 ;
      RECT 76.8 3.77 77.6 4.07 ;
      RECT 76.815 3.725 77.115 4.085 ;
      RECT 76.46 3.075 76.79 3.405 ;
      RECT 76.46 3.09 77.26 3.39 ;
      RECT 76.545 3.065 76.845 3.39 ;
      RECT 75.78 4.155 76.11 4.485 ;
      RECT 73.74 4.155 74.07 4.485 ;
      RECT 73.74 4.17 76.11 4.47 ;
      RECT 75.43 3.415 75.76 3.745 ;
      RECT 74.97 3.43 75.77 3.73 ;
      RECT 75.1 2.225 75.43 2.555 ;
      RECT 74.63 2.24 75.43 2.54 ;
      RECT 75.09 2.235 75.43 2.54 ;
      RECT 54.28 7.435 60.295 7.735 ;
      RECT 59.995 5.805 60.295 7.735 ;
      RECT 58.94 5.785 59.24 7.735 ;
      RECT 57.91 6.48 58.21 7.735 ;
      RECT 54.28 7.035 54.58 7.735 ;
      RECT 53.145 7 53.515 7.37 ;
      RECT 53.145 7.035 54.58 7.335 ;
      RECT 57.88 6.48 58.21 6.81 ;
      RECT 57.41 6.495 58.21 6.795 ;
      RECT 57.79 6.455 58.09 6.795 ;
      RECT 59.92 5.805 60.295 6.17 ;
      RECT 59.985 5.765 60.285 6.17 ;
      RECT 58.9 5.785 59.24 6.135 ;
      RECT 58.915 5.745 59.215 6.135 ;
      RECT 58.89 5.79 59.24 6.12 ;
      RECT 59.92 5.805 60.73 6.105 ;
      RECT 58.42 5.805 59.24 6.105 ;
      RECT 59.93 5.79 60.285 6.17 ;
      RECT 59.58 3.755 59.91 4.085 ;
      RECT 59.58 3.77 60.38 4.07 ;
      RECT 59.595 3.725 59.895 4.085 ;
      RECT 59.24 3.075 59.57 3.405 ;
      RECT 59.24 3.09 60.04 3.39 ;
      RECT 59.325 3.065 59.625 3.39 ;
      RECT 58.56 4.155 58.89 4.485 ;
      RECT 56.52 4.155 56.85 4.485 ;
      RECT 56.52 4.17 58.89 4.47 ;
      RECT 58.21 3.415 58.54 3.745 ;
      RECT 57.75 3.43 58.55 3.73 ;
      RECT 57.88 2.225 58.21 2.555 ;
      RECT 57.41 2.24 58.21 2.54 ;
      RECT 57.87 2.235 58.21 2.54 ;
      RECT 37.06 7.435 43.075 7.735 ;
      RECT 42.775 5.805 43.075 7.735 ;
      RECT 41.72 5.785 42.02 7.735 ;
      RECT 40.69 6.48 40.99 7.735 ;
      RECT 37.06 7.035 37.36 7.735 ;
      RECT 35.925 7 36.295 7.37 ;
      RECT 35.925 7.035 37.36 7.335 ;
      RECT 40.66 6.48 40.99 6.81 ;
      RECT 40.19 6.495 40.99 6.795 ;
      RECT 40.57 6.455 40.87 6.795 ;
      RECT 42.7 5.805 43.075 6.17 ;
      RECT 42.765 5.765 43.065 6.17 ;
      RECT 41.68 5.785 42.02 6.135 ;
      RECT 41.695 5.745 41.995 6.135 ;
      RECT 41.67 5.79 42.02 6.12 ;
      RECT 42.7 5.805 43.51 6.105 ;
      RECT 41.2 5.805 42.02 6.105 ;
      RECT 42.71 5.79 43.065 6.17 ;
      RECT 42.36 3.755 42.69 4.085 ;
      RECT 42.36 3.77 43.16 4.07 ;
      RECT 42.375 3.725 42.675 4.085 ;
      RECT 42.02 3.075 42.35 3.405 ;
      RECT 42.02 3.09 42.82 3.39 ;
      RECT 42.105 3.065 42.405 3.39 ;
      RECT 41.34 4.155 41.67 4.485 ;
      RECT 39.3 4.155 39.63 4.485 ;
      RECT 39.3 4.17 41.67 4.47 ;
      RECT 40.99 3.415 41.32 3.745 ;
      RECT 40.53 3.43 41.33 3.73 ;
      RECT 40.66 2.225 40.99 2.555 ;
      RECT 40.19 2.24 40.99 2.54 ;
      RECT 40.65 2.235 40.99 2.54 ;
      RECT 19.84 7.435 25.855 7.735 ;
      RECT 25.555 5.805 25.855 7.735 ;
      RECT 24.5 5.785 24.8 7.735 ;
      RECT 23.47 6.48 23.77 7.735 ;
      RECT 19.84 7.035 20.14 7.735 ;
      RECT 18.705 7 19.075 7.37 ;
      RECT 18.705 7.035 20.14 7.335 ;
      RECT 23.44 6.48 23.77 6.81 ;
      RECT 22.97 6.495 23.77 6.795 ;
      RECT 23.35 6.455 23.65 6.795 ;
      RECT 25.48 5.805 25.855 6.17 ;
      RECT 25.545 5.765 25.845 6.17 ;
      RECT 24.46 5.785 24.8 6.135 ;
      RECT 24.475 5.745 24.775 6.135 ;
      RECT 24.45 5.79 24.8 6.12 ;
      RECT 25.48 5.805 26.29 6.105 ;
      RECT 23.98 5.805 24.8 6.105 ;
      RECT 25.49 5.79 25.845 6.17 ;
      RECT 25.14 3.755 25.47 4.085 ;
      RECT 25.14 3.77 25.94 4.07 ;
      RECT 25.155 3.725 25.455 4.085 ;
      RECT 24.8 3.075 25.13 3.405 ;
      RECT 24.8 3.09 25.6 3.39 ;
      RECT 24.885 3.065 25.185 3.39 ;
      RECT 24.12 4.155 24.45 4.485 ;
      RECT 22.08 4.155 22.41 4.485 ;
      RECT 22.08 4.17 24.45 4.47 ;
      RECT 23.77 3.415 24.1 3.745 ;
      RECT 23.31 3.43 24.11 3.73 ;
      RECT 23.44 2.225 23.77 2.555 ;
      RECT 22.97 2.24 23.77 2.54 ;
      RECT 23.43 2.235 23.77 2.54 ;
      RECT 2.62 7.435 8.635 7.735 ;
      RECT 8.335 5.805 8.635 7.735 ;
      RECT 7.28 5.785 7.58 7.735 ;
      RECT 6.25 6.48 6.55 7.735 ;
      RECT 2.62 7.035 2.92 7.735 ;
      RECT 1.485 7 1.855 7.37 ;
      RECT 1.485 7.035 2.92 7.335 ;
      RECT 6.22 6.48 6.55 6.81 ;
      RECT 5.75 6.495 6.55 6.795 ;
      RECT 6.13 6.455 6.43 6.795 ;
      RECT 8.26 5.805 8.635 6.17 ;
      RECT 8.325 5.765 8.625 6.17 ;
      RECT 7.24 5.785 7.58 6.135 ;
      RECT 7.255 5.745 7.555 6.135 ;
      RECT 7.23 5.79 7.58 6.12 ;
      RECT 8.26 5.805 9.07 6.105 ;
      RECT 6.76 5.805 7.58 6.105 ;
      RECT 8.27 5.79 8.625 6.17 ;
      RECT 7.92 3.755 8.25 4.085 ;
      RECT 7.92 3.77 8.72 4.07 ;
      RECT 7.935 3.725 8.235 4.085 ;
      RECT 7.58 3.075 7.91 3.405 ;
      RECT 7.58 3.09 8.38 3.39 ;
      RECT 7.665 3.065 7.965 3.39 ;
      RECT 6.9 4.155 7.23 4.485 ;
      RECT 4.86 4.155 5.19 4.485 ;
      RECT 4.86 4.17 7.23 4.47 ;
      RECT 6.55 3.415 6.88 3.745 ;
      RECT 6.09 3.43 6.89 3.73 ;
      RECT 6.22 2.225 6.55 2.555 ;
      RECT 5.75 2.24 6.55 2.54 ;
      RECT 6.21 2.235 6.55 2.54 ;
    LAYER via2 ;
      RECT 77.215 5.855 77.415 6.055 ;
      RECT 76.865 3.82 77.065 4.02 ;
      RECT 76.525 3.14 76.725 3.34 ;
      RECT 76.175 5.855 76.375 6.055 ;
      RECT 75.845 4.22 76.045 4.42 ;
      RECT 75.495 3.48 75.695 3.68 ;
      RECT 75.165 2.29 75.365 2.49 ;
      RECT 75.165 6.545 75.365 6.745 ;
      RECT 73.805 4.22 74.005 4.42 ;
      RECT 70.45 7.085 70.65 7.285 ;
      RECT 59.995 5.855 60.195 6.055 ;
      RECT 59.645 3.82 59.845 4.02 ;
      RECT 59.305 3.14 59.505 3.34 ;
      RECT 58.955 5.855 59.155 6.055 ;
      RECT 58.625 4.22 58.825 4.42 ;
      RECT 58.275 3.48 58.475 3.68 ;
      RECT 57.945 2.29 58.145 2.49 ;
      RECT 57.945 6.545 58.145 6.745 ;
      RECT 56.585 4.22 56.785 4.42 ;
      RECT 53.23 7.085 53.43 7.285 ;
      RECT 42.775 5.855 42.975 6.055 ;
      RECT 42.425 3.82 42.625 4.02 ;
      RECT 42.085 3.14 42.285 3.34 ;
      RECT 41.735 5.855 41.935 6.055 ;
      RECT 41.405 4.22 41.605 4.42 ;
      RECT 41.055 3.48 41.255 3.68 ;
      RECT 40.725 2.29 40.925 2.49 ;
      RECT 40.725 6.545 40.925 6.745 ;
      RECT 39.365 4.22 39.565 4.42 ;
      RECT 36.01 7.085 36.21 7.285 ;
      RECT 25.555 5.855 25.755 6.055 ;
      RECT 25.205 3.82 25.405 4.02 ;
      RECT 24.865 3.14 25.065 3.34 ;
      RECT 24.515 5.855 24.715 6.055 ;
      RECT 24.185 4.22 24.385 4.42 ;
      RECT 23.835 3.48 24.035 3.68 ;
      RECT 23.505 2.29 23.705 2.49 ;
      RECT 23.505 6.545 23.705 6.745 ;
      RECT 22.145 4.22 22.345 4.42 ;
      RECT 18.79 7.085 18.99 7.285 ;
      RECT 8.335 5.855 8.535 6.055 ;
      RECT 7.985 3.82 8.185 4.02 ;
      RECT 7.645 3.14 7.845 3.34 ;
      RECT 7.295 5.855 7.495 6.055 ;
      RECT 6.965 4.22 7.165 4.42 ;
      RECT 6.615 3.48 6.815 3.68 ;
      RECT 6.285 2.29 6.485 2.49 ;
      RECT 6.285 6.545 6.485 6.745 ;
      RECT 4.925 4.22 5.125 4.42 ;
      RECT 1.57 7.085 1.77 7.285 ;
    LAYER met2 ;
      RECT -2.21 8.6 85.1 8.77 ;
      RECT 84.93 7.3 85.1 8.77 ;
      RECT -2.21 6.255 -2.04 8.77 ;
      RECT 84.895 7.3 85.22 7.625 ;
      RECT -2.265 6.255 -1.985 6.595 ;
      RECT 81.74 6.28 82.06 6.605 ;
      RECT 81.77 5.695 81.94 6.605 ;
      RECT 81.77 5.695 81.945 6.045 ;
      RECT 81.77 5.695 82.745 5.87 ;
      RECT 82.57 1.965 82.745 5.87 ;
      RECT 76.485 3.055 76.765 3.425 ;
      RECT 76.555 2.345 76.73 3.425 ;
      RECT 76.555 2.345 79.775 2.52 ;
      RECT 79.6 2.025 79.775 2.52 ;
      RECT 80.07 1.995 80.395 2.32 ;
      RECT 82.515 1.965 82.865 2.315 ;
      RECT 79.6 2.025 82.865 2.195 ;
      RECT 70.89 8.29 81.585 8.46 ;
      RECT 81.425 2.395 81.585 8.46 ;
      RECT 70.89 6.545 71.06 8.46 ;
      RECT 82.54 6.655 82.865 6.98 ;
      RECT 67.71 6.655 68.035 6.98 ;
      RECT 81.425 6.745 82.865 6.915 ;
      RECT 70.84 6.545 71.12 6.885 ;
      RECT 67.71 6.685 71.12 6.855 ;
      RECT 81.74 2.365 82.06 2.685 ;
      RECT 81.425 2.395 82.06 2.565 ;
      RECT 78.195 6.48 78.455 6.8 ;
      RECT 78.255 2.74 78.395 6.8 ;
      RECT 78.195 2.74 78.455 3.06 ;
      RECT 77.515 4.78 77.775 5.1 ;
      RECT 77.575 3.76 77.715 5.1 ;
      RECT 77.515 3.76 77.775 4.08 ;
      RECT 76.495 6.48 76.755 6.8 ;
      RECT 76.555 5.21 76.695 6.8 ;
      RECT 75.875 5.21 76.695 5.35 ;
      RECT 75.875 2.74 76.015 5.35 ;
      RECT 75.805 4.135 76.085 4.505 ;
      RECT 75.815 2.74 76.075 3.06 ;
      RECT 73.765 4.135 74.045 4.505 ;
      RECT 73.835 2.4 73.975 4.505 ;
      RECT 73.775 2.4 74.035 2.72 ;
      RECT 73.095 4.78 73.355 5.1 ;
      RECT 73.155 2.74 73.295 5.1 ;
      RECT 73.095 2.74 73.355 3.06 ;
      RECT 64.52 6.28 64.84 6.605 ;
      RECT 64.55 5.695 64.72 6.605 ;
      RECT 64.55 5.695 64.725 6.045 ;
      RECT 64.55 5.695 65.525 5.87 ;
      RECT 65.35 1.965 65.525 5.87 ;
      RECT 59.265 3.055 59.545 3.425 ;
      RECT 59.335 2.345 59.51 3.425 ;
      RECT 59.335 2.345 62.555 2.52 ;
      RECT 62.38 2.025 62.555 2.52 ;
      RECT 62.85 1.995 63.175 2.32 ;
      RECT 65.295 1.965 65.645 2.315 ;
      RECT 62.38 2.025 65.645 2.195 ;
      RECT 53.67 8.29 64.365 8.46 ;
      RECT 64.205 2.395 64.365 8.46 ;
      RECT 53.67 6.545 53.84 8.46 ;
      RECT 65.32 6.655 65.645 6.98 ;
      RECT 50.49 6.655 50.815 6.98 ;
      RECT 64.205 6.745 65.645 6.915 ;
      RECT 53.62 6.545 53.9 6.885 ;
      RECT 50.49 6.685 53.9 6.855 ;
      RECT 64.52 2.365 64.84 2.685 ;
      RECT 64.205 2.395 64.84 2.565 ;
      RECT 60.975 6.48 61.235 6.8 ;
      RECT 61.035 2.74 61.175 6.8 ;
      RECT 60.975 2.74 61.235 3.06 ;
      RECT 60.295 4.78 60.555 5.1 ;
      RECT 60.355 3.76 60.495 5.1 ;
      RECT 60.295 3.76 60.555 4.08 ;
      RECT 59.275 6.48 59.535 6.8 ;
      RECT 59.335 5.21 59.475 6.8 ;
      RECT 58.655 5.21 59.475 5.35 ;
      RECT 58.655 2.74 58.795 5.35 ;
      RECT 58.585 4.135 58.865 4.505 ;
      RECT 58.595 2.74 58.855 3.06 ;
      RECT 56.545 4.135 56.825 4.505 ;
      RECT 56.615 2.4 56.755 4.505 ;
      RECT 56.555 2.4 56.815 2.72 ;
      RECT 55.875 4.78 56.135 5.1 ;
      RECT 55.935 2.74 56.075 5.1 ;
      RECT 55.875 2.74 56.135 3.06 ;
      RECT 47.3 6.28 47.62 6.605 ;
      RECT 47.33 5.695 47.5 6.605 ;
      RECT 47.33 5.695 47.505 6.045 ;
      RECT 47.33 5.695 48.305 5.87 ;
      RECT 48.13 1.965 48.305 5.87 ;
      RECT 42.045 3.055 42.325 3.425 ;
      RECT 42.115 2.345 42.29 3.425 ;
      RECT 42.115 2.345 45.335 2.52 ;
      RECT 45.16 2.025 45.335 2.52 ;
      RECT 45.63 1.995 45.955 2.32 ;
      RECT 48.075 1.965 48.425 2.315 ;
      RECT 45.16 2.025 48.425 2.195 ;
      RECT 36.45 8.29 47.145 8.46 ;
      RECT 46.985 2.395 47.145 8.46 ;
      RECT 36.45 6.545 36.62 8.46 ;
      RECT 48.1 6.655 48.425 6.98 ;
      RECT 33.27 6.655 33.595 6.98 ;
      RECT 46.985 6.745 48.425 6.915 ;
      RECT 36.4 6.545 36.68 6.885 ;
      RECT 33.27 6.685 36.69 6.855 ;
      RECT 47.3 2.365 47.62 2.685 ;
      RECT 46.985 2.395 47.62 2.565 ;
      RECT 43.755 6.48 44.015 6.8 ;
      RECT 43.815 2.74 43.955 6.8 ;
      RECT 43.755 2.74 44.015 3.06 ;
      RECT 43.075 4.78 43.335 5.1 ;
      RECT 43.135 3.76 43.275 5.1 ;
      RECT 43.075 3.76 43.335 4.08 ;
      RECT 42.055 6.48 42.315 6.8 ;
      RECT 42.115 5.21 42.255 6.8 ;
      RECT 41.435 5.21 42.255 5.35 ;
      RECT 41.435 2.74 41.575 5.35 ;
      RECT 41.365 4.135 41.645 4.505 ;
      RECT 41.375 2.74 41.635 3.06 ;
      RECT 39.325 4.135 39.605 4.505 ;
      RECT 39.395 2.4 39.535 4.505 ;
      RECT 39.335 2.4 39.595 2.72 ;
      RECT 38.655 4.78 38.915 5.1 ;
      RECT 38.715 2.74 38.855 5.1 ;
      RECT 38.655 2.74 38.915 3.06 ;
      RECT 30.08 6.28 30.4 6.605 ;
      RECT 30.11 5.695 30.28 6.605 ;
      RECT 30.11 5.695 30.285 6.045 ;
      RECT 30.11 5.695 31.085 5.87 ;
      RECT 30.91 1.965 31.085 5.87 ;
      RECT 24.825 3.055 25.105 3.425 ;
      RECT 24.895 2.345 25.07 3.425 ;
      RECT 24.895 2.345 28.115 2.52 ;
      RECT 27.94 2.025 28.115 2.52 ;
      RECT 28.41 1.995 28.735 2.32 ;
      RECT 30.855 1.965 31.205 2.315 ;
      RECT 27.94 2.025 31.205 2.195 ;
      RECT 19.23 8.29 29.925 8.46 ;
      RECT 29.765 2.395 29.925 8.46 ;
      RECT 19.23 6.545 19.4 8.46 ;
      RECT 30.88 6.655 31.205 6.98 ;
      RECT 16.05 6.655 16.375 6.98 ;
      RECT 29.765 6.745 31.205 6.915 ;
      RECT 19.18 6.545 19.46 6.885 ;
      RECT 16.05 6.685 19.46 6.855 ;
      RECT 30.08 2.365 30.4 2.685 ;
      RECT 29.765 2.395 30.4 2.565 ;
      RECT 26.535 6.48 26.795 6.8 ;
      RECT 26.595 2.74 26.735 6.8 ;
      RECT 26.535 2.74 26.795 3.06 ;
      RECT 25.855 4.78 26.115 5.1 ;
      RECT 25.915 3.76 26.055 5.1 ;
      RECT 25.855 3.76 26.115 4.08 ;
      RECT 24.835 6.48 25.095 6.8 ;
      RECT 24.895 5.21 25.035 6.8 ;
      RECT 24.215 5.21 25.035 5.35 ;
      RECT 24.215 2.74 24.355 5.35 ;
      RECT 24.145 4.135 24.425 4.505 ;
      RECT 24.155 2.74 24.415 3.06 ;
      RECT 22.105 4.135 22.385 4.505 ;
      RECT 22.175 2.4 22.315 4.505 ;
      RECT 22.115 2.4 22.375 2.72 ;
      RECT 21.435 4.78 21.695 5.1 ;
      RECT 21.495 2.74 21.635 5.1 ;
      RECT 21.435 2.74 21.695 3.06 ;
      RECT 12.86 6.28 13.18 6.605 ;
      RECT 12.89 5.695 13.06 6.605 ;
      RECT 12.89 5.695 13.065 6.045 ;
      RECT 12.89 5.695 13.865 5.87 ;
      RECT 13.69 1.965 13.865 5.87 ;
      RECT 7.605 3.055 7.885 3.425 ;
      RECT 7.675 2.345 7.85 3.425 ;
      RECT 7.675 2.345 10.895 2.52 ;
      RECT 10.72 2.025 10.895 2.52 ;
      RECT 11.19 1.995 11.515 2.32 ;
      RECT 13.635 1.965 13.985 2.315 ;
      RECT 10.72 2.025 13.985 2.195 ;
      RECT 2.01 8.29 12.705 8.46 ;
      RECT 12.545 2.395 12.705 8.46 ;
      RECT 2.01 6.545 2.18 8.46 ;
      RECT -1.89 6.995 -1.61 7.335 ;
      RECT -1.89 7.06 -0.68 7.23 ;
      RECT -0.85 6.685 -0.68 7.23 ;
      RECT 13.66 6.655 13.985 6.98 ;
      RECT 12.545 6.745 13.985 6.915 ;
      RECT 1.96 6.545 2.24 6.885 ;
      RECT -0.85 6.685 2.24 6.855 ;
      RECT 12.86 2.365 13.18 2.685 ;
      RECT 12.545 2.395 13.18 2.565 ;
      RECT 9.315 6.48 9.575 6.8 ;
      RECT 9.375 2.74 9.515 6.8 ;
      RECT 9.315 2.74 9.575 3.06 ;
      RECT 8.635 4.78 8.895 5.1 ;
      RECT 8.695 3.76 8.835 5.1 ;
      RECT 8.635 3.76 8.895 4.08 ;
      RECT 7.615 6.48 7.875 6.8 ;
      RECT 7.675 5.21 7.815 6.8 ;
      RECT 6.995 5.21 7.815 5.35 ;
      RECT 6.995 2.74 7.135 5.35 ;
      RECT 6.925 4.135 7.205 4.505 ;
      RECT 6.935 2.74 7.195 3.06 ;
      RECT 4.885 4.135 5.165 4.505 ;
      RECT 4.955 2.4 5.095 4.505 ;
      RECT 4.895 2.4 5.155 2.72 ;
      RECT 4.215 4.78 4.475 5.1 ;
      RECT 4.275 2.74 4.415 5.1 ;
      RECT 4.215 2.74 4.475 3.06 ;
      RECT 77.175 5.77 77.455 6.14 ;
      RECT 76.825 3.735 77.105 4.105 ;
      RECT 76.135 5.77 76.415 6.14 ;
      RECT 75.455 3.395 75.735 3.765 ;
      RECT 75.125 2.205 75.405 2.575 ;
      RECT 75.125 6.46 75.405 6.83 ;
      RECT 70.365 7 70.735 7.37 ;
      RECT 59.955 5.77 60.235 6.14 ;
      RECT 59.605 3.735 59.885 4.105 ;
      RECT 58.915 5.77 59.195 6.14 ;
      RECT 58.235 3.395 58.515 3.765 ;
      RECT 57.905 2.205 58.185 2.575 ;
      RECT 57.905 6.46 58.185 6.83 ;
      RECT 53.145 7 53.515 7.37 ;
      RECT 42.735 5.77 43.015 6.14 ;
      RECT 42.385 3.735 42.665 4.105 ;
      RECT 41.695 5.77 41.975 6.14 ;
      RECT 41.015 3.395 41.295 3.765 ;
      RECT 40.685 2.205 40.965 2.575 ;
      RECT 40.685 6.46 40.965 6.83 ;
      RECT 35.925 7 36.295 7.37 ;
      RECT 25.515 5.77 25.795 6.14 ;
      RECT 25.165 3.735 25.445 4.105 ;
      RECT 24.475 5.77 24.755 6.14 ;
      RECT 23.795 3.395 24.075 3.765 ;
      RECT 23.465 2.205 23.745 2.575 ;
      RECT 23.465 6.46 23.745 6.83 ;
      RECT 18.705 7 19.075 7.37 ;
      RECT 8.295 5.77 8.575 6.14 ;
      RECT 7.945 3.735 8.225 4.105 ;
      RECT 7.255 5.77 7.535 6.14 ;
      RECT 6.575 3.395 6.855 3.765 ;
      RECT 6.245 2.205 6.525 2.575 ;
      RECT 6.245 6.46 6.525 6.83 ;
      RECT 1.485 7 1.855 7.37 ;
    LAYER via1 ;
      RECT 84.985 7.385 85.135 7.535 ;
      RECT 82.63 6.74 82.78 6.89 ;
      RECT 82.615 2.065 82.765 2.215 ;
      RECT 81.825 2.45 81.975 2.6 ;
      RECT 81.825 6.37 81.975 6.52 ;
      RECT 80.16 2.08 80.31 2.23 ;
      RECT 78.25 2.825 78.4 2.975 ;
      RECT 78.25 6.565 78.4 6.715 ;
      RECT 77.57 3.845 77.72 3.995 ;
      RECT 77.57 4.865 77.72 5.015 ;
      RECT 77.23 5.885 77.38 6.035 ;
      RECT 76.89 3.845 77.04 3.995 ;
      RECT 76.55 3.165 76.7 3.315 ;
      RECT 76.55 6.565 76.7 6.715 ;
      RECT 76.2 5.885 76.35 6.035 ;
      RECT 75.87 2.825 76.02 2.975 ;
      RECT 75.53 3.505 75.68 3.655 ;
      RECT 75.19 2.315 75.34 2.465 ;
      RECT 75.19 6.565 75.34 6.715 ;
      RECT 73.83 2.485 73.98 2.635 ;
      RECT 73.15 2.825 73.3 2.975 ;
      RECT 73.15 4.865 73.3 5.015 ;
      RECT 70.905 6.64 71.055 6.79 ;
      RECT 70.475 7.11 70.625 7.26 ;
      RECT 67.8 6.74 67.95 6.89 ;
      RECT 65.41 6.74 65.56 6.89 ;
      RECT 65.395 2.065 65.545 2.215 ;
      RECT 64.605 2.45 64.755 2.6 ;
      RECT 64.605 6.37 64.755 6.52 ;
      RECT 62.94 2.08 63.09 2.23 ;
      RECT 61.03 2.825 61.18 2.975 ;
      RECT 61.03 6.565 61.18 6.715 ;
      RECT 60.35 3.845 60.5 3.995 ;
      RECT 60.35 4.865 60.5 5.015 ;
      RECT 60.01 5.885 60.16 6.035 ;
      RECT 59.67 3.845 59.82 3.995 ;
      RECT 59.33 3.165 59.48 3.315 ;
      RECT 59.33 6.565 59.48 6.715 ;
      RECT 58.98 5.885 59.13 6.035 ;
      RECT 58.65 2.825 58.8 2.975 ;
      RECT 58.31 3.505 58.46 3.655 ;
      RECT 57.97 2.315 58.12 2.465 ;
      RECT 57.97 6.565 58.12 6.715 ;
      RECT 56.61 2.485 56.76 2.635 ;
      RECT 55.93 2.825 56.08 2.975 ;
      RECT 55.93 4.865 56.08 5.015 ;
      RECT 53.685 6.64 53.835 6.79 ;
      RECT 53.255 7.11 53.405 7.26 ;
      RECT 50.58 6.74 50.73 6.89 ;
      RECT 48.19 6.74 48.34 6.89 ;
      RECT 48.175 2.065 48.325 2.215 ;
      RECT 47.385 2.45 47.535 2.6 ;
      RECT 47.385 6.37 47.535 6.52 ;
      RECT 45.72 2.08 45.87 2.23 ;
      RECT 43.81 2.825 43.96 2.975 ;
      RECT 43.81 6.565 43.96 6.715 ;
      RECT 43.13 3.845 43.28 3.995 ;
      RECT 43.13 4.865 43.28 5.015 ;
      RECT 42.79 5.885 42.94 6.035 ;
      RECT 42.45 3.845 42.6 3.995 ;
      RECT 42.11 3.165 42.26 3.315 ;
      RECT 42.11 6.565 42.26 6.715 ;
      RECT 41.76 5.885 41.91 6.035 ;
      RECT 41.43 2.825 41.58 2.975 ;
      RECT 41.09 3.505 41.24 3.655 ;
      RECT 40.75 2.315 40.9 2.465 ;
      RECT 40.75 6.565 40.9 6.715 ;
      RECT 39.39 2.485 39.54 2.635 ;
      RECT 38.71 2.825 38.86 2.975 ;
      RECT 38.71 4.865 38.86 5.015 ;
      RECT 36.465 6.64 36.615 6.79 ;
      RECT 36.035 7.11 36.185 7.26 ;
      RECT 33.36 6.74 33.51 6.89 ;
      RECT 30.97 6.74 31.12 6.89 ;
      RECT 30.955 2.065 31.105 2.215 ;
      RECT 30.165 2.45 30.315 2.6 ;
      RECT 30.165 6.37 30.315 6.52 ;
      RECT 28.5 2.08 28.65 2.23 ;
      RECT 26.59 2.825 26.74 2.975 ;
      RECT 26.59 6.565 26.74 6.715 ;
      RECT 25.91 3.845 26.06 3.995 ;
      RECT 25.91 4.865 26.06 5.015 ;
      RECT 25.57 5.885 25.72 6.035 ;
      RECT 25.23 3.845 25.38 3.995 ;
      RECT 24.89 3.165 25.04 3.315 ;
      RECT 24.89 6.565 25.04 6.715 ;
      RECT 24.54 5.885 24.69 6.035 ;
      RECT 24.21 2.825 24.36 2.975 ;
      RECT 23.87 3.505 24.02 3.655 ;
      RECT 23.53 2.315 23.68 2.465 ;
      RECT 23.53 6.565 23.68 6.715 ;
      RECT 22.17 2.485 22.32 2.635 ;
      RECT 21.49 2.825 21.64 2.975 ;
      RECT 21.49 4.865 21.64 5.015 ;
      RECT 19.245 6.64 19.395 6.79 ;
      RECT 18.815 7.11 18.965 7.26 ;
      RECT 16.14 6.74 16.29 6.89 ;
      RECT 13.75 6.74 13.9 6.89 ;
      RECT 13.735 2.065 13.885 2.215 ;
      RECT 12.945 2.45 13.095 2.6 ;
      RECT 12.945 6.37 13.095 6.52 ;
      RECT 11.28 2.08 11.43 2.23 ;
      RECT 9.37 2.825 9.52 2.975 ;
      RECT 9.37 6.565 9.52 6.715 ;
      RECT 8.69 3.845 8.84 3.995 ;
      RECT 8.69 4.865 8.84 5.015 ;
      RECT 8.35 5.885 8.5 6.035 ;
      RECT 8.01 3.845 8.16 3.995 ;
      RECT 7.67 3.165 7.82 3.315 ;
      RECT 7.67 6.565 7.82 6.715 ;
      RECT 7.32 5.885 7.47 6.035 ;
      RECT 6.99 2.825 7.14 2.975 ;
      RECT 6.65 3.505 6.8 3.655 ;
      RECT 6.31 2.315 6.46 2.465 ;
      RECT 6.31 6.565 6.46 6.715 ;
      RECT 4.95 2.485 5.1 2.635 ;
      RECT 4.27 2.825 4.42 2.975 ;
      RECT 4.27 4.865 4.42 5.015 ;
      RECT 2.025 6.64 2.175 6.79 ;
      RECT 1.595 7.11 1.745 7.26 ;
      RECT -1.825 7.09 -1.675 7.24 ;
      RECT -2.2 6.35 -2.05 6.5 ;
    LAYER met1 ;
      RECT 84.865 7.77 85.155 8 ;
      RECT 84.925 6.29 85.095 8 ;
      RECT 84.895 7.3 85.22 7.625 ;
      RECT 84.865 6.29 85.155 6.52 ;
      RECT 84.46 2.395 84.565 2.965 ;
      RECT 84.46 2.73 84.785 2.96 ;
      RECT 84.46 2.76 84.955 2.93 ;
      RECT 84.46 2.395 84.65 2.96 ;
      RECT 83.875 2.36 84.165 2.59 ;
      RECT 83.875 2.395 84.65 2.565 ;
      RECT 83.935 0.88 84.105 2.59 ;
      RECT 83.875 0.88 84.165 1.11 ;
      RECT 83.875 7.77 84.165 8 ;
      RECT 83.935 6.29 84.105 8 ;
      RECT 83.875 6.29 84.165 6.52 ;
      RECT 83.875 6.325 84.73 6.485 ;
      RECT 84.56 5.92 84.73 6.485 ;
      RECT 83.875 6.32 84.27 6.485 ;
      RECT 84.495 5.92 84.785 6.15 ;
      RECT 84.495 5.95 84.955 6.12 ;
      RECT 83.505 2.73 83.795 2.96 ;
      RECT 83.505 2.76 83.965 2.93 ;
      RECT 83.57 1.655 83.735 2.96 ;
      RECT 82.085 1.625 82.375 1.855 ;
      RECT 82.085 1.655 83.735 1.825 ;
      RECT 82.145 0.885 82.315 1.855 ;
      RECT 82.085 0.885 82.375 1.115 ;
      RECT 82.085 7.765 82.375 7.995 ;
      RECT 82.145 7.025 82.315 7.995 ;
      RECT 82.145 7.12 83.735 7.29 ;
      RECT 83.565 5.92 83.735 7.29 ;
      RECT 82.085 7.025 82.375 7.255 ;
      RECT 83.505 5.92 83.795 6.15 ;
      RECT 83.505 5.95 83.965 6.12 ;
      RECT 82.515 1.965 82.865 2.315 ;
      RECT 82.345 2.025 82.865 2.195 ;
      RECT 82.54 6.655 82.865 6.98 ;
      RECT 82.515 6.655 82.865 6.885 ;
      RECT 82.345 6.685 82.865 6.855 ;
      RECT 81.74 2.365 82.06 2.685 ;
      RECT 81.71 2.365 82.06 2.595 ;
      RECT 81.425 2.395 82.06 2.565 ;
      RECT 81.74 6.28 82.06 6.605 ;
      RECT 81.71 6.285 82.06 6.515 ;
      RECT 81.54 6.315 82.06 6.485 ;
      RECT 77.485 3.79 77.805 4.05 ;
      RECT 78.52 3.805 78.81 4.035 ;
      RECT 77.485 3.85 78.81 3.99 ;
      RECT 77.145 5.83 77.465 6.09 ;
      RECT 78.52 5.845 78.81 6.075 ;
      RECT 78.595 5.55 78.735 6.075 ;
      RECT 77.235 5.55 77.375 6.09 ;
      RECT 77.235 5.55 78.735 5.69 ;
      RECT 78.165 2.77 78.485 3.03 ;
      RECT 77.89 2.83 78.485 2.97 ;
      RECT 75.105 6.51 75.425 6.77 ;
      RECT 74.1 6.525 74.39 6.755 ;
      RECT 74.1 6.57 76.015 6.71 ;
      RECT 75.875 6.23 76.015 6.71 ;
      RECT 75.875 6.23 77.885 6.37 ;
      RECT 77.745 5.845 77.885 6.37 ;
      RECT 77.67 5.845 77.96 6.075 ;
      RECT 77.485 4.81 77.805 5.07 ;
      RECT 75.34 4.825 75.63 5.055 ;
      RECT 75.34 4.87 77.805 5.01 ;
      RECT 76.805 3.79 77.125 4.05 ;
      RECT 74.44 3.805 74.73 4.035 ;
      RECT 74.44 3.85 77.125 3.99 ;
      RECT 76.465 6.51 76.785 6.77 ;
      RECT 76.465 6.57 77.06 6.71 ;
      RECT 76.465 3.11 76.785 3.37 ;
      RECT 76.19 3.17 76.785 3.31 ;
      RECT 75.785 2.77 76.105 3.03 ;
      RECT 75.51 2.83 76.105 2.97 ;
      RECT 75.445 3.45 75.765 3.71 ;
      RECT 72.57 3.465 72.86 3.695 ;
      RECT 72.57 3.51 75.765 3.65 ;
      RECT 75.025 2.79 75.165 3.65 ;
      RECT 74.95 2.79 75.24 3.02 ;
      RECT 75.105 2.26 75.425 2.52 ;
      RECT 75.105 2.275 75.61 2.505 ;
      RECT 75.015 2.32 75.61 2.46 ;
      RECT 74.44 2.79 74.73 3.02 ;
      RECT 73.835 2.835 74.73 2.975 ;
      RECT 73.835 2.43 73.975 2.975 ;
      RECT 73.745 2.43 74.065 2.69 ;
      RECT 73.065 2.77 73.385 3.03 ;
      RECT 72.79 2.83 73.385 2.97 ;
      RECT 73.065 4.81 73.385 5.07 ;
      RECT 72.79 4.87 73.385 5.01 ;
      RECT 70.83 6.575 71.12 6.885 ;
      RECT 70.66 6.685 71.15 6.855 ;
      RECT 70.81 6.575 71.15 6.855 ;
      RECT 70.4 7.765 70.69 7.995 ;
      RECT 70.46 6.995 70.63 7.995 ;
      RECT 70.365 6.995 70.735 7.37 ;
      RECT 67.645 7.77 67.935 8 ;
      RECT 67.705 6.29 67.875 8 ;
      RECT 67.705 6.655 68.035 6.98 ;
      RECT 67.645 6.29 67.935 6.52 ;
      RECT 67.24 2.395 67.345 2.965 ;
      RECT 67.24 2.73 67.565 2.96 ;
      RECT 67.24 2.76 67.735 2.93 ;
      RECT 67.24 2.395 67.43 2.96 ;
      RECT 66.655 2.36 66.945 2.59 ;
      RECT 66.655 2.395 67.43 2.565 ;
      RECT 66.715 0.88 66.885 2.59 ;
      RECT 66.655 0.88 66.945 1.11 ;
      RECT 66.655 7.77 66.945 8 ;
      RECT 66.715 6.29 66.885 8 ;
      RECT 66.655 6.29 66.945 6.52 ;
      RECT 66.655 6.325 67.51 6.485 ;
      RECT 67.34 5.92 67.51 6.485 ;
      RECT 66.655 6.32 67.05 6.485 ;
      RECT 67.275 5.92 67.565 6.15 ;
      RECT 67.275 5.95 67.735 6.12 ;
      RECT 66.285 2.73 66.575 2.96 ;
      RECT 66.285 2.76 66.745 2.93 ;
      RECT 66.35 1.655 66.515 2.96 ;
      RECT 64.865 1.625 65.155 1.855 ;
      RECT 64.865 1.655 66.515 1.825 ;
      RECT 64.925 0.885 65.095 1.855 ;
      RECT 64.865 0.885 65.155 1.115 ;
      RECT 64.865 7.765 65.155 7.995 ;
      RECT 64.925 7.025 65.095 7.995 ;
      RECT 64.925 7.12 66.515 7.29 ;
      RECT 66.345 5.92 66.515 7.29 ;
      RECT 64.865 7.025 65.155 7.255 ;
      RECT 66.285 5.92 66.575 6.15 ;
      RECT 66.285 5.95 66.745 6.12 ;
      RECT 65.295 1.965 65.645 2.315 ;
      RECT 65.125 2.025 65.645 2.195 ;
      RECT 65.32 6.655 65.645 6.98 ;
      RECT 65.295 6.655 65.645 6.885 ;
      RECT 65.125 6.685 65.645 6.855 ;
      RECT 64.52 2.365 64.84 2.685 ;
      RECT 64.49 2.365 64.84 2.595 ;
      RECT 64.205 2.395 64.84 2.565 ;
      RECT 64.52 6.28 64.84 6.605 ;
      RECT 64.49 6.285 64.84 6.515 ;
      RECT 64.32 6.315 64.84 6.485 ;
      RECT 60.265 3.79 60.585 4.05 ;
      RECT 61.3 3.805 61.59 4.035 ;
      RECT 60.265 3.85 61.59 3.99 ;
      RECT 59.925 5.83 60.245 6.09 ;
      RECT 61.3 5.845 61.59 6.075 ;
      RECT 61.375 5.55 61.515 6.075 ;
      RECT 60.015 5.55 60.155 6.09 ;
      RECT 60.015 5.55 61.515 5.69 ;
      RECT 60.945 2.77 61.265 3.03 ;
      RECT 60.67 2.83 61.265 2.97 ;
      RECT 57.885 6.51 58.205 6.77 ;
      RECT 56.88 6.525 57.17 6.755 ;
      RECT 56.88 6.57 58.795 6.71 ;
      RECT 58.655 6.23 58.795 6.71 ;
      RECT 58.655 6.23 60.665 6.37 ;
      RECT 60.525 5.845 60.665 6.37 ;
      RECT 60.45 5.845 60.74 6.075 ;
      RECT 60.265 4.81 60.585 5.07 ;
      RECT 58.12 4.825 58.41 5.055 ;
      RECT 58.12 4.87 60.585 5.01 ;
      RECT 59.585 3.79 59.905 4.05 ;
      RECT 57.22 3.805 57.51 4.035 ;
      RECT 57.22 3.85 59.905 3.99 ;
      RECT 59.245 6.51 59.565 6.77 ;
      RECT 59.245 6.57 59.84 6.71 ;
      RECT 59.245 3.11 59.565 3.37 ;
      RECT 58.97 3.17 59.565 3.31 ;
      RECT 58.565 2.77 58.885 3.03 ;
      RECT 58.29 2.83 58.885 2.97 ;
      RECT 58.225 3.45 58.545 3.71 ;
      RECT 55.35 3.465 55.64 3.695 ;
      RECT 55.35 3.51 58.545 3.65 ;
      RECT 57.805 2.79 57.945 3.65 ;
      RECT 57.73 2.79 58.02 3.02 ;
      RECT 57.885 2.26 58.205 2.52 ;
      RECT 57.885 2.275 58.39 2.505 ;
      RECT 57.795 2.32 58.39 2.46 ;
      RECT 57.22 2.79 57.51 3.02 ;
      RECT 56.615 2.835 57.51 2.975 ;
      RECT 56.615 2.43 56.755 2.975 ;
      RECT 56.525 2.43 56.845 2.69 ;
      RECT 55.845 2.77 56.165 3.03 ;
      RECT 55.57 2.83 56.165 2.97 ;
      RECT 55.845 4.81 56.165 5.07 ;
      RECT 55.57 4.87 56.165 5.01 ;
      RECT 53.61 6.575 53.9 6.885 ;
      RECT 53.44 6.685 53.93 6.855 ;
      RECT 53.59 6.575 53.93 6.855 ;
      RECT 53.18 7.765 53.47 7.995 ;
      RECT 53.24 6.995 53.41 7.995 ;
      RECT 53.145 6.995 53.515 7.37 ;
      RECT 50.425 7.77 50.715 8 ;
      RECT 50.485 6.29 50.655 8 ;
      RECT 50.485 6.655 50.815 6.98 ;
      RECT 50.425 6.29 50.715 6.52 ;
      RECT 50.02 2.395 50.125 2.965 ;
      RECT 50.02 2.73 50.345 2.96 ;
      RECT 50.02 2.76 50.515 2.93 ;
      RECT 50.02 2.395 50.21 2.96 ;
      RECT 49.435 2.36 49.725 2.59 ;
      RECT 49.435 2.395 50.21 2.565 ;
      RECT 49.495 0.88 49.665 2.59 ;
      RECT 49.435 0.88 49.725 1.11 ;
      RECT 49.435 7.77 49.725 8 ;
      RECT 49.495 6.29 49.665 8 ;
      RECT 49.435 6.29 49.725 6.52 ;
      RECT 49.435 6.325 50.29 6.485 ;
      RECT 50.12 5.92 50.29 6.485 ;
      RECT 49.435 6.32 49.83 6.485 ;
      RECT 50.055 5.92 50.345 6.15 ;
      RECT 50.055 5.95 50.515 6.12 ;
      RECT 49.065 2.73 49.355 2.96 ;
      RECT 49.065 2.76 49.525 2.93 ;
      RECT 49.13 1.655 49.295 2.96 ;
      RECT 47.645 1.625 47.935 1.855 ;
      RECT 47.645 1.655 49.295 1.825 ;
      RECT 47.705 0.885 47.875 1.855 ;
      RECT 47.645 0.885 47.935 1.115 ;
      RECT 47.645 7.765 47.935 7.995 ;
      RECT 47.705 7.025 47.875 7.995 ;
      RECT 47.705 7.12 49.295 7.29 ;
      RECT 49.125 5.92 49.295 7.29 ;
      RECT 47.645 7.025 47.935 7.255 ;
      RECT 49.065 5.92 49.355 6.15 ;
      RECT 49.065 5.95 49.525 6.12 ;
      RECT 48.075 1.965 48.425 2.315 ;
      RECT 47.905 2.025 48.425 2.195 ;
      RECT 48.1 6.655 48.425 6.98 ;
      RECT 48.075 6.655 48.425 6.885 ;
      RECT 47.905 6.685 48.425 6.855 ;
      RECT 47.3 2.365 47.62 2.685 ;
      RECT 47.27 2.365 47.62 2.595 ;
      RECT 46.985 2.395 47.62 2.565 ;
      RECT 47.3 6.28 47.62 6.605 ;
      RECT 47.27 6.285 47.62 6.515 ;
      RECT 47.1 6.315 47.62 6.485 ;
      RECT 43.045 3.79 43.365 4.05 ;
      RECT 44.08 3.805 44.37 4.035 ;
      RECT 43.045 3.85 44.37 3.99 ;
      RECT 42.705 5.83 43.025 6.09 ;
      RECT 44.08 5.845 44.37 6.075 ;
      RECT 44.155 5.55 44.295 6.075 ;
      RECT 42.795 5.55 42.935 6.09 ;
      RECT 42.795 5.55 44.295 5.69 ;
      RECT 43.725 2.77 44.045 3.03 ;
      RECT 43.45 2.83 44.045 2.97 ;
      RECT 40.665 6.51 40.985 6.77 ;
      RECT 39.66 6.525 39.95 6.755 ;
      RECT 39.66 6.57 41.575 6.71 ;
      RECT 41.435 6.23 41.575 6.71 ;
      RECT 41.435 6.23 43.445 6.37 ;
      RECT 43.305 5.845 43.445 6.37 ;
      RECT 43.23 5.845 43.52 6.075 ;
      RECT 43.045 4.81 43.365 5.07 ;
      RECT 40.9 4.825 41.19 5.055 ;
      RECT 40.9 4.87 43.365 5.01 ;
      RECT 42.365 3.79 42.685 4.05 ;
      RECT 40 3.805 40.29 4.035 ;
      RECT 40 3.85 42.685 3.99 ;
      RECT 42.025 6.51 42.345 6.77 ;
      RECT 42.025 6.57 42.62 6.71 ;
      RECT 42.025 3.11 42.345 3.37 ;
      RECT 41.75 3.17 42.345 3.31 ;
      RECT 41.345 2.77 41.665 3.03 ;
      RECT 41.07 2.83 41.665 2.97 ;
      RECT 41.005 3.45 41.325 3.71 ;
      RECT 38.13 3.465 38.42 3.695 ;
      RECT 38.13 3.51 41.325 3.65 ;
      RECT 40.585 2.79 40.725 3.65 ;
      RECT 40.51 2.79 40.8 3.02 ;
      RECT 40.665 2.26 40.985 2.52 ;
      RECT 40.665 2.275 41.17 2.505 ;
      RECT 40.575 2.32 41.17 2.46 ;
      RECT 40 2.79 40.29 3.02 ;
      RECT 39.395 2.835 40.29 2.975 ;
      RECT 39.395 2.43 39.535 2.975 ;
      RECT 39.305 2.43 39.625 2.69 ;
      RECT 38.625 2.77 38.945 3.03 ;
      RECT 38.35 2.83 38.945 2.97 ;
      RECT 38.625 4.81 38.945 5.07 ;
      RECT 38.35 4.87 38.945 5.01 ;
      RECT 36.39 6.575 36.68 6.885 ;
      RECT 36.22 6.685 36.71 6.855 ;
      RECT 36.37 6.575 36.71 6.855 ;
      RECT 35.96 7.765 36.25 7.995 ;
      RECT 36.02 6.995 36.19 7.995 ;
      RECT 35.925 6.995 36.295 7.37 ;
      RECT 33.205 7.77 33.495 8 ;
      RECT 33.265 6.29 33.435 8 ;
      RECT 33.265 6.655 33.595 6.98 ;
      RECT 33.205 6.29 33.495 6.52 ;
      RECT 32.8 2.395 32.905 2.965 ;
      RECT 32.8 2.73 33.125 2.96 ;
      RECT 32.8 2.76 33.295 2.93 ;
      RECT 32.8 2.395 32.99 2.96 ;
      RECT 32.215 2.36 32.505 2.59 ;
      RECT 32.215 2.395 32.99 2.565 ;
      RECT 32.275 0.88 32.445 2.59 ;
      RECT 32.215 0.88 32.505 1.11 ;
      RECT 32.215 7.77 32.505 8 ;
      RECT 32.275 6.29 32.445 8 ;
      RECT 32.215 6.29 32.505 6.52 ;
      RECT 32.215 6.325 33.07 6.485 ;
      RECT 32.9 5.92 33.07 6.485 ;
      RECT 32.215 6.32 32.61 6.485 ;
      RECT 32.835 5.92 33.125 6.15 ;
      RECT 32.835 5.95 33.295 6.12 ;
      RECT 31.845 2.73 32.135 2.96 ;
      RECT 31.845 2.76 32.305 2.93 ;
      RECT 31.91 1.655 32.075 2.96 ;
      RECT 30.425 1.625 30.715 1.855 ;
      RECT 30.425 1.655 32.075 1.825 ;
      RECT 30.485 0.885 30.655 1.855 ;
      RECT 30.425 0.885 30.715 1.115 ;
      RECT 30.425 7.765 30.715 7.995 ;
      RECT 30.485 7.025 30.655 7.995 ;
      RECT 30.485 7.12 32.075 7.29 ;
      RECT 31.905 5.92 32.075 7.29 ;
      RECT 30.425 7.025 30.715 7.255 ;
      RECT 31.845 5.92 32.135 6.15 ;
      RECT 31.845 5.95 32.305 6.12 ;
      RECT 30.855 1.965 31.205 2.315 ;
      RECT 30.685 2.025 31.205 2.195 ;
      RECT 30.88 6.655 31.205 6.98 ;
      RECT 30.855 6.655 31.205 6.885 ;
      RECT 30.685 6.685 31.205 6.855 ;
      RECT 30.08 2.365 30.4 2.685 ;
      RECT 30.05 2.365 30.4 2.595 ;
      RECT 29.765 2.395 30.4 2.565 ;
      RECT 30.08 6.28 30.4 6.605 ;
      RECT 30.05 6.285 30.4 6.515 ;
      RECT 29.88 6.315 30.4 6.485 ;
      RECT 25.825 3.79 26.145 4.05 ;
      RECT 26.86 3.805 27.15 4.035 ;
      RECT 25.825 3.85 27.15 3.99 ;
      RECT 25.485 5.83 25.805 6.09 ;
      RECT 26.86 5.845 27.15 6.075 ;
      RECT 26.935 5.55 27.075 6.075 ;
      RECT 25.575 5.55 25.715 6.09 ;
      RECT 25.575 5.55 27.075 5.69 ;
      RECT 26.505 2.77 26.825 3.03 ;
      RECT 26.23 2.83 26.825 2.97 ;
      RECT 23.445 6.51 23.765 6.77 ;
      RECT 22.44 6.525 22.73 6.755 ;
      RECT 22.44 6.57 24.355 6.71 ;
      RECT 24.215 6.23 24.355 6.71 ;
      RECT 24.215 6.23 26.225 6.37 ;
      RECT 26.085 5.845 26.225 6.37 ;
      RECT 26.01 5.845 26.3 6.075 ;
      RECT 25.825 4.81 26.145 5.07 ;
      RECT 23.68 4.825 23.97 5.055 ;
      RECT 23.68 4.87 26.145 5.01 ;
      RECT 25.145 3.79 25.465 4.05 ;
      RECT 22.78 3.805 23.07 4.035 ;
      RECT 22.78 3.85 25.465 3.99 ;
      RECT 24.805 6.51 25.125 6.77 ;
      RECT 24.805 6.57 25.4 6.71 ;
      RECT 24.805 3.11 25.125 3.37 ;
      RECT 24.53 3.17 25.125 3.31 ;
      RECT 24.125 2.77 24.445 3.03 ;
      RECT 23.85 2.83 24.445 2.97 ;
      RECT 23.785 3.45 24.105 3.71 ;
      RECT 20.91 3.465 21.2 3.695 ;
      RECT 20.91 3.51 24.105 3.65 ;
      RECT 23.365 2.79 23.505 3.65 ;
      RECT 23.29 2.79 23.58 3.02 ;
      RECT 23.445 2.26 23.765 2.52 ;
      RECT 23.445 2.275 23.95 2.505 ;
      RECT 23.355 2.32 23.95 2.46 ;
      RECT 22.78 2.79 23.07 3.02 ;
      RECT 22.175 2.835 23.07 2.975 ;
      RECT 22.175 2.43 22.315 2.975 ;
      RECT 22.085 2.43 22.405 2.69 ;
      RECT 21.405 2.77 21.725 3.03 ;
      RECT 21.13 2.83 21.725 2.97 ;
      RECT 21.405 4.81 21.725 5.07 ;
      RECT 21.13 4.87 21.725 5.01 ;
      RECT 19.17 6.575 19.46 6.885 ;
      RECT 19 6.685 19.49 6.855 ;
      RECT 19.15 6.575 19.49 6.855 ;
      RECT 18.74 7.765 19.03 7.995 ;
      RECT 18.8 6.995 18.97 7.995 ;
      RECT 18.705 6.995 19.075 7.37 ;
      RECT 15.985 7.77 16.275 8 ;
      RECT 16.045 6.29 16.215 8 ;
      RECT 16.045 6.655 16.375 6.98 ;
      RECT 15.985 6.29 16.275 6.52 ;
      RECT 15.58 2.395 15.685 2.965 ;
      RECT 15.58 2.73 15.905 2.96 ;
      RECT 15.58 2.76 16.075 2.93 ;
      RECT 15.58 2.395 15.77 2.96 ;
      RECT 14.995 2.36 15.285 2.59 ;
      RECT 14.995 2.395 15.77 2.565 ;
      RECT 15.055 0.88 15.225 2.59 ;
      RECT 14.995 0.88 15.285 1.11 ;
      RECT 14.995 7.77 15.285 8 ;
      RECT 15.055 6.29 15.225 8 ;
      RECT 14.995 6.29 15.285 6.52 ;
      RECT 14.995 6.325 15.85 6.485 ;
      RECT 15.68 5.92 15.85 6.485 ;
      RECT 14.995 6.32 15.39 6.485 ;
      RECT 15.615 5.92 15.905 6.15 ;
      RECT 15.615 5.95 16.075 6.12 ;
      RECT 14.625 2.73 14.915 2.96 ;
      RECT 14.625 2.76 15.085 2.93 ;
      RECT 14.69 1.655 14.855 2.96 ;
      RECT 13.205 1.625 13.495 1.855 ;
      RECT 13.205 1.655 14.855 1.825 ;
      RECT 13.265 0.885 13.435 1.855 ;
      RECT 13.205 0.885 13.495 1.115 ;
      RECT 13.205 7.765 13.495 7.995 ;
      RECT 13.265 7.025 13.435 7.995 ;
      RECT 13.265 7.12 14.855 7.29 ;
      RECT 14.685 5.92 14.855 7.29 ;
      RECT 13.205 7.025 13.495 7.255 ;
      RECT 14.625 5.92 14.915 6.15 ;
      RECT 14.625 5.95 15.085 6.12 ;
      RECT 13.635 1.965 13.985 2.315 ;
      RECT 13.465 2.025 13.985 2.195 ;
      RECT 13.66 6.655 13.985 6.98 ;
      RECT 13.635 6.655 13.985 6.885 ;
      RECT 13.465 6.685 13.985 6.855 ;
      RECT 12.86 2.365 13.18 2.685 ;
      RECT 12.83 2.365 13.18 2.595 ;
      RECT 12.545 2.395 13.18 2.565 ;
      RECT 12.86 6.28 13.18 6.605 ;
      RECT 12.83 6.285 13.18 6.515 ;
      RECT 12.66 6.315 13.18 6.485 ;
      RECT 8.605 3.79 8.925 4.05 ;
      RECT 9.64 3.805 9.93 4.035 ;
      RECT 8.605 3.85 9.93 3.99 ;
      RECT 8.265 5.83 8.585 6.09 ;
      RECT 9.64 5.845 9.93 6.075 ;
      RECT 9.715 5.55 9.855 6.075 ;
      RECT 8.355 5.55 8.495 6.09 ;
      RECT 8.355 5.55 9.855 5.69 ;
      RECT 9.285 2.77 9.605 3.03 ;
      RECT 9.01 2.83 9.605 2.97 ;
      RECT 6.225 6.51 6.545 6.77 ;
      RECT 5.22 6.525 5.51 6.755 ;
      RECT 5.22 6.57 7.135 6.71 ;
      RECT 6.995 6.23 7.135 6.71 ;
      RECT 6.995 6.23 9.005 6.37 ;
      RECT 8.865 5.845 9.005 6.37 ;
      RECT 8.79 5.845 9.08 6.075 ;
      RECT 8.605 4.81 8.925 5.07 ;
      RECT 6.46 4.825 6.75 5.055 ;
      RECT 6.46 4.87 8.925 5.01 ;
      RECT 7.925 3.79 8.245 4.05 ;
      RECT 5.56 3.805 5.85 4.035 ;
      RECT 5.56 3.85 8.245 3.99 ;
      RECT 7.585 6.51 7.905 6.77 ;
      RECT 7.585 6.57 8.18 6.71 ;
      RECT 7.585 3.11 7.905 3.37 ;
      RECT 7.31 3.17 7.905 3.31 ;
      RECT 6.905 2.77 7.225 3.03 ;
      RECT 6.63 2.83 7.225 2.97 ;
      RECT 6.565 3.45 6.885 3.71 ;
      RECT 3.69 3.465 3.98 3.695 ;
      RECT 3.69 3.51 6.885 3.65 ;
      RECT 6.145 2.79 6.285 3.65 ;
      RECT 6.07 2.79 6.36 3.02 ;
      RECT 6.225 2.26 6.545 2.52 ;
      RECT 6.225 2.275 6.73 2.505 ;
      RECT 6.135 2.32 6.73 2.46 ;
      RECT 5.56 2.79 5.85 3.02 ;
      RECT 4.955 2.835 5.85 2.975 ;
      RECT 4.955 2.43 5.095 2.975 ;
      RECT 4.865 2.43 5.185 2.69 ;
      RECT 4.185 2.77 4.505 3.03 ;
      RECT 3.91 2.83 4.505 2.97 ;
      RECT 4.185 4.81 4.505 5.07 ;
      RECT 3.91 4.87 4.505 5.01 ;
      RECT 1.95 6.575 2.24 6.885 ;
      RECT 1.78 6.685 2.27 6.855 ;
      RECT 1.93 6.575 2.27 6.855 ;
      RECT 1.52 7.765 1.81 7.995 ;
      RECT 1.58 6.995 1.75 7.995 ;
      RECT 1.485 6.995 1.855 7.37 ;
      RECT -1.89 7.765 -1.6 7.995 ;
      RECT -1.83 7.025 -1.66 7.995 ;
      RECT -1.92 7.025 -1.58 7.305 ;
      RECT -2.295 6.285 -1.955 6.565 ;
      RECT -2.435 6.315 -1.955 6.485 ;
      RECT 80.07 1.995 80.395 2.32 ;
      RECT 77.84 6.51 78.485 6.77 ;
      RECT 75.79 5.83 76.435 6.09 ;
      RECT 62.85 1.995 63.175 2.32 ;
      RECT 60.62 6.51 61.265 6.77 ;
      RECT 58.57 5.83 59.215 6.09 ;
      RECT 45.63 1.995 45.955 2.32 ;
      RECT 43.4 6.51 44.045 6.77 ;
      RECT 41.35 5.83 41.995 6.09 ;
      RECT 28.41 1.995 28.735 2.32 ;
      RECT 26.18 6.51 26.825 6.77 ;
      RECT 24.13 5.83 24.775 6.09 ;
      RECT 11.19 1.995 11.515 2.32 ;
      RECT 8.96 6.51 9.605 6.77 ;
      RECT 6.91 5.83 7.555 6.09 ;
    LAYER mcon ;
      RECT 84.925 6.32 85.095 6.49 ;
      RECT 84.93 6.315 85.1 6.485 ;
      RECT 67.705 6.32 67.875 6.49 ;
      RECT 67.71 6.315 67.88 6.485 ;
      RECT 50.485 6.32 50.655 6.49 ;
      RECT 50.49 6.315 50.66 6.485 ;
      RECT 33.265 6.32 33.435 6.49 ;
      RECT 33.27 6.315 33.44 6.485 ;
      RECT 16.045 6.32 16.215 6.49 ;
      RECT 16.05 6.315 16.22 6.485 ;
      RECT 84.925 7.8 85.095 7.97 ;
      RECT 84.555 2.76 84.725 2.93 ;
      RECT 84.555 5.95 84.725 6.12 ;
      RECT 83.935 0.91 84.105 1.08 ;
      RECT 83.935 2.39 84.105 2.56 ;
      RECT 83.935 6.32 84.105 6.49 ;
      RECT 83.935 7.8 84.105 7.97 ;
      RECT 83.565 2.76 83.735 2.93 ;
      RECT 83.565 5.95 83.735 6.12 ;
      RECT 82.575 2.025 82.745 2.195 ;
      RECT 82.575 6.685 82.745 6.855 ;
      RECT 82.145 0.915 82.315 1.085 ;
      RECT 82.145 1.655 82.315 1.825 ;
      RECT 82.145 7.055 82.315 7.225 ;
      RECT 82.145 7.795 82.315 7.965 ;
      RECT 81.77 2.395 81.94 2.565 ;
      RECT 81.77 6.315 81.94 6.485 ;
      RECT 78.58 3.835 78.75 4.005 ;
      RECT 78.58 5.875 78.75 6.045 ;
      RECT 78.24 2.815 78.41 2.985 ;
      RECT 77.9 6.555 78.07 6.725 ;
      RECT 77.73 5.875 77.9 6.045 ;
      RECT 77.22 5.875 77.39 6.045 ;
      RECT 76.54 3.155 76.71 3.325 ;
      RECT 76.54 6.555 76.71 6.725 ;
      RECT 75.86 2.815 76.03 2.985 ;
      RECT 75.85 5.875 76.02 6.045 ;
      RECT 75.4 4.855 75.57 5.025 ;
      RECT 75.38 2.305 75.55 2.475 ;
      RECT 75.01 2.82 75.18 2.99 ;
      RECT 74.5 2.82 74.67 2.99 ;
      RECT 74.5 3.835 74.67 4.005 ;
      RECT 74.16 6.555 74.33 6.725 ;
      RECT 73.14 2.815 73.31 2.985 ;
      RECT 73.14 4.855 73.31 5.025 ;
      RECT 72.63 3.495 72.8 3.665 ;
      RECT 70.89 6.685 71.06 6.855 ;
      RECT 70.46 7.055 70.63 7.225 ;
      RECT 70.46 7.795 70.63 7.965 ;
      RECT 67.705 7.8 67.875 7.97 ;
      RECT 67.335 2.76 67.505 2.93 ;
      RECT 67.335 5.95 67.505 6.12 ;
      RECT 66.715 0.91 66.885 1.08 ;
      RECT 66.715 2.39 66.885 2.56 ;
      RECT 66.715 6.32 66.885 6.49 ;
      RECT 66.715 7.8 66.885 7.97 ;
      RECT 66.345 2.76 66.515 2.93 ;
      RECT 66.345 5.95 66.515 6.12 ;
      RECT 65.355 2.025 65.525 2.195 ;
      RECT 65.355 6.685 65.525 6.855 ;
      RECT 64.925 0.915 65.095 1.085 ;
      RECT 64.925 1.655 65.095 1.825 ;
      RECT 64.925 7.055 65.095 7.225 ;
      RECT 64.925 7.795 65.095 7.965 ;
      RECT 64.55 2.395 64.72 2.565 ;
      RECT 64.55 6.315 64.72 6.485 ;
      RECT 61.36 3.835 61.53 4.005 ;
      RECT 61.36 5.875 61.53 6.045 ;
      RECT 61.02 2.815 61.19 2.985 ;
      RECT 60.68 6.555 60.85 6.725 ;
      RECT 60.51 5.875 60.68 6.045 ;
      RECT 60 5.875 60.17 6.045 ;
      RECT 59.32 3.155 59.49 3.325 ;
      RECT 59.32 6.555 59.49 6.725 ;
      RECT 58.64 2.815 58.81 2.985 ;
      RECT 58.63 5.875 58.8 6.045 ;
      RECT 58.18 4.855 58.35 5.025 ;
      RECT 58.16 2.305 58.33 2.475 ;
      RECT 57.79 2.82 57.96 2.99 ;
      RECT 57.28 2.82 57.45 2.99 ;
      RECT 57.28 3.835 57.45 4.005 ;
      RECT 56.94 6.555 57.11 6.725 ;
      RECT 55.92 2.815 56.09 2.985 ;
      RECT 55.92 4.855 56.09 5.025 ;
      RECT 55.41 3.495 55.58 3.665 ;
      RECT 53.67 6.685 53.84 6.855 ;
      RECT 53.24 7.055 53.41 7.225 ;
      RECT 53.24 7.795 53.41 7.965 ;
      RECT 50.485 7.8 50.655 7.97 ;
      RECT 50.115 2.76 50.285 2.93 ;
      RECT 50.115 5.95 50.285 6.12 ;
      RECT 49.495 0.91 49.665 1.08 ;
      RECT 49.495 2.39 49.665 2.56 ;
      RECT 49.495 6.32 49.665 6.49 ;
      RECT 49.495 7.8 49.665 7.97 ;
      RECT 49.125 2.76 49.295 2.93 ;
      RECT 49.125 5.95 49.295 6.12 ;
      RECT 48.135 2.025 48.305 2.195 ;
      RECT 48.135 6.685 48.305 6.855 ;
      RECT 47.705 0.915 47.875 1.085 ;
      RECT 47.705 1.655 47.875 1.825 ;
      RECT 47.705 7.055 47.875 7.225 ;
      RECT 47.705 7.795 47.875 7.965 ;
      RECT 47.33 2.395 47.5 2.565 ;
      RECT 47.33 6.315 47.5 6.485 ;
      RECT 44.14 3.835 44.31 4.005 ;
      RECT 44.14 5.875 44.31 6.045 ;
      RECT 43.8 2.815 43.97 2.985 ;
      RECT 43.46 6.555 43.63 6.725 ;
      RECT 43.29 5.875 43.46 6.045 ;
      RECT 42.78 5.875 42.95 6.045 ;
      RECT 42.1 3.155 42.27 3.325 ;
      RECT 42.1 6.555 42.27 6.725 ;
      RECT 41.42 2.815 41.59 2.985 ;
      RECT 41.41 5.875 41.58 6.045 ;
      RECT 40.96 4.855 41.13 5.025 ;
      RECT 40.94 2.305 41.11 2.475 ;
      RECT 40.57 2.82 40.74 2.99 ;
      RECT 40.06 2.82 40.23 2.99 ;
      RECT 40.06 3.835 40.23 4.005 ;
      RECT 39.72 6.555 39.89 6.725 ;
      RECT 38.7 2.815 38.87 2.985 ;
      RECT 38.7 4.855 38.87 5.025 ;
      RECT 38.19 3.495 38.36 3.665 ;
      RECT 36.45 6.685 36.62 6.855 ;
      RECT 36.02 7.055 36.19 7.225 ;
      RECT 36.02 7.795 36.19 7.965 ;
      RECT 33.265 7.8 33.435 7.97 ;
      RECT 32.895 2.76 33.065 2.93 ;
      RECT 32.895 5.95 33.065 6.12 ;
      RECT 32.275 0.91 32.445 1.08 ;
      RECT 32.275 2.39 32.445 2.56 ;
      RECT 32.275 6.32 32.445 6.49 ;
      RECT 32.275 7.8 32.445 7.97 ;
      RECT 31.905 2.76 32.075 2.93 ;
      RECT 31.905 5.95 32.075 6.12 ;
      RECT 30.915 2.025 31.085 2.195 ;
      RECT 30.915 6.685 31.085 6.855 ;
      RECT 30.485 0.915 30.655 1.085 ;
      RECT 30.485 1.655 30.655 1.825 ;
      RECT 30.485 7.055 30.655 7.225 ;
      RECT 30.485 7.795 30.655 7.965 ;
      RECT 30.11 2.395 30.28 2.565 ;
      RECT 30.11 6.315 30.28 6.485 ;
      RECT 26.92 3.835 27.09 4.005 ;
      RECT 26.92 5.875 27.09 6.045 ;
      RECT 26.58 2.815 26.75 2.985 ;
      RECT 26.24 6.555 26.41 6.725 ;
      RECT 26.07 5.875 26.24 6.045 ;
      RECT 25.56 5.875 25.73 6.045 ;
      RECT 24.88 3.155 25.05 3.325 ;
      RECT 24.88 6.555 25.05 6.725 ;
      RECT 24.2 2.815 24.37 2.985 ;
      RECT 24.19 5.875 24.36 6.045 ;
      RECT 23.74 4.855 23.91 5.025 ;
      RECT 23.72 2.305 23.89 2.475 ;
      RECT 23.35 2.82 23.52 2.99 ;
      RECT 22.84 2.82 23.01 2.99 ;
      RECT 22.84 3.835 23.01 4.005 ;
      RECT 22.5 6.555 22.67 6.725 ;
      RECT 21.48 2.815 21.65 2.985 ;
      RECT 21.48 4.855 21.65 5.025 ;
      RECT 20.97 3.495 21.14 3.665 ;
      RECT 19.23 6.685 19.4 6.855 ;
      RECT 18.8 7.055 18.97 7.225 ;
      RECT 18.8 7.795 18.97 7.965 ;
      RECT 16.045 7.8 16.215 7.97 ;
      RECT 15.675 2.76 15.845 2.93 ;
      RECT 15.675 5.95 15.845 6.12 ;
      RECT 15.055 0.91 15.225 1.08 ;
      RECT 15.055 2.39 15.225 2.56 ;
      RECT 15.055 6.32 15.225 6.49 ;
      RECT 15.055 7.8 15.225 7.97 ;
      RECT 14.685 2.76 14.855 2.93 ;
      RECT 14.685 5.95 14.855 6.12 ;
      RECT 13.695 2.025 13.865 2.195 ;
      RECT 13.695 6.685 13.865 6.855 ;
      RECT 13.265 0.915 13.435 1.085 ;
      RECT 13.265 1.655 13.435 1.825 ;
      RECT 13.265 7.055 13.435 7.225 ;
      RECT 13.265 7.795 13.435 7.965 ;
      RECT 12.89 2.395 13.06 2.565 ;
      RECT 12.89 6.315 13.06 6.485 ;
      RECT 9.7 3.835 9.87 4.005 ;
      RECT 9.7 5.875 9.87 6.045 ;
      RECT 9.36 2.815 9.53 2.985 ;
      RECT 9.02 6.555 9.19 6.725 ;
      RECT 8.85 5.875 9.02 6.045 ;
      RECT 8.34 5.875 8.51 6.045 ;
      RECT 7.66 3.155 7.83 3.325 ;
      RECT 7.66 6.555 7.83 6.725 ;
      RECT 6.98 2.815 7.15 2.985 ;
      RECT 6.97 5.875 7.14 6.045 ;
      RECT 6.52 4.855 6.69 5.025 ;
      RECT 6.5 2.305 6.67 2.475 ;
      RECT 6.13 2.82 6.3 2.99 ;
      RECT 5.62 2.82 5.79 2.99 ;
      RECT 5.62 3.835 5.79 4.005 ;
      RECT 5.28 6.555 5.45 6.725 ;
      RECT 4.26 2.815 4.43 2.985 ;
      RECT 4.26 4.855 4.43 5.025 ;
      RECT 3.75 3.495 3.92 3.665 ;
      RECT 2.01 6.685 2.18 6.855 ;
      RECT 1.58 7.055 1.75 7.225 ;
      RECT 1.58 7.795 1.75 7.965 ;
      RECT -1.83 7.055 -1.66 7.225 ;
      RECT -1.83 7.795 -1.66 7.965 ;
      RECT -2.205 6.315 -2.035 6.485 ;
    LAYER li1 ;
      RECT 84.925 5.02 85.095 6.49 ;
      RECT 84.925 6.315 85.1 6.485 ;
      RECT 84.555 1.74 84.725 2.93 ;
      RECT 84.555 1.74 85.025 1.91 ;
      RECT 84.555 6.97 85.025 7.14 ;
      RECT 84.555 5.95 84.725 7.14 ;
      RECT 83.565 1.74 83.735 2.93 ;
      RECT 83.565 1.74 84.035 1.91 ;
      RECT 83.565 6.97 84.035 7.14 ;
      RECT 83.565 5.95 83.735 7.14 ;
      RECT 81.715 2.635 81.885 3.865 ;
      RECT 81.77 0.855 81.94 2.805 ;
      RECT 81.715 0.575 81.885 1.025 ;
      RECT 81.715 7.855 81.885 8.305 ;
      RECT 81.77 6.075 81.94 8.025 ;
      RECT 81.715 5.015 81.885 6.245 ;
      RECT 81.195 0.575 81.365 3.865 ;
      RECT 81.195 2.075 81.6 2.405 ;
      RECT 81.195 1.235 81.6 1.565 ;
      RECT 81.195 5.015 81.365 8.305 ;
      RECT 81.195 7.315 81.6 7.645 ;
      RECT 81.195 6.475 81.6 6.805 ;
      RECT 78.93 3.495 79.31 4.175 ;
      RECT 79.14 2.365 79.31 4.175 ;
      RECT 77.06 2.365 77.29 3.035 ;
      RECT 77.06 2.365 79.31 2.535 ;
      RECT 78.59 2.045 78.76 2.535 ;
      RECT 78.58 3.155 78.75 4.005 ;
      RECT 77.665 3.155 78.97 3.325 ;
      RECT 78.725 2.705 78.97 3.325 ;
      RECT 77.665 2.785 77.835 3.325 ;
      RECT 77.46 2.785 77.835 2.955 ;
      RECT 77.64 6.265 78.335 6.895 ;
      RECT 78.165 4.685 78.335 6.895 ;
      RECT 78.07 4.685 78.4 5.665 ;
      RECT 77.67 3.495 78 4.175 ;
      RECT 76.76 3.495 77.16 4.175 ;
      RECT 76.76 3.495 78 3.665 ;
      RECT 76.26 3.075 76.58 4.175 ;
      RECT 76.26 3.075 76.71 3.325 ;
      RECT 76.26 3.075 76.89 3.245 ;
      RECT 76.72 2.025 76.89 3.245 ;
      RECT 76.72 2.025 77.675 2.195 ;
      RECT 76.26 6.265 76.955 6.895 ;
      RECT 76.785 4.685 76.955 6.895 ;
      RECT 76.69 4.685 77.02 5.665 ;
      RECT 76.28 5.825 76.615 6.075 ;
      RECT 75.735 5.825 76.07 6.075 ;
      RECT 75.735 5.875 76.615 6.045 ;
      RECT 75.395 6.265 76.09 6.895 ;
      RECT 75.395 4.685 75.565 6.895 ;
      RECT 75.33 4.685 75.66 5.665 ;
      RECT 74.89 3.205 75.22 4.16 ;
      RECT 74.89 3.205 75.57 3.375 ;
      RECT 75.4 1.965 75.57 3.375 ;
      RECT 75.31 1.965 75.64 2.605 ;
      RECT 74.37 3.205 74.7 4.16 ;
      RECT 74.02 3.205 74.7 3.375 ;
      RECT 74.02 1.965 74.19 3.375 ;
      RECT 73.95 1.965 74.28 2.605 ;
      RECT 74.16 5.875 74.33 6.725 ;
      RECT 73.435 5.825 73.77 6.075 ;
      RECT 73.435 5.875 74.33 6.045 ;
      RECT 73.5 2.785 73.85 3.035 ;
      RECT 72.98 2.785 73.31 3.035 ;
      RECT 72.98 2.815 73.85 2.985 ;
      RECT 73.095 6.265 73.79 6.895 ;
      RECT 73.095 4.685 73.265 6.895 ;
      RECT 73.03 4.685 73.36 5.665 ;
      RECT 72.56 3.195 72.89 4.175 ;
      RECT 72.56 1.965 72.81 4.175 ;
      RECT 72.56 1.965 72.89 2.595 ;
      RECT 69.51 5.015 69.68 8.305 ;
      RECT 69.51 7.315 69.915 7.645 ;
      RECT 69.51 6.475 69.915 6.805 ;
      RECT 67.705 5.02 67.875 6.49 ;
      RECT 67.705 6.315 67.88 6.485 ;
      RECT 67.335 1.74 67.505 2.93 ;
      RECT 67.335 1.74 67.805 1.91 ;
      RECT 67.335 6.97 67.805 7.14 ;
      RECT 67.335 5.95 67.505 7.14 ;
      RECT 66.345 1.74 66.515 2.93 ;
      RECT 66.345 1.74 66.815 1.91 ;
      RECT 66.345 6.97 66.815 7.14 ;
      RECT 66.345 5.95 66.515 7.14 ;
      RECT 64.495 2.635 64.665 3.865 ;
      RECT 64.55 0.855 64.72 2.805 ;
      RECT 64.495 0.575 64.665 1.025 ;
      RECT 64.495 7.855 64.665 8.305 ;
      RECT 64.55 6.075 64.72 8.025 ;
      RECT 64.495 5.015 64.665 6.245 ;
      RECT 63.975 0.575 64.145 3.865 ;
      RECT 63.975 2.075 64.38 2.405 ;
      RECT 63.975 1.235 64.38 1.565 ;
      RECT 63.975 5.015 64.145 8.305 ;
      RECT 63.975 7.315 64.38 7.645 ;
      RECT 63.975 6.475 64.38 6.805 ;
      RECT 61.71 3.495 62.09 4.175 ;
      RECT 61.92 2.365 62.09 4.175 ;
      RECT 59.84 2.365 60.07 3.035 ;
      RECT 59.84 2.365 62.09 2.535 ;
      RECT 61.37 2.045 61.54 2.535 ;
      RECT 61.36 3.155 61.53 4.005 ;
      RECT 60.445 3.155 61.75 3.325 ;
      RECT 61.505 2.705 61.75 3.325 ;
      RECT 60.445 2.785 60.615 3.325 ;
      RECT 60.24 2.785 60.615 2.955 ;
      RECT 60.42 6.265 61.115 6.895 ;
      RECT 60.945 4.685 61.115 6.895 ;
      RECT 60.85 4.685 61.18 5.665 ;
      RECT 60.45 3.495 60.78 4.175 ;
      RECT 59.54 3.495 59.94 4.175 ;
      RECT 59.54 3.495 60.78 3.665 ;
      RECT 59.04 3.075 59.36 4.175 ;
      RECT 59.04 3.075 59.49 3.325 ;
      RECT 59.04 3.075 59.67 3.245 ;
      RECT 59.5 2.025 59.67 3.245 ;
      RECT 59.5 2.025 60.455 2.195 ;
      RECT 59.04 6.265 59.735 6.895 ;
      RECT 59.565 4.685 59.735 6.895 ;
      RECT 59.47 4.685 59.8 5.665 ;
      RECT 59.06 5.825 59.395 6.075 ;
      RECT 58.515 5.825 58.85 6.075 ;
      RECT 58.515 5.875 59.395 6.045 ;
      RECT 58.175 6.265 58.87 6.895 ;
      RECT 58.175 4.685 58.345 6.895 ;
      RECT 58.11 4.685 58.44 5.665 ;
      RECT 57.67 3.205 58 4.16 ;
      RECT 57.67 3.205 58.35 3.375 ;
      RECT 58.18 1.965 58.35 3.375 ;
      RECT 58.09 1.965 58.42 2.605 ;
      RECT 57.15 3.205 57.48 4.16 ;
      RECT 56.8 3.205 57.48 3.375 ;
      RECT 56.8 1.965 56.97 3.375 ;
      RECT 56.73 1.965 57.06 2.605 ;
      RECT 56.94 5.875 57.11 6.725 ;
      RECT 56.215 5.825 56.55 6.075 ;
      RECT 56.215 5.875 57.11 6.045 ;
      RECT 56.28 2.785 56.63 3.035 ;
      RECT 55.76 2.785 56.09 3.035 ;
      RECT 55.76 2.815 56.63 2.985 ;
      RECT 55.875 6.265 56.57 6.895 ;
      RECT 55.875 4.685 56.045 6.895 ;
      RECT 55.81 4.685 56.14 5.665 ;
      RECT 55.34 3.195 55.67 4.175 ;
      RECT 55.34 1.965 55.59 4.175 ;
      RECT 55.34 1.965 55.67 2.595 ;
      RECT 52.29 5.015 52.46 8.305 ;
      RECT 52.29 7.315 52.695 7.645 ;
      RECT 52.29 6.475 52.695 6.805 ;
      RECT 50.485 5.02 50.655 6.49 ;
      RECT 50.485 6.315 50.66 6.485 ;
      RECT 50.115 1.74 50.285 2.93 ;
      RECT 50.115 1.74 50.585 1.91 ;
      RECT 50.115 6.97 50.585 7.14 ;
      RECT 50.115 5.95 50.285 7.14 ;
      RECT 49.125 1.74 49.295 2.93 ;
      RECT 49.125 1.74 49.595 1.91 ;
      RECT 49.125 6.97 49.595 7.14 ;
      RECT 49.125 5.95 49.295 7.14 ;
      RECT 47.275 2.635 47.445 3.865 ;
      RECT 47.33 0.855 47.5 2.805 ;
      RECT 47.275 0.575 47.445 1.025 ;
      RECT 47.275 7.855 47.445 8.305 ;
      RECT 47.33 6.075 47.5 8.025 ;
      RECT 47.275 5.015 47.445 6.245 ;
      RECT 46.755 0.575 46.925 3.865 ;
      RECT 46.755 2.075 47.16 2.405 ;
      RECT 46.755 1.235 47.16 1.565 ;
      RECT 46.755 5.015 46.925 8.305 ;
      RECT 46.755 7.315 47.16 7.645 ;
      RECT 46.755 6.475 47.16 6.805 ;
      RECT 44.49 3.495 44.87 4.175 ;
      RECT 44.7 2.365 44.87 4.175 ;
      RECT 42.62 2.365 42.85 3.035 ;
      RECT 42.62 2.365 44.87 2.535 ;
      RECT 44.15 2.045 44.32 2.535 ;
      RECT 44.14 3.155 44.31 4.005 ;
      RECT 43.225 3.155 44.53 3.325 ;
      RECT 44.285 2.705 44.53 3.325 ;
      RECT 43.225 2.785 43.395 3.325 ;
      RECT 43.02 2.785 43.395 2.955 ;
      RECT 43.2 6.265 43.895 6.895 ;
      RECT 43.725 4.685 43.895 6.895 ;
      RECT 43.63 4.685 43.96 5.665 ;
      RECT 43.23 3.495 43.56 4.175 ;
      RECT 42.32 3.495 42.72 4.175 ;
      RECT 42.32 3.495 43.56 3.665 ;
      RECT 41.82 3.075 42.14 4.175 ;
      RECT 41.82 3.075 42.27 3.325 ;
      RECT 41.82 3.075 42.45 3.245 ;
      RECT 42.28 2.025 42.45 3.245 ;
      RECT 42.28 2.025 43.235 2.195 ;
      RECT 41.82 6.265 42.515 6.895 ;
      RECT 42.345 4.685 42.515 6.895 ;
      RECT 42.25 4.685 42.58 5.665 ;
      RECT 41.84 5.825 42.175 6.075 ;
      RECT 41.295 5.825 41.63 6.075 ;
      RECT 41.295 5.875 42.175 6.045 ;
      RECT 40.955 6.265 41.65 6.895 ;
      RECT 40.955 4.685 41.125 6.895 ;
      RECT 40.89 4.685 41.22 5.665 ;
      RECT 40.45 3.205 40.78 4.16 ;
      RECT 40.45 3.205 41.13 3.375 ;
      RECT 40.96 1.965 41.13 3.375 ;
      RECT 40.87 1.965 41.2 2.605 ;
      RECT 39.93 3.205 40.26 4.16 ;
      RECT 39.58 3.205 40.26 3.375 ;
      RECT 39.58 1.965 39.75 3.375 ;
      RECT 39.51 1.965 39.84 2.605 ;
      RECT 39.72 5.875 39.89 6.725 ;
      RECT 38.995 5.825 39.33 6.075 ;
      RECT 38.995 5.875 39.89 6.045 ;
      RECT 39.06 2.785 39.41 3.035 ;
      RECT 38.54 2.785 38.87 3.035 ;
      RECT 38.54 2.815 39.41 2.985 ;
      RECT 38.655 6.265 39.35 6.895 ;
      RECT 38.655 4.685 38.825 6.895 ;
      RECT 38.59 4.685 38.92 5.665 ;
      RECT 38.12 3.195 38.45 4.175 ;
      RECT 38.12 1.965 38.37 4.175 ;
      RECT 38.12 1.965 38.45 2.595 ;
      RECT 35.07 5.015 35.24 8.305 ;
      RECT 35.07 7.315 35.475 7.645 ;
      RECT 35.07 6.475 35.475 6.805 ;
      RECT 33.265 5.02 33.435 6.49 ;
      RECT 33.265 6.315 33.44 6.485 ;
      RECT 32.895 1.74 33.065 2.93 ;
      RECT 32.895 1.74 33.365 1.91 ;
      RECT 32.895 6.97 33.365 7.14 ;
      RECT 32.895 5.95 33.065 7.14 ;
      RECT 31.905 1.74 32.075 2.93 ;
      RECT 31.905 1.74 32.375 1.91 ;
      RECT 31.905 6.97 32.375 7.14 ;
      RECT 31.905 5.95 32.075 7.14 ;
      RECT 30.055 2.635 30.225 3.865 ;
      RECT 30.11 0.855 30.28 2.805 ;
      RECT 30.055 0.575 30.225 1.025 ;
      RECT 30.055 7.855 30.225 8.305 ;
      RECT 30.11 6.075 30.28 8.025 ;
      RECT 30.055 5.015 30.225 6.245 ;
      RECT 29.535 0.575 29.705 3.865 ;
      RECT 29.535 2.075 29.94 2.405 ;
      RECT 29.535 1.235 29.94 1.565 ;
      RECT 29.535 5.015 29.705 8.305 ;
      RECT 29.535 7.315 29.94 7.645 ;
      RECT 29.535 6.475 29.94 6.805 ;
      RECT 27.27 3.495 27.65 4.175 ;
      RECT 27.48 2.365 27.65 4.175 ;
      RECT 25.4 2.365 25.63 3.035 ;
      RECT 25.4 2.365 27.65 2.535 ;
      RECT 26.93 2.045 27.1 2.535 ;
      RECT 26.92 3.155 27.09 4.005 ;
      RECT 26.005 3.155 27.31 3.325 ;
      RECT 27.065 2.705 27.31 3.325 ;
      RECT 26.005 2.785 26.175 3.325 ;
      RECT 25.8 2.785 26.175 2.955 ;
      RECT 25.98 6.265 26.675 6.895 ;
      RECT 26.505 4.685 26.675 6.895 ;
      RECT 26.41 4.685 26.74 5.665 ;
      RECT 26.01 3.495 26.34 4.175 ;
      RECT 25.1 3.495 25.5 4.175 ;
      RECT 25.1 3.495 26.34 3.665 ;
      RECT 24.6 3.075 24.92 4.175 ;
      RECT 24.6 3.075 25.05 3.325 ;
      RECT 24.6 3.075 25.23 3.245 ;
      RECT 25.06 2.025 25.23 3.245 ;
      RECT 25.06 2.025 26.015 2.195 ;
      RECT 24.6 6.265 25.295 6.895 ;
      RECT 25.125 4.685 25.295 6.895 ;
      RECT 25.03 4.685 25.36 5.665 ;
      RECT 24.62 5.825 24.955 6.075 ;
      RECT 24.075 5.825 24.41 6.075 ;
      RECT 24.075 5.875 24.955 6.045 ;
      RECT 23.735 6.265 24.43 6.895 ;
      RECT 23.735 4.685 23.905 6.895 ;
      RECT 23.67 4.685 24 5.665 ;
      RECT 23.23 3.205 23.56 4.16 ;
      RECT 23.23 3.205 23.91 3.375 ;
      RECT 23.74 1.965 23.91 3.375 ;
      RECT 23.65 1.965 23.98 2.605 ;
      RECT 22.71 3.205 23.04 4.16 ;
      RECT 22.36 3.205 23.04 3.375 ;
      RECT 22.36 1.965 22.53 3.375 ;
      RECT 22.29 1.965 22.62 2.605 ;
      RECT 22.5 5.875 22.67 6.725 ;
      RECT 21.775 5.825 22.11 6.075 ;
      RECT 21.775 5.875 22.67 6.045 ;
      RECT 21.84 2.785 22.19 3.035 ;
      RECT 21.32 2.785 21.65 3.035 ;
      RECT 21.32 2.815 22.19 2.985 ;
      RECT 21.435 6.265 22.13 6.895 ;
      RECT 21.435 4.685 21.605 6.895 ;
      RECT 21.37 4.685 21.7 5.665 ;
      RECT 20.9 3.195 21.23 4.175 ;
      RECT 20.9 1.965 21.15 4.175 ;
      RECT 20.9 1.965 21.23 2.595 ;
      RECT 17.85 5.015 18.02 8.305 ;
      RECT 17.85 7.315 18.255 7.645 ;
      RECT 17.85 6.475 18.255 6.805 ;
      RECT 16.045 5.02 16.215 6.49 ;
      RECT 16.045 6.315 16.22 6.485 ;
      RECT 15.675 1.74 15.845 2.93 ;
      RECT 15.675 1.74 16.145 1.91 ;
      RECT 15.675 6.97 16.145 7.14 ;
      RECT 15.675 5.95 15.845 7.14 ;
      RECT 14.685 1.74 14.855 2.93 ;
      RECT 14.685 1.74 15.155 1.91 ;
      RECT 14.685 6.97 15.155 7.14 ;
      RECT 14.685 5.95 14.855 7.14 ;
      RECT 12.835 2.635 13.005 3.865 ;
      RECT 12.89 0.855 13.06 2.805 ;
      RECT 12.835 0.575 13.005 1.025 ;
      RECT 12.835 7.855 13.005 8.305 ;
      RECT 12.89 6.075 13.06 8.025 ;
      RECT 12.835 5.015 13.005 6.245 ;
      RECT 12.315 0.575 12.485 3.865 ;
      RECT 12.315 2.075 12.72 2.405 ;
      RECT 12.315 1.235 12.72 1.565 ;
      RECT 12.315 5.015 12.485 8.305 ;
      RECT 12.315 7.315 12.72 7.645 ;
      RECT 12.315 6.475 12.72 6.805 ;
      RECT 10.05 3.495 10.43 4.175 ;
      RECT 10.26 2.365 10.43 4.175 ;
      RECT 8.18 2.365 8.41 3.035 ;
      RECT 8.18 2.365 10.43 2.535 ;
      RECT 9.71 2.045 9.88 2.535 ;
      RECT 9.7 3.155 9.87 4.005 ;
      RECT 8.785 3.155 10.09 3.325 ;
      RECT 9.845 2.705 10.09 3.325 ;
      RECT 8.785 2.785 8.955 3.325 ;
      RECT 8.58 2.785 8.955 2.955 ;
      RECT 8.76 6.265 9.455 6.895 ;
      RECT 9.285 4.685 9.455 6.895 ;
      RECT 9.19 4.685 9.52 5.665 ;
      RECT 8.79 3.495 9.12 4.175 ;
      RECT 7.88 3.495 8.28 4.175 ;
      RECT 7.88 3.495 9.12 3.665 ;
      RECT 7.38 3.075 7.7 4.175 ;
      RECT 7.38 3.075 7.83 3.325 ;
      RECT 7.38 3.075 8.01 3.245 ;
      RECT 7.84 2.025 8.01 3.245 ;
      RECT 7.84 2.025 8.795 2.195 ;
      RECT 7.38 6.265 8.075 6.895 ;
      RECT 7.905 4.685 8.075 6.895 ;
      RECT 7.81 4.685 8.14 5.665 ;
      RECT 7.4 5.825 7.735 6.075 ;
      RECT 6.855 5.825 7.19 6.075 ;
      RECT 6.855 5.875 7.735 6.045 ;
      RECT 6.515 6.265 7.21 6.895 ;
      RECT 6.515 4.685 6.685 6.895 ;
      RECT 6.45 4.685 6.78 5.665 ;
      RECT 6.01 3.205 6.34 4.16 ;
      RECT 6.01 3.205 6.69 3.375 ;
      RECT 6.52 1.965 6.69 3.375 ;
      RECT 6.43 1.965 6.76 2.605 ;
      RECT 5.49 3.205 5.82 4.16 ;
      RECT 5.14 3.205 5.82 3.375 ;
      RECT 5.14 1.965 5.31 3.375 ;
      RECT 5.07 1.965 5.4 2.605 ;
      RECT 5.28 5.875 5.45 6.725 ;
      RECT 4.555 5.825 4.89 6.075 ;
      RECT 4.555 5.875 5.45 6.045 ;
      RECT 4.62 2.785 4.97 3.035 ;
      RECT 4.1 2.785 4.43 3.035 ;
      RECT 4.1 2.815 4.97 2.985 ;
      RECT 4.215 6.265 4.91 6.895 ;
      RECT 4.215 4.685 4.385 6.895 ;
      RECT 4.15 4.685 4.48 5.665 ;
      RECT 3.68 3.195 4.01 4.175 ;
      RECT 3.68 1.965 3.93 4.175 ;
      RECT 3.68 1.965 4.01 2.595 ;
      RECT 0.63 5.015 0.8 8.305 ;
      RECT 0.63 7.315 1.035 7.645 ;
      RECT 0.63 6.475 1.035 6.805 ;
      RECT -2.26 7.855 -2.09 8.305 ;
      RECT -2.205 6.075 -2.035 8.025 ;
      RECT -2.26 5.015 -2.09 6.245 ;
      RECT -2.78 5.015 -2.61 8.305 ;
      RECT -2.78 7.315 -2.375 7.645 ;
      RECT -2.78 6.475 -2.375 6.805 ;
      RECT 84.925 7.8 85.095 8.31 ;
      RECT 83.935 0.57 84.105 1.08 ;
      RECT 83.935 2.39 84.105 3.86 ;
      RECT 83.935 5.02 84.105 6.49 ;
      RECT 83.935 7.8 84.105 8.31 ;
      RECT 82.575 0.575 82.745 3.865 ;
      RECT 82.575 5.015 82.745 8.305 ;
      RECT 82.145 0.575 82.315 1.085 ;
      RECT 82.145 1.655 82.315 3.865 ;
      RECT 82.145 5.015 82.315 7.225 ;
      RECT 82.145 7.795 82.315 8.305 ;
      RECT 78.505 5.825 78.84 6.095 ;
      RECT 78.005 2.785 78.555 2.985 ;
      RECT 77.66 5.825 77.995 6.075 ;
      RECT 77.125 5.825 77.46 6.095 ;
      RECT 75.74 2.785 76.09 3.035 ;
      RECT 74.88 2.785 75.23 3.035 ;
      RECT 74.36 2.785 74.71 3.035 ;
      RECT 70.89 5.015 71.06 8.305 ;
      RECT 70.46 5.015 70.63 7.225 ;
      RECT 70.46 7.795 70.63 8.305 ;
      RECT 67.705 7.8 67.875 8.31 ;
      RECT 66.715 0.57 66.885 1.08 ;
      RECT 66.715 2.39 66.885 3.86 ;
      RECT 66.715 5.02 66.885 6.49 ;
      RECT 66.715 7.8 66.885 8.31 ;
      RECT 65.355 0.575 65.525 3.865 ;
      RECT 65.355 5.015 65.525 8.305 ;
      RECT 64.925 0.575 65.095 1.085 ;
      RECT 64.925 1.655 65.095 3.865 ;
      RECT 64.925 5.015 65.095 7.225 ;
      RECT 64.925 7.795 65.095 8.305 ;
      RECT 61.285 5.825 61.62 6.095 ;
      RECT 60.785 2.785 61.335 2.985 ;
      RECT 60.44 5.825 60.775 6.075 ;
      RECT 59.905 5.825 60.24 6.095 ;
      RECT 58.52 2.785 58.87 3.035 ;
      RECT 57.66 2.785 58.01 3.035 ;
      RECT 57.14 2.785 57.49 3.035 ;
      RECT 53.67 5.015 53.84 8.305 ;
      RECT 53.24 5.015 53.41 7.225 ;
      RECT 53.24 7.795 53.41 8.305 ;
      RECT 50.485 7.8 50.655 8.31 ;
      RECT 49.495 0.57 49.665 1.08 ;
      RECT 49.495 2.39 49.665 3.86 ;
      RECT 49.495 5.02 49.665 6.49 ;
      RECT 49.495 7.8 49.665 8.31 ;
      RECT 48.135 0.575 48.305 3.865 ;
      RECT 48.135 5.015 48.305 8.305 ;
      RECT 47.705 0.575 47.875 1.085 ;
      RECT 47.705 1.655 47.875 3.865 ;
      RECT 47.705 5.015 47.875 7.225 ;
      RECT 47.705 7.795 47.875 8.305 ;
      RECT 44.065 5.825 44.4 6.095 ;
      RECT 43.565 2.785 44.115 2.985 ;
      RECT 43.22 5.825 43.555 6.075 ;
      RECT 42.685 5.825 43.02 6.095 ;
      RECT 41.3 2.785 41.65 3.035 ;
      RECT 40.44 2.785 40.79 3.035 ;
      RECT 39.92 2.785 40.27 3.035 ;
      RECT 36.45 5.015 36.62 8.305 ;
      RECT 36.02 5.015 36.19 7.225 ;
      RECT 36.02 7.795 36.19 8.305 ;
      RECT 33.265 7.8 33.435 8.31 ;
      RECT 32.275 0.57 32.445 1.08 ;
      RECT 32.275 2.39 32.445 3.86 ;
      RECT 32.275 5.02 32.445 6.49 ;
      RECT 32.275 7.8 32.445 8.31 ;
      RECT 30.915 0.575 31.085 3.865 ;
      RECT 30.915 5.015 31.085 8.305 ;
      RECT 30.485 0.575 30.655 1.085 ;
      RECT 30.485 1.655 30.655 3.865 ;
      RECT 30.485 5.015 30.655 7.225 ;
      RECT 30.485 7.795 30.655 8.305 ;
      RECT 26.845 5.825 27.18 6.095 ;
      RECT 26.345 2.785 26.895 2.985 ;
      RECT 26 5.825 26.335 6.075 ;
      RECT 25.465 5.825 25.8 6.095 ;
      RECT 24.08 2.785 24.43 3.035 ;
      RECT 23.22 2.785 23.57 3.035 ;
      RECT 22.7 2.785 23.05 3.035 ;
      RECT 19.23 5.015 19.4 8.305 ;
      RECT 18.8 5.015 18.97 7.225 ;
      RECT 18.8 7.795 18.97 8.305 ;
      RECT 16.045 7.8 16.215 8.31 ;
      RECT 15.055 0.57 15.225 1.08 ;
      RECT 15.055 2.39 15.225 3.86 ;
      RECT 15.055 5.02 15.225 6.49 ;
      RECT 15.055 7.8 15.225 8.31 ;
      RECT 13.695 0.575 13.865 3.865 ;
      RECT 13.695 5.015 13.865 8.305 ;
      RECT 13.265 0.575 13.435 1.085 ;
      RECT 13.265 1.655 13.435 3.865 ;
      RECT 13.265 5.015 13.435 7.225 ;
      RECT 13.265 7.795 13.435 8.305 ;
      RECT 9.625 5.825 9.96 6.095 ;
      RECT 9.125 2.785 9.675 2.985 ;
      RECT 8.78 5.825 9.115 6.075 ;
      RECT 8.245 5.825 8.58 6.095 ;
      RECT 6.86 2.785 7.21 3.035 ;
      RECT 6 2.785 6.35 3.035 ;
      RECT 5.48 2.785 5.83 3.035 ;
      RECT 2.01 5.015 2.18 8.305 ;
      RECT 1.58 5.015 1.75 7.225 ;
      RECT 1.58 7.795 1.75 8.305 ;
      RECT -1.83 5.015 -1.66 7.225 ;
      RECT -1.83 7.795 -1.66 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2ct_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2ct_8_b0r2
  CLASS BLOCK ;
  ORIGIN 3.43 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ct_8_b0r2 ;
  SIZE 88.9 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 16.05 0.915 16.22 1.085 ;
        RECT 16.045 0.91 16.215 1.08 ;
        RECT 16.045 2.39 16.215 2.56 ;
      LAYER li1 ;
        RECT 16.05 0.915 16.22 1.085 ;
        RECT 16.045 0.57 16.215 1.08 ;
        RECT 16.045 2.39 16.215 3.86 ;
      LAYER met1 ;
        RECT 15.985 2.36 16.275 2.59 ;
        RECT 15.985 0.88 16.275 1.11 ;
        RECT 16.045 0.88 16.215 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 33.27 0.915 33.44 1.085 ;
        RECT 33.265 0.91 33.435 1.08 ;
        RECT 33.265 2.39 33.435 2.56 ;
      LAYER li1 ;
        RECT 33.27 0.915 33.44 1.085 ;
        RECT 33.265 0.57 33.435 1.08 ;
        RECT 33.265 2.39 33.435 3.86 ;
      LAYER met1 ;
        RECT 33.205 2.36 33.495 2.59 ;
        RECT 33.205 0.88 33.495 1.11 ;
        RECT 33.265 0.88 33.435 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 50.49 0.915 50.66 1.085 ;
        RECT 50.485 0.91 50.655 1.08 ;
        RECT 50.485 2.39 50.655 2.56 ;
      LAYER li1 ;
        RECT 50.49 0.915 50.66 1.085 ;
        RECT 50.485 0.57 50.655 1.08 ;
        RECT 50.485 2.39 50.655 3.86 ;
      LAYER met1 ;
        RECT 50.425 2.36 50.715 2.59 ;
        RECT 50.425 0.88 50.715 1.11 ;
        RECT 50.485 0.88 50.655 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 67.71 0.915 67.88 1.085 ;
        RECT 67.705 0.91 67.875 1.08 ;
        RECT 67.705 2.39 67.875 2.56 ;
      LAYER li1 ;
        RECT 67.71 0.915 67.88 1.085 ;
        RECT 67.705 0.57 67.875 1.08 ;
        RECT 67.705 2.39 67.875 3.86 ;
      LAYER met1 ;
        RECT 67.645 2.36 67.935 2.59 ;
        RECT 67.645 0.88 67.935 1.11 ;
        RECT 67.705 0.88 67.875 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 84.93 0.915 85.1 1.085 ;
        RECT 84.925 0.91 85.095 1.08 ;
        RECT 84.925 2.39 85.095 2.56 ;
      LAYER li1 ;
        RECT 84.93 0.915 85.1 1.085 ;
        RECT 84.925 0.57 85.095 1.08 ;
        RECT 84.925 2.39 85.095 3.86 ;
      LAYER met1 ;
        RECT 84.865 2.36 85.155 2.59 ;
        RECT 84.865 0.88 85.155 1.11 ;
        RECT 84.925 0.88 85.095 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 11.895 1.66 12.065 2.935 ;
        RECT 11.895 5.94 12.065 7.22 ;
        RECT 11.885 5.94 12.065 6.18 ;
        RECT 0.21 5.945 0.38 7.22 ;
      LAYER met2 ;
        RECT 11.815 5.855 12.14 6.18 ;
        RECT 11.815 3.495 12.14 3.82 ;
        RECT 2.515 7.55 12.065 7.72 ;
        RECT 11.895 5.855 12.065 7.72 ;
        RECT 11.885 3.495 12.055 6.18 ;
        RECT 2.46 5.86 2.74 6.2 ;
        RECT 2.515 5.86 2.685 7.72 ;
      LAYER met1 ;
        RECT 11.835 2.765 12.295 2.935 ;
        RECT 11.815 3.495 12.14 3.82 ;
        RECT 11.835 2.735 12.125 2.965 ;
        RECT 11.895 2.735 12.065 3.82 ;
        RECT 11.815 5.945 12.295 6.115 ;
        RECT 11.815 5.855 12.14 6.18 ;
        RECT 2.43 5.89 2.77 6.17 ;
        RECT 0.15 5.945 2.77 6.115 ;
        RECT 0.15 5.915 0.44 6.145 ;
      LAYER via1 ;
        RECT 2.525 5.955 2.675 6.105 ;
        RECT 11.905 5.94 12.055 6.09 ;
        RECT 11.905 3.58 12.055 3.73 ;
      LAYER mcon ;
        RECT 0.21 5.945 0.38 6.115 ;
        RECT 11.895 5.945 12.065 6.115 ;
        RECT 11.895 2.765 12.065 2.935 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 29.115 1.66 29.285 2.935 ;
        RECT 29.115 5.94 29.285 7.22 ;
        RECT 29.105 5.94 29.285 6.18 ;
        RECT 17.43 5.945 17.6 7.22 ;
      LAYER met2 ;
        RECT 29.035 5.855 29.36 6.18 ;
        RECT 29.035 3.495 29.36 3.82 ;
        RECT 19.735 7.55 29.285 7.72 ;
        RECT 29.115 5.855 29.285 7.72 ;
        RECT 29.105 3.495 29.275 6.18 ;
        RECT 19.68 5.86 19.96 6.2 ;
        RECT 19.735 5.86 19.905 7.72 ;
      LAYER met1 ;
        RECT 29.055 2.765 29.515 2.935 ;
        RECT 29.035 3.495 29.36 3.82 ;
        RECT 29.055 2.735 29.345 2.965 ;
        RECT 29.115 2.735 29.285 3.82 ;
        RECT 29.035 5.945 29.515 6.115 ;
        RECT 29.035 5.855 29.36 6.18 ;
        RECT 19.65 5.89 19.99 6.17 ;
        RECT 17.37 5.945 19.99 6.115 ;
        RECT 17.37 5.915 17.66 6.145 ;
      LAYER via1 ;
        RECT 19.745 5.955 19.895 6.105 ;
        RECT 29.125 5.94 29.275 6.09 ;
        RECT 29.125 3.58 29.275 3.73 ;
      LAYER mcon ;
        RECT 17.43 5.945 17.6 6.115 ;
        RECT 29.115 5.945 29.285 6.115 ;
        RECT 29.115 2.765 29.285 2.935 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 46.335 1.66 46.505 2.935 ;
        RECT 46.335 5.94 46.505 7.22 ;
        RECT 46.325 5.94 46.505 6.18 ;
        RECT 34.65 5.945 34.82 7.22 ;
      LAYER met2 ;
        RECT 46.255 5.855 46.58 6.18 ;
        RECT 46.255 3.495 46.58 3.82 ;
        RECT 36.955 7.55 46.505 7.72 ;
        RECT 46.335 5.855 46.505 7.72 ;
        RECT 46.325 3.495 46.495 6.18 ;
        RECT 36.9 5.86 37.18 6.2 ;
        RECT 36.955 5.86 37.125 7.72 ;
      LAYER met1 ;
        RECT 46.275 2.765 46.735 2.935 ;
        RECT 46.255 3.495 46.58 3.82 ;
        RECT 46.275 2.735 46.565 2.965 ;
        RECT 46.335 2.735 46.505 3.82 ;
        RECT 46.255 5.945 46.735 6.115 ;
        RECT 46.255 5.855 46.58 6.18 ;
        RECT 36.87 5.89 37.21 6.17 ;
        RECT 34.59 5.945 37.21 6.115 ;
        RECT 34.59 5.915 34.88 6.145 ;
      LAYER via1 ;
        RECT 36.965 5.955 37.115 6.105 ;
        RECT 46.345 5.94 46.495 6.09 ;
        RECT 46.345 3.58 46.495 3.73 ;
      LAYER mcon ;
        RECT 34.65 5.945 34.82 6.115 ;
        RECT 46.335 5.945 46.505 6.115 ;
        RECT 46.335 2.765 46.505 2.935 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 63.555 1.66 63.725 2.935 ;
        RECT 63.555 5.94 63.725 7.22 ;
        RECT 63.545 5.94 63.725 6.18 ;
        RECT 51.87 5.945 52.04 7.22 ;
      LAYER met2 ;
        RECT 63.475 5.855 63.8 6.18 ;
        RECT 63.475 3.495 63.8 3.82 ;
        RECT 54.175 7.55 63.725 7.72 ;
        RECT 63.555 5.855 63.725 7.72 ;
        RECT 63.545 3.495 63.715 6.18 ;
        RECT 54.12 5.86 54.4 6.2 ;
        RECT 54.175 5.86 54.345 7.72 ;
      LAYER met1 ;
        RECT 63.495 2.765 63.955 2.935 ;
        RECT 63.475 3.495 63.8 3.82 ;
        RECT 63.495 2.735 63.785 2.965 ;
        RECT 63.555 2.735 63.725 3.82 ;
        RECT 63.475 5.945 63.955 6.115 ;
        RECT 63.475 5.855 63.8 6.18 ;
        RECT 54.09 5.89 54.43 6.17 ;
        RECT 51.81 5.945 54.43 6.115 ;
        RECT 51.81 5.915 52.1 6.145 ;
      LAYER via1 ;
        RECT 54.185 5.955 54.335 6.105 ;
        RECT 63.565 5.94 63.715 6.09 ;
        RECT 63.565 3.58 63.715 3.73 ;
      LAYER mcon ;
        RECT 51.87 5.945 52.04 6.115 ;
        RECT 63.555 5.945 63.725 6.115 ;
        RECT 63.555 2.765 63.725 2.935 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 80.775 1.66 80.945 2.935 ;
        RECT 80.775 5.94 80.945 7.22 ;
        RECT 80.765 5.94 80.945 6.18 ;
        RECT 69.09 5.945 69.26 7.22 ;
      LAYER met2 ;
        RECT 80.695 5.855 81.02 6.18 ;
        RECT 80.695 3.495 81.02 3.82 ;
        RECT 71.395 7.55 80.945 7.72 ;
        RECT 80.775 5.855 80.945 7.72 ;
        RECT 80.765 3.495 80.935 6.18 ;
        RECT 71.34 5.86 71.62 6.2 ;
        RECT 71.395 5.86 71.565 7.72 ;
      LAYER met1 ;
        RECT 80.715 2.765 81.175 2.935 ;
        RECT 80.695 3.495 81.02 3.82 ;
        RECT 80.715 2.735 81.005 2.965 ;
        RECT 80.775 2.735 80.945 3.82 ;
        RECT 80.695 5.945 81.175 6.115 ;
        RECT 80.695 5.855 81.02 6.18 ;
        RECT 71.31 5.89 71.65 6.17 ;
        RECT 69.03 5.945 71.65 6.115 ;
        RECT 69.03 5.915 69.32 6.145 ;
      LAYER via1 ;
        RECT 71.405 5.955 71.555 6.105 ;
        RECT 80.785 5.94 80.935 6.09 ;
        RECT 80.785 3.58 80.935 3.73 ;
      LAYER mcon ;
        RECT 69.09 5.945 69.26 6.115 ;
        RECT 80.775 5.945 80.945 6.115 ;
        RECT 80.775 2.765 80.945 2.935 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT -3.2 5.945 -3.03 7.22 ;
      LAYER met1 ;
        RECT -3.26 5.945 -2.8 6.115 ;
        RECT -3.26 5.915 -2.97 6.145 ;
      LAYER mcon ;
        RECT -3.2 5.945 -3.03 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 79.485 4.135 85.47 4.745 ;
        RECT 83.335 4.13 85.315 4.75 ;
        RECT 84.495 3.4 84.665 5.48 ;
        RECT 83.505 3.4 83.675 5.48 ;
        RECT 80.765 3.405 80.935 5.475 ;
        RECT -3.43 4.345 85.47 4.515 ;
        RECT 79.48 4.135 85.47 4.515 ;
        RECT 78.57 4.345 78.85 5.655 ;
        RECT 78.17 3.495 78.34 4.515 ;
        RECT 77.64 4.345 77.9 5.655 ;
        RECT 77.33 3.835 77.5 4.515 ;
        RECT 77.19 4.345 77.47 5.655 ;
        RECT 76.26 4.345 76.52 5.655 ;
        RECT 75.83 4.345 76.09 5.655 ;
        RECT 75.75 3.205 76.08 4.515 ;
        RECT 74.88 4.345 75.16 5.655 ;
        RECT 73.51 3.205 73.84 4.515 ;
        RECT 73.53 3.205 73.79 5.655 ;
        RECT 73.06 3.205 73.29 4.515 ;
        RECT 72.58 4.345 72.86 5.655 ;
        RECT 62.265 4.345 72.41 4.74 ;
        RECT 62.26 4.135 72.39 4.515 ;
        RECT 72.18 3.205 72.39 4.74 ;
        RECT 68.245 4.13 72.39 4.74 ;
        RECT 68.905 4.13 71.655 4.745 ;
        RECT 69.08 4.13 69.25 5.475 ;
        RECT 62.265 4.135 68.25 4.745 ;
        RECT 66.115 4.13 68.095 4.75 ;
        RECT 67.275 3.4 67.445 5.48 ;
        RECT 66.285 3.4 66.455 5.48 ;
        RECT 63.545 3.405 63.715 5.475 ;
        RECT 61.35 4.345 61.63 5.655 ;
        RECT 60.95 3.495 61.12 4.515 ;
        RECT 60.42 4.345 60.68 5.655 ;
        RECT 60.11 3.835 60.28 4.515 ;
        RECT 59.97 4.345 60.25 5.655 ;
        RECT 59.04 4.345 59.3 5.655 ;
        RECT 58.61 4.345 58.87 5.655 ;
        RECT 58.53 3.205 58.86 4.515 ;
        RECT 57.66 4.345 57.94 5.655 ;
        RECT 56.29 3.205 56.62 4.515 ;
        RECT 56.31 3.205 56.57 5.655 ;
        RECT 55.84 3.205 56.07 4.515 ;
        RECT 55.36 4.345 55.64 5.655 ;
        RECT 45.045 4.345 55.19 4.74 ;
        RECT 45.04 4.135 55.17 4.515 ;
        RECT 54.96 3.205 55.17 4.74 ;
        RECT 51.025 4.13 55.17 4.74 ;
        RECT 51.685 4.13 54.435 4.745 ;
        RECT 51.86 4.13 52.03 5.475 ;
        RECT 45.045 4.135 51.03 4.745 ;
        RECT 48.895 4.13 50.875 4.75 ;
        RECT 50.055 3.4 50.225 5.48 ;
        RECT 49.065 3.4 49.235 5.48 ;
        RECT 46.325 3.405 46.495 5.475 ;
        RECT 44.13 4.345 44.41 5.655 ;
        RECT 43.73 3.495 43.9 4.515 ;
        RECT 43.2 4.345 43.46 5.655 ;
        RECT 42.89 3.835 43.06 4.515 ;
        RECT 42.75 4.345 43.03 5.655 ;
        RECT 41.82 4.345 42.08 5.655 ;
        RECT 41.39 4.345 41.65 5.655 ;
        RECT 41.31 3.205 41.64 4.515 ;
        RECT 40.44 4.345 40.72 5.655 ;
        RECT 39.07 3.205 39.4 4.515 ;
        RECT 39.09 3.205 39.35 5.655 ;
        RECT 38.62 3.205 38.85 4.515 ;
        RECT 38.14 4.345 38.42 5.655 ;
        RECT 27.825 4.345 37.97 4.74 ;
        RECT 27.82 4.135 37.95 4.515 ;
        RECT 37.74 3.205 37.95 4.74 ;
        RECT 33.805 4.13 37.95 4.74 ;
        RECT 34.465 4.13 37.215 4.745 ;
        RECT 34.64 4.13 34.81 5.475 ;
        RECT 27.825 4.135 33.81 4.745 ;
        RECT 31.675 4.13 33.655 4.75 ;
        RECT 32.835 3.4 33.005 5.48 ;
        RECT 31.845 3.4 32.015 5.48 ;
        RECT 29.105 3.405 29.275 5.475 ;
        RECT 26.91 4.345 27.19 5.655 ;
        RECT 26.51 3.495 26.68 4.515 ;
        RECT 25.98 4.345 26.24 5.655 ;
        RECT 25.67 3.835 25.84 4.515 ;
        RECT 25.53 4.345 25.81 5.655 ;
        RECT 24.6 4.345 24.86 5.655 ;
        RECT 24.17 4.345 24.43 5.655 ;
        RECT 24.09 3.205 24.42 4.515 ;
        RECT 23.22 4.345 23.5 5.655 ;
        RECT 21.85 3.205 22.18 4.515 ;
        RECT 21.87 3.205 22.13 5.655 ;
        RECT 21.4 3.205 21.63 4.515 ;
        RECT 20.92 4.345 21.2 5.655 ;
        RECT 10.605 4.345 20.75 4.74 ;
        RECT 10.6 4.135 20.73 4.515 ;
        RECT 20.52 3.205 20.73 4.74 ;
        RECT 16.585 4.13 20.73 4.74 ;
        RECT 17.245 4.13 19.995 4.745 ;
        RECT 17.42 4.13 17.59 5.475 ;
        RECT 10.605 4.135 16.59 4.745 ;
        RECT 14.455 4.13 16.435 4.75 ;
        RECT 15.615 3.4 15.785 5.48 ;
        RECT 14.625 3.4 14.795 5.48 ;
        RECT 11.885 3.405 12.055 5.475 ;
        RECT 9.69 4.345 9.97 5.655 ;
        RECT 9.29 3.495 9.46 4.515 ;
        RECT 8.76 4.345 9.02 5.655 ;
        RECT 8.45 3.835 8.62 4.515 ;
        RECT 8.31 4.345 8.59 5.655 ;
        RECT 7.38 4.345 7.64 5.655 ;
        RECT 6.95 4.345 7.21 5.655 ;
        RECT 6.87 3.205 7.2 4.515 ;
        RECT 6 4.345 6.28 5.655 ;
        RECT 4.63 3.205 4.96 4.515 ;
        RECT 4.65 3.205 4.91 5.655 ;
        RECT 4.18 3.205 4.41 4.515 ;
        RECT 3.7 4.345 3.98 5.655 ;
        RECT -3.43 4.345 3.53 4.74 ;
        RECT -3.43 4.13 3.51 4.74 ;
        RECT 3.3 3.205 3.51 4.74 ;
        RECT 0.025 4.13 2.775 4.745 ;
        RECT 0.2 4.13 0.37 5.475 ;
        RECT -3.385 4.13 -0.635 4.745 ;
        RECT -1.4 4.13 -1.23 8.305 ;
        RECT -3.21 4.13 -3.04 5.475 ;
      LAYER met1 ;
        RECT 79.485 4.135 85.47 4.745 ;
        RECT 83.335 4.13 85.315 4.75 ;
        RECT -3.43 4.19 85.47 4.67 ;
        RECT 79.48 4.135 85.47 4.67 ;
        RECT 62.265 4.19 72.41 4.74 ;
        RECT 62.26 4.135 72.39 4.67 ;
        RECT 68.245 4.13 72.39 4.74 ;
        RECT 68.905 4.13 71.655 4.745 ;
        RECT 62.265 4.135 68.25 4.745 ;
        RECT 66.115 4.13 68.095 4.75 ;
        RECT 45.045 4.19 55.19 4.74 ;
        RECT 45.04 4.135 55.17 4.67 ;
        RECT 51.025 4.13 55.17 4.74 ;
        RECT 51.685 4.13 54.435 4.745 ;
        RECT 45.045 4.135 51.03 4.745 ;
        RECT 48.895 4.13 50.875 4.75 ;
        RECT 27.825 4.19 37.97 4.74 ;
        RECT 27.82 4.135 37.95 4.67 ;
        RECT 33.805 4.13 37.95 4.74 ;
        RECT 34.465 4.13 37.215 4.745 ;
        RECT 27.825 4.135 33.81 4.745 ;
        RECT 31.675 4.13 33.655 4.75 ;
        RECT 10.605 4.19 20.75 4.74 ;
        RECT 10.6 4.135 20.73 4.67 ;
        RECT 16.585 4.13 20.73 4.74 ;
        RECT 17.245 4.13 19.995 4.745 ;
        RECT 10.605 4.135 16.59 4.745 ;
        RECT 14.455 4.13 16.435 4.75 ;
        RECT -3.43 4.19 3.53 4.74 ;
        RECT -3.43 4.13 3.51 4.74 ;
        RECT 0.025 4.13 2.775 4.745 ;
        RECT -3.385 4.13 -0.635 4.745 ;
        RECT -1.46 6.655 -1.17 6.885 ;
        RECT -1.63 6.685 -1.17 6.855 ;
      LAYER mcon ;
        RECT -1.4 6.685 -1.23 6.855 ;
        RECT -1.09 4.545 -0.92 4.715 ;
        RECT 2.32 4.545 2.49 4.715 ;
        RECT 3.3 4.345 3.47 4.515 ;
        RECT 3.76 4.345 3.93 4.515 ;
        RECT 4.22 4.345 4.39 4.515 ;
        RECT 4.68 4.345 4.85 4.515 ;
        RECT 5.14 4.345 5.31 4.515 ;
        RECT 5.6 4.345 5.77 4.515 ;
        RECT 6.06 4.345 6.23 4.515 ;
        RECT 6.52 4.345 6.69 4.515 ;
        RECT 6.98 4.345 7.15 4.515 ;
        RECT 7.44 4.345 7.61 4.515 ;
        RECT 7.9 4.345 8.07 4.515 ;
        RECT 8.36 4.345 8.53 4.515 ;
        RECT 8.82 4.345 8.99 4.515 ;
        RECT 9.28 4.345 9.45 4.515 ;
        RECT 9.74 4.345 9.91 4.515 ;
        RECT 10.2 4.345 10.37 4.515 ;
        RECT 14.005 4.545 14.175 4.715 ;
        RECT 14.005 4.165 14.175 4.335 ;
        RECT 14.705 4.55 14.875 4.72 ;
        RECT 14.705 4.16 14.875 4.33 ;
        RECT 15.695 4.55 15.865 4.72 ;
        RECT 15.695 4.16 15.865 4.33 ;
        RECT 19.54 4.545 19.71 4.715 ;
        RECT 20.52 4.345 20.69 4.515 ;
        RECT 20.98 4.345 21.15 4.515 ;
        RECT 21.44 4.345 21.61 4.515 ;
        RECT 21.9 4.345 22.07 4.515 ;
        RECT 22.36 4.345 22.53 4.515 ;
        RECT 22.82 4.345 22.99 4.515 ;
        RECT 23.28 4.345 23.45 4.515 ;
        RECT 23.74 4.345 23.91 4.515 ;
        RECT 24.2 4.345 24.37 4.515 ;
        RECT 24.66 4.345 24.83 4.515 ;
        RECT 25.12 4.345 25.29 4.515 ;
        RECT 25.58 4.345 25.75 4.515 ;
        RECT 26.04 4.345 26.21 4.515 ;
        RECT 26.5 4.345 26.67 4.515 ;
        RECT 26.96 4.345 27.13 4.515 ;
        RECT 27.42 4.345 27.59 4.515 ;
        RECT 31.225 4.545 31.395 4.715 ;
        RECT 31.225 4.165 31.395 4.335 ;
        RECT 31.925 4.55 32.095 4.72 ;
        RECT 31.925 4.16 32.095 4.33 ;
        RECT 32.915 4.55 33.085 4.72 ;
        RECT 32.915 4.16 33.085 4.33 ;
        RECT 36.76 4.545 36.93 4.715 ;
        RECT 37.74 4.345 37.91 4.515 ;
        RECT 38.2 4.345 38.37 4.515 ;
        RECT 38.66 4.345 38.83 4.515 ;
        RECT 39.12 4.345 39.29 4.515 ;
        RECT 39.58 4.345 39.75 4.515 ;
        RECT 40.04 4.345 40.21 4.515 ;
        RECT 40.5 4.345 40.67 4.515 ;
        RECT 40.96 4.345 41.13 4.515 ;
        RECT 41.42 4.345 41.59 4.515 ;
        RECT 41.88 4.345 42.05 4.515 ;
        RECT 42.34 4.345 42.51 4.515 ;
        RECT 42.8 4.345 42.97 4.515 ;
        RECT 43.26 4.345 43.43 4.515 ;
        RECT 43.72 4.345 43.89 4.515 ;
        RECT 44.18 4.345 44.35 4.515 ;
        RECT 44.64 4.345 44.81 4.515 ;
        RECT 48.445 4.545 48.615 4.715 ;
        RECT 48.445 4.165 48.615 4.335 ;
        RECT 49.145 4.55 49.315 4.72 ;
        RECT 49.145 4.16 49.315 4.33 ;
        RECT 50.135 4.55 50.305 4.72 ;
        RECT 50.135 4.16 50.305 4.33 ;
        RECT 53.98 4.545 54.15 4.715 ;
        RECT 54.96 4.345 55.13 4.515 ;
        RECT 55.42 4.345 55.59 4.515 ;
        RECT 55.88 4.345 56.05 4.515 ;
        RECT 56.34 4.345 56.51 4.515 ;
        RECT 56.8 4.345 56.97 4.515 ;
        RECT 57.26 4.345 57.43 4.515 ;
        RECT 57.72 4.345 57.89 4.515 ;
        RECT 58.18 4.345 58.35 4.515 ;
        RECT 58.64 4.345 58.81 4.515 ;
        RECT 59.1 4.345 59.27 4.515 ;
        RECT 59.56 4.345 59.73 4.515 ;
        RECT 60.02 4.345 60.19 4.515 ;
        RECT 60.48 4.345 60.65 4.515 ;
        RECT 60.94 4.345 61.11 4.515 ;
        RECT 61.4 4.345 61.57 4.515 ;
        RECT 61.86 4.345 62.03 4.515 ;
        RECT 65.665 4.545 65.835 4.715 ;
        RECT 65.665 4.165 65.835 4.335 ;
        RECT 66.365 4.55 66.535 4.72 ;
        RECT 66.365 4.16 66.535 4.33 ;
        RECT 67.355 4.55 67.525 4.72 ;
        RECT 67.355 4.16 67.525 4.33 ;
        RECT 71.2 4.545 71.37 4.715 ;
        RECT 72.18 4.345 72.35 4.515 ;
        RECT 72.64 4.345 72.81 4.515 ;
        RECT 73.1 4.345 73.27 4.515 ;
        RECT 73.56 4.345 73.73 4.515 ;
        RECT 74.02 4.345 74.19 4.515 ;
        RECT 74.48 4.345 74.65 4.515 ;
        RECT 74.94 4.345 75.11 4.515 ;
        RECT 75.4 4.345 75.57 4.515 ;
        RECT 75.86 4.345 76.03 4.515 ;
        RECT 76.32 4.345 76.49 4.515 ;
        RECT 76.78 4.345 76.95 4.515 ;
        RECT 77.24 4.345 77.41 4.515 ;
        RECT 77.7 4.345 77.87 4.515 ;
        RECT 78.16 4.345 78.33 4.515 ;
        RECT 78.62 4.345 78.79 4.515 ;
        RECT 79.08 4.345 79.25 4.515 ;
        RECT 82.885 4.545 83.055 4.715 ;
        RECT 82.885 4.165 83.055 4.335 ;
        RECT 83.585 4.55 83.755 4.72 ;
        RECT 83.585 4.16 83.755 4.33 ;
        RECT 84.575 4.55 84.745 4.72 ;
        RECT 84.575 4.16 84.745 4.33 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 74.42 5.79 74.75 6.12 ;
        RECT 73.95 5.805 74.75 6.105 ;
        RECT 57.2 5.79 57.53 6.12 ;
        RECT 56.73 5.805 57.53 6.105 ;
        RECT 39.98 5.79 40.31 6.12 ;
        RECT 39.51 5.805 40.31 6.105 ;
        RECT 22.76 5.79 23.09 6.12 ;
        RECT 22.29 5.805 23.09 6.105 ;
        RECT 5.54 5.79 5.87 6.12 ;
        RECT 5.07 5.805 5.87 6.105 ;
      LAYER li1 ;
        RECT 85.29 0 85.47 0.305 ;
        RECT -3.43 0 85.47 0.3 ;
        RECT 84.495 0 84.665 0.93 ;
        RECT 83.505 0 83.675 0.93 ;
        RECT 68.07 0 83.34 0.305 ;
        RECT 80.765 0 80.935 0.935 ;
        RECT 72.035 0 79.69 1.795 ;
        RECT 78.93 0 79.26 2.185 ;
        RECT 78.09 0 78.42 2.185 ;
        RECT 76.26 0 76.55 2.63 ;
        RECT 75.81 0 76.08 2.605 ;
        RECT 74.9 0 75.14 2.605 ;
        RECT 74.45 0 74.69 2.605 ;
        RECT 73.51 0 73.78 2.605 ;
        RECT 73.06 0 73.29 2.615 ;
        RECT 72.18 0 72.39 2.615 ;
        RECT 72.03 0 79.69 1.635 ;
        RECT 67.275 0 67.445 0.93 ;
        RECT 66.285 0 66.455 0.93 ;
        RECT 50.85 0 66.12 0.305 ;
        RECT 63.545 0 63.715 0.935 ;
        RECT 54.815 0 62.47 1.795 ;
        RECT 61.71 0 62.04 2.185 ;
        RECT 60.87 0 61.2 2.185 ;
        RECT 59.04 0 59.33 2.63 ;
        RECT 58.59 0 58.86 2.605 ;
        RECT 57.68 0 57.92 2.605 ;
        RECT 57.23 0 57.47 2.605 ;
        RECT 56.29 0 56.56 2.605 ;
        RECT 55.84 0 56.07 2.615 ;
        RECT 54.96 0 55.17 2.615 ;
        RECT 54.81 0 62.47 1.635 ;
        RECT 50.055 0 50.225 0.93 ;
        RECT 49.065 0 49.235 0.93 ;
        RECT 33.63 0 48.9 0.305 ;
        RECT 46.325 0 46.495 0.935 ;
        RECT 37.595 0 45.25 1.795 ;
        RECT 44.49 0 44.82 2.185 ;
        RECT 43.65 0 43.98 2.185 ;
        RECT 41.82 0 42.11 2.63 ;
        RECT 41.37 0 41.64 2.605 ;
        RECT 40.46 0 40.7 2.605 ;
        RECT 40.01 0 40.25 2.605 ;
        RECT 39.07 0 39.34 2.605 ;
        RECT 38.62 0 38.85 2.615 ;
        RECT 37.74 0 37.95 2.615 ;
        RECT 37.59 0 45.25 1.635 ;
        RECT 32.835 0 33.005 0.93 ;
        RECT 31.845 0 32.015 0.93 ;
        RECT 16.41 0 31.68 0.305 ;
        RECT 29.105 0 29.275 0.935 ;
        RECT 20.375 0 28.03 1.795 ;
        RECT 27.27 0 27.6 2.185 ;
        RECT 26.43 0 26.76 2.185 ;
        RECT 24.6 0 24.89 2.63 ;
        RECT 24.15 0 24.42 2.605 ;
        RECT 23.24 0 23.48 2.605 ;
        RECT 22.79 0 23.03 2.605 ;
        RECT 21.85 0 22.12 2.605 ;
        RECT 21.4 0 21.63 2.615 ;
        RECT 20.52 0 20.73 2.615 ;
        RECT 20.37 0 28.03 1.635 ;
        RECT 15.615 0 15.785 0.93 ;
        RECT 14.625 0 14.795 0.93 ;
        RECT -3.43 0 14.46 0.305 ;
        RECT 11.885 0 12.055 0.935 ;
        RECT 3.155 0 10.81 1.795 ;
        RECT 10.05 0 10.38 2.185 ;
        RECT 9.21 0 9.54 2.185 ;
        RECT 7.38 0 7.67 2.63 ;
        RECT 6.93 0 7.2 2.605 ;
        RECT 6.02 0 6.26 2.605 ;
        RECT 5.57 0 5.81 2.605 ;
        RECT 4.63 0 4.9 2.605 ;
        RECT 4.18 0 4.41 2.615 ;
        RECT 3.3 0 3.51 2.615 ;
        RECT 3.15 0 10.81 1.635 ;
        RECT -3.43 8.58 85.47 8.88 ;
        RECT 85.29 8.575 85.47 8.88 ;
        RECT 84.495 7.95 84.665 8.88 ;
        RECT 83.505 7.95 83.675 8.88 ;
        RECT 68.07 8.575 83.34 8.88 ;
        RECT 80.765 7.945 80.935 8.88 ;
        RECT 72.305 7.18 79.505 8.88 ;
        RECT 72.035 7.065 79.395 7.235 ;
        RECT 78.54 6.265 78.85 8.88 ;
        RECT 77.16 6.265 77.47 8.88 ;
        RECT 74.89 5.825 75.225 6.095 ;
        RECT 74.88 6.265 75.19 8.88 ;
        RECT 74.5 5.875 75.225 6.045 ;
        RECT 74.51 5.875 74.68 8.88 ;
        RECT 72.58 6.265 72.89 8.88 ;
        RECT 69.08 7.945 69.25 8.88 ;
        RECT 67.275 7.95 67.445 8.88 ;
        RECT 66.285 7.95 66.455 8.88 ;
        RECT 50.85 8.575 66.12 8.88 ;
        RECT 63.545 7.945 63.715 8.88 ;
        RECT 55.085 7.18 62.285 8.88 ;
        RECT 54.815 7.065 62.175 7.235 ;
        RECT 61.32 6.265 61.63 8.88 ;
        RECT 59.94 6.265 60.25 8.88 ;
        RECT 57.67 5.825 58.005 6.095 ;
        RECT 57.66 6.265 57.97 8.88 ;
        RECT 57.28 5.875 58.005 6.045 ;
        RECT 57.29 5.875 57.46 8.88 ;
        RECT 55.36 6.265 55.67 8.88 ;
        RECT 51.86 7.945 52.03 8.88 ;
        RECT 50.055 7.95 50.225 8.88 ;
        RECT 49.065 7.95 49.235 8.88 ;
        RECT 33.63 8.575 48.9 8.88 ;
        RECT 46.325 7.945 46.495 8.88 ;
        RECT 37.865 7.18 45.065 8.88 ;
        RECT 37.595 7.065 44.955 7.235 ;
        RECT 44.1 6.265 44.41 8.88 ;
        RECT 42.72 6.265 43.03 8.88 ;
        RECT 40.45 5.825 40.785 6.095 ;
        RECT 40.44 6.265 40.75 8.88 ;
        RECT 40.06 5.875 40.785 6.045 ;
        RECT 40.07 5.875 40.24 8.88 ;
        RECT 38.14 6.265 38.45 8.88 ;
        RECT 34.64 7.945 34.81 8.88 ;
        RECT 32.835 7.95 33.005 8.88 ;
        RECT 31.845 7.95 32.015 8.88 ;
        RECT 16.41 8.575 31.68 8.88 ;
        RECT 29.105 7.945 29.275 8.88 ;
        RECT 20.645 7.18 27.845 8.88 ;
        RECT 20.375 7.065 27.735 7.235 ;
        RECT 26.88 6.265 27.19 8.88 ;
        RECT 25.5 6.265 25.81 8.88 ;
        RECT 23.23 5.825 23.565 6.095 ;
        RECT 23.22 6.265 23.53 8.88 ;
        RECT 22.84 5.875 23.565 6.045 ;
        RECT 22.85 5.875 23.02 8.88 ;
        RECT 20.92 6.265 21.23 8.88 ;
        RECT 17.42 7.945 17.59 8.88 ;
        RECT 15.615 7.95 15.785 8.88 ;
        RECT 14.625 7.95 14.795 8.88 ;
        RECT -3.43 8.575 14.46 8.88 ;
        RECT 11.885 7.945 12.055 8.88 ;
        RECT 3.425 7.18 10.625 8.88 ;
        RECT 3.155 7.065 10.515 7.235 ;
        RECT 9.66 6.265 9.97 8.88 ;
        RECT 8.28 6.265 8.59 8.88 ;
        RECT 6.01 5.825 6.345 6.095 ;
        RECT 6 6.265 6.31 8.88 ;
        RECT 5.62 5.875 6.345 6.045 ;
        RECT 5.63 5.875 5.8 8.88 ;
        RECT 3.7 6.265 4.01 8.88 ;
        RECT 0.2 7.945 0.37 8.88 ;
        RECT -3.21 7.945 -3.04 8.88 ;
        RECT 72.59 5.825 72.925 6.095 ;
        RECT 72.12 5.875 72.925 6.045 ;
        RECT 70.085 6.075 70.255 8.025 ;
        RECT 70.03 7.855 70.2 8.305 ;
        RECT 70.03 5.015 70.2 6.245 ;
        RECT 55.37 5.825 55.705 6.095 ;
        RECT 54.9 5.875 55.705 6.045 ;
        RECT 52.865 6.075 53.035 8.025 ;
        RECT 52.81 7.855 52.98 8.305 ;
        RECT 52.81 5.015 52.98 6.245 ;
        RECT 38.15 5.825 38.485 6.095 ;
        RECT 37.68 5.875 38.485 6.045 ;
        RECT 35.645 6.075 35.815 8.025 ;
        RECT 35.59 7.855 35.76 8.305 ;
        RECT 35.59 5.015 35.76 6.245 ;
        RECT 20.93 5.825 21.265 6.095 ;
        RECT 20.46 5.875 21.265 6.045 ;
        RECT 18.425 6.075 18.595 8.025 ;
        RECT 18.37 7.855 18.54 8.305 ;
        RECT 18.37 5.015 18.54 6.245 ;
        RECT 3.71 5.825 4.045 6.095 ;
        RECT 3.24 5.875 4.045 6.045 ;
        RECT 1.205 6.075 1.375 8.025 ;
        RECT 1.15 7.855 1.32 8.305 ;
        RECT 1.15 5.015 1.32 6.245 ;
      LAYER met2 ;
        RECT 74.445 5.77 74.725 6.14 ;
        RECT 57.225 5.77 57.505 6.14 ;
        RECT 40.005 5.77 40.285 6.14 ;
        RECT 22.785 5.77 23.065 6.14 ;
        RECT 5.565 5.77 5.845 6.14 ;
      LAYER met1 ;
        RECT 85.29 0 85.47 0.305 ;
        RECT -3.43 0 85.47 0.3 ;
        RECT 68.07 0 83.34 0.305 ;
        RECT 72.035 0 79.69 1.795 ;
        RECT 72.035 0 79.395 1.95 ;
        RECT 72.03 0 79.69 1.635 ;
        RECT 50.85 0 66.12 0.305 ;
        RECT 54.815 0 62.47 1.795 ;
        RECT 54.815 0 62.175 1.95 ;
        RECT 54.81 0 62.47 1.635 ;
        RECT 33.63 0 48.9 0.305 ;
        RECT 37.595 0 45.25 1.795 ;
        RECT 37.595 0 44.955 1.95 ;
        RECT 37.59 0 45.25 1.635 ;
        RECT 16.41 0 31.68 0.305 ;
        RECT 20.375 0 28.03 1.795 ;
        RECT 20.375 0 27.735 1.95 ;
        RECT 20.37 0 28.03 1.635 ;
        RECT -3.43 0 14.46 0.305 ;
        RECT 3.155 0 10.81 1.795 ;
        RECT 3.155 0 10.515 1.95 ;
        RECT 3.15 0 10.81 1.635 ;
        RECT -3.43 8.58 85.47 8.88 ;
        RECT 85.29 8.575 85.47 8.88 ;
        RECT 68.07 8.575 83.34 8.88 ;
        RECT 72.305 7.18 79.505 8.88 ;
        RECT 72.035 6.91 79.395 7.39 ;
        RECT 70.025 6.285 70.315 6.515 ;
        RECT 69.625 6.315 70.315 6.485 ;
        RECT 69.625 6.315 69.795 8.88 ;
        RECT 50.85 8.575 66.12 8.88 ;
        RECT 55.085 7.18 62.285 8.88 ;
        RECT 54.815 6.91 62.175 7.39 ;
        RECT 52.805 6.285 53.095 6.515 ;
        RECT 52.405 6.315 53.095 6.485 ;
        RECT 52.405 6.315 52.575 8.88 ;
        RECT 33.63 8.575 48.9 8.88 ;
        RECT 37.865 7.18 45.065 8.88 ;
        RECT 37.595 6.91 44.955 7.39 ;
        RECT 35.585 6.285 35.875 6.515 ;
        RECT 35.185 6.315 35.875 6.485 ;
        RECT 35.185 6.315 35.355 8.88 ;
        RECT 16.41 8.575 31.68 8.88 ;
        RECT 20.645 7.18 27.845 8.88 ;
        RECT 20.375 6.91 27.735 7.39 ;
        RECT 18.365 6.285 18.655 6.515 ;
        RECT 17.965 6.315 18.655 6.485 ;
        RECT 17.965 6.315 18.135 8.88 ;
        RECT -3.43 8.575 14.46 8.88 ;
        RECT 3.425 7.18 10.625 8.88 ;
        RECT 3.155 6.91 10.515 7.39 ;
        RECT 1.145 6.285 1.435 6.515 ;
        RECT 0.745 6.315 1.435 6.485 ;
        RECT 0.745 6.315 0.915 8.88 ;
        RECT 74.425 5.83 74.745 6.09 ;
        RECT 72.06 5.89 74.745 6.03 ;
        RECT 72.06 5.845 72.35 6.075 ;
        RECT 57.205 5.83 57.525 6.09 ;
        RECT 54.84 5.89 57.525 6.03 ;
        RECT 54.84 5.845 55.13 6.075 ;
        RECT 39.985 5.83 40.305 6.09 ;
        RECT 37.62 5.89 40.305 6.03 ;
        RECT 37.62 5.845 37.91 6.075 ;
        RECT 22.765 5.83 23.085 6.09 ;
        RECT 20.4 5.89 23.085 6.03 ;
        RECT 20.4 5.845 20.69 6.075 ;
        RECT 5.545 5.83 5.865 6.09 ;
        RECT 3.18 5.89 5.865 6.03 ;
        RECT 3.18 5.845 3.47 6.075 ;
      LAYER via2 ;
        RECT 5.605 5.855 5.805 6.055 ;
        RECT 22.825 5.855 23.025 6.055 ;
        RECT 40.045 5.855 40.245 6.055 ;
        RECT 57.265 5.855 57.465 6.055 ;
        RECT 74.485 5.855 74.685 6.055 ;
      LAYER via1 ;
        RECT 5.63 5.885 5.78 6.035 ;
        RECT 22.85 5.885 23 6.035 ;
        RECT 40.07 5.885 40.22 6.035 ;
        RECT 57.29 5.885 57.44 6.035 ;
        RECT 74.51 5.885 74.66 6.035 ;
      LAYER mcon ;
        RECT -3.13 8.605 -2.96 8.775 ;
        RECT -2.45 8.605 -2.28 8.775 ;
        RECT -1.77 8.605 -1.6 8.775 ;
        RECT -1.09 8.605 -0.92 8.775 ;
        RECT 0.28 8.605 0.45 8.775 ;
        RECT 0.96 8.605 1.13 8.775 ;
        RECT 1.205 6.315 1.375 6.485 ;
        RECT 1.64 8.605 1.81 8.775 ;
        RECT 2.32 8.605 2.49 8.775 ;
        RECT 3.24 5.875 3.41 6.045 ;
        RECT 3.3 7.065 3.47 7.235 ;
        RECT 3.3 1.625 3.47 1.795 ;
        RECT 3.76 7.065 3.93 7.235 ;
        RECT 3.76 1.625 3.93 1.795 ;
        RECT 4.22 7.065 4.39 7.235 ;
        RECT 4.22 1.625 4.39 1.795 ;
        RECT 4.68 7.065 4.85 7.235 ;
        RECT 4.68 1.625 4.85 1.795 ;
        RECT 5.14 7.065 5.31 7.235 ;
        RECT 5.14 1.625 5.31 1.795 ;
        RECT 5.6 7.065 5.77 7.235 ;
        RECT 5.6 1.625 5.77 1.795 ;
        RECT 5.62 5.875 5.79 6.045 ;
        RECT 6.06 7.065 6.23 7.235 ;
        RECT 6.06 1.625 6.23 1.795 ;
        RECT 6.52 7.065 6.69 7.235 ;
        RECT 6.52 1.625 6.69 1.795 ;
        RECT 6.98 7.065 7.15 7.235 ;
        RECT 6.98 1.625 7.15 1.795 ;
        RECT 7.44 7.065 7.61 7.235 ;
        RECT 7.44 1.625 7.61 1.795 ;
        RECT 7.9 7.065 8.07 7.235 ;
        RECT 7.9 1.625 8.07 1.795 ;
        RECT 8.36 7.065 8.53 7.235 ;
        RECT 8.36 1.625 8.53 1.795 ;
        RECT 8.82 7.065 8.99 7.235 ;
        RECT 8.82 1.625 8.99 1.795 ;
        RECT 9.28 7.065 9.45 7.235 ;
        RECT 9.28 1.625 9.45 1.795 ;
        RECT 9.74 7.065 9.91 7.235 ;
        RECT 9.74 1.625 9.91 1.795 ;
        RECT 10.2 7.065 10.37 7.235 ;
        RECT 10.2 1.625 10.37 1.795 ;
        RECT 11.965 8.605 12.135 8.775 ;
        RECT 11.965 0.105 12.135 0.275 ;
        RECT 12.645 8.605 12.815 8.775 ;
        RECT 12.645 0.105 12.815 0.275 ;
        RECT 13.325 8.605 13.495 8.775 ;
        RECT 13.325 0.105 13.495 0.275 ;
        RECT 14.005 8.605 14.175 8.775 ;
        RECT 14.005 0.105 14.175 0.275 ;
        RECT 14.705 8.61 14.875 8.78 ;
        RECT 14.705 0.1 14.875 0.27 ;
        RECT 15.695 8.61 15.865 8.78 ;
        RECT 15.695 0.1 15.865 0.27 ;
        RECT 17.5 8.605 17.67 8.775 ;
        RECT 18.18 8.605 18.35 8.775 ;
        RECT 18.425 6.315 18.595 6.485 ;
        RECT 18.86 8.605 19.03 8.775 ;
        RECT 19.54 8.605 19.71 8.775 ;
        RECT 20.46 5.875 20.63 6.045 ;
        RECT 20.52 7.065 20.69 7.235 ;
        RECT 20.52 1.625 20.69 1.795 ;
        RECT 20.98 7.065 21.15 7.235 ;
        RECT 20.98 1.625 21.15 1.795 ;
        RECT 21.44 7.065 21.61 7.235 ;
        RECT 21.44 1.625 21.61 1.795 ;
        RECT 21.9 7.065 22.07 7.235 ;
        RECT 21.9 1.625 22.07 1.795 ;
        RECT 22.36 7.065 22.53 7.235 ;
        RECT 22.36 1.625 22.53 1.795 ;
        RECT 22.82 7.065 22.99 7.235 ;
        RECT 22.82 1.625 22.99 1.795 ;
        RECT 22.84 5.875 23.01 6.045 ;
        RECT 23.28 7.065 23.45 7.235 ;
        RECT 23.28 1.625 23.45 1.795 ;
        RECT 23.74 7.065 23.91 7.235 ;
        RECT 23.74 1.625 23.91 1.795 ;
        RECT 24.2 7.065 24.37 7.235 ;
        RECT 24.2 1.625 24.37 1.795 ;
        RECT 24.66 7.065 24.83 7.235 ;
        RECT 24.66 1.625 24.83 1.795 ;
        RECT 25.12 7.065 25.29 7.235 ;
        RECT 25.12 1.625 25.29 1.795 ;
        RECT 25.58 7.065 25.75 7.235 ;
        RECT 25.58 1.625 25.75 1.795 ;
        RECT 26.04 7.065 26.21 7.235 ;
        RECT 26.04 1.625 26.21 1.795 ;
        RECT 26.5 7.065 26.67 7.235 ;
        RECT 26.5 1.625 26.67 1.795 ;
        RECT 26.96 7.065 27.13 7.235 ;
        RECT 26.96 1.625 27.13 1.795 ;
        RECT 27.42 7.065 27.59 7.235 ;
        RECT 27.42 1.625 27.59 1.795 ;
        RECT 29.185 8.605 29.355 8.775 ;
        RECT 29.185 0.105 29.355 0.275 ;
        RECT 29.865 8.605 30.035 8.775 ;
        RECT 29.865 0.105 30.035 0.275 ;
        RECT 30.545 8.605 30.715 8.775 ;
        RECT 30.545 0.105 30.715 0.275 ;
        RECT 31.225 8.605 31.395 8.775 ;
        RECT 31.225 0.105 31.395 0.275 ;
        RECT 31.925 8.61 32.095 8.78 ;
        RECT 31.925 0.1 32.095 0.27 ;
        RECT 32.915 8.61 33.085 8.78 ;
        RECT 32.915 0.1 33.085 0.27 ;
        RECT 34.72 8.605 34.89 8.775 ;
        RECT 35.4 8.605 35.57 8.775 ;
        RECT 35.645 6.315 35.815 6.485 ;
        RECT 36.08 8.605 36.25 8.775 ;
        RECT 36.76 8.605 36.93 8.775 ;
        RECT 37.68 5.875 37.85 6.045 ;
        RECT 37.74 7.065 37.91 7.235 ;
        RECT 37.74 1.625 37.91 1.795 ;
        RECT 38.2 7.065 38.37 7.235 ;
        RECT 38.2 1.625 38.37 1.795 ;
        RECT 38.66 7.065 38.83 7.235 ;
        RECT 38.66 1.625 38.83 1.795 ;
        RECT 39.12 7.065 39.29 7.235 ;
        RECT 39.12 1.625 39.29 1.795 ;
        RECT 39.58 7.065 39.75 7.235 ;
        RECT 39.58 1.625 39.75 1.795 ;
        RECT 40.04 7.065 40.21 7.235 ;
        RECT 40.04 1.625 40.21 1.795 ;
        RECT 40.06 5.875 40.23 6.045 ;
        RECT 40.5 7.065 40.67 7.235 ;
        RECT 40.5 1.625 40.67 1.795 ;
        RECT 40.96 7.065 41.13 7.235 ;
        RECT 40.96 1.625 41.13 1.795 ;
        RECT 41.42 7.065 41.59 7.235 ;
        RECT 41.42 1.625 41.59 1.795 ;
        RECT 41.88 7.065 42.05 7.235 ;
        RECT 41.88 1.625 42.05 1.795 ;
        RECT 42.34 7.065 42.51 7.235 ;
        RECT 42.34 1.625 42.51 1.795 ;
        RECT 42.8 7.065 42.97 7.235 ;
        RECT 42.8 1.625 42.97 1.795 ;
        RECT 43.26 7.065 43.43 7.235 ;
        RECT 43.26 1.625 43.43 1.795 ;
        RECT 43.72 7.065 43.89 7.235 ;
        RECT 43.72 1.625 43.89 1.795 ;
        RECT 44.18 7.065 44.35 7.235 ;
        RECT 44.18 1.625 44.35 1.795 ;
        RECT 44.64 7.065 44.81 7.235 ;
        RECT 44.64 1.625 44.81 1.795 ;
        RECT 46.405 8.605 46.575 8.775 ;
        RECT 46.405 0.105 46.575 0.275 ;
        RECT 47.085 8.605 47.255 8.775 ;
        RECT 47.085 0.105 47.255 0.275 ;
        RECT 47.765 8.605 47.935 8.775 ;
        RECT 47.765 0.105 47.935 0.275 ;
        RECT 48.445 8.605 48.615 8.775 ;
        RECT 48.445 0.105 48.615 0.275 ;
        RECT 49.145 8.61 49.315 8.78 ;
        RECT 49.145 0.1 49.315 0.27 ;
        RECT 50.135 8.61 50.305 8.78 ;
        RECT 50.135 0.1 50.305 0.27 ;
        RECT 51.94 8.605 52.11 8.775 ;
        RECT 52.62 8.605 52.79 8.775 ;
        RECT 52.865 6.315 53.035 6.485 ;
        RECT 53.3 8.605 53.47 8.775 ;
        RECT 53.98 8.605 54.15 8.775 ;
        RECT 54.9 5.875 55.07 6.045 ;
        RECT 54.96 7.065 55.13 7.235 ;
        RECT 54.96 1.625 55.13 1.795 ;
        RECT 55.42 7.065 55.59 7.235 ;
        RECT 55.42 1.625 55.59 1.795 ;
        RECT 55.88 7.065 56.05 7.235 ;
        RECT 55.88 1.625 56.05 1.795 ;
        RECT 56.34 7.065 56.51 7.235 ;
        RECT 56.34 1.625 56.51 1.795 ;
        RECT 56.8 7.065 56.97 7.235 ;
        RECT 56.8 1.625 56.97 1.795 ;
        RECT 57.26 7.065 57.43 7.235 ;
        RECT 57.26 1.625 57.43 1.795 ;
        RECT 57.28 5.875 57.45 6.045 ;
        RECT 57.72 7.065 57.89 7.235 ;
        RECT 57.72 1.625 57.89 1.795 ;
        RECT 58.18 7.065 58.35 7.235 ;
        RECT 58.18 1.625 58.35 1.795 ;
        RECT 58.64 7.065 58.81 7.235 ;
        RECT 58.64 1.625 58.81 1.795 ;
        RECT 59.1 7.065 59.27 7.235 ;
        RECT 59.1 1.625 59.27 1.795 ;
        RECT 59.56 7.065 59.73 7.235 ;
        RECT 59.56 1.625 59.73 1.795 ;
        RECT 60.02 7.065 60.19 7.235 ;
        RECT 60.02 1.625 60.19 1.795 ;
        RECT 60.48 7.065 60.65 7.235 ;
        RECT 60.48 1.625 60.65 1.795 ;
        RECT 60.94 7.065 61.11 7.235 ;
        RECT 60.94 1.625 61.11 1.795 ;
        RECT 61.4 7.065 61.57 7.235 ;
        RECT 61.4 1.625 61.57 1.795 ;
        RECT 61.86 7.065 62.03 7.235 ;
        RECT 61.86 1.625 62.03 1.795 ;
        RECT 63.625 8.605 63.795 8.775 ;
        RECT 63.625 0.105 63.795 0.275 ;
        RECT 64.305 8.605 64.475 8.775 ;
        RECT 64.305 0.105 64.475 0.275 ;
        RECT 64.985 8.605 65.155 8.775 ;
        RECT 64.985 0.105 65.155 0.275 ;
        RECT 65.665 8.605 65.835 8.775 ;
        RECT 65.665 0.105 65.835 0.275 ;
        RECT 66.365 8.61 66.535 8.78 ;
        RECT 66.365 0.1 66.535 0.27 ;
        RECT 67.355 8.61 67.525 8.78 ;
        RECT 67.355 0.1 67.525 0.27 ;
        RECT 69.16 8.605 69.33 8.775 ;
        RECT 69.84 8.605 70.01 8.775 ;
        RECT 70.085 6.315 70.255 6.485 ;
        RECT 70.52 8.605 70.69 8.775 ;
        RECT 71.2 8.605 71.37 8.775 ;
        RECT 72.12 5.875 72.29 6.045 ;
        RECT 72.18 7.065 72.35 7.235 ;
        RECT 72.18 1.625 72.35 1.795 ;
        RECT 72.64 7.065 72.81 7.235 ;
        RECT 72.64 1.625 72.81 1.795 ;
        RECT 73.1 7.065 73.27 7.235 ;
        RECT 73.1 1.625 73.27 1.795 ;
        RECT 73.56 7.065 73.73 7.235 ;
        RECT 73.56 1.625 73.73 1.795 ;
        RECT 74.02 7.065 74.19 7.235 ;
        RECT 74.02 1.625 74.19 1.795 ;
        RECT 74.48 7.065 74.65 7.235 ;
        RECT 74.48 1.625 74.65 1.795 ;
        RECT 74.5 5.875 74.67 6.045 ;
        RECT 74.94 7.065 75.11 7.235 ;
        RECT 74.94 1.625 75.11 1.795 ;
        RECT 75.4 7.065 75.57 7.235 ;
        RECT 75.4 1.625 75.57 1.795 ;
        RECT 75.86 7.065 76.03 7.235 ;
        RECT 75.86 1.625 76.03 1.795 ;
        RECT 76.32 7.065 76.49 7.235 ;
        RECT 76.32 1.625 76.49 1.795 ;
        RECT 76.78 7.065 76.95 7.235 ;
        RECT 76.78 1.625 76.95 1.795 ;
        RECT 77.24 7.065 77.41 7.235 ;
        RECT 77.24 1.625 77.41 1.795 ;
        RECT 77.7 7.065 77.87 7.235 ;
        RECT 77.7 1.625 77.87 1.795 ;
        RECT 78.16 7.065 78.33 7.235 ;
        RECT 78.16 1.625 78.33 1.795 ;
        RECT 78.62 7.065 78.79 7.235 ;
        RECT 78.62 1.625 78.79 1.795 ;
        RECT 79.08 7.065 79.25 7.235 ;
        RECT 79.08 1.625 79.25 1.795 ;
        RECT 80.845 8.605 81.015 8.775 ;
        RECT 80.845 0.105 81.015 0.275 ;
        RECT 81.525 8.605 81.695 8.775 ;
        RECT 81.525 0.105 81.695 0.275 ;
        RECT 82.205 8.605 82.375 8.775 ;
        RECT 82.205 0.105 82.375 0.275 ;
        RECT 82.885 8.605 83.055 8.775 ;
        RECT 82.885 0.105 83.055 0.275 ;
        RECT 83.585 8.61 83.755 8.78 ;
        RECT 83.585 0.1 83.755 0.27 ;
        RECT 84.575 8.61 84.745 8.78 ;
        RECT 84.575 0.1 84.745 0.27 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 71.5 7.435 77.515 7.735 ;
      RECT 77.215 5.805 77.515 7.735 ;
      RECT 76.16 5.785 76.46 7.735 ;
      RECT 75.13 6.48 75.43 7.735 ;
      RECT 71.5 7.035 71.8 7.735 ;
      RECT 70.365 7 70.735 7.37 ;
      RECT 70.365 7.035 71.8 7.335 ;
      RECT 75.1 6.48 75.43 6.81 ;
      RECT 74.63 6.495 75.43 6.795 ;
      RECT 75.01 6.455 75.31 6.795 ;
      RECT 77.14 5.805 77.515 6.17 ;
      RECT 77.205 5.765 77.505 6.17 ;
      RECT 76.12 5.785 76.46 6.135 ;
      RECT 76.135 5.745 76.435 6.135 ;
      RECT 76.11 5.79 76.46 6.12 ;
      RECT 77.14 5.805 77.95 6.105 ;
      RECT 75.64 5.805 76.46 6.105 ;
      RECT 77.15 5.79 77.505 6.17 ;
      RECT 76.8 3.755 77.13 4.085 ;
      RECT 76.8 3.77 77.6 4.07 ;
      RECT 76.815 3.725 77.115 4.085 ;
      RECT 76.46 3.075 76.79 3.405 ;
      RECT 76.46 3.09 77.26 3.39 ;
      RECT 76.545 3.065 76.845 3.39 ;
      RECT 75.78 4.155 76.11 4.485 ;
      RECT 73.74 4.155 74.07 4.485 ;
      RECT 73.74 4.17 76.11 4.47 ;
      RECT 75.43 3.415 75.76 3.745 ;
      RECT 74.97 3.43 75.77 3.73 ;
      RECT 75.1 2.225 75.43 2.555 ;
      RECT 74.63 2.24 75.43 2.54 ;
      RECT 75.09 2.235 75.43 2.54 ;
      RECT 54.28 7.435 60.295 7.735 ;
      RECT 59.995 5.805 60.295 7.735 ;
      RECT 58.94 5.785 59.24 7.735 ;
      RECT 57.91 6.48 58.21 7.735 ;
      RECT 54.28 7.035 54.58 7.735 ;
      RECT 53.145 7 53.515 7.37 ;
      RECT 53.145 7.035 54.58 7.335 ;
      RECT 57.88 6.48 58.21 6.81 ;
      RECT 57.41 6.495 58.21 6.795 ;
      RECT 57.79 6.455 58.09 6.795 ;
      RECT 59.92 5.805 60.295 6.17 ;
      RECT 59.985 5.765 60.285 6.17 ;
      RECT 58.9 5.785 59.24 6.135 ;
      RECT 58.915 5.745 59.215 6.135 ;
      RECT 58.89 5.79 59.24 6.12 ;
      RECT 59.92 5.805 60.73 6.105 ;
      RECT 58.42 5.805 59.24 6.105 ;
      RECT 59.93 5.79 60.285 6.17 ;
      RECT 59.58 3.755 59.91 4.085 ;
      RECT 59.58 3.77 60.38 4.07 ;
      RECT 59.595 3.725 59.895 4.085 ;
      RECT 59.24 3.075 59.57 3.405 ;
      RECT 59.24 3.09 60.04 3.39 ;
      RECT 59.325 3.065 59.625 3.39 ;
      RECT 58.56 4.155 58.89 4.485 ;
      RECT 56.52 4.155 56.85 4.485 ;
      RECT 56.52 4.17 58.89 4.47 ;
      RECT 58.21 3.415 58.54 3.745 ;
      RECT 57.75 3.43 58.55 3.73 ;
      RECT 57.88 2.225 58.21 2.555 ;
      RECT 57.41 2.24 58.21 2.54 ;
      RECT 57.87 2.235 58.21 2.54 ;
      RECT 37.06 7.435 43.075 7.735 ;
      RECT 42.775 5.805 43.075 7.735 ;
      RECT 41.72 5.785 42.02 7.735 ;
      RECT 40.69 6.48 40.99 7.735 ;
      RECT 37.06 7.035 37.36 7.735 ;
      RECT 35.925 7 36.295 7.37 ;
      RECT 35.925 7.035 37.36 7.335 ;
      RECT 40.66 6.48 40.99 6.81 ;
      RECT 40.19 6.495 40.99 6.795 ;
      RECT 40.57 6.455 40.87 6.795 ;
      RECT 42.7 5.805 43.075 6.17 ;
      RECT 42.765 5.765 43.065 6.17 ;
      RECT 41.68 5.785 42.02 6.135 ;
      RECT 41.695 5.745 41.995 6.135 ;
      RECT 41.67 5.79 42.02 6.12 ;
      RECT 42.7 5.805 43.51 6.105 ;
      RECT 41.2 5.805 42.02 6.105 ;
      RECT 42.71 5.79 43.065 6.17 ;
      RECT 42.36 3.755 42.69 4.085 ;
      RECT 42.36 3.77 43.16 4.07 ;
      RECT 42.375 3.725 42.675 4.085 ;
      RECT 42.02 3.075 42.35 3.405 ;
      RECT 42.02 3.09 42.82 3.39 ;
      RECT 42.105 3.065 42.405 3.39 ;
      RECT 41.34 4.155 41.67 4.485 ;
      RECT 39.3 4.155 39.63 4.485 ;
      RECT 39.3 4.17 41.67 4.47 ;
      RECT 40.99 3.415 41.32 3.745 ;
      RECT 40.53 3.43 41.33 3.73 ;
      RECT 40.66 2.225 40.99 2.555 ;
      RECT 40.19 2.24 40.99 2.54 ;
      RECT 40.65 2.235 40.99 2.54 ;
      RECT 19.84 7.435 25.855 7.735 ;
      RECT 25.555 5.805 25.855 7.735 ;
      RECT 24.5 5.785 24.8 7.735 ;
      RECT 23.47 6.48 23.77 7.735 ;
      RECT 19.84 7.035 20.14 7.735 ;
      RECT 18.705 7 19.075 7.37 ;
      RECT 18.705 7.035 20.14 7.335 ;
      RECT 23.44 6.48 23.77 6.81 ;
      RECT 22.97 6.495 23.77 6.795 ;
      RECT 23.35 6.455 23.65 6.795 ;
      RECT 25.48 5.805 25.855 6.17 ;
      RECT 25.545 5.765 25.845 6.17 ;
      RECT 24.46 5.785 24.8 6.135 ;
      RECT 24.475 5.745 24.775 6.135 ;
      RECT 24.45 5.79 24.8 6.12 ;
      RECT 25.48 5.805 26.29 6.105 ;
      RECT 23.98 5.805 24.8 6.105 ;
      RECT 25.49 5.79 25.845 6.17 ;
      RECT 25.14 3.755 25.47 4.085 ;
      RECT 25.14 3.77 25.94 4.07 ;
      RECT 25.155 3.725 25.455 4.085 ;
      RECT 24.8 3.075 25.13 3.405 ;
      RECT 24.8 3.09 25.6 3.39 ;
      RECT 24.885 3.065 25.185 3.39 ;
      RECT 24.12 4.155 24.45 4.485 ;
      RECT 22.08 4.155 22.41 4.485 ;
      RECT 22.08 4.17 24.45 4.47 ;
      RECT 23.77 3.415 24.1 3.745 ;
      RECT 23.31 3.43 24.11 3.73 ;
      RECT 23.44 2.225 23.77 2.555 ;
      RECT 22.97 2.24 23.77 2.54 ;
      RECT 23.43 2.235 23.77 2.54 ;
      RECT 2.62 7.435 8.635 7.735 ;
      RECT 8.335 5.805 8.635 7.735 ;
      RECT 7.28 5.785 7.58 7.735 ;
      RECT 6.25 6.48 6.55 7.735 ;
      RECT 2.62 7.035 2.92 7.735 ;
      RECT 1.485 7 1.855 7.37 ;
      RECT 1.485 7.035 2.92 7.335 ;
      RECT 6.22 6.48 6.55 6.81 ;
      RECT 5.75 6.495 6.55 6.795 ;
      RECT 6.13 6.455 6.43 6.795 ;
      RECT 8.26 5.805 8.635 6.17 ;
      RECT 8.325 5.765 8.625 6.17 ;
      RECT 7.24 5.785 7.58 6.135 ;
      RECT 7.255 5.745 7.555 6.135 ;
      RECT 7.23 5.79 7.58 6.12 ;
      RECT 8.26 5.805 9.07 6.105 ;
      RECT 6.76 5.805 7.58 6.105 ;
      RECT 8.27 5.79 8.625 6.17 ;
      RECT 7.92 3.755 8.25 4.085 ;
      RECT 7.92 3.77 8.72 4.07 ;
      RECT 7.935 3.725 8.235 4.085 ;
      RECT 7.58 3.075 7.91 3.405 ;
      RECT 7.58 3.09 8.38 3.39 ;
      RECT 7.665 3.065 7.965 3.39 ;
      RECT 6.9 4.155 7.23 4.485 ;
      RECT 4.86 4.155 5.19 4.485 ;
      RECT 4.86 4.17 7.23 4.47 ;
      RECT 6.55 3.415 6.88 3.745 ;
      RECT 6.09 3.43 6.89 3.73 ;
      RECT 6.22 2.225 6.55 2.555 ;
      RECT 5.75 2.24 6.55 2.54 ;
      RECT 6.21 2.235 6.55 2.54 ;
    LAYER via2 ;
      RECT 77.215 5.855 77.415 6.055 ;
      RECT 76.865 3.82 77.065 4.02 ;
      RECT 76.525 3.14 76.725 3.34 ;
      RECT 76.175 5.855 76.375 6.055 ;
      RECT 75.845 4.22 76.045 4.42 ;
      RECT 75.495 3.48 75.695 3.68 ;
      RECT 75.165 2.29 75.365 2.49 ;
      RECT 75.165 6.545 75.365 6.745 ;
      RECT 73.805 4.22 74.005 4.42 ;
      RECT 70.45 7.085 70.65 7.285 ;
      RECT 59.995 5.855 60.195 6.055 ;
      RECT 59.645 3.82 59.845 4.02 ;
      RECT 59.305 3.14 59.505 3.34 ;
      RECT 58.955 5.855 59.155 6.055 ;
      RECT 58.625 4.22 58.825 4.42 ;
      RECT 58.275 3.48 58.475 3.68 ;
      RECT 57.945 2.29 58.145 2.49 ;
      RECT 57.945 6.545 58.145 6.745 ;
      RECT 56.585 4.22 56.785 4.42 ;
      RECT 53.23 7.085 53.43 7.285 ;
      RECT 42.775 5.855 42.975 6.055 ;
      RECT 42.425 3.82 42.625 4.02 ;
      RECT 42.085 3.14 42.285 3.34 ;
      RECT 41.735 5.855 41.935 6.055 ;
      RECT 41.405 4.22 41.605 4.42 ;
      RECT 41.055 3.48 41.255 3.68 ;
      RECT 40.725 2.29 40.925 2.49 ;
      RECT 40.725 6.545 40.925 6.745 ;
      RECT 39.365 4.22 39.565 4.42 ;
      RECT 36.01 7.085 36.21 7.285 ;
      RECT 25.555 5.855 25.755 6.055 ;
      RECT 25.205 3.82 25.405 4.02 ;
      RECT 24.865 3.14 25.065 3.34 ;
      RECT 24.515 5.855 24.715 6.055 ;
      RECT 24.185 4.22 24.385 4.42 ;
      RECT 23.835 3.48 24.035 3.68 ;
      RECT 23.505 2.29 23.705 2.49 ;
      RECT 23.505 6.545 23.705 6.745 ;
      RECT 22.145 4.22 22.345 4.42 ;
      RECT 18.79 7.085 18.99 7.285 ;
      RECT 8.335 5.855 8.535 6.055 ;
      RECT 7.985 3.82 8.185 4.02 ;
      RECT 7.645 3.14 7.845 3.34 ;
      RECT 7.295 5.855 7.495 6.055 ;
      RECT 6.965 4.22 7.165 4.42 ;
      RECT 6.615 3.48 6.815 3.68 ;
      RECT 6.285 2.29 6.485 2.49 ;
      RECT 6.285 6.545 6.485 6.745 ;
      RECT 4.925 4.22 5.125 4.42 ;
      RECT 1.57 7.085 1.77 7.285 ;
    LAYER met2 ;
      RECT -2.22 8.6 85.1 8.77 ;
      RECT 84.93 7.3 85.1 8.77 ;
      RECT -2.22 6.255 -2.05 8.77 ;
      RECT 84.895 7.3 85.22 7.625 ;
      RECT -2.265 6.255 -1.985 6.595 ;
      RECT 81.74 6.28 82.06 6.605 ;
      RECT 81.77 5.695 81.94 6.605 ;
      RECT 81.77 5.695 81.945 6.045 ;
      RECT 81.77 5.695 82.745 5.87 ;
      RECT 82.57 1.965 82.745 5.87 ;
      RECT 75.125 2.205 75.405 2.575 ;
      RECT 75.125 2.345 79.775 2.52 ;
      RECT 79.6 2.025 79.775 2.52 ;
      RECT 80.07 1.995 80.395 2.32 ;
      RECT 82.515 1.965 82.865 2.315 ;
      RECT 79.6 2.025 82.865 2.195 ;
      RECT 70.89 8.29 81.585 8.46 ;
      RECT 81.425 2.395 81.585 8.46 ;
      RECT 70.89 6.545 71.06 8.46 ;
      RECT 82.54 6.655 82.865 6.98 ;
      RECT 67.71 6.655 68.035 6.98 ;
      RECT 81.425 6.745 82.865 6.915 ;
      RECT 70.84 6.545 71.12 6.885 ;
      RECT 67.71 6.685 71.12 6.855 ;
      RECT 81.74 2.365 82.06 2.685 ;
      RECT 81.425 2.395 82.06 2.565 ;
      RECT 78.195 6.48 78.455 6.8 ;
      RECT 78.255 2.74 78.395 6.8 ;
      RECT 78.195 2.74 78.455 3.06 ;
      RECT 77.515 4.78 77.775 5.1 ;
      RECT 77.575 3.76 77.715 5.1 ;
      RECT 77.515 3.76 77.775 4.08 ;
      RECT 76.495 6.48 76.755 6.8 ;
      RECT 76.555 5.21 76.695 6.8 ;
      RECT 75.875 5.21 76.695 5.35 ;
      RECT 75.875 2.74 76.015 5.35 ;
      RECT 75.805 4.135 76.085 4.505 ;
      RECT 75.815 2.74 76.075 3.06 ;
      RECT 73.765 4.135 74.045 4.505 ;
      RECT 73.835 2.4 73.975 4.505 ;
      RECT 73.775 2.4 74.035 2.72 ;
      RECT 73.095 4.78 73.355 5.1 ;
      RECT 73.155 2.74 73.295 5.1 ;
      RECT 73.095 2.74 73.355 3.06 ;
      RECT 64.52 6.28 64.84 6.605 ;
      RECT 64.55 5.695 64.72 6.605 ;
      RECT 64.55 5.695 64.725 6.045 ;
      RECT 64.55 5.695 65.525 5.87 ;
      RECT 65.35 1.965 65.525 5.87 ;
      RECT 57.905 2.205 58.185 2.575 ;
      RECT 57.905 2.345 62.555 2.52 ;
      RECT 62.38 2.025 62.555 2.52 ;
      RECT 62.85 1.995 63.175 2.32 ;
      RECT 65.295 1.965 65.645 2.315 ;
      RECT 62.38 2.025 65.645 2.195 ;
      RECT 53.67 8.29 64.365 8.46 ;
      RECT 64.205 2.395 64.365 8.46 ;
      RECT 53.67 6.545 53.84 8.46 ;
      RECT 65.32 6.655 65.645 6.98 ;
      RECT 50.49 6.655 50.815 6.98 ;
      RECT 64.205 6.745 65.645 6.915 ;
      RECT 53.62 6.545 53.9 6.885 ;
      RECT 50.49 6.685 53.9 6.855 ;
      RECT 64.52 2.365 64.84 2.685 ;
      RECT 64.205 2.395 64.84 2.565 ;
      RECT 60.975 6.48 61.235 6.8 ;
      RECT 61.035 2.74 61.175 6.8 ;
      RECT 60.975 2.74 61.235 3.06 ;
      RECT 60.295 4.78 60.555 5.1 ;
      RECT 60.355 3.76 60.495 5.1 ;
      RECT 60.295 3.76 60.555 4.08 ;
      RECT 59.275 6.48 59.535 6.8 ;
      RECT 59.335 5.21 59.475 6.8 ;
      RECT 58.655 5.21 59.475 5.35 ;
      RECT 58.655 2.74 58.795 5.35 ;
      RECT 58.585 4.135 58.865 4.505 ;
      RECT 58.595 2.74 58.855 3.06 ;
      RECT 56.545 4.135 56.825 4.505 ;
      RECT 56.615 2.4 56.755 4.505 ;
      RECT 56.555 2.4 56.815 2.72 ;
      RECT 55.875 4.78 56.135 5.1 ;
      RECT 55.935 2.74 56.075 5.1 ;
      RECT 55.875 2.74 56.135 3.06 ;
      RECT 47.3 6.28 47.62 6.605 ;
      RECT 47.33 5.695 47.5 6.605 ;
      RECT 47.33 5.695 47.505 6.045 ;
      RECT 47.33 5.695 48.305 5.87 ;
      RECT 48.13 1.965 48.305 5.87 ;
      RECT 40.685 2.205 40.965 2.575 ;
      RECT 40.685 2.345 45.335 2.52 ;
      RECT 45.16 2.025 45.335 2.52 ;
      RECT 45.63 1.995 45.955 2.32 ;
      RECT 48.075 1.965 48.425 2.315 ;
      RECT 45.16 2.025 48.425 2.195 ;
      RECT 36.45 8.29 47.145 8.46 ;
      RECT 46.985 2.395 47.145 8.46 ;
      RECT 36.45 6.545 36.62 8.46 ;
      RECT 48.1 6.655 48.425 6.98 ;
      RECT 33.27 6.655 33.595 6.98 ;
      RECT 46.985 6.745 48.425 6.915 ;
      RECT 36.4 6.545 36.68 6.885 ;
      RECT 33.27 6.685 36.69 6.855 ;
      RECT 47.3 2.365 47.62 2.685 ;
      RECT 46.985 2.395 47.62 2.565 ;
      RECT 43.755 6.48 44.015 6.8 ;
      RECT 43.815 2.74 43.955 6.8 ;
      RECT 43.755 2.74 44.015 3.06 ;
      RECT 43.075 4.78 43.335 5.1 ;
      RECT 43.135 3.76 43.275 5.1 ;
      RECT 43.075 3.76 43.335 4.08 ;
      RECT 42.055 6.48 42.315 6.8 ;
      RECT 42.115 5.21 42.255 6.8 ;
      RECT 41.435 5.21 42.255 5.35 ;
      RECT 41.435 2.74 41.575 5.35 ;
      RECT 41.365 4.135 41.645 4.505 ;
      RECT 41.375 2.74 41.635 3.06 ;
      RECT 39.325 4.135 39.605 4.505 ;
      RECT 39.395 2.4 39.535 4.505 ;
      RECT 39.335 2.4 39.595 2.72 ;
      RECT 38.655 4.78 38.915 5.1 ;
      RECT 38.715 2.74 38.855 5.1 ;
      RECT 38.655 2.74 38.915 3.06 ;
      RECT 30.08 6.28 30.4 6.605 ;
      RECT 30.11 5.695 30.28 6.605 ;
      RECT 30.11 5.695 30.285 6.045 ;
      RECT 30.11 5.695 31.085 5.87 ;
      RECT 30.91 1.965 31.085 5.87 ;
      RECT 23.465 2.205 23.745 2.575 ;
      RECT 23.465 2.345 28.115 2.52 ;
      RECT 27.94 2.025 28.115 2.52 ;
      RECT 28.41 1.995 28.735 2.32 ;
      RECT 30.855 1.965 31.205 2.315 ;
      RECT 27.94 2.025 31.205 2.195 ;
      RECT 19.23 8.29 29.925 8.46 ;
      RECT 29.765 2.395 29.925 8.46 ;
      RECT 19.23 6.545 19.4 8.46 ;
      RECT 30.88 6.655 31.205 6.98 ;
      RECT 16.05 6.655 16.375 6.98 ;
      RECT 29.765 6.745 31.205 6.915 ;
      RECT 19.18 6.545 19.46 6.885 ;
      RECT 16.05 6.685 19.46 6.855 ;
      RECT 30.08 2.365 30.4 2.685 ;
      RECT 29.765 2.395 30.4 2.565 ;
      RECT 26.535 6.48 26.795 6.8 ;
      RECT 26.595 2.74 26.735 6.8 ;
      RECT 26.535 2.74 26.795 3.06 ;
      RECT 25.855 4.78 26.115 5.1 ;
      RECT 25.915 3.76 26.055 5.1 ;
      RECT 25.855 3.76 26.115 4.08 ;
      RECT 24.835 6.48 25.095 6.8 ;
      RECT 24.895 5.21 25.035 6.8 ;
      RECT 24.215 5.21 25.035 5.35 ;
      RECT 24.215 2.74 24.355 5.35 ;
      RECT 24.145 4.135 24.425 4.505 ;
      RECT 24.155 2.74 24.415 3.06 ;
      RECT 22.105 4.135 22.385 4.505 ;
      RECT 22.175 2.4 22.315 4.505 ;
      RECT 22.115 2.4 22.375 2.72 ;
      RECT 21.435 4.78 21.695 5.1 ;
      RECT 21.495 2.74 21.635 5.1 ;
      RECT 21.435 2.74 21.695 3.06 ;
      RECT 12.86 6.28 13.18 6.605 ;
      RECT 12.89 5.695 13.06 6.605 ;
      RECT 12.89 5.695 13.065 6.045 ;
      RECT 12.89 5.695 13.865 5.87 ;
      RECT 13.69 1.965 13.865 5.87 ;
      RECT 6.245 2.205 6.525 2.575 ;
      RECT 6.245 2.345 10.895 2.52 ;
      RECT 10.72 2.025 10.895 2.52 ;
      RECT 11.19 1.995 11.515 2.32 ;
      RECT 13.635 1.965 13.985 2.315 ;
      RECT 10.72 2.025 13.985 2.195 ;
      RECT 2.01 8.29 12.705 8.46 ;
      RECT 12.545 2.395 12.705 8.46 ;
      RECT 2.01 6.545 2.18 8.46 ;
      RECT -1.89 6.995 -1.61 7.335 ;
      RECT -1.89 7.06 -0.685 7.23 ;
      RECT -0.855 6.685 -0.685 7.23 ;
      RECT 13.66 6.655 13.985 6.98 ;
      RECT 12.545 6.745 13.985 6.915 ;
      RECT 1.96 6.545 2.24 6.885 ;
      RECT -0.855 6.685 2.24 6.855 ;
      RECT 12.86 2.365 13.18 2.685 ;
      RECT 12.545 2.395 13.18 2.565 ;
      RECT 9.315 6.48 9.575 6.8 ;
      RECT 9.375 2.74 9.515 6.8 ;
      RECT 9.315 2.74 9.575 3.06 ;
      RECT 8.635 4.78 8.895 5.1 ;
      RECT 8.695 3.76 8.835 5.1 ;
      RECT 8.635 3.76 8.895 4.08 ;
      RECT 7.615 6.48 7.875 6.8 ;
      RECT 7.675 5.21 7.815 6.8 ;
      RECT 6.995 5.21 7.815 5.35 ;
      RECT 6.995 2.74 7.135 5.35 ;
      RECT 6.925 4.135 7.205 4.505 ;
      RECT 6.935 2.74 7.195 3.06 ;
      RECT 4.885 4.135 5.165 4.505 ;
      RECT 4.955 2.4 5.095 4.505 ;
      RECT 4.895 2.4 5.155 2.72 ;
      RECT 4.215 4.78 4.475 5.1 ;
      RECT 4.275 2.74 4.415 5.1 ;
      RECT 4.215 2.74 4.475 3.06 ;
      RECT 77.175 5.77 77.455 6.14 ;
      RECT 76.825 3.735 77.105 4.105 ;
      RECT 76.485 3.055 76.765 3.425 ;
      RECT 76.135 5.77 76.415 6.14 ;
      RECT 75.455 3.395 75.735 3.765 ;
      RECT 75.125 6.46 75.405 6.83 ;
      RECT 70.365 7 70.735 7.37 ;
      RECT 59.955 5.77 60.235 6.14 ;
      RECT 59.605 3.735 59.885 4.105 ;
      RECT 59.265 3.055 59.545 3.425 ;
      RECT 58.915 5.77 59.195 6.14 ;
      RECT 58.235 3.395 58.515 3.765 ;
      RECT 57.905 6.46 58.185 6.83 ;
      RECT 53.145 7 53.515 7.37 ;
      RECT 42.735 5.77 43.015 6.14 ;
      RECT 42.385 3.735 42.665 4.105 ;
      RECT 42.045 3.055 42.325 3.425 ;
      RECT 41.695 5.77 41.975 6.14 ;
      RECT 41.015 3.395 41.295 3.765 ;
      RECT 40.685 6.46 40.965 6.83 ;
      RECT 35.925 7 36.295 7.37 ;
      RECT 25.515 5.77 25.795 6.14 ;
      RECT 25.165 3.735 25.445 4.105 ;
      RECT 24.825 3.055 25.105 3.425 ;
      RECT 24.475 5.77 24.755 6.14 ;
      RECT 23.795 3.395 24.075 3.765 ;
      RECT 23.465 6.46 23.745 6.83 ;
      RECT 18.705 7 19.075 7.37 ;
      RECT 8.295 5.77 8.575 6.14 ;
      RECT 7.945 3.735 8.225 4.105 ;
      RECT 7.605 3.055 7.885 3.425 ;
      RECT 7.255 5.77 7.535 6.14 ;
      RECT 6.575 3.395 6.855 3.765 ;
      RECT 6.245 6.46 6.525 6.83 ;
      RECT 1.485 7 1.855 7.37 ;
    LAYER via1 ;
      RECT 84.985 7.385 85.135 7.535 ;
      RECT 82.63 6.74 82.78 6.89 ;
      RECT 82.615 2.065 82.765 2.215 ;
      RECT 81.825 2.45 81.975 2.6 ;
      RECT 81.825 6.37 81.975 6.52 ;
      RECT 80.16 2.08 80.31 2.23 ;
      RECT 78.25 2.825 78.4 2.975 ;
      RECT 78.25 6.565 78.4 6.715 ;
      RECT 77.57 3.845 77.72 3.995 ;
      RECT 77.57 4.865 77.72 5.015 ;
      RECT 77.23 5.885 77.38 6.035 ;
      RECT 76.89 3.845 77.04 3.995 ;
      RECT 76.55 3.165 76.7 3.315 ;
      RECT 76.55 6.565 76.7 6.715 ;
      RECT 76.2 5.885 76.35 6.035 ;
      RECT 75.87 2.825 76.02 2.975 ;
      RECT 75.53 3.505 75.68 3.655 ;
      RECT 75.19 2.315 75.34 2.465 ;
      RECT 75.19 6.565 75.34 6.715 ;
      RECT 73.83 2.485 73.98 2.635 ;
      RECT 73.15 2.825 73.3 2.975 ;
      RECT 73.15 4.865 73.3 5.015 ;
      RECT 70.905 6.64 71.055 6.79 ;
      RECT 70.475 7.11 70.625 7.26 ;
      RECT 67.8 6.74 67.95 6.89 ;
      RECT 65.41 6.74 65.56 6.89 ;
      RECT 65.395 2.065 65.545 2.215 ;
      RECT 64.605 2.45 64.755 2.6 ;
      RECT 64.605 6.37 64.755 6.52 ;
      RECT 62.94 2.08 63.09 2.23 ;
      RECT 61.03 2.825 61.18 2.975 ;
      RECT 61.03 6.565 61.18 6.715 ;
      RECT 60.35 3.845 60.5 3.995 ;
      RECT 60.35 4.865 60.5 5.015 ;
      RECT 60.01 5.885 60.16 6.035 ;
      RECT 59.67 3.845 59.82 3.995 ;
      RECT 59.33 3.165 59.48 3.315 ;
      RECT 59.33 6.565 59.48 6.715 ;
      RECT 58.98 5.885 59.13 6.035 ;
      RECT 58.65 2.825 58.8 2.975 ;
      RECT 58.31 3.505 58.46 3.655 ;
      RECT 57.97 2.315 58.12 2.465 ;
      RECT 57.97 6.565 58.12 6.715 ;
      RECT 56.61 2.485 56.76 2.635 ;
      RECT 55.93 2.825 56.08 2.975 ;
      RECT 55.93 4.865 56.08 5.015 ;
      RECT 53.685 6.64 53.835 6.79 ;
      RECT 53.255 7.11 53.405 7.26 ;
      RECT 50.58 6.74 50.73 6.89 ;
      RECT 48.19 6.74 48.34 6.89 ;
      RECT 48.175 2.065 48.325 2.215 ;
      RECT 47.385 2.45 47.535 2.6 ;
      RECT 47.385 6.37 47.535 6.52 ;
      RECT 45.72 2.08 45.87 2.23 ;
      RECT 43.81 2.825 43.96 2.975 ;
      RECT 43.81 6.565 43.96 6.715 ;
      RECT 43.13 3.845 43.28 3.995 ;
      RECT 43.13 4.865 43.28 5.015 ;
      RECT 42.79 5.885 42.94 6.035 ;
      RECT 42.45 3.845 42.6 3.995 ;
      RECT 42.11 3.165 42.26 3.315 ;
      RECT 42.11 6.565 42.26 6.715 ;
      RECT 41.76 5.885 41.91 6.035 ;
      RECT 41.43 2.825 41.58 2.975 ;
      RECT 41.09 3.505 41.24 3.655 ;
      RECT 40.75 2.315 40.9 2.465 ;
      RECT 40.75 6.565 40.9 6.715 ;
      RECT 39.39 2.485 39.54 2.635 ;
      RECT 38.71 2.825 38.86 2.975 ;
      RECT 38.71 4.865 38.86 5.015 ;
      RECT 36.465 6.64 36.615 6.79 ;
      RECT 36.035 7.11 36.185 7.26 ;
      RECT 33.36 6.74 33.51 6.89 ;
      RECT 30.97 6.74 31.12 6.89 ;
      RECT 30.955 2.065 31.105 2.215 ;
      RECT 30.165 2.45 30.315 2.6 ;
      RECT 30.165 6.37 30.315 6.52 ;
      RECT 28.5 2.08 28.65 2.23 ;
      RECT 26.59 2.825 26.74 2.975 ;
      RECT 26.59 6.565 26.74 6.715 ;
      RECT 25.91 3.845 26.06 3.995 ;
      RECT 25.91 4.865 26.06 5.015 ;
      RECT 25.57 5.885 25.72 6.035 ;
      RECT 25.23 3.845 25.38 3.995 ;
      RECT 24.89 3.165 25.04 3.315 ;
      RECT 24.89 6.565 25.04 6.715 ;
      RECT 24.54 5.885 24.69 6.035 ;
      RECT 24.21 2.825 24.36 2.975 ;
      RECT 23.87 3.505 24.02 3.655 ;
      RECT 23.53 2.315 23.68 2.465 ;
      RECT 23.53 6.565 23.68 6.715 ;
      RECT 22.17 2.485 22.32 2.635 ;
      RECT 21.49 2.825 21.64 2.975 ;
      RECT 21.49 4.865 21.64 5.015 ;
      RECT 19.245 6.64 19.395 6.79 ;
      RECT 18.815 7.11 18.965 7.26 ;
      RECT 16.14 6.74 16.29 6.89 ;
      RECT 13.75 6.74 13.9 6.89 ;
      RECT 13.735 2.065 13.885 2.215 ;
      RECT 12.945 2.45 13.095 2.6 ;
      RECT 12.945 6.37 13.095 6.52 ;
      RECT 11.28 2.08 11.43 2.23 ;
      RECT 9.37 2.825 9.52 2.975 ;
      RECT 9.37 6.565 9.52 6.715 ;
      RECT 8.69 3.845 8.84 3.995 ;
      RECT 8.69 4.865 8.84 5.015 ;
      RECT 8.35 5.885 8.5 6.035 ;
      RECT 8.01 3.845 8.16 3.995 ;
      RECT 7.67 3.165 7.82 3.315 ;
      RECT 7.67 6.565 7.82 6.715 ;
      RECT 7.32 5.885 7.47 6.035 ;
      RECT 6.99 2.825 7.14 2.975 ;
      RECT 6.65 3.505 6.8 3.655 ;
      RECT 6.31 2.315 6.46 2.465 ;
      RECT 6.31 6.565 6.46 6.715 ;
      RECT 4.95 2.485 5.1 2.635 ;
      RECT 4.27 2.825 4.42 2.975 ;
      RECT 4.27 4.865 4.42 5.015 ;
      RECT 2.025 6.64 2.175 6.79 ;
      RECT 1.595 7.11 1.745 7.26 ;
      RECT -1.825 7.09 -1.675 7.24 ;
      RECT -2.2 6.35 -2.05 6.5 ;
    LAYER met1 ;
      RECT 84.865 7.77 85.155 8 ;
      RECT 84.925 6.29 85.095 8 ;
      RECT 84.895 7.3 85.22 7.625 ;
      RECT 84.865 6.29 85.155 6.52 ;
      RECT 84.46 2.395 84.565 2.965 ;
      RECT 84.46 2.73 84.785 2.96 ;
      RECT 84.46 2.76 84.955 2.93 ;
      RECT 84.46 2.395 84.65 2.96 ;
      RECT 83.875 2.36 84.165 2.59 ;
      RECT 83.875 2.395 84.65 2.565 ;
      RECT 83.935 0.88 84.105 2.59 ;
      RECT 83.875 0.88 84.165 1.11 ;
      RECT 83.875 7.77 84.165 8 ;
      RECT 83.935 6.29 84.105 8 ;
      RECT 83.875 6.29 84.165 6.52 ;
      RECT 83.875 6.325 84.73 6.485 ;
      RECT 84.56 5.92 84.73 6.485 ;
      RECT 83.875 6.32 84.27 6.485 ;
      RECT 84.495 5.92 84.785 6.15 ;
      RECT 84.495 5.95 84.955 6.12 ;
      RECT 83.505 2.73 83.795 2.96 ;
      RECT 83.505 2.76 83.965 2.93 ;
      RECT 83.57 1.655 83.735 2.96 ;
      RECT 82.085 1.625 82.375 1.855 ;
      RECT 82.085 1.655 83.735 1.825 ;
      RECT 82.145 0.885 82.315 1.855 ;
      RECT 82.085 0.885 82.375 1.115 ;
      RECT 82.085 7.765 82.375 7.995 ;
      RECT 82.145 7.025 82.315 7.995 ;
      RECT 82.145 7.12 83.735 7.29 ;
      RECT 83.565 5.92 83.735 7.29 ;
      RECT 82.085 7.025 82.375 7.255 ;
      RECT 83.505 5.92 83.795 6.15 ;
      RECT 83.505 5.95 83.965 6.12 ;
      RECT 82.515 1.965 82.865 2.315 ;
      RECT 82.345 2.025 82.865 2.195 ;
      RECT 82.54 6.655 82.865 6.98 ;
      RECT 82.515 6.655 82.865 6.885 ;
      RECT 82.345 6.685 82.865 6.855 ;
      RECT 81.74 2.365 82.06 2.685 ;
      RECT 81.71 2.365 82.06 2.595 ;
      RECT 81.425 2.395 82.06 2.565 ;
      RECT 81.74 6.28 82.06 6.605 ;
      RECT 81.71 6.285 82.06 6.515 ;
      RECT 81.54 6.315 82.06 6.485 ;
      RECT 77.485 3.79 77.805 4.05 ;
      RECT 78.52 3.805 78.81 4.035 ;
      RECT 77.485 3.85 78.81 3.99 ;
      RECT 77.145 5.83 77.465 6.09 ;
      RECT 78.52 5.845 78.81 6.075 ;
      RECT 78.595 5.55 78.735 6.075 ;
      RECT 77.235 5.55 77.375 6.09 ;
      RECT 77.235 5.55 78.735 5.69 ;
      RECT 78.165 2.77 78.485 3.03 ;
      RECT 77.89 2.83 78.485 2.97 ;
      RECT 75.105 6.51 75.425 6.77 ;
      RECT 74.1 6.525 74.39 6.755 ;
      RECT 74.1 6.57 76.015 6.71 ;
      RECT 75.875 6.23 76.015 6.71 ;
      RECT 75.875 6.23 77.885 6.37 ;
      RECT 77.745 5.845 77.885 6.37 ;
      RECT 77.67 5.845 77.96 6.075 ;
      RECT 77.485 4.81 77.805 5.07 ;
      RECT 75.34 4.825 75.63 5.055 ;
      RECT 75.34 4.87 77.805 5.01 ;
      RECT 76.805 3.79 77.125 4.05 ;
      RECT 74.44 3.805 74.73 4.035 ;
      RECT 74.44 3.85 77.125 3.99 ;
      RECT 76.465 6.51 76.785 6.77 ;
      RECT 76.465 6.57 77.06 6.71 ;
      RECT 76.465 3.11 76.785 3.37 ;
      RECT 76.19 3.17 76.785 3.31 ;
      RECT 75.785 2.77 76.105 3.03 ;
      RECT 75.51 2.83 76.105 2.97 ;
      RECT 75.445 3.45 75.765 3.71 ;
      RECT 72.57 3.465 72.86 3.695 ;
      RECT 72.57 3.51 75.765 3.65 ;
      RECT 75.025 2.79 75.165 3.65 ;
      RECT 74.95 2.79 75.24 3.02 ;
      RECT 75.105 2.26 75.425 2.52 ;
      RECT 75.105 2.275 75.61 2.505 ;
      RECT 75.015 2.32 75.61 2.46 ;
      RECT 74.44 2.79 74.73 3.02 ;
      RECT 73.835 2.835 74.73 2.975 ;
      RECT 73.835 2.43 73.975 2.975 ;
      RECT 73.745 2.43 74.065 2.69 ;
      RECT 73.065 2.77 73.385 3.03 ;
      RECT 72.79 2.83 73.385 2.97 ;
      RECT 73.065 4.81 73.385 5.07 ;
      RECT 72.79 4.87 73.385 5.01 ;
      RECT 70.83 6.575 71.12 6.885 ;
      RECT 70.66 6.685 71.15 6.855 ;
      RECT 70.81 6.575 71.15 6.855 ;
      RECT 70.4 7.765 70.69 7.995 ;
      RECT 70.46 6.995 70.63 7.995 ;
      RECT 70.365 6.995 70.735 7.37 ;
      RECT 67.645 7.77 67.935 8 ;
      RECT 67.705 6.29 67.875 8 ;
      RECT 67.705 6.655 68.035 6.98 ;
      RECT 67.645 6.29 67.935 6.52 ;
      RECT 67.24 2.395 67.345 2.965 ;
      RECT 67.24 2.73 67.565 2.96 ;
      RECT 67.24 2.76 67.735 2.93 ;
      RECT 67.24 2.395 67.43 2.96 ;
      RECT 66.655 2.36 66.945 2.59 ;
      RECT 66.655 2.395 67.43 2.565 ;
      RECT 66.715 0.88 66.885 2.59 ;
      RECT 66.655 0.88 66.945 1.11 ;
      RECT 66.655 7.77 66.945 8 ;
      RECT 66.715 6.29 66.885 8 ;
      RECT 66.655 6.29 66.945 6.52 ;
      RECT 66.655 6.325 67.51 6.485 ;
      RECT 67.34 5.92 67.51 6.485 ;
      RECT 66.655 6.32 67.05 6.485 ;
      RECT 67.275 5.92 67.565 6.15 ;
      RECT 67.275 5.95 67.735 6.12 ;
      RECT 66.285 2.73 66.575 2.96 ;
      RECT 66.285 2.76 66.745 2.93 ;
      RECT 66.35 1.655 66.515 2.96 ;
      RECT 64.865 1.625 65.155 1.855 ;
      RECT 64.865 1.655 66.515 1.825 ;
      RECT 64.925 0.885 65.095 1.855 ;
      RECT 64.865 0.885 65.155 1.115 ;
      RECT 64.865 7.765 65.155 7.995 ;
      RECT 64.925 7.025 65.095 7.995 ;
      RECT 64.925 7.12 66.515 7.29 ;
      RECT 66.345 5.92 66.515 7.29 ;
      RECT 64.865 7.025 65.155 7.255 ;
      RECT 66.285 5.92 66.575 6.15 ;
      RECT 66.285 5.95 66.745 6.12 ;
      RECT 65.295 1.965 65.645 2.315 ;
      RECT 65.125 2.025 65.645 2.195 ;
      RECT 65.32 6.655 65.645 6.98 ;
      RECT 65.295 6.655 65.645 6.885 ;
      RECT 65.125 6.685 65.645 6.855 ;
      RECT 64.52 2.365 64.84 2.685 ;
      RECT 64.49 2.365 64.84 2.595 ;
      RECT 64.205 2.395 64.84 2.565 ;
      RECT 64.52 6.28 64.84 6.605 ;
      RECT 64.49 6.285 64.84 6.515 ;
      RECT 64.32 6.315 64.84 6.485 ;
      RECT 60.265 3.79 60.585 4.05 ;
      RECT 61.3 3.805 61.59 4.035 ;
      RECT 60.265 3.85 61.59 3.99 ;
      RECT 59.925 5.83 60.245 6.09 ;
      RECT 61.3 5.845 61.59 6.075 ;
      RECT 61.375 5.55 61.515 6.075 ;
      RECT 60.015 5.55 60.155 6.09 ;
      RECT 60.015 5.55 61.515 5.69 ;
      RECT 60.945 2.77 61.265 3.03 ;
      RECT 60.67 2.83 61.265 2.97 ;
      RECT 57.885 6.51 58.205 6.77 ;
      RECT 56.88 6.525 57.17 6.755 ;
      RECT 56.88 6.57 58.795 6.71 ;
      RECT 58.655 6.23 58.795 6.71 ;
      RECT 58.655 6.23 60.665 6.37 ;
      RECT 60.525 5.845 60.665 6.37 ;
      RECT 60.45 5.845 60.74 6.075 ;
      RECT 60.265 4.81 60.585 5.07 ;
      RECT 58.12 4.825 58.41 5.055 ;
      RECT 58.12 4.87 60.585 5.01 ;
      RECT 59.585 3.79 59.905 4.05 ;
      RECT 57.22 3.805 57.51 4.035 ;
      RECT 57.22 3.85 59.905 3.99 ;
      RECT 59.245 6.51 59.565 6.77 ;
      RECT 59.245 6.57 59.84 6.71 ;
      RECT 59.245 3.11 59.565 3.37 ;
      RECT 58.97 3.17 59.565 3.31 ;
      RECT 58.565 2.77 58.885 3.03 ;
      RECT 58.29 2.83 58.885 2.97 ;
      RECT 58.225 3.45 58.545 3.71 ;
      RECT 55.35 3.465 55.64 3.695 ;
      RECT 55.35 3.51 58.545 3.65 ;
      RECT 57.805 2.79 57.945 3.65 ;
      RECT 57.73 2.79 58.02 3.02 ;
      RECT 57.885 2.26 58.205 2.52 ;
      RECT 57.885 2.275 58.39 2.505 ;
      RECT 57.795 2.32 58.39 2.46 ;
      RECT 57.22 2.79 57.51 3.02 ;
      RECT 56.615 2.835 57.51 2.975 ;
      RECT 56.615 2.43 56.755 2.975 ;
      RECT 56.525 2.43 56.845 2.69 ;
      RECT 55.845 2.77 56.165 3.03 ;
      RECT 55.57 2.83 56.165 2.97 ;
      RECT 55.845 4.81 56.165 5.07 ;
      RECT 55.57 4.87 56.165 5.01 ;
      RECT 53.61 6.575 53.9 6.885 ;
      RECT 53.44 6.685 53.93 6.855 ;
      RECT 53.59 6.575 53.93 6.855 ;
      RECT 53.18 7.765 53.47 7.995 ;
      RECT 53.24 6.995 53.41 7.995 ;
      RECT 53.145 6.995 53.515 7.37 ;
      RECT 50.425 7.77 50.715 8 ;
      RECT 50.485 6.29 50.655 8 ;
      RECT 50.485 6.655 50.815 6.98 ;
      RECT 50.425 6.29 50.715 6.52 ;
      RECT 50.02 2.395 50.125 2.965 ;
      RECT 50.02 2.73 50.345 2.96 ;
      RECT 50.02 2.76 50.515 2.93 ;
      RECT 50.02 2.395 50.21 2.96 ;
      RECT 49.435 2.36 49.725 2.59 ;
      RECT 49.435 2.395 50.21 2.565 ;
      RECT 49.495 0.88 49.665 2.59 ;
      RECT 49.435 0.88 49.725 1.11 ;
      RECT 49.435 7.77 49.725 8 ;
      RECT 49.495 6.29 49.665 8 ;
      RECT 49.435 6.29 49.725 6.52 ;
      RECT 49.435 6.325 50.29 6.485 ;
      RECT 50.12 5.92 50.29 6.485 ;
      RECT 49.435 6.32 49.83 6.485 ;
      RECT 50.055 5.92 50.345 6.15 ;
      RECT 50.055 5.95 50.515 6.12 ;
      RECT 49.065 2.73 49.355 2.96 ;
      RECT 49.065 2.76 49.525 2.93 ;
      RECT 49.13 1.655 49.295 2.96 ;
      RECT 47.645 1.625 47.935 1.855 ;
      RECT 47.645 1.655 49.295 1.825 ;
      RECT 47.705 0.885 47.875 1.855 ;
      RECT 47.645 0.885 47.935 1.115 ;
      RECT 47.645 7.765 47.935 7.995 ;
      RECT 47.705 7.025 47.875 7.995 ;
      RECT 47.705 7.12 49.295 7.29 ;
      RECT 49.125 5.92 49.295 7.29 ;
      RECT 47.645 7.025 47.935 7.255 ;
      RECT 49.065 5.92 49.355 6.15 ;
      RECT 49.065 5.95 49.525 6.12 ;
      RECT 48.075 1.965 48.425 2.315 ;
      RECT 47.905 2.025 48.425 2.195 ;
      RECT 48.1 6.655 48.425 6.98 ;
      RECT 48.075 6.655 48.425 6.885 ;
      RECT 47.905 6.685 48.425 6.855 ;
      RECT 47.3 2.365 47.62 2.685 ;
      RECT 47.27 2.365 47.62 2.595 ;
      RECT 46.985 2.395 47.62 2.565 ;
      RECT 47.3 6.28 47.62 6.605 ;
      RECT 47.27 6.285 47.62 6.515 ;
      RECT 47.1 6.315 47.62 6.485 ;
      RECT 43.045 3.79 43.365 4.05 ;
      RECT 44.08 3.805 44.37 4.035 ;
      RECT 43.045 3.85 44.37 3.99 ;
      RECT 42.705 5.83 43.025 6.09 ;
      RECT 44.08 5.845 44.37 6.075 ;
      RECT 44.155 5.55 44.295 6.075 ;
      RECT 42.795 5.55 42.935 6.09 ;
      RECT 42.795 5.55 44.295 5.69 ;
      RECT 43.725 2.77 44.045 3.03 ;
      RECT 43.45 2.83 44.045 2.97 ;
      RECT 40.665 6.51 40.985 6.77 ;
      RECT 39.66 6.525 39.95 6.755 ;
      RECT 39.66 6.57 41.575 6.71 ;
      RECT 41.435 6.23 41.575 6.71 ;
      RECT 41.435 6.23 43.445 6.37 ;
      RECT 43.305 5.845 43.445 6.37 ;
      RECT 43.23 5.845 43.52 6.075 ;
      RECT 43.045 4.81 43.365 5.07 ;
      RECT 40.9 4.825 41.19 5.055 ;
      RECT 40.9 4.87 43.365 5.01 ;
      RECT 42.365 3.79 42.685 4.05 ;
      RECT 40 3.805 40.29 4.035 ;
      RECT 40 3.85 42.685 3.99 ;
      RECT 42.025 6.51 42.345 6.77 ;
      RECT 42.025 6.57 42.62 6.71 ;
      RECT 42.025 3.11 42.345 3.37 ;
      RECT 41.75 3.17 42.345 3.31 ;
      RECT 41.345 2.77 41.665 3.03 ;
      RECT 41.07 2.83 41.665 2.97 ;
      RECT 41.005 3.45 41.325 3.71 ;
      RECT 38.13 3.465 38.42 3.695 ;
      RECT 38.13 3.51 41.325 3.65 ;
      RECT 40.585 2.79 40.725 3.65 ;
      RECT 40.51 2.79 40.8 3.02 ;
      RECT 40.665 2.26 40.985 2.52 ;
      RECT 40.665 2.275 41.17 2.505 ;
      RECT 40.575 2.32 41.17 2.46 ;
      RECT 40 2.79 40.29 3.02 ;
      RECT 39.395 2.835 40.29 2.975 ;
      RECT 39.395 2.43 39.535 2.975 ;
      RECT 39.305 2.43 39.625 2.69 ;
      RECT 38.625 2.77 38.945 3.03 ;
      RECT 38.35 2.83 38.945 2.97 ;
      RECT 38.625 4.81 38.945 5.07 ;
      RECT 38.35 4.87 38.945 5.01 ;
      RECT 36.39 6.575 36.68 6.885 ;
      RECT 36.22 6.685 36.71 6.855 ;
      RECT 36.37 6.575 36.71 6.855 ;
      RECT 35.96 7.765 36.25 7.995 ;
      RECT 36.02 6.995 36.19 7.995 ;
      RECT 35.925 6.995 36.295 7.37 ;
      RECT 33.205 7.77 33.495 8 ;
      RECT 33.265 6.29 33.435 8 ;
      RECT 33.265 6.655 33.595 6.98 ;
      RECT 33.205 6.29 33.495 6.52 ;
      RECT 32.8 2.395 32.905 2.965 ;
      RECT 32.8 2.73 33.125 2.96 ;
      RECT 32.8 2.76 33.295 2.93 ;
      RECT 32.8 2.395 32.99 2.96 ;
      RECT 32.215 2.36 32.505 2.59 ;
      RECT 32.215 2.395 32.99 2.565 ;
      RECT 32.275 0.88 32.445 2.59 ;
      RECT 32.215 0.88 32.505 1.11 ;
      RECT 32.215 7.77 32.505 8 ;
      RECT 32.275 6.29 32.445 8 ;
      RECT 32.215 6.29 32.505 6.52 ;
      RECT 32.215 6.325 33.07 6.485 ;
      RECT 32.9 5.92 33.07 6.485 ;
      RECT 32.215 6.32 32.61 6.485 ;
      RECT 32.835 5.92 33.125 6.15 ;
      RECT 32.835 5.95 33.295 6.12 ;
      RECT 31.845 2.73 32.135 2.96 ;
      RECT 31.845 2.76 32.305 2.93 ;
      RECT 31.91 1.655 32.075 2.96 ;
      RECT 30.425 1.625 30.715 1.855 ;
      RECT 30.425 1.655 32.075 1.825 ;
      RECT 30.485 0.885 30.655 1.855 ;
      RECT 30.425 0.885 30.715 1.115 ;
      RECT 30.425 7.765 30.715 7.995 ;
      RECT 30.485 7.025 30.655 7.995 ;
      RECT 30.485 7.12 32.075 7.29 ;
      RECT 31.905 5.92 32.075 7.29 ;
      RECT 30.425 7.025 30.715 7.255 ;
      RECT 31.845 5.92 32.135 6.15 ;
      RECT 31.845 5.95 32.305 6.12 ;
      RECT 30.855 1.965 31.205 2.315 ;
      RECT 30.685 2.025 31.205 2.195 ;
      RECT 30.88 6.655 31.205 6.98 ;
      RECT 30.855 6.655 31.205 6.885 ;
      RECT 30.685 6.685 31.205 6.855 ;
      RECT 30.08 2.365 30.4 2.685 ;
      RECT 30.05 2.365 30.4 2.595 ;
      RECT 29.765 2.395 30.4 2.565 ;
      RECT 30.08 6.28 30.4 6.605 ;
      RECT 30.05 6.285 30.4 6.515 ;
      RECT 29.88 6.315 30.4 6.485 ;
      RECT 25.825 3.79 26.145 4.05 ;
      RECT 26.86 3.805 27.15 4.035 ;
      RECT 25.825 3.85 27.15 3.99 ;
      RECT 25.485 5.83 25.805 6.09 ;
      RECT 26.86 5.845 27.15 6.075 ;
      RECT 26.935 5.55 27.075 6.075 ;
      RECT 25.575 5.55 25.715 6.09 ;
      RECT 25.575 5.55 27.075 5.69 ;
      RECT 26.505 2.77 26.825 3.03 ;
      RECT 26.23 2.83 26.825 2.97 ;
      RECT 23.445 6.51 23.765 6.77 ;
      RECT 22.44 6.525 22.73 6.755 ;
      RECT 22.44 6.57 24.355 6.71 ;
      RECT 24.215 6.23 24.355 6.71 ;
      RECT 24.215 6.23 26.225 6.37 ;
      RECT 26.085 5.845 26.225 6.37 ;
      RECT 26.01 5.845 26.3 6.075 ;
      RECT 25.825 4.81 26.145 5.07 ;
      RECT 23.68 4.825 23.97 5.055 ;
      RECT 23.68 4.87 26.145 5.01 ;
      RECT 25.145 3.79 25.465 4.05 ;
      RECT 22.78 3.805 23.07 4.035 ;
      RECT 22.78 3.85 25.465 3.99 ;
      RECT 24.805 6.51 25.125 6.77 ;
      RECT 24.805 6.57 25.4 6.71 ;
      RECT 24.805 3.11 25.125 3.37 ;
      RECT 24.53 3.17 25.125 3.31 ;
      RECT 24.125 2.77 24.445 3.03 ;
      RECT 23.85 2.83 24.445 2.97 ;
      RECT 23.785 3.45 24.105 3.71 ;
      RECT 20.91 3.465 21.2 3.695 ;
      RECT 20.91 3.51 24.105 3.65 ;
      RECT 23.365 2.79 23.505 3.65 ;
      RECT 23.29 2.79 23.58 3.02 ;
      RECT 23.445 2.26 23.765 2.52 ;
      RECT 23.445 2.275 23.95 2.505 ;
      RECT 23.355 2.32 23.95 2.46 ;
      RECT 22.78 2.79 23.07 3.02 ;
      RECT 22.175 2.835 23.07 2.975 ;
      RECT 22.175 2.43 22.315 2.975 ;
      RECT 22.085 2.43 22.405 2.69 ;
      RECT 21.405 2.77 21.725 3.03 ;
      RECT 21.13 2.83 21.725 2.97 ;
      RECT 21.405 4.81 21.725 5.07 ;
      RECT 21.13 4.87 21.725 5.01 ;
      RECT 19.17 6.575 19.46 6.885 ;
      RECT 19 6.685 19.49 6.855 ;
      RECT 19.15 6.575 19.49 6.855 ;
      RECT 18.74 7.765 19.03 7.995 ;
      RECT 18.8 6.995 18.97 7.995 ;
      RECT 18.705 6.995 19.075 7.37 ;
      RECT 15.985 7.77 16.275 8 ;
      RECT 16.045 6.29 16.215 8 ;
      RECT 16.045 6.655 16.375 6.98 ;
      RECT 15.985 6.29 16.275 6.52 ;
      RECT 15.58 2.395 15.685 2.965 ;
      RECT 15.58 2.73 15.905 2.96 ;
      RECT 15.58 2.76 16.075 2.93 ;
      RECT 15.58 2.395 15.77 2.96 ;
      RECT 14.995 2.36 15.285 2.59 ;
      RECT 14.995 2.395 15.77 2.565 ;
      RECT 15.055 0.88 15.225 2.59 ;
      RECT 14.995 0.88 15.285 1.11 ;
      RECT 14.995 7.77 15.285 8 ;
      RECT 15.055 6.29 15.225 8 ;
      RECT 14.995 6.29 15.285 6.52 ;
      RECT 14.995 6.325 15.85 6.485 ;
      RECT 15.68 5.92 15.85 6.485 ;
      RECT 14.995 6.32 15.39 6.485 ;
      RECT 15.615 5.92 15.905 6.15 ;
      RECT 15.615 5.95 16.075 6.12 ;
      RECT 14.625 2.73 14.915 2.96 ;
      RECT 14.625 2.76 15.085 2.93 ;
      RECT 14.69 1.655 14.855 2.96 ;
      RECT 13.205 1.625 13.495 1.855 ;
      RECT 13.205 1.655 14.855 1.825 ;
      RECT 13.265 0.885 13.435 1.855 ;
      RECT 13.205 0.885 13.495 1.115 ;
      RECT 13.205 7.765 13.495 7.995 ;
      RECT 13.265 7.025 13.435 7.995 ;
      RECT 13.265 7.12 14.855 7.29 ;
      RECT 14.685 5.92 14.855 7.29 ;
      RECT 13.205 7.025 13.495 7.255 ;
      RECT 14.625 5.92 14.915 6.15 ;
      RECT 14.625 5.95 15.085 6.12 ;
      RECT 13.635 1.965 13.985 2.315 ;
      RECT 13.465 2.025 13.985 2.195 ;
      RECT 13.66 6.655 13.985 6.98 ;
      RECT 13.635 6.655 13.985 6.885 ;
      RECT 13.465 6.685 13.985 6.855 ;
      RECT 12.86 2.365 13.18 2.685 ;
      RECT 12.83 2.365 13.18 2.595 ;
      RECT 12.545 2.395 13.18 2.565 ;
      RECT 12.86 6.28 13.18 6.605 ;
      RECT 12.83 6.285 13.18 6.515 ;
      RECT 12.66 6.315 13.18 6.485 ;
      RECT 8.605 3.79 8.925 4.05 ;
      RECT 9.64 3.805 9.93 4.035 ;
      RECT 8.605 3.85 9.93 3.99 ;
      RECT 8.265 5.83 8.585 6.09 ;
      RECT 9.64 5.845 9.93 6.075 ;
      RECT 9.715 5.55 9.855 6.075 ;
      RECT 8.355 5.55 8.495 6.09 ;
      RECT 8.355 5.55 9.855 5.69 ;
      RECT 9.285 2.77 9.605 3.03 ;
      RECT 9.01 2.83 9.605 2.97 ;
      RECT 6.225 6.51 6.545 6.77 ;
      RECT 5.22 6.525 5.51 6.755 ;
      RECT 5.22 6.57 7.135 6.71 ;
      RECT 6.995 6.23 7.135 6.71 ;
      RECT 6.995 6.23 9.005 6.37 ;
      RECT 8.865 5.845 9.005 6.37 ;
      RECT 8.79 5.845 9.08 6.075 ;
      RECT 8.605 4.81 8.925 5.07 ;
      RECT 6.46 4.825 6.75 5.055 ;
      RECT 6.46 4.87 8.925 5.01 ;
      RECT 7.925 3.79 8.245 4.05 ;
      RECT 5.56 3.805 5.85 4.035 ;
      RECT 5.56 3.85 8.245 3.99 ;
      RECT 7.585 6.51 7.905 6.77 ;
      RECT 7.585 6.57 8.18 6.71 ;
      RECT 7.585 3.11 7.905 3.37 ;
      RECT 7.31 3.17 7.905 3.31 ;
      RECT 6.905 2.77 7.225 3.03 ;
      RECT 6.63 2.83 7.225 2.97 ;
      RECT 6.565 3.45 6.885 3.71 ;
      RECT 3.69 3.465 3.98 3.695 ;
      RECT 3.69 3.51 6.885 3.65 ;
      RECT 6.145 2.79 6.285 3.65 ;
      RECT 6.07 2.79 6.36 3.02 ;
      RECT 6.225 2.26 6.545 2.52 ;
      RECT 6.225 2.275 6.73 2.505 ;
      RECT 6.135 2.32 6.73 2.46 ;
      RECT 5.56 2.79 5.85 3.02 ;
      RECT 4.955 2.835 5.85 2.975 ;
      RECT 4.955 2.43 5.095 2.975 ;
      RECT 4.865 2.43 5.185 2.69 ;
      RECT 4.185 2.77 4.505 3.03 ;
      RECT 3.91 2.83 4.505 2.97 ;
      RECT 4.185 4.81 4.505 5.07 ;
      RECT 3.91 4.87 4.505 5.01 ;
      RECT 1.95 6.575 2.24 6.885 ;
      RECT 1.78 6.685 2.27 6.855 ;
      RECT 1.93 6.575 2.27 6.855 ;
      RECT 1.52 7.765 1.81 7.995 ;
      RECT 1.58 6.995 1.75 7.995 ;
      RECT 1.485 6.995 1.855 7.37 ;
      RECT -1.89 7.765 -1.6 7.995 ;
      RECT -1.83 7.025 -1.66 7.995 ;
      RECT -1.92 7.025 -1.58 7.305 ;
      RECT -2.295 6.285 -1.955 6.565 ;
      RECT -2.435 6.315 -1.955 6.485 ;
      RECT 80.07 1.995 80.395 2.32 ;
      RECT 77.84 6.51 78.485 6.77 ;
      RECT 75.79 5.83 76.435 6.09 ;
      RECT 62.85 1.995 63.175 2.32 ;
      RECT 60.62 6.51 61.265 6.77 ;
      RECT 58.57 5.83 59.215 6.09 ;
      RECT 45.63 1.995 45.955 2.32 ;
      RECT 43.4 6.51 44.045 6.77 ;
      RECT 41.35 5.83 41.995 6.09 ;
      RECT 28.41 1.995 28.735 2.32 ;
      RECT 26.18 6.51 26.825 6.77 ;
      RECT 24.13 5.83 24.775 6.09 ;
      RECT 11.19 1.995 11.515 2.32 ;
      RECT 8.96 6.51 9.605 6.77 ;
      RECT 6.91 5.83 7.555 6.09 ;
    LAYER mcon ;
      RECT 84.925 6.32 85.095 6.49 ;
      RECT 84.93 6.315 85.1 6.485 ;
      RECT 67.705 6.32 67.875 6.49 ;
      RECT 67.71 6.315 67.88 6.485 ;
      RECT 50.485 6.32 50.655 6.49 ;
      RECT 50.49 6.315 50.66 6.485 ;
      RECT 33.265 6.32 33.435 6.49 ;
      RECT 33.27 6.315 33.44 6.485 ;
      RECT 16.045 6.32 16.215 6.49 ;
      RECT 16.05 6.315 16.22 6.485 ;
      RECT 84.925 7.8 85.095 7.97 ;
      RECT 84.555 2.76 84.725 2.93 ;
      RECT 84.555 5.95 84.725 6.12 ;
      RECT 83.935 0.91 84.105 1.08 ;
      RECT 83.935 2.39 84.105 2.56 ;
      RECT 83.935 6.32 84.105 6.49 ;
      RECT 83.935 7.8 84.105 7.97 ;
      RECT 83.565 2.76 83.735 2.93 ;
      RECT 83.565 5.95 83.735 6.12 ;
      RECT 82.575 2.025 82.745 2.195 ;
      RECT 82.575 6.685 82.745 6.855 ;
      RECT 82.145 0.915 82.315 1.085 ;
      RECT 82.145 1.655 82.315 1.825 ;
      RECT 82.145 7.055 82.315 7.225 ;
      RECT 82.145 7.795 82.315 7.965 ;
      RECT 81.77 2.395 81.94 2.565 ;
      RECT 81.77 6.315 81.94 6.485 ;
      RECT 78.58 3.835 78.75 4.005 ;
      RECT 78.58 5.875 78.75 6.045 ;
      RECT 78.24 2.815 78.41 2.985 ;
      RECT 77.9 6.555 78.07 6.725 ;
      RECT 77.73 5.875 77.9 6.045 ;
      RECT 77.22 5.875 77.39 6.045 ;
      RECT 76.54 3.155 76.71 3.325 ;
      RECT 76.54 6.555 76.71 6.725 ;
      RECT 75.86 2.815 76.03 2.985 ;
      RECT 75.85 5.875 76.02 6.045 ;
      RECT 75.4 4.855 75.57 5.025 ;
      RECT 75.38 2.305 75.55 2.475 ;
      RECT 75.01 2.82 75.18 2.99 ;
      RECT 74.5 2.82 74.67 2.99 ;
      RECT 74.5 3.835 74.67 4.005 ;
      RECT 74.16 6.555 74.33 6.725 ;
      RECT 73.14 2.815 73.31 2.985 ;
      RECT 73.14 4.855 73.31 5.025 ;
      RECT 72.63 3.495 72.8 3.665 ;
      RECT 70.89 6.685 71.06 6.855 ;
      RECT 70.46 7.055 70.63 7.225 ;
      RECT 70.46 7.795 70.63 7.965 ;
      RECT 67.705 7.8 67.875 7.97 ;
      RECT 67.335 2.76 67.505 2.93 ;
      RECT 67.335 5.95 67.505 6.12 ;
      RECT 66.715 0.91 66.885 1.08 ;
      RECT 66.715 2.39 66.885 2.56 ;
      RECT 66.715 6.32 66.885 6.49 ;
      RECT 66.715 7.8 66.885 7.97 ;
      RECT 66.345 2.76 66.515 2.93 ;
      RECT 66.345 5.95 66.515 6.12 ;
      RECT 65.355 2.025 65.525 2.195 ;
      RECT 65.355 6.685 65.525 6.855 ;
      RECT 64.925 0.915 65.095 1.085 ;
      RECT 64.925 1.655 65.095 1.825 ;
      RECT 64.925 7.055 65.095 7.225 ;
      RECT 64.925 7.795 65.095 7.965 ;
      RECT 64.55 2.395 64.72 2.565 ;
      RECT 64.55 6.315 64.72 6.485 ;
      RECT 61.36 3.835 61.53 4.005 ;
      RECT 61.36 5.875 61.53 6.045 ;
      RECT 61.02 2.815 61.19 2.985 ;
      RECT 60.68 6.555 60.85 6.725 ;
      RECT 60.51 5.875 60.68 6.045 ;
      RECT 60 5.875 60.17 6.045 ;
      RECT 59.32 3.155 59.49 3.325 ;
      RECT 59.32 6.555 59.49 6.725 ;
      RECT 58.64 2.815 58.81 2.985 ;
      RECT 58.63 5.875 58.8 6.045 ;
      RECT 58.18 4.855 58.35 5.025 ;
      RECT 58.16 2.305 58.33 2.475 ;
      RECT 57.79 2.82 57.96 2.99 ;
      RECT 57.28 2.82 57.45 2.99 ;
      RECT 57.28 3.835 57.45 4.005 ;
      RECT 56.94 6.555 57.11 6.725 ;
      RECT 55.92 2.815 56.09 2.985 ;
      RECT 55.92 4.855 56.09 5.025 ;
      RECT 55.41 3.495 55.58 3.665 ;
      RECT 53.67 6.685 53.84 6.855 ;
      RECT 53.24 7.055 53.41 7.225 ;
      RECT 53.24 7.795 53.41 7.965 ;
      RECT 50.485 7.8 50.655 7.97 ;
      RECT 50.115 2.76 50.285 2.93 ;
      RECT 50.115 5.95 50.285 6.12 ;
      RECT 49.495 0.91 49.665 1.08 ;
      RECT 49.495 2.39 49.665 2.56 ;
      RECT 49.495 6.32 49.665 6.49 ;
      RECT 49.495 7.8 49.665 7.97 ;
      RECT 49.125 2.76 49.295 2.93 ;
      RECT 49.125 5.95 49.295 6.12 ;
      RECT 48.135 2.025 48.305 2.195 ;
      RECT 48.135 6.685 48.305 6.855 ;
      RECT 47.705 0.915 47.875 1.085 ;
      RECT 47.705 1.655 47.875 1.825 ;
      RECT 47.705 7.055 47.875 7.225 ;
      RECT 47.705 7.795 47.875 7.965 ;
      RECT 47.33 2.395 47.5 2.565 ;
      RECT 47.33 6.315 47.5 6.485 ;
      RECT 44.14 3.835 44.31 4.005 ;
      RECT 44.14 5.875 44.31 6.045 ;
      RECT 43.8 2.815 43.97 2.985 ;
      RECT 43.46 6.555 43.63 6.725 ;
      RECT 43.29 5.875 43.46 6.045 ;
      RECT 42.78 5.875 42.95 6.045 ;
      RECT 42.1 3.155 42.27 3.325 ;
      RECT 42.1 6.555 42.27 6.725 ;
      RECT 41.42 2.815 41.59 2.985 ;
      RECT 41.41 5.875 41.58 6.045 ;
      RECT 40.96 4.855 41.13 5.025 ;
      RECT 40.94 2.305 41.11 2.475 ;
      RECT 40.57 2.82 40.74 2.99 ;
      RECT 40.06 2.82 40.23 2.99 ;
      RECT 40.06 3.835 40.23 4.005 ;
      RECT 39.72 6.555 39.89 6.725 ;
      RECT 38.7 2.815 38.87 2.985 ;
      RECT 38.7 4.855 38.87 5.025 ;
      RECT 38.19 3.495 38.36 3.665 ;
      RECT 36.45 6.685 36.62 6.855 ;
      RECT 36.02 7.055 36.19 7.225 ;
      RECT 36.02 7.795 36.19 7.965 ;
      RECT 33.265 7.8 33.435 7.97 ;
      RECT 32.895 2.76 33.065 2.93 ;
      RECT 32.895 5.95 33.065 6.12 ;
      RECT 32.275 0.91 32.445 1.08 ;
      RECT 32.275 2.39 32.445 2.56 ;
      RECT 32.275 6.32 32.445 6.49 ;
      RECT 32.275 7.8 32.445 7.97 ;
      RECT 31.905 2.76 32.075 2.93 ;
      RECT 31.905 5.95 32.075 6.12 ;
      RECT 30.915 2.025 31.085 2.195 ;
      RECT 30.915 6.685 31.085 6.855 ;
      RECT 30.485 0.915 30.655 1.085 ;
      RECT 30.485 1.655 30.655 1.825 ;
      RECT 30.485 7.055 30.655 7.225 ;
      RECT 30.485 7.795 30.655 7.965 ;
      RECT 30.11 2.395 30.28 2.565 ;
      RECT 30.11 6.315 30.28 6.485 ;
      RECT 26.92 3.835 27.09 4.005 ;
      RECT 26.92 5.875 27.09 6.045 ;
      RECT 26.58 2.815 26.75 2.985 ;
      RECT 26.24 6.555 26.41 6.725 ;
      RECT 26.07 5.875 26.24 6.045 ;
      RECT 25.56 5.875 25.73 6.045 ;
      RECT 24.88 3.155 25.05 3.325 ;
      RECT 24.88 6.555 25.05 6.725 ;
      RECT 24.2 2.815 24.37 2.985 ;
      RECT 24.19 5.875 24.36 6.045 ;
      RECT 23.74 4.855 23.91 5.025 ;
      RECT 23.72 2.305 23.89 2.475 ;
      RECT 23.35 2.82 23.52 2.99 ;
      RECT 22.84 2.82 23.01 2.99 ;
      RECT 22.84 3.835 23.01 4.005 ;
      RECT 22.5 6.555 22.67 6.725 ;
      RECT 21.48 2.815 21.65 2.985 ;
      RECT 21.48 4.855 21.65 5.025 ;
      RECT 20.97 3.495 21.14 3.665 ;
      RECT 19.23 6.685 19.4 6.855 ;
      RECT 18.8 7.055 18.97 7.225 ;
      RECT 18.8 7.795 18.97 7.965 ;
      RECT 16.045 7.8 16.215 7.97 ;
      RECT 15.675 2.76 15.845 2.93 ;
      RECT 15.675 5.95 15.845 6.12 ;
      RECT 15.055 0.91 15.225 1.08 ;
      RECT 15.055 2.39 15.225 2.56 ;
      RECT 15.055 6.32 15.225 6.49 ;
      RECT 15.055 7.8 15.225 7.97 ;
      RECT 14.685 2.76 14.855 2.93 ;
      RECT 14.685 5.95 14.855 6.12 ;
      RECT 13.695 2.025 13.865 2.195 ;
      RECT 13.695 6.685 13.865 6.855 ;
      RECT 13.265 0.915 13.435 1.085 ;
      RECT 13.265 1.655 13.435 1.825 ;
      RECT 13.265 7.055 13.435 7.225 ;
      RECT 13.265 7.795 13.435 7.965 ;
      RECT 12.89 2.395 13.06 2.565 ;
      RECT 12.89 6.315 13.06 6.485 ;
      RECT 9.7 3.835 9.87 4.005 ;
      RECT 9.7 5.875 9.87 6.045 ;
      RECT 9.36 2.815 9.53 2.985 ;
      RECT 9.02 6.555 9.19 6.725 ;
      RECT 8.85 5.875 9.02 6.045 ;
      RECT 8.34 5.875 8.51 6.045 ;
      RECT 7.66 3.155 7.83 3.325 ;
      RECT 7.66 6.555 7.83 6.725 ;
      RECT 6.98 2.815 7.15 2.985 ;
      RECT 6.97 5.875 7.14 6.045 ;
      RECT 6.52 4.855 6.69 5.025 ;
      RECT 6.5 2.305 6.67 2.475 ;
      RECT 6.13 2.82 6.3 2.99 ;
      RECT 5.62 2.82 5.79 2.99 ;
      RECT 5.62 3.835 5.79 4.005 ;
      RECT 5.28 6.555 5.45 6.725 ;
      RECT 4.26 2.815 4.43 2.985 ;
      RECT 4.26 4.855 4.43 5.025 ;
      RECT 3.75 3.495 3.92 3.665 ;
      RECT 2.01 6.685 2.18 6.855 ;
      RECT 1.58 7.055 1.75 7.225 ;
      RECT 1.58 7.795 1.75 7.965 ;
      RECT -1.83 7.055 -1.66 7.225 ;
      RECT -1.83 7.795 -1.66 7.965 ;
      RECT -2.205 6.315 -2.035 6.485 ;
    LAYER li1 ;
      RECT 84.925 5.02 85.095 6.49 ;
      RECT 84.925 6.315 85.1 6.485 ;
      RECT 84.555 1.74 84.725 2.93 ;
      RECT 84.555 1.74 85.025 1.91 ;
      RECT 84.555 6.97 85.025 7.14 ;
      RECT 84.555 5.95 84.725 7.14 ;
      RECT 83.565 1.74 83.735 2.93 ;
      RECT 83.565 1.74 84.035 1.91 ;
      RECT 83.565 6.97 84.035 7.14 ;
      RECT 83.565 5.95 83.735 7.14 ;
      RECT 81.715 2.635 81.885 3.865 ;
      RECT 81.77 0.855 81.94 2.805 ;
      RECT 81.715 0.575 81.885 1.025 ;
      RECT 81.715 7.855 81.885 8.305 ;
      RECT 81.77 6.075 81.94 8.025 ;
      RECT 81.715 5.015 81.885 6.245 ;
      RECT 81.195 0.575 81.365 3.865 ;
      RECT 81.195 2.075 81.6 2.405 ;
      RECT 81.195 1.235 81.6 1.565 ;
      RECT 81.195 5.015 81.365 8.305 ;
      RECT 81.195 7.315 81.6 7.645 ;
      RECT 81.195 6.475 81.6 6.805 ;
      RECT 78.93 3.495 79.31 4.175 ;
      RECT 79.14 2.365 79.31 4.175 ;
      RECT 77.06 2.365 77.29 3.035 ;
      RECT 77.06 2.365 79.31 2.535 ;
      RECT 78.59 2.045 78.76 2.535 ;
      RECT 78.58 3.155 78.75 4.005 ;
      RECT 77.665 3.155 78.97 3.325 ;
      RECT 78.725 2.705 78.97 3.325 ;
      RECT 77.665 2.785 77.835 3.325 ;
      RECT 77.46 2.785 77.835 2.955 ;
      RECT 77.64 6.265 78.335 6.895 ;
      RECT 78.165 4.685 78.335 6.895 ;
      RECT 78.07 4.685 78.4 5.665 ;
      RECT 77.67 3.495 78 4.175 ;
      RECT 76.76 3.495 77.16 4.175 ;
      RECT 76.76 3.495 78 3.665 ;
      RECT 76.26 3.075 76.58 4.175 ;
      RECT 76.26 3.075 76.71 3.325 ;
      RECT 76.26 3.075 76.89 3.245 ;
      RECT 76.72 2.025 76.89 3.245 ;
      RECT 76.72 2.025 77.675 2.195 ;
      RECT 76.26 6.265 76.955 6.895 ;
      RECT 76.785 4.685 76.955 6.895 ;
      RECT 76.69 4.685 77.02 5.665 ;
      RECT 76.28 5.825 76.615 6.075 ;
      RECT 75.735 5.825 76.07 6.075 ;
      RECT 75.735 5.875 76.615 6.045 ;
      RECT 75.395 6.265 76.09 6.895 ;
      RECT 75.395 4.685 75.565 6.895 ;
      RECT 75.33 4.685 75.66 5.665 ;
      RECT 74.89 3.205 75.22 4.16 ;
      RECT 74.89 3.205 75.57 3.375 ;
      RECT 75.4 1.965 75.57 3.375 ;
      RECT 75.31 1.965 75.64 2.605 ;
      RECT 74.37 3.205 74.7 4.16 ;
      RECT 74.02 3.205 74.7 3.375 ;
      RECT 74.02 1.965 74.19 3.375 ;
      RECT 73.95 1.965 74.28 2.605 ;
      RECT 74.16 5.875 74.33 6.725 ;
      RECT 73.435 5.825 73.77 6.075 ;
      RECT 73.435 5.875 74.33 6.045 ;
      RECT 73.5 2.785 73.85 3.035 ;
      RECT 72.98 2.785 73.31 3.035 ;
      RECT 72.98 2.815 73.85 2.985 ;
      RECT 73.095 6.265 73.79 6.895 ;
      RECT 73.095 4.685 73.265 6.895 ;
      RECT 73.03 4.685 73.36 5.665 ;
      RECT 72.56 3.195 72.89 4.175 ;
      RECT 72.56 1.965 72.81 4.175 ;
      RECT 72.56 1.965 72.89 2.595 ;
      RECT 69.51 5.015 69.68 8.305 ;
      RECT 69.51 7.315 69.915 7.645 ;
      RECT 69.51 6.475 69.915 6.805 ;
      RECT 67.705 5.02 67.875 6.49 ;
      RECT 67.705 6.315 67.88 6.485 ;
      RECT 67.335 1.74 67.505 2.93 ;
      RECT 67.335 1.74 67.805 1.91 ;
      RECT 67.335 6.97 67.805 7.14 ;
      RECT 67.335 5.95 67.505 7.14 ;
      RECT 66.345 1.74 66.515 2.93 ;
      RECT 66.345 1.74 66.815 1.91 ;
      RECT 66.345 6.97 66.815 7.14 ;
      RECT 66.345 5.95 66.515 7.14 ;
      RECT 64.495 2.635 64.665 3.865 ;
      RECT 64.55 0.855 64.72 2.805 ;
      RECT 64.495 0.575 64.665 1.025 ;
      RECT 64.495 7.855 64.665 8.305 ;
      RECT 64.55 6.075 64.72 8.025 ;
      RECT 64.495 5.015 64.665 6.245 ;
      RECT 63.975 0.575 64.145 3.865 ;
      RECT 63.975 2.075 64.38 2.405 ;
      RECT 63.975 1.235 64.38 1.565 ;
      RECT 63.975 5.015 64.145 8.305 ;
      RECT 63.975 7.315 64.38 7.645 ;
      RECT 63.975 6.475 64.38 6.805 ;
      RECT 61.71 3.495 62.09 4.175 ;
      RECT 61.92 2.365 62.09 4.175 ;
      RECT 59.84 2.365 60.07 3.035 ;
      RECT 59.84 2.365 62.09 2.535 ;
      RECT 61.37 2.045 61.54 2.535 ;
      RECT 61.36 3.155 61.53 4.005 ;
      RECT 60.445 3.155 61.75 3.325 ;
      RECT 61.505 2.705 61.75 3.325 ;
      RECT 60.445 2.785 60.615 3.325 ;
      RECT 60.24 2.785 60.615 2.955 ;
      RECT 60.42 6.265 61.115 6.895 ;
      RECT 60.945 4.685 61.115 6.895 ;
      RECT 60.85 4.685 61.18 5.665 ;
      RECT 60.45 3.495 60.78 4.175 ;
      RECT 59.54 3.495 59.94 4.175 ;
      RECT 59.54 3.495 60.78 3.665 ;
      RECT 59.04 3.075 59.36 4.175 ;
      RECT 59.04 3.075 59.49 3.325 ;
      RECT 59.04 3.075 59.67 3.245 ;
      RECT 59.5 2.025 59.67 3.245 ;
      RECT 59.5 2.025 60.455 2.195 ;
      RECT 59.04 6.265 59.735 6.895 ;
      RECT 59.565 4.685 59.735 6.895 ;
      RECT 59.47 4.685 59.8 5.665 ;
      RECT 59.06 5.825 59.395 6.075 ;
      RECT 58.515 5.825 58.85 6.075 ;
      RECT 58.515 5.875 59.395 6.045 ;
      RECT 58.175 6.265 58.87 6.895 ;
      RECT 58.175 4.685 58.345 6.895 ;
      RECT 58.11 4.685 58.44 5.665 ;
      RECT 57.67 3.205 58 4.16 ;
      RECT 57.67 3.205 58.35 3.375 ;
      RECT 58.18 1.965 58.35 3.375 ;
      RECT 58.09 1.965 58.42 2.605 ;
      RECT 57.15 3.205 57.48 4.16 ;
      RECT 56.8 3.205 57.48 3.375 ;
      RECT 56.8 1.965 56.97 3.375 ;
      RECT 56.73 1.965 57.06 2.605 ;
      RECT 56.94 5.875 57.11 6.725 ;
      RECT 56.215 5.825 56.55 6.075 ;
      RECT 56.215 5.875 57.11 6.045 ;
      RECT 56.28 2.785 56.63 3.035 ;
      RECT 55.76 2.785 56.09 3.035 ;
      RECT 55.76 2.815 56.63 2.985 ;
      RECT 55.875 6.265 56.57 6.895 ;
      RECT 55.875 4.685 56.045 6.895 ;
      RECT 55.81 4.685 56.14 5.665 ;
      RECT 55.34 3.195 55.67 4.175 ;
      RECT 55.34 1.965 55.59 4.175 ;
      RECT 55.34 1.965 55.67 2.595 ;
      RECT 52.29 5.015 52.46 8.305 ;
      RECT 52.29 7.315 52.695 7.645 ;
      RECT 52.29 6.475 52.695 6.805 ;
      RECT 50.485 5.02 50.655 6.49 ;
      RECT 50.485 6.315 50.66 6.485 ;
      RECT 50.115 1.74 50.285 2.93 ;
      RECT 50.115 1.74 50.585 1.91 ;
      RECT 50.115 6.97 50.585 7.14 ;
      RECT 50.115 5.95 50.285 7.14 ;
      RECT 49.125 1.74 49.295 2.93 ;
      RECT 49.125 1.74 49.595 1.91 ;
      RECT 49.125 6.97 49.595 7.14 ;
      RECT 49.125 5.95 49.295 7.14 ;
      RECT 47.275 2.635 47.445 3.865 ;
      RECT 47.33 0.855 47.5 2.805 ;
      RECT 47.275 0.575 47.445 1.025 ;
      RECT 47.275 7.855 47.445 8.305 ;
      RECT 47.33 6.075 47.5 8.025 ;
      RECT 47.275 5.015 47.445 6.245 ;
      RECT 46.755 0.575 46.925 3.865 ;
      RECT 46.755 2.075 47.16 2.405 ;
      RECT 46.755 1.235 47.16 1.565 ;
      RECT 46.755 5.015 46.925 8.305 ;
      RECT 46.755 7.315 47.16 7.645 ;
      RECT 46.755 6.475 47.16 6.805 ;
      RECT 44.49 3.495 44.87 4.175 ;
      RECT 44.7 2.365 44.87 4.175 ;
      RECT 42.62 2.365 42.85 3.035 ;
      RECT 42.62 2.365 44.87 2.535 ;
      RECT 44.15 2.045 44.32 2.535 ;
      RECT 44.14 3.155 44.31 4.005 ;
      RECT 43.225 3.155 44.53 3.325 ;
      RECT 44.285 2.705 44.53 3.325 ;
      RECT 43.225 2.785 43.395 3.325 ;
      RECT 43.02 2.785 43.395 2.955 ;
      RECT 43.2 6.265 43.895 6.895 ;
      RECT 43.725 4.685 43.895 6.895 ;
      RECT 43.63 4.685 43.96 5.665 ;
      RECT 43.23 3.495 43.56 4.175 ;
      RECT 42.32 3.495 42.72 4.175 ;
      RECT 42.32 3.495 43.56 3.665 ;
      RECT 41.82 3.075 42.14 4.175 ;
      RECT 41.82 3.075 42.27 3.325 ;
      RECT 41.82 3.075 42.45 3.245 ;
      RECT 42.28 2.025 42.45 3.245 ;
      RECT 42.28 2.025 43.235 2.195 ;
      RECT 41.82 6.265 42.515 6.895 ;
      RECT 42.345 4.685 42.515 6.895 ;
      RECT 42.25 4.685 42.58 5.665 ;
      RECT 41.84 5.825 42.175 6.075 ;
      RECT 41.295 5.825 41.63 6.075 ;
      RECT 41.295 5.875 42.175 6.045 ;
      RECT 40.955 6.265 41.65 6.895 ;
      RECT 40.955 4.685 41.125 6.895 ;
      RECT 40.89 4.685 41.22 5.665 ;
      RECT 40.45 3.205 40.78 4.16 ;
      RECT 40.45 3.205 41.13 3.375 ;
      RECT 40.96 1.965 41.13 3.375 ;
      RECT 40.87 1.965 41.2 2.605 ;
      RECT 39.93 3.205 40.26 4.16 ;
      RECT 39.58 3.205 40.26 3.375 ;
      RECT 39.58 1.965 39.75 3.375 ;
      RECT 39.51 1.965 39.84 2.605 ;
      RECT 39.72 5.875 39.89 6.725 ;
      RECT 38.995 5.825 39.33 6.075 ;
      RECT 38.995 5.875 39.89 6.045 ;
      RECT 39.06 2.785 39.41 3.035 ;
      RECT 38.54 2.785 38.87 3.035 ;
      RECT 38.54 2.815 39.41 2.985 ;
      RECT 38.655 6.265 39.35 6.895 ;
      RECT 38.655 4.685 38.825 6.895 ;
      RECT 38.59 4.685 38.92 5.665 ;
      RECT 38.12 3.195 38.45 4.175 ;
      RECT 38.12 1.965 38.37 4.175 ;
      RECT 38.12 1.965 38.45 2.595 ;
      RECT 35.07 5.015 35.24 8.305 ;
      RECT 35.07 7.315 35.475 7.645 ;
      RECT 35.07 6.475 35.475 6.805 ;
      RECT 33.265 5.02 33.435 6.49 ;
      RECT 33.265 6.315 33.44 6.485 ;
      RECT 32.895 1.74 33.065 2.93 ;
      RECT 32.895 1.74 33.365 1.91 ;
      RECT 32.895 6.97 33.365 7.14 ;
      RECT 32.895 5.95 33.065 7.14 ;
      RECT 31.905 1.74 32.075 2.93 ;
      RECT 31.905 1.74 32.375 1.91 ;
      RECT 31.905 6.97 32.375 7.14 ;
      RECT 31.905 5.95 32.075 7.14 ;
      RECT 30.055 2.635 30.225 3.865 ;
      RECT 30.11 0.855 30.28 2.805 ;
      RECT 30.055 0.575 30.225 1.025 ;
      RECT 30.055 7.855 30.225 8.305 ;
      RECT 30.11 6.075 30.28 8.025 ;
      RECT 30.055 5.015 30.225 6.245 ;
      RECT 29.535 0.575 29.705 3.865 ;
      RECT 29.535 2.075 29.94 2.405 ;
      RECT 29.535 1.235 29.94 1.565 ;
      RECT 29.535 5.015 29.705 8.305 ;
      RECT 29.535 7.315 29.94 7.645 ;
      RECT 29.535 6.475 29.94 6.805 ;
      RECT 27.27 3.495 27.65 4.175 ;
      RECT 27.48 2.365 27.65 4.175 ;
      RECT 25.4 2.365 25.63 3.035 ;
      RECT 25.4 2.365 27.65 2.535 ;
      RECT 26.93 2.045 27.1 2.535 ;
      RECT 26.92 3.155 27.09 4.005 ;
      RECT 26.005 3.155 27.31 3.325 ;
      RECT 27.065 2.705 27.31 3.325 ;
      RECT 26.005 2.785 26.175 3.325 ;
      RECT 25.8 2.785 26.175 2.955 ;
      RECT 25.98 6.265 26.675 6.895 ;
      RECT 26.505 4.685 26.675 6.895 ;
      RECT 26.41 4.685 26.74 5.665 ;
      RECT 26.01 3.495 26.34 4.175 ;
      RECT 25.1 3.495 25.5 4.175 ;
      RECT 25.1 3.495 26.34 3.665 ;
      RECT 24.6 3.075 24.92 4.175 ;
      RECT 24.6 3.075 25.05 3.325 ;
      RECT 24.6 3.075 25.23 3.245 ;
      RECT 25.06 2.025 25.23 3.245 ;
      RECT 25.06 2.025 26.015 2.195 ;
      RECT 24.6 6.265 25.295 6.895 ;
      RECT 25.125 4.685 25.295 6.895 ;
      RECT 25.03 4.685 25.36 5.665 ;
      RECT 24.62 5.825 24.955 6.075 ;
      RECT 24.075 5.825 24.41 6.075 ;
      RECT 24.075 5.875 24.955 6.045 ;
      RECT 23.735 6.265 24.43 6.895 ;
      RECT 23.735 4.685 23.905 6.895 ;
      RECT 23.67 4.685 24 5.665 ;
      RECT 23.23 3.205 23.56 4.16 ;
      RECT 23.23 3.205 23.91 3.375 ;
      RECT 23.74 1.965 23.91 3.375 ;
      RECT 23.65 1.965 23.98 2.605 ;
      RECT 22.71 3.205 23.04 4.16 ;
      RECT 22.36 3.205 23.04 3.375 ;
      RECT 22.36 1.965 22.53 3.375 ;
      RECT 22.29 1.965 22.62 2.605 ;
      RECT 22.5 5.875 22.67 6.725 ;
      RECT 21.775 5.825 22.11 6.075 ;
      RECT 21.775 5.875 22.67 6.045 ;
      RECT 21.84 2.785 22.19 3.035 ;
      RECT 21.32 2.785 21.65 3.035 ;
      RECT 21.32 2.815 22.19 2.985 ;
      RECT 21.435 6.265 22.13 6.895 ;
      RECT 21.435 4.685 21.605 6.895 ;
      RECT 21.37 4.685 21.7 5.665 ;
      RECT 20.9 3.195 21.23 4.175 ;
      RECT 20.9 1.965 21.15 4.175 ;
      RECT 20.9 1.965 21.23 2.595 ;
      RECT 17.85 5.015 18.02 8.305 ;
      RECT 17.85 7.315 18.255 7.645 ;
      RECT 17.85 6.475 18.255 6.805 ;
      RECT 16.045 5.02 16.215 6.49 ;
      RECT 16.045 6.315 16.22 6.485 ;
      RECT 15.675 1.74 15.845 2.93 ;
      RECT 15.675 1.74 16.145 1.91 ;
      RECT 15.675 6.97 16.145 7.14 ;
      RECT 15.675 5.95 15.845 7.14 ;
      RECT 14.685 1.74 14.855 2.93 ;
      RECT 14.685 1.74 15.155 1.91 ;
      RECT 14.685 6.97 15.155 7.14 ;
      RECT 14.685 5.95 14.855 7.14 ;
      RECT 12.835 2.635 13.005 3.865 ;
      RECT 12.89 0.855 13.06 2.805 ;
      RECT 12.835 0.575 13.005 1.025 ;
      RECT 12.835 7.855 13.005 8.305 ;
      RECT 12.89 6.075 13.06 8.025 ;
      RECT 12.835 5.015 13.005 6.245 ;
      RECT 12.315 0.575 12.485 3.865 ;
      RECT 12.315 2.075 12.72 2.405 ;
      RECT 12.315 1.235 12.72 1.565 ;
      RECT 12.315 5.015 12.485 8.305 ;
      RECT 12.315 7.315 12.72 7.645 ;
      RECT 12.315 6.475 12.72 6.805 ;
      RECT 10.05 3.495 10.43 4.175 ;
      RECT 10.26 2.365 10.43 4.175 ;
      RECT 8.18 2.365 8.41 3.035 ;
      RECT 8.18 2.365 10.43 2.535 ;
      RECT 9.71 2.045 9.88 2.535 ;
      RECT 9.7 3.155 9.87 4.005 ;
      RECT 8.785 3.155 10.09 3.325 ;
      RECT 9.845 2.705 10.09 3.325 ;
      RECT 8.785 2.785 8.955 3.325 ;
      RECT 8.58 2.785 8.955 2.955 ;
      RECT 8.76 6.265 9.455 6.895 ;
      RECT 9.285 4.685 9.455 6.895 ;
      RECT 9.19 4.685 9.52 5.665 ;
      RECT 8.79 3.495 9.12 4.175 ;
      RECT 7.88 3.495 8.28 4.175 ;
      RECT 7.88 3.495 9.12 3.665 ;
      RECT 7.38 3.075 7.7 4.175 ;
      RECT 7.38 3.075 7.83 3.325 ;
      RECT 7.38 3.075 8.01 3.245 ;
      RECT 7.84 2.025 8.01 3.245 ;
      RECT 7.84 2.025 8.795 2.195 ;
      RECT 7.38 6.265 8.075 6.895 ;
      RECT 7.905 4.685 8.075 6.895 ;
      RECT 7.81 4.685 8.14 5.665 ;
      RECT 7.4 5.825 7.735 6.075 ;
      RECT 6.855 5.825 7.19 6.075 ;
      RECT 6.855 5.875 7.735 6.045 ;
      RECT 6.515 6.265 7.21 6.895 ;
      RECT 6.515 4.685 6.685 6.895 ;
      RECT 6.45 4.685 6.78 5.665 ;
      RECT 6.01 3.205 6.34 4.16 ;
      RECT 6.01 3.205 6.69 3.375 ;
      RECT 6.52 1.965 6.69 3.375 ;
      RECT 6.43 1.965 6.76 2.605 ;
      RECT 5.49 3.205 5.82 4.16 ;
      RECT 5.14 3.205 5.82 3.375 ;
      RECT 5.14 1.965 5.31 3.375 ;
      RECT 5.07 1.965 5.4 2.605 ;
      RECT 5.28 5.875 5.45 6.725 ;
      RECT 4.555 5.825 4.89 6.075 ;
      RECT 4.555 5.875 5.45 6.045 ;
      RECT 4.62 2.785 4.97 3.035 ;
      RECT 4.1 2.785 4.43 3.035 ;
      RECT 4.1 2.815 4.97 2.985 ;
      RECT 4.215 6.265 4.91 6.895 ;
      RECT 4.215 4.685 4.385 6.895 ;
      RECT 4.15 4.685 4.48 5.665 ;
      RECT 3.68 3.195 4.01 4.175 ;
      RECT 3.68 1.965 3.93 4.175 ;
      RECT 3.68 1.965 4.01 2.595 ;
      RECT 0.63 5.015 0.8 8.305 ;
      RECT 0.63 7.315 1.035 7.645 ;
      RECT 0.63 6.475 1.035 6.805 ;
      RECT -2.26 7.855 -2.09 8.305 ;
      RECT -2.205 6.075 -2.035 8.025 ;
      RECT -2.26 5.015 -2.09 6.245 ;
      RECT -2.78 5.015 -2.61 8.305 ;
      RECT -2.78 7.315 -2.375 7.645 ;
      RECT -2.78 6.475 -2.375 6.805 ;
      RECT 84.925 7.8 85.095 8.31 ;
      RECT 83.935 0.57 84.105 1.08 ;
      RECT 83.935 2.39 84.105 3.86 ;
      RECT 83.935 5.02 84.105 6.49 ;
      RECT 83.935 7.8 84.105 8.31 ;
      RECT 82.575 0.575 82.745 3.865 ;
      RECT 82.575 5.015 82.745 8.305 ;
      RECT 82.145 0.575 82.315 1.085 ;
      RECT 82.145 1.655 82.315 3.865 ;
      RECT 82.145 5.015 82.315 7.225 ;
      RECT 82.145 7.795 82.315 8.305 ;
      RECT 78.505 5.825 78.84 6.095 ;
      RECT 78.005 2.785 78.555 2.985 ;
      RECT 77.66 5.825 77.995 6.075 ;
      RECT 77.125 5.825 77.46 6.095 ;
      RECT 75.74 2.785 76.09 3.035 ;
      RECT 74.88 2.785 75.23 3.035 ;
      RECT 74.36 2.785 74.71 3.035 ;
      RECT 70.89 5.015 71.06 8.305 ;
      RECT 70.46 5.015 70.63 7.225 ;
      RECT 70.46 7.795 70.63 8.305 ;
      RECT 67.705 7.8 67.875 8.31 ;
      RECT 66.715 0.57 66.885 1.08 ;
      RECT 66.715 2.39 66.885 3.86 ;
      RECT 66.715 5.02 66.885 6.49 ;
      RECT 66.715 7.8 66.885 8.31 ;
      RECT 65.355 0.575 65.525 3.865 ;
      RECT 65.355 5.015 65.525 8.305 ;
      RECT 64.925 0.575 65.095 1.085 ;
      RECT 64.925 1.655 65.095 3.865 ;
      RECT 64.925 5.015 65.095 7.225 ;
      RECT 64.925 7.795 65.095 8.305 ;
      RECT 61.285 5.825 61.62 6.095 ;
      RECT 60.785 2.785 61.335 2.985 ;
      RECT 60.44 5.825 60.775 6.075 ;
      RECT 59.905 5.825 60.24 6.095 ;
      RECT 58.52 2.785 58.87 3.035 ;
      RECT 57.66 2.785 58.01 3.035 ;
      RECT 57.14 2.785 57.49 3.035 ;
      RECT 53.67 5.015 53.84 8.305 ;
      RECT 53.24 5.015 53.41 7.225 ;
      RECT 53.24 7.795 53.41 8.305 ;
      RECT 50.485 7.8 50.655 8.31 ;
      RECT 49.495 0.57 49.665 1.08 ;
      RECT 49.495 2.39 49.665 3.86 ;
      RECT 49.495 5.02 49.665 6.49 ;
      RECT 49.495 7.8 49.665 8.31 ;
      RECT 48.135 0.575 48.305 3.865 ;
      RECT 48.135 5.015 48.305 8.305 ;
      RECT 47.705 0.575 47.875 1.085 ;
      RECT 47.705 1.655 47.875 3.865 ;
      RECT 47.705 5.015 47.875 7.225 ;
      RECT 47.705 7.795 47.875 8.305 ;
      RECT 44.065 5.825 44.4 6.095 ;
      RECT 43.565 2.785 44.115 2.985 ;
      RECT 43.22 5.825 43.555 6.075 ;
      RECT 42.685 5.825 43.02 6.095 ;
      RECT 41.3 2.785 41.65 3.035 ;
      RECT 40.44 2.785 40.79 3.035 ;
      RECT 39.92 2.785 40.27 3.035 ;
      RECT 36.45 5.015 36.62 8.305 ;
      RECT 36.02 5.015 36.19 7.225 ;
      RECT 36.02 7.795 36.19 8.305 ;
      RECT 33.265 7.8 33.435 8.31 ;
      RECT 32.275 0.57 32.445 1.08 ;
      RECT 32.275 2.39 32.445 3.86 ;
      RECT 32.275 5.02 32.445 6.49 ;
      RECT 32.275 7.8 32.445 8.31 ;
      RECT 30.915 0.575 31.085 3.865 ;
      RECT 30.915 5.015 31.085 8.305 ;
      RECT 30.485 0.575 30.655 1.085 ;
      RECT 30.485 1.655 30.655 3.865 ;
      RECT 30.485 5.015 30.655 7.225 ;
      RECT 30.485 7.795 30.655 8.305 ;
      RECT 26.845 5.825 27.18 6.095 ;
      RECT 26.345 2.785 26.895 2.985 ;
      RECT 26 5.825 26.335 6.075 ;
      RECT 25.465 5.825 25.8 6.095 ;
      RECT 24.08 2.785 24.43 3.035 ;
      RECT 23.22 2.785 23.57 3.035 ;
      RECT 22.7 2.785 23.05 3.035 ;
      RECT 19.23 5.015 19.4 8.305 ;
      RECT 18.8 5.015 18.97 7.225 ;
      RECT 18.8 7.795 18.97 8.305 ;
      RECT 16.045 7.8 16.215 8.31 ;
      RECT 15.055 0.57 15.225 1.08 ;
      RECT 15.055 2.39 15.225 3.86 ;
      RECT 15.055 5.02 15.225 6.49 ;
      RECT 15.055 7.8 15.225 8.31 ;
      RECT 13.695 0.575 13.865 3.865 ;
      RECT 13.695 5.015 13.865 8.305 ;
      RECT 13.265 0.575 13.435 1.085 ;
      RECT 13.265 1.655 13.435 3.865 ;
      RECT 13.265 5.015 13.435 7.225 ;
      RECT 13.265 7.795 13.435 8.305 ;
      RECT 9.625 5.825 9.96 6.095 ;
      RECT 9.125 2.785 9.675 2.985 ;
      RECT 8.78 5.825 9.115 6.075 ;
      RECT 8.245 5.825 8.58 6.095 ;
      RECT 6.86 2.785 7.21 3.035 ;
      RECT 6 2.785 6.35 3.035 ;
      RECT 5.48 2.785 5.83 3.035 ;
      RECT 2.01 5.015 2.18 8.305 ;
      RECT 1.58 5.015 1.75 7.225 ;
      RECT 1.58 7.795 1.75 8.305 ;
      RECT -1.83 5.015 -1.66 7.225 ;
      RECT -1.83 7.795 -1.66 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2ct_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2ea_8_b0r1
  CLASS BLOCK ;
  ORIGIN 3.275 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ea_8_b0r1 ;
  SIZE 84.425 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 15.31 0.915 15.48 1.085 ;
        RECT 15.305 0.91 15.475 1.08 ;
        RECT 15.305 2.39 15.475 2.56 ;
      LAYER li1 ;
        RECT 15.31 0.915 15.48 1.085 ;
        RECT 15.305 0.57 15.475 1.08 ;
        RECT 15.305 2.39 15.475 3.86 ;
      LAYER met1 ;
        RECT 15.245 2.36 15.535 2.59 ;
        RECT 15.245 0.88 15.535 1.11 ;
        RECT 15.305 0.88 15.475 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 31.635 0.915 31.805 1.085 ;
        RECT 31.63 0.91 31.8 1.08 ;
        RECT 31.63 2.39 31.8 2.56 ;
      LAYER li1 ;
        RECT 31.635 0.915 31.805 1.085 ;
        RECT 31.63 0.57 31.8 1.08 ;
        RECT 31.63 2.39 31.8 3.86 ;
      LAYER met1 ;
        RECT 31.57 2.36 31.86 2.59 ;
        RECT 31.57 0.88 31.86 1.11 ;
        RECT 31.63 0.88 31.8 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 47.96 0.915 48.13 1.085 ;
        RECT 47.955 0.91 48.125 1.08 ;
        RECT 47.955 2.39 48.125 2.56 ;
      LAYER li1 ;
        RECT 47.96 0.915 48.13 1.085 ;
        RECT 47.955 0.57 48.125 1.08 ;
        RECT 47.955 2.39 48.125 3.86 ;
      LAYER met1 ;
        RECT 47.895 2.36 48.185 2.59 ;
        RECT 47.895 0.88 48.185 1.11 ;
        RECT 47.955 0.88 48.125 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 64.285 0.915 64.455 1.085 ;
        RECT 64.28 0.91 64.45 1.08 ;
        RECT 64.28 2.39 64.45 2.56 ;
      LAYER li1 ;
        RECT 64.285 0.915 64.455 1.085 ;
        RECT 64.28 0.57 64.45 1.08 ;
        RECT 64.28 2.39 64.45 3.86 ;
      LAYER met1 ;
        RECT 64.22 2.36 64.51 2.59 ;
        RECT 64.22 0.88 64.51 1.11 ;
        RECT 64.28 0.88 64.45 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 80.61 0.915 80.78 1.085 ;
        RECT 80.605 0.91 80.775 1.08 ;
        RECT 80.605 2.39 80.775 2.56 ;
      LAYER li1 ;
        RECT 80.61 0.915 80.78 1.085 ;
        RECT 80.605 0.57 80.775 1.08 ;
        RECT 80.605 2.39 80.775 3.86 ;
      LAYER met1 ;
        RECT 80.545 2.36 80.835 2.59 ;
        RECT 80.545 0.88 80.835 1.11 ;
        RECT 80.605 0.88 80.775 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 11.155 1.66 11.325 2.935 ;
        RECT 11.155 5.945 11.325 7.22 ;
        RECT 5.54 5.945 5.71 7.22 ;
      LAYER met2 ;
        RECT 11.08 2.705 11.42 3.055 ;
        RECT 11.07 5.84 11.41 6.19 ;
        RECT 11.155 2.705 11.325 6.19 ;
      LAYER met1 ;
        RECT 11.08 2.765 11.555 2.935 ;
        RECT 11.08 2.705 11.42 3.055 ;
        RECT 5.48 5.945 11.555 6.115 ;
        RECT 11.07 5.84 11.41 6.19 ;
        RECT 5.48 5.915 5.77 6.145 ;
      LAYER via1 ;
        RECT 11.17 5.94 11.32 6.09 ;
        RECT 11.18 2.805 11.33 2.955 ;
      LAYER mcon ;
        RECT 5.54 5.945 5.71 6.115 ;
        RECT 11.155 5.945 11.325 6.115 ;
        RECT 11.155 2.765 11.325 2.935 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 27.48 1.66 27.65 2.935 ;
        RECT 27.48 5.945 27.65 7.22 ;
        RECT 21.865 5.945 22.035 7.22 ;
      LAYER met2 ;
        RECT 27.405 2.705 27.745 3.055 ;
        RECT 27.395 5.84 27.735 6.19 ;
        RECT 27.48 2.705 27.65 6.19 ;
      LAYER met1 ;
        RECT 27.405 2.765 27.88 2.935 ;
        RECT 27.405 2.705 27.745 3.055 ;
        RECT 21.805 5.945 27.88 6.115 ;
        RECT 27.395 5.84 27.735 6.19 ;
        RECT 21.805 5.915 22.095 6.145 ;
      LAYER via1 ;
        RECT 27.495 5.94 27.645 6.09 ;
        RECT 27.505 2.805 27.655 2.955 ;
      LAYER mcon ;
        RECT 21.865 5.945 22.035 6.115 ;
        RECT 27.48 5.945 27.65 6.115 ;
        RECT 27.48 2.765 27.65 2.935 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 43.805 1.66 43.975 2.935 ;
        RECT 43.805 5.945 43.975 7.22 ;
        RECT 38.19 5.945 38.36 7.22 ;
      LAYER met2 ;
        RECT 43.73 2.705 44.07 3.055 ;
        RECT 43.72 5.84 44.06 6.19 ;
        RECT 43.805 2.705 43.975 6.19 ;
      LAYER met1 ;
        RECT 43.73 2.765 44.205 2.935 ;
        RECT 43.73 2.705 44.07 3.055 ;
        RECT 38.13 5.945 44.205 6.115 ;
        RECT 43.72 5.84 44.06 6.19 ;
        RECT 38.13 5.915 38.42 6.145 ;
      LAYER via1 ;
        RECT 43.82 5.94 43.97 6.09 ;
        RECT 43.83 2.805 43.98 2.955 ;
      LAYER mcon ;
        RECT 38.19 5.945 38.36 6.115 ;
        RECT 43.805 5.945 43.975 6.115 ;
        RECT 43.805 2.765 43.975 2.935 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 60.13 1.66 60.3 2.935 ;
        RECT 60.13 5.945 60.3 7.22 ;
        RECT 54.515 5.945 54.685 7.22 ;
      LAYER met2 ;
        RECT 60.055 2.705 60.395 3.055 ;
        RECT 60.045 5.84 60.385 6.19 ;
        RECT 60.13 2.705 60.3 6.19 ;
      LAYER met1 ;
        RECT 60.055 2.765 60.53 2.935 ;
        RECT 60.055 2.705 60.395 3.055 ;
        RECT 54.455 5.945 60.53 6.115 ;
        RECT 60.045 5.84 60.385 6.19 ;
        RECT 54.455 5.915 54.745 6.145 ;
      LAYER via1 ;
        RECT 60.145 5.94 60.295 6.09 ;
        RECT 60.155 2.805 60.305 2.955 ;
      LAYER mcon ;
        RECT 54.515 5.945 54.685 6.115 ;
        RECT 60.13 5.945 60.3 6.115 ;
        RECT 60.13 2.765 60.3 2.935 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 76.455 1.66 76.625 2.935 ;
        RECT 76.455 5.945 76.625 7.22 ;
        RECT 70.84 5.945 71.01 7.22 ;
      LAYER met2 ;
        RECT 76.38 2.705 76.72 3.055 ;
        RECT 76.37 5.84 76.71 6.19 ;
        RECT 76.455 2.705 76.625 6.19 ;
      LAYER met1 ;
        RECT 76.38 2.765 76.855 2.935 ;
        RECT 76.38 2.705 76.72 3.055 ;
        RECT 70.78 5.945 76.855 6.115 ;
        RECT 76.37 5.84 76.71 6.19 ;
        RECT 70.78 5.915 71.07 6.145 ;
      LAYER via1 ;
        RECT 76.47 5.94 76.62 6.09 ;
        RECT 76.48 2.805 76.63 2.955 ;
      LAYER mcon ;
        RECT 70.84 5.945 71.01 6.115 ;
        RECT 76.455 5.945 76.625 6.115 ;
        RECT 76.455 2.765 76.625 2.935 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT -3.04 5.945 -2.87 7.22 ;
      LAYER met1 ;
        RECT -3.1 5.945 -2.64 6.115 ;
        RECT -3.1 5.915 -2.81 6.145 ;
      LAYER mcon ;
        RECT -3.04 5.945 -2.87 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT -3.275 4.135 81.15 4.745 ;
        RECT 79.015 4.13 80.995 4.75 ;
        RECT 80.175 3.4 80.345 5.48 ;
        RECT 79.185 3.4 79.355 5.48 ;
        RECT 76.445 3.405 76.615 5.475 ;
        RECT 74.655 3.635 74.825 4.745 ;
        RECT 73.695 3.635 73.865 4.745 ;
        RECT 71.255 3.635 71.425 4.745 ;
        RECT 70.83 4.135 71 5.475 ;
        RECT 70.255 3.635 70.425 4.745 ;
        RECT 69.295 3.635 69.465 4.745 ;
        RECT 66.855 3.635 67.025 4.745 ;
        RECT 62.69 4.13 64.67 4.75 ;
        RECT 63.85 3.4 64.02 5.48 ;
        RECT 62.86 3.4 63.03 5.48 ;
        RECT 60.12 3.405 60.29 5.475 ;
        RECT 58.33 3.635 58.5 4.745 ;
        RECT 57.37 3.635 57.54 4.745 ;
        RECT 54.93 3.635 55.1 4.745 ;
        RECT 54.505 4.135 54.675 5.475 ;
        RECT 53.93 3.635 54.1 4.745 ;
        RECT 52.97 3.635 53.14 4.745 ;
        RECT 50.53 3.635 50.7 4.745 ;
        RECT 46.365 4.13 48.345 4.75 ;
        RECT 47.525 3.4 47.695 5.48 ;
        RECT 46.535 3.4 46.705 5.48 ;
        RECT 43.795 3.405 43.965 5.475 ;
        RECT 42.005 3.635 42.175 4.745 ;
        RECT 41.045 3.635 41.215 4.745 ;
        RECT 38.605 3.635 38.775 4.745 ;
        RECT 38.18 4.135 38.35 5.475 ;
        RECT 37.605 3.635 37.775 4.745 ;
        RECT 36.645 3.635 36.815 4.745 ;
        RECT 34.205 3.635 34.375 4.745 ;
        RECT 30.04 4.13 32.02 4.75 ;
        RECT 31.2 3.4 31.37 5.48 ;
        RECT 30.21 3.4 30.38 5.48 ;
        RECT 27.47 3.405 27.64 5.475 ;
        RECT 25.68 3.635 25.85 4.745 ;
        RECT 24.72 3.635 24.89 4.745 ;
        RECT 22.28 3.635 22.45 4.745 ;
        RECT 21.855 4.135 22.025 5.475 ;
        RECT 21.28 3.635 21.45 4.745 ;
        RECT 20.32 3.635 20.49 4.745 ;
        RECT 17.88 3.635 18.05 4.745 ;
        RECT 13.715 4.13 15.695 4.75 ;
        RECT 14.875 3.4 15.045 5.48 ;
        RECT 13.885 3.4 14.055 5.48 ;
        RECT 11.145 3.405 11.315 5.475 ;
        RECT 9.355 3.635 9.525 4.745 ;
        RECT 8.395 3.635 8.565 4.745 ;
        RECT 5.955 3.635 6.125 4.745 ;
        RECT 5.53 4.135 5.7 5.475 ;
        RECT 4.955 3.635 5.125 4.745 ;
        RECT 3.995 3.635 4.165 4.745 ;
        RECT 1.555 3.635 1.725 4.745 ;
        RECT -1.24 4.135 -1.07 8.305 ;
        RECT -3.05 4.135 -2.88 5.475 ;
      LAYER met1 ;
        RECT -3.275 4.135 81.15 4.745 ;
        RECT 79.015 4.13 80.995 4.75 ;
        RECT 65.565 3.98 75.225 4.745 ;
        RECT 62.69 4.13 64.67 4.75 ;
        RECT 49.24 3.98 58.9 4.745 ;
        RECT 46.365 4.13 48.345 4.75 ;
        RECT 32.915 3.98 42.575 4.745 ;
        RECT 30.04 4.13 32.02 4.75 ;
        RECT 16.59 3.98 26.25 4.745 ;
        RECT 13.715 4.13 15.695 4.75 ;
        RECT 0.265 3.98 9.925 4.745 ;
        RECT -1.3 6.655 -1.01 6.885 ;
        RECT -1.47 6.685 -1.01 6.855 ;
      LAYER mcon ;
        RECT -1.24 6.685 -1.07 6.855 ;
        RECT -0.93 4.545 -0.76 4.715 ;
        RECT 0.41 4.135 0.58 4.305 ;
        RECT 0.87 4.135 1.04 4.305 ;
        RECT 1.33 4.135 1.5 4.305 ;
        RECT 1.79 4.135 1.96 4.305 ;
        RECT 2.25 4.135 2.42 4.305 ;
        RECT 2.71 4.135 2.88 4.305 ;
        RECT 3.17 4.135 3.34 4.305 ;
        RECT 3.63 4.135 3.8 4.305 ;
        RECT 4.09 4.135 4.26 4.305 ;
        RECT 4.55 4.135 4.72 4.305 ;
        RECT 5.01 4.135 5.18 4.305 ;
        RECT 5.47 4.135 5.64 4.305 ;
        RECT 5.93 4.135 6.1 4.305 ;
        RECT 6.39 4.135 6.56 4.305 ;
        RECT 6.85 4.135 7.02 4.305 ;
        RECT 7.31 4.135 7.48 4.305 ;
        RECT 7.65 4.545 7.82 4.715 ;
        RECT 7.77 4.135 7.94 4.305 ;
        RECT 8.23 4.135 8.4 4.305 ;
        RECT 8.69 4.135 8.86 4.305 ;
        RECT 9.15 4.135 9.32 4.305 ;
        RECT 9.61 4.135 9.78 4.305 ;
        RECT 13.265 4.545 13.435 4.715 ;
        RECT 13.265 4.165 13.435 4.335 ;
        RECT 13.965 4.55 14.135 4.72 ;
        RECT 13.965 4.16 14.135 4.33 ;
        RECT 14.955 4.55 15.125 4.72 ;
        RECT 14.955 4.16 15.125 4.33 ;
        RECT 16.735 4.135 16.905 4.305 ;
        RECT 17.195 4.135 17.365 4.305 ;
        RECT 17.655 4.135 17.825 4.305 ;
        RECT 18.115 4.135 18.285 4.305 ;
        RECT 18.575 4.135 18.745 4.305 ;
        RECT 19.035 4.135 19.205 4.305 ;
        RECT 19.495 4.135 19.665 4.305 ;
        RECT 19.955 4.135 20.125 4.305 ;
        RECT 20.415 4.135 20.585 4.305 ;
        RECT 20.875 4.135 21.045 4.305 ;
        RECT 21.335 4.135 21.505 4.305 ;
        RECT 21.795 4.135 21.965 4.305 ;
        RECT 22.255 4.135 22.425 4.305 ;
        RECT 22.715 4.135 22.885 4.305 ;
        RECT 23.175 4.135 23.345 4.305 ;
        RECT 23.635 4.135 23.805 4.305 ;
        RECT 23.975 4.545 24.145 4.715 ;
        RECT 24.095 4.135 24.265 4.305 ;
        RECT 24.555 4.135 24.725 4.305 ;
        RECT 25.015 4.135 25.185 4.305 ;
        RECT 25.475 4.135 25.645 4.305 ;
        RECT 25.935 4.135 26.105 4.305 ;
        RECT 29.59 4.545 29.76 4.715 ;
        RECT 29.59 4.165 29.76 4.335 ;
        RECT 30.29 4.55 30.46 4.72 ;
        RECT 30.29 4.16 30.46 4.33 ;
        RECT 31.28 4.55 31.45 4.72 ;
        RECT 31.28 4.16 31.45 4.33 ;
        RECT 33.06 4.135 33.23 4.305 ;
        RECT 33.52 4.135 33.69 4.305 ;
        RECT 33.98 4.135 34.15 4.305 ;
        RECT 34.44 4.135 34.61 4.305 ;
        RECT 34.9 4.135 35.07 4.305 ;
        RECT 35.36 4.135 35.53 4.305 ;
        RECT 35.82 4.135 35.99 4.305 ;
        RECT 36.28 4.135 36.45 4.305 ;
        RECT 36.74 4.135 36.91 4.305 ;
        RECT 37.2 4.135 37.37 4.305 ;
        RECT 37.66 4.135 37.83 4.305 ;
        RECT 38.12 4.135 38.29 4.305 ;
        RECT 38.58 4.135 38.75 4.305 ;
        RECT 39.04 4.135 39.21 4.305 ;
        RECT 39.5 4.135 39.67 4.305 ;
        RECT 39.96 4.135 40.13 4.305 ;
        RECT 40.3 4.545 40.47 4.715 ;
        RECT 40.42 4.135 40.59 4.305 ;
        RECT 40.88 4.135 41.05 4.305 ;
        RECT 41.34 4.135 41.51 4.305 ;
        RECT 41.8 4.135 41.97 4.305 ;
        RECT 42.26 4.135 42.43 4.305 ;
        RECT 45.915 4.545 46.085 4.715 ;
        RECT 45.915 4.165 46.085 4.335 ;
        RECT 46.615 4.55 46.785 4.72 ;
        RECT 46.615 4.16 46.785 4.33 ;
        RECT 47.605 4.55 47.775 4.72 ;
        RECT 47.605 4.16 47.775 4.33 ;
        RECT 49.385 4.135 49.555 4.305 ;
        RECT 49.845 4.135 50.015 4.305 ;
        RECT 50.305 4.135 50.475 4.305 ;
        RECT 50.765 4.135 50.935 4.305 ;
        RECT 51.225 4.135 51.395 4.305 ;
        RECT 51.685 4.135 51.855 4.305 ;
        RECT 52.145 4.135 52.315 4.305 ;
        RECT 52.605 4.135 52.775 4.305 ;
        RECT 53.065 4.135 53.235 4.305 ;
        RECT 53.525 4.135 53.695 4.305 ;
        RECT 53.985 4.135 54.155 4.305 ;
        RECT 54.445 4.135 54.615 4.305 ;
        RECT 54.905 4.135 55.075 4.305 ;
        RECT 55.365 4.135 55.535 4.305 ;
        RECT 55.825 4.135 55.995 4.305 ;
        RECT 56.285 4.135 56.455 4.305 ;
        RECT 56.625 4.545 56.795 4.715 ;
        RECT 56.745 4.135 56.915 4.305 ;
        RECT 57.205 4.135 57.375 4.305 ;
        RECT 57.665 4.135 57.835 4.305 ;
        RECT 58.125 4.135 58.295 4.305 ;
        RECT 58.585 4.135 58.755 4.305 ;
        RECT 62.24 4.545 62.41 4.715 ;
        RECT 62.24 4.165 62.41 4.335 ;
        RECT 62.94 4.55 63.11 4.72 ;
        RECT 62.94 4.16 63.11 4.33 ;
        RECT 63.93 4.55 64.1 4.72 ;
        RECT 63.93 4.16 64.1 4.33 ;
        RECT 65.71 4.135 65.88 4.305 ;
        RECT 66.17 4.135 66.34 4.305 ;
        RECT 66.63 4.135 66.8 4.305 ;
        RECT 67.09 4.135 67.26 4.305 ;
        RECT 67.55 4.135 67.72 4.305 ;
        RECT 68.01 4.135 68.18 4.305 ;
        RECT 68.47 4.135 68.64 4.305 ;
        RECT 68.93 4.135 69.1 4.305 ;
        RECT 69.39 4.135 69.56 4.305 ;
        RECT 69.85 4.135 70.02 4.305 ;
        RECT 70.31 4.135 70.48 4.305 ;
        RECT 70.77 4.135 70.94 4.305 ;
        RECT 71.23 4.135 71.4 4.305 ;
        RECT 71.69 4.135 71.86 4.305 ;
        RECT 72.15 4.135 72.32 4.305 ;
        RECT 72.61 4.135 72.78 4.305 ;
        RECT 72.95 4.545 73.12 4.715 ;
        RECT 73.07 4.135 73.24 4.305 ;
        RECT 73.53 4.135 73.7 4.305 ;
        RECT 73.99 4.135 74.16 4.305 ;
        RECT 74.45 4.135 74.62 4.305 ;
        RECT 74.91 4.135 75.08 4.305 ;
        RECT 78.565 4.545 78.735 4.715 ;
        RECT 78.565 4.165 78.735 4.335 ;
        RECT 79.265 4.55 79.435 4.72 ;
        RECT 79.265 4.16 79.435 4.33 ;
        RECT 80.255 4.55 80.425 4.72 ;
        RECT 80.255 4.16 80.425 4.33 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 74.455 2.975 74.785 3.705 ;
        RECT 58.13 2.975 58.46 3.705 ;
        RECT 41.805 2.975 42.135 3.705 ;
        RECT 25.48 2.975 25.81 3.705 ;
        RECT 9.155 2.975 9.485 3.705 ;
      LAYER li1 ;
        RECT 80.97 0 81.15 0.305 ;
        RECT -3.275 0 81.15 0.3 ;
        RECT 80.175 0 80.345 0.93 ;
        RECT 79.185 0 79.355 0.93 ;
        RECT 64.645 0 79.02 0.305 ;
        RECT 76.445 0 76.615 0.935 ;
        RECT 65.565 0 75.38 1.585 ;
        RECT 73.695 0 73.865 2.085 ;
        RECT 71.735 0 71.905 2.085 ;
        RECT 71.665 0 71.905 1.595 ;
        RECT 70.115 0 70.31 1.595 ;
        RECT 69.295 0 69.465 2.085 ;
        RECT 68.335 0 68.505 2.085 ;
        RECT 67.99 0 68.185 1.595 ;
        RECT 67.815 0 67.985 2.085 ;
        RECT 66.855 0 67.025 2.085 ;
        RECT 65.895 0 66.065 2.085 ;
        RECT 65.69 0 65.885 1.595 ;
        RECT 63.85 0 64.02 0.93 ;
        RECT 62.86 0 63.03 0.93 ;
        RECT 48.32 0 62.695 0.305 ;
        RECT 60.12 0 60.29 0.935 ;
        RECT 49.24 0 59.055 1.585 ;
        RECT 57.37 0 57.54 2.085 ;
        RECT 55.41 0 55.58 2.085 ;
        RECT 55.34 0 55.58 1.595 ;
        RECT 53.79 0 53.985 1.595 ;
        RECT 52.97 0 53.14 2.085 ;
        RECT 52.01 0 52.18 2.085 ;
        RECT 51.665 0 51.86 1.595 ;
        RECT 51.49 0 51.66 2.085 ;
        RECT 50.53 0 50.7 2.085 ;
        RECT 49.57 0 49.74 2.085 ;
        RECT 49.365 0 49.56 1.595 ;
        RECT 47.525 0 47.695 0.93 ;
        RECT 46.535 0 46.705 0.93 ;
        RECT 31.995 0 46.37 0.305 ;
        RECT 43.795 0 43.965 0.935 ;
        RECT 32.915 0 42.73 1.585 ;
        RECT 41.045 0 41.215 2.085 ;
        RECT 39.085 0 39.255 2.085 ;
        RECT 39.015 0 39.255 1.595 ;
        RECT 37.465 0 37.66 1.595 ;
        RECT 36.645 0 36.815 2.085 ;
        RECT 35.685 0 35.855 2.085 ;
        RECT 35.34 0 35.535 1.595 ;
        RECT 35.165 0 35.335 2.085 ;
        RECT 34.205 0 34.375 2.085 ;
        RECT 33.245 0 33.415 2.085 ;
        RECT 33.04 0 33.235 1.595 ;
        RECT 31.2 0 31.37 0.93 ;
        RECT 30.21 0 30.38 0.93 ;
        RECT 15.67 0 30.045 0.305 ;
        RECT 27.47 0 27.64 0.935 ;
        RECT 16.59 0 26.405 1.585 ;
        RECT 24.72 0 24.89 2.085 ;
        RECT 22.76 0 22.93 2.085 ;
        RECT 22.69 0 22.93 1.595 ;
        RECT 21.14 0 21.335 1.595 ;
        RECT 20.32 0 20.49 2.085 ;
        RECT 19.36 0 19.53 2.085 ;
        RECT 19.015 0 19.21 1.595 ;
        RECT 18.84 0 19.01 2.085 ;
        RECT 17.88 0 18.05 2.085 ;
        RECT 16.92 0 17.09 2.085 ;
        RECT 16.715 0 16.91 1.595 ;
        RECT 14.875 0 15.045 0.93 ;
        RECT 13.885 0 14.055 0.93 ;
        RECT -3.275 0 13.72 0.305 ;
        RECT 11.145 0 11.315 0.935 ;
        RECT 0.265 0 10.08 1.585 ;
        RECT 8.395 0 8.565 2.085 ;
        RECT 6.435 0 6.605 2.085 ;
        RECT 6.365 0 6.605 1.595 ;
        RECT 4.815 0 5.01 1.595 ;
        RECT 3.995 0 4.165 2.085 ;
        RECT 3.035 0 3.205 2.085 ;
        RECT 2.69 0 2.885 1.595 ;
        RECT 2.515 0 2.685 2.085 ;
        RECT 1.555 0 1.725 2.085 ;
        RECT 0.595 0 0.765 2.085 ;
        RECT 0.39 0 0.585 1.595 ;
        RECT -3.275 8.58 81.15 8.88 ;
        RECT 80.97 8.575 81.15 8.88 ;
        RECT 80.175 7.95 80.345 8.88 ;
        RECT 79.185 7.95 79.355 8.88 ;
        RECT 64.645 8.575 79.02 8.88 ;
        RECT 76.445 7.945 76.615 8.88 ;
        RECT 70.83 7.945 71 8.88 ;
        RECT 63.85 7.95 64.02 8.88 ;
        RECT 62.86 7.95 63.03 8.88 ;
        RECT 48.32 8.575 62.695 8.88 ;
        RECT 60.12 7.945 60.29 8.88 ;
        RECT 54.505 7.945 54.675 8.88 ;
        RECT 47.525 7.95 47.695 8.88 ;
        RECT 46.535 7.95 46.705 8.88 ;
        RECT 31.995 8.575 46.37 8.88 ;
        RECT 43.795 7.945 43.965 8.88 ;
        RECT 38.18 7.945 38.35 8.88 ;
        RECT 31.2 7.95 31.37 8.88 ;
        RECT 30.21 7.95 30.38 8.88 ;
        RECT 15.67 8.575 30.045 8.88 ;
        RECT 27.47 7.945 27.64 8.88 ;
        RECT 21.855 7.945 22.025 8.88 ;
        RECT 14.875 7.95 15.045 8.88 ;
        RECT 13.885 7.95 14.055 8.88 ;
        RECT -3.275 8.575 13.72 8.88 ;
        RECT 11.145 7.945 11.315 8.88 ;
        RECT 5.53 7.945 5.7 8.88 ;
        RECT -3.05 7.945 -2.88 8.88 ;
        RECT 74.655 2.575 74.825 2.945 ;
        RECT 74.335 2.575 74.825 2.745 ;
        RECT 72.695 2.575 72.865 2.945 ;
        RECT 72.375 2.575 72.865 2.745 ;
        RECT 71.835 6.075 72.005 8.025 ;
        RECT 71.78 7.855 71.95 8.305 ;
        RECT 71.78 5.015 71.95 6.245 ;
        RECT 58.33 2.575 58.5 2.945 ;
        RECT 58.01 2.575 58.5 2.745 ;
        RECT 56.37 2.575 56.54 2.945 ;
        RECT 56.05 2.575 56.54 2.745 ;
        RECT 55.51 6.075 55.68 8.025 ;
        RECT 55.455 7.855 55.625 8.305 ;
        RECT 55.455 5.015 55.625 6.245 ;
        RECT 42.005 2.575 42.175 2.945 ;
        RECT 41.685 2.575 42.175 2.745 ;
        RECT 40.045 2.575 40.215 2.945 ;
        RECT 39.725 2.575 40.215 2.745 ;
        RECT 39.185 6.075 39.355 8.025 ;
        RECT 39.13 7.855 39.3 8.305 ;
        RECT 39.13 5.015 39.3 6.245 ;
        RECT 25.68 2.575 25.85 2.945 ;
        RECT 25.36 2.575 25.85 2.745 ;
        RECT 23.72 2.575 23.89 2.945 ;
        RECT 23.4 2.575 23.89 2.745 ;
        RECT 22.86 6.075 23.03 8.025 ;
        RECT 22.805 7.855 22.975 8.305 ;
        RECT 22.805 5.015 22.975 6.245 ;
        RECT 9.355 2.575 9.525 2.945 ;
        RECT 9.035 2.575 9.525 2.745 ;
        RECT 7.395 2.575 7.565 2.945 ;
        RECT 7.075 2.575 7.565 2.745 ;
        RECT 6.535 6.075 6.705 8.025 ;
        RECT 6.48 7.855 6.65 8.305 ;
        RECT 6.48 5.015 6.65 6.245 ;
      LAYER met2 ;
        RECT 74.48 2.955 74.76 3.325 ;
        RECT 74.49 2.7 74.75 3.325 ;
        RECT 58.155 2.955 58.435 3.325 ;
        RECT 58.165 2.7 58.425 3.325 ;
        RECT 41.83 2.955 42.11 3.325 ;
        RECT 41.84 2.7 42.1 3.325 ;
        RECT 25.505 2.955 25.785 3.325 ;
        RECT 25.515 2.7 25.775 3.325 ;
        RECT 9.18 2.955 9.46 3.325 ;
        RECT 9.19 2.7 9.45 3.325 ;
      LAYER met1 ;
        RECT 80.97 0 81.15 0.305 ;
        RECT -3.275 0 81.15 0.3 ;
        RECT 64.645 0 79.02 0.305 ;
        RECT 75.195 0 75.38 2.945 ;
        RECT 74.43 2.79 75.38 2.945 ;
        RECT 74.46 2.76 75.38 2.945 ;
        RECT 65.565 0 75.38 1.74 ;
        RECT 74.46 2.745 74.885 2.975 ;
        RECT 74.46 2.73 74.78 2.99 ;
        RECT 72.97 2.93 74.735 3.055 ;
        RECT 72.97 2.93 74.57 3.07 ;
        RECT 72.635 2.79 73.11 2.975 ;
        RECT 72.635 2.745 72.925 2.975 ;
        RECT 48.32 0 62.695 0.305 ;
        RECT 58.87 0 59.055 2.945 ;
        RECT 58.105 2.79 59.055 2.945 ;
        RECT 58.135 2.76 59.055 2.945 ;
        RECT 49.24 0 59.055 1.74 ;
        RECT 58.135 2.745 58.56 2.975 ;
        RECT 58.135 2.73 58.455 2.99 ;
        RECT 56.645 2.93 58.41 3.055 ;
        RECT 56.645 2.93 58.245 3.07 ;
        RECT 56.31 2.79 56.785 2.975 ;
        RECT 56.31 2.745 56.6 2.975 ;
        RECT 31.995 0 46.37 0.305 ;
        RECT 42.545 0 42.73 2.945 ;
        RECT 41.78 2.79 42.73 2.945 ;
        RECT 41.81 2.76 42.73 2.945 ;
        RECT 32.915 0 42.73 1.74 ;
        RECT 41.81 2.745 42.235 2.975 ;
        RECT 41.81 2.73 42.13 2.99 ;
        RECT 40.32 2.93 42.085 3.055 ;
        RECT 40.32 2.93 41.92 3.07 ;
        RECT 39.985 2.79 40.46 2.975 ;
        RECT 39.985 2.745 40.275 2.975 ;
        RECT 15.67 0 30.045 0.305 ;
        RECT 26.22 0 26.405 2.945 ;
        RECT 25.455 2.79 26.405 2.945 ;
        RECT 25.485 2.76 26.405 2.945 ;
        RECT 16.59 0 26.405 1.74 ;
        RECT 25.485 2.745 25.91 2.975 ;
        RECT 25.485 2.73 25.805 2.99 ;
        RECT 23.995 2.93 25.76 3.055 ;
        RECT 23.995 2.93 25.595 3.07 ;
        RECT 23.66 2.79 24.135 2.975 ;
        RECT 23.66 2.745 23.95 2.975 ;
        RECT -3.275 0 13.72 0.305 ;
        RECT 9.895 0 10.08 2.945 ;
        RECT 9.13 2.79 10.08 2.945 ;
        RECT 9.16 2.76 10.08 2.945 ;
        RECT 0.265 0 10.08 1.74 ;
        RECT 9.16 2.745 9.585 2.975 ;
        RECT 9.16 2.73 9.48 2.99 ;
        RECT 7.67 2.93 9.435 3.055 ;
        RECT 7.67 2.93 9.27 3.07 ;
        RECT 7.335 2.79 7.81 2.975 ;
        RECT 7.335 2.745 7.625 2.975 ;
        RECT -3.275 8.58 81.15 8.88 ;
        RECT 80.97 8.575 81.15 8.88 ;
        RECT 64.645 8.575 79.02 8.88 ;
        RECT 71.775 6.285 72.065 6.515 ;
        RECT 71.4 6.315 72.065 6.485 ;
        RECT 71.4 6.315 71.575 8.88 ;
        RECT 48.32 8.575 62.695 8.88 ;
        RECT 55.45 6.285 55.74 6.515 ;
        RECT 55.075 6.315 55.74 6.485 ;
        RECT 55.075 6.315 55.25 8.88 ;
        RECT 31.995 8.575 46.37 8.88 ;
        RECT 39.125 6.285 39.415 6.515 ;
        RECT 38.75 6.315 39.415 6.485 ;
        RECT 38.75 6.315 38.925 8.88 ;
        RECT 15.67 8.575 30.045 8.88 ;
        RECT 22.8 6.285 23.09 6.515 ;
        RECT 22.425 6.315 23.09 6.485 ;
        RECT 22.425 6.315 22.6 8.88 ;
        RECT -3.275 8.575 13.72 8.88 ;
        RECT 6.475 6.285 6.765 6.515 ;
        RECT 6.1 6.315 6.765 6.485 ;
        RECT 6.1 6.315 6.275 8.88 ;
      LAYER via2 ;
        RECT 9.22 3.04 9.42 3.24 ;
        RECT 25.545 3.04 25.745 3.24 ;
        RECT 41.87 3.04 42.07 3.24 ;
        RECT 58.195 3.04 58.395 3.24 ;
        RECT 74.52 3.04 74.72 3.24 ;
      LAYER via1 ;
        RECT 9.245 2.785 9.395 2.935 ;
        RECT 25.57 2.785 25.72 2.935 ;
        RECT 41.895 2.785 42.045 2.935 ;
        RECT 58.22 2.785 58.37 2.935 ;
        RECT 74.545 2.785 74.695 2.935 ;
      LAYER mcon ;
        RECT -2.97 8.605 -2.8 8.775 ;
        RECT -2.29 8.605 -2.12 8.775 ;
        RECT -1.61 8.605 -1.44 8.775 ;
        RECT -0.93 8.605 -0.76 8.775 ;
        RECT 0.41 1.415 0.58 1.585 ;
        RECT 0.87 1.415 1.04 1.585 ;
        RECT 1.33 1.415 1.5 1.585 ;
        RECT 1.79 1.415 1.96 1.585 ;
        RECT 2.25 1.415 2.42 1.585 ;
        RECT 2.71 1.415 2.88 1.585 ;
        RECT 3.17 1.415 3.34 1.585 ;
        RECT 3.63 1.415 3.8 1.585 ;
        RECT 4.09 1.415 4.26 1.585 ;
        RECT 4.55 1.415 4.72 1.585 ;
        RECT 5.01 1.415 5.18 1.585 ;
        RECT 5.47 1.415 5.64 1.585 ;
        RECT 5.61 8.605 5.78 8.775 ;
        RECT 5.93 1.415 6.1 1.585 ;
        RECT 6.29 8.605 6.46 8.775 ;
        RECT 6.39 1.415 6.56 1.585 ;
        RECT 6.535 6.315 6.705 6.485 ;
        RECT 6.85 1.415 7.02 1.585 ;
        RECT 6.97 8.605 7.14 8.775 ;
        RECT 7.31 1.415 7.48 1.585 ;
        RECT 7.395 2.775 7.565 2.945 ;
        RECT 7.65 8.605 7.82 8.775 ;
        RECT 7.77 1.415 7.94 1.585 ;
        RECT 8.23 1.415 8.4 1.585 ;
        RECT 8.69 1.415 8.86 1.585 ;
        RECT 9.15 1.415 9.32 1.585 ;
        RECT 9.355 2.775 9.525 2.945 ;
        RECT 9.61 1.415 9.78 1.585 ;
        RECT 11.225 8.605 11.395 8.775 ;
        RECT 11.225 0.105 11.395 0.275 ;
        RECT 11.905 8.605 12.075 8.775 ;
        RECT 11.905 0.105 12.075 0.275 ;
        RECT 12.585 8.605 12.755 8.775 ;
        RECT 12.585 0.105 12.755 0.275 ;
        RECT 13.265 8.605 13.435 8.775 ;
        RECT 13.265 0.105 13.435 0.275 ;
        RECT 13.965 8.61 14.135 8.78 ;
        RECT 13.965 0.1 14.135 0.27 ;
        RECT 14.955 8.61 15.125 8.78 ;
        RECT 14.955 0.1 15.125 0.27 ;
        RECT 16.735 1.415 16.905 1.585 ;
        RECT 17.195 1.415 17.365 1.585 ;
        RECT 17.655 1.415 17.825 1.585 ;
        RECT 18.115 1.415 18.285 1.585 ;
        RECT 18.575 1.415 18.745 1.585 ;
        RECT 19.035 1.415 19.205 1.585 ;
        RECT 19.495 1.415 19.665 1.585 ;
        RECT 19.955 1.415 20.125 1.585 ;
        RECT 20.415 1.415 20.585 1.585 ;
        RECT 20.875 1.415 21.045 1.585 ;
        RECT 21.335 1.415 21.505 1.585 ;
        RECT 21.795 1.415 21.965 1.585 ;
        RECT 21.935 8.605 22.105 8.775 ;
        RECT 22.255 1.415 22.425 1.585 ;
        RECT 22.615 8.605 22.785 8.775 ;
        RECT 22.715 1.415 22.885 1.585 ;
        RECT 22.86 6.315 23.03 6.485 ;
        RECT 23.175 1.415 23.345 1.585 ;
        RECT 23.295 8.605 23.465 8.775 ;
        RECT 23.635 1.415 23.805 1.585 ;
        RECT 23.72 2.775 23.89 2.945 ;
        RECT 23.975 8.605 24.145 8.775 ;
        RECT 24.095 1.415 24.265 1.585 ;
        RECT 24.555 1.415 24.725 1.585 ;
        RECT 25.015 1.415 25.185 1.585 ;
        RECT 25.475 1.415 25.645 1.585 ;
        RECT 25.68 2.775 25.85 2.945 ;
        RECT 25.935 1.415 26.105 1.585 ;
        RECT 27.55 8.605 27.72 8.775 ;
        RECT 27.55 0.105 27.72 0.275 ;
        RECT 28.23 8.605 28.4 8.775 ;
        RECT 28.23 0.105 28.4 0.275 ;
        RECT 28.91 8.605 29.08 8.775 ;
        RECT 28.91 0.105 29.08 0.275 ;
        RECT 29.59 8.605 29.76 8.775 ;
        RECT 29.59 0.105 29.76 0.275 ;
        RECT 30.29 8.61 30.46 8.78 ;
        RECT 30.29 0.1 30.46 0.27 ;
        RECT 31.28 8.61 31.45 8.78 ;
        RECT 31.28 0.1 31.45 0.27 ;
        RECT 33.06 1.415 33.23 1.585 ;
        RECT 33.52 1.415 33.69 1.585 ;
        RECT 33.98 1.415 34.15 1.585 ;
        RECT 34.44 1.415 34.61 1.585 ;
        RECT 34.9 1.415 35.07 1.585 ;
        RECT 35.36 1.415 35.53 1.585 ;
        RECT 35.82 1.415 35.99 1.585 ;
        RECT 36.28 1.415 36.45 1.585 ;
        RECT 36.74 1.415 36.91 1.585 ;
        RECT 37.2 1.415 37.37 1.585 ;
        RECT 37.66 1.415 37.83 1.585 ;
        RECT 38.12 1.415 38.29 1.585 ;
        RECT 38.26 8.605 38.43 8.775 ;
        RECT 38.58 1.415 38.75 1.585 ;
        RECT 38.94 8.605 39.11 8.775 ;
        RECT 39.04 1.415 39.21 1.585 ;
        RECT 39.185 6.315 39.355 6.485 ;
        RECT 39.5 1.415 39.67 1.585 ;
        RECT 39.62 8.605 39.79 8.775 ;
        RECT 39.96 1.415 40.13 1.585 ;
        RECT 40.045 2.775 40.215 2.945 ;
        RECT 40.3 8.605 40.47 8.775 ;
        RECT 40.42 1.415 40.59 1.585 ;
        RECT 40.88 1.415 41.05 1.585 ;
        RECT 41.34 1.415 41.51 1.585 ;
        RECT 41.8 1.415 41.97 1.585 ;
        RECT 42.005 2.775 42.175 2.945 ;
        RECT 42.26 1.415 42.43 1.585 ;
        RECT 43.875 8.605 44.045 8.775 ;
        RECT 43.875 0.105 44.045 0.275 ;
        RECT 44.555 8.605 44.725 8.775 ;
        RECT 44.555 0.105 44.725 0.275 ;
        RECT 45.235 8.605 45.405 8.775 ;
        RECT 45.235 0.105 45.405 0.275 ;
        RECT 45.915 8.605 46.085 8.775 ;
        RECT 45.915 0.105 46.085 0.275 ;
        RECT 46.615 8.61 46.785 8.78 ;
        RECT 46.615 0.1 46.785 0.27 ;
        RECT 47.605 8.61 47.775 8.78 ;
        RECT 47.605 0.1 47.775 0.27 ;
        RECT 49.385 1.415 49.555 1.585 ;
        RECT 49.845 1.415 50.015 1.585 ;
        RECT 50.305 1.415 50.475 1.585 ;
        RECT 50.765 1.415 50.935 1.585 ;
        RECT 51.225 1.415 51.395 1.585 ;
        RECT 51.685 1.415 51.855 1.585 ;
        RECT 52.145 1.415 52.315 1.585 ;
        RECT 52.605 1.415 52.775 1.585 ;
        RECT 53.065 1.415 53.235 1.585 ;
        RECT 53.525 1.415 53.695 1.585 ;
        RECT 53.985 1.415 54.155 1.585 ;
        RECT 54.445 1.415 54.615 1.585 ;
        RECT 54.585 8.605 54.755 8.775 ;
        RECT 54.905 1.415 55.075 1.585 ;
        RECT 55.265 8.605 55.435 8.775 ;
        RECT 55.365 1.415 55.535 1.585 ;
        RECT 55.51 6.315 55.68 6.485 ;
        RECT 55.825 1.415 55.995 1.585 ;
        RECT 55.945 8.605 56.115 8.775 ;
        RECT 56.285 1.415 56.455 1.585 ;
        RECT 56.37 2.775 56.54 2.945 ;
        RECT 56.625 8.605 56.795 8.775 ;
        RECT 56.745 1.415 56.915 1.585 ;
        RECT 57.205 1.415 57.375 1.585 ;
        RECT 57.665 1.415 57.835 1.585 ;
        RECT 58.125 1.415 58.295 1.585 ;
        RECT 58.33 2.775 58.5 2.945 ;
        RECT 58.585 1.415 58.755 1.585 ;
        RECT 60.2 8.605 60.37 8.775 ;
        RECT 60.2 0.105 60.37 0.275 ;
        RECT 60.88 8.605 61.05 8.775 ;
        RECT 60.88 0.105 61.05 0.275 ;
        RECT 61.56 8.605 61.73 8.775 ;
        RECT 61.56 0.105 61.73 0.275 ;
        RECT 62.24 8.605 62.41 8.775 ;
        RECT 62.24 0.105 62.41 0.275 ;
        RECT 62.94 8.61 63.11 8.78 ;
        RECT 62.94 0.1 63.11 0.27 ;
        RECT 63.93 8.61 64.1 8.78 ;
        RECT 63.93 0.1 64.1 0.27 ;
        RECT 65.71 1.415 65.88 1.585 ;
        RECT 66.17 1.415 66.34 1.585 ;
        RECT 66.63 1.415 66.8 1.585 ;
        RECT 67.09 1.415 67.26 1.585 ;
        RECT 67.55 1.415 67.72 1.585 ;
        RECT 68.01 1.415 68.18 1.585 ;
        RECT 68.47 1.415 68.64 1.585 ;
        RECT 68.93 1.415 69.1 1.585 ;
        RECT 69.39 1.415 69.56 1.585 ;
        RECT 69.85 1.415 70.02 1.585 ;
        RECT 70.31 1.415 70.48 1.585 ;
        RECT 70.77 1.415 70.94 1.585 ;
        RECT 70.91 8.605 71.08 8.775 ;
        RECT 71.23 1.415 71.4 1.585 ;
        RECT 71.59 8.605 71.76 8.775 ;
        RECT 71.69 1.415 71.86 1.585 ;
        RECT 71.835 6.315 72.005 6.485 ;
        RECT 72.15 1.415 72.32 1.585 ;
        RECT 72.27 8.605 72.44 8.775 ;
        RECT 72.61 1.415 72.78 1.585 ;
        RECT 72.695 2.775 72.865 2.945 ;
        RECT 72.95 8.605 73.12 8.775 ;
        RECT 73.07 1.415 73.24 1.585 ;
        RECT 73.53 1.415 73.7 1.585 ;
        RECT 73.99 1.415 74.16 1.585 ;
        RECT 74.45 1.415 74.62 1.585 ;
        RECT 74.655 2.775 74.825 2.945 ;
        RECT 74.91 1.415 75.08 1.585 ;
        RECT 76.525 8.605 76.695 8.775 ;
        RECT 76.525 0.105 76.695 0.275 ;
        RECT 77.205 8.605 77.375 8.775 ;
        RECT 77.205 0.105 77.375 0.275 ;
        RECT 77.885 8.605 78.055 8.775 ;
        RECT 77.885 0.105 78.055 0.275 ;
        RECT 78.565 8.605 78.735 8.775 ;
        RECT 78.565 0.105 78.735 0.275 ;
        RECT 79.265 8.61 79.435 8.78 ;
        RECT 79.265 0.1 79.435 0.27 ;
        RECT 80.255 8.61 80.425 8.78 ;
        RECT 80.255 0.1 80.425 0.27 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 72.13 7.055 72.5 7.425 ;
      RECT 72.13 7.09 74.115 7.39 ;
      RECT 73.815 2.28 74.115 7.39 ;
      RECT 70.815 2.015 71.145 2.745 ;
      RECT 69.935 2.015 70.265 2.745 ;
      RECT 73.015 2.28 74.305 2.58 ;
      RECT 73.975 1.85 74.305 2.58 ;
      RECT 69.935 2.28 72.075 2.58 ;
      RECT 71.775 1.965 72.075 2.58 ;
      RECT 73.015 1.98 73.32 2.58 ;
      RECT 71.775 1.965 73.135 2.275 ;
      RECT 70.435 3.535 70.765 3.865 ;
      RECT 69.23 3.55 70.765 3.85 ;
      RECT 69.23 2.43 69.53 3.85 ;
      RECT 68.975 2.415 69.305 2.745 ;
      RECT 55.805 7.055 56.175 7.425 ;
      RECT 55.805 7.09 57.79 7.39 ;
      RECT 57.49 2.28 57.79 7.39 ;
      RECT 54.49 2.015 54.82 2.745 ;
      RECT 53.61 2.015 53.94 2.745 ;
      RECT 56.69 2.28 57.98 2.58 ;
      RECT 57.65 1.85 57.98 2.58 ;
      RECT 53.61 2.28 55.75 2.58 ;
      RECT 55.45 1.965 55.75 2.58 ;
      RECT 56.69 1.98 56.995 2.58 ;
      RECT 55.45 1.965 56.81 2.275 ;
      RECT 54.11 3.535 54.44 3.865 ;
      RECT 52.905 3.55 54.44 3.85 ;
      RECT 52.905 2.43 53.205 3.85 ;
      RECT 52.65 2.415 52.98 2.745 ;
      RECT 39.48 7.055 39.85 7.425 ;
      RECT 39.48 7.09 41.465 7.39 ;
      RECT 41.165 2.28 41.465 7.39 ;
      RECT 38.165 2.015 38.495 2.745 ;
      RECT 37.285 2.015 37.615 2.745 ;
      RECT 40.365 2.28 41.655 2.58 ;
      RECT 41.325 1.85 41.655 2.58 ;
      RECT 37.285 2.28 39.425 2.58 ;
      RECT 39.125 1.965 39.425 2.58 ;
      RECT 40.365 1.98 40.67 2.58 ;
      RECT 39.125 1.965 40.485 2.275 ;
      RECT 37.785 3.535 38.115 3.865 ;
      RECT 36.58 3.55 38.115 3.85 ;
      RECT 36.58 2.43 36.88 3.85 ;
      RECT 36.325 2.415 36.655 2.745 ;
      RECT 23.155 7.055 23.525 7.425 ;
      RECT 23.155 7.09 25.14 7.39 ;
      RECT 24.84 2.28 25.14 7.39 ;
      RECT 21.84 2.015 22.17 2.745 ;
      RECT 20.96 2.015 21.29 2.745 ;
      RECT 24.04 2.28 25.33 2.58 ;
      RECT 25 1.85 25.33 2.58 ;
      RECT 20.96 2.28 23.1 2.58 ;
      RECT 22.8 1.965 23.1 2.58 ;
      RECT 24.04 1.98 24.345 2.58 ;
      RECT 22.8 1.965 24.16 2.275 ;
      RECT 21.46 3.535 21.79 3.865 ;
      RECT 20.255 3.55 21.79 3.85 ;
      RECT 20.255 2.43 20.555 3.85 ;
      RECT 20 2.415 20.33 2.745 ;
      RECT 6.83 7.055 7.2 7.425 ;
      RECT 6.83 7.09 8.815 7.39 ;
      RECT 8.515 2.28 8.815 7.39 ;
      RECT 5.515 2.015 5.845 2.745 ;
      RECT 4.635 2.015 4.965 2.745 ;
      RECT 7.715 2.28 9.005 2.58 ;
      RECT 8.675 1.85 9.005 2.58 ;
      RECT 4.635 2.28 6.775 2.58 ;
      RECT 6.475 1.965 6.775 2.58 ;
      RECT 7.715 1.98 8.02 2.58 ;
      RECT 6.475 1.965 7.835 2.275 ;
      RECT 5.135 3.535 5.465 3.865 ;
      RECT 3.93 3.55 5.465 3.85 ;
      RECT 3.93 2.43 4.23 3.85 ;
      RECT 3.675 2.415 4.005 2.745 ;
      RECT 72.375 2.575 72.705 3.305 ;
      RECT 68.255 2.415 68.585 3.145 ;
      RECT 67.255 1.855 67.585 2.585 ;
      RECT 65.815 2.575 66.145 3.305 ;
      RECT 56.05 2.575 56.38 3.305 ;
      RECT 51.93 2.415 52.26 3.145 ;
      RECT 50.93 1.855 51.26 2.585 ;
      RECT 49.49 2.575 49.82 3.305 ;
      RECT 39.725 2.575 40.055 3.305 ;
      RECT 35.605 2.415 35.935 3.145 ;
      RECT 34.605 1.855 34.935 2.585 ;
      RECT 33.165 2.575 33.495 3.305 ;
      RECT 23.4 2.575 23.73 3.305 ;
      RECT 19.28 2.415 19.61 3.145 ;
      RECT 18.28 1.855 18.61 2.585 ;
      RECT 16.84 2.575 17.17 3.305 ;
      RECT 7.075 2.575 7.405 3.305 ;
      RECT 2.955 2.415 3.285 3.145 ;
      RECT 1.955 1.855 2.285 2.585 ;
      RECT 0.515 2.575 0.845 3.305 ;
    LAYER via2 ;
      RECT 74.04 2.315 74.24 2.515 ;
      RECT 72.44 3.04 72.64 3.24 ;
      RECT 72.215 7.14 72.415 7.34 ;
      RECT 70.88 2.48 71.08 2.68 ;
      RECT 70.5 3.6 70.7 3.8 ;
      RECT 70 2.48 70.2 2.68 ;
      RECT 69.04 2.48 69.24 2.68 ;
      RECT 68.32 2.48 68.52 2.68 ;
      RECT 67.32 1.92 67.52 2.12 ;
      RECT 65.88 3.04 66.08 3.24 ;
      RECT 57.715 2.315 57.915 2.515 ;
      RECT 56.115 3.04 56.315 3.24 ;
      RECT 55.89 7.14 56.09 7.34 ;
      RECT 54.555 2.48 54.755 2.68 ;
      RECT 54.175 3.6 54.375 3.8 ;
      RECT 53.675 2.48 53.875 2.68 ;
      RECT 52.715 2.48 52.915 2.68 ;
      RECT 51.995 2.48 52.195 2.68 ;
      RECT 50.995 1.92 51.195 2.12 ;
      RECT 49.555 3.04 49.755 3.24 ;
      RECT 41.39 2.315 41.59 2.515 ;
      RECT 39.79 3.04 39.99 3.24 ;
      RECT 39.565 7.14 39.765 7.34 ;
      RECT 38.23 2.48 38.43 2.68 ;
      RECT 37.85 3.6 38.05 3.8 ;
      RECT 37.35 2.48 37.55 2.68 ;
      RECT 36.39 2.48 36.59 2.68 ;
      RECT 35.67 2.48 35.87 2.68 ;
      RECT 34.67 1.92 34.87 2.12 ;
      RECT 33.23 3.04 33.43 3.24 ;
      RECT 25.065 2.315 25.265 2.515 ;
      RECT 23.465 3.04 23.665 3.24 ;
      RECT 23.24 7.14 23.44 7.34 ;
      RECT 21.905 2.48 22.105 2.68 ;
      RECT 21.525 3.6 21.725 3.8 ;
      RECT 21.025 2.48 21.225 2.68 ;
      RECT 20.065 2.48 20.265 2.68 ;
      RECT 19.345 2.48 19.545 2.68 ;
      RECT 18.345 1.92 18.545 2.12 ;
      RECT 16.905 3.04 17.105 3.24 ;
      RECT 8.74 2.315 8.94 2.515 ;
      RECT 7.14 3.04 7.34 3.24 ;
      RECT 6.915 7.14 7.115 7.34 ;
      RECT 5.58 2.48 5.78 2.68 ;
      RECT 5.2 3.6 5.4 3.8 ;
      RECT 4.7 2.48 4.9 2.68 ;
      RECT 3.74 2.48 3.94 2.68 ;
      RECT 3.02 2.48 3.22 2.68 ;
      RECT 2.02 1.92 2.22 2.12 ;
      RECT 0.58 3.04 0.78 3.24 ;
    LAYER met2 ;
      RECT -2.045 8.4 80.78 8.57 ;
      RECT 80.61 7.275 80.78 8.57 ;
      RECT -2.045 6.255 -1.875 8.57 ;
      RECT 80.58 7.275 80.93 7.625 ;
      RECT -2.105 6.255 -1.815 6.605 ;
      RECT 77.42 6.22 77.74 6.545 ;
      RECT 77.45 5.695 77.62 6.545 ;
      RECT 77.45 5.695 77.625 6.045 ;
      RECT 77.45 5.695 78.425 5.87 ;
      RECT 78.25 1.965 78.425 5.87 ;
      RECT 78.195 1.965 78.545 2.315 ;
      RECT 78.22 6.655 78.545 6.98 ;
      RECT 77.105 6.745 78.545 6.915 ;
      RECT 77.105 2.395 77.265 6.915 ;
      RECT 77.42 2.365 77.74 2.685 ;
      RECT 77.105 2.395 77.74 2.565 ;
      RECT 67.28 1.835 67.56 2.205 ;
      RECT 67.315 1.29 67.485 2.205 ;
      RECT 75.89 1.29 76.06 1.815 ;
      RECT 75.8 1.46 76.14 1.81 ;
      RECT 67.315 1.29 76.06 1.46 ;
      RECT 72.52 2.395 72.8 2.765 ;
      RECT 71.45 2.42 71.71 2.74 ;
      RECT 74 2.23 74.28 2.6 ;
      RECT 74.61 2.14 74.87 2.46 ;
      RECT 71.51 1.58 71.65 2.74 ;
      RECT 72.59 1.58 72.73 2.765 ;
      RECT 73.71 2.23 74.87 2.37 ;
      RECT 73.71 1.58 73.85 2.37 ;
      RECT 71.51 1.58 73.85 1.72 ;
      RECT 71.54 3.72 73.715 3.885 ;
      RECT 73.57 2.6 73.715 3.885 ;
      RECT 70.46 3.515 70.74 3.885 ;
      RECT 70.46 3.63 71.68 3.77 ;
      RECT 73.29 2.6 73.715 2.74 ;
      RECT 73.29 2.42 73.55 2.74 ;
      RECT 66.63 4 70.29 4.14 ;
      RECT 70.15 3.185 70.29 4.14 ;
      RECT 66.63 3.07 66.77 4.14 ;
      RECT 73.17 3.26 73.43 3.58 ;
      RECT 70.15 3.185 72.68 3.325 ;
      RECT 72.4 2.955 72.68 3.325 ;
      RECT 66.63 3.07 67.08 3.325 ;
      RECT 66.8 2.955 67.08 3.325 ;
      RECT 73.17 3.07 73.37 3.58 ;
      RECT 72.4 3.07 73.37 3.21 ;
      RECT 72.97 1.86 73.11 3.21 ;
      RECT 72.91 1.86 73.17 2.18 ;
      RECT 64.23 6.655 64.58 7.005 ;
      RECT 72.785 6.61 73.135 6.96 ;
      RECT 64.23 6.685 73.135 6.885 ;
      RECT 66.81 2.42 67.07 2.74 ;
      RECT 66.81 2.51 67.85 2.65 ;
      RECT 67.71 1.72 67.85 2.65 ;
      RECT 70.47 1.86 70.73 2.18 ;
      RECT 67.71 1.72 70.67 1.86 ;
      RECT 69.85 2.7 70.11 3.02 ;
      RECT 69.85 2.7 70.17 2.93 ;
      RECT 69.96 2.395 70.24 2.765 ;
      RECT 69.55 3.26 69.87 3.58 ;
      RECT 69.55 2.14 69.69 3.58 ;
      RECT 69.49 2.14 69.75 2.46 ;
      RECT 67.05 3.54 67.31 3.86 ;
      RECT 67.05 3.63 68.73 3.77 ;
      RECT 68.59 3.35 68.73 3.77 ;
      RECT 68.59 3.35 69.03 3.58 ;
      RECT 68.77 3.26 69.03 3.58 ;
      RECT 68.09 2.42 68.49 2.93 ;
      RECT 68.28 2.395 68.56 2.765 ;
      RECT 68.03 2.42 68.56 2.74 ;
      RECT 61.095 6.22 61.415 6.545 ;
      RECT 61.125 5.695 61.295 6.545 ;
      RECT 61.125 5.695 61.3 6.045 ;
      RECT 61.125 5.695 62.1 5.87 ;
      RECT 61.925 1.965 62.1 5.87 ;
      RECT 61.87 1.965 62.22 2.315 ;
      RECT 61.895 6.655 62.22 6.98 ;
      RECT 60.78 6.745 62.22 6.915 ;
      RECT 60.78 2.395 60.94 6.915 ;
      RECT 61.095 2.365 61.415 2.685 ;
      RECT 60.78 2.395 61.415 2.565 ;
      RECT 50.955 1.835 51.235 2.205 ;
      RECT 50.99 1.29 51.16 2.205 ;
      RECT 59.565 1.29 59.735 1.815 ;
      RECT 59.475 1.46 59.815 1.81 ;
      RECT 50.99 1.29 59.735 1.46 ;
      RECT 56.195 2.395 56.475 2.765 ;
      RECT 55.125 2.42 55.385 2.74 ;
      RECT 57.675 2.23 57.955 2.6 ;
      RECT 58.285 2.14 58.545 2.46 ;
      RECT 55.185 1.58 55.325 2.74 ;
      RECT 56.265 1.58 56.405 2.765 ;
      RECT 57.385 2.23 58.545 2.37 ;
      RECT 57.385 1.58 57.525 2.37 ;
      RECT 55.185 1.58 57.525 1.72 ;
      RECT 55.215 3.72 57.39 3.885 ;
      RECT 57.245 2.6 57.39 3.885 ;
      RECT 54.135 3.515 54.415 3.885 ;
      RECT 54.135 3.63 55.355 3.77 ;
      RECT 56.965 2.6 57.39 2.74 ;
      RECT 56.965 2.42 57.225 2.74 ;
      RECT 50.305 4 53.965 4.14 ;
      RECT 53.825 3.185 53.965 4.14 ;
      RECT 50.305 3.07 50.445 4.14 ;
      RECT 56.845 3.26 57.105 3.58 ;
      RECT 53.825 3.185 56.355 3.325 ;
      RECT 56.075 2.955 56.355 3.325 ;
      RECT 50.305 3.07 50.755 3.325 ;
      RECT 50.475 2.955 50.755 3.325 ;
      RECT 56.845 3.07 57.045 3.58 ;
      RECT 56.075 3.07 57.045 3.21 ;
      RECT 56.645 1.86 56.785 3.21 ;
      RECT 56.585 1.86 56.845 2.18 ;
      RECT 47.905 6.655 48.255 7.005 ;
      RECT 56.455 6.61 56.805 6.96 ;
      RECT 47.905 6.685 56.805 6.885 ;
      RECT 50.485 2.42 50.745 2.74 ;
      RECT 50.485 2.51 51.525 2.65 ;
      RECT 51.385 1.72 51.525 2.65 ;
      RECT 54.145 1.86 54.405 2.18 ;
      RECT 51.385 1.72 54.345 1.86 ;
      RECT 53.525 2.7 53.785 3.02 ;
      RECT 53.525 2.7 53.845 2.93 ;
      RECT 53.635 2.395 53.915 2.765 ;
      RECT 53.225 3.26 53.545 3.58 ;
      RECT 53.225 2.14 53.365 3.58 ;
      RECT 53.165 2.14 53.425 2.46 ;
      RECT 50.725 3.54 50.985 3.86 ;
      RECT 50.725 3.63 52.405 3.77 ;
      RECT 52.265 3.35 52.405 3.77 ;
      RECT 52.265 3.35 52.705 3.58 ;
      RECT 52.445 3.26 52.705 3.58 ;
      RECT 51.765 2.42 52.165 2.93 ;
      RECT 51.955 2.395 52.235 2.765 ;
      RECT 51.705 2.42 52.235 2.74 ;
      RECT 44.77 6.22 45.09 6.545 ;
      RECT 44.8 5.695 44.97 6.545 ;
      RECT 44.8 5.695 44.975 6.045 ;
      RECT 44.8 5.695 45.775 5.87 ;
      RECT 45.6 1.965 45.775 5.87 ;
      RECT 45.545 1.965 45.895 2.315 ;
      RECT 45.57 6.655 45.895 6.98 ;
      RECT 44.455 6.745 45.895 6.915 ;
      RECT 44.455 2.395 44.615 6.915 ;
      RECT 44.77 2.365 45.09 2.685 ;
      RECT 44.455 2.395 45.09 2.565 ;
      RECT 34.63 1.835 34.91 2.205 ;
      RECT 34.665 1.29 34.835 2.205 ;
      RECT 43.24 1.29 43.41 1.815 ;
      RECT 43.15 1.46 43.49 1.81 ;
      RECT 34.665 1.29 43.41 1.46 ;
      RECT 39.87 2.395 40.15 2.765 ;
      RECT 38.8 2.42 39.06 2.74 ;
      RECT 41.35 2.23 41.63 2.6 ;
      RECT 41.96 2.14 42.22 2.46 ;
      RECT 38.86 1.58 39 2.74 ;
      RECT 39.94 1.58 40.08 2.765 ;
      RECT 41.06 2.23 42.22 2.37 ;
      RECT 41.06 1.58 41.2 2.37 ;
      RECT 38.86 1.58 41.2 1.72 ;
      RECT 38.89 3.72 41.065 3.885 ;
      RECT 40.92 2.6 41.065 3.885 ;
      RECT 37.81 3.515 38.09 3.885 ;
      RECT 37.81 3.63 39.03 3.77 ;
      RECT 40.64 2.6 41.065 2.74 ;
      RECT 40.64 2.42 40.9 2.74 ;
      RECT 33.98 4 37.64 4.14 ;
      RECT 37.5 3.185 37.64 4.14 ;
      RECT 33.98 3.07 34.12 4.14 ;
      RECT 40.52 3.26 40.78 3.58 ;
      RECT 37.5 3.185 40.03 3.325 ;
      RECT 39.75 2.955 40.03 3.325 ;
      RECT 33.98 3.07 34.43 3.325 ;
      RECT 34.15 2.955 34.43 3.325 ;
      RECT 40.52 3.07 40.72 3.58 ;
      RECT 39.75 3.07 40.72 3.21 ;
      RECT 40.32 1.86 40.46 3.21 ;
      RECT 40.26 1.86 40.52 2.18 ;
      RECT 31.625 6.66 31.975 7.01 ;
      RECT 40.13 6.615 40.48 6.965 ;
      RECT 31.625 6.69 40.48 6.89 ;
      RECT 34.16 2.42 34.42 2.74 ;
      RECT 34.16 2.51 35.2 2.65 ;
      RECT 35.06 1.72 35.2 2.65 ;
      RECT 37.82 1.86 38.08 2.18 ;
      RECT 35.06 1.72 38.02 1.86 ;
      RECT 37.2 2.7 37.46 3.02 ;
      RECT 37.2 2.7 37.52 2.93 ;
      RECT 37.31 2.395 37.59 2.765 ;
      RECT 36.9 3.26 37.22 3.58 ;
      RECT 36.9 2.14 37.04 3.58 ;
      RECT 36.84 2.14 37.1 2.46 ;
      RECT 34.4 3.54 34.66 3.86 ;
      RECT 34.4 3.63 36.08 3.77 ;
      RECT 35.94 3.35 36.08 3.77 ;
      RECT 35.94 3.35 36.38 3.58 ;
      RECT 36.12 3.26 36.38 3.58 ;
      RECT 35.44 2.42 35.84 2.93 ;
      RECT 35.63 2.395 35.91 2.765 ;
      RECT 35.38 2.42 35.91 2.74 ;
      RECT 28.445 6.22 28.765 6.545 ;
      RECT 28.475 5.695 28.645 6.545 ;
      RECT 28.475 5.695 28.65 6.045 ;
      RECT 28.475 5.695 29.45 5.87 ;
      RECT 29.275 1.965 29.45 5.87 ;
      RECT 29.22 1.965 29.57 2.315 ;
      RECT 29.245 6.655 29.57 6.98 ;
      RECT 28.13 6.745 29.57 6.915 ;
      RECT 28.13 2.395 28.29 6.915 ;
      RECT 28.445 2.365 28.765 2.685 ;
      RECT 28.13 2.395 28.765 2.565 ;
      RECT 18.305 1.835 18.585 2.205 ;
      RECT 18.34 1.29 18.51 2.205 ;
      RECT 26.915 1.29 27.085 1.815 ;
      RECT 26.825 1.46 27.165 1.81 ;
      RECT 18.34 1.29 27.085 1.46 ;
      RECT 23.545 2.395 23.825 2.765 ;
      RECT 22.475 2.42 22.735 2.74 ;
      RECT 25.025 2.23 25.305 2.6 ;
      RECT 25.635 2.14 25.895 2.46 ;
      RECT 22.535 1.58 22.675 2.74 ;
      RECT 23.615 1.58 23.755 2.765 ;
      RECT 24.735 2.23 25.895 2.37 ;
      RECT 24.735 1.58 24.875 2.37 ;
      RECT 22.535 1.58 24.875 1.72 ;
      RECT 22.565 3.72 24.74 3.885 ;
      RECT 24.595 2.6 24.74 3.885 ;
      RECT 21.485 3.515 21.765 3.885 ;
      RECT 21.485 3.63 22.705 3.77 ;
      RECT 24.315 2.6 24.74 2.74 ;
      RECT 24.315 2.42 24.575 2.74 ;
      RECT 17.655 4 21.315 4.14 ;
      RECT 21.175 3.185 21.315 4.14 ;
      RECT 17.655 3.07 17.795 4.14 ;
      RECT 24.195 3.26 24.455 3.58 ;
      RECT 21.175 3.185 23.705 3.325 ;
      RECT 23.425 2.955 23.705 3.325 ;
      RECT 17.655 3.07 18.105 3.325 ;
      RECT 17.825 2.955 18.105 3.325 ;
      RECT 24.195 3.07 24.395 3.58 ;
      RECT 23.425 3.07 24.395 3.21 ;
      RECT 23.995 1.86 24.135 3.21 ;
      RECT 23.935 1.86 24.195 2.18 ;
      RECT 15.3 6.655 15.65 7.005 ;
      RECT 23.805 6.61 24.155 6.96 ;
      RECT 15.3 6.685 24.155 6.885 ;
      RECT 17.835 2.42 18.095 2.74 ;
      RECT 17.835 2.51 18.875 2.65 ;
      RECT 18.735 1.72 18.875 2.65 ;
      RECT 21.495 1.86 21.755 2.18 ;
      RECT 18.735 1.72 21.695 1.86 ;
      RECT 20.875 2.7 21.135 3.02 ;
      RECT 20.875 2.7 21.195 2.93 ;
      RECT 20.985 2.395 21.265 2.765 ;
      RECT 20.575 3.26 20.895 3.58 ;
      RECT 20.575 2.14 20.715 3.58 ;
      RECT 20.515 2.14 20.775 2.46 ;
      RECT 18.075 3.54 18.335 3.86 ;
      RECT 18.075 3.63 19.755 3.77 ;
      RECT 19.615 3.35 19.755 3.77 ;
      RECT 19.615 3.35 20.055 3.58 ;
      RECT 19.795 3.26 20.055 3.58 ;
      RECT 19.115 2.42 19.515 2.93 ;
      RECT 19.305 2.395 19.585 2.765 ;
      RECT 19.055 2.42 19.585 2.74 ;
      RECT 12.12 6.22 12.44 6.545 ;
      RECT 12.15 5.695 12.32 6.545 ;
      RECT 12.15 5.695 12.325 6.045 ;
      RECT 12.15 5.695 13.125 5.87 ;
      RECT 12.95 1.965 13.125 5.87 ;
      RECT 12.895 1.965 13.245 2.315 ;
      RECT 12.92 6.655 13.245 6.98 ;
      RECT 11.805 6.745 13.245 6.915 ;
      RECT 11.805 2.395 11.965 6.915 ;
      RECT 12.12 2.365 12.44 2.685 ;
      RECT 11.805 2.395 12.44 2.565 ;
      RECT 1.98 1.835 2.26 2.205 ;
      RECT 2.015 1.29 2.185 2.205 ;
      RECT 10.59 1.29 10.76 1.815 ;
      RECT 10.5 1.46 10.84 1.81 ;
      RECT 2.015 1.29 10.76 1.46 ;
      RECT 7.22 2.395 7.5 2.765 ;
      RECT 6.15 2.42 6.41 2.74 ;
      RECT 8.7 2.23 8.98 2.6 ;
      RECT 9.31 2.14 9.57 2.46 ;
      RECT 6.21 1.58 6.35 2.74 ;
      RECT 7.29 1.58 7.43 2.765 ;
      RECT 8.41 2.23 9.57 2.37 ;
      RECT 8.41 1.58 8.55 2.37 ;
      RECT 6.21 1.58 8.55 1.72 ;
      RECT -1.73 6.995 -1.44 7.345 ;
      RECT -1.73 7.05 -0.445 7.225 ;
      RECT -0.62 6.685 -0.445 7.225 ;
      RECT 8.315 6.605 8.665 6.955 ;
      RECT -0.62 6.685 8.665 6.86 ;
      RECT 6.24 3.72 8.415 3.885 ;
      RECT 8.27 2.6 8.415 3.885 ;
      RECT 5.16 3.515 5.44 3.885 ;
      RECT 5.16 3.63 6.38 3.77 ;
      RECT 7.99 2.6 8.415 2.74 ;
      RECT 7.99 2.42 8.25 2.74 ;
      RECT 1.33 4 4.99 4.14 ;
      RECT 4.85 3.185 4.99 4.14 ;
      RECT 1.33 3.07 1.47 4.14 ;
      RECT 7.87 3.26 8.13 3.58 ;
      RECT 4.85 3.185 7.38 3.325 ;
      RECT 7.1 2.955 7.38 3.325 ;
      RECT 1.33 3.07 1.78 3.325 ;
      RECT 1.5 2.955 1.78 3.325 ;
      RECT 7.87 3.07 8.07 3.58 ;
      RECT 7.1 3.07 8.07 3.21 ;
      RECT 7.67 1.86 7.81 3.21 ;
      RECT 7.61 1.86 7.87 2.18 ;
      RECT 1.51 2.42 1.77 2.74 ;
      RECT 1.51 2.51 2.55 2.65 ;
      RECT 2.41 1.72 2.55 2.65 ;
      RECT 5.17 1.86 5.43 2.18 ;
      RECT 2.41 1.72 5.37 1.86 ;
      RECT 4.55 2.7 4.81 3.02 ;
      RECT 4.55 2.7 4.87 2.93 ;
      RECT 4.66 2.395 4.94 2.765 ;
      RECT 4.25 3.26 4.57 3.58 ;
      RECT 4.25 2.14 4.39 3.58 ;
      RECT 4.19 2.14 4.45 2.46 ;
      RECT 1.75 3.54 2.01 3.86 ;
      RECT 1.75 3.63 3.43 3.77 ;
      RECT 3.29 3.35 3.43 3.77 ;
      RECT 3.29 3.35 3.73 3.58 ;
      RECT 3.47 3.26 3.73 3.58 ;
      RECT 2.79 2.42 3.19 2.93 ;
      RECT 2.98 2.395 3.26 2.765 ;
      RECT 2.73 2.42 3.26 2.74 ;
      RECT 72.13 7.055 72.5 7.425 ;
      RECT 70.84 2.395 71.12 2.765 ;
      RECT 69 2.395 69.28 2.765 ;
      RECT 65.84 2.955 66.12 3.325 ;
      RECT 55.805 7.055 56.175 7.425 ;
      RECT 54.515 2.395 54.795 2.765 ;
      RECT 52.675 2.395 52.955 2.765 ;
      RECT 49.515 2.955 49.795 3.325 ;
      RECT 39.48 7.055 39.85 7.425 ;
      RECT 38.19 2.395 38.47 2.765 ;
      RECT 36.35 2.395 36.63 2.765 ;
      RECT 33.19 2.955 33.47 3.325 ;
      RECT 23.155 7.055 23.525 7.425 ;
      RECT 21.865 2.395 22.145 2.765 ;
      RECT 20.025 2.395 20.305 2.765 ;
      RECT 16.865 2.955 17.145 3.325 ;
      RECT 6.83 7.055 7.2 7.425 ;
      RECT 5.54 2.395 5.82 2.765 ;
      RECT 3.7 2.395 3.98 2.765 ;
      RECT 0.54 2.955 0.82 3.325 ;
    LAYER via1 ;
      RECT 80.68 7.375 80.83 7.525 ;
      RECT 78.31 6.74 78.46 6.89 ;
      RECT 78.295 2.065 78.445 2.215 ;
      RECT 77.505 2.45 77.655 2.6 ;
      RECT 77.505 6.325 77.655 6.475 ;
      RECT 75.9 1.56 76.05 1.71 ;
      RECT 74.665 2.225 74.815 2.375 ;
      RECT 73.345 2.505 73.495 2.655 ;
      RECT 73.225 3.345 73.375 3.495 ;
      RECT 72.965 1.945 73.115 2.095 ;
      RECT 72.885 6.71 73.035 6.86 ;
      RECT 72.24 7.165 72.39 7.315 ;
      RECT 71.505 2.505 71.655 2.655 ;
      RECT 70.905 2.505 71.055 2.655 ;
      RECT 70.525 1.945 70.675 2.095 ;
      RECT 69.905 2.785 70.055 2.935 ;
      RECT 69.665 3.345 69.815 3.495 ;
      RECT 69.545 2.225 69.695 2.375 ;
      RECT 69.065 2.505 69.215 2.655 ;
      RECT 68.825 3.345 68.975 3.495 ;
      RECT 68.085 2.505 68.235 2.655 ;
      RECT 67.345 1.945 67.495 2.095 ;
      RECT 67.105 3.625 67.255 3.775 ;
      RECT 66.865 2.505 67.015 2.655 ;
      RECT 66.865 3.065 67.015 3.215 ;
      RECT 65.905 3.065 66.055 3.215 ;
      RECT 64.33 6.755 64.48 6.905 ;
      RECT 61.985 6.74 62.135 6.89 ;
      RECT 61.97 2.065 62.12 2.215 ;
      RECT 61.18 2.45 61.33 2.6 ;
      RECT 61.18 6.325 61.33 6.475 ;
      RECT 59.575 1.56 59.725 1.71 ;
      RECT 58.34 2.225 58.49 2.375 ;
      RECT 57.02 2.505 57.17 2.655 ;
      RECT 56.9 3.345 57.05 3.495 ;
      RECT 56.64 1.945 56.79 2.095 ;
      RECT 56.555 6.71 56.705 6.86 ;
      RECT 55.915 7.165 56.065 7.315 ;
      RECT 55.18 2.505 55.33 2.655 ;
      RECT 54.58 2.505 54.73 2.655 ;
      RECT 54.2 1.945 54.35 2.095 ;
      RECT 53.58 2.785 53.73 2.935 ;
      RECT 53.34 3.345 53.49 3.495 ;
      RECT 53.22 2.225 53.37 2.375 ;
      RECT 52.74 2.505 52.89 2.655 ;
      RECT 52.5 3.345 52.65 3.495 ;
      RECT 51.76 2.505 51.91 2.655 ;
      RECT 51.02 1.945 51.17 2.095 ;
      RECT 50.78 3.625 50.93 3.775 ;
      RECT 50.54 2.505 50.69 2.655 ;
      RECT 50.54 3.065 50.69 3.215 ;
      RECT 49.58 3.065 49.73 3.215 ;
      RECT 48.005 6.755 48.155 6.905 ;
      RECT 45.66 6.74 45.81 6.89 ;
      RECT 45.645 2.065 45.795 2.215 ;
      RECT 44.855 2.45 45.005 2.6 ;
      RECT 44.855 6.325 45.005 6.475 ;
      RECT 43.25 1.56 43.4 1.71 ;
      RECT 42.015 2.225 42.165 2.375 ;
      RECT 40.695 2.505 40.845 2.655 ;
      RECT 40.575 3.345 40.725 3.495 ;
      RECT 40.315 1.945 40.465 2.095 ;
      RECT 40.23 6.715 40.38 6.865 ;
      RECT 39.59 7.165 39.74 7.315 ;
      RECT 38.855 2.505 39.005 2.655 ;
      RECT 38.255 2.505 38.405 2.655 ;
      RECT 37.875 1.945 38.025 2.095 ;
      RECT 37.255 2.785 37.405 2.935 ;
      RECT 37.015 3.345 37.165 3.495 ;
      RECT 36.895 2.225 37.045 2.375 ;
      RECT 36.415 2.505 36.565 2.655 ;
      RECT 36.175 3.345 36.325 3.495 ;
      RECT 35.435 2.505 35.585 2.655 ;
      RECT 34.695 1.945 34.845 2.095 ;
      RECT 34.455 3.625 34.605 3.775 ;
      RECT 34.215 2.505 34.365 2.655 ;
      RECT 34.215 3.065 34.365 3.215 ;
      RECT 33.255 3.065 33.405 3.215 ;
      RECT 31.725 6.76 31.875 6.91 ;
      RECT 29.335 6.74 29.485 6.89 ;
      RECT 29.32 2.065 29.47 2.215 ;
      RECT 28.53 2.45 28.68 2.6 ;
      RECT 28.53 6.325 28.68 6.475 ;
      RECT 26.925 1.56 27.075 1.71 ;
      RECT 25.69 2.225 25.84 2.375 ;
      RECT 24.37 2.505 24.52 2.655 ;
      RECT 24.25 3.345 24.4 3.495 ;
      RECT 23.99 1.945 24.14 2.095 ;
      RECT 23.905 6.71 24.055 6.86 ;
      RECT 23.265 7.165 23.415 7.315 ;
      RECT 22.53 2.505 22.68 2.655 ;
      RECT 21.93 2.505 22.08 2.655 ;
      RECT 21.55 1.945 21.7 2.095 ;
      RECT 20.93 2.785 21.08 2.935 ;
      RECT 20.69 3.345 20.84 3.495 ;
      RECT 20.57 2.225 20.72 2.375 ;
      RECT 20.09 2.505 20.24 2.655 ;
      RECT 19.85 3.345 20 3.495 ;
      RECT 19.11 2.505 19.26 2.655 ;
      RECT 18.37 1.945 18.52 2.095 ;
      RECT 18.13 3.625 18.28 3.775 ;
      RECT 17.89 2.505 18.04 2.655 ;
      RECT 17.89 3.065 18.04 3.215 ;
      RECT 16.93 3.065 17.08 3.215 ;
      RECT 15.4 6.755 15.55 6.905 ;
      RECT 13.01 6.74 13.16 6.89 ;
      RECT 12.995 2.065 13.145 2.215 ;
      RECT 12.205 2.45 12.355 2.6 ;
      RECT 12.205 6.325 12.355 6.475 ;
      RECT 10.6 1.56 10.75 1.71 ;
      RECT 9.365 2.225 9.515 2.375 ;
      RECT 8.415 6.705 8.565 6.855 ;
      RECT 8.045 2.505 8.195 2.655 ;
      RECT 7.925 3.345 8.075 3.495 ;
      RECT 7.665 1.945 7.815 2.095 ;
      RECT 6.94 7.165 7.09 7.315 ;
      RECT 6.205 2.505 6.355 2.655 ;
      RECT 5.605 2.505 5.755 2.655 ;
      RECT 5.225 1.945 5.375 2.095 ;
      RECT 4.605 2.785 4.755 2.935 ;
      RECT 4.365 3.345 4.515 3.495 ;
      RECT 4.245 2.225 4.395 2.375 ;
      RECT 3.765 2.505 3.915 2.655 ;
      RECT 3.525 3.345 3.675 3.495 ;
      RECT 2.785 2.505 2.935 2.655 ;
      RECT 2.045 1.945 2.195 2.095 ;
      RECT 1.805 3.625 1.955 3.775 ;
      RECT 1.565 2.505 1.715 2.655 ;
      RECT 1.565 3.065 1.715 3.215 ;
      RECT 0.605 3.065 0.755 3.215 ;
      RECT -1.66 7.095 -1.51 7.245 ;
      RECT -2.035 6.355 -1.885 6.505 ;
    LAYER met1 ;
      RECT 80.545 7.77 80.835 8 ;
      RECT 80.605 6.29 80.775 8 ;
      RECT 80.58 7.275 80.93 7.625 ;
      RECT 80.545 6.29 80.835 6.52 ;
      RECT 80.14 2.395 80.245 2.965 ;
      RECT 80.14 2.73 80.465 2.96 ;
      RECT 80.14 2.76 80.635 2.93 ;
      RECT 80.14 2.395 80.33 2.96 ;
      RECT 79.555 2.36 79.845 2.59 ;
      RECT 79.555 2.395 80.33 2.565 ;
      RECT 79.615 0.88 79.785 2.59 ;
      RECT 79.555 0.88 79.845 1.11 ;
      RECT 79.555 7.77 79.845 8 ;
      RECT 79.615 6.29 79.785 8 ;
      RECT 79.555 6.29 79.845 6.52 ;
      RECT 79.555 6.325 80.41 6.485 ;
      RECT 80.24 5.92 80.41 6.485 ;
      RECT 79.555 6.32 79.95 6.485 ;
      RECT 80.175 5.92 80.465 6.15 ;
      RECT 80.175 5.95 80.635 6.12 ;
      RECT 79.185 2.73 79.475 2.96 ;
      RECT 79.185 2.76 79.645 2.93 ;
      RECT 79.25 1.655 79.415 2.96 ;
      RECT 77.765 1.625 78.055 1.855 ;
      RECT 77.765 1.655 79.415 1.825 ;
      RECT 77.825 0.885 77.995 1.855 ;
      RECT 77.765 0.885 78.055 1.115 ;
      RECT 77.765 7.765 78.055 7.995 ;
      RECT 77.825 7.025 77.995 7.995 ;
      RECT 77.825 7.12 79.415 7.29 ;
      RECT 79.245 5.92 79.415 7.29 ;
      RECT 77.765 7.025 78.055 7.255 ;
      RECT 79.185 5.92 79.475 6.15 ;
      RECT 79.185 5.95 79.645 6.12 ;
      RECT 78.195 1.965 78.545 2.315 ;
      RECT 75.89 2.025 78.545 2.195 ;
      RECT 75.89 1.46 76.06 2.195 ;
      RECT 75.8 1.46 76.14 1.81 ;
      RECT 78.22 6.655 78.545 6.98 ;
      RECT 72.785 6.61 73.135 6.96 ;
      RECT 78.195 6.655 78.545 6.885 ;
      RECT 72.58 6.655 73.135 6.885 ;
      RECT 72.41 6.685 78.545 6.855 ;
      RECT 77.42 2.365 77.74 2.685 ;
      RECT 77.39 2.365 77.74 2.595 ;
      RECT 77.22 2.395 77.74 2.565 ;
      RECT 77.42 6.255 77.74 6.545 ;
      RECT 77.39 6.285 77.74 6.515 ;
      RECT 77.22 6.315 77.74 6.485 ;
      RECT 73.875 2.465 74.165 2.695 ;
      RECT 73.875 2.465 74.33 2.65 ;
      RECT 74.19 2.37 74.81 2.51 ;
      RECT 74.58 2.17 74.9 2.43 ;
      RECT 73.26 2.45 73.58 2.71 ;
      RECT 73.26 2.45 73.725 2.695 ;
      RECT 73.585 2.07 73.725 2.695 ;
      RECT 73.585 2.07 73.85 2.21 ;
      RECT 74.115 1.905 74.405 2.135 ;
      RECT 73.71 1.95 74.405 2.09 ;
      RECT 73.155 3.29 73.445 3.815 ;
      RECT 73.14 3.29 73.46 3.55 ;
      RECT 72.88 1.89 73.2 2.15 ;
      RECT 72.88 1.905 73.445 2.135 ;
      RECT 72.155 3.585 72.445 3.815 ;
      RECT 72.35 2.23 72.49 3.77 ;
      RECT 72.395 2.185 72.685 2.415 ;
      RECT 71.99 2.23 72.685 2.37 ;
      RECT 71.99 2.07 72.13 2.37 ;
      RECT 70.53 2.07 72.13 2.21 ;
      RECT 70.44 1.89 70.76 2.15 ;
      RECT 70.44 1.905 71.005 2.15 ;
      RECT 72.15 7.765 72.44 7.995 ;
      RECT 72.21 7.025 72.38 7.995 ;
      RECT 72.13 7.075 72.5 7.425 ;
      RECT 72.13 7.055 72.44 7.425 ;
      RECT 72.15 7.025 72.44 7.425 ;
      RECT 69.55 2.93 72.13 3.07 ;
      RECT 71.915 2.745 72.205 2.975 ;
      RECT 69.475 2.745 70.14 2.975 ;
      RECT 69.82 2.73 70.14 3.07 ;
      RECT 70.82 2.45 71.14 2.71 ;
      RECT 70.82 2.465 71.245 2.695 ;
      RECT 69.46 2.17 69.78 2.43 ;
      RECT 69.955 2.185 70.245 2.415 ;
      RECT 69.46 2.23 70.245 2.37 ;
      RECT 69.58 3.29 69.9 3.55 ;
      RECT 68.74 3.29 69.06 3.55 ;
      RECT 69.58 3.305 70.005 3.535 ;
      RECT 68.74 3.35 70.005 3.49 ;
      RECT 68.275 3.025 68.565 3.255 ;
      RECT 68.35 1.95 68.49 3.255 ;
      RECT 68 2.45 68.49 2.71 ;
      RECT 67.755 2.465 68.49 2.695 ;
      RECT 68.755 1.905 69.045 2.135 ;
      RECT 68.35 1.95 69.045 2.09 ;
      RECT 67.515 3.305 67.805 3.535 ;
      RECT 67.515 3.305 67.97 3.49 ;
      RECT 67.83 2.93 67.97 3.49 ;
      RECT 67.47 2.93 67.97 3.07 ;
      RECT 67.47 1.95 67.61 3.07 ;
      RECT 67.26 1.89 67.58 2.15 ;
      RECT 67.02 3.57 67.34 3.83 ;
      RECT 66.315 3.585 66.605 3.815 ;
      RECT 66.315 3.63 67.34 3.77 ;
      RECT 66.39 3.58 66.65 3.77 ;
      RECT 66.78 2.45 67.1 2.71 ;
      RECT 66.78 2.465 67.325 2.695 ;
      RECT 66.78 3.01 67.1 3.27 ;
      RECT 66.78 3.025 67.325 3.255 ;
      RECT 65.82 3.01 66.14 3.27 ;
      RECT 65.91 1.95 66.05 3.27 ;
      RECT 66.315 1.905 66.605 2.135 ;
      RECT 65.91 1.95 66.605 2.09 ;
      RECT 64.22 7.77 64.51 8 ;
      RECT 64.28 6.29 64.45 8 ;
      RECT 64.23 6.655 64.58 7.005 ;
      RECT 64.22 6.29 64.51 6.52 ;
      RECT 63.815 2.395 63.92 2.965 ;
      RECT 63.815 2.73 64.14 2.96 ;
      RECT 63.815 2.76 64.31 2.93 ;
      RECT 63.815 2.395 64.005 2.96 ;
      RECT 63.23 2.36 63.52 2.59 ;
      RECT 63.23 2.395 64.005 2.565 ;
      RECT 63.29 0.88 63.46 2.59 ;
      RECT 63.23 0.88 63.52 1.11 ;
      RECT 63.23 7.77 63.52 8 ;
      RECT 63.29 6.29 63.46 8 ;
      RECT 63.23 6.29 63.52 6.52 ;
      RECT 63.23 6.325 64.085 6.485 ;
      RECT 63.915 5.92 64.085 6.485 ;
      RECT 63.23 6.32 63.625 6.485 ;
      RECT 63.85 5.92 64.14 6.15 ;
      RECT 63.85 5.95 64.31 6.12 ;
      RECT 62.86 2.73 63.15 2.96 ;
      RECT 62.86 2.76 63.32 2.93 ;
      RECT 62.925 1.655 63.09 2.96 ;
      RECT 61.44 1.625 61.73 1.855 ;
      RECT 61.44 1.655 63.09 1.825 ;
      RECT 61.5 0.885 61.67 1.855 ;
      RECT 61.44 0.885 61.73 1.115 ;
      RECT 61.44 7.765 61.73 7.995 ;
      RECT 61.5 7.025 61.67 7.995 ;
      RECT 61.5 7.12 63.09 7.29 ;
      RECT 62.92 5.92 63.09 7.29 ;
      RECT 61.44 7.025 61.73 7.255 ;
      RECT 62.86 5.92 63.15 6.15 ;
      RECT 62.86 5.95 63.32 6.12 ;
      RECT 61.87 1.965 62.22 2.315 ;
      RECT 59.565 2.025 62.22 2.195 ;
      RECT 59.565 1.46 59.735 2.195 ;
      RECT 59.475 1.46 59.815 1.81 ;
      RECT 61.895 6.655 62.22 6.98 ;
      RECT 56.455 6.61 56.805 6.96 ;
      RECT 61.87 6.655 62.22 6.885 ;
      RECT 56.255 6.655 56.805 6.885 ;
      RECT 56.085 6.685 62.22 6.855 ;
      RECT 61.095 2.365 61.415 2.685 ;
      RECT 61.065 2.365 61.415 2.595 ;
      RECT 60.895 2.395 61.415 2.565 ;
      RECT 61.095 6.255 61.415 6.545 ;
      RECT 61.065 6.285 61.415 6.515 ;
      RECT 60.895 6.315 61.415 6.485 ;
      RECT 57.55 2.465 57.84 2.695 ;
      RECT 57.55 2.465 58.005 2.65 ;
      RECT 57.865 2.37 58.485 2.51 ;
      RECT 58.255 2.17 58.575 2.43 ;
      RECT 56.935 2.45 57.255 2.71 ;
      RECT 56.935 2.45 57.4 2.695 ;
      RECT 57.26 2.07 57.4 2.695 ;
      RECT 57.26 2.07 57.525 2.21 ;
      RECT 57.79 1.905 58.08 2.135 ;
      RECT 57.385 1.95 58.08 2.09 ;
      RECT 56.83 3.29 57.12 3.815 ;
      RECT 56.815 3.29 57.135 3.55 ;
      RECT 56.555 1.89 56.875 2.15 ;
      RECT 56.555 1.905 57.12 2.135 ;
      RECT 55.83 3.585 56.12 3.815 ;
      RECT 56.025 2.23 56.165 3.77 ;
      RECT 56.07 2.185 56.36 2.415 ;
      RECT 55.665 2.23 56.36 2.37 ;
      RECT 55.665 2.07 55.805 2.37 ;
      RECT 54.205 2.07 55.805 2.21 ;
      RECT 54.115 1.89 54.435 2.15 ;
      RECT 54.115 1.905 54.68 2.15 ;
      RECT 55.825 7.765 56.115 7.995 ;
      RECT 55.885 7.025 56.055 7.995 ;
      RECT 55.805 7.075 56.175 7.425 ;
      RECT 55.805 7.055 56.115 7.425 ;
      RECT 55.825 7.025 56.115 7.425 ;
      RECT 53.225 2.93 55.805 3.07 ;
      RECT 55.59 2.745 55.88 2.975 ;
      RECT 53.15 2.745 53.815 2.975 ;
      RECT 53.495 2.73 53.815 3.07 ;
      RECT 54.495 2.45 54.815 2.71 ;
      RECT 54.495 2.465 54.92 2.695 ;
      RECT 53.135 2.17 53.455 2.43 ;
      RECT 53.63 2.185 53.92 2.415 ;
      RECT 53.135 2.23 53.92 2.37 ;
      RECT 53.255 3.29 53.575 3.55 ;
      RECT 52.415 3.29 52.735 3.55 ;
      RECT 53.255 3.305 53.68 3.535 ;
      RECT 52.415 3.35 53.68 3.49 ;
      RECT 51.95 3.025 52.24 3.255 ;
      RECT 52.025 1.95 52.165 3.255 ;
      RECT 51.675 2.45 52.165 2.71 ;
      RECT 51.43 2.465 52.165 2.695 ;
      RECT 52.43 1.905 52.72 2.135 ;
      RECT 52.025 1.95 52.72 2.09 ;
      RECT 51.19 3.305 51.48 3.535 ;
      RECT 51.19 3.305 51.645 3.49 ;
      RECT 51.505 2.93 51.645 3.49 ;
      RECT 51.145 2.93 51.645 3.07 ;
      RECT 51.145 1.95 51.285 3.07 ;
      RECT 50.935 1.89 51.255 2.15 ;
      RECT 50.695 3.57 51.015 3.83 ;
      RECT 49.99 3.585 50.28 3.815 ;
      RECT 49.99 3.63 51.015 3.77 ;
      RECT 50.065 3.58 50.325 3.77 ;
      RECT 50.455 2.45 50.775 2.71 ;
      RECT 50.455 2.465 51 2.695 ;
      RECT 50.455 3.01 50.775 3.27 ;
      RECT 50.455 3.025 51 3.255 ;
      RECT 49.495 3.01 49.815 3.27 ;
      RECT 49.585 1.95 49.725 3.27 ;
      RECT 49.99 1.905 50.28 2.135 ;
      RECT 49.585 1.95 50.28 2.09 ;
      RECT 47.895 7.77 48.185 8 ;
      RECT 47.955 6.29 48.125 8 ;
      RECT 47.905 6.655 48.255 7.005 ;
      RECT 47.895 6.29 48.185 6.52 ;
      RECT 47.49 2.395 47.595 2.965 ;
      RECT 47.49 2.73 47.815 2.96 ;
      RECT 47.49 2.76 47.985 2.93 ;
      RECT 47.49 2.395 47.68 2.96 ;
      RECT 46.905 2.36 47.195 2.59 ;
      RECT 46.905 2.395 47.68 2.565 ;
      RECT 46.965 0.88 47.135 2.59 ;
      RECT 46.905 0.88 47.195 1.11 ;
      RECT 46.905 7.77 47.195 8 ;
      RECT 46.965 6.29 47.135 8 ;
      RECT 46.905 6.29 47.195 6.52 ;
      RECT 46.905 6.325 47.76 6.485 ;
      RECT 47.59 5.92 47.76 6.485 ;
      RECT 46.905 6.32 47.3 6.485 ;
      RECT 47.525 5.92 47.815 6.15 ;
      RECT 47.525 5.95 47.985 6.12 ;
      RECT 46.535 2.73 46.825 2.96 ;
      RECT 46.535 2.76 46.995 2.93 ;
      RECT 46.6 1.655 46.765 2.96 ;
      RECT 45.115 1.625 45.405 1.855 ;
      RECT 45.115 1.655 46.765 1.825 ;
      RECT 45.175 0.885 45.345 1.855 ;
      RECT 45.115 0.885 45.405 1.115 ;
      RECT 45.115 7.765 45.405 7.995 ;
      RECT 45.175 7.025 45.345 7.995 ;
      RECT 45.175 7.12 46.765 7.29 ;
      RECT 46.595 5.92 46.765 7.29 ;
      RECT 45.115 7.025 45.405 7.255 ;
      RECT 46.535 5.92 46.825 6.15 ;
      RECT 46.535 5.95 46.995 6.12 ;
      RECT 45.545 1.965 45.895 2.315 ;
      RECT 43.24 2.025 45.895 2.195 ;
      RECT 43.24 1.46 43.41 2.195 ;
      RECT 43.15 1.46 43.49 1.81 ;
      RECT 45.57 6.655 45.895 6.98 ;
      RECT 40.13 6.615 40.48 6.965 ;
      RECT 45.545 6.655 45.895 6.885 ;
      RECT 39.93 6.655 40.48 6.885 ;
      RECT 39.76 6.685 45.895 6.855 ;
      RECT 44.77 2.365 45.09 2.685 ;
      RECT 44.74 2.365 45.09 2.595 ;
      RECT 44.57 2.395 45.09 2.565 ;
      RECT 44.77 6.255 45.09 6.545 ;
      RECT 44.74 6.285 45.09 6.515 ;
      RECT 44.57 6.315 45.09 6.485 ;
      RECT 41.225 2.465 41.515 2.695 ;
      RECT 41.225 2.465 41.68 2.65 ;
      RECT 41.54 2.37 42.16 2.51 ;
      RECT 41.93 2.17 42.25 2.43 ;
      RECT 40.61 2.45 40.93 2.71 ;
      RECT 40.61 2.45 41.075 2.695 ;
      RECT 40.935 2.07 41.075 2.695 ;
      RECT 40.935 2.07 41.2 2.21 ;
      RECT 41.465 1.905 41.755 2.135 ;
      RECT 41.06 1.95 41.755 2.09 ;
      RECT 40.505 3.29 40.795 3.815 ;
      RECT 40.49 3.29 40.81 3.55 ;
      RECT 40.23 1.89 40.55 2.15 ;
      RECT 40.23 1.905 40.795 2.135 ;
      RECT 39.505 3.585 39.795 3.815 ;
      RECT 39.7 2.23 39.84 3.77 ;
      RECT 39.745 2.185 40.035 2.415 ;
      RECT 39.34 2.23 40.035 2.37 ;
      RECT 39.34 2.07 39.48 2.37 ;
      RECT 37.88 2.07 39.48 2.21 ;
      RECT 37.79 1.89 38.11 2.15 ;
      RECT 37.79 1.905 38.355 2.15 ;
      RECT 39.5 7.765 39.79 7.995 ;
      RECT 39.56 7.025 39.73 7.995 ;
      RECT 39.48 7.075 39.85 7.425 ;
      RECT 39.48 7.055 39.79 7.425 ;
      RECT 39.5 7.025 39.79 7.425 ;
      RECT 36.9 2.93 39.48 3.07 ;
      RECT 39.265 2.745 39.555 2.975 ;
      RECT 36.825 2.745 37.49 2.975 ;
      RECT 37.17 2.73 37.49 3.07 ;
      RECT 38.17 2.45 38.49 2.71 ;
      RECT 38.17 2.465 38.595 2.695 ;
      RECT 36.81 2.17 37.13 2.43 ;
      RECT 37.305 2.185 37.595 2.415 ;
      RECT 36.81 2.23 37.595 2.37 ;
      RECT 36.93 3.29 37.25 3.55 ;
      RECT 36.09 3.29 36.41 3.55 ;
      RECT 36.93 3.305 37.355 3.535 ;
      RECT 36.09 3.35 37.355 3.49 ;
      RECT 35.625 3.025 35.915 3.255 ;
      RECT 35.7 1.95 35.84 3.255 ;
      RECT 35.35 2.45 35.84 2.71 ;
      RECT 35.105 2.465 35.84 2.695 ;
      RECT 36.105 1.905 36.395 2.135 ;
      RECT 35.7 1.95 36.395 2.09 ;
      RECT 34.865 3.305 35.155 3.535 ;
      RECT 34.865 3.305 35.32 3.49 ;
      RECT 35.18 2.93 35.32 3.49 ;
      RECT 34.82 2.93 35.32 3.07 ;
      RECT 34.82 1.95 34.96 3.07 ;
      RECT 34.61 1.89 34.93 2.15 ;
      RECT 34.37 3.57 34.69 3.83 ;
      RECT 33.665 3.585 33.955 3.815 ;
      RECT 33.665 3.63 34.69 3.77 ;
      RECT 33.74 3.58 34 3.77 ;
      RECT 34.13 2.45 34.45 2.71 ;
      RECT 34.13 2.465 34.675 2.695 ;
      RECT 34.13 3.01 34.45 3.27 ;
      RECT 34.13 3.025 34.675 3.255 ;
      RECT 33.17 3.01 33.49 3.27 ;
      RECT 33.26 1.95 33.4 3.27 ;
      RECT 33.665 1.905 33.955 2.135 ;
      RECT 33.26 1.95 33.955 2.09 ;
      RECT 31.57 7.77 31.86 8 ;
      RECT 31.63 6.29 31.8 8 ;
      RECT 31.62 6.66 31.975 7.015 ;
      RECT 31.57 6.29 31.86 6.52 ;
      RECT 31.165 2.395 31.27 2.965 ;
      RECT 31.165 2.73 31.49 2.96 ;
      RECT 31.165 2.76 31.66 2.93 ;
      RECT 31.165 2.395 31.355 2.96 ;
      RECT 30.58 2.36 30.87 2.59 ;
      RECT 30.58 2.395 31.355 2.565 ;
      RECT 30.64 0.88 30.81 2.59 ;
      RECT 30.58 0.88 30.87 1.11 ;
      RECT 30.58 7.77 30.87 8 ;
      RECT 30.64 6.29 30.81 8 ;
      RECT 30.58 6.29 30.87 6.52 ;
      RECT 30.58 6.325 31.435 6.485 ;
      RECT 31.265 5.92 31.435 6.485 ;
      RECT 30.58 6.32 30.975 6.485 ;
      RECT 31.2 5.92 31.49 6.15 ;
      RECT 31.2 5.95 31.66 6.12 ;
      RECT 30.21 2.73 30.5 2.96 ;
      RECT 30.21 2.76 30.67 2.93 ;
      RECT 30.275 1.655 30.44 2.96 ;
      RECT 28.79 1.625 29.08 1.855 ;
      RECT 28.79 1.655 30.44 1.825 ;
      RECT 28.85 0.885 29.02 1.855 ;
      RECT 28.79 0.885 29.08 1.115 ;
      RECT 28.79 7.765 29.08 7.995 ;
      RECT 28.85 7.025 29.02 7.995 ;
      RECT 28.85 7.12 30.44 7.29 ;
      RECT 30.27 5.92 30.44 7.29 ;
      RECT 28.79 7.025 29.08 7.255 ;
      RECT 30.21 5.92 30.5 6.15 ;
      RECT 30.21 5.95 30.67 6.12 ;
      RECT 29.22 1.965 29.57 2.315 ;
      RECT 26.915 2.025 29.57 2.195 ;
      RECT 26.915 1.46 27.085 2.195 ;
      RECT 26.825 1.46 27.165 1.81 ;
      RECT 29.245 6.655 29.57 6.98 ;
      RECT 23.805 6.61 24.155 6.96 ;
      RECT 29.22 6.655 29.57 6.885 ;
      RECT 23.605 6.655 24.155 6.885 ;
      RECT 23.435 6.685 29.57 6.855 ;
      RECT 28.445 2.365 28.765 2.685 ;
      RECT 28.415 2.365 28.765 2.595 ;
      RECT 28.245 2.395 28.765 2.565 ;
      RECT 28.445 6.255 28.765 6.545 ;
      RECT 28.415 6.285 28.765 6.515 ;
      RECT 28.245 6.315 28.765 6.485 ;
      RECT 24.9 2.465 25.19 2.695 ;
      RECT 24.9 2.465 25.355 2.65 ;
      RECT 25.215 2.37 25.835 2.51 ;
      RECT 25.605 2.17 25.925 2.43 ;
      RECT 24.285 2.45 24.605 2.71 ;
      RECT 24.285 2.45 24.75 2.695 ;
      RECT 24.61 2.07 24.75 2.695 ;
      RECT 24.61 2.07 24.875 2.21 ;
      RECT 25.14 1.905 25.43 2.135 ;
      RECT 24.735 1.95 25.43 2.09 ;
      RECT 24.18 3.29 24.47 3.815 ;
      RECT 24.165 3.29 24.485 3.55 ;
      RECT 23.905 1.89 24.225 2.15 ;
      RECT 23.905 1.905 24.47 2.135 ;
      RECT 23.18 3.585 23.47 3.815 ;
      RECT 23.375 2.23 23.515 3.77 ;
      RECT 23.42 2.185 23.71 2.415 ;
      RECT 23.015 2.23 23.71 2.37 ;
      RECT 23.015 2.07 23.155 2.37 ;
      RECT 21.555 2.07 23.155 2.21 ;
      RECT 21.465 1.89 21.785 2.15 ;
      RECT 21.465 1.905 22.03 2.15 ;
      RECT 23.175 7.765 23.465 7.995 ;
      RECT 23.235 7.025 23.405 7.995 ;
      RECT 23.155 7.075 23.525 7.425 ;
      RECT 23.155 7.055 23.465 7.425 ;
      RECT 23.175 7.025 23.465 7.425 ;
      RECT 20.575 2.93 23.155 3.07 ;
      RECT 22.94 2.745 23.23 2.975 ;
      RECT 20.5 2.745 21.165 2.975 ;
      RECT 20.845 2.73 21.165 3.07 ;
      RECT 21.845 2.45 22.165 2.71 ;
      RECT 21.845 2.465 22.27 2.695 ;
      RECT 20.485 2.17 20.805 2.43 ;
      RECT 20.98 2.185 21.27 2.415 ;
      RECT 20.485 2.23 21.27 2.37 ;
      RECT 20.605 3.29 20.925 3.55 ;
      RECT 19.765 3.29 20.085 3.55 ;
      RECT 20.605 3.305 21.03 3.535 ;
      RECT 19.765 3.35 21.03 3.49 ;
      RECT 19.3 3.025 19.59 3.255 ;
      RECT 19.375 1.95 19.515 3.255 ;
      RECT 19.025 2.45 19.515 2.71 ;
      RECT 18.78 2.465 19.515 2.695 ;
      RECT 19.78 1.905 20.07 2.135 ;
      RECT 19.375 1.95 20.07 2.09 ;
      RECT 18.54 3.305 18.83 3.535 ;
      RECT 18.54 3.305 18.995 3.49 ;
      RECT 18.855 2.93 18.995 3.49 ;
      RECT 18.495 2.93 18.995 3.07 ;
      RECT 18.495 1.95 18.635 3.07 ;
      RECT 18.285 1.89 18.605 2.15 ;
      RECT 18.045 3.57 18.365 3.83 ;
      RECT 17.34 3.585 17.63 3.815 ;
      RECT 17.34 3.63 18.365 3.77 ;
      RECT 17.415 3.58 17.675 3.77 ;
      RECT 17.805 2.45 18.125 2.71 ;
      RECT 17.805 2.465 18.35 2.695 ;
      RECT 17.805 3.01 18.125 3.27 ;
      RECT 17.805 3.025 18.35 3.255 ;
      RECT 16.845 3.01 17.165 3.27 ;
      RECT 16.935 1.95 17.075 3.27 ;
      RECT 17.34 1.905 17.63 2.135 ;
      RECT 16.935 1.95 17.63 2.09 ;
      RECT 15.245 7.77 15.535 8 ;
      RECT 15.305 6.29 15.475 8 ;
      RECT 15.3 6.655 15.65 7.005 ;
      RECT 15.245 6.29 15.535 6.52 ;
      RECT 14.84 2.395 14.945 2.965 ;
      RECT 14.84 2.73 15.165 2.96 ;
      RECT 14.84 2.76 15.335 2.93 ;
      RECT 14.84 2.395 15.03 2.96 ;
      RECT 14.255 2.36 14.545 2.59 ;
      RECT 14.255 2.395 15.03 2.565 ;
      RECT 14.315 0.88 14.485 2.59 ;
      RECT 14.255 0.88 14.545 1.11 ;
      RECT 14.255 7.77 14.545 8 ;
      RECT 14.315 6.29 14.485 8 ;
      RECT 14.255 6.29 14.545 6.52 ;
      RECT 14.255 6.325 15.11 6.485 ;
      RECT 14.94 5.92 15.11 6.485 ;
      RECT 14.255 6.32 14.65 6.485 ;
      RECT 14.875 5.92 15.165 6.15 ;
      RECT 14.875 5.95 15.335 6.12 ;
      RECT 13.885 2.73 14.175 2.96 ;
      RECT 13.885 2.76 14.345 2.93 ;
      RECT 13.95 1.655 14.115 2.96 ;
      RECT 12.465 1.625 12.755 1.855 ;
      RECT 12.465 1.655 14.115 1.825 ;
      RECT 12.525 0.885 12.695 1.855 ;
      RECT 12.465 0.885 12.755 1.115 ;
      RECT 12.465 7.765 12.755 7.995 ;
      RECT 12.525 7.025 12.695 7.995 ;
      RECT 12.525 7.12 14.115 7.29 ;
      RECT 13.945 5.92 14.115 7.29 ;
      RECT 12.465 7.025 12.755 7.255 ;
      RECT 13.885 5.92 14.175 6.15 ;
      RECT 13.885 5.95 14.345 6.12 ;
      RECT 12.895 1.965 13.245 2.315 ;
      RECT 10.59 2.025 13.245 2.195 ;
      RECT 10.59 1.46 10.76 2.195 ;
      RECT 10.5 1.46 10.84 1.81 ;
      RECT 12.92 6.655 13.245 6.98 ;
      RECT 8.315 6.605 8.665 6.955 ;
      RECT 12.895 6.655 13.245 6.885 ;
      RECT 7.28 6.655 7.57 6.885 ;
      RECT 7.11 6.685 13.245 6.855 ;
      RECT 12.12 2.365 12.44 2.685 ;
      RECT 12.09 2.365 12.44 2.595 ;
      RECT 11.92 2.395 12.44 2.565 ;
      RECT 12.12 6.255 12.44 6.545 ;
      RECT 12.09 6.285 12.44 6.515 ;
      RECT 11.92 6.315 12.44 6.485 ;
      RECT 8.575 2.465 8.865 2.695 ;
      RECT 8.575 2.465 9.03 2.65 ;
      RECT 8.89 2.37 9.51 2.51 ;
      RECT 9.28 2.17 9.6 2.43 ;
      RECT 7.96 2.45 8.28 2.71 ;
      RECT 7.96 2.45 8.425 2.695 ;
      RECT 8.285 2.07 8.425 2.695 ;
      RECT 8.285 2.07 8.55 2.21 ;
      RECT 8.815 1.905 9.105 2.135 ;
      RECT 8.41 1.95 9.105 2.09 ;
      RECT 7.855 3.29 8.145 3.815 ;
      RECT 7.84 3.29 8.16 3.55 ;
      RECT 7.58 1.89 7.9 2.15 ;
      RECT 7.58 1.905 8.145 2.135 ;
      RECT 6.855 3.585 7.145 3.815 ;
      RECT 7.05 2.23 7.19 3.77 ;
      RECT 7.095 2.185 7.385 2.415 ;
      RECT 6.69 2.23 7.385 2.37 ;
      RECT 6.69 2.07 6.83 2.37 ;
      RECT 5.23 2.07 6.83 2.21 ;
      RECT 5.14 1.89 5.46 2.15 ;
      RECT 5.14 1.905 5.705 2.15 ;
      RECT 6.85 7.765 7.14 7.995 ;
      RECT 6.91 7.025 7.08 7.995 ;
      RECT 6.83 7.075 7.2 7.425 ;
      RECT 6.83 7.055 7.14 7.425 ;
      RECT 6.85 7.025 7.14 7.425 ;
      RECT 4.25 2.93 6.83 3.07 ;
      RECT 6.615 2.745 6.905 2.975 ;
      RECT 4.175 2.745 4.84 2.975 ;
      RECT 4.52 2.73 4.84 3.07 ;
      RECT 5.52 2.45 5.84 2.71 ;
      RECT 5.52 2.465 5.945 2.695 ;
      RECT 4.16 2.17 4.48 2.43 ;
      RECT 4.655 2.185 4.945 2.415 ;
      RECT 4.16 2.23 4.945 2.37 ;
      RECT 4.28 3.29 4.6 3.55 ;
      RECT 3.44 3.29 3.76 3.55 ;
      RECT 4.28 3.305 4.705 3.535 ;
      RECT 3.44 3.35 4.705 3.49 ;
      RECT 2.975 3.025 3.265 3.255 ;
      RECT 3.05 1.95 3.19 3.255 ;
      RECT 2.7 2.45 3.19 2.71 ;
      RECT 2.455 2.465 3.19 2.695 ;
      RECT 3.455 1.905 3.745 2.135 ;
      RECT 3.05 1.95 3.745 2.09 ;
      RECT 2.215 3.305 2.505 3.535 ;
      RECT 2.215 3.305 2.67 3.49 ;
      RECT 2.53 2.93 2.67 3.49 ;
      RECT 2.17 2.93 2.67 3.07 ;
      RECT 2.17 1.95 2.31 3.07 ;
      RECT 1.96 1.89 2.28 2.15 ;
      RECT 1.72 3.57 2.04 3.83 ;
      RECT 1.015 3.585 1.305 3.815 ;
      RECT 1.015 3.63 2.04 3.77 ;
      RECT 1.09 3.58 1.35 3.77 ;
      RECT 1.48 2.45 1.8 2.71 ;
      RECT 1.48 2.465 2.025 2.695 ;
      RECT 1.48 3.01 1.8 3.27 ;
      RECT 1.48 3.025 2.025 3.255 ;
      RECT 0.52 3.01 0.84 3.27 ;
      RECT 0.61 1.95 0.75 3.27 ;
      RECT 1.015 1.905 1.305 2.135 ;
      RECT 0.61 1.95 1.305 2.09 ;
      RECT -1.73 7.765 -1.44 7.995 ;
      RECT -1.67 7.025 -1.5 7.995 ;
      RECT -1.76 7.025 -1.41 7.315 ;
      RECT -2.135 6.285 -1.785 6.575 ;
      RECT -2.275 6.315 -1.785 6.485 ;
      RECT 71.42 2.45 71.74 2.71 ;
      RECT 68.98 2.45 69.3 2.71 ;
      RECT 55.095 2.45 55.415 2.71 ;
      RECT 52.655 2.45 52.975 2.71 ;
      RECT 38.77 2.45 39.09 2.71 ;
      RECT 36.33 2.45 36.65 2.71 ;
      RECT 22.445 2.45 22.765 2.71 ;
      RECT 20.005 2.45 20.325 2.71 ;
      RECT 6.12 2.45 6.44 2.71 ;
      RECT 3.68 2.45 4 2.71 ;
    LAYER mcon ;
      RECT 80.605 6.32 80.775 6.49 ;
      RECT 80.61 6.315 80.78 6.485 ;
      RECT 64.28 6.32 64.45 6.49 ;
      RECT 64.285 6.315 64.455 6.485 ;
      RECT 47.955 6.32 48.125 6.49 ;
      RECT 47.96 6.315 48.13 6.485 ;
      RECT 31.63 6.32 31.8 6.49 ;
      RECT 31.635 6.315 31.805 6.485 ;
      RECT 15.305 6.32 15.475 6.49 ;
      RECT 15.31 6.315 15.48 6.485 ;
      RECT 80.605 7.8 80.775 7.97 ;
      RECT 80.235 2.76 80.405 2.93 ;
      RECT 80.235 5.95 80.405 6.12 ;
      RECT 79.615 0.91 79.785 1.08 ;
      RECT 79.615 2.39 79.785 2.56 ;
      RECT 79.615 6.32 79.785 6.49 ;
      RECT 79.615 7.8 79.785 7.97 ;
      RECT 79.245 2.76 79.415 2.93 ;
      RECT 79.245 5.95 79.415 6.12 ;
      RECT 78.255 2.025 78.425 2.195 ;
      RECT 78.255 6.685 78.425 6.855 ;
      RECT 77.825 0.915 77.995 1.085 ;
      RECT 77.825 1.655 77.995 1.825 ;
      RECT 77.825 7.055 77.995 7.225 ;
      RECT 77.825 7.795 77.995 7.965 ;
      RECT 77.45 2.395 77.62 2.565 ;
      RECT 77.45 6.315 77.62 6.485 ;
      RECT 74.175 1.935 74.345 2.105 ;
      RECT 73.935 2.495 74.105 2.665 ;
      RECT 73.455 2.495 73.625 2.665 ;
      RECT 73.215 1.935 73.385 2.105 ;
      RECT 73.215 3.615 73.385 3.785 ;
      RECT 72.64 6.685 72.81 6.855 ;
      RECT 72.455 2.215 72.625 2.385 ;
      RECT 72.215 3.615 72.385 3.785 ;
      RECT 72.21 7.055 72.38 7.225 ;
      RECT 72.21 7.795 72.38 7.965 ;
      RECT 71.975 2.775 72.145 2.945 ;
      RECT 71.495 2.495 71.665 2.665 ;
      RECT 71.015 2.495 71.185 2.665 ;
      RECT 70.775 1.935 70.945 2.105 ;
      RECT 70.015 2.215 70.185 2.385 ;
      RECT 69.775 3.335 69.945 3.505 ;
      RECT 69.535 2.775 69.705 2.945 ;
      RECT 69.055 2.495 69.225 2.665 ;
      RECT 68.815 1.935 68.985 2.105 ;
      RECT 68.815 3.335 68.985 3.505 ;
      RECT 68.335 3.055 68.505 3.225 ;
      RECT 67.815 2.495 67.985 2.665 ;
      RECT 67.575 3.335 67.745 3.505 ;
      RECT 67.335 1.935 67.505 2.105 ;
      RECT 67.095 2.495 67.265 2.665 ;
      RECT 67.095 3.055 67.265 3.225 ;
      RECT 66.375 1.935 66.545 2.105 ;
      RECT 66.375 3.615 66.545 3.785 ;
      RECT 65.895 3.055 66.065 3.225 ;
      RECT 64.28 7.8 64.45 7.97 ;
      RECT 63.91 2.76 64.08 2.93 ;
      RECT 63.91 5.95 64.08 6.12 ;
      RECT 63.29 0.91 63.46 1.08 ;
      RECT 63.29 2.39 63.46 2.56 ;
      RECT 63.29 6.32 63.46 6.49 ;
      RECT 63.29 7.8 63.46 7.97 ;
      RECT 62.92 2.76 63.09 2.93 ;
      RECT 62.92 5.95 63.09 6.12 ;
      RECT 61.93 2.025 62.1 2.195 ;
      RECT 61.93 6.685 62.1 6.855 ;
      RECT 61.5 0.915 61.67 1.085 ;
      RECT 61.5 1.655 61.67 1.825 ;
      RECT 61.5 7.055 61.67 7.225 ;
      RECT 61.5 7.795 61.67 7.965 ;
      RECT 61.125 2.395 61.295 2.565 ;
      RECT 61.125 6.315 61.295 6.485 ;
      RECT 57.85 1.935 58.02 2.105 ;
      RECT 57.61 2.495 57.78 2.665 ;
      RECT 57.13 2.495 57.3 2.665 ;
      RECT 56.89 1.935 57.06 2.105 ;
      RECT 56.89 3.615 57.06 3.785 ;
      RECT 56.315 6.685 56.485 6.855 ;
      RECT 56.13 2.215 56.3 2.385 ;
      RECT 55.89 3.615 56.06 3.785 ;
      RECT 55.885 7.055 56.055 7.225 ;
      RECT 55.885 7.795 56.055 7.965 ;
      RECT 55.65 2.775 55.82 2.945 ;
      RECT 55.17 2.495 55.34 2.665 ;
      RECT 54.69 2.495 54.86 2.665 ;
      RECT 54.45 1.935 54.62 2.105 ;
      RECT 53.69 2.215 53.86 2.385 ;
      RECT 53.45 3.335 53.62 3.505 ;
      RECT 53.21 2.775 53.38 2.945 ;
      RECT 52.73 2.495 52.9 2.665 ;
      RECT 52.49 1.935 52.66 2.105 ;
      RECT 52.49 3.335 52.66 3.505 ;
      RECT 52.01 3.055 52.18 3.225 ;
      RECT 51.49 2.495 51.66 2.665 ;
      RECT 51.25 3.335 51.42 3.505 ;
      RECT 51.01 1.935 51.18 2.105 ;
      RECT 50.77 2.495 50.94 2.665 ;
      RECT 50.77 3.055 50.94 3.225 ;
      RECT 50.05 1.935 50.22 2.105 ;
      RECT 50.05 3.615 50.22 3.785 ;
      RECT 49.57 3.055 49.74 3.225 ;
      RECT 47.955 7.8 48.125 7.97 ;
      RECT 47.585 2.76 47.755 2.93 ;
      RECT 47.585 5.95 47.755 6.12 ;
      RECT 46.965 0.91 47.135 1.08 ;
      RECT 46.965 2.39 47.135 2.56 ;
      RECT 46.965 6.32 47.135 6.49 ;
      RECT 46.965 7.8 47.135 7.97 ;
      RECT 46.595 2.76 46.765 2.93 ;
      RECT 46.595 5.95 46.765 6.12 ;
      RECT 45.605 2.025 45.775 2.195 ;
      RECT 45.605 6.685 45.775 6.855 ;
      RECT 45.175 0.915 45.345 1.085 ;
      RECT 45.175 1.655 45.345 1.825 ;
      RECT 45.175 7.055 45.345 7.225 ;
      RECT 45.175 7.795 45.345 7.965 ;
      RECT 44.8 2.395 44.97 2.565 ;
      RECT 44.8 6.315 44.97 6.485 ;
      RECT 41.525 1.935 41.695 2.105 ;
      RECT 41.285 2.495 41.455 2.665 ;
      RECT 40.805 2.495 40.975 2.665 ;
      RECT 40.565 1.935 40.735 2.105 ;
      RECT 40.565 3.615 40.735 3.785 ;
      RECT 39.99 6.685 40.16 6.855 ;
      RECT 39.805 2.215 39.975 2.385 ;
      RECT 39.565 3.615 39.735 3.785 ;
      RECT 39.56 7.055 39.73 7.225 ;
      RECT 39.56 7.795 39.73 7.965 ;
      RECT 39.325 2.775 39.495 2.945 ;
      RECT 38.845 2.495 39.015 2.665 ;
      RECT 38.365 2.495 38.535 2.665 ;
      RECT 38.125 1.935 38.295 2.105 ;
      RECT 37.365 2.215 37.535 2.385 ;
      RECT 37.125 3.335 37.295 3.505 ;
      RECT 36.885 2.775 37.055 2.945 ;
      RECT 36.405 2.495 36.575 2.665 ;
      RECT 36.165 1.935 36.335 2.105 ;
      RECT 36.165 3.335 36.335 3.505 ;
      RECT 35.685 3.055 35.855 3.225 ;
      RECT 35.165 2.495 35.335 2.665 ;
      RECT 34.925 3.335 35.095 3.505 ;
      RECT 34.685 1.935 34.855 2.105 ;
      RECT 34.445 2.495 34.615 2.665 ;
      RECT 34.445 3.055 34.615 3.225 ;
      RECT 33.725 1.935 33.895 2.105 ;
      RECT 33.725 3.615 33.895 3.785 ;
      RECT 33.245 3.055 33.415 3.225 ;
      RECT 31.63 7.8 31.8 7.97 ;
      RECT 31.26 2.76 31.43 2.93 ;
      RECT 31.26 5.95 31.43 6.12 ;
      RECT 30.64 0.91 30.81 1.08 ;
      RECT 30.64 2.39 30.81 2.56 ;
      RECT 30.64 6.32 30.81 6.49 ;
      RECT 30.64 7.8 30.81 7.97 ;
      RECT 30.27 2.76 30.44 2.93 ;
      RECT 30.27 5.95 30.44 6.12 ;
      RECT 29.28 2.025 29.45 2.195 ;
      RECT 29.28 6.685 29.45 6.855 ;
      RECT 28.85 0.915 29.02 1.085 ;
      RECT 28.85 1.655 29.02 1.825 ;
      RECT 28.85 7.055 29.02 7.225 ;
      RECT 28.85 7.795 29.02 7.965 ;
      RECT 28.475 2.395 28.645 2.565 ;
      RECT 28.475 6.315 28.645 6.485 ;
      RECT 25.2 1.935 25.37 2.105 ;
      RECT 24.96 2.495 25.13 2.665 ;
      RECT 24.48 2.495 24.65 2.665 ;
      RECT 24.24 1.935 24.41 2.105 ;
      RECT 24.24 3.615 24.41 3.785 ;
      RECT 23.665 6.685 23.835 6.855 ;
      RECT 23.48 2.215 23.65 2.385 ;
      RECT 23.24 3.615 23.41 3.785 ;
      RECT 23.235 7.055 23.405 7.225 ;
      RECT 23.235 7.795 23.405 7.965 ;
      RECT 23 2.775 23.17 2.945 ;
      RECT 22.52 2.495 22.69 2.665 ;
      RECT 22.04 2.495 22.21 2.665 ;
      RECT 21.8 1.935 21.97 2.105 ;
      RECT 21.04 2.215 21.21 2.385 ;
      RECT 20.8 3.335 20.97 3.505 ;
      RECT 20.56 2.775 20.73 2.945 ;
      RECT 20.08 2.495 20.25 2.665 ;
      RECT 19.84 1.935 20.01 2.105 ;
      RECT 19.84 3.335 20.01 3.505 ;
      RECT 19.36 3.055 19.53 3.225 ;
      RECT 18.84 2.495 19.01 2.665 ;
      RECT 18.6 3.335 18.77 3.505 ;
      RECT 18.36 1.935 18.53 2.105 ;
      RECT 18.12 2.495 18.29 2.665 ;
      RECT 18.12 3.055 18.29 3.225 ;
      RECT 17.4 1.935 17.57 2.105 ;
      RECT 17.4 3.615 17.57 3.785 ;
      RECT 16.92 3.055 17.09 3.225 ;
      RECT 15.305 7.8 15.475 7.97 ;
      RECT 14.935 2.76 15.105 2.93 ;
      RECT 14.935 5.95 15.105 6.12 ;
      RECT 14.315 0.91 14.485 1.08 ;
      RECT 14.315 2.39 14.485 2.56 ;
      RECT 14.315 6.32 14.485 6.49 ;
      RECT 14.315 7.8 14.485 7.97 ;
      RECT 13.945 2.76 14.115 2.93 ;
      RECT 13.945 5.95 14.115 6.12 ;
      RECT 12.955 2.025 13.125 2.195 ;
      RECT 12.955 6.685 13.125 6.855 ;
      RECT 12.525 0.915 12.695 1.085 ;
      RECT 12.525 1.655 12.695 1.825 ;
      RECT 12.525 7.055 12.695 7.225 ;
      RECT 12.525 7.795 12.695 7.965 ;
      RECT 12.15 2.395 12.32 2.565 ;
      RECT 12.15 6.315 12.32 6.485 ;
      RECT 8.875 1.935 9.045 2.105 ;
      RECT 8.635 2.495 8.805 2.665 ;
      RECT 8.155 2.495 8.325 2.665 ;
      RECT 7.915 1.935 8.085 2.105 ;
      RECT 7.915 3.615 8.085 3.785 ;
      RECT 7.34 6.685 7.51 6.855 ;
      RECT 7.155 2.215 7.325 2.385 ;
      RECT 6.915 3.615 7.085 3.785 ;
      RECT 6.91 7.055 7.08 7.225 ;
      RECT 6.91 7.795 7.08 7.965 ;
      RECT 6.675 2.775 6.845 2.945 ;
      RECT 6.195 2.495 6.365 2.665 ;
      RECT 5.715 2.495 5.885 2.665 ;
      RECT 5.475 1.935 5.645 2.105 ;
      RECT 4.715 2.215 4.885 2.385 ;
      RECT 4.475 3.335 4.645 3.505 ;
      RECT 4.235 2.775 4.405 2.945 ;
      RECT 3.755 2.495 3.925 2.665 ;
      RECT 3.515 1.935 3.685 2.105 ;
      RECT 3.515 3.335 3.685 3.505 ;
      RECT 3.035 3.055 3.205 3.225 ;
      RECT 2.515 2.495 2.685 2.665 ;
      RECT 2.275 3.335 2.445 3.505 ;
      RECT 2.035 1.935 2.205 2.105 ;
      RECT 1.795 2.495 1.965 2.665 ;
      RECT 1.795 3.055 1.965 3.225 ;
      RECT 1.075 1.935 1.245 2.105 ;
      RECT 1.075 3.615 1.245 3.785 ;
      RECT 0.595 3.055 0.765 3.225 ;
      RECT -1.67 7.055 -1.5 7.225 ;
      RECT -1.67 7.795 -1.5 7.965 ;
      RECT -2.045 6.315 -1.875 6.485 ;
    LAYER li1 ;
      RECT 80.605 5.02 80.775 6.49 ;
      RECT 80.605 6.315 80.78 6.485 ;
      RECT 80.235 1.74 80.405 2.93 ;
      RECT 80.235 1.74 80.705 1.91 ;
      RECT 80.235 6.97 80.705 7.14 ;
      RECT 80.235 5.95 80.405 7.14 ;
      RECT 79.245 1.74 79.415 2.93 ;
      RECT 79.245 1.74 79.715 1.91 ;
      RECT 79.245 6.97 79.715 7.14 ;
      RECT 79.245 5.95 79.415 7.14 ;
      RECT 77.395 2.635 77.565 3.865 ;
      RECT 77.45 0.855 77.62 2.805 ;
      RECT 77.395 0.575 77.565 1.025 ;
      RECT 77.395 7.855 77.565 8.305 ;
      RECT 77.45 6.075 77.62 8.025 ;
      RECT 77.395 5.015 77.565 6.245 ;
      RECT 76.875 0.575 77.045 3.865 ;
      RECT 76.875 2.075 77.28 2.405 ;
      RECT 76.875 1.235 77.28 1.565 ;
      RECT 76.875 5.015 77.045 8.305 ;
      RECT 76.875 7.315 77.28 7.645 ;
      RECT 76.875 6.475 77.28 6.805 ;
      RECT 74.175 1.835 74.345 2.105 ;
      RECT 74.175 1.835 74.905 2.005 ;
      RECT 74.095 3.225 74.425 3.395 ;
      RECT 73.335 3.055 74.345 3.225 ;
      RECT 73.335 2.575 73.505 3.225 ;
      RECT 73.455 2.495 73.625 2.825 ;
      RECT 72.615 3.225 72.945 3.395 ;
      RECT 70.695 3.225 71.985 3.395 ;
      RECT 71.735 3.14 72.865 3.31 ;
      RECT 72.455 2.215 72.865 2.385 ;
      RECT 72.695 1.755 72.865 2.385 ;
      RECT 71.26 5.015 71.43 8.305 ;
      RECT 71.26 7.315 71.665 7.645 ;
      RECT 71.26 6.475 71.665 6.805 ;
      RECT 69.935 2.575 71.265 2.745 ;
      RECT 71.015 2.495 71.185 2.745 ;
      RECT 70.015 2.175 70.185 2.385 ;
      RECT 70.015 2.175 70.505 2.345 ;
      RECT 68.695 3.335 68.985 3.505 ;
      RECT 68.695 2.575 68.865 3.505 ;
      RECT 68.495 2.575 68.865 2.745 ;
      RECT 67.495 2.575 67.985 2.745 ;
      RECT 67.815 2.495 67.985 2.745 ;
      RECT 67.575 3.335 67.985 3.505 ;
      RECT 67.815 3.145 67.985 3.505 ;
      RECT 66.615 3.055 67.265 3.225 ;
      RECT 66.615 2.495 66.785 3.225 ;
      RECT 66.255 3.615 66.545 3.785 ;
      RECT 66.255 2.575 66.425 3.785 ;
      RECT 66.055 2.575 66.425 2.745 ;
      RECT 64.28 5.02 64.45 6.49 ;
      RECT 64.28 6.315 64.455 6.485 ;
      RECT 63.91 1.74 64.08 2.93 ;
      RECT 63.91 1.74 64.38 1.91 ;
      RECT 63.91 6.97 64.38 7.14 ;
      RECT 63.91 5.95 64.08 7.14 ;
      RECT 62.92 1.74 63.09 2.93 ;
      RECT 62.92 1.74 63.39 1.91 ;
      RECT 62.92 6.97 63.39 7.14 ;
      RECT 62.92 5.95 63.09 7.14 ;
      RECT 61.07 2.635 61.24 3.865 ;
      RECT 61.125 0.855 61.295 2.805 ;
      RECT 61.07 0.575 61.24 1.025 ;
      RECT 61.07 7.855 61.24 8.305 ;
      RECT 61.125 6.075 61.295 8.025 ;
      RECT 61.07 5.015 61.24 6.245 ;
      RECT 60.55 0.575 60.72 3.865 ;
      RECT 60.55 2.075 60.955 2.405 ;
      RECT 60.55 1.235 60.955 1.565 ;
      RECT 60.55 5.015 60.72 8.305 ;
      RECT 60.55 7.315 60.955 7.645 ;
      RECT 60.55 6.475 60.955 6.805 ;
      RECT 57.85 1.835 58.02 2.105 ;
      RECT 57.85 1.835 58.58 2.005 ;
      RECT 57.77 3.225 58.1 3.395 ;
      RECT 57.01 3.055 58.02 3.225 ;
      RECT 57.01 2.575 57.18 3.225 ;
      RECT 57.13 2.495 57.3 2.825 ;
      RECT 56.29 3.225 56.62 3.395 ;
      RECT 54.37 3.225 55.66 3.395 ;
      RECT 55.41 3.14 56.54 3.31 ;
      RECT 56.13 2.215 56.54 2.385 ;
      RECT 56.37 1.755 56.54 2.385 ;
      RECT 54.935 5.015 55.105 8.305 ;
      RECT 54.935 7.315 55.34 7.645 ;
      RECT 54.935 6.475 55.34 6.805 ;
      RECT 53.61 2.575 54.94 2.745 ;
      RECT 54.69 2.495 54.86 2.745 ;
      RECT 53.69 2.175 53.86 2.385 ;
      RECT 53.69 2.175 54.18 2.345 ;
      RECT 52.37 3.335 52.66 3.505 ;
      RECT 52.37 2.575 52.54 3.505 ;
      RECT 52.17 2.575 52.54 2.745 ;
      RECT 51.17 2.575 51.66 2.745 ;
      RECT 51.49 2.495 51.66 2.745 ;
      RECT 51.25 3.335 51.66 3.505 ;
      RECT 51.49 3.145 51.66 3.505 ;
      RECT 50.29 3.055 50.94 3.225 ;
      RECT 50.29 2.495 50.46 3.225 ;
      RECT 49.93 3.615 50.22 3.785 ;
      RECT 49.93 2.575 50.1 3.785 ;
      RECT 49.73 2.575 50.1 2.745 ;
      RECT 47.955 5.02 48.125 6.49 ;
      RECT 47.955 6.315 48.13 6.485 ;
      RECT 47.585 1.74 47.755 2.93 ;
      RECT 47.585 1.74 48.055 1.91 ;
      RECT 47.585 6.97 48.055 7.14 ;
      RECT 47.585 5.95 47.755 7.14 ;
      RECT 46.595 1.74 46.765 2.93 ;
      RECT 46.595 1.74 47.065 1.91 ;
      RECT 46.595 6.97 47.065 7.14 ;
      RECT 46.595 5.95 46.765 7.14 ;
      RECT 44.745 2.635 44.915 3.865 ;
      RECT 44.8 0.855 44.97 2.805 ;
      RECT 44.745 0.575 44.915 1.025 ;
      RECT 44.745 7.855 44.915 8.305 ;
      RECT 44.8 6.075 44.97 8.025 ;
      RECT 44.745 5.015 44.915 6.245 ;
      RECT 44.225 0.575 44.395 3.865 ;
      RECT 44.225 2.075 44.63 2.405 ;
      RECT 44.225 1.235 44.63 1.565 ;
      RECT 44.225 5.015 44.395 8.305 ;
      RECT 44.225 7.315 44.63 7.645 ;
      RECT 44.225 6.475 44.63 6.805 ;
      RECT 41.525 1.835 41.695 2.105 ;
      RECT 41.525 1.835 42.255 2.005 ;
      RECT 41.445 3.225 41.775 3.395 ;
      RECT 40.685 3.055 41.695 3.225 ;
      RECT 40.685 2.575 40.855 3.225 ;
      RECT 40.805 2.495 40.975 2.825 ;
      RECT 39.965 3.225 40.295 3.395 ;
      RECT 38.045 3.225 39.335 3.395 ;
      RECT 39.085 3.14 40.215 3.31 ;
      RECT 39.805 2.215 40.215 2.385 ;
      RECT 40.045 1.755 40.215 2.385 ;
      RECT 38.61 5.015 38.78 8.305 ;
      RECT 38.61 7.315 39.015 7.645 ;
      RECT 38.61 6.475 39.015 6.805 ;
      RECT 37.285 2.575 38.615 2.745 ;
      RECT 38.365 2.495 38.535 2.745 ;
      RECT 37.365 2.175 37.535 2.385 ;
      RECT 37.365 2.175 37.855 2.345 ;
      RECT 36.045 3.335 36.335 3.505 ;
      RECT 36.045 2.575 36.215 3.505 ;
      RECT 35.845 2.575 36.215 2.745 ;
      RECT 34.845 2.575 35.335 2.745 ;
      RECT 35.165 2.495 35.335 2.745 ;
      RECT 34.925 3.335 35.335 3.505 ;
      RECT 35.165 3.145 35.335 3.505 ;
      RECT 33.965 3.055 34.615 3.225 ;
      RECT 33.965 2.495 34.135 3.225 ;
      RECT 33.605 3.615 33.895 3.785 ;
      RECT 33.605 2.575 33.775 3.785 ;
      RECT 33.405 2.575 33.775 2.745 ;
      RECT 31.63 5.02 31.8 6.49 ;
      RECT 31.63 6.315 31.805 6.485 ;
      RECT 31.26 1.74 31.43 2.93 ;
      RECT 31.26 1.74 31.73 1.91 ;
      RECT 31.26 6.97 31.73 7.14 ;
      RECT 31.26 5.95 31.43 7.14 ;
      RECT 30.27 1.74 30.44 2.93 ;
      RECT 30.27 1.74 30.74 1.91 ;
      RECT 30.27 6.97 30.74 7.14 ;
      RECT 30.27 5.95 30.44 7.14 ;
      RECT 28.42 2.635 28.59 3.865 ;
      RECT 28.475 0.855 28.645 2.805 ;
      RECT 28.42 0.575 28.59 1.025 ;
      RECT 28.42 7.855 28.59 8.305 ;
      RECT 28.475 6.075 28.645 8.025 ;
      RECT 28.42 5.015 28.59 6.245 ;
      RECT 27.9 0.575 28.07 3.865 ;
      RECT 27.9 2.075 28.305 2.405 ;
      RECT 27.9 1.235 28.305 1.565 ;
      RECT 27.9 5.015 28.07 8.305 ;
      RECT 27.9 7.315 28.305 7.645 ;
      RECT 27.9 6.475 28.305 6.805 ;
      RECT 25.2 1.835 25.37 2.105 ;
      RECT 25.2 1.835 25.93 2.005 ;
      RECT 25.12 3.225 25.45 3.395 ;
      RECT 24.36 3.055 25.37 3.225 ;
      RECT 24.36 2.575 24.53 3.225 ;
      RECT 24.48 2.495 24.65 2.825 ;
      RECT 23.64 3.225 23.97 3.395 ;
      RECT 21.72 3.225 23.01 3.395 ;
      RECT 22.76 3.14 23.89 3.31 ;
      RECT 23.48 2.215 23.89 2.385 ;
      RECT 23.72 1.755 23.89 2.385 ;
      RECT 22.285 5.015 22.455 8.305 ;
      RECT 22.285 7.315 22.69 7.645 ;
      RECT 22.285 6.475 22.69 6.805 ;
      RECT 20.96 2.575 22.29 2.745 ;
      RECT 22.04 2.495 22.21 2.745 ;
      RECT 21.04 2.175 21.21 2.385 ;
      RECT 21.04 2.175 21.53 2.345 ;
      RECT 19.72 3.335 20.01 3.505 ;
      RECT 19.72 2.575 19.89 3.505 ;
      RECT 19.52 2.575 19.89 2.745 ;
      RECT 18.52 2.575 19.01 2.745 ;
      RECT 18.84 2.495 19.01 2.745 ;
      RECT 18.6 3.335 19.01 3.505 ;
      RECT 18.84 3.145 19.01 3.505 ;
      RECT 17.64 3.055 18.29 3.225 ;
      RECT 17.64 2.495 17.81 3.225 ;
      RECT 17.28 3.615 17.57 3.785 ;
      RECT 17.28 2.575 17.45 3.785 ;
      RECT 17.08 2.575 17.45 2.745 ;
      RECT 15.305 5.02 15.475 6.49 ;
      RECT 15.305 6.315 15.48 6.485 ;
      RECT 14.935 1.74 15.105 2.93 ;
      RECT 14.935 1.74 15.405 1.91 ;
      RECT 14.935 6.97 15.405 7.14 ;
      RECT 14.935 5.95 15.105 7.14 ;
      RECT 13.945 1.74 14.115 2.93 ;
      RECT 13.945 1.74 14.415 1.91 ;
      RECT 13.945 6.97 14.415 7.14 ;
      RECT 13.945 5.95 14.115 7.14 ;
      RECT 12.095 2.635 12.265 3.865 ;
      RECT 12.15 0.855 12.32 2.805 ;
      RECT 12.095 0.575 12.265 1.025 ;
      RECT 12.095 7.855 12.265 8.305 ;
      RECT 12.15 6.075 12.32 8.025 ;
      RECT 12.095 5.015 12.265 6.245 ;
      RECT 11.575 0.575 11.745 3.865 ;
      RECT 11.575 2.075 11.98 2.405 ;
      RECT 11.575 1.235 11.98 1.565 ;
      RECT 11.575 5.015 11.745 8.305 ;
      RECT 11.575 7.315 11.98 7.645 ;
      RECT 11.575 6.475 11.98 6.805 ;
      RECT 8.875 1.835 9.045 2.105 ;
      RECT 8.875 1.835 9.605 2.005 ;
      RECT 8.795 3.225 9.125 3.395 ;
      RECT 8.035 3.055 9.045 3.225 ;
      RECT 8.035 2.575 8.205 3.225 ;
      RECT 8.155 2.495 8.325 2.825 ;
      RECT 7.315 3.225 7.645 3.395 ;
      RECT 5.395 3.225 6.685 3.395 ;
      RECT 6.435 3.14 7.565 3.31 ;
      RECT 7.155 2.215 7.565 2.385 ;
      RECT 7.395 1.755 7.565 2.385 ;
      RECT 5.96 5.015 6.13 8.305 ;
      RECT 5.96 7.315 6.365 7.645 ;
      RECT 5.96 6.475 6.365 6.805 ;
      RECT 4.635 2.575 5.965 2.745 ;
      RECT 5.715 2.495 5.885 2.745 ;
      RECT 4.715 2.175 4.885 2.385 ;
      RECT 4.715 2.175 5.205 2.345 ;
      RECT 3.395 3.335 3.685 3.505 ;
      RECT 3.395 2.575 3.565 3.505 ;
      RECT 3.195 2.575 3.565 2.745 ;
      RECT 2.195 2.575 2.685 2.745 ;
      RECT 2.515 2.495 2.685 2.745 ;
      RECT 2.275 3.335 2.685 3.505 ;
      RECT 2.515 3.145 2.685 3.505 ;
      RECT 1.315 3.055 1.965 3.225 ;
      RECT 1.315 2.495 1.485 3.225 ;
      RECT 0.955 3.615 1.245 3.785 ;
      RECT 0.955 2.575 1.125 3.785 ;
      RECT 0.755 2.575 1.125 2.745 ;
      RECT -2.1 7.855 -1.93 8.305 ;
      RECT -2.045 6.075 -1.875 8.025 ;
      RECT -2.1 5.015 -1.93 6.245 ;
      RECT -2.62 5.015 -2.45 8.305 ;
      RECT -2.62 7.315 -2.215 7.645 ;
      RECT -2.62 6.475 -2.215 6.805 ;
      RECT 80.605 7.8 80.775 8.31 ;
      RECT 79.615 0.57 79.785 1.08 ;
      RECT 79.615 2.39 79.785 3.86 ;
      RECT 79.615 5.02 79.785 6.49 ;
      RECT 79.615 7.8 79.785 8.31 ;
      RECT 78.255 0.575 78.425 3.865 ;
      RECT 78.255 5.015 78.425 8.305 ;
      RECT 77.825 0.575 77.995 1.085 ;
      RECT 77.825 1.655 77.995 3.865 ;
      RECT 77.825 5.015 77.995 7.225 ;
      RECT 77.825 7.795 77.995 8.305 ;
      RECT 73.935 2.495 74.105 2.825 ;
      RECT 73.215 1.755 73.385 2.105 ;
      RECT 73.215 3.485 73.385 3.815 ;
      RECT 72.64 5.015 72.81 8.305 ;
      RECT 72.215 3.485 72.385 3.815 ;
      RECT 72.21 5.015 72.38 7.225 ;
      RECT 72.21 7.795 72.38 8.305 ;
      RECT 71.975 2.495 72.145 2.945 ;
      RECT 71.495 2.495 71.665 2.825 ;
      RECT 70.775 1.755 70.945 2.105 ;
      RECT 69.775 3.145 69.945 3.505 ;
      RECT 69.535 2.495 69.705 2.945 ;
      RECT 69.055 2.495 69.225 2.825 ;
      RECT 68.815 1.755 68.985 2.105 ;
      RECT 68.335 3.055 68.505 3.475 ;
      RECT 67.335 1.755 67.505 2.105 ;
      RECT 67.095 2.495 67.265 2.825 ;
      RECT 66.375 1.755 66.545 2.105 ;
      RECT 65.895 3.055 66.065 3.475 ;
      RECT 64.28 7.8 64.45 8.31 ;
      RECT 63.29 0.57 63.46 1.08 ;
      RECT 63.29 2.39 63.46 3.86 ;
      RECT 63.29 5.02 63.46 6.49 ;
      RECT 63.29 7.8 63.46 8.31 ;
      RECT 61.93 0.575 62.1 3.865 ;
      RECT 61.93 5.015 62.1 8.305 ;
      RECT 61.5 0.575 61.67 1.085 ;
      RECT 61.5 1.655 61.67 3.865 ;
      RECT 61.5 5.015 61.67 7.225 ;
      RECT 61.5 7.795 61.67 8.305 ;
      RECT 57.61 2.495 57.78 2.825 ;
      RECT 56.89 1.755 57.06 2.105 ;
      RECT 56.89 3.485 57.06 3.815 ;
      RECT 56.315 5.015 56.485 8.305 ;
      RECT 55.89 3.485 56.06 3.815 ;
      RECT 55.885 5.015 56.055 7.225 ;
      RECT 55.885 7.795 56.055 8.305 ;
      RECT 55.65 2.495 55.82 2.945 ;
      RECT 55.17 2.495 55.34 2.825 ;
      RECT 54.45 1.755 54.62 2.105 ;
      RECT 53.45 3.145 53.62 3.505 ;
      RECT 53.21 2.495 53.38 2.945 ;
      RECT 52.73 2.495 52.9 2.825 ;
      RECT 52.49 1.755 52.66 2.105 ;
      RECT 52.01 3.055 52.18 3.475 ;
      RECT 51.01 1.755 51.18 2.105 ;
      RECT 50.77 2.495 50.94 2.825 ;
      RECT 50.05 1.755 50.22 2.105 ;
      RECT 49.57 3.055 49.74 3.475 ;
      RECT 47.955 7.8 48.125 8.31 ;
      RECT 46.965 0.57 47.135 1.08 ;
      RECT 46.965 2.39 47.135 3.86 ;
      RECT 46.965 5.02 47.135 6.49 ;
      RECT 46.965 7.8 47.135 8.31 ;
      RECT 45.605 0.575 45.775 3.865 ;
      RECT 45.605 5.015 45.775 8.305 ;
      RECT 45.175 0.575 45.345 1.085 ;
      RECT 45.175 1.655 45.345 3.865 ;
      RECT 45.175 5.015 45.345 7.225 ;
      RECT 45.175 7.795 45.345 8.305 ;
      RECT 41.285 2.495 41.455 2.825 ;
      RECT 40.565 1.755 40.735 2.105 ;
      RECT 40.565 3.485 40.735 3.815 ;
      RECT 39.99 5.015 40.16 8.305 ;
      RECT 39.565 3.485 39.735 3.815 ;
      RECT 39.56 5.015 39.73 7.225 ;
      RECT 39.56 7.795 39.73 8.305 ;
      RECT 39.325 2.495 39.495 2.945 ;
      RECT 38.845 2.495 39.015 2.825 ;
      RECT 38.125 1.755 38.295 2.105 ;
      RECT 37.125 3.145 37.295 3.505 ;
      RECT 36.885 2.495 37.055 2.945 ;
      RECT 36.405 2.495 36.575 2.825 ;
      RECT 36.165 1.755 36.335 2.105 ;
      RECT 35.685 3.055 35.855 3.475 ;
      RECT 34.685 1.755 34.855 2.105 ;
      RECT 34.445 2.495 34.615 2.825 ;
      RECT 33.725 1.755 33.895 2.105 ;
      RECT 33.245 3.055 33.415 3.475 ;
      RECT 31.63 7.8 31.8 8.31 ;
      RECT 30.64 0.57 30.81 1.08 ;
      RECT 30.64 2.39 30.81 3.86 ;
      RECT 30.64 5.02 30.81 6.49 ;
      RECT 30.64 7.8 30.81 8.31 ;
      RECT 29.28 0.575 29.45 3.865 ;
      RECT 29.28 5.015 29.45 8.305 ;
      RECT 28.85 0.575 29.02 1.085 ;
      RECT 28.85 1.655 29.02 3.865 ;
      RECT 28.85 5.015 29.02 7.225 ;
      RECT 28.85 7.795 29.02 8.305 ;
      RECT 24.96 2.495 25.13 2.825 ;
      RECT 24.24 1.755 24.41 2.105 ;
      RECT 24.24 3.485 24.41 3.815 ;
      RECT 23.665 5.015 23.835 8.305 ;
      RECT 23.24 3.485 23.41 3.815 ;
      RECT 23.235 5.015 23.405 7.225 ;
      RECT 23.235 7.795 23.405 8.305 ;
      RECT 23 2.495 23.17 2.945 ;
      RECT 22.52 2.495 22.69 2.825 ;
      RECT 21.8 1.755 21.97 2.105 ;
      RECT 20.8 3.145 20.97 3.505 ;
      RECT 20.56 2.495 20.73 2.945 ;
      RECT 20.08 2.495 20.25 2.825 ;
      RECT 19.84 1.755 20.01 2.105 ;
      RECT 19.36 3.055 19.53 3.475 ;
      RECT 18.36 1.755 18.53 2.105 ;
      RECT 18.12 2.495 18.29 2.825 ;
      RECT 17.4 1.755 17.57 2.105 ;
      RECT 16.92 3.055 17.09 3.475 ;
      RECT 15.305 7.8 15.475 8.31 ;
      RECT 14.315 0.57 14.485 1.08 ;
      RECT 14.315 2.39 14.485 3.86 ;
      RECT 14.315 5.02 14.485 6.49 ;
      RECT 14.315 7.8 14.485 8.31 ;
      RECT 12.955 0.575 13.125 3.865 ;
      RECT 12.955 5.015 13.125 8.305 ;
      RECT 12.525 0.575 12.695 1.085 ;
      RECT 12.525 1.655 12.695 3.865 ;
      RECT 12.525 5.015 12.695 7.225 ;
      RECT 12.525 7.795 12.695 8.305 ;
      RECT 8.635 2.495 8.805 2.825 ;
      RECT 7.915 1.755 8.085 2.105 ;
      RECT 7.915 3.485 8.085 3.815 ;
      RECT 7.34 5.015 7.51 8.305 ;
      RECT 6.915 3.485 7.085 3.815 ;
      RECT 6.91 5.015 7.08 7.225 ;
      RECT 6.91 7.795 7.08 8.305 ;
      RECT 6.675 2.495 6.845 2.945 ;
      RECT 6.195 2.495 6.365 2.825 ;
      RECT 5.475 1.755 5.645 2.105 ;
      RECT 4.475 3.145 4.645 3.505 ;
      RECT 4.235 2.495 4.405 2.945 ;
      RECT 3.755 2.495 3.925 2.825 ;
      RECT 3.515 1.755 3.685 2.105 ;
      RECT 3.035 3.055 3.205 3.475 ;
      RECT 2.035 1.755 2.205 2.105 ;
      RECT 1.795 2.495 1.965 2.825 ;
      RECT 1.075 1.755 1.245 2.105 ;
      RECT 0.595 3.055 0.765 3.475 ;
      RECT -1.67 5.015 -1.5 7.225 ;
      RECT -1.67 7.795 -1.5 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2ea_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2ea_8_b0r2
  CLASS BLOCK ;
  ORIGIN 3.27 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ea_8_b0r2 ;
  SIZE 84.42 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 15.31 0.915 15.48 1.085 ;
        RECT 15.305 0.91 15.475 1.08 ;
        RECT 15.305 2.39 15.475 2.56 ;
      LAYER li1 ;
        RECT 15.31 0.915 15.48 1.085 ;
        RECT 15.305 0.57 15.475 1.08 ;
        RECT 15.305 2.39 15.475 3.86 ;
      LAYER met1 ;
        RECT 15.245 2.36 15.535 2.59 ;
        RECT 15.245 0.88 15.535 1.11 ;
        RECT 15.305 0.88 15.475 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 31.635 0.915 31.805 1.085 ;
        RECT 31.63 0.91 31.8 1.08 ;
        RECT 31.63 2.39 31.8 2.56 ;
      LAYER li1 ;
        RECT 31.635 0.915 31.805 1.085 ;
        RECT 31.63 0.57 31.8 1.08 ;
        RECT 31.63 2.39 31.8 3.86 ;
      LAYER met1 ;
        RECT 31.57 2.36 31.86 2.59 ;
        RECT 31.57 0.88 31.86 1.11 ;
        RECT 31.63 0.88 31.8 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 47.96 0.915 48.13 1.085 ;
        RECT 47.955 0.91 48.125 1.08 ;
        RECT 47.955 2.39 48.125 2.56 ;
      LAYER li1 ;
        RECT 47.96 0.915 48.13 1.085 ;
        RECT 47.955 0.57 48.125 1.08 ;
        RECT 47.955 2.39 48.125 3.86 ;
      LAYER met1 ;
        RECT 47.895 2.36 48.185 2.59 ;
        RECT 47.895 0.88 48.185 1.11 ;
        RECT 47.955 0.88 48.125 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 64.285 0.915 64.455 1.085 ;
        RECT 64.28 0.91 64.45 1.08 ;
        RECT 64.28 2.39 64.45 2.56 ;
      LAYER li1 ;
        RECT 64.285 0.915 64.455 1.085 ;
        RECT 64.28 0.57 64.45 1.08 ;
        RECT 64.28 2.39 64.45 3.86 ;
      LAYER met1 ;
        RECT 64.22 2.36 64.51 2.59 ;
        RECT 64.22 0.88 64.51 1.11 ;
        RECT 64.28 0.88 64.45 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 80.61 0.915 80.78 1.085 ;
        RECT 80.605 0.91 80.775 1.08 ;
        RECT 80.605 2.39 80.775 2.56 ;
      LAYER li1 ;
        RECT 80.61 0.915 80.78 1.085 ;
        RECT 80.605 0.57 80.775 1.08 ;
        RECT 80.605 2.39 80.775 3.86 ;
      LAYER met1 ;
        RECT 80.545 2.36 80.835 2.59 ;
        RECT 80.545 0.88 80.835 1.11 ;
        RECT 80.605 0.88 80.775 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 11.155 1.66 11.325 2.935 ;
        RECT 11.155 5.945 11.325 7.22 ;
        RECT 5.54 5.945 5.71 7.22 ;
      LAYER met2 ;
        RECT 11.08 2.705 11.42 3.055 ;
        RECT 11.07 5.84 11.41 6.19 ;
        RECT 11.155 2.705 11.325 6.19 ;
      LAYER met1 ;
        RECT 11.08 2.765 11.555 2.935 ;
        RECT 11.08 2.705 11.42 3.055 ;
        RECT 5.48 5.945 11.555 6.115 ;
        RECT 11.07 5.84 11.41 6.19 ;
        RECT 5.48 5.915 5.77 6.145 ;
      LAYER via1 ;
        RECT 11.17 5.94 11.32 6.09 ;
        RECT 11.18 2.805 11.33 2.955 ;
      LAYER mcon ;
        RECT 5.54 5.945 5.71 6.115 ;
        RECT 11.155 5.945 11.325 6.115 ;
        RECT 11.155 2.765 11.325 2.935 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 27.48 1.66 27.65 2.935 ;
        RECT 27.48 5.945 27.65 7.22 ;
        RECT 21.865 5.945 22.035 7.22 ;
      LAYER met2 ;
        RECT 27.405 2.705 27.745 3.055 ;
        RECT 27.395 5.84 27.735 6.19 ;
        RECT 27.48 2.705 27.65 6.19 ;
      LAYER met1 ;
        RECT 27.405 2.765 27.88 2.935 ;
        RECT 27.405 2.705 27.745 3.055 ;
        RECT 21.805 5.945 27.88 6.115 ;
        RECT 27.395 5.84 27.735 6.19 ;
        RECT 21.805 5.915 22.095 6.145 ;
      LAYER via1 ;
        RECT 27.495 5.94 27.645 6.09 ;
        RECT 27.505 2.805 27.655 2.955 ;
      LAYER mcon ;
        RECT 21.865 5.945 22.035 6.115 ;
        RECT 27.48 5.945 27.65 6.115 ;
        RECT 27.48 2.765 27.65 2.935 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 43.805 1.66 43.975 2.935 ;
        RECT 43.805 5.945 43.975 7.22 ;
        RECT 38.19 5.945 38.36 7.22 ;
      LAYER met2 ;
        RECT 43.73 2.705 44.07 3.055 ;
        RECT 43.72 5.84 44.06 6.19 ;
        RECT 43.805 2.705 43.975 6.19 ;
      LAYER met1 ;
        RECT 43.73 2.765 44.205 2.935 ;
        RECT 43.73 2.705 44.07 3.055 ;
        RECT 38.13 5.945 44.205 6.115 ;
        RECT 43.72 5.84 44.06 6.19 ;
        RECT 38.13 5.915 38.42 6.145 ;
      LAYER via1 ;
        RECT 43.82 5.94 43.97 6.09 ;
        RECT 43.83 2.805 43.98 2.955 ;
      LAYER mcon ;
        RECT 38.19 5.945 38.36 6.115 ;
        RECT 43.805 5.945 43.975 6.115 ;
        RECT 43.805 2.765 43.975 2.935 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 60.13 1.66 60.3 2.935 ;
        RECT 60.13 5.945 60.3 7.22 ;
        RECT 54.515 5.945 54.685 7.22 ;
      LAYER met2 ;
        RECT 60.055 2.705 60.395 3.055 ;
        RECT 60.045 5.84 60.385 6.19 ;
        RECT 60.13 2.705 60.3 6.19 ;
      LAYER met1 ;
        RECT 60.055 2.765 60.53 2.935 ;
        RECT 60.055 2.705 60.395 3.055 ;
        RECT 54.455 5.945 60.53 6.115 ;
        RECT 60.045 5.84 60.385 6.19 ;
        RECT 54.455 5.915 54.745 6.145 ;
      LAYER via1 ;
        RECT 60.145 5.94 60.295 6.09 ;
        RECT 60.155 2.805 60.305 2.955 ;
      LAYER mcon ;
        RECT 54.515 5.945 54.685 6.115 ;
        RECT 60.13 5.945 60.3 6.115 ;
        RECT 60.13 2.765 60.3 2.935 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 76.455 1.66 76.625 2.935 ;
        RECT 76.455 5.945 76.625 7.22 ;
        RECT 70.84 5.945 71.01 7.22 ;
      LAYER met2 ;
        RECT 76.38 2.705 76.72 3.055 ;
        RECT 76.37 5.84 76.71 6.19 ;
        RECT 76.455 2.705 76.625 6.19 ;
      LAYER met1 ;
        RECT 76.38 2.765 76.855 2.935 ;
        RECT 76.38 2.705 76.72 3.055 ;
        RECT 70.78 5.945 76.855 6.115 ;
        RECT 76.37 5.84 76.71 6.19 ;
        RECT 70.78 5.915 71.07 6.145 ;
      LAYER via1 ;
        RECT 76.47 5.94 76.62 6.09 ;
        RECT 76.48 2.805 76.63 2.955 ;
      LAYER mcon ;
        RECT 70.84 5.945 71.01 6.115 ;
        RECT 76.455 5.945 76.625 6.115 ;
        RECT 76.455 2.765 76.625 2.935 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT -3.04 5.945 -2.87 7.22 ;
      LAYER met1 ;
        RECT -3.1 5.945 -2.64 6.115 ;
        RECT -3.1 5.915 -2.81 6.145 ;
      LAYER mcon ;
        RECT -3.04 5.945 -2.87 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT -3.27 4.135 81.15 4.745 ;
        RECT 79.015 4.13 80.995 4.75 ;
        RECT 80.175 3.4 80.345 5.48 ;
        RECT 79.185 3.4 79.355 5.48 ;
        RECT 76.445 3.405 76.615 5.475 ;
        RECT 74.655 3.635 74.825 4.745 ;
        RECT 73.695 3.635 73.865 4.745 ;
        RECT 71.255 3.635 71.425 4.745 ;
        RECT 70.83 4.135 71 5.475 ;
        RECT 70.255 3.635 70.425 4.745 ;
        RECT 69.295 3.635 69.465 4.745 ;
        RECT 66.855 3.635 67.025 4.745 ;
        RECT 62.69 4.13 64.67 4.75 ;
        RECT 63.85 3.4 64.02 5.48 ;
        RECT 62.86 3.4 63.03 5.48 ;
        RECT 60.12 3.405 60.29 5.475 ;
        RECT 58.33 3.635 58.5 4.745 ;
        RECT 57.37 3.635 57.54 4.745 ;
        RECT 54.93 3.635 55.1 4.745 ;
        RECT 54.505 4.135 54.675 5.475 ;
        RECT 53.93 3.635 54.1 4.745 ;
        RECT 52.97 3.635 53.14 4.745 ;
        RECT 50.53 3.635 50.7 4.745 ;
        RECT 46.365 4.13 48.345 4.75 ;
        RECT 47.525 3.4 47.695 5.48 ;
        RECT 46.535 3.4 46.705 5.48 ;
        RECT 43.795 3.405 43.965 5.475 ;
        RECT 42.005 3.635 42.175 4.745 ;
        RECT 41.045 3.635 41.215 4.745 ;
        RECT 38.605 3.635 38.775 4.745 ;
        RECT 38.18 4.135 38.35 5.475 ;
        RECT 37.605 3.635 37.775 4.745 ;
        RECT 36.645 3.635 36.815 4.745 ;
        RECT 34.205 3.635 34.375 4.745 ;
        RECT 30.04 4.13 32.02 4.75 ;
        RECT 31.2 3.4 31.37 5.48 ;
        RECT 30.21 3.4 30.38 5.48 ;
        RECT 27.47 3.405 27.64 5.475 ;
        RECT 25.68 3.635 25.85 4.745 ;
        RECT 24.72 3.635 24.89 4.745 ;
        RECT 22.28 3.635 22.45 4.745 ;
        RECT 21.855 4.135 22.025 5.475 ;
        RECT 21.28 3.635 21.45 4.745 ;
        RECT 20.32 3.635 20.49 4.745 ;
        RECT 17.88 3.635 18.05 4.745 ;
        RECT 13.715 4.13 15.695 4.75 ;
        RECT 14.875 3.4 15.045 5.48 ;
        RECT 13.885 3.4 14.055 5.48 ;
        RECT 11.145 3.405 11.315 5.475 ;
        RECT 9.355 3.635 9.525 4.745 ;
        RECT 8.395 3.635 8.565 4.745 ;
        RECT 5.955 3.635 6.125 4.745 ;
        RECT 5.53 4.135 5.7 5.475 ;
        RECT 4.955 3.635 5.125 4.745 ;
        RECT 3.995 3.635 4.165 4.745 ;
        RECT 1.555 3.635 1.725 4.745 ;
        RECT -1.24 4.135 -1.07 8.305 ;
        RECT -3.05 4.135 -2.88 5.475 ;
      LAYER met1 ;
        RECT -3.27 4.135 81.15 4.745 ;
        RECT 79.015 4.13 80.995 4.75 ;
        RECT 65.565 3.98 75.225 4.745 ;
        RECT 62.69 4.13 64.67 4.75 ;
        RECT 49.24 3.98 58.9 4.745 ;
        RECT 46.365 4.13 48.345 4.75 ;
        RECT 32.915 3.98 42.575 4.745 ;
        RECT 30.04 4.13 32.02 4.75 ;
        RECT 16.59 3.98 26.25 4.745 ;
        RECT 13.715 4.13 15.695 4.75 ;
        RECT 0.265 3.98 9.925 4.745 ;
        RECT -1.3 6.655 -1.01 6.885 ;
        RECT -1.47 6.685 -1.01 6.855 ;
      LAYER mcon ;
        RECT -1.24 6.685 -1.07 6.855 ;
        RECT -0.93 4.545 -0.76 4.715 ;
        RECT 0.41 4.135 0.58 4.305 ;
        RECT 0.87 4.135 1.04 4.305 ;
        RECT 1.33 4.135 1.5 4.305 ;
        RECT 1.79 4.135 1.96 4.305 ;
        RECT 2.25 4.135 2.42 4.305 ;
        RECT 2.71 4.135 2.88 4.305 ;
        RECT 3.17 4.135 3.34 4.305 ;
        RECT 3.63 4.135 3.8 4.305 ;
        RECT 4.09 4.135 4.26 4.305 ;
        RECT 4.55 4.135 4.72 4.305 ;
        RECT 5.01 4.135 5.18 4.305 ;
        RECT 5.47 4.135 5.64 4.305 ;
        RECT 5.93 4.135 6.1 4.305 ;
        RECT 6.39 4.135 6.56 4.305 ;
        RECT 6.85 4.135 7.02 4.305 ;
        RECT 7.31 4.135 7.48 4.305 ;
        RECT 7.65 4.545 7.82 4.715 ;
        RECT 7.77 4.135 7.94 4.305 ;
        RECT 8.23 4.135 8.4 4.305 ;
        RECT 8.69 4.135 8.86 4.305 ;
        RECT 9.15 4.135 9.32 4.305 ;
        RECT 9.61 4.135 9.78 4.305 ;
        RECT 13.265 4.545 13.435 4.715 ;
        RECT 13.265 4.165 13.435 4.335 ;
        RECT 13.965 4.55 14.135 4.72 ;
        RECT 13.965 4.16 14.135 4.33 ;
        RECT 14.955 4.55 15.125 4.72 ;
        RECT 14.955 4.16 15.125 4.33 ;
        RECT 16.735 4.135 16.905 4.305 ;
        RECT 17.195 4.135 17.365 4.305 ;
        RECT 17.655 4.135 17.825 4.305 ;
        RECT 18.115 4.135 18.285 4.305 ;
        RECT 18.575 4.135 18.745 4.305 ;
        RECT 19.035 4.135 19.205 4.305 ;
        RECT 19.495 4.135 19.665 4.305 ;
        RECT 19.955 4.135 20.125 4.305 ;
        RECT 20.415 4.135 20.585 4.305 ;
        RECT 20.875 4.135 21.045 4.305 ;
        RECT 21.335 4.135 21.505 4.305 ;
        RECT 21.795 4.135 21.965 4.305 ;
        RECT 22.255 4.135 22.425 4.305 ;
        RECT 22.715 4.135 22.885 4.305 ;
        RECT 23.175 4.135 23.345 4.305 ;
        RECT 23.635 4.135 23.805 4.305 ;
        RECT 23.975 4.545 24.145 4.715 ;
        RECT 24.095 4.135 24.265 4.305 ;
        RECT 24.555 4.135 24.725 4.305 ;
        RECT 25.015 4.135 25.185 4.305 ;
        RECT 25.475 4.135 25.645 4.305 ;
        RECT 25.935 4.135 26.105 4.305 ;
        RECT 29.59 4.545 29.76 4.715 ;
        RECT 29.59 4.165 29.76 4.335 ;
        RECT 30.29 4.55 30.46 4.72 ;
        RECT 30.29 4.16 30.46 4.33 ;
        RECT 31.28 4.55 31.45 4.72 ;
        RECT 31.28 4.16 31.45 4.33 ;
        RECT 33.06 4.135 33.23 4.305 ;
        RECT 33.52 4.135 33.69 4.305 ;
        RECT 33.98 4.135 34.15 4.305 ;
        RECT 34.44 4.135 34.61 4.305 ;
        RECT 34.9 4.135 35.07 4.305 ;
        RECT 35.36 4.135 35.53 4.305 ;
        RECT 35.82 4.135 35.99 4.305 ;
        RECT 36.28 4.135 36.45 4.305 ;
        RECT 36.74 4.135 36.91 4.305 ;
        RECT 37.2 4.135 37.37 4.305 ;
        RECT 37.66 4.135 37.83 4.305 ;
        RECT 38.12 4.135 38.29 4.305 ;
        RECT 38.58 4.135 38.75 4.305 ;
        RECT 39.04 4.135 39.21 4.305 ;
        RECT 39.5 4.135 39.67 4.305 ;
        RECT 39.96 4.135 40.13 4.305 ;
        RECT 40.3 4.545 40.47 4.715 ;
        RECT 40.42 4.135 40.59 4.305 ;
        RECT 40.88 4.135 41.05 4.305 ;
        RECT 41.34 4.135 41.51 4.305 ;
        RECT 41.8 4.135 41.97 4.305 ;
        RECT 42.26 4.135 42.43 4.305 ;
        RECT 45.915 4.545 46.085 4.715 ;
        RECT 45.915 4.165 46.085 4.335 ;
        RECT 46.615 4.55 46.785 4.72 ;
        RECT 46.615 4.16 46.785 4.33 ;
        RECT 47.605 4.55 47.775 4.72 ;
        RECT 47.605 4.16 47.775 4.33 ;
        RECT 49.385 4.135 49.555 4.305 ;
        RECT 49.845 4.135 50.015 4.305 ;
        RECT 50.305 4.135 50.475 4.305 ;
        RECT 50.765 4.135 50.935 4.305 ;
        RECT 51.225 4.135 51.395 4.305 ;
        RECT 51.685 4.135 51.855 4.305 ;
        RECT 52.145 4.135 52.315 4.305 ;
        RECT 52.605 4.135 52.775 4.305 ;
        RECT 53.065 4.135 53.235 4.305 ;
        RECT 53.525 4.135 53.695 4.305 ;
        RECT 53.985 4.135 54.155 4.305 ;
        RECT 54.445 4.135 54.615 4.305 ;
        RECT 54.905 4.135 55.075 4.305 ;
        RECT 55.365 4.135 55.535 4.305 ;
        RECT 55.825 4.135 55.995 4.305 ;
        RECT 56.285 4.135 56.455 4.305 ;
        RECT 56.625 4.545 56.795 4.715 ;
        RECT 56.745 4.135 56.915 4.305 ;
        RECT 57.205 4.135 57.375 4.305 ;
        RECT 57.665 4.135 57.835 4.305 ;
        RECT 58.125 4.135 58.295 4.305 ;
        RECT 58.585 4.135 58.755 4.305 ;
        RECT 62.24 4.545 62.41 4.715 ;
        RECT 62.24 4.165 62.41 4.335 ;
        RECT 62.94 4.55 63.11 4.72 ;
        RECT 62.94 4.16 63.11 4.33 ;
        RECT 63.93 4.55 64.1 4.72 ;
        RECT 63.93 4.16 64.1 4.33 ;
        RECT 65.71 4.135 65.88 4.305 ;
        RECT 66.17 4.135 66.34 4.305 ;
        RECT 66.63 4.135 66.8 4.305 ;
        RECT 67.09 4.135 67.26 4.305 ;
        RECT 67.55 4.135 67.72 4.305 ;
        RECT 68.01 4.135 68.18 4.305 ;
        RECT 68.47 4.135 68.64 4.305 ;
        RECT 68.93 4.135 69.1 4.305 ;
        RECT 69.39 4.135 69.56 4.305 ;
        RECT 69.85 4.135 70.02 4.305 ;
        RECT 70.31 4.135 70.48 4.305 ;
        RECT 70.77 4.135 70.94 4.305 ;
        RECT 71.23 4.135 71.4 4.305 ;
        RECT 71.69 4.135 71.86 4.305 ;
        RECT 72.15 4.135 72.32 4.305 ;
        RECT 72.61 4.135 72.78 4.305 ;
        RECT 72.95 4.545 73.12 4.715 ;
        RECT 73.07 4.135 73.24 4.305 ;
        RECT 73.53 4.135 73.7 4.305 ;
        RECT 73.99 4.135 74.16 4.305 ;
        RECT 74.45 4.135 74.62 4.305 ;
        RECT 74.91 4.135 75.08 4.305 ;
        RECT 78.565 4.545 78.735 4.715 ;
        RECT 78.565 4.165 78.735 4.335 ;
        RECT 79.265 4.55 79.435 4.72 ;
        RECT 79.265 4.16 79.435 4.33 ;
        RECT 80.255 4.55 80.425 4.72 ;
        RECT 80.255 4.16 80.425 4.33 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 74.455 2.975 74.785 3.705 ;
        RECT 58.13 2.975 58.46 3.705 ;
        RECT 41.805 2.975 42.135 3.705 ;
        RECT 25.48 2.975 25.81 3.705 ;
        RECT 9.155 2.975 9.485 3.705 ;
      LAYER li1 ;
        RECT 80.97 0 81.15 0.305 ;
        RECT -3.27 0 81.15 0.3 ;
        RECT 80.175 0 80.345 0.93 ;
        RECT 79.185 0 79.355 0.93 ;
        RECT 64.645 0 79.02 0.305 ;
        RECT 76.445 0 76.615 0.935 ;
        RECT 65.565 0 75.38 1.585 ;
        RECT 73.695 0 73.865 2.085 ;
        RECT 71.735 0 71.905 2.085 ;
        RECT 71.665 0 71.905 1.595 ;
        RECT 70.115 0 70.31 1.595 ;
        RECT 69.295 0 69.465 2.085 ;
        RECT 68.335 0 68.505 2.085 ;
        RECT 67.99 0 68.185 1.595 ;
        RECT 67.815 0 67.985 2.085 ;
        RECT 66.855 0 67.025 2.085 ;
        RECT 65.895 0 66.065 2.085 ;
        RECT 65.69 0 65.885 1.595 ;
        RECT 63.85 0 64.02 0.93 ;
        RECT 62.86 0 63.03 0.93 ;
        RECT 48.32 0 62.695 0.305 ;
        RECT 60.12 0 60.29 0.935 ;
        RECT 49.24 0 59.055 1.585 ;
        RECT 57.37 0 57.54 2.085 ;
        RECT 55.41 0 55.58 2.085 ;
        RECT 55.34 0 55.58 1.595 ;
        RECT 53.79 0 53.985 1.595 ;
        RECT 52.97 0 53.14 2.085 ;
        RECT 52.01 0 52.18 2.085 ;
        RECT 51.665 0 51.86 1.595 ;
        RECT 51.49 0 51.66 2.085 ;
        RECT 50.53 0 50.7 2.085 ;
        RECT 49.57 0 49.74 2.085 ;
        RECT 49.365 0 49.56 1.595 ;
        RECT 47.525 0 47.695 0.93 ;
        RECT 46.535 0 46.705 0.93 ;
        RECT 31.995 0 46.37 0.305 ;
        RECT 43.795 0 43.965 0.935 ;
        RECT 32.915 0 42.73 1.585 ;
        RECT 41.045 0 41.215 2.085 ;
        RECT 39.085 0 39.255 2.085 ;
        RECT 39.015 0 39.255 1.595 ;
        RECT 37.465 0 37.66 1.595 ;
        RECT 36.645 0 36.815 2.085 ;
        RECT 35.685 0 35.855 2.085 ;
        RECT 35.34 0 35.535 1.595 ;
        RECT 35.165 0 35.335 2.085 ;
        RECT 34.205 0 34.375 2.085 ;
        RECT 33.245 0 33.415 2.085 ;
        RECT 33.04 0 33.235 1.595 ;
        RECT 31.2 0 31.37 0.93 ;
        RECT 30.21 0 30.38 0.93 ;
        RECT 15.67 0 30.045 0.305 ;
        RECT 27.47 0 27.64 0.935 ;
        RECT 16.59 0 26.405 1.585 ;
        RECT 24.72 0 24.89 2.085 ;
        RECT 22.76 0 22.93 2.085 ;
        RECT 22.69 0 22.93 1.595 ;
        RECT 21.14 0 21.335 1.595 ;
        RECT 20.32 0 20.49 2.085 ;
        RECT 19.36 0 19.53 2.085 ;
        RECT 19.015 0 19.21 1.595 ;
        RECT 18.84 0 19.01 2.085 ;
        RECT 17.88 0 18.05 2.085 ;
        RECT 16.92 0 17.09 2.085 ;
        RECT 16.715 0 16.91 1.595 ;
        RECT 14.875 0 15.045 0.93 ;
        RECT 13.885 0 14.055 0.93 ;
        RECT -3.27 0 13.72 0.305 ;
        RECT 11.145 0 11.315 0.935 ;
        RECT 0.265 0 10.08 1.585 ;
        RECT 8.395 0 8.565 2.085 ;
        RECT 6.435 0 6.605 2.085 ;
        RECT 6.365 0 6.605 1.595 ;
        RECT 4.815 0 5.01 1.595 ;
        RECT 3.995 0 4.165 2.085 ;
        RECT 3.035 0 3.205 2.085 ;
        RECT 2.69 0 2.885 1.595 ;
        RECT 2.515 0 2.685 2.085 ;
        RECT 1.555 0 1.725 2.085 ;
        RECT 0.595 0 0.765 2.085 ;
        RECT 0.39 0 0.585 1.595 ;
        RECT -3.27 8.58 81.15 8.88 ;
        RECT 80.97 8.575 81.15 8.88 ;
        RECT 80.175 7.95 80.345 8.88 ;
        RECT 79.185 7.95 79.355 8.88 ;
        RECT 64.645 8.575 79.02 8.88 ;
        RECT 76.445 7.945 76.615 8.88 ;
        RECT 70.83 7.945 71 8.88 ;
        RECT 63.85 7.95 64.02 8.88 ;
        RECT 62.86 7.95 63.03 8.88 ;
        RECT 48.32 8.575 62.695 8.88 ;
        RECT 60.12 7.945 60.29 8.88 ;
        RECT 54.505 7.945 54.675 8.88 ;
        RECT 47.525 7.95 47.695 8.88 ;
        RECT 46.535 7.95 46.705 8.88 ;
        RECT 31.995 8.575 46.37 8.88 ;
        RECT 43.795 7.945 43.965 8.88 ;
        RECT 38.18 7.945 38.35 8.88 ;
        RECT 31.2 7.95 31.37 8.88 ;
        RECT 30.21 7.95 30.38 8.88 ;
        RECT 15.67 8.575 30.045 8.88 ;
        RECT 27.47 7.945 27.64 8.88 ;
        RECT 21.855 7.945 22.025 8.88 ;
        RECT 14.875 7.95 15.045 8.88 ;
        RECT 13.885 7.95 14.055 8.88 ;
        RECT -3.27 8.575 13.72 8.88 ;
        RECT 11.145 7.945 11.315 8.88 ;
        RECT 5.53 7.945 5.7 8.88 ;
        RECT -3.05 7.945 -2.88 8.88 ;
        RECT 74.655 2.575 74.825 2.945 ;
        RECT 74.335 2.575 74.825 2.745 ;
        RECT 72.695 2.575 72.865 2.945 ;
        RECT 72.375 2.575 72.865 2.745 ;
        RECT 71.835 6.075 72.005 8.025 ;
        RECT 71.78 7.855 71.95 8.305 ;
        RECT 71.78 5.015 71.95 6.245 ;
        RECT 58.33 2.575 58.5 2.945 ;
        RECT 58.01 2.575 58.5 2.745 ;
        RECT 56.37 2.575 56.54 2.945 ;
        RECT 56.05 2.575 56.54 2.745 ;
        RECT 55.51 6.075 55.68 8.025 ;
        RECT 55.455 7.855 55.625 8.305 ;
        RECT 55.455 5.015 55.625 6.245 ;
        RECT 42.005 2.575 42.175 2.945 ;
        RECT 41.685 2.575 42.175 2.745 ;
        RECT 40.045 2.575 40.215 2.945 ;
        RECT 39.725 2.575 40.215 2.745 ;
        RECT 39.185 6.075 39.355 8.025 ;
        RECT 39.13 7.855 39.3 8.305 ;
        RECT 39.13 5.015 39.3 6.245 ;
        RECT 25.68 2.575 25.85 2.945 ;
        RECT 25.36 2.575 25.85 2.745 ;
        RECT 23.72 2.575 23.89 2.945 ;
        RECT 23.4 2.575 23.89 2.745 ;
        RECT 22.86 6.075 23.03 8.025 ;
        RECT 22.805 7.855 22.975 8.305 ;
        RECT 22.805 5.015 22.975 6.245 ;
        RECT 9.355 2.575 9.525 2.945 ;
        RECT 9.035 2.575 9.525 2.745 ;
        RECT 7.395 2.575 7.565 2.945 ;
        RECT 7.075 2.575 7.565 2.745 ;
        RECT 6.535 6.075 6.705 8.025 ;
        RECT 6.48 7.855 6.65 8.305 ;
        RECT 6.48 5.015 6.65 6.245 ;
      LAYER met2 ;
        RECT 74.48 2.955 74.76 3.325 ;
        RECT 74.49 2.7 74.75 3.325 ;
        RECT 58.155 2.955 58.435 3.325 ;
        RECT 58.165 2.7 58.425 3.325 ;
        RECT 41.83 2.955 42.11 3.325 ;
        RECT 41.84 2.7 42.1 3.325 ;
        RECT 25.505 2.955 25.785 3.325 ;
        RECT 25.515 2.7 25.775 3.325 ;
        RECT 9.18 2.955 9.46 3.325 ;
        RECT 9.19 2.7 9.45 3.325 ;
      LAYER met1 ;
        RECT 80.97 0 81.15 0.305 ;
        RECT -3.27 0 81.15 0.3 ;
        RECT 64.645 0 79.02 0.305 ;
        RECT 75.195 0 75.38 2.945 ;
        RECT 74.43 2.79 75.38 2.945 ;
        RECT 74.46 2.76 75.38 2.945 ;
        RECT 65.565 0 75.38 1.74 ;
        RECT 74.46 2.745 74.885 2.975 ;
        RECT 74.46 2.73 74.78 2.99 ;
        RECT 72.97 2.93 74.735 3.055 ;
        RECT 72.97 2.93 74.57 3.07 ;
        RECT 72.635 2.79 73.11 2.975 ;
        RECT 72.635 2.745 72.925 2.975 ;
        RECT 48.32 0 62.695 0.305 ;
        RECT 58.87 0 59.055 2.945 ;
        RECT 58.105 2.79 59.055 2.945 ;
        RECT 58.135 2.76 59.055 2.945 ;
        RECT 49.24 0 59.055 1.74 ;
        RECT 58.135 2.745 58.56 2.975 ;
        RECT 58.135 2.73 58.455 2.99 ;
        RECT 56.645 2.93 58.41 3.055 ;
        RECT 56.645 2.93 58.245 3.07 ;
        RECT 56.31 2.79 56.785 2.975 ;
        RECT 56.31 2.745 56.6 2.975 ;
        RECT 31.995 0 46.37 0.305 ;
        RECT 42.545 0 42.73 2.945 ;
        RECT 41.78 2.79 42.73 2.945 ;
        RECT 41.81 2.76 42.73 2.945 ;
        RECT 32.915 0 42.73 1.74 ;
        RECT 41.81 2.745 42.235 2.975 ;
        RECT 41.81 2.73 42.13 2.99 ;
        RECT 40.32 2.93 42.085 3.055 ;
        RECT 40.32 2.93 41.92 3.07 ;
        RECT 39.985 2.79 40.46 2.975 ;
        RECT 39.985 2.745 40.275 2.975 ;
        RECT 15.67 0 30.045 0.305 ;
        RECT 26.22 0 26.405 2.945 ;
        RECT 25.455 2.79 26.405 2.945 ;
        RECT 25.485 2.76 26.405 2.945 ;
        RECT 16.59 0 26.405 1.74 ;
        RECT 25.485 2.745 25.91 2.975 ;
        RECT 25.485 2.73 25.805 2.99 ;
        RECT 23.995 2.93 25.76 3.055 ;
        RECT 23.995 2.93 25.595 3.07 ;
        RECT 23.66 2.79 24.135 2.975 ;
        RECT 23.66 2.745 23.95 2.975 ;
        RECT -3.27 0 13.72 0.305 ;
        RECT 9.895 0 10.08 2.945 ;
        RECT 9.13 2.79 10.08 2.945 ;
        RECT 9.16 2.76 10.08 2.945 ;
        RECT 0.265 0 10.08 1.74 ;
        RECT 9.16 2.745 9.585 2.975 ;
        RECT 9.16 2.73 9.48 2.99 ;
        RECT 7.67 2.93 9.435 3.055 ;
        RECT 7.67 2.93 9.27 3.07 ;
        RECT 7.335 2.79 7.81 2.975 ;
        RECT 7.335 2.745 7.625 2.975 ;
        RECT -3.27 8.58 81.15 8.88 ;
        RECT 80.97 8.575 81.15 8.88 ;
        RECT 64.645 8.575 79.02 8.88 ;
        RECT 71.775 6.285 72.065 6.515 ;
        RECT 71.4 6.315 72.065 6.485 ;
        RECT 71.4 6.315 71.575 8.88 ;
        RECT 48.32 8.575 62.695 8.88 ;
        RECT 55.45 6.285 55.74 6.515 ;
        RECT 55.075 6.315 55.74 6.485 ;
        RECT 55.075 6.315 55.25 8.88 ;
        RECT 31.995 8.575 46.37 8.88 ;
        RECT 39.125 6.285 39.415 6.515 ;
        RECT 38.75 6.315 39.415 6.485 ;
        RECT 38.75 6.315 38.925 8.88 ;
        RECT 15.67 8.575 30.045 8.88 ;
        RECT 22.8 6.285 23.09 6.515 ;
        RECT 22.425 6.315 23.09 6.485 ;
        RECT 22.425 6.315 22.6 8.88 ;
        RECT -3.27 8.575 13.72 8.88 ;
        RECT 6.475 6.285 6.765 6.515 ;
        RECT 6.1 6.315 6.765 6.485 ;
        RECT 6.1 6.315 6.275 8.88 ;
      LAYER via2 ;
        RECT 9.22 3.04 9.42 3.24 ;
        RECT 25.545 3.04 25.745 3.24 ;
        RECT 41.87 3.04 42.07 3.24 ;
        RECT 58.195 3.04 58.395 3.24 ;
        RECT 74.52 3.04 74.72 3.24 ;
      LAYER via1 ;
        RECT 9.245 2.785 9.395 2.935 ;
        RECT 25.57 2.785 25.72 2.935 ;
        RECT 41.895 2.785 42.045 2.935 ;
        RECT 58.22 2.785 58.37 2.935 ;
        RECT 74.545 2.785 74.695 2.935 ;
      LAYER mcon ;
        RECT -2.97 8.605 -2.8 8.775 ;
        RECT -2.29 8.605 -2.12 8.775 ;
        RECT -1.61 8.605 -1.44 8.775 ;
        RECT -0.93 8.605 -0.76 8.775 ;
        RECT 0.41 1.415 0.58 1.585 ;
        RECT 0.87 1.415 1.04 1.585 ;
        RECT 1.33 1.415 1.5 1.585 ;
        RECT 1.79 1.415 1.96 1.585 ;
        RECT 2.25 1.415 2.42 1.585 ;
        RECT 2.71 1.415 2.88 1.585 ;
        RECT 3.17 1.415 3.34 1.585 ;
        RECT 3.63 1.415 3.8 1.585 ;
        RECT 4.09 1.415 4.26 1.585 ;
        RECT 4.55 1.415 4.72 1.585 ;
        RECT 5.01 1.415 5.18 1.585 ;
        RECT 5.47 1.415 5.64 1.585 ;
        RECT 5.61 8.605 5.78 8.775 ;
        RECT 5.93 1.415 6.1 1.585 ;
        RECT 6.29 8.605 6.46 8.775 ;
        RECT 6.39 1.415 6.56 1.585 ;
        RECT 6.535 6.315 6.705 6.485 ;
        RECT 6.85 1.415 7.02 1.585 ;
        RECT 6.97 8.605 7.14 8.775 ;
        RECT 7.31 1.415 7.48 1.585 ;
        RECT 7.395 2.775 7.565 2.945 ;
        RECT 7.65 8.605 7.82 8.775 ;
        RECT 7.77 1.415 7.94 1.585 ;
        RECT 8.23 1.415 8.4 1.585 ;
        RECT 8.69 1.415 8.86 1.585 ;
        RECT 9.15 1.415 9.32 1.585 ;
        RECT 9.355 2.775 9.525 2.945 ;
        RECT 9.61 1.415 9.78 1.585 ;
        RECT 11.225 8.605 11.395 8.775 ;
        RECT 11.225 0.105 11.395 0.275 ;
        RECT 11.905 8.605 12.075 8.775 ;
        RECT 11.905 0.105 12.075 0.275 ;
        RECT 12.585 8.605 12.755 8.775 ;
        RECT 12.585 0.105 12.755 0.275 ;
        RECT 13.265 8.605 13.435 8.775 ;
        RECT 13.265 0.105 13.435 0.275 ;
        RECT 13.965 8.61 14.135 8.78 ;
        RECT 13.965 0.1 14.135 0.27 ;
        RECT 14.955 8.61 15.125 8.78 ;
        RECT 14.955 0.1 15.125 0.27 ;
        RECT 16.735 1.415 16.905 1.585 ;
        RECT 17.195 1.415 17.365 1.585 ;
        RECT 17.655 1.415 17.825 1.585 ;
        RECT 18.115 1.415 18.285 1.585 ;
        RECT 18.575 1.415 18.745 1.585 ;
        RECT 19.035 1.415 19.205 1.585 ;
        RECT 19.495 1.415 19.665 1.585 ;
        RECT 19.955 1.415 20.125 1.585 ;
        RECT 20.415 1.415 20.585 1.585 ;
        RECT 20.875 1.415 21.045 1.585 ;
        RECT 21.335 1.415 21.505 1.585 ;
        RECT 21.795 1.415 21.965 1.585 ;
        RECT 21.935 8.605 22.105 8.775 ;
        RECT 22.255 1.415 22.425 1.585 ;
        RECT 22.615 8.605 22.785 8.775 ;
        RECT 22.715 1.415 22.885 1.585 ;
        RECT 22.86 6.315 23.03 6.485 ;
        RECT 23.175 1.415 23.345 1.585 ;
        RECT 23.295 8.605 23.465 8.775 ;
        RECT 23.635 1.415 23.805 1.585 ;
        RECT 23.72 2.775 23.89 2.945 ;
        RECT 23.975 8.605 24.145 8.775 ;
        RECT 24.095 1.415 24.265 1.585 ;
        RECT 24.555 1.415 24.725 1.585 ;
        RECT 25.015 1.415 25.185 1.585 ;
        RECT 25.475 1.415 25.645 1.585 ;
        RECT 25.68 2.775 25.85 2.945 ;
        RECT 25.935 1.415 26.105 1.585 ;
        RECT 27.55 8.605 27.72 8.775 ;
        RECT 27.55 0.105 27.72 0.275 ;
        RECT 28.23 8.605 28.4 8.775 ;
        RECT 28.23 0.105 28.4 0.275 ;
        RECT 28.91 8.605 29.08 8.775 ;
        RECT 28.91 0.105 29.08 0.275 ;
        RECT 29.59 8.605 29.76 8.775 ;
        RECT 29.59 0.105 29.76 0.275 ;
        RECT 30.29 8.61 30.46 8.78 ;
        RECT 30.29 0.1 30.46 0.27 ;
        RECT 31.28 8.61 31.45 8.78 ;
        RECT 31.28 0.1 31.45 0.27 ;
        RECT 33.06 1.415 33.23 1.585 ;
        RECT 33.52 1.415 33.69 1.585 ;
        RECT 33.98 1.415 34.15 1.585 ;
        RECT 34.44 1.415 34.61 1.585 ;
        RECT 34.9 1.415 35.07 1.585 ;
        RECT 35.36 1.415 35.53 1.585 ;
        RECT 35.82 1.415 35.99 1.585 ;
        RECT 36.28 1.415 36.45 1.585 ;
        RECT 36.74 1.415 36.91 1.585 ;
        RECT 37.2 1.415 37.37 1.585 ;
        RECT 37.66 1.415 37.83 1.585 ;
        RECT 38.12 1.415 38.29 1.585 ;
        RECT 38.26 8.605 38.43 8.775 ;
        RECT 38.58 1.415 38.75 1.585 ;
        RECT 38.94 8.605 39.11 8.775 ;
        RECT 39.04 1.415 39.21 1.585 ;
        RECT 39.185 6.315 39.355 6.485 ;
        RECT 39.5 1.415 39.67 1.585 ;
        RECT 39.62 8.605 39.79 8.775 ;
        RECT 39.96 1.415 40.13 1.585 ;
        RECT 40.045 2.775 40.215 2.945 ;
        RECT 40.3 8.605 40.47 8.775 ;
        RECT 40.42 1.415 40.59 1.585 ;
        RECT 40.88 1.415 41.05 1.585 ;
        RECT 41.34 1.415 41.51 1.585 ;
        RECT 41.8 1.415 41.97 1.585 ;
        RECT 42.005 2.775 42.175 2.945 ;
        RECT 42.26 1.415 42.43 1.585 ;
        RECT 43.875 8.605 44.045 8.775 ;
        RECT 43.875 0.105 44.045 0.275 ;
        RECT 44.555 8.605 44.725 8.775 ;
        RECT 44.555 0.105 44.725 0.275 ;
        RECT 45.235 8.605 45.405 8.775 ;
        RECT 45.235 0.105 45.405 0.275 ;
        RECT 45.915 8.605 46.085 8.775 ;
        RECT 45.915 0.105 46.085 0.275 ;
        RECT 46.615 8.61 46.785 8.78 ;
        RECT 46.615 0.1 46.785 0.27 ;
        RECT 47.605 8.61 47.775 8.78 ;
        RECT 47.605 0.1 47.775 0.27 ;
        RECT 49.385 1.415 49.555 1.585 ;
        RECT 49.845 1.415 50.015 1.585 ;
        RECT 50.305 1.415 50.475 1.585 ;
        RECT 50.765 1.415 50.935 1.585 ;
        RECT 51.225 1.415 51.395 1.585 ;
        RECT 51.685 1.415 51.855 1.585 ;
        RECT 52.145 1.415 52.315 1.585 ;
        RECT 52.605 1.415 52.775 1.585 ;
        RECT 53.065 1.415 53.235 1.585 ;
        RECT 53.525 1.415 53.695 1.585 ;
        RECT 53.985 1.415 54.155 1.585 ;
        RECT 54.445 1.415 54.615 1.585 ;
        RECT 54.585 8.605 54.755 8.775 ;
        RECT 54.905 1.415 55.075 1.585 ;
        RECT 55.265 8.605 55.435 8.775 ;
        RECT 55.365 1.415 55.535 1.585 ;
        RECT 55.51 6.315 55.68 6.485 ;
        RECT 55.825 1.415 55.995 1.585 ;
        RECT 55.945 8.605 56.115 8.775 ;
        RECT 56.285 1.415 56.455 1.585 ;
        RECT 56.37 2.775 56.54 2.945 ;
        RECT 56.625 8.605 56.795 8.775 ;
        RECT 56.745 1.415 56.915 1.585 ;
        RECT 57.205 1.415 57.375 1.585 ;
        RECT 57.665 1.415 57.835 1.585 ;
        RECT 58.125 1.415 58.295 1.585 ;
        RECT 58.33 2.775 58.5 2.945 ;
        RECT 58.585 1.415 58.755 1.585 ;
        RECT 60.2 8.605 60.37 8.775 ;
        RECT 60.2 0.105 60.37 0.275 ;
        RECT 60.88 8.605 61.05 8.775 ;
        RECT 60.88 0.105 61.05 0.275 ;
        RECT 61.56 8.605 61.73 8.775 ;
        RECT 61.56 0.105 61.73 0.275 ;
        RECT 62.24 8.605 62.41 8.775 ;
        RECT 62.24 0.105 62.41 0.275 ;
        RECT 62.94 8.61 63.11 8.78 ;
        RECT 62.94 0.1 63.11 0.27 ;
        RECT 63.93 8.61 64.1 8.78 ;
        RECT 63.93 0.1 64.1 0.27 ;
        RECT 65.71 1.415 65.88 1.585 ;
        RECT 66.17 1.415 66.34 1.585 ;
        RECT 66.63 1.415 66.8 1.585 ;
        RECT 67.09 1.415 67.26 1.585 ;
        RECT 67.55 1.415 67.72 1.585 ;
        RECT 68.01 1.415 68.18 1.585 ;
        RECT 68.47 1.415 68.64 1.585 ;
        RECT 68.93 1.415 69.1 1.585 ;
        RECT 69.39 1.415 69.56 1.585 ;
        RECT 69.85 1.415 70.02 1.585 ;
        RECT 70.31 1.415 70.48 1.585 ;
        RECT 70.77 1.415 70.94 1.585 ;
        RECT 70.91 8.605 71.08 8.775 ;
        RECT 71.23 1.415 71.4 1.585 ;
        RECT 71.59 8.605 71.76 8.775 ;
        RECT 71.69 1.415 71.86 1.585 ;
        RECT 71.835 6.315 72.005 6.485 ;
        RECT 72.15 1.415 72.32 1.585 ;
        RECT 72.27 8.605 72.44 8.775 ;
        RECT 72.61 1.415 72.78 1.585 ;
        RECT 72.695 2.775 72.865 2.945 ;
        RECT 72.95 8.605 73.12 8.775 ;
        RECT 73.07 1.415 73.24 1.585 ;
        RECT 73.53 1.415 73.7 1.585 ;
        RECT 73.99 1.415 74.16 1.585 ;
        RECT 74.45 1.415 74.62 1.585 ;
        RECT 74.655 2.775 74.825 2.945 ;
        RECT 74.91 1.415 75.08 1.585 ;
        RECT 76.525 8.605 76.695 8.775 ;
        RECT 76.525 0.105 76.695 0.275 ;
        RECT 77.205 8.605 77.375 8.775 ;
        RECT 77.205 0.105 77.375 0.275 ;
        RECT 77.885 8.605 78.055 8.775 ;
        RECT 77.885 0.105 78.055 0.275 ;
        RECT 78.565 8.605 78.735 8.775 ;
        RECT 78.565 0.105 78.735 0.275 ;
        RECT 79.265 8.61 79.435 8.78 ;
        RECT 79.265 0.1 79.435 0.27 ;
        RECT 80.255 8.61 80.425 8.78 ;
        RECT 80.255 0.1 80.425 0.27 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 72.13 7.055 72.5 7.425 ;
      RECT 72.13 7.09 74.115 7.39 ;
      RECT 73.815 2.28 74.115 7.39 ;
      RECT 70.815 2.015 71.145 2.745 ;
      RECT 69.935 2.015 70.265 2.745 ;
      RECT 73.015 2.28 74.305 2.58 ;
      RECT 73.975 1.85 74.305 2.58 ;
      RECT 69.935 2.28 72.075 2.58 ;
      RECT 71.775 1.965 72.075 2.58 ;
      RECT 73.015 1.98 73.32 2.58 ;
      RECT 71.775 1.965 73.135 2.275 ;
      RECT 70.435 3.535 70.765 3.865 ;
      RECT 69.23 3.55 70.765 3.85 ;
      RECT 69.23 2.43 69.53 3.85 ;
      RECT 68.975 2.415 69.305 2.745 ;
      RECT 55.805 7.055 56.175 7.425 ;
      RECT 55.805 7.09 57.79 7.39 ;
      RECT 57.49 2.28 57.79 7.39 ;
      RECT 54.49 2.015 54.82 2.745 ;
      RECT 53.61 2.015 53.94 2.745 ;
      RECT 56.69 2.28 57.98 2.58 ;
      RECT 57.65 1.85 57.98 2.58 ;
      RECT 53.61 2.28 55.75 2.58 ;
      RECT 55.45 1.965 55.75 2.58 ;
      RECT 56.69 1.98 56.995 2.58 ;
      RECT 55.45 1.965 56.81 2.275 ;
      RECT 54.11 3.535 54.44 3.865 ;
      RECT 52.905 3.55 54.44 3.85 ;
      RECT 52.905 2.43 53.205 3.85 ;
      RECT 52.65 2.415 52.98 2.745 ;
      RECT 39.48 7.055 39.85 7.425 ;
      RECT 39.48 7.09 41.465 7.39 ;
      RECT 41.165 2.28 41.465 7.39 ;
      RECT 38.165 2.015 38.495 2.745 ;
      RECT 37.285 2.015 37.615 2.745 ;
      RECT 40.365 2.28 41.655 2.58 ;
      RECT 41.325 1.85 41.655 2.58 ;
      RECT 37.285 2.28 39.425 2.58 ;
      RECT 39.125 1.965 39.425 2.58 ;
      RECT 40.365 1.98 40.67 2.58 ;
      RECT 39.125 1.965 40.485 2.275 ;
      RECT 37.785 3.535 38.115 3.865 ;
      RECT 36.58 3.55 38.115 3.85 ;
      RECT 36.58 2.43 36.88 3.85 ;
      RECT 36.325 2.415 36.655 2.745 ;
      RECT 23.155 7.055 23.525 7.425 ;
      RECT 23.155 7.09 25.14 7.39 ;
      RECT 24.84 2.28 25.14 7.39 ;
      RECT 21.84 2.015 22.17 2.745 ;
      RECT 20.96 2.015 21.29 2.745 ;
      RECT 24.04 2.28 25.33 2.58 ;
      RECT 25 1.85 25.33 2.58 ;
      RECT 20.96 2.28 23.1 2.58 ;
      RECT 22.8 1.965 23.1 2.58 ;
      RECT 24.04 1.98 24.345 2.58 ;
      RECT 22.8 1.965 24.16 2.275 ;
      RECT 21.46 3.535 21.79 3.865 ;
      RECT 20.255 3.55 21.79 3.85 ;
      RECT 20.255 2.43 20.555 3.85 ;
      RECT 20 2.415 20.33 2.745 ;
      RECT 6.83 7.055 7.2 7.425 ;
      RECT 6.83 7.09 8.815 7.39 ;
      RECT 8.515 2.28 8.815 7.39 ;
      RECT 5.515 2.015 5.845 2.745 ;
      RECT 4.635 2.015 4.965 2.745 ;
      RECT 7.715 2.28 9.005 2.58 ;
      RECT 8.675 1.85 9.005 2.58 ;
      RECT 4.635 2.28 6.775 2.58 ;
      RECT 6.475 1.965 6.775 2.58 ;
      RECT 7.715 1.98 8.02 2.58 ;
      RECT 6.475 1.965 7.835 2.275 ;
      RECT 5.135 3.535 5.465 3.865 ;
      RECT 3.93 3.55 5.465 3.85 ;
      RECT 3.93 2.43 4.23 3.85 ;
      RECT 3.675 2.415 4.005 2.745 ;
      RECT 72.375 2.575 72.705 3.305 ;
      RECT 68.255 2.415 68.585 3.145 ;
      RECT 67.255 1.855 67.585 2.585 ;
      RECT 65.815 2.575 66.145 3.305 ;
      RECT 56.05 2.575 56.38 3.305 ;
      RECT 51.93 2.415 52.26 3.145 ;
      RECT 50.93 1.855 51.26 2.585 ;
      RECT 49.49 2.575 49.82 3.305 ;
      RECT 39.725 2.575 40.055 3.305 ;
      RECT 35.605 2.415 35.935 3.145 ;
      RECT 34.605 1.855 34.935 2.585 ;
      RECT 33.165 2.575 33.495 3.305 ;
      RECT 23.4 2.575 23.73 3.305 ;
      RECT 19.28 2.415 19.61 3.145 ;
      RECT 18.28 1.855 18.61 2.585 ;
      RECT 16.84 2.575 17.17 3.305 ;
      RECT 7.075 2.575 7.405 3.305 ;
      RECT 2.955 2.415 3.285 3.145 ;
      RECT 1.955 1.855 2.285 2.585 ;
      RECT 0.515 2.575 0.845 3.305 ;
    LAYER via2 ;
      RECT 74.04 2.315 74.24 2.515 ;
      RECT 72.44 3.04 72.64 3.24 ;
      RECT 72.215 7.14 72.415 7.34 ;
      RECT 70.88 2.48 71.08 2.68 ;
      RECT 70.5 3.6 70.7 3.8 ;
      RECT 70 2.48 70.2 2.68 ;
      RECT 69.04 2.48 69.24 2.68 ;
      RECT 68.32 2.48 68.52 2.68 ;
      RECT 67.32 1.92 67.52 2.12 ;
      RECT 65.88 3.04 66.08 3.24 ;
      RECT 57.715 2.315 57.915 2.515 ;
      RECT 56.115 3.04 56.315 3.24 ;
      RECT 55.89 7.14 56.09 7.34 ;
      RECT 54.555 2.48 54.755 2.68 ;
      RECT 54.175 3.6 54.375 3.8 ;
      RECT 53.675 2.48 53.875 2.68 ;
      RECT 52.715 2.48 52.915 2.68 ;
      RECT 51.995 2.48 52.195 2.68 ;
      RECT 50.995 1.92 51.195 2.12 ;
      RECT 49.555 3.04 49.755 3.24 ;
      RECT 41.39 2.315 41.59 2.515 ;
      RECT 39.79 3.04 39.99 3.24 ;
      RECT 39.565 7.14 39.765 7.34 ;
      RECT 38.23 2.48 38.43 2.68 ;
      RECT 37.85 3.6 38.05 3.8 ;
      RECT 37.35 2.48 37.55 2.68 ;
      RECT 36.39 2.48 36.59 2.68 ;
      RECT 35.67 2.48 35.87 2.68 ;
      RECT 34.67 1.92 34.87 2.12 ;
      RECT 33.23 3.04 33.43 3.24 ;
      RECT 25.065 2.315 25.265 2.515 ;
      RECT 23.465 3.04 23.665 3.24 ;
      RECT 23.24 7.14 23.44 7.34 ;
      RECT 21.905 2.48 22.105 2.68 ;
      RECT 21.525 3.6 21.725 3.8 ;
      RECT 21.025 2.48 21.225 2.68 ;
      RECT 20.065 2.48 20.265 2.68 ;
      RECT 19.345 2.48 19.545 2.68 ;
      RECT 18.345 1.92 18.545 2.12 ;
      RECT 16.905 3.04 17.105 3.24 ;
      RECT 8.74 2.315 8.94 2.515 ;
      RECT 7.14 3.04 7.34 3.24 ;
      RECT 6.915 7.14 7.115 7.34 ;
      RECT 5.58 2.48 5.78 2.68 ;
      RECT 5.2 3.6 5.4 3.8 ;
      RECT 4.7 2.48 4.9 2.68 ;
      RECT 3.74 2.48 3.94 2.68 ;
      RECT 3.02 2.48 3.22 2.68 ;
      RECT 2.02 1.92 2.22 2.12 ;
      RECT 0.58 3.04 0.78 3.24 ;
    LAYER met2 ;
      RECT -2.045 8.4 80.78 8.57 ;
      RECT 80.61 7.275 80.78 8.57 ;
      RECT -2.045 6.255 -1.875 8.57 ;
      RECT 80.58 7.275 80.93 7.625 ;
      RECT -2.105 6.255 -1.815 6.605 ;
      RECT 77.42 6.22 77.74 6.545 ;
      RECT 77.45 5.695 77.62 6.545 ;
      RECT 77.45 5.695 77.625 6.045 ;
      RECT 77.45 5.695 78.425 5.87 ;
      RECT 78.25 1.965 78.425 5.87 ;
      RECT 78.195 1.965 78.545 2.315 ;
      RECT 78.22 6.655 78.545 6.98 ;
      RECT 77.105 6.745 78.545 6.915 ;
      RECT 77.105 2.395 77.265 6.915 ;
      RECT 77.42 2.365 77.74 2.685 ;
      RECT 77.105 2.395 77.74 2.565 ;
      RECT 65.84 2.955 66.12 3.325 ;
      RECT 65.895 1.29 66.065 3.325 ;
      RECT 75.89 1.29 76.06 1.815 ;
      RECT 75.8 1.46 76.14 1.81 ;
      RECT 65.895 1.29 76.06 1.46 ;
      RECT 72.52 2.395 72.8 2.765 ;
      RECT 71.45 2.42 71.71 2.74 ;
      RECT 74 2.23 74.28 2.6 ;
      RECT 74.61 2.14 74.87 2.46 ;
      RECT 71.51 1.58 71.65 2.74 ;
      RECT 72.59 1.58 72.73 2.765 ;
      RECT 73.71 2.23 74.87 2.37 ;
      RECT 73.71 1.58 73.85 2.37 ;
      RECT 71.51 1.58 73.85 1.72 ;
      RECT 71.54 3.72 73.715 3.885 ;
      RECT 73.57 2.6 73.715 3.885 ;
      RECT 70.46 3.515 70.74 3.885 ;
      RECT 70.46 3.63 71.68 3.77 ;
      RECT 73.29 2.6 73.715 2.74 ;
      RECT 73.29 2.42 73.55 2.74 ;
      RECT 66.63 4 70.29 4.14 ;
      RECT 70.15 3.185 70.29 4.14 ;
      RECT 66.63 3.07 66.77 4.14 ;
      RECT 73.17 3.26 73.43 3.58 ;
      RECT 70.15 3.185 72.68 3.325 ;
      RECT 72.4 2.955 72.68 3.325 ;
      RECT 66.63 3.07 67.08 3.325 ;
      RECT 66.8 2.955 67.08 3.325 ;
      RECT 73.17 3.07 73.37 3.58 ;
      RECT 72.4 3.07 73.37 3.21 ;
      RECT 72.97 1.86 73.11 3.21 ;
      RECT 72.91 1.86 73.17 2.18 ;
      RECT 64.23 6.655 64.58 7.005 ;
      RECT 72.785 6.61 73.135 6.96 ;
      RECT 64.23 6.685 73.135 6.885 ;
      RECT 66.81 2.42 67.07 2.74 ;
      RECT 66.81 2.51 67.85 2.65 ;
      RECT 67.71 1.72 67.85 2.65 ;
      RECT 70.47 1.86 70.73 2.18 ;
      RECT 67.71 1.72 70.67 1.86 ;
      RECT 69.85 2.7 70.11 3.02 ;
      RECT 69.85 2.7 70.17 2.93 ;
      RECT 69.96 2.395 70.24 2.765 ;
      RECT 69.55 3.26 69.87 3.58 ;
      RECT 69.55 2.14 69.69 3.58 ;
      RECT 69.49 2.14 69.75 2.46 ;
      RECT 67.05 3.54 67.31 3.86 ;
      RECT 67.05 3.63 68.73 3.77 ;
      RECT 68.59 3.35 68.73 3.77 ;
      RECT 68.59 3.35 69.03 3.58 ;
      RECT 68.77 3.26 69.03 3.58 ;
      RECT 68.09 2.42 68.49 2.93 ;
      RECT 68.28 2.395 68.56 2.765 ;
      RECT 68.03 2.42 68.56 2.74 ;
      RECT 61.095 6.22 61.415 6.545 ;
      RECT 61.125 5.695 61.295 6.545 ;
      RECT 61.125 5.695 61.3 6.045 ;
      RECT 61.125 5.695 62.1 5.87 ;
      RECT 61.925 1.965 62.1 5.87 ;
      RECT 61.87 1.965 62.22 2.315 ;
      RECT 61.895 6.655 62.22 6.98 ;
      RECT 60.78 6.745 62.22 6.915 ;
      RECT 60.78 2.395 60.94 6.915 ;
      RECT 61.095 2.365 61.415 2.685 ;
      RECT 60.78 2.395 61.415 2.565 ;
      RECT 49.515 2.955 49.795 3.325 ;
      RECT 49.57 1.29 49.74 3.325 ;
      RECT 59.565 1.29 59.735 1.815 ;
      RECT 59.475 1.46 59.815 1.81 ;
      RECT 49.57 1.29 59.735 1.46 ;
      RECT 56.195 2.395 56.475 2.765 ;
      RECT 55.125 2.42 55.385 2.74 ;
      RECT 57.675 2.23 57.955 2.6 ;
      RECT 58.285 2.14 58.545 2.46 ;
      RECT 55.185 1.58 55.325 2.74 ;
      RECT 56.265 1.58 56.405 2.765 ;
      RECT 57.385 2.23 58.545 2.37 ;
      RECT 57.385 1.58 57.525 2.37 ;
      RECT 55.185 1.58 57.525 1.72 ;
      RECT 55.215 3.72 57.39 3.885 ;
      RECT 57.245 2.6 57.39 3.885 ;
      RECT 54.135 3.515 54.415 3.885 ;
      RECT 54.135 3.63 55.355 3.77 ;
      RECT 56.965 2.6 57.39 2.74 ;
      RECT 56.965 2.42 57.225 2.74 ;
      RECT 50.305 4 53.965 4.14 ;
      RECT 53.825 3.185 53.965 4.14 ;
      RECT 50.305 3.07 50.445 4.14 ;
      RECT 56.845 3.26 57.105 3.58 ;
      RECT 53.825 3.185 56.355 3.325 ;
      RECT 56.075 2.955 56.355 3.325 ;
      RECT 50.305 3.07 50.755 3.325 ;
      RECT 50.475 2.955 50.755 3.325 ;
      RECT 56.845 3.07 57.045 3.58 ;
      RECT 56.075 3.07 57.045 3.21 ;
      RECT 56.645 1.86 56.785 3.21 ;
      RECT 56.585 1.86 56.845 2.18 ;
      RECT 47.905 6.655 48.255 7.005 ;
      RECT 56.455 6.61 56.805 6.96 ;
      RECT 47.905 6.685 56.805 6.885 ;
      RECT 50.485 2.42 50.745 2.74 ;
      RECT 50.485 2.51 51.525 2.65 ;
      RECT 51.385 1.72 51.525 2.65 ;
      RECT 54.145 1.86 54.405 2.18 ;
      RECT 51.385 1.72 54.345 1.86 ;
      RECT 53.525 2.7 53.785 3.02 ;
      RECT 53.525 2.7 53.845 2.93 ;
      RECT 53.635 2.395 53.915 2.765 ;
      RECT 53.225 3.26 53.545 3.58 ;
      RECT 53.225 2.14 53.365 3.58 ;
      RECT 53.165 2.14 53.425 2.46 ;
      RECT 50.725 3.54 50.985 3.86 ;
      RECT 50.725 3.63 52.405 3.77 ;
      RECT 52.265 3.35 52.405 3.77 ;
      RECT 52.265 3.35 52.705 3.58 ;
      RECT 52.445 3.26 52.705 3.58 ;
      RECT 51.765 2.42 52.165 2.93 ;
      RECT 51.955 2.395 52.235 2.765 ;
      RECT 51.705 2.42 52.235 2.74 ;
      RECT 44.77 6.22 45.09 6.545 ;
      RECT 44.8 5.695 44.97 6.545 ;
      RECT 44.8 5.695 44.975 6.045 ;
      RECT 44.8 5.695 45.775 5.87 ;
      RECT 45.6 1.965 45.775 5.87 ;
      RECT 45.545 1.965 45.895 2.315 ;
      RECT 45.57 6.655 45.895 6.98 ;
      RECT 44.455 6.745 45.895 6.915 ;
      RECT 44.455 2.395 44.615 6.915 ;
      RECT 44.77 2.365 45.09 2.685 ;
      RECT 44.455 2.395 45.09 2.565 ;
      RECT 33.19 2.955 33.47 3.325 ;
      RECT 33.245 1.29 33.415 3.325 ;
      RECT 43.24 1.29 43.41 1.815 ;
      RECT 43.15 1.46 43.49 1.81 ;
      RECT 33.245 1.29 43.41 1.46 ;
      RECT 39.87 2.395 40.15 2.765 ;
      RECT 38.8 2.42 39.06 2.74 ;
      RECT 41.35 2.23 41.63 2.6 ;
      RECT 41.96 2.14 42.22 2.46 ;
      RECT 38.86 1.58 39 2.74 ;
      RECT 39.94 1.58 40.08 2.765 ;
      RECT 41.06 2.23 42.22 2.37 ;
      RECT 41.06 1.58 41.2 2.37 ;
      RECT 38.86 1.58 41.2 1.72 ;
      RECT 38.89 3.72 41.065 3.885 ;
      RECT 40.92 2.6 41.065 3.885 ;
      RECT 37.81 3.515 38.09 3.885 ;
      RECT 37.81 3.63 39.03 3.77 ;
      RECT 40.64 2.6 41.065 2.74 ;
      RECT 40.64 2.42 40.9 2.74 ;
      RECT 33.98 4 37.64 4.14 ;
      RECT 37.5 3.185 37.64 4.14 ;
      RECT 33.98 3.07 34.12 4.14 ;
      RECT 40.52 3.26 40.78 3.58 ;
      RECT 37.5 3.185 40.03 3.325 ;
      RECT 39.75 2.955 40.03 3.325 ;
      RECT 33.98 3.07 34.43 3.325 ;
      RECT 34.15 2.955 34.43 3.325 ;
      RECT 40.52 3.07 40.72 3.58 ;
      RECT 39.75 3.07 40.72 3.21 ;
      RECT 40.32 1.86 40.46 3.21 ;
      RECT 40.26 1.86 40.52 2.18 ;
      RECT 31.625 6.66 31.975 7.01 ;
      RECT 40.13 6.615 40.48 6.965 ;
      RECT 31.625 6.69 40.48 6.89 ;
      RECT 34.16 2.42 34.42 2.74 ;
      RECT 34.16 2.51 35.2 2.65 ;
      RECT 35.06 1.72 35.2 2.65 ;
      RECT 37.82 1.86 38.08 2.18 ;
      RECT 35.06 1.72 38.02 1.86 ;
      RECT 37.2 2.7 37.46 3.02 ;
      RECT 37.2 2.7 37.52 2.93 ;
      RECT 37.31 2.395 37.59 2.765 ;
      RECT 36.9 3.26 37.22 3.58 ;
      RECT 36.9 2.14 37.04 3.58 ;
      RECT 36.84 2.14 37.1 2.46 ;
      RECT 34.4 3.54 34.66 3.86 ;
      RECT 34.4 3.63 36.08 3.77 ;
      RECT 35.94 3.35 36.08 3.77 ;
      RECT 35.94 3.35 36.38 3.58 ;
      RECT 36.12 3.26 36.38 3.58 ;
      RECT 35.44 2.42 35.84 2.93 ;
      RECT 35.63 2.395 35.91 2.765 ;
      RECT 35.38 2.42 35.91 2.74 ;
      RECT 28.445 6.22 28.765 6.545 ;
      RECT 28.475 5.695 28.645 6.545 ;
      RECT 28.475 5.695 28.65 6.045 ;
      RECT 28.475 5.695 29.45 5.87 ;
      RECT 29.275 1.965 29.45 5.87 ;
      RECT 29.22 1.965 29.57 2.315 ;
      RECT 29.245 6.655 29.57 6.98 ;
      RECT 28.13 6.745 29.57 6.915 ;
      RECT 28.13 2.395 28.29 6.915 ;
      RECT 28.445 2.365 28.765 2.685 ;
      RECT 28.13 2.395 28.765 2.565 ;
      RECT 16.865 2.955 17.145 3.325 ;
      RECT 16.92 1.29 17.09 3.325 ;
      RECT 26.915 1.29 27.085 1.815 ;
      RECT 26.825 1.46 27.165 1.81 ;
      RECT 16.92 1.29 27.085 1.46 ;
      RECT 23.545 2.395 23.825 2.765 ;
      RECT 22.475 2.42 22.735 2.74 ;
      RECT 25.025 2.23 25.305 2.6 ;
      RECT 25.635 2.14 25.895 2.46 ;
      RECT 22.535 1.58 22.675 2.74 ;
      RECT 23.615 1.58 23.755 2.765 ;
      RECT 24.735 2.23 25.895 2.37 ;
      RECT 24.735 1.58 24.875 2.37 ;
      RECT 22.535 1.58 24.875 1.72 ;
      RECT 22.565 3.72 24.74 3.885 ;
      RECT 24.595 2.6 24.74 3.885 ;
      RECT 21.485 3.515 21.765 3.885 ;
      RECT 21.485 3.63 22.705 3.77 ;
      RECT 24.315 2.6 24.74 2.74 ;
      RECT 24.315 2.42 24.575 2.74 ;
      RECT 17.655 4 21.315 4.14 ;
      RECT 21.175 3.185 21.315 4.14 ;
      RECT 17.655 3.07 17.795 4.14 ;
      RECT 24.195 3.26 24.455 3.58 ;
      RECT 21.175 3.185 23.705 3.325 ;
      RECT 23.425 2.955 23.705 3.325 ;
      RECT 17.655 3.07 18.105 3.325 ;
      RECT 17.825 2.955 18.105 3.325 ;
      RECT 24.195 3.07 24.395 3.58 ;
      RECT 23.425 3.07 24.395 3.21 ;
      RECT 23.995 1.86 24.135 3.21 ;
      RECT 23.935 1.86 24.195 2.18 ;
      RECT 15.3 6.655 15.65 7.005 ;
      RECT 23.805 6.61 24.155 6.96 ;
      RECT 15.3 6.685 24.155 6.885 ;
      RECT 17.835 2.42 18.095 2.74 ;
      RECT 17.835 2.51 18.875 2.65 ;
      RECT 18.735 1.72 18.875 2.65 ;
      RECT 21.495 1.86 21.755 2.18 ;
      RECT 18.735 1.72 21.695 1.86 ;
      RECT 20.875 2.7 21.135 3.02 ;
      RECT 20.875 2.7 21.195 2.93 ;
      RECT 20.985 2.395 21.265 2.765 ;
      RECT 20.575 3.26 20.895 3.58 ;
      RECT 20.575 2.14 20.715 3.58 ;
      RECT 20.515 2.14 20.775 2.46 ;
      RECT 18.075 3.54 18.335 3.86 ;
      RECT 18.075 3.63 19.755 3.77 ;
      RECT 19.615 3.35 19.755 3.77 ;
      RECT 19.615 3.35 20.055 3.58 ;
      RECT 19.795 3.26 20.055 3.58 ;
      RECT 19.115 2.42 19.515 2.93 ;
      RECT 19.305 2.395 19.585 2.765 ;
      RECT 19.055 2.42 19.585 2.74 ;
      RECT 12.12 6.22 12.44 6.545 ;
      RECT 12.15 5.695 12.32 6.545 ;
      RECT 12.15 5.695 12.325 6.045 ;
      RECT 12.15 5.695 13.125 5.87 ;
      RECT 12.95 1.965 13.125 5.87 ;
      RECT 12.895 1.965 13.245 2.315 ;
      RECT 12.92 6.655 13.245 6.98 ;
      RECT 11.805 6.745 13.245 6.915 ;
      RECT 11.805 2.395 11.965 6.915 ;
      RECT 12.12 2.365 12.44 2.685 ;
      RECT 11.805 2.395 12.44 2.565 ;
      RECT 0.54 2.955 0.82 3.325 ;
      RECT 0.595 1.29 0.765 3.325 ;
      RECT 10.59 1.29 10.76 1.815 ;
      RECT 10.5 1.46 10.84 1.81 ;
      RECT 0.595 1.29 10.76 1.46 ;
      RECT 7.22 2.395 7.5 2.765 ;
      RECT 6.15 2.42 6.41 2.74 ;
      RECT 8.7 2.23 8.98 2.6 ;
      RECT 9.31 2.14 9.57 2.46 ;
      RECT 6.21 1.58 6.35 2.74 ;
      RECT 7.29 1.58 7.43 2.765 ;
      RECT 8.41 2.23 9.57 2.37 ;
      RECT 8.41 1.58 8.55 2.37 ;
      RECT 6.21 1.58 8.55 1.72 ;
      RECT -1.73 6.995 -1.44 7.345 ;
      RECT -1.73 7.05 -0.39 7.22 ;
      RECT -0.56 6.685 -0.39 7.22 ;
      RECT 8.315 6.605 8.665 6.955 ;
      RECT -0.56 6.685 8.665 6.855 ;
      RECT 6.24 3.72 8.415 3.885 ;
      RECT 8.27 2.6 8.415 3.885 ;
      RECT 5.16 3.515 5.44 3.885 ;
      RECT 5.16 3.63 6.38 3.77 ;
      RECT 7.99 2.6 8.415 2.74 ;
      RECT 7.99 2.42 8.25 2.74 ;
      RECT 1.33 4 4.99 4.14 ;
      RECT 4.85 3.185 4.99 4.14 ;
      RECT 1.33 3.07 1.47 4.14 ;
      RECT 7.87 3.26 8.13 3.58 ;
      RECT 4.85 3.185 7.38 3.325 ;
      RECT 7.1 2.955 7.38 3.325 ;
      RECT 1.33 3.07 1.78 3.325 ;
      RECT 1.5 2.955 1.78 3.325 ;
      RECT 7.87 3.07 8.07 3.58 ;
      RECT 7.1 3.07 8.07 3.21 ;
      RECT 7.67 1.86 7.81 3.21 ;
      RECT 7.61 1.86 7.87 2.18 ;
      RECT 1.51 2.42 1.77 2.74 ;
      RECT 1.51 2.51 2.55 2.65 ;
      RECT 2.41 1.72 2.55 2.65 ;
      RECT 5.17 1.86 5.43 2.18 ;
      RECT 2.41 1.72 5.37 1.86 ;
      RECT 4.55 2.7 4.81 3.02 ;
      RECT 4.55 2.7 4.87 2.93 ;
      RECT 4.66 2.395 4.94 2.765 ;
      RECT 4.25 3.26 4.57 3.58 ;
      RECT 4.25 2.14 4.39 3.58 ;
      RECT 4.19 2.14 4.45 2.46 ;
      RECT 1.75 3.54 2.01 3.86 ;
      RECT 1.75 3.63 3.43 3.77 ;
      RECT 3.29 3.35 3.43 3.77 ;
      RECT 3.29 3.35 3.73 3.58 ;
      RECT 3.47 3.26 3.73 3.58 ;
      RECT 2.79 2.42 3.19 2.93 ;
      RECT 2.98 2.395 3.26 2.765 ;
      RECT 2.73 2.42 3.26 2.74 ;
      RECT 72.13 7.055 72.5 7.425 ;
      RECT 70.84 2.395 71.12 2.765 ;
      RECT 69 2.395 69.28 2.765 ;
      RECT 67.28 1.835 67.56 2.205 ;
      RECT 55.805 7.055 56.175 7.425 ;
      RECT 54.515 2.395 54.795 2.765 ;
      RECT 52.675 2.395 52.955 2.765 ;
      RECT 50.955 1.835 51.235 2.205 ;
      RECT 39.48 7.055 39.85 7.425 ;
      RECT 38.19 2.395 38.47 2.765 ;
      RECT 36.35 2.395 36.63 2.765 ;
      RECT 34.63 1.835 34.91 2.205 ;
      RECT 23.155 7.055 23.525 7.425 ;
      RECT 21.865 2.395 22.145 2.765 ;
      RECT 20.025 2.395 20.305 2.765 ;
      RECT 18.305 1.835 18.585 2.205 ;
      RECT 6.83 7.055 7.2 7.425 ;
      RECT 5.54 2.395 5.82 2.765 ;
      RECT 3.7 2.395 3.98 2.765 ;
      RECT 1.98 1.835 2.26 2.205 ;
    LAYER via1 ;
      RECT 80.68 7.375 80.83 7.525 ;
      RECT 78.31 6.74 78.46 6.89 ;
      RECT 78.295 2.065 78.445 2.215 ;
      RECT 77.505 2.45 77.655 2.6 ;
      RECT 77.505 6.325 77.655 6.475 ;
      RECT 75.9 1.56 76.05 1.71 ;
      RECT 74.665 2.225 74.815 2.375 ;
      RECT 73.345 2.505 73.495 2.655 ;
      RECT 73.225 3.345 73.375 3.495 ;
      RECT 72.965 1.945 73.115 2.095 ;
      RECT 72.885 6.71 73.035 6.86 ;
      RECT 72.24 7.165 72.39 7.315 ;
      RECT 71.505 2.505 71.655 2.655 ;
      RECT 70.905 2.505 71.055 2.655 ;
      RECT 70.525 1.945 70.675 2.095 ;
      RECT 69.905 2.785 70.055 2.935 ;
      RECT 69.665 3.345 69.815 3.495 ;
      RECT 69.545 2.225 69.695 2.375 ;
      RECT 69.065 2.505 69.215 2.655 ;
      RECT 68.825 3.345 68.975 3.495 ;
      RECT 68.085 2.505 68.235 2.655 ;
      RECT 67.345 1.945 67.495 2.095 ;
      RECT 67.105 3.625 67.255 3.775 ;
      RECT 66.865 2.505 67.015 2.655 ;
      RECT 66.865 3.065 67.015 3.215 ;
      RECT 65.905 3.065 66.055 3.215 ;
      RECT 64.33 6.755 64.48 6.905 ;
      RECT 61.985 6.74 62.135 6.89 ;
      RECT 61.97 2.065 62.12 2.215 ;
      RECT 61.18 2.45 61.33 2.6 ;
      RECT 61.18 6.325 61.33 6.475 ;
      RECT 59.575 1.56 59.725 1.71 ;
      RECT 58.34 2.225 58.49 2.375 ;
      RECT 57.02 2.505 57.17 2.655 ;
      RECT 56.9 3.345 57.05 3.495 ;
      RECT 56.64 1.945 56.79 2.095 ;
      RECT 56.555 6.71 56.705 6.86 ;
      RECT 55.915 7.165 56.065 7.315 ;
      RECT 55.18 2.505 55.33 2.655 ;
      RECT 54.58 2.505 54.73 2.655 ;
      RECT 54.2 1.945 54.35 2.095 ;
      RECT 53.58 2.785 53.73 2.935 ;
      RECT 53.34 3.345 53.49 3.495 ;
      RECT 53.22 2.225 53.37 2.375 ;
      RECT 52.74 2.505 52.89 2.655 ;
      RECT 52.5 3.345 52.65 3.495 ;
      RECT 51.76 2.505 51.91 2.655 ;
      RECT 51.02 1.945 51.17 2.095 ;
      RECT 50.78 3.625 50.93 3.775 ;
      RECT 50.54 2.505 50.69 2.655 ;
      RECT 50.54 3.065 50.69 3.215 ;
      RECT 49.58 3.065 49.73 3.215 ;
      RECT 48.005 6.755 48.155 6.905 ;
      RECT 45.66 6.74 45.81 6.89 ;
      RECT 45.645 2.065 45.795 2.215 ;
      RECT 44.855 2.45 45.005 2.6 ;
      RECT 44.855 6.325 45.005 6.475 ;
      RECT 43.25 1.56 43.4 1.71 ;
      RECT 42.015 2.225 42.165 2.375 ;
      RECT 40.695 2.505 40.845 2.655 ;
      RECT 40.575 3.345 40.725 3.495 ;
      RECT 40.315 1.945 40.465 2.095 ;
      RECT 40.23 6.715 40.38 6.865 ;
      RECT 39.59 7.165 39.74 7.315 ;
      RECT 38.855 2.505 39.005 2.655 ;
      RECT 38.255 2.505 38.405 2.655 ;
      RECT 37.875 1.945 38.025 2.095 ;
      RECT 37.255 2.785 37.405 2.935 ;
      RECT 37.015 3.345 37.165 3.495 ;
      RECT 36.895 2.225 37.045 2.375 ;
      RECT 36.415 2.505 36.565 2.655 ;
      RECT 36.175 3.345 36.325 3.495 ;
      RECT 35.435 2.505 35.585 2.655 ;
      RECT 34.695 1.945 34.845 2.095 ;
      RECT 34.455 3.625 34.605 3.775 ;
      RECT 34.215 2.505 34.365 2.655 ;
      RECT 34.215 3.065 34.365 3.215 ;
      RECT 33.255 3.065 33.405 3.215 ;
      RECT 31.725 6.76 31.875 6.91 ;
      RECT 29.335 6.74 29.485 6.89 ;
      RECT 29.32 2.065 29.47 2.215 ;
      RECT 28.53 2.45 28.68 2.6 ;
      RECT 28.53 6.325 28.68 6.475 ;
      RECT 26.925 1.56 27.075 1.71 ;
      RECT 25.69 2.225 25.84 2.375 ;
      RECT 24.37 2.505 24.52 2.655 ;
      RECT 24.25 3.345 24.4 3.495 ;
      RECT 23.99 1.945 24.14 2.095 ;
      RECT 23.905 6.71 24.055 6.86 ;
      RECT 23.265 7.165 23.415 7.315 ;
      RECT 22.53 2.505 22.68 2.655 ;
      RECT 21.93 2.505 22.08 2.655 ;
      RECT 21.55 1.945 21.7 2.095 ;
      RECT 20.93 2.785 21.08 2.935 ;
      RECT 20.69 3.345 20.84 3.495 ;
      RECT 20.57 2.225 20.72 2.375 ;
      RECT 20.09 2.505 20.24 2.655 ;
      RECT 19.85 3.345 20 3.495 ;
      RECT 19.11 2.505 19.26 2.655 ;
      RECT 18.37 1.945 18.52 2.095 ;
      RECT 18.13 3.625 18.28 3.775 ;
      RECT 17.89 2.505 18.04 2.655 ;
      RECT 17.89 3.065 18.04 3.215 ;
      RECT 16.93 3.065 17.08 3.215 ;
      RECT 15.4 6.755 15.55 6.905 ;
      RECT 13.01 6.74 13.16 6.89 ;
      RECT 12.995 2.065 13.145 2.215 ;
      RECT 12.205 2.45 12.355 2.6 ;
      RECT 12.205 6.325 12.355 6.475 ;
      RECT 10.6 1.56 10.75 1.71 ;
      RECT 9.365 2.225 9.515 2.375 ;
      RECT 8.415 6.705 8.565 6.855 ;
      RECT 8.045 2.505 8.195 2.655 ;
      RECT 7.925 3.345 8.075 3.495 ;
      RECT 7.665 1.945 7.815 2.095 ;
      RECT 6.94 7.165 7.09 7.315 ;
      RECT 6.205 2.505 6.355 2.655 ;
      RECT 5.605 2.505 5.755 2.655 ;
      RECT 5.225 1.945 5.375 2.095 ;
      RECT 4.605 2.785 4.755 2.935 ;
      RECT 4.365 3.345 4.515 3.495 ;
      RECT 4.245 2.225 4.395 2.375 ;
      RECT 3.765 2.505 3.915 2.655 ;
      RECT 3.525 3.345 3.675 3.495 ;
      RECT 2.785 2.505 2.935 2.655 ;
      RECT 2.045 1.945 2.195 2.095 ;
      RECT 1.805 3.625 1.955 3.775 ;
      RECT 1.565 2.505 1.715 2.655 ;
      RECT 1.565 3.065 1.715 3.215 ;
      RECT 0.605 3.065 0.755 3.215 ;
      RECT -1.66 7.095 -1.51 7.245 ;
      RECT -2.035 6.355 -1.885 6.505 ;
    LAYER met1 ;
      RECT 80.545 7.77 80.835 8 ;
      RECT 80.605 6.29 80.775 8 ;
      RECT 80.58 7.275 80.93 7.625 ;
      RECT 80.545 6.29 80.835 6.52 ;
      RECT 80.14 2.395 80.245 2.965 ;
      RECT 80.14 2.73 80.465 2.96 ;
      RECT 80.14 2.76 80.635 2.93 ;
      RECT 80.14 2.395 80.33 2.96 ;
      RECT 79.555 2.36 79.845 2.59 ;
      RECT 79.555 2.395 80.33 2.565 ;
      RECT 79.615 0.88 79.785 2.59 ;
      RECT 79.555 0.88 79.845 1.11 ;
      RECT 79.555 7.77 79.845 8 ;
      RECT 79.615 6.29 79.785 8 ;
      RECT 79.555 6.29 79.845 6.52 ;
      RECT 79.555 6.325 80.41 6.485 ;
      RECT 80.24 5.92 80.41 6.485 ;
      RECT 79.555 6.32 79.95 6.485 ;
      RECT 80.175 5.92 80.465 6.15 ;
      RECT 80.175 5.95 80.635 6.12 ;
      RECT 79.185 2.73 79.475 2.96 ;
      RECT 79.185 2.76 79.645 2.93 ;
      RECT 79.25 1.655 79.415 2.96 ;
      RECT 77.765 1.625 78.055 1.855 ;
      RECT 77.765 1.655 79.415 1.825 ;
      RECT 77.825 0.885 77.995 1.855 ;
      RECT 77.765 0.885 78.055 1.115 ;
      RECT 77.765 7.765 78.055 7.995 ;
      RECT 77.825 7.025 77.995 7.995 ;
      RECT 77.825 7.12 79.415 7.29 ;
      RECT 79.245 5.92 79.415 7.29 ;
      RECT 77.765 7.025 78.055 7.255 ;
      RECT 79.185 5.92 79.475 6.15 ;
      RECT 79.185 5.95 79.645 6.12 ;
      RECT 78.195 1.965 78.545 2.315 ;
      RECT 75.89 2.025 78.545 2.195 ;
      RECT 75.89 1.46 76.06 2.195 ;
      RECT 75.8 1.46 76.14 1.81 ;
      RECT 78.22 6.655 78.545 6.98 ;
      RECT 72.785 6.61 73.135 6.96 ;
      RECT 78.195 6.655 78.545 6.885 ;
      RECT 72.58 6.655 73.135 6.885 ;
      RECT 72.41 6.685 78.545 6.855 ;
      RECT 77.42 2.365 77.74 2.685 ;
      RECT 77.39 2.365 77.74 2.595 ;
      RECT 77.22 2.395 77.74 2.565 ;
      RECT 77.42 6.255 77.74 6.545 ;
      RECT 77.39 6.285 77.74 6.515 ;
      RECT 77.22 6.315 77.74 6.485 ;
      RECT 73.875 2.465 74.165 2.695 ;
      RECT 73.875 2.465 74.33 2.65 ;
      RECT 74.19 2.37 74.81 2.51 ;
      RECT 74.58 2.17 74.9 2.43 ;
      RECT 73.26 2.45 73.58 2.71 ;
      RECT 73.26 2.45 73.725 2.695 ;
      RECT 73.585 2.07 73.725 2.695 ;
      RECT 73.585 2.07 73.85 2.21 ;
      RECT 74.115 1.905 74.405 2.135 ;
      RECT 73.71 1.95 74.405 2.09 ;
      RECT 73.155 3.29 73.445 3.815 ;
      RECT 73.14 3.29 73.46 3.55 ;
      RECT 72.88 1.89 73.2 2.15 ;
      RECT 72.88 1.905 73.445 2.135 ;
      RECT 72.155 3.585 72.445 3.815 ;
      RECT 72.35 2.23 72.49 3.77 ;
      RECT 72.395 2.185 72.685 2.415 ;
      RECT 71.99 2.23 72.685 2.37 ;
      RECT 71.99 2.07 72.13 2.37 ;
      RECT 70.53 2.07 72.13 2.21 ;
      RECT 70.44 1.89 70.76 2.15 ;
      RECT 70.44 1.905 71.005 2.15 ;
      RECT 72.15 7.765 72.44 7.995 ;
      RECT 72.21 7.025 72.38 7.995 ;
      RECT 72.13 7.075 72.5 7.425 ;
      RECT 72.13 7.055 72.44 7.425 ;
      RECT 72.15 7.025 72.44 7.425 ;
      RECT 69.55 2.93 72.13 3.07 ;
      RECT 71.915 2.745 72.205 2.975 ;
      RECT 69.475 2.745 70.14 2.975 ;
      RECT 69.82 2.73 70.14 3.07 ;
      RECT 70.82 2.45 71.14 2.71 ;
      RECT 70.82 2.465 71.245 2.695 ;
      RECT 69.46 2.17 69.78 2.43 ;
      RECT 69.955 2.185 70.245 2.415 ;
      RECT 69.46 2.23 70.245 2.37 ;
      RECT 69.58 3.29 69.9 3.55 ;
      RECT 68.74 3.29 69.06 3.55 ;
      RECT 69.58 3.305 70.005 3.535 ;
      RECT 68.74 3.35 70.005 3.49 ;
      RECT 68.275 3.025 68.565 3.255 ;
      RECT 68.35 1.95 68.49 3.255 ;
      RECT 68 2.45 68.49 2.71 ;
      RECT 67.755 2.465 68.49 2.695 ;
      RECT 68.755 1.905 69.045 2.135 ;
      RECT 68.35 1.95 69.045 2.09 ;
      RECT 67.515 3.305 67.805 3.535 ;
      RECT 67.515 3.305 67.97 3.49 ;
      RECT 67.83 2.93 67.97 3.49 ;
      RECT 67.47 2.93 67.97 3.07 ;
      RECT 67.47 1.95 67.61 3.07 ;
      RECT 67.26 1.89 67.58 2.15 ;
      RECT 67.02 3.57 67.34 3.83 ;
      RECT 66.315 3.585 66.605 3.815 ;
      RECT 66.315 3.63 67.34 3.77 ;
      RECT 66.39 3.58 66.65 3.77 ;
      RECT 66.78 2.45 67.1 2.71 ;
      RECT 66.78 2.465 67.325 2.695 ;
      RECT 66.78 3.01 67.1 3.27 ;
      RECT 66.78 3.025 67.325 3.255 ;
      RECT 65.82 3.01 66.14 3.27 ;
      RECT 65.91 1.95 66.05 3.27 ;
      RECT 66.315 1.905 66.605 2.135 ;
      RECT 65.91 1.95 66.605 2.09 ;
      RECT 64.22 7.77 64.51 8 ;
      RECT 64.28 6.29 64.45 8 ;
      RECT 64.23 6.655 64.58 7.005 ;
      RECT 64.22 6.29 64.51 6.52 ;
      RECT 63.815 2.395 63.92 2.965 ;
      RECT 63.815 2.73 64.14 2.96 ;
      RECT 63.815 2.76 64.31 2.93 ;
      RECT 63.815 2.395 64.005 2.96 ;
      RECT 63.23 2.36 63.52 2.59 ;
      RECT 63.23 2.395 64.005 2.565 ;
      RECT 63.29 0.88 63.46 2.59 ;
      RECT 63.23 0.88 63.52 1.11 ;
      RECT 63.23 7.77 63.52 8 ;
      RECT 63.29 6.29 63.46 8 ;
      RECT 63.23 6.29 63.52 6.52 ;
      RECT 63.23 6.325 64.085 6.485 ;
      RECT 63.915 5.92 64.085 6.485 ;
      RECT 63.23 6.32 63.625 6.485 ;
      RECT 63.85 5.92 64.14 6.15 ;
      RECT 63.85 5.95 64.31 6.12 ;
      RECT 62.86 2.73 63.15 2.96 ;
      RECT 62.86 2.76 63.32 2.93 ;
      RECT 62.925 1.655 63.09 2.96 ;
      RECT 61.44 1.625 61.73 1.855 ;
      RECT 61.44 1.655 63.09 1.825 ;
      RECT 61.5 0.885 61.67 1.855 ;
      RECT 61.44 0.885 61.73 1.115 ;
      RECT 61.44 7.765 61.73 7.995 ;
      RECT 61.5 7.025 61.67 7.995 ;
      RECT 61.5 7.12 63.09 7.29 ;
      RECT 62.92 5.92 63.09 7.29 ;
      RECT 61.44 7.025 61.73 7.255 ;
      RECT 62.86 5.92 63.15 6.15 ;
      RECT 62.86 5.95 63.32 6.12 ;
      RECT 61.87 1.965 62.22 2.315 ;
      RECT 59.565 2.025 62.22 2.195 ;
      RECT 59.565 1.46 59.735 2.195 ;
      RECT 59.475 1.46 59.815 1.81 ;
      RECT 61.895 6.655 62.22 6.98 ;
      RECT 56.455 6.61 56.805 6.96 ;
      RECT 61.87 6.655 62.22 6.885 ;
      RECT 56.255 6.655 56.805 6.885 ;
      RECT 56.085 6.685 62.22 6.855 ;
      RECT 61.095 2.365 61.415 2.685 ;
      RECT 61.065 2.365 61.415 2.595 ;
      RECT 60.895 2.395 61.415 2.565 ;
      RECT 61.095 6.255 61.415 6.545 ;
      RECT 61.065 6.285 61.415 6.515 ;
      RECT 60.895 6.315 61.415 6.485 ;
      RECT 57.55 2.465 57.84 2.695 ;
      RECT 57.55 2.465 58.005 2.65 ;
      RECT 57.865 2.37 58.485 2.51 ;
      RECT 58.255 2.17 58.575 2.43 ;
      RECT 56.935 2.45 57.255 2.71 ;
      RECT 56.935 2.45 57.4 2.695 ;
      RECT 57.26 2.07 57.4 2.695 ;
      RECT 57.26 2.07 57.525 2.21 ;
      RECT 57.79 1.905 58.08 2.135 ;
      RECT 57.385 1.95 58.08 2.09 ;
      RECT 56.83 3.29 57.12 3.815 ;
      RECT 56.815 3.29 57.135 3.55 ;
      RECT 56.555 1.89 56.875 2.15 ;
      RECT 56.555 1.905 57.12 2.135 ;
      RECT 55.83 3.585 56.12 3.815 ;
      RECT 56.025 2.23 56.165 3.77 ;
      RECT 56.07 2.185 56.36 2.415 ;
      RECT 55.665 2.23 56.36 2.37 ;
      RECT 55.665 2.07 55.805 2.37 ;
      RECT 54.205 2.07 55.805 2.21 ;
      RECT 54.115 1.89 54.435 2.15 ;
      RECT 54.115 1.905 54.68 2.15 ;
      RECT 55.825 7.765 56.115 7.995 ;
      RECT 55.885 7.025 56.055 7.995 ;
      RECT 55.805 7.075 56.175 7.425 ;
      RECT 55.805 7.055 56.115 7.425 ;
      RECT 55.825 7.025 56.115 7.425 ;
      RECT 53.225 2.93 55.805 3.07 ;
      RECT 55.59 2.745 55.88 2.975 ;
      RECT 53.15 2.745 53.815 2.975 ;
      RECT 53.495 2.73 53.815 3.07 ;
      RECT 54.495 2.45 54.815 2.71 ;
      RECT 54.495 2.465 54.92 2.695 ;
      RECT 53.135 2.17 53.455 2.43 ;
      RECT 53.63 2.185 53.92 2.415 ;
      RECT 53.135 2.23 53.92 2.37 ;
      RECT 53.255 3.29 53.575 3.55 ;
      RECT 52.415 3.29 52.735 3.55 ;
      RECT 53.255 3.305 53.68 3.535 ;
      RECT 52.415 3.35 53.68 3.49 ;
      RECT 51.95 3.025 52.24 3.255 ;
      RECT 52.025 1.95 52.165 3.255 ;
      RECT 51.675 2.45 52.165 2.71 ;
      RECT 51.43 2.465 52.165 2.695 ;
      RECT 52.43 1.905 52.72 2.135 ;
      RECT 52.025 1.95 52.72 2.09 ;
      RECT 51.19 3.305 51.48 3.535 ;
      RECT 51.19 3.305 51.645 3.49 ;
      RECT 51.505 2.93 51.645 3.49 ;
      RECT 51.145 2.93 51.645 3.07 ;
      RECT 51.145 1.95 51.285 3.07 ;
      RECT 50.935 1.89 51.255 2.15 ;
      RECT 50.695 3.57 51.015 3.83 ;
      RECT 49.99 3.585 50.28 3.815 ;
      RECT 49.99 3.63 51.015 3.77 ;
      RECT 50.065 3.58 50.325 3.77 ;
      RECT 50.455 2.45 50.775 2.71 ;
      RECT 50.455 2.465 51 2.695 ;
      RECT 50.455 3.01 50.775 3.27 ;
      RECT 50.455 3.025 51 3.255 ;
      RECT 49.495 3.01 49.815 3.27 ;
      RECT 49.585 1.95 49.725 3.27 ;
      RECT 49.99 1.905 50.28 2.135 ;
      RECT 49.585 1.95 50.28 2.09 ;
      RECT 47.895 7.77 48.185 8 ;
      RECT 47.955 6.29 48.125 8 ;
      RECT 47.905 6.655 48.255 7.005 ;
      RECT 47.895 6.29 48.185 6.52 ;
      RECT 47.49 2.395 47.595 2.965 ;
      RECT 47.49 2.73 47.815 2.96 ;
      RECT 47.49 2.76 47.985 2.93 ;
      RECT 47.49 2.395 47.68 2.96 ;
      RECT 46.905 2.36 47.195 2.59 ;
      RECT 46.905 2.395 47.68 2.565 ;
      RECT 46.965 0.88 47.135 2.59 ;
      RECT 46.905 0.88 47.195 1.11 ;
      RECT 46.905 7.77 47.195 8 ;
      RECT 46.965 6.29 47.135 8 ;
      RECT 46.905 6.29 47.195 6.52 ;
      RECT 46.905 6.325 47.76 6.485 ;
      RECT 47.59 5.92 47.76 6.485 ;
      RECT 46.905 6.32 47.3 6.485 ;
      RECT 47.525 5.92 47.815 6.15 ;
      RECT 47.525 5.95 47.985 6.12 ;
      RECT 46.535 2.73 46.825 2.96 ;
      RECT 46.535 2.76 46.995 2.93 ;
      RECT 46.6 1.655 46.765 2.96 ;
      RECT 45.115 1.625 45.405 1.855 ;
      RECT 45.115 1.655 46.765 1.825 ;
      RECT 45.175 0.885 45.345 1.855 ;
      RECT 45.115 0.885 45.405 1.115 ;
      RECT 45.115 7.765 45.405 7.995 ;
      RECT 45.175 7.025 45.345 7.995 ;
      RECT 45.175 7.12 46.765 7.29 ;
      RECT 46.595 5.92 46.765 7.29 ;
      RECT 45.115 7.025 45.405 7.255 ;
      RECT 46.535 5.92 46.825 6.15 ;
      RECT 46.535 5.95 46.995 6.12 ;
      RECT 45.545 1.965 45.895 2.315 ;
      RECT 43.24 2.025 45.895 2.195 ;
      RECT 43.24 1.46 43.41 2.195 ;
      RECT 43.15 1.46 43.49 1.81 ;
      RECT 45.57 6.655 45.895 6.98 ;
      RECT 40.13 6.615 40.48 6.965 ;
      RECT 45.545 6.655 45.895 6.885 ;
      RECT 39.93 6.655 40.48 6.885 ;
      RECT 39.76 6.685 45.895 6.855 ;
      RECT 44.77 2.365 45.09 2.685 ;
      RECT 44.74 2.365 45.09 2.595 ;
      RECT 44.57 2.395 45.09 2.565 ;
      RECT 44.77 6.255 45.09 6.545 ;
      RECT 44.74 6.285 45.09 6.515 ;
      RECT 44.57 6.315 45.09 6.485 ;
      RECT 41.225 2.465 41.515 2.695 ;
      RECT 41.225 2.465 41.68 2.65 ;
      RECT 41.54 2.37 42.16 2.51 ;
      RECT 41.93 2.17 42.25 2.43 ;
      RECT 40.61 2.45 40.93 2.71 ;
      RECT 40.61 2.45 41.075 2.695 ;
      RECT 40.935 2.07 41.075 2.695 ;
      RECT 40.935 2.07 41.2 2.21 ;
      RECT 41.465 1.905 41.755 2.135 ;
      RECT 41.06 1.95 41.755 2.09 ;
      RECT 40.505 3.29 40.795 3.815 ;
      RECT 40.49 3.29 40.81 3.55 ;
      RECT 40.23 1.89 40.55 2.15 ;
      RECT 40.23 1.905 40.795 2.135 ;
      RECT 39.505 3.585 39.795 3.815 ;
      RECT 39.7 2.23 39.84 3.77 ;
      RECT 39.745 2.185 40.035 2.415 ;
      RECT 39.34 2.23 40.035 2.37 ;
      RECT 39.34 2.07 39.48 2.37 ;
      RECT 37.88 2.07 39.48 2.21 ;
      RECT 37.79 1.89 38.11 2.15 ;
      RECT 37.79 1.905 38.355 2.15 ;
      RECT 39.5 7.765 39.79 7.995 ;
      RECT 39.56 7.025 39.73 7.995 ;
      RECT 39.48 7.075 39.85 7.425 ;
      RECT 39.48 7.055 39.79 7.425 ;
      RECT 39.5 7.025 39.79 7.425 ;
      RECT 36.9 2.93 39.48 3.07 ;
      RECT 39.265 2.745 39.555 2.975 ;
      RECT 36.825 2.745 37.49 2.975 ;
      RECT 37.17 2.73 37.49 3.07 ;
      RECT 38.17 2.45 38.49 2.71 ;
      RECT 38.17 2.465 38.595 2.695 ;
      RECT 36.81 2.17 37.13 2.43 ;
      RECT 37.305 2.185 37.595 2.415 ;
      RECT 36.81 2.23 37.595 2.37 ;
      RECT 36.93 3.29 37.25 3.55 ;
      RECT 36.09 3.29 36.41 3.55 ;
      RECT 36.93 3.305 37.355 3.535 ;
      RECT 36.09 3.35 37.355 3.49 ;
      RECT 35.625 3.025 35.915 3.255 ;
      RECT 35.7 1.95 35.84 3.255 ;
      RECT 35.35 2.45 35.84 2.71 ;
      RECT 35.105 2.465 35.84 2.695 ;
      RECT 36.105 1.905 36.395 2.135 ;
      RECT 35.7 1.95 36.395 2.09 ;
      RECT 34.865 3.305 35.155 3.535 ;
      RECT 34.865 3.305 35.32 3.49 ;
      RECT 35.18 2.93 35.32 3.49 ;
      RECT 34.82 2.93 35.32 3.07 ;
      RECT 34.82 1.95 34.96 3.07 ;
      RECT 34.61 1.89 34.93 2.15 ;
      RECT 34.37 3.57 34.69 3.83 ;
      RECT 33.665 3.585 33.955 3.815 ;
      RECT 33.665 3.63 34.69 3.77 ;
      RECT 33.74 3.58 34 3.77 ;
      RECT 34.13 2.45 34.45 2.71 ;
      RECT 34.13 2.465 34.675 2.695 ;
      RECT 34.13 3.01 34.45 3.27 ;
      RECT 34.13 3.025 34.675 3.255 ;
      RECT 33.17 3.01 33.49 3.27 ;
      RECT 33.26 1.95 33.4 3.27 ;
      RECT 33.665 1.905 33.955 2.135 ;
      RECT 33.26 1.95 33.955 2.09 ;
      RECT 31.57 7.77 31.86 8 ;
      RECT 31.63 6.29 31.8 8 ;
      RECT 31.62 6.66 31.975 7.015 ;
      RECT 31.57 6.29 31.86 6.52 ;
      RECT 31.165 2.395 31.27 2.965 ;
      RECT 31.165 2.73 31.49 2.96 ;
      RECT 31.165 2.76 31.66 2.93 ;
      RECT 31.165 2.395 31.355 2.96 ;
      RECT 30.58 2.36 30.87 2.59 ;
      RECT 30.58 2.395 31.355 2.565 ;
      RECT 30.64 0.88 30.81 2.59 ;
      RECT 30.58 0.88 30.87 1.11 ;
      RECT 30.58 7.77 30.87 8 ;
      RECT 30.64 6.29 30.81 8 ;
      RECT 30.58 6.29 30.87 6.52 ;
      RECT 30.58 6.325 31.435 6.485 ;
      RECT 31.265 5.92 31.435 6.485 ;
      RECT 30.58 6.32 30.975 6.485 ;
      RECT 31.2 5.92 31.49 6.15 ;
      RECT 31.2 5.95 31.66 6.12 ;
      RECT 30.21 2.73 30.5 2.96 ;
      RECT 30.21 2.76 30.67 2.93 ;
      RECT 30.275 1.655 30.44 2.96 ;
      RECT 28.79 1.625 29.08 1.855 ;
      RECT 28.79 1.655 30.44 1.825 ;
      RECT 28.85 0.885 29.02 1.855 ;
      RECT 28.79 0.885 29.08 1.115 ;
      RECT 28.79 7.765 29.08 7.995 ;
      RECT 28.85 7.025 29.02 7.995 ;
      RECT 28.85 7.12 30.44 7.29 ;
      RECT 30.27 5.92 30.44 7.29 ;
      RECT 28.79 7.025 29.08 7.255 ;
      RECT 30.21 5.92 30.5 6.15 ;
      RECT 30.21 5.95 30.67 6.12 ;
      RECT 29.22 1.965 29.57 2.315 ;
      RECT 26.915 2.025 29.57 2.195 ;
      RECT 26.915 1.46 27.085 2.195 ;
      RECT 26.825 1.46 27.165 1.81 ;
      RECT 29.245 6.655 29.57 6.98 ;
      RECT 23.805 6.61 24.155 6.96 ;
      RECT 29.22 6.655 29.57 6.885 ;
      RECT 23.605 6.655 24.155 6.885 ;
      RECT 23.435 6.685 29.57 6.855 ;
      RECT 28.445 2.365 28.765 2.685 ;
      RECT 28.415 2.365 28.765 2.595 ;
      RECT 28.245 2.395 28.765 2.565 ;
      RECT 28.445 6.255 28.765 6.545 ;
      RECT 28.415 6.285 28.765 6.515 ;
      RECT 28.245 6.315 28.765 6.485 ;
      RECT 24.9 2.465 25.19 2.695 ;
      RECT 24.9 2.465 25.355 2.65 ;
      RECT 25.215 2.37 25.835 2.51 ;
      RECT 25.605 2.17 25.925 2.43 ;
      RECT 24.285 2.45 24.605 2.71 ;
      RECT 24.285 2.45 24.75 2.695 ;
      RECT 24.61 2.07 24.75 2.695 ;
      RECT 24.61 2.07 24.875 2.21 ;
      RECT 25.14 1.905 25.43 2.135 ;
      RECT 24.735 1.95 25.43 2.09 ;
      RECT 24.18 3.29 24.47 3.815 ;
      RECT 24.165 3.29 24.485 3.55 ;
      RECT 23.905 1.89 24.225 2.15 ;
      RECT 23.905 1.905 24.47 2.135 ;
      RECT 23.18 3.585 23.47 3.815 ;
      RECT 23.375 2.23 23.515 3.77 ;
      RECT 23.42 2.185 23.71 2.415 ;
      RECT 23.015 2.23 23.71 2.37 ;
      RECT 23.015 2.07 23.155 2.37 ;
      RECT 21.555 2.07 23.155 2.21 ;
      RECT 21.465 1.89 21.785 2.15 ;
      RECT 21.465 1.905 22.03 2.15 ;
      RECT 23.175 7.765 23.465 7.995 ;
      RECT 23.235 7.025 23.405 7.995 ;
      RECT 23.155 7.075 23.525 7.425 ;
      RECT 23.155 7.055 23.465 7.425 ;
      RECT 23.175 7.025 23.465 7.425 ;
      RECT 20.575 2.93 23.155 3.07 ;
      RECT 22.94 2.745 23.23 2.975 ;
      RECT 20.5 2.745 21.165 2.975 ;
      RECT 20.845 2.73 21.165 3.07 ;
      RECT 21.845 2.45 22.165 2.71 ;
      RECT 21.845 2.465 22.27 2.695 ;
      RECT 20.485 2.17 20.805 2.43 ;
      RECT 20.98 2.185 21.27 2.415 ;
      RECT 20.485 2.23 21.27 2.37 ;
      RECT 20.605 3.29 20.925 3.55 ;
      RECT 19.765 3.29 20.085 3.55 ;
      RECT 20.605 3.305 21.03 3.535 ;
      RECT 19.765 3.35 21.03 3.49 ;
      RECT 19.3 3.025 19.59 3.255 ;
      RECT 19.375 1.95 19.515 3.255 ;
      RECT 19.025 2.45 19.515 2.71 ;
      RECT 18.78 2.465 19.515 2.695 ;
      RECT 19.78 1.905 20.07 2.135 ;
      RECT 19.375 1.95 20.07 2.09 ;
      RECT 18.54 3.305 18.83 3.535 ;
      RECT 18.54 3.305 18.995 3.49 ;
      RECT 18.855 2.93 18.995 3.49 ;
      RECT 18.495 2.93 18.995 3.07 ;
      RECT 18.495 1.95 18.635 3.07 ;
      RECT 18.285 1.89 18.605 2.15 ;
      RECT 18.045 3.57 18.365 3.83 ;
      RECT 17.34 3.585 17.63 3.815 ;
      RECT 17.34 3.63 18.365 3.77 ;
      RECT 17.415 3.58 17.675 3.77 ;
      RECT 17.805 2.45 18.125 2.71 ;
      RECT 17.805 2.465 18.35 2.695 ;
      RECT 17.805 3.01 18.125 3.27 ;
      RECT 17.805 3.025 18.35 3.255 ;
      RECT 16.845 3.01 17.165 3.27 ;
      RECT 16.935 1.95 17.075 3.27 ;
      RECT 17.34 1.905 17.63 2.135 ;
      RECT 16.935 1.95 17.63 2.09 ;
      RECT 15.245 7.77 15.535 8 ;
      RECT 15.305 6.29 15.475 8 ;
      RECT 15.3 6.655 15.65 7.005 ;
      RECT 15.245 6.29 15.535 6.52 ;
      RECT 14.84 2.395 14.945 2.965 ;
      RECT 14.84 2.73 15.165 2.96 ;
      RECT 14.84 2.76 15.335 2.93 ;
      RECT 14.84 2.395 15.03 2.96 ;
      RECT 14.255 2.36 14.545 2.59 ;
      RECT 14.255 2.395 15.03 2.565 ;
      RECT 14.315 0.88 14.485 2.59 ;
      RECT 14.255 0.88 14.545 1.11 ;
      RECT 14.255 7.77 14.545 8 ;
      RECT 14.315 6.29 14.485 8 ;
      RECT 14.255 6.29 14.545 6.52 ;
      RECT 14.255 6.325 15.11 6.485 ;
      RECT 14.94 5.92 15.11 6.485 ;
      RECT 14.255 6.32 14.65 6.485 ;
      RECT 14.875 5.92 15.165 6.15 ;
      RECT 14.875 5.95 15.335 6.12 ;
      RECT 13.885 2.73 14.175 2.96 ;
      RECT 13.885 2.76 14.345 2.93 ;
      RECT 13.95 1.655 14.115 2.96 ;
      RECT 12.465 1.625 12.755 1.855 ;
      RECT 12.465 1.655 14.115 1.825 ;
      RECT 12.525 0.885 12.695 1.855 ;
      RECT 12.465 0.885 12.755 1.115 ;
      RECT 12.465 7.765 12.755 7.995 ;
      RECT 12.525 7.025 12.695 7.995 ;
      RECT 12.525 7.12 14.115 7.29 ;
      RECT 13.945 5.92 14.115 7.29 ;
      RECT 12.465 7.025 12.755 7.255 ;
      RECT 13.885 5.92 14.175 6.15 ;
      RECT 13.885 5.95 14.345 6.12 ;
      RECT 12.895 1.965 13.245 2.315 ;
      RECT 10.59 2.025 13.245 2.195 ;
      RECT 10.59 1.46 10.76 2.195 ;
      RECT 10.5 1.46 10.84 1.81 ;
      RECT 12.92 6.655 13.245 6.98 ;
      RECT 8.315 6.605 8.665 6.955 ;
      RECT 12.895 6.655 13.245 6.885 ;
      RECT 7.28 6.655 7.57 6.885 ;
      RECT 7.11 6.685 13.245 6.855 ;
      RECT 12.12 2.365 12.44 2.685 ;
      RECT 12.09 2.365 12.44 2.595 ;
      RECT 11.92 2.395 12.44 2.565 ;
      RECT 12.12 6.255 12.44 6.545 ;
      RECT 12.09 6.285 12.44 6.515 ;
      RECT 11.92 6.315 12.44 6.485 ;
      RECT 8.575 2.465 8.865 2.695 ;
      RECT 8.575 2.465 9.03 2.65 ;
      RECT 8.89 2.37 9.51 2.51 ;
      RECT 9.28 2.17 9.6 2.43 ;
      RECT 7.96 2.45 8.28 2.71 ;
      RECT 7.96 2.45 8.425 2.695 ;
      RECT 8.285 2.07 8.425 2.695 ;
      RECT 8.285 2.07 8.55 2.21 ;
      RECT 8.815 1.905 9.105 2.135 ;
      RECT 8.41 1.95 9.105 2.09 ;
      RECT 7.855 3.29 8.145 3.815 ;
      RECT 7.84 3.29 8.16 3.55 ;
      RECT 7.58 1.89 7.9 2.15 ;
      RECT 7.58 1.905 8.145 2.135 ;
      RECT 6.855 3.585 7.145 3.815 ;
      RECT 7.05 2.23 7.19 3.77 ;
      RECT 7.095 2.185 7.385 2.415 ;
      RECT 6.69 2.23 7.385 2.37 ;
      RECT 6.69 2.07 6.83 2.37 ;
      RECT 5.23 2.07 6.83 2.21 ;
      RECT 5.14 1.89 5.46 2.15 ;
      RECT 5.14 1.905 5.705 2.15 ;
      RECT 6.85 7.765 7.14 7.995 ;
      RECT 6.91 7.025 7.08 7.995 ;
      RECT 6.83 7.075 7.2 7.425 ;
      RECT 6.83 7.055 7.14 7.425 ;
      RECT 6.85 7.025 7.14 7.425 ;
      RECT 4.25 2.93 6.83 3.07 ;
      RECT 6.615 2.745 6.905 2.975 ;
      RECT 4.175 2.745 4.84 2.975 ;
      RECT 4.52 2.73 4.84 3.07 ;
      RECT 5.52 2.45 5.84 2.71 ;
      RECT 5.52 2.465 5.945 2.695 ;
      RECT 4.16 2.17 4.48 2.43 ;
      RECT 4.655 2.185 4.945 2.415 ;
      RECT 4.16 2.23 4.945 2.37 ;
      RECT 4.28 3.29 4.6 3.55 ;
      RECT 3.44 3.29 3.76 3.55 ;
      RECT 4.28 3.305 4.705 3.535 ;
      RECT 3.44 3.35 4.705 3.49 ;
      RECT 2.975 3.025 3.265 3.255 ;
      RECT 3.05 1.95 3.19 3.255 ;
      RECT 2.7 2.45 3.19 2.71 ;
      RECT 2.455 2.465 3.19 2.695 ;
      RECT 3.455 1.905 3.745 2.135 ;
      RECT 3.05 1.95 3.745 2.09 ;
      RECT 2.215 3.305 2.505 3.535 ;
      RECT 2.215 3.305 2.67 3.49 ;
      RECT 2.53 2.93 2.67 3.49 ;
      RECT 2.17 2.93 2.67 3.07 ;
      RECT 2.17 1.95 2.31 3.07 ;
      RECT 1.96 1.89 2.28 2.15 ;
      RECT 1.72 3.57 2.04 3.83 ;
      RECT 1.015 3.585 1.305 3.815 ;
      RECT 1.015 3.63 2.04 3.77 ;
      RECT 1.09 3.58 1.35 3.77 ;
      RECT 1.48 2.45 1.8 2.71 ;
      RECT 1.48 2.465 2.025 2.695 ;
      RECT 1.48 3.01 1.8 3.27 ;
      RECT 1.48 3.025 2.025 3.255 ;
      RECT 0.52 3.01 0.84 3.27 ;
      RECT 0.61 1.95 0.75 3.27 ;
      RECT 1.015 1.905 1.305 2.135 ;
      RECT 0.61 1.95 1.305 2.09 ;
      RECT -1.73 7.765 -1.44 7.995 ;
      RECT -1.67 7.025 -1.5 7.995 ;
      RECT -1.76 7.025 -1.41 7.315 ;
      RECT -2.135 6.285 -1.785 6.575 ;
      RECT -2.275 6.315 -1.785 6.485 ;
      RECT 71.42 2.45 71.74 2.71 ;
      RECT 68.98 2.45 69.3 2.71 ;
      RECT 55.095 2.45 55.415 2.71 ;
      RECT 52.655 2.45 52.975 2.71 ;
      RECT 38.77 2.45 39.09 2.71 ;
      RECT 36.33 2.45 36.65 2.71 ;
      RECT 22.445 2.45 22.765 2.71 ;
      RECT 20.005 2.45 20.325 2.71 ;
      RECT 6.12 2.45 6.44 2.71 ;
      RECT 3.68 2.45 4 2.71 ;
    LAYER mcon ;
      RECT 80.605 6.32 80.775 6.49 ;
      RECT 80.61 6.315 80.78 6.485 ;
      RECT 64.28 6.32 64.45 6.49 ;
      RECT 64.285 6.315 64.455 6.485 ;
      RECT 47.955 6.32 48.125 6.49 ;
      RECT 47.96 6.315 48.13 6.485 ;
      RECT 31.63 6.32 31.8 6.49 ;
      RECT 31.635 6.315 31.805 6.485 ;
      RECT 15.305 6.32 15.475 6.49 ;
      RECT 15.31 6.315 15.48 6.485 ;
      RECT 80.605 7.8 80.775 7.97 ;
      RECT 80.235 2.76 80.405 2.93 ;
      RECT 80.235 5.95 80.405 6.12 ;
      RECT 79.615 0.91 79.785 1.08 ;
      RECT 79.615 2.39 79.785 2.56 ;
      RECT 79.615 6.32 79.785 6.49 ;
      RECT 79.615 7.8 79.785 7.97 ;
      RECT 79.245 2.76 79.415 2.93 ;
      RECT 79.245 5.95 79.415 6.12 ;
      RECT 78.255 2.025 78.425 2.195 ;
      RECT 78.255 6.685 78.425 6.855 ;
      RECT 77.825 0.915 77.995 1.085 ;
      RECT 77.825 1.655 77.995 1.825 ;
      RECT 77.825 7.055 77.995 7.225 ;
      RECT 77.825 7.795 77.995 7.965 ;
      RECT 77.45 2.395 77.62 2.565 ;
      RECT 77.45 6.315 77.62 6.485 ;
      RECT 74.175 1.935 74.345 2.105 ;
      RECT 73.935 2.495 74.105 2.665 ;
      RECT 73.455 2.495 73.625 2.665 ;
      RECT 73.215 1.935 73.385 2.105 ;
      RECT 73.215 3.615 73.385 3.785 ;
      RECT 72.64 6.685 72.81 6.855 ;
      RECT 72.455 2.215 72.625 2.385 ;
      RECT 72.215 3.615 72.385 3.785 ;
      RECT 72.21 7.055 72.38 7.225 ;
      RECT 72.21 7.795 72.38 7.965 ;
      RECT 71.975 2.775 72.145 2.945 ;
      RECT 71.495 2.495 71.665 2.665 ;
      RECT 71.015 2.495 71.185 2.665 ;
      RECT 70.775 1.935 70.945 2.105 ;
      RECT 70.015 2.215 70.185 2.385 ;
      RECT 69.775 3.335 69.945 3.505 ;
      RECT 69.535 2.775 69.705 2.945 ;
      RECT 69.055 2.495 69.225 2.665 ;
      RECT 68.815 1.935 68.985 2.105 ;
      RECT 68.815 3.335 68.985 3.505 ;
      RECT 68.335 3.055 68.505 3.225 ;
      RECT 67.815 2.495 67.985 2.665 ;
      RECT 67.575 3.335 67.745 3.505 ;
      RECT 67.335 1.935 67.505 2.105 ;
      RECT 67.095 2.495 67.265 2.665 ;
      RECT 67.095 3.055 67.265 3.225 ;
      RECT 66.375 1.935 66.545 2.105 ;
      RECT 66.375 3.615 66.545 3.785 ;
      RECT 65.895 3.055 66.065 3.225 ;
      RECT 64.28 7.8 64.45 7.97 ;
      RECT 63.91 2.76 64.08 2.93 ;
      RECT 63.91 5.95 64.08 6.12 ;
      RECT 63.29 0.91 63.46 1.08 ;
      RECT 63.29 2.39 63.46 2.56 ;
      RECT 63.29 6.32 63.46 6.49 ;
      RECT 63.29 7.8 63.46 7.97 ;
      RECT 62.92 2.76 63.09 2.93 ;
      RECT 62.92 5.95 63.09 6.12 ;
      RECT 61.93 2.025 62.1 2.195 ;
      RECT 61.93 6.685 62.1 6.855 ;
      RECT 61.5 0.915 61.67 1.085 ;
      RECT 61.5 1.655 61.67 1.825 ;
      RECT 61.5 7.055 61.67 7.225 ;
      RECT 61.5 7.795 61.67 7.965 ;
      RECT 61.125 2.395 61.295 2.565 ;
      RECT 61.125 6.315 61.295 6.485 ;
      RECT 57.85 1.935 58.02 2.105 ;
      RECT 57.61 2.495 57.78 2.665 ;
      RECT 57.13 2.495 57.3 2.665 ;
      RECT 56.89 1.935 57.06 2.105 ;
      RECT 56.89 3.615 57.06 3.785 ;
      RECT 56.315 6.685 56.485 6.855 ;
      RECT 56.13 2.215 56.3 2.385 ;
      RECT 55.89 3.615 56.06 3.785 ;
      RECT 55.885 7.055 56.055 7.225 ;
      RECT 55.885 7.795 56.055 7.965 ;
      RECT 55.65 2.775 55.82 2.945 ;
      RECT 55.17 2.495 55.34 2.665 ;
      RECT 54.69 2.495 54.86 2.665 ;
      RECT 54.45 1.935 54.62 2.105 ;
      RECT 53.69 2.215 53.86 2.385 ;
      RECT 53.45 3.335 53.62 3.505 ;
      RECT 53.21 2.775 53.38 2.945 ;
      RECT 52.73 2.495 52.9 2.665 ;
      RECT 52.49 1.935 52.66 2.105 ;
      RECT 52.49 3.335 52.66 3.505 ;
      RECT 52.01 3.055 52.18 3.225 ;
      RECT 51.49 2.495 51.66 2.665 ;
      RECT 51.25 3.335 51.42 3.505 ;
      RECT 51.01 1.935 51.18 2.105 ;
      RECT 50.77 2.495 50.94 2.665 ;
      RECT 50.77 3.055 50.94 3.225 ;
      RECT 50.05 1.935 50.22 2.105 ;
      RECT 50.05 3.615 50.22 3.785 ;
      RECT 49.57 3.055 49.74 3.225 ;
      RECT 47.955 7.8 48.125 7.97 ;
      RECT 47.585 2.76 47.755 2.93 ;
      RECT 47.585 5.95 47.755 6.12 ;
      RECT 46.965 0.91 47.135 1.08 ;
      RECT 46.965 2.39 47.135 2.56 ;
      RECT 46.965 6.32 47.135 6.49 ;
      RECT 46.965 7.8 47.135 7.97 ;
      RECT 46.595 2.76 46.765 2.93 ;
      RECT 46.595 5.95 46.765 6.12 ;
      RECT 45.605 2.025 45.775 2.195 ;
      RECT 45.605 6.685 45.775 6.855 ;
      RECT 45.175 0.915 45.345 1.085 ;
      RECT 45.175 1.655 45.345 1.825 ;
      RECT 45.175 7.055 45.345 7.225 ;
      RECT 45.175 7.795 45.345 7.965 ;
      RECT 44.8 2.395 44.97 2.565 ;
      RECT 44.8 6.315 44.97 6.485 ;
      RECT 41.525 1.935 41.695 2.105 ;
      RECT 41.285 2.495 41.455 2.665 ;
      RECT 40.805 2.495 40.975 2.665 ;
      RECT 40.565 1.935 40.735 2.105 ;
      RECT 40.565 3.615 40.735 3.785 ;
      RECT 39.99 6.685 40.16 6.855 ;
      RECT 39.805 2.215 39.975 2.385 ;
      RECT 39.565 3.615 39.735 3.785 ;
      RECT 39.56 7.055 39.73 7.225 ;
      RECT 39.56 7.795 39.73 7.965 ;
      RECT 39.325 2.775 39.495 2.945 ;
      RECT 38.845 2.495 39.015 2.665 ;
      RECT 38.365 2.495 38.535 2.665 ;
      RECT 38.125 1.935 38.295 2.105 ;
      RECT 37.365 2.215 37.535 2.385 ;
      RECT 37.125 3.335 37.295 3.505 ;
      RECT 36.885 2.775 37.055 2.945 ;
      RECT 36.405 2.495 36.575 2.665 ;
      RECT 36.165 1.935 36.335 2.105 ;
      RECT 36.165 3.335 36.335 3.505 ;
      RECT 35.685 3.055 35.855 3.225 ;
      RECT 35.165 2.495 35.335 2.665 ;
      RECT 34.925 3.335 35.095 3.505 ;
      RECT 34.685 1.935 34.855 2.105 ;
      RECT 34.445 2.495 34.615 2.665 ;
      RECT 34.445 3.055 34.615 3.225 ;
      RECT 33.725 1.935 33.895 2.105 ;
      RECT 33.725 3.615 33.895 3.785 ;
      RECT 33.245 3.055 33.415 3.225 ;
      RECT 31.63 7.8 31.8 7.97 ;
      RECT 31.26 2.76 31.43 2.93 ;
      RECT 31.26 5.95 31.43 6.12 ;
      RECT 30.64 0.91 30.81 1.08 ;
      RECT 30.64 2.39 30.81 2.56 ;
      RECT 30.64 6.32 30.81 6.49 ;
      RECT 30.64 7.8 30.81 7.97 ;
      RECT 30.27 2.76 30.44 2.93 ;
      RECT 30.27 5.95 30.44 6.12 ;
      RECT 29.28 2.025 29.45 2.195 ;
      RECT 29.28 6.685 29.45 6.855 ;
      RECT 28.85 0.915 29.02 1.085 ;
      RECT 28.85 1.655 29.02 1.825 ;
      RECT 28.85 7.055 29.02 7.225 ;
      RECT 28.85 7.795 29.02 7.965 ;
      RECT 28.475 2.395 28.645 2.565 ;
      RECT 28.475 6.315 28.645 6.485 ;
      RECT 25.2 1.935 25.37 2.105 ;
      RECT 24.96 2.495 25.13 2.665 ;
      RECT 24.48 2.495 24.65 2.665 ;
      RECT 24.24 1.935 24.41 2.105 ;
      RECT 24.24 3.615 24.41 3.785 ;
      RECT 23.665 6.685 23.835 6.855 ;
      RECT 23.48 2.215 23.65 2.385 ;
      RECT 23.24 3.615 23.41 3.785 ;
      RECT 23.235 7.055 23.405 7.225 ;
      RECT 23.235 7.795 23.405 7.965 ;
      RECT 23 2.775 23.17 2.945 ;
      RECT 22.52 2.495 22.69 2.665 ;
      RECT 22.04 2.495 22.21 2.665 ;
      RECT 21.8 1.935 21.97 2.105 ;
      RECT 21.04 2.215 21.21 2.385 ;
      RECT 20.8 3.335 20.97 3.505 ;
      RECT 20.56 2.775 20.73 2.945 ;
      RECT 20.08 2.495 20.25 2.665 ;
      RECT 19.84 1.935 20.01 2.105 ;
      RECT 19.84 3.335 20.01 3.505 ;
      RECT 19.36 3.055 19.53 3.225 ;
      RECT 18.84 2.495 19.01 2.665 ;
      RECT 18.6 3.335 18.77 3.505 ;
      RECT 18.36 1.935 18.53 2.105 ;
      RECT 18.12 2.495 18.29 2.665 ;
      RECT 18.12 3.055 18.29 3.225 ;
      RECT 17.4 1.935 17.57 2.105 ;
      RECT 17.4 3.615 17.57 3.785 ;
      RECT 16.92 3.055 17.09 3.225 ;
      RECT 15.305 7.8 15.475 7.97 ;
      RECT 14.935 2.76 15.105 2.93 ;
      RECT 14.935 5.95 15.105 6.12 ;
      RECT 14.315 0.91 14.485 1.08 ;
      RECT 14.315 2.39 14.485 2.56 ;
      RECT 14.315 6.32 14.485 6.49 ;
      RECT 14.315 7.8 14.485 7.97 ;
      RECT 13.945 2.76 14.115 2.93 ;
      RECT 13.945 5.95 14.115 6.12 ;
      RECT 12.955 2.025 13.125 2.195 ;
      RECT 12.955 6.685 13.125 6.855 ;
      RECT 12.525 0.915 12.695 1.085 ;
      RECT 12.525 1.655 12.695 1.825 ;
      RECT 12.525 7.055 12.695 7.225 ;
      RECT 12.525 7.795 12.695 7.965 ;
      RECT 12.15 2.395 12.32 2.565 ;
      RECT 12.15 6.315 12.32 6.485 ;
      RECT 8.875 1.935 9.045 2.105 ;
      RECT 8.635 2.495 8.805 2.665 ;
      RECT 8.155 2.495 8.325 2.665 ;
      RECT 7.915 1.935 8.085 2.105 ;
      RECT 7.915 3.615 8.085 3.785 ;
      RECT 7.34 6.685 7.51 6.855 ;
      RECT 7.155 2.215 7.325 2.385 ;
      RECT 6.915 3.615 7.085 3.785 ;
      RECT 6.91 7.055 7.08 7.225 ;
      RECT 6.91 7.795 7.08 7.965 ;
      RECT 6.675 2.775 6.845 2.945 ;
      RECT 6.195 2.495 6.365 2.665 ;
      RECT 5.715 2.495 5.885 2.665 ;
      RECT 5.475 1.935 5.645 2.105 ;
      RECT 4.715 2.215 4.885 2.385 ;
      RECT 4.475 3.335 4.645 3.505 ;
      RECT 4.235 2.775 4.405 2.945 ;
      RECT 3.755 2.495 3.925 2.665 ;
      RECT 3.515 1.935 3.685 2.105 ;
      RECT 3.515 3.335 3.685 3.505 ;
      RECT 3.035 3.055 3.205 3.225 ;
      RECT 2.515 2.495 2.685 2.665 ;
      RECT 2.275 3.335 2.445 3.505 ;
      RECT 2.035 1.935 2.205 2.105 ;
      RECT 1.795 2.495 1.965 2.665 ;
      RECT 1.795 3.055 1.965 3.225 ;
      RECT 1.075 1.935 1.245 2.105 ;
      RECT 1.075 3.615 1.245 3.785 ;
      RECT 0.595 3.055 0.765 3.225 ;
      RECT -1.67 7.055 -1.5 7.225 ;
      RECT -1.67 7.795 -1.5 7.965 ;
      RECT -2.045 6.315 -1.875 6.485 ;
    LAYER li1 ;
      RECT 80.605 5.02 80.775 6.49 ;
      RECT 80.605 6.315 80.78 6.485 ;
      RECT 80.235 1.74 80.405 2.93 ;
      RECT 80.235 1.74 80.705 1.91 ;
      RECT 80.235 6.97 80.705 7.14 ;
      RECT 80.235 5.95 80.405 7.14 ;
      RECT 79.245 1.74 79.415 2.93 ;
      RECT 79.245 1.74 79.715 1.91 ;
      RECT 79.245 6.97 79.715 7.14 ;
      RECT 79.245 5.95 79.415 7.14 ;
      RECT 77.395 2.635 77.565 3.865 ;
      RECT 77.45 0.855 77.62 2.805 ;
      RECT 77.395 0.575 77.565 1.025 ;
      RECT 77.395 7.855 77.565 8.305 ;
      RECT 77.45 6.075 77.62 8.025 ;
      RECT 77.395 5.015 77.565 6.245 ;
      RECT 76.875 0.575 77.045 3.865 ;
      RECT 76.875 2.075 77.28 2.405 ;
      RECT 76.875 1.235 77.28 1.565 ;
      RECT 76.875 5.015 77.045 8.305 ;
      RECT 76.875 7.315 77.28 7.645 ;
      RECT 76.875 6.475 77.28 6.805 ;
      RECT 74.175 1.835 74.345 2.105 ;
      RECT 74.175 1.835 74.905 2.005 ;
      RECT 74.095 3.225 74.425 3.395 ;
      RECT 73.335 3.055 74.345 3.225 ;
      RECT 73.335 2.575 73.505 3.225 ;
      RECT 73.455 2.495 73.625 2.825 ;
      RECT 72.615 3.225 72.945 3.395 ;
      RECT 70.695 3.225 71.985 3.395 ;
      RECT 71.735 3.14 72.865 3.31 ;
      RECT 72.455 2.215 72.865 2.385 ;
      RECT 72.695 1.755 72.865 2.385 ;
      RECT 71.26 5.015 71.43 8.305 ;
      RECT 71.26 7.315 71.665 7.645 ;
      RECT 71.26 6.475 71.665 6.805 ;
      RECT 69.935 2.575 71.265 2.745 ;
      RECT 71.015 2.495 71.185 2.745 ;
      RECT 70.015 2.175 70.185 2.385 ;
      RECT 70.015 2.175 70.505 2.345 ;
      RECT 68.695 3.335 68.985 3.505 ;
      RECT 68.695 2.575 68.865 3.505 ;
      RECT 68.495 2.575 68.865 2.745 ;
      RECT 67.495 2.575 67.985 2.745 ;
      RECT 67.815 2.495 67.985 2.745 ;
      RECT 67.575 3.335 67.985 3.505 ;
      RECT 67.815 3.145 67.985 3.505 ;
      RECT 66.615 3.055 67.265 3.225 ;
      RECT 66.615 2.495 66.785 3.225 ;
      RECT 66.255 3.615 66.545 3.785 ;
      RECT 66.255 2.575 66.425 3.785 ;
      RECT 66.055 2.575 66.425 2.745 ;
      RECT 64.28 5.02 64.45 6.49 ;
      RECT 64.28 6.315 64.455 6.485 ;
      RECT 63.91 1.74 64.08 2.93 ;
      RECT 63.91 1.74 64.38 1.91 ;
      RECT 63.91 6.97 64.38 7.14 ;
      RECT 63.91 5.95 64.08 7.14 ;
      RECT 62.92 1.74 63.09 2.93 ;
      RECT 62.92 1.74 63.39 1.91 ;
      RECT 62.92 6.97 63.39 7.14 ;
      RECT 62.92 5.95 63.09 7.14 ;
      RECT 61.07 2.635 61.24 3.865 ;
      RECT 61.125 0.855 61.295 2.805 ;
      RECT 61.07 0.575 61.24 1.025 ;
      RECT 61.07 7.855 61.24 8.305 ;
      RECT 61.125 6.075 61.295 8.025 ;
      RECT 61.07 5.015 61.24 6.245 ;
      RECT 60.55 0.575 60.72 3.865 ;
      RECT 60.55 2.075 60.955 2.405 ;
      RECT 60.55 1.235 60.955 1.565 ;
      RECT 60.55 5.015 60.72 8.305 ;
      RECT 60.55 7.315 60.955 7.645 ;
      RECT 60.55 6.475 60.955 6.805 ;
      RECT 57.85 1.835 58.02 2.105 ;
      RECT 57.85 1.835 58.58 2.005 ;
      RECT 57.77 3.225 58.1 3.395 ;
      RECT 57.01 3.055 58.02 3.225 ;
      RECT 57.01 2.575 57.18 3.225 ;
      RECT 57.13 2.495 57.3 2.825 ;
      RECT 56.29 3.225 56.62 3.395 ;
      RECT 54.37 3.225 55.66 3.395 ;
      RECT 55.41 3.14 56.54 3.31 ;
      RECT 56.13 2.215 56.54 2.385 ;
      RECT 56.37 1.755 56.54 2.385 ;
      RECT 54.935 5.015 55.105 8.305 ;
      RECT 54.935 7.315 55.34 7.645 ;
      RECT 54.935 6.475 55.34 6.805 ;
      RECT 53.61 2.575 54.94 2.745 ;
      RECT 54.69 2.495 54.86 2.745 ;
      RECT 53.69 2.175 53.86 2.385 ;
      RECT 53.69 2.175 54.18 2.345 ;
      RECT 52.37 3.335 52.66 3.505 ;
      RECT 52.37 2.575 52.54 3.505 ;
      RECT 52.17 2.575 52.54 2.745 ;
      RECT 51.17 2.575 51.66 2.745 ;
      RECT 51.49 2.495 51.66 2.745 ;
      RECT 51.25 3.335 51.66 3.505 ;
      RECT 51.49 3.145 51.66 3.505 ;
      RECT 50.29 3.055 50.94 3.225 ;
      RECT 50.29 2.495 50.46 3.225 ;
      RECT 49.93 3.615 50.22 3.785 ;
      RECT 49.93 2.575 50.1 3.785 ;
      RECT 49.73 2.575 50.1 2.745 ;
      RECT 47.955 5.02 48.125 6.49 ;
      RECT 47.955 6.315 48.13 6.485 ;
      RECT 47.585 1.74 47.755 2.93 ;
      RECT 47.585 1.74 48.055 1.91 ;
      RECT 47.585 6.97 48.055 7.14 ;
      RECT 47.585 5.95 47.755 7.14 ;
      RECT 46.595 1.74 46.765 2.93 ;
      RECT 46.595 1.74 47.065 1.91 ;
      RECT 46.595 6.97 47.065 7.14 ;
      RECT 46.595 5.95 46.765 7.14 ;
      RECT 44.745 2.635 44.915 3.865 ;
      RECT 44.8 0.855 44.97 2.805 ;
      RECT 44.745 0.575 44.915 1.025 ;
      RECT 44.745 7.855 44.915 8.305 ;
      RECT 44.8 6.075 44.97 8.025 ;
      RECT 44.745 5.015 44.915 6.245 ;
      RECT 44.225 0.575 44.395 3.865 ;
      RECT 44.225 2.075 44.63 2.405 ;
      RECT 44.225 1.235 44.63 1.565 ;
      RECT 44.225 5.015 44.395 8.305 ;
      RECT 44.225 7.315 44.63 7.645 ;
      RECT 44.225 6.475 44.63 6.805 ;
      RECT 41.525 1.835 41.695 2.105 ;
      RECT 41.525 1.835 42.255 2.005 ;
      RECT 41.445 3.225 41.775 3.395 ;
      RECT 40.685 3.055 41.695 3.225 ;
      RECT 40.685 2.575 40.855 3.225 ;
      RECT 40.805 2.495 40.975 2.825 ;
      RECT 39.965 3.225 40.295 3.395 ;
      RECT 38.045 3.225 39.335 3.395 ;
      RECT 39.085 3.14 40.215 3.31 ;
      RECT 39.805 2.215 40.215 2.385 ;
      RECT 40.045 1.755 40.215 2.385 ;
      RECT 38.61 5.015 38.78 8.305 ;
      RECT 38.61 7.315 39.015 7.645 ;
      RECT 38.61 6.475 39.015 6.805 ;
      RECT 37.285 2.575 38.615 2.745 ;
      RECT 38.365 2.495 38.535 2.745 ;
      RECT 37.365 2.175 37.535 2.385 ;
      RECT 37.365 2.175 37.855 2.345 ;
      RECT 36.045 3.335 36.335 3.505 ;
      RECT 36.045 2.575 36.215 3.505 ;
      RECT 35.845 2.575 36.215 2.745 ;
      RECT 34.845 2.575 35.335 2.745 ;
      RECT 35.165 2.495 35.335 2.745 ;
      RECT 34.925 3.335 35.335 3.505 ;
      RECT 35.165 3.145 35.335 3.505 ;
      RECT 33.965 3.055 34.615 3.225 ;
      RECT 33.965 2.495 34.135 3.225 ;
      RECT 33.605 3.615 33.895 3.785 ;
      RECT 33.605 2.575 33.775 3.785 ;
      RECT 33.405 2.575 33.775 2.745 ;
      RECT 31.63 5.02 31.8 6.49 ;
      RECT 31.63 6.315 31.805 6.485 ;
      RECT 31.26 1.74 31.43 2.93 ;
      RECT 31.26 1.74 31.73 1.91 ;
      RECT 31.26 6.97 31.73 7.14 ;
      RECT 31.26 5.95 31.43 7.14 ;
      RECT 30.27 1.74 30.44 2.93 ;
      RECT 30.27 1.74 30.74 1.91 ;
      RECT 30.27 6.97 30.74 7.14 ;
      RECT 30.27 5.95 30.44 7.14 ;
      RECT 28.42 2.635 28.59 3.865 ;
      RECT 28.475 0.855 28.645 2.805 ;
      RECT 28.42 0.575 28.59 1.025 ;
      RECT 28.42 7.855 28.59 8.305 ;
      RECT 28.475 6.075 28.645 8.025 ;
      RECT 28.42 5.015 28.59 6.245 ;
      RECT 27.9 0.575 28.07 3.865 ;
      RECT 27.9 2.075 28.305 2.405 ;
      RECT 27.9 1.235 28.305 1.565 ;
      RECT 27.9 5.015 28.07 8.305 ;
      RECT 27.9 7.315 28.305 7.645 ;
      RECT 27.9 6.475 28.305 6.805 ;
      RECT 25.2 1.835 25.37 2.105 ;
      RECT 25.2 1.835 25.93 2.005 ;
      RECT 25.12 3.225 25.45 3.395 ;
      RECT 24.36 3.055 25.37 3.225 ;
      RECT 24.36 2.575 24.53 3.225 ;
      RECT 24.48 2.495 24.65 2.825 ;
      RECT 23.64 3.225 23.97 3.395 ;
      RECT 21.72 3.225 23.01 3.395 ;
      RECT 22.76 3.14 23.89 3.31 ;
      RECT 23.48 2.215 23.89 2.385 ;
      RECT 23.72 1.755 23.89 2.385 ;
      RECT 22.285 5.015 22.455 8.305 ;
      RECT 22.285 7.315 22.69 7.645 ;
      RECT 22.285 6.475 22.69 6.805 ;
      RECT 20.96 2.575 22.29 2.745 ;
      RECT 22.04 2.495 22.21 2.745 ;
      RECT 21.04 2.175 21.21 2.385 ;
      RECT 21.04 2.175 21.53 2.345 ;
      RECT 19.72 3.335 20.01 3.505 ;
      RECT 19.72 2.575 19.89 3.505 ;
      RECT 19.52 2.575 19.89 2.745 ;
      RECT 18.52 2.575 19.01 2.745 ;
      RECT 18.84 2.495 19.01 2.745 ;
      RECT 18.6 3.335 19.01 3.505 ;
      RECT 18.84 3.145 19.01 3.505 ;
      RECT 17.64 3.055 18.29 3.225 ;
      RECT 17.64 2.495 17.81 3.225 ;
      RECT 17.28 3.615 17.57 3.785 ;
      RECT 17.28 2.575 17.45 3.785 ;
      RECT 17.08 2.575 17.45 2.745 ;
      RECT 15.305 5.02 15.475 6.49 ;
      RECT 15.305 6.315 15.48 6.485 ;
      RECT 14.935 1.74 15.105 2.93 ;
      RECT 14.935 1.74 15.405 1.91 ;
      RECT 14.935 6.97 15.405 7.14 ;
      RECT 14.935 5.95 15.105 7.14 ;
      RECT 13.945 1.74 14.115 2.93 ;
      RECT 13.945 1.74 14.415 1.91 ;
      RECT 13.945 6.97 14.415 7.14 ;
      RECT 13.945 5.95 14.115 7.14 ;
      RECT 12.095 2.635 12.265 3.865 ;
      RECT 12.15 0.855 12.32 2.805 ;
      RECT 12.095 0.575 12.265 1.025 ;
      RECT 12.095 7.855 12.265 8.305 ;
      RECT 12.15 6.075 12.32 8.025 ;
      RECT 12.095 5.015 12.265 6.245 ;
      RECT 11.575 0.575 11.745 3.865 ;
      RECT 11.575 2.075 11.98 2.405 ;
      RECT 11.575 1.235 11.98 1.565 ;
      RECT 11.575 5.015 11.745 8.305 ;
      RECT 11.575 7.315 11.98 7.645 ;
      RECT 11.575 6.475 11.98 6.805 ;
      RECT 8.875 1.835 9.045 2.105 ;
      RECT 8.875 1.835 9.605 2.005 ;
      RECT 8.795 3.225 9.125 3.395 ;
      RECT 8.035 3.055 9.045 3.225 ;
      RECT 8.035 2.575 8.205 3.225 ;
      RECT 8.155 2.495 8.325 2.825 ;
      RECT 7.315 3.225 7.645 3.395 ;
      RECT 5.395 3.225 6.685 3.395 ;
      RECT 6.435 3.14 7.565 3.31 ;
      RECT 7.155 2.215 7.565 2.385 ;
      RECT 7.395 1.755 7.565 2.385 ;
      RECT 5.96 5.015 6.13 8.305 ;
      RECT 5.96 7.315 6.365 7.645 ;
      RECT 5.96 6.475 6.365 6.805 ;
      RECT 4.635 2.575 5.965 2.745 ;
      RECT 5.715 2.495 5.885 2.745 ;
      RECT 4.715 2.175 4.885 2.385 ;
      RECT 4.715 2.175 5.205 2.345 ;
      RECT 3.395 3.335 3.685 3.505 ;
      RECT 3.395 2.575 3.565 3.505 ;
      RECT 3.195 2.575 3.565 2.745 ;
      RECT 2.195 2.575 2.685 2.745 ;
      RECT 2.515 2.495 2.685 2.745 ;
      RECT 2.275 3.335 2.685 3.505 ;
      RECT 2.515 3.145 2.685 3.505 ;
      RECT 1.315 3.055 1.965 3.225 ;
      RECT 1.315 2.495 1.485 3.225 ;
      RECT 0.955 3.615 1.245 3.785 ;
      RECT 0.955 2.575 1.125 3.785 ;
      RECT 0.755 2.575 1.125 2.745 ;
      RECT -2.1 7.855 -1.93 8.305 ;
      RECT -2.045 6.075 -1.875 8.025 ;
      RECT -2.1 5.015 -1.93 6.245 ;
      RECT -2.62 5.015 -2.45 8.305 ;
      RECT -2.62 7.315 -2.215 7.645 ;
      RECT -2.62 6.475 -2.215 6.805 ;
      RECT 80.605 7.8 80.775 8.31 ;
      RECT 79.615 0.57 79.785 1.08 ;
      RECT 79.615 2.39 79.785 3.86 ;
      RECT 79.615 5.02 79.785 6.49 ;
      RECT 79.615 7.8 79.785 8.31 ;
      RECT 78.255 0.575 78.425 3.865 ;
      RECT 78.255 5.015 78.425 8.305 ;
      RECT 77.825 0.575 77.995 1.085 ;
      RECT 77.825 1.655 77.995 3.865 ;
      RECT 77.825 5.015 77.995 7.225 ;
      RECT 77.825 7.795 77.995 8.305 ;
      RECT 73.935 2.495 74.105 2.825 ;
      RECT 73.215 1.755 73.385 2.105 ;
      RECT 73.215 3.485 73.385 3.815 ;
      RECT 72.64 5.015 72.81 8.305 ;
      RECT 72.215 3.485 72.385 3.815 ;
      RECT 72.21 5.015 72.38 7.225 ;
      RECT 72.21 7.795 72.38 8.305 ;
      RECT 71.975 2.495 72.145 2.945 ;
      RECT 71.495 2.495 71.665 2.825 ;
      RECT 70.775 1.755 70.945 2.105 ;
      RECT 69.775 3.145 69.945 3.505 ;
      RECT 69.535 2.495 69.705 2.945 ;
      RECT 69.055 2.495 69.225 2.825 ;
      RECT 68.815 1.755 68.985 2.105 ;
      RECT 68.335 3.055 68.505 3.475 ;
      RECT 67.335 1.755 67.505 2.105 ;
      RECT 67.095 2.495 67.265 2.825 ;
      RECT 66.375 1.755 66.545 2.105 ;
      RECT 65.895 3.055 66.065 3.475 ;
      RECT 64.28 7.8 64.45 8.31 ;
      RECT 63.29 0.57 63.46 1.08 ;
      RECT 63.29 2.39 63.46 3.86 ;
      RECT 63.29 5.02 63.46 6.49 ;
      RECT 63.29 7.8 63.46 8.31 ;
      RECT 61.93 0.575 62.1 3.865 ;
      RECT 61.93 5.015 62.1 8.305 ;
      RECT 61.5 0.575 61.67 1.085 ;
      RECT 61.5 1.655 61.67 3.865 ;
      RECT 61.5 5.015 61.67 7.225 ;
      RECT 61.5 7.795 61.67 8.305 ;
      RECT 57.61 2.495 57.78 2.825 ;
      RECT 56.89 1.755 57.06 2.105 ;
      RECT 56.89 3.485 57.06 3.815 ;
      RECT 56.315 5.015 56.485 8.305 ;
      RECT 55.89 3.485 56.06 3.815 ;
      RECT 55.885 5.015 56.055 7.225 ;
      RECT 55.885 7.795 56.055 8.305 ;
      RECT 55.65 2.495 55.82 2.945 ;
      RECT 55.17 2.495 55.34 2.825 ;
      RECT 54.45 1.755 54.62 2.105 ;
      RECT 53.45 3.145 53.62 3.505 ;
      RECT 53.21 2.495 53.38 2.945 ;
      RECT 52.73 2.495 52.9 2.825 ;
      RECT 52.49 1.755 52.66 2.105 ;
      RECT 52.01 3.055 52.18 3.475 ;
      RECT 51.01 1.755 51.18 2.105 ;
      RECT 50.77 2.495 50.94 2.825 ;
      RECT 50.05 1.755 50.22 2.105 ;
      RECT 49.57 3.055 49.74 3.475 ;
      RECT 47.955 7.8 48.125 8.31 ;
      RECT 46.965 0.57 47.135 1.08 ;
      RECT 46.965 2.39 47.135 3.86 ;
      RECT 46.965 5.02 47.135 6.49 ;
      RECT 46.965 7.8 47.135 8.31 ;
      RECT 45.605 0.575 45.775 3.865 ;
      RECT 45.605 5.015 45.775 8.305 ;
      RECT 45.175 0.575 45.345 1.085 ;
      RECT 45.175 1.655 45.345 3.865 ;
      RECT 45.175 5.015 45.345 7.225 ;
      RECT 45.175 7.795 45.345 8.305 ;
      RECT 41.285 2.495 41.455 2.825 ;
      RECT 40.565 1.755 40.735 2.105 ;
      RECT 40.565 3.485 40.735 3.815 ;
      RECT 39.99 5.015 40.16 8.305 ;
      RECT 39.565 3.485 39.735 3.815 ;
      RECT 39.56 5.015 39.73 7.225 ;
      RECT 39.56 7.795 39.73 8.305 ;
      RECT 39.325 2.495 39.495 2.945 ;
      RECT 38.845 2.495 39.015 2.825 ;
      RECT 38.125 1.755 38.295 2.105 ;
      RECT 37.125 3.145 37.295 3.505 ;
      RECT 36.885 2.495 37.055 2.945 ;
      RECT 36.405 2.495 36.575 2.825 ;
      RECT 36.165 1.755 36.335 2.105 ;
      RECT 35.685 3.055 35.855 3.475 ;
      RECT 34.685 1.755 34.855 2.105 ;
      RECT 34.445 2.495 34.615 2.825 ;
      RECT 33.725 1.755 33.895 2.105 ;
      RECT 33.245 3.055 33.415 3.475 ;
      RECT 31.63 7.8 31.8 8.31 ;
      RECT 30.64 0.57 30.81 1.08 ;
      RECT 30.64 2.39 30.81 3.86 ;
      RECT 30.64 5.02 30.81 6.49 ;
      RECT 30.64 7.8 30.81 8.31 ;
      RECT 29.28 0.575 29.45 3.865 ;
      RECT 29.28 5.015 29.45 8.305 ;
      RECT 28.85 0.575 29.02 1.085 ;
      RECT 28.85 1.655 29.02 3.865 ;
      RECT 28.85 5.015 29.02 7.225 ;
      RECT 28.85 7.795 29.02 8.305 ;
      RECT 24.96 2.495 25.13 2.825 ;
      RECT 24.24 1.755 24.41 2.105 ;
      RECT 24.24 3.485 24.41 3.815 ;
      RECT 23.665 5.015 23.835 8.305 ;
      RECT 23.24 3.485 23.41 3.815 ;
      RECT 23.235 5.015 23.405 7.225 ;
      RECT 23.235 7.795 23.405 8.305 ;
      RECT 23 2.495 23.17 2.945 ;
      RECT 22.52 2.495 22.69 2.825 ;
      RECT 21.8 1.755 21.97 2.105 ;
      RECT 20.8 3.145 20.97 3.505 ;
      RECT 20.56 2.495 20.73 2.945 ;
      RECT 20.08 2.495 20.25 2.825 ;
      RECT 19.84 1.755 20.01 2.105 ;
      RECT 19.36 3.055 19.53 3.475 ;
      RECT 18.36 1.755 18.53 2.105 ;
      RECT 18.12 2.495 18.29 2.825 ;
      RECT 17.4 1.755 17.57 2.105 ;
      RECT 16.92 3.055 17.09 3.475 ;
      RECT 15.305 7.8 15.475 8.31 ;
      RECT 14.315 0.57 14.485 1.08 ;
      RECT 14.315 2.39 14.485 3.86 ;
      RECT 14.315 5.02 14.485 6.49 ;
      RECT 14.315 7.8 14.485 8.31 ;
      RECT 12.955 0.575 13.125 3.865 ;
      RECT 12.955 5.015 13.125 8.305 ;
      RECT 12.525 0.575 12.695 1.085 ;
      RECT 12.525 1.655 12.695 3.865 ;
      RECT 12.525 5.015 12.695 7.225 ;
      RECT 12.525 7.795 12.695 8.305 ;
      RECT 8.635 2.495 8.805 2.825 ;
      RECT 7.915 1.755 8.085 2.105 ;
      RECT 7.915 3.485 8.085 3.815 ;
      RECT 7.34 5.015 7.51 8.305 ;
      RECT 6.915 3.485 7.085 3.815 ;
      RECT 6.91 5.015 7.08 7.225 ;
      RECT 6.91 7.795 7.08 8.305 ;
      RECT 6.675 2.495 6.845 2.945 ;
      RECT 6.195 2.495 6.365 2.825 ;
      RECT 5.475 1.755 5.645 2.105 ;
      RECT 4.475 3.145 4.645 3.505 ;
      RECT 4.235 2.495 4.405 2.945 ;
      RECT 3.755 2.495 3.925 2.825 ;
      RECT 3.515 1.755 3.685 2.105 ;
      RECT 3.035 3.055 3.205 3.475 ;
      RECT 2.035 1.755 2.205 2.105 ;
      RECT 1.795 2.495 1.965 2.825 ;
      RECT 1.075 1.755 1.245 2.105 ;
      RECT 0.595 3.055 0.765 3.475 ;
      RECT -1.67 5.015 -1.5 7.225 ;
      RECT -1.67 7.795 -1.5 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2ea_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2et_8_b0r1
  CLASS BLOCK ;
  ORIGIN 5.505 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2et_8_b0r1 ;
  SIZE 95.595 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 15.31 0.915 15.48 1.085 ;
        RECT 15.305 0.91 15.475 1.08 ;
        RECT 15.305 2.39 15.475 2.56 ;
      LAYER li1 ;
        RECT 15.31 0.915 15.48 1.085 ;
        RECT 15.305 0.57 15.475 1.08 ;
        RECT 15.305 2.39 15.475 3.86 ;
      LAYER met1 ;
        RECT 15.245 2.36 15.535 2.59 ;
        RECT 15.245 0.88 15.535 1.11 ;
        RECT 15.305 0.88 15.475 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 33.87 0.915 34.04 1.085 ;
        RECT 33.865 0.91 34.035 1.08 ;
        RECT 33.865 2.39 34.035 2.56 ;
      LAYER li1 ;
        RECT 33.87 0.915 34.04 1.085 ;
        RECT 33.865 0.57 34.035 1.08 ;
        RECT 33.865 2.39 34.035 3.86 ;
      LAYER met1 ;
        RECT 33.805 2.36 34.095 2.59 ;
        RECT 33.805 0.88 34.095 1.11 ;
        RECT 33.865 0.88 34.035 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 52.43 0.915 52.6 1.085 ;
        RECT 52.425 0.91 52.595 1.08 ;
        RECT 52.425 2.39 52.595 2.56 ;
      LAYER li1 ;
        RECT 52.43 0.915 52.6 1.085 ;
        RECT 52.425 0.57 52.595 1.08 ;
        RECT 52.425 2.39 52.595 3.86 ;
      LAYER met1 ;
        RECT 52.365 2.36 52.655 2.59 ;
        RECT 52.365 0.88 52.655 1.11 ;
        RECT 52.425 0.88 52.595 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 70.99 0.915 71.16 1.085 ;
        RECT 70.985 0.91 71.155 1.08 ;
        RECT 70.985 2.39 71.155 2.56 ;
      LAYER li1 ;
        RECT 70.99 0.915 71.16 1.085 ;
        RECT 70.985 0.57 71.155 1.08 ;
        RECT 70.985 2.39 71.155 3.86 ;
      LAYER met1 ;
        RECT 70.925 2.36 71.215 2.59 ;
        RECT 70.925 0.88 71.215 1.11 ;
        RECT 70.985 0.88 71.155 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 89.55 0.915 89.72 1.085 ;
        RECT 89.545 0.91 89.715 1.08 ;
        RECT 89.545 2.39 89.715 2.56 ;
      LAYER li1 ;
        RECT 89.55 0.915 89.72 1.085 ;
        RECT 89.545 0.57 89.715 1.08 ;
        RECT 89.545 2.39 89.715 3.86 ;
      LAYER met1 ;
        RECT 89.485 2.36 89.775 2.59 ;
        RECT 89.485 0.88 89.775 1.11 ;
        RECT 89.545 0.88 89.715 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 11.155 1.66 11.325 2.935 ;
        RECT 11.155 5.945 11.325 7.22 ;
        RECT 5.54 5.945 5.71 7.22 ;
      LAYER met2 ;
        RECT 11.08 2.705 11.42 3.055 ;
        RECT 11.07 5.845 11.41 6.195 ;
        RECT 11.155 2.705 11.325 6.195 ;
      LAYER met1 ;
        RECT 11.08 2.765 11.555 2.935 ;
        RECT 11.08 2.705 11.42 3.055 ;
        RECT 5.48 5.945 11.555 6.115 ;
        RECT 11.07 5.845 11.41 6.195 ;
        RECT 5.48 5.915 5.77 6.145 ;
      LAYER via1 ;
        RECT 11.17 5.945 11.32 6.095 ;
        RECT 11.18 2.805 11.33 2.955 ;
      LAYER mcon ;
        RECT 5.54 5.945 5.71 6.115 ;
        RECT 11.155 5.945 11.325 6.115 ;
        RECT 11.155 2.765 11.325 2.935 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 29.715 1.66 29.885 2.935 ;
        RECT 29.715 5.945 29.885 7.22 ;
        RECT 24.1 5.945 24.27 7.22 ;
      LAYER met2 ;
        RECT 29.64 2.705 29.98 3.055 ;
        RECT 29.63 5.845 29.97 6.195 ;
        RECT 29.715 2.705 29.885 6.195 ;
      LAYER met1 ;
        RECT 29.64 2.765 30.115 2.935 ;
        RECT 29.64 2.705 29.98 3.055 ;
        RECT 24.04 5.945 30.115 6.115 ;
        RECT 29.63 5.845 29.97 6.195 ;
        RECT 24.04 5.915 24.33 6.145 ;
      LAYER via1 ;
        RECT 29.73 5.945 29.88 6.095 ;
        RECT 29.74 2.805 29.89 2.955 ;
      LAYER mcon ;
        RECT 24.1 5.945 24.27 6.115 ;
        RECT 29.715 5.945 29.885 6.115 ;
        RECT 29.715 2.765 29.885 2.935 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 48.275 1.66 48.445 2.935 ;
        RECT 48.275 5.945 48.445 7.22 ;
        RECT 42.66 5.945 42.83 7.22 ;
      LAYER met2 ;
        RECT 48.2 2.705 48.54 3.055 ;
        RECT 48.19 5.845 48.53 6.195 ;
        RECT 48.275 2.705 48.445 6.195 ;
      LAYER met1 ;
        RECT 48.2 2.765 48.675 2.935 ;
        RECT 48.2 2.705 48.54 3.055 ;
        RECT 42.6 5.945 48.675 6.115 ;
        RECT 48.19 5.845 48.53 6.195 ;
        RECT 42.6 5.915 42.89 6.145 ;
      LAYER via1 ;
        RECT 48.29 5.945 48.44 6.095 ;
        RECT 48.3 2.805 48.45 2.955 ;
      LAYER mcon ;
        RECT 42.66 5.945 42.83 6.115 ;
        RECT 48.275 5.945 48.445 6.115 ;
        RECT 48.275 2.765 48.445 2.935 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 66.835 1.66 67.005 2.935 ;
        RECT 66.835 5.945 67.005 7.22 ;
        RECT 61.22 5.945 61.39 7.22 ;
      LAYER met2 ;
        RECT 66.76 2.705 67.1 3.055 ;
        RECT 66.75 5.845 67.09 6.195 ;
        RECT 66.835 2.705 67.005 6.195 ;
      LAYER met1 ;
        RECT 66.76 2.765 67.235 2.935 ;
        RECT 66.76 2.705 67.1 3.055 ;
        RECT 61.16 5.945 67.235 6.115 ;
        RECT 66.75 5.845 67.09 6.195 ;
        RECT 61.16 5.915 61.45 6.145 ;
      LAYER via1 ;
        RECT 66.85 5.945 67 6.095 ;
        RECT 66.86 2.805 67.01 2.955 ;
      LAYER mcon ;
        RECT 61.22 5.945 61.39 6.115 ;
        RECT 66.835 5.945 67.005 6.115 ;
        RECT 66.835 2.765 67.005 2.935 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 85.395 1.66 85.565 2.935 ;
        RECT 85.395 5.945 85.565 7.22 ;
        RECT 79.78 5.945 79.95 7.22 ;
      LAYER met2 ;
        RECT 85.32 2.705 85.66 3.055 ;
        RECT 85.31 5.845 85.65 6.195 ;
        RECT 85.395 2.705 85.565 6.195 ;
      LAYER met1 ;
        RECT 85.32 2.765 85.795 2.935 ;
        RECT 85.32 2.705 85.66 3.055 ;
        RECT 79.72 5.945 85.795 6.115 ;
        RECT 85.31 5.845 85.65 6.195 ;
        RECT 79.72 5.915 80.01 6.145 ;
      LAYER via1 ;
        RECT 85.41 5.945 85.56 6.095 ;
        RECT 85.42 2.805 85.57 2.955 ;
      LAYER mcon ;
        RECT 79.78 5.945 79.95 6.115 ;
        RECT 85.395 5.945 85.565 6.115 ;
        RECT 85.395 2.765 85.565 2.935 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT -5.275 5.945 -5.105 7.22 ;
      LAYER met1 ;
        RECT -5.335 5.945 -4.875 6.115 ;
        RECT -5.335 5.915 -5.045 6.145 ;
      LAYER mcon ;
        RECT -5.275 5.945 -5.105 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 72.275 4.135 90.09 4.745 ;
        RECT 87.955 4.13 89.935 4.75 ;
        RECT 89.115 3.4 89.285 5.48 ;
        RECT 88.125 3.4 88.295 5.48 ;
        RECT 85.385 3.405 85.555 5.475 ;
        RECT 82.365 3.635 82.535 4.745 ;
        RECT 79.925 3.635 80.095 4.745 ;
        RECT 79.77 4.135 79.94 5.475 ;
        RECT 77.965 3.635 78.135 4.745 ;
        RECT 77.005 3.635 77.175 4.745 ;
        RECT 75.045 3.635 75.215 4.745 ;
        RECT 74.045 3.635 74.215 4.745 ;
        RECT 71.53 4.145 73.995 4.75 ;
        RECT 73.085 3.635 73.255 4.75 ;
        RECT 53.715 4.135 71.53 4.745 ;
        RECT 69.395 4.13 71.375 4.75 ;
        RECT 70.555 3.4 70.725 5.48 ;
        RECT 69.565 3.4 69.735 5.48 ;
        RECT 66.825 3.405 66.995 5.475 ;
        RECT 63.805 3.635 63.975 4.745 ;
        RECT 61.365 3.635 61.535 4.745 ;
        RECT 61.21 4.135 61.38 5.475 ;
        RECT 59.405 3.635 59.575 4.745 ;
        RECT 58.445 3.635 58.615 4.745 ;
        RECT 56.485 3.635 56.655 4.745 ;
        RECT 55.485 3.635 55.655 4.745 ;
        RECT 52.97 4.145 55.435 4.75 ;
        RECT 54.525 3.635 54.695 4.75 ;
        RECT 35.155 4.135 52.97 4.745 ;
        RECT 50.835 4.13 52.815 4.75 ;
        RECT 51.995 3.4 52.165 5.48 ;
        RECT 51.005 3.4 51.175 5.48 ;
        RECT 48.265 3.405 48.435 5.475 ;
        RECT 45.245 3.635 45.415 4.745 ;
        RECT 42.805 3.635 42.975 4.745 ;
        RECT 42.65 4.135 42.82 5.475 ;
        RECT 40.845 3.635 41.015 4.745 ;
        RECT 39.885 3.635 40.055 4.745 ;
        RECT 37.925 3.635 38.095 4.745 ;
        RECT 36.925 3.635 37.095 4.745 ;
        RECT 34.41 4.145 36.875 4.75 ;
        RECT 35.965 3.635 36.135 4.75 ;
        RECT 16.595 4.135 34.41 4.745 ;
        RECT 32.275 4.13 34.255 4.75 ;
        RECT 33.435 3.4 33.605 5.48 ;
        RECT 32.445 3.4 32.615 5.48 ;
        RECT 29.705 3.405 29.875 5.475 ;
        RECT 26.685 3.635 26.855 4.745 ;
        RECT 24.245 3.635 24.415 4.745 ;
        RECT 24.09 4.135 24.26 5.475 ;
        RECT 22.285 3.635 22.455 4.745 ;
        RECT 21.325 3.635 21.495 4.745 ;
        RECT 19.365 3.635 19.535 4.745 ;
        RECT 18.365 3.635 18.535 4.745 ;
        RECT 15.85 4.145 18.315 4.75 ;
        RECT 17.405 3.635 17.575 4.75 ;
        RECT -1.965 4.135 15.85 4.745 ;
        RECT 13.715 4.13 15.695 4.75 ;
        RECT 14.875 3.4 15.045 5.48 ;
        RECT 13.885 3.4 14.055 5.48 ;
        RECT 11.145 3.405 11.315 5.475 ;
        RECT 8.125 3.635 8.295 4.745 ;
        RECT 5.685 3.635 5.855 4.745 ;
        RECT 5.53 4.135 5.7 5.475 ;
        RECT 3.725 3.635 3.895 4.745 ;
        RECT 2.765 3.635 2.935 4.745 ;
        RECT 0.805 3.635 0.975 4.745 ;
        RECT -0.195 3.635 -0.025 4.745 ;
        RECT -5.505 4.145 -0.245 4.75 ;
        RECT -1.155 3.635 -0.985 4.75 ;
        RECT -3.475 4.145 -3.305 8.305 ;
        RECT -5.285 4.145 -5.115 5.475 ;
      LAYER met1 ;
        RECT 72.275 4.135 90.09 4.745 ;
        RECT 87.955 4.13 89.935 4.75 ;
        RECT 72.275 3.98 84.235 4.745 ;
        RECT 71.53 4.145 73.995 4.75 ;
        RECT 53.715 4.135 71.53 4.745 ;
        RECT 69.395 4.13 71.375 4.75 ;
        RECT 53.715 3.98 65.675 4.745 ;
        RECT 52.97 4.145 55.435 4.75 ;
        RECT 35.155 4.135 52.97 4.745 ;
        RECT 50.835 4.13 52.815 4.75 ;
        RECT 35.155 3.98 47.115 4.745 ;
        RECT 34.41 4.145 36.875 4.75 ;
        RECT 16.595 4.135 34.41 4.745 ;
        RECT 32.275 4.13 34.255 4.75 ;
        RECT 16.595 3.98 28.555 4.745 ;
        RECT 15.85 4.145 18.315 4.75 ;
        RECT -1.965 4.135 15.85 4.745 ;
        RECT 13.715 4.13 15.695 4.75 ;
        RECT -1.965 3.98 9.995 4.745 ;
        RECT -5.505 4.145 -0.245 4.75 ;
        RECT -3.535 6.655 -3.245 6.885 ;
        RECT -3.705 6.685 -3.245 6.855 ;
      LAYER mcon ;
        RECT -3.475 6.685 -3.305 6.855 ;
        RECT -3.165 4.545 -2.995 4.715 ;
        RECT -1.82 4.135 -1.65 4.305 ;
        RECT -1.36 4.135 -1.19 4.305 ;
        RECT -0.9 4.135 -0.73 4.305 ;
        RECT -0.44 4.135 -0.27 4.305 ;
        RECT 0.02 4.135 0.19 4.305 ;
        RECT 0.48 4.135 0.65 4.305 ;
        RECT 0.94 4.135 1.11 4.305 ;
        RECT 1.4 4.135 1.57 4.305 ;
        RECT 1.86 4.135 2.03 4.305 ;
        RECT 2.32 4.135 2.49 4.305 ;
        RECT 2.78 4.135 2.95 4.305 ;
        RECT 3.24 4.135 3.41 4.305 ;
        RECT 3.7 4.135 3.87 4.305 ;
        RECT 4.16 4.135 4.33 4.305 ;
        RECT 4.62 4.135 4.79 4.305 ;
        RECT 5.08 4.135 5.25 4.305 ;
        RECT 5.54 4.135 5.71 4.305 ;
        RECT 6 4.135 6.17 4.305 ;
        RECT 6.46 4.135 6.63 4.305 ;
        RECT 6.92 4.135 7.09 4.305 ;
        RECT 7.38 4.135 7.55 4.305 ;
        RECT 7.65 4.545 7.82 4.715 ;
        RECT 7.84 4.135 8.01 4.305 ;
        RECT 8.3 4.135 8.47 4.305 ;
        RECT 8.76 4.135 8.93 4.305 ;
        RECT 9.22 4.135 9.39 4.305 ;
        RECT 9.68 4.135 9.85 4.305 ;
        RECT 13.265 4.545 13.435 4.715 ;
        RECT 13.265 4.165 13.435 4.335 ;
        RECT 13.965 4.55 14.135 4.72 ;
        RECT 13.965 4.16 14.135 4.33 ;
        RECT 14.955 4.55 15.125 4.72 ;
        RECT 14.955 4.16 15.125 4.33 ;
        RECT 16.74 4.135 16.91 4.305 ;
        RECT 17.2 4.135 17.37 4.305 ;
        RECT 17.66 4.135 17.83 4.305 ;
        RECT 18.12 4.135 18.29 4.305 ;
        RECT 18.58 4.135 18.75 4.305 ;
        RECT 19.04 4.135 19.21 4.305 ;
        RECT 19.5 4.135 19.67 4.305 ;
        RECT 19.96 4.135 20.13 4.305 ;
        RECT 20.42 4.135 20.59 4.305 ;
        RECT 20.88 4.135 21.05 4.305 ;
        RECT 21.34 4.135 21.51 4.305 ;
        RECT 21.8 4.135 21.97 4.305 ;
        RECT 22.26 4.135 22.43 4.305 ;
        RECT 22.72 4.135 22.89 4.305 ;
        RECT 23.18 4.135 23.35 4.305 ;
        RECT 23.64 4.135 23.81 4.305 ;
        RECT 24.1 4.135 24.27 4.305 ;
        RECT 24.56 4.135 24.73 4.305 ;
        RECT 25.02 4.135 25.19 4.305 ;
        RECT 25.48 4.135 25.65 4.305 ;
        RECT 25.94 4.135 26.11 4.305 ;
        RECT 26.21 4.545 26.38 4.715 ;
        RECT 26.4 4.135 26.57 4.305 ;
        RECT 26.86 4.135 27.03 4.305 ;
        RECT 27.32 4.135 27.49 4.305 ;
        RECT 27.78 4.135 27.95 4.305 ;
        RECT 28.24 4.135 28.41 4.305 ;
        RECT 31.825 4.545 31.995 4.715 ;
        RECT 31.825 4.165 31.995 4.335 ;
        RECT 32.525 4.55 32.695 4.72 ;
        RECT 32.525 4.16 32.695 4.33 ;
        RECT 33.515 4.55 33.685 4.72 ;
        RECT 33.515 4.16 33.685 4.33 ;
        RECT 35.3 4.135 35.47 4.305 ;
        RECT 35.76 4.135 35.93 4.305 ;
        RECT 36.22 4.135 36.39 4.305 ;
        RECT 36.68 4.135 36.85 4.305 ;
        RECT 37.14 4.135 37.31 4.305 ;
        RECT 37.6 4.135 37.77 4.305 ;
        RECT 38.06 4.135 38.23 4.305 ;
        RECT 38.52 4.135 38.69 4.305 ;
        RECT 38.98 4.135 39.15 4.305 ;
        RECT 39.44 4.135 39.61 4.305 ;
        RECT 39.9 4.135 40.07 4.305 ;
        RECT 40.36 4.135 40.53 4.305 ;
        RECT 40.82 4.135 40.99 4.305 ;
        RECT 41.28 4.135 41.45 4.305 ;
        RECT 41.74 4.135 41.91 4.305 ;
        RECT 42.2 4.135 42.37 4.305 ;
        RECT 42.66 4.135 42.83 4.305 ;
        RECT 43.12 4.135 43.29 4.305 ;
        RECT 43.58 4.135 43.75 4.305 ;
        RECT 44.04 4.135 44.21 4.305 ;
        RECT 44.5 4.135 44.67 4.305 ;
        RECT 44.77 4.545 44.94 4.715 ;
        RECT 44.96 4.135 45.13 4.305 ;
        RECT 45.42 4.135 45.59 4.305 ;
        RECT 45.88 4.135 46.05 4.305 ;
        RECT 46.34 4.135 46.51 4.305 ;
        RECT 46.8 4.135 46.97 4.305 ;
        RECT 50.385 4.545 50.555 4.715 ;
        RECT 50.385 4.165 50.555 4.335 ;
        RECT 51.085 4.55 51.255 4.72 ;
        RECT 51.085 4.16 51.255 4.33 ;
        RECT 52.075 4.55 52.245 4.72 ;
        RECT 52.075 4.16 52.245 4.33 ;
        RECT 53.86 4.135 54.03 4.305 ;
        RECT 54.32 4.135 54.49 4.305 ;
        RECT 54.78 4.135 54.95 4.305 ;
        RECT 55.24 4.135 55.41 4.305 ;
        RECT 55.7 4.135 55.87 4.305 ;
        RECT 56.16 4.135 56.33 4.305 ;
        RECT 56.62 4.135 56.79 4.305 ;
        RECT 57.08 4.135 57.25 4.305 ;
        RECT 57.54 4.135 57.71 4.305 ;
        RECT 58 4.135 58.17 4.305 ;
        RECT 58.46 4.135 58.63 4.305 ;
        RECT 58.92 4.135 59.09 4.305 ;
        RECT 59.38 4.135 59.55 4.305 ;
        RECT 59.84 4.135 60.01 4.305 ;
        RECT 60.3 4.135 60.47 4.305 ;
        RECT 60.76 4.135 60.93 4.305 ;
        RECT 61.22 4.135 61.39 4.305 ;
        RECT 61.68 4.135 61.85 4.305 ;
        RECT 62.14 4.135 62.31 4.305 ;
        RECT 62.6 4.135 62.77 4.305 ;
        RECT 63.06 4.135 63.23 4.305 ;
        RECT 63.33 4.545 63.5 4.715 ;
        RECT 63.52 4.135 63.69 4.305 ;
        RECT 63.98 4.135 64.15 4.305 ;
        RECT 64.44 4.135 64.61 4.305 ;
        RECT 64.9 4.135 65.07 4.305 ;
        RECT 65.36 4.135 65.53 4.305 ;
        RECT 68.945 4.545 69.115 4.715 ;
        RECT 68.945 4.165 69.115 4.335 ;
        RECT 69.645 4.55 69.815 4.72 ;
        RECT 69.645 4.16 69.815 4.33 ;
        RECT 70.635 4.55 70.805 4.72 ;
        RECT 70.635 4.16 70.805 4.33 ;
        RECT 72.42 4.135 72.59 4.305 ;
        RECT 72.88 4.135 73.05 4.305 ;
        RECT 73.34 4.135 73.51 4.305 ;
        RECT 73.8 4.135 73.97 4.305 ;
        RECT 74.26 4.135 74.43 4.305 ;
        RECT 74.72 4.135 74.89 4.305 ;
        RECT 75.18 4.135 75.35 4.305 ;
        RECT 75.64 4.135 75.81 4.305 ;
        RECT 76.1 4.135 76.27 4.305 ;
        RECT 76.56 4.135 76.73 4.305 ;
        RECT 77.02 4.135 77.19 4.305 ;
        RECT 77.48 4.135 77.65 4.305 ;
        RECT 77.94 4.135 78.11 4.305 ;
        RECT 78.4 4.135 78.57 4.305 ;
        RECT 78.86 4.135 79.03 4.305 ;
        RECT 79.32 4.135 79.49 4.305 ;
        RECT 79.78 4.135 79.95 4.305 ;
        RECT 80.24 4.135 80.41 4.305 ;
        RECT 80.7 4.135 80.87 4.305 ;
        RECT 81.16 4.135 81.33 4.305 ;
        RECT 81.62 4.135 81.79 4.305 ;
        RECT 81.89 4.545 82.06 4.715 ;
        RECT 82.08 4.135 82.25 4.305 ;
        RECT 82.54 4.135 82.71 4.305 ;
        RECT 83 4.135 83.17 4.305 ;
        RECT 83.46 4.135 83.63 4.305 ;
        RECT 83.92 4.135 84.09 4.305 ;
        RECT 87.505 4.545 87.675 4.715 ;
        RECT 87.505 4.165 87.675 4.335 ;
        RECT 88.205 4.55 88.375 4.72 ;
        RECT 88.205 4.16 88.375 4.33 ;
        RECT 89.195 4.55 89.365 4.72 ;
        RECT 89.195 4.16 89.365 4.33 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 73.89 2.415 74.62 2.745 ;
        RECT 55.33 2.415 56.06 2.745 ;
        RECT 36.77 2.415 37.5 2.745 ;
        RECT 18.21 2.415 18.94 2.745 ;
        RECT -0.35 2.415 0.38 2.745 ;
      LAYER li1 ;
        RECT 89.91 0 90.09 0.305 ;
        RECT -5.505 0 90.09 0.3 ;
        RECT 89.115 0 89.285 0.93 ;
        RECT 88.125 0 88.295 0.93 ;
        RECT 71.35 0 87.96 0.305 ;
        RECT 85.385 0 85.555 0.935 ;
        RECT 72.275 0 84.32 1.585 ;
        RECT 83.325 0 83.495 2.085 ;
        RECT 82.365 0 82.535 2.085 ;
        RECT 81.405 0 81.575 2.085 ;
        RECT 80.885 0 81.055 2.085 ;
        RECT 80.605 0 80.8 1.595 ;
        RECT 79.925 0 80.095 2.085 ;
        RECT 78.925 0 79.095 2.085 ;
        RECT 77.965 0 78.135 2.085 ;
        RECT 76.93 0 77.125 1.595 ;
        RECT 76.485 0 76.655 2.085 ;
        RECT 74.565 0 74.825 1.595 ;
        RECT 74.565 0 74.735 2.085 ;
        RECT 73.085 0 73.255 2.085 ;
        RECT 70.555 0 70.725 0.93 ;
        RECT 69.565 0 69.735 0.93 ;
        RECT 52.79 0 69.4 0.305 ;
        RECT 66.825 0 66.995 0.935 ;
        RECT 53.715 0 65.76 1.585 ;
        RECT 64.765 0 64.935 2.085 ;
        RECT 63.805 0 63.975 2.085 ;
        RECT 62.845 0 63.015 2.085 ;
        RECT 62.325 0 62.495 2.085 ;
        RECT 62.045 0 62.24 1.595 ;
        RECT 61.365 0 61.535 2.085 ;
        RECT 60.365 0 60.535 2.085 ;
        RECT 59.405 0 59.575 2.085 ;
        RECT 58.37 0 58.565 1.595 ;
        RECT 57.925 0 58.095 2.085 ;
        RECT 56.005 0 56.265 1.595 ;
        RECT 56.005 0 56.175 2.085 ;
        RECT 54.525 0 54.695 2.085 ;
        RECT 51.995 0 52.165 0.93 ;
        RECT 51.005 0 51.175 0.93 ;
        RECT 34.23 0 50.84 0.305 ;
        RECT 48.265 0 48.435 0.935 ;
        RECT 35.155 0 47.2 1.585 ;
        RECT 46.205 0 46.375 2.085 ;
        RECT 45.245 0 45.415 2.085 ;
        RECT 44.285 0 44.455 2.085 ;
        RECT 43.765 0 43.935 2.085 ;
        RECT 43.485 0 43.68 1.595 ;
        RECT 42.805 0 42.975 2.085 ;
        RECT 41.805 0 41.975 2.085 ;
        RECT 40.845 0 41.015 2.085 ;
        RECT 39.81 0 40.005 1.595 ;
        RECT 39.365 0 39.535 2.085 ;
        RECT 37.445 0 37.705 1.595 ;
        RECT 37.445 0 37.615 2.085 ;
        RECT 35.965 0 36.135 2.085 ;
        RECT 33.435 0 33.605 0.93 ;
        RECT 32.445 0 32.615 0.93 ;
        RECT 15.67 0 32.28 0.305 ;
        RECT 29.705 0 29.875 0.935 ;
        RECT 16.595 0 28.64 1.585 ;
        RECT 27.645 0 27.815 2.085 ;
        RECT 26.685 0 26.855 2.085 ;
        RECT 25.725 0 25.895 2.085 ;
        RECT 25.205 0 25.375 2.085 ;
        RECT 24.925 0 25.12 1.595 ;
        RECT 24.245 0 24.415 2.085 ;
        RECT 23.245 0 23.415 2.085 ;
        RECT 22.285 0 22.455 2.085 ;
        RECT 21.25 0 21.445 1.595 ;
        RECT 20.805 0 20.975 2.085 ;
        RECT 18.885 0 19.145 1.595 ;
        RECT 18.885 0 19.055 2.085 ;
        RECT 17.405 0 17.575 2.085 ;
        RECT 14.875 0 15.045 0.93 ;
        RECT 13.885 0 14.055 0.93 ;
        RECT -5.505 0 13.72 0.305 ;
        RECT 11.145 0 11.315 0.935 ;
        RECT -1.965 0 10.08 1.585 ;
        RECT 9.085 0 9.255 2.085 ;
        RECT 8.125 0 8.295 2.085 ;
        RECT 7.165 0 7.335 2.085 ;
        RECT 6.645 0 6.815 2.085 ;
        RECT 6.365 0 6.56 1.595 ;
        RECT 5.685 0 5.855 2.085 ;
        RECT 4.685 0 4.855 2.085 ;
        RECT 3.725 0 3.895 2.085 ;
        RECT 2.69 0 2.885 1.595 ;
        RECT 2.245 0 2.415 2.085 ;
        RECT 0.325 0 0.585 1.595 ;
        RECT 0.325 0 0.495 2.085 ;
        RECT -1.155 0 -0.985 2.085 ;
        RECT -5.505 8.58 90.09 8.88 ;
        RECT 89.91 8.575 90.09 8.88 ;
        RECT 89.115 7.95 89.285 8.88 ;
        RECT 88.125 7.95 88.295 8.88 ;
        RECT 71.35 8.575 87.96 8.88 ;
        RECT 85.385 7.945 85.555 8.88 ;
        RECT 79.77 7.945 79.94 8.88 ;
        RECT 70.555 7.95 70.725 8.88 ;
        RECT 69.565 7.95 69.735 8.88 ;
        RECT 52.79 8.575 69.4 8.88 ;
        RECT 66.825 7.945 66.995 8.88 ;
        RECT 61.21 7.945 61.38 8.88 ;
        RECT 51.995 7.95 52.165 8.88 ;
        RECT 51.005 7.95 51.175 8.88 ;
        RECT 34.23 8.575 50.84 8.88 ;
        RECT 48.265 7.945 48.435 8.88 ;
        RECT 42.65 7.945 42.82 8.88 ;
        RECT 33.435 7.95 33.605 8.88 ;
        RECT 32.445 7.95 32.615 8.88 ;
        RECT 15.67 8.575 32.28 8.88 ;
        RECT 29.705 7.945 29.875 8.88 ;
        RECT 24.09 7.945 24.26 8.88 ;
        RECT 14.875 7.95 15.045 8.88 ;
        RECT 13.885 7.95 14.055 8.88 ;
        RECT -5.505 8.575 13.72 8.88 ;
        RECT 11.145 7.945 11.315 8.88 ;
        RECT 5.53 7.945 5.7 8.88 ;
        RECT -5.285 7.945 -5.115 8.88 ;
        RECT 80.775 6.075 80.945 8.025 ;
        RECT 80.72 7.855 80.89 8.305 ;
        RECT 80.72 5.015 80.89 6.245 ;
        RECT 75.765 2.495 75.935 2.825 ;
        RECT 73.925 3.055 74.215 3.225 ;
        RECT 73.925 2.575 74.095 3.225 ;
        RECT 73.725 2.575 74.095 2.745 ;
        RECT 62.215 6.075 62.385 8.025 ;
        RECT 62.16 7.855 62.33 8.305 ;
        RECT 62.16 5.015 62.33 6.245 ;
        RECT 57.205 2.495 57.375 2.825 ;
        RECT 55.365 3.055 55.655 3.225 ;
        RECT 55.365 2.575 55.535 3.225 ;
        RECT 55.165 2.575 55.535 2.745 ;
        RECT 43.655 6.075 43.825 8.025 ;
        RECT 43.6 7.855 43.77 8.305 ;
        RECT 43.6 5.015 43.77 6.245 ;
        RECT 38.645 2.495 38.815 2.825 ;
        RECT 36.805 3.055 37.095 3.225 ;
        RECT 36.805 2.575 36.975 3.225 ;
        RECT 36.605 2.575 36.975 2.745 ;
        RECT 25.095 6.075 25.265 8.025 ;
        RECT 25.04 7.855 25.21 8.305 ;
        RECT 25.04 5.015 25.21 6.245 ;
        RECT 20.085 2.495 20.255 2.825 ;
        RECT 18.245 3.055 18.535 3.225 ;
        RECT 18.245 2.575 18.415 3.225 ;
        RECT 18.045 2.575 18.415 2.745 ;
        RECT 6.535 6.075 6.705 8.025 ;
        RECT 6.48 7.855 6.65 8.305 ;
        RECT 6.48 5.015 6.65 6.245 ;
        RECT 1.525 2.495 1.695 2.825 ;
        RECT -0.315 3.055 -0.025 3.225 ;
        RECT -0.315 2.575 -0.145 3.225 ;
        RECT -0.515 2.575 -0.145 2.745 ;
      LAYER met2 ;
        RECT 75.72 2.42 75.98 2.74 ;
        RECT 73.94 2.51 75.98 2.65 ;
        RECT 74.32 1 74.66 1.34 ;
        RECT 74.25 2.395 74.53 2.765 ;
        RECT 74.345 1 74.515 2.765 ;
        RECT 74 2.98 74.26 3.3 ;
        RECT 73.94 2.51 74.08 3.21 ;
        RECT 57.16 2.42 57.42 2.74 ;
        RECT 55.38 2.51 57.42 2.65 ;
        RECT 55.76 1 56.1 1.34 ;
        RECT 55.69 2.395 55.97 2.765 ;
        RECT 55.785 1 55.955 2.765 ;
        RECT 55.44 2.98 55.7 3.3 ;
        RECT 55.38 2.51 55.52 3.21 ;
        RECT 38.6 2.42 38.86 2.74 ;
        RECT 36.82 2.51 38.86 2.65 ;
        RECT 37.2 1 37.54 1.34 ;
        RECT 37.13 2.395 37.41 2.765 ;
        RECT 37.225 1 37.395 2.765 ;
        RECT 36.88 2.98 37.14 3.3 ;
        RECT 36.82 2.51 36.96 3.21 ;
        RECT 20.04 2.42 20.3 2.74 ;
        RECT 18.26 2.51 20.3 2.65 ;
        RECT 18.64 1 18.98 1.34 ;
        RECT 18.57 2.395 18.85 2.765 ;
        RECT 18.665 1 18.835 2.765 ;
        RECT 18.32 2.98 18.58 3.3 ;
        RECT 18.26 2.51 18.4 3.21 ;
        RECT 1.48 2.42 1.74 2.74 ;
        RECT -0.3 2.51 1.74 2.65 ;
        RECT 0.08 1 0.42 1.34 ;
        RECT 0.01 2.395 0.29 2.765 ;
        RECT 0.105 1 0.275 2.765 ;
        RECT -0.24 2.98 0.02 3.3 ;
        RECT -0.3 2.51 -0.16 3.21 ;
      LAYER met1 ;
        RECT 89.91 0 90.09 0.305 ;
        RECT -5.505 0 90.09 0.3 ;
        RECT 71.35 0 87.96 0.305 ;
        RECT 72.275 0 84.32 1.585 ;
        RECT 72.275 0 84.235 1.74 ;
        RECT 52.79 0 69.4 0.305 ;
        RECT 53.715 0 65.76 1.585 ;
        RECT 53.715 0 65.675 1.74 ;
        RECT 34.23 0 50.84 0.305 ;
        RECT 35.155 0 47.2 1.585 ;
        RECT 35.155 0 47.115 1.74 ;
        RECT 15.67 0 32.28 0.305 ;
        RECT 16.595 0 28.64 1.585 ;
        RECT 16.595 0 28.555 1.74 ;
        RECT -5.505 0 13.72 0.305 ;
        RECT -1.965 0 10.08 1.585 ;
        RECT -1.965 0 9.995 1.74 ;
        RECT -5.505 8.58 90.09 8.88 ;
        RECT 89.91 8.575 90.09 8.88 ;
        RECT 71.35 8.575 87.96 8.88 ;
        RECT 80.715 6.285 81.005 6.515 ;
        RECT 80.28 6.315 81.005 6.485 ;
        RECT 80.28 6.315 80.45 8.88 ;
        RECT 52.79 8.575 69.4 8.88 ;
        RECT 62.155 6.285 62.445 6.515 ;
        RECT 61.72 6.315 62.445 6.485 ;
        RECT 61.72 6.315 61.89 8.88 ;
        RECT 34.23 8.575 50.84 8.88 ;
        RECT 43.595 6.285 43.885 6.515 ;
        RECT 43.16 6.315 43.885 6.485 ;
        RECT 43.16 6.315 43.33 8.88 ;
        RECT 15.67 8.575 32.28 8.88 ;
        RECT 25.035 6.285 25.325 6.515 ;
        RECT 24.6 6.315 25.325 6.485 ;
        RECT 24.6 6.315 24.77 8.88 ;
        RECT -5.505 8.575 13.72 8.88 ;
        RECT 6.475 6.285 6.765 6.515 ;
        RECT 6.04 6.315 6.765 6.485 ;
        RECT 6.04 6.315 6.21 8.88 ;
        RECT 75.705 2.37 75.995 2.74 ;
        RECT 74.94 2.37 75.995 2.51 ;
        RECT 73.97 3.01 74.29 3.27 ;
        RECT 57.145 2.37 57.435 2.74 ;
        RECT 56.38 2.37 57.435 2.51 ;
        RECT 55.41 3.01 55.73 3.27 ;
        RECT 38.585 2.37 38.875 2.74 ;
        RECT 37.82 2.37 38.875 2.51 ;
        RECT 36.85 3.01 37.17 3.27 ;
        RECT 20.025 2.37 20.315 2.74 ;
        RECT 19.26 2.37 20.315 2.51 ;
        RECT 18.29 3.01 18.61 3.27 ;
        RECT 1.465 2.37 1.755 2.74 ;
        RECT 0.7 2.37 1.755 2.51 ;
        RECT -0.27 3.01 0.05 3.27 ;
      LAYER via2 ;
        RECT 0.05 2.48 0.25 2.68 ;
        RECT 18.61 2.48 18.81 2.68 ;
        RECT 37.17 2.48 37.37 2.68 ;
        RECT 55.73 2.48 55.93 2.68 ;
        RECT 74.29 2.48 74.49 2.68 ;
      LAYER via1 ;
        RECT -0.185 3.065 -0.035 3.215 ;
        RECT 0.175 1.095 0.325 1.245 ;
        RECT 1.535 2.505 1.685 2.655 ;
        RECT 18.375 3.065 18.525 3.215 ;
        RECT 18.735 1.095 18.885 1.245 ;
        RECT 20.095 2.505 20.245 2.655 ;
        RECT 36.935 3.065 37.085 3.215 ;
        RECT 37.295 1.095 37.445 1.245 ;
        RECT 38.655 2.505 38.805 2.655 ;
        RECT 55.495 3.065 55.645 3.215 ;
        RECT 55.855 1.095 56.005 1.245 ;
        RECT 57.215 2.505 57.365 2.655 ;
        RECT 74.055 3.065 74.205 3.215 ;
        RECT 74.415 1.095 74.565 1.245 ;
        RECT 75.775 2.505 75.925 2.655 ;
      LAYER mcon ;
        RECT -5.205 8.605 -5.035 8.775 ;
        RECT -4.525 8.605 -4.355 8.775 ;
        RECT -3.845 8.605 -3.675 8.775 ;
        RECT -3.165 8.605 -2.995 8.775 ;
        RECT -1.82 1.415 -1.65 1.585 ;
        RECT -1.36 1.415 -1.19 1.585 ;
        RECT -0.9 1.415 -0.73 1.585 ;
        RECT -0.44 1.415 -0.27 1.585 ;
        RECT -0.195 3.055 -0.025 3.225 ;
        RECT 0.02 1.415 0.19 1.585 ;
        RECT 0.48 1.415 0.65 1.585 ;
        RECT 0.94 1.415 1.11 1.585 ;
        RECT 1.4 1.415 1.57 1.585 ;
        RECT 1.525 2.495 1.695 2.665 ;
        RECT 1.86 1.415 2.03 1.585 ;
        RECT 2.32 1.415 2.49 1.585 ;
        RECT 2.78 1.415 2.95 1.585 ;
        RECT 3.24 1.415 3.41 1.585 ;
        RECT 3.7 1.415 3.87 1.585 ;
        RECT 4.16 1.415 4.33 1.585 ;
        RECT 4.62 1.415 4.79 1.585 ;
        RECT 5.08 1.415 5.25 1.585 ;
        RECT 5.54 1.415 5.71 1.585 ;
        RECT 5.61 8.605 5.78 8.775 ;
        RECT 6 1.415 6.17 1.585 ;
        RECT 6.29 8.605 6.46 8.775 ;
        RECT 6.46 1.415 6.63 1.585 ;
        RECT 6.535 6.315 6.705 6.485 ;
        RECT 6.92 1.415 7.09 1.585 ;
        RECT 6.97 8.605 7.14 8.775 ;
        RECT 7.38 1.415 7.55 1.585 ;
        RECT 7.65 8.605 7.82 8.775 ;
        RECT 7.84 1.415 8.01 1.585 ;
        RECT 8.3 1.415 8.47 1.585 ;
        RECT 8.76 1.415 8.93 1.585 ;
        RECT 9.22 1.415 9.39 1.585 ;
        RECT 9.68 1.415 9.85 1.585 ;
        RECT 11.225 8.605 11.395 8.775 ;
        RECT 11.225 0.105 11.395 0.275 ;
        RECT 11.905 8.605 12.075 8.775 ;
        RECT 11.905 0.105 12.075 0.275 ;
        RECT 12.585 8.605 12.755 8.775 ;
        RECT 12.585 0.105 12.755 0.275 ;
        RECT 13.265 8.605 13.435 8.775 ;
        RECT 13.265 0.105 13.435 0.275 ;
        RECT 13.965 8.61 14.135 8.78 ;
        RECT 13.965 0.1 14.135 0.27 ;
        RECT 14.955 8.61 15.125 8.78 ;
        RECT 14.955 0.1 15.125 0.27 ;
        RECT 16.74 1.415 16.91 1.585 ;
        RECT 17.2 1.415 17.37 1.585 ;
        RECT 17.66 1.415 17.83 1.585 ;
        RECT 18.12 1.415 18.29 1.585 ;
        RECT 18.365 3.055 18.535 3.225 ;
        RECT 18.58 1.415 18.75 1.585 ;
        RECT 19.04 1.415 19.21 1.585 ;
        RECT 19.5 1.415 19.67 1.585 ;
        RECT 19.96 1.415 20.13 1.585 ;
        RECT 20.085 2.495 20.255 2.665 ;
        RECT 20.42 1.415 20.59 1.585 ;
        RECT 20.88 1.415 21.05 1.585 ;
        RECT 21.34 1.415 21.51 1.585 ;
        RECT 21.8 1.415 21.97 1.585 ;
        RECT 22.26 1.415 22.43 1.585 ;
        RECT 22.72 1.415 22.89 1.585 ;
        RECT 23.18 1.415 23.35 1.585 ;
        RECT 23.64 1.415 23.81 1.585 ;
        RECT 24.1 1.415 24.27 1.585 ;
        RECT 24.17 8.605 24.34 8.775 ;
        RECT 24.56 1.415 24.73 1.585 ;
        RECT 24.85 8.605 25.02 8.775 ;
        RECT 25.02 1.415 25.19 1.585 ;
        RECT 25.095 6.315 25.265 6.485 ;
        RECT 25.48 1.415 25.65 1.585 ;
        RECT 25.53 8.605 25.7 8.775 ;
        RECT 25.94 1.415 26.11 1.585 ;
        RECT 26.21 8.605 26.38 8.775 ;
        RECT 26.4 1.415 26.57 1.585 ;
        RECT 26.86 1.415 27.03 1.585 ;
        RECT 27.32 1.415 27.49 1.585 ;
        RECT 27.78 1.415 27.95 1.585 ;
        RECT 28.24 1.415 28.41 1.585 ;
        RECT 29.785 8.605 29.955 8.775 ;
        RECT 29.785 0.105 29.955 0.275 ;
        RECT 30.465 8.605 30.635 8.775 ;
        RECT 30.465 0.105 30.635 0.275 ;
        RECT 31.145 8.605 31.315 8.775 ;
        RECT 31.145 0.105 31.315 0.275 ;
        RECT 31.825 8.605 31.995 8.775 ;
        RECT 31.825 0.105 31.995 0.275 ;
        RECT 32.525 8.61 32.695 8.78 ;
        RECT 32.525 0.1 32.695 0.27 ;
        RECT 33.515 8.61 33.685 8.78 ;
        RECT 33.515 0.1 33.685 0.27 ;
        RECT 35.3 1.415 35.47 1.585 ;
        RECT 35.76 1.415 35.93 1.585 ;
        RECT 36.22 1.415 36.39 1.585 ;
        RECT 36.68 1.415 36.85 1.585 ;
        RECT 36.925 3.055 37.095 3.225 ;
        RECT 37.14 1.415 37.31 1.585 ;
        RECT 37.6 1.415 37.77 1.585 ;
        RECT 38.06 1.415 38.23 1.585 ;
        RECT 38.52 1.415 38.69 1.585 ;
        RECT 38.645 2.495 38.815 2.665 ;
        RECT 38.98 1.415 39.15 1.585 ;
        RECT 39.44 1.415 39.61 1.585 ;
        RECT 39.9 1.415 40.07 1.585 ;
        RECT 40.36 1.415 40.53 1.585 ;
        RECT 40.82 1.415 40.99 1.585 ;
        RECT 41.28 1.415 41.45 1.585 ;
        RECT 41.74 1.415 41.91 1.585 ;
        RECT 42.2 1.415 42.37 1.585 ;
        RECT 42.66 1.415 42.83 1.585 ;
        RECT 42.73 8.605 42.9 8.775 ;
        RECT 43.12 1.415 43.29 1.585 ;
        RECT 43.41 8.605 43.58 8.775 ;
        RECT 43.58 1.415 43.75 1.585 ;
        RECT 43.655 6.315 43.825 6.485 ;
        RECT 44.04 1.415 44.21 1.585 ;
        RECT 44.09 8.605 44.26 8.775 ;
        RECT 44.5 1.415 44.67 1.585 ;
        RECT 44.77 8.605 44.94 8.775 ;
        RECT 44.96 1.415 45.13 1.585 ;
        RECT 45.42 1.415 45.59 1.585 ;
        RECT 45.88 1.415 46.05 1.585 ;
        RECT 46.34 1.415 46.51 1.585 ;
        RECT 46.8 1.415 46.97 1.585 ;
        RECT 48.345 8.605 48.515 8.775 ;
        RECT 48.345 0.105 48.515 0.275 ;
        RECT 49.025 8.605 49.195 8.775 ;
        RECT 49.025 0.105 49.195 0.275 ;
        RECT 49.705 8.605 49.875 8.775 ;
        RECT 49.705 0.105 49.875 0.275 ;
        RECT 50.385 8.605 50.555 8.775 ;
        RECT 50.385 0.105 50.555 0.275 ;
        RECT 51.085 8.61 51.255 8.78 ;
        RECT 51.085 0.1 51.255 0.27 ;
        RECT 52.075 8.61 52.245 8.78 ;
        RECT 52.075 0.1 52.245 0.27 ;
        RECT 53.86 1.415 54.03 1.585 ;
        RECT 54.32 1.415 54.49 1.585 ;
        RECT 54.78 1.415 54.95 1.585 ;
        RECT 55.24 1.415 55.41 1.585 ;
        RECT 55.485 3.055 55.655 3.225 ;
        RECT 55.7 1.415 55.87 1.585 ;
        RECT 56.16 1.415 56.33 1.585 ;
        RECT 56.62 1.415 56.79 1.585 ;
        RECT 57.08 1.415 57.25 1.585 ;
        RECT 57.205 2.495 57.375 2.665 ;
        RECT 57.54 1.415 57.71 1.585 ;
        RECT 58 1.415 58.17 1.585 ;
        RECT 58.46 1.415 58.63 1.585 ;
        RECT 58.92 1.415 59.09 1.585 ;
        RECT 59.38 1.415 59.55 1.585 ;
        RECT 59.84 1.415 60.01 1.585 ;
        RECT 60.3 1.415 60.47 1.585 ;
        RECT 60.76 1.415 60.93 1.585 ;
        RECT 61.22 1.415 61.39 1.585 ;
        RECT 61.29 8.605 61.46 8.775 ;
        RECT 61.68 1.415 61.85 1.585 ;
        RECT 61.97 8.605 62.14 8.775 ;
        RECT 62.14 1.415 62.31 1.585 ;
        RECT 62.215 6.315 62.385 6.485 ;
        RECT 62.6 1.415 62.77 1.585 ;
        RECT 62.65 8.605 62.82 8.775 ;
        RECT 63.06 1.415 63.23 1.585 ;
        RECT 63.33 8.605 63.5 8.775 ;
        RECT 63.52 1.415 63.69 1.585 ;
        RECT 63.98 1.415 64.15 1.585 ;
        RECT 64.44 1.415 64.61 1.585 ;
        RECT 64.9 1.415 65.07 1.585 ;
        RECT 65.36 1.415 65.53 1.585 ;
        RECT 66.905 8.605 67.075 8.775 ;
        RECT 66.905 0.105 67.075 0.275 ;
        RECT 67.585 8.605 67.755 8.775 ;
        RECT 67.585 0.105 67.755 0.275 ;
        RECT 68.265 8.605 68.435 8.775 ;
        RECT 68.265 0.105 68.435 0.275 ;
        RECT 68.945 8.605 69.115 8.775 ;
        RECT 68.945 0.105 69.115 0.275 ;
        RECT 69.645 8.61 69.815 8.78 ;
        RECT 69.645 0.1 69.815 0.27 ;
        RECT 70.635 8.61 70.805 8.78 ;
        RECT 70.635 0.1 70.805 0.27 ;
        RECT 72.42 1.415 72.59 1.585 ;
        RECT 72.88 1.415 73.05 1.585 ;
        RECT 73.34 1.415 73.51 1.585 ;
        RECT 73.8 1.415 73.97 1.585 ;
        RECT 74.045 3.055 74.215 3.225 ;
        RECT 74.26 1.415 74.43 1.585 ;
        RECT 74.72 1.415 74.89 1.585 ;
        RECT 75.18 1.415 75.35 1.585 ;
        RECT 75.64 1.415 75.81 1.585 ;
        RECT 75.765 2.495 75.935 2.665 ;
        RECT 76.1 1.415 76.27 1.585 ;
        RECT 76.56 1.415 76.73 1.585 ;
        RECT 77.02 1.415 77.19 1.585 ;
        RECT 77.48 1.415 77.65 1.585 ;
        RECT 77.94 1.415 78.11 1.585 ;
        RECT 78.4 1.415 78.57 1.585 ;
        RECT 78.86 1.415 79.03 1.585 ;
        RECT 79.32 1.415 79.49 1.585 ;
        RECT 79.78 1.415 79.95 1.585 ;
        RECT 79.85 8.605 80.02 8.775 ;
        RECT 80.24 1.415 80.41 1.585 ;
        RECT 80.53 8.605 80.7 8.775 ;
        RECT 80.7 1.415 80.87 1.585 ;
        RECT 80.775 6.315 80.945 6.485 ;
        RECT 81.16 1.415 81.33 1.585 ;
        RECT 81.21 8.605 81.38 8.775 ;
        RECT 81.62 1.415 81.79 1.585 ;
        RECT 81.89 8.605 82.06 8.775 ;
        RECT 82.08 1.415 82.25 1.585 ;
        RECT 82.54 1.415 82.71 1.585 ;
        RECT 83 1.415 83.17 1.585 ;
        RECT 83.46 1.415 83.63 1.585 ;
        RECT 83.92 1.415 84.09 1.585 ;
        RECT 85.465 8.605 85.635 8.775 ;
        RECT 85.465 0.105 85.635 0.275 ;
        RECT 86.145 8.605 86.315 8.775 ;
        RECT 86.145 0.105 86.315 0.275 ;
        RECT 86.825 8.605 86.995 8.775 ;
        RECT 86.825 0.105 86.995 0.275 ;
        RECT 87.505 8.605 87.675 8.775 ;
        RECT 87.505 0.105 87.675 0.275 ;
        RECT 88.205 8.61 88.375 8.78 ;
        RECT 88.205 0.1 88.375 0.27 ;
        RECT 89.195 8.61 89.365 8.78 ;
        RECT 89.195 0.1 89.365 0.27 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 81.58 3.535 82.135 3.865 ;
      RECT 81.58 1.87 81.88 3.865 ;
      RECT 77.645 2.975 78.2 3.305 ;
      RECT 77.9 1.87 78.2 3.305 ;
      RECT 77.9 1.87 81.88 2.17 ;
      RECT 81.05 7.055 81.425 7.425 ;
      RECT 81.05 7.095 82.055 7.395 ;
      RECT 81.755 4.405 82.055 7.395 ;
      RECT 71.925 4.405 82.055 4.705 ;
      RECT 76.43 2.415 76.73 4.705 ;
      RECT 74.995 2.975 75.295 4.705 ;
      RECT 71.925 2.42 72.225 4.705 ;
      RECT 74.965 2.975 75.695 3.305 ;
      RECT 76.405 2.415 77.135 2.745 ;
      RECT 72.855 2.415 73.585 2.745 ;
      RECT 71.925 2.42 73.585 2.72 ;
      RECT 63.02 3.535 63.575 3.865 ;
      RECT 63.02 1.87 63.32 3.865 ;
      RECT 59.085 2.975 59.64 3.305 ;
      RECT 59.34 1.87 59.64 3.305 ;
      RECT 59.34 1.87 63.32 2.17 ;
      RECT 62.49 7.055 62.865 7.425 ;
      RECT 62.49 7.095 63.495 7.395 ;
      RECT 63.195 4.405 63.495 7.395 ;
      RECT 53.365 4.405 63.495 4.705 ;
      RECT 57.87 2.415 58.17 4.705 ;
      RECT 56.435 2.975 56.735 4.705 ;
      RECT 53.365 2.42 53.665 4.705 ;
      RECT 56.405 2.975 57.135 3.305 ;
      RECT 57.845 2.415 58.575 2.745 ;
      RECT 54.295 2.415 55.025 2.745 ;
      RECT 53.365 2.42 55.025 2.72 ;
      RECT 44.46 3.535 45.015 3.865 ;
      RECT 44.46 1.87 44.76 3.865 ;
      RECT 40.525 2.975 41.08 3.305 ;
      RECT 40.78 1.87 41.08 3.305 ;
      RECT 40.78 1.87 44.76 2.17 ;
      RECT 43.93 7.055 44.305 7.425 ;
      RECT 43.93 7.095 44.935 7.395 ;
      RECT 44.635 4.405 44.935 7.395 ;
      RECT 34.805 4.405 44.935 4.705 ;
      RECT 39.31 2.415 39.61 4.705 ;
      RECT 37.875 2.975 38.175 4.705 ;
      RECT 34.805 2.42 35.105 4.705 ;
      RECT 37.845 2.975 38.575 3.305 ;
      RECT 39.285 2.415 40.015 2.745 ;
      RECT 35.735 2.415 36.465 2.745 ;
      RECT 34.805 2.42 36.465 2.72 ;
      RECT 25.9 3.535 26.455 3.865 ;
      RECT 25.9 1.87 26.2 3.865 ;
      RECT 21.965 2.975 22.52 3.305 ;
      RECT 22.22 1.87 22.52 3.305 ;
      RECT 22.22 1.87 26.2 2.17 ;
      RECT 25.37 7.055 25.745 7.425 ;
      RECT 25.37 7.095 26.375 7.395 ;
      RECT 26.075 4.405 26.375 7.395 ;
      RECT 16.245 4.405 26.375 4.705 ;
      RECT 20.75 2.415 21.05 4.705 ;
      RECT 19.315 2.975 19.615 4.705 ;
      RECT 16.245 2.42 16.545 4.705 ;
      RECT 19.285 2.975 20.015 3.305 ;
      RECT 20.725 2.415 21.455 2.745 ;
      RECT 17.175 2.415 17.905 2.745 ;
      RECT 16.245 2.42 17.905 2.72 ;
      RECT 7.34 3.535 7.895 3.865 ;
      RECT 7.34 1.87 7.64 3.865 ;
      RECT 3.405 2.975 3.96 3.305 ;
      RECT 3.66 1.87 3.96 3.305 ;
      RECT 3.66 1.87 7.64 2.17 ;
      RECT 6.81 7.055 7.185 7.425 ;
      RECT 6.81 7.095 7.815 7.395 ;
      RECT 7.515 4.405 7.815 7.395 ;
      RECT -5.505 4.145 -0.245 4.75 ;
      RECT -5.505 4.405 7.815 4.705 ;
      RECT 2.19 2.415 2.49 4.705 ;
      RECT 0.755 2.975 1.055 4.705 ;
      RECT -2.315 2.42 -2.015 4.75 ;
      RECT 0.725 2.975 1.455 3.305 ;
      RECT 2.165 2.415 2.895 2.745 ;
      RECT -1.385 2.415 -0.655 2.745 ;
      RECT -2.315 2.42 -0.655 2.72 ;
      RECT 82.765 1.855 83.495 2.185 ;
      RECT 80.545 3.535 81.275 3.865 ;
      RECT 78.845 3.535 79.575 3.865 ;
      RECT 72.525 3.535 73.255 3.865 ;
      RECT 64.205 1.855 64.935 2.185 ;
      RECT 61.985 3.535 62.715 3.865 ;
      RECT 60.285 3.535 61.015 3.865 ;
      RECT 53.965 3.535 54.695 3.865 ;
      RECT 45.645 1.855 46.375 2.185 ;
      RECT 43.425 3.535 44.155 3.865 ;
      RECT 41.725 3.535 42.455 3.865 ;
      RECT 35.405 3.535 36.135 3.865 ;
      RECT 27.085 1.855 27.815 2.185 ;
      RECT 24.865 3.535 25.595 3.865 ;
      RECT 23.165 3.535 23.895 3.865 ;
      RECT 16.845 3.535 17.575 3.865 ;
      RECT 8.525 1.855 9.255 2.185 ;
      RECT 6.305 3.535 7.035 3.865 ;
      RECT 4.605 3.535 5.335 3.865 ;
      RECT -1.715 3.535 -0.985 3.865 ;
    LAYER via2 ;
      RECT 82.83 1.92 83.03 2.12 ;
      RECT 81.87 3.6 82.07 3.8 ;
      RECT 81.135 7.14 81.335 7.34 ;
      RECT 80.87 3.6 81.07 3.8 ;
      RECT 78.91 3.6 79.11 3.8 ;
      RECT 77.71 3.04 77.91 3.24 ;
      RECT 76.47 2.48 76.67 2.68 ;
      RECT 75.03 3.04 75.23 3.24 ;
      RECT 73.07 2.48 73.27 2.68 ;
      RECT 72.59 3.6 72.79 3.8 ;
      RECT 64.27 1.92 64.47 2.12 ;
      RECT 63.31 3.6 63.51 3.8 ;
      RECT 62.575 7.14 62.775 7.34 ;
      RECT 62.31 3.6 62.51 3.8 ;
      RECT 60.35 3.6 60.55 3.8 ;
      RECT 59.15 3.04 59.35 3.24 ;
      RECT 57.91 2.48 58.11 2.68 ;
      RECT 56.47 3.04 56.67 3.24 ;
      RECT 54.51 2.48 54.71 2.68 ;
      RECT 54.03 3.6 54.23 3.8 ;
      RECT 45.71 1.92 45.91 2.12 ;
      RECT 44.75 3.6 44.95 3.8 ;
      RECT 44.015 7.14 44.215 7.34 ;
      RECT 43.75 3.6 43.95 3.8 ;
      RECT 41.79 3.6 41.99 3.8 ;
      RECT 40.59 3.04 40.79 3.24 ;
      RECT 39.35 2.48 39.55 2.68 ;
      RECT 37.91 3.04 38.11 3.24 ;
      RECT 35.95 2.48 36.15 2.68 ;
      RECT 35.47 3.6 35.67 3.8 ;
      RECT 27.15 1.92 27.35 2.12 ;
      RECT 26.19 3.6 26.39 3.8 ;
      RECT 25.455 7.14 25.655 7.34 ;
      RECT 25.19 3.6 25.39 3.8 ;
      RECT 23.23 3.6 23.43 3.8 ;
      RECT 22.03 3.04 22.23 3.24 ;
      RECT 20.79 2.48 20.99 2.68 ;
      RECT 19.35 3.04 19.55 3.24 ;
      RECT 17.39 2.48 17.59 2.68 ;
      RECT 16.91 3.6 17.11 3.8 ;
      RECT 8.59 1.92 8.79 2.12 ;
      RECT 7.63 3.6 7.83 3.8 ;
      RECT 6.895 7.14 7.095 7.34 ;
      RECT 6.63 3.6 6.83 3.8 ;
      RECT 4.67 3.6 4.87 3.8 ;
      RECT 3.47 3.04 3.67 3.24 ;
      RECT 2.23 2.48 2.43 2.68 ;
      RECT 0.79 3.04 0.99 3.24 ;
      RECT -1.17 2.48 -0.97 2.68 ;
      RECT -1.65 3.6 -1.45 3.8 ;
    LAYER met2 ;
      RECT -4.275 8.4 89.72 8.57 ;
      RECT 89.55 7.275 89.72 8.57 ;
      RECT -4.275 6.255 -4.105 8.57 ;
      RECT 89.52 7.275 89.87 7.625 ;
      RECT -4.34 6.255 -4.05 6.605 ;
      RECT 86.36 6.22 86.68 6.545 ;
      RECT 86.39 5.695 86.56 6.545 ;
      RECT 86.39 5.695 86.565 6.045 ;
      RECT 86.39 5.695 87.365 5.87 ;
      RECT 87.19 1.965 87.365 5.87 ;
      RECT 87.135 1.965 87.485 2.315 ;
      RECT 87.16 6.655 87.485 6.98 ;
      RECT 86.045 6.745 87.485 6.915 ;
      RECT 86.045 2.395 86.205 6.915 ;
      RECT 86.36 2.365 86.68 2.685 ;
      RECT 86.045 2.395 86.68 2.565 ;
      RECT 80.88 4.135 85.015 4.325 ;
      RECT 84.845 3.145 85.015 4.325 ;
      RECT 84.825 3.15 85.015 4.325 ;
      RECT 80.88 3.515 81.07 4.325 ;
      RECT 80.83 3.515 81.11 3.885 ;
      RECT 84.755 3.15 85.095 3.5 ;
      RECT 70.935 6.655 71.285 7.005 ;
      RECT 81.72 6.61 82.07 6.96 ;
      RECT 70.935 6.685 82.07 6.885 ;
      RECT 81.36 2.98 81.62 3.3 ;
      RECT 81.42 1.86 81.56 3.3 ;
      RECT 81.36 1.86 81.62 2.18 ;
      RECT 80.36 3.54 80.62 3.86 ;
      RECT 80.36 2.955 80.56 3.86 ;
      RECT 80.3 1.86 80.44 3.49 ;
      RECT 80.3 2.955 80.8 3.325 ;
      RECT 80.24 1.86 80.5 2.18 ;
      RECT 79.88 3.54 80.14 3.86 ;
      RECT 79.94 1.95 80.08 3.86 ;
      RECT 79.64 1.95 80.08 2.18 ;
      RECT 79.64 1.86 79.9 2.18 ;
      RECT 79.4 2.42 79.66 2.74 ;
      RECT 78.82 2.51 79.66 2.65 ;
      RECT 78.82 1.57 78.96 2.65 ;
      RECT 75.48 1.86 75.74 2.18 ;
      RECT 75.48 1.95 76.52 2.09 ;
      RECT 76.38 1.57 76.52 2.09 ;
      RECT 76.38 1.57 78.96 1.71 ;
      RECT 78.87 3.515 79.15 3.885 ;
      RECT 78.94 3.07 79.08 3.885 ;
      RECT 78.75 2.955 79.03 3.325 ;
      RECT 78.46 3.07 79.08 3.21 ;
      RECT 78.46 1.86 78.6 3.21 ;
      RECT 78.4 1.86 78.66 2.18 ;
      RECT 77.67 2.955 77.95 3.325 ;
      RECT 77.74 1.86 77.88 3.325 ;
      RECT 77.68 1.86 77.94 2.18 ;
      RECT 77.32 3.54 77.58 3.86 ;
      RECT 77.38 1.95 77.52 3.86 ;
      RECT 76.96 1.86 77.22 2.18 ;
      RECT 76.96 1.95 77.52 2.09 ;
      RECT 74.99 2.955 75.27 3.325 ;
      RECT 76.96 2.98 77.22 3.3 ;
      RECT 74.64 2.98 75.27 3.3 ;
      RECT 74.64 3.07 77.22 3.21 ;
      RECT 76.43 2.395 76.71 2.765 ;
      RECT 76.43 2.42 76.96 2.74 ;
      RECT 73.52 2.98 73.78 3.3 ;
      RECT 73.58 1.86 73.72 3.3 ;
      RECT 73.52 1.86 73.78 2.18 ;
      RECT 72.55 3.515 72.83 3.885 ;
      RECT 72.56 3.26 72.82 3.885 ;
      RECT 67.8 6.22 68.12 6.545 ;
      RECT 67.83 5.695 68 6.545 ;
      RECT 67.83 5.695 68.005 6.045 ;
      RECT 67.83 5.695 68.805 5.87 ;
      RECT 68.63 1.965 68.805 5.87 ;
      RECT 68.575 1.965 68.925 2.315 ;
      RECT 68.6 6.655 68.925 6.98 ;
      RECT 67.485 6.745 68.925 6.915 ;
      RECT 67.485 2.395 67.645 6.915 ;
      RECT 67.8 2.365 68.12 2.685 ;
      RECT 67.485 2.395 68.12 2.565 ;
      RECT 62.32 4.135 66.455 4.325 ;
      RECT 66.285 3.145 66.455 4.325 ;
      RECT 66.265 3.15 66.455 4.325 ;
      RECT 62.32 3.515 62.51 4.325 ;
      RECT 62.27 3.515 62.55 3.885 ;
      RECT 66.195 3.15 66.535 3.5 ;
      RECT 52.375 6.655 52.725 7.005 ;
      RECT 63.16 6.61 63.51 6.96 ;
      RECT 52.375 6.685 63.51 6.885 ;
      RECT 62.8 2.98 63.06 3.3 ;
      RECT 62.86 1.86 63 3.3 ;
      RECT 62.8 1.86 63.06 2.18 ;
      RECT 61.8 3.54 62.06 3.86 ;
      RECT 61.8 2.955 62 3.86 ;
      RECT 61.74 1.86 61.88 3.49 ;
      RECT 61.74 2.955 62.24 3.325 ;
      RECT 61.68 1.86 61.94 2.18 ;
      RECT 61.32 3.54 61.58 3.86 ;
      RECT 61.38 1.95 61.52 3.86 ;
      RECT 61.08 1.95 61.52 2.18 ;
      RECT 61.08 1.86 61.34 2.18 ;
      RECT 60.84 2.42 61.1 2.74 ;
      RECT 60.26 2.51 61.1 2.65 ;
      RECT 60.26 1.57 60.4 2.65 ;
      RECT 56.92 1.86 57.18 2.18 ;
      RECT 56.92 1.95 57.96 2.09 ;
      RECT 57.82 1.57 57.96 2.09 ;
      RECT 57.82 1.57 60.4 1.71 ;
      RECT 60.31 3.515 60.59 3.885 ;
      RECT 60.38 3.07 60.52 3.885 ;
      RECT 60.19 2.955 60.47 3.325 ;
      RECT 59.9 3.07 60.52 3.21 ;
      RECT 59.9 1.86 60.04 3.21 ;
      RECT 59.84 1.86 60.1 2.18 ;
      RECT 59.11 2.955 59.39 3.325 ;
      RECT 59.18 1.86 59.32 3.325 ;
      RECT 59.12 1.86 59.38 2.18 ;
      RECT 58.76 3.54 59.02 3.86 ;
      RECT 58.82 1.95 58.96 3.86 ;
      RECT 58.4 1.86 58.66 2.18 ;
      RECT 58.4 1.95 58.96 2.09 ;
      RECT 56.43 2.955 56.71 3.325 ;
      RECT 58.4 2.98 58.66 3.3 ;
      RECT 56.08 2.98 56.71 3.3 ;
      RECT 56.08 3.07 58.66 3.21 ;
      RECT 57.87 2.395 58.15 2.765 ;
      RECT 57.87 2.42 58.4 2.74 ;
      RECT 54.96 2.98 55.22 3.3 ;
      RECT 55.02 1.86 55.16 3.3 ;
      RECT 54.96 1.86 55.22 2.18 ;
      RECT 53.99 3.515 54.27 3.885 ;
      RECT 54 3.26 54.26 3.885 ;
      RECT 49.24 6.22 49.56 6.545 ;
      RECT 49.27 5.695 49.44 6.545 ;
      RECT 49.27 5.695 49.445 6.045 ;
      RECT 49.27 5.695 50.245 5.87 ;
      RECT 50.07 1.965 50.245 5.87 ;
      RECT 50.015 1.965 50.365 2.315 ;
      RECT 50.04 6.655 50.365 6.98 ;
      RECT 48.925 6.745 50.365 6.915 ;
      RECT 48.925 2.395 49.085 6.915 ;
      RECT 49.24 2.365 49.56 2.685 ;
      RECT 48.925 2.395 49.56 2.565 ;
      RECT 43.76 4.135 47.895 4.325 ;
      RECT 47.725 3.145 47.895 4.325 ;
      RECT 47.705 3.15 47.895 4.325 ;
      RECT 43.76 3.515 43.95 4.325 ;
      RECT 43.71 3.515 43.99 3.885 ;
      RECT 47.635 3.15 47.975 3.5 ;
      RECT 33.86 6.66 34.21 7.01 ;
      RECT 44.6 6.615 44.95 6.965 ;
      RECT 33.86 6.69 44.95 6.89 ;
      RECT 44.24 2.98 44.5 3.3 ;
      RECT 44.3 1.86 44.44 3.3 ;
      RECT 44.24 1.86 44.5 2.18 ;
      RECT 43.24 3.54 43.5 3.86 ;
      RECT 43.24 2.955 43.44 3.86 ;
      RECT 43.18 1.86 43.32 3.49 ;
      RECT 43.18 2.955 43.68 3.325 ;
      RECT 43.12 1.86 43.38 2.18 ;
      RECT 42.76 3.54 43.02 3.86 ;
      RECT 42.82 1.95 42.96 3.86 ;
      RECT 42.52 1.95 42.96 2.18 ;
      RECT 42.52 1.86 42.78 2.18 ;
      RECT 42.28 2.42 42.54 2.74 ;
      RECT 41.7 2.51 42.54 2.65 ;
      RECT 41.7 1.57 41.84 2.65 ;
      RECT 38.36 1.86 38.62 2.18 ;
      RECT 38.36 1.95 39.4 2.09 ;
      RECT 39.26 1.57 39.4 2.09 ;
      RECT 39.26 1.57 41.84 1.71 ;
      RECT 41.75 3.515 42.03 3.885 ;
      RECT 41.82 3.07 41.96 3.885 ;
      RECT 41.63 2.955 41.91 3.325 ;
      RECT 41.34 3.07 41.96 3.21 ;
      RECT 41.34 1.86 41.48 3.21 ;
      RECT 41.28 1.86 41.54 2.18 ;
      RECT 40.55 2.955 40.83 3.325 ;
      RECT 40.62 1.86 40.76 3.325 ;
      RECT 40.56 1.86 40.82 2.18 ;
      RECT 40.2 3.54 40.46 3.86 ;
      RECT 40.26 1.95 40.4 3.86 ;
      RECT 39.84 1.86 40.1 2.18 ;
      RECT 39.84 1.95 40.4 2.09 ;
      RECT 37.87 2.955 38.15 3.325 ;
      RECT 39.84 2.98 40.1 3.3 ;
      RECT 37.52 2.98 38.15 3.3 ;
      RECT 37.52 3.07 40.1 3.21 ;
      RECT 39.31 2.395 39.59 2.765 ;
      RECT 39.31 2.42 39.84 2.74 ;
      RECT 36.4 2.98 36.66 3.3 ;
      RECT 36.46 1.86 36.6 3.3 ;
      RECT 36.4 1.86 36.66 2.18 ;
      RECT 35.43 3.515 35.71 3.885 ;
      RECT 35.44 3.26 35.7 3.885 ;
      RECT 30.68 6.22 31 6.545 ;
      RECT 30.71 5.695 30.88 6.545 ;
      RECT 30.71 5.695 30.885 6.045 ;
      RECT 30.71 5.695 31.685 5.87 ;
      RECT 31.51 1.965 31.685 5.87 ;
      RECT 31.455 1.965 31.805 2.315 ;
      RECT 31.48 6.655 31.805 6.98 ;
      RECT 30.365 6.745 31.805 6.915 ;
      RECT 30.365 2.395 30.525 6.915 ;
      RECT 30.68 2.365 31 2.685 ;
      RECT 30.365 2.395 31 2.565 ;
      RECT 25.2 4.135 29.335 4.325 ;
      RECT 29.165 3.145 29.335 4.325 ;
      RECT 29.145 3.15 29.335 4.325 ;
      RECT 25.2 3.515 25.39 4.325 ;
      RECT 25.15 3.515 25.43 3.885 ;
      RECT 29.075 3.15 29.415 3.5 ;
      RECT 15.3 6.655 15.65 7.005 ;
      RECT 26.045 6.61 26.395 6.96 ;
      RECT 15.3 6.685 26.395 6.885 ;
      RECT 25.68 2.98 25.94 3.3 ;
      RECT 25.74 1.86 25.88 3.3 ;
      RECT 25.68 1.86 25.94 2.18 ;
      RECT 24.68 3.54 24.94 3.86 ;
      RECT 24.68 2.955 24.88 3.86 ;
      RECT 24.62 1.86 24.76 3.49 ;
      RECT 24.62 2.955 25.12 3.325 ;
      RECT 24.56 1.86 24.82 2.18 ;
      RECT 24.2 3.54 24.46 3.86 ;
      RECT 24.26 1.95 24.4 3.86 ;
      RECT 23.96 1.95 24.4 2.18 ;
      RECT 23.96 1.86 24.22 2.18 ;
      RECT 23.72 2.42 23.98 2.74 ;
      RECT 23.14 2.51 23.98 2.65 ;
      RECT 23.14 1.57 23.28 2.65 ;
      RECT 19.8 1.86 20.06 2.18 ;
      RECT 19.8 1.95 20.84 2.09 ;
      RECT 20.7 1.57 20.84 2.09 ;
      RECT 20.7 1.57 23.28 1.71 ;
      RECT 23.19 3.515 23.47 3.885 ;
      RECT 23.26 3.07 23.4 3.885 ;
      RECT 23.07 2.955 23.35 3.325 ;
      RECT 22.78 3.07 23.4 3.21 ;
      RECT 22.78 1.86 22.92 3.21 ;
      RECT 22.72 1.86 22.98 2.18 ;
      RECT 21.99 2.955 22.27 3.325 ;
      RECT 22.06 1.86 22.2 3.325 ;
      RECT 22 1.86 22.26 2.18 ;
      RECT 21.64 3.54 21.9 3.86 ;
      RECT 21.7 1.95 21.84 3.86 ;
      RECT 21.28 1.86 21.54 2.18 ;
      RECT 21.28 1.95 21.84 2.09 ;
      RECT 19.31 2.955 19.59 3.325 ;
      RECT 21.28 2.98 21.54 3.3 ;
      RECT 18.96 2.98 19.59 3.3 ;
      RECT 18.96 3.07 21.54 3.21 ;
      RECT 20.75 2.395 21.03 2.765 ;
      RECT 20.75 2.42 21.28 2.74 ;
      RECT 17.84 2.98 18.1 3.3 ;
      RECT 17.9 1.86 18.04 3.3 ;
      RECT 17.84 1.86 18.1 2.18 ;
      RECT 16.87 3.515 17.15 3.885 ;
      RECT 16.88 3.26 17.14 3.885 ;
      RECT 12.12 6.22 12.44 6.545 ;
      RECT 12.15 5.695 12.32 6.545 ;
      RECT 12.15 5.695 12.325 6.045 ;
      RECT 12.15 5.695 13.125 5.87 ;
      RECT 12.95 1.965 13.125 5.87 ;
      RECT 12.895 1.965 13.245 2.315 ;
      RECT 12.92 6.655 13.245 6.98 ;
      RECT 11.805 6.745 13.245 6.915 ;
      RECT 11.805 2.395 11.965 6.915 ;
      RECT 12.12 2.365 12.44 2.685 ;
      RECT 11.805 2.395 12.44 2.565 ;
      RECT 6.64 4.135 10.775 4.325 ;
      RECT 10.605 3.145 10.775 4.325 ;
      RECT 10.585 3.15 10.775 4.325 ;
      RECT 6.64 3.515 6.83 4.325 ;
      RECT 6.59 3.515 6.87 3.885 ;
      RECT 10.515 3.15 10.855 3.5 ;
      RECT -3.965 6.995 -3.675 7.345 ;
      RECT -3.965 7.05 -2.65 7.22 ;
      RECT -2.82 6.685 -2.65 7.22 ;
      RECT 7.485 6.605 7.835 6.955 ;
      RECT -2.82 6.685 7.835 6.855 ;
      RECT 7.12 2.98 7.38 3.3 ;
      RECT 7.18 1.86 7.32 3.3 ;
      RECT 7.12 1.86 7.38 2.18 ;
      RECT 6.12 3.54 6.38 3.86 ;
      RECT 6.12 2.955 6.32 3.86 ;
      RECT 6.06 1.86 6.2 3.49 ;
      RECT 6.06 2.955 6.56 3.325 ;
      RECT 6 1.86 6.26 2.18 ;
      RECT 5.64 3.54 5.9 3.86 ;
      RECT 5.7 1.95 5.84 3.86 ;
      RECT 5.4 1.95 5.84 2.18 ;
      RECT 5.4 1.86 5.66 2.18 ;
      RECT 5.16 2.42 5.42 2.74 ;
      RECT 4.58 2.51 5.42 2.65 ;
      RECT 4.58 1.57 4.72 2.65 ;
      RECT 1.24 1.86 1.5 2.18 ;
      RECT 1.24 1.95 2.28 2.09 ;
      RECT 2.14 1.57 2.28 2.09 ;
      RECT 2.14 1.57 4.72 1.71 ;
      RECT 4.63 3.515 4.91 3.885 ;
      RECT 4.7 3.07 4.84 3.885 ;
      RECT 4.51 2.955 4.79 3.325 ;
      RECT 4.22 3.07 4.84 3.21 ;
      RECT 4.22 1.86 4.36 3.21 ;
      RECT 4.16 1.86 4.42 2.18 ;
      RECT 3.43 2.955 3.71 3.325 ;
      RECT 3.5 1.86 3.64 3.325 ;
      RECT 3.44 1.86 3.7 2.18 ;
      RECT 3.08 3.54 3.34 3.86 ;
      RECT 3.14 1.95 3.28 3.86 ;
      RECT 2.72 1.86 2.98 2.18 ;
      RECT 2.72 1.95 3.28 2.09 ;
      RECT 0.75 2.955 1.03 3.325 ;
      RECT 2.72 2.98 2.98 3.3 ;
      RECT 0.4 2.98 1.03 3.3 ;
      RECT 0.4 3.07 2.98 3.21 ;
      RECT 2.19 2.395 2.47 2.765 ;
      RECT 2.19 2.42 2.72 2.74 ;
      RECT -0.72 2.98 -0.46 3.3 ;
      RECT -0.66 1.86 -0.52 3.3 ;
      RECT -0.72 1.86 -0.46 2.18 ;
      RECT -1.69 3.515 -1.41 3.885 ;
      RECT -1.68 3.26 -1.42 3.885 ;
      RECT 82.79 1.835 83.07 2.205 ;
      RECT 81.83 3.515 82.11 3.885 ;
      RECT 81.05 7.055 81.425 7.425 ;
      RECT 73.03 2.395 73.31 2.765 ;
      RECT 64.23 1.835 64.51 2.205 ;
      RECT 63.27 3.515 63.55 3.885 ;
      RECT 62.49 7.055 62.865 7.425 ;
      RECT 54.47 2.395 54.75 2.765 ;
      RECT 45.67 1.835 45.95 2.205 ;
      RECT 44.71 3.515 44.99 3.885 ;
      RECT 43.93 7.055 44.305 7.425 ;
      RECT 35.91 2.395 36.19 2.765 ;
      RECT 27.11 1.835 27.39 2.205 ;
      RECT 26.15 3.515 26.43 3.885 ;
      RECT 25.37 7.055 25.745 7.425 ;
      RECT 17.35 2.395 17.63 2.765 ;
      RECT 8.55 1.835 8.83 2.205 ;
      RECT 7.59 3.515 7.87 3.885 ;
      RECT 6.81 7.055 7.185 7.425 ;
      RECT -1.21 2.395 -0.93 2.765 ;
    LAYER via1 ;
      RECT 89.62 7.375 89.77 7.525 ;
      RECT 87.25 6.74 87.4 6.89 ;
      RECT 87.235 2.065 87.385 2.215 ;
      RECT 86.445 2.45 86.595 2.6 ;
      RECT 86.445 6.325 86.595 6.475 ;
      RECT 84.855 3.25 85.005 3.4 ;
      RECT 82.855 1.945 83.005 2.095 ;
      RECT 81.895 3.625 82.045 3.775 ;
      RECT 81.82 6.71 81.97 6.86 ;
      RECT 81.415 1.945 81.565 2.095 ;
      RECT 81.415 3.065 81.565 3.215 ;
      RECT 81.16 7.165 81.31 7.315 ;
      RECT 80.895 3.625 81.045 3.775 ;
      RECT 80.415 3.625 80.565 3.775 ;
      RECT 80.295 1.945 80.445 2.095 ;
      RECT 79.935 3.625 80.085 3.775 ;
      RECT 79.695 1.945 79.845 2.095 ;
      RECT 79.455 2.505 79.605 2.655 ;
      RECT 78.935 3.625 79.085 3.775 ;
      RECT 78.455 1.945 78.605 2.095 ;
      RECT 77.735 1.945 77.885 2.095 ;
      RECT 77.735 3.065 77.885 3.215 ;
      RECT 77.375 3.625 77.525 3.775 ;
      RECT 77.015 1.945 77.165 2.095 ;
      RECT 77.015 3.065 77.165 3.215 ;
      RECT 76.755 2.505 76.905 2.655 ;
      RECT 75.535 1.945 75.685 2.095 ;
      RECT 74.695 3.065 74.845 3.215 ;
      RECT 73.575 1.945 73.725 2.095 ;
      RECT 73.575 3.065 73.725 3.215 ;
      RECT 73.095 2.505 73.245 2.655 ;
      RECT 72.615 3.345 72.765 3.495 ;
      RECT 71.035 6.755 71.185 6.905 ;
      RECT 68.69 6.74 68.84 6.89 ;
      RECT 68.675 2.065 68.825 2.215 ;
      RECT 67.885 2.45 68.035 2.6 ;
      RECT 67.885 6.325 68.035 6.475 ;
      RECT 66.295 3.25 66.445 3.4 ;
      RECT 64.295 1.945 64.445 2.095 ;
      RECT 63.335 3.625 63.485 3.775 ;
      RECT 63.26 6.71 63.41 6.86 ;
      RECT 62.855 1.945 63.005 2.095 ;
      RECT 62.855 3.065 63.005 3.215 ;
      RECT 62.6 7.165 62.75 7.315 ;
      RECT 62.335 3.625 62.485 3.775 ;
      RECT 61.855 3.625 62.005 3.775 ;
      RECT 61.735 1.945 61.885 2.095 ;
      RECT 61.375 3.625 61.525 3.775 ;
      RECT 61.135 1.945 61.285 2.095 ;
      RECT 60.895 2.505 61.045 2.655 ;
      RECT 60.375 3.625 60.525 3.775 ;
      RECT 59.895 1.945 60.045 2.095 ;
      RECT 59.175 1.945 59.325 2.095 ;
      RECT 59.175 3.065 59.325 3.215 ;
      RECT 58.815 3.625 58.965 3.775 ;
      RECT 58.455 1.945 58.605 2.095 ;
      RECT 58.455 3.065 58.605 3.215 ;
      RECT 58.195 2.505 58.345 2.655 ;
      RECT 56.975 1.945 57.125 2.095 ;
      RECT 56.135 3.065 56.285 3.215 ;
      RECT 55.015 1.945 55.165 2.095 ;
      RECT 55.015 3.065 55.165 3.215 ;
      RECT 54.535 2.505 54.685 2.655 ;
      RECT 54.055 3.345 54.205 3.495 ;
      RECT 52.475 6.755 52.625 6.905 ;
      RECT 50.13 6.74 50.28 6.89 ;
      RECT 50.115 2.065 50.265 2.215 ;
      RECT 49.325 2.45 49.475 2.6 ;
      RECT 49.325 6.325 49.475 6.475 ;
      RECT 47.735 3.25 47.885 3.4 ;
      RECT 45.735 1.945 45.885 2.095 ;
      RECT 44.775 3.625 44.925 3.775 ;
      RECT 44.7 6.715 44.85 6.865 ;
      RECT 44.295 1.945 44.445 2.095 ;
      RECT 44.295 3.065 44.445 3.215 ;
      RECT 44.04 7.165 44.19 7.315 ;
      RECT 43.775 3.625 43.925 3.775 ;
      RECT 43.295 3.625 43.445 3.775 ;
      RECT 43.175 1.945 43.325 2.095 ;
      RECT 42.815 3.625 42.965 3.775 ;
      RECT 42.575 1.945 42.725 2.095 ;
      RECT 42.335 2.505 42.485 2.655 ;
      RECT 41.815 3.625 41.965 3.775 ;
      RECT 41.335 1.945 41.485 2.095 ;
      RECT 40.615 1.945 40.765 2.095 ;
      RECT 40.615 3.065 40.765 3.215 ;
      RECT 40.255 3.625 40.405 3.775 ;
      RECT 39.895 1.945 40.045 2.095 ;
      RECT 39.895 3.065 40.045 3.215 ;
      RECT 39.635 2.505 39.785 2.655 ;
      RECT 38.415 1.945 38.565 2.095 ;
      RECT 37.575 3.065 37.725 3.215 ;
      RECT 36.455 1.945 36.605 2.095 ;
      RECT 36.455 3.065 36.605 3.215 ;
      RECT 35.975 2.505 36.125 2.655 ;
      RECT 35.495 3.345 35.645 3.495 ;
      RECT 33.96 6.76 34.11 6.91 ;
      RECT 31.57 6.74 31.72 6.89 ;
      RECT 31.555 2.065 31.705 2.215 ;
      RECT 30.765 2.45 30.915 2.6 ;
      RECT 30.765 6.325 30.915 6.475 ;
      RECT 29.175 3.25 29.325 3.4 ;
      RECT 27.175 1.945 27.325 2.095 ;
      RECT 26.215 3.625 26.365 3.775 ;
      RECT 26.145 6.71 26.295 6.86 ;
      RECT 25.735 1.945 25.885 2.095 ;
      RECT 25.735 3.065 25.885 3.215 ;
      RECT 25.48 7.165 25.63 7.315 ;
      RECT 25.215 3.625 25.365 3.775 ;
      RECT 24.735 3.625 24.885 3.775 ;
      RECT 24.615 1.945 24.765 2.095 ;
      RECT 24.255 3.625 24.405 3.775 ;
      RECT 24.015 1.945 24.165 2.095 ;
      RECT 23.775 2.505 23.925 2.655 ;
      RECT 23.255 3.625 23.405 3.775 ;
      RECT 22.775 1.945 22.925 2.095 ;
      RECT 22.055 1.945 22.205 2.095 ;
      RECT 22.055 3.065 22.205 3.215 ;
      RECT 21.695 3.625 21.845 3.775 ;
      RECT 21.335 1.945 21.485 2.095 ;
      RECT 21.335 3.065 21.485 3.215 ;
      RECT 21.075 2.505 21.225 2.655 ;
      RECT 19.855 1.945 20.005 2.095 ;
      RECT 19.015 3.065 19.165 3.215 ;
      RECT 17.895 1.945 18.045 2.095 ;
      RECT 17.895 3.065 18.045 3.215 ;
      RECT 17.415 2.505 17.565 2.655 ;
      RECT 16.935 3.345 17.085 3.495 ;
      RECT 15.4 6.755 15.55 6.905 ;
      RECT 13.01 6.74 13.16 6.89 ;
      RECT 12.995 2.065 13.145 2.215 ;
      RECT 12.205 2.45 12.355 2.6 ;
      RECT 12.205 6.325 12.355 6.475 ;
      RECT 10.615 3.25 10.765 3.4 ;
      RECT 8.615 1.945 8.765 2.095 ;
      RECT 7.655 3.625 7.805 3.775 ;
      RECT 7.585 6.705 7.735 6.855 ;
      RECT 7.175 1.945 7.325 2.095 ;
      RECT 7.175 3.065 7.325 3.215 ;
      RECT 6.92 7.165 7.07 7.315 ;
      RECT 6.655 3.625 6.805 3.775 ;
      RECT 6.175 3.625 6.325 3.775 ;
      RECT 6.055 1.945 6.205 2.095 ;
      RECT 5.695 3.625 5.845 3.775 ;
      RECT 5.455 1.945 5.605 2.095 ;
      RECT 5.215 2.505 5.365 2.655 ;
      RECT 4.695 3.625 4.845 3.775 ;
      RECT 4.215 1.945 4.365 2.095 ;
      RECT 3.495 1.945 3.645 2.095 ;
      RECT 3.495 3.065 3.645 3.215 ;
      RECT 3.135 3.625 3.285 3.775 ;
      RECT 2.775 1.945 2.925 2.095 ;
      RECT 2.775 3.065 2.925 3.215 ;
      RECT 2.515 2.505 2.665 2.655 ;
      RECT 1.295 1.945 1.445 2.095 ;
      RECT 0.455 3.065 0.605 3.215 ;
      RECT -0.665 1.945 -0.515 2.095 ;
      RECT -0.665 3.065 -0.515 3.215 ;
      RECT -1.145 2.505 -0.995 2.655 ;
      RECT -1.625 3.345 -1.475 3.495 ;
      RECT -3.895 7.095 -3.745 7.245 ;
      RECT -4.27 6.355 -4.12 6.505 ;
    LAYER met1 ;
      RECT 89.485 7.77 89.775 8 ;
      RECT 89.545 6.29 89.715 8 ;
      RECT 89.52 7.275 89.87 7.625 ;
      RECT 89.485 6.29 89.775 6.52 ;
      RECT 89.08 2.395 89.185 2.965 ;
      RECT 89.08 2.73 89.405 2.96 ;
      RECT 89.08 2.76 89.575 2.93 ;
      RECT 89.08 2.395 89.27 2.96 ;
      RECT 88.495 2.36 88.785 2.59 ;
      RECT 88.495 2.395 89.27 2.565 ;
      RECT 88.555 0.88 88.725 2.59 ;
      RECT 88.495 0.88 88.785 1.11 ;
      RECT 88.495 7.77 88.785 8 ;
      RECT 88.555 6.29 88.725 8 ;
      RECT 88.495 6.29 88.785 6.52 ;
      RECT 88.495 6.325 89.35 6.485 ;
      RECT 89.18 5.92 89.35 6.485 ;
      RECT 88.495 6.32 88.89 6.485 ;
      RECT 89.115 5.92 89.405 6.15 ;
      RECT 89.115 5.95 89.575 6.12 ;
      RECT 88.125 2.73 88.415 2.96 ;
      RECT 88.125 2.76 88.585 2.93 ;
      RECT 88.19 1.655 88.355 2.96 ;
      RECT 86.705 1.625 86.995 1.855 ;
      RECT 86.705 1.655 88.355 1.825 ;
      RECT 86.765 0.885 86.935 1.855 ;
      RECT 86.705 0.885 86.995 1.115 ;
      RECT 86.705 7.765 86.995 7.995 ;
      RECT 86.765 7.025 86.935 7.995 ;
      RECT 86.765 7.12 88.355 7.29 ;
      RECT 88.185 5.92 88.355 7.29 ;
      RECT 86.705 7.025 86.995 7.255 ;
      RECT 88.125 5.92 88.415 6.15 ;
      RECT 88.125 5.95 88.585 6.12 ;
      RECT 84.755 3.15 85.095 3.5 ;
      RECT 84.845 2.025 85.015 3.5 ;
      RECT 87.135 1.965 87.485 2.315 ;
      RECT 84.845 2.025 87.485 2.195 ;
      RECT 87.16 6.655 87.485 6.98 ;
      RECT 81.72 6.61 82.07 6.96 ;
      RECT 87.135 6.655 87.485 6.885 ;
      RECT 81.52 6.655 82.07 6.885 ;
      RECT 81.35 6.685 87.485 6.855 ;
      RECT 86.36 2.365 86.68 2.685 ;
      RECT 86.33 2.365 86.68 2.595 ;
      RECT 86.16 2.395 86.68 2.565 ;
      RECT 86.36 6.255 86.68 6.545 ;
      RECT 86.33 6.285 86.68 6.515 ;
      RECT 86.16 6.315 86.68 6.485 ;
      RECT 81.81 3.57 82.13 3.83 ;
      RECT 83.1 2.745 83.24 3.605 ;
      RECT 81.9 3.465 83.24 3.605 ;
      RECT 81.9 3.025 82.04 3.83 ;
      RECT 81.825 3.025 82.115 3.255 ;
      RECT 83.025 2.745 83.315 2.975 ;
      RECT 82.545 3.025 82.835 3.255 ;
      RECT 82.74 1.95 82.88 3.21 ;
      RECT 82.77 1.89 83.09 2.15 ;
      RECT 79.37 2.45 79.69 2.71 ;
      RECT 82.065 2.465 82.355 2.695 ;
      RECT 79.46 2.37 82.28 2.51 ;
      RECT 81.33 1.89 81.65 2.15 ;
      RECT 81.825 1.905 82.115 2.135 ;
      RECT 81.33 1.95 82.115 2.09 ;
      RECT 81.33 3.01 81.65 3.27 ;
      RECT 81.33 2.79 81.56 3.27 ;
      RECT 80.825 2.745 81.115 2.975 ;
      RECT 80.825 2.79 81.56 2.93 ;
      RECT 81.09 7.765 81.38 7.995 ;
      RECT 81.15 7.025 81.32 7.995 ;
      RECT 81.05 7.055 81.43 7.425 ;
      RECT 81.09 7.025 81.38 7.425 ;
      RECT 79.85 3.57 80.17 3.83 ;
      RECT 79.385 3.585 79.675 3.815 ;
      RECT 79.385 3.63 80.17 3.77 ;
      RECT 78.145 2.465 78.435 2.695 ;
      RECT 78.145 2.51 79.08 2.65 ;
      RECT 78.94 1.95 79.08 2.65 ;
      RECT 79.61 1.89 79.93 2.15 ;
      RECT 79.385 1.905 79.93 2.135 ;
      RECT 78.94 1.95 79.93 2.09 ;
      RECT 77.29 3.57 77.61 3.83 ;
      RECT 77.29 3.63 78.36 3.77 ;
      RECT 78.22 3.07 78.36 3.77 ;
      RECT 79.385 3.025 79.675 3.255 ;
      RECT 78.22 3.07 79.675 3.21 ;
      RECT 77.65 1.89 77.97 2.15 ;
      RECT 77.425 1.905 77.97 2.135 ;
      RECT 76.67 2.45 76.99 2.71 ;
      RECT 77.665 2.465 77.955 2.695 ;
      RECT 76.425 2.465 76.99 2.695 ;
      RECT 76.425 2.51 77.955 2.65 ;
      RECT 75.945 3.025 76.235 3.255 ;
      RECT 76.14 1.95 76.28 3.21 ;
      RECT 76.93 1.89 77.25 2.15 ;
      RECT 75.945 1.905 76.235 2.135 ;
      RECT 75.945 1.95 77.25 2.09 ;
      RECT 75.54 3.465 76.64 3.605 ;
      RECT 76.425 3.305 76.715 3.535 ;
      RECT 75.465 3.305 75.755 3.535 ;
      RECT 75.45 1.89 75.77 2.15 ;
      RECT 73.49 1.89 73.81 2.15 ;
      RECT 73.49 1.95 75.77 2.09 ;
      RECT 74.61 3.01 74.93 3.27 ;
      RECT 74.61 3.01 75.44 3.15 ;
      RECT 75.225 2.745 75.44 3.15 ;
      RECT 75.225 2.745 75.515 2.975 ;
      RECT 73.01 2.45 73.33 2.71 ;
      RECT 74.42 2.465 74.71 2.695 ;
      RECT 73.01 2.465 73.555 2.695 ;
      RECT 73.01 2.55 73.96 2.69 ;
      RECT 73.82 2.37 73.96 2.69 ;
      RECT 74.32 2.465 74.71 2.65 ;
      RECT 73.82 2.37 74.46 2.51 ;
      RECT 72.53 3.26 72.85 3.675 ;
      RECT 72.61 1.905 72.765 3.675 ;
      RECT 72.545 1.905 72.835 2.135 ;
      RECT 70.925 7.77 71.215 8 ;
      RECT 70.985 6.29 71.155 8 ;
      RECT 70.935 6.655 71.285 7.005 ;
      RECT 70.925 6.29 71.215 6.52 ;
      RECT 70.52 2.395 70.625 2.965 ;
      RECT 70.52 2.73 70.845 2.96 ;
      RECT 70.52 2.76 71.015 2.93 ;
      RECT 70.52 2.395 70.71 2.96 ;
      RECT 69.935 2.36 70.225 2.59 ;
      RECT 69.935 2.395 70.71 2.565 ;
      RECT 69.995 0.88 70.165 2.59 ;
      RECT 69.935 0.88 70.225 1.11 ;
      RECT 69.935 7.77 70.225 8 ;
      RECT 69.995 6.29 70.165 8 ;
      RECT 69.935 6.29 70.225 6.52 ;
      RECT 69.935 6.325 70.79 6.485 ;
      RECT 70.62 5.92 70.79 6.485 ;
      RECT 69.935 6.32 70.33 6.485 ;
      RECT 70.555 5.92 70.845 6.15 ;
      RECT 70.555 5.95 71.015 6.12 ;
      RECT 69.565 2.73 69.855 2.96 ;
      RECT 69.565 2.76 70.025 2.93 ;
      RECT 69.63 1.655 69.795 2.96 ;
      RECT 68.145 1.625 68.435 1.855 ;
      RECT 68.145 1.655 69.795 1.825 ;
      RECT 68.205 0.885 68.375 1.855 ;
      RECT 68.145 0.885 68.435 1.115 ;
      RECT 68.145 7.765 68.435 7.995 ;
      RECT 68.205 7.025 68.375 7.995 ;
      RECT 68.205 7.12 69.795 7.29 ;
      RECT 69.625 5.92 69.795 7.29 ;
      RECT 68.145 7.025 68.435 7.255 ;
      RECT 69.565 5.92 69.855 6.15 ;
      RECT 69.565 5.95 70.025 6.12 ;
      RECT 66.195 3.15 66.535 3.5 ;
      RECT 66.285 2.025 66.455 3.5 ;
      RECT 68.575 1.965 68.925 2.315 ;
      RECT 66.285 2.025 68.925 2.195 ;
      RECT 68.6 6.655 68.925 6.98 ;
      RECT 63.16 6.61 63.51 6.96 ;
      RECT 68.575 6.655 68.925 6.885 ;
      RECT 62.96 6.655 63.51 6.885 ;
      RECT 62.79 6.685 68.925 6.855 ;
      RECT 67.8 2.365 68.12 2.685 ;
      RECT 67.77 2.365 68.12 2.595 ;
      RECT 67.6 2.395 68.12 2.565 ;
      RECT 67.8 6.255 68.12 6.545 ;
      RECT 67.77 6.285 68.12 6.515 ;
      RECT 67.6 6.315 68.12 6.485 ;
      RECT 63.25 3.57 63.57 3.83 ;
      RECT 64.54 2.745 64.68 3.605 ;
      RECT 63.34 3.465 64.68 3.605 ;
      RECT 63.34 3.025 63.48 3.83 ;
      RECT 63.265 3.025 63.555 3.255 ;
      RECT 64.465 2.745 64.755 2.975 ;
      RECT 63.985 3.025 64.275 3.255 ;
      RECT 64.18 1.95 64.32 3.21 ;
      RECT 64.21 1.89 64.53 2.15 ;
      RECT 60.81 2.45 61.13 2.71 ;
      RECT 63.505 2.465 63.795 2.695 ;
      RECT 60.9 2.37 63.72 2.51 ;
      RECT 62.77 1.89 63.09 2.15 ;
      RECT 63.265 1.905 63.555 2.135 ;
      RECT 62.77 1.95 63.555 2.09 ;
      RECT 62.77 3.01 63.09 3.27 ;
      RECT 62.77 2.79 63 3.27 ;
      RECT 62.265 2.745 62.555 2.975 ;
      RECT 62.265 2.79 63 2.93 ;
      RECT 62.53 7.765 62.82 7.995 ;
      RECT 62.59 7.025 62.76 7.995 ;
      RECT 62.49 7.055 62.87 7.425 ;
      RECT 62.53 7.025 62.82 7.425 ;
      RECT 61.29 3.57 61.61 3.83 ;
      RECT 60.825 3.585 61.115 3.815 ;
      RECT 60.825 3.63 61.61 3.77 ;
      RECT 59.585 2.465 59.875 2.695 ;
      RECT 59.585 2.51 60.52 2.65 ;
      RECT 60.38 1.95 60.52 2.65 ;
      RECT 61.05 1.89 61.37 2.15 ;
      RECT 60.825 1.905 61.37 2.135 ;
      RECT 60.38 1.95 61.37 2.09 ;
      RECT 58.73 3.57 59.05 3.83 ;
      RECT 58.73 3.63 59.8 3.77 ;
      RECT 59.66 3.07 59.8 3.77 ;
      RECT 60.825 3.025 61.115 3.255 ;
      RECT 59.66 3.07 61.115 3.21 ;
      RECT 59.09 1.89 59.41 2.15 ;
      RECT 58.865 1.905 59.41 2.135 ;
      RECT 58.11 2.45 58.43 2.71 ;
      RECT 59.105 2.465 59.395 2.695 ;
      RECT 57.865 2.465 58.43 2.695 ;
      RECT 57.865 2.51 59.395 2.65 ;
      RECT 57.385 3.025 57.675 3.255 ;
      RECT 57.58 1.95 57.72 3.21 ;
      RECT 58.37 1.89 58.69 2.15 ;
      RECT 57.385 1.905 57.675 2.135 ;
      RECT 57.385 1.95 58.69 2.09 ;
      RECT 56.98 3.465 58.08 3.605 ;
      RECT 57.865 3.305 58.155 3.535 ;
      RECT 56.905 3.305 57.195 3.535 ;
      RECT 56.89 1.89 57.21 2.15 ;
      RECT 54.93 1.89 55.25 2.15 ;
      RECT 54.93 1.95 57.21 2.09 ;
      RECT 56.05 3.01 56.37 3.27 ;
      RECT 56.05 3.01 56.88 3.15 ;
      RECT 56.665 2.745 56.88 3.15 ;
      RECT 56.665 2.745 56.955 2.975 ;
      RECT 54.45 2.45 54.77 2.71 ;
      RECT 55.86 2.465 56.15 2.695 ;
      RECT 54.45 2.465 54.995 2.695 ;
      RECT 54.45 2.55 55.4 2.69 ;
      RECT 55.26 2.37 55.4 2.69 ;
      RECT 55.76 2.465 56.15 2.65 ;
      RECT 55.26 2.37 55.9 2.51 ;
      RECT 53.97 3.26 54.29 3.675 ;
      RECT 54.05 1.905 54.205 3.675 ;
      RECT 53.985 1.905 54.275 2.135 ;
      RECT 52.365 7.77 52.655 8 ;
      RECT 52.425 6.29 52.595 8 ;
      RECT 52.375 6.655 52.725 7.005 ;
      RECT 52.365 6.29 52.655 6.52 ;
      RECT 51.96 2.395 52.065 2.965 ;
      RECT 51.96 2.73 52.285 2.96 ;
      RECT 51.96 2.76 52.455 2.93 ;
      RECT 51.96 2.395 52.15 2.96 ;
      RECT 51.375 2.36 51.665 2.59 ;
      RECT 51.375 2.395 52.15 2.565 ;
      RECT 51.435 0.88 51.605 2.59 ;
      RECT 51.375 0.88 51.665 1.11 ;
      RECT 51.375 7.77 51.665 8 ;
      RECT 51.435 6.29 51.605 8 ;
      RECT 51.375 6.29 51.665 6.52 ;
      RECT 51.375 6.325 52.23 6.485 ;
      RECT 52.06 5.92 52.23 6.485 ;
      RECT 51.375 6.32 51.77 6.485 ;
      RECT 51.995 5.92 52.285 6.15 ;
      RECT 51.995 5.95 52.455 6.12 ;
      RECT 51.005 2.73 51.295 2.96 ;
      RECT 51.005 2.76 51.465 2.93 ;
      RECT 51.07 1.655 51.235 2.96 ;
      RECT 49.585 1.625 49.875 1.855 ;
      RECT 49.585 1.655 51.235 1.825 ;
      RECT 49.645 0.885 49.815 1.855 ;
      RECT 49.585 0.885 49.875 1.115 ;
      RECT 49.585 7.765 49.875 7.995 ;
      RECT 49.645 7.025 49.815 7.995 ;
      RECT 49.645 7.12 51.235 7.29 ;
      RECT 51.065 5.92 51.235 7.29 ;
      RECT 49.585 7.025 49.875 7.255 ;
      RECT 51.005 5.92 51.295 6.15 ;
      RECT 51.005 5.95 51.465 6.12 ;
      RECT 47.635 3.15 47.975 3.5 ;
      RECT 47.725 2.025 47.895 3.5 ;
      RECT 50.015 1.965 50.365 2.315 ;
      RECT 47.725 2.025 50.365 2.195 ;
      RECT 50.04 6.655 50.365 6.98 ;
      RECT 44.6 6.615 44.95 6.965 ;
      RECT 50.015 6.655 50.365 6.885 ;
      RECT 44.4 6.655 44.95 6.885 ;
      RECT 44.23 6.685 50.365 6.855 ;
      RECT 49.24 2.365 49.56 2.685 ;
      RECT 49.21 2.365 49.56 2.595 ;
      RECT 49.04 2.395 49.56 2.565 ;
      RECT 49.24 6.255 49.56 6.545 ;
      RECT 49.21 6.285 49.56 6.515 ;
      RECT 49.04 6.315 49.56 6.485 ;
      RECT 44.69 3.57 45.01 3.83 ;
      RECT 45.98 2.745 46.12 3.605 ;
      RECT 44.78 3.465 46.12 3.605 ;
      RECT 44.78 3.025 44.92 3.83 ;
      RECT 44.705 3.025 44.995 3.255 ;
      RECT 45.905 2.745 46.195 2.975 ;
      RECT 45.425 3.025 45.715 3.255 ;
      RECT 45.62 1.95 45.76 3.21 ;
      RECT 45.65 1.89 45.97 2.15 ;
      RECT 42.25 2.45 42.57 2.71 ;
      RECT 44.945 2.465 45.235 2.695 ;
      RECT 42.34 2.37 45.16 2.51 ;
      RECT 44.21 1.89 44.53 2.15 ;
      RECT 44.705 1.905 44.995 2.135 ;
      RECT 44.21 1.95 44.995 2.09 ;
      RECT 44.21 3.01 44.53 3.27 ;
      RECT 44.21 2.79 44.44 3.27 ;
      RECT 43.705 2.745 43.995 2.975 ;
      RECT 43.705 2.79 44.44 2.93 ;
      RECT 43.97 7.765 44.26 7.995 ;
      RECT 44.03 7.025 44.2 7.995 ;
      RECT 43.93 7.055 44.31 7.425 ;
      RECT 43.97 7.025 44.26 7.425 ;
      RECT 42.73 3.57 43.05 3.83 ;
      RECT 42.265 3.585 42.555 3.815 ;
      RECT 42.265 3.63 43.05 3.77 ;
      RECT 41.025 2.465 41.315 2.695 ;
      RECT 41.025 2.51 41.96 2.65 ;
      RECT 41.82 1.95 41.96 2.65 ;
      RECT 42.49 1.89 42.81 2.15 ;
      RECT 42.265 1.905 42.81 2.135 ;
      RECT 41.82 1.95 42.81 2.09 ;
      RECT 40.17 3.57 40.49 3.83 ;
      RECT 40.17 3.63 41.24 3.77 ;
      RECT 41.1 3.07 41.24 3.77 ;
      RECT 42.265 3.025 42.555 3.255 ;
      RECT 41.1 3.07 42.555 3.21 ;
      RECT 40.53 1.89 40.85 2.15 ;
      RECT 40.305 1.905 40.85 2.135 ;
      RECT 39.55 2.45 39.87 2.71 ;
      RECT 40.545 2.465 40.835 2.695 ;
      RECT 39.305 2.465 39.87 2.695 ;
      RECT 39.305 2.51 40.835 2.65 ;
      RECT 38.825 3.025 39.115 3.255 ;
      RECT 39.02 1.95 39.16 3.21 ;
      RECT 39.81 1.89 40.13 2.15 ;
      RECT 38.825 1.905 39.115 2.135 ;
      RECT 38.825 1.95 40.13 2.09 ;
      RECT 38.42 3.465 39.52 3.605 ;
      RECT 39.305 3.305 39.595 3.535 ;
      RECT 38.345 3.305 38.635 3.535 ;
      RECT 38.33 1.89 38.65 2.15 ;
      RECT 36.37 1.89 36.69 2.15 ;
      RECT 36.37 1.95 38.65 2.09 ;
      RECT 37.49 3.01 37.81 3.27 ;
      RECT 37.49 3.01 38.32 3.15 ;
      RECT 38.105 2.745 38.32 3.15 ;
      RECT 38.105 2.745 38.395 2.975 ;
      RECT 35.89 2.45 36.21 2.71 ;
      RECT 37.3 2.465 37.59 2.695 ;
      RECT 35.89 2.465 36.435 2.695 ;
      RECT 35.89 2.55 36.84 2.69 ;
      RECT 36.7 2.37 36.84 2.69 ;
      RECT 37.2 2.465 37.59 2.65 ;
      RECT 36.7 2.37 37.34 2.51 ;
      RECT 35.41 3.26 35.73 3.675 ;
      RECT 35.49 1.905 35.645 3.675 ;
      RECT 35.425 1.905 35.715 2.135 ;
      RECT 33.805 7.77 34.095 8 ;
      RECT 33.865 6.29 34.035 8 ;
      RECT 33.855 6.66 34.21 7.015 ;
      RECT 33.805 6.29 34.095 6.52 ;
      RECT 33.4 2.395 33.505 2.965 ;
      RECT 33.4 2.73 33.725 2.96 ;
      RECT 33.4 2.76 33.895 2.93 ;
      RECT 33.4 2.395 33.59 2.96 ;
      RECT 32.815 2.36 33.105 2.59 ;
      RECT 32.815 2.395 33.59 2.565 ;
      RECT 32.875 0.88 33.045 2.59 ;
      RECT 32.815 0.88 33.105 1.11 ;
      RECT 32.815 7.77 33.105 8 ;
      RECT 32.875 6.29 33.045 8 ;
      RECT 32.815 6.29 33.105 6.52 ;
      RECT 32.815 6.325 33.67 6.485 ;
      RECT 33.5 5.92 33.67 6.485 ;
      RECT 32.815 6.32 33.21 6.485 ;
      RECT 33.435 5.92 33.725 6.15 ;
      RECT 33.435 5.95 33.895 6.12 ;
      RECT 32.445 2.73 32.735 2.96 ;
      RECT 32.445 2.76 32.905 2.93 ;
      RECT 32.51 1.655 32.675 2.96 ;
      RECT 31.025 1.625 31.315 1.855 ;
      RECT 31.025 1.655 32.675 1.825 ;
      RECT 31.085 0.885 31.255 1.855 ;
      RECT 31.025 0.885 31.315 1.115 ;
      RECT 31.025 7.765 31.315 7.995 ;
      RECT 31.085 7.025 31.255 7.995 ;
      RECT 31.085 7.12 32.675 7.29 ;
      RECT 32.505 5.92 32.675 7.29 ;
      RECT 31.025 7.025 31.315 7.255 ;
      RECT 32.445 5.92 32.735 6.15 ;
      RECT 32.445 5.95 32.905 6.12 ;
      RECT 29.075 3.15 29.415 3.5 ;
      RECT 29.165 2.025 29.335 3.5 ;
      RECT 31.455 1.965 31.805 2.315 ;
      RECT 29.165 2.025 31.805 2.195 ;
      RECT 31.48 6.655 31.805 6.98 ;
      RECT 26.045 6.61 26.395 6.96 ;
      RECT 31.455 6.655 31.805 6.885 ;
      RECT 25.84 6.655 26.395 6.885 ;
      RECT 25.67 6.685 31.805 6.855 ;
      RECT 30.68 2.365 31 2.685 ;
      RECT 30.65 2.365 31 2.595 ;
      RECT 30.48 2.395 31 2.565 ;
      RECT 30.68 6.255 31 6.545 ;
      RECT 30.65 6.285 31 6.515 ;
      RECT 30.48 6.315 31 6.485 ;
      RECT 26.13 3.57 26.45 3.83 ;
      RECT 27.42 2.745 27.56 3.605 ;
      RECT 26.22 3.465 27.56 3.605 ;
      RECT 26.22 3.025 26.36 3.83 ;
      RECT 26.145 3.025 26.435 3.255 ;
      RECT 27.345 2.745 27.635 2.975 ;
      RECT 26.865 3.025 27.155 3.255 ;
      RECT 27.06 1.95 27.2 3.21 ;
      RECT 27.09 1.89 27.41 2.15 ;
      RECT 23.69 2.45 24.01 2.71 ;
      RECT 26.385 2.465 26.675 2.695 ;
      RECT 23.78 2.37 26.6 2.51 ;
      RECT 25.65 1.89 25.97 2.15 ;
      RECT 26.145 1.905 26.435 2.135 ;
      RECT 25.65 1.95 26.435 2.09 ;
      RECT 25.65 3.01 25.97 3.27 ;
      RECT 25.65 2.79 25.88 3.27 ;
      RECT 25.145 2.745 25.435 2.975 ;
      RECT 25.145 2.79 25.88 2.93 ;
      RECT 25.41 7.765 25.7 7.995 ;
      RECT 25.47 7.025 25.64 7.995 ;
      RECT 25.37 7.055 25.75 7.425 ;
      RECT 25.41 7.025 25.7 7.425 ;
      RECT 24.17 3.57 24.49 3.83 ;
      RECT 23.705 3.585 23.995 3.815 ;
      RECT 23.705 3.63 24.49 3.77 ;
      RECT 22.465 2.465 22.755 2.695 ;
      RECT 22.465 2.51 23.4 2.65 ;
      RECT 23.26 1.95 23.4 2.65 ;
      RECT 23.93 1.89 24.25 2.15 ;
      RECT 23.705 1.905 24.25 2.135 ;
      RECT 23.26 1.95 24.25 2.09 ;
      RECT 21.61 3.57 21.93 3.83 ;
      RECT 21.61 3.63 22.68 3.77 ;
      RECT 22.54 3.07 22.68 3.77 ;
      RECT 23.705 3.025 23.995 3.255 ;
      RECT 22.54 3.07 23.995 3.21 ;
      RECT 21.97 1.89 22.29 2.15 ;
      RECT 21.745 1.905 22.29 2.135 ;
      RECT 20.99 2.45 21.31 2.71 ;
      RECT 21.985 2.465 22.275 2.695 ;
      RECT 20.745 2.465 21.31 2.695 ;
      RECT 20.745 2.51 22.275 2.65 ;
      RECT 20.265 3.025 20.555 3.255 ;
      RECT 20.46 1.95 20.6 3.21 ;
      RECT 21.25 1.89 21.57 2.15 ;
      RECT 20.265 1.905 20.555 2.135 ;
      RECT 20.265 1.95 21.57 2.09 ;
      RECT 19.86 3.465 20.96 3.605 ;
      RECT 20.745 3.305 21.035 3.535 ;
      RECT 19.785 3.305 20.075 3.535 ;
      RECT 19.77 1.89 20.09 2.15 ;
      RECT 17.81 1.89 18.13 2.15 ;
      RECT 17.81 1.95 20.09 2.09 ;
      RECT 18.93 3.01 19.25 3.27 ;
      RECT 18.93 3.01 19.76 3.15 ;
      RECT 19.545 2.745 19.76 3.15 ;
      RECT 19.545 2.745 19.835 2.975 ;
      RECT 17.33 2.45 17.65 2.71 ;
      RECT 18.74 2.465 19.03 2.695 ;
      RECT 17.33 2.465 17.875 2.695 ;
      RECT 17.33 2.55 18.28 2.69 ;
      RECT 18.14 2.37 18.28 2.69 ;
      RECT 18.64 2.465 19.03 2.65 ;
      RECT 18.14 2.37 18.78 2.51 ;
      RECT 16.85 3.26 17.17 3.675 ;
      RECT 16.93 1.905 17.085 3.675 ;
      RECT 16.865 1.905 17.155 2.135 ;
      RECT 15.245 7.77 15.535 8 ;
      RECT 15.305 6.29 15.475 8 ;
      RECT 15.3 6.655 15.65 7.005 ;
      RECT 15.245 6.29 15.535 6.52 ;
      RECT 14.84 2.395 14.945 2.965 ;
      RECT 14.84 2.73 15.165 2.96 ;
      RECT 14.84 2.76 15.335 2.93 ;
      RECT 14.84 2.395 15.03 2.96 ;
      RECT 14.255 2.36 14.545 2.59 ;
      RECT 14.255 2.395 15.03 2.565 ;
      RECT 14.315 0.88 14.485 2.59 ;
      RECT 14.255 0.88 14.545 1.11 ;
      RECT 14.255 7.77 14.545 8 ;
      RECT 14.315 6.29 14.485 8 ;
      RECT 14.255 6.29 14.545 6.52 ;
      RECT 14.255 6.325 15.11 6.485 ;
      RECT 14.94 5.92 15.11 6.485 ;
      RECT 14.255 6.32 14.65 6.485 ;
      RECT 14.875 5.92 15.165 6.15 ;
      RECT 14.875 5.95 15.335 6.12 ;
      RECT 13.885 2.73 14.175 2.96 ;
      RECT 13.885 2.76 14.345 2.93 ;
      RECT 13.95 1.655 14.115 2.96 ;
      RECT 12.465 1.625 12.755 1.855 ;
      RECT 12.465 1.655 14.115 1.825 ;
      RECT 12.525 0.885 12.695 1.855 ;
      RECT 12.465 0.885 12.755 1.115 ;
      RECT 12.465 7.765 12.755 7.995 ;
      RECT 12.525 7.025 12.695 7.995 ;
      RECT 12.525 7.12 14.115 7.29 ;
      RECT 13.945 5.92 14.115 7.29 ;
      RECT 12.465 7.025 12.755 7.255 ;
      RECT 13.885 5.92 14.175 6.15 ;
      RECT 13.885 5.95 14.345 6.12 ;
      RECT 10.515 3.15 10.855 3.5 ;
      RECT 10.605 2.025 10.775 3.5 ;
      RECT 12.895 1.965 13.245 2.315 ;
      RECT 10.605 2.025 13.245 2.195 ;
      RECT 12.92 6.655 13.245 6.98 ;
      RECT 7.485 6.605 7.835 6.955 ;
      RECT 12.895 6.655 13.245 6.885 ;
      RECT 7.28 6.655 7.835 6.885 ;
      RECT 7.11 6.685 13.245 6.855 ;
      RECT 12.12 2.365 12.44 2.685 ;
      RECT 12.09 2.365 12.44 2.595 ;
      RECT 11.92 2.395 12.44 2.565 ;
      RECT 12.12 6.255 12.44 6.545 ;
      RECT 12.09 6.285 12.44 6.515 ;
      RECT 11.92 6.315 12.44 6.485 ;
      RECT 7.57 3.57 7.89 3.83 ;
      RECT 8.86 2.745 9 3.605 ;
      RECT 7.66 3.465 9 3.605 ;
      RECT 7.66 3.025 7.8 3.83 ;
      RECT 7.585 3.025 7.875 3.255 ;
      RECT 8.785 2.745 9.075 2.975 ;
      RECT 8.305 3.025 8.595 3.255 ;
      RECT 8.5 1.95 8.64 3.21 ;
      RECT 8.53 1.89 8.85 2.15 ;
      RECT 5.13 2.45 5.45 2.71 ;
      RECT 7.825 2.465 8.115 2.695 ;
      RECT 5.22 2.37 8.04 2.51 ;
      RECT 7.09 1.89 7.41 2.15 ;
      RECT 7.585 1.905 7.875 2.135 ;
      RECT 7.09 1.95 7.875 2.09 ;
      RECT 7.09 3.01 7.41 3.27 ;
      RECT 7.09 2.79 7.32 3.27 ;
      RECT 6.585 2.745 6.875 2.975 ;
      RECT 6.585 2.79 7.32 2.93 ;
      RECT 6.85 7.765 7.14 7.995 ;
      RECT 6.91 7.025 7.08 7.995 ;
      RECT 6.81 7.055 7.19 7.425 ;
      RECT 6.85 7.025 7.14 7.425 ;
      RECT 5.61 3.57 5.93 3.83 ;
      RECT 5.145 3.585 5.435 3.815 ;
      RECT 5.145 3.63 5.93 3.77 ;
      RECT 3.905 2.465 4.195 2.695 ;
      RECT 3.905 2.51 4.84 2.65 ;
      RECT 4.7 1.95 4.84 2.65 ;
      RECT 5.37 1.89 5.69 2.15 ;
      RECT 5.145 1.905 5.69 2.135 ;
      RECT 4.7 1.95 5.69 2.09 ;
      RECT 3.05 3.57 3.37 3.83 ;
      RECT 3.05 3.63 4.12 3.77 ;
      RECT 3.98 3.07 4.12 3.77 ;
      RECT 5.145 3.025 5.435 3.255 ;
      RECT 3.98 3.07 5.435 3.21 ;
      RECT 3.41 1.89 3.73 2.15 ;
      RECT 3.185 1.905 3.73 2.135 ;
      RECT 2.43 2.45 2.75 2.71 ;
      RECT 3.425 2.465 3.715 2.695 ;
      RECT 2.185 2.465 2.75 2.695 ;
      RECT 2.185 2.51 3.715 2.65 ;
      RECT 1.705 3.025 1.995 3.255 ;
      RECT 1.9 1.95 2.04 3.21 ;
      RECT 2.69 1.89 3.01 2.15 ;
      RECT 1.705 1.905 1.995 2.135 ;
      RECT 1.705 1.95 3.01 2.09 ;
      RECT 1.3 3.465 2.4 3.605 ;
      RECT 2.185 3.305 2.475 3.535 ;
      RECT 1.225 3.305 1.515 3.535 ;
      RECT 1.21 1.89 1.53 2.15 ;
      RECT -0.75 1.89 -0.43 2.15 ;
      RECT -0.75 1.95 1.53 2.09 ;
      RECT 0.37 3.01 0.69 3.27 ;
      RECT 0.37 3.01 1.2 3.15 ;
      RECT 0.985 2.745 1.2 3.15 ;
      RECT 0.985 2.745 1.275 2.975 ;
      RECT -1.23 2.45 -0.91 2.71 ;
      RECT 0.18 2.465 0.47 2.695 ;
      RECT -1.23 2.465 -0.685 2.695 ;
      RECT -1.23 2.55 -0.28 2.69 ;
      RECT -0.42 2.37 -0.28 2.69 ;
      RECT 0.08 2.465 0.47 2.65 ;
      RECT -0.42 2.37 0.22 2.51 ;
      RECT -1.71 3.26 -1.39 3.675 ;
      RECT -1.63 1.905 -1.475 3.675 ;
      RECT -1.695 1.905 -1.405 2.135 ;
      RECT -3.965 7.765 -3.675 7.995 ;
      RECT -3.905 7.025 -3.735 7.995 ;
      RECT -3.995 7.025 -3.645 7.315 ;
      RECT -4.37 6.285 -4.02 6.575 ;
      RECT -4.51 6.315 -4.02 6.485 ;
      RECT 80.81 3.57 81.13 3.83 ;
      RECT 80.21 1.89 80.89 2.15 ;
      RECT 80.33 3.57 80.65 3.83 ;
      RECT 78.85 3.57 79.17 3.83 ;
      RECT 78.37 1.89 78.69 2.15 ;
      RECT 77.65 3.01 77.97 3.27 ;
      RECT 76.93 3.01 77.25 3.27 ;
      RECT 73.49 3.01 73.81 3.27 ;
      RECT 62.25 3.57 62.57 3.83 ;
      RECT 61.65 1.89 62.33 2.15 ;
      RECT 61.77 3.57 62.09 3.83 ;
      RECT 60.29 3.57 60.61 3.83 ;
      RECT 59.81 1.89 60.13 2.15 ;
      RECT 59.09 3.01 59.41 3.27 ;
      RECT 58.37 3.01 58.69 3.27 ;
      RECT 54.93 3.01 55.25 3.27 ;
      RECT 43.69 3.57 44.01 3.83 ;
      RECT 43.09 1.89 43.77 2.15 ;
      RECT 43.21 3.57 43.53 3.83 ;
      RECT 41.73 3.57 42.05 3.83 ;
      RECT 41.25 1.89 41.57 2.15 ;
      RECT 40.53 3.01 40.85 3.27 ;
      RECT 39.81 3.01 40.13 3.27 ;
      RECT 36.37 3.01 36.69 3.27 ;
      RECT 25.13 3.57 25.45 3.83 ;
      RECT 24.53 1.89 25.21 2.15 ;
      RECT 24.65 3.57 24.97 3.83 ;
      RECT 23.17 3.57 23.49 3.83 ;
      RECT 22.69 1.89 23.01 2.15 ;
      RECT 21.97 3.01 22.29 3.27 ;
      RECT 21.25 3.01 21.57 3.27 ;
      RECT 17.81 3.01 18.13 3.27 ;
      RECT 6.57 3.57 6.89 3.83 ;
      RECT 5.97 1.89 6.65 2.15 ;
      RECT 6.09 3.57 6.41 3.83 ;
      RECT 4.61 3.57 4.93 3.83 ;
      RECT 4.13 1.89 4.45 2.15 ;
      RECT 3.41 3.01 3.73 3.27 ;
      RECT 2.69 3.01 3.01 3.27 ;
      RECT -0.75 3.01 -0.43 3.27 ;
    LAYER mcon ;
      RECT 89.545 6.32 89.715 6.49 ;
      RECT 89.55 6.315 89.72 6.485 ;
      RECT 70.985 6.32 71.155 6.49 ;
      RECT 70.99 6.315 71.16 6.485 ;
      RECT 52.425 6.32 52.595 6.49 ;
      RECT 52.43 6.315 52.6 6.485 ;
      RECT 33.865 6.32 34.035 6.49 ;
      RECT 33.87 6.315 34.04 6.485 ;
      RECT 15.305 6.32 15.475 6.49 ;
      RECT 15.31 6.315 15.48 6.485 ;
      RECT 89.545 7.8 89.715 7.97 ;
      RECT 89.175 2.76 89.345 2.93 ;
      RECT 89.175 5.95 89.345 6.12 ;
      RECT 88.555 0.91 88.725 1.08 ;
      RECT 88.555 2.39 88.725 2.56 ;
      RECT 88.555 6.32 88.725 6.49 ;
      RECT 88.555 7.8 88.725 7.97 ;
      RECT 88.185 2.76 88.355 2.93 ;
      RECT 88.185 5.95 88.355 6.12 ;
      RECT 87.195 2.025 87.365 2.195 ;
      RECT 87.195 6.685 87.365 6.855 ;
      RECT 86.765 0.915 86.935 1.085 ;
      RECT 86.765 1.655 86.935 1.825 ;
      RECT 86.765 7.055 86.935 7.225 ;
      RECT 86.765 7.795 86.935 7.965 ;
      RECT 86.39 2.395 86.56 2.565 ;
      RECT 86.39 6.315 86.56 6.485 ;
      RECT 83.085 2.775 83.255 2.945 ;
      RECT 82.845 1.935 83.015 2.105 ;
      RECT 82.605 3.055 82.775 3.225 ;
      RECT 82.125 2.495 82.295 2.665 ;
      RECT 81.885 1.935 82.055 2.105 ;
      RECT 81.885 3.055 82.055 3.225 ;
      RECT 81.885 3.615 82.055 3.785 ;
      RECT 81.58 6.685 81.75 6.855 ;
      RECT 81.405 3.055 81.575 3.225 ;
      RECT 81.15 7.055 81.32 7.225 ;
      RECT 81.15 7.795 81.32 7.965 ;
      RECT 80.885 2.775 81.055 2.945 ;
      RECT 80.885 3.615 81.055 3.785 ;
      RECT 80.405 1.935 80.575 2.105 ;
      RECT 80.405 3.615 80.575 3.785 ;
      RECT 79.445 1.935 79.615 2.105 ;
      RECT 79.445 2.495 79.615 2.665 ;
      RECT 79.445 3.055 79.615 3.225 ;
      RECT 79.445 3.615 79.615 3.785 ;
      RECT 78.925 3.615 79.095 3.785 ;
      RECT 78.445 1.935 78.615 2.105 ;
      RECT 78.205 2.495 78.375 2.665 ;
      RECT 77.725 2.495 77.895 2.665 ;
      RECT 77.725 3.055 77.895 3.225 ;
      RECT 77.485 1.935 77.655 2.105 ;
      RECT 77.005 3.055 77.175 3.225 ;
      RECT 76.485 2.495 76.655 2.665 ;
      RECT 76.485 3.335 76.655 3.505 ;
      RECT 76.005 1.935 76.175 2.105 ;
      RECT 76.005 3.055 76.175 3.225 ;
      RECT 75.525 3.335 75.695 3.505 ;
      RECT 75.285 2.775 75.455 2.945 ;
      RECT 74.48 2.495 74.65 2.665 ;
      RECT 73.565 1.935 73.735 2.105 ;
      RECT 73.565 3.055 73.735 3.225 ;
      RECT 73.325 2.495 73.495 2.665 ;
      RECT 72.605 1.935 72.775 2.105 ;
      RECT 72.605 3.475 72.775 3.645 ;
      RECT 70.985 7.8 71.155 7.97 ;
      RECT 70.615 2.76 70.785 2.93 ;
      RECT 70.615 5.95 70.785 6.12 ;
      RECT 69.995 0.91 70.165 1.08 ;
      RECT 69.995 2.39 70.165 2.56 ;
      RECT 69.995 6.32 70.165 6.49 ;
      RECT 69.995 7.8 70.165 7.97 ;
      RECT 69.625 2.76 69.795 2.93 ;
      RECT 69.625 5.95 69.795 6.12 ;
      RECT 68.635 2.025 68.805 2.195 ;
      RECT 68.635 6.685 68.805 6.855 ;
      RECT 68.205 0.915 68.375 1.085 ;
      RECT 68.205 1.655 68.375 1.825 ;
      RECT 68.205 7.055 68.375 7.225 ;
      RECT 68.205 7.795 68.375 7.965 ;
      RECT 67.83 2.395 68 2.565 ;
      RECT 67.83 6.315 68 6.485 ;
      RECT 64.525 2.775 64.695 2.945 ;
      RECT 64.285 1.935 64.455 2.105 ;
      RECT 64.045 3.055 64.215 3.225 ;
      RECT 63.565 2.495 63.735 2.665 ;
      RECT 63.325 1.935 63.495 2.105 ;
      RECT 63.325 3.055 63.495 3.225 ;
      RECT 63.325 3.615 63.495 3.785 ;
      RECT 63.02 6.685 63.19 6.855 ;
      RECT 62.845 3.055 63.015 3.225 ;
      RECT 62.59 7.055 62.76 7.225 ;
      RECT 62.59 7.795 62.76 7.965 ;
      RECT 62.325 2.775 62.495 2.945 ;
      RECT 62.325 3.615 62.495 3.785 ;
      RECT 61.845 1.935 62.015 2.105 ;
      RECT 61.845 3.615 62.015 3.785 ;
      RECT 60.885 1.935 61.055 2.105 ;
      RECT 60.885 2.495 61.055 2.665 ;
      RECT 60.885 3.055 61.055 3.225 ;
      RECT 60.885 3.615 61.055 3.785 ;
      RECT 60.365 3.615 60.535 3.785 ;
      RECT 59.885 1.935 60.055 2.105 ;
      RECT 59.645 2.495 59.815 2.665 ;
      RECT 59.165 2.495 59.335 2.665 ;
      RECT 59.165 3.055 59.335 3.225 ;
      RECT 58.925 1.935 59.095 2.105 ;
      RECT 58.445 3.055 58.615 3.225 ;
      RECT 57.925 2.495 58.095 2.665 ;
      RECT 57.925 3.335 58.095 3.505 ;
      RECT 57.445 1.935 57.615 2.105 ;
      RECT 57.445 3.055 57.615 3.225 ;
      RECT 56.965 3.335 57.135 3.505 ;
      RECT 56.725 2.775 56.895 2.945 ;
      RECT 55.92 2.495 56.09 2.665 ;
      RECT 55.005 1.935 55.175 2.105 ;
      RECT 55.005 3.055 55.175 3.225 ;
      RECT 54.765 2.495 54.935 2.665 ;
      RECT 54.045 1.935 54.215 2.105 ;
      RECT 54.045 3.475 54.215 3.645 ;
      RECT 52.425 7.8 52.595 7.97 ;
      RECT 52.055 2.76 52.225 2.93 ;
      RECT 52.055 5.95 52.225 6.12 ;
      RECT 51.435 0.91 51.605 1.08 ;
      RECT 51.435 2.39 51.605 2.56 ;
      RECT 51.435 6.32 51.605 6.49 ;
      RECT 51.435 7.8 51.605 7.97 ;
      RECT 51.065 2.76 51.235 2.93 ;
      RECT 51.065 5.95 51.235 6.12 ;
      RECT 50.075 2.025 50.245 2.195 ;
      RECT 50.075 6.685 50.245 6.855 ;
      RECT 49.645 0.915 49.815 1.085 ;
      RECT 49.645 1.655 49.815 1.825 ;
      RECT 49.645 7.055 49.815 7.225 ;
      RECT 49.645 7.795 49.815 7.965 ;
      RECT 49.27 2.395 49.44 2.565 ;
      RECT 49.27 6.315 49.44 6.485 ;
      RECT 45.965 2.775 46.135 2.945 ;
      RECT 45.725 1.935 45.895 2.105 ;
      RECT 45.485 3.055 45.655 3.225 ;
      RECT 45.005 2.495 45.175 2.665 ;
      RECT 44.765 1.935 44.935 2.105 ;
      RECT 44.765 3.055 44.935 3.225 ;
      RECT 44.765 3.615 44.935 3.785 ;
      RECT 44.46 6.685 44.63 6.855 ;
      RECT 44.285 3.055 44.455 3.225 ;
      RECT 44.03 7.055 44.2 7.225 ;
      RECT 44.03 7.795 44.2 7.965 ;
      RECT 43.765 2.775 43.935 2.945 ;
      RECT 43.765 3.615 43.935 3.785 ;
      RECT 43.285 1.935 43.455 2.105 ;
      RECT 43.285 3.615 43.455 3.785 ;
      RECT 42.325 1.935 42.495 2.105 ;
      RECT 42.325 2.495 42.495 2.665 ;
      RECT 42.325 3.055 42.495 3.225 ;
      RECT 42.325 3.615 42.495 3.785 ;
      RECT 41.805 3.615 41.975 3.785 ;
      RECT 41.325 1.935 41.495 2.105 ;
      RECT 41.085 2.495 41.255 2.665 ;
      RECT 40.605 2.495 40.775 2.665 ;
      RECT 40.605 3.055 40.775 3.225 ;
      RECT 40.365 1.935 40.535 2.105 ;
      RECT 39.885 3.055 40.055 3.225 ;
      RECT 39.365 2.495 39.535 2.665 ;
      RECT 39.365 3.335 39.535 3.505 ;
      RECT 38.885 1.935 39.055 2.105 ;
      RECT 38.885 3.055 39.055 3.225 ;
      RECT 38.405 3.335 38.575 3.505 ;
      RECT 38.165 2.775 38.335 2.945 ;
      RECT 37.36 2.495 37.53 2.665 ;
      RECT 36.445 1.935 36.615 2.105 ;
      RECT 36.445 3.055 36.615 3.225 ;
      RECT 36.205 2.495 36.375 2.665 ;
      RECT 35.485 1.935 35.655 2.105 ;
      RECT 35.485 3.475 35.655 3.645 ;
      RECT 33.865 7.8 34.035 7.97 ;
      RECT 33.495 2.76 33.665 2.93 ;
      RECT 33.495 5.95 33.665 6.12 ;
      RECT 32.875 0.91 33.045 1.08 ;
      RECT 32.875 2.39 33.045 2.56 ;
      RECT 32.875 6.32 33.045 6.49 ;
      RECT 32.875 7.8 33.045 7.97 ;
      RECT 32.505 2.76 32.675 2.93 ;
      RECT 32.505 5.95 32.675 6.12 ;
      RECT 31.515 2.025 31.685 2.195 ;
      RECT 31.515 6.685 31.685 6.855 ;
      RECT 31.085 0.915 31.255 1.085 ;
      RECT 31.085 1.655 31.255 1.825 ;
      RECT 31.085 7.055 31.255 7.225 ;
      RECT 31.085 7.795 31.255 7.965 ;
      RECT 30.71 2.395 30.88 2.565 ;
      RECT 30.71 6.315 30.88 6.485 ;
      RECT 27.405 2.775 27.575 2.945 ;
      RECT 27.165 1.935 27.335 2.105 ;
      RECT 26.925 3.055 27.095 3.225 ;
      RECT 26.445 2.495 26.615 2.665 ;
      RECT 26.205 1.935 26.375 2.105 ;
      RECT 26.205 3.055 26.375 3.225 ;
      RECT 26.205 3.615 26.375 3.785 ;
      RECT 25.9 6.685 26.07 6.855 ;
      RECT 25.725 3.055 25.895 3.225 ;
      RECT 25.47 7.055 25.64 7.225 ;
      RECT 25.47 7.795 25.64 7.965 ;
      RECT 25.205 2.775 25.375 2.945 ;
      RECT 25.205 3.615 25.375 3.785 ;
      RECT 24.725 1.935 24.895 2.105 ;
      RECT 24.725 3.615 24.895 3.785 ;
      RECT 23.765 1.935 23.935 2.105 ;
      RECT 23.765 2.495 23.935 2.665 ;
      RECT 23.765 3.055 23.935 3.225 ;
      RECT 23.765 3.615 23.935 3.785 ;
      RECT 23.245 3.615 23.415 3.785 ;
      RECT 22.765 1.935 22.935 2.105 ;
      RECT 22.525 2.495 22.695 2.665 ;
      RECT 22.045 2.495 22.215 2.665 ;
      RECT 22.045 3.055 22.215 3.225 ;
      RECT 21.805 1.935 21.975 2.105 ;
      RECT 21.325 3.055 21.495 3.225 ;
      RECT 20.805 2.495 20.975 2.665 ;
      RECT 20.805 3.335 20.975 3.505 ;
      RECT 20.325 1.935 20.495 2.105 ;
      RECT 20.325 3.055 20.495 3.225 ;
      RECT 19.845 3.335 20.015 3.505 ;
      RECT 19.605 2.775 19.775 2.945 ;
      RECT 18.8 2.495 18.97 2.665 ;
      RECT 17.885 1.935 18.055 2.105 ;
      RECT 17.885 3.055 18.055 3.225 ;
      RECT 17.645 2.495 17.815 2.665 ;
      RECT 16.925 1.935 17.095 2.105 ;
      RECT 16.925 3.475 17.095 3.645 ;
      RECT 15.305 7.8 15.475 7.97 ;
      RECT 14.935 2.76 15.105 2.93 ;
      RECT 14.935 5.95 15.105 6.12 ;
      RECT 14.315 0.91 14.485 1.08 ;
      RECT 14.315 2.39 14.485 2.56 ;
      RECT 14.315 6.32 14.485 6.49 ;
      RECT 14.315 7.8 14.485 7.97 ;
      RECT 13.945 2.76 14.115 2.93 ;
      RECT 13.945 5.95 14.115 6.12 ;
      RECT 12.955 2.025 13.125 2.195 ;
      RECT 12.955 6.685 13.125 6.855 ;
      RECT 12.525 0.915 12.695 1.085 ;
      RECT 12.525 1.655 12.695 1.825 ;
      RECT 12.525 7.055 12.695 7.225 ;
      RECT 12.525 7.795 12.695 7.965 ;
      RECT 12.15 2.395 12.32 2.565 ;
      RECT 12.15 6.315 12.32 6.485 ;
      RECT 8.845 2.775 9.015 2.945 ;
      RECT 8.605 1.935 8.775 2.105 ;
      RECT 8.365 3.055 8.535 3.225 ;
      RECT 7.885 2.495 8.055 2.665 ;
      RECT 7.645 1.935 7.815 2.105 ;
      RECT 7.645 3.055 7.815 3.225 ;
      RECT 7.645 3.615 7.815 3.785 ;
      RECT 7.34 6.685 7.51 6.855 ;
      RECT 7.165 3.055 7.335 3.225 ;
      RECT 6.91 7.055 7.08 7.225 ;
      RECT 6.91 7.795 7.08 7.965 ;
      RECT 6.645 2.775 6.815 2.945 ;
      RECT 6.645 3.615 6.815 3.785 ;
      RECT 6.165 1.935 6.335 2.105 ;
      RECT 6.165 3.615 6.335 3.785 ;
      RECT 5.205 1.935 5.375 2.105 ;
      RECT 5.205 2.495 5.375 2.665 ;
      RECT 5.205 3.055 5.375 3.225 ;
      RECT 5.205 3.615 5.375 3.785 ;
      RECT 4.685 3.615 4.855 3.785 ;
      RECT 4.205 1.935 4.375 2.105 ;
      RECT 3.965 2.495 4.135 2.665 ;
      RECT 3.485 2.495 3.655 2.665 ;
      RECT 3.485 3.055 3.655 3.225 ;
      RECT 3.245 1.935 3.415 2.105 ;
      RECT 2.765 3.055 2.935 3.225 ;
      RECT 2.245 2.495 2.415 2.665 ;
      RECT 2.245 3.335 2.415 3.505 ;
      RECT 1.765 1.935 1.935 2.105 ;
      RECT 1.765 3.055 1.935 3.225 ;
      RECT 1.285 3.335 1.455 3.505 ;
      RECT 1.045 2.775 1.215 2.945 ;
      RECT 0.24 2.495 0.41 2.665 ;
      RECT -0.675 1.935 -0.505 2.105 ;
      RECT -0.675 3.055 -0.505 3.225 ;
      RECT -0.915 2.495 -0.745 2.665 ;
      RECT -1.635 1.935 -1.465 2.105 ;
      RECT -1.635 3.475 -1.465 3.645 ;
      RECT -3.905 7.055 -3.735 7.225 ;
      RECT -3.905 7.795 -3.735 7.965 ;
      RECT -4.28 6.315 -4.11 6.485 ;
    LAYER li1 ;
      RECT 89.545 5.02 89.715 6.49 ;
      RECT 89.545 6.315 89.72 6.485 ;
      RECT 89.175 1.74 89.345 2.93 ;
      RECT 89.175 1.74 89.645 1.91 ;
      RECT 89.175 6.97 89.645 7.14 ;
      RECT 89.175 5.95 89.345 7.14 ;
      RECT 88.185 1.74 88.355 2.93 ;
      RECT 88.185 1.74 88.655 1.91 ;
      RECT 88.185 6.97 88.655 7.14 ;
      RECT 88.185 5.95 88.355 7.14 ;
      RECT 86.335 2.635 86.505 3.865 ;
      RECT 86.39 0.855 86.56 2.805 ;
      RECT 86.335 0.575 86.505 1.025 ;
      RECT 86.335 7.855 86.505 8.305 ;
      RECT 86.39 6.075 86.56 8.025 ;
      RECT 86.335 5.015 86.505 6.245 ;
      RECT 85.815 0.575 85.985 3.865 ;
      RECT 85.815 2.075 86.22 2.405 ;
      RECT 85.815 1.235 86.22 1.565 ;
      RECT 85.815 5.015 85.985 8.305 ;
      RECT 85.815 7.315 86.22 7.645 ;
      RECT 85.815 6.475 86.22 6.805 ;
      RECT 82.605 3.225 83.575 3.395 ;
      RECT 82.605 3.055 82.775 3.395 ;
      RECT 82.125 2.495 82.295 2.825 ;
      RECT 82.125 2.575 82.855 2.745 ;
      RECT 81.765 3.615 82.055 3.785 ;
      RECT 81.765 2.575 81.935 3.785 ;
      RECT 81.765 3.055 82.055 3.225 ;
      RECT 81.565 2.575 81.935 2.745 ;
      RECT 80.885 2.675 81.055 2.945 ;
      RECT 80.645 2.675 81.055 2.845 ;
      RECT 80.565 2.575 80.895 2.745 ;
      RECT 80.405 3.615 81.055 3.785 ;
      RECT 80.885 3.145 81.055 3.785 ;
      RECT 80.765 3.225 81.055 3.785 ;
      RECT 80.2 5.015 80.37 8.305 ;
      RECT 80.2 7.315 80.605 7.645 ;
      RECT 80.2 6.475 80.605 6.805 ;
      RECT 79.445 2.915 79.615 3.225 ;
      RECT 79.445 2.915 80.335 3.085 ;
      RECT 80.165 2.495 80.335 3.085 ;
      RECT 79.445 2.575 79.935 2.745 ;
      RECT 79.445 2.495 79.615 2.745 ;
      RECT 77.405 3.225 77.895 3.395 ;
      RECT 78.565 2.575 78.735 3.225 ;
      RECT 77.725 3.055 78.735 3.225 ;
      RECT 78.685 2.495 78.855 2.825 ;
      RECT 77.485 1.835 77.655 2.105 ;
      RECT 76.925 1.835 77.655 2.005 ;
      RECT 77.005 2.575 77.175 3.225 ;
      RECT 77.005 2.575 77.495 2.745 ;
      RECT 76.165 2.575 76.655 2.745 ;
      RECT 76.485 2.495 76.655 2.745 ;
      RECT 76.005 1.835 76.175 2.105 ;
      RECT 75.445 1.835 76.175 2.005 ;
      RECT 75.525 3.225 75.695 3.505 ;
      RECT 74.485 3.225 75.775 3.395 ;
      RECT 74.48 2.575 75.055 2.745 ;
      RECT 74.48 2.495 74.65 2.745 ;
      RECT 73.565 1.835 73.735 2.105 ;
      RECT 73.565 1.835 74.295 2.005 ;
      RECT 73.565 3.055 73.735 3.475 ;
      RECT 72.945 3.14 73.735 3.31 ;
      RECT 72.945 2.915 73.115 3.31 ;
      RECT 72.845 2.495 73.015 3.085 ;
      RECT 72.605 2.575 73.015 2.845 ;
      RECT 70.985 5.02 71.155 6.49 ;
      RECT 70.985 6.315 71.16 6.485 ;
      RECT 70.615 1.74 70.785 2.93 ;
      RECT 70.615 1.74 71.085 1.91 ;
      RECT 70.615 6.97 71.085 7.14 ;
      RECT 70.615 5.95 70.785 7.14 ;
      RECT 69.625 1.74 69.795 2.93 ;
      RECT 69.625 1.74 70.095 1.91 ;
      RECT 69.625 6.97 70.095 7.14 ;
      RECT 69.625 5.95 69.795 7.14 ;
      RECT 67.775 2.635 67.945 3.865 ;
      RECT 67.83 0.855 68 2.805 ;
      RECT 67.775 0.575 67.945 1.025 ;
      RECT 67.775 7.855 67.945 8.305 ;
      RECT 67.83 6.075 68 8.025 ;
      RECT 67.775 5.015 67.945 6.245 ;
      RECT 67.255 0.575 67.425 3.865 ;
      RECT 67.255 2.075 67.66 2.405 ;
      RECT 67.255 1.235 67.66 1.565 ;
      RECT 67.255 5.015 67.425 8.305 ;
      RECT 67.255 7.315 67.66 7.645 ;
      RECT 67.255 6.475 67.66 6.805 ;
      RECT 64.045 3.225 65.015 3.395 ;
      RECT 64.045 3.055 64.215 3.395 ;
      RECT 63.565 2.495 63.735 2.825 ;
      RECT 63.565 2.575 64.295 2.745 ;
      RECT 63.205 3.615 63.495 3.785 ;
      RECT 63.205 2.575 63.375 3.785 ;
      RECT 63.205 3.055 63.495 3.225 ;
      RECT 63.005 2.575 63.375 2.745 ;
      RECT 62.325 2.675 62.495 2.945 ;
      RECT 62.085 2.675 62.495 2.845 ;
      RECT 62.005 2.575 62.335 2.745 ;
      RECT 61.845 3.615 62.495 3.785 ;
      RECT 62.325 3.145 62.495 3.785 ;
      RECT 62.205 3.225 62.495 3.785 ;
      RECT 61.64 5.015 61.81 8.305 ;
      RECT 61.64 7.315 62.045 7.645 ;
      RECT 61.64 6.475 62.045 6.805 ;
      RECT 60.885 2.915 61.055 3.225 ;
      RECT 60.885 2.915 61.775 3.085 ;
      RECT 61.605 2.495 61.775 3.085 ;
      RECT 60.885 2.575 61.375 2.745 ;
      RECT 60.885 2.495 61.055 2.745 ;
      RECT 58.845 3.225 59.335 3.395 ;
      RECT 60.005 2.575 60.175 3.225 ;
      RECT 59.165 3.055 60.175 3.225 ;
      RECT 60.125 2.495 60.295 2.825 ;
      RECT 58.925 1.835 59.095 2.105 ;
      RECT 58.365 1.835 59.095 2.005 ;
      RECT 58.445 2.575 58.615 3.225 ;
      RECT 58.445 2.575 58.935 2.745 ;
      RECT 57.605 2.575 58.095 2.745 ;
      RECT 57.925 2.495 58.095 2.745 ;
      RECT 57.445 1.835 57.615 2.105 ;
      RECT 56.885 1.835 57.615 2.005 ;
      RECT 56.965 3.225 57.135 3.505 ;
      RECT 55.925 3.225 57.215 3.395 ;
      RECT 55.92 2.575 56.495 2.745 ;
      RECT 55.92 2.495 56.09 2.745 ;
      RECT 55.005 1.835 55.175 2.105 ;
      RECT 55.005 1.835 55.735 2.005 ;
      RECT 55.005 3.055 55.175 3.475 ;
      RECT 54.385 3.14 55.175 3.31 ;
      RECT 54.385 2.915 54.555 3.31 ;
      RECT 54.285 2.495 54.455 3.085 ;
      RECT 54.045 2.575 54.455 2.845 ;
      RECT 52.425 5.02 52.595 6.49 ;
      RECT 52.425 6.315 52.6 6.485 ;
      RECT 52.055 1.74 52.225 2.93 ;
      RECT 52.055 1.74 52.525 1.91 ;
      RECT 52.055 6.97 52.525 7.14 ;
      RECT 52.055 5.95 52.225 7.14 ;
      RECT 51.065 1.74 51.235 2.93 ;
      RECT 51.065 1.74 51.535 1.91 ;
      RECT 51.065 6.97 51.535 7.14 ;
      RECT 51.065 5.95 51.235 7.14 ;
      RECT 49.215 2.635 49.385 3.865 ;
      RECT 49.27 0.855 49.44 2.805 ;
      RECT 49.215 0.575 49.385 1.025 ;
      RECT 49.215 7.855 49.385 8.305 ;
      RECT 49.27 6.075 49.44 8.025 ;
      RECT 49.215 5.015 49.385 6.245 ;
      RECT 48.695 0.575 48.865 3.865 ;
      RECT 48.695 2.075 49.1 2.405 ;
      RECT 48.695 1.235 49.1 1.565 ;
      RECT 48.695 5.015 48.865 8.305 ;
      RECT 48.695 7.315 49.1 7.645 ;
      RECT 48.695 6.475 49.1 6.805 ;
      RECT 45.485 3.225 46.455 3.395 ;
      RECT 45.485 3.055 45.655 3.395 ;
      RECT 45.005 2.495 45.175 2.825 ;
      RECT 45.005 2.575 45.735 2.745 ;
      RECT 44.645 3.615 44.935 3.785 ;
      RECT 44.645 2.575 44.815 3.785 ;
      RECT 44.645 3.055 44.935 3.225 ;
      RECT 44.445 2.575 44.815 2.745 ;
      RECT 43.765 2.675 43.935 2.945 ;
      RECT 43.525 2.675 43.935 2.845 ;
      RECT 43.445 2.575 43.775 2.745 ;
      RECT 43.285 3.615 43.935 3.785 ;
      RECT 43.765 3.145 43.935 3.785 ;
      RECT 43.645 3.225 43.935 3.785 ;
      RECT 43.08 5.015 43.25 8.305 ;
      RECT 43.08 7.315 43.485 7.645 ;
      RECT 43.08 6.475 43.485 6.805 ;
      RECT 42.325 2.915 42.495 3.225 ;
      RECT 42.325 2.915 43.215 3.085 ;
      RECT 43.045 2.495 43.215 3.085 ;
      RECT 42.325 2.575 42.815 2.745 ;
      RECT 42.325 2.495 42.495 2.745 ;
      RECT 40.285 3.225 40.775 3.395 ;
      RECT 41.445 2.575 41.615 3.225 ;
      RECT 40.605 3.055 41.615 3.225 ;
      RECT 41.565 2.495 41.735 2.825 ;
      RECT 40.365 1.835 40.535 2.105 ;
      RECT 39.805 1.835 40.535 2.005 ;
      RECT 39.885 2.575 40.055 3.225 ;
      RECT 39.885 2.575 40.375 2.745 ;
      RECT 39.045 2.575 39.535 2.745 ;
      RECT 39.365 2.495 39.535 2.745 ;
      RECT 38.885 1.835 39.055 2.105 ;
      RECT 38.325 1.835 39.055 2.005 ;
      RECT 38.405 3.225 38.575 3.505 ;
      RECT 37.365 3.225 38.655 3.395 ;
      RECT 37.36 2.575 37.935 2.745 ;
      RECT 37.36 2.495 37.53 2.745 ;
      RECT 36.445 1.835 36.615 2.105 ;
      RECT 36.445 1.835 37.175 2.005 ;
      RECT 36.445 3.055 36.615 3.475 ;
      RECT 35.825 3.14 36.615 3.31 ;
      RECT 35.825 2.915 35.995 3.31 ;
      RECT 35.725 2.495 35.895 3.085 ;
      RECT 35.485 2.575 35.895 2.845 ;
      RECT 33.865 5.02 34.035 6.49 ;
      RECT 33.865 6.315 34.04 6.485 ;
      RECT 33.495 1.74 33.665 2.93 ;
      RECT 33.495 1.74 33.965 1.91 ;
      RECT 33.495 6.97 33.965 7.14 ;
      RECT 33.495 5.95 33.665 7.14 ;
      RECT 32.505 1.74 32.675 2.93 ;
      RECT 32.505 1.74 32.975 1.91 ;
      RECT 32.505 6.97 32.975 7.14 ;
      RECT 32.505 5.95 32.675 7.14 ;
      RECT 30.655 2.635 30.825 3.865 ;
      RECT 30.71 0.855 30.88 2.805 ;
      RECT 30.655 0.575 30.825 1.025 ;
      RECT 30.655 7.855 30.825 8.305 ;
      RECT 30.71 6.075 30.88 8.025 ;
      RECT 30.655 5.015 30.825 6.245 ;
      RECT 30.135 0.575 30.305 3.865 ;
      RECT 30.135 2.075 30.54 2.405 ;
      RECT 30.135 1.235 30.54 1.565 ;
      RECT 30.135 5.015 30.305 8.305 ;
      RECT 30.135 7.315 30.54 7.645 ;
      RECT 30.135 6.475 30.54 6.805 ;
      RECT 26.925 3.225 27.895 3.395 ;
      RECT 26.925 3.055 27.095 3.395 ;
      RECT 26.445 2.495 26.615 2.825 ;
      RECT 26.445 2.575 27.175 2.745 ;
      RECT 26.085 3.615 26.375 3.785 ;
      RECT 26.085 2.575 26.255 3.785 ;
      RECT 26.085 3.055 26.375 3.225 ;
      RECT 25.885 2.575 26.255 2.745 ;
      RECT 25.205 2.675 25.375 2.945 ;
      RECT 24.965 2.675 25.375 2.845 ;
      RECT 24.885 2.575 25.215 2.745 ;
      RECT 24.725 3.615 25.375 3.785 ;
      RECT 25.205 3.145 25.375 3.785 ;
      RECT 25.085 3.225 25.375 3.785 ;
      RECT 24.52 5.015 24.69 8.305 ;
      RECT 24.52 7.315 24.925 7.645 ;
      RECT 24.52 6.475 24.925 6.805 ;
      RECT 23.765 2.915 23.935 3.225 ;
      RECT 23.765 2.915 24.655 3.085 ;
      RECT 24.485 2.495 24.655 3.085 ;
      RECT 23.765 2.575 24.255 2.745 ;
      RECT 23.765 2.495 23.935 2.745 ;
      RECT 21.725 3.225 22.215 3.395 ;
      RECT 22.885 2.575 23.055 3.225 ;
      RECT 22.045 3.055 23.055 3.225 ;
      RECT 23.005 2.495 23.175 2.825 ;
      RECT 21.805 1.835 21.975 2.105 ;
      RECT 21.245 1.835 21.975 2.005 ;
      RECT 21.325 2.575 21.495 3.225 ;
      RECT 21.325 2.575 21.815 2.745 ;
      RECT 20.485 2.575 20.975 2.745 ;
      RECT 20.805 2.495 20.975 2.745 ;
      RECT 20.325 1.835 20.495 2.105 ;
      RECT 19.765 1.835 20.495 2.005 ;
      RECT 19.845 3.225 20.015 3.505 ;
      RECT 18.805 3.225 20.095 3.395 ;
      RECT 18.8 2.575 19.375 2.745 ;
      RECT 18.8 2.495 18.97 2.745 ;
      RECT 17.885 1.835 18.055 2.105 ;
      RECT 17.885 1.835 18.615 2.005 ;
      RECT 17.885 3.055 18.055 3.475 ;
      RECT 17.265 3.14 18.055 3.31 ;
      RECT 17.265 2.915 17.435 3.31 ;
      RECT 17.165 2.495 17.335 3.085 ;
      RECT 16.925 2.575 17.335 2.845 ;
      RECT 15.305 5.02 15.475 6.49 ;
      RECT 15.305 6.315 15.48 6.485 ;
      RECT 14.935 1.74 15.105 2.93 ;
      RECT 14.935 1.74 15.405 1.91 ;
      RECT 14.935 6.97 15.405 7.14 ;
      RECT 14.935 5.95 15.105 7.14 ;
      RECT 13.945 1.74 14.115 2.93 ;
      RECT 13.945 1.74 14.415 1.91 ;
      RECT 13.945 6.97 14.415 7.14 ;
      RECT 13.945 5.95 14.115 7.14 ;
      RECT 12.095 2.635 12.265 3.865 ;
      RECT 12.15 0.855 12.32 2.805 ;
      RECT 12.095 0.575 12.265 1.025 ;
      RECT 12.095 7.855 12.265 8.305 ;
      RECT 12.15 6.075 12.32 8.025 ;
      RECT 12.095 5.015 12.265 6.245 ;
      RECT 11.575 0.575 11.745 3.865 ;
      RECT 11.575 2.075 11.98 2.405 ;
      RECT 11.575 1.235 11.98 1.565 ;
      RECT 11.575 5.015 11.745 8.305 ;
      RECT 11.575 7.315 11.98 7.645 ;
      RECT 11.575 6.475 11.98 6.805 ;
      RECT 8.365 3.225 9.335 3.395 ;
      RECT 8.365 3.055 8.535 3.395 ;
      RECT 7.885 2.495 8.055 2.825 ;
      RECT 7.885 2.575 8.615 2.745 ;
      RECT 7.525 3.615 7.815 3.785 ;
      RECT 7.525 2.575 7.695 3.785 ;
      RECT 7.525 3.055 7.815 3.225 ;
      RECT 7.325 2.575 7.695 2.745 ;
      RECT 6.645 2.675 6.815 2.945 ;
      RECT 6.405 2.675 6.815 2.845 ;
      RECT 6.325 2.575 6.655 2.745 ;
      RECT 6.165 3.615 6.815 3.785 ;
      RECT 6.645 3.145 6.815 3.785 ;
      RECT 6.525 3.225 6.815 3.785 ;
      RECT 5.96 5.015 6.13 8.305 ;
      RECT 5.96 7.315 6.365 7.645 ;
      RECT 5.96 6.475 6.365 6.805 ;
      RECT 5.205 2.915 5.375 3.225 ;
      RECT 5.205 2.915 6.095 3.085 ;
      RECT 5.925 2.495 6.095 3.085 ;
      RECT 5.205 2.575 5.695 2.745 ;
      RECT 5.205 2.495 5.375 2.745 ;
      RECT 3.165 3.225 3.655 3.395 ;
      RECT 4.325 2.575 4.495 3.225 ;
      RECT 3.485 3.055 4.495 3.225 ;
      RECT 4.445 2.495 4.615 2.825 ;
      RECT 3.245 1.835 3.415 2.105 ;
      RECT 2.685 1.835 3.415 2.005 ;
      RECT 2.765 2.575 2.935 3.225 ;
      RECT 2.765 2.575 3.255 2.745 ;
      RECT 1.925 2.575 2.415 2.745 ;
      RECT 2.245 2.495 2.415 2.745 ;
      RECT 1.765 1.835 1.935 2.105 ;
      RECT 1.205 1.835 1.935 2.005 ;
      RECT 1.285 3.225 1.455 3.505 ;
      RECT 0.245 3.225 1.535 3.395 ;
      RECT 0.24 2.575 0.815 2.745 ;
      RECT 0.24 2.495 0.41 2.745 ;
      RECT -0.675 1.835 -0.505 2.105 ;
      RECT -0.675 1.835 0.055 2.005 ;
      RECT -0.675 3.055 -0.505 3.475 ;
      RECT -1.295 3.14 -0.505 3.31 ;
      RECT -1.295 2.915 -1.125 3.31 ;
      RECT -1.395 2.495 -1.225 3.085 ;
      RECT -1.635 2.575 -1.225 2.845 ;
      RECT -4.335 7.855 -4.165 8.305 ;
      RECT -4.28 6.075 -4.11 8.025 ;
      RECT -4.335 5.015 -4.165 6.245 ;
      RECT -4.855 5.015 -4.685 8.305 ;
      RECT -4.855 7.315 -4.45 7.645 ;
      RECT -4.855 6.475 -4.45 6.805 ;
      RECT 89.545 7.8 89.715 8.31 ;
      RECT 88.555 0.57 88.725 1.08 ;
      RECT 88.555 2.39 88.725 3.86 ;
      RECT 88.555 5.02 88.725 6.49 ;
      RECT 88.555 7.8 88.725 8.31 ;
      RECT 87.195 0.575 87.365 3.865 ;
      RECT 87.195 5.015 87.365 8.305 ;
      RECT 86.765 0.575 86.935 1.085 ;
      RECT 86.765 1.655 86.935 3.865 ;
      RECT 86.765 5.015 86.935 7.225 ;
      RECT 86.765 7.795 86.935 8.305 ;
      RECT 83.085 2.495 83.255 2.945 ;
      RECT 82.845 1.755 83.015 2.105 ;
      RECT 81.885 1.755 82.055 2.105 ;
      RECT 81.58 5.015 81.75 8.305 ;
      RECT 81.405 3.055 81.575 3.475 ;
      RECT 81.15 5.015 81.32 7.225 ;
      RECT 81.15 7.795 81.32 8.305 ;
      RECT 80.405 1.755 80.575 2.105 ;
      RECT 79.445 1.755 79.615 2.105 ;
      RECT 79.445 3.485 79.615 3.815 ;
      RECT 78.925 3.145 79.095 3.785 ;
      RECT 78.445 1.755 78.615 2.105 ;
      RECT 78.205 2.495 78.375 2.825 ;
      RECT 77.725 2.495 77.895 2.825 ;
      RECT 76.485 3.145 76.655 3.505 ;
      RECT 76.005 3.055 76.175 3.475 ;
      RECT 75.285 2.495 75.455 2.945 ;
      RECT 73.325 2.495 73.495 2.825 ;
      RECT 72.605 1.755 72.775 2.105 ;
      RECT 72.605 3.285 72.775 3.645 ;
      RECT 70.985 7.8 71.155 8.31 ;
      RECT 69.995 0.57 70.165 1.08 ;
      RECT 69.995 2.39 70.165 3.86 ;
      RECT 69.995 5.02 70.165 6.49 ;
      RECT 69.995 7.8 70.165 8.31 ;
      RECT 68.635 0.575 68.805 3.865 ;
      RECT 68.635 5.015 68.805 8.305 ;
      RECT 68.205 0.575 68.375 1.085 ;
      RECT 68.205 1.655 68.375 3.865 ;
      RECT 68.205 5.015 68.375 7.225 ;
      RECT 68.205 7.795 68.375 8.305 ;
      RECT 64.525 2.495 64.695 2.945 ;
      RECT 64.285 1.755 64.455 2.105 ;
      RECT 63.325 1.755 63.495 2.105 ;
      RECT 63.02 5.015 63.19 8.305 ;
      RECT 62.845 3.055 63.015 3.475 ;
      RECT 62.59 5.015 62.76 7.225 ;
      RECT 62.59 7.795 62.76 8.305 ;
      RECT 61.845 1.755 62.015 2.105 ;
      RECT 60.885 1.755 61.055 2.105 ;
      RECT 60.885 3.485 61.055 3.815 ;
      RECT 60.365 3.145 60.535 3.785 ;
      RECT 59.885 1.755 60.055 2.105 ;
      RECT 59.645 2.495 59.815 2.825 ;
      RECT 59.165 2.495 59.335 2.825 ;
      RECT 57.925 3.145 58.095 3.505 ;
      RECT 57.445 3.055 57.615 3.475 ;
      RECT 56.725 2.495 56.895 2.945 ;
      RECT 54.765 2.495 54.935 2.825 ;
      RECT 54.045 1.755 54.215 2.105 ;
      RECT 54.045 3.285 54.215 3.645 ;
      RECT 52.425 7.8 52.595 8.31 ;
      RECT 51.435 0.57 51.605 1.08 ;
      RECT 51.435 2.39 51.605 3.86 ;
      RECT 51.435 5.02 51.605 6.49 ;
      RECT 51.435 7.8 51.605 8.31 ;
      RECT 50.075 0.575 50.245 3.865 ;
      RECT 50.075 5.015 50.245 8.305 ;
      RECT 49.645 0.575 49.815 1.085 ;
      RECT 49.645 1.655 49.815 3.865 ;
      RECT 49.645 5.015 49.815 7.225 ;
      RECT 49.645 7.795 49.815 8.305 ;
      RECT 45.965 2.495 46.135 2.945 ;
      RECT 45.725 1.755 45.895 2.105 ;
      RECT 44.765 1.755 44.935 2.105 ;
      RECT 44.46 5.015 44.63 8.305 ;
      RECT 44.285 3.055 44.455 3.475 ;
      RECT 44.03 5.015 44.2 7.225 ;
      RECT 44.03 7.795 44.2 8.305 ;
      RECT 43.285 1.755 43.455 2.105 ;
      RECT 42.325 1.755 42.495 2.105 ;
      RECT 42.325 3.485 42.495 3.815 ;
      RECT 41.805 3.145 41.975 3.785 ;
      RECT 41.325 1.755 41.495 2.105 ;
      RECT 41.085 2.495 41.255 2.825 ;
      RECT 40.605 2.495 40.775 2.825 ;
      RECT 39.365 3.145 39.535 3.505 ;
      RECT 38.885 3.055 39.055 3.475 ;
      RECT 38.165 2.495 38.335 2.945 ;
      RECT 36.205 2.495 36.375 2.825 ;
      RECT 35.485 1.755 35.655 2.105 ;
      RECT 35.485 3.285 35.655 3.645 ;
      RECT 33.865 7.8 34.035 8.31 ;
      RECT 32.875 0.57 33.045 1.08 ;
      RECT 32.875 2.39 33.045 3.86 ;
      RECT 32.875 5.02 33.045 6.49 ;
      RECT 32.875 7.8 33.045 8.31 ;
      RECT 31.515 0.575 31.685 3.865 ;
      RECT 31.515 5.015 31.685 8.305 ;
      RECT 31.085 0.575 31.255 1.085 ;
      RECT 31.085 1.655 31.255 3.865 ;
      RECT 31.085 5.015 31.255 7.225 ;
      RECT 31.085 7.795 31.255 8.305 ;
      RECT 27.405 2.495 27.575 2.945 ;
      RECT 27.165 1.755 27.335 2.105 ;
      RECT 26.205 1.755 26.375 2.105 ;
      RECT 25.9 5.015 26.07 8.305 ;
      RECT 25.725 3.055 25.895 3.475 ;
      RECT 25.47 5.015 25.64 7.225 ;
      RECT 25.47 7.795 25.64 8.305 ;
      RECT 24.725 1.755 24.895 2.105 ;
      RECT 23.765 1.755 23.935 2.105 ;
      RECT 23.765 3.485 23.935 3.815 ;
      RECT 23.245 3.145 23.415 3.785 ;
      RECT 22.765 1.755 22.935 2.105 ;
      RECT 22.525 2.495 22.695 2.825 ;
      RECT 22.045 2.495 22.215 2.825 ;
      RECT 20.805 3.145 20.975 3.505 ;
      RECT 20.325 3.055 20.495 3.475 ;
      RECT 19.605 2.495 19.775 2.945 ;
      RECT 17.645 2.495 17.815 2.825 ;
      RECT 16.925 1.755 17.095 2.105 ;
      RECT 16.925 3.285 17.095 3.645 ;
      RECT 15.305 7.8 15.475 8.31 ;
      RECT 14.315 0.57 14.485 1.08 ;
      RECT 14.315 2.39 14.485 3.86 ;
      RECT 14.315 5.02 14.485 6.49 ;
      RECT 14.315 7.8 14.485 8.31 ;
      RECT 12.955 0.575 13.125 3.865 ;
      RECT 12.955 5.015 13.125 8.305 ;
      RECT 12.525 0.575 12.695 1.085 ;
      RECT 12.525 1.655 12.695 3.865 ;
      RECT 12.525 5.015 12.695 7.225 ;
      RECT 12.525 7.795 12.695 8.305 ;
      RECT 8.845 2.495 9.015 2.945 ;
      RECT 8.605 1.755 8.775 2.105 ;
      RECT 7.645 1.755 7.815 2.105 ;
      RECT 7.34 5.015 7.51 8.305 ;
      RECT 7.165 3.055 7.335 3.475 ;
      RECT 6.91 5.015 7.08 7.225 ;
      RECT 6.91 7.795 7.08 8.305 ;
      RECT 6.165 1.755 6.335 2.105 ;
      RECT 5.205 1.755 5.375 2.105 ;
      RECT 5.205 3.485 5.375 3.815 ;
      RECT 4.685 3.145 4.855 3.785 ;
      RECT 4.205 1.755 4.375 2.105 ;
      RECT 3.965 2.495 4.135 2.825 ;
      RECT 3.485 2.495 3.655 2.825 ;
      RECT 2.245 3.145 2.415 3.505 ;
      RECT 1.765 3.055 1.935 3.475 ;
      RECT 1.045 2.495 1.215 2.945 ;
      RECT -0.915 2.495 -0.745 2.825 ;
      RECT -1.635 1.755 -1.465 2.105 ;
      RECT -1.635 3.285 -1.465 3.645 ;
      RECT -3.905 5.015 -3.735 7.225 ;
      RECT -3.905 7.795 -3.735 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2et_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2et_8_b0r2
  CLASS BLOCK ;
  ORIGIN 5.505 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2et_8_b0r2 ;
  SIZE 95.595 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 15.31 0.915 15.48 1.085 ;
        RECT 15.305 0.91 15.475 1.08 ;
        RECT 15.305 2.39 15.475 2.56 ;
      LAYER li1 ;
        RECT 15.31 0.915 15.48 1.085 ;
        RECT 15.305 0.57 15.475 1.08 ;
        RECT 15.305 2.39 15.475 3.86 ;
      LAYER met1 ;
        RECT 15.245 2.36 15.535 2.59 ;
        RECT 15.245 0.88 15.535 1.11 ;
        RECT 15.305 0.88 15.475 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 33.87 0.915 34.04 1.085 ;
        RECT 33.865 0.91 34.035 1.08 ;
        RECT 33.865 2.39 34.035 2.56 ;
      LAYER li1 ;
        RECT 33.87 0.915 34.04 1.085 ;
        RECT 33.865 0.57 34.035 1.08 ;
        RECT 33.865 2.39 34.035 3.86 ;
      LAYER met1 ;
        RECT 33.805 2.36 34.095 2.59 ;
        RECT 33.805 0.88 34.095 1.11 ;
        RECT 33.865 0.88 34.035 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 52.43 0.915 52.6 1.085 ;
        RECT 52.425 0.91 52.595 1.08 ;
        RECT 52.425 2.39 52.595 2.56 ;
      LAYER li1 ;
        RECT 52.43 0.915 52.6 1.085 ;
        RECT 52.425 0.57 52.595 1.08 ;
        RECT 52.425 2.39 52.595 3.86 ;
      LAYER met1 ;
        RECT 52.365 2.36 52.655 2.59 ;
        RECT 52.365 0.88 52.655 1.11 ;
        RECT 52.425 0.88 52.595 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 70.99 0.915 71.16 1.085 ;
        RECT 70.985 0.91 71.155 1.08 ;
        RECT 70.985 2.39 71.155 2.56 ;
      LAYER li1 ;
        RECT 70.99 0.915 71.16 1.085 ;
        RECT 70.985 0.57 71.155 1.08 ;
        RECT 70.985 2.39 71.155 3.86 ;
      LAYER met1 ;
        RECT 70.925 2.36 71.215 2.59 ;
        RECT 70.925 0.88 71.215 1.11 ;
        RECT 70.985 0.88 71.155 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 89.55 0.915 89.72 1.085 ;
        RECT 89.545 0.91 89.715 1.08 ;
        RECT 89.545 2.39 89.715 2.56 ;
      LAYER li1 ;
        RECT 89.55 0.915 89.72 1.085 ;
        RECT 89.545 0.57 89.715 1.08 ;
        RECT 89.545 2.39 89.715 3.86 ;
      LAYER met1 ;
        RECT 89.485 2.36 89.775 2.59 ;
        RECT 89.485 0.88 89.775 1.11 ;
        RECT 89.545 0.88 89.715 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 11.155 1.66 11.325 2.935 ;
        RECT 11.155 5.945 11.325 7.22 ;
        RECT 5.54 5.945 5.71 7.22 ;
      LAYER met2 ;
        RECT 11.08 2.705 11.42 3.055 ;
        RECT 11.07 5.845 11.41 6.195 ;
        RECT 11.155 2.705 11.325 6.195 ;
      LAYER met1 ;
        RECT 11.08 2.765 11.555 2.935 ;
        RECT 11.08 2.705 11.42 3.055 ;
        RECT 5.48 5.945 11.555 6.115 ;
        RECT 11.07 5.845 11.41 6.195 ;
        RECT 5.48 5.915 5.77 6.145 ;
      LAYER via1 ;
        RECT 11.17 5.945 11.32 6.095 ;
        RECT 11.18 2.805 11.33 2.955 ;
      LAYER mcon ;
        RECT 5.54 5.945 5.71 6.115 ;
        RECT 11.155 5.945 11.325 6.115 ;
        RECT 11.155 2.765 11.325 2.935 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 29.715 1.66 29.885 2.935 ;
        RECT 29.715 5.945 29.885 7.22 ;
        RECT 24.1 5.945 24.27 7.22 ;
      LAYER met2 ;
        RECT 29.64 2.705 29.98 3.055 ;
        RECT 29.63 5.845 29.97 6.195 ;
        RECT 29.715 2.705 29.885 6.195 ;
      LAYER met1 ;
        RECT 29.64 2.765 30.115 2.935 ;
        RECT 29.64 2.705 29.98 3.055 ;
        RECT 24.04 5.945 30.115 6.115 ;
        RECT 29.63 5.845 29.97 6.195 ;
        RECT 24.04 5.915 24.33 6.145 ;
      LAYER via1 ;
        RECT 29.73 5.945 29.88 6.095 ;
        RECT 29.74 2.805 29.89 2.955 ;
      LAYER mcon ;
        RECT 24.1 5.945 24.27 6.115 ;
        RECT 29.715 5.945 29.885 6.115 ;
        RECT 29.715 2.765 29.885 2.935 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 48.275 1.66 48.445 2.935 ;
        RECT 48.275 5.945 48.445 7.22 ;
        RECT 42.66 5.945 42.83 7.22 ;
      LAYER met2 ;
        RECT 48.2 2.705 48.54 3.055 ;
        RECT 48.19 5.845 48.53 6.195 ;
        RECT 48.275 2.705 48.445 6.195 ;
      LAYER met1 ;
        RECT 48.2 2.765 48.675 2.935 ;
        RECT 48.2 2.705 48.54 3.055 ;
        RECT 42.6 5.945 48.675 6.115 ;
        RECT 48.19 5.845 48.53 6.195 ;
        RECT 42.6 5.915 42.89 6.145 ;
      LAYER via1 ;
        RECT 48.29 5.945 48.44 6.095 ;
        RECT 48.3 2.805 48.45 2.955 ;
      LAYER mcon ;
        RECT 42.66 5.945 42.83 6.115 ;
        RECT 48.275 5.945 48.445 6.115 ;
        RECT 48.275 2.765 48.445 2.935 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 66.835 1.66 67.005 2.935 ;
        RECT 66.835 5.945 67.005 7.22 ;
        RECT 61.22 5.945 61.39 7.22 ;
      LAYER met2 ;
        RECT 66.76 2.705 67.1 3.055 ;
        RECT 66.75 5.845 67.09 6.195 ;
        RECT 66.835 2.705 67.005 6.195 ;
      LAYER met1 ;
        RECT 66.76 2.765 67.235 2.935 ;
        RECT 66.76 2.705 67.1 3.055 ;
        RECT 61.16 5.945 67.235 6.115 ;
        RECT 66.75 5.845 67.09 6.195 ;
        RECT 61.16 5.915 61.45 6.145 ;
      LAYER via1 ;
        RECT 66.85 5.945 67 6.095 ;
        RECT 66.86 2.805 67.01 2.955 ;
      LAYER mcon ;
        RECT 61.22 5.945 61.39 6.115 ;
        RECT 66.835 5.945 67.005 6.115 ;
        RECT 66.835 2.765 67.005 2.935 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER li1 ;
        RECT 85.395 1.66 85.565 2.935 ;
        RECT 85.395 5.945 85.565 7.22 ;
        RECT 79.78 5.945 79.95 7.22 ;
      LAYER met2 ;
        RECT 85.32 2.705 85.66 3.055 ;
        RECT 85.31 5.845 85.65 6.195 ;
        RECT 85.395 2.705 85.565 6.195 ;
      LAYER met1 ;
        RECT 85.32 2.765 85.795 2.935 ;
        RECT 85.32 2.705 85.66 3.055 ;
        RECT 79.72 5.945 85.795 6.115 ;
        RECT 85.31 5.845 85.65 6.195 ;
        RECT 79.72 5.915 80.01 6.145 ;
      LAYER via1 ;
        RECT 85.41 5.945 85.56 6.095 ;
        RECT 85.42 2.805 85.57 2.955 ;
      LAYER mcon ;
        RECT 79.78 5.945 79.95 6.115 ;
        RECT 85.395 5.945 85.565 6.115 ;
        RECT 85.395 2.765 85.565 2.935 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT -5.275 5.945 -5.105 7.22 ;
      LAYER met1 ;
        RECT -5.365 5.945 -4.875 6.115 ;
        RECT -5.365 5.905 -5.025 6.165 ;
      LAYER mcon ;
        RECT -5.275 5.945 -5.105 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 72.275 4.135 90.09 4.745 ;
        RECT 87.955 4.13 89.935 4.75 ;
        RECT 89.115 3.4 89.285 5.48 ;
        RECT 88.125 3.4 88.295 5.48 ;
        RECT 85.385 3.405 85.555 5.475 ;
        RECT 82.365 3.635 82.535 4.745 ;
        RECT 79.925 3.635 80.095 4.745 ;
        RECT 79.77 4.135 79.94 5.475 ;
        RECT 77.965 3.635 78.135 4.745 ;
        RECT 77.005 3.635 77.175 4.745 ;
        RECT 75.045 3.635 75.215 4.745 ;
        RECT 74.045 3.635 74.215 4.745 ;
        RECT 71.53 4.145 73.995 4.75 ;
        RECT 73.085 3.635 73.255 4.75 ;
        RECT 53.715 4.135 71.53 4.745 ;
        RECT 69.395 4.13 71.375 4.75 ;
        RECT 70.555 3.4 70.725 5.48 ;
        RECT 69.565 3.4 69.735 5.48 ;
        RECT 66.825 3.405 66.995 5.475 ;
        RECT 63.805 3.635 63.975 4.745 ;
        RECT 61.365 3.635 61.535 4.745 ;
        RECT 61.21 4.135 61.38 5.475 ;
        RECT 59.405 3.635 59.575 4.745 ;
        RECT 58.445 3.635 58.615 4.745 ;
        RECT 56.485 3.635 56.655 4.745 ;
        RECT 55.485 3.635 55.655 4.745 ;
        RECT 52.97 4.145 55.435 4.75 ;
        RECT 54.525 3.635 54.695 4.75 ;
        RECT 35.155 4.135 52.97 4.745 ;
        RECT 50.835 4.13 52.815 4.75 ;
        RECT 51.995 3.4 52.165 5.48 ;
        RECT 51.005 3.4 51.175 5.48 ;
        RECT 48.265 3.405 48.435 5.475 ;
        RECT 45.245 3.635 45.415 4.745 ;
        RECT 42.805 3.635 42.975 4.745 ;
        RECT 42.65 4.135 42.82 5.475 ;
        RECT 40.845 3.635 41.015 4.745 ;
        RECT 39.885 3.635 40.055 4.745 ;
        RECT 37.925 3.635 38.095 4.745 ;
        RECT 36.925 3.635 37.095 4.745 ;
        RECT 34.41 4.145 36.875 4.75 ;
        RECT 35.965 3.635 36.135 4.75 ;
        RECT 16.595 4.135 34.41 4.745 ;
        RECT 32.275 4.13 34.255 4.75 ;
        RECT 33.435 3.4 33.605 5.48 ;
        RECT 32.445 3.4 32.615 5.48 ;
        RECT 29.705 3.405 29.875 5.475 ;
        RECT 26.685 3.635 26.855 4.745 ;
        RECT 24.245 3.635 24.415 4.745 ;
        RECT 24.09 4.135 24.26 5.475 ;
        RECT 22.285 3.635 22.455 4.745 ;
        RECT 21.325 3.635 21.495 4.745 ;
        RECT 19.365 3.635 19.535 4.745 ;
        RECT 18.365 3.635 18.535 4.745 ;
        RECT 15.85 4.145 18.315 4.75 ;
        RECT 17.405 3.635 17.575 4.75 ;
        RECT -1.965 4.135 15.85 4.745 ;
        RECT 13.715 4.13 15.695 4.75 ;
        RECT 14.875 3.4 15.045 5.48 ;
        RECT 13.885 3.4 14.055 5.48 ;
        RECT 11.145 3.405 11.315 5.475 ;
        RECT 8.125 3.635 8.295 4.745 ;
        RECT 5.685 3.635 5.855 4.745 ;
        RECT 5.53 4.135 5.7 5.475 ;
        RECT 3.725 3.635 3.895 4.745 ;
        RECT 2.765 3.635 2.935 4.745 ;
        RECT 0.805 3.635 0.975 4.745 ;
        RECT -0.195 3.635 -0.025 4.745 ;
        RECT -5.505 4.145 -0.245 4.75 ;
        RECT -1.155 3.635 -0.985 4.75 ;
        RECT -3.475 4.145 -3.305 8.305 ;
        RECT -5.285 4.145 -5.115 5.475 ;
      LAYER met1 ;
        RECT 72.275 4.135 90.09 4.745 ;
        RECT 87.955 4.13 89.935 4.75 ;
        RECT 72.275 3.98 84.235 4.745 ;
        RECT 71.53 4.145 73.995 4.75 ;
        RECT 53.715 4.135 71.53 4.745 ;
        RECT 69.395 4.13 71.375 4.75 ;
        RECT 53.715 3.98 65.675 4.745 ;
        RECT 52.97 4.145 55.435 4.75 ;
        RECT 35.155 4.135 52.97 4.745 ;
        RECT 50.835 4.13 52.815 4.75 ;
        RECT 35.155 3.98 47.115 4.745 ;
        RECT 34.41 4.145 36.875 4.75 ;
        RECT 16.595 4.135 34.41 4.745 ;
        RECT 32.275 4.13 34.255 4.75 ;
        RECT 16.595 3.98 28.555 4.745 ;
        RECT 15.85 4.145 18.315 4.75 ;
        RECT -1.965 4.135 15.85 4.745 ;
        RECT 13.715 4.13 15.695 4.75 ;
        RECT -1.965 3.98 9.995 4.745 ;
        RECT -5.505 4.145 -0.245 4.75 ;
        RECT -3.535 6.655 -3.245 6.885 ;
        RECT -3.705 6.685 -3.245 6.855 ;
      LAYER mcon ;
        RECT -3.475 6.685 -3.305 6.855 ;
        RECT -3.165 4.545 -2.995 4.715 ;
        RECT -1.82 4.135 -1.65 4.305 ;
        RECT -1.36 4.135 -1.19 4.305 ;
        RECT -0.9 4.135 -0.73 4.305 ;
        RECT -0.44 4.135 -0.27 4.305 ;
        RECT 0.02 4.135 0.19 4.305 ;
        RECT 0.48 4.135 0.65 4.305 ;
        RECT 0.94 4.135 1.11 4.305 ;
        RECT 1.4 4.135 1.57 4.305 ;
        RECT 1.86 4.135 2.03 4.305 ;
        RECT 2.32 4.135 2.49 4.305 ;
        RECT 2.78 4.135 2.95 4.305 ;
        RECT 3.24 4.135 3.41 4.305 ;
        RECT 3.7 4.135 3.87 4.305 ;
        RECT 4.16 4.135 4.33 4.305 ;
        RECT 4.62 4.135 4.79 4.305 ;
        RECT 5.08 4.135 5.25 4.305 ;
        RECT 5.54 4.135 5.71 4.305 ;
        RECT 6 4.135 6.17 4.305 ;
        RECT 6.46 4.135 6.63 4.305 ;
        RECT 6.92 4.135 7.09 4.305 ;
        RECT 7.38 4.135 7.55 4.305 ;
        RECT 7.65 4.545 7.82 4.715 ;
        RECT 7.84 4.135 8.01 4.305 ;
        RECT 8.3 4.135 8.47 4.305 ;
        RECT 8.76 4.135 8.93 4.305 ;
        RECT 9.22 4.135 9.39 4.305 ;
        RECT 9.68 4.135 9.85 4.305 ;
        RECT 13.265 4.545 13.435 4.715 ;
        RECT 13.265 4.165 13.435 4.335 ;
        RECT 13.965 4.55 14.135 4.72 ;
        RECT 13.965 4.16 14.135 4.33 ;
        RECT 14.955 4.55 15.125 4.72 ;
        RECT 14.955 4.16 15.125 4.33 ;
        RECT 16.74 4.135 16.91 4.305 ;
        RECT 17.2 4.135 17.37 4.305 ;
        RECT 17.66 4.135 17.83 4.305 ;
        RECT 18.12 4.135 18.29 4.305 ;
        RECT 18.58 4.135 18.75 4.305 ;
        RECT 19.04 4.135 19.21 4.305 ;
        RECT 19.5 4.135 19.67 4.305 ;
        RECT 19.96 4.135 20.13 4.305 ;
        RECT 20.42 4.135 20.59 4.305 ;
        RECT 20.88 4.135 21.05 4.305 ;
        RECT 21.34 4.135 21.51 4.305 ;
        RECT 21.8 4.135 21.97 4.305 ;
        RECT 22.26 4.135 22.43 4.305 ;
        RECT 22.72 4.135 22.89 4.305 ;
        RECT 23.18 4.135 23.35 4.305 ;
        RECT 23.64 4.135 23.81 4.305 ;
        RECT 24.1 4.135 24.27 4.305 ;
        RECT 24.56 4.135 24.73 4.305 ;
        RECT 25.02 4.135 25.19 4.305 ;
        RECT 25.48 4.135 25.65 4.305 ;
        RECT 25.94 4.135 26.11 4.305 ;
        RECT 26.21 4.545 26.38 4.715 ;
        RECT 26.4 4.135 26.57 4.305 ;
        RECT 26.86 4.135 27.03 4.305 ;
        RECT 27.32 4.135 27.49 4.305 ;
        RECT 27.78 4.135 27.95 4.305 ;
        RECT 28.24 4.135 28.41 4.305 ;
        RECT 31.825 4.545 31.995 4.715 ;
        RECT 31.825 4.165 31.995 4.335 ;
        RECT 32.525 4.55 32.695 4.72 ;
        RECT 32.525 4.16 32.695 4.33 ;
        RECT 33.515 4.55 33.685 4.72 ;
        RECT 33.515 4.16 33.685 4.33 ;
        RECT 35.3 4.135 35.47 4.305 ;
        RECT 35.76 4.135 35.93 4.305 ;
        RECT 36.22 4.135 36.39 4.305 ;
        RECT 36.68 4.135 36.85 4.305 ;
        RECT 37.14 4.135 37.31 4.305 ;
        RECT 37.6 4.135 37.77 4.305 ;
        RECT 38.06 4.135 38.23 4.305 ;
        RECT 38.52 4.135 38.69 4.305 ;
        RECT 38.98 4.135 39.15 4.305 ;
        RECT 39.44 4.135 39.61 4.305 ;
        RECT 39.9 4.135 40.07 4.305 ;
        RECT 40.36 4.135 40.53 4.305 ;
        RECT 40.82 4.135 40.99 4.305 ;
        RECT 41.28 4.135 41.45 4.305 ;
        RECT 41.74 4.135 41.91 4.305 ;
        RECT 42.2 4.135 42.37 4.305 ;
        RECT 42.66 4.135 42.83 4.305 ;
        RECT 43.12 4.135 43.29 4.305 ;
        RECT 43.58 4.135 43.75 4.305 ;
        RECT 44.04 4.135 44.21 4.305 ;
        RECT 44.5 4.135 44.67 4.305 ;
        RECT 44.77 4.545 44.94 4.715 ;
        RECT 44.96 4.135 45.13 4.305 ;
        RECT 45.42 4.135 45.59 4.305 ;
        RECT 45.88 4.135 46.05 4.305 ;
        RECT 46.34 4.135 46.51 4.305 ;
        RECT 46.8 4.135 46.97 4.305 ;
        RECT 50.385 4.545 50.555 4.715 ;
        RECT 50.385 4.165 50.555 4.335 ;
        RECT 51.085 4.55 51.255 4.72 ;
        RECT 51.085 4.16 51.255 4.33 ;
        RECT 52.075 4.55 52.245 4.72 ;
        RECT 52.075 4.16 52.245 4.33 ;
        RECT 53.86 4.135 54.03 4.305 ;
        RECT 54.32 4.135 54.49 4.305 ;
        RECT 54.78 4.135 54.95 4.305 ;
        RECT 55.24 4.135 55.41 4.305 ;
        RECT 55.7 4.135 55.87 4.305 ;
        RECT 56.16 4.135 56.33 4.305 ;
        RECT 56.62 4.135 56.79 4.305 ;
        RECT 57.08 4.135 57.25 4.305 ;
        RECT 57.54 4.135 57.71 4.305 ;
        RECT 58 4.135 58.17 4.305 ;
        RECT 58.46 4.135 58.63 4.305 ;
        RECT 58.92 4.135 59.09 4.305 ;
        RECT 59.38 4.135 59.55 4.305 ;
        RECT 59.84 4.135 60.01 4.305 ;
        RECT 60.3 4.135 60.47 4.305 ;
        RECT 60.76 4.135 60.93 4.305 ;
        RECT 61.22 4.135 61.39 4.305 ;
        RECT 61.68 4.135 61.85 4.305 ;
        RECT 62.14 4.135 62.31 4.305 ;
        RECT 62.6 4.135 62.77 4.305 ;
        RECT 63.06 4.135 63.23 4.305 ;
        RECT 63.33 4.545 63.5 4.715 ;
        RECT 63.52 4.135 63.69 4.305 ;
        RECT 63.98 4.135 64.15 4.305 ;
        RECT 64.44 4.135 64.61 4.305 ;
        RECT 64.9 4.135 65.07 4.305 ;
        RECT 65.36 4.135 65.53 4.305 ;
        RECT 68.945 4.545 69.115 4.715 ;
        RECT 68.945 4.165 69.115 4.335 ;
        RECT 69.645 4.55 69.815 4.72 ;
        RECT 69.645 4.16 69.815 4.33 ;
        RECT 70.635 4.55 70.805 4.72 ;
        RECT 70.635 4.16 70.805 4.33 ;
        RECT 72.42 4.135 72.59 4.305 ;
        RECT 72.88 4.135 73.05 4.305 ;
        RECT 73.34 4.135 73.51 4.305 ;
        RECT 73.8 4.135 73.97 4.305 ;
        RECT 74.26 4.135 74.43 4.305 ;
        RECT 74.72 4.135 74.89 4.305 ;
        RECT 75.18 4.135 75.35 4.305 ;
        RECT 75.64 4.135 75.81 4.305 ;
        RECT 76.1 4.135 76.27 4.305 ;
        RECT 76.56 4.135 76.73 4.305 ;
        RECT 77.02 4.135 77.19 4.305 ;
        RECT 77.48 4.135 77.65 4.305 ;
        RECT 77.94 4.135 78.11 4.305 ;
        RECT 78.4 4.135 78.57 4.305 ;
        RECT 78.86 4.135 79.03 4.305 ;
        RECT 79.32 4.135 79.49 4.305 ;
        RECT 79.78 4.135 79.95 4.305 ;
        RECT 80.24 4.135 80.41 4.305 ;
        RECT 80.7 4.135 80.87 4.305 ;
        RECT 81.16 4.135 81.33 4.305 ;
        RECT 81.62 4.135 81.79 4.305 ;
        RECT 81.89 4.545 82.06 4.715 ;
        RECT 82.08 4.135 82.25 4.305 ;
        RECT 82.54 4.135 82.71 4.305 ;
        RECT 83 4.135 83.17 4.305 ;
        RECT 83.46 4.135 83.63 4.305 ;
        RECT 83.92 4.135 84.09 4.305 ;
        RECT 87.505 4.545 87.675 4.715 ;
        RECT 87.505 4.165 87.675 4.335 ;
        RECT 88.205 4.55 88.375 4.72 ;
        RECT 88.205 4.16 88.375 4.33 ;
        RECT 89.195 4.55 89.365 4.72 ;
        RECT 89.195 4.16 89.365 4.33 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 73.89 2.415 74.62 2.745 ;
        RECT 55.33 2.415 56.06 2.745 ;
        RECT 36.77 2.415 37.5 2.745 ;
        RECT 18.21 2.415 18.94 2.745 ;
        RECT -0.35 2.415 0.38 2.745 ;
      LAYER li1 ;
        RECT 89.91 0 90.09 0.305 ;
        RECT -5.505 0 90.09 0.3 ;
        RECT 89.115 0 89.285 0.93 ;
        RECT 88.125 0 88.295 0.93 ;
        RECT 71.35 0 87.96 0.305 ;
        RECT 85.385 0 85.555 0.935 ;
        RECT 72.275 0 84.32 1.585 ;
        RECT 83.325 0 83.495 2.085 ;
        RECT 82.365 0 82.535 2.085 ;
        RECT 81.405 0 81.575 2.085 ;
        RECT 80.885 0 81.055 2.085 ;
        RECT 80.605 0 80.8 1.595 ;
        RECT 79.925 0 80.095 2.085 ;
        RECT 78.925 0 79.095 2.085 ;
        RECT 77.965 0 78.135 2.085 ;
        RECT 76.93 0 77.125 1.595 ;
        RECT 76.485 0 76.655 2.085 ;
        RECT 74.565 0 74.825 1.595 ;
        RECT 74.565 0 74.735 2.085 ;
        RECT 73.085 0 73.255 2.085 ;
        RECT 70.555 0 70.725 0.93 ;
        RECT 69.565 0 69.735 0.93 ;
        RECT 52.79 0 69.4 0.305 ;
        RECT 66.825 0 66.995 0.935 ;
        RECT 53.715 0 65.76 1.585 ;
        RECT 64.765 0 64.935 2.085 ;
        RECT 63.805 0 63.975 2.085 ;
        RECT 62.845 0 63.015 2.085 ;
        RECT 62.325 0 62.495 2.085 ;
        RECT 62.045 0 62.24 1.595 ;
        RECT 61.365 0 61.535 2.085 ;
        RECT 60.365 0 60.535 2.085 ;
        RECT 59.405 0 59.575 2.085 ;
        RECT 58.37 0 58.565 1.595 ;
        RECT 57.925 0 58.095 2.085 ;
        RECT 56.005 0 56.265 1.595 ;
        RECT 56.005 0 56.175 2.085 ;
        RECT 54.525 0 54.695 2.085 ;
        RECT 51.995 0 52.165 0.93 ;
        RECT 51.005 0 51.175 0.93 ;
        RECT 34.23 0 50.84 0.305 ;
        RECT 48.265 0 48.435 0.935 ;
        RECT 35.155 0 47.2 1.585 ;
        RECT 46.205 0 46.375 2.085 ;
        RECT 45.245 0 45.415 2.085 ;
        RECT 44.285 0 44.455 2.085 ;
        RECT 43.765 0 43.935 2.085 ;
        RECT 43.485 0 43.68 1.595 ;
        RECT 42.805 0 42.975 2.085 ;
        RECT 41.805 0 41.975 2.085 ;
        RECT 40.845 0 41.015 2.085 ;
        RECT 39.81 0 40.005 1.595 ;
        RECT 39.365 0 39.535 2.085 ;
        RECT 37.445 0 37.705 1.595 ;
        RECT 37.445 0 37.615 2.085 ;
        RECT 35.965 0 36.135 2.085 ;
        RECT 33.435 0 33.605 0.93 ;
        RECT 32.445 0 32.615 0.93 ;
        RECT 15.67 0 32.28 0.305 ;
        RECT 29.705 0 29.875 0.935 ;
        RECT 16.595 0 28.64 1.585 ;
        RECT 27.645 0 27.815 2.085 ;
        RECT 26.685 0 26.855 2.085 ;
        RECT 25.725 0 25.895 2.085 ;
        RECT 25.205 0 25.375 2.085 ;
        RECT 24.925 0 25.12 1.595 ;
        RECT 24.245 0 24.415 2.085 ;
        RECT 23.245 0 23.415 2.085 ;
        RECT 22.285 0 22.455 2.085 ;
        RECT 21.25 0 21.445 1.595 ;
        RECT 20.805 0 20.975 2.085 ;
        RECT 18.885 0 19.145 1.595 ;
        RECT 18.885 0 19.055 2.085 ;
        RECT 17.405 0 17.575 2.085 ;
        RECT 14.875 0 15.045 0.93 ;
        RECT 13.885 0 14.055 0.93 ;
        RECT -5.505 0 13.72 0.305 ;
        RECT 11.145 0 11.315 0.935 ;
        RECT -1.965 0 10.08 1.585 ;
        RECT 9.085 0 9.255 2.085 ;
        RECT 8.125 0 8.295 2.085 ;
        RECT 7.165 0 7.335 2.085 ;
        RECT 6.645 0 6.815 2.085 ;
        RECT 6.365 0 6.56 1.595 ;
        RECT 5.685 0 5.855 2.085 ;
        RECT 4.685 0 4.855 2.085 ;
        RECT 3.725 0 3.895 2.085 ;
        RECT 2.69 0 2.885 1.595 ;
        RECT 2.245 0 2.415 2.085 ;
        RECT 0.325 0 0.585 1.595 ;
        RECT 0.325 0 0.495 2.085 ;
        RECT -1.155 0 -0.985 2.085 ;
        RECT -5.505 8.58 90.09 8.88 ;
        RECT 89.91 8.575 90.09 8.88 ;
        RECT 89.115 7.95 89.285 8.88 ;
        RECT 88.125 7.95 88.295 8.88 ;
        RECT 71.35 8.575 87.96 8.88 ;
        RECT 85.385 7.945 85.555 8.88 ;
        RECT 79.77 7.945 79.94 8.88 ;
        RECT 70.555 7.95 70.725 8.88 ;
        RECT 69.565 7.95 69.735 8.88 ;
        RECT 52.79 8.575 69.4 8.88 ;
        RECT 66.825 7.945 66.995 8.88 ;
        RECT 61.21 7.945 61.38 8.88 ;
        RECT 51.995 7.95 52.165 8.88 ;
        RECT 51.005 7.95 51.175 8.88 ;
        RECT 34.23 8.575 50.84 8.88 ;
        RECT 48.265 7.945 48.435 8.88 ;
        RECT 42.65 7.945 42.82 8.88 ;
        RECT 33.435 7.95 33.605 8.88 ;
        RECT 32.445 7.95 32.615 8.88 ;
        RECT 15.67 8.575 32.28 8.88 ;
        RECT 29.705 7.945 29.875 8.88 ;
        RECT 24.09 7.945 24.26 8.88 ;
        RECT 14.875 7.95 15.045 8.88 ;
        RECT 13.885 7.95 14.055 8.88 ;
        RECT -5.505 8.575 13.72 8.88 ;
        RECT 11.145 7.945 11.315 8.88 ;
        RECT 5.53 7.945 5.7 8.88 ;
        RECT -5.285 7.945 -5.115 8.88 ;
        RECT 80.775 6.075 80.945 8.025 ;
        RECT 80.72 7.855 80.89 8.305 ;
        RECT 80.72 5.015 80.89 6.245 ;
        RECT 75.765 2.495 75.935 2.825 ;
        RECT 73.925 3.055 74.215 3.225 ;
        RECT 73.925 2.575 74.095 3.225 ;
        RECT 73.725 2.575 74.095 2.745 ;
        RECT 62.215 6.075 62.385 8.025 ;
        RECT 62.16 7.855 62.33 8.305 ;
        RECT 62.16 5.015 62.33 6.245 ;
        RECT 57.205 2.495 57.375 2.825 ;
        RECT 55.365 3.055 55.655 3.225 ;
        RECT 55.365 2.575 55.535 3.225 ;
        RECT 55.165 2.575 55.535 2.745 ;
        RECT 43.655 6.075 43.825 8.025 ;
        RECT 43.6 7.855 43.77 8.305 ;
        RECT 43.6 5.015 43.77 6.245 ;
        RECT 38.645 2.495 38.815 2.825 ;
        RECT 36.805 3.055 37.095 3.225 ;
        RECT 36.805 2.575 36.975 3.225 ;
        RECT 36.605 2.575 36.975 2.745 ;
        RECT 25.095 6.075 25.265 8.025 ;
        RECT 25.04 7.855 25.21 8.305 ;
        RECT 25.04 5.015 25.21 6.245 ;
        RECT 20.085 2.495 20.255 2.825 ;
        RECT 18.245 3.055 18.535 3.225 ;
        RECT 18.245 2.575 18.415 3.225 ;
        RECT 18.045 2.575 18.415 2.745 ;
        RECT 6.535 6.075 6.705 8.025 ;
        RECT 6.48 7.855 6.65 8.305 ;
        RECT 6.48 5.015 6.65 6.245 ;
        RECT 1.525 2.495 1.695 2.825 ;
        RECT -0.315 3.055 -0.025 3.225 ;
        RECT -0.315 2.575 -0.145 3.225 ;
        RECT -0.515 2.575 -0.145 2.745 ;
      LAYER met2 ;
        RECT 75.72 2.42 75.98 2.74 ;
        RECT 73.94 2.51 75.98 2.65 ;
        RECT 74.32 1 74.66 1.34 ;
        RECT 74.25 2.395 74.53 2.765 ;
        RECT 74.345 1 74.515 2.765 ;
        RECT 74 2.98 74.26 3.3 ;
        RECT 73.94 2.51 74.08 3.21 ;
        RECT 57.16 2.42 57.42 2.74 ;
        RECT 55.38 2.51 57.42 2.65 ;
        RECT 55.76 1 56.1 1.34 ;
        RECT 55.69 2.395 55.97 2.765 ;
        RECT 55.785 1 55.955 2.765 ;
        RECT 55.44 2.98 55.7 3.3 ;
        RECT 55.38 2.51 55.52 3.21 ;
        RECT 38.6 2.42 38.86 2.74 ;
        RECT 36.82 2.51 38.86 2.65 ;
        RECT 37.2 1 37.54 1.34 ;
        RECT 37.13 2.395 37.41 2.765 ;
        RECT 37.225 1 37.395 2.765 ;
        RECT 36.88 2.98 37.14 3.3 ;
        RECT 36.82 2.51 36.96 3.21 ;
        RECT 20.04 2.42 20.3 2.74 ;
        RECT 18.26 2.51 20.3 2.65 ;
        RECT 18.64 1 18.98 1.34 ;
        RECT 18.57 2.395 18.85 2.765 ;
        RECT 18.665 1 18.835 2.765 ;
        RECT 18.32 2.98 18.58 3.3 ;
        RECT 18.26 2.51 18.4 3.21 ;
        RECT 1.48 2.42 1.74 2.74 ;
        RECT -0.3 2.51 1.74 2.65 ;
        RECT 0.08 1 0.42 1.34 ;
        RECT 0.01 2.395 0.29 2.765 ;
        RECT 0.105 1 0.275 2.765 ;
        RECT -0.24 2.98 0.02 3.3 ;
        RECT -0.3 2.51 -0.16 3.21 ;
      LAYER met1 ;
        RECT 89.91 0 90.09 0.305 ;
        RECT -5.505 0 90.09 0.3 ;
        RECT 71.35 0 87.96 0.305 ;
        RECT 72.275 0 84.32 1.585 ;
        RECT 72.275 0 84.235 1.74 ;
        RECT 52.79 0 69.4 0.305 ;
        RECT 53.715 0 65.76 1.585 ;
        RECT 53.715 0 65.675 1.74 ;
        RECT 34.23 0 50.84 0.305 ;
        RECT 35.155 0 47.2 1.585 ;
        RECT 35.155 0 47.115 1.74 ;
        RECT 15.67 0 32.28 0.305 ;
        RECT 16.595 0 28.64 1.585 ;
        RECT 16.595 0 28.555 1.74 ;
        RECT -5.505 0 13.72 0.305 ;
        RECT -1.965 0 10.08 1.585 ;
        RECT -1.965 0 9.995 1.74 ;
        RECT -5.505 8.58 90.09 8.88 ;
        RECT 89.91 8.575 90.09 8.88 ;
        RECT 71.35 8.575 87.96 8.88 ;
        RECT 80.715 6.285 81.005 6.515 ;
        RECT 80.28 6.315 81.005 6.485 ;
        RECT 80.28 6.315 80.45 8.88 ;
        RECT 52.79 8.575 69.4 8.88 ;
        RECT 62.155 6.285 62.445 6.515 ;
        RECT 61.72 6.315 62.445 6.485 ;
        RECT 61.72 6.315 61.89 8.88 ;
        RECT 34.23 8.575 50.84 8.88 ;
        RECT 43.595 6.285 43.885 6.515 ;
        RECT 43.16 6.315 43.885 6.485 ;
        RECT 43.16 6.315 43.33 8.88 ;
        RECT 15.67 8.575 32.28 8.88 ;
        RECT 25.035 6.285 25.325 6.515 ;
        RECT 24.6 6.315 25.325 6.485 ;
        RECT 24.6 6.315 24.77 8.88 ;
        RECT -5.505 8.575 13.72 8.88 ;
        RECT 6.475 6.285 6.765 6.515 ;
        RECT 6.04 6.315 6.765 6.485 ;
        RECT 6.04 6.315 6.21 8.88 ;
        RECT 75.705 2.37 75.995 2.74 ;
        RECT 74.94 2.37 75.995 2.51 ;
        RECT 73.97 3.01 74.29 3.27 ;
        RECT 57.145 2.37 57.435 2.74 ;
        RECT 56.38 2.37 57.435 2.51 ;
        RECT 55.41 3.01 55.73 3.27 ;
        RECT 38.585 2.37 38.875 2.74 ;
        RECT 37.82 2.37 38.875 2.51 ;
        RECT 36.85 3.01 37.17 3.27 ;
        RECT 20.025 2.37 20.315 2.74 ;
        RECT 19.26 2.37 20.315 2.51 ;
        RECT 18.29 3.01 18.61 3.27 ;
        RECT 1.465 2.37 1.755 2.74 ;
        RECT 0.7 2.37 1.755 2.51 ;
        RECT -0.27 3.01 0.05 3.27 ;
      LAYER via2 ;
        RECT 0.05 2.48 0.25 2.68 ;
        RECT 18.61 2.48 18.81 2.68 ;
        RECT 37.17 2.48 37.37 2.68 ;
        RECT 55.73 2.48 55.93 2.68 ;
        RECT 74.29 2.48 74.49 2.68 ;
      LAYER via1 ;
        RECT -0.185 3.065 -0.035 3.215 ;
        RECT 0.175 1.095 0.325 1.245 ;
        RECT 1.535 2.505 1.685 2.655 ;
        RECT 18.375 3.065 18.525 3.215 ;
        RECT 18.735 1.095 18.885 1.245 ;
        RECT 20.095 2.505 20.245 2.655 ;
        RECT 36.935 3.065 37.085 3.215 ;
        RECT 37.295 1.095 37.445 1.245 ;
        RECT 38.655 2.505 38.805 2.655 ;
        RECT 55.495 3.065 55.645 3.215 ;
        RECT 55.855 1.095 56.005 1.245 ;
        RECT 57.215 2.505 57.365 2.655 ;
        RECT 74.055 3.065 74.205 3.215 ;
        RECT 74.415 1.095 74.565 1.245 ;
        RECT 75.775 2.505 75.925 2.655 ;
      LAYER mcon ;
        RECT -5.205 8.605 -5.035 8.775 ;
        RECT -4.525 8.605 -4.355 8.775 ;
        RECT -3.845 8.605 -3.675 8.775 ;
        RECT -3.165 8.605 -2.995 8.775 ;
        RECT -1.82 1.415 -1.65 1.585 ;
        RECT -1.36 1.415 -1.19 1.585 ;
        RECT -0.9 1.415 -0.73 1.585 ;
        RECT -0.44 1.415 -0.27 1.585 ;
        RECT -0.195 3.055 -0.025 3.225 ;
        RECT 0.02 1.415 0.19 1.585 ;
        RECT 0.48 1.415 0.65 1.585 ;
        RECT 0.94 1.415 1.11 1.585 ;
        RECT 1.4 1.415 1.57 1.585 ;
        RECT 1.525 2.495 1.695 2.665 ;
        RECT 1.86 1.415 2.03 1.585 ;
        RECT 2.32 1.415 2.49 1.585 ;
        RECT 2.78 1.415 2.95 1.585 ;
        RECT 3.24 1.415 3.41 1.585 ;
        RECT 3.7 1.415 3.87 1.585 ;
        RECT 4.16 1.415 4.33 1.585 ;
        RECT 4.62 1.415 4.79 1.585 ;
        RECT 5.08 1.415 5.25 1.585 ;
        RECT 5.54 1.415 5.71 1.585 ;
        RECT 5.61 8.605 5.78 8.775 ;
        RECT 6 1.415 6.17 1.585 ;
        RECT 6.29 8.605 6.46 8.775 ;
        RECT 6.46 1.415 6.63 1.585 ;
        RECT 6.535 6.315 6.705 6.485 ;
        RECT 6.92 1.415 7.09 1.585 ;
        RECT 6.97 8.605 7.14 8.775 ;
        RECT 7.38 1.415 7.55 1.585 ;
        RECT 7.65 8.605 7.82 8.775 ;
        RECT 7.84 1.415 8.01 1.585 ;
        RECT 8.3 1.415 8.47 1.585 ;
        RECT 8.76 1.415 8.93 1.585 ;
        RECT 9.22 1.415 9.39 1.585 ;
        RECT 9.68 1.415 9.85 1.585 ;
        RECT 11.225 8.605 11.395 8.775 ;
        RECT 11.225 0.105 11.395 0.275 ;
        RECT 11.905 8.605 12.075 8.775 ;
        RECT 11.905 0.105 12.075 0.275 ;
        RECT 12.585 8.605 12.755 8.775 ;
        RECT 12.585 0.105 12.755 0.275 ;
        RECT 13.265 8.605 13.435 8.775 ;
        RECT 13.265 0.105 13.435 0.275 ;
        RECT 13.965 8.61 14.135 8.78 ;
        RECT 13.965 0.1 14.135 0.27 ;
        RECT 14.955 8.61 15.125 8.78 ;
        RECT 14.955 0.1 15.125 0.27 ;
        RECT 16.74 1.415 16.91 1.585 ;
        RECT 17.2 1.415 17.37 1.585 ;
        RECT 17.66 1.415 17.83 1.585 ;
        RECT 18.12 1.415 18.29 1.585 ;
        RECT 18.365 3.055 18.535 3.225 ;
        RECT 18.58 1.415 18.75 1.585 ;
        RECT 19.04 1.415 19.21 1.585 ;
        RECT 19.5 1.415 19.67 1.585 ;
        RECT 19.96 1.415 20.13 1.585 ;
        RECT 20.085 2.495 20.255 2.665 ;
        RECT 20.42 1.415 20.59 1.585 ;
        RECT 20.88 1.415 21.05 1.585 ;
        RECT 21.34 1.415 21.51 1.585 ;
        RECT 21.8 1.415 21.97 1.585 ;
        RECT 22.26 1.415 22.43 1.585 ;
        RECT 22.72 1.415 22.89 1.585 ;
        RECT 23.18 1.415 23.35 1.585 ;
        RECT 23.64 1.415 23.81 1.585 ;
        RECT 24.1 1.415 24.27 1.585 ;
        RECT 24.17 8.605 24.34 8.775 ;
        RECT 24.56 1.415 24.73 1.585 ;
        RECT 24.85 8.605 25.02 8.775 ;
        RECT 25.02 1.415 25.19 1.585 ;
        RECT 25.095 6.315 25.265 6.485 ;
        RECT 25.48 1.415 25.65 1.585 ;
        RECT 25.53 8.605 25.7 8.775 ;
        RECT 25.94 1.415 26.11 1.585 ;
        RECT 26.21 8.605 26.38 8.775 ;
        RECT 26.4 1.415 26.57 1.585 ;
        RECT 26.86 1.415 27.03 1.585 ;
        RECT 27.32 1.415 27.49 1.585 ;
        RECT 27.78 1.415 27.95 1.585 ;
        RECT 28.24 1.415 28.41 1.585 ;
        RECT 29.785 8.605 29.955 8.775 ;
        RECT 29.785 0.105 29.955 0.275 ;
        RECT 30.465 8.605 30.635 8.775 ;
        RECT 30.465 0.105 30.635 0.275 ;
        RECT 31.145 8.605 31.315 8.775 ;
        RECT 31.145 0.105 31.315 0.275 ;
        RECT 31.825 8.605 31.995 8.775 ;
        RECT 31.825 0.105 31.995 0.275 ;
        RECT 32.525 8.61 32.695 8.78 ;
        RECT 32.525 0.1 32.695 0.27 ;
        RECT 33.515 8.61 33.685 8.78 ;
        RECT 33.515 0.1 33.685 0.27 ;
        RECT 35.3 1.415 35.47 1.585 ;
        RECT 35.76 1.415 35.93 1.585 ;
        RECT 36.22 1.415 36.39 1.585 ;
        RECT 36.68 1.415 36.85 1.585 ;
        RECT 36.925 3.055 37.095 3.225 ;
        RECT 37.14 1.415 37.31 1.585 ;
        RECT 37.6 1.415 37.77 1.585 ;
        RECT 38.06 1.415 38.23 1.585 ;
        RECT 38.52 1.415 38.69 1.585 ;
        RECT 38.645 2.495 38.815 2.665 ;
        RECT 38.98 1.415 39.15 1.585 ;
        RECT 39.44 1.415 39.61 1.585 ;
        RECT 39.9 1.415 40.07 1.585 ;
        RECT 40.36 1.415 40.53 1.585 ;
        RECT 40.82 1.415 40.99 1.585 ;
        RECT 41.28 1.415 41.45 1.585 ;
        RECT 41.74 1.415 41.91 1.585 ;
        RECT 42.2 1.415 42.37 1.585 ;
        RECT 42.66 1.415 42.83 1.585 ;
        RECT 42.73 8.605 42.9 8.775 ;
        RECT 43.12 1.415 43.29 1.585 ;
        RECT 43.41 8.605 43.58 8.775 ;
        RECT 43.58 1.415 43.75 1.585 ;
        RECT 43.655 6.315 43.825 6.485 ;
        RECT 44.04 1.415 44.21 1.585 ;
        RECT 44.09 8.605 44.26 8.775 ;
        RECT 44.5 1.415 44.67 1.585 ;
        RECT 44.77 8.605 44.94 8.775 ;
        RECT 44.96 1.415 45.13 1.585 ;
        RECT 45.42 1.415 45.59 1.585 ;
        RECT 45.88 1.415 46.05 1.585 ;
        RECT 46.34 1.415 46.51 1.585 ;
        RECT 46.8 1.415 46.97 1.585 ;
        RECT 48.345 8.605 48.515 8.775 ;
        RECT 48.345 0.105 48.515 0.275 ;
        RECT 49.025 8.605 49.195 8.775 ;
        RECT 49.025 0.105 49.195 0.275 ;
        RECT 49.705 8.605 49.875 8.775 ;
        RECT 49.705 0.105 49.875 0.275 ;
        RECT 50.385 8.605 50.555 8.775 ;
        RECT 50.385 0.105 50.555 0.275 ;
        RECT 51.085 8.61 51.255 8.78 ;
        RECT 51.085 0.1 51.255 0.27 ;
        RECT 52.075 8.61 52.245 8.78 ;
        RECT 52.075 0.1 52.245 0.27 ;
        RECT 53.86 1.415 54.03 1.585 ;
        RECT 54.32 1.415 54.49 1.585 ;
        RECT 54.78 1.415 54.95 1.585 ;
        RECT 55.24 1.415 55.41 1.585 ;
        RECT 55.485 3.055 55.655 3.225 ;
        RECT 55.7 1.415 55.87 1.585 ;
        RECT 56.16 1.415 56.33 1.585 ;
        RECT 56.62 1.415 56.79 1.585 ;
        RECT 57.08 1.415 57.25 1.585 ;
        RECT 57.205 2.495 57.375 2.665 ;
        RECT 57.54 1.415 57.71 1.585 ;
        RECT 58 1.415 58.17 1.585 ;
        RECT 58.46 1.415 58.63 1.585 ;
        RECT 58.92 1.415 59.09 1.585 ;
        RECT 59.38 1.415 59.55 1.585 ;
        RECT 59.84 1.415 60.01 1.585 ;
        RECT 60.3 1.415 60.47 1.585 ;
        RECT 60.76 1.415 60.93 1.585 ;
        RECT 61.22 1.415 61.39 1.585 ;
        RECT 61.29 8.605 61.46 8.775 ;
        RECT 61.68 1.415 61.85 1.585 ;
        RECT 61.97 8.605 62.14 8.775 ;
        RECT 62.14 1.415 62.31 1.585 ;
        RECT 62.215 6.315 62.385 6.485 ;
        RECT 62.6 1.415 62.77 1.585 ;
        RECT 62.65 8.605 62.82 8.775 ;
        RECT 63.06 1.415 63.23 1.585 ;
        RECT 63.33 8.605 63.5 8.775 ;
        RECT 63.52 1.415 63.69 1.585 ;
        RECT 63.98 1.415 64.15 1.585 ;
        RECT 64.44 1.415 64.61 1.585 ;
        RECT 64.9 1.415 65.07 1.585 ;
        RECT 65.36 1.415 65.53 1.585 ;
        RECT 66.905 8.605 67.075 8.775 ;
        RECT 66.905 0.105 67.075 0.275 ;
        RECT 67.585 8.605 67.755 8.775 ;
        RECT 67.585 0.105 67.755 0.275 ;
        RECT 68.265 8.605 68.435 8.775 ;
        RECT 68.265 0.105 68.435 0.275 ;
        RECT 68.945 8.605 69.115 8.775 ;
        RECT 68.945 0.105 69.115 0.275 ;
        RECT 69.645 8.61 69.815 8.78 ;
        RECT 69.645 0.1 69.815 0.27 ;
        RECT 70.635 8.61 70.805 8.78 ;
        RECT 70.635 0.1 70.805 0.27 ;
        RECT 72.42 1.415 72.59 1.585 ;
        RECT 72.88 1.415 73.05 1.585 ;
        RECT 73.34 1.415 73.51 1.585 ;
        RECT 73.8 1.415 73.97 1.585 ;
        RECT 74.045 3.055 74.215 3.225 ;
        RECT 74.26 1.415 74.43 1.585 ;
        RECT 74.72 1.415 74.89 1.585 ;
        RECT 75.18 1.415 75.35 1.585 ;
        RECT 75.64 1.415 75.81 1.585 ;
        RECT 75.765 2.495 75.935 2.665 ;
        RECT 76.1 1.415 76.27 1.585 ;
        RECT 76.56 1.415 76.73 1.585 ;
        RECT 77.02 1.415 77.19 1.585 ;
        RECT 77.48 1.415 77.65 1.585 ;
        RECT 77.94 1.415 78.11 1.585 ;
        RECT 78.4 1.415 78.57 1.585 ;
        RECT 78.86 1.415 79.03 1.585 ;
        RECT 79.32 1.415 79.49 1.585 ;
        RECT 79.78 1.415 79.95 1.585 ;
        RECT 79.85 8.605 80.02 8.775 ;
        RECT 80.24 1.415 80.41 1.585 ;
        RECT 80.53 8.605 80.7 8.775 ;
        RECT 80.7 1.415 80.87 1.585 ;
        RECT 80.775 6.315 80.945 6.485 ;
        RECT 81.16 1.415 81.33 1.585 ;
        RECT 81.21 8.605 81.38 8.775 ;
        RECT 81.62 1.415 81.79 1.585 ;
        RECT 81.89 8.605 82.06 8.775 ;
        RECT 82.08 1.415 82.25 1.585 ;
        RECT 82.54 1.415 82.71 1.585 ;
        RECT 83 1.415 83.17 1.585 ;
        RECT 83.46 1.415 83.63 1.585 ;
        RECT 83.92 1.415 84.09 1.585 ;
        RECT 85.465 8.605 85.635 8.775 ;
        RECT 85.465 0.105 85.635 0.275 ;
        RECT 86.145 8.605 86.315 8.775 ;
        RECT 86.145 0.105 86.315 0.275 ;
        RECT 86.825 8.605 86.995 8.775 ;
        RECT 86.825 0.105 86.995 0.275 ;
        RECT 87.505 8.605 87.675 8.775 ;
        RECT 87.505 0.105 87.675 0.275 ;
        RECT 88.205 8.61 88.375 8.78 ;
        RECT 88.205 0.1 88.375 0.27 ;
        RECT 89.195 8.61 89.365 8.78 ;
        RECT 89.195 0.1 89.365 0.27 ;
    END
  END vssd1
  OBS
    LAYER met3 ;
      RECT 81.58 3.535 82.135 3.865 ;
      RECT 81.58 1.87 81.88 3.865 ;
      RECT 77.645 2.975 78.2 3.305 ;
      RECT 77.9 1.87 78.2 3.305 ;
      RECT 77.9 1.87 81.88 2.17 ;
      RECT 81.05 7.055 81.425 7.425 ;
      RECT 81.05 7.095 82.055 7.395 ;
      RECT 81.755 4.405 82.055 7.395 ;
      RECT 71.925 4.405 82.055 4.705 ;
      RECT 76.43 2.415 76.73 4.705 ;
      RECT 74.995 2.975 75.295 4.705 ;
      RECT 71.925 2.42 72.225 4.705 ;
      RECT 74.965 2.975 75.695 3.305 ;
      RECT 76.405 2.415 77.135 2.745 ;
      RECT 72.855 2.415 73.585 2.745 ;
      RECT 71.925 2.42 73.585 2.72 ;
      RECT 63.02 3.535 63.575 3.865 ;
      RECT 63.02 1.87 63.32 3.865 ;
      RECT 59.085 2.975 59.64 3.305 ;
      RECT 59.34 1.87 59.64 3.305 ;
      RECT 59.34 1.87 63.32 2.17 ;
      RECT 62.49 7.055 62.865 7.425 ;
      RECT 62.49 7.095 63.495 7.395 ;
      RECT 63.195 4.405 63.495 7.395 ;
      RECT 53.365 4.405 63.495 4.705 ;
      RECT 57.87 2.415 58.17 4.705 ;
      RECT 56.435 2.975 56.735 4.705 ;
      RECT 53.365 2.42 53.665 4.705 ;
      RECT 56.405 2.975 57.135 3.305 ;
      RECT 57.845 2.415 58.575 2.745 ;
      RECT 54.295 2.415 55.025 2.745 ;
      RECT 53.365 2.42 55.025 2.72 ;
      RECT 44.46 3.535 45.015 3.865 ;
      RECT 44.46 1.87 44.76 3.865 ;
      RECT 40.525 2.975 41.08 3.305 ;
      RECT 40.78 1.87 41.08 3.305 ;
      RECT 40.78 1.87 44.76 2.17 ;
      RECT 43.93 7.055 44.305 7.425 ;
      RECT 43.93 7.095 44.935 7.395 ;
      RECT 44.635 4.405 44.935 7.395 ;
      RECT 34.805 4.405 44.935 4.705 ;
      RECT 39.31 2.415 39.61 4.705 ;
      RECT 37.875 2.975 38.175 4.705 ;
      RECT 34.805 2.42 35.105 4.705 ;
      RECT 37.845 2.975 38.575 3.305 ;
      RECT 39.285 2.415 40.015 2.745 ;
      RECT 35.735 2.415 36.465 2.745 ;
      RECT 34.805 2.42 36.465 2.72 ;
      RECT 25.9 3.535 26.455 3.865 ;
      RECT 25.9 1.87 26.2 3.865 ;
      RECT 21.965 2.975 22.52 3.305 ;
      RECT 22.22 1.87 22.52 3.305 ;
      RECT 22.22 1.87 26.2 2.17 ;
      RECT 25.37 7.055 25.745 7.425 ;
      RECT 25.37 7.095 26.375 7.395 ;
      RECT 26.075 4.405 26.375 7.395 ;
      RECT 16.245 4.405 26.375 4.705 ;
      RECT 20.75 2.415 21.05 4.705 ;
      RECT 19.315 2.975 19.615 4.705 ;
      RECT 16.245 2.42 16.545 4.705 ;
      RECT 19.285 2.975 20.015 3.305 ;
      RECT 20.725 2.415 21.455 2.745 ;
      RECT 17.175 2.415 17.905 2.745 ;
      RECT 16.245 2.42 17.905 2.72 ;
      RECT 7.34 3.535 7.895 3.865 ;
      RECT 7.34 1.87 7.64 3.865 ;
      RECT 3.405 2.975 3.96 3.305 ;
      RECT 3.66 1.87 3.96 3.305 ;
      RECT 3.66 1.87 7.64 2.17 ;
      RECT 6.81 7.055 7.185 7.425 ;
      RECT 6.81 7.095 7.815 7.395 ;
      RECT 7.515 4.405 7.815 7.395 ;
      RECT -2.315 4.405 7.815 4.705 ;
      RECT 2.19 2.415 2.49 4.705 ;
      RECT 0.755 2.975 1.055 4.705 ;
      RECT -2.315 2.42 -2.015 4.705 ;
      RECT 0.725 2.975 1.455 3.305 ;
      RECT 2.165 2.415 2.895 2.745 ;
      RECT -1.385 2.415 -0.655 2.745 ;
      RECT -2.315 2.42 -0.655 2.72 ;
      RECT 82.765 1.855 83.495 2.185 ;
      RECT 80.545 3.535 81.275 3.865 ;
      RECT 78.845 3.535 79.575 3.865 ;
      RECT 72.525 3.535 73.255 3.865 ;
      RECT 64.205 1.855 64.935 2.185 ;
      RECT 61.985 3.535 62.715 3.865 ;
      RECT 60.285 3.535 61.015 3.865 ;
      RECT 53.965 3.535 54.695 3.865 ;
      RECT 45.645 1.855 46.375 2.185 ;
      RECT 43.425 3.535 44.155 3.865 ;
      RECT 41.725 3.535 42.455 3.865 ;
      RECT 35.405 3.535 36.135 3.865 ;
      RECT 27.085 1.855 27.815 2.185 ;
      RECT 24.865 3.535 25.595 3.865 ;
      RECT 23.165 3.535 23.895 3.865 ;
      RECT 16.845 3.535 17.575 3.865 ;
      RECT 8.525 1.855 9.255 2.185 ;
      RECT 6.305 3.535 7.035 3.865 ;
      RECT 4.605 3.535 5.335 3.865 ;
      RECT -1.715 3.535 -0.985 3.865 ;
    LAYER via2 ;
      RECT 82.83 1.92 83.03 2.12 ;
      RECT 81.87 3.6 82.07 3.8 ;
      RECT 81.135 7.14 81.335 7.34 ;
      RECT 80.87 3.6 81.07 3.8 ;
      RECT 78.91 3.6 79.11 3.8 ;
      RECT 77.71 3.04 77.91 3.24 ;
      RECT 76.47 2.48 76.67 2.68 ;
      RECT 75.03 3.04 75.23 3.24 ;
      RECT 73.07 2.48 73.27 2.68 ;
      RECT 72.59 3.6 72.79 3.8 ;
      RECT 64.27 1.92 64.47 2.12 ;
      RECT 63.31 3.6 63.51 3.8 ;
      RECT 62.575 7.14 62.775 7.34 ;
      RECT 62.31 3.6 62.51 3.8 ;
      RECT 60.35 3.6 60.55 3.8 ;
      RECT 59.15 3.04 59.35 3.24 ;
      RECT 57.91 2.48 58.11 2.68 ;
      RECT 56.47 3.04 56.67 3.24 ;
      RECT 54.51 2.48 54.71 2.68 ;
      RECT 54.03 3.6 54.23 3.8 ;
      RECT 45.71 1.92 45.91 2.12 ;
      RECT 44.75 3.6 44.95 3.8 ;
      RECT 44.015 7.14 44.215 7.34 ;
      RECT 43.75 3.6 43.95 3.8 ;
      RECT 41.79 3.6 41.99 3.8 ;
      RECT 40.59 3.04 40.79 3.24 ;
      RECT 39.35 2.48 39.55 2.68 ;
      RECT 37.91 3.04 38.11 3.24 ;
      RECT 35.95 2.48 36.15 2.68 ;
      RECT 35.47 3.6 35.67 3.8 ;
      RECT 27.15 1.92 27.35 2.12 ;
      RECT 26.19 3.6 26.39 3.8 ;
      RECT 25.455 7.14 25.655 7.34 ;
      RECT 25.19 3.6 25.39 3.8 ;
      RECT 23.23 3.6 23.43 3.8 ;
      RECT 22.03 3.04 22.23 3.24 ;
      RECT 20.79 2.48 20.99 2.68 ;
      RECT 19.35 3.04 19.55 3.24 ;
      RECT 17.39 2.48 17.59 2.68 ;
      RECT 16.91 3.6 17.11 3.8 ;
      RECT 8.59 1.92 8.79 2.12 ;
      RECT 7.63 3.6 7.83 3.8 ;
      RECT 6.895 7.14 7.095 7.34 ;
      RECT 6.63 3.6 6.83 3.8 ;
      RECT 4.67 3.6 4.87 3.8 ;
      RECT 3.47 3.04 3.67 3.24 ;
      RECT 2.23 2.48 2.43 2.68 ;
      RECT 0.79 3.04 0.99 3.24 ;
      RECT -1.17 2.48 -0.97 2.68 ;
      RECT -1.65 3.6 -1.45 3.8 ;
    LAYER met2 ;
      RECT -4.28 8.4 89.72 8.57 ;
      RECT 89.55 7.275 89.72 8.57 ;
      RECT -4.28 6.255 -4.11 8.57 ;
      RECT 89.52 7.275 89.87 7.625 ;
      RECT -4.34 6.255 -4.05 6.605 ;
      RECT 86.36 6.22 86.68 6.545 ;
      RECT 86.39 5.695 86.56 6.545 ;
      RECT 86.39 5.695 86.565 6.045 ;
      RECT 86.39 5.695 87.365 5.87 ;
      RECT 87.19 1.965 87.365 5.87 ;
      RECT 87.135 1.965 87.485 2.315 ;
      RECT 87.16 6.655 87.485 6.98 ;
      RECT 86.045 6.745 87.485 6.915 ;
      RECT 86.045 2.395 86.205 6.915 ;
      RECT 86.36 2.365 86.68 2.685 ;
      RECT 86.045 2.395 86.68 2.565 ;
      RECT 78.925 4.135 85.015 4.325 ;
      RECT 84.845 3.145 85.015 4.325 ;
      RECT 84.825 3.15 85.015 4.325 ;
      RECT 78.925 3.515 79.095 4.325 ;
      RECT 78.87 3.515 79.15 3.885 ;
      RECT 78.94 3.07 79.08 4.325 ;
      RECT 84.755 3.15 85.095 3.5 ;
      RECT 78.75 2.955 79.03 3.325 ;
      RECT 78.46 3.07 79.08 3.21 ;
      RECT 78.46 1.86 78.6 3.21 ;
      RECT 78.4 1.86 78.66 2.18 ;
      RECT 70.935 6.655 71.285 7.005 ;
      RECT 81.72 6.61 82.07 6.96 ;
      RECT 70.935 6.685 82.07 6.885 ;
      RECT 81.36 2.98 81.62 3.3 ;
      RECT 81.42 1.86 81.56 3.3 ;
      RECT 81.36 1.86 81.62 2.18 ;
      RECT 80.36 3.54 80.62 3.86 ;
      RECT 80.36 2.955 80.56 3.86 ;
      RECT 80.3 1.86 80.44 3.49 ;
      RECT 80.3 2.955 80.8 3.325 ;
      RECT 80.24 1.86 80.5 2.18 ;
      RECT 79.88 3.54 80.14 3.86 ;
      RECT 79.94 1.95 80.08 3.86 ;
      RECT 79.64 1.95 80.08 2.18 ;
      RECT 79.64 1.86 79.9 2.18 ;
      RECT 79.4 2.42 79.66 2.74 ;
      RECT 78.82 2.51 79.66 2.65 ;
      RECT 78.82 1.57 78.96 2.65 ;
      RECT 75.48 1.86 75.74 2.18 ;
      RECT 75.48 1.95 76.52 2.09 ;
      RECT 76.38 1.57 76.52 2.09 ;
      RECT 76.38 1.57 78.96 1.71 ;
      RECT 77.67 2.955 77.95 3.325 ;
      RECT 77.74 1.86 77.88 3.325 ;
      RECT 77.68 1.86 77.94 2.18 ;
      RECT 77.32 3.54 77.58 3.86 ;
      RECT 77.38 1.95 77.52 3.86 ;
      RECT 76.96 1.86 77.22 2.18 ;
      RECT 76.96 1.95 77.52 2.09 ;
      RECT 74.99 2.955 75.27 3.325 ;
      RECT 76.96 2.98 77.22 3.3 ;
      RECT 74.64 2.98 75.27 3.3 ;
      RECT 74.64 3.07 77.22 3.21 ;
      RECT 76.43 2.395 76.71 2.765 ;
      RECT 76.43 2.42 76.96 2.74 ;
      RECT 73.52 2.98 73.78 3.3 ;
      RECT 73.58 1.86 73.72 3.3 ;
      RECT 73.52 1.86 73.78 2.18 ;
      RECT 72.55 3.515 72.83 3.885 ;
      RECT 72.56 3.26 72.82 3.885 ;
      RECT 67.8 6.22 68.12 6.545 ;
      RECT 67.83 5.695 68 6.545 ;
      RECT 67.83 5.695 68.005 6.045 ;
      RECT 67.83 5.695 68.805 5.87 ;
      RECT 68.63 1.965 68.805 5.87 ;
      RECT 68.575 1.965 68.925 2.315 ;
      RECT 68.6 6.655 68.925 6.98 ;
      RECT 67.485 6.745 68.925 6.915 ;
      RECT 67.485 2.395 67.645 6.915 ;
      RECT 67.8 2.365 68.12 2.685 ;
      RECT 67.485 2.395 68.12 2.565 ;
      RECT 60.365 4.135 66.455 4.325 ;
      RECT 66.285 3.145 66.455 4.325 ;
      RECT 66.265 3.15 66.455 4.325 ;
      RECT 60.365 3.515 60.535 4.325 ;
      RECT 60.31 3.515 60.59 3.885 ;
      RECT 60.38 3.07 60.52 4.325 ;
      RECT 66.195 3.15 66.535 3.5 ;
      RECT 60.19 2.955 60.47 3.325 ;
      RECT 59.9 3.07 60.52 3.21 ;
      RECT 59.9 1.86 60.04 3.21 ;
      RECT 59.84 1.86 60.1 2.18 ;
      RECT 52.375 6.655 52.725 7.005 ;
      RECT 63.16 6.61 63.51 6.96 ;
      RECT 52.375 6.685 63.51 6.885 ;
      RECT 62.8 2.98 63.06 3.3 ;
      RECT 62.86 1.86 63 3.3 ;
      RECT 62.8 1.86 63.06 2.18 ;
      RECT 61.8 3.54 62.06 3.86 ;
      RECT 61.8 2.955 62 3.86 ;
      RECT 61.74 1.86 61.88 3.49 ;
      RECT 61.74 2.955 62.24 3.325 ;
      RECT 61.68 1.86 61.94 2.18 ;
      RECT 61.32 3.54 61.58 3.86 ;
      RECT 61.38 1.95 61.52 3.86 ;
      RECT 61.08 1.95 61.52 2.18 ;
      RECT 61.08 1.86 61.34 2.18 ;
      RECT 60.84 2.42 61.1 2.74 ;
      RECT 60.26 2.51 61.1 2.65 ;
      RECT 60.26 1.57 60.4 2.65 ;
      RECT 56.92 1.86 57.18 2.18 ;
      RECT 56.92 1.95 57.96 2.09 ;
      RECT 57.82 1.57 57.96 2.09 ;
      RECT 57.82 1.57 60.4 1.71 ;
      RECT 59.11 2.955 59.39 3.325 ;
      RECT 59.18 1.86 59.32 3.325 ;
      RECT 59.12 1.86 59.38 2.18 ;
      RECT 58.76 3.54 59.02 3.86 ;
      RECT 58.82 1.95 58.96 3.86 ;
      RECT 58.4 1.86 58.66 2.18 ;
      RECT 58.4 1.95 58.96 2.09 ;
      RECT 56.43 2.955 56.71 3.325 ;
      RECT 58.4 2.98 58.66 3.3 ;
      RECT 56.08 2.98 56.71 3.3 ;
      RECT 56.08 3.07 58.66 3.21 ;
      RECT 57.87 2.395 58.15 2.765 ;
      RECT 57.87 2.42 58.4 2.74 ;
      RECT 54.96 2.98 55.22 3.3 ;
      RECT 55.02 1.86 55.16 3.3 ;
      RECT 54.96 1.86 55.22 2.18 ;
      RECT 53.99 3.515 54.27 3.885 ;
      RECT 54 3.26 54.26 3.885 ;
      RECT 49.24 6.22 49.56 6.545 ;
      RECT 49.27 5.695 49.44 6.545 ;
      RECT 49.27 5.695 49.445 6.045 ;
      RECT 49.27 5.695 50.245 5.87 ;
      RECT 50.07 1.965 50.245 5.87 ;
      RECT 50.015 1.965 50.365 2.315 ;
      RECT 50.04 6.655 50.365 6.98 ;
      RECT 48.925 6.745 50.365 6.915 ;
      RECT 48.925 2.395 49.085 6.915 ;
      RECT 49.24 2.365 49.56 2.685 ;
      RECT 48.925 2.395 49.56 2.565 ;
      RECT 41.805 4.135 47.895 4.325 ;
      RECT 47.725 3.145 47.895 4.325 ;
      RECT 47.705 3.15 47.895 4.325 ;
      RECT 41.805 3.515 41.975 4.325 ;
      RECT 41.75 3.515 42.03 3.885 ;
      RECT 41.82 3.07 41.96 4.325 ;
      RECT 47.635 3.15 47.975 3.5 ;
      RECT 41.63 2.955 41.91 3.325 ;
      RECT 41.34 3.07 41.96 3.21 ;
      RECT 41.34 1.86 41.48 3.21 ;
      RECT 41.28 1.86 41.54 2.18 ;
      RECT 33.86 6.66 34.21 7.01 ;
      RECT 44.6 6.615 44.95 6.965 ;
      RECT 33.86 6.69 44.95 6.89 ;
      RECT 44.24 2.98 44.5 3.3 ;
      RECT 44.3 1.86 44.44 3.3 ;
      RECT 44.24 1.86 44.5 2.18 ;
      RECT 43.24 3.54 43.5 3.86 ;
      RECT 43.24 2.955 43.44 3.86 ;
      RECT 43.18 1.86 43.32 3.49 ;
      RECT 43.18 2.955 43.68 3.325 ;
      RECT 43.12 1.86 43.38 2.18 ;
      RECT 42.76 3.54 43.02 3.86 ;
      RECT 42.82 1.95 42.96 3.86 ;
      RECT 42.52 1.95 42.96 2.18 ;
      RECT 42.52 1.86 42.78 2.18 ;
      RECT 42.28 2.42 42.54 2.74 ;
      RECT 41.7 2.51 42.54 2.65 ;
      RECT 41.7 1.57 41.84 2.65 ;
      RECT 38.36 1.86 38.62 2.18 ;
      RECT 38.36 1.95 39.4 2.09 ;
      RECT 39.26 1.57 39.4 2.09 ;
      RECT 39.26 1.57 41.84 1.71 ;
      RECT 40.55 2.955 40.83 3.325 ;
      RECT 40.62 1.86 40.76 3.325 ;
      RECT 40.56 1.86 40.82 2.18 ;
      RECT 40.2 3.54 40.46 3.86 ;
      RECT 40.26 1.95 40.4 3.86 ;
      RECT 39.84 1.86 40.1 2.18 ;
      RECT 39.84 1.95 40.4 2.09 ;
      RECT 37.87 2.955 38.15 3.325 ;
      RECT 39.84 2.98 40.1 3.3 ;
      RECT 37.52 2.98 38.15 3.3 ;
      RECT 37.52 3.07 40.1 3.21 ;
      RECT 39.31 2.395 39.59 2.765 ;
      RECT 39.31 2.42 39.84 2.74 ;
      RECT 36.4 2.98 36.66 3.3 ;
      RECT 36.46 1.86 36.6 3.3 ;
      RECT 36.4 1.86 36.66 2.18 ;
      RECT 35.43 3.515 35.71 3.885 ;
      RECT 35.44 3.26 35.7 3.885 ;
      RECT 30.68 6.22 31 6.545 ;
      RECT 30.71 5.695 30.88 6.545 ;
      RECT 30.71 5.695 30.885 6.045 ;
      RECT 30.71 5.695 31.685 5.87 ;
      RECT 31.51 1.965 31.685 5.87 ;
      RECT 31.455 1.965 31.805 2.315 ;
      RECT 31.48 6.655 31.805 6.98 ;
      RECT 30.365 6.745 31.805 6.915 ;
      RECT 30.365 2.395 30.525 6.915 ;
      RECT 30.68 2.365 31 2.685 ;
      RECT 30.365 2.395 31 2.565 ;
      RECT 23.245 4.135 29.335 4.325 ;
      RECT 29.165 3.145 29.335 4.325 ;
      RECT 29.145 3.15 29.335 4.325 ;
      RECT 23.245 3.515 23.415 4.325 ;
      RECT 23.19 3.515 23.47 3.885 ;
      RECT 23.26 3.07 23.4 4.325 ;
      RECT 29.075 3.15 29.415 3.5 ;
      RECT 23.07 2.955 23.35 3.325 ;
      RECT 22.78 3.07 23.4 3.21 ;
      RECT 22.78 1.86 22.92 3.21 ;
      RECT 22.72 1.86 22.98 2.18 ;
      RECT 15.3 6.655 15.65 7.005 ;
      RECT 26.045 6.61 26.395 6.96 ;
      RECT 15.3 6.685 26.395 6.885 ;
      RECT 25.68 2.98 25.94 3.3 ;
      RECT 25.74 1.86 25.88 3.3 ;
      RECT 25.68 1.86 25.94 2.18 ;
      RECT 24.68 3.54 24.94 3.86 ;
      RECT 24.68 2.955 24.88 3.86 ;
      RECT 24.62 1.86 24.76 3.49 ;
      RECT 24.62 2.955 25.12 3.325 ;
      RECT 24.56 1.86 24.82 2.18 ;
      RECT 24.2 3.54 24.46 3.86 ;
      RECT 24.26 1.95 24.4 3.86 ;
      RECT 23.96 1.95 24.4 2.18 ;
      RECT 23.96 1.86 24.22 2.18 ;
      RECT 23.72 2.42 23.98 2.74 ;
      RECT 23.14 2.51 23.98 2.65 ;
      RECT 23.14 1.57 23.28 2.65 ;
      RECT 19.8 1.86 20.06 2.18 ;
      RECT 19.8 1.95 20.84 2.09 ;
      RECT 20.7 1.57 20.84 2.09 ;
      RECT 20.7 1.57 23.28 1.71 ;
      RECT 21.99 2.955 22.27 3.325 ;
      RECT 22.06 1.86 22.2 3.325 ;
      RECT 22 1.86 22.26 2.18 ;
      RECT 21.64 3.54 21.9 3.86 ;
      RECT 21.7 1.95 21.84 3.86 ;
      RECT 21.28 1.86 21.54 2.18 ;
      RECT 21.28 1.95 21.84 2.09 ;
      RECT 19.31 2.955 19.59 3.325 ;
      RECT 21.28 2.98 21.54 3.3 ;
      RECT 18.96 2.98 19.59 3.3 ;
      RECT 18.96 3.07 21.54 3.21 ;
      RECT 20.75 2.395 21.03 2.765 ;
      RECT 20.75 2.42 21.28 2.74 ;
      RECT 17.84 2.98 18.1 3.3 ;
      RECT 17.9 1.86 18.04 3.3 ;
      RECT 17.84 1.86 18.1 2.18 ;
      RECT 16.87 3.515 17.15 3.885 ;
      RECT 16.88 3.26 17.14 3.885 ;
      RECT 12.12 6.22 12.44 6.545 ;
      RECT 12.15 5.695 12.32 6.545 ;
      RECT 12.15 5.695 12.325 6.045 ;
      RECT 12.15 5.695 13.125 5.87 ;
      RECT 12.95 1.965 13.125 5.87 ;
      RECT 12.895 1.965 13.245 2.315 ;
      RECT 12.92 6.655 13.245 6.98 ;
      RECT 11.805 6.745 13.245 6.915 ;
      RECT 11.805 2.395 11.965 6.915 ;
      RECT 12.12 2.365 12.44 2.685 ;
      RECT 11.805 2.395 12.44 2.565 ;
      RECT 4.685 4.135 10.775 4.325 ;
      RECT 10.605 3.145 10.775 4.325 ;
      RECT 10.585 3.15 10.775 4.325 ;
      RECT 4.685 3.515 4.855 4.325 ;
      RECT 4.63 3.515 4.91 3.885 ;
      RECT 4.7 3.07 4.84 4.325 ;
      RECT 10.515 3.15 10.855 3.5 ;
      RECT 4.51 2.955 4.79 3.325 ;
      RECT 4.22 3.07 4.84 3.21 ;
      RECT 4.22 1.86 4.36 3.21 ;
      RECT 4.16 1.86 4.42 2.18 ;
      RECT -3.965 6.995 -3.675 7.345 ;
      RECT -3.965 7.055 -2.775 7.225 ;
      RECT -2.945 6.685 -2.775 7.225 ;
      RECT 7.485 6.605 7.835 6.955 ;
      RECT -2.945 6.685 7.835 6.855 ;
      RECT 7.12 2.98 7.38 3.3 ;
      RECT 7.18 1.86 7.32 3.3 ;
      RECT 7.12 1.86 7.38 2.18 ;
      RECT 6.12 3.54 6.38 3.86 ;
      RECT 6.12 2.955 6.32 3.86 ;
      RECT 6.06 1.86 6.2 3.49 ;
      RECT 6.06 2.955 6.56 3.325 ;
      RECT 6 1.86 6.26 2.18 ;
      RECT 5.64 3.54 5.9 3.86 ;
      RECT 5.7 1.95 5.84 3.86 ;
      RECT 5.4 1.95 5.84 2.18 ;
      RECT 5.4 1.86 5.66 2.18 ;
      RECT 5.16 2.42 5.42 2.74 ;
      RECT 4.58 2.51 5.42 2.65 ;
      RECT 4.58 1.57 4.72 2.65 ;
      RECT 1.24 1.86 1.5 2.18 ;
      RECT 1.24 1.95 2.28 2.09 ;
      RECT 2.14 1.57 2.28 2.09 ;
      RECT 2.14 1.57 4.72 1.71 ;
      RECT 3.43 2.955 3.71 3.325 ;
      RECT 3.5 1.86 3.64 3.325 ;
      RECT 3.44 1.86 3.7 2.18 ;
      RECT 3.08 3.54 3.34 3.86 ;
      RECT 3.14 1.95 3.28 3.86 ;
      RECT 2.72 1.86 2.98 2.18 ;
      RECT 2.72 1.95 3.28 2.09 ;
      RECT 0.75 2.955 1.03 3.325 ;
      RECT 2.72 2.98 2.98 3.3 ;
      RECT 0.4 2.98 1.03 3.3 ;
      RECT 0.4 3.07 2.98 3.21 ;
      RECT 2.19 2.395 2.47 2.765 ;
      RECT 2.19 2.42 2.72 2.74 ;
      RECT -0.72 2.98 -0.46 3.3 ;
      RECT -0.66 1.86 -0.52 3.3 ;
      RECT -0.72 1.86 -0.46 2.18 ;
      RECT -1.69 3.515 -1.41 3.885 ;
      RECT -1.68 3.26 -1.42 3.885 ;
      RECT 82.79 1.835 83.07 2.205 ;
      RECT 81.83 3.515 82.11 3.885 ;
      RECT 81.05 7.055 81.425 7.425 ;
      RECT 80.83 3.515 81.11 3.885 ;
      RECT 73.03 2.395 73.31 2.765 ;
      RECT 64.23 1.835 64.51 2.205 ;
      RECT 63.27 3.515 63.55 3.885 ;
      RECT 62.49 7.055 62.865 7.425 ;
      RECT 62.27 3.515 62.55 3.885 ;
      RECT 54.47 2.395 54.75 2.765 ;
      RECT 45.67 1.835 45.95 2.205 ;
      RECT 44.71 3.515 44.99 3.885 ;
      RECT 43.93 7.055 44.305 7.425 ;
      RECT 43.71 3.515 43.99 3.885 ;
      RECT 35.91 2.395 36.19 2.765 ;
      RECT 27.11 1.835 27.39 2.205 ;
      RECT 26.15 3.515 26.43 3.885 ;
      RECT 25.37 7.055 25.745 7.425 ;
      RECT 25.15 3.515 25.43 3.885 ;
      RECT 17.35 2.395 17.63 2.765 ;
      RECT 8.55 1.835 8.83 2.205 ;
      RECT 7.59 3.515 7.87 3.885 ;
      RECT 6.81 7.055 7.185 7.425 ;
      RECT 6.59 3.515 6.87 3.885 ;
      RECT -1.21 2.395 -0.93 2.765 ;
    LAYER via1 ;
      RECT 89.62 7.375 89.77 7.525 ;
      RECT 87.25 6.74 87.4 6.89 ;
      RECT 87.235 2.065 87.385 2.215 ;
      RECT 86.445 2.45 86.595 2.6 ;
      RECT 86.445 6.325 86.595 6.475 ;
      RECT 84.855 3.25 85.005 3.4 ;
      RECT 82.855 1.945 83.005 2.095 ;
      RECT 81.895 3.625 82.045 3.775 ;
      RECT 81.82 6.71 81.97 6.86 ;
      RECT 81.415 1.945 81.565 2.095 ;
      RECT 81.415 3.065 81.565 3.215 ;
      RECT 81.16 7.165 81.31 7.315 ;
      RECT 80.895 3.625 81.045 3.775 ;
      RECT 80.415 3.625 80.565 3.775 ;
      RECT 80.295 1.945 80.445 2.095 ;
      RECT 79.935 3.625 80.085 3.775 ;
      RECT 79.695 1.945 79.845 2.095 ;
      RECT 79.455 2.505 79.605 2.655 ;
      RECT 78.935 3.625 79.085 3.775 ;
      RECT 78.455 1.945 78.605 2.095 ;
      RECT 77.735 1.945 77.885 2.095 ;
      RECT 77.735 3.065 77.885 3.215 ;
      RECT 77.375 3.625 77.525 3.775 ;
      RECT 77.015 1.945 77.165 2.095 ;
      RECT 77.015 3.065 77.165 3.215 ;
      RECT 76.755 2.505 76.905 2.655 ;
      RECT 75.535 1.945 75.685 2.095 ;
      RECT 74.695 3.065 74.845 3.215 ;
      RECT 73.575 1.945 73.725 2.095 ;
      RECT 73.575 3.065 73.725 3.215 ;
      RECT 73.095 2.505 73.245 2.655 ;
      RECT 72.615 3.345 72.765 3.495 ;
      RECT 71.035 6.755 71.185 6.905 ;
      RECT 68.69 6.74 68.84 6.89 ;
      RECT 68.675 2.065 68.825 2.215 ;
      RECT 67.885 2.45 68.035 2.6 ;
      RECT 67.885 6.325 68.035 6.475 ;
      RECT 66.295 3.25 66.445 3.4 ;
      RECT 64.295 1.945 64.445 2.095 ;
      RECT 63.335 3.625 63.485 3.775 ;
      RECT 63.26 6.71 63.41 6.86 ;
      RECT 62.855 1.945 63.005 2.095 ;
      RECT 62.855 3.065 63.005 3.215 ;
      RECT 62.6 7.165 62.75 7.315 ;
      RECT 62.335 3.625 62.485 3.775 ;
      RECT 61.855 3.625 62.005 3.775 ;
      RECT 61.735 1.945 61.885 2.095 ;
      RECT 61.375 3.625 61.525 3.775 ;
      RECT 61.135 1.945 61.285 2.095 ;
      RECT 60.895 2.505 61.045 2.655 ;
      RECT 60.375 3.625 60.525 3.775 ;
      RECT 59.895 1.945 60.045 2.095 ;
      RECT 59.175 1.945 59.325 2.095 ;
      RECT 59.175 3.065 59.325 3.215 ;
      RECT 58.815 3.625 58.965 3.775 ;
      RECT 58.455 1.945 58.605 2.095 ;
      RECT 58.455 3.065 58.605 3.215 ;
      RECT 58.195 2.505 58.345 2.655 ;
      RECT 56.975 1.945 57.125 2.095 ;
      RECT 56.135 3.065 56.285 3.215 ;
      RECT 55.015 1.945 55.165 2.095 ;
      RECT 55.015 3.065 55.165 3.215 ;
      RECT 54.535 2.505 54.685 2.655 ;
      RECT 54.055 3.345 54.205 3.495 ;
      RECT 52.475 6.755 52.625 6.905 ;
      RECT 50.13 6.74 50.28 6.89 ;
      RECT 50.115 2.065 50.265 2.215 ;
      RECT 49.325 2.45 49.475 2.6 ;
      RECT 49.325 6.325 49.475 6.475 ;
      RECT 47.735 3.25 47.885 3.4 ;
      RECT 45.735 1.945 45.885 2.095 ;
      RECT 44.775 3.625 44.925 3.775 ;
      RECT 44.7 6.715 44.85 6.865 ;
      RECT 44.295 1.945 44.445 2.095 ;
      RECT 44.295 3.065 44.445 3.215 ;
      RECT 44.04 7.165 44.19 7.315 ;
      RECT 43.775 3.625 43.925 3.775 ;
      RECT 43.295 3.625 43.445 3.775 ;
      RECT 43.175 1.945 43.325 2.095 ;
      RECT 42.815 3.625 42.965 3.775 ;
      RECT 42.575 1.945 42.725 2.095 ;
      RECT 42.335 2.505 42.485 2.655 ;
      RECT 41.815 3.625 41.965 3.775 ;
      RECT 41.335 1.945 41.485 2.095 ;
      RECT 40.615 1.945 40.765 2.095 ;
      RECT 40.615 3.065 40.765 3.215 ;
      RECT 40.255 3.625 40.405 3.775 ;
      RECT 39.895 1.945 40.045 2.095 ;
      RECT 39.895 3.065 40.045 3.215 ;
      RECT 39.635 2.505 39.785 2.655 ;
      RECT 38.415 1.945 38.565 2.095 ;
      RECT 37.575 3.065 37.725 3.215 ;
      RECT 36.455 1.945 36.605 2.095 ;
      RECT 36.455 3.065 36.605 3.215 ;
      RECT 35.975 2.505 36.125 2.655 ;
      RECT 35.495 3.345 35.645 3.495 ;
      RECT 33.96 6.76 34.11 6.91 ;
      RECT 31.57 6.74 31.72 6.89 ;
      RECT 31.555 2.065 31.705 2.215 ;
      RECT 30.765 2.45 30.915 2.6 ;
      RECT 30.765 6.325 30.915 6.475 ;
      RECT 29.175 3.25 29.325 3.4 ;
      RECT 27.175 1.945 27.325 2.095 ;
      RECT 26.215 3.625 26.365 3.775 ;
      RECT 26.145 6.71 26.295 6.86 ;
      RECT 25.735 1.945 25.885 2.095 ;
      RECT 25.735 3.065 25.885 3.215 ;
      RECT 25.48 7.165 25.63 7.315 ;
      RECT 25.215 3.625 25.365 3.775 ;
      RECT 24.735 3.625 24.885 3.775 ;
      RECT 24.615 1.945 24.765 2.095 ;
      RECT 24.255 3.625 24.405 3.775 ;
      RECT 24.015 1.945 24.165 2.095 ;
      RECT 23.775 2.505 23.925 2.655 ;
      RECT 23.255 3.625 23.405 3.775 ;
      RECT 22.775 1.945 22.925 2.095 ;
      RECT 22.055 1.945 22.205 2.095 ;
      RECT 22.055 3.065 22.205 3.215 ;
      RECT 21.695 3.625 21.845 3.775 ;
      RECT 21.335 1.945 21.485 2.095 ;
      RECT 21.335 3.065 21.485 3.215 ;
      RECT 21.075 2.505 21.225 2.655 ;
      RECT 19.855 1.945 20.005 2.095 ;
      RECT 19.015 3.065 19.165 3.215 ;
      RECT 17.895 1.945 18.045 2.095 ;
      RECT 17.895 3.065 18.045 3.215 ;
      RECT 17.415 2.505 17.565 2.655 ;
      RECT 16.935 3.345 17.085 3.495 ;
      RECT 15.4 6.755 15.55 6.905 ;
      RECT 13.01 6.74 13.16 6.89 ;
      RECT 12.995 2.065 13.145 2.215 ;
      RECT 12.205 2.45 12.355 2.6 ;
      RECT 12.205 6.325 12.355 6.475 ;
      RECT 10.615 3.25 10.765 3.4 ;
      RECT 8.615 1.945 8.765 2.095 ;
      RECT 7.655 3.625 7.805 3.775 ;
      RECT 7.585 6.705 7.735 6.855 ;
      RECT 7.175 1.945 7.325 2.095 ;
      RECT 7.175 3.065 7.325 3.215 ;
      RECT 6.92 7.165 7.07 7.315 ;
      RECT 6.655 3.625 6.805 3.775 ;
      RECT 6.175 3.625 6.325 3.775 ;
      RECT 6.055 1.945 6.205 2.095 ;
      RECT 5.695 3.625 5.845 3.775 ;
      RECT 5.455 1.945 5.605 2.095 ;
      RECT 5.215 2.505 5.365 2.655 ;
      RECT 4.695 3.625 4.845 3.775 ;
      RECT 4.215 1.945 4.365 2.095 ;
      RECT 3.495 1.945 3.645 2.095 ;
      RECT 3.495 3.065 3.645 3.215 ;
      RECT 3.135 3.625 3.285 3.775 ;
      RECT 2.775 1.945 2.925 2.095 ;
      RECT 2.775 3.065 2.925 3.215 ;
      RECT 2.515 2.505 2.665 2.655 ;
      RECT 1.295 1.945 1.445 2.095 ;
      RECT 0.455 3.065 0.605 3.215 ;
      RECT -0.665 1.945 -0.515 2.095 ;
      RECT -0.665 3.065 -0.515 3.215 ;
      RECT -1.145 2.505 -0.995 2.655 ;
      RECT -1.625 3.345 -1.475 3.495 ;
      RECT -3.895 7.095 -3.745 7.245 ;
      RECT -4.27 6.355 -4.12 6.505 ;
    LAYER met1 ;
      RECT 89.485 7.77 89.775 8 ;
      RECT 89.545 6.29 89.715 8 ;
      RECT 89.52 7.275 89.87 7.625 ;
      RECT 89.485 6.29 89.775 6.52 ;
      RECT 89.08 2.395 89.185 2.965 ;
      RECT 89.08 2.73 89.405 2.96 ;
      RECT 89.08 2.76 89.575 2.93 ;
      RECT 89.08 2.395 89.27 2.96 ;
      RECT 88.495 2.36 88.785 2.59 ;
      RECT 88.495 2.395 89.27 2.565 ;
      RECT 88.555 0.88 88.725 2.59 ;
      RECT 88.495 0.88 88.785 1.11 ;
      RECT 88.495 7.77 88.785 8 ;
      RECT 88.555 6.29 88.725 8 ;
      RECT 88.495 6.29 88.785 6.52 ;
      RECT 88.495 6.325 89.35 6.485 ;
      RECT 89.18 5.92 89.35 6.485 ;
      RECT 88.495 6.32 88.89 6.485 ;
      RECT 89.115 5.92 89.405 6.15 ;
      RECT 89.115 5.95 89.575 6.12 ;
      RECT 88.125 2.73 88.415 2.96 ;
      RECT 88.125 2.76 88.585 2.93 ;
      RECT 88.19 1.655 88.355 2.96 ;
      RECT 86.705 1.625 86.995 1.855 ;
      RECT 86.705 1.655 88.355 1.825 ;
      RECT 86.765 0.885 86.935 1.855 ;
      RECT 86.705 0.885 86.995 1.115 ;
      RECT 86.705 7.765 86.995 7.995 ;
      RECT 86.765 7.025 86.935 7.995 ;
      RECT 86.765 7.12 88.355 7.29 ;
      RECT 88.185 5.92 88.355 7.29 ;
      RECT 86.705 7.025 86.995 7.255 ;
      RECT 88.125 5.92 88.415 6.15 ;
      RECT 88.125 5.95 88.585 6.12 ;
      RECT 84.755 3.15 85.095 3.5 ;
      RECT 84.845 2.025 85.015 3.5 ;
      RECT 87.135 1.965 87.485 2.315 ;
      RECT 84.845 2.025 87.485 2.195 ;
      RECT 87.16 6.655 87.485 6.98 ;
      RECT 81.72 6.61 82.07 6.96 ;
      RECT 87.135 6.655 87.485 6.885 ;
      RECT 81.52 6.655 82.07 6.885 ;
      RECT 81.35 6.685 87.485 6.855 ;
      RECT 86.36 2.365 86.68 2.685 ;
      RECT 86.33 2.365 86.68 2.595 ;
      RECT 86.16 2.395 86.68 2.565 ;
      RECT 86.36 6.255 86.68 6.545 ;
      RECT 86.33 6.285 86.68 6.515 ;
      RECT 86.16 6.315 86.68 6.485 ;
      RECT 81.81 3.57 82.13 3.83 ;
      RECT 83.1 2.745 83.24 3.605 ;
      RECT 81.9 3.465 83.24 3.605 ;
      RECT 81.9 3.025 82.04 3.83 ;
      RECT 81.825 3.025 82.115 3.255 ;
      RECT 83.025 2.745 83.315 2.975 ;
      RECT 82.545 3.025 82.835 3.255 ;
      RECT 82.74 1.95 82.88 3.21 ;
      RECT 82.77 1.89 83.09 2.15 ;
      RECT 79.37 2.45 79.69 2.71 ;
      RECT 82.065 2.465 82.355 2.695 ;
      RECT 79.46 2.37 82.28 2.51 ;
      RECT 81.33 1.89 81.65 2.15 ;
      RECT 81.825 1.905 82.115 2.135 ;
      RECT 81.33 1.95 82.115 2.09 ;
      RECT 81.33 3.01 81.65 3.27 ;
      RECT 81.33 2.79 81.56 3.27 ;
      RECT 80.825 2.745 81.115 2.975 ;
      RECT 80.825 2.79 81.56 2.93 ;
      RECT 81.09 7.765 81.38 7.995 ;
      RECT 81.15 7.025 81.32 7.995 ;
      RECT 81.05 7.055 81.43 7.425 ;
      RECT 81.09 7.025 81.38 7.425 ;
      RECT 79.85 3.57 80.17 3.83 ;
      RECT 79.385 3.585 79.675 3.815 ;
      RECT 79.385 3.63 80.17 3.77 ;
      RECT 78.145 2.465 78.435 2.695 ;
      RECT 78.145 2.51 79.08 2.65 ;
      RECT 78.94 1.95 79.08 2.65 ;
      RECT 79.61 1.89 79.93 2.15 ;
      RECT 79.385 1.905 79.93 2.135 ;
      RECT 78.94 1.95 79.93 2.09 ;
      RECT 77.29 3.57 77.61 3.83 ;
      RECT 77.29 3.63 78.36 3.77 ;
      RECT 78.22 3.07 78.36 3.77 ;
      RECT 79.385 3.025 79.675 3.255 ;
      RECT 78.22 3.07 79.675 3.21 ;
      RECT 77.65 1.89 77.97 2.15 ;
      RECT 77.425 1.905 77.97 2.135 ;
      RECT 76.67 2.45 76.99 2.71 ;
      RECT 77.665 2.465 77.955 2.695 ;
      RECT 76.425 2.465 76.99 2.695 ;
      RECT 76.425 2.51 77.955 2.65 ;
      RECT 75.945 3.025 76.235 3.255 ;
      RECT 76.14 1.95 76.28 3.21 ;
      RECT 76.93 1.89 77.25 2.15 ;
      RECT 75.945 1.905 76.235 2.135 ;
      RECT 75.945 1.95 77.25 2.09 ;
      RECT 75.54 3.465 76.64 3.605 ;
      RECT 76.425 3.305 76.715 3.535 ;
      RECT 75.465 3.305 75.755 3.535 ;
      RECT 75.45 1.89 75.77 2.15 ;
      RECT 73.49 1.89 73.81 2.15 ;
      RECT 73.49 1.95 75.77 2.09 ;
      RECT 74.61 3.01 74.93 3.27 ;
      RECT 74.61 3.01 75.44 3.15 ;
      RECT 75.225 2.745 75.44 3.15 ;
      RECT 75.225 2.745 75.515 2.975 ;
      RECT 73.01 2.45 73.33 2.71 ;
      RECT 74.42 2.465 74.71 2.695 ;
      RECT 73.01 2.465 73.555 2.695 ;
      RECT 73.01 2.55 73.96 2.69 ;
      RECT 73.82 2.37 73.96 2.69 ;
      RECT 74.32 2.465 74.71 2.65 ;
      RECT 73.82 2.37 74.46 2.51 ;
      RECT 72.53 3.26 72.85 3.675 ;
      RECT 72.61 1.905 72.765 3.675 ;
      RECT 72.545 1.905 72.835 2.135 ;
      RECT 70.925 7.77 71.215 8 ;
      RECT 70.985 6.29 71.155 8 ;
      RECT 70.935 6.655 71.285 7.005 ;
      RECT 70.925 6.29 71.215 6.52 ;
      RECT 70.52 2.395 70.625 2.965 ;
      RECT 70.52 2.73 70.845 2.96 ;
      RECT 70.52 2.76 71.015 2.93 ;
      RECT 70.52 2.395 70.71 2.96 ;
      RECT 69.935 2.36 70.225 2.59 ;
      RECT 69.935 2.395 70.71 2.565 ;
      RECT 69.995 0.88 70.165 2.59 ;
      RECT 69.935 0.88 70.225 1.11 ;
      RECT 69.935 7.77 70.225 8 ;
      RECT 69.995 6.29 70.165 8 ;
      RECT 69.935 6.29 70.225 6.52 ;
      RECT 69.935 6.325 70.79 6.485 ;
      RECT 70.62 5.92 70.79 6.485 ;
      RECT 69.935 6.32 70.33 6.485 ;
      RECT 70.555 5.92 70.845 6.15 ;
      RECT 70.555 5.95 71.015 6.12 ;
      RECT 69.565 2.73 69.855 2.96 ;
      RECT 69.565 2.76 70.025 2.93 ;
      RECT 69.63 1.655 69.795 2.96 ;
      RECT 68.145 1.625 68.435 1.855 ;
      RECT 68.145 1.655 69.795 1.825 ;
      RECT 68.205 0.885 68.375 1.855 ;
      RECT 68.145 0.885 68.435 1.115 ;
      RECT 68.145 7.765 68.435 7.995 ;
      RECT 68.205 7.025 68.375 7.995 ;
      RECT 68.205 7.12 69.795 7.29 ;
      RECT 69.625 5.92 69.795 7.29 ;
      RECT 68.145 7.025 68.435 7.255 ;
      RECT 69.565 5.92 69.855 6.15 ;
      RECT 69.565 5.95 70.025 6.12 ;
      RECT 66.195 3.15 66.535 3.5 ;
      RECT 66.285 2.025 66.455 3.5 ;
      RECT 68.575 1.965 68.925 2.315 ;
      RECT 66.285 2.025 68.925 2.195 ;
      RECT 68.6 6.655 68.925 6.98 ;
      RECT 63.16 6.61 63.51 6.96 ;
      RECT 68.575 6.655 68.925 6.885 ;
      RECT 62.96 6.655 63.51 6.885 ;
      RECT 62.79 6.685 68.925 6.855 ;
      RECT 67.8 2.365 68.12 2.685 ;
      RECT 67.77 2.365 68.12 2.595 ;
      RECT 67.6 2.395 68.12 2.565 ;
      RECT 67.8 6.255 68.12 6.545 ;
      RECT 67.77 6.285 68.12 6.515 ;
      RECT 67.6 6.315 68.12 6.485 ;
      RECT 63.25 3.57 63.57 3.83 ;
      RECT 64.54 2.745 64.68 3.605 ;
      RECT 63.34 3.465 64.68 3.605 ;
      RECT 63.34 3.025 63.48 3.83 ;
      RECT 63.265 3.025 63.555 3.255 ;
      RECT 64.465 2.745 64.755 2.975 ;
      RECT 63.985 3.025 64.275 3.255 ;
      RECT 64.18 1.95 64.32 3.21 ;
      RECT 64.21 1.89 64.53 2.15 ;
      RECT 60.81 2.45 61.13 2.71 ;
      RECT 63.505 2.465 63.795 2.695 ;
      RECT 60.9 2.37 63.72 2.51 ;
      RECT 62.77 1.89 63.09 2.15 ;
      RECT 63.265 1.905 63.555 2.135 ;
      RECT 62.77 1.95 63.555 2.09 ;
      RECT 62.77 3.01 63.09 3.27 ;
      RECT 62.77 2.79 63 3.27 ;
      RECT 62.265 2.745 62.555 2.975 ;
      RECT 62.265 2.79 63 2.93 ;
      RECT 62.53 7.765 62.82 7.995 ;
      RECT 62.59 7.025 62.76 7.995 ;
      RECT 62.49 7.055 62.87 7.425 ;
      RECT 62.53 7.025 62.82 7.425 ;
      RECT 61.29 3.57 61.61 3.83 ;
      RECT 60.825 3.585 61.115 3.815 ;
      RECT 60.825 3.63 61.61 3.77 ;
      RECT 59.585 2.465 59.875 2.695 ;
      RECT 59.585 2.51 60.52 2.65 ;
      RECT 60.38 1.95 60.52 2.65 ;
      RECT 61.05 1.89 61.37 2.15 ;
      RECT 60.825 1.905 61.37 2.135 ;
      RECT 60.38 1.95 61.37 2.09 ;
      RECT 58.73 3.57 59.05 3.83 ;
      RECT 58.73 3.63 59.8 3.77 ;
      RECT 59.66 3.07 59.8 3.77 ;
      RECT 60.825 3.025 61.115 3.255 ;
      RECT 59.66 3.07 61.115 3.21 ;
      RECT 59.09 1.89 59.41 2.15 ;
      RECT 58.865 1.905 59.41 2.135 ;
      RECT 58.11 2.45 58.43 2.71 ;
      RECT 59.105 2.465 59.395 2.695 ;
      RECT 57.865 2.465 58.43 2.695 ;
      RECT 57.865 2.51 59.395 2.65 ;
      RECT 57.385 3.025 57.675 3.255 ;
      RECT 57.58 1.95 57.72 3.21 ;
      RECT 58.37 1.89 58.69 2.15 ;
      RECT 57.385 1.905 57.675 2.135 ;
      RECT 57.385 1.95 58.69 2.09 ;
      RECT 56.98 3.465 58.08 3.605 ;
      RECT 57.865 3.305 58.155 3.535 ;
      RECT 56.905 3.305 57.195 3.535 ;
      RECT 56.89 1.89 57.21 2.15 ;
      RECT 54.93 1.89 55.25 2.15 ;
      RECT 54.93 1.95 57.21 2.09 ;
      RECT 56.05 3.01 56.37 3.27 ;
      RECT 56.05 3.01 56.88 3.15 ;
      RECT 56.665 2.745 56.88 3.15 ;
      RECT 56.665 2.745 56.955 2.975 ;
      RECT 54.45 2.45 54.77 2.71 ;
      RECT 55.86 2.465 56.15 2.695 ;
      RECT 54.45 2.465 54.995 2.695 ;
      RECT 54.45 2.55 55.4 2.69 ;
      RECT 55.26 2.37 55.4 2.69 ;
      RECT 55.76 2.465 56.15 2.65 ;
      RECT 55.26 2.37 55.9 2.51 ;
      RECT 53.97 3.26 54.29 3.675 ;
      RECT 54.05 1.905 54.205 3.675 ;
      RECT 53.985 1.905 54.275 2.135 ;
      RECT 52.365 7.77 52.655 8 ;
      RECT 52.425 6.29 52.595 8 ;
      RECT 52.375 6.655 52.725 7.005 ;
      RECT 52.365 6.29 52.655 6.52 ;
      RECT 51.96 2.395 52.065 2.965 ;
      RECT 51.96 2.73 52.285 2.96 ;
      RECT 51.96 2.76 52.455 2.93 ;
      RECT 51.96 2.395 52.15 2.96 ;
      RECT 51.375 2.36 51.665 2.59 ;
      RECT 51.375 2.395 52.15 2.565 ;
      RECT 51.435 0.88 51.605 2.59 ;
      RECT 51.375 0.88 51.665 1.11 ;
      RECT 51.375 7.77 51.665 8 ;
      RECT 51.435 6.29 51.605 8 ;
      RECT 51.375 6.29 51.665 6.52 ;
      RECT 51.375 6.325 52.23 6.485 ;
      RECT 52.06 5.92 52.23 6.485 ;
      RECT 51.375 6.32 51.77 6.485 ;
      RECT 51.995 5.92 52.285 6.15 ;
      RECT 51.995 5.95 52.455 6.12 ;
      RECT 51.005 2.73 51.295 2.96 ;
      RECT 51.005 2.76 51.465 2.93 ;
      RECT 51.07 1.655 51.235 2.96 ;
      RECT 49.585 1.625 49.875 1.855 ;
      RECT 49.585 1.655 51.235 1.825 ;
      RECT 49.645 0.885 49.815 1.855 ;
      RECT 49.585 0.885 49.875 1.115 ;
      RECT 49.585 7.765 49.875 7.995 ;
      RECT 49.645 7.025 49.815 7.995 ;
      RECT 49.645 7.12 51.235 7.29 ;
      RECT 51.065 5.92 51.235 7.29 ;
      RECT 49.585 7.025 49.875 7.255 ;
      RECT 51.005 5.92 51.295 6.15 ;
      RECT 51.005 5.95 51.465 6.12 ;
      RECT 47.635 3.15 47.975 3.5 ;
      RECT 47.725 2.025 47.895 3.5 ;
      RECT 50.015 1.965 50.365 2.315 ;
      RECT 47.725 2.025 50.365 2.195 ;
      RECT 50.04 6.655 50.365 6.98 ;
      RECT 44.6 6.615 44.95 6.965 ;
      RECT 50.015 6.655 50.365 6.885 ;
      RECT 44.4 6.655 44.95 6.885 ;
      RECT 44.23 6.685 50.365 6.855 ;
      RECT 49.24 2.365 49.56 2.685 ;
      RECT 49.21 2.365 49.56 2.595 ;
      RECT 49.04 2.395 49.56 2.565 ;
      RECT 49.24 6.255 49.56 6.545 ;
      RECT 49.21 6.285 49.56 6.515 ;
      RECT 49.04 6.315 49.56 6.485 ;
      RECT 44.69 3.57 45.01 3.83 ;
      RECT 45.98 2.745 46.12 3.605 ;
      RECT 44.78 3.465 46.12 3.605 ;
      RECT 44.78 3.025 44.92 3.83 ;
      RECT 44.705 3.025 44.995 3.255 ;
      RECT 45.905 2.745 46.195 2.975 ;
      RECT 45.425 3.025 45.715 3.255 ;
      RECT 45.62 1.95 45.76 3.21 ;
      RECT 45.65 1.89 45.97 2.15 ;
      RECT 42.25 2.45 42.57 2.71 ;
      RECT 44.945 2.465 45.235 2.695 ;
      RECT 42.34 2.37 45.16 2.51 ;
      RECT 44.21 1.89 44.53 2.15 ;
      RECT 44.705 1.905 44.995 2.135 ;
      RECT 44.21 1.95 44.995 2.09 ;
      RECT 44.21 3.01 44.53 3.27 ;
      RECT 44.21 2.79 44.44 3.27 ;
      RECT 43.705 2.745 43.995 2.975 ;
      RECT 43.705 2.79 44.44 2.93 ;
      RECT 43.97 7.765 44.26 7.995 ;
      RECT 44.03 7.025 44.2 7.995 ;
      RECT 43.93 7.055 44.31 7.425 ;
      RECT 43.97 7.025 44.26 7.425 ;
      RECT 42.73 3.57 43.05 3.83 ;
      RECT 42.265 3.585 42.555 3.815 ;
      RECT 42.265 3.63 43.05 3.77 ;
      RECT 41.025 2.465 41.315 2.695 ;
      RECT 41.025 2.51 41.96 2.65 ;
      RECT 41.82 1.95 41.96 2.65 ;
      RECT 42.49 1.89 42.81 2.15 ;
      RECT 42.265 1.905 42.81 2.135 ;
      RECT 41.82 1.95 42.81 2.09 ;
      RECT 40.17 3.57 40.49 3.83 ;
      RECT 40.17 3.63 41.24 3.77 ;
      RECT 41.1 3.07 41.24 3.77 ;
      RECT 42.265 3.025 42.555 3.255 ;
      RECT 41.1 3.07 42.555 3.21 ;
      RECT 40.53 1.89 40.85 2.15 ;
      RECT 40.305 1.905 40.85 2.135 ;
      RECT 39.55 2.45 39.87 2.71 ;
      RECT 40.545 2.465 40.835 2.695 ;
      RECT 39.305 2.465 39.87 2.695 ;
      RECT 39.305 2.51 40.835 2.65 ;
      RECT 38.825 3.025 39.115 3.255 ;
      RECT 39.02 1.95 39.16 3.21 ;
      RECT 39.81 1.89 40.13 2.15 ;
      RECT 38.825 1.905 39.115 2.135 ;
      RECT 38.825 1.95 40.13 2.09 ;
      RECT 38.42 3.465 39.52 3.605 ;
      RECT 39.305 3.305 39.595 3.535 ;
      RECT 38.345 3.305 38.635 3.535 ;
      RECT 38.33 1.89 38.65 2.15 ;
      RECT 36.37 1.89 36.69 2.15 ;
      RECT 36.37 1.95 38.65 2.09 ;
      RECT 37.49 3.01 37.81 3.27 ;
      RECT 37.49 3.01 38.32 3.15 ;
      RECT 38.105 2.745 38.32 3.15 ;
      RECT 38.105 2.745 38.395 2.975 ;
      RECT 35.89 2.45 36.21 2.71 ;
      RECT 37.3 2.465 37.59 2.695 ;
      RECT 35.89 2.465 36.435 2.695 ;
      RECT 35.89 2.55 36.84 2.69 ;
      RECT 36.7 2.37 36.84 2.69 ;
      RECT 37.2 2.465 37.59 2.65 ;
      RECT 36.7 2.37 37.34 2.51 ;
      RECT 35.41 3.26 35.73 3.675 ;
      RECT 35.49 1.905 35.645 3.675 ;
      RECT 35.425 1.905 35.715 2.135 ;
      RECT 33.805 7.77 34.095 8 ;
      RECT 33.865 6.29 34.035 8 ;
      RECT 33.855 6.66 34.21 7.015 ;
      RECT 33.805 6.29 34.095 6.52 ;
      RECT 33.4 2.395 33.505 2.965 ;
      RECT 33.4 2.73 33.725 2.96 ;
      RECT 33.4 2.76 33.895 2.93 ;
      RECT 33.4 2.395 33.59 2.96 ;
      RECT 32.815 2.36 33.105 2.59 ;
      RECT 32.815 2.395 33.59 2.565 ;
      RECT 32.875 0.88 33.045 2.59 ;
      RECT 32.815 0.88 33.105 1.11 ;
      RECT 32.815 7.77 33.105 8 ;
      RECT 32.875 6.29 33.045 8 ;
      RECT 32.815 6.29 33.105 6.52 ;
      RECT 32.815 6.325 33.67 6.485 ;
      RECT 33.5 5.92 33.67 6.485 ;
      RECT 32.815 6.32 33.21 6.485 ;
      RECT 33.435 5.92 33.725 6.15 ;
      RECT 33.435 5.95 33.895 6.12 ;
      RECT 32.445 2.73 32.735 2.96 ;
      RECT 32.445 2.76 32.905 2.93 ;
      RECT 32.51 1.655 32.675 2.96 ;
      RECT 31.025 1.625 31.315 1.855 ;
      RECT 31.025 1.655 32.675 1.825 ;
      RECT 31.085 0.885 31.255 1.855 ;
      RECT 31.025 0.885 31.315 1.115 ;
      RECT 31.025 7.765 31.315 7.995 ;
      RECT 31.085 7.025 31.255 7.995 ;
      RECT 31.085 7.12 32.675 7.29 ;
      RECT 32.505 5.92 32.675 7.29 ;
      RECT 31.025 7.025 31.315 7.255 ;
      RECT 32.445 5.92 32.735 6.15 ;
      RECT 32.445 5.95 32.905 6.12 ;
      RECT 29.075 3.15 29.415 3.5 ;
      RECT 29.165 2.025 29.335 3.5 ;
      RECT 31.455 1.965 31.805 2.315 ;
      RECT 29.165 2.025 31.805 2.195 ;
      RECT 31.48 6.655 31.805 6.98 ;
      RECT 26.045 6.61 26.395 6.96 ;
      RECT 31.455 6.655 31.805 6.885 ;
      RECT 25.84 6.655 26.395 6.885 ;
      RECT 25.67 6.685 31.805 6.855 ;
      RECT 30.68 2.365 31 2.685 ;
      RECT 30.65 2.365 31 2.595 ;
      RECT 30.48 2.395 31 2.565 ;
      RECT 30.68 6.255 31 6.545 ;
      RECT 30.65 6.285 31 6.515 ;
      RECT 30.48 6.315 31 6.485 ;
      RECT 26.13 3.57 26.45 3.83 ;
      RECT 27.42 2.745 27.56 3.605 ;
      RECT 26.22 3.465 27.56 3.605 ;
      RECT 26.22 3.025 26.36 3.83 ;
      RECT 26.145 3.025 26.435 3.255 ;
      RECT 27.345 2.745 27.635 2.975 ;
      RECT 26.865 3.025 27.155 3.255 ;
      RECT 27.06 1.95 27.2 3.21 ;
      RECT 27.09 1.89 27.41 2.15 ;
      RECT 23.69 2.45 24.01 2.71 ;
      RECT 26.385 2.465 26.675 2.695 ;
      RECT 23.78 2.37 26.6 2.51 ;
      RECT 25.65 1.89 25.97 2.15 ;
      RECT 26.145 1.905 26.435 2.135 ;
      RECT 25.65 1.95 26.435 2.09 ;
      RECT 25.65 3.01 25.97 3.27 ;
      RECT 25.65 2.79 25.88 3.27 ;
      RECT 25.145 2.745 25.435 2.975 ;
      RECT 25.145 2.79 25.88 2.93 ;
      RECT 25.41 7.765 25.7 7.995 ;
      RECT 25.47 7.025 25.64 7.995 ;
      RECT 25.37 7.055 25.75 7.425 ;
      RECT 25.41 7.025 25.7 7.425 ;
      RECT 24.17 3.57 24.49 3.83 ;
      RECT 23.705 3.585 23.995 3.815 ;
      RECT 23.705 3.63 24.49 3.77 ;
      RECT 22.465 2.465 22.755 2.695 ;
      RECT 22.465 2.51 23.4 2.65 ;
      RECT 23.26 1.95 23.4 2.65 ;
      RECT 23.93 1.89 24.25 2.15 ;
      RECT 23.705 1.905 24.25 2.135 ;
      RECT 23.26 1.95 24.25 2.09 ;
      RECT 21.61 3.57 21.93 3.83 ;
      RECT 21.61 3.63 22.68 3.77 ;
      RECT 22.54 3.07 22.68 3.77 ;
      RECT 23.705 3.025 23.995 3.255 ;
      RECT 22.54 3.07 23.995 3.21 ;
      RECT 21.97 1.89 22.29 2.15 ;
      RECT 21.745 1.905 22.29 2.135 ;
      RECT 20.99 2.45 21.31 2.71 ;
      RECT 21.985 2.465 22.275 2.695 ;
      RECT 20.745 2.465 21.31 2.695 ;
      RECT 20.745 2.51 22.275 2.65 ;
      RECT 20.265 3.025 20.555 3.255 ;
      RECT 20.46 1.95 20.6 3.21 ;
      RECT 21.25 1.89 21.57 2.15 ;
      RECT 20.265 1.905 20.555 2.135 ;
      RECT 20.265 1.95 21.57 2.09 ;
      RECT 19.86 3.465 20.96 3.605 ;
      RECT 20.745 3.305 21.035 3.535 ;
      RECT 19.785 3.305 20.075 3.535 ;
      RECT 19.77 1.89 20.09 2.15 ;
      RECT 17.81 1.89 18.13 2.15 ;
      RECT 17.81 1.95 20.09 2.09 ;
      RECT 18.93 3.01 19.25 3.27 ;
      RECT 18.93 3.01 19.76 3.15 ;
      RECT 19.545 2.745 19.76 3.15 ;
      RECT 19.545 2.745 19.835 2.975 ;
      RECT 17.33 2.45 17.65 2.71 ;
      RECT 18.74 2.465 19.03 2.695 ;
      RECT 17.33 2.465 17.875 2.695 ;
      RECT 17.33 2.55 18.28 2.69 ;
      RECT 18.14 2.37 18.28 2.69 ;
      RECT 18.64 2.465 19.03 2.65 ;
      RECT 18.14 2.37 18.78 2.51 ;
      RECT 16.85 3.26 17.17 3.675 ;
      RECT 16.93 1.905 17.085 3.675 ;
      RECT 16.865 1.905 17.155 2.135 ;
      RECT 15.245 7.77 15.535 8 ;
      RECT 15.305 6.29 15.475 8 ;
      RECT 15.3 6.655 15.65 7.005 ;
      RECT 15.245 6.29 15.535 6.52 ;
      RECT 14.84 2.395 14.945 2.965 ;
      RECT 14.84 2.73 15.165 2.96 ;
      RECT 14.84 2.76 15.335 2.93 ;
      RECT 14.84 2.395 15.03 2.96 ;
      RECT 14.255 2.36 14.545 2.59 ;
      RECT 14.255 2.395 15.03 2.565 ;
      RECT 14.315 0.88 14.485 2.59 ;
      RECT 14.255 0.88 14.545 1.11 ;
      RECT 14.255 7.77 14.545 8 ;
      RECT 14.315 6.29 14.485 8 ;
      RECT 14.255 6.29 14.545 6.52 ;
      RECT 14.255 6.325 15.11 6.485 ;
      RECT 14.94 5.92 15.11 6.485 ;
      RECT 14.255 6.32 14.65 6.485 ;
      RECT 14.875 5.92 15.165 6.15 ;
      RECT 14.875 5.95 15.335 6.12 ;
      RECT 13.885 2.73 14.175 2.96 ;
      RECT 13.885 2.76 14.345 2.93 ;
      RECT 13.95 1.655 14.115 2.96 ;
      RECT 12.465 1.625 12.755 1.855 ;
      RECT 12.465 1.655 14.115 1.825 ;
      RECT 12.525 0.885 12.695 1.855 ;
      RECT 12.465 0.885 12.755 1.115 ;
      RECT 12.465 7.765 12.755 7.995 ;
      RECT 12.525 7.025 12.695 7.995 ;
      RECT 12.525 7.12 14.115 7.29 ;
      RECT 13.945 5.92 14.115 7.29 ;
      RECT 12.465 7.025 12.755 7.255 ;
      RECT 13.885 5.92 14.175 6.15 ;
      RECT 13.885 5.95 14.345 6.12 ;
      RECT 10.515 3.15 10.855 3.5 ;
      RECT 10.605 2.025 10.775 3.5 ;
      RECT 12.895 1.965 13.245 2.315 ;
      RECT 10.605 2.025 13.245 2.195 ;
      RECT 12.92 6.655 13.245 6.98 ;
      RECT 7.485 6.605 7.835 6.955 ;
      RECT 12.895 6.655 13.245 6.885 ;
      RECT 7.28 6.655 7.835 6.885 ;
      RECT 7.11 6.685 13.245 6.855 ;
      RECT 12.12 2.365 12.44 2.685 ;
      RECT 12.09 2.365 12.44 2.595 ;
      RECT 11.92 2.395 12.44 2.565 ;
      RECT 12.12 6.255 12.44 6.545 ;
      RECT 12.09 6.285 12.44 6.515 ;
      RECT 11.92 6.315 12.44 6.485 ;
      RECT 7.57 3.57 7.89 3.83 ;
      RECT 8.86 2.745 9 3.605 ;
      RECT 7.66 3.465 9 3.605 ;
      RECT 7.66 3.025 7.8 3.83 ;
      RECT 7.585 3.025 7.875 3.255 ;
      RECT 8.785 2.745 9.075 2.975 ;
      RECT 8.305 3.025 8.595 3.255 ;
      RECT 8.5 1.95 8.64 3.21 ;
      RECT 8.53 1.89 8.85 2.15 ;
      RECT 5.13 2.45 5.45 2.71 ;
      RECT 7.825 2.465 8.115 2.695 ;
      RECT 5.22 2.37 8.04 2.51 ;
      RECT 7.09 1.89 7.41 2.15 ;
      RECT 7.585 1.905 7.875 2.135 ;
      RECT 7.09 1.95 7.875 2.09 ;
      RECT 7.09 3.01 7.41 3.27 ;
      RECT 7.09 2.79 7.32 3.27 ;
      RECT 6.585 2.745 6.875 2.975 ;
      RECT 6.585 2.79 7.32 2.93 ;
      RECT 6.85 7.765 7.14 7.995 ;
      RECT 6.91 7.025 7.08 7.995 ;
      RECT 6.81 7.055 7.19 7.425 ;
      RECT 6.85 7.025 7.14 7.425 ;
      RECT 5.61 3.57 5.93 3.83 ;
      RECT 5.145 3.585 5.435 3.815 ;
      RECT 5.145 3.63 5.93 3.77 ;
      RECT 3.905 2.465 4.195 2.695 ;
      RECT 3.905 2.51 4.84 2.65 ;
      RECT 4.7 1.95 4.84 2.65 ;
      RECT 5.37 1.89 5.69 2.15 ;
      RECT 5.145 1.905 5.69 2.135 ;
      RECT 4.7 1.95 5.69 2.09 ;
      RECT 3.05 3.57 3.37 3.83 ;
      RECT 3.05 3.63 4.12 3.77 ;
      RECT 3.98 3.07 4.12 3.77 ;
      RECT 5.145 3.025 5.435 3.255 ;
      RECT 3.98 3.07 5.435 3.21 ;
      RECT 3.41 1.89 3.73 2.15 ;
      RECT 3.185 1.905 3.73 2.135 ;
      RECT 2.43 2.45 2.75 2.71 ;
      RECT 3.425 2.465 3.715 2.695 ;
      RECT 2.185 2.465 2.75 2.695 ;
      RECT 2.185 2.51 3.715 2.65 ;
      RECT 1.705 3.025 1.995 3.255 ;
      RECT 1.9 1.95 2.04 3.21 ;
      RECT 2.69 1.89 3.01 2.15 ;
      RECT 1.705 1.905 1.995 2.135 ;
      RECT 1.705 1.95 3.01 2.09 ;
      RECT 1.3 3.465 2.4 3.605 ;
      RECT 2.185 3.305 2.475 3.535 ;
      RECT 1.225 3.305 1.515 3.535 ;
      RECT 1.21 1.89 1.53 2.15 ;
      RECT -0.75 1.89 -0.43 2.15 ;
      RECT -0.75 1.95 1.53 2.09 ;
      RECT 0.37 3.01 0.69 3.27 ;
      RECT 0.37 3.01 1.2 3.15 ;
      RECT 0.985 2.745 1.2 3.15 ;
      RECT 0.985 2.745 1.275 2.975 ;
      RECT -1.23 2.45 -0.91 2.71 ;
      RECT 0.18 2.465 0.47 2.695 ;
      RECT -1.23 2.465 -0.685 2.695 ;
      RECT -1.23 2.55 -0.28 2.69 ;
      RECT -0.42 2.37 -0.28 2.69 ;
      RECT 0.08 2.465 0.47 2.65 ;
      RECT -0.42 2.37 0.22 2.51 ;
      RECT -1.71 3.26 -1.39 3.675 ;
      RECT -1.63 1.905 -1.475 3.675 ;
      RECT -1.695 1.905 -1.405 2.135 ;
      RECT -3.965 7.765 -3.675 7.995 ;
      RECT -3.905 7.025 -3.735 7.995 ;
      RECT -3.995 7.025 -3.645 7.315 ;
      RECT -4.37 6.285 -4.02 6.575 ;
      RECT -4.51 6.315 -4.02 6.485 ;
      RECT 80.81 3.57 81.13 3.83 ;
      RECT 80.21 1.89 80.89 2.15 ;
      RECT 80.33 3.57 80.65 3.83 ;
      RECT 78.85 3.57 79.17 3.83 ;
      RECT 78.37 1.89 78.69 2.15 ;
      RECT 77.65 3.01 77.97 3.27 ;
      RECT 76.93 3.01 77.25 3.27 ;
      RECT 73.49 3.01 73.81 3.27 ;
      RECT 62.25 3.57 62.57 3.83 ;
      RECT 61.65 1.89 62.33 2.15 ;
      RECT 61.77 3.57 62.09 3.83 ;
      RECT 60.29 3.57 60.61 3.83 ;
      RECT 59.81 1.89 60.13 2.15 ;
      RECT 59.09 3.01 59.41 3.27 ;
      RECT 58.37 3.01 58.69 3.27 ;
      RECT 54.93 3.01 55.25 3.27 ;
      RECT 43.69 3.57 44.01 3.83 ;
      RECT 43.09 1.89 43.77 2.15 ;
      RECT 43.21 3.57 43.53 3.83 ;
      RECT 41.73 3.57 42.05 3.83 ;
      RECT 41.25 1.89 41.57 2.15 ;
      RECT 40.53 3.01 40.85 3.27 ;
      RECT 39.81 3.01 40.13 3.27 ;
      RECT 36.37 3.01 36.69 3.27 ;
      RECT 25.13 3.57 25.45 3.83 ;
      RECT 24.53 1.89 25.21 2.15 ;
      RECT 24.65 3.57 24.97 3.83 ;
      RECT 23.17 3.57 23.49 3.83 ;
      RECT 22.69 1.89 23.01 2.15 ;
      RECT 21.97 3.01 22.29 3.27 ;
      RECT 21.25 3.01 21.57 3.27 ;
      RECT 17.81 3.01 18.13 3.27 ;
      RECT 6.57 3.57 6.89 3.83 ;
      RECT 5.97 1.89 6.65 2.15 ;
      RECT 6.09 3.57 6.41 3.83 ;
      RECT 4.61 3.57 4.93 3.83 ;
      RECT 4.13 1.89 4.45 2.15 ;
      RECT 3.41 3.01 3.73 3.27 ;
      RECT 2.69 3.01 3.01 3.27 ;
      RECT -0.75 3.01 -0.43 3.27 ;
    LAYER mcon ;
      RECT 89.545 6.32 89.715 6.49 ;
      RECT 89.55 6.315 89.72 6.485 ;
      RECT 70.985 6.32 71.155 6.49 ;
      RECT 70.99 6.315 71.16 6.485 ;
      RECT 52.425 6.32 52.595 6.49 ;
      RECT 52.43 6.315 52.6 6.485 ;
      RECT 33.865 6.32 34.035 6.49 ;
      RECT 33.87 6.315 34.04 6.485 ;
      RECT 15.305 6.32 15.475 6.49 ;
      RECT 15.31 6.315 15.48 6.485 ;
      RECT 89.545 7.8 89.715 7.97 ;
      RECT 89.175 2.76 89.345 2.93 ;
      RECT 89.175 5.95 89.345 6.12 ;
      RECT 88.555 0.91 88.725 1.08 ;
      RECT 88.555 2.39 88.725 2.56 ;
      RECT 88.555 6.32 88.725 6.49 ;
      RECT 88.555 7.8 88.725 7.97 ;
      RECT 88.185 2.76 88.355 2.93 ;
      RECT 88.185 5.95 88.355 6.12 ;
      RECT 87.195 2.025 87.365 2.195 ;
      RECT 87.195 6.685 87.365 6.855 ;
      RECT 86.765 0.915 86.935 1.085 ;
      RECT 86.765 1.655 86.935 1.825 ;
      RECT 86.765 7.055 86.935 7.225 ;
      RECT 86.765 7.795 86.935 7.965 ;
      RECT 86.39 2.395 86.56 2.565 ;
      RECT 86.39 6.315 86.56 6.485 ;
      RECT 83.085 2.775 83.255 2.945 ;
      RECT 82.845 1.935 83.015 2.105 ;
      RECT 82.605 3.055 82.775 3.225 ;
      RECT 82.125 2.495 82.295 2.665 ;
      RECT 81.885 1.935 82.055 2.105 ;
      RECT 81.885 3.055 82.055 3.225 ;
      RECT 81.885 3.615 82.055 3.785 ;
      RECT 81.58 6.685 81.75 6.855 ;
      RECT 81.405 3.055 81.575 3.225 ;
      RECT 81.15 7.055 81.32 7.225 ;
      RECT 81.15 7.795 81.32 7.965 ;
      RECT 80.885 2.775 81.055 2.945 ;
      RECT 80.885 3.615 81.055 3.785 ;
      RECT 80.405 1.935 80.575 2.105 ;
      RECT 80.405 3.615 80.575 3.785 ;
      RECT 79.445 1.935 79.615 2.105 ;
      RECT 79.445 2.495 79.615 2.665 ;
      RECT 79.445 3.055 79.615 3.225 ;
      RECT 79.445 3.615 79.615 3.785 ;
      RECT 78.925 3.615 79.095 3.785 ;
      RECT 78.445 1.935 78.615 2.105 ;
      RECT 78.205 2.495 78.375 2.665 ;
      RECT 77.725 2.495 77.895 2.665 ;
      RECT 77.725 3.055 77.895 3.225 ;
      RECT 77.485 1.935 77.655 2.105 ;
      RECT 77.005 3.055 77.175 3.225 ;
      RECT 76.485 2.495 76.655 2.665 ;
      RECT 76.485 3.335 76.655 3.505 ;
      RECT 76.005 1.935 76.175 2.105 ;
      RECT 76.005 3.055 76.175 3.225 ;
      RECT 75.525 3.335 75.695 3.505 ;
      RECT 75.285 2.775 75.455 2.945 ;
      RECT 74.48 2.495 74.65 2.665 ;
      RECT 73.565 1.935 73.735 2.105 ;
      RECT 73.565 3.055 73.735 3.225 ;
      RECT 73.325 2.495 73.495 2.665 ;
      RECT 72.605 1.935 72.775 2.105 ;
      RECT 72.605 3.475 72.775 3.645 ;
      RECT 70.985 7.8 71.155 7.97 ;
      RECT 70.615 2.76 70.785 2.93 ;
      RECT 70.615 5.95 70.785 6.12 ;
      RECT 69.995 0.91 70.165 1.08 ;
      RECT 69.995 2.39 70.165 2.56 ;
      RECT 69.995 6.32 70.165 6.49 ;
      RECT 69.995 7.8 70.165 7.97 ;
      RECT 69.625 2.76 69.795 2.93 ;
      RECT 69.625 5.95 69.795 6.12 ;
      RECT 68.635 2.025 68.805 2.195 ;
      RECT 68.635 6.685 68.805 6.855 ;
      RECT 68.205 0.915 68.375 1.085 ;
      RECT 68.205 1.655 68.375 1.825 ;
      RECT 68.205 7.055 68.375 7.225 ;
      RECT 68.205 7.795 68.375 7.965 ;
      RECT 67.83 2.395 68 2.565 ;
      RECT 67.83 6.315 68 6.485 ;
      RECT 64.525 2.775 64.695 2.945 ;
      RECT 64.285 1.935 64.455 2.105 ;
      RECT 64.045 3.055 64.215 3.225 ;
      RECT 63.565 2.495 63.735 2.665 ;
      RECT 63.325 1.935 63.495 2.105 ;
      RECT 63.325 3.055 63.495 3.225 ;
      RECT 63.325 3.615 63.495 3.785 ;
      RECT 63.02 6.685 63.19 6.855 ;
      RECT 62.845 3.055 63.015 3.225 ;
      RECT 62.59 7.055 62.76 7.225 ;
      RECT 62.59 7.795 62.76 7.965 ;
      RECT 62.325 2.775 62.495 2.945 ;
      RECT 62.325 3.615 62.495 3.785 ;
      RECT 61.845 1.935 62.015 2.105 ;
      RECT 61.845 3.615 62.015 3.785 ;
      RECT 60.885 1.935 61.055 2.105 ;
      RECT 60.885 2.495 61.055 2.665 ;
      RECT 60.885 3.055 61.055 3.225 ;
      RECT 60.885 3.615 61.055 3.785 ;
      RECT 60.365 3.615 60.535 3.785 ;
      RECT 59.885 1.935 60.055 2.105 ;
      RECT 59.645 2.495 59.815 2.665 ;
      RECT 59.165 2.495 59.335 2.665 ;
      RECT 59.165 3.055 59.335 3.225 ;
      RECT 58.925 1.935 59.095 2.105 ;
      RECT 58.445 3.055 58.615 3.225 ;
      RECT 57.925 2.495 58.095 2.665 ;
      RECT 57.925 3.335 58.095 3.505 ;
      RECT 57.445 1.935 57.615 2.105 ;
      RECT 57.445 3.055 57.615 3.225 ;
      RECT 56.965 3.335 57.135 3.505 ;
      RECT 56.725 2.775 56.895 2.945 ;
      RECT 55.92 2.495 56.09 2.665 ;
      RECT 55.005 1.935 55.175 2.105 ;
      RECT 55.005 3.055 55.175 3.225 ;
      RECT 54.765 2.495 54.935 2.665 ;
      RECT 54.045 1.935 54.215 2.105 ;
      RECT 54.045 3.475 54.215 3.645 ;
      RECT 52.425 7.8 52.595 7.97 ;
      RECT 52.055 2.76 52.225 2.93 ;
      RECT 52.055 5.95 52.225 6.12 ;
      RECT 51.435 0.91 51.605 1.08 ;
      RECT 51.435 2.39 51.605 2.56 ;
      RECT 51.435 6.32 51.605 6.49 ;
      RECT 51.435 7.8 51.605 7.97 ;
      RECT 51.065 2.76 51.235 2.93 ;
      RECT 51.065 5.95 51.235 6.12 ;
      RECT 50.075 2.025 50.245 2.195 ;
      RECT 50.075 6.685 50.245 6.855 ;
      RECT 49.645 0.915 49.815 1.085 ;
      RECT 49.645 1.655 49.815 1.825 ;
      RECT 49.645 7.055 49.815 7.225 ;
      RECT 49.645 7.795 49.815 7.965 ;
      RECT 49.27 2.395 49.44 2.565 ;
      RECT 49.27 6.315 49.44 6.485 ;
      RECT 45.965 2.775 46.135 2.945 ;
      RECT 45.725 1.935 45.895 2.105 ;
      RECT 45.485 3.055 45.655 3.225 ;
      RECT 45.005 2.495 45.175 2.665 ;
      RECT 44.765 1.935 44.935 2.105 ;
      RECT 44.765 3.055 44.935 3.225 ;
      RECT 44.765 3.615 44.935 3.785 ;
      RECT 44.46 6.685 44.63 6.855 ;
      RECT 44.285 3.055 44.455 3.225 ;
      RECT 44.03 7.055 44.2 7.225 ;
      RECT 44.03 7.795 44.2 7.965 ;
      RECT 43.765 2.775 43.935 2.945 ;
      RECT 43.765 3.615 43.935 3.785 ;
      RECT 43.285 1.935 43.455 2.105 ;
      RECT 43.285 3.615 43.455 3.785 ;
      RECT 42.325 1.935 42.495 2.105 ;
      RECT 42.325 2.495 42.495 2.665 ;
      RECT 42.325 3.055 42.495 3.225 ;
      RECT 42.325 3.615 42.495 3.785 ;
      RECT 41.805 3.615 41.975 3.785 ;
      RECT 41.325 1.935 41.495 2.105 ;
      RECT 41.085 2.495 41.255 2.665 ;
      RECT 40.605 2.495 40.775 2.665 ;
      RECT 40.605 3.055 40.775 3.225 ;
      RECT 40.365 1.935 40.535 2.105 ;
      RECT 39.885 3.055 40.055 3.225 ;
      RECT 39.365 2.495 39.535 2.665 ;
      RECT 39.365 3.335 39.535 3.505 ;
      RECT 38.885 1.935 39.055 2.105 ;
      RECT 38.885 3.055 39.055 3.225 ;
      RECT 38.405 3.335 38.575 3.505 ;
      RECT 38.165 2.775 38.335 2.945 ;
      RECT 37.36 2.495 37.53 2.665 ;
      RECT 36.445 1.935 36.615 2.105 ;
      RECT 36.445 3.055 36.615 3.225 ;
      RECT 36.205 2.495 36.375 2.665 ;
      RECT 35.485 1.935 35.655 2.105 ;
      RECT 35.485 3.475 35.655 3.645 ;
      RECT 33.865 7.8 34.035 7.97 ;
      RECT 33.495 2.76 33.665 2.93 ;
      RECT 33.495 5.95 33.665 6.12 ;
      RECT 32.875 0.91 33.045 1.08 ;
      RECT 32.875 2.39 33.045 2.56 ;
      RECT 32.875 6.32 33.045 6.49 ;
      RECT 32.875 7.8 33.045 7.97 ;
      RECT 32.505 2.76 32.675 2.93 ;
      RECT 32.505 5.95 32.675 6.12 ;
      RECT 31.515 2.025 31.685 2.195 ;
      RECT 31.515 6.685 31.685 6.855 ;
      RECT 31.085 0.915 31.255 1.085 ;
      RECT 31.085 1.655 31.255 1.825 ;
      RECT 31.085 7.055 31.255 7.225 ;
      RECT 31.085 7.795 31.255 7.965 ;
      RECT 30.71 2.395 30.88 2.565 ;
      RECT 30.71 6.315 30.88 6.485 ;
      RECT 27.405 2.775 27.575 2.945 ;
      RECT 27.165 1.935 27.335 2.105 ;
      RECT 26.925 3.055 27.095 3.225 ;
      RECT 26.445 2.495 26.615 2.665 ;
      RECT 26.205 1.935 26.375 2.105 ;
      RECT 26.205 3.055 26.375 3.225 ;
      RECT 26.205 3.615 26.375 3.785 ;
      RECT 25.9 6.685 26.07 6.855 ;
      RECT 25.725 3.055 25.895 3.225 ;
      RECT 25.47 7.055 25.64 7.225 ;
      RECT 25.47 7.795 25.64 7.965 ;
      RECT 25.205 2.775 25.375 2.945 ;
      RECT 25.205 3.615 25.375 3.785 ;
      RECT 24.725 1.935 24.895 2.105 ;
      RECT 24.725 3.615 24.895 3.785 ;
      RECT 23.765 1.935 23.935 2.105 ;
      RECT 23.765 2.495 23.935 2.665 ;
      RECT 23.765 3.055 23.935 3.225 ;
      RECT 23.765 3.615 23.935 3.785 ;
      RECT 23.245 3.615 23.415 3.785 ;
      RECT 22.765 1.935 22.935 2.105 ;
      RECT 22.525 2.495 22.695 2.665 ;
      RECT 22.045 2.495 22.215 2.665 ;
      RECT 22.045 3.055 22.215 3.225 ;
      RECT 21.805 1.935 21.975 2.105 ;
      RECT 21.325 3.055 21.495 3.225 ;
      RECT 20.805 2.495 20.975 2.665 ;
      RECT 20.805 3.335 20.975 3.505 ;
      RECT 20.325 1.935 20.495 2.105 ;
      RECT 20.325 3.055 20.495 3.225 ;
      RECT 19.845 3.335 20.015 3.505 ;
      RECT 19.605 2.775 19.775 2.945 ;
      RECT 18.8 2.495 18.97 2.665 ;
      RECT 17.885 1.935 18.055 2.105 ;
      RECT 17.885 3.055 18.055 3.225 ;
      RECT 17.645 2.495 17.815 2.665 ;
      RECT 16.925 1.935 17.095 2.105 ;
      RECT 16.925 3.475 17.095 3.645 ;
      RECT 15.305 7.8 15.475 7.97 ;
      RECT 14.935 2.76 15.105 2.93 ;
      RECT 14.935 5.95 15.105 6.12 ;
      RECT 14.315 0.91 14.485 1.08 ;
      RECT 14.315 2.39 14.485 2.56 ;
      RECT 14.315 6.32 14.485 6.49 ;
      RECT 14.315 7.8 14.485 7.97 ;
      RECT 13.945 2.76 14.115 2.93 ;
      RECT 13.945 5.95 14.115 6.12 ;
      RECT 12.955 2.025 13.125 2.195 ;
      RECT 12.955 6.685 13.125 6.855 ;
      RECT 12.525 0.915 12.695 1.085 ;
      RECT 12.525 1.655 12.695 1.825 ;
      RECT 12.525 7.055 12.695 7.225 ;
      RECT 12.525 7.795 12.695 7.965 ;
      RECT 12.15 2.395 12.32 2.565 ;
      RECT 12.15 6.315 12.32 6.485 ;
      RECT 8.845 2.775 9.015 2.945 ;
      RECT 8.605 1.935 8.775 2.105 ;
      RECT 8.365 3.055 8.535 3.225 ;
      RECT 7.885 2.495 8.055 2.665 ;
      RECT 7.645 1.935 7.815 2.105 ;
      RECT 7.645 3.055 7.815 3.225 ;
      RECT 7.645 3.615 7.815 3.785 ;
      RECT 7.34 6.685 7.51 6.855 ;
      RECT 7.165 3.055 7.335 3.225 ;
      RECT 6.91 7.055 7.08 7.225 ;
      RECT 6.91 7.795 7.08 7.965 ;
      RECT 6.645 2.775 6.815 2.945 ;
      RECT 6.645 3.615 6.815 3.785 ;
      RECT 6.165 1.935 6.335 2.105 ;
      RECT 6.165 3.615 6.335 3.785 ;
      RECT 5.205 1.935 5.375 2.105 ;
      RECT 5.205 2.495 5.375 2.665 ;
      RECT 5.205 3.055 5.375 3.225 ;
      RECT 5.205 3.615 5.375 3.785 ;
      RECT 4.685 3.615 4.855 3.785 ;
      RECT 4.205 1.935 4.375 2.105 ;
      RECT 3.965 2.495 4.135 2.665 ;
      RECT 3.485 2.495 3.655 2.665 ;
      RECT 3.485 3.055 3.655 3.225 ;
      RECT 3.245 1.935 3.415 2.105 ;
      RECT 2.765 3.055 2.935 3.225 ;
      RECT 2.245 2.495 2.415 2.665 ;
      RECT 2.245 3.335 2.415 3.505 ;
      RECT 1.765 1.935 1.935 2.105 ;
      RECT 1.765 3.055 1.935 3.225 ;
      RECT 1.285 3.335 1.455 3.505 ;
      RECT 1.045 2.775 1.215 2.945 ;
      RECT 0.24 2.495 0.41 2.665 ;
      RECT -0.675 1.935 -0.505 2.105 ;
      RECT -0.675 3.055 -0.505 3.225 ;
      RECT -0.915 2.495 -0.745 2.665 ;
      RECT -1.635 1.935 -1.465 2.105 ;
      RECT -1.635 3.475 -1.465 3.645 ;
      RECT -3.905 7.055 -3.735 7.225 ;
      RECT -3.905 7.795 -3.735 7.965 ;
      RECT -4.28 6.315 -4.11 6.485 ;
    LAYER li1 ;
      RECT 89.545 5.02 89.715 6.49 ;
      RECT 89.545 6.315 89.72 6.485 ;
      RECT 89.175 1.74 89.345 2.93 ;
      RECT 89.175 1.74 89.645 1.91 ;
      RECT 89.175 6.97 89.645 7.14 ;
      RECT 89.175 5.95 89.345 7.14 ;
      RECT 88.185 1.74 88.355 2.93 ;
      RECT 88.185 1.74 88.655 1.91 ;
      RECT 88.185 6.97 88.655 7.14 ;
      RECT 88.185 5.95 88.355 7.14 ;
      RECT 86.335 2.635 86.505 3.865 ;
      RECT 86.39 0.855 86.56 2.805 ;
      RECT 86.335 0.575 86.505 1.025 ;
      RECT 86.335 7.855 86.505 8.305 ;
      RECT 86.39 6.075 86.56 8.025 ;
      RECT 86.335 5.015 86.505 6.245 ;
      RECT 85.815 0.575 85.985 3.865 ;
      RECT 85.815 2.075 86.22 2.405 ;
      RECT 85.815 1.235 86.22 1.565 ;
      RECT 85.815 5.015 85.985 8.305 ;
      RECT 85.815 7.315 86.22 7.645 ;
      RECT 85.815 6.475 86.22 6.805 ;
      RECT 82.605 3.225 83.575 3.395 ;
      RECT 82.605 3.055 82.775 3.395 ;
      RECT 82.125 2.495 82.295 2.825 ;
      RECT 82.125 2.575 82.855 2.745 ;
      RECT 81.765 3.615 82.055 3.785 ;
      RECT 81.765 2.575 81.935 3.785 ;
      RECT 81.765 3.055 82.055 3.225 ;
      RECT 81.565 2.575 81.935 2.745 ;
      RECT 80.885 2.675 81.055 2.945 ;
      RECT 80.645 2.675 81.055 2.845 ;
      RECT 80.565 2.575 80.895 2.745 ;
      RECT 80.405 3.615 81.055 3.785 ;
      RECT 80.885 3.145 81.055 3.785 ;
      RECT 80.765 3.225 81.055 3.785 ;
      RECT 80.2 5.015 80.37 8.305 ;
      RECT 80.2 7.315 80.605 7.645 ;
      RECT 80.2 6.475 80.605 6.805 ;
      RECT 79.445 2.915 79.615 3.225 ;
      RECT 79.445 2.915 80.335 3.085 ;
      RECT 80.165 2.495 80.335 3.085 ;
      RECT 79.445 2.575 79.935 2.745 ;
      RECT 79.445 2.495 79.615 2.745 ;
      RECT 77.405 3.225 77.895 3.395 ;
      RECT 78.565 2.575 78.735 3.225 ;
      RECT 77.725 3.055 78.735 3.225 ;
      RECT 78.685 2.495 78.855 2.825 ;
      RECT 77.485 1.835 77.655 2.105 ;
      RECT 76.925 1.835 77.655 2.005 ;
      RECT 77.005 2.575 77.175 3.225 ;
      RECT 77.005 2.575 77.495 2.745 ;
      RECT 76.165 2.575 76.655 2.745 ;
      RECT 76.485 2.495 76.655 2.745 ;
      RECT 76.005 1.835 76.175 2.105 ;
      RECT 75.445 1.835 76.175 2.005 ;
      RECT 75.525 3.225 75.695 3.505 ;
      RECT 74.485 3.225 75.775 3.395 ;
      RECT 74.48 2.575 75.055 2.745 ;
      RECT 74.48 2.495 74.65 2.745 ;
      RECT 73.565 1.835 73.735 2.105 ;
      RECT 73.565 1.835 74.295 2.005 ;
      RECT 73.565 3.055 73.735 3.475 ;
      RECT 72.945 3.14 73.735 3.31 ;
      RECT 72.945 2.915 73.115 3.31 ;
      RECT 72.845 2.495 73.015 3.085 ;
      RECT 72.605 2.575 73.015 2.845 ;
      RECT 70.985 5.02 71.155 6.49 ;
      RECT 70.985 6.315 71.16 6.485 ;
      RECT 70.615 1.74 70.785 2.93 ;
      RECT 70.615 1.74 71.085 1.91 ;
      RECT 70.615 6.97 71.085 7.14 ;
      RECT 70.615 5.95 70.785 7.14 ;
      RECT 69.625 1.74 69.795 2.93 ;
      RECT 69.625 1.74 70.095 1.91 ;
      RECT 69.625 6.97 70.095 7.14 ;
      RECT 69.625 5.95 69.795 7.14 ;
      RECT 67.775 2.635 67.945 3.865 ;
      RECT 67.83 0.855 68 2.805 ;
      RECT 67.775 0.575 67.945 1.025 ;
      RECT 67.775 7.855 67.945 8.305 ;
      RECT 67.83 6.075 68 8.025 ;
      RECT 67.775 5.015 67.945 6.245 ;
      RECT 67.255 0.575 67.425 3.865 ;
      RECT 67.255 2.075 67.66 2.405 ;
      RECT 67.255 1.235 67.66 1.565 ;
      RECT 67.255 5.015 67.425 8.305 ;
      RECT 67.255 7.315 67.66 7.645 ;
      RECT 67.255 6.475 67.66 6.805 ;
      RECT 64.045 3.225 65.015 3.395 ;
      RECT 64.045 3.055 64.215 3.395 ;
      RECT 63.565 2.495 63.735 2.825 ;
      RECT 63.565 2.575 64.295 2.745 ;
      RECT 63.205 3.615 63.495 3.785 ;
      RECT 63.205 2.575 63.375 3.785 ;
      RECT 63.205 3.055 63.495 3.225 ;
      RECT 63.005 2.575 63.375 2.745 ;
      RECT 62.325 2.675 62.495 2.945 ;
      RECT 62.085 2.675 62.495 2.845 ;
      RECT 62.005 2.575 62.335 2.745 ;
      RECT 61.845 3.615 62.495 3.785 ;
      RECT 62.325 3.145 62.495 3.785 ;
      RECT 62.205 3.225 62.495 3.785 ;
      RECT 61.64 5.015 61.81 8.305 ;
      RECT 61.64 7.315 62.045 7.645 ;
      RECT 61.64 6.475 62.045 6.805 ;
      RECT 60.885 2.915 61.055 3.225 ;
      RECT 60.885 2.915 61.775 3.085 ;
      RECT 61.605 2.495 61.775 3.085 ;
      RECT 60.885 2.575 61.375 2.745 ;
      RECT 60.885 2.495 61.055 2.745 ;
      RECT 58.845 3.225 59.335 3.395 ;
      RECT 60.005 2.575 60.175 3.225 ;
      RECT 59.165 3.055 60.175 3.225 ;
      RECT 60.125 2.495 60.295 2.825 ;
      RECT 58.925 1.835 59.095 2.105 ;
      RECT 58.365 1.835 59.095 2.005 ;
      RECT 58.445 2.575 58.615 3.225 ;
      RECT 58.445 2.575 58.935 2.745 ;
      RECT 57.605 2.575 58.095 2.745 ;
      RECT 57.925 2.495 58.095 2.745 ;
      RECT 57.445 1.835 57.615 2.105 ;
      RECT 56.885 1.835 57.615 2.005 ;
      RECT 56.965 3.225 57.135 3.505 ;
      RECT 55.925 3.225 57.215 3.395 ;
      RECT 55.92 2.575 56.495 2.745 ;
      RECT 55.92 2.495 56.09 2.745 ;
      RECT 55.005 1.835 55.175 2.105 ;
      RECT 55.005 1.835 55.735 2.005 ;
      RECT 55.005 3.055 55.175 3.475 ;
      RECT 54.385 3.14 55.175 3.31 ;
      RECT 54.385 2.915 54.555 3.31 ;
      RECT 54.285 2.495 54.455 3.085 ;
      RECT 54.045 2.575 54.455 2.845 ;
      RECT 52.425 5.02 52.595 6.49 ;
      RECT 52.425 6.315 52.6 6.485 ;
      RECT 52.055 1.74 52.225 2.93 ;
      RECT 52.055 1.74 52.525 1.91 ;
      RECT 52.055 6.97 52.525 7.14 ;
      RECT 52.055 5.95 52.225 7.14 ;
      RECT 51.065 1.74 51.235 2.93 ;
      RECT 51.065 1.74 51.535 1.91 ;
      RECT 51.065 6.97 51.535 7.14 ;
      RECT 51.065 5.95 51.235 7.14 ;
      RECT 49.215 2.635 49.385 3.865 ;
      RECT 49.27 0.855 49.44 2.805 ;
      RECT 49.215 0.575 49.385 1.025 ;
      RECT 49.215 7.855 49.385 8.305 ;
      RECT 49.27 6.075 49.44 8.025 ;
      RECT 49.215 5.015 49.385 6.245 ;
      RECT 48.695 0.575 48.865 3.865 ;
      RECT 48.695 2.075 49.1 2.405 ;
      RECT 48.695 1.235 49.1 1.565 ;
      RECT 48.695 5.015 48.865 8.305 ;
      RECT 48.695 7.315 49.1 7.645 ;
      RECT 48.695 6.475 49.1 6.805 ;
      RECT 45.485 3.225 46.455 3.395 ;
      RECT 45.485 3.055 45.655 3.395 ;
      RECT 45.005 2.495 45.175 2.825 ;
      RECT 45.005 2.575 45.735 2.745 ;
      RECT 44.645 3.615 44.935 3.785 ;
      RECT 44.645 2.575 44.815 3.785 ;
      RECT 44.645 3.055 44.935 3.225 ;
      RECT 44.445 2.575 44.815 2.745 ;
      RECT 43.765 2.675 43.935 2.945 ;
      RECT 43.525 2.675 43.935 2.845 ;
      RECT 43.445 2.575 43.775 2.745 ;
      RECT 43.285 3.615 43.935 3.785 ;
      RECT 43.765 3.145 43.935 3.785 ;
      RECT 43.645 3.225 43.935 3.785 ;
      RECT 43.08 5.015 43.25 8.305 ;
      RECT 43.08 7.315 43.485 7.645 ;
      RECT 43.08 6.475 43.485 6.805 ;
      RECT 42.325 2.915 42.495 3.225 ;
      RECT 42.325 2.915 43.215 3.085 ;
      RECT 43.045 2.495 43.215 3.085 ;
      RECT 42.325 2.575 42.815 2.745 ;
      RECT 42.325 2.495 42.495 2.745 ;
      RECT 40.285 3.225 40.775 3.395 ;
      RECT 41.445 2.575 41.615 3.225 ;
      RECT 40.605 3.055 41.615 3.225 ;
      RECT 41.565 2.495 41.735 2.825 ;
      RECT 40.365 1.835 40.535 2.105 ;
      RECT 39.805 1.835 40.535 2.005 ;
      RECT 39.885 2.575 40.055 3.225 ;
      RECT 39.885 2.575 40.375 2.745 ;
      RECT 39.045 2.575 39.535 2.745 ;
      RECT 39.365 2.495 39.535 2.745 ;
      RECT 38.885 1.835 39.055 2.105 ;
      RECT 38.325 1.835 39.055 2.005 ;
      RECT 38.405 3.225 38.575 3.505 ;
      RECT 37.365 3.225 38.655 3.395 ;
      RECT 37.36 2.575 37.935 2.745 ;
      RECT 37.36 2.495 37.53 2.745 ;
      RECT 36.445 1.835 36.615 2.105 ;
      RECT 36.445 1.835 37.175 2.005 ;
      RECT 36.445 3.055 36.615 3.475 ;
      RECT 35.825 3.14 36.615 3.31 ;
      RECT 35.825 2.915 35.995 3.31 ;
      RECT 35.725 2.495 35.895 3.085 ;
      RECT 35.485 2.575 35.895 2.845 ;
      RECT 33.865 5.02 34.035 6.49 ;
      RECT 33.865 6.315 34.04 6.485 ;
      RECT 33.495 1.74 33.665 2.93 ;
      RECT 33.495 1.74 33.965 1.91 ;
      RECT 33.495 6.97 33.965 7.14 ;
      RECT 33.495 5.95 33.665 7.14 ;
      RECT 32.505 1.74 32.675 2.93 ;
      RECT 32.505 1.74 32.975 1.91 ;
      RECT 32.505 6.97 32.975 7.14 ;
      RECT 32.505 5.95 32.675 7.14 ;
      RECT 30.655 2.635 30.825 3.865 ;
      RECT 30.71 0.855 30.88 2.805 ;
      RECT 30.655 0.575 30.825 1.025 ;
      RECT 30.655 7.855 30.825 8.305 ;
      RECT 30.71 6.075 30.88 8.025 ;
      RECT 30.655 5.015 30.825 6.245 ;
      RECT 30.135 0.575 30.305 3.865 ;
      RECT 30.135 2.075 30.54 2.405 ;
      RECT 30.135 1.235 30.54 1.565 ;
      RECT 30.135 5.015 30.305 8.305 ;
      RECT 30.135 7.315 30.54 7.645 ;
      RECT 30.135 6.475 30.54 6.805 ;
      RECT 26.925 3.225 27.895 3.395 ;
      RECT 26.925 3.055 27.095 3.395 ;
      RECT 26.445 2.495 26.615 2.825 ;
      RECT 26.445 2.575 27.175 2.745 ;
      RECT 26.085 3.615 26.375 3.785 ;
      RECT 26.085 2.575 26.255 3.785 ;
      RECT 26.085 3.055 26.375 3.225 ;
      RECT 25.885 2.575 26.255 2.745 ;
      RECT 25.205 2.675 25.375 2.945 ;
      RECT 24.965 2.675 25.375 2.845 ;
      RECT 24.885 2.575 25.215 2.745 ;
      RECT 24.725 3.615 25.375 3.785 ;
      RECT 25.205 3.145 25.375 3.785 ;
      RECT 25.085 3.225 25.375 3.785 ;
      RECT 24.52 5.015 24.69 8.305 ;
      RECT 24.52 7.315 24.925 7.645 ;
      RECT 24.52 6.475 24.925 6.805 ;
      RECT 23.765 2.915 23.935 3.225 ;
      RECT 23.765 2.915 24.655 3.085 ;
      RECT 24.485 2.495 24.655 3.085 ;
      RECT 23.765 2.575 24.255 2.745 ;
      RECT 23.765 2.495 23.935 2.745 ;
      RECT 21.725 3.225 22.215 3.395 ;
      RECT 22.885 2.575 23.055 3.225 ;
      RECT 22.045 3.055 23.055 3.225 ;
      RECT 23.005 2.495 23.175 2.825 ;
      RECT 21.805 1.835 21.975 2.105 ;
      RECT 21.245 1.835 21.975 2.005 ;
      RECT 21.325 2.575 21.495 3.225 ;
      RECT 21.325 2.575 21.815 2.745 ;
      RECT 20.485 2.575 20.975 2.745 ;
      RECT 20.805 2.495 20.975 2.745 ;
      RECT 20.325 1.835 20.495 2.105 ;
      RECT 19.765 1.835 20.495 2.005 ;
      RECT 19.845 3.225 20.015 3.505 ;
      RECT 18.805 3.225 20.095 3.395 ;
      RECT 18.8 2.575 19.375 2.745 ;
      RECT 18.8 2.495 18.97 2.745 ;
      RECT 17.885 1.835 18.055 2.105 ;
      RECT 17.885 1.835 18.615 2.005 ;
      RECT 17.885 3.055 18.055 3.475 ;
      RECT 17.265 3.14 18.055 3.31 ;
      RECT 17.265 2.915 17.435 3.31 ;
      RECT 17.165 2.495 17.335 3.085 ;
      RECT 16.925 2.575 17.335 2.845 ;
      RECT 15.305 5.02 15.475 6.49 ;
      RECT 15.305 6.315 15.48 6.485 ;
      RECT 14.935 1.74 15.105 2.93 ;
      RECT 14.935 1.74 15.405 1.91 ;
      RECT 14.935 6.97 15.405 7.14 ;
      RECT 14.935 5.95 15.105 7.14 ;
      RECT 13.945 1.74 14.115 2.93 ;
      RECT 13.945 1.74 14.415 1.91 ;
      RECT 13.945 6.97 14.415 7.14 ;
      RECT 13.945 5.95 14.115 7.14 ;
      RECT 12.095 2.635 12.265 3.865 ;
      RECT 12.15 0.855 12.32 2.805 ;
      RECT 12.095 0.575 12.265 1.025 ;
      RECT 12.095 7.855 12.265 8.305 ;
      RECT 12.15 6.075 12.32 8.025 ;
      RECT 12.095 5.015 12.265 6.245 ;
      RECT 11.575 0.575 11.745 3.865 ;
      RECT 11.575 2.075 11.98 2.405 ;
      RECT 11.575 1.235 11.98 1.565 ;
      RECT 11.575 5.015 11.745 8.305 ;
      RECT 11.575 7.315 11.98 7.645 ;
      RECT 11.575 6.475 11.98 6.805 ;
      RECT 8.365 3.225 9.335 3.395 ;
      RECT 8.365 3.055 8.535 3.395 ;
      RECT 7.885 2.495 8.055 2.825 ;
      RECT 7.885 2.575 8.615 2.745 ;
      RECT 7.525 3.615 7.815 3.785 ;
      RECT 7.525 2.575 7.695 3.785 ;
      RECT 7.525 3.055 7.815 3.225 ;
      RECT 7.325 2.575 7.695 2.745 ;
      RECT 6.645 2.675 6.815 2.945 ;
      RECT 6.405 2.675 6.815 2.845 ;
      RECT 6.325 2.575 6.655 2.745 ;
      RECT 6.165 3.615 6.815 3.785 ;
      RECT 6.645 3.145 6.815 3.785 ;
      RECT 6.525 3.225 6.815 3.785 ;
      RECT 5.96 5.015 6.13 8.305 ;
      RECT 5.96 7.315 6.365 7.645 ;
      RECT 5.96 6.475 6.365 6.805 ;
      RECT 5.205 2.915 5.375 3.225 ;
      RECT 5.205 2.915 6.095 3.085 ;
      RECT 5.925 2.495 6.095 3.085 ;
      RECT 5.205 2.575 5.695 2.745 ;
      RECT 5.205 2.495 5.375 2.745 ;
      RECT 3.165 3.225 3.655 3.395 ;
      RECT 4.325 2.575 4.495 3.225 ;
      RECT 3.485 3.055 4.495 3.225 ;
      RECT 4.445 2.495 4.615 2.825 ;
      RECT 3.245 1.835 3.415 2.105 ;
      RECT 2.685 1.835 3.415 2.005 ;
      RECT 2.765 2.575 2.935 3.225 ;
      RECT 2.765 2.575 3.255 2.745 ;
      RECT 1.925 2.575 2.415 2.745 ;
      RECT 2.245 2.495 2.415 2.745 ;
      RECT 1.765 1.835 1.935 2.105 ;
      RECT 1.205 1.835 1.935 2.005 ;
      RECT 1.285 3.225 1.455 3.505 ;
      RECT 0.245 3.225 1.535 3.395 ;
      RECT 0.24 2.575 0.815 2.745 ;
      RECT 0.24 2.495 0.41 2.745 ;
      RECT -0.675 1.835 -0.505 2.105 ;
      RECT -0.675 1.835 0.055 2.005 ;
      RECT -0.675 3.055 -0.505 3.475 ;
      RECT -1.295 3.14 -0.505 3.31 ;
      RECT -1.295 2.915 -1.125 3.31 ;
      RECT -1.395 2.495 -1.225 3.085 ;
      RECT -1.635 2.575 -1.225 2.845 ;
      RECT -4.335 7.855 -4.165 8.305 ;
      RECT -4.28 6.075 -4.11 8.025 ;
      RECT -4.335 5.015 -4.165 6.245 ;
      RECT -4.855 5.015 -4.685 8.305 ;
      RECT -4.855 7.315 -4.45 7.645 ;
      RECT -4.855 6.475 -4.45 6.805 ;
      RECT 89.545 7.8 89.715 8.31 ;
      RECT 88.555 0.57 88.725 1.08 ;
      RECT 88.555 2.39 88.725 3.86 ;
      RECT 88.555 5.02 88.725 6.49 ;
      RECT 88.555 7.8 88.725 8.31 ;
      RECT 87.195 0.575 87.365 3.865 ;
      RECT 87.195 5.015 87.365 8.305 ;
      RECT 86.765 0.575 86.935 1.085 ;
      RECT 86.765 1.655 86.935 3.865 ;
      RECT 86.765 5.015 86.935 7.225 ;
      RECT 86.765 7.795 86.935 8.305 ;
      RECT 83.085 2.495 83.255 2.945 ;
      RECT 82.845 1.755 83.015 2.105 ;
      RECT 81.885 1.755 82.055 2.105 ;
      RECT 81.58 5.015 81.75 8.305 ;
      RECT 81.405 3.055 81.575 3.475 ;
      RECT 81.15 5.015 81.32 7.225 ;
      RECT 81.15 7.795 81.32 8.305 ;
      RECT 80.405 1.755 80.575 2.105 ;
      RECT 79.445 1.755 79.615 2.105 ;
      RECT 79.445 3.485 79.615 3.815 ;
      RECT 78.925 3.145 79.095 3.785 ;
      RECT 78.445 1.755 78.615 2.105 ;
      RECT 78.205 2.495 78.375 2.825 ;
      RECT 77.725 2.495 77.895 2.825 ;
      RECT 76.485 3.145 76.655 3.505 ;
      RECT 76.005 3.055 76.175 3.475 ;
      RECT 75.285 2.495 75.455 2.945 ;
      RECT 73.325 2.495 73.495 2.825 ;
      RECT 72.605 1.755 72.775 2.105 ;
      RECT 72.605 3.285 72.775 3.645 ;
      RECT 70.985 7.8 71.155 8.31 ;
      RECT 69.995 0.57 70.165 1.08 ;
      RECT 69.995 2.39 70.165 3.86 ;
      RECT 69.995 5.02 70.165 6.49 ;
      RECT 69.995 7.8 70.165 8.31 ;
      RECT 68.635 0.575 68.805 3.865 ;
      RECT 68.635 5.015 68.805 8.305 ;
      RECT 68.205 0.575 68.375 1.085 ;
      RECT 68.205 1.655 68.375 3.865 ;
      RECT 68.205 5.015 68.375 7.225 ;
      RECT 68.205 7.795 68.375 8.305 ;
      RECT 64.525 2.495 64.695 2.945 ;
      RECT 64.285 1.755 64.455 2.105 ;
      RECT 63.325 1.755 63.495 2.105 ;
      RECT 63.02 5.015 63.19 8.305 ;
      RECT 62.845 3.055 63.015 3.475 ;
      RECT 62.59 5.015 62.76 7.225 ;
      RECT 62.59 7.795 62.76 8.305 ;
      RECT 61.845 1.755 62.015 2.105 ;
      RECT 60.885 1.755 61.055 2.105 ;
      RECT 60.885 3.485 61.055 3.815 ;
      RECT 60.365 3.145 60.535 3.785 ;
      RECT 59.885 1.755 60.055 2.105 ;
      RECT 59.645 2.495 59.815 2.825 ;
      RECT 59.165 2.495 59.335 2.825 ;
      RECT 57.925 3.145 58.095 3.505 ;
      RECT 57.445 3.055 57.615 3.475 ;
      RECT 56.725 2.495 56.895 2.945 ;
      RECT 54.765 2.495 54.935 2.825 ;
      RECT 54.045 1.755 54.215 2.105 ;
      RECT 54.045 3.285 54.215 3.645 ;
      RECT 52.425 7.8 52.595 8.31 ;
      RECT 51.435 0.57 51.605 1.08 ;
      RECT 51.435 2.39 51.605 3.86 ;
      RECT 51.435 5.02 51.605 6.49 ;
      RECT 51.435 7.8 51.605 8.31 ;
      RECT 50.075 0.575 50.245 3.865 ;
      RECT 50.075 5.015 50.245 8.305 ;
      RECT 49.645 0.575 49.815 1.085 ;
      RECT 49.645 1.655 49.815 3.865 ;
      RECT 49.645 5.015 49.815 7.225 ;
      RECT 49.645 7.795 49.815 8.305 ;
      RECT 45.965 2.495 46.135 2.945 ;
      RECT 45.725 1.755 45.895 2.105 ;
      RECT 44.765 1.755 44.935 2.105 ;
      RECT 44.46 5.015 44.63 8.305 ;
      RECT 44.285 3.055 44.455 3.475 ;
      RECT 44.03 5.015 44.2 7.225 ;
      RECT 44.03 7.795 44.2 8.305 ;
      RECT 43.285 1.755 43.455 2.105 ;
      RECT 42.325 1.755 42.495 2.105 ;
      RECT 42.325 3.485 42.495 3.815 ;
      RECT 41.805 3.145 41.975 3.785 ;
      RECT 41.325 1.755 41.495 2.105 ;
      RECT 41.085 2.495 41.255 2.825 ;
      RECT 40.605 2.495 40.775 2.825 ;
      RECT 39.365 3.145 39.535 3.505 ;
      RECT 38.885 3.055 39.055 3.475 ;
      RECT 38.165 2.495 38.335 2.945 ;
      RECT 36.205 2.495 36.375 2.825 ;
      RECT 35.485 1.755 35.655 2.105 ;
      RECT 35.485 3.285 35.655 3.645 ;
      RECT 33.865 7.8 34.035 8.31 ;
      RECT 32.875 0.57 33.045 1.08 ;
      RECT 32.875 2.39 33.045 3.86 ;
      RECT 32.875 5.02 33.045 6.49 ;
      RECT 32.875 7.8 33.045 8.31 ;
      RECT 31.515 0.575 31.685 3.865 ;
      RECT 31.515 5.015 31.685 8.305 ;
      RECT 31.085 0.575 31.255 1.085 ;
      RECT 31.085 1.655 31.255 3.865 ;
      RECT 31.085 5.015 31.255 7.225 ;
      RECT 31.085 7.795 31.255 8.305 ;
      RECT 27.405 2.495 27.575 2.945 ;
      RECT 27.165 1.755 27.335 2.105 ;
      RECT 26.205 1.755 26.375 2.105 ;
      RECT 25.9 5.015 26.07 8.305 ;
      RECT 25.725 3.055 25.895 3.475 ;
      RECT 25.47 5.015 25.64 7.225 ;
      RECT 25.47 7.795 25.64 8.305 ;
      RECT 24.725 1.755 24.895 2.105 ;
      RECT 23.765 1.755 23.935 2.105 ;
      RECT 23.765 3.485 23.935 3.815 ;
      RECT 23.245 3.145 23.415 3.785 ;
      RECT 22.765 1.755 22.935 2.105 ;
      RECT 22.525 2.495 22.695 2.825 ;
      RECT 22.045 2.495 22.215 2.825 ;
      RECT 20.805 3.145 20.975 3.505 ;
      RECT 20.325 3.055 20.495 3.475 ;
      RECT 19.605 2.495 19.775 2.945 ;
      RECT 17.645 2.495 17.815 2.825 ;
      RECT 16.925 1.755 17.095 2.105 ;
      RECT 16.925 3.285 17.095 3.645 ;
      RECT 15.305 7.8 15.475 8.31 ;
      RECT 14.315 0.57 14.485 1.08 ;
      RECT 14.315 2.39 14.485 3.86 ;
      RECT 14.315 5.02 14.485 6.49 ;
      RECT 14.315 7.8 14.485 8.31 ;
      RECT 12.955 0.575 13.125 3.865 ;
      RECT 12.955 5.015 13.125 8.305 ;
      RECT 12.525 0.575 12.695 1.085 ;
      RECT 12.525 1.655 12.695 3.865 ;
      RECT 12.525 5.015 12.695 7.225 ;
      RECT 12.525 7.795 12.695 8.305 ;
      RECT 8.845 2.495 9.015 2.945 ;
      RECT 8.605 1.755 8.775 2.105 ;
      RECT 7.645 1.755 7.815 2.105 ;
      RECT 7.34 5.015 7.51 8.305 ;
      RECT 7.165 3.055 7.335 3.475 ;
      RECT 6.91 5.015 7.08 7.225 ;
      RECT 6.91 7.795 7.08 8.305 ;
      RECT 6.165 1.755 6.335 2.105 ;
      RECT 5.205 1.755 5.375 2.105 ;
      RECT 5.205 3.485 5.375 3.815 ;
      RECT 4.685 3.145 4.855 3.785 ;
      RECT 4.205 1.755 4.375 2.105 ;
      RECT 3.965 2.495 4.135 2.825 ;
      RECT 3.485 2.495 3.655 2.825 ;
      RECT 2.245 3.145 2.415 3.505 ;
      RECT 1.765 3.055 1.935 3.475 ;
      RECT 1.045 2.495 1.215 2.945 ;
      RECT -0.915 2.495 -0.745 2.825 ;
      RECT -1.635 1.755 -1.465 2.105 ;
      RECT -1.635 3.285 -1.465 3.645 ;
      RECT -3.905 5.015 -3.735 7.225 ;
      RECT -3.905 7.795 -3.735 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2et_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2xa_8_b0r1
  CLASS BLOCK ;
  ORIGIN 2.8 -0.005 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2xa_8_b0r1 ;
  SIZE 79.1 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 14.72 0.92 14.89 1.09 ;
        RECT 14.715 0.915 14.885 1.085 ;
        RECT 14.715 2.395 14.885 2.565 ;
      LAYER li1 ;
        RECT 14.72 0.92 14.89 1.09 ;
        RECT 14.715 0.575 14.885 1.085 ;
        RECT 14.715 2.395 14.885 3.865 ;
      LAYER met1 ;
        RECT 14.655 2.365 14.945 2.595 ;
        RECT 14.655 0.885 14.945 1.115 ;
        RECT 14.715 0.885 14.885 2.595 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 29.98 0.92 30.15 1.09 ;
        RECT 29.975 0.915 30.145 1.085 ;
        RECT 29.975 2.395 30.145 2.565 ;
      LAYER li1 ;
        RECT 29.98 0.92 30.15 1.09 ;
        RECT 29.975 0.575 30.145 1.085 ;
        RECT 29.975 2.395 30.145 3.865 ;
      LAYER met1 ;
        RECT 29.915 2.365 30.205 2.595 ;
        RECT 29.915 0.885 30.205 1.115 ;
        RECT 29.975 0.885 30.145 2.595 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 45.24 0.92 45.41 1.09 ;
        RECT 45.235 0.915 45.405 1.085 ;
        RECT 45.235 2.395 45.405 2.565 ;
      LAYER li1 ;
        RECT 45.24 0.92 45.41 1.09 ;
        RECT 45.235 0.575 45.405 1.085 ;
        RECT 45.235 2.395 45.405 3.865 ;
      LAYER met1 ;
        RECT 45.175 2.365 45.465 2.595 ;
        RECT 45.175 0.885 45.465 1.115 ;
        RECT 45.235 0.885 45.405 2.595 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 60.5 0.92 60.67 1.09 ;
        RECT 60.495 0.915 60.665 1.085 ;
        RECT 60.495 2.395 60.665 2.565 ;
      LAYER li1 ;
        RECT 60.5 0.92 60.67 1.09 ;
        RECT 60.495 0.575 60.665 1.085 ;
        RECT 60.495 2.395 60.665 3.865 ;
      LAYER met1 ;
        RECT 60.435 2.365 60.725 2.595 ;
        RECT 60.435 0.885 60.725 1.115 ;
        RECT 60.495 0.885 60.665 2.595 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 75.76 0.92 75.93 1.09 ;
        RECT 75.755 0.915 75.925 1.085 ;
        RECT 75.755 2.395 75.925 2.565 ;
      LAYER li1 ;
        RECT 75.76 0.92 75.93 1.09 ;
        RECT 75.755 0.575 75.925 1.085 ;
        RECT 75.755 2.395 75.925 3.865 ;
      LAYER met1 ;
        RECT 75.695 2.365 75.985 2.595 ;
        RECT 75.695 0.885 75.985 1.115 ;
        RECT 75.755 0.885 75.925 2.595 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 10.485 5.865 10.825 6.215 ;
        RECT 10.485 2.71 10.825 3.06 ;
        RECT 10.565 2.71 10.735 6.215 ;
      LAYER li1 ;
        RECT 10.565 1.665 10.735 2.94 ;
        RECT 10.565 5.95 10.735 7.225 ;
        RECT 4.95 5.95 5.12 7.225 ;
      LAYER met1 ;
        RECT 10.485 2.77 10.965 2.94 ;
        RECT 10.485 2.71 10.825 3.06 ;
        RECT 4.89 5.95 10.965 6.12 ;
        RECT 10.485 5.865 10.825 6.215 ;
        RECT 4.89 5.92 5.18 6.15 ;
      LAYER via1 ;
        RECT 10.585 5.965 10.735 6.115 ;
        RECT 10.585 2.81 10.735 2.96 ;
      LAYER mcon ;
        RECT 4.95 5.95 5.12 6.12 ;
        RECT 10.565 5.95 10.735 6.12 ;
        RECT 10.565 2.77 10.735 2.94 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 25.745 5.865 26.085 6.215 ;
        RECT 25.745 2.71 26.085 3.06 ;
        RECT 25.825 2.71 25.995 6.215 ;
      LAYER li1 ;
        RECT 25.825 1.665 25.995 2.94 ;
        RECT 25.825 5.95 25.995 7.225 ;
        RECT 20.21 5.95 20.38 7.225 ;
      LAYER met1 ;
        RECT 25.745 2.77 26.225 2.94 ;
        RECT 25.745 2.71 26.085 3.06 ;
        RECT 20.15 5.95 26.225 6.12 ;
        RECT 25.745 5.865 26.085 6.215 ;
        RECT 20.15 5.92 20.44 6.15 ;
      LAYER via1 ;
        RECT 25.845 5.965 25.995 6.115 ;
        RECT 25.845 2.81 25.995 2.96 ;
      LAYER mcon ;
        RECT 20.21 5.95 20.38 6.12 ;
        RECT 25.825 5.95 25.995 6.12 ;
        RECT 25.825 2.77 25.995 2.94 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 41.005 5.865 41.345 6.215 ;
        RECT 41.005 2.71 41.345 3.06 ;
        RECT 41.085 2.71 41.255 6.215 ;
      LAYER li1 ;
        RECT 41.085 1.665 41.255 2.94 ;
        RECT 41.085 5.95 41.255 7.225 ;
        RECT 35.47 5.95 35.64 7.225 ;
      LAYER met1 ;
        RECT 41.005 2.77 41.485 2.94 ;
        RECT 41.005 2.71 41.345 3.06 ;
        RECT 35.41 5.95 41.485 6.12 ;
        RECT 41.005 5.865 41.345 6.215 ;
        RECT 35.41 5.92 35.7 6.15 ;
      LAYER via1 ;
        RECT 41.105 5.965 41.255 6.115 ;
        RECT 41.105 2.81 41.255 2.96 ;
      LAYER mcon ;
        RECT 35.47 5.95 35.64 6.12 ;
        RECT 41.085 5.95 41.255 6.12 ;
        RECT 41.085 2.77 41.255 2.94 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 56.265 5.865 56.605 6.215 ;
        RECT 56.265 2.71 56.605 3.06 ;
        RECT 56.345 2.71 56.515 6.215 ;
      LAYER li1 ;
        RECT 56.345 1.665 56.515 2.94 ;
        RECT 56.345 5.95 56.515 7.225 ;
        RECT 50.73 5.95 50.9 7.225 ;
      LAYER met1 ;
        RECT 56.265 2.77 56.745 2.94 ;
        RECT 56.265 2.71 56.605 3.06 ;
        RECT 50.67 5.95 56.745 6.12 ;
        RECT 56.265 5.865 56.605 6.215 ;
        RECT 50.67 5.92 50.96 6.15 ;
      LAYER via1 ;
        RECT 56.365 5.965 56.515 6.115 ;
        RECT 56.365 2.81 56.515 2.96 ;
      LAYER mcon ;
        RECT 50.73 5.95 50.9 6.12 ;
        RECT 56.345 5.95 56.515 6.12 ;
        RECT 56.345 2.77 56.515 2.94 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 71.525 5.865 71.865 6.215 ;
        RECT 71.525 2.71 71.865 3.06 ;
        RECT 71.605 2.71 71.775 6.215 ;
      LAYER li1 ;
        RECT 71.605 1.665 71.775 2.94 ;
        RECT 71.605 5.95 71.775 7.225 ;
        RECT 65.99 5.95 66.16 7.225 ;
      LAYER met1 ;
        RECT 71.525 2.77 72.005 2.94 ;
        RECT 71.525 2.71 71.865 3.06 ;
        RECT 65.93 5.95 72.005 6.12 ;
        RECT 71.525 5.865 71.865 6.215 ;
        RECT 65.93 5.92 66.22 6.15 ;
      LAYER via1 ;
        RECT 71.625 5.965 71.775 6.115 ;
        RECT 71.625 2.81 71.775 2.96 ;
      LAYER mcon ;
        RECT 65.99 5.95 66.16 6.12 ;
        RECT 71.605 5.95 71.775 6.12 ;
        RECT 71.605 2.77 71.775 2.94 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT -2.565 5.95 -2.395 7.225 ;
      LAYER met1 ;
        RECT -2.625 5.95 -2.165 6.12 ;
        RECT -2.625 5.92 -2.335 6.15 ;
      LAYER mcon ;
        RECT -2.565 5.95 -2.395 6.12 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT -2.75 4.145 76.3 4.75 ;
        RECT 61.79 4.14 76.3 4.75 ;
        RECT 74.165 4.135 76.145 4.755 ;
        RECT 75.325 3.405 75.495 5.485 ;
        RECT 74.335 3.405 74.505 5.485 ;
        RECT 71.595 3.41 71.765 5.48 ;
        RECT 68.82 3.64 68.99 4.75 ;
        RECT 66.9 3.64 67.07 4.75 ;
        RECT 65.98 4.14 66.15 5.48 ;
        RECT 65.96 3.64 66.13 4.75 ;
        RECT 64.5 3.64 64.67 4.75 ;
        RECT 62.58 3.64 62.75 4.75 ;
        RECT 46.53 4.14 61.04 4.75 ;
        RECT 58.905 4.135 60.885 4.755 ;
        RECT 60.065 3.405 60.235 5.485 ;
        RECT 59.075 3.405 59.245 5.485 ;
        RECT 56.335 3.41 56.505 5.48 ;
        RECT 53.56 3.64 53.73 4.75 ;
        RECT 51.64 3.64 51.81 4.75 ;
        RECT 50.72 4.14 50.89 5.48 ;
        RECT 50.7 3.64 50.87 4.75 ;
        RECT 49.24 3.64 49.41 4.75 ;
        RECT 47.32 3.64 47.49 4.75 ;
        RECT 31.27 4.14 45.78 4.75 ;
        RECT 43.645 4.135 45.625 4.755 ;
        RECT 44.805 3.405 44.975 5.485 ;
        RECT 43.815 3.405 43.985 5.485 ;
        RECT 41.075 3.41 41.245 5.48 ;
        RECT 38.3 3.64 38.47 4.75 ;
        RECT 36.38 3.64 36.55 4.75 ;
        RECT 35.46 4.14 35.63 5.48 ;
        RECT 35.44 3.64 35.61 4.75 ;
        RECT 33.98 3.64 34.15 4.75 ;
        RECT 32.06 3.64 32.23 4.75 ;
        RECT 16.01 4.14 30.52 4.75 ;
        RECT 28.385 4.135 30.365 4.755 ;
        RECT 29.545 3.405 29.715 5.485 ;
        RECT 28.555 3.405 28.725 5.485 ;
        RECT 25.815 3.41 25.985 5.48 ;
        RECT 23.04 3.64 23.21 4.75 ;
        RECT 21.12 3.64 21.29 4.75 ;
        RECT 20.2 4.14 20.37 5.48 ;
        RECT 20.18 3.64 20.35 4.75 ;
        RECT 18.72 3.64 18.89 4.75 ;
        RECT 16.8 3.64 16.97 4.75 ;
        RECT 0.75 4.14 15.26 4.75 ;
        RECT 13.125 4.135 15.105 4.755 ;
        RECT 14.285 3.405 14.455 5.485 ;
        RECT 13.295 3.405 13.465 5.485 ;
        RECT 10.555 3.41 10.725 5.48 ;
        RECT 7.78 3.64 7.95 4.75 ;
        RECT 5.86 3.64 6.03 4.75 ;
        RECT 4.94 4.14 5.11 5.48 ;
        RECT 4.92 3.64 5.09 4.75 ;
        RECT 3.46 3.64 3.63 4.75 ;
        RECT 1.54 3.64 1.71 4.75 ;
        RECT -0.765 4.145 -0.595 8.31 ;
        RECT -2.575 4.145 -2.405 5.48 ;
      LAYER met1 ;
        RECT -2.75 4.145 76.3 4.75 ;
        RECT 61.79 4.14 76.3 4.75 ;
        RECT 74.165 4.135 76.145 4.755 ;
        RECT 61.79 3.985 70.53 4.75 ;
        RECT 46.53 4.14 61.04 4.75 ;
        RECT 58.905 4.135 60.885 4.755 ;
        RECT 46.53 3.985 55.27 4.75 ;
        RECT 31.27 4.14 45.78 4.75 ;
        RECT 43.645 4.135 45.625 4.755 ;
        RECT 31.27 3.985 40.01 4.75 ;
        RECT 16.01 4.14 30.52 4.75 ;
        RECT 28.385 4.135 30.365 4.755 ;
        RECT 16.01 3.985 24.75 4.75 ;
        RECT 0.75 4.14 15.26 4.75 ;
        RECT 13.125 4.135 15.105 4.755 ;
        RECT 0.75 3.985 9.49 4.75 ;
        RECT -0.825 6.66 -0.535 6.89 ;
        RECT -0.995 6.69 -0.535 6.86 ;
      LAYER mcon ;
        RECT -0.765 6.69 -0.595 6.86 ;
        RECT -0.455 4.55 -0.285 4.72 ;
        RECT 0.895 4.14 1.065 4.31 ;
        RECT 1.355 4.14 1.525 4.31 ;
        RECT 1.815 4.14 1.985 4.31 ;
        RECT 2.275 4.14 2.445 4.31 ;
        RECT 2.735 4.14 2.905 4.31 ;
        RECT 3.195 4.14 3.365 4.31 ;
        RECT 3.655 4.14 3.825 4.31 ;
        RECT 4.115 4.14 4.285 4.31 ;
        RECT 4.575 4.14 4.745 4.31 ;
        RECT 5.035 4.14 5.205 4.31 ;
        RECT 5.495 4.14 5.665 4.31 ;
        RECT 5.955 4.14 6.125 4.31 ;
        RECT 6.415 4.14 6.585 4.31 ;
        RECT 6.875 4.14 7.045 4.31 ;
        RECT 7.06 4.55 7.23 4.72 ;
        RECT 7.335 4.14 7.505 4.31 ;
        RECT 7.795 4.14 7.965 4.31 ;
        RECT 8.255 4.14 8.425 4.31 ;
        RECT 8.715 4.14 8.885 4.31 ;
        RECT 9.175 4.14 9.345 4.31 ;
        RECT 12.675 4.55 12.845 4.72 ;
        RECT 12.675 4.17 12.845 4.34 ;
        RECT 13.375 4.555 13.545 4.725 ;
        RECT 13.375 4.165 13.545 4.335 ;
        RECT 14.365 4.555 14.535 4.725 ;
        RECT 14.365 4.165 14.535 4.335 ;
        RECT 16.155 4.14 16.325 4.31 ;
        RECT 16.615 4.14 16.785 4.31 ;
        RECT 17.075 4.14 17.245 4.31 ;
        RECT 17.535 4.14 17.705 4.31 ;
        RECT 17.995 4.14 18.165 4.31 ;
        RECT 18.455 4.14 18.625 4.31 ;
        RECT 18.915 4.14 19.085 4.31 ;
        RECT 19.375 4.14 19.545 4.31 ;
        RECT 19.835 4.14 20.005 4.31 ;
        RECT 20.295 4.14 20.465 4.31 ;
        RECT 20.755 4.14 20.925 4.31 ;
        RECT 21.215 4.14 21.385 4.31 ;
        RECT 21.675 4.14 21.845 4.31 ;
        RECT 22.135 4.14 22.305 4.31 ;
        RECT 22.32 4.55 22.49 4.72 ;
        RECT 22.595 4.14 22.765 4.31 ;
        RECT 23.055 4.14 23.225 4.31 ;
        RECT 23.515 4.14 23.685 4.31 ;
        RECT 23.975 4.14 24.145 4.31 ;
        RECT 24.435 4.14 24.605 4.31 ;
        RECT 27.935 4.55 28.105 4.72 ;
        RECT 27.935 4.17 28.105 4.34 ;
        RECT 28.635 4.555 28.805 4.725 ;
        RECT 28.635 4.165 28.805 4.335 ;
        RECT 29.625 4.555 29.795 4.725 ;
        RECT 29.625 4.165 29.795 4.335 ;
        RECT 31.415 4.14 31.585 4.31 ;
        RECT 31.875 4.14 32.045 4.31 ;
        RECT 32.335 4.14 32.505 4.31 ;
        RECT 32.795 4.14 32.965 4.31 ;
        RECT 33.255 4.14 33.425 4.31 ;
        RECT 33.715 4.14 33.885 4.31 ;
        RECT 34.175 4.14 34.345 4.31 ;
        RECT 34.635 4.14 34.805 4.31 ;
        RECT 35.095 4.14 35.265 4.31 ;
        RECT 35.555 4.14 35.725 4.31 ;
        RECT 36.015 4.14 36.185 4.31 ;
        RECT 36.475 4.14 36.645 4.31 ;
        RECT 36.935 4.14 37.105 4.31 ;
        RECT 37.395 4.14 37.565 4.31 ;
        RECT 37.58 4.55 37.75 4.72 ;
        RECT 37.855 4.14 38.025 4.31 ;
        RECT 38.315 4.14 38.485 4.31 ;
        RECT 38.775 4.14 38.945 4.31 ;
        RECT 39.235 4.14 39.405 4.31 ;
        RECT 39.695 4.14 39.865 4.31 ;
        RECT 43.195 4.55 43.365 4.72 ;
        RECT 43.195 4.17 43.365 4.34 ;
        RECT 43.895 4.555 44.065 4.725 ;
        RECT 43.895 4.165 44.065 4.335 ;
        RECT 44.885 4.555 45.055 4.725 ;
        RECT 44.885 4.165 45.055 4.335 ;
        RECT 46.675 4.14 46.845 4.31 ;
        RECT 47.135 4.14 47.305 4.31 ;
        RECT 47.595 4.14 47.765 4.31 ;
        RECT 48.055 4.14 48.225 4.31 ;
        RECT 48.515 4.14 48.685 4.31 ;
        RECT 48.975 4.14 49.145 4.31 ;
        RECT 49.435 4.14 49.605 4.31 ;
        RECT 49.895 4.14 50.065 4.31 ;
        RECT 50.355 4.14 50.525 4.31 ;
        RECT 50.815 4.14 50.985 4.31 ;
        RECT 51.275 4.14 51.445 4.31 ;
        RECT 51.735 4.14 51.905 4.31 ;
        RECT 52.195 4.14 52.365 4.31 ;
        RECT 52.655 4.14 52.825 4.31 ;
        RECT 52.84 4.55 53.01 4.72 ;
        RECT 53.115 4.14 53.285 4.31 ;
        RECT 53.575 4.14 53.745 4.31 ;
        RECT 54.035 4.14 54.205 4.31 ;
        RECT 54.495 4.14 54.665 4.31 ;
        RECT 54.955 4.14 55.125 4.31 ;
        RECT 58.455 4.55 58.625 4.72 ;
        RECT 58.455 4.17 58.625 4.34 ;
        RECT 59.155 4.555 59.325 4.725 ;
        RECT 59.155 4.165 59.325 4.335 ;
        RECT 60.145 4.555 60.315 4.725 ;
        RECT 60.145 4.165 60.315 4.335 ;
        RECT 61.935 4.14 62.105 4.31 ;
        RECT 62.395 4.14 62.565 4.31 ;
        RECT 62.855 4.14 63.025 4.31 ;
        RECT 63.315 4.14 63.485 4.31 ;
        RECT 63.775 4.14 63.945 4.31 ;
        RECT 64.235 4.14 64.405 4.31 ;
        RECT 64.695 4.14 64.865 4.31 ;
        RECT 65.155 4.14 65.325 4.31 ;
        RECT 65.615 4.14 65.785 4.31 ;
        RECT 66.075 4.14 66.245 4.31 ;
        RECT 66.535 4.14 66.705 4.31 ;
        RECT 66.995 4.14 67.165 4.31 ;
        RECT 67.455 4.14 67.625 4.31 ;
        RECT 67.915 4.14 68.085 4.31 ;
        RECT 68.1 4.55 68.27 4.72 ;
        RECT 68.375 4.14 68.545 4.31 ;
        RECT 68.835 4.14 69.005 4.31 ;
        RECT 69.295 4.14 69.465 4.31 ;
        RECT 69.755 4.14 69.925 4.31 ;
        RECT 70.215 4.14 70.385 4.31 ;
        RECT 73.715 4.55 73.885 4.72 ;
        RECT 73.715 4.17 73.885 4.34 ;
        RECT 74.415 4.555 74.585 4.725 ;
        RECT 74.415 4.165 74.585 4.335 ;
        RECT 75.405 4.555 75.575 4.725 ;
        RECT 75.405 4.165 75.575 4.335 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 62.62 1.86 63.35 2.19 ;
        RECT 47.36 1.86 48.09 2.19 ;
        RECT 32.1 1.86 32.83 2.19 ;
        RECT 16.84 1.86 17.57 2.19 ;
        RECT 1.58 1.86 2.31 2.19 ;
      LAYER met2 ;
        RECT 62.765 1.865 63.155 2.185 ;
        RECT 62.765 1.84 63.045 2.21 ;
        RECT 47.505 1.865 47.895 2.185 ;
        RECT 47.505 1.84 47.785 2.21 ;
        RECT 32.245 1.865 32.635 2.185 ;
        RECT 32.245 1.84 32.525 2.21 ;
        RECT 16.985 1.865 17.375 2.185 ;
        RECT 16.985 1.84 17.265 2.21 ;
        RECT 1.725 1.865 2.115 2.185 ;
        RECT 1.725 1.84 2.005 2.21 ;
      LAYER li1 ;
        RECT 76.12 0.005 76.3 0.31 ;
        RECT -2.75 0.005 76.3 0.305 ;
        RECT 75.325 0.005 75.495 0.935 ;
        RECT 74.335 0.005 74.505 0.935 ;
        RECT 60.86 0.005 74.17 0.31 ;
        RECT 71.595 0.005 71.765 0.94 ;
        RECT 61.79 0.005 70.53 1.59 ;
        RECT 69.76 0.005 69.93 2.09 ;
        RECT 68.82 0.005 68.99 2.09 ;
        RECT 67.86 0.005 68.03 2.09 ;
        RECT 66.815 0.005 67.01 1.6 ;
        RECT 65.94 0.005 66.11 2.09 ;
        RECT 64.98 0.005 65.15 2.09 ;
        RECT 63.06 0.005 63.335 1.6 ;
        RECT 63.06 0.005 63.23 2.09 ;
        RECT 60.065 0.005 60.235 0.935 ;
        RECT 59.075 0.005 59.245 0.935 ;
        RECT 45.6 0.005 58.91 0.31 ;
        RECT 56.335 0.005 56.505 0.94 ;
        RECT 46.53 0.005 55.27 1.59 ;
        RECT 54.5 0.005 54.67 2.09 ;
        RECT 53.56 0.005 53.73 2.09 ;
        RECT 52.6 0.005 52.77 2.09 ;
        RECT 51.555 0.005 51.75 1.6 ;
        RECT 50.68 0.005 50.85 2.09 ;
        RECT 49.72 0.005 49.89 2.09 ;
        RECT 47.8 0.005 48.075 1.6 ;
        RECT 47.8 0.005 47.97 2.09 ;
        RECT 44.805 0.005 44.975 0.935 ;
        RECT 43.815 0.005 43.985 0.935 ;
        RECT 30.34 0.005 43.65 0.31 ;
        RECT 41.075 0.005 41.245 0.94 ;
        RECT 31.27 0.005 40.01 1.59 ;
        RECT 39.24 0.005 39.41 2.09 ;
        RECT 38.3 0.005 38.47 2.09 ;
        RECT 37.34 0.005 37.51 2.09 ;
        RECT 36.295 0.005 36.49 1.6 ;
        RECT 35.42 0.005 35.59 2.09 ;
        RECT 34.46 0.005 34.63 2.09 ;
        RECT 32.54 0.005 32.815 1.6 ;
        RECT 32.54 0.005 32.71 2.09 ;
        RECT 29.545 0.005 29.715 0.935 ;
        RECT 28.555 0.005 28.725 0.935 ;
        RECT 15.08 0.005 28.39 0.31 ;
        RECT 25.815 0.005 25.985 0.94 ;
        RECT 16.01 0.005 24.75 1.59 ;
        RECT 23.98 0.005 24.15 2.09 ;
        RECT 23.04 0.005 23.21 2.09 ;
        RECT 22.08 0.005 22.25 2.09 ;
        RECT 21.035 0.005 21.23 1.6 ;
        RECT 20.16 0.005 20.33 2.09 ;
        RECT 19.2 0.005 19.37 2.09 ;
        RECT 17.28 0.005 17.555 1.6 ;
        RECT 17.28 0.005 17.45 2.09 ;
        RECT 14.285 0.005 14.455 0.935 ;
        RECT 13.295 0.005 13.465 0.935 ;
        RECT -2.75 0.005 13.13 0.31 ;
        RECT 10.555 0.005 10.725 0.94 ;
        RECT 0.75 0.005 9.49 1.59 ;
        RECT 8.72 0.005 8.89 2.09 ;
        RECT 7.78 0.005 7.95 2.09 ;
        RECT 6.82 0.005 6.99 2.09 ;
        RECT 5.775 0.005 5.97 1.6 ;
        RECT 4.9 0.005 5.07 2.09 ;
        RECT 3.94 0.005 4.11 2.09 ;
        RECT 2.02 0.005 2.295 1.6 ;
        RECT 2.02 0.005 2.19 2.09 ;
        RECT -2.75 8.585 76.3 8.885 ;
        RECT 76.12 8.58 76.3 8.885 ;
        RECT 75.325 7.955 75.495 8.885 ;
        RECT 74.335 7.955 74.505 8.885 ;
        RECT 60.86 8.58 74.17 8.885 ;
        RECT 71.595 7.95 71.765 8.885 ;
        RECT 65.98 7.95 66.15 8.885 ;
        RECT 60.065 7.955 60.235 8.885 ;
        RECT 59.075 7.955 59.245 8.885 ;
        RECT 45.6 8.58 58.91 8.885 ;
        RECT 56.335 7.95 56.505 8.885 ;
        RECT 50.72 7.95 50.89 8.885 ;
        RECT 44.805 7.955 44.975 8.885 ;
        RECT 43.815 7.955 43.985 8.885 ;
        RECT 30.34 8.58 43.65 8.885 ;
        RECT 41.075 7.95 41.245 8.885 ;
        RECT 35.46 7.95 35.63 8.885 ;
        RECT 29.545 7.955 29.715 8.885 ;
        RECT 28.555 7.955 28.725 8.885 ;
        RECT 15.08 8.58 28.39 8.885 ;
        RECT 25.815 7.95 25.985 8.885 ;
        RECT 20.2 7.95 20.37 8.885 ;
        RECT 14.285 7.955 14.455 8.885 ;
        RECT 13.295 7.955 13.465 8.885 ;
        RECT -2.75 8.58 13.13 8.885 ;
        RECT 10.555 7.95 10.725 8.885 ;
        RECT 4.94 7.95 5.11 8.885 ;
        RECT -2.575 7.95 -2.405 8.885 ;
        RECT 66.985 6.08 67.155 8.03 ;
        RECT 66.93 7.86 67.1 8.31 ;
        RECT 66.93 5.02 67.1 6.25 ;
        RECT 63.66 2.58 64.03 2.75 ;
        RECT 63.66 1.94 63.83 2.75 ;
        RECT 63.54 1.94 63.83 2.11 ;
        RECT 62.34 2.5 62.51 2.95 ;
        RECT 51.725 6.08 51.895 8.03 ;
        RECT 51.67 7.86 51.84 8.31 ;
        RECT 51.67 5.02 51.84 6.25 ;
        RECT 48.4 2.58 48.77 2.75 ;
        RECT 48.4 1.94 48.57 2.75 ;
        RECT 48.28 1.94 48.57 2.11 ;
        RECT 47.08 2.5 47.25 2.95 ;
        RECT 36.465 6.08 36.635 8.03 ;
        RECT 36.41 7.86 36.58 8.31 ;
        RECT 36.41 5.02 36.58 6.25 ;
        RECT 33.14 2.58 33.51 2.75 ;
        RECT 33.14 1.94 33.31 2.75 ;
        RECT 33.02 1.94 33.31 2.11 ;
        RECT 31.82 2.5 31.99 2.95 ;
        RECT 21.205 6.08 21.375 8.03 ;
        RECT 21.15 7.86 21.32 8.31 ;
        RECT 21.15 5.02 21.32 6.25 ;
        RECT 17.88 2.58 18.25 2.75 ;
        RECT 17.88 1.94 18.05 2.75 ;
        RECT 17.76 1.94 18.05 2.11 ;
        RECT 16.56 2.5 16.73 2.95 ;
        RECT 5.945 6.08 6.115 8.03 ;
        RECT 5.89 7.86 6.06 8.31 ;
        RECT 5.89 5.02 6.06 6.25 ;
        RECT 2.62 2.58 2.99 2.75 ;
        RECT 2.62 1.94 2.79 2.75 ;
        RECT 2.5 1.94 2.79 2.11 ;
        RECT 1.3 2.5 1.47 2.95 ;
      LAYER met1 ;
        RECT 76.12 0.005 76.3 0.31 ;
        RECT -2.75 0.005 76.3 0.305 ;
        RECT 60.86 0.005 74.17 0.31 ;
        RECT 61.79 0.005 70.53 1.745 ;
        RECT 63.48 1.91 63.77 2.14 ;
        RECT 62.595 1.955 63.77 2.095 ;
        RECT 62.775 1.895 63.185 2.155 ;
        RECT 62.775 0.005 63.065 2.155 ;
        RECT 62.355 2.375 62.975 2.515 ;
        RECT 62.835 0.005 62.975 2.515 ;
        RECT 62.595 1.955 62.975 2.215 ;
        RECT 62.28 2.75 62.57 2.98 ;
        RECT 62.355 2.375 62.495 2.98 ;
        RECT 45.6 0.005 58.91 0.31 ;
        RECT 46.53 0.005 55.27 1.745 ;
        RECT 48.22 1.91 48.51 2.14 ;
        RECT 47.335 1.955 48.51 2.095 ;
        RECT 47.515 1.895 47.925 2.155 ;
        RECT 47.515 0.005 47.805 2.155 ;
        RECT 47.095 2.375 47.715 2.515 ;
        RECT 47.575 0.005 47.715 2.515 ;
        RECT 47.335 1.955 47.715 2.215 ;
        RECT 47.02 2.75 47.31 2.98 ;
        RECT 47.095 2.375 47.235 2.98 ;
        RECT 30.34 0.005 43.65 0.31 ;
        RECT 31.27 0.005 40.01 1.745 ;
        RECT 32.96 1.91 33.25 2.14 ;
        RECT 32.075 1.955 33.25 2.095 ;
        RECT 32.255 1.895 32.665 2.155 ;
        RECT 32.255 0.005 32.545 2.155 ;
        RECT 31.835 2.375 32.455 2.515 ;
        RECT 32.315 0.005 32.455 2.515 ;
        RECT 32.075 1.955 32.455 2.215 ;
        RECT 31.76 2.75 32.05 2.98 ;
        RECT 31.835 2.375 31.975 2.98 ;
        RECT 15.08 0.005 28.39 0.31 ;
        RECT 16.01 0.005 24.75 1.745 ;
        RECT 17.7 1.91 17.99 2.14 ;
        RECT 16.815 1.955 17.99 2.095 ;
        RECT 16.995 1.895 17.405 2.155 ;
        RECT 16.995 0.005 17.285 2.155 ;
        RECT 16.575 2.375 17.195 2.515 ;
        RECT 17.055 0.005 17.195 2.515 ;
        RECT 16.815 1.955 17.195 2.215 ;
        RECT 16.5 2.75 16.79 2.98 ;
        RECT 16.575 2.375 16.715 2.98 ;
        RECT -2.75 0.005 13.13 0.31 ;
        RECT 0.75 0.005 9.49 1.745 ;
        RECT 2.44 1.91 2.73 2.14 ;
        RECT 1.555 1.955 2.73 2.095 ;
        RECT 1.735 1.895 2.145 2.155 ;
        RECT 1.735 0.005 2.025 2.155 ;
        RECT 1.315 2.375 1.935 2.515 ;
        RECT 1.795 0.005 1.935 2.515 ;
        RECT 1.555 1.955 1.935 2.215 ;
        RECT 1.24 2.75 1.53 2.98 ;
        RECT 1.315 2.375 1.455 2.98 ;
        RECT -2.75 8.585 76.3 8.885 ;
        RECT 76.12 8.58 76.3 8.885 ;
        RECT 60.86 8.58 74.17 8.885 ;
        RECT 66.925 6.29 67.215 6.52 ;
        RECT 66.76 6.32 66.93 8.885 ;
        RECT 66.755 6.32 67.215 6.49 ;
        RECT 45.6 8.58 58.91 8.885 ;
        RECT 51.665 6.29 51.955 6.52 ;
        RECT 51.5 6.32 51.67 8.885 ;
        RECT 51.495 6.32 51.955 6.49 ;
        RECT 30.34 8.58 43.65 8.885 ;
        RECT 36.405 6.29 36.695 6.52 ;
        RECT 36.24 6.32 36.41 8.885 ;
        RECT 36.235 6.32 36.695 6.49 ;
        RECT 15.08 8.58 28.39 8.885 ;
        RECT 21.145 6.29 21.435 6.52 ;
        RECT 20.98 6.32 21.15 8.885 ;
        RECT 20.975 6.32 21.435 6.49 ;
        RECT -2.75 8.58 13.13 8.885 ;
        RECT 5.885 6.29 6.175 6.52 ;
        RECT 5.72 6.32 5.89 8.885 ;
        RECT 5.715 6.32 6.175 6.49 ;
      LAYER via2 ;
        RECT 1.765 1.925 1.965 2.125 ;
        RECT 17.025 1.925 17.225 2.125 ;
        RECT 32.285 1.925 32.485 2.125 ;
        RECT 47.545 1.925 47.745 2.125 ;
        RECT 62.805 1.925 63.005 2.125 ;
      LAYER via1 ;
        RECT 1.91 1.95 2.06 2.1 ;
        RECT 17.17 1.95 17.32 2.1 ;
        RECT 32.43 1.95 32.58 2.1 ;
        RECT 47.69 1.95 47.84 2.1 ;
        RECT 62.95 1.95 63.1 2.1 ;
      LAYER mcon ;
        RECT -2.495 8.61 -2.325 8.78 ;
        RECT -1.815 8.61 -1.645 8.78 ;
        RECT -1.135 8.61 -0.965 8.78 ;
        RECT -0.455 8.61 -0.285 8.78 ;
        RECT 0.895 1.42 1.065 1.59 ;
        RECT 1.3 2.78 1.47 2.95 ;
        RECT 1.355 1.42 1.525 1.59 ;
        RECT 1.815 1.42 1.985 1.59 ;
        RECT 2.275 1.42 2.445 1.59 ;
        RECT 2.5 1.94 2.67 2.11 ;
        RECT 2.735 1.42 2.905 1.59 ;
        RECT 3.195 1.42 3.365 1.59 ;
        RECT 3.655 1.42 3.825 1.59 ;
        RECT 4.115 1.42 4.285 1.59 ;
        RECT 4.575 1.42 4.745 1.59 ;
        RECT 5.02 8.61 5.19 8.78 ;
        RECT 5.035 1.42 5.205 1.59 ;
        RECT 5.495 1.42 5.665 1.59 ;
        RECT 5.7 8.61 5.87 8.78 ;
        RECT 5.945 6.32 6.115 6.49 ;
        RECT 5.955 1.42 6.125 1.59 ;
        RECT 6.38 8.61 6.55 8.78 ;
        RECT 6.415 1.42 6.585 1.59 ;
        RECT 6.875 1.42 7.045 1.59 ;
        RECT 7.06 8.61 7.23 8.78 ;
        RECT 7.335 1.42 7.505 1.59 ;
        RECT 7.795 1.42 7.965 1.59 ;
        RECT 8.255 1.42 8.425 1.59 ;
        RECT 8.715 1.42 8.885 1.59 ;
        RECT 9.175 1.42 9.345 1.59 ;
        RECT 10.635 8.61 10.805 8.78 ;
        RECT 10.635 0.11 10.805 0.28 ;
        RECT 11.315 8.61 11.485 8.78 ;
        RECT 11.315 0.11 11.485 0.28 ;
        RECT 11.995 8.61 12.165 8.78 ;
        RECT 11.995 0.11 12.165 0.28 ;
        RECT 12.675 8.61 12.845 8.78 ;
        RECT 12.675 0.11 12.845 0.28 ;
        RECT 13.375 8.615 13.545 8.785 ;
        RECT 13.375 0.105 13.545 0.275 ;
        RECT 14.365 8.615 14.535 8.785 ;
        RECT 14.365 0.105 14.535 0.275 ;
        RECT 16.155 1.42 16.325 1.59 ;
        RECT 16.56 2.78 16.73 2.95 ;
        RECT 16.615 1.42 16.785 1.59 ;
        RECT 17.075 1.42 17.245 1.59 ;
        RECT 17.535 1.42 17.705 1.59 ;
        RECT 17.76 1.94 17.93 2.11 ;
        RECT 17.995 1.42 18.165 1.59 ;
        RECT 18.455 1.42 18.625 1.59 ;
        RECT 18.915 1.42 19.085 1.59 ;
        RECT 19.375 1.42 19.545 1.59 ;
        RECT 19.835 1.42 20.005 1.59 ;
        RECT 20.28 8.61 20.45 8.78 ;
        RECT 20.295 1.42 20.465 1.59 ;
        RECT 20.755 1.42 20.925 1.59 ;
        RECT 20.96 8.61 21.13 8.78 ;
        RECT 21.205 6.32 21.375 6.49 ;
        RECT 21.215 1.42 21.385 1.59 ;
        RECT 21.64 8.61 21.81 8.78 ;
        RECT 21.675 1.42 21.845 1.59 ;
        RECT 22.135 1.42 22.305 1.59 ;
        RECT 22.32 8.61 22.49 8.78 ;
        RECT 22.595 1.42 22.765 1.59 ;
        RECT 23.055 1.42 23.225 1.59 ;
        RECT 23.515 1.42 23.685 1.59 ;
        RECT 23.975 1.42 24.145 1.59 ;
        RECT 24.435 1.42 24.605 1.59 ;
        RECT 25.895 8.61 26.065 8.78 ;
        RECT 25.895 0.11 26.065 0.28 ;
        RECT 26.575 8.61 26.745 8.78 ;
        RECT 26.575 0.11 26.745 0.28 ;
        RECT 27.255 8.61 27.425 8.78 ;
        RECT 27.255 0.11 27.425 0.28 ;
        RECT 27.935 8.61 28.105 8.78 ;
        RECT 27.935 0.11 28.105 0.28 ;
        RECT 28.635 8.615 28.805 8.785 ;
        RECT 28.635 0.105 28.805 0.275 ;
        RECT 29.625 8.615 29.795 8.785 ;
        RECT 29.625 0.105 29.795 0.275 ;
        RECT 31.415 1.42 31.585 1.59 ;
        RECT 31.82 2.78 31.99 2.95 ;
        RECT 31.875 1.42 32.045 1.59 ;
        RECT 32.335 1.42 32.505 1.59 ;
        RECT 32.795 1.42 32.965 1.59 ;
        RECT 33.02 1.94 33.19 2.11 ;
        RECT 33.255 1.42 33.425 1.59 ;
        RECT 33.715 1.42 33.885 1.59 ;
        RECT 34.175 1.42 34.345 1.59 ;
        RECT 34.635 1.42 34.805 1.59 ;
        RECT 35.095 1.42 35.265 1.59 ;
        RECT 35.54 8.61 35.71 8.78 ;
        RECT 35.555 1.42 35.725 1.59 ;
        RECT 36.015 1.42 36.185 1.59 ;
        RECT 36.22 8.61 36.39 8.78 ;
        RECT 36.465 6.32 36.635 6.49 ;
        RECT 36.475 1.42 36.645 1.59 ;
        RECT 36.9 8.61 37.07 8.78 ;
        RECT 36.935 1.42 37.105 1.59 ;
        RECT 37.395 1.42 37.565 1.59 ;
        RECT 37.58 8.61 37.75 8.78 ;
        RECT 37.855 1.42 38.025 1.59 ;
        RECT 38.315 1.42 38.485 1.59 ;
        RECT 38.775 1.42 38.945 1.59 ;
        RECT 39.235 1.42 39.405 1.59 ;
        RECT 39.695 1.42 39.865 1.59 ;
        RECT 41.155 8.61 41.325 8.78 ;
        RECT 41.155 0.11 41.325 0.28 ;
        RECT 41.835 8.61 42.005 8.78 ;
        RECT 41.835 0.11 42.005 0.28 ;
        RECT 42.515 8.61 42.685 8.78 ;
        RECT 42.515 0.11 42.685 0.28 ;
        RECT 43.195 8.61 43.365 8.78 ;
        RECT 43.195 0.11 43.365 0.28 ;
        RECT 43.895 8.615 44.065 8.785 ;
        RECT 43.895 0.105 44.065 0.275 ;
        RECT 44.885 8.615 45.055 8.785 ;
        RECT 44.885 0.105 45.055 0.275 ;
        RECT 46.675 1.42 46.845 1.59 ;
        RECT 47.08 2.78 47.25 2.95 ;
        RECT 47.135 1.42 47.305 1.59 ;
        RECT 47.595 1.42 47.765 1.59 ;
        RECT 48.055 1.42 48.225 1.59 ;
        RECT 48.28 1.94 48.45 2.11 ;
        RECT 48.515 1.42 48.685 1.59 ;
        RECT 48.975 1.42 49.145 1.59 ;
        RECT 49.435 1.42 49.605 1.59 ;
        RECT 49.895 1.42 50.065 1.59 ;
        RECT 50.355 1.42 50.525 1.59 ;
        RECT 50.8 8.61 50.97 8.78 ;
        RECT 50.815 1.42 50.985 1.59 ;
        RECT 51.275 1.42 51.445 1.59 ;
        RECT 51.48 8.61 51.65 8.78 ;
        RECT 51.725 6.32 51.895 6.49 ;
        RECT 51.735 1.42 51.905 1.59 ;
        RECT 52.16 8.61 52.33 8.78 ;
        RECT 52.195 1.42 52.365 1.59 ;
        RECT 52.655 1.42 52.825 1.59 ;
        RECT 52.84 8.61 53.01 8.78 ;
        RECT 53.115 1.42 53.285 1.59 ;
        RECT 53.575 1.42 53.745 1.59 ;
        RECT 54.035 1.42 54.205 1.59 ;
        RECT 54.495 1.42 54.665 1.59 ;
        RECT 54.955 1.42 55.125 1.59 ;
        RECT 56.415 8.61 56.585 8.78 ;
        RECT 56.415 0.11 56.585 0.28 ;
        RECT 57.095 8.61 57.265 8.78 ;
        RECT 57.095 0.11 57.265 0.28 ;
        RECT 57.775 8.61 57.945 8.78 ;
        RECT 57.775 0.11 57.945 0.28 ;
        RECT 58.455 8.61 58.625 8.78 ;
        RECT 58.455 0.11 58.625 0.28 ;
        RECT 59.155 8.615 59.325 8.785 ;
        RECT 59.155 0.105 59.325 0.275 ;
        RECT 60.145 8.615 60.315 8.785 ;
        RECT 60.145 0.105 60.315 0.275 ;
        RECT 61.935 1.42 62.105 1.59 ;
        RECT 62.34 2.78 62.51 2.95 ;
        RECT 62.395 1.42 62.565 1.59 ;
        RECT 62.855 1.42 63.025 1.59 ;
        RECT 63.315 1.42 63.485 1.59 ;
        RECT 63.54 1.94 63.71 2.11 ;
        RECT 63.775 1.42 63.945 1.59 ;
        RECT 64.235 1.42 64.405 1.59 ;
        RECT 64.695 1.42 64.865 1.59 ;
        RECT 65.155 1.42 65.325 1.59 ;
        RECT 65.615 1.42 65.785 1.59 ;
        RECT 66.06 8.61 66.23 8.78 ;
        RECT 66.075 1.42 66.245 1.59 ;
        RECT 66.535 1.42 66.705 1.59 ;
        RECT 66.74 8.61 66.91 8.78 ;
        RECT 66.985 6.32 67.155 6.49 ;
        RECT 66.995 1.42 67.165 1.59 ;
        RECT 67.42 8.61 67.59 8.78 ;
        RECT 67.455 1.42 67.625 1.59 ;
        RECT 67.915 1.42 68.085 1.59 ;
        RECT 68.1 8.61 68.27 8.78 ;
        RECT 68.375 1.42 68.545 1.59 ;
        RECT 68.835 1.42 69.005 1.59 ;
        RECT 69.295 1.42 69.465 1.59 ;
        RECT 69.755 1.42 69.925 1.59 ;
        RECT 70.215 1.42 70.385 1.59 ;
        RECT 71.675 8.61 71.845 8.78 ;
        RECT 71.675 0.11 71.845 0.28 ;
        RECT 72.355 8.61 72.525 8.78 ;
        RECT 72.355 0.11 72.525 0.28 ;
        RECT 73.035 8.61 73.205 8.78 ;
        RECT 73.035 0.11 73.205 0.28 ;
        RECT 73.715 8.61 73.885 8.78 ;
        RECT 73.715 0.11 73.885 0.28 ;
        RECT 74.415 8.615 74.585 8.785 ;
        RECT 74.415 0.105 74.585 0.275 ;
        RECT 75.405 8.615 75.575 8.785 ;
        RECT 75.405 0.105 75.575 0.275 ;
    END
  END vssd1
  OBS
    LAYER met4 ;
      RECT 63.94 2.98 64.27 3.31 ;
      RECT 63.955 2.505 64.27 3.31 ;
      RECT 66.1 2.49 66.43 2.845 ;
      RECT 63.955 2.505 66.43 2.805 ;
      RECT 48.68 2.98 49.01 3.31 ;
      RECT 48.695 2.505 49.01 3.31 ;
      RECT 50.84 2.49 51.17 2.845 ;
      RECT 48.695 2.505 51.17 2.805 ;
      RECT 33.42 2.98 33.75 3.31 ;
      RECT 33.435 2.505 33.75 3.31 ;
      RECT 35.58 2.49 35.91 2.845 ;
      RECT 33.435 2.505 35.91 2.805 ;
      RECT 18.16 2.98 18.49 3.31 ;
      RECT 18.175 2.505 18.49 3.31 ;
      RECT 20.32 2.49 20.65 2.845 ;
      RECT 18.175 2.505 20.65 2.805 ;
      RECT 2.9 2.98 3.23 3.31 ;
      RECT 2.915 2.505 3.23 3.31 ;
      RECT 5.06 2.49 5.39 2.845 ;
      RECT 2.915 2.505 5.39 2.805 ;
    LAYER via3 ;
      RECT 66.165 2.58 66.365 2.78 ;
      RECT 64.005 3.045 64.205 3.245 ;
      RECT 50.905 2.58 51.105 2.78 ;
      RECT 48.745 3.045 48.945 3.245 ;
      RECT 35.645 2.58 35.845 2.78 ;
      RECT 33.485 3.045 33.685 3.245 ;
      RECT 20.385 2.58 20.585 2.78 ;
      RECT 18.225 3.045 18.425 3.245 ;
      RECT 5.125 2.58 5.325 2.78 ;
      RECT 2.965 3.045 3.165 3.245 ;
    LAYER met3 ;
      RECT 67.26 7.06 67.63 7.43 ;
      RECT 67.295 4.48 67.595 7.43 ;
      RECT 65.855 4.48 67.595 4.78 ;
      RECT 63.06 4.26 66.155 4.56 ;
      RECT 65.855 2.52 66.155 4.78 ;
      RECT 63.06 2.98 63.36 4.56 ;
      RECT 66.58 3.515 66.91 3.87 ;
      RECT 64.675 3.555 66.91 3.855 ;
      RECT 64.675 2.42 64.975 3.855 ;
      RECT 62.755 2.98 63.485 3.31 ;
      RECT 65.65 2.525 66.43 2.87 ;
      RECT 66.125 2.49 66.43 2.87 ;
      RECT 64.66 2.42 64.99 2.75 ;
      RECT 63.945 2.42 64.265 3.335 ;
      RECT 63.945 2.42 64.275 2.955 ;
      RECT 52 7.06 52.37 7.43 ;
      RECT 52.035 4.48 52.335 7.43 ;
      RECT 50.595 4.48 52.335 4.78 ;
      RECT 47.8 4.26 50.895 4.56 ;
      RECT 50.595 2.52 50.895 4.78 ;
      RECT 47.8 2.98 48.1 4.56 ;
      RECT 51.32 3.515 51.65 3.87 ;
      RECT 49.415 3.555 51.65 3.855 ;
      RECT 49.415 2.42 49.715 3.855 ;
      RECT 47.495 2.98 48.225 3.31 ;
      RECT 50.39 2.525 51.17 2.87 ;
      RECT 50.865 2.49 51.17 2.87 ;
      RECT 49.4 2.42 49.73 2.75 ;
      RECT 48.685 2.42 49.005 3.335 ;
      RECT 48.685 2.42 49.015 2.955 ;
      RECT 36.74 7.06 37.11 7.43 ;
      RECT 36.775 4.48 37.075 7.43 ;
      RECT 35.335 4.48 37.075 4.78 ;
      RECT 32.54 4.26 35.635 4.56 ;
      RECT 35.335 2.52 35.635 4.78 ;
      RECT 32.54 2.98 32.84 4.56 ;
      RECT 36.06 3.515 36.39 3.87 ;
      RECT 34.155 3.555 36.39 3.855 ;
      RECT 34.155 2.42 34.455 3.855 ;
      RECT 32.235 2.98 32.965 3.31 ;
      RECT 35.13 2.525 35.91 2.87 ;
      RECT 35.605 2.49 35.91 2.87 ;
      RECT 34.14 2.42 34.47 2.75 ;
      RECT 33.425 2.42 33.745 3.335 ;
      RECT 33.425 2.42 33.755 2.955 ;
      RECT 21.48 7.06 21.85 7.43 ;
      RECT 21.515 4.48 21.815 7.43 ;
      RECT 20.075 4.48 21.815 4.78 ;
      RECT 17.28 4.26 20.375 4.56 ;
      RECT 20.075 2.52 20.375 4.78 ;
      RECT 17.28 2.98 17.58 4.56 ;
      RECT 20.8 3.515 21.13 3.87 ;
      RECT 18.895 3.555 21.13 3.855 ;
      RECT 18.895 2.42 19.195 3.855 ;
      RECT 16.975 2.98 17.705 3.31 ;
      RECT 19.87 2.525 20.65 2.87 ;
      RECT 20.345 2.49 20.65 2.87 ;
      RECT 18.88 2.42 19.21 2.75 ;
      RECT 18.165 2.42 18.485 3.335 ;
      RECT 18.165 2.42 18.495 2.955 ;
      RECT 6.22 7.06 6.59 7.43 ;
      RECT 6.255 4.48 6.555 7.43 ;
      RECT 4.815 4.48 6.555 4.78 ;
      RECT 2.02 4.26 5.115 4.56 ;
      RECT 4.815 2.52 5.115 4.78 ;
      RECT 2.02 2.98 2.32 4.56 ;
      RECT 5.54 3.515 5.87 3.87 ;
      RECT 3.635 3.555 5.87 3.855 ;
      RECT 3.635 2.42 3.935 3.855 ;
      RECT 1.715 2.98 2.445 3.31 ;
      RECT 4.61 2.525 5.39 2.87 ;
      RECT 5.085 2.49 5.39 2.87 ;
      RECT 3.62 2.42 3.95 2.75 ;
      RECT 2.905 2.42 3.225 3.335 ;
      RECT 2.905 2.42 3.235 2.955 ;
      RECT 69.5 1.86 70.23 2.19 ;
      RECT 67.81 1.875 68.54 2.205 ;
      RECT 66.775 1.86 67.505 2.21 ;
      RECT 65.225 1.885 65.955 2.215 ;
      RECT 54.24 1.86 54.97 2.19 ;
      RECT 52.55 1.875 53.28 2.205 ;
      RECT 51.515 1.86 52.245 2.21 ;
      RECT 49.965 1.885 50.695 2.215 ;
      RECT 38.98 1.86 39.71 2.19 ;
      RECT 37.29 1.875 38.02 2.205 ;
      RECT 36.255 1.86 36.985 2.21 ;
      RECT 34.705 1.885 35.435 2.215 ;
      RECT 23.72 1.86 24.45 2.19 ;
      RECT 22.03 1.875 22.76 2.205 ;
      RECT 20.995 1.86 21.725 2.21 ;
      RECT 19.445 1.885 20.175 2.215 ;
      RECT 8.46 1.86 9.19 2.19 ;
      RECT 6.77 1.875 7.5 2.205 ;
      RECT 5.735 1.86 6.465 2.21 ;
      RECT 4.185 1.885 4.915 2.215 ;
    LAYER via2 ;
      RECT 69.735 1.925 69.935 2.125 ;
      RECT 67.875 1.94 68.075 2.14 ;
      RECT 67.345 7.145 67.545 7.345 ;
      RECT 66.855 1.945 67.055 2.145 ;
      RECT 66.645 3.58 66.845 3.78 ;
      RECT 66.165 2.58 66.365 2.78 ;
      RECT 65.415 1.95 65.615 2.15 ;
      RECT 64.725 2.485 64.925 2.685 ;
      RECT 64.01 2.485 64.21 2.685 ;
      RECT 63.045 3.045 63.245 3.245 ;
      RECT 54.475 1.925 54.675 2.125 ;
      RECT 52.615 1.94 52.815 2.14 ;
      RECT 52.085 7.145 52.285 7.345 ;
      RECT 51.595 1.945 51.795 2.145 ;
      RECT 51.385 3.58 51.585 3.78 ;
      RECT 50.905 2.58 51.105 2.78 ;
      RECT 50.155 1.95 50.355 2.15 ;
      RECT 49.465 2.485 49.665 2.685 ;
      RECT 48.75 2.485 48.95 2.685 ;
      RECT 47.785 3.045 47.985 3.245 ;
      RECT 39.215 1.925 39.415 2.125 ;
      RECT 37.355 1.94 37.555 2.14 ;
      RECT 36.825 7.145 37.025 7.345 ;
      RECT 36.335 1.945 36.535 2.145 ;
      RECT 36.125 3.58 36.325 3.78 ;
      RECT 35.645 2.58 35.845 2.78 ;
      RECT 34.895 1.95 35.095 2.15 ;
      RECT 34.205 2.485 34.405 2.685 ;
      RECT 33.49 2.485 33.69 2.685 ;
      RECT 32.525 3.045 32.725 3.245 ;
      RECT 23.955 1.925 24.155 2.125 ;
      RECT 22.095 1.94 22.295 2.14 ;
      RECT 21.565 7.145 21.765 7.345 ;
      RECT 21.075 1.945 21.275 2.145 ;
      RECT 20.865 3.58 21.065 3.78 ;
      RECT 20.385 2.58 20.585 2.78 ;
      RECT 19.635 1.95 19.835 2.15 ;
      RECT 18.945 2.485 19.145 2.685 ;
      RECT 18.23 2.485 18.43 2.685 ;
      RECT 17.265 3.045 17.465 3.245 ;
      RECT 8.695 1.925 8.895 2.125 ;
      RECT 6.835 1.94 7.035 2.14 ;
      RECT 6.305 7.145 6.505 7.345 ;
      RECT 5.815 1.945 6.015 2.145 ;
      RECT 5.605 3.58 5.805 3.78 ;
      RECT 5.125 2.58 5.325 2.78 ;
      RECT 4.375 1.95 4.575 2.15 ;
      RECT 3.685 2.485 3.885 2.685 ;
      RECT 2.97 2.485 3.17 2.685 ;
      RECT 2.005 3.045 2.205 3.245 ;
    LAYER met2 ;
      RECT -1.57 8.405 75.93 8.575 ;
      RECT 75.76 7.28 75.93 8.575 ;
      RECT -1.57 6.26 -1.4 8.575 ;
      RECT 75.73 7.28 76.08 7.63 ;
      RECT -1.63 6.26 -1.34 6.61 ;
      RECT 72.57 6.225 72.89 6.55 ;
      RECT 72.6 5.7 72.77 6.55 ;
      RECT 72.6 5.7 72.775 6.05 ;
      RECT 72.6 5.7 73.575 5.875 ;
      RECT 73.4 1.97 73.575 5.875 ;
      RECT 73.345 1.97 73.695 2.32 ;
      RECT 73.37 6.66 73.695 6.985 ;
      RECT 72.255 6.75 73.695 6.92 ;
      RECT 72.255 2.4 72.415 6.92 ;
      RECT 72.57 2.37 72.89 2.69 ;
      RECT 72.255 2.4 72.89 2.57 ;
      RECT 69.705 3.545 69.965 3.865 ;
      RECT 69.765 1.84 69.905 3.865 ;
      RECT 70.965 2.705 71.305 3.055 ;
      RECT 70.34 2.775 71.305 2.975 ;
      RECT 70.34 1.945 70.54 2.975 ;
      RECT 69.59 2.4 69.905 2.77 ;
      RECT 71.055 2.7 71.225 3.055 ;
      RECT 69.66 1.955 69.905 2.77 ;
      RECT 69.695 1.84 69.975 2.21 ;
      RECT 69.695 1.945 70.54 2.145 ;
      RECT 69.015 2.425 69.275 2.745 ;
      RECT 68.355 2.515 69.275 2.655 ;
      RECT 68.355 1.575 68.495 2.655 ;
      RECT 64.815 1.865 65.075 2.185 ;
      RECT 64.995 1.575 65.135 2.095 ;
      RECT 64.995 1.575 68.495 1.715 ;
      RECT 60.445 6.66 60.795 7.01 ;
      RECT 67.93 6.615 68.28 6.965 ;
      RECT 60.445 6.69 68.28 6.89 ;
      RECT 67.845 3.265 68.105 3.585 ;
      RECT 67.905 1.855 68.045 3.585 ;
      RECT 67.835 1.855 68.115 2.225 ;
      RECT 65.235 4.015 67.67 4.155 ;
      RECT 67.53 2.705 67.67 4.155 ;
      RECT 65.235 3.635 65.375 4.155 ;
      RECT 64.935 3.635 65.375 3.865 ;
      RECT 62.595 3.635 65.375 3.775 ;
      RECT 64.935 3.545 65.195 3.865 ;
      RECT 62.595 3.355 62.735 3.775 ;
      RECT 62.085 3.265 62.345 3.585 ;
      RECT 62.085 3.355 62.735 3.495 ;
      RECT 62.145 1.865 62.285 3.585 ;
      RECT 67.47 2.705 67.73 3.025 ;
      RECT 62.085 1.865 62.345 2.185 ;
      RECT 67.095 3.545 67.355 3.865 ;
      RECT 67.155 1.955 67.295 3.865 ;
      RECT 66.815 1.955 67.295 2.23 ;
      RECT 66.615 1.86 67.095 2.205 ;
      RECT 66.605 3.495 66.885 3.865 ;
      RECT 66.675 2.4 66.815 3.865 ;
      RECT 66.615 2.4 66.875 3.025 ;
      RECT 66.605 2.4 66.885 2.77 ;
      RECT 65.535 3.545 65.795 3.865 ;
      RECT 65.535 3.355 65.735 3.865 ;
      RECT 65.34 3.355 65.735 3.495 ;
      RECT 65.34 1.865 65.48 3.495 ;
      RECT 65.34 1.865 65.655 2.235 ;
      RECT 65.28 1.865 65.655 2.185 ;
      RECT 63.005 2.96 63.285 3.33 ;
      RECT 64.455 2.985 64.715 3.305 ;
      RECT 62.835 3.075 64.715 3.215 ;
      RECT 62.835 2.96 63.285 3.215 ;
      RECT 62.775 2.4 63.035 3.025 ;
      RECT 62.765 2.4 63.045 2.77 ;
      RECT 63.845 2.4 64.255 2.77 ;
      RECT 63.255 2.425 63.515 2.745 ;
      RECT 63.255 2.515 64.255 2.655 ;
      RECT 57.31 6.225 57.63 6.55 ;
      RECT 57.34 5.7 57.51 6.55 ;
      RECT 57.34 5.7 57.515 6.05 ;
      RECT 57.34 5.7 58.315 5.875 ;
      RECT 58.14 1.97 58.315 5.875 ;
      RECT 58.085 1.97 58.435 2.32 ;
      RECT 58.11 6.66 58.435 6.985 ;
      RECT 56.995 6.75 58.435 6.92 ;
      RECT 56.995 2.4 57.155 6.92 ;
      RECT 57.31 2.37 57.63 2.69 ;
      RECT 56.995 2.4 57.63 2.57 ;
      RECT 54.445 3.545 54.705 3.865 ;
      RECT 54.505 1.84 54.645 3.865 ;
      RECT 55.705 2.705 56.045 3.055 ;
      RECT 55.08 2.775 56.045 2.975 ;
      RECT 55.08 1.945 55.28 2.975 ;
      RECT 54.33 2.4 54.645 2.77 ;
      RECT 55.795 2.7 55.965 3.055 ;
      RECT 54.4 1.955 54.645 2.77 ;
      RECT 54.435 1.84 54.715 2.21 ;
      RECT 54.435 1.945 55.28 2.145 ;
      RECT 53.755 2.425 54.015 2.745 ;
      RECT 53.095 2.515 54.015 2.655 ;
      RECT 53.095 1.575 53.235 2.655 ;
      RECT 49.555 1.865 49.815 2.185 ;
      RECT 49.735 1.575 49.875 2.095 ;
      RECT 49.735 1.575 53.235 1.715 ;
      RECT 45.185 6.66 45.535 7.01 ;
      RECT 52.675 6.615 53.025 6.965 ;
      RECT 45.185 6.69 53.025 6.89 ;
      RECT 52.585 3.265 52.845 3.585 ;
      RECT 52.645 1.855 52.785 3.585 ;
      RECT 52.575 1.855 52.855 2.225 ;
      RECT 49.975 4.015 52.41 4.155 ;
      RECT 52.27 2.705 52.41 4.155 ;
      RECT 49.975 3.635 50.115 4.155 ;
      RECT 49.675 3.635 50.115 3.865 ;
      RECT 47.335 3.635 50.115 3.775 ;
      RECT 49.675 3.545 49.935 3.865 ;
      RECT 47.335 3.355 47.475 3.775 ;
      RECT 46.825 3.265 47.085 3.585 ;
      RECT 46.825 3.355 47.475 3.495 ;
      RECT 46.885 1.865 47.025 3.585 ;
      RECT 52.21 2.705 52.47 3.025 ;
      RECT 46.825 1.865 47.085 2.185 ;
      RECT 51.835 3.545 52.095 3.865 ;
      RECT 51.895 1.955 52.035 3.865 ;
      RECT 51.555 1.955 52.035 2.23 ;
      RECT 51.355 1.86 51.835 2.205 ;
      RECT 51.345 3.495 51.625 3.865 ;
      RECT 51.415 2.4 51.555 3.865 ;
      RECT 51.355 2.4 51.615 3.025 ;
      RECT 51.345 2.4 51.625 2.77 ;
      RECT 50.275 3.545 50.535 3.865 ;
      RECT 50.275 3.355 50.475 3.865 ;
      RECT 50.08 3.355 50.475 3.495 ;
      RECT 50.08 1.865 50.22 3.495 ;
      RECT 50.08 1.865 50.395 2.235 ;
      RECT 50.02 1.865 50.395 2.185 ;
      RECT 47.745 2.96 48.025 3.33 ;
      RECT 49.195 2.985 49.455 3.305 ;
      RECT 47.575 3.075 49.455 3.215 ;
      RECT 47.575 2.96 48.025 3.215 ;
      RECT 47.515 2.4 47.775 3.025 ;
      RECT 47.505 2.4 47.785 2.77 ;
      RECT 48.585 2.4 48.995 2.77 ;
      RECT 47.995 2.425 48.255 2.745 ;
      RECT 47.995 2.515 48.995 2.655 ;
      RECT 42.05 6.225 42.37 6.55 ;
      RECT 42.08 5.7 42.25 6.55 ;
      RECT 42.08 5.7 42.255 6.05 ;
      RECT 42.08 5.7 43.055 5.875 ;
      RECT 42.88 1.97 43.055 5.875 ;
      RECT 42.825 1.97 43.175 2.32 ;
      RECT 42.85 6.66 43.175 6.985 ;
      RECT 41.735 6.75 43.175 6.92 ;
      RECT 41.735 2.4 41.895 6.92 ;
      RECT 42.05 2.37 42.37 2.69 ;
      RECT 41.735 2.4 42.37 2.57 ;
      RECT 39.185 3.545 39.445 3.865 ;
      RECT 39.245 1.84 39.385 3.865 ;
      RECT 40.445 2.705 40.785 3.055 ;
      RECT 39.82 2.775 40.785 2.975 ;
      RECT 39.82 1.945 40.02 2.975 ;
      RECT 39.07 2.4 39.385 2.77 ;
      RECT 40.535 2.7 40.705 3.055 ;
      RECT 39.14 1.955 39.385 2.77 ;
      RECT 39.175 1.84 39.455 2.21 ;
      RECT 39.175 1.945 40.02 2.145 ;
      RECT 38.495 2.425 38.755 2.745 ;
      RECT 37.835 2.515 38.755 2.655 ;
      RECT 37.835 1.575 37.975 2.655 ;
      RECT 34.295 1.865 34.555 2.185 ;
      RECT 34.475 1.575 34.615 2.095 ;
      RECT 34.475 1.575 37.975 1.715 ;
      RECT 29.97 6.665 30.32 7.015 ;
      RECT 37.41 6.62 37.76 6.97 ;
      RECT 29.97 6.695 37.76 6.895 ;
      RECT 37.325 3.265 37.585 3.585 ;
      RECT 37.385 1.855 37.525 3.585 ;
      RECT 37.315 1.855 37.595 2.225 ;
      RECT 34.715 4.015 37.15 4.155 ;
      RECT 37.01 2.705 37.15 4.155 ;
      RECT 34.715 3.635 34.855 4.155 ;
      RECT 34.415 3.635 34.855 3.865 ;
      RECT 32.075 3.635 34.855 3.775 ;
      RECT 34.415 3.545 34.675 3.865 ;
      RECT 32.075 3.355 32.215 3.775 ;
      RECT 31.565 3.265 31.825 3.585 ;
      RECT 31.565 3.355 32.215 3.495 ;
      RECT 31.625 1.865 31.765 3.585 ;
      RECT 36.95 2.705 37.21 3.025 ;
      RECT 31.565 1.865 31.825 2.185 ;
      RECT 36.575 3.545 36.835 3.865 ;
      RECT 36.635 1.955 36.775 3.865 ;
      RECT 36.295 1.955 36.775 2.23 ;
      RECT 36.095 1.86 36.575 2.205 ;
      RECT 36.085 3.495 36.365 3.865 ;
      RECT 36.155 2.4 36.295 3.865 ;
      RECT 36.095 2.4 36.355 3.025 ;
      RECT 36.085 2.4 36.365 2.77 ;
      RECT 35.015 3.545 35.275 3.865 ;
      RECT 35.015 3.355 35.215 3.865 ;
      RECT 34.82 3.355 35.215 3.495 ;
      RECT 34.82 1.865 34.96 3.495 ;
      RECT 34.82 1.865 35.135 2.235 ;
      RECT 34.76 1.865 35.135 2.185 ;
      RECT 32.485 2.96 32.765 3.33 ;
      RECT 33.935 2.985 34.195 3.305 ;
      RECT 32.315 3.075 34.195 3.215 ;
      RECT 32.315 2.96 32.765 3.215 ;
      RECT 32.255 2.4 32.515 3.025 ;
      RECT 32.245 2.4 32.525 2.77 ;
      RECT 33.325 2.4 33.735 2.77 ;
      RECT 32.735 2.425 32.995 2.745 ;
      RECT 32.735 2.515 33.735 2.655 ;
      RECT 26.79 6.225 27.11 6.55 ;
      RECT 26.82 5.7 26.99 6.55 ;
      RECT 26.82 5.7 26.995 6.05 ;
      RECT 26.82 5.7 27.795 5.875 ;
      RECT 27.62 1.97 27.795 5.875 ;
      RECT 27.565 1.97 27.915 2.32 ;
      RECT 27.59 6.66 27.915 6.985 ;
      RECT 26.475 6.75 27.915 6.92 ;
      RECT 26.475 2.4 26.635 6.92 ;
      RECT 26.79 2.37 27.11 2.69 ;
      RECT 26.475 2.4 27.11 2.57 ;
      RECT 23.925 3.545 24.185 3.865 ;
      RECT 23.985 1.84 24.125 3.865 ;
      RECT 25.185 2.705 25.525 3.055 ;
      RECT 24.56 2.775 25.525 2.975 ;
      RECT 24.56 1.945 24.76 2.975 ;
      RECT 23.81 2.4 24.125 2.77 ;
      RECT 25.275 2.7 25.445 3.055 ;
      RECT 23.88 1.955 24.125 2.77 ;
      RECT 23.915 1.84 24.195 2.21 ;
      RECT 23.915 1.945 24.76 2.145 ;
      RECT 23.235 2.425 23.495 2.745 ;
      RECT 22.575 2.515 23.495 2.655 ;
      RECT 22.575 1.575 22.715 2.655 ;
      RECT 19.035 1.865 19.295 2.185 ;
      RECT 19.215 1.575 19.355 2.095 ;
      RECT 19.215 1.575 22.715 1.715 ;
      RECT 14.71 6.66 15.06 7.01 ;
      RECT 22.15 6.615 22.5 6.965 ;
      RECT 14.71 6.69 22.5 6.89 ;
      RECT 22.065 3.265 22.325 3.585 ;
      RECT 22.125 1.855 22.265 3.585 ;
      RECT 22.055 1.855 22.335 2.225 ;
      RECT 19.455 4.015 21.89 4.155 ;
      RECT 21.75 2.705 21.89 4.155 ;
      RECT 19.455 3.635 19.595 4.155 ;
      RECT 19.155 3.635 19.595 3.865 ;
      RECT 16.815 3.635 19.595 3.775 ;
      RECT 19.155 3.545 19.415 3.865 ;
      RECT 16.815 3.355 16.955 3.775 ;
      RECT 16.305 3.265 16.565 3.585 ;
      RECT 16.305 3.355 16.955 3.495 ;
      RECT 16.365 1.865 16.505 3.585 ;
      RECT 21.69 2.705 21.95 3.025 ;
      RECT 16.305 1.865 16.565 2.185 ;
      RECT 21.315 3.545 21.575 3.865 ;
      RECT 21.375 1.955 21.515 3.865 ;
      RECT 21.035 1.955 21.515 2.23 ;
      RECT 20.835 1.86 21.315 2.205 ;
      RECT 20.825 3.495 21.105 3.865 ;
      RECT 20.895 2.4 21.035 3.865 ;
      RECT 20.835 2.4 21.095 3.025 ;
      RECT 20.825 2.4 21.105 2.77 ;
      RECT 19.755 3.545 20.015 3.865 ;
      RECT 19.755 3.355 19.955 3.865 ;
      RECT 19.56 3.355 19.955 3.495 ;
      RECT 19.56 1.865 19.7 3.495 ;
      RECT 19.56 1.865 19.875 2.235 ;
      RECT 19.5 1.865 19.875 2.185 ;
      RECT 17.225 2.96 17.505 3.33 ;
      RECT 18.675 2.985 18.935 3.305 ;
      RECT 17.055 3.075 18.935 3.215 ;
      RECT 17.055 2.96 17.505 3.215 ;
      RECT 16.995 2.4 17.255 3.025 ;
      RECT 16.985 2.4 17.265 2.77 ;
      RECT 18.065 2.4 18.475 2.77 ;
      RECT 17.475 2.425 17.735 2.745 ;
      RECT 17.475 2.515 18.475 2.655 ;
      RECT 11.53 6.225 11.85 6.55 ;
      RECT 11.56 5.7 11.73 6.55 ;
      RECT 11.56 5.7 11.735 6.05 ;
      RECT 11.56 5.7 12.535 5.875 ;
      RECT 12.36 1.97 12.535 5.875 ;
      RECT 12.305 1.97 12.655 2.32 ;
      RECT 12.33 6.66 12.655 6.985 ;
      RECT 11.215 6.75 12.655 6.92 ;
      RECT 11.215 2.4 11.375 6.92 ;
      RECT 11.53 2.37 11.85 2.69 ;
      RECT 11.215 2.4 11.85 2.57 ;
      RECT 8.665 3.545 8.925 3.865 ;
      RECT 8.725 1.84 8.865 3.865 ;
      RECT 9.925 2.705 10.265 3.055 ;
      RECT 9.3 2.775 10.265 2.975 ;
      RECT 9.3 1.945 9.5 2.975 ;
      RECT 8.55 2.4 8.865 2.77 ;
      RECT 10.015 2.7 10.185 3.055 ;
      RECT 8.62 1.955 8.865 2.77 ;
      RECT 8.655 1.84 8.935 2.21 ;
      RECT 8.655 1.945 9.5 2.145 ;
      RECT 7.975 2.425 8.235 2.745 ;
      RECT 7.315 2.515 8.235 2.655 ;
      RECT 7.315 1.575 7.455 2.655 ;
      RECT 3.775 1.865 4.035 2.185 ;
      RECT 3.955 1.575 4.095 2.095 ;
      RECT 3.955 1.575 7.455 1.715 ;
      RECT -1.255 7 -0.965 7.35 ;
      RECT -1.255 7.07 -0.035 7.24 ;
      RECT -0.205 6.69 -0.035 7.24 ;
      RECT 6.89 6.61 7.24 6.96 ;
      RECT -0.205 6.69 7.24 6.86 ;
      RECT 6.805 3.265 7.065 3.585 ;
      RECT 6.865 1.855 7.005 3.585 ;
      RECT 6.795 1.855 7.075 2.225 ;
      RECT 4.195 4.015 6.63 4.155 ;
      RECT 6.49 2.705 6.63 4.155 ;
      RECT 4.195 3.635 4.335 4.155 ;
      RECT 3.895 3.635 4.335 3.865 ;
      RECT 1.555 3.635 4.335 3.775 ;
      RECT 3.895 3.545 4.155 3.865 ;
      RECT 1.555 3.355 1.695 3.775 ;
      RECT 1.045 3.265 1.305 3.585 ;
      RECT 1.045 3.355 1.695 3.495 ;
      RECT 1.105 1.865 1.245 3.585 ;
      RECT 6.43 2.705 6.69 3.025 ;
      RECT 1.045 1.865 1.305 2.185 ;
      RECT 6.055 3.545 6.315 3.865 ;
      RECT 6.115 1.955 6.255 3.865 ;
      RECT 5.775 1.955 6.255 2.23 ;
      RECT 5.575 1.86 6.055 2.205 ;
      RECT 5.565 3.495 5.845 3.865 ;
      RECT 5.635 2.4 5.775 3.865 ;
      RECT 5.575 2.4 5.835 3.025 ;
      RECT 5.565 2.4 5.845 2.77 ;
      RECT 4.495 3.545 4.755 3.865 ;
      RECT 4.495 3.355 4.695 3.865 ;
      RECT 4.3 3.355 4.695 3.495 ;
      RECT 4.3 1.865 4.44 3.495 ;
      RECT 4.3 1.865 4.615 2.235 ;
      RECT 4.24 1.865 4.615 2.185 ;
      RECT 1.965 2.96 2.245 3.33 ;
      RECT 3.415 2.985 3.675 3.305 ;
      RECT 1.795 3.075 3.675 3.215 ;
      RECT 1.795 2.96 2.245 3.215 ;
      RECT 1.735 2.4 1.995 3.025 ;
      RECT 1.725 2.4 2.005 2.77 ;
      RECT 2.805 2.4 3.215 2.77 ;
      RECT 2.215 2.425 2.475 2.745 ;
      RECT 2.215 2.515 3.215 2.655 ;
      RECT 67.26 7.06 67.63 7.43 ;
      RECT 66.125 2.4 66.405 2.865 ;
      RECT 65.885 1.865 66.165 2.21 ;
      RECT 64.685 2.4 64.965 2.77 ;
      RECT 62.125 1.22 62.495 1.225 ;
      RECT 52 7.06 52.37 7.43 ;
      RECT 50.865 2.4 51.145 2.865 ;
      RECT 50.625 1.865 50.905 2.21 ;
      RECT 49.425 2.4 49.705 2.77 ;
      RECT 46.865 1.22 47.235 1.225 ;
      RECT 36.74 7.06 37.11 7.43 ;
      RECT 35.605 2.4 35.885 2.865 ;
      RECT 35.365 1.865 35.645 2.21 ;
      RECT 34.165 2.4 34.445 2.77 ;
      RECT 31.605 1.22 31.975 1.225 ;
      RECT 21.48 7.06 21.85 7.43 ;
      RECT 20.345 2.4 20.625 2.865 ;
      RECT 20.105 1.865 20.385 2.21 ;
      RECT 18.905 2.4 19.185 2.77 ;
      RECT 16.345 1.22 16.715 1.225 ;
      RECT 6.22 7.06 6.59 7.43 ;
      RECT 5.085 2.4 5.365 2.865 ;
      RECT 4.845 1.865 5.125 2.21 ;
      RECT 3.645 2.4 3.925 2.77 ;
      RECT 1.085 1.22 1.455 1.225 ;
    LAYER via1 ;
      RECT 75.83 7.38 75.98 7.53 ;
      RECT 73.46 6.745 73.61 6.895 ;
      RECT 73.445 2.07 73.595 2.22 ;
      RECT 72.655 2.455 72.805 2.605 ;
      RECT 72.655 6.33 72.805 6.48 ;
      RECT 71.065 2.805 71.215 2.955 ;
      RECT 69.76 1.95 69.91 2.1 ;
      RECT 69.76 3.63 69.91 3.78 ;
      RECT 69.07 2.51 69.22 2.66 ;
      RECT 68.03 6.715 68.18 6.865 ;
      RECT 67.9 1.95 68.05 2.1 ;
      RECT 67.9 3.35 68.05 3.5 ;
      RECT 67.525 2.79 67.675 2.94 ;
      RECT 67.37 7.17 67.52 7.32 ;
      RECT 67.15 3.63 67.3 3.78 ;
      RECT 66.67 1.95 66.82 2.1 ;
      RECT 66.67 2.79 66.82 2.94 ;
      RECT 66.19 2.51 66.34 2.66 ;
      RECT 65.95 1.95 66.1 2.1 ;
      RECT 65.59 3.63 65.74 3.78 ;
      RECT 65.335 1.95 65.485 2.1 ;
      RECT 64.99 3.63 65.14 3.78 ;
      RECT 64.87 1.95 65.02 2.1 ;
      RECT 64.75 2.51 64.9 2.66 ;
      RECT 64.51 3.07 64.66 3.22 ;
      RECT 63.31 2.51 63.46 2.66 ;
      RECT 62.83 2.79 62.98 2.94 ;
      RECT 62.14 1.95 62.29 2.1 ;
      RECT 62.14 3.35 62.29 3.5 ;
      RECT 60.545 6.76 60.695 6.91 ;
      RECT 58.2 6.745 58.35 6.895 ;
      RECT 58.185 2.07 58.335 2.22 ;
      RECT 57.395 2.455 57.545 2.605 ;
      RECT 57.395 6.33 57.545 6.48 ;
      RECT 55.805 2.805 55.955 2.955 ;
      RECT 54.5 1.95 54.65 2.1 ;
      RECT 54.5 3.63 54.65 3.78 ;
      RECT 53.81 2.51 53.96 2.66 ;
      RECT 52.775 6.715 52.925 6.865 ;
      RECT 52.64 1.95 52.79 2.1 ;
      RECT 52.64 3.35 52.79 3.5 ;
      RECT 52.265 2.79 52.415 2.94 ;
      RECT 52.11 7.17 52.26 7.32 ;
      RECT 51.89 3.63 52.04 3.78 ;
      RECT 51.41 1.95 51.56 2.1 ;
      RECT 51.41 2.79 51.56 2.94 ;
      RECT 50.93 2.51 51.08 2.66 ;
      RECT 50.69 1.95 50.84 2.1 ;
      RECT 50.33 3.63 50.48 3.78 ;
      RECT 50.075 1.95 50.225 2.1 ;
      RECT 49.73 3.63 49.88 3.78 ;
      RECT 49.61 1.95 49.76 2.1 ;
      RECT 49.49 2.51 49.64 2.66 ;
      RECT 49.25 3.07 49.4 3.22 ;
      RECT 48.05 2.51 48.2 2.66 ;
      RECT 47.57 2.79 47.72 2.94 ;
      RECT 46.88 1.95 47.03 2.1 ;
      RECT 46.88 3.35 47.03 3.5 ;
      RECT 45.285 6.76 45.435 6.91 ;
      RECT 42.94 6.745 43.09 6.895 ;
      RECT 42.925 2.07 43.075 2.22 ;
      RECT 42.135 2.455 42.285 2.605 ;
      RECT 42.135 6.33 42.285 6.48 ;
      RECT 40.545 2.805 40.695 2.955 ;
      RECT 39.24 1.95 39.39 2.1 ;
      RECT 39.24 3.63 39.39 3.78 ;
      RECT 38.55 2.51 38.7 2.66 ;
      RECT 37.51 6.72 37.66 6.87 ;
      RECT 37.38 1.95 37.53 2.1 ;
      RECT 37.38 3.35 37.53 3.5 ;
      RECT 37.005 2.79 37.155 2.94 ;
      RECT 36.85 7.17 37 7.32 ;
      RECT 36.63 3.63 36.78 3.78 ;
      RECT 36.15 1.95 36.3 2.1 ;
      RECT 36.15 2.79 36.3 2.94 ;
      RECT 35.67 2.51 35.82 2.66 ;
      RECT 35.43 1.95 35.58 2.1 ;
      RECT 35.07 3.63 35.22 3.78 ;
      RECT 34.815 1.95 34.965 2.1 ;
      RECT 34.47 3.63 34.62 3.78 ;
      RECT 34.35 1.95 34.5 2.1 ;
      RECT 34.23 2.51 34.38 2.66 ;
      RECT 33.99 3.07 34.14 3.22 ;
      RECT 32.79 2.51 32.94 2.66 ;
      RECT 32.31 2.79 32.46 2.94 ;
      RECT 31.62 1.95 31.77 2.1 ;
      RECT 31.62 3.35 31.77 3.5 ;
      RECT 30.07 6.765 30.22 6.915 ;
      RECT 27.68 6.745 27.83 6.895 ;
      RECT 27.665 2.07 27.815 2.22 ;
      RECT 26.875 2.455 27.025 2.605 ;
      RECT 26.875 6.33 27.025 6.48 ;
      RECT 25.285 2.805 25.435 2.955 ;
      RECT 23.98 1.95 24.13 2.1 ;
      RECT 23.98 3.63 24.13 3.78 ;
      RECT 23.29 2.51 23.44 2.66 ;
      RECT 22.25 6.715 22.4 6.865 ;
      RECT 22.12 1.95 22.27 2.1 ;
      RECT 22.12 3.35 22.27 3.5 ;
      RECT 21.745 2.79 21.895 2.94 ;
      RECT 21.59 7.17 21.74 7.32 ;
      RECT 21.37 3.63 21.52 3.78 ;
      RECT 20.89 1.95 21.04 2.1 ;
      RECT 20.89 2.79 21.04 2.94 ;
      RECT 20.41 2.51 20.56 2.66 ;
      RECT 20.17 1.95 20.32 2.1 ;
      RECT 19.81 3.63 19.96 3.78 ;
      RECT 19.555 1.95 19.705 2.1 ;
      RECT 19.21 3.63 19.36 3.78 ;
      RECT 19.09 1.95 19.24 2.1 ;
      RECT 18.97 2.51 19.12 2.66 ;
      RECT 18.73 3.07 18.88 3.22 ;
      RECT 17.53 2.51 17.68 2.66 ;
      RECT 17.05 2.79 17.2 2.94 ;
      RECT 16.36 1.95 16.51 2.1 ;
      RECT 16.36 3.35 16.51 3.5 ;
      RECT 14.81 6.76 14.96 6.91 ;
      RECT 12.42 6.745 12.57 6.895 ;
      RECT 12.405 2.07 12.555 2.22 ;
      RECT 11.615 2.455 11.765 2.605 ;
      RECT 11.615 6.33 11.765 6.48 ;
      RECT 10.025 2.805 10.175 2.955 ;
      RECT 8.72 1.95 8.87 2.1 ;
      RECT 8.72 3.63 8.87 3.78 ;
      RECT 8.03 2.51 8.18 2.66 ;
      RECT 6.99 6.71 7.14 6.86 ;
      RECT 6.86 1.95 7.01 2.1 ;
      RECT 6.86 3.35 7.01 3.5 ;
      RECT 6.485 2.79 6.635 2.94 ;
      RECT 6.33 7.17 6.48 7.32 ;
      RECT 6.11 3.63 6.26 3.78 ;
      RECT 5.63 1.95 5.78 2.1 ;
      RECT 5.63 2.79 5.78 2.94 ;
      RECT 5.15 2.51 5.3 2.66 ;
      RECT 4.91 1.95 5.06 2.1 ;
      RECT 4.55 3.63 4.7 3.78 ;
      RECT 4.295 1.95 4.445 2.1 ;
      RECT 3.95 3.63 4.1 3.78 ;
      RECT 3.83 1.95 3.98 2.1 ;
      RECT 3.71 2.51 3.86 2.66 ;
      RECT 3.47 3.07 3.62 3.22 ;
      RECT 2.27 2.51 2.42 2.66 ;
      RECT 1.79 2.79 1.94 2.94 ;
      RECT 1.1 1.95 1.25 2.1 ;
      RECT 1.1 3.35 1.25 3.5 ;
      RECT -1.185 7.1 -1.035 7.25 ;
      RECT -1.56 6.36 -1.41 6.51 ;
    LAYER met1 ;
      RECT 75.695 7.775 75.985 8.005 ;
      RECT 75.755 6.295 75.925 8.005 ;
      RECT 75.73 7.28 76.08 7.63 ;
      RECT 75.695 6.295 75.985 6.525 ;
      RECT 75.29 2.4 75.395 2.97 ;
      RECT 75.29 2.735 75.615 2.965 ;
      RECT 75.29 2.765 75.785 2.935 ;
      RECT 75.29 2.4 75.48 2.965 ;
      RECT 74.705 2.365 74.995 2.595 ;
      RECT 74.705 2.4 75.48 2.57 ;
      RECT 74.765 0.885 74.935 2.595 ;
      RECT 74.705 0.885 74.995 1.115 ;
      RECT 74.705 7.775 74.995 8.005 ;
      RECT 74.765 6.295 74.935 8.005 ;
      RECT 74.705 6.295 74.995 6.525 ;
      RECT 74.705 6.33 75.56 6.49 ;
      RECT 75.39 5.925 75.56 6.49 ;
      RECT 74.705 6.325 75.1 6.49 ;
      RECT 75.325 5.925 75.615 6.155 ;
      RECT 75.325 5.955 75.785 6.125 ;
      RECT 74.335 2.735 74.625 2.965 ;
      RECT 74.335 2.765 74.795 2.935 ;
      RECT 74.4 1.66 74.565 2.965 ;
      RECT 72.915 1.63 73.205 1.86 ;
      RECT 72.915 1.66 74.565 1.83 ;
      RECT 72.975 0.89 73.145 1.86 ;
      RECT 72.915 0.89 73.205 1.12 ;
      RECT 72.915 7.77 73.205 8 ;
      RECT 72.975 7.03 73.145 8 ;
      RECT 72.975 7.125 74.565 7.295 ;
      RECT 74.395 5.925 74.565 7.295 ;
      RECT 72.915 7.03 73.205 7.26 ;
      RECT 74.335 5.925 74.625 6.155 ;
      RECT 74.335 5.955 74.795 6.125 ;
      RECT 70.965 2.705 71.305 3.055 ;
      RECT 71.055 2.03 71.225 3.055 ;
      RECT 73.345 1.97 73.695 2.32 ;
      RECT 71.055 2.03 73.695 2.2 ;
      RECT 73.37 6.66 73.695 6.985 ;
      RECT 67.93 6.615 68.28 6.965 ;
      RECT 73.345 6.66 73.695 6.89 ;
      RECT 67.73 6.66 68.28 6.89 ;
      RECT 67.56 6.69 73.695 6.86 ;
      RECT 72.57 2.37 72.89 2.69 ;
      RECT 72.54 2.37 72.89 2.6 ;
      RECT 72.37 2.4 72.89 2.57 ;
      RECT 72.57 6.26 72.89 6.55 ;
      RECT 72.54 6.29 72.89 6.52 ;
      RECT 72.37 6.32 72.89 6.49 ;
      RECT 69.675 1.895 69.995 2.155 ;
      RECT 69.24 1.91 69.53 2.14 ;
      RECT 69.24 1.955 69.995 2.095 ;
      RECT 69.675 3.575 69.995 3.835 ;
      RECT 69.24 3.59 69.53 3.82 ;
      RECT 69.24 3.635 69.995 3.775 ;
      RECT 69 3.03 69.29 3.26 ;
      RECT 69 3.075 69.575 3.215 ;
      RECT 69.435 2.935 69.695 3.075 ;
      RECT 69.48 2.75 69.77 2.98 ;
      RECT 67.635 2.935 68.735 3.075 ;
      RECT 67.44 2.735 67.76 2.995 ;
      RECT 68.52 2.75 68.81 2.98 ;
      RECT 67.44 2.75 67.85 2.995 ;
      RECT 67.815 1.895 68.135 2.155 ;
      RECT 68.28 1.91 68.57 2.14 ;
      RECT 67.815 1.955 68.57 2.095 ;
      RECT 65.115 3.16 67.295 3.3 ;
      RECT 67.155 2.17 67.295 3.3 ;
      RECT 65.115 3.075 66.41 3.3 ;
      RECT 66.12 3.03 66.41 3.3 ;
      RECT 65.115 2.795 65.45 3.3 ;
      RECT 65.16 2.75 65.45 3.3 ;
      RECT 68.04 2.47 68.33 2.7 ;
      RECT 67.155 2.375 68.255 2.515 ;
      RECT 67.08 2.17 67.37 2.42 ;
      RECT 67.3 7.77 67.59 8 ;
      RECT 67.36 7.03 67.53 8 ;
      RECT 67.26 7.06 67.63 7.43 ;
      RECT 67.3 7.03 67.59 7.43 ;
      RECT 67.065 3.575 67.385 3.835 ;
      RECT 67.065 3.59 67.58 3.82 ;
      RECT 65.64 2.47 65.93 2.7 ;
      RECT 65.79 2.075 65.93 2.7 ;
      RECT 65.79 2.075 66.095 2.215 ;
      RECT 66.585 1.895 66.905 2.155 ;
      RECT 65.865 1.895 66.185 2.155 ;
      RECT 66.36 1.91 66.905 2.14 ;
      RECT 65.865 1.955 66.905 2.095 ;
      RECT 65.505 3.575 65.825 3.835 ;
      RECT 65.4 3.59 65.825 3.82 ;
      RECT 63.48 3.03 63.77 3.26 ;
      RECT 63.48 3.03 63.935 3.215 ;
      RECT 63.795 2.555 63.935 3.215 ;
      RECT 63.915 1.955 64.055 2.695 ;
      RECT 64.785 1.895 65.105 2.155 ;
      RECT 63.96 1.91 64.25 2.14 ;
      RECT 63.915 1.955 65.105 2.095 ;
      RECT 64.665 2.455 64.985 2.715 ;
      RECT 64.2 2.47 64.49 2.7 ;
      RECT 64.2 2.515 64.985 2.655 ;
      RECT 64.425 3.015 64.745 3.275 ;
      RECT 64.425 3.03 64.97 3.26 ;
      RECT 63.96 3.59 64.25 3.82 ;
      RECT 63.075 3.47 64.175 3.61 ;
      RECT 63 3.31 63.29 3.54 ;
      RECT 60.435 7.775 60.725 8.005 ;
      RECT 60.495 6.295 60.665 8.005 ;
      RECT 60.445 6.66 60.795 7.01 ;
      RECT 60.435 6.295 60.725 6.525 ;
      RECT 60.03 2.4 60.135 2.97 ;
      RECT 60.03 2.735 60.355 2.965 ;
      RECT 60.03 2.765 60.525 2.935 ;
      RECT 60.03 2.4 60.22 2.965 ;
      RECT 59.445 2.365 59.735 2.595 ;
      RECT 59.445 2.4 60.22 2.57 ;
      RECT 59.505 0.885 59.675 2.595 ;
      RECT 59.445 0.885 59.735 1.115 ;
      RECT 59.445 7.775 59.735 8.005 ;
      RECT 59.505 6.295 59.675 8.005 ;
      RECT 59.445 6.295 59.735 6.525 ;
      RECT 59.445 6.33 60.3 6.49 ;
      RECT 60.13 5.925 60.3 6.49 ;
      RECT 59.445 6.325 59.84 6.49 ;
      RECT 60.065 5.925 60.355 6.155 ;
      RECT 60.065 5.955 60.525 6.125 ;
      RECT 59.075 2.735 59.365 2.965 ;
      RECT 59.075 2.765 59.535 2.935 ;
      RECT 59.14 1.66 59.305 2.965 ;
      RECT 57.655 1.63 57.945 1.86 ;
      RECT 57.655 1.66 59.305 1.83 ;
      RECT 57.715 0.89 57.885 1.86 ;
      RECT 57.655 0.89 57.945 1.12 ;
      RECT 57.655 7.77 57.945 8 ;
      RECT 57.715 7.03 57.885 8 ;
      RECT 57.715 7.125 59.305 7.295 ;
      RECT 59.135 5.925 59.305 7.295 ;
      RECT 57.655 7.03 57.945 7.26 ;
      RECT 59.075 5.925 59.365 6.155 ;
      RECT 59.075 5.955 59.535 6.125 ;
      RECT 55.705 2.705 56.045 3.055 ;
      RECT 55.795 2.03 55.965 3.055 ;
      RECT 58.085 1.97 58.435 2.32 ;
      RECT 55.795 2.03 58.435 2.2 ;
      RECT 58.11 6.66 58.435 6.985 ;
      RECT 52.675 6.615 53.025 6.965 ;
      RECT 58.085 6.66 58.435 6.89 ;
      RECT 52.47 6.66 53.025 6.89 ;
      RECT 52.3 6.69 58.435 6.86 ;
      RECT 57.31 2.37 57.63 2.69 ;
      RECT 57.28 2.37 57.63 2.6 ;
      RECT 57.11 2.4 57.63 2.57 ;
      RECT 57.31 6.26 57.63 6.55 ;
      RECT 57.28 6.29 57.63 6.52 ;
      RECT 57.11 6.32 57.63 6.49 ;
      RECT 54.415 1.895 54.735 2.155 ;
      RECT 53.98 1.91 54.27 2.14 ;
      RECT 53.98 1.955 54.735 2.095 ;
      RECT 54.415 3.575 54.735 3.835 ;
      RECT 53.98 3.59 54.27 3.82 ;
      RECT 53.98 3.635 54.735 3.775 ;
      RECT 53.74 3.03 54.03 3.26 ;
      RECT 53.74 3.075 54.315 3.215 ;
      RECT 54.175 2.935 54.435 3.075 ;
      RECT 54.22 2.75 54.51 2.98 ;
      RECT 52.375 2.935 53.475 3.075 ;
      RECT 52.18 2.735 52.5 2.995 ;
      RECT 53.26 2.75 53.55 2.98 ;
      RECT 52.18 2.75 52.59 2.995 ;
      RECT 52.555 1.895 52.875 2.155 ;
      RECT 53.02 1.91 53.31 2.14 ;
      RECT 52.555 1.955 53.31 2.095 ;
      RECT 49.855 3.16 52.035 3.3 ;
      RECT 51.895 2.17 52.035 3.3 ;
      RECT 49.855 3.075 51.15 3.3 ;
      RECT 50.86 3.03 51.15 3.3 ;
      RECT 49.855 2.795 50.19 3.3 ;
      RECT 49.9 2.75 50.19 3.3 ;
      RECT 52.78 2.47 53.07 2.7 ;
      RECT 51.895 2.375 52.995 2.515 ;
      RECT 51.82 2.17 52.11 2.42 ;
      RECT 52.04 7.77 52.33 8 ;
      RECT 52.1 7.03 52.27 8 ;
      RECT 52 7.06 52.37 7.43 ;
      RECT 52.04 7.03 52.33 7.43 ;
      RECT 51.805 3.575 52.125 3.835 ;
      RECT 51.805 3.59 52.32 3.82 ;
      RECT 50.38 2.47 50.67 2.7 ;
      RECT 50.53 2.075 50.67 2.7 ;
      RECT 50.53 2.075 50.835 2.215 ;
      RECT 51.325 1.895 51.645 2.155 ;
      RECT 50.605 1.895 50.925 2.155 ;
      RECT 51.1 1.91 51.645 2.14 ;
      RECT 50.605 1.955 51.645 2.095 ;
      RECT 50.245 3.575 50.565 3.835 ;
      RECT 50.14 3.59 50.565 3.82 ;
      RECT 48.22 3.03 48.51 3.26 ;
      RECT 48.22 3.03 48.675 3.215 ;
      RECT 48.535 2.555 48.675 3.215 ;
      RECT 48.655 1.955 48.795 2.695 ;
      RECT 49.525 1.895 49.845 2.155 ;
      RECT 48.7 1.91 48.99 2.14 ;
      RECT 48.655 1.955 49.845 2.095 ;
      RECT 49.405 2.455 49.725 2.715 ;
      RECT 48.94 2.47 49.23 2.7 ;
      RECT 48.94 2.515 49.725 2.655 ;
      RECT 49.165 3.015 49.485 3.275 ;
      RECT 49.165 3.03 49.71 3.26 ;
      RECT 48.7 3.59 48.99 3.82 ;
      RECT 47.815 3.47 48.915 3.61 ;
      RECT 47.74 3.31 48.03 3.54 ;
      RECT 45.175 7.775 45.465 8.005 ;
      RECT 45.235 6.295 45.405 8.005 ;
      RECT 45.185 6.66 45.535 7.01 ;
      RECT 45.175 6.295 45.465 6.525 ;
      RECT 44.77 2.4 44.875 2.97 ;
      RECT 44.77 2.735 45.095 2.965 ;
      RECT 44.77 2.765 45.265 2.935 ;
      RECT 44.77 2.4 44.96 2.965 ;
      RECT 44.185 2.365 44.475 2.595 ;
      RECT 44.185 2.4 44.96 2.57 ;
      RECT 44.245 0.885 44.415 2.595 ;
      RECT 44.185 0.885 44.475 1.115 ;
      RECT 44.185 7.775 44.475 8.005 ;
      RECT 44.245 6.295 44.415 8.005 ;
      RECT 44.185 6.295 44.475 6.525 ;
      RECT 44.185 6.33 45.04 6.49 ;
      RECT 44.87 5.925 45.04 6.49 ;
      RECT 44.185 6.325 44.58 6.49 ;
      RECT 44.805 5.925 45.095 6.155 ;
      RECT 44.805 5.955 45.265 6.125 ;
      RECT 43.815 2.735 44.105 2.965 ;
      RECT 43.815 2.765 44.275 2.935 ;
      RECT 43.88 1.66 44.045 2.965 ;
      RECT 42.395 1.63 42.685 1.86 ;
      RECT 42.395 1.66 44.045 1.83 ;
      RECT 42.455 0.89 42.625 1.86 ;
      RECT 42.395 0.89 42.685 1.12 ;
      RECT 42.395 7.77 42.685 8 ;
      RECT 42.455 7.03 42.625 8 ;
      RECT 42.455 7.125 44.045 7.295 ;
      RECT 43.875 5.925 44.045 7.295 ;
      RECT 42.395 7.03 42.685 7.26 ;
      RECT 43.815 5.925 44.105 6.155 ;
      RECT 43.815 5.955 44.275 6.125 ;
      RECT 40.445 2.705 40.785 3.055 ;
      RECT 40.535 2.03 40.705 3.055 ;
      RECT 42.825 1.97 43.175 2.32 ;
      RECT 40.535 2.03 43.175 2.2 ;
      RECT 42.85 6.66 43.175 6.985 ;
      RECT 37.41 6.62 37.76 6.97 ;
      RECT 42.825 6.66 43.175 6.89 ;
      RECT 37.21 6.66 37.76 6.89 ;
      RECT 37.04 6.69 43.175 6.86 ;
      RECT 42.05 2.37 42.37 2.69 ;
      RECT 42.02 2.37 42.37 2.6 ;
      RECT 41.85 2.4 42.37 2.57 ;
      RECT 42.05 6.26 42.37 6.55 ;
      RECT 42.02 6.29 42.37 6.52 ;
      RECT 41.85 6.32 42.37 6.49 ;
      RECT 39.155 1.895 39.475 2.155 ;
      RECT 38.72 1.91 39.01 2.14 ;
      RECT 38.72 1.955 39.475 2.095 ;
      RECT 39.155 3.575 39.475 3.835 ;
      RECT 38.72 3.59 39.01 3.82 ;
      RECT 38.72 3.635 39.475 3.775 ;
      RECT 38.48 3.03 38.77 3.26 ;
      RECT 38.48 3.075 39.055 3.215 ;
      RECT 38.915 2.935 39.175 3.075 ;
      RECT 38.96 2.75 39.25 2.98 ;
      RECT 37.115 2.935 38.215 3.075 ;
      RECT 36.92 2.735 37.24 2.995 ;
      RECT 38 2.75 38.29 2.98 ;
      RECT 36.92 2.75 37.33 2.995 ;
      RECT 37.295 1.895 37.615 2.155 ;
      RECT 37.76 1.91 38.05 2.14 ;
      RECT 37.295 1.955 38.05 2.095 ;
      RECT 34.595 3.16 36.775 3.3 ;
      RECT 36.635 2.17 36.775 3.3 ;
      RECT 34.595 3.075 35.89 3.3 ;
      RECT 35.6 3.03 35.89 3.3 ;
      RECT 34.595 2.795 34.93 3.3 ;
      RECT 34.64 2.75 34.93 3.3 ;
      RECT 37.52 2.47 37.81 2.7 ;
      RECT 36.635 2.375 37.735 2.515 ;
      RECT 36.56 2.17 36.85 2.42 ;
      RECT 36.78 7.77 37.07 8 ;
      RECT 36.84 7.03 37.01 8 ;
      RECT 36.74 7.06 37.11 7.43 ;
      RECT 36.78 7.03 37.07 7.43 ;
      RECT 36.545 3.575 36.865 3.835 ;
      RECT 36.545 3.59 37.06 3.82 ;
      RECT 35.12 2.47 35.41 2.7 ;
      RECT 35.27 2.075 35.41 2.7 ;
      RECT 35.27 2.075 35.575 2.215 ;
      RECT 36.065 1.895 36.385 2.155 ;
      RECT 35.345 1.895 35.665 2.155 ;
      RECT 35.84 1.91 36.385 2.14 ;
      RECT 35.345 1.955 36.385 2.095 ;
      RECT 34.985 3.575 35.305 3.835 ;
      RECT 34.88 3.59 35.305 3.82 ;
      RECT 32.96 3.03 33.25 3.26 ;
      RECT 32.96 3.03 33.415 3.215 ;
      RECT 33.275 2.555 33.415 3.215 ;
      RECT 33.395 1.955 33.535 2.695 ;
      RECT 34.265 1.895 34.585 2.155 ;
      RECT 33.44 1.91 33.73 2.14 ;
      RECT 33.395 1.955 34.585 2.095 ;
      RECT 34.145 2.455 34.465 2.715 ;
      RECT 33.68 2.47 33.97 2.7 ;
      RECT 33.68 2.515 34.465 2.655 ;
      RECT 33.905 3.015 34.225 3.275 ;
      RECT 33.905 3.03 34.45 3.26 ;
      RECT 33.44 3.59 33.73 3.82 ;
      RECT 32.555 3.47 33.655 3.61 ;
      RECT 32.48 3.31 32.77 3.54 ;
      RECT 29.915 7.775 30.205 8.005 ;
      RECT 29.975 6.295 30.145 8.005 ;
      RECT 29.965 6.665 30.32 7.02 ;
      RECT 29.915 6.295 30.205 6.525 ;
      RECT 29.51 2.4 29.615 2.97 ;
      RECT 29.51 2.735 29.835 2.965 ;
      RECT 29.51 2.765 30.005 2.935 ;
      RECT 29.51 2.4 29.7 2.965 ;
      RECT 28.925 2.365 29.215 2.595 ;
      RECT 28.925 2.4 29.7 2.57 ;
      RECT 28.985 0.885 29.155 2.595 ;
      RECT 28.925 0.885 29.215 1.115 ;
      RECT 28.925 7.775 29.215 8.005 ;
      RECT 28.985 6.295 29.155 8.005 ;
      RECT 28.925 6.295 29.215 6.525 ;
      RECT 28.925 6.33 29.78 6.49 ;
      RECT 29.61 5.925 29.78 6.49 ;
      RECT 28.925 6.325 29.32 6.49 ;
      RECT 29.545 5.925 29.835 6.155 ;
      RECT 29.545 5.955 30.005 6.125 ;
      RECT 28.555 2.735 28.845 2.965 ;
      RECT 28.555 2.765 29.015 2.935 ;
      RECT 28.62 1.66 28.785 2.965 ;
      RECT 27.135 1.63 27.425 1.86 ;
      RECT 27.135 1.66 28.785 1.83 ;
      RECT 27.195 0.89 27.365 1.86 ;
      RECT 27.135 0.89 27.425 1.12 ;
      RECT 27.135 7.77 27.425 8 ;
      RECT 27.195 7.03 27.365 8 ;
      RECT 27.195 7.125 28.785 7.295 ;
      RECT 28.615 5.925 28.785 7.295 ;
      RECT 27.135 7.03 27.425 7.26 ;
      RECT 28.555 5.925 28.845 6.155 ;
      RECT 28.555 5.955 29.015 6.125 ;
      RECT 25.185 2.705 25.525 3.055 ;
      RECT 25.275 2.03 25.445 3.055 ;
      RECT 27.565 1.97 27.915 2.32 ;
      RECT 25.275 2.03 27.915 2.2 ;
      RECT 27.59 6.66 27.915 6.985 ;
      RECT 22.15 6.615 22.5 6.965 ;
      RECT 27.565 6.66 27.915 6.89 ;
      RECT 21.95 6.66 22.5 6.89 ;
      RECT 21.78 6.69 27.915 6.86 ;
      RECT 26.79 2.37 27.11 2.69 ;
      RECT 26.76 2.37 27.11 2.6 ;
      RECT 26.59 2.4 27.11 2.57 ;
      RECT 26.79 6.26 27.11 6.55 ;
      RECT 26.76 6.29 27.11 6.52 ;
      RECT 26.59 6.32 27.11 6.49 ;
      RECT 23.895 1.895 24.215 2.155 ;
      RECT 23.46 1.91 23.75 2.14 ;
      RECT 23.46 1.955 24.215 2.095 ;
      RECT 23.895 3.575 24.215 3.835 ;
      RECT 23.46 3.59 23.75 3.82 ;
      RECT 23.46 3.635 24.215 3.775 ;
      RECT 23.22 3.03 23.51 3.26 ;
      RECT 23.22 3.075 23.795 3.215 ;
      RECT 23.655 2.935 23.915 3.075 ;
      RECT 23.7 2.75 23.99 2.98 ;
      RECT 21.855 2.935 22.955 3.075 ;
      RECT 21.66 2.735 21.98 2.995 ;
      RECT 22.74 2.75 23.03 2.98 ;
      RECT 21.66 2.75 22.07 2.995 ;
      RECT 22.035 1.895 22.355 2.155 ;
      RECT 22.5 1.91 22.79 2.14 ;
      RECT 22.035 1.955 22.79 2.095 ;
      RECT 19.335 3.16 21.515 3.3 ;
      RECT 21.375 2.17 21.515 3.3 ;
      RECT 19.335 3.075 20.63 3.3 ;
      RECT 20.34 3.03 20.63 3.3 ;
      RECT 19.335 2.795 19.67 3.3 ;
      RECT 19.38 2.75 19.67 3.3 ;
      RECT 22.26 2.47 22.55 2.7 ;
      RECT 21.375 2.375 22.475 2.515 ;
      RECT 21.3 2.17 21.59 2.42 ;
      RECT 21.52 7.77 21.81 8 ;
      RECT 21.58 7.03 21.75 8 ;
      RECT 21.48 7.06 21.85 7.43 ;
      RECT 21.52 7.03 21.81 7.43 ;
      RECT 21.285 3.575 21.605 3.835 ;
      RECT 21.285 3.59 21.8 3.82 ;
      RECT 19.86 2.47 20.15 2.7 ;
      RECT 20.01 2.075 20.15 2.7 ;
      RECT 20.01 2.075 20.315 2.215 ;
      RECT 20.805 1.895 21.125 2.155 ;
      RECT 20.085 1.895 20.405 2.155 ;
      RECT 20.58 1.91 21.125 2.14 ;
      RECT 20.085 1.955 21.125 2.095 ;
      RECT 19.725 3.575 20.045 3.835 ;
      RECT 19.62 3.59 20.045 3.82 ;
      RECT 17.7 3.03 17.99 3.26 ;
      RECT 17.7 3.03 18.155 3.215 ;
      RECT 18.015 2.555 18.155 3.215 ;
      RECT 18.135 1.955 18.275 2.695 ;
      RECT 19.005 1.895 19.325 2.155 ;
      RECT 18.18 1.91 18.47 2.14 ;
      RECT 18.135 1.955 19.325 2.095 ;
      RECT 18.885 2.455 19.205 2.715 ;
      RECT 18.42 2.47 18.71 2.7 ;
      RECT 18.42 2.515 19.205 2.655 ;
      RECT 18.645 3.015 18.965 3.275 ;
      RECT 18.645 3.03 19.19 3.26 ;
      RECT 18.18 3.59 18.47 3.82 ;
      RECT 17.295 3.47 18.395 3.61 ;
      RECT 17.22 3.31 17.51 3.54 ;
      RECT 14.655 7.775 14.945 8.005 ;
      RECT 14.715 6.295 14.885 8.005 ;
      RECT 14.71 6.66 15.06 7.01 ;
      RECT 14.655 6.295 14.945 6.525 ;
      RECT 14.25 2.4 14.355 2.97 ;
      RECT 14.25 2.735 14.575 2.965 ;
      RECT 14.25 2.765 14.745 2.935 ;
      RECT 14.25 2.4 14.44 2.965 ;
      RECT 13.665 2.365 13.955 2.595 ;
      RECT 13.665 2.4 14.44 2.57 ;
      RECT 13.725 0.885 13.895 2.595 ;
      RECT 13.665 0.885 13.955 1.115 ;
      RECT 13.665 7.775 13.955 8.005 ;
      RECT 13.725 6.295 13.895 8.005 ;
      RECT 13.665 6.295 13.955 6.525 ;
      RECT 13.665 6.33 14.52 6.49 ;
      RECT 14.35 5.925 14.52 6.49 ;
      RECT 13.665 6.325 14.06 6.49 ;
      RECT 14.285 5.925 14.575 6.155 ;
      RECT 14.285 5.955 14.745 6.125 ;
      RECT 13.295 2.735 13.585 2.965 ;
      RECT 13.295 2.765 13.755 2.935 ;
      RECT 13.36 1.66 13.525 2.965 ;
      RECT 11.875 1.63 12.165 1.86 ;
      RECT 11.875 1.66 13.525 1.83 ;
      RECT 11.935 0.89 12.105 1.86 ;
      RECT 11.875 0.89 12.165 1.12 ;
      RECT 11.875 7.77 12.165 8 ;
      RECT 11.935 7.03 12.105 8 ;
      RECT 11.935 7.125 13.525 7.295 ;
      RECT 13.355 5.925 13.525 7.295 ;
      RECT 11.875 7.03 12.165 7.26 ;
      RECT 13.295 5.925 13.585 6.155 ;
      RECT 13.295 5.955 13.755 6.125 ;
      RECT 9.925 2.705 10.265 3.055 ;
      RECT 10.015 2.03 10.185 3.055 ;
      RECT 12.305 1.97 12.655 2.32 ;
      RECT 10.015 2.03 12.655 2.2 ;
      RECT 12.33 6.66 12.655 6.985 ;
      RECT 6.89 6.61 7.24 6.96 ;
      RECT 12.305 6.66 12.655 6.89 ;
      RECT 6.69 6.66 7.24 6.89 ;
      RECT 6.52 6.69 12.655 6.86 ;
      RECT 11.53 2.37 11.85 2.69 ;
      RECT 11.5 2.37 11.85 2.6 ;
      RECT 11.33 2.4 11.85 2.57 ;
      RECT 11.53 6.26 11.85 6.55 ;
      RECT 11.5 6.29 11.85 6.52 ;
      RECT 11.33 6.32 11.85 6.49 ;
      RECT 8.635 1.895 8.955 2.155 ;
      RECT 8.2 1.91 8.49 2.14 ;
      RECT 8.2 1.955 8.955 2.095 ;
      RECT 8.635 3.575 8.955 3.835 ;
      RECT 8.2 3.59 8.49 3.82 ;
      RECT 8.2 3.635 8.955 3.775 ;
      RECT 7.96 3.03 8.25 3.26 ;
      RECT 7.96 3.075 8.535 3.215 ;
      RECT 8.395 2.935 8.655 3.075 ;
      RECT 8.44 2.75 8.73 2.98 ;
      RECT 6.595 2.935 7.695 3.075 ;
      RECT 6.4 2.735 6.72 2.995 ;
      RECT 7.48 2.75 7.77 2.98 ;
      RECT 6.4 2.75 6.81 2.995 ;
      RECT 6.775 1.895 7.095 2.155 ;
      RECT 7.24 1.91 7.53 2.14 ;
      RECT 6.775 1.955 7.53 2.095 ;
      RECT 4.075 3.16 6.255 3.3 ;
      RECT 6.115 2.17 6.255 3.3 ;
      RECT 4.075 3.075 5.37 3.3 ;
      RECT 5.08 3.03 5.37 3.3 ;
      RECT 4.075 2.795 4.41 3.3 ;
      RECT 4.12 2.75 4.41 3.3 ;
      RECT 7 2.47 7.29 2.7 ;
      RECT 6.115 2.375 7.215 2.515 ;
      RECT 6.04 2.17 6.33 2.42 ;
      RECT 6.26 7.77 6.55 8 ;
      RECT 6.32 7.03 6.49 8 ;
      RECT 6.22 7.06 6.59 7.43 ;
      RECT 6.26 7.03 6.55 7.43 ;
      RECT 6.025 3.575 6.345 3.835 ;
      RECT 6.025 3.59 6.54 3.82 ;
      RECT 4.6 2.47 4.89 2.7 ;
      RECT 4.75 2.075 4.89 2.7 ;
      RECT 4.75 2.075 5.055 2.215 ;
      RECT 5.545 1.895 5.865 2.155 ;
      RECT 4.825 1.895 5.145 2.155 ;
      RECT 5.32 1.91 5.865 2.14 ;
      RECT 4.825 1.955 5.865 2.095 ;
      RECT 4.465 3.575 4.785 3.835 ;
      RECT 4.36 3.59 4.785 3.82 ;
      RECT 2.44 3.03 2.73 3.26 ;
      RECT 2.44 3.03 2.895 3.215 ;
      RECT 2.755 2.555 2.895 3.215 ;
      RECT 2.875 1.955 3.015 2.695 ;
      RECT 3.745 1.895 4.065 2.155 ;
      RECT 2.92 1.91 3.21 2.14 ;
      RECT 2.875 1.955 4.065 2.095 ;
      RECT 3.625 2.455 3.945 2.715 ;
      RECT 3.16 2.47 3.45 2.7 ;
      RECT 3.16 2.515 3.945 2.655 ;
      RECT 3.385 3.015 3.705 3.275 ;
      RECT 3.385 3.03 3.93 3.26 ;
      RECT 2.92 3.59 3.21 3.82 ;
      RECT 2.035 3.47 3.135 3.61 ;
      RECT 1.96 3.31 2.25 3.54 ;
      RECT -1.255 7.77 -0.965 8 ;
      RECT -1.195 7.03 -1.025 8 ;
      RECT -1.285 7.03 -0.935 7.32 ;
      RECT -1.66 6.29 -1.31 6.58 ;
      RECT -1.8 6.32 -1.31 6.49 ;
      RECT 68.985 2.455 69.305 2.715 ;
      RECT 67.815 3.295 68.135 3.555 ;
      RECT 66.585 2.735 66.905 2.995 ;
      RECT 66.105 2.455 66.425 2.715 ;
      RECT 65.25 1.895 65.65 2.155 ;
      RECT 64.905 3.575 65.225 3.835 ;
      RECT 63.225 2.455 63.545 2.715 ;
      RECT 62.745 2.735 63.065 2.995 ;
      RECT 62.055 1.895 62.375 2.155 ;
      RECT 62.055 3.295 62.375 3.555 ;
      RECT 53.725 2.455 54.045 2.715 ;
      RECT 52.555 3.295 52.875 3.555 ;
      RECT 51.325 2.735 51.645 2.995 ;
      RECT 50.845 2.455 51.165 2.715 ;
      RECT 49.99 1.895 50.39 2.155 ;
      RECT 49.645 3.575 49.965 3.835 ;
      RECT 47.965 2.455 48.285 2.715 ;
      RECT 47.485 2.735 47.805 2.995 ;
      RECT 46.795 1.895 47.115 2.155 ;
      RECT 46.795 3.295 47.115 3.555 ;
      RECT 38.465 2.455 38.785 2.715 ;
      RECT 37.295 3.295 37.615 3.555 ;
      RECT 36.065 2.735 36.385 2.995 ;
      RECT 35.585 2.455 35.905 2.715 ;
      RECT 34.73 1.895 35.13 2.155 ;
      RECT 34.385 3.575 34.705 3.835 ;
      RECT 32.705 2.455 33.025 2.715 ;
      RECT 32.225 2.735 32.545 2.995 ;
      RECT 31.535 1.895 31.855 2.155 ;
      RECT 31.535 3.295 31.855 3.555 ;
      RECT 23.205 2.455 23.525 2.715 ;
      RECT 22.035 3.295 22.355 3.555 ;
      RECT 20.805 2.735 21.125 2.995 ;
      RECT 20.325 2.455 20.645 2.715 ;
      RECT 19.47 1.895 19.87 2.155 ;
      RECT 19.125 3.575 19.445 3.835 ;
      RECT 17.445 2.455 17.765 2.715 ;
      RECT 16.965 2.735 17.285 2.995 ;
      RECT 16.275 1.895 16.595 2.155 ;
      RECT 16.275 3.295 16.595 3.555 ;
      RECT 7.945 2.455 8.265 2.715 ;
      RECT 6.775 3.295 7.095 3.555 ;
      RECT 5.545 2.735 5.865 2.995 ;
      RECT 5.065 2.455 5.385 2.715 ;
      RECT 4.21 1.895 4.61 2.155 ;
      RECT 3.865 3.575 4.185 3.835 ;
      RECT 2.185 2.455 2.505 2.715 ;
      RECT 1.705 2.735 2.025 2.995 ;
      RECT 1.015 1.895 1.335 2.155 ;
      RECT 1.015 3.295 1.335 3.555 ;
    LAYER mcon ;
      RECT 75.755 6.325 75.925 6.495 ;
      RECT 75.76 6.32 75.93 6.49 ;
      RECT 60.495 6.325 60.665 6.495 ;
      RECT 60.5 6.32 60.67 6.49 ;
      RECT 45.235 6.325 45.405 6.495 ;
      RECT 45.24 6.32 45.41 6.49 ;
      RECT 29.975 6.325 30.145 6.495 ;
      RECT 29.98 6.32 30.15 6.49 ;
      RECT 14.715 6.325 14.885 6.495 ;
      RECT 14.72 6.32 14.89 6.49 ;
      RECT 75.755 7.805 75.925 7.975 ;
      RECT 75.385 2.765 75.555 2.935 ;
      RECT 75.385 5.955 75.555 6.125 ;
      RECT 74.765 0.915 74.935 1.085 ;
      RECT 74.765 2.395 74.935 2.565 ;
      RECT 74.765 6.325 74.935 6.495 ;
      RECT 74.765 7.805 74.935 7.975 ;
      RECT 74.395 2.765 74.565 2.935 ;
      RECT 74.395 5.955 74.565 6.125 ;
      RECT 73.405 2.03 73.575 2.2 ;
      RECT 73.405 6.69 73.575 6.86 ;
      RECT 72.975 0.92 73.145 1.09 ;
      RECT 72.975 1.66 73.145 1.83 ;
      RECT 72.975 7.06 73.145 7.23 ;
      RECT 72.975 7.8 73.145 7.97 ;
      RECT 72.6 2.4 72.77 2.57 ;
      RECT 72.6 6.32 72.77 6.49 ;
      RECT 69.54 2.78 69.71 2.95 ;
      RECT 69.3 1.94 69.47 2.11 ;
      RECT 69.3 3.62 69.47 3.79 ;
      RECT 69.06 2.5 69.23 2.67 ;
      RECT 69.06 3.06 69.23 3.23 ;
      RECT 68.58 2.78 68.75 2.95 ;
      RECT 68.34 1.94 68.51 2.11 ;
      RECT 68.1 2.5 68.27 2.67 ;
      RECT 67.89 3.34 68.06 3.51 ;
      RECT 67.79 6.69 67.96 6.86 ;
      RECT 67.62 2.78 67.79 2.95 ;
      RECT 67.36 7.06 67.53 7.23 ;
      RECT 67.36 7.8 67.53 7.97 ;
      RECT 67.35 3.62 67.52 3.79 ;
      RECT 67.14 2.2 67.31 2.37 ;
      RECT 66.66 2.78 66.83 2.95 ;
      RECT 66.42 1.94 66.59 2.11 ;
      RECT 66.18 2.5 66.35 2.67 ;
      RECT 66.18 3.06 66.35 3.23 ;
      RECT 65.7 2.5 65.87 2.67 ;
      RECT 65.46 3.62 65.63 3.79 ;
      RECT 65.42 1.94 65.59 2.11 ;
      RECT 65.22 2.78 65.39 2.95 ;
      RECT 64.98 3.62 65.15 3.79 ;
      RECT 64.74 3.06 64.91 3.23 ;
      RECT 64.26 2.5 64.43 2.67 ;
      RECT 64.02 1.94 64.19 2.11 ;
      RECT 64.02 3.62 64.19 3.79 ;
      RECT 63.54 3.06 63.71 3.23 ;
      RECT 63.3 2.5 63.47 2.67 ;
      RECT 63.06 3.34 63.23 3.51 ;
      RECT 62.82 2.78 62.99 2.95 ;
      RECT 62.13 1.94 62.3 2.11 ;
      RECT 62.13 3.34 62.3 3.51 ;
      RECT 60.495 7.805 60.665 7.975 ;
      RECT 60.125 2.765 60.295 2.935 ;
      RECT 60.125 5.955 60.295 6.125 ;
      RECT 59.505 0.915 59.675 1.085 ;
      RECT 59.505 2.395 59.675 2.565 ;
      RECT 59.505 6.325 59.675 6.495 ;
      RECT 59.505 7.805 59.675 7.975 ;
      RECT 59.135 2.765 59.305 2.935 ;
      RECT 59.135 5.955 59.305 6.125 ;
      RECT 58.145 2.03 58.315 2.2 ;
      RECT 58.145 6.69 58.315 6.86 ;
      RECT 57.715 0.92 57.885 1.09 ;
      RECT 57.715 1.66 57.885 1.83 ;
      RECT 57.715 7.06 57.885 7.23 ;
      RECT 57.715 7.8 57.885 7.97 ;
      RECT 57.34 2.4 57.51 2.57 ;
      RECT 57.34 6.32 57.51 6.49 ;
      RECT 54.28 2.78 54.45 2.95 ;
      RECT 54.04 1.94 54.21 2.11 ;
      RECT 54.04 3.62 54.21 3.79 ;
      RECT 53.8 2.5 53.97 2.67 ;
      RECT 53.8 3.06 53.97 3.23 ;
      RECT 53.32 2.78 53.49 2.95 ;
      RECT 53.08 1.94 53.25 2.11 ;
      RECT 52.84 2.5 53.01 2.67 ;
      RECT 52.63 3.34 52.8 3.51 ;
      RECT 52.53 6.69 52.7 6.86 ;
      RECT 52.36 2.78 52.53 2.95 ;
      RECT 52.1 7.06 52.27 7.23 ;
      RECT 52.1 7.8 52.27 7.97 ;
      RECT 52.09 3.62 52.26 3.79 ;
      RECT 51.88 2.2 52.05 2.37 ;
      RECT 51.4 2.78 51.57 2.95 ;
      RECT 51.16 1.94 51.33 2.11 ;
      RECT 50.92 2.5 51.09 2.67 ;
      RECT 50.92 3.06 51.09 3.23 ;
      RECT 50.44 2.5 50.61 2.67 ;
      RECT 50.2 3.62 50.37 3.79 ;
      RECT 50.16 1.94 50.33 2.11 ;
      RECT 49.96 2.78 50.13 2.95 ;
      RECT 49.72 3.62 49.89 3.79 ;
      RECT 49.48 3.06 49.65 3.23 ;
      RECT 49 2.5 49.17 2.67 ;
      RECT 48.76 1.94 48.93 2.11 ;
      RECT 48.76 3.62 48.93 3.79 ;
      RECT 48.28 3.06 48.45 3.23 ;
      RECT 48.04 2.5 48.21 2.67 ;
      RECT 47.8 3.34 47.97 3.51 ;
      RECT 47.56 2.78 47.73 2.95 ;
      RECT 46.87 1.94 47.04 2.11 ;
      RECT 46.87 3.34 47.04 3.51 ;
      RECT 45.235 7.805 45.405 7.975 ;
      RECT 44.865 2.765 45.035 2.935 ;
      RECT 44.865 5.955 45.035 6.125 ;
      RECT 44.245 0.915 44.415 1.085 ;
      RECT 44.245 2.395 44.415 2.565 ;
      RECT 44.245 6.325 44.415 6.495 ;
      RECT 44.245 7.805 44.415 7.975 ;
      RECT 43.875 2.765 44.045 2.935 ;
      RECT 43.875 5.955 44.045 6.125 ;
      RECT 42.885 2.03 43.055 2.2 ;
      RECT 42.885 6.69 43.055 6.86 ;
      RECT 42.455 0.92 42.625 1.09 ;
      RECT 42.455 1.66 42.625 1.83 ;
      RECT 42.455 7.06 42.625 7.23 ;
      RECT 42.455 7.8 42.625 7.97 ;
      RECT 42.08 2.4 42.25 2.57 ;
      RECT 42.08 6.32 42.25 6.49 ;
      RECT 39.02 2.78 39.19 2.95 ;
      RECT 38.78 1.94 38.95 2.11 ;
      RECT 38.78 3.62 38.95 3.79 ;
      RECT 38.54 2.5 38.71 2.67 ;
      RECT 38.54 3.06 38.71 3.23 ;
      RECT 38.06 2.78 38.23 2.95 ;
      RECT 37.82 1.94 37.99 2.11 ;
      RECT 37.58 2.5 37.75 2.67 ;
      RECT 37.37 3.34 37.54 3.51 ;
      RECT 37.27 6.69 37.44 6.86 ;
      RECT 37.1 2.78 37.27 2.95 ;
      RECT 36.84 7.06 37.01 7.23 ;
      RECT 36.84 7.8 37.01 7.97 ;
      RECT 36.83 3.62 37 3.79 ;
      RECT 36.62 2.2 36.79 2.37 ;
      RECT 36.14 2.78 36.31 2.95 ;
      RECT 35.9 1.94 36.07 2.11 ;
      RECT 35.66 2.5 35.83 2.67 ;
      RECT 35.66 3.06 35.83 3.23 ;
      RECT 35.18 2.5 35.35 2.67 ;
      RECT 34.94 3.62 35.11 3.79 ;
      RECT 34.9 1.94 35.07 2.11 ;
      RECT 34.7 2.78 34.87 2.95 ;
      RECT 34.46 3.62 34.63 3.79 ;
      RECT 34.22 3.06 34.39 3.23 ;
      RECT 33.74 2.5 33.91 2.67 ;
      RECT 33.5 1.94 33.67 2.11 ;
      RECT 33.5 3.62 33.67 3.79 ;
      RECT 33.02 3.06 33.19 3.23 ;
      RECT 32.78 2.5 32.95 2.67 ;
      RECT 32.54 3.34 32.71 3.51 ;
      RECT 32.3 2.78 32.47 2.95 ;
      RECT 31.61 1.94 31.78 2.11 ;
      RECT 31.61 3.34 31.78 3.51 ;
      RECT 29.975 7.805 30.145 7.975 ;
      RECT 29.605 2.765 29.775 2.935 ;
      RECT 29.605 5.955 29.775 6.125 ;
      RECT 28.985 0.915 29.155 1.085 ;
      RECT 28.985 2.395 29.155 2.565 ;
      RECT 28.985 6.325 29.155 6.495 ;
      RECT 28.985 7.805 29.155 7.975 ;
      RECT 28.615 2.765 28.785 2.935 ;
      RECT 28.615 5.955 28.785 6.125 ;
      RECT 27.625 2.03 27.795 2.2 ;
      RECT 27.625 6.69 27.795 6.86 ;
      RECT 27.195 0.92 27.365 1.09 ;
      RECT 27.195 1.66 27.365 1.83 ;
      RECT 27.195 7.06 27.365 7.23 ;
      RECT 27.195 7.8 27.365 7.97 ;
      RECT 26.82 2.4 26.99 2.57 ;
      RECT 26.82 6.32 26.99 6.49 ;
      RECT 23.76 2.78 23.93 2.95 ;
      RECT 23.52 1.94 23.69 2.11 ;
      RECT 23.52 3.62 23.69 3.79 ;
      RECT 23.28 2.5 23.45 2.67 ;
      RECT 23.28 3.06 23.45 3.23 ;
      RECT 22.8 2.78 22.97 2.95 ;
      RECT 22.56 1.94 22.73 2.11 ;
      RECT 22.32 2.5 22.49 2.67 ;
      RECT 22.11 3.34 22.28 3.51 ;
      RECT 22.01 6.69 22.18 6.86 ;
      RECT 21.84 2.78 22.01 2.95 ;
      RECT 21.58 7.06 21.75 7.23 ;
      RECT 21.58 7.8 21.75 7.97 ;
      RECT 21.57 3.62 21.74 3.79 ;
      RECT 21.36 2.2 21.53 2.37 ;
      RECT 20.88 2.78 21.05 2.95 ;
      RECT 20.64 1.94 20.81 2.11 ;
      RECT 20.4 2.5 20.57 2.67 ;
      RECT 20.4 3.06 20.57 3.23 ;
      RECT 19.92 2.5 20.09 2.67 ;
      RECT 19.68 3.62 19.85 3.79 ;
      RECT 19.64 1.94 19.81 2.11 ;
      RECT 19.44 2.78 19.61 2.95 ;
      RECT 19.2 3.62 19.37 3.79 ;
      RECT 18.96 3.06 19.13 3.23 ;
      RECT 18.48 2.5 18.65 2.67 ;
      RECT 18.24 1.94 18.41 2.11 ;
      RECT 18.24 3.62 18.41 3.79 ;
      RECT 17.76 3.06 17.93 3.23 ;
      RECT 17.52 2.5 17.69 2.67 ;
      RECT 17.28 3.34 17.45 3.51 ;
      RECT 17.04 2.78 17.21 2.95 ;
      RECT 16.35 1.94 16.52 2.11 ;
      RECT 16.35 3.34 16.52 3.51 ;
      RECT 14.715 7.805 14.885 7.975 ;
      RECT 14.345 2.765 14.515 2.935 ;
      RECT 14.345 5.955 14.515 6.125 ;
      RECT 13.725 0.915 13.895 1.085 ;
      RECT 13.725 2.395 13.895 2.565 ;
      RECT 13.725 6.325 13.895 6.495 ;
      RECT 13.725 7.805 13.895 7.975 ;
      RECT 13.355 2.765 13.525 2.935 ;
      RECT 13.355 5.955 13.525 6.125 ;
      RECT 12.365 2.03 12.535 2.2 ;
      RECT 12.365 6.69 12.535 6.86 ;
      RECT 11.935 0.92 12.105 1.09 ;
      RECT 11.935 1.66 12.105 1.83 ;
      RECT 11.935 7.06 12.105 7.23 ;
      RECT 11.935 7.8 12.105 7.97 ;
      RECT 11.56 2.4 11.73 2.57 ;
      RECT 11.56 6.32 11.73 6.49 ;
      RECT 8.5 2.78 8.67 2.95 ;
      RECT 8.26 1.94 8.43 2.11 ;
      RECT 8.26 3.62 8.43 3.79 ;
      RECT 8.02 2.5 8.19 2.67 ;
      RECT 8.02 3.06 8.19 3.23 ;
      RECT 7.54 2.78 7.71 2.95 ;
      RECT 7.3 1.94 7.47 2.11 ;
      RECT 7.06 2.5 7.23 2.67 ;
      RECT 6.85 3.34 7.02 3.51 ;
      RECT 6.75 6.69 6.92 6.86 ;
      RECT 6.58 2.78 6.75 2.95 ;
      RECT 6.32 7.06 6.49 7.23 ;
      RECT 6.32 7.8 6.49 7.97 ;
      RECT 6.31 3.62 6.48 3.79 ;
      RECT 6.1 2.2 6.27 2.37 ;
      RECT 5.62 2.78 5.79 2.95 ;
      RECT 5.38 1.94 5.55 2.11 ;
      RECT 5.14 2.5 5.31 2.67 ;
      RECT 5.14 3.06 5.31 3.23 ;
      RECT 4.66 2.5 4.83 2.67 ;
      RECT 4.42 3.62 4.59 3.79 ;
      RECT 4.38 1.94 4.55 2.11 ;
      RECT 4.18 2.78 4.35 2.95 ;
      RECT 3.94 3.62 4.11 3.79 ;
      RECT 3.7 3.06 3.87 3.23 ;
      RECT 3.22 2.5 3.39 2.67 ;
      RECT 2.98 1.94 3.15 2.11 ;
      RECT 2.98 3.62 3.15 3.79 ;
      RECT 2.5 3.06 2.67 3.23 ;
      RECT 2.26 2.5 2.43 2.67 ;
      RECT 2.02 3.34 2.19 3.51 ;
      RECT 1.78 2.78 1.95 2.95 ;
      RECT 1.09 1.94 1.26 2.11 ;
      RECT 1.09 3.34 1.26 3.51 ;
      RECT -1.195 7.06 -1.025 7.23 ;
      RECT -1.195 7.8 -1.025 7.97 ;
      RECT -1.57 6.32 -1.4 6.49 ;
    LAYER li1 ;
      RECT 75.755 5.025 75.925 6.495 ;
      RECT 75.755 6.32 75.93 6.49 ;
      RECT 75.385 1.745 75.555 2.935 ;
      RECT 75.385 1.745 75.855 1.915 ;
      RECT 75.385 6.975 75.855 7.145 ;
      RECT 75.385 5.955 75.555 7.145 ;
      RECT 74.395 1.745 74.565 2.935 ;
      RECT 74.395 1.745 74.865 1.915 ;
      RECT 74.395 6.975 74.865 7.145 ;
      RECT 74.395 5.955 74.565 7.145 ;
      RECT 72.545 2.64 72.715 3.87 ;
      RECT 72.6 0.86 72.77 2.81 ;
      RECT 72.545 0.58 72.715 1.03 ;
      RECT 72.545 7.86 72.715 8.31 ;
      RECT 72.6 6.08 72.77 8.03 ;
      RECT 72.545 5.02 72.715 6.25 ;
      RECT 72.025 0.58 72.195 3.87 ;
      RECT 72.025 2.08 72.43 2.41 ;
      RECT 72.025 1.24 72.43 1.57 ;
      RECT 72.025 5.02 72.195 8.31 ;
      RECT 72.025 7.32 72.43 7.65 ;
      RECT 72.025 6.48 72.43 6.81 ;
      RECT 69.3 3.62 69.815 3.79 ;
      RECT 69.645 3.23 69.815 3.79 ;
      RECT 69.75 3.15 69.92 3.48 ;
      RECT 69.54 2.54 69.815 2.95 ;
      RECT 69.42 2.54 69.815 2.75 ;
      RECT 67.89 3.15 68.06 3.51 ;
      RECT 67.89 3.23 69.23 3.4 ;
      RECT 69.06 3.06 69.23 3.4 ;
      RECT 67.62 2.58 67.79 2.95 ;
      RECT 67.14 2.58 67.79 2.85 ;
      RECT 67.06 2.58 67.87 2.75 ;
      RECT 66.42 1.82 66.59 2.11 ;
      RECT 66.42 1.82 67.66 1.99 ;
      RECT 67.14 2.16 67.31 2.37 ;
      RECT 66.78 2.16 67.31 2.33 ;
      RECT 66.41 5.02 66.58 8.31 ;
      RECT 66.41 7.32 66.815 7.65 ;
      RECT 66.41 6.48 66.815 6.81 ;
      RECT 66.18 3.23 66.67 3.4 ;
      RECT 66.18 3.06 66.35 3.4 ;
      RECT 65.46 3.23 65.63 3.79 ;
      RECT 65.35 3.23 65.68 3.4 ;
      RECT 65.42 1.84 65.59 2.11 ;
      RECT 65.46 1.76 65.63 2.09 ;
      RECT 65.325 1.84 65.63 2.06 ;
      RECT 63.9 3.23 64.19 3.79 ;
      RECT 64.02 3.15 64.19 3.79 ;
      RECT 60.495 5.025 60.665 6.495 ;
      RECT 60.495 6.32 60.67 6.49 ;
      RECT 60.125 1.745 60.295 2.935 ;
      RECT 60.125 1.745 60.595 1.915 ;
      RECT 60.125 6.975 60.595 7.145 ;
      RECT 60.125 5.955 60.295 7.145 ;
      RECT 59.135 1.745 59.305 2.935 ;
      RECT 59.135 1.745 59.605 1.915 ;
      RECT 59.135 6.975 59.605 7.145 ;
      RECT 59.135 5.955 59.305 7.145 ;
      RECT 57.285 2.64 57.455 3.87 ;
      RECT 57.34 0.86 57.51 2.81 ;
      RECT 57.285 0.58 57.455 1.03 ;
      RECT 57.285 7.86 57.455 8.31 ;
      RECT 57.34 6.08 57.51 8.03 ;
      RECT 57.285 5.02 57.455 6.25 ;
      RECT 56.765 0.58 56.935 3.87 ;
      RECT 56.765 2.08 57.17 2.41 ;
      RECT 56.765 1.24 57.17 1.57 ;
      RECT 56.765 5.02 56.935 8.31 ;
      RECT 56.765 7.32 57.17 7.65 ;
      RECT 56.765 6.48 57.17 6.81 ;
      RECT 54.04 3.62 54.555 3.79 ;
      RECT 54.385 3.23 54.555 3.79 ;
      RECT 54.49 3.15 54.66 3.48 ;
      RECT 54.28 2.54 54.555 2.95 ;
      RECT 54.16 2.54 54.555 2.75 ;
      RECT 52.63 3.15 52.8 3.51 ;
      RECT 52.63 3.23 53.97 3.4 ;
      RECT 53.8 3.06 53.97 3.4 ;
      RECT 52.36 2.58 52.53 2.95 ;
      RECT 51.88 2.58 52.53 2.85 ;
      RECT 51.8 2.58 52.61 2.75 ;
      RECT 51.16 1.82 51.33 2.11 ;
      RECT 51.16 1.82 52.4 1.99 ;
      RECT 51.88 2.16 52.05 2.37 ;
      RECT 51.52 2.16 52.05 2.33 ;
      RECT 51.15 5.02 51.32 8.31 ;
      RECT 51.15 7.32 51.555 7.65 ;
      RECT 51.15 6.48 51.555 6.81 ;
      RECT 50.92 3.23 51.41 3.4 ;
      RECT 50.92 3.06 51.09 3.4 ;
      RECT 50.2 3.23 50.37 3.79 ;
      RECT 50.09 3.23 50.42 3.4 ;
      RECT 50.16 1.84 50.33 2.11 ;
      RECT 50.2 1.76 50.37 2.09 ;
      RECT 50.065 1.84 50.37 2.06 ;
      RECT 48.64 3.23 48.93 3.79 ;
      RECT 48.76 3.15 48.93 3.79 ;
      RECT 45.235 5.025 45.405 6.495 ;
      RECT 45.235 6.32 45.41 6.49 ;
      RECT 44.865 1.745 45.035 2.935 ;
      RECT 44.865 1.745 45.335 1.915 ;
      RECT 44.865 6.975 45.335 7.145 ;
      RECT 44.865 5.955 45.035 7.145 ;
      RECT 43.875 1.745 44.045 2.935 ;
      RECT 43.875 1.745 44.345 1.915 ;
      RECT 43.875 6.975 44.345 7.145 ;
      RECT 43.875 5.955 44.045 7.145 ;
      RECT 42.025 2.64 42.195 3.87 ;
      RECT 42.08 0.86 42.25 2.81 ;
      RECT 42.025 0.58 42.195 1.03 ;
      RECT 42.025 7.86 42.195 8.31 ;
      RECT 42.08 6.08 42.25 8.03 ;
      RECT 42.025 5.02 42.195 6.25 ;
      RECT 41.505 0.58 41.675 3.87 ;
      RECT 41.505 2.08 41.91 2.41 ;
      RECT 41.505 1.24 41.91 1.57 ;
      RECT 41.505 5.02 41.675 8.31 ;
      RECT 41.505 7.32 41.91 7.65 ;
      RECT 41.505 6.48 41.91 6.81 ;
      RECT 38.78 3.62 39.295 3.79 ;
      RECT 39.125 3.23 39.295 3.79 ;
      RECT 39.23 3.15 39.4 3.48 ;
      RECT 39.02 2.54 39.295 2.95 ;
      RECT 38.9 2.54 39.295 2.75 ;
      RECT 37.37 3.15 37.54 3.51 ;
      RECT 37.37 3.23 38.71 3.4 ;
      RECT 38.54 3.06 38.71 3.4 ;
      RECT 37.1 2.58 37.27 2.95 ;
      RECT 36.62 2.58 37.27 2.85 ;
      RECT 36.54 2.58 37.35 2.75 ;
      RECT 35.9 1.82 36.07 2.11 ;
      RECT 35.9 1.82 37.14 1.99 ;
      RECT 36.62 2.16 36.79 2.37 ;
      RECT 36.26 2.16 36.79 2.33 ;
      RECT 35.89 5.02 36.06 8.31 ;
      RECT 35.89 7.32 36.295 7.65 ;
      RECT 35.89 6.48 36.295 6.81 ;
      RECT 35.66 3.23 36.15 3.4 ;
      RECT 35.66 3.06 35.83 3.4 ;
      RECT 34.94 3.23 35.11 3.79 ;
      RECT 34.83 3.23 35.16 3.4 ;
      RECT 34.9 1.84 35.07 2.11 ;
      RECT 34.94 1.76 35.11 2.09 ;
      RECT 34.805 1.84 35.11 2.06 ;
      RECT 33.38 3.23 33.67 3.79 ;
      RECT 33.5 3.15 33.67 3.79 ;
      RECT 29.975 5.025 30.145 6.495 ;
      RECT 29.975 6.32 30.15 6.49 ;
      RECT 29.605 1.745 29.775 2.935 ;
      RECT 29.605 1.745 30.075 1.915 ;
      RECT 29.605 6.975 30.075 7.145 ;
      RECT 29.605 5.955 29.775 7.145 ;
      RECT 28.615 1.745 28.785 2.935 ;
      RECT 28.615 1.745 29.085 1.915 ;
      RECT 28.615 6.975 29.085 7.145 ;
      RECT 28.615 5.955 28.785 7.145 ;
      RECT 26.765 2.64 26.935 3.87 ;
      RECT 26.82 0.86 26.99 2.81 ;
      RECT 26.765 0.58 26.935 1.03 ;
      RECT 26.765 7.86 26.935 8.31 ;
      RECT 26.82 6.08 26.99 8.03 ;
      RECT 26.765 5.02 26.935 6.25 ;
      RECT 26.245 0.58 26.415 3.87 ;
      RECT 26.245 2.08 26.65 2.41 ;
      RECT 26.245 1.24 26.65 1.57 ;
      RECT 26.245 5.02 26.415 8.31 ;
      RECT 26.245 7.32 26.65 7.65 ;
      RECT 26.245 6.48 26.65 6.81 ;
      RECT 23.52 3.62 24.035 3.79 ;
      RECT 23.865 3.23 24.035 3.79 ;
      RECT 23.97 3.15 24.14 3.48 ;
      RECT 23.76 2.54 24.035 2.95 ;
      RECT 23.64 2.54 24.035 2.75 ;
      RECT 22.11 3.15 22.28 3.51 ;
      RECT 22.11 3.23 23.45 3.4 ;
      RECT 23.28 3.06 23.45 3.4 ;
      RECT 21.84 2.58 22.01 2.95 ;
      RECT 21.36 2.58 22.01 2.85 ;
      RECT 21.28 2.58 22.09 2.75 ;
      RECT 20.64 1.82 20.81 2.11 ;
      RECT 20.64 1.82 21.88 1.99 ;
      RECT 21.36 2.16 21.53 2.37 ;
      RECT 21 2.16 21.53 2.33 ;
      RECT 20.63 5.02 20.8 8.31 ;
      RECT 20.63 7.32 21.035 7.65 ;
      RECT 20.63 6.48 21.035 6.81 ;
      RECT 20.4 3.23 20.89 3.4 ;
      RECT 20.4 3.06 20.57 3.4 ;
      RECT 19.68 3.23 19.85 3.79 ;
      RECT 19.57 3.23 19.9 3.4 ;
      RECT 19.64 1.84 19.81 2.11 ;
      RECT 19.68 1.76 19.85 2.09 ;
      RECT 19.545 1.84 19.85 2.06 ;
      RECT 18.12 3.23 18.41 3.79 ;
      RECT 18.24 3.15 18.41 3.79 ;
      RECT 14.715 5.025 14.885 6.495 ;
      RECT 14.715 6.32 14.89 6.49 ;
      RECT 14.345 1.745 14.515 2.935 ;
      RECT 14.345 1.745 14.815 1.915 ;
      RECT 14.345 6.975 14.815 7.145 ;
      RECT 14.345 5.955 14.515 7.145 ;
      RECT 13.355 1.745 13.525 2.935 ;
      RECT 13.355 1.745 13.825 1.915 ;
      RECT 13.355 6.975 13.825 7.145 ;
      RECT 13.355 5.955 13.525 7.145 ;
      RECT 11.505 2.64 11.675 3.87 ;
      RECT 11.56 0.86 11.73 2.81 ;
      RECT 11.505 0.58 11.675 1.03 ;
      RECT 11.505 7.86 11.675 8.31 ;
      RECT 11.56 6.08 11.73 8.03 ;
      RECT 11.505 5.02 11.675 6.25 ;
      RECT 10.985 0.58 11.155 3.87 ;
      RECT 10.985 2.08 11.39 2.41 ;
      RECT 10.985 1.24 11.39 1.57 ;
      RECT 10.985 5.02 11.155 8.31 ;
      RECT 10.985 7.32 11.39 7.65 ;
      RECT 10.985 6.48 11.39 6.81 ;
      RECT 8.26 3.62 8.775 3.79 ;
      RECT 8.605 3.23 8.775 3.79 ;
      RECT 8.71 3.15 8.88 3.48 ;
      RECT 8.5 2.54 8.775 2.95 ;
      RECT 8.38 2.54 8.775 2.75 ;
      RECT 6.85 3.15 7.02 3.51 ;
      RECT 6.85 3.23 8.19 3.4 ;
      RECT 8.02 3.06 8.19 3.4 ;
      RECT 6.58 2.58 6.75 2.95 ;
      RECT 6.1 2.58 6.75 2.85 ;
      RECT 6.02 2.58 6.83 2.75 ;
      RECT 5.38 1.82 5.55 2.11 ;
      RECT 5.38 1.82 6.62 1.99 ;
      RECT 6.1 2.16 6.27 2.37 ;
      RECT 5.74 2.16 6.27 2.33 ;
      RECT 5.37 5.02 5.54 8.31 ;
      RECT 5.37 7.32 5.775 7.65 ;
      RECT 5.37 6.48 5.775 6.81 ;
      RECT 5.14 3.23 5.63 3.4 ;
      RECT 5.14 3.06 5.31 3.4 ;
      RECT 4.42 3.23 4.59 3.79 ;
      RECT 4.31 3.23 4.64 3.4 ;
      RECT 4.38 1.84 4.55 2.11 ;
      RECT 4.42 1.76 4.59 2.09 ;
      RECT 4.285 1.84 4.59 2.06 ;
      RECT 2.86 3.23 3.15 3.79 ;
      RECT 2.98 3.15 3.15 3.79 ;
      RECT -1.625 7.86 -1.455 8.31 ;
      RECT -1.57 6.08 -1.4 8.03 ;
      RECT -1.625 5.02 -1.455 6.25 ;
      RECT -2.145 5.02 -1.975 8.31 ;
      RECT -2.145 7.32 -1.74 7.65 ;
      RECT -2.145 6.48 -1.74 6.81 ;
      RECT 75.755 7.805 75.925 8.315 ;
      RECT 74.765 0.575 74.935 1.085 ;
      RECT 74.765 2.395 74.935 3.865 ;
      RECT 74.765 5.025 74.935 6.495 ;
      RECT 74.765 7.805 74.935 8.315 ;
      RECT 73.405 0.58 73.575 3.87 ;
      RECT 73.405 5.02 73.575 8.31 ;
      RECT 72.975 0.58 73.145 1.09 ;
      RECT 72.975 1.66 73.145 3.87 ;
      RECT 72.975 5.02 73.145 7.23 ;
      RECT 72.975 7.8 73.145 8.31 ;
      RECT 69.3 1.76 69.47 2.11 ;
      RECT 69.06 2.5 69.23 2.83 ;
      RECT 68.58 2.5 68.75 2.95 ;
      RECT 68.34 1.76 68.51 2.11 ;
      RECT 68.1 2.5 68.27 2.83 ;
      RECT 67.79 5.02 67.96 8.31 ;
      RECT 67.36 5.02 67.53 7.23 ;
      RECT 67.36 7.8 67.53 8.31 ;
      RECT 67.35 3.49 67.52 3.82 ;
      RECT 66.66 2.5 66.83 2.95 ;
      RECT 66.18 2.5 66.35 2.83 ;
      RECT 65.7 2.5 65.87 2.83 ;
      RECT 65.22 2.5 65.39 2.95 ;
      RECT 64.98 3.49 65.15 3.82 ;
      RECT 64.74 2.5 64.91 3.23 ;
      RECT 64.26 2.5 64.43 2.83 ;
      RECT 64.02 1.76 64.19 2.11 ;
      RECT 63.54 3.06 63.71 3.48 ;
      RECT 63.3 2.5 63.47 2.83 ;
      RECT 63.06 3.15 63.23 3.51 ;
      RECT 62.82 2.5 62.99 2.95 ;
      RECT 62.13 1.76 62.3 2.11 ;
      RECT 62.13 3.15 62.3 3.51 ;
      RECT 60.495 7.805 60.665 8.315 ;
      RECT 59.505 0.575 59.675 1.085 ;
      RECT 59.505 2.395 59.675 3.865 ;
      RECT 59.505 5.025 59.675 6.495 ;
      RECT 59.505 7.805 59.675 8.315 ;
      RECT 58.145 0.58 58.315 3.87 ;
      RECT 58.145 5.02 58.315 8.31 ;
      RECT 57.715 0.58 57.885 1.09 ;
      RECT 57.715 1.66 57.885 3.87 ;
      RECT 57.715 5.02 57.885 7.23 ;
      RECT 57.715 7.8 57.885 8.31 ;
      RECT 54.04 1.76 54.21 2.11 ;
      RECT 53.8 2.5 53.97 2.83 ;
      RECT 53.32 2.5 53.49 2.95 ;
      RECT 53.08 1.76 53.25 2.11 ;
      RECT 52.84 2.5 53.01 2.83 ;
      RECT 52.53 5.02 52.7 8.31 ;
      RECT 52.1 5.02 52.27 7.23 ;
      RECT 52.1 7.8 52.27 8.31 ;
      RECT 52.09 3.49 52.26 3.82 ;
      RECT 51.4 2.5 51.57 2.95 ;
      RECT 50.92 2.5 51.09 2.83 ;
      RECT 50.44 2.5 50.61 2.83 ;
      RECT 49.96 2.5 50.13 2.95 ;
      RECT 49.72 3.49 49.89 3.82 ;
      RECT 49.48 2.5 49.65 3.23 ;
      RECT 49 2.5 49.17 2.83 ;
      RECT 48.76 1.76 48.93 2.11 ;
      RECT 48.28 3.06 48.45 3.48 ;
      RECT 48.04 2.5 48.21 2.83 ;
      RECT 47.8 3.15 47.97 3.51 ;
      RECT 47.56 2.5 47.73 2.95 ;
      RECT 46.87 1.76 47.04 2.11 ;
      RECT 46.87 3.15 47.04 3.51 ;
      RECT 45.235 7.805 45.405 8.315 ;
      RECT 44.245 0.575 44.415 1.085 ;
      RECT 44.245 2.395 44.415 3.865 ;
      RECT 44.245 5.025 44.415 6.495 ;
      RECT 44.245 7.805 44.415 8.315 ;
      RECT 42.885 0.58 43.055 3.87 ;
      RECT 42.885 5.02 43.055 8.31 ;
      RECT 42.455 0.58 42.625 1.09 ;
      RECT 42.455 1.66 42.625 3.87 ;
      RECT 42.455 5.02 42.625 7.23 ;
      RECT 42.455 7.8 42.625 8.31 ;
      RECT 38.78 1.76 38.95 2.11 ;
      RECT 38.54 2.5 38.71 2.83 ;
      RECT 38.06 2.5 38.23 2.95 ;
      RECT 37.82 1.76 37.99 2.11 ;
      RECT 37.58 2.5 37.75 2.83 ;
      RECT 37.27 5.02 37.44 8.31 ;
      RECT 36.84 5.02 37.01 7.23 ;
      RECT 36.84 7.8 37.01 8.31 ;
      RECT 36.83 3.49 37 3.82 ;
      RECT 36.14 2.5 36.31 2.95 ;
      RECT 35.66 2.5 35.83 2.83 ;
      RECT 35.18 2.5 35.35 2.83 ;
      RECT 34.7 2.5 34.87 2.95 ;
      RECT 34.46 3.49 34.63 3.82 ;
      RECT 34.22 2.5 34.39 3.23 ;
      RECT 33.74 2.5 33.91 2.83 ;
      RECT 33.5 1.76 33.67 2.11 ;
      RECT 33.02 3.06 33.19 3.48 ;
      RECT 32.78 2.5 32.95 2.83 ;
      RECT 32.54 3.15 32.71 3.51 ;
      RECT 32.3 2.5 32.47 2.95 ;
      RECT 31.61 1.76 31.78 2.11 ;
      RECT 31.61 3.15 31.78 3.51 ;
      RECT 29.975 7.805 30.145 8.315 ;
      RECT 28.985 0.575 29.155 1.085 ;
      RECT 28.985 2.395 29.155 3.865 ;
      RECT 28.985 5.025 29.155 6.495 ;
      RECT 28.985 7.805 29.155 8.315 ;
      RECT 27.625 0.58 27.795 3.87 ;
      RECT 27.625 5.02 27.795 8.31 ;
      RECT 27.195 0.58 27.365 1.09 ;
      RECT 27.195 1.66 27.365 3.87 ;
      RECT 27.195 5.02 27.365 7.23 ;
      RECT 27.195 7.8 27.365 8.31 ;
      RECT 23.52 1.76 23.69 2.11 ;
      RECT 23.28 2.5 23.45 2.83 ;
      RECT 22.8 2.5 22.97 2.95 ;
      RECT 22.56 1.76 22.73 2.11 ;
      RECT 22.32 2.5 22.49 2.83 ;
      RECT 22.01 5.02 22.18 8.31 ;
      RECT 21.58 5.02 21.75 7.23 ;
      RECT 21.58 7.8 21.75 8.31 ;
      RECT 21.57 3.49 21.74 3.82 ;
      RECT 20.88 2.5 21.05 2.95 ;
      RECT 20.4 2.5 20.57 2.83 ;
      RECT 19.92 2.5 20.09 2.83 ;
      RECT 19.44 2.5 19.61 2.95 ;
      RECT 19.2 3.49 19.37 3.82 ;
      RECT 18.96 2.5 19.13 3.23 ;
      RECT 18.48 2.5 18.65 2.83 ;
      RECT 18.24 1.76 18.41 2.11 ;
      RECT 17.76 3.06 17.93 3.48 ;
      RECT 17.52 2.5 17.69 2.83 ;
      RECT 17.28 3.15 17.45 3.51 ;
      RECT 17.04 2.5 17.21 2.95 ;
      RECT 16.35 1.76 16.52 2.11 ;
      RECT 16.35 3.15 16.52 3.51 ;
      RECT 14.715 7.805 14.885 8.315 ;
      RECT 13.725 0.575 13.895 1.085 ;
      RECT 13.725 2.395 13.895 3.865 ;
      RECT 13.725 5.025 13.895 6.495 ;
      RECT 13.725 7.805 13.895 8.315 ;
      RECT 12.365 0.58 12.535 3.87 ;
      RECT 12.365 5.02 12.535 8.31 ;
      RECT 11.935 0.58 12.105 1.09 ;
      RECT 11.935 1.66 12.105 3.87 ;
      RECT 11.935 5.02 12.105 7.23 ;
      RECT 11.935 7.8 12.105 8.31 ;
      RECT 8.26 1.76 8.43 2.11 ;
      RECT 8.02 2.5 8.19 2.83 ;
      RECT 7.54 2.5 7.71 2.95 ;
      RECT 7.3 1.76 7.47 2.11 ;
      RECT 7.06 2.5 7.23 2.83 ;
      RECT 6.75 5.02 6.92 8.31 ;
      RECT 6.32 5.02 6.49 7.23 ;
      RECT 6.32 7.8 6.49 8.31 ;
      RECT 6.31 3.49 6.48 3.82 ;
      RECT 5.62 2.5 5.79 2.95 ;
      RECT 5.14 2.5 5.31 2.83 ;
      RECT 4.66 2.5 4.83 2.83 ;
      RECT 4.18 2.5 4.35 2.95 ;
      RECT 3.94 3.49 4.11 3.82 ;
      RECT 3.7 2.5 3.87 3.23 ;
      RECT 3.22 2.5 3.39 2.83 ;
      RECT 2.98 1.76 3.15 2.11 ;
      RECT 2.5 3.06 2.67 3.48 ;
      RECT 2.26 2.5 2.43 2.83 ;
      RECT 2.02 3.15 2.19 3.51 ;
      RECT 1.78 2.5 1.95 2.95 ;
      RECT 1.09 1.76 1.26 2.11 ;
      RECT 1.09 3.15 1.26 3.51 ;
      RECT -1.195 5.02 -1.025 7.23 ;
      RECT -1.195 7.8 -1.025 8.31 ;
  END
END sky130_osu_ring_oscillator_mpr2xa_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2xa_8_b0r2
  CLASS BLOCK ;
  ORIGIN 2.795 -0.005 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2xa_8_b0r2 ;
  SIZE 79.095 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 14.72 0.92 14.89 1.09 ;
        RECT 14.715 0.915 14.885 1.085 ;
        RECT 14.715 2.395 14.885 2.565 ;
      LAYER li1 ;
        RECT 14.72 0.92 14.89 1.09 ;
        RECT 14.715 0.575 14.885 1.085 ;
        RECT 14.715 2.395 14.885 3.865 ;
      LAYER met1 ;
        RECT 14.655 2.365 14.945 2.595 ;
        RECT 14.655 0.885 14.945 1.115 ;
        RECT 14.715 0.885 14.885 2.595 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 29.98 0.92 30.15 1.09 ;
        RECT 29.975 0.915 30.145 1.085 ;
        RECT 29.975 2.395 30.145 2.565 ;
      LAYER li1 ;
        RECT 29.98 0.92 30.15 1.09 ;
        RECT 29.975 0.575 30.145 1.085 ;
        RECT 29.975 2.395 30.145 3.865 ;
      LAYER met1 ;
        RECT 29.915 2.365 30.205 2.595 ;
        RECT 29.915 0.885 30.205 1.115 ;
        RECT 29.975 0.885 30.145 2.595 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 45.24 0.92 45.41 1.09 ;
        RECT 45.235 0.915 45.405 1.085 ;
        RECT 45.235 2.395 45.405 2.565 ;
      LAYER li1 ;
        RECT 45.24 0.92 45.41 1.09 ;
        RECT 45.235 0.575 45.405 1.085 ;
        RECT 45.235 2.395 45.405 3.865 ;
      LAYER met1 ;
        RECT 45.175 2.365 45.465 2.595 ;
        RECT 45.175 0.885 45.465 1.115 ;
        RECT 45.235 0.885 45.405 2.595 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 60.5 0.92 60.67 1.09 ;
        RECT 60.495 0.915 60.665 1.085 ;
        RECT 60.495 2.395 60.665 2.565 ;
      LAYER li1 ;
        RECT 60.5 0.92 60.67 1.09 ;
        RECT 60.495 0.575 60.665 1.085 ;
        RECT 60.495 2.395 60.665 3.865 ;
      LAYER met1 ;
        RECT 60.435 2.365 60.725 2.595 ;
        RECT 60.435 0.885 60.725 1.115 ;
        RECT 60.495 0.885 60.665 2.595 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 75.76 0.92 75.93 1.09 ;
        RECT 75.755 0.915 75.925 1.085 ;
        RECT 75.755 2.395 75.925 2.565 ;
      LAYER li1 ;
        RECT 75.76 0.92 75.93 1.09 ;
        RECT 75.755 0.575 75.925 1.085 ;
        RECT 75.755 2.395 75.925 3.865 ;
      LAYER met1 ;
        RECT 75.695 2.365 75.985 2.595 ;
        RECT 75.695 0.885 75.985 1.115 ;
        RECT 75.755 0.885 75.925 2.595 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 10.485 5.865 10.825 6.215 ;
        RECT 10.485 2.71 10.825 3.06 ;
        RECT 10.565 2.71 10.735 6.215 ;
      LAYER li1 ;
        RECT 10.565 1.665 10.735 2.94 ;
        RECT 10.565 5.95 10.735 7.225 ;
        RECT 4.95 5.95 5.12 7.225 ;
      LAYER met1 ;
        RECT 10.485 2.77 10.965 2.94 ;
        RECT 10.485 2.71 10.825 3.06 ;
        RECT 4.89 5.95 10.965 6.12 ;
        RECT 10.485 5.865 10.825 6.215 ;
        RECT 4.89 5.92 5.18 6.15 ;
      LAYER via1 ;
        RECT 10.585 5.965 10.735 6.115 ;
        RECT 10.585 2.81 10.735 2.96 ;
      LAYER mcon ;
        RECT 4.95 5.95 5.12 6.12 ;
        RECT 10.565 5.95 10.735 6.12 ;
        RECT 10.565 2.77 10.735 2.94 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 25.745 5.865 26.085 6.215 ;
        RECT 25.745 2.71 26.085 3.06 ;
        RECT 25.825 2.71 25.995 6.215 ;
      LAYER li1 ;
        RECT 25.825 1.665 25.995 2.94 ;
        RECT 25.825 5.95 25.995 7.225 ;
        RECT 20.21 5.95 20.38 7.225 ;
      LAYER met1 ;
        RECT 25.745 2.77 26.225 2.94 ;
        RECT 25.745 2.71 26.085 3.06 ;
        RECT 20.15 5.95 26.225 6.12 ;
        RECT 25.745 5.865 26.085 6.215 ;
        RECT 20.15 5.92 20.44 6.15 ;
      LAYER via1 ;
        RECT 25.845 5.965 25.995 6.115 ;
        RECT 25.845 2.81 25.995 2.96 ;
      LAYER mcon ;
        RECT 20.21 5.95 20.38 6.12 ;
        RECT 25.825 5.95 25.995 6.12 ;
        RECT 25.825 2.77 25.995 2.94 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 41.005 5.865 41.345 6.215 ;
        RECT 41.005 2.71 41.345 3.06 ;
        RECT 41.085 2.71 41.255 6.215 ;
      LAYER li1 ;
        RECT 41.085 1.665 41.255 2.94 ;
        RECT 41.085 5.95 41.255 7.225 ;
        RECT 35.47 5.95 35.64 7.225 ;
      LAYER met1 ;
        RECT 41.005 2.77 41.485 2.94 ;
        RECT 41.005 2.71 41.345 3.06 ;
        RECT 35.41 5.95 41.485 6.12 ;
        RECT 41.005 5.865 41.345 6.215 ;
        RECT 35.41 5.92 35.7 6.15 ;
      LAYER via1 ;
        RECT 41.105 5.965 41.255 6.115 ;
        RECT 41.105 2.81 41.255 2.96 ;
      LAYER mcon ;
        RECT 35.47 5.95 35.64 6.12 ;
        RECT 41.085 5.95 41.255 6.12 ;
        RECT 41.085 2.77 41.255 2.94 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 56.265 5.865 56.605 6.215 ;
        RECT 56.265 2.71 56.605 3.06 ;
        RECT 56.345 2.71 56.515 6.215 ;
      LAYER li1 ;
        RECT 56.345 1.665 56.515 2.94 ;
        RECT 56.345 5.95 56.515 7.225 ;
        RECT 50.73 5.95 50.9 7.225 ;
      LAYER met1 ;
        RECT 56.265 2.77 56.745 2.94 ;
        RECT 56.265 2.71 56.605 3.06 ;
        RECT 50.67 5.95 56.745 6.12 ;
        RECT 56.265 5.865 56.605 6.215 ;
        RECT 50.67 5.92 50.96 6.15 ;
      LAYER via1 ;
        RECT 56.365 5.965 56.515 6.115 ;
        RECT 56.365 2.81 56.515 2.96 ;
      LAYER mcon ;
        RECT 50.73 5.95 50.9 6.12 ;
        RECT 56.345 5.95 56.515 6.12 ;
        RECT 56.345 2.77 56.515 2.94 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 71.525 5.865 71.865 6.215 ;
        RECT 71.525 2.71 71.865 3.06 ;
        RECT 71.605 2.71 71.775 6.215 ;
      LAYER li1 ;
        RECT 71.605 1.665 71.775 2.94 ;
        RECT 71.605 5.95 71.775 7.225 ;
        RECT 65.99 5.95 66.16 7.225 ;
      LAYER met1 ;
        RECT 71.525 2.77 72.005 2.94 ;
        RECT 71.525 2.71 71.865 3.06 ;
        RECT 65.93 5.95 72.005 6.12 ;
        RECT 71.525 5.865 71.865 6.215 ;
        RECT 65.93 5.92 66.22 6.15 ;
      LAYER via1 ;
        RECT 71.625 5.965 71.775 6.115 ;
        RECT 71.625 2.81 71.775 2.96 ;
      LAYER mcon ;
        RECT 65.99 5.95 66.16 6.12 ;
        RECT 71.605 5.95 71.775 6.12 ;
        RECT 71.605 2.77 71.775 2.94 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT -2.565 5.95 -2.395 7.225 ;
      LAYER met1 ;
        RECT -2.625 5.95 -2.165 6.12 ;
        RECT -2.625 5.92 -2.335 6.15 ;
      LAYER mcon ;
        RECT -2.565 5.95 -2.395 6.12 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT -2.795 4.145 76.3 4.75 ;
        RECT 61.79 4.14 76.3 4.75 ;
        RECT 74.165 4.135 76.145 4.755 ;
        RECT 75.325 3.405 75.495 5.485 ;
        RECT 74.335 3.405 74.505 5.485 ;
        RECT 71.595 3.41 71.765 5.48 ;
        RECT 68.82 3.64 68.99 4.75 ;
        RECT 66.9 3.64 67.07 4.75 ;
        RECT 65.98 4.14 66.15 5.48 ;
        RECT 65.96 3.64 66.13 4.75 ;
        RECT 64.5 3.64 64.67 4.75 ;
        RECT 62.58 3.64 62.75 4.75 ;
        RECT 46.53 4.14 61.04 4.75 ;
        RECT 58.905 4.135 60.885 4.755 ;
        RECT 60.065 3.405 60.235 5.485 ;
        RECT 59.075 3.405 59.245 5.485 ;
        RECT 56.335 3.41 56.505 5.48 ;
        RECT 53.56 3.64 53.73 4.75 ;
        RECT 51.64 3.64 51.81 4.75 ;
        RECT 50.72 4.14 50.89 5.48 ;
        RECT 50.7 3.64 50.87 4.75 ;
        RECT 49.24 3.64 49.41 4.75 ;
        RECT 47.32 3.64 47.49 4.75 ;
        RECT 31.27 4.14 45.78 4.75 ;
        RECT 43.645 4.135 45.625 4.755 ;
        RECT 44.805 3.405 44.975 5.485 ;
        RECT 43.815 3.405 43.985 5.485 ;
        RECT 41.075 3.41 41.245 5.48 ;
        RECT 38.3 3.64 38.47 4.75 ;
        RECT 36.38 3.64 36.55 4.75 ;
        RECT 35.46 4.14 35.63 5.48 ;
        RECT 35.44 3.64 35.61 4.75 ;
        RECT 33.98 3.64 34.15 4.75 ;
        RECT 32.06 3.64 32.23 4.75 ;
        RECT 16.01 4.14 30.52 4.75 ;
        RECT 28.385 4.135 30.365 4.755 ;
        RECT 29.545 3.405 29.715 5.485 ;
        RECT 28.555 3.405 28.725 5.485 ;
        RECT 25.815 3.41 25.985 5.48 ;
        RECT 23.04 3.64 23.21 4.75 ;
        RECT 21.12 3.64 21.29 4.75 ;
        RECT 20.2 4.14 20.37 5.48 ;
        RECT 20.18 3.64 20.35 4.75 ;
        RECT 18.72 3.64 18.89 4.75 ;
        RECT 16.8 3.64 16.97 4.75 ;
        RECT 0.75 4.14 15.26 4.75 ;
        RECT 13.125 4.135 15.105 4.755 ;
        RECT 14.285 3.405 14.455 5.485 ;
        RECT 13.295 3.405 13.465 5.485 ;
        RECT 10.555 3.41 10.725 5.48 ;
        RECT 7.78 3.64 7.95 4.75 ;
        RECT 5.86 3.64 6.03 4.75 ;
        RECT 4.94 4.14 5.11 5.48 ;
        RECT 4.92 3.64 5.09 4.75 ;
        RECT 3.46 3.64 3.63 4.75 ;
        RECT 1.54 3.64 1.71 4.75 ;
        RECT -0.765 4.145 -0.595 8.31 ;
        RECT -2.575 4.145 -2.405 5.48 ;
      LAYER met1 ;
        RECT -2.795 4.145 76.3 4.75 ;
        RECT 61.79 4.14 76.3 4.75 ;
        RECT 74.165 4.135 76.145 4.755 ;
        RECT 61.79 3.985 70.53 4.75 ;
        RECT 46.53 4.14 61.04 4.75 ;
        RECT 58.905 4.135 60.885 4.755 ;
        RECT 46.53 3.985 55.27 4.75 ;
        RECT 31.27 4.14 45.78 4.75 ;
        RECT 43.645 4.135 45.625 4.755 ;
        RECT 31.27 3.985 40.01 4.75 ;
        RECT 16.01 4.14 30.52 4.75 ;
        RECT 28.385 4.135 30.365 4.755 ;
        RECT 16.01 3.985 24.75 4.75 ;
        RECT 0.75 4.14 15.26 4.75 ;
        RECT 13.125 4.135 15.105 4.755 ;
        RECT 0.75 3.985 9.49 4.75 ;
        RECT -0.825 6.66 -0.535 6.89 ;
        RECT -0.995 6.69 -0.535 6.86 ;
      LAYER mcon ;
        RECT -0.765 6.69 -0.595 6.86 ;
        RECT -0.455 4.55 -0.285 4.72 ;
        RECT 0.895 4.14 1.065 4.31 ;
        RECT 1.355 4.14 1.525 4.31 ;
        RECT 1.815 4.14 1.985 4.31 ;
        RECT 2.275 4.14 2.445 4.31 ;
        RECT 2.735 4.14 2.905 4.31 ;
        RECT 3.195 4.14 3.365 4.31 ;
        RECT 3.655 4.14 3.825 4.31 ;
        RECT 4.115 4.14 4.285 4.31 ;
        RECT 4.575 4.14 4.745 4.31 ;
        RECT 5.035 4.14 5.205 4.31 ;
        RECT 5.495 4.14 5.665 4.31 ;
        RECT 5.955 4.14 6.125 4.31 ;
        RECT 6.415 4.14 6.585 4.31 ;
        RECT 6.875 4.14 7.045 4.31 ;
        RECT 7.06 4.55 7.23 4.72 ;
        RECT 7.335 4.14 7.505 4.31 ;
        RECT 7.795 4.14 7.965 4.31 ;
        RECT 8.255 4.14 8.425 4.31 ;
        RECT 8.715 4.14 8.885 4.31 ;
        RECT 9.175 4.14 9.345 4.31 ;
        RECT 12.675 4.55 12.845 4.72 ;
        RECT 12.675 4.17 12.845 4.34 ;
        RECT 13.375 4.555 13.545 4.725 ;
        RECT 13.375 4.165 13.545 4.335 ;
        RECT 14.365 4.555 14.535 4.725 ;
        RECT 14.365 4.165 14.535 4.335 ;
        RECT 16.155 4.14 16.325 4.31 ;
        RECT 16.615 4.14 16.785 4.31 ;
        RECT 17.075 4.14 17.245 4.31 ;
        RECT 17.535 4.14 17.705 4.31 ;
        RECT 17.995 4.14 18.165 4.31 ;
        RECT 18.455 4.14 18.625 4.31 ;
        RECT 18.915 4.14 19.085 4.31 ;
        RECT 19.375 4.14 19.545 4.31 ;
        RECT 19.835 4.14 20.005 4.31 ;
        RECT 20.295 4.14 20.465 4.31 ;
        RECT 20.755 4.14 20.925 4.31 ;
        RECT 21.215 4.14 21.385 4.31 ;
        RECT 21.675 4.14 21.845 4.31 ;
        RECT 22.135 4.14 22.305 4.31 ;
        RECT 22.32 4.55 22.49 4.72 ;
        RECT 22.595 4.14 22.765 4.31 ;
        RECT 23.055 4.14 23.225 4.31 ;
        RECT 23.515 4.14 23.685 4.31 ;
        RECT 23.975 4.14 24.145 4.31 ;
        RECT 24.435 4.14 24.605 4.31 ;
        RECT 27.935 4.55 28.105 4.72 ;
        RECT 27.935 4.17 28.105 4.34 ;
        RECT 28.635 4.555 28.805 4.725 ;
        RECT 28.635 4.165 28.805 4.335 ;
        RECT 29.625 4.555 29.795 4.725 ;
        RECT 29.625 4.165 29.795 4.335 ;
        RECT 31.415 4.14 31.585 4.31 ;
        RECT 31.875 4.14 32.045 4.31 ;
        RECT 32.335 4.14 32.505 4.31 ;
        RECT 32.795 4.14 32.965 4.31 ;
        RECT 33.255 4.14 33.425 4.31 ;
        RECT 33.715 4.14 33.885 4.31 ;
        RECT 34.175 4.14 34.345 4.31 ;
        RECT 34.635 4.14 34.805 4.31 ;
        RECT 35.095 4.14 35.265 4.31 ;
        RECT 35.555 4.14 35.725 4.31 ;
        RECT 36.015 4.14 36.185 4.31 ;
        RECT 36.475 4.14 36.645 4.31 ;
        RECT 36.935 4.14 37.105 4.31 ;
        RECT 37.395 4.14 37.565 4.31 ;
        RECT 37.58 4.55 37.75 4.72 ;
        RECT 37.855 4.14 38.025 4.31 ;
        RECT 38.315 4.14 38.485 4.31 ;
        RECT 38.775 4.14 38.945 4.31 ;
        RECT 39.235 4.14 39.405 4.31 ;
        RECT 39.695 4.14 39.865 4.31 ;
        RECT 43.195 4.55 43.365 4.72 ;
        RECT 43.195 4.17 43.365 4.34 ;
        RECT 43.895 4.555 44.065 4.725 ;
        RECT 43.895 4.165 44.065 4.335 ;
        RECT 44.885 4.555 45.055 4.725 ;
        RECT 44.885 4.165 45.055 4.335 ;
        RECT 46.675 4.14 46.845 4.31 ;
        RECT 47.135 4.14 47.305 4.31 ;
        RECT 47.595 4.14 47.765 4.31 ;
        RECT 48.055 4.14 48.225 4.31 ;
        RECT 48.515 4.14 48.685 4.31 ;
        RECT 48.975 4.14 49.145 4.31 ;
        RECT 49.435 4.14 49.605 4.31 ;
        RECT 49.895 4.14 50.065 4.31 ;
        RECT 50.355 4.14 50.525 4.31 ;
        RECT 50.815 4.14 50.985 4.31 ;
        RECT 51.275 4.14 51.445 4.31 ;
        RECT 51.735 4.14 51.905 4.31 ;
        RECT 52.195 4.14 52.365 4.31 ;
        RECT 52.655 4.14 52.825 4.31 ;
        RECT 52.84 4.55 53.01 4.72 ;
        RECT 53.115 4.14 53.285 4.31 ;
        RECT 53.575 4.14 53.745 4.31 ;
        RECT 54.035 4.14 54.205 4.31 ;
        RECT 54.495 4.14 54.665 4.31 ;
        RECT 54.955 4.14 55.125 4.31 ;
        RECT 58.455 4.55 58.625 4.72 ;
        RECT 58.455 4.17 58.625 4.34 ;
        RECT 59.155 4.555 59.325 4.725 ;
        RECT 59.155 4.165 59.325 4.335 ;
        RECT 60.145 4.555 60.315 4.725 ;
        RECT 60.145 4.165 60.315 4.335 ;
        RECT 61.935 4.14 62.105 4.31 ;
        RECT 62.395 4.14 62.565 4.31 ;
        RECT 62.855 4.14 63.025 4.31 ;
        RECT 63.315 4.14 63.485 4.31 ;
        RECT 63.775 4.14 63.945 4.31 ;
        RECT 64.235 4.14 64.405 4.31 ;
        RECT 64.695 4.14 64.865 4.31 ;
        RECT 65.155 4.14 65.325 4.31 ;
        RECT 65.615 4.14 65.785 4.31 ;
        RECT 66.075 4.14 66.245 4.31 ;
        RECT 66.535 4.14 66.705 4.31 ;
        RECT 66.995 4.14 67.165 4.31 ;
        RECT 67.455 4.14 67.625 4.31 ;
        RECT 67.915 4.14 68.085 4.31 ;
        RECT 68.1 4.55 68.27 4.72 ;
        RECT 68.375 4.14 68.545 4.31 ;
        RECT 68.835 4.14 69.005 4.31 ;
        RECT 69.295 4.14 69.465 4.31 ;
        RECT 69.755 4.14 69.925 4.31 ;
        RECT 70.215 4.14 70.385 4.31 ;
        RECT 73.715 4.55 73.885 4.72 ;
        RECT 73.715 4.17 73.885 4.34 ;
        RECT 74.415 4.555 74.585 4.725 ;
        RECT 74.415 4.165 74.585 4.335 ;
        RECT 75.405 4.555 75.575 4.725 ;
        RECT 75.405 4.165 75.575 4.335 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met3 ;
        RECT 62.62 1.86 63.35 2.19 ;
        RECT 47.36 1.86 48.09 2.19 ;
        RECT 32.1 1.86 32.83 2.19 ;
        RECT 16.84 1.86 17.57 2.19 ;
        RECT 1.58 1.86 2.31 2.19 ;
      LAYER met2 ;
        RECT 62.765 1.865 63.155 2.185 ;
        RECT 62.765 1.84 63.045 2.21 ;
        RECT 47.505 1.865 47.895 2.185 ;
        RECT 47.505 1.84 47.785 2.21 ;
        RECT 32.245 1.865 32.635 2.185 ;
        RECT 32.245 1.84 32.525 2.21 ;
        RECT 16.985 1.865 17.375 2.185 ;
        RECT 16.985 1.84 17.265 2.21 ;
        RECT 1.725 1.865 2.115 2.185 ;
        RECT 1.725 1.84 2.005 2.21 ;
      LAYER li1 ;
        RECT 76.12 0.005 76.3 0.31 ;
        RECT -2.795 0.005 76.3 0.305 ;
        RECT 75.325 0.005 75.495 0.935 ;
        RECT 74.335 0.005 74.505 0.935 ;
        RECT 60.86 0.005 74.17 0.31 ;
        RECT 71.595 0.005 71.765 0.94 ;
        RECT 61.79 0.005 70.53 1.59 ;
        RECT 69.76 0.005 69.93 2.09 ;
        RECT 68.82 0.005 68.99 2.09 ;
        RECT 67.86 0.005 68.03 2.09 ;
        RECT 66.815 0.005 67.01 1.6 ;
        RECT 65.94 0.005 66.11 2.09 ;
        RECT 64.98 0.005 65.15 2.09 ;
        RECT 63.06 0.005 63.335 1.6 ;
        RECT 63.06 0.005 63.23 2.09 ;
        RECT 60.065 0.005 60.235 0.935 ;
        RECT 59.075 0.005 59.245 0.935 ;
        RECT 45.6 0.005 58.91 0.31 ;
        RECT 56.335 0.005 56.505 0.94 ;
        RECT 46.53 0.005 55.27 1.59 ;
        RECT 54.5 0.005 54.67 2.09 ;
        RECT 53.56 0.005 53.73 2.09 ;
        RECT 52.6 0.005 52.77 2.09 ;
        RECT 51.555 0.005 51.75 1.6 ;
        RECT 50.68 0.005 50.85 2.09 ;
        RECT 49.72 0.005 49.89 2.09 ;
        RECT 47.8 0.005 48.075 1.6 ;
        RECT 47.8 0.005 47.97 2.09 ;
        RECT 44.805 0.005 44.975 0.935 ;
        RECT 43.815 0.005 43.985 0.935 ;
        RECT 30.34 0.005 43.65 0.31 ;
        RECT 41.075 0.005 41.245 0.94 ;
        RECT 31.27 0.005 40.01 1.59 ;
        RECT 39.24 0.005 39.41 2.09 ;
        RECT 38.3 0.005 38.47 2.09 ;
        RECT 37.34 0.005 37.51 2.09 ;
        RECT 36.295 0.005 36.49 1.6 ;
        RECT 35.42 0.005 35.59 2.09 ;
        RECT 34.46 0.005 34.63 2.09 ;
        RECT 32.54 0.005 32.815 1.6 ;
        RECT 32.54 0.005 32.71 2.09 ;
        RECT 29.545 0.005 29.715 0.935 ;
        RECT 28.555 0.005 28.725 0.935 ;
        RECT 15.08 0.005 28.39 0.31 ;
        RECT 25.815 0.005 25.985 0.94 ;
        RECT 16.01 0.005 24.75 1.59 ;
        RECT 23.98 0.005 24.15 2.09 ;
        RECT 23.04 0.005 23.21 2.09 ;
        RECT 22.08 0.005 22.25 2.09 ;
        RECT 21.035 0.005 21.23 1.6 ;
        RECT 20.16 0.005 20.33 2.09 ;
        RECT 19.2 0.005 19.37 2.09 ;
        RECT 17.28 0.005 17.555 1.6 ;
        RECT 17.28 0.005 17.45 2.09 ;
        RECT 14.285 0.005 14.455 0.935 ;
        RECT 13.295 0.005 13.465 0.935 ;
        RECT -2.795 0.005 13.13 0.31 ;
        RECT 10.555 0.005 10.725 0.94 ;
        RECT 0.75 0.005 9.49 1.59 ;
        RECT 8.72 0.005 8.89 2.09 ;
        RECT 7.78 0.005 7.95 2.09 ;
        RECT 6.82 0.005 6.99 2.09 ;
        RECT 5.775 0.005 5.97 1.6 ;
        RECT 4.9 0.005 5.07 2.09 ;
        RECT 3.94 0.005 4.11 2.09 ;
        RECT 2.02 0.005 2.295 1.6 ;
        RECT 2.02 0.005 2.19 2.09 ;
        RECT -2.795 8.585 76.3 8.885 ;
        RECT 76.12 8.58 76.3 8.885 ;
        RECT 75.325 7.955 75.495 8.885 ;
        RECT 74.335 7.955 74.505 8.885 ;
        RECT 60.86 8.58 74.17 8.885 ;
        RECT 71.595 7.95 71.765 8.885 ;
        RECT 65.98 7.95 66.15 8.885 ;
        RECT 60.065 7.955 60.235 8.885 ;
        RECT 59.075 7.955 59.245 8.885 ;
        RECT 45.6 8.58 58.91 8.885 ;
        RECT 56.335 7.95 56.505 8.885 ;
        RECT 50.72 7.95 50.89 8.885 ;
        RECT 44.805 7.955 44.975 8.885 ;
        RECT 43.815 7.955 43.985 8.885 ;
        RECT 30.34 8.58 43.65 8.885 ;
        RECT 41.075 7.95 41.245 8.885 ;
        RECT 35.46 7.95 35.63 8.885 ;
        RECT 29.545 7.955 29.715 8.885 ;
        RECT 28.555 7.955 28.725 8.885 ;
        RECT 15.08 8.58 28.39 8.885 ;
        RECT 25.815 7.95 25.985 8.885 ;
        RECT 20.2 7.95 20.37 8.885 ;
        RECT 14.285 7.955 14.455 8.885 ;
        RECT 13.295 7.955 13.465 8.885 ;
        RECT -2.795 8.58 13.13 8.885 ;
        RECT 10.555 7.95 10.725 8.885 ;
        RECT 4.94 7.95 5.11 8.885 ;
        RECT -2.575 7.95 -2.405 8.885 ;
        RECT 66.985 6.08 67.155 8.03 ;
        RECT 66.93 7.86 67.1 8.31 ;
        RECT 66.93 5.02 67.1 6.25 ;
        RECT 63.66 2.58 64.03 2.75 ;
        RECT 63.66 1.94 63.83 2.75 ;
        RECT 63.54 1.94 63.83 2.11 ;
        RECT 62.34 2.5 62.51 2.95 ;
        RECT 51.725 6.08 51.895 8.03 ;
        RECT 51.67 7.86 51.84 8.31 ;
        RECT 51.67 5.02 51.84 6.25 ;
        RECT 48.4 2.58 48.77 2.75 ;
        RECT 48.4 1.94 48.57 2.75 ;
        RECT 48.28 1.94 48.57 2.11 ;
        RECT 47.08 2.5 47.25 2.95 ;
        RECT 36.465 6.08 36.635 8.03 ;
        RECT 36.41 7.86 36.58 8.31 ;
        RECT 36.41 5.02 36.58 6.25 ;
        RECT 33.14 2.58 33.51 2.75 ;
        RECT 33.14 1.94 33.31 2.75 ;
        RECT 33.02 1.94 33.31 2.11 ;
        RECT 31.82 2.5 31.99 2.95 ;
        RECT 21.205 6.08 21.375 8.03 ;
        RECT 21.15 7.86 21.32 8.31 ;
        RECT 21.15 5.02 21.32 6.25 ;
        RECT 17.88 2.58 18.25 2.75 ;
        RECT 17.88 1.94 18.05 2.75 ;
        RECT 17.76 1.94 18.05 2.11 ;
        RECT 16.56 2.5 16.73 2.95 ;
        RECT 5.945 6.08 6.115 8.03 ;
        RECT 5.89 7.86 6.06 8.31 ;
        RECT 5.89 5.02 6.06 6.25 ;
        RECT 2.62 2.58 2.99 2.75 ;
        RECT 2.62 1.94 2.79 2.75 ;
        RECT 2.5 1.94 2.79 2.11 ;
        RECT 1.3 2.5 1.47 2.95 ;
      LAYER met1 ;
        RECT 76.12 0.005 76.3 0.31 ;
        RECT -2.795 0.005 76.3 0.305 ;
        RECT 60.86 0.005 74.17 0.31 ;
        RECT 61.79 0.005 70.53 1.745 ;
        RECT 63.48 1.91 63.77 2.14 ;
        RECT 62.595 1.955 63.77 2.095 ;
        RECT 62.775 1.895 63.185 2.155 ;
        RECT 62.775 0.005 63.065 2.155 ;
        RECT 62.355 2.375 62.975 2.515 ;
        RECT 62.835 0.005 62.975 2.515 ;
        RECT 62.595 1.955 62.975 2.215 ;
        RECT 62.28 2.75 62.57 2.98 ;
        RECT 62.355 2.375 62.495 2.98 ;
        RECT 45.6 0.005 58.91 0.31 ;
        RECT 46.53 0.005 55.27 1.745 ;
        RECT 48.22 1.91 48.51 2.14 ;
        RECT 47.335 1.955 48.51 2.095 ;
        RECT 47.515 1.895 47.925 2.155 ;
        RECT 47.515 0.005 47.805 2.155 ;
        RECT 47.095 2.375 47.715 2.515 ;
        RECT 47.575 0.005 47.715 2.515 ;
        RECT 47.335 1.955 47.715 2.215 ;
        RECT 47.02 2.75 47.31 2.98 ;
        RECT 47.095 2.375 47.235 2.98 ;
        RECT 30.34 0.005 43.65 0.31 ;
        RECT 31.27 0.005 40.01 1.745 ;
        RECT 32.96 1.91 33.25 2.14 ;
        RECT 32.075 1.955 33.25 2.095 ;
        RECT 32.255 1.895 32.665 2.155 ;
        RECT 32.255 0.005 32.545 2.155 ;
        RECT 31.835 2.375 32.455 2.515 ;
        RECT 32.315 0.005 32.455 2.515 ;
        RECT 32.075 1.955 32.455 2.215 ;
        RECT 31.76 2.75 32.05 2.98 ;
        RECT 31.835 2.375 31.975 2.98 ;
        RECT 15.08 0.005 28.39 0.31 ;
        RECT 16.01 0.005 24.75 1.745 ;
        RECT 17.7 1.91 17.99 2.14 ;
        RECT 16.815 1.955 17.99 2.095 ;
        RECT 16.995 1.895 17.405 2.155 ;
        RECT 16.995 0.005 17.285 2.155 ;
        RECT 16.575 2.375 17.195 2.515 ;
        RECT 17.055 0.005 17.195 2.515 ;
        RECT 16.815 1.955 17.195 2.215 ;
        RECT 16.5 2.75 16.79 2.98 ;
        RECT 16.575 2.375 16.715 2.98 ;
        RECT -2.795 0.005 13.13 0.31 ;
        RECT 0.75 0.005 9.49 1.745 ;
        RECT 2.44 1.91 2.73 2.14 ;
        RECT 1.555 1.955 2.73 2.095 ;
        RECT 1.735 1.895 2.145 2.155 ;
        RECT 1.735 0.005 2.025 2.155 ;
        RECT 1.315 2.375 1.935 2.515 ;
        RECT 1.795 0.005 1.935 2.515 ;
        RECT 1.555 1.955 1.935 2.215 ;
        RECT 1.24 2.75 1.53 2.98 ;
        RECT 1.315 2.375 1.455 2.98 ;
        RECT -2.795 8.585 76.3 8.885 ;
        RECT 76.12 8.58 76.3 8.885 ;
        RECT 60.86 8.58 74.17 8.885 ;
        RECT 66.925 6.29 67.215 6.52 ;
        RECT 66.76 6.32 66.93 8.885 ;
        RECT 66.755 6.32 67.215 6.49 ;
        RECT 45.6 8.58 58.91 8.885 ;
        RECT 51.665 6.29 51.955 6.52 ;
        RECT 51.5 6.32 51.67 8.885 ;
        RECT 51.495 6.32 51.955 6.49 ;
        RECT 30.34 8.58 43.65 8.885 ;
        RECT 36.405 6.29 36.695 6.52 ;
        RECT 36.24 6.32 36.41 8.885 ;
        RECT 36.235 6.32 36.695 6.49 ;
        RECT 15.08 8.58 28.39 8.885 ;
        RECT 21.145 6.29 21.435 6.52 ;
        RECT 20.98 6.32 21.15 8.885 ;
        RECT 20.975 6.32 21.435 6.49 ;
        RECT -2.795 8.58 13.13 8.885 ;
        RECT 5.885 6.29 6.175 6.52 ;
        RECT 5.72 6.32 5.89 8.885 ;
        RECT 5.715 6.32 6.175 6.49 ;
      LAYER via2 ;
        RECT 1.765 1.925 1.965 2.125 ;
        RECT 17.025 1.925 17.225 2.125 ;
        RECT 32.285 1.925 32.485 2.125 ;
        RECT 47.545 1.925 47.745 2.125 ;
        RECT 62.805 1.925 63.005 2.125 ;
      LAYER via1 ;
        RECT 1.91 1.95 2.06 2.1 ;
        RECT 17.17 1.95 17.32 2.1 ;
        RECT 32.43 1.95 32.58 2.1 ;
        RECT 47.69 1.95 47.84 2.1 ;
        RECT 62.95 1.95 63.1 2.1 ;
      LAYER mcon ;
        RECT -2.495 8.61 -2.325 8.78 ;
        RECT -1.815 8.61 -1.645 8.78 ;
        RECT -1.135 8.61 -0.965 8.78 ;
        RECT -0.455 8.61 -0.285 8.78 ;
        RECT 0.895 1.42 1.065 1.59 ;
        RECT 1.3 2.78 1.47 2.95 ;
        RECT 1.355 1.42 1.525 1.59 ;
        RECT 1.815 1.42 1.985 1.59 ;
        RECT 2.275 1.42 2.445 1.59 ;
        RECT 2.5 1.94 2.67 2.11 ;
        RECT 2.735 1.42 2.905 1.59 ;
        RECT 3.195 1.42 3.365 1.59 ;
        RECT 3.655 1.42 3.825 1.59 ;
        RECT 4.115 1.42 4.285 1.59 ;
        RECT 4.575 1.42 4.745 1.59 ;
        RECT 5.02 8.61 5.19 8.78 ;
        RECT 5.035 1.42 5.205 1.59 ;
        RECT 5.495 1.42 5.665 1.59 ;
        RECT 5.7 8.61 5.87 8.78 ;
        RECT 5.945 6.32 6.115 6.49 ;
        RECT 5.955 1.42 6.125 1.59 ;
        RECT 6.38 8.61 6.55 8.78 ;
        RECT 6.415 1.42 6.585 1.59 ;
        RECT 6.875 1.42 7.045 1.59 ;
        RECT 7.06 8.61 7.23 8.78 ;
        RECT 7.335 1.42 7.505 1.59 ;
        RECT 7.795 1.42 7.965 1.59 ;
        RECT 8.255 1.42 8.425 1.59 ;
        RECT 8.715 1.42 8.885 1.59 ;
        RECT 9.175 1.42 9.345 1.59 ;
        RECT 10.635 8.61 10.805 8.78 ;
        RECT 10.635 0.11 10.805 0.28 ;
        RECT 11.315 8.61 11.485 8.78 ;
        RECT 11.315 0.11 11.485 0.28 ;
        RECT 11.995 8.61 12.165 8.78 ;
        RECT 11.995 0.11 12.165 0.28 ;
        RECT 12.675 8.61 12.845 8.78 ;
        RECT 12.675 0.11 12.845 0.28 ;
        RECT 13.375 8.615 13.545 8.785 ;
        RECT 13.375 0.105 13.545 0.275 ;
        RECT 14.365 8.615 14.535 8.785 ;
        RECT 14.365 0.105 14.535 0.275 ;
        RECT 16.155 1.42 16.325 1.59 ;
        RECT 16.56 2.78 16.73 2.95 ;
        RECT 16.615 1.42 16.785 1.59 ;
        RECT 17.075 1.42 17.245 1.59 ;
        RECT 17.535 1.42 17.705 1.59 ;
        RECT 17.76 1.94 17.93 2.11 ;
        RECT 17.995 1.42 18.165 1.59 ;
        RECT 18.455 1.42 18.625 1.59 ;
        RECT 18.915 1.42 19.085 1.59 ;
        RECT 19.375 1.42 19.545 1.59 ;
        RECT 19.835 1.42 20.005 1.59 ;
        RECT 20.28 8.61 20.45 8.78 ;
        RECT 20.295 1.42 20.465 1.59 ;
        RECT 20.755 1.42 20.925 1.59 ;
        RECT 20.96 8.61 21.13 8.78 ;
        RECT 21.205 6.32 21.375 6.49 ;
        RECT 21.215 1.42 21.385 1.59 ;
        RECT 21.64 8.61 21.81 8.78 ;
        RECT 21.675 1.42 21.845 1.59 ;
        RECT 22.135 1.42 22.305 1.59 ;
        RECT 22.32 8.61 22.49 8.78 ;
        RECT 22.595 1.42 22.765 1.59 ;
        RECT 23.055 1.42 23.225 1.59 ;
        RECT 23.515 1.42 23.685 1.59 ;
        RECT 23.975 1.42 24.145 1.59 ;
        RECT 24.435 1.42 24.605 1.59 ;
        RECT 25.895 8.61 26.065 8.78 ;
        RECT 25.895 0.11 26.065 0.28 ;
        RECT 26.575 8.61 26.745 8.78 ;
        RECT 26.575 0.11 26.745 0.28 ;
        RECT 27.255 8.61 27.425 8.78 ;
        RECT 27.255 0.11 27.425 0.28 ;
        RECT 27.935 8.61 28.105 8.78 ;
        RECT 27.935 0.11 28.105 0.28 ;
        RECT 28.635 8.615 28.805 8.785 ;
        RECT 28.635 0.105 28.805 0.275 ;
        RECT 29.625 8.615 29.795 8.785 ;
        RECT 29.625 0.105 29.795 0.275 ;
        RECT 31.415 1.42 31.585 1.59 ;
        RECT 31.82 2.78 31.99 2.95 ;
        RECT 31.875 1.42 32.045 1.59 ;
        RECT 32.335 1.42 32.505 1.59 ;
        RECT 32.795 1.42 32.965 1.59 ;
        RECT 33.02 1.94 33.19 2.11 ;
        RECT 33.255 1.42 33.425 1.59 ;
        RECT 33.715 1.42 33.885 1.59 ;
        RECT 34.175 1.42 34.345 1.59 ;
        RECT 34.635 1.42 34.805 1.59 ;
        RECT 35.095 1.42 35.265 1.59 ;
        RECT 35.54 8.61 35.71 8.78 ;
        RECT 35.555 1.42 35.725 1.59 ;
        RECT 36.015 1.42 36.185 1.59 ;
        RECT 36.22 8.61 36.39 8.78 ;
        RECT 36.465 6.32 36.635 6.49 ;
        RECT 36.475 1.42 36.645 1.59 ;
        RECT 36.9 8.61 37.07 8.78 ;
        RECT 36.935 1.42 37.105 1.59 ;
        RECT 37.395 1.42 37.565 1.59 ;
        RECT 37.58 8.61 37.75 8.78 ;
        RECT 37.855 1.42 38.025 1.59 ;
        RECT 38.315 1.42 38.485 1.59 ;
        RECT 38.775 1.42 38.945 1.59 ;
        RECT 39.235 1.42 39.405 1.59 ;
        RECT 39.695 1.42 39.865 1.59 ;
        RECT 41.155 8.61 41.325 8.78 ;
        RECT 41.155 0.11 41.325 0.28 ;
        RECT 41.835 8.61 42.005 8.78 ;
        RECT 41.835 0.11 42.005 0.28 ;
        RECT 42.515 8.61 42.685 8.78 ;
        RECT 42.515 0.11 42.685 0.28 ;
        RECT 43.195 8.61 43.365 8.78 ;
        RECT 43.195 0.11 43.365 0.28 ;
        RECT 43.895 8.615 44.065 8.785 ;
        RECT 43.895 0.105 44.065 0.275 ;
        RECT 44.885 8.615 45.055 8.785 ;
        RECT 44.885 0.105 45.055 0.275 ;
        RECT 46.675 1.42 46.845 1.59 ;
        RECT 47.08 2.78 47.25 2.95 ;
        RECT 47.135 1.42 47.305 1.59 ;
        RECT 47.595 1.42 47.765 1.59 ;
        RECT 48.055 1.42 48.225 1.59 ;
        RECT 48.28 1.94 48.45 2.11 ;
        RECT 48.515 1.42 48.685 1.59 ;
        RECT 48.975 1.42 49.145 1.59 ;
        RECT 49.435 1.42 49.605 1.59 ;
        RECT 49.895 1.42 50.065 1.59 ;
        RECT 50.355 1.42 50.525 1.59 ;
        RECT 50.8 8.61 50.97 8.78 ;
        RECT 50.815 1.42 50.985 1.59 ;
        RECT 51.275 1.42 51.445 1.59 ;
        RECT 51.48 8.61 51.65 8.78 ;
        RECT 51.725 6.32 51.895 6.49 ;
        RECT 51.735 1.42 51.905 1.59 ;
        RECT 52.16 8.61 52.33 8.78 ;
        RECT 52.195 1.42 52.365 1.59 ;
        RECT 52.655 1.42 52.825 1.59 ;
        RECT 52.84 8.61 53.01 8.78 ;
        RECT 53.115 1.42 53.285 1.59 ;
        RECT 53.575 1.42 53.745 1.59 ;
        RECT 54.035 1.42 54.205 1.59 ;
        RECT 54.495 1.42 54.665 1.59 ;
        RECT 54.955 1.42 55.125 1.59 ;
        RECT 56.415 8.61 56.585 8.78 ;
        RECT 56.415 0.11 56.585 0.28 ;
        RECT 57.095 8.61 57.265 8.78 ;
        RECT 57.095 0.11 57.265 0.28 ;
        RECT 57.775 8.61 57.945 8.78 ;
        RECT 57.775 0.11 57.945 0.28 ;
        RECT 58.455 8.61 58.625 8.78 ;
        RECT 58.455 0.11 58.625 0.28 ;
        RECT 59.155 8.615 59.325 8.785 ;
        RECT 59.155 0.105 59.325 0.275 ;
        RECT 60.145 8.615 60.315 8.785 ;
        RECT 60.145 0.105 60.315 0.275 ;
        RECT 61.935 1.42 62.105 1.59 ;
        RECT 62.34 2.78 62.51 2.95 ;
        RECT 62.395 1.42 62.565 1.59 ;
        RECT 62.855 1.42 63.025 1.59 ;
        RECT 63.315 1.42 63.485 1.59 ;
        RECT 63.54 1.94 63.71 2.11 ;
        RECT 63.775 1.42 63.945 1.59 ;
        RECT 64.235 1.42 64.405 1.59 ;
        RECT 64.695 1.42 64.865 1.59 ;
        RECT 65.155 1.42 65.325 1.59 ;
        RECT 65.615 1.42 65.785 1.59 ;
        RECT 66.06 8.61 66.23 8.78 ;
        RECT 66.075 1.42 66.245 1.59 ;
        RECT 66.535 1.42 66.705 1.59 ;
        RECT 66.74 8.61 66.91 8.78 ;
        RECT 66.985 6.32 67.155 6.49 ;
        RECT 66.995 1.42 67.165 1.59 ;
        RECT 67.42 8.61 67.59 8.78 ;
        RECT 67.455 1.42 67.625 1.59 ;
        RECT 67.915 1.42 68.085 1.59 ;
        RECT 68.1 8.61 68.27 8.78 ;
        RECT 68.375 1.42 68.545 1.59 ;
        RECT 68.835 1.42 69.005 1.59 ;
        RECT 69.295 1.42 69.465 1.59 ;
        RECT 69.755 1.42 69.925 1.59 ;
        RECT 70.215 1.42 70.385 1.59 ;
        RECT 71.675 8.61 71.845 8.78 ;
        RECT 71.675 0.11 71.845 0.28 ;
        RECT 72.355 8.61 72.525 8.78 ;
        RECT 72.355 0.11 72.525 0.28 ;
        RECT 73.035 8.61 73.205 8.78 ;
        RECT 73.035 0.11 73.205 0.28 ;
        RECT 73.715 8.61 73.885 8.78 ;
        RECT 73.715 0.11 73.885 0.28 ;
        RECT 74.415 8.615 74.585 8.785 ;
        RECT 74.415 0.105 74.585 0.275 ;
        RECT 75.405 8.615 75.575 8.785 ;
        RECT 75.405 0.105 75.575 0.275 ;
    END
  END vssd1
  OBS
    LAYER met4 ;
      RECT 63.94 2.98 64.27 3.31 ;
      RECT 63.955 2.505 64.27 3.31 ;
      RECT 66.1 2.49 66.43 2.845 ;
      RECT 63.955 2.505 66.43 2.805 ;
      RECT 48.68 2.98 49.01 3.31 ;
      RECT 48.695 2.505 49.01 3.31 ;
      RECT 50.84 2.49 51.17 2.845 ;
      RECT 48.695 2.505 51.17 2.805 ;
      RECT 33.42 2.98 33.75 3.31 ;
      RECT 33.435 2.505 33.75 3.31 ;
      RECT 35.58 2.49 35.91 2.845 ;
      RECT 33.435 2.505 35.91 2.805 ;
      RECT 18.16 2.98 18.49 3.31 ;
      RECT 18.175 2.505 18.49 3.31 ;
      RECT 20.32 2.49 20.65 2.845 ;
      RECT 18.175 2.505 20.65 2.805 ;
      RECT 2.9 2.98 3.23 3.31 ;
      RECT 2.915 2.505 3.23 3.31 ;
      RECT 5.06 2.49 5.39 2.845 ;
      RECT 2.915 2.505 5.39 2.805 ;
    LAYER via3 ;
      RECT 66.165 2.58 66.365 2.78 ;
      RECT 64.005 3.045 64.205 3.245 ;
      RECT 50.905 2.58 51.105 2.78 ;
      RECT 48.745 3.045 48.945 3.245 ;
      RECT 35.645 2.58 35.845 2.78 ;
      RECT 33.485 3.045 33.685 3.245 ;
      RECT 20.385 2.58 20.585 2.78 ;
      RECT 18.225 3.045 18.425 3.245 ;
      RECT 5.125 2.58 5.325 2.78 ;
      RECT 2.965 3.045 3.165 3.245 ;
    LAYER met3 ;
      RECT 70.965 1.11 71.305 3.07 ;
      RECT 65.225 1.885 65.955 2.215 ;
      RECT 65.375 1.11 65.675 2.215 ;
      RECT 65.375 1.11 71.305 1.41 ;
      RECT 67.26 7.06 67.63 7.43 ;
      RECT 67.295 4.48 67.595 7.43 ;
      RECT 65.855 4.48 67.595 4.78 ;
      RECT 63.06 4.26 66.155 4.56 ;
      RECT 65.855 2.52 66.155 4.78 ;
      RECT 63.06 2.98 63.36 4.56 ;
      RECT 66.58 3.515 66.91 3.87 ;
      RECT 64.675 3.555 66.91 3.855 ;
      RECT 64.675 2.42 64.975 3.855 ;
      RECT 62.755 2.98 63.485 3.31 ;
      RECT 65.65 2.525 66.43 2.87 ;
      RECT 66.125 2.49 66.43 2.87 ;
      RECT 64.66 2.42 64.99 2.75 ;
      RECT 63.945 2.42 64.265 3.335 ;
      RECT 63.945 2.42 64.275 2.955 ;
      RECT 55.705 1.11 56.045 3.07 ;
      RECT 49.965 1.885 50.695 2.215 ;
      RECT 50.115 1.11 50.415 2.215 ;
      RECT 50.115 1.11 56.045 1.41 ;
      RECT 52 7.06 52.37 7.43 ;
      RECT 52.035 4.48 52.335 7.43 ;
      RECT 50.595 4.48 52.335 4.78 ;
      RECT 47.8 4.26 50.895 4.56 ;
      RECT 50.595 2.52 50.895 4.78 ;
      RECT 47.8 2.98 48.1 4.56 ;
      RECT 51.32 3.515 51.65 3.87 ;
      RECT 49.415 3.555 51.65 3.855 ;
      RECT 49.415 2.42 49.715 3.855 ;
      RECT 47.495 2.98 48.225 3.31 ;
      RECT 50.39 2.525 51.17 2.87 ;
      RECT 50.865 2.49 51.17 2.87 ;
      RECT 49.4 2.42 49.73 2.75 ;
      RECT 48.685 2.42 49.005 3.335 ;
      RECT 48.685 2.42 49.015 2.955 ;
      RECT 40.445 1.11 40.785 3.07 ;
      RECT 34.705 1.885 35.435 2.215 ;
      RECT 34.855 1.11 35.155 2.215 ;
      RECT 34.855 1.11 40.785 1.41 ;
      RECT 36.74 7.06 37.11 7.43 ;
      RECT 36.775 4.48 37.075 7.43 ;
      RECT 35.335 4.48 37.075 4.78 ;
      RECT 32.54 4.26 35.635 4.56 ;
      RECT 35.335 2.52 35.635 4.78 ;
      RECT 32.54 2.98 32.84 4.56 ;
      RECT 36.06 3.515 36.39 3.87 ;
      RECT 34.155 3.555 36.39 3.855 ;
      RECT 34.155 2.42 34.455 3.855 ;
      RECT 32.235 2.98 32.965 3.31 ;
      RECT 35.13 2.525 35.91 2.87 ;
      RECT 35.605 2.49 35.91 2.87 ;
      RECT 34.14 2.42 34.47 2.75 ;
      RECT 33.425 2.42 33.745 3.335 ;
      RECT 33.425 2.42 33.755 2.955 ;
      RECT 25.185 1.11 25.525 3.07 ;
      RECT 19.445 1.885 20.175 2.215 ;
      RECT 19.595 1.11 19.895 2.215 ;
      RECT 19.595 1.11 25.525 1.41 ;
      RECT 21.48 7.06 21.85 7.43 ;
      RECT 21.515 4.48 21.815 7.43 ;
      RECT 20.075 4.48 21.815 4.78 ;
      RECT 17.28 4.26 20.375 4.56 ;
      RECT 20.075 2.52 20.375 4.78 ;
      RECT 17.28 2.98 17.58 4.56 ;
      RECT 20.8 3.515 21.13 3.87 ;
      RECT 18.895 3.555 21.13 3.855 ;
      RECT 18.895 2.42 19.195 3.855 ;
      RECT 16.975 2.98 17.705 3.31 ;
      RECT 19.87 2.525 20.65 2.87 ;
      RECT 20.345 2.49 20.65 2.87 ;
      RECT 18.88 2.42 19.21 2.75 ;
      RECT 18.165 2.42 18.485 3.335 ;
      RECT 18.165 2.42 18.495 2.955 ;
      RECT 9.925 1.11 10.265 3.07 ;
      RECT 4.185 1.885 4.915 2.215 ;
      RECT 4.335 1.11 4.635 2.215 ;
      RECT 4.335 1.11 10.265 1.41 ;
      RECT 6.22 7.06 6.59 7.43 ;
      RECT 6.255 4.48 6.555 7.43 ;
      RECT 4.815 4.48 6.555 4.78 ;
      RECT 2.02 4.26 5.115 4.56 ;
      RECT 4.815 2.52 5.115 4.78 ;
      RECT 2.02 2.98 2.32 4.56 ;
      RECT 5.54 3.515 5.87 3.87 ;
      RECT 3.635 3.555 5.87 3.855 ;
      RECT 3.635 2.42 3.935 3.855 ;
      RECT 1.715 2.98 2.445 3.31 ;
      RECT 4.61 2.525 5.39 2.87 ;
      RECT 5.085 2.49 5.39 2.87 ;
      RECT 3.62 2.42 3.95 2.75 ;
      RECT 2.905 2.42 3.225 3.335 ;
      RECT 2.905 2.42 3.235 2.955 ;
      RECT 69.5 1.86 70.23 2.19 ;
      RECT 67.81 1.875 68.54 2.205 ;
      RECT 66.775 1.86 67.505 2.21 ;
      RECT 54.24 1.86 54.97 2.19 ;
      RECT 52.55 1.875 53.28 2.205 ;
      RECT 51.515 1.86 52.245 2.21 ;
      RECT 38.98 1.86 39.71 2.19 ;
      RECT 37.29 1.875 38.02 2.205 ;
      RECT 36.255 1.86 36.985 2.21 ;
      RECT 23.72 1.86 24.45 2.19 ;
      RECT 22.03 1.875 22.76 2.205 ;
      RECT 20.995 1.86 21.725 2.21 ;
      RECT 8.46 1.86 9.19 2.19 ;
      RECT 6.77 1.875 7.5 2.205 ;
      RECT 5.735 1.86 6.465 2.21 ;
    LAYER via2 ;
      RECT 71.04 2.78 71.24 2.98 ;
      RECT 69.735 1.925 69.935 2.125 ;
      RECT 67.875 1.94 68.075 2.14 ;
      RECT 67.345 7.145 67.545 7.345 ;
      RECT 66.855 1.945 67.055 2.145 ;
      RECT 66.645 3.58 66.845 3.78 ;
      RECT 66.165 2.58 66.365 2.78 ;
      RECT 65.415 1.95 65.615 2.15 ;
      RECT 64.725 2.485 64.925 2.685 ;
      RECT 64.01 2.485 64.21 2.685 ;
      RECT 63.045 3.045 63.245 3.245 ;
      RECT 55.78 2.78 55.98 2.98 ;
      RECT 54.475 1.925 54.675 2.125 ;
      RECT 52.615 1.94 52.815 2.14 ;
      RECT 52.085 7.145 52.285 7.345 ;
      RECT 51.595 1.945 51.795 2.145 ;
      RECT 51.385 3.58 51.585 3.78 ;
      RECT 50.905 2.58 51.105 2.78 ;
      RECT 50.155 1.95 50.355 2.15 ;
      RECT 49.465 2.485 49.665 2.685 ;
      RECT 48.75 2.485 48.95 2.685 ;
      RECT 47.785 3.045 47.985 3.245 ;
      RECT 40.52 2.78 40.72 2.98 ;
      RECT 39.215 1.925 39.415 2.125 ;
      RECT 37.355 1.94 37.555 2.14 ;
      RECT 36.825 7.145 37.025 7.345 ;
      RECT 36.335 1.945 36.535 2.145 ;
      RECT 36.125 3.58 36.325 3.78 ;
      RECT 35.645 2.58 35.845 2.78 ;
      RECT 34.895 1.95 35.095 2.15 ;
      RECT 34.205 2.485 34.405 2.685 ;
      RECT 33.49 2.485 33.69 2.685 ;
      RECT 32.525 3.045 32.725 3.245 ;
      RECT 25.26 2.78 25.46 2.98 ;
      RECT 23.955 1.925 24.155 2.125 ;
      RECT 22.095 1.94 22.295 2.14 ;
      RECT 21.565 7.145 21.765 7.345 ;
      RECT 21.075 1.945 21.275 2.145 ;
      RECT 20.865 3.58 21.065 3.78 ;
      RECT 20.385 2.58 20.585 2.78 ;
      RECT 19.635 1.95 19.835 2.15 ;
      RECT 18.945 2.485 19.145 2.685 ;
      RECT 18.23 2.485 18.43 2.685 ;
      RECT 17.265 3.045 17.465 3.245 ;
      RECT 10 2.78 10.2 2.98 ;
      RECT 8.695 1.925 8.895 2.125 ;
      RECT 6.835 1.94 7.035 2.14 ;
      RECT 6.305 7.145 6.505 7.345 ;
      RECT 5.815 1.945 6.015 2.145 ;
      RECT 5.605 3.58 5.805 3.78 ;
      RECT 5.125 2.58 5.325 2.78 ;
      RECT 4.375 1.95 4.575 2.15 ;
      RECT 3.685 2.485 3.885 2.685 ;
      RECT 2.97 2.485 3.17 2.685 ;
      RECT 2.005 3.045 2.205 3.245 ;
    LAYER met2 ;
      RECT -1.565 8.405 75.93 8.575 ;
      RECT 75.76 7.28 75.93 8.575 ;
      RECT -1.565 6.26 -1.395 8.575 ;
      RECT 75.73 7.28 76.08 7.63 ;
      RECT -1.63 6.26 -1.34 6.61 ;
      RECT 72.57 6.225 72.89 6.55 ;
      RECT 72.6 5.7 72.77 6.55 ;
      RECT 72.6 5.7 72.775 6.05 ;
      RECT 72.6 5.7 73.575 5.875 ;
      RECT 73.4 1.97 73.575 5.875 ;
      RECT 73.345 1.97 73.695 2.32 ;
      RECT 73.37 6.66 73.695 6.985 ;
      RECT 72.255 6.75 73.695 6.92 ;
      RECT 72.255 2.4 72.415 6.92 ;
      RECT 72.57 2.37 72.89 2.69 ;
      RECT 72.255 2.4 72.89 2.57 ;
      RECT 70.995 2.69 71.285 3.07 ;
      RECT 70.965 2.705 71.305 3.055 ;
      RECT 69.705 3.545 69.965 3.865 ;
      RECT 69.765 1.84 69.905 3.865 ;
      RECT 69.59 2.4 69.905 2.77 ;
      RECT 69.66 1.955 69.905 2.77 ;
      RECT 69.695 1.84 69.975 2.21 ;
      RECT 69.015 2.425 69.275 2.745 ;
      RECT 68.355 2.515 69.275 2.655 ;
      RECT 68.355 1.575 68.495 2.655 ;
      RECT 64.815 1.865 65.075 2.185 ;
      RECT 64.995 1.575 65.135 2.095 ;
      RECT 64.995 1.575 68.495 1.715 ;
      RECT 60.445 6.66 60.795 7.01 ;
      RECT 67.93 6.615 68.28 6.965 ;
      RECT 60.445 6.69 68.28 6.89 ;
      RECT 67.845 3.265 68.105 3.585 ;
      RECT 67.905 1.855 68.045 3.585 ;
      RECT 67.835 1.855 68.115 2.225 ;
      RECT 65.235 4.015 67.67 4.155 ;
      RECT 67.53 2.705 67.67 4.155 ;
      RECT 65.235 3.635 65.375 4.155 ;
      RECT 64.935 3.635 65.375 3.865 ;
      RECT 62.595 3.635 65.375 3.775 ;
      RECT 64.935 3.545 65.195 3.865 ;
      RECT 62.595 3.355 62.735 3.775 ;
      RECT 62.085 3.265 62.345 3.585 ;
      RECT 62.085 3.355 62.735 3.495 ;
      RECT 62.145 1.865 62.285 3.585 ;
      RECT 67.47 2.705 67.73 3.025 ;
      RECT 62.085 1.865 62.345 2.185 ;
      RECT 67.095 3.545 67.355 3.865 ;
      RECT 67.155 1.955 67.295 3.865 ;
      RECT 66.815 1.955 67.295 2.23 ;
      RECT 66.615 1.86 67.095 2.205 ;
      RECT 66.605 3.495 66.885 3.865 ;
      RECT 66.675 2.4 66.815 3.865 ;
      RECT 66.615 2.4 66.875 3.025 ;
      RECT 66.605 2.4 66.885 2.77 ;
      RECT 65.535 3.545 65.795 3.865 ;
      RECT 65.535 3.355 65.735 3.865 ;
      RECT 65.34 3.355 65.735 3.495 ;
      RECT 65.34 1.865 65.48 3.495 ;
      RECT 65.34 1.865 65.655 2.235 ;
      RECT 65.28 1.865 65.655 2.185 ;
      RECT 63.005 2.96 63.285 3.33 ;
      RECT 64.455 2.985 64.715 3.305 ;
      RECT 62.835 3.075 64.715 3.215 ;
      RECT 62.835 2.96 63.285 3.215 ;
      RECT 62.775 2.4 63.035 3.025 ;
      RECT 62.765 2.4 63.045 2.77 ;
      RECT 63.845 2.4 64.255 2.77 ;
      RECT 63.255 2.425 63.515 2.745 ;
      RECT 63.255 2.515 64.255 2.655 ;
      RECT 57.31 6.225 57.63 6.55 ;
      RECT 57.34 5.7 57.51 6.55 ;
      RECT 57.34 5.7 57.515 6.05 ;
      RECT 57.34 5.7 58.315 5.875 ;
      RECT 58.14 1.97 58.315 5.875 ;
      RECT 58.085 1.97 58.435 2.32 ;
      RECT 58.11 6.66 58.435 6.985 ;
      RECT 56.995 6.75 58.435 6.92 ;
      RECT 56.995 2.4 57.155 6.92 ;
      RECT 57.31 2.37 57.63 2.69 ;
      RECT 56.995 2.4 57.63 2.57 ;
      RECT 55.735 2.69 56.025 3.07 ;
      RECT 55.705 2.705 56.045 3.055 ;
      RECT 54.445 3.545 54.705 3.865 ;
      RECT 54.505 1.84 54.645 3.865 ;
      RECT 54.33 2.4 54.645 2.77 ;
      RECT 54.4 1.955 54.645 2.77 ;
      RECT 54.435 1.84 54.715 2.21 ;
      RECT 53.755 2.425 54.015 2.745 ;
      RECT 53.095 2.515 54.015 2.655 ;
      RECT 53.095 1.575 53.235 2.655 ;
      RECT 49.555 1.865 49.815 2.185 ;
      RECT 49.735 1.575 49.875 2.095 ;
      RECT 49.735 1.575 53.235 1.715 ;
      RECT 45.185 6.66 45.535 7.01 ;
      RECT 52.675 6.615 53.025 6.965 ;
      RECT 45.185 6.69 53.025 6.89 ;
      RECT 52.585 3.265 52.845 3.585 ;
      RECT 52.645 1.855 52.785 3.585 ;
      RECT 52.575 1.855 52.855 2.225 ;
      RECT 49.975 4.015 52.41 4.155 ;
      RECT 52.27 2.705 52.41 4.155 ;
      RECT 49.975 3.635 50.115 4.155 ;
      RECT 49.675 3.635 50.115 3.865 ;
      RECT 47.335 3.635 50.115 3.775 ;
      RECT 49.675 3.545 49.935 3.865 ;
      RECT 47.335 3.355 47.475 3.775 ;
      RECT 46.825 3.265 47.085 3.585 ;
      RECT 46.825 3.355 47.475 3.495 ;
      RECT 46.885 1.865 47.025 3.585 ;
      RECT 52.21 2.705 52.47 3.025 ;
      RECT 46.825 1.865 47.085 2.185 ;
      RECT 51.835 3.545 52.095 3.865 ;
      RECT 51.895 1.955 52.035 3.865 ;
      RECT 51.555 1.955 52.035 2.23 ;
      RECT 51.355 1.86 51.835 2.205 ;
      RECT 51.345 3.495 51.625 3.865 ;
      RECT 51.415 2.4 51.555 3.865 ;
      RECT 51.355 2.4 51.615 3.025 ;
      RECT 51.345 2.4 51.625 2.77 ;
      RECT 50.275 3.545 50.535 3.865 ;
      RECT 50.275 3.355 50.475 3.865 ;
      RECT 50.08 3.355 50.475 3.495 ;
      RECT 50.08 1.865 50.22 3.495 ;
      RECT 50.08 1.865 50.395 2.235 ;
      RECT 50.02 1.865 50.395 2.185 ;
      RECT 47.745 2.96 48.025 3.33 ;
      RECT 49.195 2.985 49.455 3.305 ;
      RECT 47.575 3.075 49.455 3.215 ;
      RECT 47.575 2.96 48.025 3.215 ;
      RECT 47.515 2.4 47.775 3.025 ;
      RECT 47.505 2.4 47.785 2.77 ;
      RECT 48.585 2.4 48.995 2.77 ;
      RECT 47.995 2.425 48.255 2.745 ;
      RECT 47.995 2.515 48.995 2.655 ;
      RECT 42.05 6.225 42.37 6.55 ;
      RECT 42.08 5.7 42.25 6.55 ;
      RECT 42.08 5.7 42.255 6.05 ;
      RECT 42.08 5.7 43.055 5.875 ;
      RECT 42.88 1.97 43.055 5.875 ;
      RECT 42.825 1.97 43.175 2.32 ;
      RECT 42.85 6.66 43.175 6.985 ;
      RECT 41.735 6.75 43.175 6.92 ;
      RECT 41.735 2.4 41.895 6.92 ;
      RECT 42.05 2.37 42.37 2.69 ;
      RECT 41.735 2.4 42.37 2.57 ;
      RECT 40.475 2.69 40.765 3.07 ;
      RECT 40.445 2.705 40.785 3.055 ;
      RECT 39.185 3.545 39.445 3.865 ;
      RECT 39.245 1.84 39.385 3.865 ;
      RECT 39.07 2.4 39.385 2.77 ;
      RECT 39.14 1.955 39.385 2.77 ;
      RECT 39.175 1.84 39.455 2.21 ;
      RECT 38.495 2.425 38.755 2.745 ;
      RECT 37.835 2.515 38.755 2.655 ;
      RECT 37.835 1.575 37.975 2.655 ;
      RECT 34.295 1.865 34.555 2.185 ;
      RECT 34.475 1.575 34.615 2.095 ;
      RECT 34.475 1.575 37.975 1.715 ;
      RECT 29.97 6.665 30.32 7.015 ;
      RECT 37.41 6.62 37.76 6.97 ;
      RECT 29.97 6.695 37.76 6.895 ;
      RECT 37.325 3.265 37.585 3.585 ;
      RECT 37.385 1.855 37.525 3.585 ;
      RECT 37.315 1.855 37.595 2.225 ;
      RECT 34.715 4.015 37.15 4.155 ;
      RECT 37.01 2.705 37.15 4.155 ;
      RECT 34.715 3.635 34.855 4.155 ;
      RECT 34.415 3.635 34.855 3.865 ;
      RECT 32.075 3.635 34.855 3.775 ;
      RECT 34.415 3.545 34.675 3.865 ;
      RECT 32.075 3.355 32.215 3.775 ;
      RECT 31.565 3.265 31.825 3.585 ;
      RECT 31.565 3.355 32.215 3.495 ;
      RECT 31.625 1.865 31.765 3.585 ;
      RECT 36.95 2.705 37.21 3.025 ;
      RECT 31.565 1.865 31.825 2.185 ;
      RECT 36.575 3.545 36.835 3.865 ;
      RECT 36.635 1.955 36.775 3.865 ;
      RECT 36.295 1.955 36.775 2.23 ;
      RECT 36.095 1.86 36.575 2.205 ;
      RECT 36.085 3.495 36.365 3.865 ;
      RECT 36.155 2.4 36.295 3.865 ;
      RECT 36.095 2.4 36.355 3.025 ;
      RECT 36.085 2.4 36.365 2.77 ;
      RECT 35.015 3.545 35.275 3.865 ;
      RECT 35.015 3.355 35.215 3.865 ;
      RECT 34.82 3.355 35.215 3.495 ;
      RECT 34.82 1.865 34.96 3.495 ;
      RECT 34.82 1.865 35.135 2.235 ;
      RECT 34.76 1.865 35.135 2.185 ;
      RECT 32.485 2.96 32.765 3.33 ;
      RECT 33.935 2.985 34.195 3.305 ;
      RECT 32.315 3.075 34.195 3.215 ;
      RECT 32.315 2.96 32.765 3.215 ;
      RECT 32.255 2.4 32.515 3.025 ;
      RECT 32.245 2.4 32.525 2.77 ;
      RECT 33.325 2.4 33.735 2.77 ;
      RECT 32.735 2.425 32.995 2.745 ;
      RECT 32.735 2.515 33.735 2.655 ;
      RECT 26.79 6.225 27.11 6.55 ;
      RECT 26.82 5.7 26.99 6.55 ;
      RECT 26.82 5.7 26.995 6.05 ;
      RECT 26.82 5.7 27.795 5.875 ;
      RECT 27.62 1.97 27.795 5.875 ;
      RECT 27.565 1.97 27.915 2.32 ;
      RECT 27.59 6.66 27.915 6.985 ;
      RECT 26.475 6.75 27.915 6.92 ;
      RECT 26.475 2.4 26.635 6.92 ;
      RECT 26.79 2.37 27.11 2.69 ;
      RECT 26.475 2.4 27.11 2.57 ;
      RECT 25.215 2.69 25.505 3.07 ;
      RECT 25.185 2.705 25.525 3.055 ;
      RECT 23.925 3.545 24.185 3.865 ;
      RECT 23.985 1.84 24.125 3.865 ;
      RECT 23.81 2.4 24.125 2.77 ;
      RECT 23.88 1.955 24.125 2.77 ;
      RECT 23.915 1.84 24.195 2.21 ;
      RECT 23.235 2.425 23.495 2.745 ;
      RECT 22.575 2.515 23.495 2.655 ;
      RECT 22.575 1.575 22.715 2.655 ;
      RECT 19.035 1.865 19.295 2.185 ;
      RECT 19.215 1.575 19.355 2.095 ;
      RECT 19.215 1.575 22.715 1.715 ;
      RECT 14.71 6.66 15.06 7.01 ;
      RECT 22.15 6.615 22.5 6.965 ;
      RECT 14.71 6.69 22.5 6.89 ;
      RECT 22.065 3.265 22.325 3.585 ;
      RECT 22.125 1.855 22.265 3.585 ;
      RECT 22.055 1.855 22.335 2.225 ;
      RECT 19.455 4.015 21.89 4.155 ;
      RECT 21.75 2.705 21.89 4.155 ;
      RECT 19.455 3.635 19.595 4.155 ;
      RECT 19.155 3.635 19.595 3.865 ;
      RECT 16.815 3.635 19.595 3.775 ;
      RECT 19.155 3.545 19.415 3.865 ;
      RECT 16.815 3.355 16.955 3.775 ;
      RECT 16.305 3.265 16.565 3.585 ;
      RECT 16.305 3.355 16.955 3.495 ;
      RECT 16.365 1.865 16.505 3.585 ;
      RECT 21.69 2.705 21.95 3.025 ;
      RECT 16.305 1.865 16.565 2.185 ;
      RECT 21.315 3.545 21.575 3.865 ;
      RECT 21.375 1.955 21.515 3.865 ;
      RECT 21.035 1.955 21.515 2.23 ;
      RECT 20.835 1.86 21.315 2.205 ;
      RECT 20.825 3.495 21.105 3.865 ;
      RECT 20.895 2.4 21.035 3.865 ;
      RECT 20.835 2.4 21.095 3.025 ;
      RECT 20.825 2.4 21.105 2.77 ;
      RECT 19.755 3.545 20.015 3.865 ;
      RECT 19.755 3.355 19.955 3.865 ;
      RECT 19.56 3.355 19.955 3.495 ;
      RECT 19.56 1.865 19.7 3.495 ;
      RECT 19.56 1.865 19.875 2.235 ;
      RECT 19.5 1.865 19.875 2.185 ;
      RECT 17.225 2.96 17.505 3.33 ;
      RECT 18.675 2.985 18.935 3.305 ;
      RECT 17.055 3.075 18.935 3.215 ;
      RECT 17.055 2.96 17.505 3.215 ;
      RECT 16.995 2.4 17.255 3.025 ;
      RECT 16.985 2.4 17.265 2.77 ;
      RECT 18.065 2.4 18.475 2.77 ;
      RECT 17.475 2.425 17.735 2.745 ;
      RECT 17.475 2.515 18.475 2.655 ;
      RECT 11.53 6.225 11.85 6.55 ;
      RECT 11.56 5.7 11.73 6.55 ;
      RECT 11.56 5.7 11.735 6.05 ;
      RECT 11.56 5.7 12.535 5.875 ;
      RECT 12.36 1.97 12.535 5.875 ;
      RECT 12.305 1.97 12.655 2.32 ;
      RECT 12.33 6.66 12.655 6.985 ;
      RECT 11.215 6.75 12.655 6.92 ;
      RECT 11.215 2.4 11.375 6.92 ;
      RECT 11.53 2.37 11.85 2.69 ;
      RECT 11.215 2.4 11.85 2.57 ;
      RECT 9.955 2.69 10.245 3.07 ;
      RECT 9.925 2.705 10.265 3.055 ;
      RECT 8.665 3.545 8.925 3.865 ;
      RECT 8.725 1.84 8.865 3.865 ;
      RECT 8.55 2.4 8.865 2.77 ;
      RECT 8.62 1.955 8.865 2.77 ;
      RECT 8.655 1.84 8.935 2.21 ;
      RECT 7.975 2.425 8.235 2.745 ;
      RECT 7.315 2.515 8.235 2.655 ;
      RECT 7.315 1.575 7.455 2.655 ;
      RECT 3.775 1.865 4.035 2.185 ;
      RECT 3.955 1.575 4.095 2.095 ;
      RECT 3.955 1.575 7.455 1.715 ;
      RECT -1.255 7 -0.965 7.35 ;
      RECT -1.255 7.055 0 7.225 ;
      RECT -0.17 6.69 0 7.225 ;
      RECT 6.89 6.61 7.24 6.96 ;
      RECT -0.17 6.69 7.24 6.86 ;
      RECT 6.805 3.265 7.065 3.585 ;
      RECT 6.865 1.855 7.005 3.585 ;
      RECT 6.795 1.855 7.075 2.225 ;
      RECT 4.195 4.015 6.63 4.155 ;
      RECT 6.49 2.705 6.63 4.155 ;
      RECT 4.195 3.635 4.335 4.155 ;
      RECT 3.895 3.635 4.335 3.865 ;
      RECT 1.555 3.635 4.335 3.775 ;
      RECT 3.895 3.545 4.155 3.865 ;
      RECT 1.555 3.355 1.695 3.775 ;
      RECT 1.045 3.265 1.305 3.585 ;
      RECT 1.045 3.355 1.695 3.495 ;
      RECT 1.105 1.865 1.245 3.585 ;
      RECT 6.43 2.705 6.69 3.025 ;
      RECT 1.045 1.865 1.305 2.185 ;
      RECT 6.055 3.545 6.315 3.865 ;
      RECT 6.115 1.955 6.255 3.865 ;
      RECT 5.775 1.955 6.255 2.23 ;
      RECT 5.575 1.86 6.055 2.205 ;
      RECT 5.565 3.495 5.845 3.865 ;
      RECT 5.635 2.4 5.775 3.865 ;
      RECT 5.575 2.4 5.835 3.025 ;
      RECT 5.565 2.4 5.845 2.77 ;
      RECT 4.495 3.545 4.755 3.865 ;
      RECT 4.495 3.355 4.695 3.865 ;
      RECT 4.3 3.355 4.695 3.495 ;
      RECT 4.3 1.865 4.44 3.495 ;
      RECT 4.3 1.865 4.615 2.235 ;
      RECT 4.24 1.865 4.615 2.185 ;
      RECT 1.965 2.96 2.245 3.33 ;
      RECT 3.415 2.985 3.675 3.305 ;
      RECT 1.795 3.075 3.675 3.215 ;
      RECT 1.795 2.96 2.245 3.215 ;
      RECT 1.735 2.4 1.995 3.025 ;
      RECT 1.725 2.4 2.005 2.77 ;
      RECT 2.805 2.4 3.215 2.77 ;
      RECT 2.215 2.425 2.475 2.745 ;
      RECT 2.215 2.515 3.215 2.655 ;
      RECT 67.26 7.06 67.63 7.43 ;
      RECT 66.125 2.4 66.405 2.865 ;
      RECT 65.885 1.865 66.165 2.21 ;
      RECT 64.685 2.4 64.965 2.77 ;
      RECT 62.125 1.22 62.495 1.225 ;
      RECT 52 7.06 52.37 7.43 ;
      RECT 50.865 2.4 51.145 2.865 ;
      RECT 50.625 1.865 50.905 2.21 ;
      RECT 49.425 2.4 49.705 2.77 ;
      RECT 46.865 1.22 47.235 1.225 ;
      RECT 36.74 7.06 37.11 7.43 ;
      RECT 35.605 2.4 35.885 2.865 ;
      RECT 35.365 1.865 35.645 2.21 ;
      RECT 34.165 2.4 34.445 2.77 ;
      RECT 31.605 1.22 31.975 1.225 ;
      RECT 21.48 7.06 21.85 7.43 ;
      RECT 20.345 2.4 20.625 2.865 ;
      RECT 20.105 1.865 20.385 2.21 ;
      RECT 18.905 2.4 19.185 2.77 ;
      RECT 16.345 1.22 16.715 1.225 ;
      RECT 6.22 7.06 6.59 7.43 ;
      RECT 5.085 2.4 5.365 2.865 ;
      RECT 4.845 1.865 5.125 2.21 ;
      RECT 3.645 2.4 3.925 2.77 ;
      RECT 1.085 1.22 1.455 1.225 ;
    LAYER via1 ;
      RECT 75.83 7.38 75.98 7.53 ;
      RECT 73.46 6.745 73.61 6.895 ;
      RECT 73.445 2.07 73.595 2.22 ;
      RECT 72.655 2.455 72.805 2.605 ;
      RECT 72.655 6.33 72.805 6.48 ;
      RECT 71.065 2.805 71.215 2.955 ;
      RECT 69.76 1.95 69.91 2.1 ;
      RECT 69.76 3.63 69.91 3.78 ;
      RECT 69.07 2.51 69.22 2.66 ;
      RECT 68.03 6.715 68.18 6.865 ;
      RECT 67.9 1.95 68.05 2.1 ;
      RECT 67.9 3.35 68.05 3.5 ;
      RECT 67.525 2.79 67.675 2.94 ;
      RECT 67.37 7.17 67.52 7.32 ;
      RECT 67.15 3.63 67.3 3.78 ;
      RECT 66.67 1.95 66.82 2.1 ;
      RECT 66.67 2.79 66.82 2.94 ;
      RECT 66.19 2.51 66.34 2.66 ;
      RECT 65.95 1.95 66.1 2.1 ;
      RECT 65.59 3.63 65.74 3.78 ;
      RECT 65.335 1.95 65.485 2.1 ;
      RECT 64.99 3.63 65.14 3.78 ;
      RECT 64.87 1.95 65.02 2.1 ;
      RECT 64.75 2.51 64.9 2.66 ;
      RECT 64.51 3.07 64.66 3.22 ;
      RECT 63.31 2.51 63.46 2.66 ;
      RECT 62.83 2.79 62.98 2.94 ;
      RECT 62.14 1.95 62.29 2.1 ;
      RECT 62.14 3.35 62.29 3.5 ;
      RECT 60.545 6.76 60.695 6.91 ;
      RECT 58.2 6.745 58.35 6.895 ;
      RECT 58.185 2.07 58.335 2.22 ;
      RECT 57.395 2.455 57.545 2.605 ;
      RECT 57.395 6.33 57.545 6.48 ;
      RECT 55.805 2.805 55.955 2.955 ;
      RECT 54.5 1.95 54.65 2.1 ;
      RECT 54.5 3.63 54.65 3.78 ;
      RECT 53.81 2.51 53.96 2.66 ;
      RECT 52.775 6.715 52.925 6.865 ;
      RECT 52.64 1.95 52.79 2.1 ;
      RECT 52.64 3.35 52.79 3.5 ;
      RECT 52.265 2.79 52.415 2.94 ;
      RECT 52.11 7.17 52.26 7.32 ;
      RECT 51.89 3.63 52.04 3.78 ;
      RECT 51.41 1.95 51.56 2.1 ;
      RECT 51.41 2.79 51.56 2.94 ;
      RECT 50.93 2.51 51.08 2.66 ;
      RECT 50.69 1.95 50.84 2.1 ;
      RECT 50.33 3.63 50.48 3.78 ;
      RECT 50.075 1.95 50.225 2.1 ;
      RECT 49.73 3.63 49.88 3.78 ;
      RECT 49.61 1.95 49.76 2.1 ;
      RECT 49.49 2.51 49.64 2.66 ;
      RECT 49.25 3.07 49.4 3.22 ;
      RECT 48.05 2.51 48.2 2.66 ;
      RECT 47.57 2.79 47.72 2.94 ;
      RECT 46.88 1.95 47.03 2.1 ;
      RECT 46.88 3.35 47.03 3.5 ;
      RECT 45.285 6.76 45.435 6.91 ;
      RECT 42.94 6.745 43.09 6.895 ;
      RECT 42.925 2.07 43.075 2.22 ;
      RECT 42.135 2.455 42.285 2.605 ;
      RECT 42.135 6.33 42.285 6.48 ;
      RECT 40.545 2.805 40.695 2.955 ;
      RECT 39.24 1.95 39.39 2.1 ;
      RECT 39.24 3.63 39.39 3.78 ;
      RECT 38.55 2.51 38.7 2.66 ;
      RECT 37.51 6.72 37.66 6.87 ;
      RECT 37.38 1.95 37.53 2.1 ;
      RECT 37.38 3.35 37.53 3.5 ;
      RECT 37.005 2.79 37.155 2.94 ;
      RECT 36.85 7.17 37 7.32 ;
      RECT 36.63 3.63 36.78 3.78 ;
      RECT 36.15 1.95 36.3 2.1 ;
      RECT 36.15 2.79 36.3 2.94 ;
      RECT 35.67 2.51 35.82 2.66 ;
      RECT 35.43 1.95 35.58 2.1 ;
      RECT 35.07 3.63 35.22 3.78 ;
      RECT 34.815 1.95 34.965 2.1 ;
      RECT 34.47 3.63 34.62 3.78 ;
      RECT 34.35 1.95 34.5 2.1 ;
      RECT 34.23 2.51 34.38 2.66 ;
      RECT 33.99 3.07 34.14 3.22 ;
      RECT 32.79 2.51 32.94 2.66 ;
      RECT 32.31 2.79 32.46 2.94 ;
      RECT 31.62 1.95 31.77 2.1 ;
      RECT 31.62 3.35 31.77 3.5 ;
      RECT 30.07 6.765 30.22 6.915 ;
      RECT 27.68 6.745 27.83 6.895 ;
      RECT 27.665 2.07 27.815 2.22 ;
      RECT 26.875 2.455 27.025 2.605 ;
      RECT 26.875 6.33 27.025 6.48 ;
      RECT 25.285 2.805 25.435 2.955 ;
      RECT 23.98 1.95 24.13 2.1 ;
      RECT 23.98 3.63 24.13 3.78 ;
      RECT 23.29 2.51 23.44 2.66 ;
      RECT 22.25 6.715 22.4 6.865 ;
      RECT 22.12 1.95 22.27 2.1 ;
      RECT 22.12 3.35 22.27 3.5 ;
      RECT 21.745 2.79 21.895 2.94 ;
      RECT 21.59 7.17 21.74 7.32 ;
      RECT 21.37 3.63 21.52 3.78 ;
      RECT 20.89 1.95 21.04 2.1 ;
      RECT 20.89 2.79 21.04 2.94 ;
      RECT 20.41 2.51 20.56 2.66 ;
      RECT 20.17 1.95 20.32 2.1 ;
      RECT 19.81 3.63 19.96 3.78 ;
      RECT 19.555 1.95 19.705 2.1 ;
      RECT 19.21 3.63 19.36 3.78 ;
      RECT 19.09 1.95 19.24 2.1 ;
      RECT 18.97 2.51 19.12 2.66 ;
      RECT 18.73 3.07 18.88 3.22 ;
      RECT 17.53 2.51 17.68 2.66 ;
      RECT 17.05 2.79 17.2 2.94 ;
      RECT 16.36 1.95 16.51 2.1 ;
      RECT 16.36 3.35 16.51 3.5 ;
      RECT 14.81 6.76 14.96 6.91 ;
      RECT 12.42 6.745 12.57 6.895 ;
      RECT 12.405 2.07 12.555 2.22 ;
      RECT 11.615 2.455 11.765 2.605 ;
      RECT 11.615 6.33 11.765 6.48 ;
      RECT 10.025 2.805 10.175 2.955 ;
      RECT 8.72 1.95 8.87 2.1 ;
      RECT 8.72 3.63 8.87 3.78 ;
      RECT 8.03 2.51 8.18 2.66 ;
      RECT 6.99 6.71 7.14 6.86 ;
      RECT 6.86 1.95 7.01 2.1 ;
      RECT 6.86 3.35 7.01 3.5 ;
      RECT 6.485 2.79 6.635 2.94 ;
      RECT 6.33 7.17 6.48 7.32 ;
      RECT 6.11 3.63 6.26 3.78 ;
      RECT 5.63 1.95 5.78 2.1 ;
      RECT 5.63 2.79 5.78 2.94 ;
      RECT 5.15 2.51 5.3 2.66 ;
      RECT 4.91 1.95 5.06 2.1 ;
      RECT 4.55 3.63 4.7 3.78 ;
      RECT 4.295 1.95 4.445 2.1 ;
      RECT 3.95 3.63 4.1 3.78 ;
      RECT 3.83 1.95 3.98 2.1 ;
      RECT 3.71 2.51 3.86 2.66 ;
      RECT 3.47 3.07 3.62 3.22 ;
      RECT 2.27 2.51 2.42 2.66 ;
      RECT 1.79 2.79 1.94 2.94 ;
      RECT 1.1 1.95 1.25 2.1 ;
      RECT 1.1 3.35 1.25 3.5 ;
      RECT -1.185 7.1 -1.035 7.25 ;
      RECT -1.56 6.36 -1.41 6.51 ;
    LAYER met1 ;
      RECT 75.695 7.775 75.985 8.005 ;
      RECT 75.755 6.295 75.925 8.005 ;
      RECT 75.73 7.28 76.08 7.63 ;
      RECT 75.695 6.295 75.985 6.525 ;
      RECT 75.29 2.4 75.395 2.97 ;
      RECT 75.29 2.735 75.615 2.965 ;
      RECT 75.29 2.765 75.785 2.935 ;
      RECT 75.29 2.4 75.48 2.965 ;
      RECT 74.705 2.365 74.995 2.595 ;
      RECT 74.705 2.4 75.48 2.57 ;
      RECT 74.765 0.885 74.935 2.595 ;
      RECT 74.705 0.885 74.995 1.115 ;
      RECT 74.705 7.775 74.995 8.005 ;
      RECT 74.765 6.295 74.935 8.005 ;
      RECT 74.705 6.295 74.995 6.525 ;
      RECT 74.705 6.33 75.56 6.49 ;
      RECT 75.39 5.925 75.56 6.49 ;
      RECT 74.705 6.325 75.1 6.49 ;
      RECT 75.325 5.925 75.615 6.155 ;
      RECT 75.325 5.955 75.785 6.125 ;
      RECT 74.335 2.735 74.625 2.965 ;
      RECT 74.335 2.765 74.795 2.935 ;
      RECT 74.4 1.66 74.565 2.965 ;
      RECT 72.915 1.63 73.205 1.86 ;
      RECT 72.915 1.66 74.565 1.83 ;
      RECT 72.975 0.89 73.145 1.86 ;
      RECT 72.915 0.89 73.205 1.12 ;
      RECT 72.915 7.77 73.205 8 ;
      RECT 72.975 7.03 73.145 8 ;
      RECT 72.975 7.125 74.565 7.295 ;
      RECT 74.395 5.925 74.565 7.295 ;
      RECT 72.915 7.03 73.205 7.26 ;
      RECT 74.335 5.925 74.625 6.155 ;
      RECT 74.335 5.955 74.795 6.125 ;
      RECT 70.965 2.705 71.305 3.055 ;
      RECT 71.055 2.03 71.225 3.055 ;
      RECT 73.345 1.97 73.695 2.32 ;
      RECT 71.055 2.03 73.695 2.2 ;
      RECT 73.37 6.66 73.695 6.985 ;
      RECT 67.93 6.615 68.28 6.965 ;
      RECT 73.345 6.66 73.695 6.89 ;
      RECT 67.73 6.66 68.28 6.89 ;
      RECT 67.56 6.69 73.695 6.86 ;
      RECT 72.57 2.37 72.89 2.69 ;
      RECT 72.54 2.37 72.89 2.6 ;
      RECT 72.37 2.4 72.89 2.57 ;
      RECT 72.57 6.26 72.89 6.55 ;
      RECT 72.54 6.29 72.89 6.52 ;
      RECT 72.37 6.32 72.89 6.49 ;
      RECT 69.675 1.895 69.995 2.155 ;
      RECT 69.24 1.91 69.53 2.14 ;
      RECT 69.24 1.955 69.995 2.095 ;
      RECT 69.675 3.575 69.995 3.835 ;
      RECT 69.24 3.59 69.53 3.82 ;
      RECT 69.24 3.635 69.995 3.775 ;
      RECT 69 3.03 69.29 3.26 ;
      RECT 69 3.075 69.575 3.215 ;
      RECT 69.435 2.935 69.695 3.075 ;
      RECT 69.48 2.75 69.77 2.98 ;
      RECT 67.635 2.935 68.735 3.075 ;
      RECT 67.44 2.735 67.76 2.995 ;
      RECT 68.52 2.75 68.81 2.98 ;
      RECT 67.44 2.75 67.85 2.995 ;
      RECT 67.815 1.895 68.135 2.155 ;
      RECT 68.28 1.91 68.57 2.14 ;
      RECT 67.815 1.955 68.57 2.095 ;
      RECT 65.115 3.16 67.295 3.3 ;
      RECT 67.155 2.17 67.295 3.3 ;
      RECT 65.115 3.075 66.41 3.3 ;
      RECT 66.12 3.03 66.41 3.3 ;
      RECT 65.115 2.795 65.45 3.3 ;
      RECT 65.16 2.75 65.45 3.3 ;
      RECT 68.04 2.47 68.33 2.7 ;
      RECT 67.155 2.375 68.255 2.515 ;
      RECT 67.08 2.17 67.37 2.42 ;
      RECT 67.3 7.77 67.59 8 ;
      RECT 67.36 7.03 67.53 8 ;
      RECT 67.26 7.06 67.63 7.43 ;
      RECT 67.3 7.03 67.59 7.43 ;
      RECT 67.065 3.575 67.385 3.835 ;
      RECT 67.065 3.59 67.58 3.82 ;
      RECT 65.64 2.47 65.93 2.7 ;
      RECT 65.79 2.075 65.93 2.7 ;
      RECT 65.79 2.075 66.095 2.215 ;
      RECT 66.585 1.895 66.905 2.155 ;
      RECT 65.865 1.895 66.185 2.155 ;
      RECT 66.36 1.91 66.905 2.14 ;
      RECT 65.865 1.955 66.905 2.095 ;
      RECT 65.505 3.575 65.825 3.835 ;
      RECT 65.4 3.59 65.825 3.82 ;
      RECT 63.48 3.03 63.77 3.26 ;
      RECT 63.48 3.03 63.935 3.215 ;
      RECT 63.795 2.555 63.935 3.215 ;
      RECT 63.915 1.955 64.055 2.695 ;
      RECT 64.785 1.895 65.105 2.155 ;
      RECT 63.96 1.91 64.25 2.14 ;
      RECT 63.915 1.955 65.105 2.095 ;
      RECT 64.665 2.455 64.985 2.715 ;
      RECT 64.2 2.47 64.49 2.7 ;
      RECT 64.2 2.515 64.985 2.655 ;
      RECT 64.425 3.015 64.745 3.275 ;
      RECT 64.425 3.03 64.97 3.26 ;
      RECT 63.96 3.59 64.25 3.82 ;
      RECT 63.075 3.47 64.175 3.61 ;
      RECT 63 3.31 63.29 3.54 ;
      RECT 60.435 7.775 60.725 8.005 ;
      RECT 60.495 6.295 60.665 8.005 ;
      RECT 60.445 6.66 60.795 7.01 ;
      RECT 60.435 6.295 60.725 6.525 ;
      RECT 60.03 2.4 60.135 2.97 ;
      RECT 60.03 2.735 60.355 2.965 ;
      RECT 60.03 2.765 60.525 2.935 ;
      RECT 60.03 2.4 60.22 2.965 ;
      RECT 59.445 2.365 59.735 2.595 ;
      RECT 59.445 2.4 60.22 2.57 ;
      RECT 59.505 0.885 59.675 2.595 ;
      RECT 59.445 0.885 59.735 1.115 ;
      RECT 59.445 7.775 59.735 8.005 ;
      RECT 59.505 6.295 59.675 8.005 ;
      RECT 59.445 6.295 59.735 6.525 ;
      RECT 59.445 6.33 60.3 6.49 ;
      RECT 60.13 5.925 60.3 6.49 ;
      RECT 59.445 6.325 59.84 6.49 ;
      RECT 60.065 5.925 60.355 6.155 ;
      RECT 60.065 5.955 60.525 6.125 ;
      RECT 59.075 2.735 59.365 2.965 ;
      RECT 59.075 2.765 59.535 2.935 ;
      RECT 59.14 1.66 59.305 2.965 ;
      RECT 57.655 1.63 57.945 1.86 ;
      RECT 57.655 1.66 59.305 1.83 ;
      RECT 57.715 0.89 57.885 1.86 ;
      RECT 57.655 0.89 57.945 1.12 ;
      RECT 57.655 7.77 57.945 8 ;
      RECT 57.715 7.03 57.885 8 ;
      RECT 57.715 7.125 59.305 7.295 ;
      RECT 59.135 5.925 59.305 7.295 ;
      RECT 57.655 7.03 57.945 7.26 ;
      RECT 59.075 5.925 59.365 6.155 ;
      RECT 59.075 5.955 59.535 6.125 ;
      RECT 55.705 2.705 56.045 3.055 ;
      RECT 55.795 2.03 55.965 3.055 ;
      RECT 58.085 1.97 58.435 2.32 ;
      RECT 55.795 2.03 58.435 2.2 ;
      RECT 58.11 6.66 58.435 6.985 ;
      RECT 52.675 6.615 53.025 6.965 ;
      RECT 58.085 6.66 58.435 6.89 ;
      RECT 52.47 6.66 53.025 6.89 ;
      RECT 52.3 6.69 58.435 6.86 ;
      RECT 57.31 2.37 57.63 2.69 ;
      RECT 57.28 2.37 57.63 2.6 ;
      RECT 57.11 2.4 57.63 2.57 ;
      RECT 57.31 6.26 57.63 6.55 ;
      RECT 57.28 6.29 57.63 6.52 ;
      RECT 57.11 6.32 57.63 6.49 ;
      RECT 54.415 1.895 54.735 2.155 ;
      RECT 53.98 1.91 54.27 2.14 ;
      RECT 53.98 1.955 54.735 2.095 ;
      RECT 54.415 3.575 54.735 3.835 ;
      RECT 53.98 3.59 54.27 3.82 ;
      RECT 53.98 3.635 54.735 3.775 ;
      RECT 53.74 3.03 54.03 3.26 ;
      RECT 53.74 3.075 54.315 3.215 ;
      RECT 54.175 2.935 54.435 3.075 ;
      RECT 54.22 2.75 54.51 2.98 ;
      RECT 52.375 2.935 53.475 3.075 ;
      RECT 52.18 2.735 52.5 2.995 ;
      RECT 53.26 2.75 53.55 2.98 ;
      RECT 52.18 2.75 52.59 2.995 ;
      RECT 52.555 1.895 52.875 2.155 ;
      RECT 53.02 1.91 53.31 2.14 ;
      RECT 52.555 1.955 53.31 2.095 ;
      RECT 49.855 3.16 52.035 3.3 ;
      RECT 51.895 2.17 52.035 3.3 ;
      RECT 49.855 3.075 51.15 3.3 ;
      RECT 50.86 3.03 51.15 3.3 ;
      RECT 49.855 2.795 50.19 3.3 ;
      RECT 49.9 2.75 50.19 3.3 ;
      RECT 52.78 2.47 53.07 2.7 ;
      RECT 51.895 2.375 52.995 2.515 ;
      RECT 51.82 2.17 52.11 2.42 ;
      RECT 52.04 7.77 52.33 8 ;
      RECT 52.1 7.03 52.27 8 ;
      RECT 52 7.06 52.37 7.43 ;
      RECT 52.04 7.03 52.33 7.43 ;
      RECT 51.805 3.575 52.125 3.835 ;
      RECT 51.805 3.59 52.32 3.82 ;
      RECT 50.38 2.47 50.67 2.7 ;
      RECT 50.53 2.075 50.67 2.7 ;
      RECT 50.53 2.075 50.835 2.215 ;
      RECT 51.325 1.895 51.645 2.155 ;
      RECT 50.605 1.895 50.925 2.155 ;
      RECT 51.1 1.91 51.645 2.14 ;
      RECT 50.605 1.955 51.645 2.095 ;
      RECT 50.245 3.575 50.565 3.835 ;
      RECT 50.14 3.59 50.565 3.82 ;
      RECT 48.22 3.03 48.51 3.26 ;
      RECT 48.22 3.03 48.675 3.215 ;
      RECT 48.535 2.555 48.675 3.215 ;
      RECT 48.655 1.955 48.795 2.695 ;
      RECT 49.525 1.895 49.845 2.155 ;
      RECT 48.7 1.91 48.99 2.14 ;
      RECT 48.655 1.955 49.845 2.095 ;
      RECT 49.405 2.455 49.725 2.715 ;
      RECT 48.94 2.47 49.23 2.7 ;
      RECT 48.94 2.515 49.725 2.655 ;
      RECT 49.165 3.015 49.485 3.275 ;
      RECT 49.165 3.03 49.71 3.26 ;
      RECT 48.7 3.59 48.99 3.82 ;
      RECT 47.815 3.47 48.915 3.61 ;
      RECT 47.74 3.31 48.03 3.54 ;
      RECT 45.175 7.775 45.465 8.005 ;
      RECT 45.235 6.295 45.405 8.005 ;
      RECT 45.185 6.66 45.535 7.01 ;
      RECT 45.175 6.295 45.465 6.525 ;
      RECT 44.77 2.4 44.875 2.97 ;
      RECT 44.77 2.735 45.095 2.965 ;
      RECT 44.77 2.765 45.265 2.935 ;
      RECT 44.77 2.4 44.96 2.965 ;
      RECT 44.185 2.365 44.475 2.595 ;
      RECT 44.185 2.4 44.96 2.57 ;
      RECT 44.245 0.885 44.415 2.595 ;
      RECT 44.185 0.885 44.475 1.115 ;
      RECT 44.185 7.775 44.475 8.005 ;
      RECT 44.245 6.295 44.415 8.005 ;
      RECT 44.185 6.295 44.475 6.525 ;
      RECT 44.185 6.33 45.04 6.49 ;
      RECT 44.87 5.925 45.04 6.49 ;
      RECT 44.185 6.325 44.58 6.49 ;
      RECT 44.805 5.925 45.095 6.155 ;
      RECT 44.805 5.955 45.265 6.125 ;
      RECT 43.815 2.735 44.105 2.965 ;
      RECT 43.815 2.765 44.275 2.935 ;
      RECT 43.88 1.66 44.045 2.965 ;
      RECT 42.395 1.63 42.685 1.86 ;
      RECT 42.395 1.66 44.045 1.83 ;
      RECT 42.455 0.89 42.625 1.86 ;
      RECT 42.395 0.89 42.685 1.12 ;
      RECT 42.395 7.77 42.685 8 ;
      RECT 42.455 7.03 42.625 8 ;
      RECT 42.455 7.125 44.045 7.295 ;
      RECT 43.875 5.925 44.045 7.295 ;
      RECT 42.395 7.03 42.685 7.26 ;
      RECT 43.815 5.925 44.105 6.155 ;
      RECT 43.815 5.955 44.275 6.125 ;
      RECT 40.445 2.705 40.785 3.055 ;
      RECT 40.535 2.03 40.705 3.055 ;
      RECT 42.825 1.97 43.175 2.32 ;
      RECT 40.535 2.03 43.175 2.2 ;
      RECT 42.85 6.66 43.175 6.985 ;
      RECT 37.41 6.62 37.76 6.97 ;
      RECT 42.825 6.66 43.175 6.89 ;
      RECT 37.21 6.66 37.76 6.89 ;
      RECT 37.04 6.69 43.175 6.86 ;
      RECT 42.05 2.37 42.37 2.69 ;
      RECT 42.02 2.37 42.37 2.6 ;
      RECT 41.85 2.4 42.37 2.57 ;
      RECT 42.05 6.26 42.37 6.55 ;
      RECT 42.02 6.29 42.37 6.52 ;
      RECT 41.85 6.32 42.37 6.49 ;
      RECT 39.155 1.895 39.475 2.155 ;
      RECT 38.72 1.91 39.01 2.14 ;
      RECT 38.72 1.955 39.475 2.095 ;
      RECT 39.155 3.575 39.475 3.835 ;
      RECT 38.72 3.59 39.01 3.82 ;
      RECT 38.72 3.635 39.475 3.775 ;
      RECT 38.48 3.03 38.77 3.26 ;
      RECT 38.48 3.075 39.055 3.215 ;
      RECT 38.915 2.935 39.175 3.075 ;
      RECT 38.96 2.75 39.25 2.98 ;
      RECT 37.115 2.935 38.215 3.075 ;
      RECT 36.92 2.735 37.24 2.995 ;
      RECT 38 2.75 38.29 2.98 ;
      RECT 36.92 2.75 37.33 2.995 ;
      RECT 37.295 1.895 37.615 2.155 ;
      RECT 37.76 1.91 38.05 2.14 ;
      RECT 37.295 1.955 38.05 2.095 ;
      RECT 34.595 3.16 36.775 3.3 ;
      RECT 36.635 2.17 36.775 3.3 ;
      RECT 34.595 3.075 35.89 3.3 ;
      RECT 35.6 3.03 35.89 3.3 ;
      RECT 34.595 2.795 34.93 3.3 ;
      RECT 34.64 2.75 34.93 3.3 ;
      RECT 37.52 2.47 37.81 2.7 ;
      RECT 36.635 2.375 37.735 2.515 ;
      RECT 36.56 2.17 36.85 2.42 ;
      RECT 36.78 7.77 37.07 8 ;
      RECT 36.84 7.03 37.01 8 ;
      RECT 36.74 7.06 37.11 7.43 ;
      RECT 36.78 7.03 37.07 7.43 ;
      RECT 36.545 3.575 36.865 3.835 ;
      RECT 36.545 3.59 37.06 3.82 ;
      RECT 35.12 2.47 35.41 2.7 ;
      RECT 35.27 2.075 35.41 2.7 ;
      RECT 35.27 2.075 35.575 2.215 ;
      RECT 36.065 1.895 36.385 2.155 ;
      RECT 35.345 1.895 35.665 2.155 ;
      RECT 35.84 1.91 36.385 2.14 ;
      RECT 35.345 1.955 36.385 2.095 ;
      RECT 34.985 3.575 35.305 3.835 ;
      RECT 34.88 3.59 35.305 3.82 ;
      RECT 32.96 3.03 33.25 3.26 ;
      RECT 32.96 3.03 33.415 3.215 ;
      RECT 33.275 2.555 33.415 3.215 ;
      RECT 33.395 1.955 33.535 2.695 ;
      RECT 34.265 1.895 34.585 2.155 ;
      RECT 33.44 1.91 33.73 2.14 ;
      RECT 33.395 1.955 34.585 2.095 ;
      RECT 34.145 2.455 34.465 2.715 ;
      RECT 33.68 2.47 33.97 2.7 ;
      RECT 33.68 2.515 34.465 2.655 ;
      RECT 33.905 3.015 34.225 3.275 ;
      RECT 33.905 3.03 34.45 3.26 ;
      RECT 33.44 3.59 33.73 3.82 ;
      RECT 32.555 3.47 33.655 3.61 ;
      RECT 32.48 3.31 32.77 3.54 ;
      RECT 29.915 7.775 30.205 8.005 ;
      RECT 29.975 6.295 30.145 8.005 ;
      RECT 29.965 6.665 30.32 7.02 ;
      RECT 29.915 6.295 30.205 6.525 ;
      RECT 29.51 2.4 29.615 2.97 ;
      RECT 29.51 2.735 29.835 2.965 ;
      RECT 29.51 2.765 30.005 2.935 ;
      RECT 29.51 2.4 29.7 2.965 ;
      RECT 28.925 2.365 29.215 2.595 ;
      RECT 28.925 2.4 29.7 2.57 ;
      RECT 28.985 0.885 29.155 2.595 ;
      RECT 28.925 0.885 29.215 1.115 ;
      RECT 28.925 7.775 29.215 8.005 ;
      RECT 28.985 6.295 29.155 8.005 ;
      RECT 28.925 6.295 29.215 6.525 ;
      RECT 28.925 6.33 29.78 6.49 ;
      RECT 29.61 5.925 29.78 6.49 ;
      RECT 28.925 6.325 29.32 6.49 ;
      RECT 29.545 5.925 29.835 6.155 ;
      RECT 29.545 5.955 30.005 6.125 ;
      RECT 28.555 2.735 28.845 2.965 ;
      RECT 28.555 2.765 29.015 2.935 ;
      RECT 28.62 1.66 28.785 2.965 ;
      RECT 27.135 1.63 27.425 1.86 ;
      RECT 27.135 1.66 28.785 1.83 ;
      RECT 27.195 0.89 27.365 1.86 ;
      RECT 27.135 0.89 27.425 1.12 ;
      RECT 27.135 7.77 27.425 8 ;
      RECT 27.195 7.03 27.365 8 ;
      RECT 27.195 7.125 28.785 7.295 ;
      RECT 28.615 5.925 28.785 7.295 ;
      RECT 27.135 7.03 27.425 7.26 ;
      RECT 28.555 5.925 28.845 6.155 ;
      RECT 28.555 5.955 29.015 6.125 ;
      RECT 25.185 2.705 25.525 3.055 ;
      RECT 25.275 2.03 25.445 3.055 ;
      RECT 27.565 1.97 27.915 2.32 ;
      RECT 25.275 2.03 27.915 2.2 ;
      RECT 27.59 6.66 27.915 6.985 ;
      RECT 22.15 6.615 22.5 6.965 ;
      RECT 27.565 6.66 27.915 6.89 ;
      RECT 21.95 6.66 22.5 6.89 ;
      RECT 21.78 6.69 27.915 6.86 ;
      RECT 26.79 2.37 27.11 2.69 ;
      RECT 26.76 2.37 27.11 2.6 ;
      RECT 26.59 2.4 27.11 2.57 ;
      RECT 26.79 6.26 27.11 6.55 ;
      RECT 26.76 6.29 27.11 6.52 ;
      RECT 26.59 6.32 27.11 6.49 ;
      RECT 23.895 1.895 24.215 2.155 ;
      RECT 23.46 1.91 23.75 2.14 ;
      RECT 23.46 1.955 24.215 2.095 ;
      RECT 23.895 3.575 24.215 3.835 ;
      RECT 23.46 3.59 23.75 3.82 ;
      RECT 23.46 3.635 24.215 3.775 ;
      RECT 23.22 3.03 23.51 3.26 ;
      RECT 23.22 3.075 23.795 3.215 ;
      RECT 23.655 2.935 23.915 3.075 ;
      RECT 23.7 2.75 23.99 2.98 ;
      RECT 21.855 2.935 22.955 3.075 ;
      RECT 21.66 2.735 21.98 2.995 ;
      RECT 22.74 2.75 23.03 2.98 ;
      RECT 21.66 2.75 22.07 2.995 ;
      RECT 22.035 1.895 22.355 2.155 ;
      RECT 22.5 1.91 22.79 2.14 ;
      RECT 22.035 1.955 22.79 2.095 ;
      RECT 19.335 3.16 21.515 3.3 ;
      RECT 21.375 2.17 21.515 3.3 ;
      RECT 19.335 3.075 20.63 3.3 ;
      RECT 20.34 3.03 20.63 3.3 ;
      RECT 19.335 2.795 19.67 3.3 ;
      RECT 19.38 2.75 19.67 3.3 ;
      RECT 22.26 2.47 22.55 2.7 ;
      RECT 21.375 2.375 22.475 2.515 ;
      RECT 21.3 2.17 21.59 2.42 ;
      RECT 21.52 7.77 21.81 8 ;
      RECT 21.58 7.03 21.75 8 ;
      RECT 21.48 7.06 21.85 7.43 ;
      RECT 21.52 7.03 21.81 7.43 ;
      RECT 21.285 3.575 21.605 3.835 ;
      RECT 21.285 3.59 21.8 3.82 ;
      RECT 19.86 2.47 20.15 2.7 ;
      RECT 20.01 2.075 20.15 2.7 ;
      RECT 20.01 2.075 20.315 2.215 ;
      RECT 20.805 1.895 21.125 2.155 ;
      RECT 20.085 1.895 20.405 2.155 ;
      RECT 20.58 1.91 21.125 2.14 ;
      RECT 20.085 1.955 21.125 2.095 ;
      RECT 19.725 3.575 20.045 3.835 ;
      RECT 19.62 3.59 20.045 3.82 ;
      RECT 17.7 3.03 17.99 3.26 ;
      RECT 17.7 3.03 18.155 3.215 ;
      RECT 18.015 2.555 18.155 3.215 ;
      RECT 18.135 1.955 18.275 2.695 ;
      RECT 19.005 1.895 19.325 2.155 ;
      RECT 18.18 1.91 18.47 2.14 ;
      RECT 18.135 1.955 19.325 2.095 ;
      RECT 18.885 2.455 19.205 2.715 ;
      RECT 18.42 2.47 18.71 2.7 ;
      RECT 18.42 2.515 19.205 2.655 ;
      RECT 18.645 3.015 18.965 3.275 ;
      RECT 18.645 3.03 19.19 3.26 ;
      RECT 18.18 3.59 18.47 3.82 ;
      RECT 17.295 3.47 18.395 3.61 ;
      RECT 17.22 3.31 17.51 3.54 ;
      RECT 14.655 7.775 14.945 8.005 ;
      RECT 14.715 6.295 14.885 8.005 ;
      RECT 14.71 6.66 15.06 7.01 ;
      RECT 14.655 6.295 14.945 6.525 ;
      RECT 14.25 2.4 14.355 2.97 ;
      RECT 14.25 2.735 14.575 2.965 ;
      RECT 14.25 2.765 14.745 2.935 ;
      RECT 14.25 2.4 14.44 2.965 ;
      RECT 13.665 2.365 13.955 2.595 ;
      RECT 13.665 2.4 14.44 2.57 ;
      RECT 13.725 0.885 13.895 2.595 ;
      RECT 13.665 0.885 13.955 1.115 ;
      RECT 13.665 7.775 13.955 8.005 ;
      RECT 13.725 6.295 13.895 8.005 ;
      RECT 13.665 6.295 13.955 6.525 ;
      RECT 13.665 6.33 14.52 6.49 ;
      RECT 14.35 5.925 14.52 6.49 ;
      RECT 13.665 6.325 14.06 6.49 ;
      RECT 14.285 5.925 14.575 6.155 ;
      RECT 14.285 5.955 14.745 6.125 ;
      RECT 13.295 2.735 13.585 2.965 ;
      RECT 13.295 2.765 13.755 2.935 ;
      RECT 13.36 1.66 13.525 2.965 ;
      RECT 11.875 1.63 12.165 1.86 ;
      RECT 11.875 1.66 13.525 1.83 ;
      RECT 11.935 0.89 12.105 1.86 ;
      RECT 11.875 0.89 12.165 1.12 ;
      RECT 11.875 7.77 12.165 8 ;
      RECT 11.935 7.03 12.105 8 ;
      RECT 11.935 7.125 13.525 7.295 ;
      RECT 13.355 5.925 13.525 7.295 ;
      RECT 11.875 7.03 12.165 7.26 ;
      RECT 13.295 5.925 13.585 6.155 ;
      RECT 13.295 5.955 13.755 6.125 ;
      RECT 9.925 2.705 10.265 3.055 ;
      RECT 10.015 2.03 10.185 3.055 ;
      RECT 12.305 1.97 12.655 2.32 ;
      RECT 10.015 2.03 12.655 2.2 ;
      RECT 12.33 6.66 12.655 6.985 ;
      RECT 6.89 6.61 7.24 6.96 ;
      RECT 12.305 6.66 12.655 6.89 ;
      RECT 6.69 6.66 7.24 6.89 ;
      RECT 6.52 6.69 12.655 6.86 ;
      RECT 11.53 2.37 11.85 2.69 ;
      RECT 11.5 2.37 11.85 2.6 ;
      RECT 11.33 2.4 11.85 2.57 ;
      RECT 11.53 6.26 11.85 6.55 ;
      RECT 11.5 6.29 11.85 6.52 ;
      RECT 11.33 6.32 11.85 6.49 ;
      RECT 8.635 1.895 8.955 2.155 ;
      RECT 8.2 1.91 8.49 2.14 ;
      RECT 8.2 1.955 8.955 2.095 ;
      RECT 8.635 3.575 8.955 3.835 ;
      RECT 8.2 3.59 8.49 3.82 ;
      RECT 8.2 3.635 8.955 3.775 ;
      RECT 7.96 3.03 8.25 3.26 ;
      RECT 7.96 3.075 8.535 3.215 ;
      RECT 8.395 2.935 8.655 3.075 ;
      RECT 8.44 2.75 8.73 2.98 ;
      RECT 6.595 2.935 7.695 3.075 ;
      RECT 6.4 2.735 6.72 2.995 ;
      RECT 7.48 2.75 7.77 2.98 ;
      RECT 6.4 2.75 6.81 2.995 ;
      RECT 6.775 1.895 7.095 2.155 ;
      RECT 7.24 1.91 7.53 2.14 ;
      RECT 6.775 1.955 7.53 2.095 ;
      RECT 4.075 3.16 6.255 3.3 ;
      RECT 6.115 2.17 6.255 3.3 ;
      RECT 4.075 3.075 5.37 3.3 ;
      RECT 5.08 3.03 5.37 3.3 ;
      RECT 4.075 2.795 4.41 3.3 ;
      RECT 4.12 2.75 4.41 3.3 ;
      RECT 7 2.47 7.29 2.7 ;
      RECT 6.115 2.375 7.215 2.515 ;
      RECT 6.04 2.17 6.33 2.42 ;
      RECT 6.26 7.77 6.55 8 ;
      RECT 6.32 7.03 6.49 8 ;
      RECT 6.22 7.06 6.59 7.43 ;
      RECT 6.26 7.03 6.55 7.43 ;
      RECT 6.025 3.575 6.345 3.835 ;
      RECT 6.025 3.59 6.54 3.82 ;
      RECT 4.6 2.47 4.89 2.7 ;
      RECT 4.75 2.075 4.89 2.7 ;
      RECT 4.75 2.075 5.055 2.215 ;
      RECT 5.545 1.895 5.865 2.155 ;
      RECT 4.825 1.895 5.145 2.155 ;
      RECT 5.32 1.91 5.865 2.14 ;
      RECT 4.825 1.955 5.865 2.095 ;
      RECT 4.465 3.575 4.785 3.835 ;
      RECT 4.36 3.59 4.785 3.82 ;
      RECT 2.44 3.03 2.73 3.26 ;
      RECT 2.44 3.03 2.895 3.215 ;
      RECT 2.755 2.555 2.895 3.215 ;
      RECT 2.875 1.955 3.015 2.695 ;
      RECT 3.745 1.895 4.065 2.155 ;
      RECT 2.92 1.91 3.21 2.14 ;
      RECT 2.875 1.955 4.065 2.095 ;
      RECT 3.625 2.455 3.945 2.715 ;
      RECT 3.16 2.47 3.45 2.7 ;
      RECT 3.16 2.515 3.945 2.655 ;
      RECT 3.385 3.015 3.705 3.275 ;
      RECT 3.385 3.03 3.93 3.26 ;
      RECT 2.92 3.59 3.21 3.82 ;
      RECT 2.035 3.47 3.135 3.61 ;
      RECT 1.96 3.31 2.25 3.54 ;
      RECT -1.255 7.77 -0.965 8 ;
      RECT -1.195 7.03 -1.025 8 ;
      RECT -1.285 7.03 -0.935 7.32 ;
      RECT -1.66 6.29 -1.31 6.58 ;
      RECT -1.8 6.32 -1.31 6.49 ;
      RECT 68.985 2.455 69.305 2.715 ;
      RECT 67.815 3.295 68.135 3.555 ;
      RECT 66.585 2.735 66.905 2.995 ;
      RECT 66.105 2.455 66.425 2.715 ;
      RECT 65.25 1.895 65.65 2.155 ;
      RECT 64.905 3.575 65.225 3.835 ;
      RECT 63.225 2.455 63.545 2.715 ;
      RECT 62.745 2.735 63.065 2.995 ;
      RECT 62.055 1.895 62.375 2.155 ;
      RECT 62.055 3.295 62.375 3.555 ;
      RECT 53.725 2.455 54.045 2.715 ;
      RECT 52.555 3.295 52.875 3.555 ;
      RECT 51.325 2.735 51.645 2.995 ;
      RECT 50.845 2.455 51.165 2.715 ;
      RECT 49.99 1.895 50.39 2.155 ;
      RECT 49.645 3.575 49.965 3.835 ;
      RECT 47.965 2.455 48.285 2.715 ;
      RECT 47.485 2.735 47.805 2.995 ;
      RECT 46.795 1.895 47.115 2.155 ;
      RECT 46.795 3.295 47.115 3.555 ;
      RECT 38.465 2.455 38.785 2.715 ;
      RECT 37.295 3.295 37.615 3.555 ;
      RECT 36.065 2.735 36.385 2.995 ;
      RECT 35.585 2.455 35.905 2.715 ;
      RECT 34.73 1.895 35.13 2.155 ;
      RECT 34.385 3.575 34.705 3.835 ;
      RECT 32.705 2.455 33.025 2.715 ;
      RECT 32.225 2.735 32.545 2.995 ;
      RECT 31.535 1.895 31.855 2.155 ;
      RECT 31.535 3.295 31.855 3.555 ;
      RECT 23.205 2.455 23.525 2.715 ;
      RECT 22.035 3.295 22.355 3.555 ;
      RECT 20.805 2.735 21.125 2.995 ;
      RECT 20.325 2.455 20.645 2.715 ;
      RECT 19.47 1.895 19.87 2.155 ;
      RECT 19.125 3.575 19.445 3.835 ;
      RECT 17.445 2.455 17.765 2.715 ;
      RECT 16.965 2.735 17.285 2.995 ;
      RECT 16.275 1.895 16.595 2.155 ;
      RECT 16.275 3.295 16.595 3.555 ;
      RECT 7.945 2.455 8.265 2.715 ;
      RECT 6.775 3.295 7.095 3.555 ;
      RECT 5.545 2.735 5.865 2.995 ;
      RECT 5.065 2.455 5.385 2.715 ;
      RECT 4.21 1.895 4.61 2.155 ;
      RECT 3.865 3.575 4.185 3.835 ;
      RECT 2.185 2.455 2.505 2.715 ;
      RECT 1.705 2.735 2.025 2.995 ;
      RECT 1.015 1.895 1.335 2.155 ;
      RECT 1.015 3.295 1.335 3.555 ;
    LAYER mcon ;
      RECT 75.755 6.325 75.925 6.495 ;
      RECT 75.76 6.32 75.93 6.49 ;
      RECT 60.495 6.325 60.665 6.495 ;
      RECT 60.5 6.32 60.67 6.49 ;
      RECT 45.235 6.325 45.405 6.495 ;
      RECT 45.24 6.32 45.41 6.49 ;
      RECT 29.975 6.325 30.145 6.495 ;
      RECT 29.98 6.32 30.15 6.49 ;
      RECT 14.715 6.325 14.885 6.495 ;
      RECT 14.72 6.32 14.89 6.49 ;
      RECT 75.755 7.805 75.925 7.975 ;
      RECT 75.385 2.765 75.555 2.935 ;
      RECT 75.385 5.955 75.555 6.125 ;
      RECT 74.765 0.915 74.935 1.085 ;
      RECT 74.765 2.395 74.935 2.565 ;
      RECT 74.765 6.325 74.935 6.495 ;
      RECT 74.765 7.805 74.935 7.975 ;
      RECT 74.395 2.765 74.565 2.935 ;
      RECT 74.395 5.955 74.565 6.125 ;
      RECT 73.405 2.03 73.575 2.2 ;
      RECT 73.405 6.69 73.575 6.86 ;
      RECT 72.975 0.92 73.145 1.09 ;
      RECT 72.975 1.66 73.145 1.83 ;
      RECT 72.975 7.06 73.145 7.23 ;
      RECT 72.975 7.8 73.145 7.97 ;
      RECT 72.6 2.4 72.77 2.57 ;
      RECT 72.6 6.32 72.77 6.49 ;
      RECT 69.54 2.78 69.71 2.95 ;
      RECT 69.3 1.94 69.47 2.11 ;
      RECT 69.3 3.62 69.47 3.79 ;
      RECT 69.06 2.5 69.23 2.67 ;
      RECT 69.06 3.06 69.23 3.23 ;
      RECT 68.58 2.78 68.75 2.95 ;
      RECT 68.34 1.94 68.51 2.11 ;
      RECT 68.1 2.5 68.27 2.67 ;
      RECT 67.89 3.34 68.06 3.51 ;
      RECT 67.79 6.69 67.96 6.86 ;
      RECT 67.62 2.78 67.79 2.95 ;
      RECT 67.36 7.06 67.53 7.23 ;
      RECT 67.36 7.8 67.53 7.97 ;
      RECT 67.35 3.62 67.52 3.79 ;
      RECT 67.14 2.2 67.31 2.37 ;
      RECT 66.66 2.78 66.83 2.95 ;
      RECT 66.42 1.94 66.59 2.11 ;
      RECT 66.18 2.5 66.35 2.67 ;
      RECT 66.18 3.06 66.35 3.23 ;
      RECT 65.7 2.5 65.87 2.67 ;
      RECT 65.46 3.62 65.63 3.79 ;
      RECT 65.42 1.94 65.59 2.11 ;
      RECT 65.22 2.78 65.39 2.95 ;
      RECT 64.98 3.62 65.15 3.79 ;
      RECT 64.74 3.06 64.91 3.23 ;
      RECT 64.26 2.5 64.43 2.67 ;
      RECT 64.02 1.94 64.19 2.11 ;
      RECT 64.02 3.62 64.19 3.79 ;
      RECT 63.54 3.06 63.71 3.23 ;
      RECT 63.3 2.5 63.47 2.67 ;
      RECT 63.06 3.34 63.23 3.51 ;
      RECT 62.82 2.78 62.99 2.95 ;
      RECT 62.13 1.94 62.3 2.11 ;
      RECT 62.13 3.34 62.3 3.51 ;
      RECT 60.495 7.805 60.665 7.975 ;
      RECT 60.125 2.765 60.295 2.935 ;
      RECT 60.125 5.955 60.295 6.125 ;
      RECT 59.505 0.915 59.675 1.085 ;
      RECT 59.505 2.395 59.675 2.565 ;
      RECT 59.505 6.325 59.675 6.495 ;
      RECT 59.505 7.805 59.675 7.975 ;
      RECT 59.135 2.765 59.305 2.935 ;
      RECT 59.135 5.955 59.305 6.125 ;
      RECT 58.145 2.03 58.315 2.2 ;
      RECT 58.145 6.69 58.315 6.86 ;
      RECT 57.715 0.92 57.885 1.09 ;
      RECT 57.715 1.66 57.885 1.83 ;
      RECT 57.715 7.06 57.885 7.23 ;
      RECT 57.715 7.8 57.885 7.97 ;
      RECT 57.34 2.4 57.51 2.57 ;
      RECT 57.34 6.32 57.51 6.49 ;
      RECT 54.28 2.78 54.45 2.95 ;
      RECT 54.04 1.94 54.21 2.11 ;
      RECT 54.04 3.62 54.21 3.79 ;
      RECT 53.8 2.5 53.97 2.67 ;
      RECT 53.8 3.06 53.97 3.23 ;
      RECT 53.32 2.78 53.49 2.95 ;
      RECT 53.08 1.94 53.25 2.11 ;
      RECT 52.84 2.5 53.01 2.67 ;
      RECT 52.63 3.34 52.8 3.51 ;
      RECT 52.53 6.69 52.7 6.86 ;
      RECT 52.36 2.78 52.53 2.95 ;
      RECT 52.1 7.06 52.27 7.23 ;
      RECT 52.1 7.8 52.27 7.97 ;
      RECT 52.09 3.62 52.26 3.79 ;
      RECT 51.88 2.2 52.05 2.37 ;
      RECT 51.4 2.78 51.57 2.95 ;
      RECT 51.16 1.94 51.33 2.11 ;
      RECT 50.92 2.5 51.09 2.67 ;
      RECT 50.92 3.06 51.09 3.23 ;
      RECT 50.44 2.5 50.61 2.67 ;
      RECT 50.2 3.62 50.37 3.79 ;
      RECT 50.16 1.94 50.33 2.11 ;
      RECT 49.96 2.78 50.13 2.95 ;
      RECT 49.72 3.62 49.89 3.79 ;
      RECT 49.48 3.06 49.65 3.23 ;
      RECT 49 2.5 49.17 2.67 ;
      RECT 48.76 1.94 48.93 2.11 ;
      RECT 48.76 3.62 48.93 3.79 ;
      RECT 48.28 3.06 48.45 3.23 ;
      RECT 48.04 2.5 48.21 2.67 ;
      RECT 47.8 3.34 47.97 3.51 ;
      RECT 47.56 2.78 47.73 2.95 ;
      RECT 46.87 1.94 47.04 2.11 ;
      RECT 46.87 3.34 47.04 3.51 ;
      RECT 45.235 7.805 45.405 7.975 ;
      RECT 44.865 2.765 45.035 2.935 ;
      RECT 44.865 5.955 45.035 6.125 ;
      RECT 44.245 0.915 44.415 1.085 ;
      RECT 44.245 2.395 44.415 2.565 ;
      RECT 44.245 6.325 44.415 6.495 ;
      RECT 44.245 7.805 44.415 7.975 ;
      RECT 43.875 2.765 44.045 2.935 ;
      RECT 43.875 5.955 44.045 6.125 ;
      RECT 42.885 2.03 43.055 2.2 ;
      RECT 42.885 6.69 43.055 6.86 ;
      RECT 42.455 0.92 42.625 1.09 ;
      RECT 42.455 1.66 42.625 1.83 ;
      RECT 42.455 7.06 42.625 7.23 ;
      RECT 42.455 7.8 42.625 7.97 ;
      RECT 42.08 2.4 42.25 2.57 ;
      RECT 42.08 6.32 42.25 6.49 ;
      RECT 39.02 2.78 39.19 2.95 ;
      RECT 38.78 1.94 38.95 2.11 ;
      RECT 38.78 3.62 38.95 3.79 ;
      RECT 38.54 2.5 38.71 2.67 ;
      RECT 38.54 3.06 38.71 3.23 ;
      RECT 38.06 2.78 38.23 2.95 ;
      RECT 37.82 1.94 37.99 2.11 ;
      RECT 37.58 2.5 37.75 2.67 ;
      RECT 37.37 3.34 37.54 3.51 ;
      RECT 37.27 6.69 37.44 6.86 ;
      RECT 37.1 2.78 37.27 2.95 ;
      RECT 36.84 7.06 37.01 7.23 ;
      RECT 36.84 7.8 37.01 7.97 ;
      RECT 36.83 3.62 37 3.79 ;
      RECT 36.62 2.2 36.79 2.37 ;
      RECT 36.14 2.78 36.31 2.95 ;
      RECT 35.9 1.94 36.07 2.11 ;
      RECT 35.66 2.5 35.83 2.67 ;
      RECT 35.66 3.06 35.83 3.23 ;
      RECT 35.18 2.5 35.35 2.67 ;
      RECT 34.94 3.62 35.11 3.79 ;
      RECT 34.9 1.94 35.07 2.11 ;
      RECT 34.7 2.78 34.87 2.95 ;
      RECT 34.46 3.62 34.63 3.79 ;
      RECT 34.22 3.06 34.39 3.23 ;
      RECT 33.74 2.5 33.91 2.67 ;
      RECT 33.5 1.94 33.67 2.11 ;
      RECT 33.5 3.62 33.67 3.79 ;
      RECT 33.02 3.06 33.19 3.23 ;
      RECT 32.78 2.5 32.95 2.67 ;
      RECT 32.54 3.34 32.71 3.51 ;
      RECT 32.3 2.78 32.47 2.95 ;
      RECT 31.61 1.94 31.78 2.11 ;
      RECT 31.61 3.34 31.78 3.51 ;
      RECT 29.975 7.805 30.145 7.975 ;
      RECT 29.605 2.765 29.775 2.935 ;
      RECT 29.605 5.955 29.775 6.125 ;
      RECT 28.985 0.915 29.155 1.085 ;
      RECT 28.985 2.395 29.155 2.565 ;
      RECT 28.985 6.325 29.155 6.495 ;
      RECT 28.985 7.805 29.155 7.975 ;
      RECT 28.615 2.765 28.785 2.935 ;
      RECT 28.615 5.955 28.785 6.125 ;
      RECT 27.625 2.03 27.795 2.2 ;
      RECT 27.625 6.69 27.795 6.86 ;
      RECT 27.195 0.92 27.365 1.09 ;
      RECT 27.195 1.66 27.365 1.83 ;
      RECT 27.195 7.06 27.365 7.23 ;
      RECT 27.195 7.8 27.365 7.97 ;
      RECT 26.82 2.4 26.99 2.57 ;
      RECT 26.82 6.32 26.99 6.49 ;
      RECT 23.76 2.78 23.93 2.95 ;
      RECT 23.52 1.94 23.69 2.11 ;
      RECT 23.52 3.62 23.69 3.79 ;
      RECT 23.28 2.5 23.45 2.67 ;
      RECT 23.28 3.06 23.45 3.23 ;
      RECT 22.8 2.78 22.97 2.95 ;
      RECT 22.56 1.94 22.73 2.11 ;
      RECT 22.32 2.5 22.49 2.67 ;
      RECT 22.11 3.34 22.28 3.51 ;
      RECT 22.01 6.69 22.18 6.86 ;
      RECT 21.84 2.78 22.01 2.95 ;
      RECT 21.58 7.06 21.75 7.23 ;
      RECT 21.58 7.8 21.75 7.97 ;
      RECT 21.57 3.62 21.74 3.79 ;
      RECT 21.36 2.2 21.53 2.37 ;
      RECT 20.88 2.78 21.05 2.95 ;
      RECT 20.64 1.94 20.81 2.11 ;
      RECT 20.4 2.5 20.57 2.67 ;
      RECT 20.4 3.06 20.57 3.23 ;
      RECT 19.92 2.5 20.09 2.67 ;
      RECT 19.68 3.62 19.85 3.79 ;
      RECT 19.64 1.94 19.81 2.11 ;
      RECT 19.44 2.78 19.61 2.95 ;
      RECT 19.2 3.62 19.37 3.79 ;
      RECT 18.96 3.06 19.13 3.23 ;
      RECT 18.48 2.5 18.65 2.67 ;
      RECT 18.24 1.94 18.41 2.11 ;
      RECT 18.24 3.62 18.41 3.79 ;
      RECT 17.76 3.06 17.93 3.23 ;
      RECT 17.52 2.5 17.69 2.67 ;
      RECT 17.28 3.34 17.45 3.51 ;
      RECT 17.04 2.78 17.21 2.95 ;
      RECT 16.35 1.94 16.52 2.11 ;
      RECT 16.35 3.34 16.52 3.51 ;
      RECT 14.715 7.805 14.885 7.975 ;
      RECT 14.345 2.765 14.515 2.935 ;
      RECT 14.345 5.955 14.515 6.125 ;
      RECT 13.725 0.915 13.895 1.085 ;
      RECT 13.725 2.395 13.895 2.565 ;
      RECT 13.725 6.325 13.895 6.495 ;
      RECT 13.725 7.805 13.895 7.975 ;
      RECT 13.355 2.765 13.525 2.935 ;
      RECT 13.355 5.955 13.525 6.125 ;
      RECT 12.365 2.03 12.535 2.2 ;
      RECT 12.365 6.69 12.535 6.86 ;
      RECT 11.935 0.92 12.105 1.09 ;
      RECT 11.935 1.66 12.105 1.83 ;
      RECT 11.935 7.06 12.105 7.23 ;
      RECT 11.935 7.8 12.105 7.97 ;
      RECT 11.56 2.4 11.73 2.57 ;
      RECT 11.56 6.32 11.73 6.49 ;
      RECT 8.5 2.78 8.67 2.95 ;
      RECT 8.26 1.94 8.43 2.11 ;
      RECT 8.26 3.62 8.43 3.79 ;
      RECT 8.02 2.5 8.19 2.67 ;
      RECT 8.02 3.06 8.19 3.23 ;
      RECT 7.54 2.78 7.71 2.95 ;
      RECT 7.3 1.94 7.47 2.11 ;
      RECT 7.06 2.5 7.23 2.67 ;
      RECT 6.85 3.34 7.02 3.51 ;
      RECT 6.75 6.69 6.92 6.86 ;
      RECT 6.58 2.78 6.75 2.95 ;
      RECT 6.32 7.06 6.49 7.23 ;
      RECT 6.32 7.8 6.49 7.97 ;
      RECT 6.31 3.62 6.48 3.79 ;
      RECT 6.1 2.2 6.27 2.37 ;
      RECT 5.62 2.78 5.79 2.95 ;
      RECT 5.38 1.94 5.55 2.11 ;
      RECT 5.14 2.5 5.31 2.67 ;
      RECT 5.14 3.06 5.31 3.23 ;
      RECT 4.66 2.5 4.83 2.67 ;
      RECT 4.42 3.62 4.59 3.79 ;
      RECT 4.38 1.94 4.55 2.11 ;
      RECT 4.18 2.78 4.35 2.95 ;
      RECT 3.94 3.62 4.11 3.79 ;
      RECT 3.7 3.06 3.87 3.23 ;
      RECT 3.22 2.5 3.39 2.67 ;
      RECT 2.98 1.94 3.15 2.11 ;
      RECT 2.98 3.62 3.15 3.79 ;
      RECT 2.5 3.06 2.67 3.23 ;
      RECT 2.26 2.5 2.43 2.67 ;
      RECT 2.02 3.34 2.19 3.51 ;
      RECT 1.78 2.78 1.95 2.95 ;
      RECT 1.09 1.94 1.26 2.11 ;
      RECT 1.09 3.34 1.26 3.51 ;
      RECT -1.195 7.06 -1.025 7.23 ;
      RECT -1.195 7.8 -1.025 7.97 ;
      RECT -1.57 6.32 -1.4 6.49 ;
    LAYER li1 ;
      RECT 75.755 5.025 75.925 6.495 ;
      RECT 75.755 6.32 75.93 6.49 ;
      RECT 75.385 1.745 75.555 2.935 ;
      RECT 75.385 1.745 75.855 1.915 ;
      RECT 75.385 6.975 75.855 7.145 ;
      RECT 75.385 5.955 75.555 7.145 ;
      RECT 74.395 1.745 74.565 2.935 ;
      RECT 74.395 1.745 74.865 1.915 ;
      RECT 74.395 6.975 74.865 7.145 ;
      RECT 74.395 5.955 74.565 7.145 ;
      RECT 72.545 2.64 72.715 3.87 ;
      RECT 72.6 0.86 72.77 2.81 ;
      RECT 72.545 0.58 72.715 1.03 ;
      RECT 72.545 7.86 72.715 8.31 ;
      RECT 72.6 6.08 72.77 8.03 ;
      RECT 72.545 5.02 72.715 6.25 ;
      RECT 72.025 0.58 72.195 3.87 ;
      RECT 72.025 2.08 72.43 2.41 ;
      RECT 72.025 1.24 72.43 1.57 ;
      RECT 72.025 5.02 72.195 8.31 ;
      RECT 72.025 7.32 72.43 7.65 ;
      RECT 72.025 6.48 72.43 6.81 ;
      RECT 69.3 3.62 69.815 3.79 ;
      RECT 69.645 3.23 69.815 3.79 ;
      RECT 69.75 3.15 69.92 3.48 ;
      RECT 69.54 2.54 69.815 2.95 ;
      RECT 69.42 2.54 69.815 2.75 ;
      RECT 67.89 3.15 68.06 3.51 ;
      RECT 67.89 3.23 69.23 3.4 ;
      RECT 69.06 3.06 69.23 3.4 ;
      RECT 67.62 2.58 67.79 2.95 ;
      RECT 67.14 2.58 67.79 2.85 ;
      RECT 67.06 2.58 67.87 2.75 ;
      RECT 66.42 1.82 66.59 2.11 ;
      RECT 66.42 1.82 67.66 1.99 ;
      RECT 67.14 2.16 67.31 2.37 ;
      RECT 66.78 2.16 67.31 2.33 ;
      RECT 66.41 5.02 66.58 8.31 ;
      RECT 66.41 7.32 66.815 7.65 ;
      RECT 66.41 6.48 66.815 6.81 ;
      RECT 66.18 3.23 66.67 3.4 ;
      RECT 66.18 3.06 66.35 3.4 ;
      RECT 65.46 3.23 65.63 3.79 ;
      RECT 65.35 3.23 65.68 3.4 ;
      RECT 65.42 1.84 65.59 2.11 ;
      RECT 65.46 1.76 65.63 2.09 ;
      RECT 65.325 1.84 65.63 2.06 ;
      RECT 63.9 3.23 64.19 3.79 ;
      RECT 64.02 3.15 64.19 3.79 ;
      RECT 60.495 5.025 60.665 6.495 ;
      RECT 60.495 6.32 60.67 6.49 ;
      RECT 60.125 1.745 60.295 2.935 ;
      RECT 60.125 1.745 60.595 1.915 ;
      RECT 60.125 6.975 60.595 7.145 ;
      RECT 60.125 5.955 60.295 7.145 ;
      RECT 59.135 1.745 59.305 2.935 ;
      RECT 59.135 1.745 59.605 1.915 ;
      RECT 59.135 6.975 59.605 7.145 ;
      RECT 59.135 5.955 59.305 7.145 ;
      RECT 57.285 2.64 57.455 3.87 ;
      RECT 57.34 0.86 57.51 2.81 ;
      RECT 57.285 0.58 57.455 1.03 ;
      RECT 57.285 7.86 57.455 8.31 ;
      RECT 57.34 6.08 57.51 8.03 ;
      RECT 57.285 5.02 57.455 6.25 ;
      RECT 56.765 0.58 56.935 3.87 ;
      RECT 56.765 2.08 57.17 2.41 ;
      RECT 56.765 1.24 57.17 1.57 ;
      RECT 56.765 5.02 56.935 8.31 ;
      RECT 56.765 7.32 57.17 7.65 ;
      RECT 56.765 6.48 57.17 6.81 ;
      RECT 54.04 3.62 54.555 3.79 ;
      RECT 54.385 3.23 54.555 3.79 ;
      RECT 54.49 3.15 54.66 3.48 ;
      RECT 54.28 2.54 54.555 2.95 ;
      RECT 54.16 2.54 54.555 2.75 ;
      RECT 52.63 3.15 52.8 3.51 ;
      RECT 52.63 3.23 53.97 3.4 ;
      RECT 53.8 3.06 53.97 3.4 ;
      RECT 52.36 2.58 52.53 2.95 ;
      RECT 51.88 2.58 52.53 2.85 ;
      RECT 51.8 2.58 52.61 2.75 ;
      RECT 51.16 1.82 51.33 2.11 ;
      RECT 51.16 1.82 52.4 1.99 ;
      RECT 51.88 2.16 52.05 2.37 ;
      RECT 51.52 2.16 52.05 2.33 ;
      RECT 51.15 5.02 51.32 8.31 ;
      RECT 51.15 7.32 51.555 7.65 ;
      RECT 51.15 6.48 51.555 6.81 ;
      RECT 50.92 3.23 51.41 3.4 ;
      RECT 50.92 3.06 51.09 3.4 ;
      RECT 50.2 3.23 50.37 3.79 ;
      RECT 50.09 3.23 50.42 3.4 ;
      RECT 50.16 1.84 50.33 2.11 ;
      RECT 50.2 1.76 50.37 2.09 ;
      RECT 50.065 1.84 50.37 2.06 ;
      RECT 48.64 3.23 48.93 3.79 ;
      RECT 48.76 3.15 48.93 3.79 ;
      RECT 45.235 5.025 45.405 6.495 ;
      RECT 45.235 6.32 45.41 6.49 ;
      RECT 44.865 1.745 45.035 2.935 ;
      RECT 44.865 1.745 45.335 1.915 ;
      RECT 44.865 6.975 45.335 7.145 ;
      RECT 44.865 5.955 45.035 7.145 ;
      RECT 43.875 1.745 44.045 2.935 ;
      RECT 43.875 1.745 44.345 1.915 ;
      RECT 43.875 6.975 44.345 7.145 ;
      RECT 43.875 5.955 44.045 7.145 ;
      RECT 42.025 2.64 42.195 3.87 ;
      RECT 42.08 0.86 42.25 2.81 ;
      RECT 42.025 0.58 42.195 1.03 ;
      RECT 42.025 7.86 42.195 8.31 ;
      RECT 42.08 6.08 42.25 8.03 ;
      RECT 42.025 5.02 42.195 6.25 ;
      RECT 41.505 0.58 41.675 3.87 ;
      RECT 41.505 2.08 41.91 2.41 ;
      RECT 41.505 1.24 41.91 1.57 ;
      RECT 41.505 5.02 41.675 8.31 ;
      RECT 41.505 7.32 41.91 7.65 ;
      RECT 41.505 6.48 41.91 6.81 ;
      RECT 38.78 3.62 39.295 3.79 ;
      RECT 39.125 3.23 39.295 3.79 ;
      RECT 39.23 3.15 39.4 3.48 ;
      RECT 39.02 2.54 39.295 2.95 ;
      RECT 38.9 2.54 39.295 2.75 ;
      RECT 37.37 3.15 37.54 3.51 ;
      RECT 37.37 3.23 38.71 3.4 ;
      RECT 38.54 3.06 38.71 3.4 ;
      RECT 37.1 2.58 37.27 2.95 ;
      RECT 36.62 2.58 37.27 2.85 ;
      RECT 36.54 2.58 37.35 2.75 ;
      RECT 35.9 1.82 36.07 2.11 ;
      RECT 35.9 1.82 37.14 1.99 ;
      RECT 36.62 2.16 36.79 2.37 ;
      RECT 36.26 2.16 36.79 2.33 ;
      RECT 35.89 5.02 36.06 8.31 ;
      RECT 35.89 7.32 36.295 7.65 ;
      RECT 35.89 6.48 36.295 6.81 ;
      RECT 35.66 3.23 36.15 3.4 ;
      RECT 35.66 3.06 35.83 3.4 ;
      RECT 34.94 3.23 35.11 3.79 ;
      RECT 34.83 3.23 35.16 3.4 ;
      RECT 34.9 1.84 35.07 2.11 ;
      RECT 34.94 1.76 35.11 2.09 ;
      RECT 34.805 1.84 35.11 2.06 ;
      RECT 33.38 3.23 33.67 3.79 ;
      RECT 33.5 3.15 33.67 3.79 ;
      RECT 29.975 5.025 30.145 6.495 ;
      RECT 29.975 6.32 30.15 6.49 ;
      RECT 29.605 1.745 29.775 2.935 ;
      RECT 29.605 1.745 30.075 1.915 ;
      RECT 29.605 6.975 30.075 7.145 ;
      RECT 29.605 5.955 29.775 7.145 ;
      RECT 28.615 1.745 28.785 2.935 ;
      RECT 28.615 1.745 29.085 1.915 ;
      RECT 28.615 6.975 29.085 7.145 ;
      RECT 28.615 5.955 28.785 7.145 ;
      RECT 26.765 2.64 26.935 3.87 ;
      RECT 26.82 0.86 26.99 2.81 ;
      RECT 26.765 0.58 26.935 1.03 ;
      RECT 26.765 7.86 26.935 8.31 ;
      RECT 26.82 6.08 26.99 8.03 ;
      RECT 26.765 5.02 26.935 6.25 ;
      RECT 26.245 0.58 26.415 3.87 ;
      RECT 26.245 2.08 26.65 2.41 ;
      RECT 26.245 1.24 26.65 1.57 ;
      RECT 26.245 5.02 26.415 8.31 ;
      RECT 26.245 7.32 26.65 7.65 ;
      RECT 26.245 6.48 26.65 6.81 ;
      RECT 23.52 3.62 24.035 3.79 ;
      RECT 23.865 3.23 24.035 3.79 ;
      RECT 23.97 3.15 24.14 3.48 ;
      RECT 23.76 2.54 24.035 2.95 ;
      RECT 23.64 2.54 24.035 2.75 ;
      RECT 22.11 3.15 22.28 3.51 ;
      RECT 22.11 3.23 23.45 3.4 ;
      RECT 23.28 3.06 23.45 3.4 ;
      RECT 21.84 2.58 22.01 2.95 ;
      RECT 21.36 2.58 22.01 2.85 ;
      RECT 21.28 2.58 22.09 2.75 ;
      RECT 20.64 1.82 20.81 2.11 ;
      RECT 20.64 1.82 21.88 1.99 ;
      RECT 21.36 2.16 21.53 2.37 ;
      RECT 21 2.16 21.53 2.33 ;
      RECT 20.63 5.02 20.8 8.31 ;
      RECT 20.63 7.32 21.035 7.65 ;
      RECT 20.63 6.48 21.035 6.81 ;
      RECT 20.4 3.23 20.89 3.4 ;
      RECT 20.4 3.06 20.57 3.4 ;
      RECT 19.68 3.23 19.85 3.79 ;
      RECT 19.57 3.23 19.9 3.4 ;
      RECT 19.64 1.84 19.81 2.11 ;
      RECT 19.68 1.76 19.85 2.09 ;
      RECT 19.545 1.84 19.85 2.06 ;
      RECT 18.12 3.23 18.41 3.79 ;
      RECT 18.24 3.15 18.41 3.79 ;
      RECT 14.715 5.025 14.885 6.495 ;
      RECT 14.715 6.32 14.89 6.49 ;
      RECT 14.345 1.745 14.515 2.935 ;
      RECT 14.345 1.745 14.815 1.915 ;
      RECT 14.345 6.975 14.815 7.145 ;
      RECT 14.345 5.955 14.515 7.145 ;
      RECT 13.355 1.745 13.525 2.935 ;
      RECT 13.355 1.745 13.825 1.915 ;
      RECT 13.355 6.975 13.825 7.145 ;
      RECT 13.355 5.955 13.525 7.145 ;
      RECT 11.505 2.64 11.675 3.87 ;
      RECT 11.56 0.86 11.73 2.81 ;
      RECT 11.505 0.58 11.675 1.03 ;
      RECT 11.505 7.86 11.675 8.31 ;
      RECT 11.56 6.08 11.73 8.03 ;
      RECT 11.505 5.02 11.675 6.25 ;
      RECT 10.985 0.58 11.155 3.87 ;
      RECT 10.985 2.08 11.39 2.41 ;
      RECT 10.985 1.24 11.39 1.57 ;
      RECT 10.985 5.02 11.155 8.31 ;
      RECT 10.985 7.32 11.39 7.65 ;
      RECT 10.985 6.48 11.39 6.81 ;
      RECT 8.26 3.62 8.775 3.79 ;
      RECT 8.605 3.23 8.775 3.79 ;
      RECT 8.71 3.15 8.88 3.48 ;
      RECT 8.5 2.54 8.775 2.95 ;
      RECT 8.38 2.54 8.775 2.75 ;
      RECT 6.85 3.15 7.02 3.51 ;
      RECT 6.85 3.23 8.19 3.4 ;
      RECT 8.02 3.06 8.19 3.4 ;
      RECT 6.58 2.58 6.75 2.95 ;
      RECT 6.1 2.58 6.75 2.85 ;
      RECT 6.02 2.58 6.83 2.75 ;
      RECT 5.38 1.82 5.55 2.11 ;
      RECT 5.38 1.82 6.62 1.99 ;
      RECT 6.1 2.16 6.27 2.37 ;
      RECT 5.74 2.16 6.27 2.33 ;
      RECT 5.37 5.02 5.54 8.31 ;
      RECT 5.37 7.32 5.775 7.65 ;
      RECT 5.37 6.48 5.775 6.81 ;
      RECT 5.14 3.23 5.63 3.4 ;
      RECT 5.14 3.06 5.31 3.4 ;
      RECT 4.42 3.23 4.59 3.79 ;
      RECT 4.31 3.23 4.64 3.4 ;
      RECT 4.38 1.84 4.55 2.11 ;
      RECT 4.42 1.76 4.59 2.09 ;
      RECT 4.285 1.84 4.59 2.06 ;
      RECT 2.86 3.23 3.15 3.79 ;
      RECT 2.98 3.15 3.15 3.79 ;
      RECT -1.625 7.86 -1.455 8.31 ;
      RECT -1.57 6.08 -1.4 8.03 ;
      RECT -1.625 5.02 -1.455 6.25 ;
      RECT -2.145 5.02 -1.975 8.31 ;
      RECT -2.145 7.32 -1.74 7.65 ;
      RECT -2.145 6.48 -1.74 6.81 ;
      RECT 75.755 7.805 75.925 8.315 ;
      RECT 74.765 0.575 74.935 1.085 ;
      RECT 74.765 2.395 74.935 3.865 ;
      RECT 74.765 5.025 74.935 6.495 ;
      RECT 74.765 7.805 74.935 8.315 ;
      RECT 73.405 0.58 73.575 3.87 ;
      RECT 73.405 5.02 73.575 8.31 ;
      RECT 72.975 0.58 73.145 1.09 ;
      RECT 72.975 1.66 73.145 3.87 ;
      RECT 72.975 5.02 73.145 7.23 ;
      RECT 72.975 7.8 73.145 8.31 ;
      RECT 69.3 1.76 69.47 2.11 ;
      RECT 69.06 2.5 69.23 2.83 ;
      RECT 68.58 2.5 68.75 2.95 ;
      RECT 68.34 1.76 68.51 2.11 ;
      RECT 68.1 2.5 68.27 2.83 ;
      RECT 67.79 5.02 67.96 8.31 ;
      RECT 67.36 5.02 67.53 7.23 ;
      RECT 67.36 7.8 67.53 8.31 ;
      RECT 67.35 3.49 67.52 3.82 ;
      RECT 66.66 2.5 66.83 2.95 ;
      RECT 66.18 2.5 66.35 2.83 ;
      RECT 65.7 2.5 65.87 2.83 ;
      RECT 65.22 2.5 65.39 2.95 ;
      RECT 64.98 3.49 65.15 3.82 ;
      RECT 64.74 2.5 64.91 3.23 ;
      RECT 64.26 2.5 64.43 2.83 ;
      RECT 64.02 1.76 64.19 2.11 ;
      RECT 63.54 3.06 63.71 3.48 ;
      RECT 63.3 2.5 63.47 2.83 ;
      RECT 63.06 3.15 63.23 3.51 ;
      RECT 62.82 2.5 62.99 2.95 ;
      RECT 62.13 1.76 62.3 2.11 ;
      RECT 62.13 3.15 62.3 3.51 ;
      RECT 60.495 7.805 60.665 8.315 ;
      RECT 59.505 0.575 59.675 1.085 ;
      RECT 59.505 2.395 59.675 3.865 ;
      RECT 59.505 5.025 59.675 6.495 ;
      RECT 59.505 7.805 59.675 8.315 ;
      RECT 58.145 0.58 58.315 3.87 ;
      RECT 58.145 5.02 58.315 8.31 ;
      RECT 57.715 0.58 57.885 1.09 ;
      RECT 57.715 1.66 57.885 3.87 ;
      RECT 57.715 5.02 57.885 7.23 ;
      RECT 57.715 7.8 57.885 8.31 ;
      RECT 54.04 1.76 54.21 2.11 ;
      RECT 53.8 2.5 53.97 2.83 ;
      RECT 53.32 2.5 53.49 2.95 ;
      RECT 53.08 1.76 53.25 2.11 ;
      RECT 52.84 2.5 53.01 2.83 ;
      RECT 52.53 5.02 52.7 8.31 ;
      RECT 52.1 5.02 52.27 7.23 ;
      RECT 52.1 7.8 52.27 8.31 ;
      RECT 52.09 3.49 52.26 3.82 ;
      RECT 51.4 2.5 51.57 2.95 ;
      RECT 50.92 2.5 51.09 2.83 ;
      RECT 50.44 2.5 50.61 2.83 ;
      RECT 49.96 2.5 50.13 2.95 ;
      RECT 49.72 3.49 49.89 3.82 ;
      RECT 49.48 2.5 49.65 3.23 ;
      RECT 49 2.5 49.17 2.83 ;
      RECT 48.76 1.76 48.93 2.11 ;
      RECT 48.28 3.06 48.45 3.48 ;
      RECT 48.04 2.5 48.21 2.83 ;
      RECT 47.8 3.15 47.97 3.51 ;
      RECT 47.56 2.5 47.73 2.95 ;
      RECT 46.87 1.76 47.04 2.11 ;
      RECT 46.87 3.15 47.04 3.51 ;
      RECT 45.235 7.805 45.405 8.315 ;
      RECT 44.245 0.575 44.415 1.085 ;
      RECT 44.245 2.395 44.415 3.865 ;
      RECT 44.245 5.025 44.415 6.495 ;
      RECT 44.245 7.805 44.415 8.315 ;
      RECT 42.885 0.58 43.055 3.87 ;
      RECT 42.885 5.02 43.055 8.31 ;
      RECT 42.455 0.58 42.625 1.09 ;
      RECT 42.455 1.66 42.625 3.87 ;
      RECT 42.455 5.02 42.625 7.23 ;
      RECT 42.455 7.8 42.625 8.31 ;
      RECT 38.78 1.76 38.95 2.11 ;
      RECT 38.54 2.5 38.71 2.83 ;
      RECT 38.06 2.5 38.23 2.95 ;
      RECT 37.82 1.76 37.99 2.11 ;
      RECT 37.58 2.5 37.75 2.83 ;
      RECT 37.27 5.02 37.44 8.31 ;
      RECT 36.84 5.02 37.01 7.23 ;
      RECT 36.84 7.8 37.01 8.31 ;
      RECT 36.83 3.49 37 3.82 ;
      RECT 36.14 2.5 36.31 2.95 ;
      RECT 35.66 2.5 35.83 2.83 ;
      RECT 35.18 2.5 35.35 2.83 ;
      RECT 34.7 2.5 34.87 2.95 ;
      RECT 34.46 3.49 34.63 3.82 ;
      RECT 34.22 2.5 34.39 3.23 ;
      RECT 33.74 2.5 33.91 2.83 ;
      RECT 33.5 1.76 33.67 2.11 ;
      RECT 33.02 3.06 33.19 3.48 ;
      RECT 32.78 2.5 32.95 2.83 ;
      RECT 32.54 3.15 32.71 3.51 ;
      RECT 32.3 2.5 32.47 2.95 ;
      RECT 31.61 1.76 31.78 2.11 ;
      RECT 31.61 3.15 31.78 3.51 ;
      RECT 29.975 7.805 30.145 8.315 ;
      RECT 28.985 0.575 29.155 1.085 ;
      RECT 28.985 2.395 29.155 3.865 ;
      RECT 28.985 5.025 29.155 6.495 ;
      RECT 28.985 7.805 29.155 8.315 ;
      RECT 27.625 0.58 27.795 3.87 ;
      RECT 27.625 5.02 27.795 8.31 ;
      RECT 27.195 0.58 27.365 1.09 ;
      RECT 27.195 1.66 27.365 3.87 ;
      RECT 27.195 5.02 27.365 7.23 ;
      RECT 27.195 7.8 27.365 8.31 ;
      RECT 23.52 1.76 23.69 2.11 ;
      RECT 23.28 2.5 23.45 2.83 ;
      RECT 22.8 2.5 22.97 2.95 ;
      RECT 22.56 1.76 22.73 2.11 ;
      RECT 22.32 2.5 22.49 2.83 ;
      RECT 22.01 5.02 22.18 8.31 ;
      RECT 21.58 5.02 21.75 7.23 ;
      RECT 21.58 7.8 21.75 8.31 ;
      RECT 21.57 3.49 21.74 3.82 ;
      RECT 20.88 2.5 21.05 2.95 ;
      RECT 20.4 2.5 20.57 2.83 ;
      RECT 19.92 2.5 20.09 2.83 ;
      RECT 19.44 2.5 19.61 2.95 ;
      RECT 19.2 3.49 19.37 3.82 ;
      RECT 18.96 2.5 19.13 3.23 ;
      RECT 18.48 2.5 18.65 2.83 ;
      RECT 18.24 1.76 18.41 2.11 ;
      RECT 17.76 3.06 17.93 3.48 ;
      RECT 17.52 2.5 17.69 2.83 ;
      RECT 17.28 3.15 17.45 3.51 ;
      RECT 17.04 2.5 17.21 2.95 ;
      RECT 16.35 1.76 16.52 2.11 ;
      RECT 16.35 3.15 16.52 3.51 ;
      RECT 14.715 7.805 14.885 8.315 ;
      RECT 13.725 0.575 13.895 1.085 ;
      RECT 13.725 2.395 13.895 3.865 ;
      RECT 13.725 5.025 13.895 6.495 ;
      RECT 13.725 7.805 13.895 8.315 ;
      RECT 12.365 0.58 12.535 3.87 ;
      RECT 12.365 5.02 12.535 8.31 ;
      RECT 11.935 0.58 12.105 1.09 ;
      RECT 11.935 1.66 12.105 3.87 ;
      RECT 11.935 5.02 12.105 7.23 ;
      RECT 11.935 7.8 12.105 8.31 ;
      RECT 8.26 1.76 8.43 2.11 ;
      RECT 8.02 2.5 8.19 2.83 ;
      RECT 7.54 2.5 7.71 2.95 ;
      RECT 7.3 1.76 7.47 2.11 ;
      RECT 7.06 2.5 7.23 2.83 ;
      RECT 6.75 5.02 6.92 8.31 ;
      RECT 6.32 5.02 6.49 7.23 ;
      RECT 6.32 7.8 6.49 8.31 ;
      RECT 6.31 3.49 6.48 3.82 ;
      RECT 5.62 2.5 5.79 2.95 ;
      RECT 5.14 2.5 5.31 2.83 ;
      RECT 4.66 2.5 4.83 2.83 ;
      RECT 4.18 2.5 4.35 2.95 ;
      RECT 3.94 3.49 4.11 3.82 ;
      RECT 3.7 2.5 3.87 3.23 ;
      RECT 3.22 2.5 3.39 2.83 ;
      RECT 2.98 1.76 3.15 2.11 ;
      RECT 2.5 3.06 2.67 3.48 ;
      RECT 2.26 2.5 2.43 2.83 ;
      RECT 2.02 3.15 2.19 3.51 ;
      RECT 1.78 2.5 1.95 2.95 ;
      RECT 1.09 1.76 1.26 2.11 ;
      RECT 1.09 3.15 1.26 3.51 ;
      RECT -1.195 5.02 -1.025 7.23 ;
      RECT -1.195 7.8 -1.025 8.31 ;
  END
END sky130_osu_ring_oscillator_mpr2xa_8_b0r2

MACRO sky130_osu_ring_oscillator_mpr2ya_8_b0r1
  CLASS BLOCK ;
  ORIGIN -1.495 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ya_8_b0r1 ;
  SIZE 79.095 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 19.01 0.915 19.18 1.085 ;
        RECT 19.005 0.91 19.175 1.08 ;
        RECT 19.005 2.39 19.175 2.56 ;
      LAYER li1 ;
        RECT 19.01 0.915 19.18 1.085 ;
        RECT 19.005 0.57 19.175 1.08 ;
        RECT 19.005 2.39 19.175 3.86 ;
      LAYER met1 ;
        RECT 18.945 2.36 19.235 2.59 ;
        RECT 18.945 0.88 19.235 1.11 ;
        RECT 19.005 0.88 19.175 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 34.27 0.915 34.44 1.085 ;
        RECT 34.265 0.91 34.435 1.08 ;
        RECT 34.265 2.39 34.435 2.56 ;
      LAYER li1 ;
        RECT 34.27 0.915 34.44 1.085 ;
        RECT 34.265 0.57 34.435 1.08 ;
        RECT 34.265 2.39 34.435 3.86 ;
      LAYER met1 ;
        RECT 34.205 2.36 34.495 2.59 ;
        RECT 34.205 0.88 34.495 1.11 ;
        RECT 34.265 0.88 34.435 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 49.53 0.915 49.7 1.085 ;
        RECT 49.525 0.91 49.695 1.08 ;
        RECT 49.525 2.39 49.695 2.56 ;
      LAYER li1 ;
        RECT 49.53 0.915 49.7 1.085 ;
        RECT 49.525 0.57 49.695 1.08 ;
        RECT 49.525 2.39 49.695 3.86 ;
      LAYER met1 ;
        RECT 49.465 2.36 49.755 2.59 ;
        RECT 49.465 0.88 49.755 1.11 ;
        RECT 49.525 0.88 49.695 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 64.79 0.915 64.96 1.085 ;
        RECT 64.785 0.91 64.955 1.08 ;
        RECT 64.785 2.39 64.955 2.56 ;
      LAYER li1 ;
        RECT 64.79 0.915 64.96 1.085 ;
        RECT 64.785 0.57 64.955 1.08 ;
        RECT 64.785 2.39 64.955 3.86 ;
      LAYER met1 ;
        RECT 64.725 2.36 65.015 2.59 ;
        RECT 64.725 0.88 65.015 1.11 ;
        RECT 64.785 0.88 64.955 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 80.05 0.915 80.22 1.085 ;
        RECT 80.045 0.91 80.215 1.08 ;
        RECT 80.045 2.39 80.215 2.56 ;
      LAYER li1 ;
        RECT 80.05 0.915 80.22 1.085 ;
        RECT 80.045 0.57 80.215 1.08 ;
        RECT 80.045 2.39 80.215 3.86 ;
      LAYER met1 ;
        RECT 79.985 2.36 80.275 2.59 ;
        RECT 79.985 0.88 80.275 1.11 ;
        RECT 80.045 0.88 80.215 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 14.775 2.705 15.115 3.055 ;
        RECT 14.77 5.86 15.11 6.21 ;
        RECT 14.85 2.705 15.025 6.21 ;
      LAYER li1 ;
        RECT 14.855 1.66 15.025 2.935 ;
        RECT 14.855 5.945 15.025 7.22 ;
        RECT 9.22 5.945 9.39 7.22 ;
      LAYER met1 ;
        RECT 14.775 2.765 15.255 2.935 ;
        RECT 14.775 2.705 15.115 3.055 ;
        RECT 9.16 5.945 15.255 6.115 ;
        RECT 14.77 5.86 15.11 6.21 ;
        RECT 9.16 5.915 9.45 6.145 ;
      LAYER via1 ;
        RECT 14.87 5.96 15.02 6.11 ;
        RECT 14.875 2.805 15.025 2.955 ;
      LAYER mcon ;
        RECT 9.22 5.945 9.39 6.115 ;
        RECT 14.855 5.945 15.025 6.115 ;
        RECT 14.855 2.765 15.025 2.935 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 30.035 2.705 30.375 3.055 ;
        RECT 30.03 5.86 30.37 6.21 ;
        RECT 30.11 2.705 30.285 6.21 ;
      LAYER li1 ;
        RECT 30.115 1.66 30.285 2.935 ;
        RECT 30.115 5.945 30.285 7.22 ;
        RECT 24.48 5.945 24.65 7.22 ;
      LAYER met1 ;
        RECT 30.035 2.765 30.515 2.935 ;
        RECT 30.035 2.705 30.375 3.055 ;
        RECT 24.42 5.945 30.515 6.115 ;
        RECT 30.03 5.86 30.37 6.21 ;
        RECT 24.42 5.915 24.71 6.145 ;
      LAYER via1 ;
        RECT 30.13 5.96 30.28 6.11 ;
        RECT 30.135 2.805 30.285 2.955 ;
      LAYER mcon ;
        RECT 24.48 5.945 24.65 6.115 ;
        RECT 30.115 5.945 30.285 6.115 ;
        RECT 30.115 2.765 30.285 2.935 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 45.295 2.705 45.635 3.055 ;
        RECT 45.29 5.86 45.63 6.21 ;
        RECT 45.37 2.705 45.545 6.21 ;
      LAYER li1 ;
        RECT 45.375 1.66 45.545 2.935 ;
        RECT 45.375 5.945 45.545 7.22 ;
        RECT 39.74 5.945 39.91 7.22 ;
      LAYER met1 ;
        RECT 45.295 2.765 45.775 2.935 ;
        RECT 45.295 2.705 45.635 3.055 ;
        RECT 39.68 5.945 45.775 6.115 ;
        RECT 45.29 5.86 45.63 6.21 ;
        RECT 39.68 5.915 39.97 6.145 ;
      LAYER via1 ;
        RECT 45.39 5.96 45.54 6.11 ;
        RECT 45.395 2.805 45.545 2.955 ;
      LAYER mcon ;
        RECT 39.74 5.945 39.91 6.115 ;
        RECT 45.375 5.945 45.545 6.115 ;
        RECT 45.375 2.765 45.545 2.935 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 60.555 2.705 60.895 3.055 ;
        RECT 60.55 5.86 60.89 6.21 ;
        RECT 60.63 2.705 60.805 6.21 ;
      LAYER li1 ;
        RECT 60.635 1.66 60.805 2.935 ;
        RECT 60.635 5.945 60.805 7.22 ;
        RECT 55 5.945 55.17 7.22 ;
      LAYER met1 ;
        RECT 60.555 2.765 61.035 2.935 ;
        RECT 60.555 2.705 60.895 3.055 ;
        RECT 54.94 5.945 61.035 6.115 ;
        RECT 60.55 5.86 60.89 6.21 ;
        RECT 54.94 5.915 55.23 6.145 ;
      LAYER via1 ;
        RECT 60.65 5.96 60.8 6.11 ;
        RECT 60.655 2.805 60.805 2.955 ;
      LAYER mcon ;
        RECT 55 5.945 55.17 6.115 ;
        RECT 60.635 5.945 60.805 6.115 ;
        RECT 60.635 2.765 60.805 2.935 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 75.815 2.705 76.155 3.055 ;
        RECT 75.81 5.86 76.15 6.21 ;
        RECT 75.89 2.705 76.065 6.21 ;
      LAYER li1 ;
        RECT 75.895 1.66 76.065 2.935 ;
        RECT 75.895 5.945 76.065 7.22 ;
        RECT 70.26 5.945 70.43 7.22 ;
      LAYER met1 ;
        RECT 75.815 2.765 76.295 2.935 ;
        RECT 75.815 2.705 76.155 3.055 ;
        RECT 70.2 5.945 76.295 6.115 ;
        RECT 75.81 5.86 76.15 6.21 ;
        RECT 70.2 5.915 70.49 6.145 ;
      LAYER via1 ;
        RECT 75.91 5.96 76.06 6.11 ;
        RECT 75.915 2.805 76.065 2.955 ;
      LAYER mcon ;
        RECT 70.26 5.945 70.43 6.115 ;
        RECT 75.895 5.945 76.065 6.115 ;
        RECT 75.895 2.765 76.065 2.935 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 1.725 5.945 1.895 7.22 ;
      LAYER met1 ;
        RECT 1.665 5.945 2.125 6.115 ;
        RECT 1.665 5.915 1.955 6.145 ;
      LAYER mcon ;
        RECT 1.725 5.945 1.895 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.495 4.14 80.59 4.745 ;
        RECT 66.08 4.135 80.59 4.745 ;
        RECT 78.455 4.13 80.435 4.75 ;
        RECT 79.615 3.4 79.785 5.48 ;
        RECT 78.625 3.4 78.795 5.48 ;
        RECT 75.885 3.405 76.055 5.475 ;
        RECT 73.11 3.635 73.28 4.745 ;
        RECT 71.19 3.635 71.36 4.745 ;
        RECT 70.25 3.635 70.42 5.475 ;
        RECT 68.79 3.635 68.96 4.745 ;
        RECT 66.87 3.635 67.04 4.745 ;
        RECT 50.82 4.135 65.33 4.745 ;
        RECT 63.195 4.13 65.175 4.75 ;
        RECT 64.355 3.4 64.525 5.48 ;
        RECT 63.365 3.4 63.535 5.48 ;
        RECT 60.625 3.405 60.795 5.475 ;
        RECT 57.85 3.635 58.02 4.745 ;
        RECT 55.93 3.635 56.1 4.745 ;
        RECT 54.99 3.635 55.16 5.475 ;
        RECT 53.53 3.635 53.7 4.745 ;
        RECT 51.61 3.635 51.78 4.745 ;
        RECT 35.56 4.135 50.07 4.745 ;
        RECT 47.935 4.13 49.915 4.75 ;
        RECT 49.095 3.4 49.265 5.48 ;
        RECT 48.105 3.4 48.275 5.48 ;
        RECT 45.365 3.405 45.535 5.475 ;
        RECT 42.59 3.635 42.76 4.745 ;
        RECT 40.67 3.635 40.84 4.745 ;
        RECT 39.73 3.635 39.9 5.475 ;
        RECT 38.27 3.635 38.44 4.745 ;
        RECT 36.35 3.635 36.52 4.745 ;
        RECT 20.3 4.135 34.81 4.745 ;
        RECT 32.675 4.13 34.655 4.75 ;
        RECT 33.835 3.4 34.005 5.48 ;
        RECT 32.845 3.4 33.015 5.48 ;
        RECT 30.105 3.405 30.275 5.475 ;
        RECT 27.33 3.635 27.5 4.745 ;
        RECT 25.41 3.635 25.58 4.745 ;
        RECT 24.47 3.635 24.64 5.475 ;
        RECT 23.01 3.635 23.18 4.745 ;
        RECT 21.09 3.635 21.26 4.745 ;
        RECT 5.04 4.135 19.55 4.745 ;
        RECT 17.415 4.13 19.395 4.75 ;
        RECT 18.575 3.4 18.745 5.48 ;
        RECT 17.585 3.4 17.755 5.48 ;
        RECT 14.845 3.405 15.015 5.475 ;
        RECT 12.07 3.635 12.24 4.745 ;
        RECT 10.15 3.635 10.32 4.745 ;
        RECT 9.21 3.635 9.38 5.475 ;
        RECT 7.75 3.635 7.92 4.745 ;
        RECT 5.83 3.635 6 4.745 ;
        RECT 3.525 4.14 3.695 8.305 ;
        RECT 1.715 4.14 1.885 5.475 ;
      LAYER met1 ;
        RECT 1.495 4.14 80.59 4.745 ;
        RECT 66.08 4.135 80.59 4.745 ;
        RECT 78.455 4.13 80.435 4.75 ;
        RECT 66.08 3.98 74.82 4.745 ;
        RECT 50.82 4.135 65.33 4.745 ;
        RECT 63.195 4.13 65.175 4.75 ;
        RECT 50.82 3.98 59.56 4.745 ;
        RECT 35.56 4.135 50.07 4.745 ;
        RECT 47.935 4.13 49.915 4.75 ;
        RECT 35.56 3.98 44.3 4.745 ;
        RECT 20.3 4.135 34.81 4.745 ;
        RECT 32.675 4.13 34.655 4.75 ;
        RECT 20.3 3.98 29.04 4.745 ;
        RECT 5.04 4.135 19.55 4.745 ;
        RECT 17.415 4.13 19.395 4.75 ;
        RECT 5.04 3.98 13.78 4.745 ;
        RECT 3.465 6.655 3.755 6.885 ;
        RECT 3.295 6.685 3.755 6.855 ;
      LAYER mcon ;
        RECT 3.525 6.685 3.695 6.855 ;
        RECT 3.835 4.545 4.005 4.715 ;
        RECT 5.185 4.135 5.355 4.305 ;
        RECT 5.645 4.135 5.815 4.305 ;
        RECT 6.105 4.135 6.275 4.305 ;
        RECT 6.565 4.135 6.735 4.305 ;
        RECT 7.025 4.135 7.195 4.305 ;
        RECT 7.485 4.135 7.655 4.305 ;
        RECT 7.945 4.135 8.115 4.305 ;
        RECT 8.405 4.135 8.575 4.305 ;
        RECT 8.865 4.135 9.035 4.305 ;
        RECT 9.325 4.135 9.495 4.305 ;
        RECT 9.785 4.135 9.955 4.305 ;
        RECT 10.245 4.135 10.415 4.305 ;
        RECT 10.705 4.135 10.875 4.305 ;
        RECT 11.165 4.135 11.335 4.305 ;
        RECT 11.33 4.545 11.5 4.715 ;
        RECT 11.625 4.135 11.795 4.305 ;
        RECT 12.085 4.135 12.255 4.305 ;
        RECT 12.545 4.135 12.715 4.305 ;
        RECT 13.005 4.135 13.175 4.305 ;
        RECT 13.465 4.135 13.635 4.305 ;
        RECT 16.965 4.545 17.135 4.715 ;
        RECT 16.965 4.165 17.135 4.335 ;
        RECT 17.665 4.55 17.835 4.72 ;
        RECT 17.665 4.16 17.835 4.33 ;
        RECT 18.655 4.55 18.825 4.72 ;
        RECT 18.655 4.16 18.825 4.33 ;
        RECT 20.445 4.135 20.615 4.305 ;
        RECT 20.905 4.135 21.075 4.305 ;
        RECT 21.365 4.135 21.535 4.305 ;
        RECT 21.825 4.135 21.995 4.305 ;
        RECT 22.285 4.135 22.455 4.305 ;
        RECT 22.745 4.135 22.915 4.305 ;
        RECT 23.205 4.135 23.375 4.305 ;
        RECT 23.665 4.135 23.835 4.305 ;
        RECT 24.125 4.135 24.295 4.305 ;
        RECT 24.585 4.135 24.755 4.305 ;
        RECT 25.045 4.135 25.215 4.305 ;
        RECT 25.505 4.135 25.675 4.305 ;
        RECT 25.965 4.135 26.135 4.305 ;
        RECT 26.425 4.135 26.595 4.305 ;
        RECT 26.59 4.545 26.76 4.715 ;
        RECT 26.885 4.135 27.055 4.305 ;
        RECT 27.345 4.135 27.515 4.305 ;
        RECT 27.805 4.135 27.975 4.305 ;
        RECT 28.265 4.135 28.435 4.305 ;
        RECT 28.725 4.135 28.895 4.305 ;
        RECT 32.225 4.545 32.395 4.715 ;
        RECT 32.225 4.165 32.395 4.335 ;
        RECT 32.925 4.55 33.095 4.72 ;
        RECT 32.925 4.16 33.095 4.33 ;
        RECT 33.915 4.55 34.085 4.72 ;
        RECT 33.915 4.16 34.085 4.33 ;
        RECT 35.705 4.135 35.875 4.305 ;
        RECT 36.165 4.135 36.335 4.305 ;
        RECT 36.625 4.135 36.795 4.305 ;
        RECT 37.085 4.135 37.255 4.305 ;
        RECT 37.545 4.135 37.715 4.305 ;
        RECT 38.005 4.135 38.175 4.305 ;
        RECT 38.465 4.135 38.635 4.305 ;
        RECT 38.925 4.135 39.095 4.305 ;
        RECT 39.385 4.135 39.555 4.305 ;
        RECT 39.845 4.135 40.015 4.305 ;
        RECT 40.305 4.135 40.475 4.305 ;
        RECT 40.765 4.135 40.935 4.305 ;
        RECT 41.225 4.135 41.395 4.305 ;
        RECT 41.685 4.135 41.855 4.305 ;
        RECT 41.85 4.545 42.02 4.715 ;
        RECT 42.145 4.135 42.315 4.305 ;
        RECT 42.605 4.135 42.775 4.305 ;
        RECT 43.065 4.135 43.235 4.305 ;
        RECT 43.525 4.135 43.695 4.305 ;
        RECT 43.985 4.135 44.155 4.305 ;
        RECT 47.485 4.545 47.655 4.715 ;
        RECT 47.485 4.165 47.655 4.335 ;
        RECT 48.185 4.55 48.355 4.72 ;
        RECT 48.185 4.16 48.355 4.33 ;
        RECT 49.175 4.55 49.345 4.72 ;
        RECT 49.175 4.16 49.345 4.33 ;
        RECT 50.965 4.135 51.135 4.305 ;
        RECT 51.425 4.135 51.595 4.305 ;
        RECT 51.885 4.135 52.055 4.305 ;
        RECT 52.345 4.135 52.515 4.305 ;
        RECT 52.805 4.135 52.975 4.305 ;
        RECT 53.265 4.135 53.435 4.305 ;
        RECT 53.725 4.135 53.895 4.305 ;
        RECT 54.185 4.135 54.355 4.305 ;
        RECT 54.645 4.135 54.815 4.305 ;
        RECT 55.105 4.135 55.275 4.305 ;
        RECT 55.565 4.135 55.735 4.305 ;
        RECT 56.025 4.135 56.195 4.305 ;
        RECT 56.485 4.135 56.655 4.305 ;
        RECT 56.945 4.135 57.115 4.305 ;
        RECT 57.11 4.545 57.28 4.715 ;
        RECT 57.405 4.135 57.575 4.305 ;
        RECT 57.865 4.135 58.035 4.305 ;
        RECT 58.325 4.135 58.495 4.305 ;
        RECT 58.785 4.135 58.955 4.305 ;
        RECT 59.245 4.135 59.415 4.305 ;
        RECT 62.745 4.545 62.915 4.715 ;
        RECT 62.745 4.165 62.915 4.335 ;
        RECT 63.445 4.55 63.615 4.72 ;
        RECT 63.445 4.16 63.615 4.33 ;
        RECT 64.435 4.55 64.605 4.72 ;
        RECT 64.435 4.16 64.605 4.33 ;
        RECT 66.225 4.135 66.395 4.305 ;
        RECT 66.685 4.135 66.855 4.305 ;
        RECT 67.145 4.135 67.315 4.305 ;
        RECT 67.605 4.135 67.775 4.305 ;
        RECT 68.065 4.135 68.235 4.305 ;
        RECT 68.525 4.135 68.695 4.305 ;
        RECT 68.985 4.135 69.155 4.305 ;
        RECT 69.445 4.135 69.615 4.305 ;
        RECT 69.905 4.135 70.075 4.305 ;
        RECT 70.365 4.135 70.535 4.305 ;
        RECT 70.825 4.135 70.995 4.305 ;
        RECT 71.285 4.135 71.455 4.305 ;
        RECT 71.745 4.135 71.915 4.305 ;
        RECT 72.205 4.135 72.375 4.305 ;
        RECT 72.37 4.545 72.54 4.715 ;
        RECT 72.665 4.135 72.835 4.305 ;
        RECT 73.125 4.135 73.295 4.305 ;
        RECT 73.585 4.135 73.755 4.305 ;
        RECT 74.045 4.135 74.215 4.305 ;
        RECT 74.505 4.135 74.675 4.305 ;
        RECT 78.005 4.545 78.175 4.715 ;
        RECT 78.005 4.165 78.175 4.335 ;
        RECT 78.705 4.55 78.875 4.72 ;
        RECT 78.705 4.16 78.875 4.33 ;
        RECT 79.695 4.55 79.865 4.72 ;
        RECT 79.695 4.16 79.865 4.33 ;
    END
  END vccd1
  OBS
    LAYER met3 ;
      RECT 71.53 7.055 71.9 7.425 ;
      RECT 71.565 4.27 71.865 7.425 ;
      RECT 67.375 4.27 71.865 4.57 ;
      RECT 70.555 1.855 70.855 4.57 ;
      RECT 67.375 2.435 67.675 4.57 ;
      RECT 70.51 2.76 70.855 3.49 ;
      RECT 67.27 2.015 67.6 2.745 ;
      RECT 70.15 1.855 70.88 2.185 ;
      RECT 56.27 7.055 56.64 7.425 ;
      RECT 56.305 4.27 56.605 7.425 ;
      RECT 52.115 4.27 56.605 4.57 ;
      RECT 55.295 1.855 55.595 4.57 ;
      RECT 52.115 2.435 52.415 4.57 ;
      RECT 55.25 2.76 55.595 3.49 ;
      RECT 52.01 2.015 52.34 2.745 ;
      RECT 54.89 1.855 55.62 2.185 ;
      RECT 41.01 7.055 41.38 7.425 ;
      RECT 41.045 4.27 41.345 7.425 ;
      RECT 36.855 4.27 41.345 4.57 ;
      RECT 40.035 1.855 40.335 4.57 ;
      RECT 36.855 2.435 37.155 4.57 ;
      RECT 39.99 2.76 40.335 3.49 ;
      RECT 36.75 2.015 37.08 2.745 ;
      RECT 39.63 1.855 40.36 2.185 ;
      RECT 25.75 7.055 26.12 7.425 ;
      RECT 25.785 4.27 26.085 7.425 ;
      RECT 21.595 4.27 26.085 4.57 ;
      RECT 24.775 1.855 25.075 4.57 ;
      RECT 21.595 2.435 21.895 4.57 ;
      RECT 24.73 2.76 25.075 3.49 ;
      RECT 21.49 2.015 21.82 2.745 ;
      RECT 24.37 1.855 25.1 2.185 ;
      RECT 10.49 7.055 10.86 7.425 ;
      RECT 10.525 4.27 10.825 7.425 ;
      RECT 6.335 4.27 10.825 4.57 ;
      RECT 9.515 1.855 9.815 4.57 ;
      RECT 6.335 2.435 6.635 4.57 ;
      RECT 9.47 2.76 9.815 3.49 ;
      RECT 6.23 2.015 6.56 2.745 ;
      RECT 9.11 1.855 9.84 2.185 ;
      RECT 73.63 2.015 73.96 2.745 ;
      RECT 72.43 2.88 72.76 3.61 ;
      RECT 71.59 1.855 72.32 2.185 ;
      RECT 69.19 1.855 69.52 2.585 ;
      RECT 67.99 2.015 68.32 2.745 ;
      RECT 58.37 2.015 58.7 2.745 ;
      RECT 57.17 2.88 57.5 3.61 ;
      RECT 56.33 1.855 57.06 2.185 ;
      RECT 53.93 1.855 54.26 2.585 ;
      RECT 52.73 2.015 53.06 2.745 ;
      RECT 43.11 2.015 43.44 2.745 ;
      RECT 41.91 2.88 42.24 3.61 ;
      RECT 41.07 1.855 41.8 2.185 ;
      RECT 38.67 1.855 39 2.585 ;
      RECT 37.47 2.015 37.8 2.745 ;
      RECT 27.85 2.015 28.18 2.745 ;
      RECT 26.65 2.88 26.98 3.61 ;
      RECT 25.81 1.855 26.54 2.185 ;
      RECT 23.41 1.855 23.74 2.585 ;
      RECT 22.21 2.015 22.54 2.745 ;
      RECT 12.59 2.015 12.92 2.745 ;
      RECT 11.39 2.88 11.72 3.61 ;
      RECT 10.55 1.855 11.28 2.185 ;
      RECT 8.15 1.855 8.48 2.585 ;
      RECT 6.95 2.015 7.28 2.745 ;
    LAYER via2 ;
      RECT 73.695 2.48 73.895 2.68 ;
      RECT 72.495 3.04 72.695 3.24 ;
      RECT 71.655 1.92 71.855 2.12 ;
      RECT 71.615 7.14 71.815 7.34 ;
      RECT 70.575 2.825 70.775 3.025 ;
      RECT 70.215 1.92 70.415 2.12 ;
      RECT 69.255 1.92 69.455 2.12 ;
      RECT 68.055 2.48 68.255 2.68 ;
      RECT 67.335 2.48 67.535 2.68 ;
      RECT 58.435 2.48 58.635 2.68 ;
      RECT 57.235 3.04 57.435 3.24 ;
      RECT 56.395 1.92 56.595 2.12 ;
      RECT 56.355 7.14 56.555 7.34 ;
      RECT 55.315 2.825 55.515 3.025 ;
      RECT 54.955 1.92 55.155 2.12 ;
      RECT 53.995 1.92 54.195 2.12 ;
      RECT 52.795 2.48 52.995 2.68 ;
      RECT 52.075 2.48 52.275 2.68 ;
      RECT 43.175 2.48 43.375 2.68 ;
      RECT 41.975 3.04 42.175 3.24 ;
      RECT 41.135 1.92 41.335 2.12 ;
      RECT 41.095 7.14 41.295 7.34 ;
      RECT 40.055 2.825 40.255 3.025 ;
      RECT 39.695 1.92 39.895 2.12 ;
      RECT 38.735 1.92 38.935 2.12 ;
      RECT 37.535 2.48 37.735 2.68 ;
      RECT 36.815 2.48 37.015 2.68 ;
      RECT 27.915 2.48 28.115 2.68 ;
      RECT 26.715 3.04 26.915 3.24 ;
      RECT 25.875 1.92 26.075 2.12 ;
      RECT 25.835 7.14 26.035 7.34 ;
      RECT 24.795 2.825 24.995 3.025 ;
      RECT 24.435 1.92 24.635 2.12 ;
      RECT 23.475 1.92 23.675 2.12 ;
      RECT 22.275 2.48 22.475 2.68 ;
      RECT 21.555 2.48 21.755 2.68 ;
      RECT 12.655 2.48 12.855 2.68 ;
      RECT 11.455 3.04 11.655 3.24 ;
      RECT 10.615 1.92 10.815 2.12 ;
      RECT 10.575 7.14 10.775 7.34 ;
      RECT 9.535 2.825 9.735 3.025 ;
      RECT 9.175 1.92 9.375 2.12 ;
      RECT 8.215 1.92 8.415 2.12 ;
      RECT 7.015 2.48 7.215 2.68 ;
      RECT 6.295 2.48 6.495 2.68 ;
    LAYER met2 ;
      RECT 2.725 8.4 80.22 8.57 ;
      RECT 80.05 7.275 80.22 8.57 ;
      RECT 2.725 6.255 2.895 8.57 ;
      RECT 80.02 7.275 80.37 7.625 ;
      RECT 2.66 6.255 2.95 6.605 ;
      RECT 76.86 6.22 77.18 6.545 ;
      RECT 76.89 5.695 77.06 6.545 ;
      RECT 76.89 5.695 77.065 6.045 ;
      RECT 76.89 5.695 77.865 5.87 ;
      RECT 77.69 1.965 77.865 5.87 ;
      RECT 77.635 1.965 77.985 2.315 ;
      RECT 77.66 6.655 77.985 6.98 ;
      RECT 76.545 6.745 77.985 6.915 ;
      RECT 76.545 2.395 76.705 6.915 ;
      RECT 76.86 2.365 77.18 2.685 ;
      RECT 76.545 2.395 77.18 2.565 ;
      RECT 75.255 2.705 75.595 3.055 ;
      RECT 74.65 2.77 75.595 2.97 ;
      RECT 74.65 2.765 74.865 2.97 ;
      RECT 74.665 2.34 74.865 2.97 ;
      RECT 73.655 2.34 73.935 2.72 ;
      RECT 75.345 2.7 75.515 3.055 ;
      RECT 73.65 2.34 73.935 2.673 ;
      RECT 73.63 2.34 73.935 2.65 ;
      RECT 73.62 2.34 73.935 2.63 ;
      RECT 73.61 2.34 73.935 2.615 ;
      RECT 73.585 2.34 73.935 2.588 ;
      RECT 73.575 2.34 73.935 2.563 ;
      RECT 73.53 2.295 73.81 2.555 ;
      RECT 73.53 2.34 74.865 2.54 ;
      RECT 73.53 2.335 73.855 2.555 ;
      RECT 73.53 2.327 73.85 2.555 ;
      RECT 73.53 2.317 73.845 2.555 ;
      RECT 73.53 2.305 73.84 2.555 ;
      RECT 72.455 3 72.735 3.28 ;
      RECT 72.455 3 72.77 3.26 ;
      RECT 64.735 6.655 65.085 7.005 ;
      RECT 72.2 6.61 72.55 6.96 ;
      RECT 64.735 6.685 72.55 6.885 ;
      RECT 72.49 2.42 72.54 2.68 ;
      RECT 72.28 2.42 72.285 2.68 ;
      RECT 71.475 1.975 71.505 2.235 ;
      RECT 71.245 1.975 71.32 2.235 ;
      RECT 72.465 2.37 72.49 2.68 ;
      RECT 72.46 2.327 72.465 2.68 ;
      RECT 72.455 2.31 72.46 2.68 ;
      RECT 72.45 2.297 72.455 2.68 ;
      RECT 72.375 2.18 72.45 2.68 ;
      RECT 72.33 1.997 72.375 2.68 ;
      RECT 72.325 1.925 72.33 2.68 ;
      RECT 72.31 1.9 72.325 2.68 ;
      RECT 72.285 1.862 72.31 2.68 ;
      RECT 72.275 1.842 72.285 2.402 ;
      RECT 72.26 1.834 72.275 2.357 ;
      RECT 72.255 1.826 72.26 2.328 ;
      RECT 72.25 1.823 72.255 2.308 ;
      RECT 72.245 1.82 72.25 2.288 ;
      RECT 72.24 1.817 72.245 2.268 ;
      RECT 72.21 1.806 72.24 2.205 ;
      RECT 72.19 1.791 72.21 2.12 ;
      RECT 72.185 1.783 72.19 2.083 ;
      RECT 72.175 1.777 72.185 2.05 ;
      RECT 72.16 1.769 72.175 2.01 ;
      RECT 72.155 1.762 72.16 1.97 ;
      RECT 72.15 1.759 72.155 1.948 ;
      RECT 72.145 1.756 72.15 1.935 ;
      RECT 72.14 1.755 72.145 1.925 ;
      RECT 72.125 1.749 72.14 1.915 ;
      RECT 72.1 1.736 72.125 1.9 ;
      RECT 72.05 1.711 72.1 1.871 ;
      RECT 72.035 1.69 72.05 1.846 ;
      RECT 72.025 1.683 72.035 1.835 ;
      RECT 71.97 1.664 72.025 1.808 ;
      RECT 71.945 1.642 71.97 1.781 ;
      RECT 71.94 1.635 71.945 1.776 ;
      RECT 71.925 1.635 71.94 1.774 ;
      RECT 71.9 1.627 71.925 1.77 ;
      RECT 71.885 1.625 71.9 1.766 ;
      RECT 71.855 1.625 71.885 1.763 ;
      RECT 71.845 1.625 71.855 1.758 ;
      RECT 71.8 1.625 71.845 1.756 ;
      RECT 71.771 1.625 71.8 1.757 ;
      RECT 71.685 1.625 71.771 1.759 ;
      RECT 71.671 1.626 71.685 1.761 ;
      RECT 71.585 1.627 71.671 1.763 ;
      RECT 71.57 1.628 71.585 1.773 ;
      RECT 71.565 1.629 71.57 1.782 ;
      RECT 71.545 1.632 71.565 1.792 ;
      RECT 71.53 1.64 71.545 1.807 ;
      RECT 71.51 1.658 71.53 1.822 ;
      RECT 71.5 1.67 71.51 1.845 ;
      RECT 71.49 1.679 71.5 1.875 ;
      RECT 71.475 1.691 71.49 1.92 ;
      RECT 71.42 1.724 71.475 2.235 ;
      RECT 71.415 1.752 71.42 2.235 ;
      RECT 71.395 1.767 71.415 2.235 ;
      RECT 71.36 1.827 71.395 2.235 ;
      RECT 71.358 1.877 71.36 2.235 ;
      RECT 71.355 1.885 71.358 2.235 ;
      RECT 71.345 1.9 71.355 2.235 ;
      RECT 71.34 1.912 71.345 2.235 ;
      RECT 71.33 1.937 71.34 2.235 ;
      RECT 71.32 1.965 71.33 2.235 ;
      RECT 69.225 3.47 69.275 3.73 ;
      RECT 72.135 3.02 72.195 3.28 ;
      RECT 72.12 3.02 72.135 3.29 ;
      RECT 72.101 3.02 72.12 3.323 ;
      RECT 72.015 3.02 72.101 3.448 ;
      RECT 71.935 3.02 72.015 3.63 ;
      RECT 71.93 3.257 71.935 3.715 ;
      RECT 71.905 3.327 71.93 3.743 ;
      RECT 71.9 3.397 71.905 3.77 ;
      RECT 71.88 3.469 71.9 3.792 ;
      RECT 71.875 3.536 71.88 3.815 ;
      RECT 71.865 3.565 71.875 3.83 ;
      RECT 71.855 3.587 71.865 3.847 ;
      RECT 71.85 3.597 71.855 3.858 ;
      RECT 71.845 3.605 71.85 3.866 ;
      RECT 71.835 3.613 71.845 3.878 ;
      RECT 71.83 3.625 71.835 3.888 ;
      RECT 71.825 3.633 71.83 3.893 ;
      RECT 71.805 3.651 71.825 3.903 ;
      RECT 71.8 3.668 71.805 3.91 ;
      RECT 71.795 3.676 71.8 3.911 ;
      RECT 71.79 3.687 71.795 3.913 ;
      RECT 71.75 3.725 71.79 3.923 ;
      RECT 71.745 3.76 71.75 3.934 ;
      RECT 71.74 3.765 71.745 3.937 ;
      RECT 71.715 3.775 71.74 3.944 ;
      RECT 71.705 3.789 71.715 3.953 ;
      RECT 71.685 3.801 71.705 3.956 ;
      RECT 71.635 3.82 71.685 3.96 ;
      RECT 71.59 3.835 71.635 3.965 ;
      RECT 71.525 3.838 71.59 3.971 ;
      RECT 71.51 3.836 71.525 3.978 ;
      RECT 71.48 3.835 71.51 3.978 ;
      RECT 71.441 3.834 71.48 3.974 ;
      RECT 71.355 3.831 71.441 3.97 ;
      RECT 71.338 3.829 71.355 3.967 ;
      RECT 71.252 3.827 71.338 3.964 ;
      RECT 71.166 3.824 71.252 3.958 ;
      RECT 71.08 3.82 71.166 3.953 ;
      RECT 71.002 3.817 71.08 3.949 ;
      RECT 70.916 3.814 71.002 3.947 ;
      RECT 70.83 3.811 70.916 3.944 ;
      RECT 70.772 3.809 70.83 3.941 ;
      RECT 70.686 3.806 70.772 3.939 ;
      RECT 70.6 3.802 70.686 3.937 ;
      RECT 70.514 3.799 70.6 3.934 ;
      RECT 70.428 3.795 70.514 3.932 ;
      RECT 70.342 3.791 70.428 3.929 ;
      RECT 70.256 3.788 70.342 3.927 ;
      RECT 70.17 3.784 70.256 3.924 ;
      RECT 70.084 3.781 70.17 3.922 ;
      RECT 69.998 3.777 70.084 3.919 ;
      RECT 69.912 3.774 69.998 3.917 ;
      RECT 69.826 3.77 69.912 3.914 ;
      RECT 69.74 3.767 69.826 3.912 ;
      RECT 69.73 3.765 69.74 3.908 ;
      RECT 69.725 3.765 69.73 3.906 ;
      RECT 69.685 3.76 69.725 3.9 ;
      RECT 69.671 3.751 69.685 3.893 ;
      RECT 69.585 3.721 69.671 3.878 ;
      RECT 69.565 3.687 69.585 3.863 ;
      RECT 69.495 3.656 69.565 3.85 ;
      RECT 69.49 3.631 69.495 3.839 ;
      RECT 69.485 3.625 69.49 3.837 ;
      RECT 69.416 3.47 69.485 3.825 ;
      RECT 69.33 3.47 69.416 3.799 ;
      RECT 69.305 3.47 69.33 3.778 ;
      RECT 69.3 3.47 69.305 3.768 ;
      RECT 69.295 3.47 69.3 3.76 ;
      RECT 69.275 3.47 69.295 3.743 ;
      RECT 71.695 2.04 71.955 2.3 ;
      RECT 71.68 2.04 71.955 2.203 ;
      RECT 71.65 2.04 71.955 2.178 ;
      RECT 71.615 1.88 71.895 2.16 ;
      RECT 71.585 3.37 71.645 3.63 ;
      RECT 70.61 2.06 70.665 2.32 ;
      RECT 71.545 3.327 71.585 3.63 ;
      RECT 71.516 3.248 71.545 3.63 ;
      RECT 71.43 3.12 71.516 3.63 ;
      RECT 71.41 3 71.43 3.63 ;
      RECT 71.385 2.951 71.41 3.63 ;
      RECT 71.38 2.916 71.385 3.48 ;
      RECT 71.35 2.876 71.38 3.418 ;
      RECT 71.325 2.813 71.35 3.333 ;
      RECT 71.315 2.775 71.325 3.27 ;
      RECT 71.3 2.75 71.315 3.231 ;
      RECT 71.257 2.708 71.3 3.137 ;
      RECT 71.255 2.681 71.257 3.064 ;
      RECT 71.25 2.676 71.255 3.055 ;
      RECT 71.245 2.669 71.25 3.03 ;
      RECT 71.24 2.663 71.245 3.015 ;
      RECT 71.235 2.657 71.24 3.003 ;
      RECT 71.225 2.648 71.235 2.985 ;
      RECT 71.22 2.639 71.225 2.963 ;
      RECT 71.195 2.62 71.22 2.913 ;
      RECT 71.19 2.601 71.195 2.863 ;
      RECT 71.175 2.587 71.19 2.823 ;
      RECT 71.17 2.573 71.175 2.79 ;
      RECT 71.165 2.566 71.17 2.783 ;
      RECT 71.15 2.553 71.165 2.775 ;
      RECT 71.105 2.515 71.15 2.748 ;
      RECT 71.075 2.468 71.105 2.713 ;
      RECT 71.055 2.437 71.075 2.69 ;
      RECT 70.975 2.37 71.055 2.643 ;
      RECT 70.945 2.3 70.975 2.59 ;
      RECT 70.94 2.277 70.945 2.573 ;
      RECT 70.91 2.255 70.94 2.558 ;
      RECT 70.88 2.214 70.91 2.53 ;
      RECT 70.875 2.189 70.88 2.515 ;
      RECT 70.87 2.183 70.875 2.508 ;
      RECT 70.86 2.06 70.87 2.5 ;
      RECT 70.85 2.06 70.86 2.493 ;
      RECT 70.845 2.06 70.85 2.485 ;
      RECT 70.825 2.06 70.845 2.473 ;
      RECT 70.775 2.06 70.825 2.443 ;
      RECT 70.72 2.06 70.775 2.393 ;
      RECT 70.69 2.06 70.72 2.353 ;
      RECT 70.665 2.06 70.69 2.33 ;
      RECT 70.535 2.785 70.815 3.065 ;
      RECT 70.5 2.7 70.76 2.96 ;
      RECT 70.5 2.782 70.77 2.96 ;
      RECT 68.7 2.155 68.705 2.64 ;
      RECT 68.59 2.34 68.595 2.64 ;
      RECT 68.5 2.38 68.565 2.64 ;
      RECT 70.175 1.88 70.265 2.51 ;
      RECT 70.14 1.93 70.145 2.51 ;
      RECT 70.085 1.955 70.095 2.51 ;
      RECT 70.04 1.955 70.05 2.51 ;
      RECT 70.41 1.88 70.455 2.16 ;
      RECT 69.26 1.61 69.46 1.75 ;
      RECT 70.376 1.88 70.41 2.172 ;
      RECT 70.29 1.88 70.376 2.212 ;
      RECT 70.275 1.88 70.29 2.253 ;
      RECT 70.27 1.88 70.275 2.273 ;
      RECT 70.265 1.88 70.27 2.293 ;
      RECT 70.145 1.922 70.175 2.51 ;
      RECT 70.095 1.942 70.14 2.51 ;
      RECT 70.08 1.957 70.085 2.51 ;
      RECT 70.05 1.957 70.08 2.51 ;
      RECT 70.005 1.942 70.04 2.51 ;
      RECT 70 1.93 70.005 2.29 ;
      RECT 69.995 1.927 70 2.27 ;
      RECT 69.98 1.917 69.995 2.223 ;
      RECT 69.975 1.91 69.98 2.186 ;
      RECT 69.97 1.907 69.975 2.169 ;
      RECT 69.955 1.897 69.97 2.125 ;
      RECT 69.95 1.888 69.955 2.085 ;
      RECT 69.945 1.884 69.95 2.07 ;
      RECT 69.935 1.878 69.945 2.053 ;
      RECT 69.895 1.859 69.935 2.028 ;
      RECT 69.89 1.841 69.895 2.008 ;
      RECT 69.88 1.835 69.89 2.003 ;
      RECT 69.85 1.819 69.88 1.99 ;
      RECT 69.835 1.801 69.85 1.973 ;
      RECT 69.82 1.789 69.835 1.96 ;
      RECT 69.815 1.781 69.82 1.953 ;
      RECT 69.785 1.767 69.815 1.94 ;
      RECT 69.78 1.752 69.785 1.928 ;
      RECT 69.77 1.746 69.78 1.92 ;
      RECT 69.75 1.734 69.77 1.908 ;
      RECT 69.74 1.722 69.75 1.895 ;
      RECT 69.71 1.706 69.74 1.88 ;
      RECT 69.69 1.686 69.71 1.863 ;
      RECT 69.685 1.676 69.69 1.853 ;
      RECT 69.66 1.664 69.685 1.84 ;
      RECT 69.655 1.652 69.66 1.828 ;
      RECT 69.65 1.647 69.655 1.824 ;
      RECT 69.635 1.64 69.65 1.816 ;
      RECT 69.625 1.627 69.635 1.806 ;
      RECT 69.62 1.625 69.625 1.8 ;
      RECT 69.595 1.618 69.62 1.789 ;
      RECT 69.59 1.611 69.595 1.778 ;
      RECT 69.565 1.61 69.59 1.765 ;
      RECT 69.546 1.61 69.565 1.755 ;
      RECT 69.46 1.61 69.546 1.752 ;
      RECT 69.23 1.61 69.26 1.755 ;
      RECT 69.19 1.617 69.23 1.768 ;
      RECT 69.165 1.627 69.19 1.781 ;
      RECT 69.15 1.636 69.165 1.791 ;
      RECT 69.12 1.641 69.15 1.81 ;
      RECT 69.115 1.647 69.12 1.828 ;
      RECT 69.095 1.657 69.115 1.843 ;
      RECT 69.085 1.67 69.095 1.863 ;
      RECT 69.07 1.682 69.085 1.88 ;
      RECT 69.065 1.692 69.07 1.89 ;
      RECT 69.06 1.697 69.065 1.895 ;
      RECT 69.05 1.705 69.06 1.908 ;
      RECT 69 1.737 69.05 1.945 ;
      RECT 68.985 1.772 69 1.986 ;
      RECT 68.98 1.782 68.985 2.001 ;
      RECT 68.975 1.787 68.98 2.008 ;
      RECT 68.95 1.803 68.975 2.028 ;
      RECT 68.935 1.824 68.95 2.053 ;
      RECT 68.91 1.845 68.935 2.078 ;
      RECT 68.9 1.864 68.91 2.101 ;
      RECT 68.875 1.882 68.9 2.124 ;
      RECT 68.86 1.902 68.875 2.148 ;
      RECT 68.855 1.912 68.86 2.16 ;
      RECT 68.84 1.924 68.855 2.18 ;
      RECT 68.83 1.939 68.84 2.22 ;
      RECT 68.825 1.947 68.83 2.248 ;
      RECT 68.815 1.957 68.825 2.268 ;
      RECT 68.81 1.97 68.815 2.293 ;
      RECT 68.805 1.983 68.81 2.313 ;
      RECT 68.8 1.989 68.805 2.335 ;
      RECT 68.79 1.998 68.8 2.355 ;
      RECT 68.785 2.018 68.79 2.378 ;
      RECT 68.78 2.024 68.785 2.398 ;
      RECT 68.775 2.031 68.78 2.42 ;
      RECT 68.77 2.042 68.775 2.433 ;
      RECT 68.76 2.052 68.77 2.458 ;
      RECT 68.74 2.077 68.76 2.64 ;
      RECT 68.71 2.117 68.74 2.64 ;
      RECT 68.705 2.147 68.71 2.64 ;
      RECT 68.68 2.175 68.7 2.64 ;
      RECT 68.65 2.22 68.68 2.64 ;
      RECT 68.645 2.247 68.65 2.64 ;
      RECT 68.625 2.265 68.645 2.64 ;
      RECT 68.615 2.29 68.625 2.64 ;
      RECT 68.61 2.302 68.615 2.64 ;
      RECT 68.595 2.325 68.61 2.64 ;
      RECT 68.575 2.352 68.59 2.64 ;
      RECT 68.565 2.375 68.575 2.64 ;
      RECT 70.355 3.26 70.435 3.52 ;
      RECT 69.59 2.48 69.66 2.74 ;
      RECT 70.321 3.227 70.355 3.52 ;
      RECT 70.235 3.13 70.321 3.52 ;
      RECT 70.215 3.042 70.235 3.52 ;
      RECT 70.205 3.012 70.215 3.52 ;
      RECT 70.195 2.992 70.205 3.52 ;
      RECT 70.175 2.979 70.195 3.52 ;
      RECT 70.16 2.969 70.175 3.348 ;
      RECT 70.155 2.962 70.16 3.303 ;
      RECT 70.145 2.956 70.155 3.293 ;
      RECT 70.135 2.948 70.145 3.275 ;
      RECT 70.13 2.942 70.135 3.263 ;
      RECT 70.12 2.937 70.13 3.25 ;
      RECT 70.1 2.927 70.12 3.223 ;
      RECT 70.06 2.906 70.1 3.175 ;
      RECT 70.045 2.887 70.06 3.133 ;
      RECT 70.02 2.873 70.045 3.103 ;
      RECT 70.01 2.861 70.02 3.07 ;
      RECT 70.005 2.856 70.01 3.06 ;
      RECT 69.975 2.842 70.005 3.04 ;
      RECT 69.965 2.826 69.975 3.013 ;
      RECT 69.96 2.821 69.965 3.003 ;
      RECT 69.935 2.812 69.96 2.983 ;
      RECT 69.925 2.8 69.935 2.963 ;
      RECT 69.855 2.768 69.925 2.938 ;
      RECT 69.85 2.737 69.855 2.915 ;
      RECT 69.801 2.48 69.85 2.898 ;
      RECT 69.715 2.48 69.801 2.857 ;
      RECT 69.66 2.48 69.715 2.785 ;
      RECT 69.75 3.265 69.91 3.525 ;
      RECT 69.275 1.88 69.325 2.565 ;
      RECT 69.065 2.305 69.1 2.565 ;
      RECT 69.38 1.88 69.385 2.34 ;
      RECT 69.47 1.88 69.495 2.16 ;
      RECT 69.745 3.262 69.75 3.525 ;
      RECT 69.71 3.25 69.745 3.525 ;
      RECT 69.65 3.223 69.71 3.525 ;
      RECT 69.645 3.206 69.65 3.379 ;
      RECT 69.64 3.203 69.645 3.366 ;
      RECT 69.62 3.196 69.64 3.353 ;
      RECT 69.585 3.179 69.62 3.335 ;
      RECT 69.545 3.158 69.585 3.315 ;
      RECT 69.54 3.146 69.545 3.303 ;
      RECT 69.5 3.132 69.54 3.289 ;
      RECT 69.48 3.115 69.5 3.271 ;
      RECT 69.47 3.107 69.48 3.263 ;
      RECT 69.455 1.88 69.47 2.178 ;
      RECT 69.44 3.097 69.47 3.25 ;
      RECT 69.425 1.88 69.455 2.223 ;
      RECT 69.43 3.087 69.44 3.237 ;
      RECT 69.4 3.072 69.43 3.224 ;
      RECT 69.385 1.88 69.425 2.29 ;
      RECT 69.385 3.04 69.4 3.21 ;
      RECT 69.38 3.012 69.385 3.204 ;
      RECT 69.375 1.88 69.38 2.345 ;
      RECT 69.365 2.982 69.38 3.198 ;
      RECT 69.37 1.88 69.375 2.358 ;
      RECT 69.36 1.88 69.37 2.378 ;
      RECT 69.325 2.895 69.365 3.183 ;
      RECT 69.325 1.88 69.36 2.418 ;
      RECT 69.32 2.827 69.325 3.171 ;
      RECT 69.305 2.782 69.32 3.166 ;
      RECT 69.3 2.72 69.305 3.161 ;
      RECT 69.275 2.627 69.3 3.154 ;
      RECT 69.27 1.88 69.275 3.146 ;
      RECT 69.255 1.88 69.27 3.133 ;
      RECT 69.235 1.88 69.255 3.09 ;
      RECT 69.225 1.88 69.235 3.04 ;
      RECT 69.22 1.88 69.225 3.013 ;
      RECT 69.215 1.88 69.22 2.991 ;
      RECT 69.21 2.106 69.215 2.974 ;
      RECT 69.205 2.128 69.21 2.952 ;
      RECT 69.2 2.17 69.205 2.935 ;
      RECT 69.17 2.22 69.2 2.879 ;
      RECT 69.165 2.247 69.17 2.821 ;
      RECT 69.15 2.265 69.165 2.785 ;
      RECT 69.145 2.283 69.15 2.749 ;
      RECT 69.139 2.29 69.145 2.73 ;
      RECT 69.135 2.297 69.139 2.713 ;
      RECT 69.13 2.302 69.135 2.682 ;
      RECT 69.12 2.305 69.13 2.657 ;
      RECT 69.11 2.305 69.12 2.623 ;
      RECT 69.105 2.305 69.11 2.6 ;
      RECT 69.1 2.305 69.105 2.58 ;
      RECT 68.015 2.44 68.295 2.72 ;
      RECT 68.015 2.44 68.315 2.615 ;
      RECT 68.105 2.33 68.365 2.59 ;
      RECT 68.07 2.425 68.365 2.59 ;
      RECT 68.195 0.945 68.36 2.59 ;
      RECT 68.095 0.945 68.465 1.315 ;
      RECT 67.72 3.47 67.98 3.73 ;
      RECT 67.74 3.397 67.92 3.73 ;
      RECT 67.74 3.14 67.915 3.73 ;
      RECT 67.74 2.932 67.905 3.73 ;
      RECT 67.745 2.85 67.905 3.73 ;
      RECT 67.745 2.615 67.895 3.73 ;
      RECT 67.745 2.462 67.89 3.73 ;
      RECT 67.75 2.447 67.89 3.73 ;
      RECT 67.8 2.162 67.89 3.73 ;
      RECT 67.755 2.397 67.89 3.73 ;
      RECT 67.785 2.215 67.89 3.73 ;
      RECT 67.77 2.327 67.89 3.73 ;
      RECT 67.775 2.285 67.89 3.73 ;
      RECT 67.77 2.327 67.905 2.39 ;
      RECT 67.805 1.915 67.91 2.335 ;
      RECT 67.805 1.915 67.925 2.318 ;
      RECT 67.805 1.915 67.96 2.28 ;
      RECT 67.8 2.162 68.01 2.213 ;
      RECT 67.805 1.915 68.065 2.175 ;
      RECT 67.065 2.62 67.325 2.88 ;
      RECT 67.065 2.62 67.335 2.838 ;
      RECT 67.065 2.62 67.421 2.809 ;
      RECT 67.065 2.62 67.49 2.761 ;
      RECT 67.065 2.62 67.525 2.73 ;
      RECT 67.295 2.44 67.575 2.72 ;
      RECT 67.13 2.605 67.575 2.72 ;
      RECT 67.22 2.482 67.325 2.88 ;
      RECT 67.15 2.545 67.575 2.72 ;
      RECT 61.6 6.22 61.92 6.545 ;
      RECT 61.63 5.695 61.8 6.545 ;
      RECT 61.63 5.695 61.805 6.045 ;
      RECT 61.63 5.695 62.605 5.87 ;
      RECT 62.43 1.965 62.605 5.87 ;
      RECT 62.375 1.965 62.725 2.315 ;
      RECT 62.4 6.655 62.725 6.98 ;
      RECT 61.285 6.745 62.725 6.915 ;
      RECT 61.285 2.395 61.445 6.915 ;
      RECT 61.6 2.365 61.92 2.685 ;
      RECT 61.285 2.395 61.92 2.565 ;
      RECT 59.995 2.705 60.335 3.055 ;
      RECT 59.39 2.77 60.335 2.97 ;
      RECT 59.39 2.765 59.605 2.97 ;
      RECT 59.405 2.34 59.605 2.97 ;
      RECT 58.395 2.34 58.675 2.72 ;
      RECT 60.085 2.7 60.255 3.055 ;
      RECT 58.39 2.34 58.675 2.673 ;
      RECT 58.37 2.34 58.675 2.65 ;
      RECT 58.36 2.34 58.675 2.63 ;
      RECT 58.35 2.34 58.675 2.615 ;
      RECT 58.325 2.34 58.675 2.588 ;
      RECT 58.315 2.34 58.675 2.563 ;
      RECT 58.27 2.295 58.55 2.555 ;
      RECT 58.27 2.34 59.605 2.54 ;
      RECT 58.27 2.335 58.595 2.555 ;
      RECT 58.27 2.327 58.59 2.555 ;
      RECT 58.27 2.317 58.585 2.555 ;
      RECT 58.27 2.305 58.58 2.555 ;
      RECT 57.195 3 57.475 3.28 ;
      RECT 57.195 3 57.51 3.26 ;
      RECT 49.475 6.655 49.825 7.005 ;
      RECT 56.94 6.61 57.29 6.96 ;
      RECT 49.475 6.685 57.29 6.885 ;
      RECT 57.23 2.42 57.28 2.68 ;
      RECT 57.02 2.42 57.025 2.68 ;
      RECT 56.215 1.975 56.245 2.235 ;
      RECT 55.985 1.975 56.06 2.235 ;
      RECT 57.205 2.37 57.23 2.68 ;
      RECT 57.2 2.327 57.205 2.68 ;
      RECT 57.195 2.31 57.2 2.68 ;
      RECT 57.19 2.297 57.195 2.68 ;
      RECT 57.115 2.18 57.19 2.68 ;
      RECT 57.07 1.997 57.115 2.68 ;
      RECT 57.065 1.925 57.07 2.68 ;
      RECT 57.05 1.9 57.065 2.68 ;
      RECT 57.025 1.862 57.05 2.68 ;
      RECT 57.015 1.842 57.025 2.402 ;
      RECT 57 1.834 57.015 2.357 ;
      RECT 56.995 1.826 57 2.328 ;
      RECT 56.99 1.823 56.995 2.308 ;
      RECT 56.985 1.82 56.99 2.288 ;
      RECT 56.98 1.817 56.985 2.268 ;
      RECT 56.95 1.806 56.98 2.205 ;
      RECT 56.93 1.791 56.95 2.12 ;
      RECT 56.925 1.783 56.93 2.083 ;
      RECT 56.915 1.777 56.925 2.05 ;
      RECT 56.9 1.769 56.915 2.01 ;
      RECT 56.895 1.762 56.9 1.97 ;
      RECT 56.89 1.759 56.895 1.948 ;
      RECT 56.885 1.756 56.89 1.935 ;
      RECT 56.88 1.755 56.885 1.925 ;
      RECT 56.865 1.749 56.88 1.915 ;
      RECT 56.84 1.736 56.865 1.9 ;
      RECT 56.79 1.711 56.84 1.871 ;
      RECT 56.775 1.69 56.79 1.846 ;
      RECT 56.765 1.683 56.775 1.835 ;
      RECT 56.71 1.664 56.765 1.808 ;
      RECT 56.685 1.642 56.71 1.781 ;
      RECT 56.68 1.635 56.685 1.776 ;
      RECT 56.665 1.635 56.68 1.774 ;
      RECT 56.64 1.627 56.665 1.77 ;
      RECT 56.625 1.625 56.64 1.766 ;
      RECT 56.595 1.625 56.625 1.763 ;
      RECT 56.585 1.625 56.595 1.758 ;
      RECT 56.54 1.625 56.585 1.756 ;
      RECT 56.511 1.625 56.54 1.757 ;
      RECT 56.425 1.625 56.511 1.759 ;
      RECT 56.411 1.626 56.425 1.761 ;
      RECT 56.325 1.627 56.411 1.763 ;
      RECT 56.31 1.628 56.325 1.773 ;
      RECT 56.305 1.629 56.31 1.782 ;
      RECT 56.285 1.632 56.305 1.792 ;
      RECT 56.27 1.64 56.285 1.807 ;
      RECT 56.25 1.658 56.27 1.822 ;
      RECT 56.24 1.67 56.25 1.845 ;
      RECT 56.23 1.679 56.24 1.875 ;
      RECT 56.215 1.691 56.23 1.92 ;
      RECT 56.16 1.724 56.215 2.235 ;
      RECT 56.155 1.752 56.16 2.235 ;
      RECT 56.135 1.767 56.155 2.235 ;
      RECT 56.1 1.827 56.135 2.235 ;
      RECT 56.098 1.877 56.1 2.235 ;
      RECT 56.095 1.885 56.098 2.235 ;
      RECT 56.085 1.9 56.095 2.235 ;
      RECT 56.08 1.912 56.085 2.235 ;
      RECT 56.07 1.937 56.08 2.235 ;
      RECT 56.06 1.965 56.07 2.235 ;
      RECT 53.965 3.47 54.015 3.73 ;
      RECT 56.875 3.02 56.935 3.28 ;
      RECT 56.86 3.02 56.875 3.29 ;
      RECT 56.841 3.02 56.86 3.323 ;
      RECT 56.755 3.02 56.841 3.448 ;
      RECT 56.675 3.02 56.755 3.63 ;
      RECT 56.67 3.257 56.675 3.715 ;
      RECT 56.645 3.327 56.67 3.743 ;
      RECT 56.64 3.397 56.645 3.77 ;
      RECT 56.62 3.469 56.64 3.792 ;
      RECT 56.615 3.536 56.62 3.815 ;
      RECT 56.605 3.565 56.615 3.83 ;
      RECT 56.595 3.587 56.605 3.847 ;
      RECT 56.59 3.597 56.595 3.858 ;
      RECT 56.585 3.605 56.59 3.866 ;
      RECT 56.575 3.613 56.585 3.878 ;
      RECT 56.57 3.625 56.575 3.888 ;
      RECT 56.565 3.633 56.57 3.893 ;
      RECT 56.545 3.651 56.565 3.903 ;
      RECT 56.54 3.668 56.545 3.91 ;
      RECT 56.535 3.676 56.54 3.911 ;
      RECT 56.53 3.687 56.535 3.913 ;
      RECT 56.49 3.725 56.53 3.923 ;
      RECT 56.485 3.76 56.49 3.934 ;
      RECT 56.48 3.765 56.485 3.937 ;
      RECT 56.455 3.775 56.48 3.944 ;
      RECT 56.445 3.789 56.455 3.953 ;
      RECT 56.425 3.801 56.445 3.956 ;
      RECT 56.375 3.82 56.425 3.96 ;
      RECT 56.33 3.835 56.375 3.965 ;
      RECT 56.265 3.838 56.33 3.971 ;
      RECT 56.25 3.836 56.265 3.978 ;
      RECT 56.22 3.835 56.25 3.978 ;
      RECT 56.181 3.834 56.22 3.974 ;
      RECT 56.095 3.831 56.181 3.97 ;
      RECT 56.078 3.829 56.095 3.967 ;
      RECT 55.992 3.827 56.078 3.964 ;
      RECT 55.906 3.824 55.992 3.958 ;
      RECT 55.82 3.82 55.906 3.953 ;
      RECT 55.742 3.817 55.82 3.949 ;
      RECT 55.656 3.814 55.742 3.947 ;
      RECT 55.57 3.811 55.656 3.944 ;
      RECT 55.512 3.809 55.57 3.941 ;
      RECT 55.426 3.806 55.512 3.939 ;
      RECT 55.34 3.802 55.426 3.937 ;
      RECT 55.254 3.799 55.34 3.934 ;
      RECT 55.168 3.795 55.254 3.932 ;
      RECT 55.082 3.791 55.168 3.929 ;
      RECT 54.996 3.788 55.082 3.927 ;
      RECT 54.91 3.784 54.996 3.924 ;
      RECT 54.824 3.781 54.91 3.922 ;
      RECT 54.738 3.777 54.824 3.919 ;
      RECT 54.652 3.774 54.738 3.917 ;
      RECT 54.566 3.77 54.652 3.914 ;
      RECT 54.48 3.767 54.566 3.912 ;
      RECT 54.47 3.765 54.48 3.908 ;
      RECT 54.465 3.765 54.47 3.906 ;
      RECT 54.425 3.76 54.465 3.9 ;
      RECT 54.411 3.751 54.425 3.893 ;
      RECT 54.325 3.721 54.411 3.878 ;
      RECT 54.305 3.687 54.325 3.863 ;
      RECT 54.235 3.656 54.305 3.85 ;
      RECT 54.23 3.631 54.235 3.839 ;
      RECT 54.225 3.625 54.23 3.837 ;
      RECT 54.156 3.47 54.225 3.825 ;
      RECT 54.07 3.47 54.156 3.799 ;
      RECT 54.045 3.47 54.07 3.778 ;
      RECT 54.04 3.47 54.045 3.768 ;
      RECT 54.035 3.47 54.04 3.76 ;
      RECT 54.015 3.47 54.035 3.743 ;
      RECT 56.435 2.04 56.695 2.3 ;
      RECT 56.42 2.04 56.695 2.203 ;
      RECT 56.39 2.04 56.695 2.178 ;
      RECT 56.355 1.88 56.635 2.16 ;
      RECT 56.325 3.37 56.385 3.63 ;
      RECT 55.35 2.06 55.405 2.32 ;
      RECT 56.285 3.327 56.325 3.63 ;
      RECT 56.256 3.248 56.285 3.63 ;
      RECT 56.17 3.12 56.256 3.63 ;
      RECT 56.15 3 56.17 3.63 ;
      RECT 56.125 2.951 56.15 3.63 ;
      RECT 56.12 2.916 56.125 3.48 ;
      RECT 56.09 2.876 56.12 3.418 ;
      RECT 56.065 2.813 56.09 3.333 ;
      RECT 56.055 2.775 56.065 3.27 ;
      RECT 56.04 2.75 56.055 3.231 ;
      RECT 55.997 2.708 56.04 3.137 ;
      RECT 55.995 2.681 55.997 3.064 ;
      RECT 55.99 2.676 55.995 3.055 ;
      RECT 55.985 2.669 55.99 3.03 ;
      RECT 55.98 2.663 55.985 3.015 ;
      RECT 55.975 2.657 55.98 3.003 ;
      RECT 55.965 2.648 55.975 2.985 ;
      RECT 55.96 2.639 55.965 2.963 ;
      RECT 55.935 2.62 55.96 2.913 ;
      RECT 55.93 2.601 55.935 2.863 ;
      RECT 55.915 2.587 55.93 2.823 ;
      RECT 55.91 2.573 55.915 2.79 ;
      RECT 55.905 2.566 55.91 2.783 ;
      RECT 55.89 2.553 55.905 2.775 ;
      RECT 55.845 2.515 55.89 2.748 ;
      RECT 55.815 2.468 55.845 2.713 ;
      RECT 55.795 2.437 55.815 2.69 ;
      RECT 55.715 2.37 55.795 2.643 ;
      RECT 55.685 2.3 55.715 2.59 ;
      RECT 55.68 2.277 55.685 2.573 ;
      RECT 55.65 2.255 55.68 2.558 ;
      RECT 55.62 2.214 55.65 2.53 ;
      RECT 55.615 2.189 55.62 2.515 ;
      RECT 55.61 2.183 55.615 2.508 ;
      RECT 55.6 2.06 55.61 2.5 ;
      RECT 55.59 2.06 55.6 2.493 ;
      RECT 55.585 2.06 55.59 2.485 ;
      RECT 55.565 2.06 55.585 2.473 ;
      RECT 55.515 2.06 55.565 2.443 ;
      RECT 55.46 2.06 55.515 2.393 ;
      RECT 55.43 2.06 55.46 2.353 ;
      RECT 55.405 2.06 55.43 2.33 ;
      RECT 55.275 2.785 55.555 3.065 ;
      RECT 55.24 2.7 55.5 2.96 ;
      RECT 55.24 2.782 55.51 2.96 ;
      RECT 53.44 2.155 53.445 2.64 ;
      RECT 53.33 2.34 53.335 2.64 ;
      RECT 53.24 2.38 53.305 2.64 ;
      RECT 54.915 1.88 55.005 2.51 ;
      RECT 54.88 1.93 54.885 2.51 ;
      RECT 54.825 1.955 54.835 2.51 ;
      RECT 54.78 1.955 54.79 2.51 ;
      RECT 55.15 1.88 55.195 2.16 ;
      RECT 54 1.61 54.2 1.75 ;
      RECT 55.116 1.88 55.15 2.172 ;
      RECT 55.03 1.88 55.116 2.212 ;
      RECT 55.015 1.88 55.03 2.253 ;
      RECT 55.01 1.88 55.015 2.273 ;
      RECT 55.005 1.88 55.01 2.293 ;
      RECT 54.885 1.922 54.915 2.51 ;
      RECT 54.835 1.942 54.88 2.51 ;
      RECT 54.82 1.957 54.825 2.51 ;
      RECT 54.79 1.957 54.82 2.51 ;
      RECT 54.745 1.942 54.78 2.51 ;
      RECT 54.74 1.93 54.745 2.29 ;
      RECT 54.735 1.927 54.74 2.27 ;
      RECT 54.72 1.917 54.735 2.223 ;
      RECT 54.715 1.91 54.72 2.186 ;
      RECT 54.71 1.907 54.715 2.169 ;
      RECT 54.695 1.897 54.71 2.125 ;
      RECT 54.69 1.888 54.695 2.085 ;
      RECT 54.685 1.884 54.69 2.07 ;
      RECT 54.675 1.878 54.685 2.053 ;
      RECT 54.635 1.859 54.675 2.028 ;
      RECT 54.63 1.841 54.635 2.008 ;
      RECT 54.62 1.835 54.63 2.003 ;
      RECT 54.59 1.819 54.62 1.99 ;
      RECT 54.575 1.801 54.59 1.973 ;
      RECT 54.56 1.789 54.575 1.96 ;
      RECT 54.555 1.781 54.56 1.953 ;
      RECT 54.525 1.767 54.555 1.94 ;
      RECT 54.52 1.752 54.525 1.928 ;
      RECT 54.51 1.746 54.52 1.92 ;
      RECT 54.49 1.734 54.51 1.908 ;
      RECT 54.48 1.722 54.49 1.895 ;
      RECT 54.45 1.706 54.48 1.88 ;
      RECT 54.43 1.686 54.45 1.863 ;
      RECT 54.425 1.676 54.43 1.853 ;
      RECT 54.4 1.664 54.425 1.84 ;
      RECT 54.395 1.652 54.4 1.828 ;
      RECT 54.39 1.647 54.395 1.824 ;
      RECT 54.375 1.64 54.39 1.816 ;
      RECT 54.365 1.627 54.375 1.806 ;
      RECT 54.36 1.625 54.365 1.8 ;
      RECT 54.335 1.618 54.36 1.789 ;
      RECT 54.33 1.611 54.335 1.778 ;
      RECT 54.305 1.61 54.33 1.765 ;
      RECT 54.286 1.61 54.305 1.755 ;
      RECT 54.2 1.61 54.286 1.752 ;
      RECT 53.97 1.61 54 1.755 ;
      RECT 53.93 1.617 53.97 1.768 ;
      RECT 53.905 1.627 53.93 1.781 ;
      RECT 53.89 1.636 53.905 1.791 ;
      RECT 53.86 1.641 53.89 1.81 ;
      RECT 53.855 1.647 53.86 1.828 ;
      RECT 53.835 1.657 53.855 1.843 ;
      RECT 53.825 1.67 53.835 1.863 ;
      RECT 53.81 1.682 53.825 1.88 ;
      RECT 53.805 1.692 53.81 1.89 ;
      RECT 53.8 1.697 53.805 1.895 ;
      RECT 53.79 1.705 53.8 1.908 ;
      RECT 53.74 1.737 53.79 1.945 ;
      RECT 53.725 1.772 53.74 1.986 ;
      RECT 53.72 1.782 53.725 2.001 ;
      RECT 53.715 1.787 53.72 2.008 ;
      RECT 53.69 1.803 53.715 2.028 ;
      RECT 53.675 1.824 53.69 2.053 ;
      RECT 53.65 1.845 53.675 2.078 ;
      RECT 53.64 1.864 53.65 2.101 ;
      RECT 53.615 1.882 53.64 2.124 ;
      RECT 53.6 1.902 53.615 2.148 ;
      RECT 53.595 1.912 53.6 2.16 ;
      RECT 53.58 1.924 53.595 2.18 ;
      RECT 53.57 1.939 53.58 2.22 ;
      RECT 53.565 1.947 53.57 2.248 ;
      RECT 53.555 1.957 53.565 2.268 ;
      RECT 53.55 1.97 53.555 2.293 ;
      RECT 53.545 1.983 53.55 2.313 ;
      RECT 53.54 1.989 53.545 2.335 ;
      RECT 53.53 1.998 53.54 2.355 ;
      RECT 53.525 2.018 53.53 2.378 ;
      RECT 53.52 2.024 53.525 2.398 ;
      RECT 53.515 2.031 53.52 2.42 ;
      RECT 53.51 2.042 53.515 2.433 ;
      RECT 53.5 2.052 53.51 2.458 ;
      RECT 53.48 2.077 53.5 2.64 ;
      RECT 53.45 2.117 53.48 2.64 ;
      RECT 53.445 2.147 53.45 2.64 ;
      RECT 53.42 2.175 53.44 2.64 ;
      RECT 53.39 2.22 53.42 2.64 ;
      RECT 53.385 2.247 53.39 2.64 ;
      RECT 53.365 2.265 53.385 2.64 ;
      RECT 53.355 2.29 53.365 2.64 ;
      RECT 53.35 2.302 53.355 2.64 ;
      RECT 53.335 2.325 53.35 2.64 ;
      RECT 53.315 2.352 53.33 2.64 ;
      RECT 53.305 2.375 53.315 2.64 ;
      RECT 55.095 3.26 55.175 3.52 ;
      RECT 54.33 2.48 54.4 2.74 ;
      RECT 55.061 3.227 55.095 3.52 ;
      RECT 54.975 3.13 55.061 3.52 ;
      RECT 54.955 3.042 54.975 3.52 ;
      RECT 54.945 3.012 54.955 3.52 ;
      RECT 54.935 2.992 54.945 3.52 ;
      RECT 54.915 2.979 54.935 3.52 ;
      RECT 54.9 2.969 54.915 3.348 ;
      RECT 54.895 2.962 54.9 3.303 ;
      RECT 54.885 2.956 54.895 3.293 ;
      RECT 54.875 2.948 54.885 3.275 ;
      RECT 54.87 2.942 54.875 3.263 ;
      RECT 54.86 2.937 54.87 3.25 ;
      RECT 54.84 2.927 54.86 3.223 ;
      RECT 54.8 2.906 54.84 3.175 ;
      RECT 54.785 2.887 54.8 3.133 ;
      RECT 54.76 2.873 54.785 3.103 ;
      RECT 54.75 2.861 54.76 3.07 ;
      RECT 54.745 2.856 54.75 3.06 ;
      RECT 54.715 2.842 54.745 3.04 ;
      RECT 54.705 2.826 54.715 3.013 ;
      RECT 54.7 2.821 54.705 3.003 ;
      RECT 54.675 2.812 54.7 2.983 ;
      RECT 54.665 2.8 54.675 2.963 ;
      RECT 54.595 2.768 54.665 2.938 ;
      RECT 54.59 2.737 54.595 2.915 ;
      RECT 54.541 2.48 54.59 2.898 ;
      RECT 54.455 2.48 54.541 2.857 ;
      RECT 54.4 2.48 54.455 2.785 ;
      RECT 54.49 3.265 54.65 3.525 ;
      RECT 54.015 1.88 54.065 2.565 ;
      RECT 53.805 2.305 53.84 2.565 ;
      RECT 54.12 1.88 54.125 2.34 ;
      RECT 54.21 1.88 54.235 2.16 ;
      RECT 54.485 3.262 54.49 3.525 ;
      RECT 54.45 3.25 54.485 3.525 ;
      RECT 54.39 3.223 54.45 3.525 ;
      RECT 54.385 3.206 54.39 3.379 ;
      RECT 54.38 3.203 54.385 3.366 ;
      RECT 54.36 3.196 54.38 3.353 ;
      RECT 54.325 3.179 54.36 3.335 ;
      RECT 54.285 3.158 54.325 3.315 ;
      RECT 54.28 3.146 54.285 3.303 ;
      RECT 54.24 3.132 54.28 3.289 ;
      RECT 54.22 3.115 54.24 3.271 ;
      RECT 54.21 3.107 54.22 3.263 ;
      RECT 54.195 1.88 54.21 2.178 ;
      RECT 54.18 3.097 54.21 3.25 ;
      RECT 54.165 1.88 54.195 2.223 ;
      RECT 54.17 3.087 54.18 3.237 ;
      RECT 54.14 3.072 54.17 3.224 ;
      RECT 54.125 1.88 54.165 2.29 ;
      RECT 54.125 3.04 54.14 3.21 ;
      RECT 54.12 3.012 54.125 3.204 ;
      RECT 54.115 1.88 54.12 2.345 ;
      RECT 54.105 2.982 54.12 3.198 ;
      RECT 54.11 1.88 54.115 2.358 ;
      RECT 54.1 1.88 54.11 2.378 ;
      RECT 54.065 2.895 54.105 3.183 ;
      RECT 54.065 1.88 54.1 2.418 ;
      RECT 54.06 2.827 54.065 3.171 ;
      RECT 54.045 2.782 54.06 3.166 ;
      RECT 54.04 2.72 54.045 3.161 ;
      RECT 54.015 2.627 54.04 3.154 ;
      RECT 54.01 1.88 54.015 3.146 ;
      RECT 53.995 1.88 54.01 3.133 ;
      RECT 53.975 1.88 53.995 3.09 ;
      RECT 53.965 1.88 53.975 3.04 ;
      RECT 53.96 1.88 53.965 3.013 ;
      RECT 53.955 1.88 53.96 2.991 ;
      RECT 53.95 2.106 53.955 2.974 ;
      RECT 53.945 2.128 53.95 2.952 ;
      RECT 53.94 2.17 53.945 2.935 ;
      RECT 53.91 2.22 53.94 2.879 ;
      RECT 53.905 2.247 53.91 2.821 ;
      RECT 53.89 2.265 53.905 2.785 ;
      RECT 53.885 2.283 53.89 2.749 ;
      RECT 53.879 2.29 53.885 2.73 ;
      RECT 53.875 2.297 53.879 2.713 ;
      RECT 53.87 2.302 53.875 2.682 ;
      RECT 53.86 2.305 53.87 2.657 ;
      RECT 53.85 2.305 53.86 2.623 ;
      RECT 53.845 2.305 53.85 2.6 ;
      RECT 53.84 2.305 53.845 2.58 ;
      RECT 52.755 2.44 53.035 2.72 ;
      RECT 52.755 2.44 53.055 2.615 ;
      RECT 52.845 2.33 53.105 2.59 ;
      RECT 52.81 2.425 53.105 2.59 ;
      RECT 52.935 0.945 53.1 2.59 ;
      RECT 52.835 0.945 53.205 1.315 ;
      RECT 52.46 3.47 52.72 3.73 ;
      RECT 52.48 3.397 52.66 3.73 ;
      RECT 52.48 3.14 52.655 3.73 ;
      RECT 52.48 2.932 52.645 3.73 ;
      RECT 52.485 2.85 52.645 3.73 ;
      RECT 52.485 2.615 52.635 3.73 ;
      RECT 52.485 2.462 52.63 3.73 ;
      RECT 52.49 2.447 52.63 3.73 ;
      RECT 52.54 2.162 52.63 3.73 ;
      RECT 52.495 2.397 52.63 3.73 ;
      RECT 52.525 2.215 52.63 3.73 ;
      RECT 52.51 2.327 52.63 3.73 ;
      RECT 52.515 2.285 52.63 3.73 ;
      RECT 52.51 2.327 52.645 2.39 ;
      RECT 52.545 1.915 52.65 2.335 ;
      RECT 52.545 1.915 52.665 2.318 ;
      RECT 52.545 1.915 52.7 2.28 ;
      RECT 52.54 2.162 52.75 2.213 ;
      RECT 52.545 1.915 52.805 2.175 ;
      RECT 51.805 2.62 52.065 2.88 ;
      RECT 51.805 2.62 52.075 2.838 ;
      RECT 51.805 2.62 52.161 2.809 ;
      RECT 51.805 2.62 52.23 2.761 ;
      RECT 51.805 2.62 52.265 2.73 ;
      RECT 52.035 2.44 52.315 2.72 ;
      RECT 51.87 2.605 52.315 2.72 ;
      RECT 51.96 2.482 52.065 2.88 ;
      RECT 51.89 2.545 52.315 2.72 ;
      RECT 46.34 6.22 46.66 6.545 ;
      RECT 46.37 5.695 46.54 6.545 ;
      RECT 46.37 5.695 46.545 6.045 ;
      RECT 46.37 5.695 47.345 5.87 ;
      RECT 47.17 1.965 47.345 5.87 ;
      RECT 47.115 1.965 47.465 2.315 ;
      RECT 47.14 6.655 47.465 6.98 ;
      RECT 46.025 6.745 47.465 6.915 ;
      RECT 46.025 2.395 46.185 6.915 ;
      RECT 46.34 2.365 46.66 2.685 ;
      RECT 46.025 2.395 46.66 2.565 ;
      RECT 44.735 2.705 45.075 3.055 ;
      RECT 44.13 2.77 45.075 2.97 ;
      RECT 44.13 2.765 44.345 2.97 ;
      RECT 44.145 2.34 44.345 2.97 ;
      RECT 43.135 2.34 43.415 2.72 ;
      RECT 44.825 2.7 44.995 3.055 ;
      RECT 43.13 2.34 43.415 2.673 ;
      RECT 43.11 2.34 43.415 2.65 ;
      RECT 43.1 2.34 43.415 2.63 ;
      RECT 43.09 2.34 43.415 2.615 ;
      RECT 43.065 2.34 43.415 2.588 ;
      RECT 43.055 2.34 43.415 2.563 ;
      RECT 43.01 2.295 43.29 2.555 ;
      RECT 43.01 2.34 44.345 2.54 ;
      RECT 43.01 2.335 43.335 2.555 ;
      RECT 43.01 2.327 43.33 2.555 ;
      RECT 43.01 2.317 43.325 2.555 ;
      RECT 43.01 2.305 43.32 2.555 ;
      RECT 41.935 3 42.215 3.28 ;
      RECT 41.935 3 42.25 3.26 ;
      RECT 34.26 6.66 34.61 7.01 ;
      RECT 41.68 6.615 42.03 6.965 ;
      RECT 34.26 6.69 42.03 6.89 ;
      RECT 41.97 2.42 42.02 2.68 ;
      RECT 41.76 2.42 41.765 2.68 ;
      RECT 40.955 1.975 40.985 2.235 ;
      RECT 40.725 1.975 40.8 2.235 ;
      RECT 41.945 2.37 41.97 2.68 ;
      RECT 41.94 2.327 41.945 2.68 ;
      RECT 41.935 2.31 41.94 2.68 ;
      RECT 41.93 2.297 41.935 2.68 ;
      RECT 41.855 2.18 41.93 2.68 ;
      RECT 41.81 1.997 41.855 2.68 ;
      RECT 41.805 1.925 41.81 2.68 ;
      RECT 41.79 1.9 41.805 2.68 ;
      RECT 41.765 1.862 41.79 2.68 ;
      RECT 41.755 1.842 41.765 2.402 ;
      RECT 41.74 1.834 41.755 2.357 ;
      RECT 41.735 1.826 41.74 2.328 ;
      RECT 41.73 1.823 41.735 2.308 ;
      RECT 41.725 1.82 41.73 2.288 ;
      RECT 41.72 1.817 41.725 2.268 ;
      RECT 41.69 1.806 41.72 2.205 ;
      RECT 41.67 1.791 41.69 2.12 ;
      RECT 41.665 1.783 41.67 2.083 ;
      RECT 41.655 1.777 41.665 2.05 ;
      RECT 41.64 1.769 41.655 2.01 ;
      RECT 41.635 1.762 41.64 1.97 ;
      RECT 41.63 1.759 41.635 1.948 ;
      RECT 41.625 1.756 41.63 1.935 ;
      RECT 41.62 1.755 41.625 1.925 ;
      RECT 41.605 1.749 41.62 1.915 ;
      RECT 41.58 1.736 41.605 1.9 ;
      RECT 41.53 1.711 41.58 1.871 ;
      RECT 41.515 1.69 41.53 1.846 ;
      RECT 41.505 1.683 41.515 1.835 ;
      RECT 41.45 1.664 41.505 1.808 ;
      RECT 41.425 1.642 41.45 1.781 ;
      RECT 41.42 1.635 41.425 1.776 ;
      RECT 41.405 1.635 41.42 1.774 ;
      RECT 41.38 1.627 41.405 1.77 ;
      RECT 41.365 1.625 41.38 1.766 ;
      RECT 41.335 1.625 41.365 1.763 ;
      RECT 41.325 1.625 41.335 1.758 ;
      RECT 41.28 1.625 41.325 1.756 ;
      RECT 41.251 1.625 41.28 1.757 ;
      RECT 41.165 1.625 41.251 1.759 ;
      RECT 41.151 1.626 41.165 1.761 ;
      RECT 41.065 1.627 41.151 1.763 ;
      RECT 41.05 1.628 41.065 1.773 ;
      RECT 41.045 1.629 41.05 1.782 ;
      RECT 41.025 1.632 41.045 1.792 ;
      RECT 41.01 1.64 41.025 1.807 ;
      RECT 40.99 1.658 41.01 1.822 ;
      RECT 40.98 1.67 40.99 1.845 ;
      RECT 40.97 1.679 40.98 1.875 ;
      RECT 40.955 1.691 40.97 1.92 ;
      RECT 40.9 1.724 40.955 2.235 ;
      RECT 40.895 1.752 40.9 2.235 ;
      RECT 40.875 1.767 40.895 2.235 ;
      RECT 40.84 1.827 40.875 2.235 ;
      RECT 40.838 1.877 40.84 2.235 ;
      RECT 40.835 1.885 40.838 2.235 ;
      RECT 40.825 1.9 40.835 2.235 ;
      RECT 40.82 1.912 40.825 2.235 ;
      RECT 40.81 1.937 40.82 2.235 ;
      RECT 40.8 1.965 40.81 2.235 ;
      RECT 38.705 3.47 38.755 3.73 ;
      RECT 41.615 3.02 41.675 3.28 ;
      RECT 41.6 3.02 41.615 3.29 ;
      RECT 41.581 3.02 41.6 3.323 ;
      RECT 41.495 3.02 41.581 3.448 ;
      RECT 41.415 3.02 41.495 3.63 ;
      RECT 41.41 3.257 41.415 3.715 ;
      RECT 41.385 3.327 41.41 3.743 ;
      RECT 41.38 3.397 41.385 3.77 ;
      RECT 41.36 3.469 41.38 3.792 ;
      RECT 41.355 3.536 41.36 3.815 ;
      RECT 41.345 3.565 41.355 3.83 ;
      RECT 41.335 3.587 41.345 3.847 ;
      RECT 41.33 3.597 41.335 3.858 ;
      RECT 41.325 3.605 41.33 3.866 ;
      RECT 41.315 3.613 41.325 3.878 ;
      RECT 41.31 3.625 41.315 3.888 ;
      RECT 41.305 3.633 41.31 3.893 ;
      RECT 41.285 3.651 41.305 3.903 ;
      RECT 41.28 3.668 41.285 3.91 ;
      RECT 41.275 3.676 41.28 3.911 ;
      RECT 41.27 3.687 41.275 3.913 ;
      RECT 41.23 3.725 41.27 3.923 ;
      RECT 41.225 3.76 41.23 3.934 ;
      RECT 41.22 3.765 41.225 3.937 ;
      RECT 41.195 3.775 41.22 3.944 ;
      RECT 41.185 3.789 41.195 3.953 ;
      RECT 41.165 3.801 41.185 3.956 ;
      RECT 41.115 3.82 41.165 3.96 ;
      RECT 41.07 3.835 41.115 3.965 ;
      RECT 41.005 3.838 41.07 3.971 ;
      RECT 40.99 3.836 41.005 3.978 ;
      RECT 40.96 3.835 40.99 3.978 ;
      RECT 40.921 3.834 40.96 3.974 ;
      RECT 40.835 3.831 40.921 3.97 ;
      RECT 40.818 3.829 40.835 3.967 ;
      RECT 40.732 3.827 40.818 3.964 ;
      RECT 40.646 3.824 40.732 3.958 ;
      RECT 40.56 3.82 40.646 3.953 ;
      RECT 40.482 3.817 40.56 3.949 ;
      RECT 40.396 3.814 40.482 3.947 ;
      RECT 40.31 3.811 40.396 3.944 ;
      RECT 40.252 3.809 40.31 3.941 ;
      RECT 40.166 3.806 40.252 3.939 ;
      RECT 40.08 3.802 40.166 3.937 ;
      RECT 39.994 3.799 40.08 3.934 ;
      RECT 39.908 3.795 39.994 3.932 ;
      RECT 39.822 3.791 39.908 3.929 ;
      RECT 39.736 3.788 39.822 3.927 ;
      RECT 39.65 3.784 39.736 3.924 ;
      RECT 39.564 3.781 39.65 3.922 ;
      RECT 39.478 3.777 39.564 3.919 ;
      RECT 39.392 3.774 39.478 3.917 ;
      RECT 39.306 3.77 39.392 3.914 ;
      RECT 39.22 3.767 39.306 3.912 ;
      RECT 39.21 3.765 39.22 3.908 ;
      RECT 39.205 3.765 39.21 3.906 ;
      RECT 39.165 3.76 39.205 3.9 ;
      RECT 39.151 3.751 39.165 3.893 ;
      RECT 39.065 3.721 39.151 3.878 ;
      RECT 39.045 3.687 39.065 3.863 ;
      RECT 38.975 3.656 39.045 3.85 ;
      RECT 38.97 3.631 38.975 3.839 ;
      RECT 38.965 3.625 38.97 3.837 ;
      RECT 38.896 3.47 38.965 3.825 ;
      RECT 38.81 3.47 38.896 3.799 ;
      RECT 38.785 3.47 38.81 3.778 ;
      RECT 38.78 3.47 38.785 3.768 ;
      RECT 38.775 3.47 38.78 3.76 ;
      RECT 38.755 3.47 38.775 3.743 ;
      RECT 41.175 2.04 41.435 2.3 ;
      RECT 41.16 2.04 41.435 2.203 ;
      RECT 41.13 2.04 41.435 2.178 ;
      RECT 41.095 1.88 41.375 2.16 ;
      RECT 41.065 3.37 41.125 3.63 ;
      RECT 40.09 2.06 40.145 2.32 ;
      RECT 41.025 3.327 41.065 3.63 ;
      RECT 40.996 3.248 41.025 3.63 ;
      RECT 40.91 3.12 40.996 3.63 ;
      RECT 40.89 3 40.91 3.63 ;
      RECT 40.865 2.951 40.89 3.63 ;
      RECT 40.86 2.916 40.865 3.48 ;
      RECT 40.83 2.876 40.86 3.418 ;
      RECT 40.805 2.813 40.83 3.333 ;
      RECT 40.795 2.775 40.805 3.27 ;
      RECT 40.78 2.75 40.795 3.231 ;
      RECT 40.737 2.708 40.78 3.137 ;
      RECT 40.735 2.681 40.737 3.064 ;
      RECT 40.73 2.676 40.735 3.055 ;
      RECT 40.725 2.669 40.73 3.03 ;
      RECT 40.72 2.663 40.725 3.015 ;
      RECT 40.715 2.657 40.72 3.003 ;
      RECT 40.705 2.648 40.715 2.985 ;
      RECT 40.7 2.639 40.705 2.963 ;
      RECT 40.675 2.62 40.7 2.913 ;
      RECT 40.67 2.601 40.675 2.863 ;
      RECT 40.655 2.587 40.67 2.823 ;
      RECT 40.65 2.573 40.655 2.79 ;
      RECT 40.645 2.566 40.65 2.783 ;
      RECT 40.63 2.553 40.645 2.775 ;
      RECT 40.585 2.515 40.63 2.748 ;
      RECT 40.555 2.468 40.585 2.713 ;
      RECT 40.535 2.437 40.555 2.69 ;
      RECT 40.455 2.37 40.535 2.643 ;
      RECT 40.425 2.3 40.455 2.59 ;
      RECT 40.42 2.277 40.425 2.573 ;
      RECT 40.39 2.255 40.42 2.558 ;
      RECT 40.36 2.214 40.39 2.53 ;
      RECT 40.355 2.189 40.36 2.515 ;
      RECT 40.35 2.183 40.355 2.508 ;
      RECT 40.34 2.06 40.35 2.5 ;
      RECT 40.33 2.06 40.34 2.493 ;
      RECT 40.325 2.06 40.33 2.485 ;
      RECT 40.305 2.06 40.325 2.473 ;
      RECT 40.255 2.06 40.305 2.443 ;
      RECT 40.2 2.06 40.255 2.393 ;
      RECT 40.17 2.06 40.2 2.353 ;
      RECT 40.145 2.06 40.17 2.33 ;
      RECT 40.015 2.785 40.295 3.065 ;
      RECT 39.98 2.7 40.24 2.96 ;
      RECT 39.98 2.782 40.25 2.96 ;
      RECT 38.18 2.155 38.185 2.64 ;
      RECT 38.07 2.34 38.075 2.64 ;
      RECT 37.98 2.38 38.045 2.64 ;
      RECT 39.655 1.88 39.745 2.51 ;
      RECT 39.62 1.93 39.625 2.51 ;
      RECT 39.565 1.955 39.575 2.51 ;
      RECT 39.52 1.955 39.53 2.51 ;
      RECT 39.89 1.88 39.935 2.16 ;
      RECT 38.74 1.61 38.94 1.75 ;
      RECT 39.856 1.88 39.89 2.172 ;
      RECT 39.77 1.88 39.856 2.212 ;
      RECT 39.755 1.88 39.77 2.253 ;
      RECT 39.75 1.88 39.755 2.273 ;
      RECT 39.745 1.88 39.75 2.293 ;
      RECT 39.625 1.922 39.655 2.51 ;
      RECT 39.575 1.942 39.62 2.51 ;
      RECT 39.56 1.957 39.565 2.51 ;
      RECT 39.53 1.957 39.56 2.51 ;
      RECT 39.485 1.942 39.52 2.51 ;
      RECT 39.48 1.93 39.485 2.29 ;
      RECT 39.475 1.927 39.48 2.27 ;
      RECT 39.46 1.917 39.475 2.223 ;
      RECT 39.455 1.91 39.46 2.186 ;
      RECT 39.45 1.907 39.455 2.169 ;
      RECT 39.435 1.897 39.45 2.125 ;
      RECT 39.43 1.888 39.435 2.085 ;
      RECT 39.425 1.884 39.43 2.07 ;
      RECT 39.415 1.878 39.425 2.053 ;
      RECT 39.375 1.859 39.415 2.028 ;
      RECT 39.37 1.841 39.375 2.008 ;
      RECT 39.36 1.835 39.37 2.003 ;
      RECT 39.33 1.819 39.36 1.99 ;
      RECT 39.315 1.801 39.33 1.973 ;
      RECT 39.3 1.789 39.315 1.96 ;
      RECT 39.295 1.781 39.3 1.953 ;
      RECT 39.265 1.767 39.295 1.94 ;
      RECT 39.26 1.752 39.265 1.928 ;
      RECT 39.25 1.746 39.26 1.92 ;
      RECT 39.23 1.734 39.25 1.908 ;
      RECT 39.22 1.722 39.23 1.895 ;
      RECT 39.19 1.706 39.22 1.88 ;
      RECT 39.17 1.686 39.19 1.863 ;
      RECT 39.165 1.676 39.17 1.853 ;
      RECT 39.14 1.664 39.165 1.84 ;
      RECT 39.135 1.652 39.14 1.828 ;
      RECT 39.13 1.647 39.135 1.824 ;
      RECT 39.115 1.64 39.13 1.816 ;
      RECT 39.105 1.627 39.115 1.806 ;
      RECT 39.1 1.625 39.105 1.8 ;
      RECT 39.075 1.618 39.1 1.789 ;
      RECT 39.07 1.611 39.075 1.778 ;
      RECT 39.045 1.61 39.07 1.765 ;
      RECT 39.026 1.61 39.045 1.755 ;
      RECT 38.94 1.61 39.026 1.752 ;
      RECT 38.71 1.61 38.74 1.755 ;
      RECT 38.67 1.617 38.71 1.768 ;
      RECT 38.645 1.627 38.67 1.781 ;
      RECT 38.63 1.636 38.645 1.791 ;
      RECT 38.6 1.641 38.63 1.81 ;
      RECT 38.595 1.647 38.6 1.828 ;
      RECT 38.575 1.657 38.595 1.843 ;
      RECT 38.565 1.67 38.575 1.863 ;
      RECT 38.55 1.682 38.565 1.88 ;
      RECT 38.545 1.692 38.55 1.89 ;
      RECT 38.54 1.697 38.545 1.895 ;
      RECT 38.53 1.705 38.54 1.908 ;
      RECT 38.48 1.737 38.53 1.945 ;
      RECT 38.465 1.772 38.48 1.986 ;
      RECT 38.46 1.782 38.465 2.001 ;
      RECT 38.455 1.787 38.46 2.008 ;
      RECT 38.43 1.803 38.455 2.028 ;
      RECT 38.415 1.824 38.43 2.053 ;
      RECT 38.39 1.845 38.415 2.078 ;
      RECT 38.38 1.864 38.39 2.101 ;
      RECT 38.355 1.882 38.38 2.124 ;
      RECT 38.34 1.902 38.355 2.148 ;
      RECT 38.335 1.912 38.34 2.16 ;
      RECT 38.32 1.924 38.335 2.18 ;
      RECT 38.31 1.939 38.32 2.22 ;
      RECT 38.305 1.947 38.31 2.248 ;
      RECT 38.295 1.957 38.305 2.268 ;
      RECT 38.29 1.97 38.295 2.293 ;
      RECT 38.285 1.983 38.29 2.313 ;
      RECT 38.28 1.989 38.285 2.335 ;
      RECT 38.27 1.998 38.28 2.355 ;
      RECT 38.265 2.018 38.27 2.378 ;
      RECT 38.26 2.024 38.265 2.398 ;
      RECT 38.255 2.031 38.26 2.42 ;
      RECT 38.25 2.042 38.255 2.433 ;
      RECT 38.24 2.052 38.25 2.458 ;
      RECT 38.22 2.077 38.24 2.64 ;
      RECT 38.19 2.117 38.22 2.64 ;
      RECT 38.185 2.147 38.19 2.64 ;
      RECT 38.16 2.175 38.18 2.64 ;
      RECT 38.13 2.22 38.16 2.64 ;
      RECT 38.125 2.247 38.13 2.64 ;
      RECT 38.105 2.265 38.125 2.64 ;
      RECT 38.095 2.29 38.105 2.64 ;
      RECT 38.09 2.302 38.095 2.64 ;
      RECT 38.075 2.325 38.09 2.64 ;
      RECT 38.055 2.352 38.07 2.64 ;
      RECT 38.045 2.375 38.055 2.64 ;
      RECT 39.835 3.26 39.915 3.52 ;
      RECT 39.07 2.48 39.14 2.74 ;
      RECT 39.801 3.227 39.835 3.52 ;
      RECT 39.715 3.13 39.801 3.52 ;
      RECT 39.695 3.042 39.715 3.52 ;
      RECT 39.685 3.012 39.695 3.52 ;
      RECT 39.675 2.992 39.685 3.52 ;
      RECT 39.655 2.979 39.675 3.52 ;
      RECT 39.64 2.969 39.655 3.348 ;
      RECT 39.635 2.962 39.64 3.303 ;
      RECT 39.625 2.956 39.635 3.293 ;
      RECT 39.615 2.948 39.625 3.275 ;
      RECT 39.61 2.942 39.615 3.263 ;
      RECT 39.6 2.937 39.61 3.25 ;
      RECT 39.58 2.927 39.6 3.223 ;
      RECT 39.54 2.906 39.58 3.175 ;
      RECT 39.525 2.887 39.54 3.133 ;
      RECT 39.5 2.873 39.525 3.103 ;
      RECT 39.49 2.861 39.5 3.07 ;
      RECT 39.485 2.856 39.49 3.06 ;
      RECT 39.455 2.842 39.485 3.04 ;
      RECT 39.445 2.826 39.455 3.013 ;
      RECT 39.44 2.821 39.445 3.003 ;
      RECT 39.415 2.812 39.44 2.983 ;
      RECT 39.405 2.8 39.415 2.963 ;
      RECT 39.335 2.768 39.405 2.938 ;
      RECT 39.33 2.737 39.335 2.915 ;
      RECT 39.281 2.48 39.33 2.898 ;
      RECT 39.195 2.48 39.281 2.857 ;
      RECT 39.14 2.48 39.195 2.785 ;
      RECT 39.23 3.265 39.39 3.525 ;
      RECT 38.755 1.88 38.805 2.565 ;
      RECT 38.545 2.305 38.58 2.565 ;
      RECT 38.86 1.88 38.865 2.34 ;
      RECT 38.95 1.88 38.975 2.16 ;
      RECT 39.225 3.262 39.23 3.525 ;
      RECT 39.19 3.25 39.225 3.525 ;
      RECT 39.13 3.223 39.19 3.525 ;
      RECT 39.125 3.206 39.13 3.379 ;
      RECT 39.12 3.203 39.125 3.366 ;
      RECT 39.1 3.196 39.12 3.353 ;
      RECT 39.065 3.179 39.1 3.335 ;
      RECT 39.025 3.158 39.065 3.315 ;
      RECT 39.02 3.146 39.025 3.303 ;
      RECT 38.98 3.132 39.02 3.289 ;
      RECT 38.96 3.115 38.98 3.271 ;
      RECT 38.95 3.107 38.96 3.263 ;
      RECT 38.935 1.88 38.95 2.178 ;
      RECT 38.92 3.097 38.95 3.25 ;
      RECT 38.905 1.88 38.935 2.223 ;
      RECT 38.91 3.087 38.92 3.237 ;
      RECT 38.88 3.072 38.91 3.224 ;
      RECT 38.865 1.88 38.905 2.29 ;
      RECT 38.865 3.04 38.88 3.21 ;
      RECT 38.86 3.012 38.865 3.204 ;
      RECT 38.855 1.88 38.86 2.345 ;
      RECT 38.845 2.982 38.86 3.198 ;
      RECT 38.85 1.88 38.855 2.358 ;
      RECT 38.84 1.88 38.85 2.378 ;
      RECT 38.805 2.895 38.845 3.183 ;
      RECT 38.805 1.88 38.84 2.418 ;
      RECT 38.8 2.827 38.805 3.171 ;
      RECT 38.785 2.782 38.8 3.166 ;
      RECT 38.78 2.72 38.785 3.161 ;
      RECT 38.755 2.627 38.78 3.154 ;
      RECT 38.75 1.88 38.755 3.146 ;
      RECT 38.735 1.88 38.75 3.133 ;
      RECT 38.715 1.88 38.735 3.09 ;
      RECT 38.705 1.88 38.715 3.04 ;
      RECT 38.7 1.88 38.705 3.013 ;
      RECT 38.695 1.88 38.7 2.991 ;
      RECT 38.69 2.106 38.695 2.974 ;
      RECT 38.685 2.128 38.69 2.952 ;
      RECT 38.68 2.17 38.685 2.935 ;
      RECT 38.65 2.22 38.68 2.879 ;
      RECT 38.645 2.247 38.65 2.821 ;
      RECT 38.63 2.265 38.645 2.785 ;
      RECT 38.625 2.283 38.63 2.749 ;
      RECT 38.619 2.29 38.625 2.73 ;
      RECT 38.615 2.297 38.619 2.713 ;
      RECT 38.61 2.302 38.615 2.682 ;
      RECT 38.6 2.305 38.61 2.657 ;
      RECT 38.59 2.305 38.6 2.623 ;
      RECT 38.585 2.305 38.59 2.6 ;
      RECT 38.58 2.305 38.585 2.58 ;
      RECT 37.495 2.44 37.775 2.72 ;
      RECT 37.495 2.44 37.795 2.615 ;
      RECT 37.585 2.33 37.845 2.59 ;
      RECT 37.55 2.425 37.845 2.59 ;
      RECT 37.675 0.945 37.84 2.59 ;
      RECT 37.575 0.945 37.945 1.315 ;
      RECT 37.2 3.47 37.46 3.73 ;
      RECT 37.22 3.397 37.4 3.73 ;
      RECT 37.22 3.14 37.395 3.73 ;
      RECT 37.22 2.932 37.385 3.73 ;
      RECT 37.225 2.85 37.385 3.73 ;
      RECT 37.225 2.615 37.375 3.73 ;
      RECT 37.225 2.462 37.37 3.73 ;
      RECT 37.23 2.447 37.37 3.73 ;
      RECT 37.28 2.162 37.37 3.73 ;
      RECT 37.235 2.397 37.37 3.73 ;
      RECT 37.265 2.215 37.37 3.73 ;
      RECT 37.25 2.327 37.37 3.73 ;
      RECT 37.255 2.285 37.37 3.73 ;
      RECT 37.25 2.327 37.385 2.39 ;
      RECT 37.285 1.915 37.39 2.335 ;
      RECT 37.285 1.915 37.405 2.318 ;
      RECT 37.285 1.915 37.44 2.28 ;
      RECT 37.28 2.162 37.49 2.213 ;
      RECT 37.285 1.915 37.545 2.175 ;
      RECT 36.545 2.62 36.805 2.88 ;
      RECT 36.545 2.62 36.815 2.838 ;
      RECT 36.545 2.62 36.901 2.809 ;
      RECT 36.545 2.62 36.97 2.761 ;
      RECT 36.545 2.62 37.005 2.73 ;
      RECT 36.775 2.44 37.055 2.72 ;
      RECT 36.61 2.605 37.055 2.72 ;
      RECT 36.7 2.482 36.805 2.88 ;
      RECT 36.63 2.545 37.055 2.72 ;
      RECT 31.08 6.22 31.4 6.545 ;
      RECT 31.11 5.695 31.28 6.545 ;
      RECT 31.11 5.695 31.285 6.045 ;
      RECT 31.11 5.695 32.085 5.87 ;
      RECT 31.91 1.965 32.085 5.87 ;
      RECT 31.855 1.965 32.205 2.315 ;
      RECT 31.88 6.655 32.205 6.98 ;
      RECT 30.765 6.745 32.205 6.915 ;
      RECT 30.765 2.395 30.925 6.915 ;
      RECT 31.08 2.365 31.4 2.685 ;
      RECT 30.765 2.395 31.4 2.565 ;
      RECT 29.475 2.705 29.815 3.055 ;
      RECT 28.87 2.77 29.815 2.97 ;
      RECT 28.87 2.765 29.085 2.97 ;
      RECT 28.885 2.34 29.085 2.97 ;
      RECT 27.875 2.34 28.155 2.72 ;
      RECT 29.565 2.7 29.735 3.055 ;
      RECT 27.87 2.34 28.155 2.673 ;
      RECT 27.85 2.34 28.155 2.65 ;
      RECT 27.84 2.34 28.155 2.63 ;
      RECT 27.83 2.34 28.155 2.615 ;
      RECT 27.805 2.34 28.155 2.588 ;
      RECT 27.795 2.34 28.155 2.563 ;
      RECT 27.75 2.295 28.03 2.555 ;
      RECT 27.75 2.34 29.085 2.54 ;
      RECT 27.75 2.335 28.075 2.555 ;
      RECT 27.75 2.327 28.07 2.555 ;
      RECT 27.75 2.317 28.065 2.555 ;
      RECT 27.75 2.305 28.06 2.555 ;
      RECT 26.675 3 26.955 3.28 ;
      RECT 26.675 3 26.99 3.26 ;
      RECT 19 6.655 19.35 7.005 ;
      RECT 26.42 6.61 26.77 6.96 ;
      RECT 19 6.685 26.77 6.885 ;
      RECT 26.71 2.42 26.76 2.68 ;
      RECT 26.5 2.42 26.505 2.68 ;
      RECT 25.695 1.975 25.725 2.235 ;
      RECT 25.465 1.975 25.54 2.235 ;
      RECT 26.685 2.37 26.71 2.68 ;
      RECT 26.68 2.327 26.685 2.68 ;
      RECT 26.675 2.31 26.68 2.68 ;
      RECT 26.67 2.297 26.675 2.68 ;
      RECT 26.595 2.18 26.67 2.68 ;
      RECT 26.55 1.997 26.595 2.68 ;
      RECT 26.545 1.925 26.55 2.68 ;
      RECT 26.53 1.9 26.545 2.68 ;
      RECT 26.505 1.862 26.53 2.68 ;
      RECT 26.495 1.842 26.505 2.402 ;
      RECT 26.48 1.834 26.495 2.357 ;
      RECT 26.475 1.826 26.48 2.328 ;
      RECT 26.47 1.823 26.475 2.308 ;
      RECT 26.465 1.82 26.47 2.288 ;
      RECT 26.46 1.817 26.465 2.268 ;
      RECT 26.43 1.806 26.46 2.205 ;
      RECT 26.41 1.791 26.43 2.12 ;
      RECT 26.405 1.783 26.41 2.083 ;
      RECT 26.395 1.777 26.405 2.05 ;
      RECT 26.38 1.769 26.395 2.01 ;
      RECT 26.375 1.762 26.38 1.97 ;
      RECT 26.37 1.759 26.375 1.948 ;
      RECT 26.365 1.756 26.37 1.935 ;
      RECT 26.36 1.755 26.365 1.925 ;
      RECT 26.345 1.749 26.36 1.915 ;
      RECT 26.32 1.736 26.345 1.9 ;
      RECT 26.27 1.711 26.32 1.871 ;
      RECT 26.255 1.69 26.27 1.846 ;
      RECT 26.245 1.683 26.255 1.835 ;
      RECT 26.19 1.664 26.245 1.808 ;
      RECT 26.165 1.642 26.19 1.781 ;
      RECT 26.16 1.635 26.165 1.776 ;
      RECT 26.145 1.635 26.16 1.774 ;
      RECT 26.12 1.627 26.145 1.77 ;
      RECT 26.105 1.625 26.12 1.766 ;
      RECT 26.075 1.625 26.105 1.763 ;
      RECT 26.065 1.625 26.075 1.758 ;
      RECT 26.02 1.625 26.065 1.756 ;
      RECT 25.991 1.625 26.02 1.757 ;
      RECT 25.905 1.625 25.991 1.759 ;
      RECT 25.891 1.626 25.905 1.761 ;
      RECT 25.805 1.627 25.891 1.763 ;
      RECT 25.79 1.628 25.805 1.773 ;
      RECT 25.785 1.629 25.79 1.782 ;
      RECT 25.765 1.632 25.785 1.792 ;
      RECT 25.75 1.64 25.765 1.807 ;
      RECT 25.73 1.658 25.75 1.822 ;
      RECT 25.72 1.67 25.73 1.845 ;
      RECT 25.71 1.679 25.72 1.875 ;
      RECT 25.695 1.691 25.71 1.92 ;
      RECT 25.64 1.724 25.695 2.235 ;
      RECT 25.635 1.752 25.64 2.235 ;
      RECT 25.615 1.767 25.635 2.235 ;
      RECT 25.58 1.827 25.615 2.235 ;
      RECT 25.578 1.877 25.58 2.235 ;
      RECT 25.575 1.885 25.578 2.235 ;
      RECT 25.565 1.9 25.575 2.235 ;
      RECT 25.56 1.912 25.565 2.235 ;
      RECT 25.55 1.937 25.56 2.235 ;
      RECT 25.54 1.965 25.55 2.235 ;
      RECT 23.445 3.47 23.495 3.73 ;
      RECT 26.355 3.02 26.415 3.28 ;
      RECT 26.34 3.02 26.355 3.29 ;
      RECT 26.321 3.02 26.34 3.323 ;
      RECT 26.235 3.02 26.321 3.448 ;
      RECT 26.155 3.02 26.235 3.63 ;
      RECT 26.15 3.257 26.155 3.715 ;
      RECT 26.125 3.327 26.15 3.743 ;
      RECT 26.12 3.397 26.125 3.77 ;
      RECT 26.1 3.469 26.12 3.792 ;
      RECT 26.095 3.536 26.1 3.815 ;
      RECT 26.085 3.565 26.095 3.83 ;
      RECT 26.075 3.587 26.085 3.847 ;
      RECT 26.07 3.597 26.075 3.858 ;
      RECT 26.065 3.605 26.07 3.866 ;
      RECT 26.055 3.613 26.065 3.878 ;
      RECT 26.05 3.625 26.055 3.888 ;
      RECT 26.045 3.633 26.05 3.893 ;
      RECT 26.025 3.651 26.045 3.903 ;
      RECT 26.02 3.668 26.025 3.91 ;
      RECT 26.015 3.676 26.02 3.911 ;
      RECT 26.01 3.687 26.015 3.913 ;
      RECT 25.97 3.725 26.01 3.923 ;
      RECT 25.965 3.76 25.97 3.934 ;
      RECT 25.96 3.765 25.965 3.937 ;
      RECT 25.935 3.775 25.96 3.944 ;
      RECT 25.925 3.789 25.935 3.953 ;
      RECT 25.905 3.801 25.925 3.956 ;
      RECT 25.855 3.82 25.905 3.96 ;
      RECT 25.81 3.835 25.855 3.965 ;
      RECT 25.745 3.838 25.81 3.971 ;
      RECT 25.73 3.836 25.745 3.978 ;
      RECT 25.7 3.835 25.73 3.978 ;
      RECT 25.661 3.834 25.7 3.974 ;
      RECT 25.575 3.831 25.661 3.97 ;
      RECT 25.558 3.829 25.575 3.967 ;
      RECT 25.472 3.827 25.558 3.964 ;
      RECT 25.386 3.824 25.472 3.958 ;
      RECT 25.3 3.82 25.386 3.953 ;
      RECT 25.222 3.817 25.3 3.949 ;
      RECT 25.136 3.814 25.222 3.947 ;
      RECT 25.05 3.811 25.136 3.944 ;
      RECT 24.992 3.809 25.05 3.941 ;
      RECT 24.906 3.806 24.992 3.939 ;
      RECT 24.82 3.802 24.906 3.937 ;
      RECT 24.734 3.799 24.82 3.934 ;
      RECT 24.648 3.795 24.734 3.932 ;
      RECT 24.562 3.791 24.648 3.929 ;
      RECT 24.476 3.788 24.562 3.927 ;
      RECT 24.39 3.784 24.476 3.924 ;
      RECT 24.304 3.781 24.39 3.922 ;
      RECT 24.218 3.777 24.304 3.919 ;
      RECT 24.132 3.774 24.218 3.917 ;
      RECT 24.046 3.77 24.132 3.914 ;
      RECT 23.96 3.767 24.046 3.912 ;
      RECT 23.95 3.765 23.96 3.908 ;
      RECT 23.945 3.765 23.95 3.906 ;
      RECT 23.905 3.76 23.945 3.9 ;
      RECT 23.891 3.751 23.905 3.893 ;
      RECT 23.805 3.721 23.891 3.878 ;
      RECT 23.785 3.687 23.805 3.863 ;
      RECT 23.715 3.656 23.785 3.85 ;
      RECT 23.71 3.631 23.715 3.839 ;
      RECT 23.705 3.625 23.71 3.837 ;
      RECT 23.636 3.47 23.705 3.825 ;
      RECT 23.55 3.47 23.636 3.799 ;
      RECT 23.525 3.47 23.55 3.778 ;
      RECT 23.52 3.47 23.525 3.768 ;
      RECT 23.515 3.47 23.52 3.76 ;
      RECT 23.495 3.47 23.515 3.743 ;
      RECT 25.915 2.04 26.175 2.3 ;
      RECT 25.9 2.04 26.175 2.203 ;
      RECT 25.87 2.04 26.175 2.178 ;
      RECT 25.835 1.88 26.115 2.16 ;
      RECT 25.805 3.37 25.865 3.63 ;
      RECT 24.83 2.06 24.885 2.32 ;
      RECT 25.765 3.327 25.805 3.63 ;
      RECT 25.736 3.248 25.765 3.63 ;
      RECT 25.65 3.12 25.736 3.63 ;
      RECT 25.63 3 25.65 3.63 ;
      RECT 25.605 2.951 25.63 3.63 ;
      RECT 25.6 2.916 25.605 3.48 ;
      RECT 25.57 2.876 25.6 3.418 ;
      RECT 25.545 2.813 25.57 3.333 ;
      RECT 25.535 2.775 25.545 3.27 ;
      RECT 25.52 2.75 25.535 3.231 ;
      RECT 25.477 2.708 25.52 3.137 ;
      RECT 25.475 2.681 25.477 3.064 ;
      RECT 25.47 2.676 25.475 3.055 ;
      RECT 25.465 2.669 25.47 3.03 ;
      RECT 25.46 2.663 25.465 3.015 ;
      RECT 25.455 2.657 25.46 3.003 ;
      RECT 25.445 2.648 25.455 2.985 ;
      RECT 25.44 2.639 25.445 2.963 ;
      RECT 25.415 2.62 25.44 2.913 ;
      RECT 25.41 2.601 25.415 2.863 ;
      RECT 25.395 2.587 25.41 2.823 ;
      RECT 25.39 2.573 25.395 2.79 ;
      RECT 25.385 2.566 25.39 2.783 ;
      RECT 25.37 2.553 25.385 2.775 ;
      RECT 25.325 2.515 25.37 2.748 ;
      RECT 25.295 2.468 25.325 2.713 ;
      RECT 25.275 2.437 25.295 2.69 ;
      RECT 25.195 2.37 25.275 2.643 ;
      RECT 25.165 2.3 25.195 2.59 ;
      RECT 25.16 2.277 25.165 2.573 ;
      RECT 25.13 2.255 25.16 2.558 ;
      RECT 25.1 2.214 25.13 2.53 ;
      RECT 25.095 2.189 25.1 2.515 ;
      RECT 25.09 2.183 25.095 2.508 ;
      RECT 25.08 2.06 25.09 2.5 ;
      RECT 25.07 2.06 25.08 2.493 ;
      RECT 25.065 2.06 25.07 2.485 ;
      RECT 25.045 2.06 25.065 2.473 ;
      RECT 24.995 2.06 25.045 2.443 ;
      RECT 24.94 2.06 24.995 2.393 ;
      RECT 24.91 2.06 24.94 2.353 ;
      RECT 24.885 2.06 24.91 2.33 ;
      RECT 24.755 2.785 25.035 3.065 ;
      RECT 24.72 2.7 24.98 2.96 ;
      RECT 24.72 2.782 24.99 2.96 ;
      RECT 22.92 2.155 22.925 2.64 ;
      RECT 22.81 2.34 22.815 2.64 ;
      RECT 22.72 2.38 22.785 2.64 ;
      RECT 24.395 1.88 24.485 2.51 ;
      RECT 24.36 1.93 24.365 2.51 ;
      RECT 24.305 1.955 24.315 2.51 ;
      RECT 24.26 1.955 24.27 2.51 ;
      RECT 24.63 1.88 24.675 2.16 ;
      RECT 23.48 1.61 23.68 1.75 ;
      RECT 24.596 1.88 24.63 2.172 ;
      RECT 24.51 1.88 24.596 2.212 ;
      RECT 24.495 1.88 24.51 2.253 ;
      RECT 24.49 1.88 24.495 2.273 ;
      RECT 24.485 1.88 24.49 2.293 ;
      RECT 24.365 1.922 24.395 2.51 ;
      RECT 24.315 1.942 24.36 2.51 ;
      RECT 24.3 1.957 24.305 2.51 ;
      RECT 24.27 1.957 24.3 2.51 ;
      RECT 24.225 1.942 24.26 2.51 ;
      RECT 24.22 1.93 24.225 2.29 ;
      RECT 24.215 1.927 24.22 2.27 ;
      RECT 24.2 1.917 24.215 2.223 ;
      RECT 24.195 1.91 24.2 2.186 ;
      RECT 24.19 1.907 24.195 2.169 ;
      RECT 24.175 1.897 24.19 2.125 ;
      RECT 24.17 1.888 24.175 2.085 ;
      RECT 24.165 1.884 24.17 2.07 ;
      RECT 24.155 1.878 24.165 2.053 ;
      RECT 24.115 1.859 24.155 2.028 ;
      RECT 24.11 1.841 24.115 2.008 ;
      RECT 24.1 1.835 24.11 2.003 ;
      RECT 24.07 1.819 24.1 1.99 ;
      RECT 24.055 1.801 24.07 1.973 ;
      RECT 24.04 1.789 24.055 1.96 ;
      RECT 24.035 1.781 24.04 1.953 ;
      RECT 24.005 1.767 24.035 1.94 ;
      RECT 24 1.752 24.005 1.928 ;
      RECT 23.99 1.746 24 1.92 ;
      RECT 23.97 1.734 23.99 1.908 ;
      RECT 23.96 1.722 23.97 1.895 ;
      RECT 23.93 1.706 23.96 1.88 ;
      RECT 23.91 1.686 23.93 1.863 ;
      RECT 23.905 1.676 23.91 1.853 ;
      RECT 23.88 1.664 23.905 1.84 ;
      RECT 23.875 1.652 23.88 1.828 ;
      RECT 23.87 1.647 23.875 1.824 ;
      RECT 23.855 1.64 23.87 1.816 ;
      RECT 23.845 1.627 23.855 1.806 ;
      RECT 23.84 1.625 23.845 1.8 ;
      RECT 23.815 1.618 23.84 1.789 ;
      RECT 23.81 1.611 23.815 1.778 ;
      RECT 23.785 1.61 23.81 1.765 ;
      RECT 23.766 1.61 23.785 1.755 ;
      RECT 23.68 1.61 23.766 1.752 ;
      RECT 23.45 1.61 23.48 1.755 ;
      RECT 23.41 1.617 23.45 1.768 ;
      RECT 23.385 1.627 23.41 1.781 ;
      RECT 23.37 1.636 23.385 1.791 ;
      RECT 23.34 1.641 23.37 1.81 ;
      RECT 23.335 1.647 23.34 1.828 ;
      RECT 23.315 1.657 23.335 1.843 ;
      RECT 23.305 1.67 23.315 1.863 ;
      RECT 23.29 1.682 23.305 1.88 ;
      RECT 23.285 1.692 23.29 1.89 ;
      RECT 23.28 1.697 23.285 1.895 ;
      RECT 23.27 1.705 23.28 1.908 ;
      RECT 23.22 1.737 23.27 1.945 ;
      RECT 23.205 1.772 23.22 1.986 ;
      RECT 23.2 1.782 23.205 2.001 ;
      RECT 23.195 1.787 23.2 2.008 ;
      RECT 23.17 1.803 23.195 2.028 ;
      RECT 23.155 1.824 23.17 2.053 ;
      RECT 23.13 1.845 23.155 2.078 ;
      RECT 23.12 1.864 23.13 2.101 ;
      RECT 23.095 1.882 23.12 2.124 ;
      RECT 23.08 1.902 23.095 2.148 ;
      RECT 23.075 1.912 23.08 2.16 ;
      RECT 23.06 1.924 23.075 2.18 ;
      RECT 23.05 1.939 23.06 2.22 ;
      RECT 23.045 1.947 23.05 2.248 ;
      RECT 23.035 1.957 23.045 2.268 ;
      RECT 23.03 1.97 23.035 2.293 ;
      RECT 23.025 1.983 23.03 2.313 ;
      RECT 23.02 1.989 23.025 2.335 ;
      RECT 23.01 1.998 23.02 2.355 ;
      RECT 23.005 2.018 23.01 2.378 ;
      RECT 23 2.024 23.005 2.398 ;
      RECT 22.995 2.031 23 2.42 ;
      RECT 22.99 2.042 22.995 2.433 ;
      RECT 22.98 2.052 22.99 2.458 ;
      RECT 22.96 2.077 22.98 2.64 ;
      RECT 22.93 2.117 22.96 2.64 ;
      RECT 22.925 2.147 22.93 2.64 ;
      RECT 22.9 2.175 22.92 2.64 ;
      RECT 22.87 2.22 22.9 2.64 ;
      RECT 22.865 2.247 22.87 2.64 ;
      RECT 22.845 2.265 22.865 2.64 ;
      RECT 22.835 2.29 22.845 2.64 ;
      RECT 22.83 2.302 22.835 2.64 ;
      RECT 22.815 2.325 22.83 2.64 ;
      RECT 22.795 2.352 22.81 2.64 ;
      RECT 22.785 2.375 22.795 2.64 ;
      RECT 24.575 3.26 24.655 3.52 ;
      RECT 23.81 2.48 23.88 2.74 ;
      RECT 24.541 3.227 24.575 3.52 ;
      RECT 24.455 3.13 24.541 3.52 ;
      RECT 24.435 3.042 24.455 3.52 ;
      RECT 24.425 3.012 24.435 3.52 ;
      RECT 24.415 2.992 24.425 3.52 ;
      RECT 24.395 2.979 24.415 3.52 ;
      RECT 24.38 2.969 24.395 3.348 ;
      RECT 24.375 2.962 24.38 3.303 ;
      RECT 24.365 2.956 24.375 3.293 ;
      RECT 24.355 2.948 24.365 3.275 ;
      RECT 24.35 2.942 24.355 3.263 ;
      RECT 24.34 2.937 24.35 3.25 ;
      RECT 24.32 2.927 24.34 3.223 ;
      RECT 24.28 2.906 24.32 3.175 ;
      RECT 24.265 2.887 24.28 3.133 ;
      RECT 24.24 2.873 24.265 3.103 ;
      RECT 24.23 2.861 24.24 3.07 ;
      RECT 24.225 2.856 24.23 3.06 ;
      RECT 24.195 2.842 24.225 3.04 ;
      RECT 24.185 2.826 24.195 3.013 ;
      RECT 24.18 2.821 24.185 3.003 ;
      RECT 24.155 2.812 24.18 2.983 ;
      RECT 24.145 2.8 24.155 2.963 ;
      RECT 24.075 2.768 24.145 2.938 ;
      RECT 24.07 2.737 24.075 2.915 ;
      RECT 24.021 2.48 24.07 2.898 ;
      RECT 23.935 2.48 24.021 2.857 ;
      RECT 23.88 2.48 23.935 2.785 ;
      RECT 23.97 3.265 24.13 3.525 ;
      RECT 23.495 1.88 23.545 2.565 ;
      RECT 23.285 2.305 23.32 2.565 ;
      RECT 23.6 1.88 23.605 2.34 ;
      RECT 23.69 1.88 23.715 2.16 ;
      RECT 23.965 3.262 23.97 3.525 ;
      RECT 23.93 3.25 23.965 3.525 ;
      RECT 23.87 3.223 23.93 3.525 ;
      RECT 23.865 3.206 23.87 3.379 ;
      RECT 23.86 3.203 23.865 3.366 ;
      RECT 23.84 3.196 23.86 3.353 ;
      RECT 23.805 3.179 23.84 3.335 ;
      RECT 23.765 3.158 23.805 3.315 ;
      RECT 23.76 3.146 23.765 3.303 ;
      RECT 23.72 3.132 23.76 3.289 ;
      RECT 23.7 3.115 23.72 3.271 ;
      RECT 23.69 3.107 23.7 3.263 ;
      RECT 23.675 1.88 23.69 2.178 ;
      RECT 23.66 3.097 23.69 3.25 ;
      RECT 23.645 1.88 23.675 2.223 ;
      RECT 23.65 3.087 23.66 3.237 ;
      RECT 23.62 3.072 23.65 3.224 ;
      RECT 23.605 1.88 23.645 2.29 ;
      RECT 23.605 3.04 23.62 3.21 ;
      RECT 23.6 3.012 23.605 3.204 ;
      RECT 23.595 1.88 23.6 2.345 ;
      RECT 23.585 2.982 23.6 3.198 ;
      RECT 23.59 1.88 23.595 2.358 ;
      RECT 23.58 1.88 23.59 2.378 ;
      RECT 23.545 2.895 23.585 3.183 ;
      RECT 23.545 1.88 23.58 2.418 ;
      RECT 23.54 2.827 23.545 3.171 ;
      RECT 23.525 2.782 23.54 3.166 ;
      RECT 23.52 2.72 23.525 3.161 ;
      RECT 23.495 2.627 23.52 3.154 ;
      RECT 23.49 1.88 23.495 3.146 ;
      RECT 23.475 1.88 23.49 3.133 ;
      RECT 23.455 1.88 23.475 3.09 ;
      RECT 23.445 1.88 23.455 3.04 ;
      RECT 23.44 1.88 23.445 3.013 ;
      RECT 23.435 1.88 23.44 2.991 ;
      RECT 23.43 2.106 23.435 2.974 ;
      RECT 23.425 2.128 23.43 2.952 ;
      RECT 23.42 2.17 23.425 2.935 ;
      RECT 23.39 2.22 23.42 2.879 ;
      RECT 23.385 2.247 23.39 2.821 ;
      RECT 23.37 2.265 23.385 2.785 ;
      RECT 23.365 2.283 23.37 2.749 ;
      RECT 23.359 2.29 23.365 2.73 ;
      RECT 23.355 2.297 23.359 2.713 ;
      RECT 23.35 2.302 23.355 2.682 ;
      RECT 23.34 2.305 23.35 2.657 ;
      RECT 23.33 2.305 23.34 2.623 ;
      RECT 23.325 2.305 23.33 2.6 ;
      RECT 23.32 2.305 23.325 2.58 ;
      RECT 22.235 2.44 22.515 2.72 ;
      RECT 22.235 2.44 22.535 2.615 ;
      RECT 22.325 2.33 22.585 2.59 ;
      RECT 22.29 2.425 22.585 2.59 ;
      RECT 22.415 0.945 22.58 2.59 ;
      RECT 22.315 0.945 22.685 1.315 ;
      RECT 21.94 3.47 22.2 3.73 ;
      RECT 21.96 3.397 22.14 3.73 ;
      RECT 21.96 3.14 22.135 3.73 ;
      RECT 21.96 2.932 22.125 3.73 ;
      RECT 21.965 2.85 22.125 3.73 ;
      RECT 21.965 2.615 22.115 3.73 ;
      RECT 21.965 2.462 22.11 3.73 ;
      RECT 21.97 2.447 22.11 3.73 ;
      RECT 22.02 2.162 22.11 3.73 ;
      RECT 21.975 2.397 22.11 3.73 ;
      RECT 22.005 2.215 22.11 3.73 ;
      RECT 21.99 2.327 22.11 3.73 ;
      RECT 21.995 2.285 22.11 3.73 ;
      RECT 21.99 2.327 22.125 2.39 ;
      RECT 22.025 1.915 22.13 2.335 ;
      RECT 22.025 1.915 22.145 2.318 ;
      RECT 22.025 1.915 22.18 2.28 ;
      RECT 22.02 2.162 22.23 2.213 ;
      RECT 22.025 1.915 22.285 2.175 ;
      RECT 21.285 2.62 21.545 2.88 ;
      RECT 21.285 2.62 21.555 2.838 ;
      RECT 21.285 2.62 21.641 2.809 ;
      RECT 21.285 2.62 21.71 2.761 ;
      RECT 21.285 2.62 21.745 2.73 ;
      RECT 21.515 2.44 21.795 2.72 ;
      RECT 21.35 2.605 21.795 2.72 ;
      RECT 21.44 2.482 21.545 2.88 ;
      RECT 21.37 2.545 21.795 2.72 ;
      RECT 15.82 6.22 16.14 6.545 ;
      RECT 15.85 5.695 16.02 6.545 ;
      RECT 15.85 5.695 16.025 6.045 ;
      RECT 15.85 5.695 16.825 5.87 ;
      RECT 16.65 1.965 16.825 5.87 ;
      RECT 16.595 1.965 16.945 2.315 ;
      RECT 16.62 6.655 16.945 6.98 ;
      RECT 15.505 6.745 16.945 6.915 ;
      RECT 15.505 2.395 15.665 6.915 ;
      RECT 15.82 2.365 16.14 2.685 ;
      RECT 15.505 2.395 16.14 2.565 ;
      RECT 14.215 2.705 14.555 3.055 ;
      RECT 13.61 2.77 14.555 2.97 ;
      RECT 13.61 2.765 13.825 2.97 ;
      RECT 13.625 2.34 13.825 2.97 ;
      RECT 12.615 2.34 12.895 2.72 ;
      RECT 14.305 2.7 14.475 3.055 ;
      RECT 12.61 2.34 12.895 2.673 ;
      RECT 12.59 2.34 12.895 2.65 ;
      RECT 12.58 2.34 12.895 2.63 ;
      RECT 12.57 2.34 12.895 2.615 ;
      RECT 12.545 2.34 12.895 2.588 ;
      RECT 12.535 2.34 12.895 2.563 ;
      RECT 12.49 2.295 12.77 2.555 ;
      RECT 12.49 2.34 13.825 2.54 ;
      RECT 12.49 2.335 12.815 2.555 ;
      RECT 12.49 2.327 12.81 2.555 ;
      RECT 12.49 2.317 12.805 2.555 ;
      RECT 12.49 2.305 12.8 2.555 ;
      RECT 11.415 3 11.695 3.28 ;
      RECT 11.415 3 11.73 3.26 ;
      RECT 3.035 6.995 3.325 7.345 ;
      RECT 3.035 7.055 4.365 7.225 ;
      RECT 4.195 6.685 4.365 7.225 ;
      RECT 11.16 6.605 11.51 6.955 ;
      RECT 4.195 6.685 11.51 6.855 ;
      RECT 11.45 2.42 11.5 2.68 ;
      RECT 11.24 2.42 11.245 2.68 ;
      RECT 10.435 1.975 10.465 2.235 ;
      RECT 10.205 1.975 10.28 2.235 ;
      RECT 11.425 2.37 11.45 2.68 ;
      RECT 11.42 2.327 11.425 2.68 ;
      RECT 11.415 2.31 11.42 2.68 ;
      RECT 11.41 2.297 11.415 2.68 ;
      RECT 11.335 2.18 11.41 2.68 ;
      RECT 11.29 1.997 11.335 2.68 ;
      RECT 11.285 1.925 11.29 2.68 ;
      RECT 11.27 1.9 11.285 2.68 ;
      RECT 11.245 1.862 11.27 2.68 ;
      RECT 11.235 1.842 11.245 2.402 ;
      RECT 11.22 1.834 11.235 2.357 ;
      RECT 11.215 1.826 11.22 2.328 ;
      RECT 11.21 1.823 11.215 2.308 ;
      RECT 11.205 1.82 11.21 2.288 ;
      RECT 11.2 1.817 11.205 2.268 ;
      RECT 11.17 1.806 11.2 2.205 ;
      RECT 11.15 1.791 11.17 2.12 ;
      RECT 11.145 1.783 11.15 2.083 ;
      RECT 11.135 1.777 11.145 2.05 ;
      RECT 11.12 1.769 11.135 2.01 ;
      RECT 11.115 1.762 11.12 1.97 ;
      RECT 11.11 1.759 11.115 1.948 ;
      RECT 11.105 1.756 11.11 1.935 ;
      RECT 11.1 1.755 11.105 1.925 ;
      RECT 11.085 1.749 11.1 1.915 ;
      RECT 11.06 1.736 11.085 1.9 ;
      RECT 11.01 1.711 11.06 1.871 ;
      RECT 10.995 1.69 11.01 1.846 ;
      RECT 10.985 1.683 10.995 1.835 ;
      RECT 10.93 1.664 10.985 1.808 ;
      RECT 10.905 1.642 10.93 1.781 ;
      RECT 10.9 1.635 10.905 1.776 ;
      RECT 10.885 1.635 10.9 1.774 ;
      RECT 10.86 1.627 10.885 1.77 ;
      RECT 10.845 1.625 10.86 1.766 ;
      RECT 10.815 1.625 10.845 1.763 ;
      RECT 10.805 1.625 10.815 1.758 ;
      RECT 10.76 1.625 10.805 1.756 ;
      RECT 10.731 1.625 10.76 1.757 ;
      RECT 10.645 1.625 10.731 1.759 ;
      RECT 10.631 1.626 10.645 1.761 ;
      RECT 10.545 1.627 10.631 1.763 ;
      RECT 10.53 1.628 10.545 1.773 ;
      RECT 10.525 1.629 10.53 1.782 ;
      RECT 10.505 1.632 10.525 1.792 ;
      RECT 10.49 1.64 10.505 1.807 ;
      RECT 10.47 1.658 10.49 1.822 ;
      RECT 10.46 1.67 10.47 1.845 ;
      RECT 10.45 1.679 10.46 1.875 ;
      RECT 10.435 1.691 10.45 1.92 ;
      RECT 10.38 1.724 10.435 2.235 ;
      RECT 10.375 1.752 10.38 2.235 ;
      RECT 10.355 1.767 10.375 2.235 ;
      RECT 10.32 1.827 10.355 2.235 ;
      RECT 10.318 1.877 10.32 2.235 ;
      RECT 10.315 1.885 10.318 2.235 ;
      RECT 10.305 1.9 10.315 2.235 ;
      RECT 10.3 1.912 10.305 2.235 ;
      RECT 10.29 1.937 10.3 2.235 ;
      RECT 10.28 1.965 10.29 2.235 ;
      RECT 8.185 3.47 8.235 3.73 ;
      RECT 11.095 3.02 11.155 3.28 ;
      RECT 11.08 3.02 11.095 3.29 ;
      RECT 11.061 3.02 11.08 3.323 ;
      RECT 10.975 3.02 11.061 3.448 ;
      RECT 10.895 3.02 10.975 3.63 ;
      RECT 10.89 3.257 10.895 3.715 ;
      RECT 10.865 3.327 10.89 3.743 ;
      RECT 10.86 3.397 10.865 3.77 ;
      RECT 10.84 3.469 10.86 3.792 ;
      RECT 10.835 3.536 10.84 3.815 ;
      RECT 10.825 3.565 10.835 3.83 ;
      RECT 10.815 3.587 10.825 3.847 ;
      RECT 10.81 3.597 10.815 3.858 ;
      RECT 10.805 3.605 10.81 3.866 ;
      RECT 10.795 3.613 10.805 3.878 ;
      RECT 10.79 3.625 10.795 3.888 ;
      RECT 10.785 3.633 10.79 3.893 ;
      RECT 10.765 3.651 10.785 3.903 ;
      RECT 10.76 3.668 10.765 3.91 ;
      RECT 10.755 3.676 10.76 3.911 ;
      RECT 10.75 3.687 10.755 3.913 ;
      RECT 10.71 3.725 10.75 3.923 ;
      RECT 10.705 3.76 10.71 3.934 ;
      RECT 10.7 3.765 10.705 3.937 ;
      RECT 10.675 3.775 10.7 3.944 ;
      RECT 10.665 3.789 10.675 3.953 ;
      RECT 10.645 3.801 10.665 3.956 ;
      RECT 10.595 3.82 10.645 3.96 ;
      RECT 10.55 3.835 10.595 3.965 ;
      RECT 10.485 3.838 10.55 3.971 ;
      RECT 10.47 3.836 10.485 3.978 ;
      RECT 10.44 3.835 10.47 3.978 ;
      RECT 10.401 3.834 10.44 3.974 ;
      RECT 10.315 3.831 10.401 3.97 ;
      RECT 10.298 3.829 10.315 3.967 ;
      RECT 10.212 3.827 10.298 3.964 ;
      RECT 10.126 3.824 10.212 3.958 ;
      RECT 10.04 3.82 10.126 3.953 ;
      RECT 9.962 3.817 10.04 3.949 ;
      RECT 9.876 3.814 9.962 3.947 ;
      RECT 9.79 3.811 9.876 3.944 ;
      RECT 9.732 3.809 9.79 3.941 ;
      RECT 9.646 3.806 9.732 3.939 ;
      RECT 9.56 3.802 9.646 3.937 ;
      RECT 9.474 3.799 9.56 3.934 ;
      RECT 9.388 3.795 9.474 3.932 ;
      RECT 9.302 3.791 9.388 3.929 ;
      RECT 9.216 3.788 9.302 3.927 ;
      RECT 9.13 3.784 9.216 3.924 ;
      RECT 9.044 3.781 9.13 3.922 ;
      RECT 8.958 3.777 9.044 3.919 ;
      RECT 8.872 3.774 8.958 3.917 ;
      RECT 8.786 3.77 8.872 3.914 ;
      RECT 8.7 3.767 8.786 3.912 ;
      RECT 8.69 3.765 8.7 3.908 ;
      RECT 8.685 3.765 8.69 3.906 ;
      RECT 8.645 3.76 8.685 3.9 ;
      RECT 8.631 3.751 8.645 3.893 ;
      RECT 8.545 3.721 8.631 3.878 ;
      RECT 8.525 3.687 8.545 3.863 ;
      RECT 8.455 3.656 8.525 3.85 ;
      RECT 8.45 3.631 8.455 3.839 ;
      RECT 8.445 3.625 8.45 3.837 ;
      RECT 8.376 3.47 8.445 3.825 ;
      RECT 8.29 3.47 8.376 3.799 ;
      RECT 8.265 3.47 8.29 3.778 ;
      RECT 8.26 3.47 8.265 3.768 ;
      RECT 8.255 3.47 8.26 3.76 ;
      RECT 8.235 3.47 8.255 3.743 ;
      RECT 10.655 2.04 10.915 2.3 ;
      RECT 10.64 2.04 10.915 2.203 ;
      RECT 10.61 2.04 10.915 2.178 ;
      RECT 10.575 1.88 10.855 2.16 ;
      RECT 10.545 3.37 10.605 3.63 ;
      RECT 9.57 2.06 9.625 2.32 ;
      RECT 10.505 3.327 10.545 3.63 ;
      RECT 10.476 3.248 10.505 3.63 ;
      RECT 10.39 3.12 10.476 3.63 ;
      RECT 10.37 3 10.39 3.63 ;
      RECT 10.345 2.951 10.37 3.63 ;
      RECT 10.34 2.916 10.345 3.48 ;
      RECT 10.31 2.876 10.34 3.418 ;
      RECT 10.285 2.813 10.31 3.333 ;
      RECT 10.275 2.775 10.285 3.27 ;
      RECT 10.26 2.75 10.275 3.231 ;
      RECT 10.217 2.708 10.26 3.137 ;
      RECT 10.215 2.681 10.217 3.064 ;
      RECT 10.21 2.676 10.215 3.055 ;
      RECT 10.205 2.669 10.21 3.03 ;
      RECT 10.2 2.663 10.205 3.015 ;
      RECT 10.195 2.657 10.2 3.003 ;
      RECT 10.185 2.648 10.195 2.985 ;
      RECT 10.18 2.639 10.185 2.963 ;
      RECT 10.155 2.62 10.18 2.913 ;
      RECT 10.15 2.601 10.155 2.863 ;
      RECT 10.135 2.587 10.15 2.823 ;
      RECT 10.13 2.573 10.135 2.79 ;
      RECT 10.125 2.566 10.13 2.783 ;
      RECT 10.11 2.553 10.125 2.775 ;
      RECT 10.065 2.515 10.11 2.748 ;
      RECT 10.035 2.468 10.065 2.713 ;
      RECT 10.015 2.437 10.035 2.69 ;
      RECT 9.935 2.37 10.015 2.643 ;
      RECT 9.905 2.3 9.935 2.59 ;
      RECT 9.9 2.277 9.905 2.573 ;
      RECT 9.87 2.255 9.9 2.558 ;
      RECT 9.84 2.214 9.87 2.53 ;
      RECT 9.835 2.189 9.84 2.515 ;
      RECT 9.83 2.183 9.835 2.508 ;
      RECT 9.82 2.06 9.83 2.5 ;
      RECT 9.81 2.06 9.82 2.493 ;
      RECT 9.805 2.06 9.81 2.485 ;
      RECT 9.785 2.06 9.805 2.473 ;
      RECT 9.735 2.06 9.785 2.443 ;
      RECT 9.68 2.06 9.735 2.393 ;
      RECT 9.65 2.06 9.68 2.353 ;
      RECT 9.625 2.06 9.65 2.33 ;
      RECT 9.495 2.785 9.775 3.065 ;
      RECT 9.46 2.7 9.72 2.96 ;
      RECT 9.46 2.782 9.73 2.96 ;
      RECT 7.66 2.155 7.665 2.64 ;
      RECT 7.55 2.34 7.555 2.64 ;
      RECT 7.46 2.38 7.525 2.64 ;
      RECT 9.135 1.88 9.225 2.51 ;
      RECT 9.1 1.93 9.105 2.51 ;
      RECT 9.045 1.955 9.055 2.51 ;
      RECT 9 1.955 9.01 2.51 ;
      RECT 9.37 1.88 9.415 2.16 ;
      RECT 8.22 1.61 8.42 1.75 ;
      RECT 9.336 1.88 9.37 2.172 ;
      RECT 9.25 1.88 9.336 2.212 ;
      RECT 9.235 1.88 9.25 2.253 ;
      RECT 9.23 1.88 9.235 2.273 ;
      RECT 9.225 1.88 9.23 2.293 ;
      RECT 9.105 1.922 9.135 2.51 ;
      RECT 9.055 1.942 9.1 2.51 ;
      RECT 9.04 1.957 9.045 2.51 ;
      RECT 9.01 1.957 9.04 2.51 ;
      RECT 8.965 1.942 9 2.51 ;
      RECT 8.96 1.93 8.965 2.29 ;
      RECT 8.955 1.927 8.96 2.27 ;
      RECT 8.94 1.917 8.955 2.223 ;
      RECT 8.935 1.91 8.94 2.186 ;
      RECT 8.93 1.907 8.935 2.169 ;
      RECT 8.915 1.897 8.93 2.125 ;
      RECT 8.91 1.888 8.915 2.085 ;
      RECT 8.905 1.884 8.91 2.07 ;
      RECT 8.895 1.878 8.905 2.053 ;
      RECT 8.855 1.859 8.895 2.028 ;
      RECT 8.85 1.841 8.855 2.008 ;
      RECT 8.84 1.835 8.85 2.003 ;
      RECT 8.81 1.819 8.84 1.99 ;
      RECT 8.795 1.801 8.81 1.973 ;
      RECT 8.78 1.789 8.795 1.96 ;
      RECT 8.775 1.781 8.78 1.953 ;
      RECT 8.745 1.767 8.775 1.94 ;
      RECT 8.74 1.752 8.745 1.928 ;
      RECT 8.73 1.746 8.74 1.92 ;
      RECT 8.71 1.734 8.73 1.908 ;
      RECT 8.7 1.722 8.71 1.895 ;
      RECT 8.67 1.706 8.7 1.88 ;
      RECT 8.65 1.686 8.67 1.863 ;
      RECT 8.645 1.676 8.65 1.853 ;
      RECT 8.62 1.664 8.645 1.84 ;
      RECT 8.615 1.652 8.62 1.828 ;
      RECT 8.61 1.647 8.615 1.824 ;
      RECT 8.595 1.64 8.61 1.816 ;
      RECT 8.585 1.627 8.595 1.806 ;
      RECT 8.58 1.625 8.585 1.8 ;
      RECT 8.555 1.618 8.58 1.789 ;
      RECT 8.55 1.611 8.555 1.778 ;
      RECT 8.525 1.61 8.55 1.765 ;
      RECT 8.506 1.61 8.525 1.755 ;
      RECT 8.42 1.61 8.506 1.752 ;
      RECT 8.19 1.61 8.22 1.755 ;
      RECT 8.15 1.617 8.19 1.768 ;
      RECT 8.125 1.627 8.15 1.781 ;
      RECT 8.11 1.636 8.125 1.791 ;
      RECT 8.08 1.641 8.11 1.81 ;
      RECT 8.075 1.647 8.08 1.828 ;
      RECT 8.055 1.657 8.075 1.843 ;
      RECT 8.045 1.67 8.055 1.863 ;
      RECT 8.03 1.682 8.045 1.88 ;
      RECT 8.025 1.692 8.03 1.89 ;
      RECT 8.02 1.697 8.025 1.895 ;
      RECT 8.01 1.705 8.02 1.908 ;
      RECT 7.96 1.737 8.01 1.945 ;
      RECT 7.945 1.772 7.96 1.986 ;
      RECT 7.94 1.782 7.945 2.001 ;
      RECT 7.935 1.787 7.94 2.008 ;
      RECT 7.91 1.803 7.935 2.028 ;
      RECT 7.895 1.824 7.91 2.053 ;
      RECT 7.87 1.845 7.895 2.078 ;
      RECT 7.86 1.864 7.87 2.101 ;
      RECT 7.835 1.882 7.86 2.124 ;
      RECT 7.82 1.902 7.835 2.148 ;
      RECT 7.815 1.912 7.82 2.16 ;
      RECT 7.8 1.924 7.815 2.18 ;
      RECT 7.79 1.939 7.8 2.22 ;
      RECT 7.785 1.947 7.79 2.248 ;
      RECT 7.775 1.957 7.785 2.268 ;
      RECT 7.77 1.97 7.775 2.293 ;
      RECT 7.765 1.983 7.77 2.313 ;
      RECT 7.76 1.989 7.765 2.335 ;
      RECT 7.75 1.998 7.76 2.355 ;
      RECT 7.745 2.018 7.75 2.378 ;
      RECT 7.74 2.024 7.745 2.398 ;
      RECT 7.735 2.031 7.74 2.42 ;
      RECT 7.73 2.042 7.735 2.433 ;
      RECT 7.72 2.052 7.73 2.458 ;
      RECT 7.7 2.077 7.72 2.64 ;
      RECT 7.67 2.117 7.7 2.64 ;
      RECT 7.665 2.147 7.67 2.64 ;
      RECT 7.64 2.175 7.66 2.64 ;
      RECT 7.61 2.22 7.64 2.64 ;
      RECT 7.605 2.247 7.61 2.64 ;
      RECT 7.585 2.265 7.605 2.64 ;
      RECT 7.575 2.29 7.585 2.64 ;
      RECT 7.57 2.302 7.575 2.64 ;
      RECT 7.555 2.325 7.57 2.64 ;
      RECT 7.535 2.352 7.55 2.64 ;
      RECT 7.525 2.375 7.535 2.64 ;
      RECT 9.315 3.26 9.395 3.52 ;
      RECT 8.55 2.48 8.62 2.74 ;
      RECT 9.281 3.227 9.315 3.52 ;
      RECT 9.195 3.13 9.281 3.52 ;
      RECT 9.175 3.042 9.195 3.52 ;
      RECT 9.165 3.012 9.175 3.52 ;
      RECT 9.155 2.992 9.165 3.52 ;
      RECT 9.135 2.979 9.155 3.52 ;
      RECT 9.12 2.969 9.135 3.348 ;
      RECT 9.115 2.962 9.12 3.303 ;
      RECT 9.105 2.956 9.115 3.293 ;
      RECT 9.095 2.948 9.105 3.275 ;
      RECT 9.09 2.942 9.095 3.263 ;
      RECT 9.08 2.937 9.09 3.25 ;
      RECT 9.06 2.927 9.08 3.223 ;
      RECT 9.02 2.906 9.06 3.175 ;
      RECT 9.005 2.887 9.02 3.133 ;
      RECT 8.98 2.873 9.005 3.103 ;
      RECT 8.97 2.861 8.98 3.07 ;
      RECT 8.965 2.856 8.97 3.06 ;
      RECT 8.935 2.842 8.965 3.04 ;
      RECT 8.925 2.826 8.935 3.013 ;
      RECT 8.92 2.821 8.925 3.003 ;
      RECT 8.895 2.812 8.92 2.983 ;
      RECT 8.885 2.8 8.895 2.963 ;
      RECT 8.815 2.768 8.885 2.938 ;
      RECT 8.81 2.737 8.815 2.915 ;
      RECT 8.761 2.48 8.81 2.898 ;
      RECT 8.675 2.48 8.761 2.857 ;
      RECT 8.62 2.48 8.675 2.785 ;
      RECT 8.71 3.265 8.87 3.525 ;
      RECT 8.235 1.88 8.285 2.565 ;
      RECT 8.025 2.305 8.06 2.565 ;
      RECT 8.34 1.88 8.345 2.34 ;
      RECT 8.43 1.88 8.455 2.16 ;
      RECT 8.705 3.262 8.71 3.525 ;
      RECT 8.67 3.25 8.705 3.525 ;
      RECT 8.61 3.223 8.67 3.525 ;
      RECT 8.605 3.206 8.61 3.379 ;
      RECT 8.6 3.203 8.605 3.366 ;
      RECT 8.58 3.196 8.6 3.353 ;
      RECT 8.545 3.179 8.58 3.335 ;
      RECT 8.505 3.158 8.545 3.315 ;
      RECT 8.5 3.146 8.505 3.303 ;
      RECT 8.46 3.132 8.5 3.289 ;
      RECT 8.44 3.115 8.46 3.271 ;
      RECT 8.43 3.107 8.44 3.263 ;
      RECT 8.415 1.88 8.43 2.178 ;
      RECT 8.4 3.097 8.43 3.25 ;
      RECT 8.385 1.88 8.415 2.223 ;
      RECT 8.39 3.087 8.4 3.237 ;
      RECT 8.36 3.072 8.39 3.224 ;
      RECT 8.345 1.88 8.385 2.29 ;
      RECT 8.345 3.04 8.36 3.21 ;
      RECT 8.34 3.012 8.345 3.204 ;
      RECT 8.335 1.88 8.34 2.345 ;
      RECT 8.325 2.982 8.34 3.198 ;
      RECT 8.33 1.88 8.335 2.358 ;
      RECT 8.32 1.88 8.33 2.378 ;
      RECT 8.285 2.895 8.325 3.183 ;
      RECT 8.285 1.88 8.32 2.418 ;
      RECT 8.28 2.827 8.285 3.171 ;
      RECT 8.265 2.782 8.28 3.166 ;
      RECT 8.26 2.72 8.265 3.161 ;
      RECT 8.235 2.627 8.26 3.154 ;
      RECT 8.23 1.88 8.235 3.146 ;
      RECT 8.215 1.88 8.23 3.133 ;
      RECT 8.195 1.88 8.215 3.09 ;
      RECT 8.185 1.88 8.195 3.04 ;
      RECT 8.18 1.88 8.185 3.013 ;
      RECT 8.175 1.88 8.18 2.991 ;
      RECT 8.17 2.106 8.175 2.974 ;
      RECT 8.165 2.128 8.17 2.952 ;
      RECT 8.16 2.17 8.165 2.935 ;
      RECT 8.13 2.22 8.16 2.879 ;
      RECT 8.125 2.247 8.13 2.821 ;
      RECT 8.11 2.265 8.125 2.785 ;
      RECT 8.105 2.283 8.11 2.749 ;
      RECT 8.099 2.29 8.105 2.73 ;
      RECT 8.095 2.297 8.099 2.713 ;
      RECT 8.09 2.302 8.095 2.682 ;
      RECT 8.08 2.305 8.09 2.657 ;
      RECT 8.07 2.305 8.08 2.623 ;
      RECT 8.065 2.305 8.07 2.6 ;
      RECT 8.06 2.305 8.065 2.58 ;
      RECT 6.975 2.44 7.255 2.72 ;
      RECT 6.975 2.44 7.275 2.615 ;
      RECT 7.065 2.33 7.325 2.59 ;
      RECT 7.03 2.425 7.325 2.59 ;
      RECT 7.155 0.945 7.32 2.59 ;
      RECT 7.055 0.945 7.425 1.315 ;
      RECT 6.68 3.47 6.94 3.73 ;
      RECT 6.7 3.397 6.88 3.73 ;
      RECT 6.7 3.14 6.875 3.73 ;
      RECT 6.7 2.932 6.865 3.73 ;
      RECT 6.705 2.85 6.865 3.73 ;
      RECT 6.705 2.615 6.855 3.73 ;
      RECT 6.705 2.462 6.85 3.73 ;
      RECT 6.71 2.447 6.85 3.73 ;
      RECT 6.76 2.162 6.85 3.73 ;
      RECT 6.715 2.397 6.85 3.73 ;
      RECT 6.745 2.215 6.85 3.73 ;
      RECT 6.73 2.327 6.85 3.73 ;
      RECT 6.735 2.285 6.85 3.73 ;
      RECT 6.73 2.327 6.865 2.39 ;
      RECT 6.765 1.915 6.87 2.335 ;
      RECT 6.765 1.915 6.885 2.318 ;
      RECT 6.765 1.915 6.92 2.28 ;
      RECT 6.76 2.162 6.97 2.213 ;
      RECT 6.765 1.915 7.025 2.175 ;
      RECT 6.025 2.62 6.285 2.88 ;
      RECT 6.025 2.62 6.295 2.838 ;
      RECT 6.025 2.62 6.381 2.809 ;
      RECT 6.025 2.62 6.45 2.761 ;
      RECT 6.025 2.62 6.485 2.73 ;
      RECT 6.255 2.44 6.535 2.72 ;
      RECT 6.09 2.605 6.535 2.72 ;
      RECT 6.18 2.482 6.285 2.88 ;
      RECT 6.11 2.545 6.535 2.72 ;
      RECT 71.53 7.055 71.9 7.425 ;
      RECT 56.27 7.055 56.64 7.425 ;
      RECT 41.01 7.055 41.38 7.425 ;
      RECT 25.75 7.055 26.12 7.425 ;
      RECT 10.49 7.055 10.86 7.425 ;
    LAYER via1 ;
      RECT 80.12 7.375 80.27 7.525 ;
      RECT 77.75 6.74 77.9 6.89 ;
      RECT 77.735 2.065 77.885 2.215 ;
      RECT 76.945 2.45 77.095 2.6 ;
      RECT 76.945 6.325 77.095 6.475 ;
      RECT 75.355 2.805 75.505 2.955 ;
      RECT 73.585 2.35 73.735 2.5 ;
      RECT 72.565 3.055 72.715 3.205 ;
      RECT 72.335 2.475 72.485 2.625 ;
      RECT 72.3 6.71 72.45 6.86 ;
      RECT 71.99 3.075 72.14 3.225 ;
      RECT 71.75 2.095 71.9 2.245 ;
      RECT 71.64 7.165 71.79 7.315 ;
      RECT 71.44 3.425 71.59 3.575 ;
      RECT 71.3 2.03 71.45 2.18 ;
      RECT 70.665 2.115 70.815 2.265 ;
      RECT 70.555 2.755 70.705 2.905 ;
      RECT 70.23 3.315 70.38 3.465 ;
      RECT 70.06 2.305 70.21 2.455 ;
      RECT 69.705 3.32 69.855 3.47 ;
      RECT 69.645 2.535 69.795 2.685 ;
      RECT 69.28 3.525 69.43 3.675 ;
      RECT 69.12 2.36 69.27 2.51 ;
      RECT 68.555 2.435 68.705 2.585 ;
      RECT 68.205 1.055 68.355 1.205 ;
      RECT 68.16 2.385 68.31 2.535 ;
      RECT 67.86 1.97 68.01 2.12 ;
      RECT 67.775 3.525 67.925 3.675 ;
      RECT 67.12 2.675 67.27 2.825 ;
      RECT 64.835 6.755 64.985 6.905 ;
      RECT 62.49 6.74 62.64 6.89 ;
      RECT 62.475 2.065 62.625 2.215 ;
      RECT 61.685 2.45 61.835 2.6 ;
      RECT 61.685 6.325 61.835 6.475 ;
      RECT 60.095 2.805 60.245 2.955 ;
      RECT 58.325 2.35 58.475 2.5 ;
      RECT 57.305 3.055 57.455 3.205 ;
      RECT 57.075 2.475 57.225 2.625 ;
      RECT 57.04 6.71 57.19 6.86 ;
      RECT 56.73 3.075 56.88 3.225 ;
      RECT 56.49 2.095 56.64 2.245 ;
      RECT 56.38 7.165 56.53 7.315 ;
      RECT 56.18 3.425 56.33 3.575 ;
      RECT 56.04 2.03 56.19 2.18 ;
      RECT 55.405 2.115 55.555 2.265 ;
      RECT 55.295 2.755 55.445 2.905 ;
      RECT 54.97 3.315 55.12 3.465 ;
      RECT 54.8 2.305 54.95 2.455 ;
      RECT 54.445 3.32 54.595 3.47 ;
      RECT 54.385 2.535 54.535 2.685 ;
      RECT 54.02 3.525 54.17 3.675 ;
      RECT 53.86 2.36 54.01 2.51 ;
      RECT 53.295 2.435 53.445 2.585 ;
      RECT 52.945 1.055 53.095 1.205 ;
      RECT 52.9 2.385 53.05 2.535 ;
      RECT 52.6 1.97 52.75 2.12 ;
      RECT 52.515 3.525 52.665 3.675 ;
      RECT 51.86 2.675 52.01 2.825 ;
      RECT 49.575 6.755 49.725 6.905 ;
      RECT 47.23 6.74 47.38 6.89 ;
      RECT 47.215 2.065 47.365 2.215 ;
      RECT 46.425 2.45 46.575 2.6 ;
      RECT 46.425 6.325 46.575 6.475 ;
      RECT 44.835 2.805 44.985 2.955 ;
      RECT 43.065 2.35 43.215 2.5 ;
      RECT 42.045 3.055 42.195 3.205 ;
      RECT 41.815 2.475 41.965 2.625 ;
      RECT 41.78 6.715 41.93 6.865 ;
      RECT 41.47 3.075 41.62 3.225 ;
      RECT 41.23 2.095 41.38 2.245 ;
      RECT 41.12 7.165 41.27 7.315 ;
      RECT 40.92 3.425 41.07 3.575 ;
      RECT 40.78 2.03 40.93 2.18 ;
      RECT 40.145 2.115 40.295 2.265 ;
      RECT 40.035 2.755 40.185 2.905 ;
      RECT 39.71 3.315 39.86 3.465 ;
      RECT 39.54 2.305 39.69 2.455 ;
      RECT 39.185 3.32 39.335 3.47 ;
      RECT 39.125 2.535 39.275 2.685 ;
      RECT 38.76 3.525 38.91 3.675 ;
      RECT 38.6 2.36 38.75 2.51 ;
      RECT 38.035 2.435 38.185 2.585 ;
      RECT 37.685 1.055 37.835 1.205 ;
      RECT 37.64 2.385 37.79 2.535 ;
      RECT 37.34 1.97 37.49 2.12 ;
      RECT 37.255 3.525 37.405 3.675 ;
      RECT 36.6 2.675 36.75 2.825 ;
      RECT 34.36 6.76 34.51 6.91 ;
      RECT 31.97 6.74 32.12 6.89 ;
      RECT 31.955 2.065 32.105 2.215 ;
      RECT 31.165 2.45 31.315 2.6 ;
      RECT 31.165 6.325 31.315 6.475 ;
      RECT 29.575 2.805 29.725 2.955 ;
      RECT 27.805 2.35 27.955 2.5 ;
      RECT 26.785 3.055 26.935 3.205 ;
      RECT 26.555 2.475 26.705 2.625 ;
      RECT 26.52 6.71 26.67 6.86 ;
      RECT 26.21 3.075 26.36 3.225 ;
      RECT 25.97 2.095 26.12 2.245 ;
      RECT 25.86 7.165 26.01 7.315 ;
      RECT 25.66 3.425 25.81 3.575 ;
      RECT 25.52 2.03 25.67 2.18 ;
      RECT 24.885 2.115 25.035 2.265 ;
      RECT 24.775 2.755 24.925 2.905 ;
      RECT 24.45 3.315 24.6 3.465 ;
      RECT 24.28 2.305 24.43 2.455 ;
      RECT 23.925 3.32 24.075 3.47 ;
      RECT 23.865 2.535 24.015 2.685 ;
      RECT 23.5 3.525 23.65 3.675 ;
      RECT 23.34 2.36 23.49 2.51 ;
      RECT 22.775 2.435 22.925 2.585 ;
      RECT 22.425 1.055 22.575 1.205 ;
      RECT 22.38 2.385 22.53 2.535 ;
      RECT 22.08 1.97 22.23 2.12 ;
      RECT 21.995 3.525 22.145 3.675 ;
      RECT 21.34 2.675 21.49 2.825 ;
      RECT 19.1 6.755 19.25 6.905 ;
      RECT 16.71 6.74 16.86 6.89 ;
      RECT 16.695 2.065 16.845 2.215 ;
      RECT 15.905 2.45 16.055 2.6 ;
      RECT 15.905 6.325 16.055 6.475 ;
      RECT 14.315 2.805 14.465 2.955 ;
      RECT 12.545 2.35 12.695 2.5 ;
      RECT 11.525 3.055 11.675 3.205 ;
      RECT 11.295 2.475 11.445 2.625 ;
      RECT 11.26 6.705 11.41 6.855 ;
      RECT 10.95 3.075 11.1 3.225 ;
      RECT 10.71 2.095 10.86 2.245 ;
      RECT 10.6 7.165 10.75 7.315 ;
      RECT 10.4 3.425 10.55 3.575 ;
      RECT 10.26 2.03 10.41 2.18 ;
      RECT 9.625 2.115 9.775 2.265 ;
      RECT 9.515 2.755 9.665 2.905 ;
      RECT 9.19 3.315 9.34 3.465 ;
      RECT 9.02 2.305 9.17 2.455 ;
      RECT 8.665 3.32 8.815 3.47 ;
      RECT 8.605 2.535 8.755 2.685 ;
      RECT 8.24 3.525 8.39 3.675 ;
      RECT 8.08 2.36 8.23 2.51 ;
      RECT 7.515 2.435 7.665 2.585 ;
      RECT 7.165 1.055 7.315 1.205 ;
      RECT 7.12 2.385 7.27 2.535 ;
      RECT 6.82 1.97 6.97 2.12 ;
      RECT 6.735 3.525 6.885 3.675 ;
      RECT 6.08 2.675 6.23 2.825 ;
      RECT 3.105 7.095 3.255 7.245 ;
      RECT 2.73 6.355 2.88 6.505 ;
    LAYER met1 ;
      RECT 66.08 0 74.82 1.74 ;
      RECT 50.82 0 59.56 1.74 ;
      RECT 35.56 0 44.3 1.74 ;
      RECT 20.3 0 29.04 1.74 ;
      RECT 5.04 0 13.78 1.74 ;
      RECT 80.41 0 80.59 0.305 ;
      RECT 65.15 0 78.46 0.305 ;
      RECT 49.89 0 63.2 0.305 ;
      RECT 34.63 0 47.94 0.305 ;
      RECT 19.37 0 32.68 0.305 ;
      RECT 1.495 0 17.42 0.305 ;
      RECT 1.495 0 80.59 0.3 ;
      RECT 1.495 8.58 80.59 8.88 ;
      RECT 80.41 8.575 80.59 8.88 ;
      RECT 65.15 8.575 78.46 8.88 ;
      RECT 49.89 8.575 63.2 8.88 ;
      RECT 34.63 8.575 47.94 8.88 ;
      RECT 19.37 8.575 32.68 8.88 ;
      RECT 1.495 8.575 17.42 8.88 ;
      RECT 71.025 6.315 71.195 8.88 ;
      RECT 55.765 6.315 55.935 8.88 ;
      RECT 40.505 6.315 40.675 8.88 ;
      RECT 25.245 6.315 25.415 8.88 ;
      RECT 9.985 6.315 10.155 8.88 ;
      RECT 71.195 6.285 71.485 6.515 ;
      RECT 55.935 6.285 56.225 6.515 ;
      RECT 40.675 6.285 40.965 6.515 ;
      RECT 25.415 6.285 25.705 6.515 ;
      RECT 10.155 6.285 10.445 6.515 ;
      RECT 79.985 7.77 80.275 8 ;
      RECT 80.045 6.29 80.215 8 ;
      RECT 80.02 7.275 80.37 7.625 ;
      RECT 79.985 6.29 80.275 6.52 ;
      RECT 79.58 2.395 79.685 2.965 ;
      RECT 79.58 2.73 79.905 2.96 ;
      RECT 79.58 2.76 80.075 2.93 ;
      RECT 79.58 2.395 79.77 2.96 ;
      RECT 78.995 2.36 79.285 2.59 ;
      RECT 78.995 2.395 79.77 2.565 ;
      RECT 79.055 0.88 79.225 2.59 ;
      RECT 78.995 0.88 79.285 1.11 ;
      RECT 78.995 7.77 79.285 8 ;
      RECT 79.055 6.29 79.225 8 ;
      RECT 78.995 6.29 79.285 6.52 ;
      RECT 78.995 6.325 79.85 6.485 ;
      RECT 79.68 5.92 79.85 6.485 ;
      RECT 78.995 6.32 79.39 6.485 ;
      RECT 79.615 5.92 79.905 6.15 ;
      RECT 79.615 5.95 80.075 6.12 ;
      RECT 78.625 2.73 78.915 2.96 ;
      RECT 78.625 2.76 79.085 2.93 ;
      RECT 78.69 1.655 78.855 2.96 ;
      RECT 77.205 1.625 77.495 1.855 ;
      RECT 77.205 1.655 78.855 1.825 ;
      RECT 77.265 0.885 77.435 1.855 ;
      RECT 77.205 0.885 77.495 1.115 ;
      RECT 77.205 7.765 77.495 7.995 ;
      RECT 77.265 7.025 77.435 7.995 ;
      RECT 77.265 7.12 78.855 7.29 ;
      RECT 78.685 5.92 78.855 7.29 ;
      RECT 77.205 7.025 77.495 7.255 ;
      RECT 78.625 5.92 78.915 6.15 ;
      RECT 78.625 5.95 79.085 6.12 ;
      RECT 75.255 2.705 75.595 3.055 ;
      RECT 75.345 2.025 75.515 3.055 ;
      RECT 77.635 1.965 77.985 2.315 ;
      RECT 75.345 2.025 77.985 2.195 ;
      RECT 77.66 6.655 77.985 6.98 ;
      RECT 72.2 6.61 72.55 6.96 ;
      RECT 77.635 6.655 77.985 6.885 ;
      RECT 72 6.655 72.55 6.885 ;
      RECT 71.83 6.685 77.985 6.855 ;
      RECT 76.86 2.365 77.18 2.685 ;
      RECT 76.83 2.365 77.18 2.595 ;
      RECT 76.66 2.395 77.18 2.565 ;
      RECT 76.86 6.255 77.18 6.545 ;
      RECT 76.83 6.285 77.18 6.515 ;
      RECT 76.66 6.315 77.18 6.485 ;
      RECT 72.55 2.985 72.7 3.26 ;
      RECT 73.09 2.065 73.095 2.285 ;
      RECT 74.24 2.265 74.255 2.463 ;
      RECT 74.205 2.257 74.24 2.47 ;
      RECT 74.175 2.25 74.205 2.47 ;
      RECT 74.12 2.215 74.175 2.47 ;
      RECT 74.055 2.152 74.12 2.47 ;
      RECT 74.05 2.117 74.055 2.468 ;
      RECT 74.045 2.112 74.05 2.46 ;
      RECT 74.04 2.107 74.045 2.446 ;
      RECT 74.035 2.104 74.04 2.439 ;
      RECT 73.99 2.094 74.035 2.39 ;
      RECT 73.97 2.081 73.99 2.325 ;
      RECT 73.965 2.076 73.97 2.298 ;
      RECT 73.96 2.075 73.965 2.291 ;
      RECT 73.955 2.074 73.96 2.284 ;
      RECT 73.87 2.059 73.955 2.23 ;
      RECT 73.84 2.04 73.87 2.18 ;
      RECT 73.76 2.023 73.84 2.165 ;
      RECT 73.725 2.01 73.76 2.15 ;
      RECT 73.717 2.01 73.725 2.145 ;
      RECT 73.631 2.011 73.717 2.145 ;
      RECT 73.545 2.013 73.631 2.145 ;
      RECT 73.52 2.014 73.545 2.149 ;
      RECT 73.445 2.02 73.52 2.164 ;
      RECT 73.362 2.032 73.445 2.188 ;
      RECT 73.276 2.045 73.362 2.214 ;
      RECT 73.19 2.058 73.276 2.24 ;
      RECT 73.155 2.067 73.19 2.259 ;
      RECT 73.105 2.067 73.155 2.272 ;
      RECT 73.095 2.065 73.105 2.283 ;
      RECT 73.08 2.062 73.09 2.285 ;
      RECT 73.065 2.054 73.08 2.293 ;
      RECT 73.05 2.046 73.065 2.313 ;
      RECT 73.045 2.041 73.05 2.37 ;
      RECT 73.03 2.036 73.045 2.443 ;
      RECT 73.025 2.031 73.03 2.485 ;
      RECT 73.02 2.029 73.025 2.513 ;
      RECT 73.015 2.027 73.02 2.535 ;
      RECT 73.005 2.023 73.015 2.578 ;
      RECT 73 2.02 73.005 2.603 ;
      RECT 72.995 2.018 73 2.623 ;
      RECT 72.99 2.016 72.995 2.647 ;
      RECT 72.985 2.012 72.99 2.67 ;
      RECT 72.98 2.008 72.985 2.693 ;
      RECT 72.945 1.998 72.98 2.8 ;
      RECT 72.94 1.988 72.945 2.898 ;
      RECT 72.935 1.986 72.94 2.925 ;
      RECT 72.93 1.985 72.935 2.945 ;
      RECT 72.925 1.977 72.93 2.965 ;
      RECT 72.92 1.972 72.925 3 ;
      RECT 72.915 1.97 72.92 3.018 ;
      RECT 72.91 1.97 72.915 3.043 ;
      RECT 72.905 1.97 72.91 3.065 ;
      RECT 72.87 1.97 72.905 3.108 ;
      RECT 72.845 1.97 72.87 3.137 ;
      RECT 72.835 1.97 72.845 2.323 ;
      RECT 72.838 2.38 72.845 3.147 ;
      RECT 72.835 2.437 72.838 3.15 ;
      RECT 72.83 1.97 72.835 2.295 ;
      RECT 72.83 2.487 72.835 3.153 ;
      RECT 72.82 1.97 72.83 2.285 ;
      RECT 72.825 2.54 72.83 3.156 ;
      RECT 72.82 2.625 72.825 3.16 ;
      RECT 72.81 1.97 72.82 2.273 ;
      RECT 72.815 2.672 72.82 3.164 ;
      RECT 72.81 2.747 72.815 3.168 ;
      RECT 72.775 1.97 72.81 2.248 ;
      RECT 72.8 2.83 72.81 3.173 ;
      RECT 72.79 2.897 72.8 3.18 ;
      RECT 72.785 2.925 72.79 3.185 ;
      RECT 72.775 2.938 72.785 3.191 ;
      RECT 72.73 1.97 72.775 2.205 ;
      RECT 72.77 2.943 72.775 3.198 ;
      RECT 72.73 2.96 72.77 3.26 ;
      RECT 72.725 1.972 72.73 2.178 ;
      RECT 72.7 2.98 72.73 3.26 ;
      RECT 72.72 1.977 72.725 2.15 ;
      RECT 72.51 2.989 72.55 3.26 ;
      RECT 72.485 2.997 72.51 3.23 ;
      RECT 72.44 3.005 72.485 3.23 ;
      RECT 72.425 3.01 72.44 3.225 ;
      RECT 72.415 3.01 72.425 3.219 ;
      RECT 72.405 3.017 72.415 3.216 ;
      RECT 72.4 3.055 72.405 3.205 ;
      RECT 72.395 3.117 72.4 3.183 ;
      RECT 73.665 2.992 73.85 3.215 ;
      RECT 73.665 3.007 73.855 3.211 ;
      RECT 73.655 2.28 73.74 3.21 ;
      RECT 73.655 3.007 73.86 3.204 ;
      RECT 73.65 3.015 73.86 3.203 ;
      RECT 73.855 2.735 74.175 3.055 ;
      RECT 73.65 2.907 73.82 2.998 ;
      RECT 73.645 2.907 73.82 2.98 ;
      RECT 73.635 2.715 73.77 2.955 ;
      RECT 73.63 2.715 73.77 2.9 ;
      RECT 73.59 2.295 73.76 2.8 ;
      RECT 73.575 2.295 73.76 2.67 ;
      RECT 73.57 2.295 73.76 2.623 ;
      RECT 73.565 2.295 73.76 2.603 ;
      RECT 73.56 2.295 73.76 2.578 ;
      RECT 73.53 2.295 73.79 2.555 ;
      RECT 73.54 2.292 73.75 2.555 ;
      RECT 73.665 2.287 73.75 3.215 ;
      RECT 73.55 2.28 73.74 2.555 ;
      RECT 73.545 2.285 73.74 2.555 ;
      RECT 72.375 2.497 72.56 2.71 ;
      RECT 72.375 2.505 72.57 2.703 ;
      RECT 72.355 2.505 72.57 2.7 ;
      RECT 72.35 2.505 72.57 2.685 ;
      RECT 72.28 2.42 72.54 2.68 ;
      RECT 72.28 2.565 72.575 2.593 ;
      RECT 71.935 3.02 72.195 3.28 ;
      RECT 71.96 2.965 72.155 3.28 ;
      RECT 71.955 2.714 72.135 3.008 ;
      RECT 71.955 2.72 72.145 3.008 ;
      RECT 71.935 2.722 72.145 2.953 ;
      RECT 71.93 2.732 72.145 2.82 ;
      RECT 71.96 2.712 72.135 3.28 ;
      RECT 72.046 2.71 72.135 3.28 ;
      RECT 71.905 1.93 71.94 2.3 ;
      RECT 71.695 2.04 71.7 2.3 ;
      RECT 71.94 1.937 71.955 2.3 ;
      RECT 71.83 1.93 71.905 2.378 ;
      RECT 71.82 1.93 71.83 2.463 ;
      RECT 71.795 1.93 71.82 2.498 ;
      RECT 71.755 1.93 71.795 2.566 ;
      RECT 71.745 1.937 71.755 2.618 ;
      RECT 71.715 2.04 71.745 2.659 ;
      RECT 71.71 2.04 71.715 2.698 ;
      RECT 71.7 2.04 71.71 2.718 ;
      RECT 71.695 2.335 71.7 2.755 ;
      RECT 71.69 2.352 71.695 2.775 ;
      RECT 71.675 2.415 71.69 2.815 ;
      RECT 71.67 2.458 71.675 2.85 ;
      RECT 71.665 2.466 71.67 2.863 ;
      RECT 71.655 2.48 71.665 2.885 ;
      RECT 71.63 2.515 71.655 2.95 ;
      RECT 71.62 2.55 71.63 3.013 ;
      RECT 71.6 2.58 71.62 3.074 ;
      RECT 71.585 2.616 71.6 3.141 ;
      RECT 71.575 2.644 71.585 3.18 ;
      RECT 71.565 2.666 71.575 3.2 ;
      RECT 71.56 2.676 71.565 3.211 ;
      RECT 71.555 2.685 71.56 3.214 ;
      RECT 71.545 2.703 71.555 3.218 ;
      RECT 71.535 2.721 71.545 3.219 ;
      RECT 71.51 2.76 71.535 3.216 ;
      RECT 71.49 2.802 71.51 3.213 ;
      RECT 71.475 2.84 71.49 3.212 ;
      RECT 71.44 2.875 71.475 3.209 ;
      RECT 71.435 2.897 71.44 3.207 ;
      RECT 71.37 2.937 71.435 3.204 ;
      RECT 71.365 2.977 71.37 3.2 ;
      RECT 71.35 2.987 71.365 3.191 ;
      RECT 71.34 3.107 71.35 3.176 ;
      RECT 71.82 3.52 71.83 3.78 ;
      RECT 71.82 3.523 71.84 3.779 ;
      RECT 71.81 3.513 71.82 3.778 ;
      RECT 71.8 3.528 71.88 3.774 ;
      RECT 71.785 3.507 71.8 3.772 ;
      RECT 71.76 3.532 71.885 3.768 ;
      RECT 71.745 3.492 71.76 3.763 ;
      RECT 71.745 3.534 71.895 3.762 ;
      RECT 71.745 3.542 71.91 3.755 ;
      RECT 71.685 3.479 71.745 3.745 ;
      RECT 71.675 3.466 71.685 3.727 ;
      RECT 71.65 3.456 71.675 3.717 ;
      RECT 71.645 3.446 71.65 3.709 ;
      RECT 71.58 3.542 71.91 3.691 ;
      RECT 71.495 3.542 71.91 3.653 ;
      RECT 71.385 3.37 71.645 3.63 ;
      RECT 71.76 3.5 71.785 3.768 ;
      RECT 71.8 3.51 71.81 3.774 ;
      RECT 71.385 3.518 71.825 3.63 ;
      RECT 71.57 7.765 71.86 7.995 ;
      RECT 71.63 7.025 71.8 7.995 ;
      RECT 71.53 7.055 71.9 7.425 ;
      RECT 71.57 7.025 71.86 7.425 ;
      RECT 70.6 3.275 70.63 3.575 ;
      RECT 70.375 3.26 70.38 3.535 ;
      RECT 70.175 3.26 70.33 3.52 ;
      RECT 71.475 1.975 71.505 2.235 ;
      RECT 71.465 1.975 71.475 2.343 ;
      RECT 71.445 1.975 71.465 2.353 ;
      RECT 71.43 1.975 71.445 2.365 ;
      RECT 71.375 1.975 71.43 2.415 ;
      RECT 71.36 1.975 71.375 2.463 ;
      RECT 71.33 1.975 71.36 2.498 ;
      RECT 71.275 1.975 71.33 2.56 ;
      RECT 71.255 1.975 71.275 2.628 ;
      RECT 71.25 1.975 71.255 2.658 ;
      RECT 71.245 1.975 71.25 2.67 ;
      RECT 71.24 2.092 71.245 2.688 ;
      RECT 71.22 2.11 71.24 2.713 ;
      RECT 71.2 2.137 71.22 2.763 ;
      RECT 71.195 2.157 71.2 2.794 ;
      RECT 71.19 2.165 71.195 2.811 ;
      RECT 71.175 2.191 71.19 2.84 ;
      RECT 71.16 2.233 71.175 2.875 ;
      RECT 71.155 2.262 71.16 2.898 ;
      RECT 71.15 2.277 71.155 2.911 ;
      RECT 71.145 2.3 71.15 2.922 ;
      RECT 71.135 2.32 71.145 2.94 ;
      RECT 71.125 2.35 71.135 2.963 ;
      RECT 71.12 2.372 71.125 2.983 ;
      RECT 71.115 2.387 71.12 2.998 ;
      RECT 71.1 2.417 71.115 3.025 ;
      RECT 71.095 2.447 71.1 3.051 ;
      RECT 71.09 2.465 71.095 3.063 ;
      RECT 71.08 2.495 71.09 3.082 ;
      RECT 71.07 2.52 71.08 3.107 ;
      RECT 71.065 2.54 71.07 3.126 ;
      RECT 71.06 2.557 71.065 3.139 ;
      RECT 71.05 2.583 71.06 3.158 ;
      RECT 71.04 2.621 71.05 3.185 ;
      RECT 71.035 2.647 71.04 3.205 ;
      RECT 71.03 2.657 71.035 3.215 ;
      RECT 71.025 2.67 71.03 3.23 ;
      RECT 71.02 2.685 71.025 3.24 ;
      RECT 71.015 2.707 71.02 3.255 ;
      RECT 71.01 2.725 71.015 3.266 ;
      RECT 71.005 2.735 71.01 3.277 ;
      RECT 71 2.743 71.005 3.289 ;
      RECT 70.995 2.751 71 3.3 ;
      RECT 70.99 2.777 70.995 3.313 ;
      RECT 70.98 2.805 70.99 3.326 ;
      RECT 70.975 2.835 70.98 3.335 ;
      RECT 70.97 2.85 70.975 3.342 ;
      RECT 70.955 2.875 70.97 3.349 ;
      RECT 70.95 2.897 70.955 3.355 ;
      RECT 70.945 2.922 70.95 3.358 ;
      RECT 70.936 2.95 70.945 3.362 ;
      RECT 70.93 2.967 70.936 3.367 ;
      RECT 70.925 2.985 70.93 3.371 ;
      RECT 70.92 2.997 70.925 3.374 ;
      RECT 70.915 3.018 70.92 3.378 ;
      RECT 70.91 3.036 70.915 3.381 ;
      RECT 70.905 3.05 70.91 3.384 ;
      RECT 70.9 3.067 70.905 3.387 ;
      RECT 70.895 3.08 70.9 3.39 ;
      RECT 70.87 3.117 70.895 3.398 ;
      RECT 70.865 3.162 70.87 3.407 ;
      RECT 70.86 3.19 70.865 3.41 ;
      RECT 70.85 3.21 70.86 3.414 ;
      RECT 70.845 3.23 70.85 3.419 ;
      RECT 70.84 3.245 70.845 3.422 ;
      RECT 70.82 3.255 70.84 3.429 ;
      RECT 70.755 3.262 70.82 3.455 ;
      RECT 70.72 3.265 70.755 3.483 ;
      RECT 70.705 3.268 70.72 3.498 ;
      RECT 70.695 3.269 70.705 3.513 ;
      RECT 70.685 3.27 70.695 3.53 ;
      RECT 70.68 3.27 70.685 3.545 ;
      RECT 70.675 3.27 70.68 3.553 ;
      RECT 70.66 3.271 70.675 3.568 ;
      RECT 70.63 3.273 70.66 3.575 ;
      RECT 70.52 3.28 70.6 3.575 ;
      RECT 70.475 3.285 70.52 3.575 ;
      RECT 70.465 3.286 70.475 3.565 ;
      RECT 70.455 3.287 70.465 3.558 ;
      RECT 70.435 3.289 70.455 3.553 ;
      RECT 70.425 3.26 70.435 3.548 ;
      RECT 70.38 3.26 70.425 3.54 ;
      RECT 70.35 3.26 70.375 3.53 ;
      RECT 70.33 3.26 70.35 3.523 ;
      RECT 70.61 2.06 70.87 2.32 ;
      RECT 70.49 2.075 70.5 2.24 ;
      RECT 70.475 2.075 70.48 2.235 ;
      RECT 67.84 1.915 68.025 2.205 ;
      RECT 69.655 2.04 69.67 2.195 ;
      RECT 67.805 1.915 67.83 2.175 ;
      RECT 70.22 1.965 70.225 2.107 ;
      RECT 70.135 1.96 70.16 2.1 ;
      RECT 70.535 2.077 70.61 2.27 ;
      RECT 70.52 2.075 70.535 2.253 ;
      RECT 70.5 2.075 70.52 2.245 ;
      RECT 70.48 2.075 70.49 2.238 ;
      RECT 70.435 2.07 70.475 2.228 ;
      RECT 70.395 2.045 70.435 2.213 ;
      RECT 70.38 2.02 70.395 2.203 ;
      RECT 70.375 2.014 70.38 2.201 ;
      RECT 70.34 2.006 70.375 2.184 ;
      RECT 70.335 1.999 70.34 2.172 ;
      RECT 70.315 1.994 70.335 2.16 ;
      RECT 70.305 1.988 70.315 2.145 ;
      RECT 70.285 1.983 70.305 2.13 ;
      RECT 70.275 1.978 70.285 2.123 ;
      RECT 70.27 1.976 70.275 2.118 ;
      RECT 70.265 1.975 70.27 2.115 ;
      RECT 70.225 1.97 70.265 2.111 ;
      RECT 70.205 1.964 70.22 2.106 ;
      RECT 70.17 1.961 70.205 2.103 ;
      RECT 70.16 1.96 70.17 2.101 ;
      RECT 70.1 1.96 70.135 2.098 ;
      RECT 70.055 1.96 70.1 2.098 ;
      RECT 70.005 1.96 70.055 2.101 ;
      RECT 69.99 1.962 70.005 2.103 ;
      RECT 69.975 1.965 69.99 2.104 ;
      RECT 69.965 1.97 69.975 2.105 ;
      RECT 69.935 1.975 69.965 2.11 ;
      RECT 69.925 1.981 69.935 2.118 ;
      RECT 69.915 1.983 69.925 2.122 ;
      RECT 69.905 1.987 69.915 2.126 ;
      RECT 69.88 1.993 69.905 2.134 ;
      RECT 69.87 1.998 69.88 2.142 ;
      RECT 69.855 2.002 69.87 2.146 ;
      RECT 69.82 2.008 69.855 2.154 ;
      RECT 69.8 2.013 69.82 2.164 ;
      RECT 69.77 2.02 69.8 2.173 ;
      RECT 69.725 2.029 69.77 2.187 ;
      RECT 69.72 2.034 69.725 2.198 ;
      RECT 69.7 2.037 69.72 2.199 ;
      RECT 69.67 2.04 69.7 2.197 ;
      RECT 69.635 2.04 69.655 2.193 ;
      RECT 69.565 2.04 69.635 2.184 ;
      RECT 69.55 2.037 69.565 2.176 ;
      RECT 69.51 2.03 69.55 2.171 ;
      RECT 69.485 2.02 69.51 2.164 ;
      RECT 69.48 2.014 69.485 2.161 ;
      RECT 69.44 2.008 69.48 2.158 ;
      RECT 69.425 2.001 69.44 2.153 ;
      RECT 69.405 1.997 69.425 2.148 ;
      RECT 69.39 1.992 69.405 2.144 ;
      RECT 69.375 1.987 69.39 2.142 ;
      RECT 69.36 1.983 69.375 2.141 ;
      RECT 69.345 1.981 69.36 2.137 ;
      RECT 69.335 1.979 69.345 2.132 ;
      RECT 69.32 1.976 69.335 2.128 ;
      RECT 69.31 1.974 69.32 2.123 ;
      RECT 69.29 1.971 69.31 2.119 ;
      RECT 69.245 1.97 69.29 2.117 ;
      RECT 69.185 1.972 69.245 2.118 ;
      RECT 69.165 1.974 69.185 2.12 ;
      RECT 69.135 1.977 69.165 2.121 ;
      RECT 69.085 1.982 69.135 2.123 ;
      RECT 69.08 1.985 69.085 2.125 ;
      RECT 69.07 1.987 69.08 2.128 ;
      RECT 69.065 1.989 69.07 2.131 ;
      RECT 69.015 1.992 69.065 2.138 ;
      RECT 68.995 1.996 69.015 2.15 ;
      RECT 68.985 1.999 68.995 2.156 ;
      RECT 68.975 2 68.985 2.159 ;
      RECT 68.936 2.003 68.975 2.161 ;
      RECT 68.85 2.01 68.936 2.164 ;
      RECT 68.776 2.02 68.85 2.168 ;
      RECT 68.69 2.031 68.776 2.173 ;
      RECT 68.675 2.038 68.69 2.175 ;
      RECT 68.62 2.042 68.675 2.176 ;
      RECT 68.606 2.045 68.62 2.178 ;
      RECT 68.52 2.045 68.606 2.18 ;
      RECT 68.48 2.042 68.52 2.183 ;
      RECT 68.456 2.038 68.48 2.185 ;
      RECT 68.37 2.028 68.456 2.188 ;
      RECT 68.34 2.017 68.37 2.189 ;
      RECT 68.321 2.013 68.34 2.188 ;
      RECT 68.235 2.006 68.321 2.185 ;
      RECT 68.175 1.995 68.235 2.182 ;
      RECT 68.155 1.987 68.175 2.18 ;
      RECT 68.12 1.982 68.155 2.179 ;
      RECT 68.095 1.977 68.12 2.178 ;
      RECT 68.065 1.972 68.095 2.177 ;
      RECT 68.04 1.915 68.065 2.176 ;
      RECT 68.025 1.915 68.04 2.2 ;
      RECT 67.83 1.915 67.84 2.2 ;
      RECT 69.605 2.935 69.61 3.075 ;
      RECT 69.265 2.935 69.3 3.073 ;
      RECT 68.84 2.92 68.855 3.065 ;
      RECT 70.67 2.7 70.76 2.96 ;
      RECT 70.5 2.565 70.6 2.96 ;
      RECT 67.535 2.54 67.615 2.75 ;
      RECT 70.625 2.677 70.67 2.96 ;
      RECT 70.615 2.647 70.625 2.96 ;
      RECT 70.6 2.57 70.615 2.96 ;
      RECT 70.415 2.565 70.5 2.925 ;
      RECT 70.41 2.567 70.415 2.92 ;
      RECT 70.405 2.572 70.41 2.92 ;
      RECT 70.37 2.672 70.405 2.92 ;
      RECT 70.36 2.7 70.37 2.92 ;
      RECT 70.35 2.715 70.36 2.92 ;
      RECT 70.34 2.727 70.35 2.92 ;
      RECT 70.335 2.737 70.34 2.92 ;
      RECT 70.32 2.747 70.335 2.922 ;
      RECT 70.315 2.762 70.32 2.924 ;
      RECT 70.3 2.775 70.315 2.926 ;
      RECT 70.295 2.79 70.3 2.929 ;
      RECT 70.275 2.8 70.295 2.933 ;
      RECT 70.26 2.81 70.275 2.936 ;
      RECT 70.225 2.817 70.26 2.941 ;
      RECT 70.181 2.824 70.225 2.949 ;
      RECT 70.095 2.836 70.181 2.962 ;
      RECT 70.07 2.847 70.095 2.973 ;
      RECT 70.04 2.852 70.07 2.978 ;
      RECT 70.005 2.857 70.04 2.986 ;
      RECT 69.975 2.862 70.005 2.993 ;
      RECT 69.95 2.867 69.975 2.998 ;
      RECT 69.885 2.874 69.95 3.007 ;
      RECT 69.815 2.887 69.885 3.023 ;
      RECT 69.785 2.897 69.815 3.035 ;
      RECT 69.76 2.902 69.785 3.042 ;
      RECT 69.705 2.909 69.76 3.05 ;
      RECT 69.7 2.916 69.705 3.055 ;
      RECT 69.695 2.918 69.7 3.056 ;
      RECT 69.68 2.92 69.695 3.058 ;
      RECT 69.675 2.92 69.68 3.061 ;
      RECT 69.61 2.927 69.675 3.068 ;
      RECT 69.575 2.937 69.605 3.078 ;
      RECT 69.558 2.94 69.575 3.08 ;
      RECT 69.472 2.939 69.558 3.079 ;
      RECT 69.386 2.937 69.472 3.076 ;
      RECT 69.3 2.936 69.386 3.074 ;
      RECT 69.199 2.934 69.265 3.073 ;
      RECT 69.113 2.931 69.199 3.071 ;
      RECT 69.027 2.927 69.113 3.069 ;
      RECT 68.941 2.924 69.027 3.068 ;
      RECT 68.855 2.921 68.941 3.066 ;
      RECT 68.755 2.92 68.84 3.063 ;
      RECT 68.705 2.918 68.755 3.061 ;
      RECT 68.685 2.915 68.705 3.059 ;
      RECT 68.665 2.913 68.685 3.056 ;
      RECT 68.64 2.909 68.665 3.053 ;
      RECT 68.595 2.903 68.64 3.048 ;
      RECT 68.555 2.897 68.595 3.04 ;
      RECT 68.53 2.892 68.555 3.033 ;
      RECT 68.475 2.885 68.53 3.025 ;
      RECT 68.451 2.878 68.475 3.018 ;
      RECT 68.365 2.869 68.451 3.008 ;
      RECT 68.335 2.861 68.365 2.998 ;
      RECT 68.305 2.857 68.335 2.993 ;
      RECT 68.3 2.854 68.305 2.99 ;
      RECT 68.295 2.853 68.3 2.99 ;
      RECT 68.22 2.846 68.295 2.983 ;
      RECT 68.181 2.837 68.22 2.972 ;
      RECT 68.095 2.827 68.181 2.96 ;
      RECT 68.055 2.817 68.095 2.948 ;
      RECT 68.016 2.812 68.055 2.941 ;
      RECT 67.93 2.802 68.016 2.93 ;
      RECT 67.89 2.79 67.93 2.919 ;
      RECT 67.855 2.775 67.89 2.912 ;
      RECT 67.845 2.765 67.855 2.909 ;
      RECT 67.825 2.75 67.845 2.907 ;
      RECT 67.795 2.72 67.825 2.903 ;
      RECT 67.785 2.7 67.795 2.898 ;
      RECT 67.78 2.692 67.785 2.895 ;
      RECT 67.775 2.685 67.78 2.893 ;
      RECT 67.76 2.672 67.775 2.886 ;
      RECT 67.755 2.662 67.76 2.878 ;
      RECT 67.75 2.655 67.755 2.873 ;
      RECT 67.745 2.65 67.75 2.869 ;
      RECT 67.73 2.637 67.745 2.861 ;
      RECT 67.725 2.547 67.73 2.85 ;
      RECT 67.72 2.542 67.725 2.843 ;
      RECT 67.645 2.54 67.72 2.803 ;
      RECT 67.615 2.54 67.645 2.758 ;
      RECT 67.52 2.545 67.535 2.745 ;
      RECT 70.005 2.25 70.265 2.51 ;
      RECT 69.99 2.238 70.17 2.475 ;
      RECT 69.985 2.239 70.17 2.473 ;
      RECT 69.97 2.243 70.18 2.463 ;
      RECT 69.965 2.248 70.185 2.433 ;
      RECT 69.97 2.245 70.185 2.463 ;
      RECT 69.985 2.24 70.18 2.473 ;
      RECT 70.005 2.237 70.17 2.51 ;
      RECT 70.005 2.236 70.16 2.51 ;
      RECT 70.03 2.235 70.16 2.51 ;
      RECT 69.59 2.48 69.85 2.74 ;
      RECT 69.465 2.525 69.85 2.735 ;
      RECT 69.455 2.53 69.85 2.73 ;
      RECT 69.47 3.47 69.485 3.78 ;
      RECT 68.065 3.24 68.075 3.37 ;
      RECT 67.845 3.235 67.95 3.37 ;
      RECT 67.76 3.24 67.81 3.37 ;
      RECT 66.31 1.975 66.315 3.08 ;
      RECT 69.565 3.562 69.57 3.698 ;
      RECT 69.56 3.557 69.565 3.758 ;
      RECT 69.555 3.555 69.56 3.771 ;
      RECT 69.54 3.552 69.555 3.773 ;
      RECT 69.535 3.547 69.54 3.775 ;
      RECT 69.53 3.543 69.535 3.778 ;
      RECT 69.515 3.538 69.53 3.78 ;
      RECT 69.485 3.53 69.515 3.78 ;
      RECT 69.446 3.47 69.47 3.78 ;
      RECT 69.36 3.47 69.446 3.777 ;
      RECT 69.33 3.47 69.36 3.77 ;
      RECT 69.305 3.47 69.33 3.763 ;
      RECT 69.28 3.47 69.305 3.755 ;
      RECT 69.265 3.47 69.28 3.748 ;
      RECT 69.24 3.47 69.265 3.74 ;
      RECT 69.225 3.47 69.24 3.733 ;
      RECT 69.185 3.48 69.225 3.722 ;
      RECT 69.175 3.475 69.185 3.712 ;
      RECT 69.171 3.474 69.175 3.709 ;
      RECT 69.085 3.466 69.171 3.692 ;
      RECT 69.052 3.455 69.085 3.669 ;
      RECT 68.966 3.444 69.052 3.647 ;
      RECT 68.88 3.428 68.966 3.616 ;
      RECT 68.81 3.413 68.88 3.588 ;
      RECT 68.8 3.406 68.81 3.575 ;
      RECT 68.77 3.403 68.8 3.565 ;
      RECT 68.745 3.399 68.77 3.558 ;
      RECT 68.73 3.396 68.745 3.553 ;
      RECT 68.725 3.395 68.73 3.548 ;
      RECT 68.695 3.39 68.725 3.541 ;
      RECT 68.69 3.385 68.695 3.536 ;
      RECT 68.675 3.382 68.69 3.531 ;
      RECT 68.67 3.377 68.675 3.526 ;
      RECT 68.65 3.372 68.67 3.523 ;
      RECT 68.635 3.367 68.65 3.515 ;
      RECT 68.62 3.361 68.635 3.51 ;
      RECT 68.59 3.352 68.62 3.503 ;
      RECT 68.585 3.345 68.59 3.495 ;
      RECT 68.58 3.343 68.585 3.493 ;
      RECT 68.575 3.342 68.58 3.49 ;
      RECT 68.535 3.335 68.575 3.483 ;
      RECT 68.521 3.325 68.535 3.473 ;
      RECT 68.47 3.314 68.521 3.461 ;
      RECT 68.445 3.3 68.47 3.447 ;
      RECT 68.42 3.289 68.445 3.439 ;
      RECT 68.4 3.278 68.42 3.433 ;
      RECT 68.39 3.272 68.4 3.428 ;
      RECT 68.385 3.27 68.39 3.424 ;
      RECT 68.365 3.265 68.385 3.419 ;
      RECT 68.335 3.255 68.365 3.409 ;
      RECT 68.33 3.247 68.335 3.402 ;
      RECT 68.315 3.245 68.33 3.398 ;
      RECT 68.295 3.245 68.315 3.393 ;
      RECT 68.29 3.244 68.295 3.391 ;
      RECT 68.285 3.244 68.29 3.388 ;
      RECT 68.245 3.243 68.285 3.383 ;
      RECT 68.22 3.242 68.245 3.378 ;
      RECT 68.16 3.241 68.22 3.375 ;
      RECT 68.075 3.24 68.16 3.373 ;
      RECT 68.036 3.239 68.065 3.37 ;
      RECT 67.95 3.237 68.036 3.37 ;
      RECT 67.81 3.237 67.845 3.37 ;
      RECT 67.72 3.241 67.76 3.373 ;
      RECT 67.705 3.244 67.72 3.38 ;
      RECT 67.695 3.245 67.705 3.387 ;
      RECT 67.67 3.248 67.695 3.392 ;
      RECT 67.665 3.25 67.67 3.395 ;
      RECT 67.615 3.252 67.665 3.396 ;
      RECT 67.576 3.256 67.615 3.398 ;
      RECT 67.49 3.258 67.576 3.401 ;
      RECT 67.472 3.26 67.49 3.403 ;
      RECT 67.386 3.263 67.472 3.405 ;
      RECT 67.3 3.267 67.386 3.408 ;
      RECT 67.263 3.271 67.3 3.411 ;
      RECT 67.177 3.274 67.263 3.414 ;
      RECT 67.091 3.278 67.177 3.417 ;
      RECT 67.005 3.283 67.091 3.421 ;
      RECT 66.985 3.285 67.005 3.424 ;
      RECT 66.965 3.284 66.985 3.425 ;
      RECT 66.916 3.281 66.965 3.426 ;
      RECT 66.83 3.276 66.916 3.429 ;
      RECT 66.78 3.271 66.83 3.431 ;
      RECT 66.756 3.269 66.78 3.432 ;
      RECT 66.67 3.264 66.756 3.434 ;
      RECT 66.645 3.26 66.67 3.433 ;
      RECT 66.635 3.257 66.645 3.431 ;
      RECT 66.625 3.25 66.635 3.428 ;
      RECT 66.62 3.23 66.625 3.423 ;
      RECT 66.61 3.2 66.62 3.418 ;
      RECT 66.595 3.07 66.61 3.409 ;
      RECT 66.59 3.062 66.595 3.402 ;
      RECT 66.57 3.055 66.59 3.394 ;
      RECT 66.565 3.037 66.57 3.386 ;
      RECT 66.555 3.017 66.565 3.381 ;
      RECT 66.55 2.99 66.555 3.377 ;
      RECT 66.545 2.967 66.55 3.374 ;
      RECT 66.525 2.925 66.545 3.366 ;
      RECT 66.49 2.84 66.525 3.35 ;
      RECT 66.485 2.772 66.49 3.338 ;
      RECT 66.47 2.742 66.485 3.332 ;
      RECT 66.465 1.987 66.47 2.233 ;
      RECT 66.455 2.712 66.47 3.323 ;
      RECT 66.46 1.982 66.465 2.265 ;
      RECT 66.455 1.977 66.46 2.308 ;
      RECT 66.45 1.975 66.455 2.343 ;
      RECT 66.435 2.675 66.455 3.313 ;
      RECT 66.445 1.975 66.45 2.38 ;
      RECT 66.43 1.975 66.445 2.478 ;
      RECT 66.43 2.648 66.435 3.306 ;
      RECT 66.425 1.975 66.43 2.553 ;
      RECT 66.425 2.636 66.43 3.303 ;
      RECT 66.42 1.975 66.425 2.585 ;
      RECT 66.42 2.615 66.425 3.3 ;
      RECT 66.415 1.975 66.42 3.297 ;
      RECT 66.38 1.975 66.415 3.283 ;
      RECT 66.365 1.975 66.38 3.265 ;
      RECT 66.345 1.975 66.365 3.255 ;
      RECT 66.32 1.975 66.345 3.238 ;
      RECT 66.315 1.975 66.32 3.188 ;
      RECT 66.305 1.975 66.31 3.018 ;
      RECT 66.3 1.975 66.305 2.925 ;
      RECT 66.295 1.975 66.3 2.838 ;
      RECT 66.29 1.975 66.295 2.77 ;
      RECT 66.285 1.975 66.29 2.713 ;
      RECT 66.275 1.975 66.285 2.608 ;
      RECT 66.27 1.975 66.275 2.48 ;
      RECT 66.265 1.975 66.27 2.398 ;
      RECT 66.26 1.977 66.265 2.315 ;
      RECT 66.255 1.982 66.26 2.248 ;
      RECT 66.25 1.987 66.255 2.175 ;
      RECT 69.065 2.305 69.325 2.565 ;
      RECT 69.085 2.272 69.295 2.565 ;
      RECT 69.085 2.27 69.285 2.565 ;
      RECT 69.095 2.257 69.285 2.565 ;
      RECT 69.095 2.255 69.21 2.565 ;
      RECT 68.57 2.38 68.745 2.66 ;
      RECT 68.565 2.38 68.745 2.658 ;
      RECT 68.565 2.38 68.76 2.655 ;
      RECT 68.555 2.38 68.76 2.653 ;
      RECT 68.5 2.38 68.76 2.64 ;
      RECT 68.5 2.455 68.765 2.618 ;
      RECT 68.045 2.392 68.065 2.635 ;
      RECT 68.045 2.392 68.105 2.634 ;
      RECT 68.04 2.394 68.105 2.633 ;
      RECT 68.04 2.394 68.191 2.632 ;
      RECT 68.04 2.394 68.26 2.631 ;
      RECT 68.04 2.394 68.28 2.623 ;
      RECT 68.02 2.397 68.28 2.621 ;
      RECT 68.005 2.407 68.28 2.606 ;
      RECT 68.005 2.407 68.295 2.605 ;
      RECT 68 2.416 68.295 2.597 ;
      RECT 68 2.416 68.3 2.593 ;
      RECT 68.105 2.33 68.365 2.59 ;
      RECT 67.995 2.418 68.365 2.475 ;
      RECT 68.065 2.385 68.365 2.59 ;
      RECT 68.03 3.578 68.035 3.785 ;
      RECT 67.98 3.572 68.03 3.784 ;
      RECT 67.947 3.586 68.04 3.783 ;
      RECT 67.861 3.586 68.04 3.782 ;
      RECT 67.775 3.586 68.04 3.781 ;
      RECT 67.775 3.685 68.045 3.778 ;
      RECT 67.77 3.685 68.045 3.773 ;
      RECT 67.765 3.685 68.045 3.755 ;
      RECT 67.76 3.685 68.045 3.738 ;
      RECT 67.72 3.47 67.98 3.73 ;
      RECT 67.18 2.62 67.266 3.034 ;
      RECT 67.18 2.62 67.305 3.031 ;
      RECT 67.18 2.62 67.325 3.021 ;
      RECT 67.135 2.62 67.325 3.018 ;
      RECT 67.135 2.772 67.335 3.008 ;
      RECT 67.135 2.793 67.34 3.002 ;
      RECT 67.135 2.811 67.345 2.998 ;
      RECT 67.135 2.831 67.355 2.993 ;
      RECT 67.11 2.831 67.355 2.99 ;
      RECT 67.1 2.831 67.355 2.968 ;
      RECT 67.1 2.847 67.36 2.938 ;
      RECT 67.065 2.62 67.325 2.925 ;
      RECT 67.065 2.859 67.365 2.88 ;
      RECT 64.725 7.77 65.015 8 ;
      RECT 64.785 6.29 64.955 8 ;
      RECT 64.735 6.655 65.085 7.005 ;
      RECT 64.725 6.29 65.015 6.52 ;
      RECT 64.32 2.395 64.425 2.965 ;
      RECT 64.32 2.73 64.645 2.96 ;
      RECT 64.32 2.76 64.815 2.93 ;
      RECT 64.32 2.395 64.51 2.96 ;
      RECT 63.735 2.36 64.025 2.59 ;
      RECT 63.735 2.395 64.51 2.565 ;
      RECT 63.795 0.88 63.965 2.59 ;
      RECT 63.735 0.88 64.025 1.11 ;
      RECT 63.735 7.77 64.025 8 ;
      RECT 63.795 6.29 63.965 8 ;
      RECT 63.735 6.29 64.025 6.52 ;
      RECT 63.735 6.325 64.59 6.485 ;
      RECT 64.42 5.92 64.59 6.485 ;
      RECT 63.735 6.32 64.13 6.485 ;
      RECT 64.355 5.92 64.645 6.15 ;
      RECT 64.355 5.95 64.815 6.12 ;
      RECT 63.365 2.73 63.655 2.96 ;
      RECT 63.365 2.76 63.825 2.93 ;
      RECT 63.43 1.655 63.595 2.96 ;
      RECT 61.945 1.625 62.235 1.855 ;
      RECT 61.945 1.655 63.595 1.825 ;
      RECT 62.005 0.885 62.175 1.855 ;
      RECT 61.945 0.885 62.235 1.115 ;
      RECT 61.945 7.765 62.235 7.995 ;
      RECT 62.005 7.025 62.175 7.995 ;
      RECT 62.005 7.12 63.595 7.29 ;
      RECT 63.425 5.92 63.595 7.29 ;
      RECT 61.945 7.025 62.235 7.255 ;
      RECT 63.365 5.92 63.655 6.15 ;
      RECT 63.365 5.95 63.825 6.12 ;
      RECT 59.995 2.705 60.335 3.055 ;
      RECT 60.085 2.025 60.255 3.055 ;
      RECT 62.375 1.965 62.725 2.315 ;
      RECT 60.085 2.025 62.725 2.195 ;
      RECT 62.4 6.655 62.725 6.98 ;
      RECT 56.94 6.61 57.29 6.96 ;
      RECT 62.375 6.655 62.725 6.885 ;
      RECT 56.74 6.655 57.29 6.885 ;
      RECT 56.57 6.685 62.725 6.855 ;
      RECT 61.6 2.365 61.92 2.685 ;
      RECT 61.57 2.365 61.92 2.595 ;
      RECT 61.4 2.395 61.92 2.565 ;
      RECT 61.6 6.255 61.92 6.545 ;
      RECT 61.57 6.285 61.92 6.515 ;
      RECT 61.4 6.315 61.92 6.485 ;
      RECT 57.29 2.985 57.44 3.26 ;
      RECT 57.83 2.065 57.835 2.285 ;
      RECT 58.98 2.265 58.995 2.463 ;
      RECT 58.945 2.257 58.98 2.47 ;
      RECT 58.915 2.25 58.945 2.47 ;
      RECT 58.86 2.215 58.915 2.47 ;
      RECT 58.795 2.152 58.86 2.47 ;
      RECT 58.79 2.117 58.795 2.468 ;
      RECT 58.785 2.112 58.79 2.46 ;
      RECT 58.78 2.107 58.785 2.446 ;
      RECT 58.775 2.104 58.78 2.439 ;
      RECT 58.73 2.094 58.775 2.39 ;
      RECT 58.71 2.081 58.73 2.325 ;
      RECT 58.705 2.076 58.71 2.298 ;
      RECT 58.7 2.075 58.705 2.291 ;
      RECT 58.695 2.074 58.7 2.284 ;
      RECT 58.61 2.059 58.695 2.23 ;
      RECT 58.58 2.04 58.61 2.18 ;
      RECT 58.5 2.023 58.58 2.165 ;
      RECT 58.465 2.01 58.5 2.15 ;
      RECT 58.457 2.01 58.465 2.145 ;
      RECT 58.371 2.011 58.457 2.145 ;
      RECT 58.285 2.013 58.371 2.145 ;
      RECT 58.26 2.014 58.285 2.149 ;
      RECT 58.185 2.02 58.26 2.164 ;
      RECT 58.102 2.032 58.185 2.188 ;
      RECT 58.016 2.045 58.102 2.214 ;
      RECT 57.93 2.058 58.016 2.24 ;
      RECT 57.895 2.067 57.93 2.259 ;
      RECT 57.845 2.067 57.895 2.272 ;
      RECT 57.835 2.065 57.845 2.283 ;
      RECT 57.82 2.062 57.83 2.285 ;
      RECT 57.805 2.054 57.82 2.293 ;
      RECT 57.79 2.046 57.805 2.313 ;
      RECT 57.785 2.041 57.79 2.37 ;
      RECT 57.77 2.036 57.785 2.443 ;
      RECT 57.765 2.031 57.77 2.485 ;
      RECT 57.76 2.029 57.765 2.513 ;
      RECT 57.755 2.027 57.76 2.535 ;
      RECT 57.745 2.023 57.755 2.578 ;
      RECT 57.74 2.02 57.745 2.603 ;
      RECT 57.735 2.018 57.74 2.623 ;
      RECT 57.73 2.016 57.735 2.647 ;
      RECT 57.725 2.012 57.73 2.67 ;
      RECT 57.72 2.008 57.725 2.693 ;
      RECT 57.685 1.998 57.72 2.8 ;
      RECT 57.68 1.988 57.685 2.898 ;
      RECT 57.675 1.986 57.68 2.925 ;
      RECT 57.67 1.985 57.675 2.945 ;
      RECT 57.665 1.977 57.67 2.965 ;
      RECT 57.66 1.972 57.665 3 ;
      RECT 57.655 1.97 57.66 3.018 ;
      RECT 57.65 1.97 57.655 3.043 ;
      RECT 57.645 1.97 57.65 3.065 ;
      RECT 57.61 1.97 57.645 3.108 ;
      RECT 57.585 1.97 57.61 3.137 ;
      RECT 57.575 1.97 57.585 2.323 ;
      RECT 57.578 2.38 57.585 3.147 ;
      RECT 57.575 2.437 57.578 3.15 ;
      RECT 57.57 1.97 57.575 2.295 ;
      RECT 57.57 2.487 57.575 3.153 ;
      RECT 57.56 1.97 57.57 2.285 ;
      RECT 57.565 2.54 57.57 3.156 ;
      RECT 57.56 2.625 57.565 3.16 ;
      RECT 57.55 1.97 57.56 2.273 ;
      RECT 57.555 2.672 57.56 3.164 ;
      RECT 57.55 2.747 57.555 3.168 ;
      RECT 57.515 1.97 57.55 2.248 ;
      RECT 57.54 2.83 57.55 3.173 ;
      RECT 57.53 2.897 57.54 3.18 ;
      RECT 57.525 2.925 57.53 3.185 ;
      RECT 57.515 2.938 57.525 3.191 ;
      RECT 57.47 1.97 57.515 2.205 ;
      RECT 57.51 2.943 57.515 3.198 ;
      RECT 57.47 2.96 57.51 3.26 ;
      RECT 57.465 1.972 57.47 2.178 ;
      RECT 57.44 2.98 57.47 3.26 ;
      RECT 57.46 1.977 57.465 2.15 ;
      RECT 57.25 2.989 57.29 3.26 ;
      RECT 57.225 2.997 57.25 3.23 ;
      RECT 57.18 3.005 57.225 3.23 ;
      RECT 57.165 3.01 57.18 3.225 ;
      RECT 57.155 3.01 57.165 3.219 ;
      RECT 57.145 3.017 57.155 3.216 ;
      RECT 57.14 3.055 57.145 3.205 ;
      RECT 57.135 3.117 57.14 3.183 ;
      RECT 58.405 2.992 58.59 3.215 ;
      RECT 58.405 3.007 58.595 3.211 ;
      RECT 58.395 2.28 58.48 3.21 ;
      RECT 58.395 3.007 58.6 3.204 ;
      RECT 58.39 3.015 58.6 3.203 ;
      RECT 58.595 2.735 58.915 3.055 ;
      RECT 58.39 2.907 58.56 2.998 ;
      RECT 58.385 2.907 58.56 2.98 ;
      RECT 58.375 2.715 58.51 2.955 ;
      RECT 58.37 2.715 58.51 2.9 ;
      RECT 58.33 2.295 58.5 2.8 ;
      RECT 58.315 2.295 58.5 2.67 ;
      RECT 58.31 2.295 58.5 2.623 ;
      RECT 58.305 2.295 58.5 2.603 ;
      RECT 58.3 2.295 58.5 2.578 ;
      RECT 58.27 2.295 58.53 2.555 ;
      RECT 58.28 2.292 58.49 2.555 ;
      RECT 58.405 2.287 58.49 3.215 ;
      RECT 58.29 2.28 58.48 2.555 ;
      RECT 58.285 2.285 58.48 2.555 ;
      RECT 57.115 2.497 57.3 2.71 ;
      RECT 57.115 2.505 57.31 2.703 ;
      RECT 57.095 2.505 57.31 2.7 ;
      RECT 57.09 2.505 57.31 2.685 ;
      RECT 57.02 2.42 57.28 2.68 ;
      RECT 57.02 2.565 57.315 2.593 ;
      RECT 56.675 3.02 56.935 3.28 ;
      RECT 56.7 2.965 56.895 3.28 ;
      RECT 56.695 2.714 56.875 3.008 ;
      RECT 56.695 2.72 56.885 3.008 ;
      RECT 56.675 2.722 56.885 2.953 ;
      RECT 56.67 2.732 56.885 2.82 ;
      RECT 56.7 2.712 56.875 3.28 ;
      RECT 56.786 2.71 56.875 3.28 ;
      RECT 56.645 1.93 56.68 2.3 ;
      RECT 56.435 2.04 56.44 2.3 ;
      RECT 56.68 1.937 56.695 2.3 ;
      RECT 56.57 1.93 56.645 2.378 ;
      RECT 56.56 1.93 56.57 2.463 ;
      RECT 56.535 1.93 56.56 2.498 ;
      RECT 56.495 1.93 56.535 2.566 ;
      RECT 56.485 1.937 56.495 2.618 ;
      RECT 56.455 2.04 56.485 2.659 ;
      RECT 56.45 2.04 56.455 2.698 ;
      RECT 56.44 2.04 56.45 2.718 ;
      RECT 56.435 2.335 56.44 2.755 ;
      RECT 56.43 2.352 56.435 2.775 ;
      RECT 56.415 2.415 56.43 2.815 ;
      RECT 56.41 2.458 56.415 2.85 ;
      RECT 56.405 2.466 56.41 2.863 ;
      RECT 56.395 2.48 56.405 2.885 ;
      RECT 56.37 2.515 56.395 2.95 ;
      RECT 56.36 2.55 56.37 3.013 ;
      RECT 56.34 2.58 56.36 3.074 ;
      RECT 56.325 2.616 56.34 3.141 ;
      RECT 56.315 2.644 56.325 3.18 ;
      RECT 56.305 2.666 56.315 3.2 ;
      RECT 56.3 2.676 56.305 3.211 ;
      RECT 56.295 2.685 56.3 3.214 ;
      RECT 56.285 2.703 56.295 3.218 ;
      RECT 56.275 2.721 56.285 3.219 ;
      RECT 56.25 2.76 56.275 3.216 ;
      RECT 56.23 2.802 56.25 3.213 ;
      RECT 56.215 2.84 56.23 3.212 ;
      RECT 56.18 2.875 56.215 3.209 ;
      RECT 56.175 2.897 56.18 3.207 ;
      RECT 56.11 2.937 56.175 3.204 ;
      RECT 56.105 2.977 56.11 3.2 ;
      RECT 56.09 2.987 56.105 3.191 ;
      RECT 56.08 3.107 56.09 3.176 ;
      RECT 56.56 3.52 56.57 3.78 ;
      RECT 56.56 3.523 56.58 3.779 ;
      RECT 56.55 3.513 56.56 3.778 ;
      RECT 56.54 3.528 56.62 3.774 ;
      RECT 56.525 3.507 56.54 3.772 ;
      RECT 56.5 3.532 56.625 3.768 ;
      RECT 56.485 3.492 56.5 3.763 ;
      RECT 56.485 3.534 56.635 3.762 ;
      RECT 56.485 3.542 56.65 3.755 ;
      RECT 56.425 3.479 56.485 3.745 ;
      RECT 56.415 3.466 56.425 3.727 ;
      RECT 56.39 3.456 56.415 3.717 ;
      RECT 56.385 3.446 56.39 3.709 ;
      RECT 56.32 3.542 56.65 3.691 ;
      RECT 56.235 3.542 56.65 3.653 ;
      RECT 56.125 3.37 56.385 3.63 ;
      RECT 56.5 3.5 56.525 3.768 ;
      RECT 56.54 3.51 56.55 3.774 ;
      RECT 56.125 3.518 56.565 3.63 ;
      RECT 56.31 7.765 56.6 7.995 ;
      RECT 56.37 7.025 56.54 7.995 ;
      RECT 56.27 7.055 56.64 7.425 ;
      RECT 56.31 7.025 56.6 7.425 ;
      RECT 55.34 3.275 55.37 3.575 ;
      RECT 55.115 3.26 55.12 3.535 ;
      RECT 54.915 3.26 55.07 3.52 ;
      RECT 56.215 1.975 56.245 2.235 ;
      RECT 56.205 1.975 56.215 2.343 ;
      RECT 56.185 1.975 56.205 2.353 ;
      RECT 56.17 1.975 56.185 2.365 ;
      RECT 56.115 1.975 56.17 2.415 ;
      RECT 56.1 1.975 56.115 2.463 ;
      RECT 56.07 1.975 56.1 2.498 ;
      RECT 56.015 1.975 56.07 2.56 ;
      RECT 55.995 1.975 56.015 2.628 ;
      RECT 55.99 1.975 55.995 2.658 ;
      RECT 55.985 1.975 55.99 2.67 ;
      RECT 55.98 2.092 55.985 2.688 ;
      RECT 55.96 2.11 55.98 2.713 ;
      RECT 55.94 2.137 55.96 2.763 ;
      RECT 55.935 2.157 55.94 2.794 ;
      RECT 55.93 2.165 55.935 2.811 ;
      RECT 55.915 2.191 55.93 2.84 ;
      RECT 55.9 2.233 55.915 2.875 ;
      RECT 55.895 2.262 55.9 2.898 ;
      RECT 55.89 2.277 55.895 2.911 ;
      RECT 55.885 2.3 55.89 2.922 ;
      RECT 55.875 2.32 55.885 2.94 ;
      RECT 55.865 2.35 55.875 2.963 ;
      RECT 55.86 2.372 55.865 2.983 ;
      RECT 55.855 2.387 55.86 2.998 ;
      RECT 55.84 2.417 55.855 3.025 ;
      RECT 55.835 2.447 55.84 3.051 ;
      RECT 55.83 2.465 55.835 3.063 ;
      RECT 55.82 2.495 55.83 3.082 ;
      RECT 55.81 2.52 55.82 3.107 ;
      RECT 55.805 2.54 55.81 3.126 ;
      RECT 55.8 2.557 55.805 3.139 ;
      RECT 55.79 2.583 55.8 3.158 ;
      RECT 55.78 2.621 55.79 3.185 ;
      RECT 55.775 2.647 55.78 3.205 ;
      RECT 55.77 2.657 55.775 3.215 ;
      RECT 55.765 2.67 55.77 3.23 ;
      RECT 55.76 2.685 55.765 3.24 ;
      RECT 55.755 2.707 55.76 3.255 ;
      RECT 55.75 2.725 55.755 3.266 ;
      RECT 55.745 2.735 55.75 3.277 ;
      RECT 55.74 2.743 55.745 3.289 ;
      RECT 55.735 2.751 55.74 3.3 ;
      RECT 55.73 2.777 55.735 3.313 ;
      RECT 55.72 2.805 55.73 3.326 ;
      RECT 55.715 2.835 55.72 3.335 ;
      RECT 55.71 2.85 55.715 3.342 ;
      RECT 55.695 2.875 55.71 3.349 ;
      RECT 55.69 2.897 55.695 3.355 ;
      RECT 55.685 2.922 55.69 3.358 ;
      RECT 55.676 2.95 55.685 3.362 ;
      RECT 55.67 2.967 55.676 3.367 ;
      RECT 55.665 2.985 55.67 3.371 ;
      RECT 55.66 2.997 55.665 3.374 ;
      RECT 55.655 3.018 55.66 3.378 ;
      RECT 55.65 3.036 55.655 3.381 ;
      RECT 55.645 3.05 55.65 3.384 ;
      RECT 55.64 3.067 55.645 3.387 ;
      RECT 55.635 3.08 55.64 3.39 ;
      RECT 55.61 3.117 55.635 3.398 ;
      RECT 55.605 3.162 55.61 3.407 ;
      RECT 55.6 3.19 55.605 3.41 ;
      RECT 55.59 3.21 55.6 3.414 ;
      RECT 55.585 3.23 55.59 3.419 ;
      RECT 55.58 3.245 55.585 3.422 ;
      RECT 55.56 3.255 55.58 3.429 ;
      RECT 55.495 3.262 55.56 3.455 ;
      RECT 55.46 3.265 55.495 3.483 ;
      RECT 55.445 3.268 55.46 3.498 ;
      RECT 55.435 3.269 55.445 3.513 ;
      RECT 55.425 3.27 55.435 3.53 ;
      RECT 55.42 3.27 55.425 3.545 ;
      RECT 55.415 3.27 55.42 3.553 ;
      RECT 55.4 3.271 55.415 3.568 ;
      RECT 55.37 3.273 55.4 3.575 ;
      RECT 55.26 3.28 55.34 3.575 ;
      RECT 55.215 3.285 55.26 3.575 ;
      RECT 55.205 3.286 55.215 3.565 ;
      RECT 55.195 3.287 55.205 3.558 ;
      RECT 55.175 3.289 55.195 3.553 ;
      RECT 55.165 3.26 55.175 3.548 ;
      RECT 55.12 3.26 55.165 3.54 ;
      RECT 55.09 3.26 55.115 3.53 ;
      RECT 55.07 3.26 55.09 3.523 ;
      RECT 55.35 2.06 55.61 2.32 ;
      RECT 55.23 2.075 55.24 2.24 ;
      RECT 55.215 2.075 55.22 2.235 ;
      RECT 52.58 1.915 52.765 2.205 ;
      RECT 54.395 2.04 54.41 2.195 ;
      RECT 52.545 1.915 52.57 2.175 ;
      RECT 54.96 1.965 54.965 2.107 ;
      RECT 54.875 1.96 54.9 2.1 ;
      RECT 55.275 2.077 55.35 2.27 ;
      RECT 55.26 2.075 55.275 2.253 ;
      RECT 55.24 2.075 55.26 2.245 ;
      RECT 55.22 2.075 55.23 2.238 ;
      RECT 55.175 2.07 55.215 2.228 ;
      RECT 55.135 2.045 55.175 2.213 ;
      RECT 55.12 2.02 55.135 2.203 ;
      RECT 55.115 2.014 55.12 2.201 ;
      RECT 55.08 2.006 55.115 2.184 ;
      RECT 55.075 1.999 55.08 2.172 ;
      RECT 55.055 1.994 55.075 2.16 ;
      RECT 55.045 1.988 55.055 2.145 ;
      RECT 55.025 1.983 55.045 2.13 ;
      RECT 55.015 1.978 55.025 2.123 ;
      RECT 55.01 1.976 55.015 2.118 ;
      RECT 55.005 1.975 55.01 2.115 ;
      RECT 54.965 1.97 55.005 2.111 ;
      RECT 54.945 1.964 54.96 2.106 ;
      RECT 54.91 1.961 54.945 2.103 ;
      RECT 54.9 1.96 54.91 2.101 ;
      RECT 54.84 1.96 54.875 2.098 ;
      RECT 54.795 1.96 54.84 2.098 ;
      RECT 54.745 1.96 54.795 2.101 ;
      RECT 54.73 1.962 54.745 2.103 ;
      RECT 54.715 1.965 54.73 2.104 ;
      RECT 54.705 1.97 54.715 2.105 ;
      RECT 54.675 1.975 54.705 2.11 ;
      RECT 54.665 1.981 54.675 2.118 ;
      RECT 54.655 1.983 54.665 2.122 ;
      RECT 54.645 1.987 54.655 2.126 ;
      RECT 54.62 1.993 54.645 2.134 ;
      RECT 54.61 1.998 54.62 2.142 ;
      RECT 54.595 2.002 54.61 2.146 ;
      RECT 54.56 2.008 54.595 2.154 ;
      RECT 54.54 2.013 54.56 2.164 ;
      RECT 54.51 2.02 54.54 2.173 ;
      RECT 54.465 2.029 54.51 2.187 ;
      RECT 54.46 2.034 54.465 2.198 ;
      RECT 54.44 2.037 54.46 2.199 ;
      RECT 54.41 2.04 54.44 2.197 ;
      RECT 54.375 2.04 54.395 2.193 ;
      RECT 54.305 2.04 54.375 2.184 ;
      RECT 54.29 2.037 54.305 2.176 ;
      RECT 54.25 2.03 54.29 2.171 ;
      RECT 54.225 2.02 54.25 2.164 ;
      RECT 54.22 2.014 54.225 2.161 ;
      RECT 54.18 2.008 54.22 2.158 ;
      RECT 54.165 2.001 54.18 2.153 ;
      RECT 54.145 1.997 54.165 2.148 ;
      RECT 54.13 1.992 54.145 2.144 ;
      RECT 54.115 1.987 54.13 2.142 ;
      RECT 54.1 1.983 54.115 2.141 ;
      RECT 54.085 1.981 54.1 2.137 ;
      RECT 54.075 1.979 54.085 2.132 ;
      RECT 54.06 1.976 54.075 2.128 ;
      RECT 54.05 1.974 54.06 2.123 ;
      RECT 54.03 1.971 54.05 2.119 ;
      RECT 53.985 1.97 54.03 2.117 ;
      RECT 53.925 1.972 53.985 2.118 ;
      RECT 53.905 1.974 53.925 2.12 ;
      RECT 53.875 1.977 53.905 2.121 ;
      RECT 53.825 1.982 53.875 2.123 ;
      RECT 53.82 1.985 53.825 2.125 ;
      RECT 53.81 1.987 53.82 2.128 ;
      RECT 53.805 1.989 53.81 2.131 ;
      RECT 53.755 1.992 53.805 2.138 ;
      RECT 53.735 1.996 53.755 2.15 ;
      RECT 53.725 1.999 53.735 2.156 ;
      RECT 53.715 2 53.725 2.159 ;
      RECT 53.676 2.003 53.715 2.161 ;
      RECT 53.59 2.01 53.676 2.164 ;
      RECT 53.516 2.02 53.59 2.168 ;
      RECT 53.43 2.031 53.516 2.173 ;
      RECT 53.415 2.038 53.43 2.175 ;
      RECT 53.36 2.042 53.415 2.176 ;
      RECT 53.346 2.045 53.36 2.178 ;
      RECT 53.26 2.045 53.346 2.18 ;
      RECT 53.22 2.042 53.26 2.183 ;
      RECT 53.196 2.038 53.22 2.185 ;
      RECT 53.11 2.028 53.196 2.188 ;
      RECT 53.08 2.017 53.11 2.189 ;
      RECT 53.061 2.013 53.08 2.188 ;
      RECT 52.975 2.006 53.061 2.185 ;
      RECT 52.915 1.995 52.975 2.182 ;
      RECT 52.895 1.987 52.915 2.18 ;
      RECT 52.86 1.982 52.895 2.179 ;
      RECT 52.835 1.977 52.86 2.178 ;
      RECT 52.805 1.972 52.835 2.177 ;
      RECT 52.78 1.915 52.805 2.176 ;
      RECT 52.765 1.915 52.78 2.2 ;
      RECT 52.57 1.915 52.58 2.2 ;
      RECT 54.345 2.935 54.35 3.075 ;
      RECT 54.005 2.935 54.04 3.073 ;
      RECT 53.58 2.92 53.595 3.065 ;
      RECT 55.41 2.7 55.5 2.96 ;
      RECT 55.24 2.565 55.34 2.96 ;
      RECT 52.275 2.54 52.355 2.75 ;
      RECT 55.365 2.677 55.41 2.96 ;
      RECT 55.355 2.647 55.365 2.96 ;
      RECT 55.34 2.57 55.355 2.96 ;
      RECT 55.155 2.565 55.24 2.925 ;
      RECT 55.15 2.567 55.155 2.92 ;
      RECT 55.145 2.572 55.15 2.92 ;
      RECT 55.11 2.672 55.145 2.92 ;
      RECT 55.1 2.7 55.11 2.92 ;
      RECT 55.09 2.715 55.1 2.92 ;
      RECT 55.08 2.727 55.09 2.92 ;
      RECT 55.075 2.737 55.08 2.92 ;
      RECT 55.06 2.747 55.075 2.922 ;
      RECT 55.055 2.762 55.06 2.924 ;
      RECT 55.04 2.775 55.055 2.926 ;
      RECT 55.035 2.79 55.04 2.929 ;
      RECT 55.015 2.8 55.035 2.933 ;
      RECT 55 2.81 55.015 2.936 ;
      RECT 54.965 2.817 55 2.941 ;
      RECT 54.921 2.824 54.965 2.949 ;
      RECT 54.835 2.836 54.921 2.962 ;
      RECT 54.81 2.847 54.835 2.973 ;
      RECT 54.78 2.852 54.81 2.978 ;
      RECT 54.745 2.857 54.78 2.986 ;
      RECT 54.715 2.862 54.745 2.993 ;
      RECT 54.69 2.867 54.715 2.998 ;
      RECT 54.625 2.874 54.69 3.007 ;
      RECT 54.555 2.887 54.625 3.023 ;
      RECT 54.525 2.897 54.555 3.035 ;
      RECT 54.5 2.902 54.525 3.042 ;
      RECT 54.445 2.909 54.5 3.05 ;
      RECT 54.44 2.916 54.445 3.055 ;
      RECT 54.435 2.918 54.44 3.056 ;
      RECT 54.42 2.92 54.435 3.058 ;
      RECT 54.415 2.92 54.42 3.061 ;
      RECT 54.35 2.927 54.415 3.068 ;
      RECT 54.315 2.937 54.345 3.078 ;
      RECT 54.298 2.94 54.315 3.08 ;
      RECT 54.212 2.939 54.298 3.079 ;
      RECT 54.126 2.937 54.212 3.076 ;
      RECT 54.04 2.936 54.126 3.074 ;
      RECT 53.939 2.934 54.005 3.073 ;
      RECT 53.853 2.931 53.939 3.071 ;
      RECT 53.767 2.927 53.853 3.069 ;
      RECT 53.681 2.924 53.767 3.068 ;
      RECT 53.595 2.921 53.681 3.066 ;
      RECT 53.495 2.92 53.58 3.063 ;
      RECT 53.445 2.918 53.495 3.061 ;
      RECT 53.425 2.915 53.445 3.059 ;
      RECT 53.405 2.913 53.425 3.056 ;
      RECT 53.38 2.909 53.405 3.053 ;
      RECT 53.335 2.903 53.38 3.048 ;
      RECT 53.295 2.897 53.335 3.04 ;
      RECT 53.27 2.892 53.295 3.033 ;
      RECT 53.215 2.885 53.27 3.025 ;
      RECT 53.191 2.878 53.215 3.018 ;
      RECT 53.105 2.869 53.191 3.008 ;
      RECT 53.075 2.861 53.105 2.998 ;
      RECT 53.045 2.857 53.075 2.993 ;
      RECT 53.04 2.854 53.045 2.99 ;
      RECT 53.035 2.853 53.04 2.99 ;
      RECT 52.96 2.846 53.035 2.983 ;
      RECT 52.921 2.837 52.96 2.972 ;
      RECT 52.835 2.827 52.921 2.96 ;
      RECT 52.795 2.817 52.835 2.948 ;
      RECT 52.756 2.812 52.795 2.941 ;
      RECT 52.67 2.802 52.756 2.93 ;
      RECT 52.63 2.79 52.67 2.919 ;
      RECT 52.595 2.775 52.63 2.912 ;
      RECT 52.585 2.765 52.595 2.909 ;
      RECT 52.565 2.75 52.585 2.907 ;
      RECT 52.535 2.72 52.565 2.903 ;
      RECT 52.525 2.7 52.535 2.898 ;
      RECT 52.52 2.692 52.525 2.895 ;
      RECT 52.515 2.685 52.52 2.893 ;
      RECT 52.5 2.672 52.515 2.886 ;
      RECT 52.495 2.662 52.5 2.878 ;
      RECT 52.49 2.655 52.495 2.873 ;
      RECT 52.485 2.65 52.49 2.869 ;
      RECT 52.47 2.637 52.485 2.861 ;
      RECT 52.465 2.547 52.47 2.85 ;
      RECT 52.46 2.542 52.465 2.843 ;
      RECT 52.385 2.54 52.46 2.803 ;
      RECT 52.355 2.54 52.385 2.758 ;
      RECT 52.26 2.545 52.275 2.745 ;
      RECT 54.745 2.25 55.005 2.51 ;
      RECT 54.73 2.238 54.91 2.475 ;
      RECT 54.725 2.239 54.91 2.473 ;
      RECT 54.71 2.243 54.92 2.463 ;
      RECT 54.705 2.248 54.925 2.433 ;
      RECT 54.71 2.245 54.925 2.463 ;
      RECT 54.725 2.24 54.92 2.473 ;
      RECT 54.745 2.237 54.91 2.51 ;
      RECT 54.745 2.236 54.9 2.51 ;
      RECT 54.77 2.235 54.9 2.51 ;
      RECT 54.33 2.48 54.59 2.74 ;
      RECT 54.205 2.525 54.59 2.735 ;
      RECT 54.195 2.53 54.59 2.73 ;
      RECT 54.21 3.47 54.225 3.78 ;
      RECT 52.805 3.24 52.815 3.37 ;
      RECT 52.585 3.235 52.69 3.37 ;
      RECT 52.5 3.24 52.55 3.37 ;
      RECT 51.05 1.975 51.055 3.08 ;
      RECT 54.305 3.562 54.31 3.698 ;
      RECT 54.3 3.557 54.305 3.758 ;
      RECT 54.295 3.555 54.3 3.771 ;
      RECT 54.28 3.552 54.295 3.773 ;
      RECT 54.275 3.547 54.28 3.775 ;
      RECT 54.27 3.543 54.275 3.778 ;
      RECT 54.255 3.538 54.27 3.78 ;
      RECT 54.225 3.53 54.255 3.78 ;
      RECT 54.186 3.47 54.21 3.78 ;
      RECT 54.1 3.47 54.186 3.777 ;
      RECT 54.07 3.47 54.1 3.77 ;
      RECT 54.045 3.47 54.07 3.763 ;
      RECT 54.02 3.47 54.045 3.755 ;
      RECT 54.005 3.47 54.02 3.748 ;
      RECT 53.98 3.47 54.005 3.74 ;
      RECT 53.965 3.47 53.98 3.733 ;
      RECT 53.925 3.48 53.965 3.722 ;
      RECT 53.915 3.475 53.925 3.712 ;
      RECT 53.911 3.474 53.915 3.709 ;
      RECT 53.825 3.466 53.911 3.692 ;
      RECT 53.792 3.455 53.825 3.669 ;
      RECT 53.706 3.444 53.792 3.647 ;
      RECT 53.62 3.428 53.706 3.616 ;
      RECT 53.55 3.413 53.62 3.588 ;
      RECT 53.54 3.406 53.55 3.575 ;
      RECT 53.51 3.403 53.54 3.565 ;
      RECT 53.485 3.399 53.51 3.558 ;
      RECT 53.47 3.396 53.485 3.553 ;
      RECT 53.465 3.395 53.47 3.548 ;
      RECT 53.435 3.39 53.465 3.541 ;
      RECT 53.43 3.385 53.435 3.536 ;
      RECT 53.415 3.382 53.43 3.531 ;
      RECT 53.41 3.377 53.415 3.526 ;
      RECT 53.39 3.372 53.41 3.523 ;
      RECT 53.375 3.367 53.39 3.515 ;
      RECT 53.36 3.361 53.375 3.51 ;
      RECT 53.33 3.352 53.36 3.503 ;
      RECT 53.325 3.345 53.33 3.495 ;
      RECT 53.32 3.343 53.325 3.493 ;
      RECT 53.315 3.342 53.32 3.49 ;
      RECT 53.275 3.335 53.315 3.483 ;
      RECT 53.261 3.325 53.275 3.473 ;
      RECT 53.21 3.314 53.261 3.461 ;
      RECT 53.185 3.3 53.21 3.447 ;
      RECT 53.16 3.289 53.185 3.439 ;
      RECT 53.14 3.278 53.16 3.433 ;
      RECT 53.13 3.272 53.14 3.428 ;
      RECT 53.125 3.27 53.13 3.424 ;
      RECT 53.105 3.265 53.125 3.419 ;
      RECT 53.075 3.255 53.105 3.409 ;
      RECT 53.07 3.247 53.075 3.402 ;
      RECT 53.055 3.245 53.07 3.398 ;
      RECT 53.035 3.245 53.055 3.393 ;
      RECT 53.03 3.244 53.035 3.391 ;
      RECT 53.025 3.244 53.03 3.388 ;
      RECT 52.985 3.243 53.025 3.383 ;
      RECT 52.96 3.242 52.985 3.378 ;
      RECT 52.9 3.241 52.96 3.375 ;
      RECT 52.815 3.24 52.9 3.373 ;
      RECT 52.776 3.239 52.805 3.37 ;
      RECT 52.69 3.237 52.776 3.37 ;
      RECT 52.55 3.237 52.585 3.37 ;
      RECT 52.46 3.241 52.5 3.373 ;
      RECT 52.445 3.244 52.46 3.38 ;
      RECT 52.435 3.245 52.445 3.387 ;
      RECT 52.41 3.248 52.435 3.392 ;
      RECT 52.405 3.25 52.41 3.395 ;
      RECT 52.355 3.252 52.405 3.396 ;
      RECT 52.316 3.256 52.355 3.398 ;
      RECT 52.23 3.258 52.316 3.401 ;
      RECT 52.212 3.26 52.23 3.403 ;
      RECT 52.126 3.263 52.212 3.405 ;
      RECT 52.04 3.267 52.126 3.408 ;
      RECT 52.003 3.271 52.04 3.411 ;
      RECT 51.917 3.274 52.003 3.414 ;
      RECT 51.831 3.278 51.917 3.417 ;
      RECT 51.745 3.283 51.831 3.421 ;
      RECT 51.725 3.285 51.745 3.424 ;
      RECT 51.705 3.284 51.725 3.425 ;
      RECT 51.656 3.281 51.705 3.426 ;
      RECT 51.57 3.276 51.656 3.429 ;
      RECT 51.52 3.271 51.57 3.431 ;
      RECT 51.496 3.269 51.52 3.432 ;
      RECT 51.41 3.264 51.496 3.434 ;
      RECT 51.385 3.26 51.41 3.433 ;
      RECT 51.375 3.257 51.385 3.431 ;
      RECT 51.365 3.25 51.375 3.428 ;
      RECT 51.36 3.23 51.365 3.423 ;
      RECT 51.35 3.2 51.36 3.418 ;
      RECT 51.335 3.07 51.35 3.409 ;
      RECT 51.33 3.062 51.335 3.402 ;
      RECT 51.31 3.055 51.33 3.394 ;
      RECT 51.305 3.037 51.31 3.386 ;
      RECT 51.295 3.017 51.305 3.381 ;
      RECT 51.29 2.99 51.295 3.377 ;
      RECT 51.285 2.967 51.29 3.374 ;
      RECT 51.265 2.925 51.285 3.366 ;
      RECT 51.23 2.84 51.265 3.35 ;
      RECT 51.225 2.772 51.23 3.338 ;
      RECT 51.21 2.742 51.225 3.332 ;
      RECT 51.205 1.987 51.21 2.233 ;
      RECT 51.195 2.712 51.21 3.323 ;
      RECT 51.2 1.982 51.205 2.265 ;
      RECT 51.195 1.977 51.2 2.308 ;
      RECT 51.19 1.975 51.195 2.343 ;
      RECT 51.175 2.675 51.195 3.313 ;
      RECT 51.185 1.975 51.19 2.38 ;
      RECT 51.17 1.975 51.185 2.478 ;
      RECT 51.17 2.648 51.175 3.306 ;
      RECT 51.165 1.975 51.17 2.553 ;
      RECT 51.165 2.636 51.17 3.303 ;
      RECT 51.16 1.975 51.165 2.585 ;
      RECT 51.16 2.615 51.165 3.3 ;
      RECT 51.155 1.975 51.16 3.297 ;
      RECT 51.12 1.975 51.155 3.283 ;
      RECT 51.105 1.975 51.12 3.265 ;
      RECT 51.085 1.975 51.105 3.255 ;
      RECT 51.06 1.975 51.085 3.238 ;
      RECT 51.055 1.975 51.06 3.188 ;
      RECT 51.045 1.975 51.05 3.018 ;
      RECT 51.04 1.975 51.045 2.925 ;
      RECT 51.035 1.975 51.04 2.838 ;
      RECT 51.03 1.975 51.035 2.77 ;
      RECT 51.025 1.975 51.03 2.713 ;
      RECT 51.015 1.975 51.025 2.608 ;
      RECT 51.01 1.975 51.015 2.48 ;
      RECT 51.005 1.975 51.01 2.398 ;
      RECT 51 1.977 51.005 2.315 ;
      RECT 50.995 1.982 51 2.248 ;
      RECT 50.99 1.987 50.995 2.175 ;
      RECT 53.805 2.305 54.065 2.565 ;
      RECT 53.825 2.272 54.035 2.565 ;
      RECT 53.825 2.27 54.025 2.565 ;
      RECT 53.835 2.257 54.025 2.565 ;
      RECT 53.835 2.255 53.95 2.565 ;
      RECT 53.31 2.38 53.485 2.66 ;
      RECT 53.305 2.38 53.485 2.658 ;
      RECT 53.305 2.38 53.5 2.655 ;
      RECT 53.295 2.38 53.5 2.653 ;
      RECT 53.24 2.38 53.5 2.64 ;
      RECT 53.24 2.455 53.505 2.618 ;
      RECT 52.785 2.392 52.805 2.635 ;
      RECT 52.785 2.392 52.845 2.634 ;
      RECT 52.78 2.394 52.845 2.633 ;
      RECT 52.78 2.394 52.931 2.632 ;
      RECT 52.78 2.394 53 2.631 ;
      RECT 52.78 2.394 53.02 2.623 ;
      RECT 52.76 2.397 53.02 2.621 ;
      RECT 52.745 2.407 53.02 2.606 ;
      RECT 52.745 2.407 53.035 2.605 ;
      RECT 52.74 2.416 53.035 2.597 ;
      RECT 52.74 2.416 53.04 2.593 ;
      RECT 52.845 2.33 53.105 2.59 ;
      RECT 52.735 2.418 53.105 2.475 ;
      RECT 52.805 2.385 53.105 2.59 ;
      RECT 52.77 3.578 52.775 3.785 ;
      RECT 52.72 3.572 52.77 3.784 ;
      RECT 52.687 3.586 52.78 3.783 ;
      RECT 52.601 3.586 52.78 3.782 ;
      RECT 52.515 3.586 52.78 3.781 ;
      RECT 52.515 3.685 52.785 3.778 ;
      RECT 52.51 3.685 52.785 3.773 ;
      RECT 52.505 3.685 52.785 3.755 ;
      RECT 52.5 3.685 52.785 3.738 ;
      RECT 52.46 3.47 52.72 3.73 ;
      RECT 51.92 2.62 52.006 3.034 ;
      RECT 51.92 2.62 52.045 3.031 ;
      RECT 51.92 2.62 52.065 3.021 ;
      RECT 51.875 2.62 52.065 3.018 ;
      RECT 51.875 2.772 52.075 3.008 ;
      RECT 51.875 2.793 52.08 3.002 ;
      RECT 51.875 2.811 52.085 2.998 ;
      RECT 51.875 2.831 52.095 2.993 ;
      RECT 51.85 2.831 52.095 2.99 ;
      RECT 51.84 2.831 52.095 2.968 ;
      RECT 51.84 2.847 52.1 2.938 ;
      RECT 51.805 2.62 52.065 2.925 ;
      RECT 51.805 2.859 52.105 2.88 ;
      RECT 49.465 7.77 49.755 8 ;
      RECT 49.525 6.29 49.695 8 ;
      RECT 49.475 6.655 49.825 7.005 ;
      RECT 49.465 6.29 49.755 6.52 ;
      RECT 49.06 2.395 49.165 2.965 ;
      RECT 49.06 2.73 49.385 2.96 ;
      RECT 49.06 2.76 49.555 2.93 ;
      RECT 49.06 2.395 49.25 2.96 ;
      RECT 48.475 2.36 48.765 2.59 ;
      RECT 48.475 2.395 49.25 2.565 ;
      RECT 48.535 0.88 48.705 2.59 ;
      RECT 48.475 0.88 48.765 1.11 ;
      RECT 48.475 7.77 48.765 8 ;
      RECT 48.535 6.29 48.705 8 ;
      RECT 48.475 6.29 48.765 6.52 ;
      RECT 48.475 6.325 49.33 6.485 ;
      RECT 49.16 5.92 49.33 6.485 ;
      RECT 48.475 6.32 48.87 6.485 ;
      RECT 49.095 5.92 49.385 6.15 ;
      RECT 49.095 5.95 49.555 6.12 ;
      RECT 48.105 2.73 48.395 2.96 ;
      RECT 48.105 2.76 48.565 2.93 ;
      RECT 48.17 1.655 48.335 2.96 ;
      RECT 46.685 1.625 46.975 1.855 ;
      RECT 46.685 1.655 48.335 1.825 ;
      RECT 46.745 0.885 46.915 1.855 ;
      RECT 46.685 0.885 46.975 1.115 ;
      RECT 46.685 7.765 46.975 7.995 ;
      RECT 46.745 7.025 46.915 7.995 ;
      RECT 46.745 7.12 48.335 7.29 ;
      RECT 48.165 5.92 48.335 7.29 ;
      RECT 46.685 7.025 46.975 7.255 ;
      RECT 48.105 5.92 48.395 6.15 ;
      RECT 48.105 5.95 48.565 6.12 ;
      RECT 44.735 2.705 45.075 3.055 ;
      RECT 44.825 2.025 44.995 3.055 ;
      RECT 47.115 1.965 47.465 2.315 ;
      RECT 44.825 2.025 47.465 2.195 ;
      RECT 47.14 6.655 47.465 6.98 ;
      RECT 41.68 6.615 42.03 6.965 ;
      RECT 47.115 6.655 47.465 6.885 ;
      RECT 41.48 6.655 42.03 6.885 ;
      RECT 41.31 6.685 47.465 6.855 ;
      RECT 46.34 2.365 46.66 2.685 ;
      RECT 46.31 2.365 46.66 2.595 ;
      RECT 46.14 2.395 46.66 2.565 ;
      RECT 46.34 6.255 46.66 6.545 ;
      RECT 46.31 6.285 46.66 6.515 ;
      RECT 46.14 6.315 46.66 6.485 ;
      RECT 42.03 2.985 42.18 3.26 ;
      RECT 42.57 2.065 42.575 2.285 ;
      RECT 43.72 2.265 43.735 2.463 ;
      RECT 43.685 2.257 43.72 2.47 ;
      RECT 43.655 2.25 43.685 2.47 ;
      RECT 43.6 2.215 43.655 2.47 ;
      RECT 43.535 2.152 43.6 2.47 ;
      RECT 43.53 2.117 43.535 2.468 ;
      RECT 43.525 2.112 43.53 2.46 ;
      RECT 43.52 2.107 43.525 2.446 ;
      RECT 43.515 2.104 43.52 2.439 ;
      RECT 43.47 2.094 43.515 2.39 ;
      RECT 43.45 2.081 43.47 2.325 ;
      RECT 43.445 2.076 43.45 2.298 ;
      RECT 43.44 2.075 43.445 2.291 ;
      RECT 43.435 2.074 43.44 2.284 ;
      RECT 43.35 2.059 43.435 2.23 ;
      RECT 43.32 2.04 43.35 2.18 ;
      RECT 43.24 2.023 43.32 2.165 ;
      RECT 43.205 2.01 43.24 2.15 ;
      RECT 43.197 2.01 43.205 2.145 ;
      RECT 43.111 2.011 43.197 2.145 ;
      RECT 43.025 2.013 43.111 2.145 ;
      RECT 43 2.014 43.025 2.149 ;
      RECT 42.925 2.02 43 2.164 ;
      RECT 42.842 2.032 42.925 2.188 ;
      RECT 42.756 2.045 42.842 2.214 ;
      RECT 42.67 2.058 42.756 2.24 ;
      RECT 42.635 2.067 42.67 2.259 ;
      RECT 42.585 2.067 42.635 2.272 ;
      RECT 42.575 2.065 42.585 2.283 ;
      RECT 42.56 2.062 42.57 2.285 ;
      RECT 42.545 2.054 42.56 2.293 ;
      RECT 42.53 2.046 42.545 2.313 ;
      RECT 42.525 2.041 42.53 2.37 ;
      RECT 42.51 2.036 42.525 2.443 ;
      RECT 42.505 2.031 42.51 2.485 ;
      RECT 42.5 2.029 42.505 2.513 ;
      RECT 42.495 2.027 42.5 2.535 ;
      RECT 42.485 2.023 42.495 2.578 ;
      RECT 42.48 2.02 42.485 2.603 ;
      RECT 42.475 2.018 42.48 2.623 ;
      RECT 42.47 2.016 42.475 2.647 ;
      RECT 42.465 2.012 42.47 2.67 ;
      RECT 42.46 2.008 42.465 2.693 ;
      RECT 42.425 1.998 42.46 2.8 ;
      RECT 42.42 1.988 42.425 2.898 ;
      RECT 42.415 1.986 42.42 2.925 ;
      RECT 42.41 1.985 42.415 2.945 ;
      RECT 42.405 1.977 42.41 2.965 ;
      RECT 42.4 1.972 42.405 3 ;
      RECT 42.395 1.97 42.4 3.018 ;
      RECT 42.39 1.97 42.395 3.043 ;
      RECT 42.385 1.97 42.39 3.065 ;
      RECT 42.35 1.97 42.385 3.108 ;
      RECT 42.325 1.97 42.35 3.137 ;
      RECT 42.315 1.97 42.325 2.323 ;
      RECT 42.318 2.38 42.325 3.147 ;
      RECT 42.315 2.437 42.318 3.15 ;
      RECT 42.31 1.97 42.315 2.295 ;
      RECT 42.31 2.487 42.315 3.153 ;
      RECT 42.3 1.97 42.31 2.285 ;
      RECT 42.305 2.54 42.31 3.156 ;
      RECT 42.3 2.625 42.305 3.16 ;
      RECT 42.29 1.97 42.3 2.273 ;
      RECT 42.295 2.672 42.3 3.164 ;
      RECT 42.29 2.747 42.295 3.168 ;
      RECT 42.255 1.97 42.29 2.248 ;
      RECT 42.28 2.83 42.29 3.173 ;
      RECT 42.27 2.897 42.28 3.18 ;
      RECT 42.265 2.925 42.27 3.185 ;
      RECT 42.255 2.938 42.265 3.191 ;
      RECT 42.21 1.97 42.255 2.205 ;
      RECT 42.25 2.943 42.255 3.198 ;
      RECT 42.21 2.96 42.25 3.26 ;
      RECT 42.205 1.972 42.21 2.178 ;
      RECT 42.18 2.98 42.21 3.26 ;
      RECT 42.2 1.977 42.205 2.15 ;
      RECT 41.99 2.989 42.03 3.26 ;
      RECT 41.965 2.997 41.99 3.23 ;
      RECT 41.92 3.005 41.965 3.23 ;
      RECT 41.905 3.01 41.92 3.225 ;
      RECT 41.895 3.01 41.905 3.219 ;
      RECT 41.885 3.017 41.895 3.216 ;
      RECT 41.88 3.055 41.885 3.205 ;
      RECT 41.875 3.117 41.88 3.183 ;
      RECT 43.145 2.992 43.33 3.215 ;
      RECT 43.145 3.007 43.335 3.211 ;
      RECT 43.135 2.28 43.22 3.21 ;
      RECT 43.135 3.007 43.34 3.204 ;
      RECT 43.13 3.015 43.34 3.203 ;
      RECT 43.335 2.735 43.655 3.055 ;
      RECT 43.13 2.907 43.3 2.998 ;
      RECT 43.125 2.907 43.3 2.98 ;
      RECT 43.115 2.715 43.25 2.955 ;
      RECT 43.11 2.715 43.25 2.9 ;
      RECT 43.07 2.295 43.24 2.8 ;
      RECT 43.055 2.295 43.24 2.67 ;
      RECT 43.05 2.295 43.24 2.623 ;
      RECT 43.045 2.295 43.24 2.603 ;
      RECT 43.04 2.295 43.24 2.578 ;
      RECT 43.01 2.295 43.27 2.555 ;
      RECT 43.02 2.292 43.23 2.555 ;
      RECT 43.145 2.287 43.23 3.215 ;
      RECT 43.03 2.28 43.22 2.555 ;
      RECT 43.025 2.285 43.22 2.555 ;
      RECT 41.855 2.497 42.04 2.71 ;
      RECT 41.855 2.505 42.05 2.703 ;
      RECT 41.835 2.505 42.05 2.7 ;
      RECT 41.83 2.505 42.05 2.685 ;
      RECT 41.76 2.42 42.02 2.68 ;
      RECT 41.76 2.565 42.055 2.593 ;
      RECT 41.415 3.02 41.675 3.28 ;
      RECT 41.44 2.965 41.635 3.28 ;
      RECT 41.435 2.714 41.615 3.008 ;
      RECT 41.435 2.72 41.625 3.008 ;
      RECT 41.415 2.722 41.625 2.953 ;
      RECT 41.41 2.732 41.625 2.82 ;
      RECT 41.44 2.712 41.615 3.28 ;
      RECT 41.526 2.71 41.615 3.28 ;
      RECT 41.385 1.93 41.42 2.3 ;
      RECT 41.175 2.04 41.18 2.3 ;
      RECT 41.42 1.937 41.435 2.3 ;
      RECT 41.31 1.93 41.385 2.378 ;
      RECT 41.3 1.93 41.31 2.463 ;
      RECT 41.275 1.93 41.3 2.498 ;
      RECT 41.235 1.93 41.275 2.566 ;
      RECT 41.225 1.937 41.235 2.618 ;
      RECT 41.195 2.04 41.225 2.659 ;
      RECT 41.19 2.04 41.195 2.698 ;
      RECT 41.18 2.04 41.19 2.718 ;
      RECT 41.175 2.335 41.18 2.755 ;
      RECT 41.17 2.352 41.175 2.775 ;
      RECT 41.155 2.415 41.17 2.815 ;
      RECT 41.15 2.458 41.155 2.85 ;
      RECT 41.145 2.466 41.15 2.863 ;
      RECT 41.135 2.48 41.145 2.885 ;
      RECT 41.11 2.515 41.135 2.95 ;
      RECT 41.1 2.55 41.11 3.013 ;
      RECT 41.08 2.58 41.1 3.074 ;
      RECT 41.065 2.616 41.08 3.141 ;
      RECT 41.055 2.644 41.065 3.18 ;
      RECT 41.045 2.666 41.055 3.2 ;
      RECT 41.04 2.676 41.045 3.211 ;
      RECT 41.035 2.685 41.04 3.214 ;
      RECT 41.025 2.703 41.035 3.218 ;
      RECT 41.015 2.721 41.025 3.219 ;
      RECT 40.99 2.76 41.015 3.216 ;
      RECT 40.97 2.802 40.99 3.213 ;
      RECT 40.955 2.84 40.97 3.212 ;
      RECT 40.92 2.875 40.955 3.209 ;
      RECT 40.915 2.897 40.92 3.207 ;
      RECT 40.85 2.937 40.915 3.204 ;
      RECT 40.845 2.977 40.85 3.2 ;
      RECT 40.83 2.987 40.845 3.191 ;
      RECT 40.82 3.107 40.83 3.176 ;
      RECT 41.3 3.52 41.31 3.78 ;
      RECT 41.3 3.523 41.32 3.779 ;
      RECT 41.29 3.513 41.3 3.778 ;
      RECT 41.28 3.528 41.36 3.774 ;
      RECT 41.265 3.507 41.28 3.772 ;
      RECT 41.24 3.532 41.365 3.768 ;
      RECT 41.225 3.492 41.24 3.763 ;
      RECT 41.225 3.534 41.375 3.762 ;
      RECT 41.225 3.542 41.39 3.755 ;
      RECT 41.165 3.479 41.225 3.745 ;
      RECT 41.155 3.466 41.165 3.727 ;
      RECT 41.13 3.456 41.155 3.717 ;
      RECT 41.125 3.446 41.13 3.709 ;
      RECT 41.06 3.542 41.39 3.691 ;
      RECT 40.975 3.542 41.39 3.653 ;
      RECT 40.865 3.37 41.125 3.63 ;
      RECT 41.24 3.5 41.265 3.768 ;
      RECT 41.28 3.51 41.29 3.774 ;
      RECT 40.865 3.518 41.305 3.63 ;
      RECT 41.05 7.765 41.34 7.995 ;
      RECT 41.11 7.025 41.28 7.995 ;
      RECT 41.01 7.055 41.38 7.425 ;
      RECT 41.05 7.025 41.34 7.425 ;
      RECT 40.08 3.275 40.11 3.575 ;
      RECT 39.855 3.26 39.86 3.535 ;
      RECT 39.655 3.26 39.81 3.52 ;
      RECT 40.955 1.975 40.985 2.235 ;
      RECT 40.945 1.975 40.955 2.343 ;
      RECT 40.925 1.975 40.945 2.353 ;
      RECT 40.91 1.975 40.925 2.365 ;
      RECT 40.855 1.975 40.91 2.415 ;
      RECT 40.84 1.975 40.855 2.463 ;
      RECT 40.81 1.975 40.84 2.498 ;
      RECT 40.755 1.975 40.81 2.56 ;
      RECT 40.735 1.975 40.755 2.628 ;
      RECT 40.73 1.975 40.735 2.658 ;
      RECT 40.725 1.975 40.73 2.67 ;
      RECT 40.72 2.092 40.725 2.688 ;
      RECT 40.7 2.11 40.72 2.713 ;
      RECT 40.68 2.137 40.7 2.763 ;
      RECT 40.675 2.157 40.68 2.794 ;
      RECT 40.67 2.165 40.675 2.811 ;
      RECT 40.655 2.191 40.67 2.84 ;
      RECT 40.64 2.233 40.655 2.875 ;
      RECT 40.635 2.262 40.64 2.898 ;
      RECT 40.63 2.277 40.635 2.911 ;
      RECT 40.625 2.3 40.63 2.922 ;
      RECT 40.615 2.32 40.625 2.94 ;
      RECT 40.605 2.35 40.615 2.963 ;
      RECT 40.6 2.372 40.605 2.983 ;
      RECT 40.595 2.387 40.6 2.998 ;
      RECT 40.58 2.417 40.595 3.025 ;
      RECT 40.575 2.447 40.58 3.051 ;
      RECT 40.57 2.465 40.575 3.063 ;
      RECT 40.56 2.495 40.57 3.082 ;
      RECT 40.55 2.52 40.56 3.107 ;
      RECT 40.545 2.54 40.55 3.126 ;
      RECT 40.54 2.557 40.545 3.139 ;
      RECT 40.53 2.583 40.54 3.158 ;
      RECT 40.52 2.621 40.53 3.185 ;
      RECT 40.515 2.647 40.52 3.205 ;
      RECT 40.51 2.657 40.515 3.215 ;
      RECT 40.505 2.67 40.51 3.23 ;
      RECT 40.5 2.685 40.505 3.24 ;
      RECT 40.495 2.707 40.5 3.255 ;
      RECT 40.49 2.725 40.495 3.266 ;
      RECT 40.485 2.735 40.49 3.277 ;
      RECT 40.48 2.743 40.485 3.289 ;
      RECT 40.475 2.751 40.48 3.3 ;
      RECT 40.47 2.777 40.475 3.313 ;
      RECT 40.46 2.805 40.47 3.326 ;
      RECT 40.455 2.835 40.46 3.335 ;
      RECT 40.45 2.85 40.455 3.342 ;
      RECT 40.435 2.875 40.45 3.349 ;
      RECT 40.43 2.897 40.435 3.355 ;
      RECT 40.425 2.922 40.43 3.358 ;
      RECT 40.416 2.95 40.425 3.362 ;
      RECT 40.41 2.967 40.416 3.367 ;
      RECT 40.405 2.985 40.41 3.371 ;
      RECT 40.4 2.997 40.405 3.374 ;
      RECT 40.395 3.018 40.4 3.378 ;
      RECT 40.39 3.036 40.395 3.381 ;
      RECT 40.385 3.05 40.39 3.384 ;
      RECT 40.38 3.067 40.385 3.387 ;
      RECT 40.375 3.08 40.38 3.39 ;
      RECT 40.35 3.117 40.375 3.398 ;
      RECT 40.345 3.162 40.35 3.407 ;
      RECT 40.34 3.19 40.345 3.41 ;
      RECT 40.33 3.21 40.34 3.414 ;
      RECT 40.325 3.23 40.33 3.419 ;
      RECT 40.32 3.245 40.325 3.422 ;
      RECT 40.3 3.255 40.32 3.429 ;
      RECT 40.235 3.262 40.3 3.455 ;
      RECT 40.2 3.265 40.235 3.483 ;
      RECT 40.185 3.268 40.2 3.498 ;
      RECT 40.175 3.269 40.185 3.513 ;
      RECT 40.165 3.27 40.175 3.53 ;
      RECT 40.16 3.27 40.165 3.545 ;
      RECT 40.155 3.27 40.16 3.553 ;
      RECT 40.14 3.271 40.155 3.568 ;
      RECT 40.11 3.273 40.14 3.575 ;
      RECT 40 3.28 40.08 3.575 ;
      RECT 39.955 3.285 40 3.575 ;
      RECT 39.945 3.286 39.955 3.565 ;
      RECT 39.935 3.287 39.945 3.558 ;
      RECT 39.915 3.289 39.935 3.553 ;
      RECT 39.905 3.26 39.915 3.548 ;
      RECT 39.86 3.26 39.905 3.54 ;
      RECT 39.83 3.26 39.855 3.53 ;
      RECT 39.81 3.26 39.83 3.523 ;
      RECT 40.09 2.06 40.35 2.32 ;
      RECT 39.97 2.075 39.98 2.24 ;
      RECT 39.955 2.075 39.96 2.235 ;
      RECT 37.32 1.915 37.505 2.205 ;
      RECT 39.135 2.04 39.15 2.195 ;
      RECT 37.285 1.915 37.31 2.175 ;
      RECT 39.7 1.965 39.705 2.107 ;
      RECT 39.615 1.96 39.64 2.1 ;
      RECT 40.015 2.077 40.09 2.27 ;
      RECT 40 2.075 40.015 2.253 ;
      RECT 39.98 2.075 40 2.245 ;
      RECT 39.96 2.075 39.97 2.238 ;
      RECT 39.915 2.07 39.955 2.228 ;
      RECT 39.875 2.045 39.915 2.213 ;
      RECT 39.86 2.02 39.875 2.203 ;
      RECT 39.855 2.014 39.86 2.201 ;
      RECT 39.82 2.006 39.855 2.184 ;
      RECT 39.815 1.999 39.82 2.172 ;
      RECT 39.795 1.994 39.815 2.16 ;
      RECT 39.785 1.988 39.795 2.145 ;
      RECT 39.765 1.983 39.785 2.13 ;
      RECT 39.755 1.978 39.765 2.123 ;
      RECT 39.75 1.976 39.755 2.118 ;
      RECT 39.745 1.975 39.75 2.115 ;
      RECT 39.705 1.97 39.745 2.111 ;
      RECT 39.685 1.964 39.7 2.106 ;
      RECT 39.65 1.961 39.685 2.103 ;
      RECT 39.64 1.96 39.65 2.101 ;
      RECT 39.58 1.96 39.615 2.098 ;
      RECT 39.535 1.96 39.58 2.098 ;
      RECT 39.485 1.96 39.535 2.101 ;
      RECT 39.47 1.962 39.485 2.103 ;
      RECT 39.455 1.965 39.47 2.104 ;
      RECT 39.445 1.97 39.455 2.105 ;
      RECT 39.415 1.975 39.445 2.11 ;
      RECT 39.405 1.981 39.415 2.118 ;
      RECT 39.395 1.983 39.405 2.122 ;
      RECT 39.385 1.987 39.395 2.126 ;
      RECT 39.36 1.993 39.385 2.134 ;
      RECT 39.35 1.998 39.36 2.142 ;
      RECT 39.335 2.002 39.35 2.146 ;
      RECT 39.3 2.008 39.335 2.154 ;
      RECT 39.28 2.013 39.3 2.164 ;
      RECT 39.25 2.02 39.28 2.173 ;
      RECT 39.205 2.029 39.25 2.187 ;
      RECT 39.2 2.034 39.205 2.198 ;
      RECT 39.18 2.037 39.2 2.199 ;
      RECT 39.15 2.04 39.18 2.197 ;
      RECT 39.115 2.04 39.135 2.193 ;
      RECT 39.045 2.04 39.115 2.184 ;
      RECT 39.03 2.037 39.045 2.176 ;
      RECT 38.99 2.03 39.03 2.171 ;
      RECT 38.965 2.02 38.99 2.164 ;
      RECT 38.96 2.014 38.965 2.161 ;
      RECT 38.92 2.008 38.96 2.158 ;
      RECT 38.905 2.001 38.92 2.153 ;
      RECT 38.885 1.997 38.905 2.148 ;
      RECT 38.87 1.992 38.885 2.144 ;
      RECT 38.855 1.987 38.87 2.142 ;
      RECT 38.84 1.983 38.855 2.141 ;
      RECT 38.825 1.981 38.84 2.137 ;
      RECT 38.815 1.979 38.825 2.132 ;
      RECT 38.8 1.976 38.815 2.128 ;
      RECT 38.79 1.974 38.8 2.123 ;
      RECT 38.77 1.971 38.79 2.119 ;
      RECT 38.725 1.97 38.77 2.117 ;
      RECT 38.665 1.972 38.725 2.118 ;
      RECT 38.645 1.974 38.665 2.12 ;
      RECT 38.615 1.977 38.645 2.121 ;
      RECT 38.565 1.982 38.615 2.123 ;
      RECT 38.56 1.985 38.565 2.125 ;
      RECT 38.55 1.987 38.56 2.128 ;
      RECT 38.545 1.989 38.55 2.131 ;
      RECT 38.495 1.992 38.545 2.138 ;
      RECT 38.475 1.996 38.495 2.15 ;
      RECT 38.465 1.999 38.475 2.156 ;
      RECT 38.455 2 38.465 2.159 ;
      RECT 38.416 2.003 38.455 2.161 ;
      RECT 38.33 2.01 38.416 2.164 ;
      RECT 38.256 2.02 38.33 2.168 ;
      RECT 38.17 2.031 38.256 2.173 ;
      RECT 38.155 2.038 38.17 2.175 ;
      RECT 38.1 2.042 38.155 2.176 ;
      RECT 38.086 2.045 38.1 2.178 ;
      RECT 38 2.045 38.086 2.18 ;
      RECT 37.96 2.042 38 2.183 ;
      RECT 37.936 2.038 37.96 2.185 ;
      RECT 37.85 2.028 37.936 2.188 ;
      RECT 37.82 2.017 37.85 2.189 ;
      RECT 37.801 2.013 37.82 2.188 ;
      RECT 37.715 2.006 37.801 2.185 ;
      RECT 37.655 1.995 37.715 2.182 ;
      RECT 37.635 1.987 37.655 2.18 ;
      RECT 37.6 1.982 37.635 2.179 ;
      RECT 37.575 1.977 37.6 2.178 ;
      RECT 37.545 1.972 37.575 2.177 ;
      RECT 37.52 1.915 37.545 2.176 ;
      RECT 37.505 1.915 37.52 2.2 ;
      RECT 37.31 1.915 37.32 2.2 ;
      RECT 39.085 2.935 39.09 3.075 ;
      RECT 38.745 2.935 38.78 3.073 ;
      RECT 38.32 2.92 38.335 3.065 ;
      RECT 40.15 2.7 40.24 2.96 ;
      RECT 39.98 2.565 40.08 2.96 ;
      RECT 37.015 2.54 37.095 2.75 ;
      RECT 40.105 2.677 40.15 2.96 ;
      RECT 40.095 2.647 40.105 2.96 ;
      RECT 40.08 2.57 40.095 2.96 ;
      RECT 39.895 2.565 39.98 2.925 ;
      RECT 39.89 2.567 39.895 2.92 ;
      RECT 39.885 2.572 39.89 2.92 ;
      RECT 39.85 2.672 39.885 2.92 ;
      RECT 39.84 2.7 39.85 2.92 ;
      RECT 39.83 2.715 39.84 2.92 ;
      RECT 39.82 2.727 39.83 2.92 ;
      RECT 39.815 2.737 39.82 2.92 ;
      RECT 39.8 2.747 39.815 2.922 ;
      RECT 39.795 2.762 39.8 2.924 ;
      RECT 39.78 2.775 39.795 2.926 ;
      RECT 39.775 2.79 39.78 2.929 ;
      RECT 39.755 2.8 39.775 2.933 ;
      RECT 39.74 2.81 39.755 2.936 ;
      RECT 39.705 2.817 39.74 2.941 ;
      RECT 39.661 2.824 39.705 2.949 ;
      RECT 39.575 2.836 39.661 2.962 ;
      RECT 39.55 2.847 39.575 2.973 ;
      RECT 39.52 2.852 39.55 2.978 ;
      RECT 39.485 2.857 39.52 2.986 ;
      RECT 39.455 2.862 39.485 2.993 ;
      RECT 39.43 2.867 39.455 2.998 ;
      RECT 39.365 2.874 39.43 3.007 ;
      RECT 39.295 2.887 39.365 3.023 ;
      RECT 39.265 2.897 39.295 3.035 ;
      RECT 39.24 2.902 39.265 3.042 ;
      RECT 39.185 2.909 39.24 3.05 ;
      RECT 39.18 2.916 39.185 3.055 ;
      RECT 39.175 2.918 39.18 3.056 ;
      RECT 39.16 2.92 39.175 3.058 ;
      RECT 39.155 2.92 39.16 3.061 ;
      RECT 39.09 2.927 39.155 3.068 ;
      RECT 39.055 2.937 39.085 3.078 ;
      RECT 39.038 2.94 39.055 3.08 ;
      RECT 38.952 2.939 39.038 3.079 ;
      RECT 38.866 2.937 38.952 3.076 ;
      RECT 38.78 2.936 38.866 3.074 ;
      RECT 38.679 2.934 38.745 3.073 ;
      RECT 38.593 2.931 38.679 3.071 ;
      RECT 38.507 2.927 38.593 3.069 ;
      RECT 38.421 2.924 38.507 3.068 ;
      RECT 38.335 2.921 38.421 3.066 ;
      RECT 38.235 2.92 38.32 3.063 ;
      RECT 38.185 2.918 38.235 3.061 ;
      RECT 38.165 2.915 38.185 3.059 ;
      RECT 38.145 2.913 38.165 3.056 ;
      RECT 38.12 2.909 38.145 3.053 ;
      RECT 38.075 2.903 38.12 3.048 ;
      RECT 38.035 2.897 38.075 3.04 ;
      RECT 38.01 2.892 38.035 3.033 ;
      RECT 37.955 2.885 38.01 3.025 ;
      RECT 37.931 2.878 37.955 3.018 ;
      RECT 37.845 2.869 37.931 3.008 ;
      RECT 37.815 2.861 37.845 2.998 ;
      RECT 37.785 2.857 37.815 2.993 ;
      RECT 37.78 2.854 37.785 2.99 ;
      RECT 37.775 2.853 37.78 2.99 ;
      RECT 37.7 2.846 37.775 2.983 ;
      RECT 37.661 2.837 37.7 2.972 ;
      RECT 37.575 2.827 37.661 2.96 ;
      RECT 37.535 2.817 37.575 2.948 ;
      RECT 37.496 2.812 37.535 2.941 ;
      RECT 37.41 2.802 37.496 2.93 ;
      RECT 37.37 2.79 37.41 2.919 ;
      RECT 37.335 2.775 37.37 2.912 ;
      RECT 37.325 2.765 37.335 2.909 ;
      RECT 37.305 2.75 37.325 2.907 ;
      RECT 37.275 2.72 37.305 2.903 ;
      RECT 37.265 2.7 37.275 2.898 ;
      RECT 37.26 2.692 37.265 2.895 ;
      RECT 37.255 2.685 37.26 2.893 ;
      RECT 37.24 2.672 37.255 2.886 ;
      RECT 37.235 2.662 37.24 2.878 ;
      RECT 37.23 2.655 37.235 2.873 ;
      RECT 37.225 2.65 37.23 2.869 ;
      RECT 37.21 2.637 37.225 2.861 ;
      RECT 37.205 2.547 37.21 2.85 ;
      RECT 37.2 2.542 37.205 2.843 ;
      RECT 37.125 2.54 37.2 2.803 ;
      RECT 37.095 2.54 37.125 2.758 ;
      RECT 37 2.545 37.015 2.745 ;
      RECT 39.485 2.25 39.745 2.51 ;
      RECT 39.47 2.238 39.65 2.475 ;
      RECT 39.465 2.239 39.65 2.473 ;
      RECT 39.45 2.243 39.66 2.463 ;
      RECT 39.445 2.248 39.665 2.433 ;
      RECT 39.45 2.245 39.665 2.463 ;
      RECT 39.465 2.24 39.66 2.473 ;
      RECT 39.485 2.237 39.65 2.51 ;
      RECT 39.485 2.236 39.64 2.51 ;
      RECT 39.51 2.235 39.64 2.51 ;
      RECT 39.07 2.48 39.33 2.74 ;
      RECT 38.945 2.525 39.33 2.735 ;
      RECT 38.935 2.53 39.33 2.73 ;
      RECT 38.95 3.47 38.965 3.78 ;
      RECT 37.545 3.24 37.555 3.37 ;
      RECT 37.325 3.235 37.43 3.37 ;
      RECT 37.24 3.24 37.29 3.37 ;
      RECT 35.79 1.975 35.795 3.08 ;
      RECT 39.045 3.562 39.05 3.698 ;
      RECT 39.04 3.557 39.045 3.758 ;
      RECT 39.035 3.555 39.04 3.771 ;
      RECT 39.02 3.552 39.035 3.773 ;
      RECT 39.015 3.547 39.02 3.775 ;
      RECT 39.01 3.543 39.015 3.778 ;
      RECT 38.995 3.538 39.01 3.78 ;
      RECT 38.965 3.53 38.995 3.78 ;
      RECT 38.926 3.47 38.95 3.78 ;
      RECT 38.84 3.47 38.926 3.777 ;
      RECT 38.81 3.47 38.84 3.77 ;
      RECT 38.785 3.47 38.81 3.763 ;
      RECT 38.76 3.47 38.785 3.755 ;
      RECT 38.745 3.47 38.76 3.748 ;
      RECT 38.72 3.47 38.745 3.74 ;
      RECT 38.705 3.47 38.72 3.733 ;
      RECT 38.665 3.48 38.705 3.722 ;
      RECT 38.655 3.475 38.665 3.712 ;
      RECT 38.651 3.474 38.655 3.709 ;
      RECT 38.565 3.466 38.651 3.692 ;
      RECT 38.532 3.455 38.565 3.669 ;
      RECT 38.446 3.444 38.532 3.647 ;
      RECT 38.36 3.428 38.446 3.616 ;
      RECT 38.29 3.413 38.36 3.588 ;
      RECT 38.28 3.406 38.29 3.575 ;
      RECT 38.25 3.403 38.28 3.565 ;
      RECT 38.225 3.399 38.25 3.558 ;
      RECT 38.21 3.396 38.225 3.553 ;
      RECT 38.205 3.395 38.21 3.548 ;
      RECT 38.175 3.39 38.205 3.541 ;
      RECT 38.17 3.385 38.175 3.536 ;
      RECT 38.155 3.382 38.17 3.531 ;
      RECT 38.15 3.377 38.155 3.526 ;
      RECT 38.13 3.372 38.15 3.523 ;
      RECT 38.115 3.367 38.13 3.515 ;
      RECT 38.1 3.361 38.115 3.51 ;
      RECT 38.07 3.352 38.1 3.503 ;
      RECT 38.065 3.345 38.07 3.495 ;
      RECT 38.06 3.343 38.065 3.493 ;
      RECT 38.055 3.342 38.06 3.49 ;
      RECT 38.015 3.335 38.055 3.483 ;
      RECT 38.001 3.325 38.015 3.473 ;
      RECT 37.95 3.314 38.001 3.461 ;
      RECT 37.925 3.3 37.95 3.447 ;
      RECT 37.9 3.289 37.925 3.439 ;
      RECT 37.88 3.278 37.9 3.433 ;
      RECT 37.87 3.272 37.88 3.428 ;
      RECT 37.865 3.27 37.87 3.424 ;
      RECT 37.845 3.265 37.865 3.419 ;
      RECT 37.815 3.255 37.845 3.409 ;
      RECT 37.81 3.247 37.815 3.402 ;
      RECT 37.795 3.245 37.81 3.398 ;
      RECT 37.775 3.245 37.795 3.393 ;
      RECT 37.77 3.244 37.775 3.391 ;
      RECT 37.765 3.244 37.77 3.388 ;
      RECT 37.725 3.243 37.765 3.383 ;
      RECT 37.7 3.242 37.725 3.378 ;
      RECT 37.64 3.241 37.7 3.375 ;
      RECT 37.555 3.24 37.64 3.373 ;
      RECT 37.516 3.239 37.545 3.37 ;
      RECT 37.43 3.237 37.516 3.37 ;
      RECT 37.29 3.237 37.325 3.37 ;
      RECT 37.2 3.241 37.24 3.373 ;
      RECT 37.185 3.244 37.2 3.38 ;
      RECT 37.175 3.245 37.185 3.387 ;
      RECT 37.15 3.248 37.175 3.392 ;
      RECT 37.145 3.25 37.15 3.395 ;
      RECT 37.095 3.252 37.145 3.396 ;
      RECT 37.056 3.256 37.095 3.398 ;
      RECT 36.97 3.258 37.056 3.401 ;
      RECT 36.952 3.26 36.97 3.403 ;
      RECT 36.866 3.263 36.952 3.405 ;
      RECT 36.78 3.267 36.866 3.408 ;
      RECT 36.743 3.271 36.78 3.411 ;
      RECT 36.657 3.274 36.743 3.414 ;
      RECT 36.571 3.278 36.657 3.417 ;
      RECT 36.485 3.283 36.571 3.421 ;
      RECT 36.465 3.285 36.485 3.424 ;
      RECT 36.445 3.284 36.465 3.425 ;
      RECT 36.396 3.281 36.445 3.426 ;
      RECT 36.31 3.276 36.396 3.429 ;
      RECT 36.26 3.271 36.31 3.431 ;
      RECT 36.236 3.269 36.26 3.432 ;
      RECT 36.15 3.264 36.236 3.434 ;
      RECT 36.125 3.26 36.15 3.433 ;
      RECT 36.115 3.257 36.125 3.431 ;
      RECT 36.105 3.25 36.115 3.428 ;
      RECT 36.1 3.23 36.105 3.423 ;
      RECT 36.09 3.2 36.1 3.418 ;
      RECT 36.075 3.07 36.09 3.409 ;
      RECT 36.07 3.062 36.075 3.402 ;
      RECT 36.05 3.055 36.07 3.394 ;
      RECT 36.045 3.037 36.05 3.386 ;
      RECT 36.035 3.017 36.045 3.381 ;
      RECT 36.03 2.99 36.035 3.377 ;
      RECT 36.025 2.967 36.03 3.374 ;
      RECT 36.005 2.925 36.025 3.366 ;
      RECT 35.97 2.84 36.005 3.35 ;
      RECT 35.965 2.772 35.97 3.338 ;
      RECT 35.95 2.742 35.965 3.332 ;
      RECT 35.945 1.987 35.95 2.233 ;
      RECT 35.935 2.712 35.95 3.323 ;
      RECT 35.94 1.982 35.945 2.265 ;
      RECT 35.935 1.977 35.94 2.308 ;
      RECT 35.93 1.975 35.935 2.343 ;
      RECT 35.915 2.675 35.935 3.313 ;
      RECT 35.925 1.975 35.93 2.38 ;
      RECT 35.91 1.975 35.925 2.478 ;
      RECT 35.91 2.648 35.915 3.306 ;
      RECT 35.905 1.975 35.91 2.553 ;
      RECT 35.905 2.636 35.91 3.303 ;
      RECT 35.9 1.975 35.905 2.585 ;
      RECT 35.9 2.615 35.905 3.3 ;
      RECT 35.895 1.975 35.9 3.297 ;
      RECT 35.86 1.975 35.895 3.283 ;
      RECT 35.845 1.975 35.86 3.265 ;
      RECT 35.825 1.975 35.845 3.255 ;
      RECT 35.8 1.975 35.825 3.238 ;
      RECT 35.795 1.975 35.8 3.188 ;
      RECT 35.785 1.975 35.79 3.018 ;
      RECT 35.78 1.975 35.785 2.925 ;
      RECT 35.775 1.975 35.78 2.838 ;
      RECT 35.77 1.975 35.775 2.77 ;
      RECT 35.765 1.975 35.77 2.713 ;
      RECT 35.755 1.975 35.765 2.608 ;
      RECT 35.75 1.975 35.755 2.48 ;
      RECT 35.745 1.975 35.75 2.398 ;
      RECT 35.74 1.977 35.745 2.315 ;
      RECT 35.735 1.982 35.74 2.248 ;
      RECT 35.73 1.987 35.735 2.175 ;
      RECT 38.545 2.305 38.805 2.565 ;
      RECT 38.565 2.272 38.775 2.565 ;
      RECT 38.565 2.27 38.765 2.565 ;
      RECT 38.575 2.257 38.765 2.565 ;
      RECT 38.575 2.255 38.69 2.565 ;
      RECT 38.05 2.38 38.225 2.66 ;
      RECT 38.045 2.38 38.225 2.658 ;
      RECT 38.045 2.38 38.24 2.655 ;
      RECT 38.035 2.38 38.24 2.653 ;
      RECT 37.98 2.38 38.24 2.64 ;
      RECT 37.98 2.455 38.245 2.618 ;
      RECT 37.525 2.392 37.545 2.635 ;
      RECT 37.525 2.392 37.585 2.634 ;
      RECT 37.52 2.394 37.585 2.633 ;
      RECT 37.52 2.394 37.671 2.632 ;
      RECT 37.52 2.394 37.74 2.631 ;
      RECT 37.52 2.394 37.76 2.623 ;
      RECT 37.5 2.397 37.76 2.621 ;
      RECT 37.485 2.407 37.76 2.606 ;
      RECT 37.485 2.407 37.775 2.605 ;
      RECT 37.48 2.416 37.775 2.597 ;
      RECT 37.48 2.416 37.78 2.593 ;
      RECT 37.585 2.33 37.845 2.59 ;
      RECT 37.475 2.418 37.845 2.475 ;
      RECT 37.545 2.385 37.845 2.59 ;
      RECT 37.51 3.578 37.515 3.785 ;
      RECT 37.46 3.572 37.51 3.784 ;
      RECT 37.427 3.586 37.52 3.783 ;
      RECT 37.341 3.586 37.52 3.782 ;
      RECT 37.255 3.586 37.52 3.781 ;
      RECT 37.255 3.685 37.525 3.778 ;
      RECT 37.25 3.685 37.525 3.773 ;
      RECT 37.245 3.685 37.525 3.755 ;
      RECT 37.24 3.685 37.525 3.738 ;
      RECT 37.2 3.47 37.46 3.73 ;
      RECT 36.66 2.62 36.746 3.034 ;
      RECT 36.66 2.62 36.785 3.031 ;
      RECT 36.66 2.62 36.805 3.021 ;
      RECT 36.615 2.62 36.805 3.018 ;
      RECT 36.615 2.772 36.815 3.008 ;
      RECT 36.615 2.793 36.82 3.002 ;
      RECT 36.615 2.811 36.825 2.998 ;
      RECT 36.615 2.831 36.835 2.993 ;
      RECT 36.59 2.831 36.835 2.99 ;
      RECT 36.58 2.831 36.835 2.968 ;
      RECT 36.58 2.847 36.84 2.938 ;
      RECT 36.545 2.62 36.805 2.925 ;
      RECT 36.545 2.859 36.845 2.88 ;
      RECT 34.205 7.77 34.495 8 ;
      RECT 34.265 6.29 34.435 8 ;
      RECT 34.255 6.66 34.61 7.015 ;
      RECT 34.205 6.29 34.495 6.52 ;
      RECT 33.8 2.395 33.905 2.965 ;
      RECT 33.8 2.73 34.125 2.96 ;
      RECT 33.8 2.76 34.295 2.93 ;
      RECT 33.8 2.395 33.99 2.96 ;
      RECT 33.215 2.36 33.505 2.59 ;
      RECT 33.215 2.395 33.99 2.565 ;
      RECT 33.275 0.88 33.445 2.59 ;
      RECT 33.215 0.88 33.505 1.11 ;
      RECT 33.215 7.77 33.505 8 ;
      RECT 33.275 6.29 33.445 8 ;
      RECT 33.215 6.29 33.505 6.52 ;
      RECT 33.215 6.325 34.07 6.485 ;
      RECT 33.9 5.92 34.07 6.485 ;
      RECT 33.215 6.32 33.61 6.485 ;
      RECT 33.835 5.92 34.125 6.15 ;
      RECT 33.835 5.95 34.295 6.12 ;
      RECT 32.845 2.73 33.135 2.96 ;
      RECT 32.845 2.76 33.305 2.93 ;
      RECT 32.91 1.655 33.075 2.96 ;
      RECT 31.425 1.625 31.715 1.855 ;
      RECT 31.425 1.655 33.075 1.825 ;
      RECT 31.485 0.885 31.655 1.855 ;
      RECT 31.425 0.885 31.715 1.115 ;
      RECT 31.425 7.765 31.715 7.995 ;
      RECT 31.485 7.025 31.655 7.995 ;
      RECT 31.485 7.12 33.075 7.29 ;
      RECT 32.905 5.92 33.075 7.29 ;
      RECT 31.425 7.025 31.715 7.255 ;
      RECT 32.845 5.92 33.135 6.15 ;
      RECT 32.845 5.95 33.305 6.12 ;
      RECT 29.475 2.705 29.815 3.055 ;
      RECT 29.565 2.025 29.735 3.055 ;
      RECT 31.855 1.965 32.205 2.315 ;
      RECT 29.565 2.025 32.205 2.195 ;
      RECT 31.88 6.655 32.205 6.98 ;
      RECT 26.42 6.61 26.77 6.96 ;
      RECT 31.855 6.655 32.205 6.885 ;
      RECT 26.22 6.655 26.77 6.885 ;
      RECT 26.05 6.685 32.205 6.855 ;
      RECT 31.08 2.365 31.4 2.685 ;
      RECT 31.05 2.365 31.4 2.595 ;
      RECT 30.88 2.395 31.4 2.565 ;
      RECT 31.08 6.255 31.4 6.545 ;
      RECT 31.05 6.285 31.4 6.515 ;
      RECT 30.88 6.315 31.4 6.485 ;
      RECT 26.77 2.985 26.92 3.26 ;
      RECT 27.31 2.065 27.315 2.285 ;
      RECT 28.46 2.265 28.475 2.463 ;
      RECT 28.425 2.257 28.46 2.47 ;
      RECT 28.395 2.25 28.425 2.47 ;
      RECT 28.34 2.215 28.395 2.47 ;
      RECT 28.275 2.152 28.34 2.47 ;
      RECT 28.27 2.117 28.275 2.468 ;
      RECT 28.265 2.112 28.27 2.46 ;
      RECT 28.26 2.107 28.265 2.446 ;
      RECT 28.255 2.104 28.26 2.439 ;
      RECT 28.21 2.094 28.255 2.39 ;
      RECT 28.19 2.081 28.21 2.325 ;
      RECT 28.185 2.076 28.19 2.298 ;
      RECT 28.18 2.075 28.185 2.291 ;
      RECT 28.175 2.074 28.18 2.284 ;
      RECT 28.09 2.059 28.175 2.23 ;
      RECT 28.06 2.04 28.09 2.18 ;
      RECT 27.98 2.023 28.06 2.165 ;
      RECT 27.945 2.01 27.98 2.15 ;
      RECT 27.937 2.01 27.945 2.145 ;
      RECT 27.851 2.011 27.937 2.145 ;
      RECT 27.765 2.013 27.851 2.145 ;
      RECT 27.74 2.014 27.765 2.149 ;
      RECT 27.665 2.02 27.74 2.164 ;
      RECT 27.582 2.032 27.665 2.188 ;
      RECT 27.496 2.045 27.582 2.214 ;
      RECT 27.41 2.058 27.496 2.24 ;
      RECT 27.375 2.067 27.41 2.259 ;
      RECT 27.325 2.067 27.375 2.272 ;
      RECT 27.315 2.065 27.325 2.283 ;
      RECT 27.3 2.062 27.31 2.285 ;
      RECT 27.285 2.054 27.3 2.293 ;
      RECT 27.27 2.046 27.285 2.313 ;
      RECT 27.265 2.041 27.27 2.37 ;
      RECT 27.25 2.036 27.265 2.443 ;
      RECT 27.245 2.031 27.25 2.485 ;
      RECT 27.24 2.029 27.245 2.513 ;
      RECT 27.235 2.027 27.24 2.535 ;
      RECT 27.225 2.023 27.235 2.578 ;
      RECT 27.22 2.02 27.225 2.603 ;
      RECT 27.215 2.018 27.22 2.623 ;
      RECT 27.21 2.016 27.215 2.647 ;
      RECT 27.205 2.012 27.21 2.67 ;
      RECT 27.2 2.008 27.205 2.693 ;
      RECT 27.165 1.998 27.2 2.8 ;
      RECT 27.16 1.988 27.165 2.898 ;
      RECT 27.155 1.986 27.16 2.925 ;
      RECT 27.15 1.985 27.155 2.945 ;
      RECT 27.145 1.977 27.15 2.965 ;
      RECT 27.14 1.972 27.145 3 ;
      RECT 27.135 1.97 27.14 3.018 ;
      RECT 27.13 1.97 27.135 3.043 ;
      RECT 27.125 1.97 27.13 3.065 ;
      RECT 27.09 1.97 27.125 3.108 ;
      RECT 27.065 1.97 27.09 3.137 ;
      RECT 27.055 1.97 27.065 2.323 ;
      RECT 27.058 2.38 27.065 3.147 ;
      RECT 27.055 2.437 27.058 3.15 ;
      RECT 27.05 1.97 27.055 2.295 ;
      RECT 27.05 2.487 27.055 3.153 ;
      RECT 27.04 1.97 27.05 2.285 ;
      RECT 27.045 2.54 27.05 3.156 ;
      RECT 27.04 2.625 27.045 3.16 ;
      RECT 27.03 1.97 27.04 2.273 ;
      RECT 27.035 2.672 27.04 3.164 ;
      RECT 27.03 2.747 27.035 3.168 ;
      RECT 26.995 1.97 27.03 2.248 ;
      RECT 27.02 2.83 27.03 3.173 ;
      RECT 27.01 2.897 27.02 3.18 ;
      RECT 27.005 2.925 27.01 3.185 ;
      RECT 26.995 2.938 27.005 3.191 ;
      RECT 26.95 1.97 26.995 2.205 ;
      RECT 26.99 2.943 26.995 3.198 ;
      RECT 26.95 2.96 26.99 3.26 ;
      RECT 26.945 1.972 26.95 2.178 ;
      RECT 26.92 2.98 26.95 3.26 ;
      RECT 26.94 1.977 26.945 2.15 ;
      RECT 26.73 2.989 26.77 3.26 ;
      RECT 26.705 2.997 26.73 3.23 ;
      RECT 26.66 3.005 26.705 3.23 ;
      RECT 26.645 3.01 26.66 3.225 ;
      RECT 26.635 3.01 26.645 3.219 ;
      RECT 26.625 3.017 26.635 3.216 ;
      RECT 26.62 3.055 26.625 3.205 ;
      RECT 26.615 3.117 26.62 3.183 ;
      RECT 27.885 2.992 28.07 3.215 ;
      RECT 27.885 3.007 28.075 3.211 ;
      RECT 27.875 2.28 27.96 3.21 ;
      RECT 27.875 3.007 28.08 3.204 ;
      RECT 27.87 3.015 28.08 3.203 ;
      RECT 28.075 2.735 28.395 3.055 ;
      RECT 27.87 2.907 28.04 2.998 ;
      RECT 27.865 2.907 28.04 2.98 ;
      RECT 27.855 2.715 27.99 2.955 ;
      RECT 27.85 2.715 27.99 2.9 ;
      RECT 27.81 2.295 27.98 2.8 ;
      RECT 27.795 2.295 27.98 2.67 ;
      RECT 27.79 2.295 27.98 2.623 ;
      RECT 27.785 2.295 27.98 2.603 ;
      RECT 27.78 2.295 27.98 2.578 ;
      RECT 27.75 2.295 28.01 2.555 ;
      RECT 27.76 2.292 27.97 2.555 ;
      RECT 27.885 2.287 27.97 3.215 ;
      RECT 27.77 2.28 27.96 2.555 ;
      RECT 27.765 2.285 27.96 2.555 ;
      RECT 26.595 2.497 26.78 2.71 ;
      RECT 26.595 2.505 26.79 2.703 ;
      RECT 26.575 2.505 26.79 2.7 ;
      RECT 26.57 2.505 26.79 2.685 ;
      RECT 26.5 2.42 26.76 2.68 ;
      RECT 26.5 2.565 26.795 2.593 ;
      RECT 26.155 3.02 26.415 3.28 ;
      RECT 26.18 2.965 26.375 3.28 ;
      RECT 26.175 2.714 26.355 3.008 ;
      RECT 26.175 2.72 26.365 3.008 ;
      RECT 26.155 2.722 26.365 2.953 ;
      RECT 26.15 2.732 26.365 2.82 ;
      RECT 26.18 2.712 26.355 3.28 ;
      RECT 26.266 2.71 26.355 3.28 ;
      RECT 26.125 1.93 26.16 2.3 ;
      RECT 25.915 2.04 25.92 2.3 ;
      RECT 26.16 1.937 26.175 2.3 ;
      RECT 26.05 1.93 26.125 2.378 ;
      RECT 26.04 1.93 26.05 2.463 ;
      RECT 26.015 1.93 26.04 2.498 ;
      RECT 25.975 1.93 26.015 2.566 ;
      RECT 25.965 1.937 25.975 2.618 ;
      RECT 25.935 2.04 25.965 2.659 ;
      RECT 25.93 2.04 25.935 2.698 ;
      RECT 25.92 2.04 25.93 2.718 ;
      RECT 25.915 2.335 25.92 2.755 ;
      RECT 25.91 2.352 25.915 2.775 ;
      RECT 25.895 2.415 25.91 2.815 ;
      RECT 25.89 2.458 25.895 2.85 ;
      RECT 25.885 2.466 25.89 2.863 ;
      RECT 25.875 2.48 25.885 2.885 ;
      RECT 25.85 2.515 25.875 2.95 ;
      RECT 25.84 2.55 25.85 3.013 ;
      RECT 25.82 2.58 25.84 3.074 ;
      RECT 25.805 2.616 25.82 3.141 ;
      RECT 25.795 2.644 25.805 3.18 ;
      RECT 25.785 2.666 25.795 3.2 ;
      RECT 25.78 2.676 25.785 3.211 ;
      RECT 25.775 2.685 25.78 3.214 ;
      RECT 25.765 2.703 25.775 3.218 ;
      RECT 25.755 2.721 25.765 3.219 ;
      RECT 25.73 2.76 25.755 3.216 ;
      RECT 25.71 2.802 25.73 3.213 ;
      RECT 25.695 2.84 25.71 3.212 ;
      RECT 25.66 2.875 25.695 3.209 ;
      RECT 25.655 2.897 25.66 3.207 ;
      RECT 25.59 2.937 25.655 3.204 ;
      RECT 25.585 2.977 25.59 3.2 ;
      RECT 25.57 2.987 25.585 3.191 ;
      RECT 25.56 3.107 25.57 3.176 ;
      RECT 26.04 3.52 26.05 3.78 ;
      RECT 26.04 3.523 26.06 3.779 ;
      RECT 26.03 3.513 26.04 3.778 ;
      RECT 26.02 3.528 26.1 3.774 ;
      RECT 26.005 3.507 26.02 3.772 ;
      RECT 25.98 3.532 26.105 3.768 ;
      RECT 25.965 3.492 25.98 3.763 ;
      RECT 25.965 3.534 26.115 3.762 ;
      RECT 25.965 3.542 26.13 3.755 ;
      RECT 25.905 3.479 25.965 3.745 ;
      RECT 25.895 3.466 25.905 3.727 ;
      RECT 25.87 3.456 25.895 3.717 ;
      RECT 25.865 3.446 25.87 3.709 ;
      RECT 25.8 3.542 26.13 3.691 ;
      RECT 25.715 3.542 26.13 3.653 ;
      RECT 25.605 3.37 25.865 3.63 ;
      RECT 25.98 3.5 26.005 3.768 ;
      RECT 26.02 3.51 26.03 3.774 ;
      RECT 25.605 3.518 26.045 3.63 ;
      RECT 25.79 7.765 26.08 7.995 ;
      RECT 25.85 7.025 26.02 7.995 ;
      RECT 25.75 7.055 26.12 7.425 ;
      RECT 25.79 7.025 26.08 7.425 ;
      RECT 24.82 3.275 24.85 3.575 ;
      RECT 24.595 3.26 24.6 3.535 ;
      RECT 24.395 3.26 24.55 3.52 ;
      RECT 25.695 1.975 25.725 2.235 ;
      RECT 25.685 1.975 25.695 2.343 ;
      RECT 25.665 1.975 25.685 2.353 ;
      RECT 25.65 1.975 25.665 2.365 ;
      RECT 25.595 1.975 25.65 2.415 ;
      RECT 25.58 1.975 25.595 2.463 ;
      RECT 25.55 1.975 25.58 2.498 ;
      RECT 25.495 1.975 25.55 2.56 ;
      RECT 25.475 1.975 25.495 2.628 ;
      RECT 25.47 1.975 25.475 2.658 ;
      RECT 25.465 1.975 25.47 2.67 ;
      RECT 25.46 2.092 25.465 2.688 ;
      RECT 25.44 2.11 25.46 2.713 ;
      RECT 25.42 2.137 25.44 2.763 ;
      RECT 25.415 2.157 25.42 2.794 ;
      RECT 25.41 2.165 25.415 2.811 ;
      RECT 25.395 2.191 25.41 2.84 ;
      RECT 25.38 2.233 25.395 2.875 ;
      RECT 25.375 2.262 25.38 2.898 ;
      RECT 25.37 2.277 25.375 2.911 ;
      RECT 25.365 2.3 25.37 2.922 ;
      RECT 25.355 2.32 25.365 2.94 ;
      RECT 25.345 2.35 25.355 2.963 ;
      RECT 25.34 2.372 25.345 2.983 ;
      RECT 25.335 2.387 25.34 2.998 ;
      RECT 25.32 2.417 25.335 3.025 ;
      RECT 25.315 2.447 25.32 3.051 ;
      RECT 25.31 2.465 25.315 3.063 ;
      RECT 25.3 2.495 25.31 3.082 ;
      RECT 25.29 2.52 25.3 3.107 ;
      RECT 25.285 2.54 25.29 3.126 ;
      RECT 25.28 2.557 25.285 3.139 ;
      RECT 25.27 2.583 25.28 3.158 ;
      RECT 25.26 2.621 25.27 3.185 ;
      RECT 25.255 2.647 25.26 3.205 ;
      RECT 25.25 2.657 25.255 3.215 ;
      RECT 25.245 2.67 25.25 3.23 ;
      RECT 25.24 2.685 25.245 3.24 ;
      RECT 25.235 2.707 25.24 3.255 ;
      RECT 25.23 2.725 25.235 3.266 ;
      RECT 25.225 2.735 25.23 3.277 ;
      RECT 25.22 2.743 25.225 3.289 ;
      RECT 25.215 2.751 25.22 3.3 ;
      RECT 25.21 2.777 25.215 3.313 ;
      RECT 25.2 2.805 25.21 3.326 ;
      RECT 25.195 2.835 25.2 3.335 ;
      RECT 25.19 2.85 25.195 3.342 ;
      RECT 25.175 2.875 25.19 3.349 ;
      RECT 25.17 2.897 25.175 3.355 ;
      RECT 25.165 2.922 25.17 3.358 ;
      RECT 25.156 2.95 25.165 3.362 ;
      RECT 25.15 2.967 25.156 3.367 ;
      RECT 25.145 2.985 25.15 3.371 ;
      RECT 25.14 2.997 25.145 3.374 ;
      RECT 25.135 3.018 25.14 3.378 ;
      RECT 25.13 3.036 25.135 3.381 ;
      RECT 25.125 3.05 25.13 3.384 ;
      RECT 25.12 3.067 25.125 3.387 ;
      RECT 25.115 3.08 25.12 3.39 ;
      RECT 25.09 3.117 25.115 3.398 ;
      RECT 25.085 3.162 25.09 3.407 ;
      RECT 25.08 3.19 25.085 3.41 ;
      RECT 25.07 3.21 25.08 3.414 ;
      RECT 25.065 3.23 25.07 3.419 ;
      RECT 25.06 3.245 25.065 3.422 ;
      RECT 25.04 3.255 25.06 3.429 ;
      RECT 24.975 3.262 25.04 3.455 ;
      RECT 24.94 3.265 24.975 3.483 ;
      RECT 24.925 3.268 24.94 3.498 ;
      RECT 24.915 3.269 24.925 3.513 ;
      RECT 24.905 3.27 24.915 3.53 ;
      RECT 24.9 3.27 24.905 3.545 ;
      RECT 24.895 3.27 24.9 3.553 ;
      RECT 24.88 3.271 24.895 3.568 ;
      RECT 24.85 3.273 24.88 3.575 ;
      RECT 24.74 3.28 24.82 3.575 ;
      RECT 24.695 3.285 24.74 3.575 ;
      RECT 24.685 3.286 24.695 3.565 ;
      RECT 24.675 3.287 24.685 3.558 ;
      RECT 24.655 3.289 24.675 3.553 ;
      RECT 24.645 3.26 24.655 3.548 ;
      RECT 24.6 3.26 24.645 3.54 ;
      RECT 24.57 3.26 24.595 3.53 ;
      RECT 24.55 3.26 24.57 3.523 ;
      RECT 24.83 2.06 25.09 2.32 ;
      RECT 24.71 2.075 24.72 2.24 ;
      RECT 24.695 2.075 24.7 2.235 ;
      RECT 22.06 1.915 22.245 2.205 ;
      RECT 23.875 2.04 23.89 2.195 ;
      RECT 22.025 1.915 22.05 2.175 ;
      RECT 24.44 1.965 24.445 2.107 ;
      RECT 24.355 1.96 24.38 2.1 ;
      RECT 24.755 2.077 24.83 2.27 ;
      RECT 24.74 2.075 24.755 2.253 ;
      RECT 24.72 2.075 24.74 2.245 ;
      RECT 24.7 2.075 24.71 2.238 ;
      RECT 24.655 2.07 24.695 2.228 ;
      RECT 24.615 2.045 24.655 2.213 ;
      RECT 24.6 2.02 24.615 2.203 ;
      RECT 24.595 2.014 24.6 2.201 ;
      RECT 24.56 2.006 24.595 2.184 ;
      RECT 24.555 1.999 24.56 2.172 ;
      RECT 24.535 1.994 24.555 2.16 ;
      RECT 24.525 1.988 24.535 2.145 ;
      RECT 24.505 1.983 24.525 2.13 ;
      RECT 24.495 1.978 24.505 2.123 ;
      RECT 24.49 1.976 24.495 2.118 ;
      RECT 24.485 1.975 24.49 2.115 ;
      RECT 24.445 1.97 24.485 2.111 ;
      RECT 24.425 1.964 24.44 2.106 ;
      RECT 24.39 1.961 24.425 2.103 ;
      RECT 24.38 1.96 24.39 2.101 ;
      RECT 24.32 1.96 24.355 2.098 ;
      RECT 24.275 1.96 24.32 2.098 ;
      RECT 24.225 1.96 24.275 2.101 ;
      RECT 24.21 1.962 24.225 2.103 ;
      RECT 24.195 1.965 24.21 2.104 ;
      RECT 24.185 1.97 24.195 2.105 ;
      RECT 24.155 1.975 24.185 2.11 ;
      RECT 24.145 1.981 24.155 2.118 ;
      RECT 24.135 1.983 24.145 2.122 ;
      RECT 24.125 1.987 24.135 2.126 ;
      RECT 24.1 1.993 24.125 2.134 ;
      RECT 24.09 1.998 24.1 2.142 ;
      RECT 24.075 2.002 24.09 2.146 ;
      RECT 24.04 2.008 24.075 2.154 ;
      RECT 24.02 2.013 24.04 2.164 ;
      RECT 23.99 2.02 24.02 2.173 ;
      RECT 23.945 2.029 23.99 2.187 ;
      RECT 23.94 2.034 23.945 2.198 ;
      RECT 23.92 2.037 23.94 2.199 ;
      RECT 23.89 2.04 23.92 2.197 ;
      RECT 23.855 2.04 23.875 2.193 ;
      RECT 23.785 2.04 23.855 2.184 ;
      RECT 23.77 2.037 23.785 2.176 ;
      RECT 23.73 2.03 23.77 2.171 ;
      RECT 23.705 2.02 23.73 2.164 ;
      RECT 23.7 2.014 23.705 2.161 ;
      RECT 23.66 2.008 23.7 2.158 ;
      RECT 23.645 2.001 23.66 2.153 ;
      RECT 23.625 1.997 23.645 2.148 ;
      RECT 23.61 1.992 23.625 2.144 ;
      RECT 23.595 1.987 23.61 2.142 ;
      RECT 23.58 1.983 23.595 2.141 ;
      RECT 23.565 1.981 23.58 2.137 ;
      RECT 23.555 1.979 23.565 2.132 ;
      RECT 23.54 1.976 23.555 2.128 ;
      RECT 23.53 1.974 23.54 2.123 ;
      RECT 23.51 1.971 23.53 2.119 ;
      RECT 23.465 1.97 23.51 2.117 ;
      RECT 23.405 1.972 23.465 2.118 ;
      RECT 23.385 1.974 23.405 2.12 ;
      RECT 23.355 1.977 23.385 2.121 ;
      RECT 23.305 1.982 23.355 2.123 ;
      RECT 23.3 1.985 23.305 2.125 ;
      RECT 23.29 1.987 23.3 2.128 ;
      RECT 23.285 1.989 23.29 2.131 ;
      RECT 23.235 1.992 23.285 2.138 ;
      RECT 23.215 1.996 23.235 2.15 ;
      RECT 23.205 1.999 23.215 2.156 ;
      RECT 23.195 2 23.205 2.159 ;
      RECT 23.156 2.003 23.195 2.161 ;
      RECT 23.07 2.01 23.156 2.164 ;
      RECT 22.996 2.02 23.07 2.168 ;
      RECT 22.91 2.031 22.996 2.173 ;
      RECT 22.895 2.038 22.91 2.175 ;
      RECT 22.84 2.042 22.895 2.176 ;
      RECT 22.826 2.045 22.84 2.178 ;
      RECT 22.74 2.045 22.826 2.18 ;
      RECT 22.7 2.042 22.74 2.183 ;
      RECT 22.676 2.038 22.7 2.185 ;
      RECT 22.59 2.028 22.676 2.188 ;
      RECT 22.56 2.017 22.59 2.189 ;
      RECT 22.541 2.013 22.56 2.188 ;
      RECT 22.455 2.006 22.541 2.185 ;
      RECT 22.395 1.995 22.455 2.182 ;
      RECT 22.375 1.987 22.395 2.18 ;
      RECT 22.34 1.982 22.375 2.179 ;
      RECT 22.315 1.977 22.34 2.178 ;
      RECT 22.285 1.972 22.315 2.177 ;
      RECT 22.26 1.915 22.285 2.176 ;
      RECT 22.245 1.915 22.26 2.2 ;
      RECT 22.05 1.915 22.06 2.2 ;
      RECT 23.825 2.935 23.83 3.075 ;
      RECT 23.485 2.935 23.52 3.073 ;
      RECT 23.06 2.92 23.075 3.065 ;
      RECT 24.89 2.7 24.98 2.96 ;
      RECT 24.72 2.565 24.82 2.96 ;
      RECT 21.755 2.54 21.835 2.75 ;
      RECT 24.845 2.677 24.89 2.96 ;
      RECT 24.835 2.647 24.845 2.96 ;
      RECT 24.82 2.57 24.835 2.96 ;
      RECT 24.635 2.565 24.72 2.925 ;
      RECT 24.63 2.567 24.635 2.92 ;
      RECT 24.625 2.572 24.63 2.92 ;
      RECT 24.59 2.672 24.625 2.92 ;
      RECT 24.58 2.7 24.59 2.92 ;
      RECT 24.57 2.715 24.58 2.92 ;
      RECT 24.56 2.727 24.57 2.92 ;
      RECT 24.555 2.737 24.56 2.92 ;
      RECT 24.54 2.747 24.555 2.922 ;
      RECT 24.535 2.762 24.54 2.924 ;
      RECT 24.52 2.775 24.535 2.926 ;
      RECT 24.515 2.79 24.52 2.929 ;
      RECT 24.495 2.8 24.515 2.933 ;
      RECT 24.48 2.81 24.495 2.936 ;
      RECT 24.445 2.817 24.48 2.941 ;
      RECT 24.401 2.824 24.445 2.949 ;
      RECT 24.315 2.836 24.401 2.962 ;
      RECT 24.29 2.847 24.315 2.973 ;
      RECT 24.26 2.852 24.29 2.978 ;
      RECT 24.225 2.857 24.26 2.986 ;
      RECT 24.195 2.862 24.225 2.993 ;
      RECT 24.17 2.867 24.195 2.998 ;
      RECT 24.105 2.874 24.17 3.007 ;
      RECT 24.035 2.887 24.105 3.023 ;
      RECT 24.005 2.897 24.035 3.035 ;
      RECT 23.98 2.902 24.005 3.042 ;
      RECT 23.925 2.909 23.98 3.05 ;
      RECT 23.92 2.916 23.925 3.055 ;
      RECT 23.915 2.918 23.92 3.056 ;
      RECT 23.9 2.92 23.915 3.058 ;
      RECT 23.895 2.92 23.9 3.061 ;
      RECT 23.83 2.927 23.895 3.068 ;
      RECT 23.795 2.937 23.825 3.078 ;
      RECT 23.778 2.94 23.795 3.08 ;
      RECT 23.692 2.939 23.778 3.079 ;
      RECT 23.606 2.937 23.692 3.076 ;
      RECT 23.52 2.936 23.606 3.074 ;
      RECT 23.419 2.934 23.485 3.073 ;
      RECT 23.333 2.931 23.419 3.071 ;
      RECT 23.247 2.927 23.333 3.069 ;
      RECT 23.161 2.924 23.247 3.068 ;
      RECT 23.075 2.921 23.161 3.066 ;
      RECT 22.975 2.92 23.06 3.063 ;
      RECT 22.925 2.918 22.975 3.061 ;
      RECT 22.905 2.915 22.925 3.059 ;
      RECT 22.885 2.913 22.905 3.056 ;
      RECT 22.86 2.909 22.885 3.053 ;
      RECT 22.815 2.903 22.86 3.048 ;
      RECT 22.775 2.897 22.815 3.04 ;
      RECT 22.75 2.892 22.775 3.033 ;
      RECT 22.695 2.885 22.75 3.025 ;
      RECT 22.671 2.878 22.695 3.018 ;
      RECT 22.585 2.869 22.671 3.008 ;
      RECT 22.555 2.861 22.585 2.998 ;
      RECT 22.525 2.857 22.555 2.993 ;
      RECT 22.52 2.854 22.525 2.99 ;
      RECT 22.515 2.853 22.52 2.99 ;
      RECT 22.44 2.846 22.515 2.983 ;
      RECT 22.401 2.837 22.44 2.972 ;
      RECT 22.315 2.827 22.401 2.96 ;
      RECT 22.275 2.817 22.315 2.948 ;
      RECT 22.236 2.812 22.275 2.941 ;
      RECT 22.15 2.802 22.236 2.93 ;
      RECT 22.11 2.79 22.15 2.919 ;
      RECT 22.075 2.775 22.11 2.912 ;
      RECT 22.065 2.765 22.075 2.909 ;
      RECT 22.045 2.75 22.065 2.907 ;
      RECT 22.015 2.72 22.045 2.903 ;
      RECT 22.005 2.7 22.015 2.898 ;
      RECT 22 2.692 22.005 2.895 ;
      RECT 21.995 2.685 22 2.893 ;
      RECT 21.98 2.672 21.995 2.886 ;
      RECT 21.975 2.662 21.98 2.878 ;
      RECT 21.97 2.655 21.975 2.873 ;
      RECT 21.965 2.65 21.97 2.869 ;
      RECT 21.95 2.637 21.965 2.861 ;
      RECT 21.945 2.547 21.95 2.85 ;
      RECT 21.94 2.542 21.945 2.843 ;
      RECT 21.865 2.54 21.94 2.803 ;
      RECT 21.835 2.54 21.865 2.758 ;
      RECT 21.74 2.545 21.755 2.745 ;
      RECT 24.225 2.25 24.485 2.51 ;
      RECT 24.21 2.238 24.39 2.475 ;
      RECT 24.205 2.239 24.39 2.473 ;
      RECT 24.19 2.243 24.4 2.463 ;
      RECT 24.185 2.248 24.405 2.433 ;
      RECT 24.19 2.245 24.405 2.463 ;
      RECT 24.205 2.24 24.4 2.473 ;
      RECT 24.225 2.237 24.39 2.51 ;
      RECT 24.225 2.236 24.38 2.51 ;
      RECT 24.25 2.235 24.38 2.51 ;
      RECT 23.81 2.48 24.07 2.74 ;
      RECT 23.685 2.525 24.07 2.735 ;
      RECT 23.675 2.53 24.07 2.73 ;
      RECT 23.69 3.47 23.705 3.78 ;
      RECT 22.285 3.24 22.295 3.37 ;
      RECT 22.065 3.235 22.17 3.37 ;
      RECT 21.98 3.24 22.03 3.37 ;
      RECT 20.53 1.975 20.535 3.08 ;
      RECT 23.785 3.562 23.79 3.698 ;
      RECT 23.78 3.557 23.785 3.758 ;
      RECT 23.775 3.555 23.78 3.771 ;
      RECT 23.76 3.552 23.775 3.773 ;
      RECT 23.755 3.547 23.76 3.775 ;
      RECT 23.75 3.543 23.755 3.778 ;
      RECT 23.735 3.538 23.75 3.78 ;
      RECT 23.705 3.53 23.735 3.78 ;
      RECT 23.666 3.47 23.69 3.78 ;
      RECT 23.58 3.47 23.666 3.777 ;
      RECT 23.55 3.47 23.58 3.77 ;
      RECT 23.525 3.47 23.55 3.763 ;
      RECT 23.5 3.47 23.525 3.755 ;
      RECT 23.485 3.47 23.5 3.748 ;
      RECT 23.46 3.47 23.485 3.74 ;
      RECT 23.445 3.47 23.46 3.733 ;
      RECT 23.405 3.48 23.445 3.722 ;
      RECT 23.395 3.475 23.405 3.712 ;
      RECT 23.391 3.474 23.395 3.709 ;
      RECT 23.305 3.466 23.391 3.692 ;
      RECT 23.272 3.455 23.305 3.669 ;
      RECT 23.186 3.444 23.272 3.647 ;
      RECT 23.1 3.428 23.186 3.616 ;
      RECT 23.03 3.413 23.1 3.588 ;
      RECT 23.02 3.406 23.03 3.575 ;
      RECT 22.99 3.403 23.02 3.565 ;
      RECT 22.965 3.399 22.99 3.558 ;
      RECT 22.95 3.396 22.965 3.553 ;
      RECT 22.945 3.395 22.95 3.548 ;
      RECT 22.915 3.39 22.945 3.541 ;
      RECT 22.91 3.385 22.915 3.536 ;
      RECT 22.895 3.382 22.91 3.531 ;
      RECT 22.89 3.377 22.895 3.526 ;
      RECT 22.87 3.372 22.89 3.523 ;
      RECT 22.855 3.367 22.87 3.515 ;
      RECT 22.84 3.361 22.855 3.51 ;
      RECT 22.81 3.352 22.84 3.503 ;
      RECT 22.805 3.345 22.81 3.495 ;
      RECT 22.8 3.343 22.805 3.493 ;
      RECT 22.795 3.342 22.8 3.49 ;
      RECT 22.755 3.335 22.795 3.483 ;
      RECT 22.741 3.325 22.755 3.473 ;
      RECT 22.69 3.314 22.741 3.461 ;
      RECT 22.665 3.3 22.69 3.447 ;
      RECT 22.64 3.289 22.665 3.439 ;
      RECT 22.62 3.278 22.64 3.433 ;
      RECT 22.61 3.272 22.62 3.428 ;
      RECT 22.605 3.27 22.61 3.424 ;
      RECT 22.585 3.265 22.605 3.419 ;
      RECT 22.555 3.255 22.585 3.409 ;
      RECT 22.55 3.247 22.555 3.402 ;
      RECT 22.535 3.245 22.55 3.398 ;
      RECT 22.515 3.245 22.535 3.393 ;
      RECT 22.51 3.244 22.515 3.391 ;
      RECT 22.505 3.244 22.51 3.388 ;
      RECT 22.465 3.243 22.505 3.383 ;
      RECT 22.44 3.242 22.465 3.378 ;
      RECT 22.38 3.241 22.44 3.375 ;
      RECT 22.295 3.24 22.38 3.373 ;
      RECT 22.256 3.239 22.285 3.37 ;
      RECT 22.17 3.237 22.256 3.37 ;
      RECT 22.03 3.237 22.065 3.37 ;
      RECT 21.94 3.241 21.98 3.373 ;
      RECT 21.925 3.244 21.94 3.38 ;
      RECT 21.915 3.245 21.925 3.387 ;
      RECT 21.89 3.248 21.915 3.392 ;
      RECT 21.885 3.25 21.89 3.395 ;
      RECT 21.835 3.252 21.885 3.396 ;
      RECT 21.796 3.256 21.835 3.398 ;
      RECT 21.71 3.258 21.796 3.401 ;
      RECT 21.692 3.26 21.71 3.403 ;
      RECT 21.606 3.263 21.692 3.405 ;
      RECT 21.52 3.267 21.606 3.408 ;
      RECT 21.483 3.271 21.52 3.411 ;
      RECT 21.397 3.274 21.483 3.414 ;
      RECT 21.311 3.278 21.397 3.417 ;
      RECT 21.225 3.283 21.311 3.421 ;
      RECT 21.205 3.285 21.225 3.424 ;
      RECT 21.185 3.284 21.205 3.425 ;
      RECT 21.136 3.281 21.185 3.426 ;
      RECT 21.05 3.276 21.136 3.429 ;
      RECT 21 3.271 21.05 3.431 ;
      RECT 20.976 3.269 21 3.432 ;
      RECT 20.89 3.264 20.976 3.434 ;
      RECT 20.865 3.26 20.89 3.433 ;
      RECT 20.855 3.257 20.865 3.431 ;
      RECT 20.845 3.25 20.855 3.428 ;
      RECT 20.84 3.23 20.845 3.423 ;
      RECT 20.83 3.2 20.84 3.418 ;
      RECT 20.815 3.07 20.83 3.409 ;
      RECT 20.81 3.062 20.815 3.402 ;
      RECT 20.79 3.055 20.81 3.394 ;
      RECT 20.785 3.037 20.79 3.386 ;
      RECT 20.775 3.017 20.785 3.381 ;
      RECT 20.77 2.99 20.775 3.377 ;
      RECT 20.765 2.967 20.77 3.374 ;
      RECT 20.745 2.925 20.765 3.366 ;
      RECT 20.71 2.84 20.745 3.35 ;
      RECT 20.705 2.772 20.71 3.338 ;
      RECT 20.69 2.742 20.705 3.332 ;
      RECT 20.685 1.987 20.69 2.233 ;
      RECT 20.675 2.712 20.69 3.323 ;
      RECT 20.68 1.982 20.685 2.265 ;
      RECT 20.675 1.977 20.68 2.308 ;
      RECT 20.67 1.975 20.675 2.343 ;
      RECT 20.655 2.675 20.675 3.313 ;
      RECT 20.665 1.975 20.67 2.38 ;
      RECT 20.65 1.975 20.665 2.478 ;
      RECT 20.65 2.648 20.655 3.306 ;
      RECT 20.645 1.975 20.65 2.553 ;
      RECT 20.645 2.636 20.65 3.303 ;
      RECT 20.64 1.975 20.645 2.585 ;
      RECT 20.64 2.615 20.645 3.3 ;
      RECT 20.635 1.975 20.64 3.297 ;
      RECT 20.6 1.975 20.635 3.283 ;
      RECT 20.585 1.975 20.6 3.265 ;
      RECT 20.565 1.975 20.585 3.255 ;
      RECT 20.54 1.975 20.565 3.238 ;
      RECT 20.535 1.975 20.54 3.188 ;
      RECT 20.525 1.975 20.53 3.018 ;
      RECT 20.52 1.975 20.525 2.925 ;
      RECT 20.515 1.975 20.52 2.838 ;
      RECT 20.51 1.975 20.515 2.77 ;
      RECT 20.505 1.975 20.51 2.713 ;
      RECT 20.495 1.975 20.505 2.608 ;
      RECT 20.49 1.975 20.495 2.48 ;
      RECT 20.485 1.975 20.49 2.398 ;
      RECT 20.48 1.977 20.485 2.315 ;
      RECT 20.475 1.982 20.48 2.248 ;
      RECT 20.47 1.987 20.475 2.175 ;
      RECT 23.285 2.305 23.545 2.565 ;
      RECT 23.305 2.272 23.515 2.565 ;
      RECT 23.305 2.27 23.505 2.565 ;
      RECT 23.315 2.257 23.505 2.565 ;
      RECT 23.315 2.255 23.43 2.565 ;
      RECT 22.79 2.38 22.965 2.66 ;
      RECT 22.785 2.38 22.965 2.658 ;
      RECT 22.785 2.38 22.98 2.655 ;
      RECT 22.775 2.38 22.98 2.653 ;
      RECT 22.72 2.38 22.98 2.64 ;
      RECT 22.72 2.455 22.985 2.618 ;
      RECT 22.265 2.392 22.285 2.635 ;
      RECT 22.265 2.392 22.325 2.634 ;
      RECT 22.26 2.394 22.325 2.633 ;
      RECT 22.26 2.394 22.411 2.632 ;
      RECT 22.26 2.394 22.48 2.631 ;
      RECT 22.26 2.394 22.5 2.623 ;
      RECT 22.24 2.397 22.5 2.621 ;
      RECT 22.225 2.407 22.5 2.606 ;
      RECT 22.225 2.407 22.515 2.605 ;
      RECT 22.22 2.416 22.515 2.597 ;
      RECT 22.22 2.416 22.52 2.593 ;
      RECT 22.325 2.33 22.585 2.59 ;
      RECT 22.215 2.418 22.585 2.475 ;
      RECT 22.285 2.385 22.585 2.59 ;
      RECT 22.25 3.578 22.255 3.785 ;
      RECT 22.2 3.572 22.25 3.784 ;
      RECT 22.167 3.586 22.26 3.783 ;
      RECT 22.081 3.586 22.26 3.782 ;
      RECT 21.995 3.586 22.26 3.781 ;
      RECT 21.995 3.685 22.265 3.778 ;
      RECT 21.99 3.685 22.265 3.773 ;
      RECT 21.985 3.685 22.265 3.755 ;
      RECT 21.98 3.685 22.265 3.738 ;
      RECT 21.94 3.47 22.2 3.73 ;
      RECT 21.4 2.62 21.486 3.034 ;
      RECT 21.4 2.62 21.525 3.031 ;
      RECT 21.4 2.62 21.545 3.021 ;
      RECT 21.355 2.62 21.545 3.018 ;
      RECT 21.355 2.772 21.555 3.008 ;
      RECT 21.355 2.793 21.56 3.002 ;
      RECT 21.355 2.811 21.565 2.998 ;
      RECT 21.355 2.831 21.575 2.993 ;
      RECT 21.33 2.831 21.575 2.99 ;
      RECT 21.32 2.831 21.575 2.968 ;
      RECT 21.32 2.847 21.58 2.938 ;
      RECT 21.285 2.62 21.545 2.925 ;
      RECT 21.285 2.859 21.585 2.88 ;
      RECT 18.945 7.77 19.235 8 ;
      RECT 19.005 6.29 19.175 8 ;
      RECT 19 6.655 19.35 7.005 ;
      RECT 18.945 6.29 19.235 6.52 ;
      RECT 18.54 2.395 18.645 2.965 ;
      RECT 18.54 2.73 18.865 2.96 ;
      RECT 18.54 2.76 19.035 2.93 ;
      RECT 18.54 2.395 18.73 2.96 ;
      RECT 17.955 2.36 18.245 2.59 ;
      RECT 17.955 2.395 18.73 2.565 ;
      RECT 18.015 0.88 18.185 2.59 ;
      RECT 17.955 0.88 18.245 1.11 ;
      RECT 17.955 7.77 18.245 8 ;
      RECT 18.015 6.29 18.185 8 ;
      RECT 17.955 6.29 18.245 6.52 ;
      RECT 17.955 6.325 18.81 6.485 ;
      RECT 18.64 5.92 18.81 6.485 ;
      RECT 17.955 6.32 18.35 6.485 ;
      RECT 18.575 5.92 18.865 6.15 ;
      RECT 18.575 5.95 19.035 6.12 ;
      RECT 17.585 2.73 17.875 2.96 ;
      RECT 17.585 2.76 18.045 2.93 ;
      RECT 17.65 1.655 17.815 2.96 ;
      RECT 16.165 1.625 16.455 1.855 ;
      RECT 16.165 1.655 17.815 1.825 ;
      RECT 16.225 0.885 16.395 1.855 ;
      RECT 16.165 0.885 16.455 1.115 ;
      RECT 16.165 7.765 16.455 7.995 ;
      RECT 16.225 7.025 16.395 7.995 ;
      RECT 16.225 7.12 17.815 7.29 ;
      RECT 17.645 5.92 17.815 7.29 ;
      RECT 16.165 7.025 16.455 7.255 ;
      RECT 17.585 5.92 17.875 6.15 ;
      RECT 17.585 5.95 18.045 6.12 ;
      RECT 14.215 2.705 14.555 3.055 ;
      RECT 14.305 2.025 14.475 3.055 ;
      RECT 16.595 1.965 16.945 2.315 ;
      RECT 14.305 2.025 16.945 2.195 ;
      RECT 16.62 6.655 16.945 6.98 ;
      RECT 11.16 6.605 11.51 6.955 ;
      RECT 16.595 6.655 16.945 6.885 ;
      RECT 10.96 6.655 11.51 6.885 ;
      RECT 10.79 6.685 16.945 6.855 ;
      RECT 15.82 2.365 16.14 2.685 ;
      RECT 15.79 2.365 16.14 2.595 ;
      RECT 15.62 2.395 16.14 2.565 ;
      RECT 15.82 6.255 16.14 6.545 ;
      RECT 15.79 6.285 16.14 6.515 ;
      RECT 15.62 6.315 16.14 6.485 ;
      RECT 11.51 2.985 11.66 3.26 ;
      RECT 12.05 2.065 12.055 2.285 ;
      RECT 13.2 2.265 13.215 2.463 ;
      RECT 13.165 2.257 13.2 2.47 ;
      RECT 13.135 2.25 13.165 2.47 ;
      RECT 13.08 2.215 13.135 2.47 ;
      RECT 13.015 2.152 13.08 2.47 ;
      RECT 13.01 2.117 13.015 2.468 ;
      RECT 13.005 2.112 13.01 2.46 ;
      RECT 13 2.107 13.005 2.446 ;
      RECT 12.995 2.104 13 2.439 ;
      RECT 12.95 2.094 12.995 2.39 ;
      RECT 12.93 2.081 12.95 2.325 ;
      RECT 12.925 2.076 12.93 2.298 ;
      RECT 12.92 2.075 12.925 2.291 ;
      RECT 12.915 2.074 12.92 2.284 ;
      RECT 12.83 2.059 12.915 2.23 ;
      RECT 12.8 2.04 12.83 2.18 ;
      RECT 12.72 2.023 12.8 2.165 ;
      RECT 12.685 2.01 12.72 2.15 ;
      RECT 12.677 2.01 12.685 2.145 ;
      RECT 12.591 2.011 12.677 2.145 ;
      RECT 12.505 2.013 12.591 2.145 ;
      RECT 12.48 2.014 12.505 2.149 ;
      RECT 12.405 2.02 12.48 2.164 ;
      RECT 12.322 2.032 12.405 2.188 ;
      RECT 12.236 2.045 12.322 2.214 ;
      RECT 12.15 2.058 12.236 2.24 ;
      RECT 12.115 2.067 12.15 2.259 ;
      RECT 12.065 2.067 12.115 2.272 ;
      RECT 12.055 2.065 12.065 2.283 ;
      RECT 12.04 2.062 12.05 2.285 ;
      RECT 12.025 2.054 12.04 2.293 ;
      RECT 12.01 2.046 12.025 2.313 ;
      RECT 12.005 2.041 12.01 2.37 ;
      RECT 11.99 2.036 12.005 2.443 ;
      RECT 11.985 2.031 11.99 2.485 ;
      RECT 11.98 2.029 11.985 2.513 ;
      RECT 11.975 2.027 11.98 2.535 ;
      RECT 11.965 2.023 11.975 2.578 ;
      RECT 11.96 2.02 11.965 2.603 ;
      RECT 11.955 2.018 11.96 2.623 ;
      RECT 11.95 2.016 11.955 2.647 ;
      RECT 11.945 2.012 11.95 2.67 ;
      RECT 11.94 2.008 11.945 2.693 ;
      RECT 11.905 1.998 11.94 2.8 ;
      RECT 11.9 1.988 11.905 2.898 ;
      RECT 11.895 1.986 11.9 2.925 ;
      RECT 11.89 1.985 11.895 2.945 ;
      RECT 11.885 1.977 11.89 2.965 ;
      RECT 11.88 1.972 11.885 3 ;
      RECT 11.875 1.97 11.88 3.018 ;
      RECT 11.87 1.97 11.875 3.043 ;
      RECT 11.865 1.97 11.87 3.065 ;
      RECT 11.83 1.97 11.865 3.108 ;
      RECT 11.805 1.97 11.83 3.137 ;
      RECT 11.795 1.97 11.805 2.323 ;
      RECT 11.798 2.38 11.805 3.147 ;
      RECT 11.795 2.437 11.798 3.15 ;
      RECT 11.79 1.97 11.795 2.295 ;
      RECT 11.79 2.487 11.795 3.153 ;
      RECT 11.78 1.97 11.79 2.285 ;
      RECT 11.785 2.54 11.79 3.156 ;
      RECT 11.78 2.625 11.785 3.16 ;
      RECT 11.77 1.97 11.78 2.273 ;
      RECT 11.775 2.672 11.78 3.164 ;
      RECT 11.77 2.747 11.775 3.168 ;
      RECT 11.735 1.97 11.77 2.248 ;
      RECT 11.76 2.83 11.77 3.173 ;
      RECT 11.75 2.897 11.76 3.18 ;
      RECT 11.745 2.925 11.75 3.185 ;
      RECT 11.735 2.938 11.745 3.191 ;
      RECT 11.69 1.97 11.735 2.205 ;
      RECT 11.73 2.943 11.735 3.198 ;
      RECT 11.69 2.96 11.73 3.26 ;
      RECT 11.685 1.972 11.69 2.178 ;
      RECT 11.66 2.98 11.69 3.26 ;
      RECT 11.68 1.977 11.685 2.15 ;
      RECT 11.47 2.989 11.51 3.26 ;
      RECT 11.445 2.997 11.47 3.23 ;
      RECT 11.4 3.005 11.445 3.23 ;
      RECT 11.385 3.01 11.4 3.225 ;
      RECT 11.375 3.01 11.385 3.219 ;
      RECT 11.365 3.017 11.375 3.216 ;
      RECT 11.36 3.055 11.365 3.205 ;
      RECT 11.355 3.117 11.36 3.183 ;
      RECT 12.625 2.992 12.81 3.215 ;
      RECT 12.625 3.007 12.815 3.211 ;
      RECT 12.615 2.28 12.7 3.21 ;
      RECT 12.615 3.007 12.82 3.204 ;
      RECT 12.61 3.015 12.82 3.203 ;
      RECT 12.815 2.735 13.135 3.055 ;
      RECT 12.61 2.907 12.78 2.998 ;
      RECT 12.605 2.907 12.78 2.98 ;
      RECT 12.595 2.715 12.73 2.955 ;
      RECT 12.59 2.715 12.73 2.9 ;
      RECT 12.55 2.295 12.72 2.8 ;
      RECT 12.535 2.295 12.72 2.67 ;
      RECT 12.53 2.295 12.72 2.623 ;
      RECT 12.525 2.295 12.72 2.603 ;
      RECT 12.52 2.295 12.72 2.578 ;
      RECT 12.49 2.295 12.75 2.555 ;
      RECT 12.5 2.292 12.71 2.555 ;
      RECT 12.625 2.287 12.71 3.215 ;
      RECT 12.51 2.28 12.7 2.555 ;
      RECT 12.505 2.285 12.7 2.555 ;
      RECT 11.335 2.497 11.52 2.71 ;
      RECT 11.335 2.505 11.53 2.703 ;
      RECT 11.315 2.505 11.53 2.7 ;
      RECT 11.31 2.505 11.53 2.685 ;
      RECT 11.24 2.42 11.5 2.68 ;
      RECT 11.24 2.565 11.535 2.593 ;
      RECT 10.895 3.02 11.155 3.28 ;
      RECT 10.92 2.965 11.115 3.28 ;
      RECT 10.915 2.714 11.095 3.008 ;
      RECT 10.915 2.72 11.105 3.008 ;
      RECT 10.895 2.722 11.105 2.953 ;
      RECT 10.89 2.732 11.105 2.82 ;
      RECT 10.92 2.712 11.095 3.28 ;
      RECT 11.006 2.71 11.095 3.28 ;
      RECT 10.865 1.93 10.9 2.3 ;
      RECT 10.655 2.04 10.66 2.3 ;
      RECT 10.9 1.937 10.915 2.3 ;
      RECT 10.79 1.93 10.865 2.378 ;
      RECT 10.78 1.93 10.79 2.463 ;
      RECT 10.755 1.93 10.78 2.498 ;
      RECT 10.715 1.93 10.755 2.566 ;
      RECT 10.705 1.937 10.715 2.618 ;
      RECT 10.675 2.04 10.705 2.659 ;
      RECT 10.67 2.04 10.675 2.698 ;
      RECT 10.66 2.04 10.67 2.718 ;
      RECT 10.655 2.335 10.66 2.755 ;
      RECT 10.65 2.352 10.655 2.775 ;
      RECT 10.635 2.415 10.65 2.815 ;
      RECT 10.63 2.458 10.635 2.85 ;
      RECT 10.625 2.466 10.63 2.863 ;
      RECT 10.615 2.48 10.625 2.885 ;
      RECT 10.59 2.515 10.615 2.95 ;
      RECT 10.58 2.55 10.59 3.013 ;
      RECT 10.56 2.58 10.58 3.074 ;
      RECT 10.545 2.616 10.56 3.141 ;
      RECT 10.535 2.644 10.545 3.18 ;
      RECT 10.525 2.666 10.535 3.2 ;
      RECT 10.52 2.676 10.525 3.211 ;
      RECT 10.515 2.685 10.52 3.214 ;
      RECT 10.505 2.703 10.515 3.218 ;
      RECT 10.495 2.721 10.505 3.219 ;
      RECT 10.47 2.76 10.495 3.216 ;
      RECT 10.45 2.802 10.47 3.213 ;
      RECT 10.435 2.84 10.45 3.212 ;
      RECT 10.4 2.875 10.435 3.209 ;
      RECT 10.395 2.897 10.4 3.207 ;
      RECT 10.33 2.937 10.395 3.204 ;
      RECT 10.325 2.977 10.33 3.2 ;
      RECT 10.31 2.987 10.325 3.191 ;
      RECT 10.3 3.107 10.31 3.176 ;
      RECT 10.78 3.52 10.79 3.78 ;
      RECT 10.78 3.523 10.8 3.779 ;
      RECT 10.77 3.513 10.78 3.778 ;
      RECT 10.76 3.528 10.84 3.774 ;
      RECT 10.745 3.507 10.76 3.772 ;
      RECT 10.72 3.532 10.845 3.768 ;
      RECT 10.705 3.492 10.72 3.763 ;
      RECT 10.705 3.534 10.855 3.762 ;
      RECT 10.705 3.542 10.87 3.755 ;
      RECT 10.645 3.479 10.705 3.745 ;
      RECT 10.635 3.466 10.645 3.727 ;
      RECT 10.61 3.456 10.635 3.717 ;
      RECT 10.605 3.446 10.61 3.709 ;
      RECT 10.54 3.542 10.87 3.691 ;
      RECT 10.455 3.542 10.87 3.653 ;
      RECT 10.345 3.37 10.605 3.63 ;
      RECT 10.72 3.5 10.745 3.768 ;
      RECT 10.76 3.51 10.77 3.774 ;
      RECT 10.345 3.518 10.785 3.63 ;
      RECT 10.53 7.765 10.82 7.995 ;
      RECT 10.59 7.025 10.76 7.995 ;
      RECT 10.49 7.055 10.86 7.425 ;
      RECT 10.53 7.025 10.82 7.425 ;
      RECT 9.56 3.275 9.59 3.575 ;
      RECT 9.335 3.26 9.34 3.535 ;
      RECT 9.135 3.26 9.29 3.52 ;
      RECT 10.435 1.975 10.465 2.235 ;
      RECT 10.425 1.975 10.435 2.343 ;
      RECT 10.405 1.975 10.425 2.353 ;
      RECT 10.39 1.975 10.405 2.365 ;
      RECT 10.335 1.975 10.39 2.415 ;
      RECT 10.32 1.975 10.335 2.463 ;
      RECT 10.29 1.975 10.32 2.498 ;
      RECT 10.235 1.975 10.29 2.56 ;
      RECT 10.215 1.975 10.235 2.628 ;
      RECT 10.21 1.975 10.215 2.658 ;
      RECT 10.205 1.975 10.21 2.67 ;
      RECT 10.2 2.092 10.205 2.688 ;
      RECT 10.18 2.11 10.2 2.713 ;
      RECT 10.16 2.137 10.18 2.763 ;
      RECT 10.155 2.157 10.16 2.794 ;
      RECT 10.15 2.165 10.155 2.811 ;
      RECT 10.135 2.191 10.15 2.84 ;
      RECT 10.12 2.233 10.135 2.875 ;
      RECT 10.115 2.262 10.12 2.898 ;
      RECT 10.11 2.277 10.115 2.911 ;
      RECT 10.105 2.3 10.11 2.922 ;
      RECT 10.095 2.32 10.105 2.94 ;
      RECT 10.085 2.35 10.095 2.963 ;
      RECT 10.08 2.372 10.085 2.983 ;
      RECT 10.075 2.387 10.08 2.998 ;
      RECT 10.06 2.417 10.075 3.025 ;
      RECT 10.055 2.447 10.06 3.051 ;
      RECT 10.05 2.465 10.055 3.063 ;
      RECT 10.04 2.495 10.05 3.082 ;
      RECT 10.03 2.52 10.04 3.107 ;
      RECT 10.025 2.54 10.03 3.126 ;
      RECT 10.02 2.557 10.025 3.139 ;
      RECT 10.01 2.583 10.02 3.158 ;
      RECT 10 2.621 10.01 3.185 ;
      RECT 9.995 2.647 10 3.205 ;
      RECT 9.99 2.657 9.995 3.215 ;
      RECT 9.985 2.67 9.99 3.23 ;
      RECT 9.98 2.685 9.985 3.24 ;
      RECT 9.975 2.707 9.98 3.255 ;
      RECT 9.97 2.725 9.975 3.266 ;
      RECT 9.965 2.735 9.97 3.277 ;
      RECT 9.96 2.743 9.965 3.289 ;
      RECT 9.955 2.751 9.96 3.3 ;
      RECT 9.95 2.777 9.955 3.313 ;
      RECT 9.94 2.805 9.95 3.326 ;
      RECT 9.935 2.835 9.94 3.335 ;
      RECT 9.93 2.85 9.935 3.342 ;
      RECT 9.915 2.875 9.93 3.349 ;
      RECT 9.91 2.897 9.915 3.355 ;
      RECT 9.905 2.922 9.91 3.358 ;
      RECT 9.896 2.95 9.905 3.362 ;
      RECT 9.89 2.967 9.896 3.367 ;
      RECT 9.885 2.985 9.89 3.371 ;
      RECT 9.88 2.997 9.885 3.374 ;
      RECT 9.875 3.018 9.88 3.378 ;
      RECT 9.87 3.036 9.875 3.381 ;
      RECT 9.865 3.05 9.87 3.384 ;
      RECT 9.86 3.067 9.865 3.387 ;
      RECT 9.855 3.08 9.86 3.39 ;
      RECT 9.83 3.117 9.855 3.398 ;
      RECT 9.825 3.162 9.83 3.407 ;
      RECT 9.82 3.19 9.825 3.41 ;
      RECT 9.81 3.21 9.82 3.414 ;
      RECT 9.805 3.23 9.81 3.419 ;
      RECT 9.8 3.245 9.805 3.422 ;
      RECT 9.78 3.255 9.8 3.429 ;
      RECT 9.715 3.262 9.78 3.455 ;
      RECT 9.68 3.265 9.715 3.483 ;
      RECT 9.665 3.268 9.68 3.498 ;
      RECT 9.655 3.269 9.665 3.513 ;
      RECT 9.645 3.27 9.655 3.53 ;
      RECT 9.64 3.27 9.645 3.545 ;
      RECT 9.635 3.27 9.64 3.553 ;
      RECT 9.62 3.271 9.635 3.568 ;
      RECT 9.59 3.273 9.62 3.575 ;
      RECT 9.48 3.28 9.56 3.575 ;
      RECT 9.435 3.285 9.48 3.575 ;
      RECT 9.425 3.286 9.435 3.565 ;
      RECT 9.415 3.287 9.425 3.558 ;
      RECT 9.395 3.289 9.415 3.553 ;
      RECT 9.385 3.26 9.395 3.548 ;
      RECT 9.34 3.26 9.385 3.54 ;
      RECT 9.31 3.26 9.335 3.53 ;
      RECT 9.29 3.26 9.31 3.523 ;
      RECT 9.57 2.06 9.83 2.32 ;
      RECT 9.45 2.075 9.46 2.24 ;
      RECT 9.435 2.075 9.44 2.235 ;
      RECT 6.8 1.915 6.985 2.205 ;
      RECT 8.615 2.04 8.63 2.195 ;
      RECT 6.765 1.915 6.79 2.175 ;
      RECT 9.18 1.965 9.185 2.107 ;
      RECT 9.095 1.96 9.12 2.1 ;
      RECT 9.495 2.077 9.57 2.27 ;
      RECT 9.48 2.075 9.495 2.253 ;
      RECT 9.46 2.075 9.48 2.245 ;
      RECT 9.44 2.075 9.45 2.238 ;
      RECT 9.395 2.07 9.435 2.228 ;
      RECT 9.355 2.045 9.395 2.213 ;
      RECT 9.34 2.02 9.355 2.203 ;
      RECT 9.335 2.014 9.34 2.201 ;
      RECT 9.3 2.006 9.335 2.184 ;
      RECT 9.295 1.999 9.3 2.172 ;
      RECT 9.275 1.994 9.295 2.16 ;
      RECT 9.265 1.988 9.275 2.145 ;
      RECT 9.245 1.983 9.265 2.13 ;
      RECT 9.235 1.978 9.245 2.123 ;
      RECT 9.23 1.976 9.235 2.118 ;
      RECT 9.225 1.975 9.23 2.115 ;
      RECT 9.185 1.97 9.225 2.111 ;
      RECT 9.165 1.964 9.18 2.106 ;
      RECT 9.13 1.961 9.165 2.103 ;
      RECT 9.12 1.96 9.13 2.101 ;
      RECT 9.06 1.96 9.095 2.098 ;
      RECT 9.015 1.96 9.06 2.098 ;
      RECT 8.965 1.96 9.015 2.101 ;
      RECT 8.95 1.962 8.965 2.103 ;
      RECT 8.935 1.965 8.95 2.104 ;
      RECT 8.925 1.97 8.935 2.105 ;
      RECT 8.895 1.975 8.925 2.11 ;
      RECT 8.885 1.981 8.895 2.118 ;
      RECT 8.875 1.983 8.885 2.122 ;
      RECT 8.865 1.987 8.875 2.126 ;
      RECT 8.84 1.993 8.865 2.134 ;
      RECT 8.83 1.998 8.84 2.142 ;
      RECT 8.815 2.002 8.83 2.146 ;
      RECT 8.78 2.008 8.815 2.154 ;
      RECT 8.76 2.013 8.78 2.164 ;
      RECT 8.73 2.02 8.76 2.173 ;
      RECT 8.685 2.029 8.73 2.187 ;
      RECT 8.68 2.034 8.685 2.198 ;
      RECT 8.66 2.037 8.68 2.199 ;
      RECT 8.63 2.04 8.66 2.197 ;
      RECT 8.595 2.04 8.615 2.193 ;
      RECT 8.525 2.04 8.595 2.184 ;
      RECT 8.51 2.037 8.525 2.176 ;
      RECT 8.47 2.03 8.51 2.171 ;
      RECT 8.445 2.02 8.47 2.164 ;
      RECT 8.44 2.014 8.445 2.161 ;
      RECT 8.4 2.008 8.44 2.158 ;
      RECT 8.385 2.001 8.4 2.153 ;
      RECT 8.365 1.997 8.385 2.148 ;
      RECT 8.35 1.992 8.365 2.144 ;
      RECT 8.335 1.987 8.35 2.142 ;
      RECT 8.32 1.983 8.335 2.141 ;
      RECT 8.305 1.981 8.32 2.137 ;
      RECT 8.295 1.979 8.305 2.132 ;
      RECT 8.28 1.976 8.295 2.128 ;
      RECT 8.27 1.974 8.28 2.123 ;
      RECT 8.25 1.971 8.27 2.119 ;
      RECT 8.205 1.97 8.25 2.117 ;
      RECT 8.145 1.972 8.205 2.118 ;
      RECT 8.125 1.974 8.145 2.12 ;
      RECT 8.095 1.977 8.125 2.121 ;
      RECT 8.045 1.982 8.095 2.123 ;
      RECT 8.04 1.985 8.045 2.125 ;
      RECT 8.03 1.987 8.04 2.128 ;
      RECT 8.025 1.989 8.03 2.131 ;
      RECT 7.975 1.992 8.025 2.138 ;
      RECT 7.955 1.996 7.975 2.15 ;
      RECT 7.945 1.999 7.955 2.156 ;
      RECT 7.935 2 7.945 2.159 ;
      RECT 7.896 2.003 7.935 2.161 ;
      RECT 7.81 2.01 7.896 2.164 ;
      RECT 7.736 2.02 7.81 2.168 ;
      RECT 7.65 2.031 7.736 2.173 ;
      RECT 7.635 2.038 7.65 2.175 ;
      RECT 7.58 2.042 7.635 2.176 ;
      RECT 7.566 2.045 7.58 2.178 ;
      RECT 7.48 2.045 7.566 2.18 ;
      RECT 7.44 2.042 7.48 2.183 ;
      RECT 7.416 2.038 7.44 2.185 ;
      RECT 7.33 2.028 7.416 2.188 ;
      RECT 7.3 2.017 7.33 2.189 ;
      RECT 7.281 2.013 7.3 2.188 ;
      RECT 7.195 2.006 7.281 2.185 ;
      RECT 7.135 1.995 7.195 2.182 ;
      RECT 7.115 1.987 7.135 2.18 ;
      RECT 7.08 1.982 7.115 2.179 ;
      RECT 7.055 1.977 7.08 2.178 ;
      RECT 7.025 1.972 7.055 2.177 ;
      RECT 7 1.915 7.025 2.176 ;
      RECT 6.985 1.915 7 2.2 ;
      RECT 6.79 1.915 6.8 2.2 ;
      RECT 8.565 2.935 8.57 3.075 ;
      RECT 8.225 2.935 8.26 3.073 ;
      RECT 7.8 2.92 7.815 3.065 ;
      RECT 9.63 2.7 9.72 2.96 ;
      RECT 9.46 2.565 9.56 2.96 ;
      RECT 6.495 2.54 6.575 2.75 ;
      RECT 9.585 2.677 9.63 2.96 ;
      RECT 9.575 2.647 9.585 2.96 ;
      RECT 9.56 2.57 9.575 2.96 ;
      RECT 9.375 2.565 9.46 2.925 ;
      RECT 9.37 2.567 9.375 2.92 ;
      RECT 9.365 2.572 9.37 2.92 ;
      RECT 9.33 2.672 9.365 2.92 ;
      RECT 9.32 2.7 9.33 2.92 ;
      RECT 9.31 2.715 9.32 2.92 ;
      RECT 9.3 2.727 9.31 2.92 ;
      RECT 9.295 2.737 9.3 2.92 ;
      RECT 9.28 2.747 9.295 2.922 ;
      RECT 9.275 2.762 9.28 2.924 ;
      RECT 9.26 2.775 9.275 2.926 ;
      RECT 9.255 2.79 9.26 2.929 ;
      RECT 9.235 2.8 9.255 2.933 ;
      RECT 9.22 2.81 9.235 2.936 ;
      RECT 9.185 2.817 9.22 2.941 ;
      RECT 9.141 2.824 9.185 2.949 ;
      RECT 9.055 2.836 9.141 2.962 ;
      RECT 9.03 2.847 9.055 2.973 ;
      RECT 9 2.852 9.03 2.978 ;
      RECT 8.965 2.857 9 2.986 ;
      RECT 8.935 2.862 8.965 2.993 ;
      RECT 8.91 2.867 8.935 2.998 ;
      RECT 8.845 2.874 8.91 3.007 ;
      RECT 8.775 2.887 8.845 3.023 ;
      RECT 8.745 2.897 8.775 3.035 ;
      RECT 8.72 2.902 8.745 3.042 ;
      RECT 8.665 2.909 8.72 3.05 ;
      RECT 8.66 2.916 8.665 3.055 ;
      RECT 8.655 2.918 8.66 3.056 ;
      RECT 8.64 2.92 8.655 3.058 ;
      RECT 8.635 2.92 8.64 3.061 ;
      RECT 8.57 2.927 8.635 3.068 ;
      RECT 8.535 2.937 8.565 3.078 ;
      RECT 8.518 2.94 8.535 3.08 ;
      RECT 8.432 2.939 8.518 3.079 ;
      RECT 8.346 2.937 8.432 3.076 ;
      RECT 8.26 2.936 8.346 3.074 ;
      RECT 8.159 2.934 8.225 3.073 ;
      RECT 8.073 2.931 8.159 3.071 ;
      RECT 7.987 2.927 8.073 3.069 ;
      RECT 7.901 2.924 7.987 3.068 ;
      RECT 7.815 2.921 7.901 3.066 ;
      RECT 7.715 2.92 7.8 3.063 ;
      RECT 7.665 2.918 7.715 3.061 ;
      RECT 7.645 2.915 7.665 3.059 ;
      RECT 7.625 2.913 7.645 3.056 ;
      RECT 7.6 2.909 7.625 3.053 ;
      RECT 7.555 2.903 7.6 3.048 ;
      RECT 7.515 2.897 7.555 3.04 ;
      RECT 7.49 2.892 7.515 3.033 ;
      RECT 7.435 2.885 7.49 3.025 ;
      RECT 7.411 2.878 7.435 3.018 ;
      RECT 7.325 2.869 7.411 3.008 ;
      RECT 7.295 2.861 7.325 2.998 ;
      RECT 7.265 2.857 7.295 2.993 ;
      RECT 7.26 2.854 7.265 2.99 ;
      RECT 7.255 2.853 7.26 2.99 ;
      RECT 7.18 2.846 7.255 2.983 ;
      RECT 7.141 2.837 7.18 2.972 ;
      RECT 7.055 2.827 7.141 2.96 ;
      RECT 7.015 2.817 7.055 2.948 ;
      RECT 6.976 2.812 7.015 2.941 ;
      RECT 6.89 2.802 6.976 2.93 ;
      RECT 6.85 2.79 6.89 2.919 ;
      RECT 6.815 2.775 6.85 2.912 ;
      RECT 6.805 2.765 6.815 2.909 ;
      RECT 6.785 2.75 6.805 2.907 ;
      RECT 6.755 2.72 6.785 2.903 ;
      RECT 6.745 2.7 6.755 2.898 ;
      RECT 6.74 2.692 6.745 2.895 ;
      RECT 6.735 2.685 6.74 2.893 ;
      RECT 6.72 2.672 6.735 2.886 ;
      RECT 6.715 2.662 6.72 2.878 ;
      RECT 6.71 2.655 6.715 2.873 ;
      RECT 6.705 2.65 6.71 2.869 ;
      RECT 6.69 2.637 6.705 2.861 ;
      RECT 6.685 2.547 6.69 2.85 ;
      RECT 6.68 2.542 6.685 2.843 ;
      RECT 6.605 2.54 6.68 2.803 ;
      RECT 6.575 2.54 6.605 2.758 ;
      RECT 6.48 2.545 6.495 2.745 ;
      RECT 8.965 2.25 9.225 2.51 ;
      RECT 8.95 2.238 9.13 2.475 ;
      RECT 8.945 2.239 9.13 2.473 ;
      RECT 8.93 2.243 9.14 2.463 ;
      RECT 8.925 2.248 9.145 2.433 ;
      RECT 8.93 2.245 9.145 2.463 ;
      RECT 8.945 2.24 9.14 2.473 ;
      RECT 8.965 2.237 9.13 2.51 ;
      RECT 8.965 2.236 9.12 2.51 ;
      RECT 8.99 2.235 9.12 2.51 ;
      RECT 8.55 2.48 8.81 2.74 ;
      RECT 8.425 2.525 8.81 2.735 ;
      RECT 8.415 2.53 8.81 2.73 ;
      RECT 8.43 3.47 8.445 3.78 ;
      RECT 7.025 3.24 7.035 3.37 ;
      RECT 6.805 3.235 6.91 3.37 ;
      RECT 6.72 3.24 6.77 3.37 ;
      RECT 5.27 1.975 5.275 3.08 ;
      RECT 8.525 3.562 8.53 3.698 ;
      RECT 8.52 3.557 8.525 3.758 ;
      RECT 8.515 3.555 8.52 3.771 ;
      RECT 8.5 3.552 8.515 3.773 ;
      RECT 8.495 3.547 8.5 3.775 ;
      RECT 8.49 3.543 8.495 3.778 ;
      RECT 8.475 3.538 8.49 3.78 ;
      RECT 8.445 3.53 8.475 3.78 ;
      RECT 8.406 3.47 8.43 3.78 ;
      RECT 8.32 3.47 8.406 3.777 ;
      RECT 8.29 3.47 8.32 3.77 ;
      RECT 8.265 3.47 8.29 3.763 ;
      RECT 8.24 3.47 8.265 3.755 ;
      RECT 8.225 3.47 8.24 3.748 ;
      RECT 8.2 3.47 8.225 3.74 ;
      RECT 8.185 3.47 8.2 3.733 ;
      RECT 8.145 3.48 8.185 3.722 ;
      RECT 8.135 3.475 8.145 3.712 ;
      RECT 8.131 3.474 8.135 3.709 ;
      RECT 8.045 3.466 8.131 3.692 ;
      RECT 8.012 3.455 8.045 3.669 ;
      RECT 7.926 3.444 8.012 3.647 ;
      RECT 7.84 3.428 7.926 3.616 ;
      RECT 7.77 3.413 7.84 3.588 ;
      RECT 7.76 3.406 7.77 3.575 ;
      RECT 7.73 3.403 7.76 3.565 ;
      RECT 7.705 3.399 7.73 3.558 ;
      RECT 7.69 3.396 7.705 3.553 ;
      RECT 7.685 3.395 7.69 3.548 ;
      RECT 7.655 3.39 7.685 3.541 ;
      RECT 7.65 3.385 7.655 3.536 ;
      RECT 7.635 3.382 7.65 3.531 ;
      RECT 7.63 3.377 7.635 3.526 ;
      RECT 7.61 3.372 7.63 3.523 ;
      RECT 7.595 3.367 7.61 3.515 ;
      RECT 7.58 3.361 7.595 3.51 ;
      RECT 7.55 3.352 7.58 3.503 ;
      RECT 7.545 3.345 7.55 3.495 ;
      RECT 7.54 3.343 7.545 3.493 ;
      RECT 7.535 3.342 7.54 3.49 ;
      RECT 7.495 3.335 7.535 3.483 ;
      RECT 7.481 3.325 7.495 3.473 ;
      RECT 7.43 3.314 7.481 3.461 ;
      RECT 7.405 3.3 7.43 3.447 ;
      RECT 7.38 3.289 7.405 3.439 ;
      RECT 7.36 3.278 7.38 3.433 ;
      RECT 7.35 3.272 7.36 3.428 ;
      RECT 7.345 3.27 7.35 3.424 ;
      RECT 7.325 3.265 7.345 3.419 ;
      RECT 7.295 3.255 7.325 3.409 ;
      RECT 7.29 3.247 7.295 3.402 ;
      RECT 7.275 3.245 7.29 3.398 ;
      RECT 7.255 3.245 7.275 3.393 ;
      RECT 7.25 3.244 7.255 3.391 ;
      RECT 7.245 3.244 7.25 3.388 ;
      RECT 7.205 3.243 7.245 3.383 ;
      RECT 7.18 3.242 7.205 3.378 ;
      RECT 7.12 3.241 7.18 3.375 ;
      RECT 7.035 3.24 7.12 3.373 ;
      RECT 6.996 3.239 7.025 3.37 ;
      RECT 6.91 3.237 6.996 3.37 ;
      RECT 6.77 3.237 6.805 3.37 ;
      RECT 6.68 3.241 6.72 3.373 ;
      RECT 6.665 3.244 6.68 3.38 ;
      RECT 6.655 3.245 6.665 3.387 ;
      RECT 6.63 3.248 6.655 3.392 ;
      RECT 6.625 3.25 6.63 3.395 ;
      RECT 6.575 3.252 6.625 3.396 ;
      RECT 6.536 3.256 6.575 3.398 ;
      RECT 6.45 3.258 6.536 3.401 ;
      RECT 6.432 3.26 6.45 3.403 ;
      RECT 6.346 3.263 6.432 3.405 ;
      RECT 6.26 3.267 6.346 3.408 ;
      RECT 6.223 3.271 6.26 3.411 ;
      RECT 6.137 3.274 6.223 3.414 ;
      RECT 6.051 3.278 6.137 3.417 ;
      RECT 5.965 3.283 6.051 3.421 ;
      RECT 5.945 3.285 5.965 3.424 ;
      RECT 5.925 3.284 5.945 3.425 ;
      RECT 5.876 3.281 5.925 3.426 ;
      RECT 5.79 3.276 5.876 3.429 ;
      RECT 5.74 3.271 5.79 3.431 ;
      RECT 5.716 3.269 5.74 3.432 ;
      RECT 5.63 3.264 5.716 3.434 ;
      RECT 5.605 3.26 5.63 3.433 ;
      RECT 5.595 3.257 5.605 3.431 ;
      RECT 5.585 3.25 5.595 3.428 ;
      RECT 5.58 3.23 5.585 3.423 ;
      RECT 5.57 3.2 5.58 3.418 ;
      RECT 5.555 3.07 5.57 3.409 ;
      RECT 5.55 3.062 5.555 3.402 ;
      RECT 5.53 3.055 5.55 3.394 ;
      RECT 5.525 3.037 5.53 3.386 ;
      RECT 5.515 3.017 5.525 3.381 ;
      RECT 5.51 2.99 5.515 3.377 ;
      RECT 5.505 2.967 5.51 3.374 ;
      RECT 5.485 2.925 5.505 3.366 ;
      RECT 5.45 2.84 5.485 3.35 ;
      RECT 5.445 2.772 5.45 3.338 ;
      RECT 5.43 2.742 5.445 3.332 ;
      RECT 5.425 1.987 5.43 2.233 ;
      RECT 5.415 2.712 5.43 3.323 ;
      RECT 5.42 1.982 5.425 2.265 ;
      RECT 5.415 1.977 5.42 2.308 ;
      RECT 5.41 1.975 5.415 2.343 ;
      RECT 5.395 2.675 5.415 3.313 ;
      RECT 5.405 1.975 5.41 2.38 ;
      RECT 5.39 1.975 5.405 2.478 ;
      RECT 5.39 2.648 5.395 3.306 ;
      RECT 5.385 1.975 5.39 2.553 ;
      RECT 5.385 2.636 5.39 3.303 ;
      RECT 5.38 1.975 5.385 2.585 ;
      RECT 5.38 2.615 5.385 3.3 ;
      RECT 5.375 1.975 5.38 3.297 ;
      RECT 5.34 1.975 5.375 3.283 ;
      RECT 5.325 1.975 5.34 3.265 ;
      RECT 5.305 1.975 5.325 3.255 ;
      RECT 5.28 1.975 5.305 3.238 ;
      RECT 5.275 1.975 5.28 3.188 ;
      RECT 5.265 1.975 5.27 3.018 ;
      RECT 5.26 1.975 5.265 2.925 ;
      RECT 5.255 1.975 5.26 2.838 ;
      RECT 5.25 1.975 5.255 2.77 ;
      RECT 5.245 1.975 5.25 2.713 ;
      RECT 5.235 1.975 5.245 2.608 ;
      RECT 5.23 1.975 5.235 2.48 ;
      RECT 5.225 1.975 5.23 2.398 ;
      RECT 5.22 1.977 5.225 2.315 ;
      RECT 5.215 1.982 5.22 2.248 ;
      RECT 5.21 1.987 5.215 2.175 ;
      RECT 8.025 2.305 8.285 2.565 ;
      RECT 8.045 2.272 8.255 2.565 ;
      RECT 8.045 2.27 8.245 2.565 ;
      RECT 8.055 2.257 8.245 2.565 ;
      RECT 8.055 2.255 8.17 2.565 ;
      RECT 7.53 2.38 7.705 2.66 ;
      RECT 7.525 2.38 7.705 2.658 ;
      RECT 7.525 2.38 7.72 2.655 ;
      RECT 7.515 2.38 7.72 2.653 ;
      RECT 7.46 2.38 7.72 2.64 ;
      RECT 7.46 2.455 7.725 2.618 ;
      RECT 7.005 2.392 7.025 2.635 ;
      RECT 7.005 2.392 7.065 2.634 ;
      RECT 7 2.394 7.065 2.633 ;
      RECT 7 2.394 7.151 2.632 ;
      RECT 7 2.394 7.22 2.631 ;
      RECT 7 2.394 7.24 2.623 ;
      RECT 6.98 2.397 7.24 2.621 ;
      RECT 6.965 2.407 7.24 2.606 ;
      RECT 6.965 2.407 7.255 2.605 ;
      RECT 6.96 2.416 7.255 2.597 ;
      RECT 6.96 2.416 7.26 2.593 ;
      RECT 7.065 2.33 7.325 2.59 ;
      RECT 6.955 2.418 7.325 2.475 ;
      RECT 7.025 2.385 7.325 2.59 ;
      RECT 6.99 3.578 6.995 3.785 ;
      RECT 6.94 3.572 6.99 3.784 ;
      RECT 6.907 3.586 7 3.783 ;
      RECT 6.821 3.586 7 3.782 ;
      RECT 6.735 3.586 7 3.781 ;
      RECT 6.735 3.685 7.005 3.778 ;
      RECT 6.73 3.685 7.005 3.773 ;
      RECT 6.725 3.685 7.005 3.755 ;
      RECT 6.72 3.685 7.005 3.738 ;
      RECT 6.68 3.47 6.94 3.73 ;
      RECT 6.14 2.62 6.226 3.034 ;
      RECT 6.14 2.62 6.265 3.031 ;
      RECT 6.14 2.62 6.285 3.021 ;
      RECT 6.095 2.62 6.285 3.018 ;
      RECT 6.095 2.772 6.295 3.008 ;
      RECT 6.095 2.793 6.3 3.002 ;
      RECT 6.095 2.811 6.305 2.998 ;
      RECT 6.095 2.831 6.315 2.993 ;
      RECT 6.07 2.831 6.315 2.99 ;
      RECT 6.06 2.831 6.315 2.968 ;
      RECT 6.06 2.847 6.32 2.938 ;
      RECT 6.025 2.62 6.285 2.925 ;
      RECT 6.025 2.859 6.325 2.88 ;
      RECT 3.035 7.765 3.325 7.995 ;
      RECT 3.095 7.025 3.265 7.995 ;
      RECT 3.005 7.025 3.355 7.315 ;
      RECT 2.63 6.285 2.98 6.575 ;
      RECT 2.49 6.315 2.98 6.485 ;
      RECT 69.65 3.265 69.91 3.525 ;
      RECT 54.39 3.265 54.65 3.525 ;
      RECT 39.13 3.265 39.39 3.525 ;
      RECT 23.87 3.265 24.13 3.525 ;
      RECT 8.61 3.265 8.87 3.525 ;
    LAYER mcon ;
      RECT 80.045 6.32 80.215 6.49 ;
      RECT 80.05 6.315 80.22 6.485 ;
      RECT 64.785 6.32 64.955 6.49 ;
      RECT 64.79 6.315 64.96 6.485 ;
      RECT 49.525 6.32 49.695 6.49 ;
      RECT 49.53 6.315 49.7 6.485 ;
      RECT 34.265 6.32 34.435 6.49 ;
      RECT 34.27 6.315 34.44 6.485 ;
      RECT 19.005 6.32 19.175 6.49 ;
      RECT 19.01 6.315 19.18 6.485 ;
      RECT 80.045 7.8 80.215 7.97 ;
      RECT 79.695 0.1 79.865 0.27 ;
      RECT 79.695 8.61 79.865 8.78 ;
      RECT 79.675 2.76 79.845 2.93 ;
      RECT 79.675 5.95 79.845 6.12 ;
      RECT 79.055 0.91 79.225 1.08 ;
      RECT 79.055 2.39 79.225 2.56 ;
      RECT 79.055 6.32 79.225 6.49 ;
      RECT 79.055 7.8 79.225 7.97 ;
      RECT 78.705 0.1 78.875 0.27 ;
      RECT 78.705 8.61 78.875 8.78 ;
      RECT 78.685 2.76 78.855 2.93 ;
      RECT 78.685 5.95 78.855 6.12 ;
      RECT 78.005 0.105 78.175 0.275 ;
      RECT 78.005 8.605 78.175 8.775 ;
      RECT 77.695 2.025 77.865 2.195 ;
      RECT 77.695 6.685 77.865 6.855 ;
      RECT 77.325 0.105 77.495 0.275 ;
      RECT 77.325 8.605 77.495 8.775 ;
      RECT 77.265 0.915 77.435 1.085 ;
      RECT 77.265 1.655 77.435 1.825 ;
      RECT 77.265 7.055 77.435 7.225 ;
      RECT 77.265 7.795 77.435 7.965 ;
      RECT 76.89 2.395 77.06 2.565 ;
      RECT 76.89 6.315 77.06 6.485 ;
      RECT 76.645 0.105 76.815 0.275 ;
      RECT 76.645 8.605 76.815 8.775 ;
      RECT 75.965 0.105 76.135 0.275 ;
      RECT 75.965 8.605 76.135 8.775 ;
      RECT 74.505 1.415 74.675 1.585 ;
      RECT 74.065 2.28 74.235 2.45 ;
      RECT 74.045 1.415 74.215 1.585 ;
      RECT 73.67 3.025 73.84 3.195 ;
      RECT 73.585 1.415 73.755 1.585 ;
      RECT 73.56 2.3 73.73 2.47 ;
      RECT 73.125 1.415 73.295 1.585 ;
      RECT 72.74 1.99 72.91 2.16 ;
      RECT 72.665 1.415 72.835 1.585 ;
      RECT 72.425 3.03 72.595 3.2 ;
      RECT 72.38 2.52 72.55 2.69 ;
      RECT 72.37 8.605 72.54 8.775 ;
      RECT 72.205 1.415 72.375 1.585 ;
      RECT 72.06 6.685 72.23 6.855 ;
      RECT 71.955 2.73 72.125 2.9 ;
      RECT 71.765 1.95 71.935 2.12 ;
      RECT 71.745 1.415 71.915 1.585 ;
      RECT 71.715 3.56 71.885 3.73 ;
      RECT 71.69 8.605 71.86 8.775 ;
      RECT 71.63 7.055 71.8 7.225 ;
      RECT 71.63 7.795 71.8 7.965 ;
      RECT 71.38 3 71.55 3.17 ;
      RECT 71.285 1.415 71.455 1.585 ;
      RECT 71.285 2.16 71.455 2.33 ;
      RECT 71.255 6.315 71.425 6.485 ;
      RECT 71.01 8.605 71.18 8.775 ;
      RECT 70.825 1.415 70.995 1.585 ;
      RECT 70.485 3.385 70.655 3.555 ;
      RECT 70.425 2.585 70.595 2.755 ;
      RECT 70.365 1.415 70.535 1.585 ;
      RECT 70.33 8.605 70.5 8.775 ;
      RECT 69.985 2.255 70.155 2.425 ;
      RECT 69.905 1.415 70.075 1.585 ;
      RECT 69.72 3.305 69.89 3.475 ;
      RECT 69.475 2.545 69.645 2.715 ;
      RECT 69.445 1.415 69.615 1.585 ;
      RECT 69.38 3.575 69.55 3.745 ;
      RECT 69.105 2.27 69.275 2.44 ;
      RECT 68.985 1.415 69.155 1.585 ;
      RECT 68.575 2.47 68.745 2.64 ;
      RECT 68.525 1.415 68.695 1.585 ;
      RECT 68.065 1.415 68.235 1.585 ;
      RECT 68.055 2.415 68.225 2.585 ;
      RECT 67.85 2.015 68.02 2.185 ;
      RECT 67.85 3.595 68.02 3.765 ;
      RECT 67.605 1.415 67.775 1.585 ;
      RECT 67.54 2.56 67.71 2.73 ;
      RECT 67.145 1.415 67.315 1.585 ;
      RECT 67.13 2.785 67.3 2.955 ;
      RECT 66.685 1.415 66.855 1.585 ;
      RECT 66.42 3.085 66.59 3.255 ;
      RECT 66.275 1.995 66.445 2.165 ;
      RECT 66.225 1.415 66.395 1.585 ;
      RECT 64.785 7.8 64.955 7.97 ;
      RECT 64.435 0.1 64.605 0.27 ;
      RECT 64.435 8.61 64.605 8.78 ;
      RECT 64.415 2.76 64.585 2.93 ;
      RECT 64.415 5.95 64.585 6.12 ;
      RECT 63.795 0.91 63.965 1.08 ;
      RECT 63.795 2.39 63.965 2.56 ;
      RECT 63.795 6.32 63.965 6.49 ;
      RECT 63.795 7.8 63.965 7.97 ;
      RECT 63.445 0.1 63.615 0.27 ;
      RECT 63.445 8.61 63.615 8.78 ;
      RECT 63.425 2.76 63.595 2.93 ;
      RECT 63.425 5.95 63.595 6.12 ;
      RECT 62.745 0.105 62.915 0.275 ;
      RECT 62.745 8.605 62.915 8.775 ;
      RECT 62.435 2.025 62.605 2.195 ;
      RECT 62.435 6.685 62.605 6.855 ;
      RECT 62.065 0.105 62.235 0.275 ;
      RECT 62.065 8.605 62.235 8.775 ;
      RECT 62.005 0.915 62.175 1.085 ;
      RECT 62.005 1.655 62.175 1.825 ;
      RECT 62.005 7.055 62.175 7.225 ;
      RECT 62.005 7.795 62.175 7.965 ;
      RECT 61.63 2.395 61.8 2.565 ;
      RECT 61.63 6.315 61.8 6.485 ;
      RECT 61.385 0.105 61.555 0.275 ;
      RECT 61.385 8.605 61.555 8.775 ;
      RECT 60.705 0.105 60.875 0.275 ;
      RECT 60.705 8.605 60.875 8.775 ;
      RECT 59.245 1.415 59.415 1.585 ;
      RECT 58.805 2.28 58.975 2.45 ;
      RECT 58.785 1.415 58.955 1.585 ;
      RECT 58.41 3.025 58.58 3.195 ;
      RECT 58.325 1.415 58.495 1.585 ;
      RECT 58.3 2.3 58.47 2.47 ;
      RECT 57.865 1.415 58.035 1.585 ;
      RECT 57.48 1.99 57.65 2.16 ;
      RECT 57.405 1.415 57.575 1.585 ;
      RECT 57.165 3.03 57.335 3.2 ;
      RECT 57.12 2.52 57.29 2.69 ;
      RECT 57.11 8.605 57.28 8.775 ;
      RECT 56.945 1.415 57.115 1.585 ;
      RECT 56.8 6.685 56.97 6.855 ;
      RECT 56.695 2.73 56.865 2.9 ;
      RECT 56.505 1.95 56.675 2.12 ;
      RECT 56.485 1.415 56.655 1.585 ;
      RECT 56.455 3.56 56.625 3.73 ;
      RECT 56.43 8.605 56.6 8.775 ;
      RECT 56.37 7.055 56.54 7.225 ;
      RECT 56.37 7.795 56.54 7.965 ;
      RECT 56.12 3 56.29 3.17 ;
      RECT 56.025 1.415 56.195 1.585 ;
      RECT 56.025 2.16 56.195 2.33 ;
      RECT 55.995 6.315 56.165 6.485 ;
      RECT 55.75 8.605 55.92 8.775 ;
      RECT 55.565 1.415 55.735 1.585 ;
      RECT 55.225 3.385 55.395 3.555 ;
      RECT 55.165 2.585 55.335 2.755 ;
      RECT 55.105 1.415 55.275 1.585 ;
      RECT 55.07 8.605 55.24 8.775 ;
      RECT 54.725 2.255 54.895 2.425 ;
      RECT 54.645 1.415 54.815 1.585 ;
      RECT 54.46 3.305 54.63 3.475 ;
      RECT 54.215 2.545 54.385 2.715 ;
      RECT 54.185 1.415 54.355 1.585 ;
      RECT 54.12 3.575 54.29 3.745 ;
      RECT 53.845 2.27 54.015 2.44 ;
      RECT 53.725 1.415 53.895 1.585 ;
      RECT 53.315 2.47 53.485 2.64 ;
      RECT 53.265 1.415 53.435 1.585 ;
      RECT 52.805 1.415 52.975 1.585 ;
      RECT 52.795 2.415 52.965 2.585 ;
      RECT 52.59 2.015 52.76 2.185 ;
      RECT 52.59 3.595 52.76 3.765 ;
      RECT 52.345 1.415 52.515 1.585 ;
      RECT 52.28 2.56 52.45 2.73 ;
      RECT 51.885 1.415 52.055 1.585 ;
      RECT 51.87 2.785 52.04 2.955 ;
      RECT 51.425 1.415 51.595 1.585 ;
      RECT 51.16 3.085 51.33 3.255 ;
      RECT 51.015 1.995 51.185 2.165 ;
      RECT 50.965 1.415 51.135 1.585 ;
      RECT 49.525 7.8 49.695 7.97 ;
      RECT 49.175 0.1 49.345 0.27 ;
      RECT 49.175 8.61 49.345 8.78 ;
      RECT 49.155 2.76 49.325 2.93 ;
      RECT 49.155 5.95 49.325 6.12 ;
      RECT 48.535 0.91 48.705 1.08 ;
      RECT 48.535 2.39 48.705 2.56 ;
      RECT 48.535 6.32 48.705 6.49 ;
      RECT 48.535 7.8 48.705 7.97 ;
      RECT 48.185 0.1 48.355 0.27 ;
      RECT 48.185 8.61 48.355 8.78 ;
      RECT 48.165 2.76 48.335 2.93 ;
      RECT 48.165 5.95 48.335 6.12 ;
      RECT 47.485 0.105 47.655 0.275 ;
      RECT 47.485 8.605 47.655 8.775 ;
      RECT 47.175 2.025 47.345 2.195 ;
      RECT 47.175 6.685 47.345 6.855 ;
      RECT 46.805 0.105 46.975 0.275 ;
      RECT 46.805 8.605 46.975 8.775 ;
      RECT 46.745 0.915 46.915 1.085 ;
      RECT 46.745 1.655 46.915 1.825 ;
      RECT 46.745 7.055 46.915 7.225 ;
      RECT 46.745 7.795 46.915 7.965 ;
      RECT 46.37 2.395 46.54 2.565 ;
      RECT 46.37 6.315 46.54 6.485 ;
      RECT 46.125 0.105 46.295 0.275 ;
      RECT 46.125 8.605 46.295 8.775 ;
      RECT 45.445 0.105 45.615 0.275 ;
      RECT 45.445 8.605 45.615 8.775 ;
      RECT 43.985 1.415 44.155 1.585 ;
      RECT 43.545 2.28 43.715 2.45 ;
      RECT 43.525 1.415 43.695 1.585 ;
      RECT 43.15 3.025 43.32 3.195 ;
      RECT 43.065 1.415 43.235 1.585 ;
      RECT 43.04 2.3 43.21 2.47 ;
      RECT 42.605 1.415 42.775 1.585 ;
      RECT 42.22 1.99 42.39 2.16 ;
      RECT 42.145 1.415 42.315 1.585 ;
      RECT 41.905 3.03 42.075 3.2 ;
      RECT 41.86 2.52 42.03 2.69 ;
      RECT 41.85 8.605 42.02 8.775 ;
      RECT 41.685 1.415 41.855 1.585 ;
      RECT 41.54 6.685 41.71 6.855 ;
      RECT 41.435 2.73 41.605 2.9 ;
      RECT 41.245 1.95 41.415 2.12 ;
      RECT 41.225 1.415 41.395 1.585 ;
      RECT 41.195 3.56 41.365 3.73 ;
      RECT 41.17 8.605 41.34 8.775 ;
      RECT 41.11 7.055 41.28 7.225 ;
      RECT 41.11 7.795 41.28 7.965 ;
      RECT 40.86 3 41.03 3.17 ;
      RECT 40.765 1.415 40.935 1.585 ;
      RECT 40.765 2.16 40.935 2.33 ;
      RECT 40.735 6.315 40.905 6.485 ;
      RECT 40.49 8.605 40.66 8.775 ;
      RECT 40.305 1.415 40.475 1.585 ;
      RECT 39.965 3.385 40.135 3.555 ;
      RECT 39.905 2.585 40.075 2.755 ;
      RECT 39.845 1.415 40.015 1.585 ;
      RECT 39.81 8.605 39.98 8.775 ;
      RECT 39.465 2.255 39.635 2.425 ;
      RECT 39.385 1.415 39.555 1.585 ;
      RECT 39.2 3.305 39.37 3.475 ;
      RECT 38.955 2.545 39.125 2.715 ;
      RECT 38.925 1.415 39.095 1.585 ;
      RECT 38.86 3.575 39.03 3.745 ;
      RECT 38.585 2.27 38.755 2.44 ;
      RECT 38.465 1.415 38.635 1.585 ;
      RECT 38.055 2.47 38.225 2.64 ;
      RECT 38.005 1.415 38.175 1.585 ;
      RECT 37.545 1.415 37.715 1.585 ;
      RECT 37.535 2.415 37.705 2.585 ;
      RECT 37.33 2.015 37.5 2.185 ;
      RECT 37.33 3.595 37.5 3.765 ;
      RECT 37.085 1.415 37.255 1.585 ;
      RECT 37.02 2.56 37.19 2.73 ;
      RECT 36.625 1.415 36.795 1.585 ;
      RECT 36.61 2.785 36.78 2.955 ;
      RECT 36.165 1.415 36.335 1.585 ;
      RECT 35.9 3.085 36.07 3.255 ;
      RECT 35.755 1.995 35.925 2.165 ;
      RECT 35.705 1.415 35.875 1.585 ;
      RECT 34.265 7.8 34.435 7.97 ;
      RECT 33.915 0.1 34.085 0.27 ;
      RECT 33.915 8.61 34.085 8.78 ;
      RECT 33.895 2.76 34.065 2.93 ;
      RECT 33.895 5.95 34.065 6.12 ;
      RECT 33.275 0.91 33.445 1.08 ;
      RECT 33.275 2.39 33.445 2.56 ;
      RECT 33.275 6.32 33.445 6.49 ;
      RECT 33.275 7.8 33.445 7.97 ;
      RECT 32.925 0.1 33.095 0.27 ;
      RECT 32.925 8.61 33.095 8.78 ;
      RECT 32.905 2.76 33.075 2.93 ;
      RECT 32.905 5.95 33.075 6.12 ;
      RECT 32.225 0.105 32.395 0.275 ;
      RECT 32.225 8.605 32.395 8.775 ;
      RECT 31.915 2.025 32.085 2.195 ;
      RECT 31.915 6.685 32.085 6.855 ;
      RECT 31.545 0.105 31.715 0.275 ;
      RECT 31.545 8.605 31.715 8.775 ;
      RECT 31.485 0.915 31.655 1.085 ;
      RECT 31.485 1.655 31.655 1.825 ;
      RECT 31.485 7.055 31.655 7.225 ;
      RECT 31.485 7.795 31.655 7.965 ;
      RECT 31.11 2.395 31.28 2.565 ;
      RECT 31.11 6.315 31.28 6.485 ;
      RECT 30.865 0.105 31.035 0.275 ;
      RECT 30.865 8.605 31.035 8.775 ;
      RECT 30.185 0.105 30.355 0.275 ;
      RECT 30.185 8.605 30.355 8.775 ;
      RECT 28.725 1.415 28.895 1.585 ;
      RECT 28.285 2.28 28.455 2.45 ;
      RECT 28.265 1.415 28.435 1.585 ;
      RECT 27.89 3.025 28.06 3.195 ;
      RECT 27.805 1.415 27.975 1.585 ;
      RECT 27.78 2.3 27.95 2.47 ;
      RECT 27.345 1.415 27.515 1.585 ;
      RECT 26.96 1.99 27.13 2.16 ;
      RECT 26.885 1.415 27.055 1.585 ;
      RECT 26.645 3.03 26.815 3.2 ;
      RECT 26.6 2.52 26.77 2.69 ;
      RECT 26.59 8.605 26.76 8.775 ;
      RECT 26.425 1.415 26.595 1.585 ;
      RECT 26.28 6.685 26.45 6.855 ;
      RECT 26.175 2.73 26.345 2.9 ;
      RECT 25.985 1.95 26.155 2.12 ;
      RECT 25.965 1.415 26.135 1.585 ;
      RECT 25.935 3.56 26.105 3.73 ;
      RECT 25.91 8.605 26.08 8.775 ;
      RECT 25.85 7.055 26.02 7.225 ;
      RECT 25.85 7.795 26.02 7.965 ;
      RECT 25.6 3 25.77 3.17 ;
      RECT 25.505 1.415 25.675 1.585 ;
      RECT 25.505 2.16 25.675 2.33 ;
      RECT 25.475 6.315 25.645 6.485 ;
      RECT 25.23 8.605 25.4 8.775 ;
      RECT 25.045 1.415 25.215 1.585 ;
      RECT 24.705 3.385 24.875 3.555 ;
      RECT 24.645 2.585 24.815 2.755 ;
      RECT 24.585 1.415 24.755 1.585 ;
      RECT 24.55 8.605 24.72 8.775 ;
      RECT 24.205 2.255 24.375 2.425 ;
      RECT 24.125 1.415 24.295 1.585 ;
      RECT 23.94 3.305 24.11 3.475 ;
      RECT 23.695 2.545 23.865 2.715 ;
      RECT 23.665 1.415 23.835 1.585 ;
      RECT 23.6 3.575 23.77 3.745 ;
      RECT 23.325 2.27 23.495 2.44 ;
      RECT 23.205 1.415 23.375 1.585 ;
      RECT 22.795 2.47 22.965 2.64 ;
      RECT 22.745 1.415 22.915 1.585 ;
      RECT 22.285 1.415 22.455 1.585 ;
      RECT 22.275 2.415 22.445 2.585 ;
      RECT 22.07 2.015 22.24 2.185 ;
      RECT 22.07 3.595 22.24 3.765 ;
      RECT 21.825 1.415 21.995 1.585 ;
      RECT 21.76 2.56 21.93 2.73 ;
      RECT 21.365 1.415 21.535 1.585 ;
      RECT 21.35 2.785 21.52 2.955 ;
      RECT 20.905 1.415 21.075 1.585 ;
      RECT 20.64 3.085 20.81 3.255 ;
      RECT 20.495 1.995 20.665 2.165 ;
      RECT 20.445 1.415 20.615 1.585 ;
      RECT 19.005 7.8 19.175 7.97 ;
      RECT 18.655 0.1 18.825 0.27 ;
      RECT 18.655 8.61 18.825 8.78 ;
      RECT 18.635 2.76 18.805 2.93 ;
      RECT 18.635 5.95 18.805 6.12 ;
      RECT 18.015 0.91 18.185 1.08 ;
      RECT 18.015 2.39 18.185 2.56 ;
      RECT 18.015 6.32 18.185 6.49 ;
      RECT 18.015 7.8 18.185 7.97 ;
      RECT 17.665 0.1 17.835 0.27 ;
      RECT 17.665 8.61 17.835 8.78 ;
      RECT 17.645 2.76 17.815 2.93 ;
      RECT 17.645 5.95 17.815 6.12 ;
      RECT 16.965 0.105 17.135 0.275 ;
      RECT 16.965 8.605 17.135 8.775 ;
      RECT 16.655 2.025 16.825 2.195 ;
      RECT 16.655 6.685 16.825 6.855 ;
      RECT 16.285 0.105 16.455 0.275 ;
      RECT 16.285 8.605 16.455 8.775 ;
      RECT 16.225 0.915 16.395 1.085 ;
      RECT 16.225 1.655 16.395 1.825 ;
      RECT 16.225 7.055 16.395 7.225 ;
      RECT 16.225 7.795 16.395 7.965 ;
      RECT 15.85 2.395 16.02 2.565 ;
      RECT 15.85 6.315 16.02 6.485 ;
      RECT 15.605 0.105 15.775 0.275 ;
      RECT 15.605 8.605 15.775 8.775 ;
      RECT 14.925 0.105 15.095 0.275 ;
      RECT 14.925 8.605 15.095 8.775 ;
      RECT 13.465 1.415 13.635 1.585 ;
      RECT 13.025 2.28 13.195 2.45 ;
      RECT 13.005 1.415 13.175 1.585 ;
      RECT 12.63 3.025 12.8 3.195 ;
      RECT 12.545 1.415 12.715 1.585 ;
      RECT 12.52 2.3 12.69 2.47 ;
      RECT 12.085 1.415 12.255 1.585 ;
      RECT 11.7 1.99 11.87 2.16 ;
      RECT 11.625 1.415 11.795 1.585 ;
      RECT 11.385 3.03 11.555 3.2 ;
      RECT 11.34 2.52 11.51 2.69 ;
      RECT 11.33 8.605 11.5 8.775 ;
      RECT 11.165 1.415 11.335 1.585 ;
      RECT 11.02 6.685 11.19 6.855 ;
      RECT 10.915 2.73 11.085 2.9 ;
      RECT 10.725 1.95 10.895 2.12 ;
      RECT 10.705 1.415 10.875 1.585 ;
      RECT 10.675 3.56 10.845 3.73 ;
      RECT 10.65 8.605 10.82 8.775 ;
      RECT 10.59 7.055 10.76 7.225 ;
      RECT 10.59 7.795 10.76 7.965 ;
      RECT 10.34 3 10.51 3.17 ;
      RECT 10.245 1.415 10.415 1.585 ;
      RECT 10.245 2.16 10.415 2.33 ;
      RECT 10.215 6.315 10.385 6.485 ;
      RECT 9.97 8.605 10.14 8.775 ;
      RECT 9.785 1.415 9.955 1.585 ;
      RECT 9.445 3.385 9.615 3.555 ;
      RECT 9.385 2.585 9.555 2.755 ;
      RECT 9.325 1.415 9.495 1.585 ;
      RECT 9.29 8.605 9.46 8.775 ;
      RECT 8.945 2.255 9.115 2.425 ;
      RECT 8.865 1.415 9.035 1.585 ;
      RECT 8.68 3.305 8.85 3.475 ;
      RECT 8.435 2.545 8.605 2.715 ;
      RECT 8.405 1.415 8.575 1.585 ;
      RECT 8.34 3.575 8.51 3.745 ;
      RECT 8.065 2.27 8.235 2.44 ;
      RECT 7.945 1.415 8.115 1.585 ;
      RECT 7.535 2.47 7.705 2.64 ;
      RECT 7.485 1.415 7.655 1.585 ;
      RECT 7.025 1.415 7.195 1.585 ;
      RECT 7.015 2.415 7.185 2.585 ;
      RECT 6.81 2.015 6.98 2.185 ;
      RECT 6.81 3.595 6.98 3.765 ;
      RECT 6.565 1.415 6.735 1.585 ;
      RECT 6.5 2.56 6.67 2.73 ;
      RECT 6.105 1.415 6.275 1.585 ;
      RECT 6.09 2.785 6.26 2.955 ;
      RECT 5.645 1.415 5.815 1.585 ;
      RECT 5.38 3.085 5.55 3.255 ;
      RECT 5.235 1.995 5.405 2.165 ;
      RECT 5.185 1.415 5.355 1.585 ;
      RECT 3.835 8.605 4.005 8.775 ;
      RECT 3.155 8.605 3.325 8.775 ;
      RECT 3.095 7.055 3.265 7.225 ;
      RECT 3.095 7.795 3.265 7.965 ;
      RECT 2.72 6.315 2.89 6.485 ;
      RECT 2.475 8.605 2.645 8.775 ;
      RECT 1.795 8.605 1.965 8.775 ;
    LAYER li1 ;
      RECT 74.05 0 74.22 2.085 ;
      RECT 73.11 0 73.28 2.085 ;
      RECT 72.15 0 72.32 2.085 ;
      RECT 70.23 0 70.4 2.085 ;
      RECT 69.27 0 69.44 2.085 ;
      RECT 67.35 0 67.52 2.085 ;
      RECT 58.79 0 58.96 2.085 ;
      RECT 57.85 0 58.02 2.085 ;
      RECT 56.89 0 57.06 2.085 ;
      RECT 54.97 0 55.14 2.085 ;
      RECT 54.01 0 54.18 2.085 ;
      RECT 52.09 0 52.26 2.085 ;
      RECT 43.53 0 43.7 2.085 ;
      RECT 42.59 0 42.76 2.085 ;
      RECT 41.63 0 41.8 2.085 ;
      RECT 39.71 0 39.88 2.085 ;
      RECT 38.75 0 38.92 2.085 ;
      RECT 36.83 0 37 2.085 ;
      RECT 28.27 0 28.44 2.085 ;
      RECT 27.33 0 27.5 2.085 ;
      RECT 26.37 0 26.54 2.085 ;
      RECT 24.45 0 24.62 2.085 ;
      RECT 23.49 0 23.66 2.085 ;
      RECT 21.57 0 21.74 2.085 ;
      RECT 13.01 0 13.18 2.085 ;
      RECT 12.07 0 12.24 2.085 ;
      RECT 11.11 0 11.28 2.085 ;
      RECT 9.19 0 9.36 2.085 ;
      RECT 8.23 0 8.4 2.085 ;
      RECT 6.31 0 6.48 2.085 ;
      RECT 71.105 0 71.3 1.595 ;
      RECT 67.35 0 67.625 1.595 ;
      RECT 55.845 0 56.04 1.595 ;
      RECT 52.09 0 52.365 1.595 ;
      RECT 40.585 0 40.78 1.595 ;
      RECT 36.83 0 37.105 1.595 ;
      RECT 25.325 0 25.52 1.595 ;
      RECT 21.57 0 21.845 1.595 ;
      RECT 10.065 0 10.26 1.595 ;
      RECT 6.31 0 6.585 1.595 ;
      RECT 66.08 0 74.82 1.585 ;
      RECT 50.82 0 59.56 1.585 ;
      RECT 35.56 0 44.3 1.585 ;
      RECT 20.3 0 29.04 1.585 ;
      RECT 5.04 0 13.78 1.585 ;
      RECT 75.885 0 76.055 0.935 ;
      RECT 60.625 0 60.795 0.935 ;
      RECT 45.365 0 45.535 0.935 ;
      RECT 30.105 0 30.275 0.935 ;
      RECT 14.845 0 15.015 0.935 ;
      RECT 79.615 0 79.785 0.93 ;
      RECT 78.625 0 78.795 0.93 ;
      RECT 64.355 0 64.525 0.93 ;
      RECT 63.365 0 63.535 0.93 ;
      RECT 49.095 0 49.265 0.93 ;
      RECT 48.105 0 48.275 0.93 ;
      RECT 33.835 0 34.005 0.93 ;
      RECT 32.845 0 33.015 0.93 ;
      RECT 18.575 0 18.745 0.93 ;
      RECT 17.585 0 17.755 0.93 ;
      RECT 80.41 0 80.59 0.305 ;
      RECT 65.15 0 78.46 0.305 ;
      RECT 49.89 0 63.2 0.305 ;
      RECT 34.63 0 47.94 0.305 ;
      RECT 19.37 0 32.68 0.305 ;
      RECT 1.495 0 17.42 0.305 ;
      RECT 1.495 0 80.59 0.3 ;
      RECT 1.495 8.58 80.59 8.88 ;
      RECT 80.41 8.575 80.59 8.88 ;
      RECT 79.615 7.95 79.785 8.88 ;
      RECT 78.625 7.95 78.795 8.88 ;
      RECT 65.15 8.575 78.46 8.88 ;
      RECT 64.355 7.95 64.525 8.88 ;
      RECT 63.365 7.95 63.535 8.88 ;
      RECT 49.89 8.575 63.2 8.88 ;
      RECT 49.095 7.95 49.265 8.88 ;
      RECT 48.105 7.95 48.275 8.88 ;
      RECT 34.63 8.575 47.94 8.88 ;
      RECT 33.835 7.95 34.005 8.88 ;
      RECT 32.845 7.95 33.015 8.88 ;
      RECT 19.37 8.575 32.68 8.88 ;
      RECT 18.575 7.95 18.745 8.88 ;
      RECT 17.585 7.95 17.755 8.88 ;
      RECT 1.495 8.575 17.42 8.88 ;
      RECT 75.885 7.945 76.055 8.88 ;
      RECT 70.25 7.945 70.42 8.88 ;
      RECT 60.625 7.945 60.795 8.88 ;
      RECT 54.99 7.945 55.16 8.88 ;
      RECT 45.365 7.945 45.535 8.88 ;
      RECT 39.73 7.945 39.9 8.88 ;
      RECT 30.105 7.945 30.275 8.88 ;
      RECT 24.47 7.945 24.64 8.88 ;
      RECT 14.845 7.945 15.015 8.88 ;
      RECT 9.21 7.945 9.38 8.88 ;
      RECT 1.715 7.945 1.885 8.88 ;
      RECT 80.045 5.02 80.215 6.49 ;
      RECT 80.045 6.315 80.22 6.485 ;
      RECT 79.675 1.74 79.845 2.93 ;
      RECT 79.675 1.74 80.145 1.91 ;
      RECT 79.675 6.97 80.145 7.14 ;
      RECT 79.675 5.95 79.845 7.14 ;
      RECT 78.685 1.74 78.855 2.93 ;
      RECT 78.685 1.74 79.155 1.91 ;
      RECT 78.685 6.97 79.155 7.14 ;
      RECT 78.685 5.95 78.855 7.14 ;
      RECT 76.835 2.635 77.005 3.865 ;
      RECT 76.89 0.855 77.06 2.805 ;
      RECT 76.835 0.575 77.005 1.025 ;
      RECT 76.835 7.855 77.005 8.305 ;
      RECT 76.89 6.075 77.06 8.025 ;
      RECT 76.835 5.015 77.005 6.245 ;
      RECT 76.315 0.575 76.485 3.865 ;
      RECT 76.315 2.075 76.72 2.405 ;
      RECT 76.315 1.235 76.72 1.565 ;
      RECT 76.315 5.015 76.485 8.305 ;
      RECT 76.315 7.315 76.72 7.645 ;
      RECT 76.315 6.475 76.72 6.805 ;
      RECT 74.24 3.126 74.245 3.298 ;
      RECT 74.235 3.119 74.24 3.388 ;
      RECT 74.23 3.113 74.235 3.407 ;
      RECT 74.21 3.107 74.23 3.417 ;
      RECT 74.195 3.102 74.21 3.425 ;
      RECT 74.158 3.096 74.195 3.423 ;
      RECT 74.072 3.082 74.158 3.419 ;
      RECT 73.986 3.064 74.072 3.414 ;
      RECT 73.9 3.045 73.986 3.408 ;
      RECT 73.87 3.033 73.9 3.404 ;
      RECT 73.85 3.027 73.87 3.403 ;
      RECT 73.785 3.025 73.85 3.401 ;
      RECT 73.77 3.025 73.785 3.393 ;
      RECT 73.755 3.025 73.77 3.38 ;
      RECT 73.75 3.025 73.755 3.37 ;
      RECT 73.735 3.025 73.75 3.348 ;
      RECT 73.72 3.025 73.735 3.315 ;
      RECT 73.715 3.025 73.72 3.293 ;
      RECT 73.705 3.025 73.715 3.275 ;
      RECT 73.69 3.025 73.705 3.253 ;
      RECT 73.67 3.025 73.69 3.215 ;
      RECT 74.02 2.31 74.055 2.749 ;
      RECT 74.02 2.31 74.06 2.748 ;
      RECT 73.965 2.37 74.06 2.747 ;
      RECT 73.83 2.542 74.06 2.746 ;
      RECT 73.94 2.42 74.06 2.746 ;
      RECT 73.83 2.542 74.085 2.736 ;
      RECT 73.885 2.487 74.165 2.653 ;
      RECT 74.06 2.281 74.065 2.744 ;
      RECT 73.915 2.457 74.205 2.53 ;
      RECT 73.93 2.44 74.06 2.746 ;
      RECT 74.065 2.28 74.235 2.468 ;
      RECT 74.055 2.283 74.235 2.468 ;
      RECT 73.56 2.16 73.73 2.47 ;
      RECT 73.56 2.16 73.735 2.443 ;
      RECT 73.56 2.16 73.74 2.42 ;
      RECT 73.56 2.16 73.75 2.37 ;
      RECT 73.555 2.265 73.75 2.34 ;
      RECT 73.59 1.835 73.76 2.313 ;
      RECT 73.59 1.835 73.775 2.234 ;
      RECT 73.58 2.045 73.775 2.234 ;
      RECT 73.59 1.845 73.785 2.149 ;
      RECT 73.52 2.587 73.525 2.79 ;
      RECT 73.51 2.575 73.52 2.9 ;
      RECT 73.485 2.575 73.51 2.94 ;
      RECT 73.405 2.575 73.485 3.025 ;
      RECT 73.395 2.575 73.405 3.095 ;
      RECT 73.37 2.575 73.395 3.118 ;
      RECT 73.35 2.575 73.37 3.153 ;
      RECT 73.305 2.585 73.35 3.196 ;
      RECT 73.295 2.597 73.305 3.233 ;
      RECT 73.275 2.611 73.295 3.253 ;
      RECT 73.265 2.629 73.275 3.269 ;
      RECT 73.25 2.655 73.265 3.279 ;
      RECT 73.235 2.696 73.25 3.293 ;
      RECT 73.225 2.731 73.235 3.303 ;
      RECT 73.22 2.747 73.225 3.308 ;
      RECT 73.21 2.762 73.22 3.313 ;
      RECT 73.19 2.805 73.21 3.323 ;
      RECT 73.17 2.842 73.19 3.336 ;
      RECT 73.135 2.865 73.17 3.354 ;
      RECT 73.125 2.879 73.135 3.37 ;
      RECT 73.105 2.889 73.125 3.38 ;
      RECT 73.1 2.898 73.105 3.388 ;
      RECT 73.09 2.905 73.1 3.395 ;
      RECT 73.08 2.912 73.09 3.403 ;
      RECT 73.065 2.922 73.08 3.411 ;
      RECT 73.055 2.936 73.065 3.421 ;
      RECT 73.045 2.948 73.055 3.433 ;
      RECT 73.03 2.97 73.045 3.446 ;
      RECT 73.02 2.992 73.03 3.457 ;
      RECT 73.01 3.012 73.02 3.466 ;
      RECT 73.005 3.027 73.01 3.473 ;
      RECT 72.975 3.06 73.005 3.487 ;
      RECT 72.965 3.095 72.975 3.502 ;
      RECT 72.96 3.102 72.965 3.508 ;
      RECT 72.94 3.117 72.96 3.515 ;
      RECT 72.935 3.132 72.94 3.523 ;
      RECT 72.93 3.141 72.935 3.528 ;
      RECT 72.915 3.147 72.93 3.535 ;
      RECT 72.91 3.153 72.915 3.543 ;
      RECT 72.905 3.157 72.91 3.55 ;
      RECT 72.9 3.161 72.905 3.56 ;
      RECT 72.89 3.166 72.9 3.57 ;
      RECT 72.87 3.177 72.89 3.598 ;
      RECT 72.855 3.189 72.87 3.625 ;
      RECT 72.835 3.202 72.855 3.65 ;
      RECT 72.815 3.217 72.835 3.674 ;
      RECT 72.8 3.232 72.815 3.689 ;
      RECT 72.795 3.243 72.8 3.698 ;
      RECT 72.73 3.288 72.795 3.708 ;
      RECT 72.695 3.347 72.73 3.721 ;
      RECT 72.69 3.37 72.695 3.727 ;
      RECT 72.685 3.377 72.69 3.729 ;
      RECT 72.67 3.387 72.685 3.732 ;
      RECT 72.64 3.412 72.67 3.736 ;
      RECT 72.635 3.43 72.64 3.74 ;
      RECT 72.63 3.437 72.635 3.741 ;
      RECT 72.61 3.445 72.63 3.745 ;
      RECT 72.6 3.452 72.61 3.749 ;
      RECT 72.556 3.463 72.6 3.756 ;
      RECT 72.47 3.491 72.556 3.772 ;
      RECT 72.41 3.515 72.47 3.79 ;
      RECT 72.365 3.525 72.41 3.804 ;
      RECT 72.306 3.533 72.365 3.818 ;
      RECT 72.22 3.54 72.306 3.837 ;
      RECT 72.195 3.545 72.22 3.852 ;
      RECT 72.115 3.548 72.195 3.855 ;
      RECT 72.035 3.552 72.115 3.842 ;
      RECT 72.026 3.555 72.035 3.827 ;
      RECT 71.94 3.555 72.026 3.812 ;
      RECT 71.88 3.557 71.94 3.789 ;
      RECT 71.876 3.56 71.88 3.779 ;
      RECT 71.79 3.56 71.876 3.764 ;
      RECT 71.715 3.56 71.79 3.74 ;
      RECT 73.03 2.569 73.04 2.745 ;
      RECT 72.985 2.536 73.03 2.745 ;
      RECT 72.94 2.487 72.985 2.745 ;
      RECT 72.91 2.457 72.94 2.746 ;
      RECT 72.905 2.44 72.91 2.747 ;
      RECT 72.88 2.42 72.905 2.748 ;
      RECT 72.865 2.395 72.88 2.749 ;
      RECT 72.86 2.382 72.865 2.75 ;
      RECT 72.855 2.376 72.86 2.748 ;
      RECT 72.85 2.368 72.855 2.742 ;
      RECT 72.825 2.36 72.85 2.722 ;
      RECT 72.805 2.349 72.825 2.693 ;
      RECT 72.775 2.334 72.805 2.664 ;
      RECT 72.755 2.32 72.775 2.636 ;
      RECT 72.745 2.314 72.755 2.615 ;
      RECT 72.74 2.311 72.745 2.598 ;
      RECT 72.735 2.308 72.74 2.583 ;
      RECT 72.72 2.303 72.735 2.548 ;
      RECT 72.715 2.299 72.72 2.515 ;
      RECT 72.695 2.294 72.715 2.491 ;
      RECT 72.665 2.286 72.695 2.456 ;
      RECT 72.65 2.28 72.665 2.433 ;
      RECT 72.61 2.273 72.65 2.418 ;
      RECT 72.585 2.265 72.61 2.398 ;
      RECT 72.565 2.26 72.585 2.388 ;
      RECT 72.53 2.254 72.565 2.383 ;
      RECT 72.485 2.245 72.53 2.382 ;
      RECT 72.455 2.241 72.485 2.384 ;
      RECT 72.37 2.249 72.455 2.388 ;
      RECT 72.3 2.26 72.37 2.41 ;
      RECT 72.287 2.266 72.3 2.433 ;
      RECT 72.201 2.273 72.287 2.455 ;
      RECT 72.115 2.285 72.201 2.492 ;
      RECT 72.115 2.662 72.125 2.9 ;
      RECT 72.11 2.291 72.115 2.515 ;
      RECT 72.105 2.547 72.115 2.9 ;
      RECT 72.105 2.292 72.11 2.52 ;
      RECT 72.1 2.293 72.105 2.9 ;
      RECT 72.076 2.295 72.1 2.901 ;
      RECT 71.99 2.303 72.076 2.903 ;
      RECT 71.97 2.317 71.99 2.906 ;
      RECT 71.965 2.345 71.97 2.907 ;
      RECT 71.96 2.357 71.965 2.908 ;
      RECT 71.955 2.372 71.96 2.909 ;
      RECT 71.945 2.402 71.955 2.91 ;
      RECT 71.94 2.44 71.945 2.908 ;
      RECT 71.935 2.46 71.94 2.903 ;
      RECT 71.92 2.495 71.935 2.888 ;
      RECT 71.91 2.547 71.92 2.868 ;
      RECT 71.905 2.577 71.91 2.856 ;
      RECT 71.89 2.59 71.905 2.839 ;
      RECT 71.865 2.594 71.89 2.806 ;
      RECT 71.85 2.592 71.865 2.783 ;
      RECT 71.835 2.591 71.85 2.78 ;
      RECT 71.775 2.589 71.835 2.778 ;
      RECT 71.765 2.587 71.775 2.773 ;
      RECT 71.725 2.586 71.765 2.77 ;
      RECT 71.655 2.583 71.725 2.768 ;
      RECT 71.6 2.581 71.655 2.763 ;
      RECT 71.53 2.575 71.6 2.758 ;
      RECT 71.521 2.575 71.53 2.755 ;
      RECT 71.435 2.575 71.521 2.75 ;
      RECT 71.43 2.575 71.435 2.745 ;
      RECT 72.735 1.81 72.91 2.16 ;
      RECT 72.735 1.825 72.92 2.158 ;
      RECT 72.71 1.775 72.855 2.155 ;
      RECT 72.69 1.776 72.855 2.148 ;
      RECT 72.68 1.777 72.865 2.143 ;
      RECT 72.65 1.778 72.865 2.13 ;
      RECT 72.6 1.779 72.865 2.106 ;
      RECT 72.595 1.781 72.865 2.091 ;
      RECT 72.595 1.847 72.925 2.085 ;
      RECT 72.575 1.788 72.88 2.065 ;
      RECT 72.565 1.797 72.89 1.92 ;
      RECT 72.575 1.792 72.89 2.065 ;
      RECT 72.595 1.782 72.88 2.091 ;
      RECT 72.18 3.107 72.35 3.395 ;
      RECT 72.175 3.125 72.36 3.39 ;
      RECT 72.14 3.133 72.425 3.31 ;
      RECT 72.14 3.133 72.511 3.3 ;
      RECT 72.14 3.133 72.565 3.246 ;
      RECT 72.425 3.03 72.595 3.214 ;
      RECT 72.14 3.185 72.6 3.202 ;
      RECT 72.125 3.155 72.595 3.198 ;
      RECT 72.385 3.037 72.425 3.349 ;
      RECT 72.265 3.074 72.595 3.214 ;
      RECT 72.36 3.049 72.385 3.375 ;
      RECT 72.35 3.056 72.595 3.214 ;
      RECT 72.481 2.52 72.55 2.779 ;
      RECT 72.481 2.575 72.555 2.778 ;
      RECT 72.395 2.575 72.555 2.777 ;
      RECT 72.39 2.575 72.56 2.77 ;
      RECT 72.38 2.52 72.55 2.765 ;
      RECT 71.76 1.819 71.935 2.12 ;
      RECT 71.745 1.807 71.76 2.105 ;
      RECT 71.715 1.806 71.745 2.058 ;
      RECT 71.715 1.824 71.94 2.053 ;
      RECT 71.7 1.808 71.76 2.018 ;
      RECT 71.695 1.83 71.95 1.918 ;
      RECT 71.695 1.813 71.846 1.918 ;
      RECT 71.695 1.815 71.85 1.918 ;
      RECT 71.7 1.811 71.846 2.018 ;
      RECT 71.805 3.047 71.81 3.395 ;
      RECT 71.795 3.037 71.805 3.401 ;
      RECT 71.76 3.027 71.795 3.403 ;
      RECT 71.722 3.022 71.76 3.407 ;
      RECT 71.636 3.015 71.722 3.414 ;
      RECT 71.55 3.005 71.636 3.424 ;
      RECT 71.505 3 71.55 3.432 ;
      RECT 71.501 3 71.505 3.436 ;
      RECT 71.415 3 71.501 3.443 ;
      RECT 71.4 3 71.415 3.443 ;
      RECT 71.39 2.998 71.4 3.415 ;
      RECT 71.38 2.994 71.39 3.358 ;
      RECT 71.36 2.988 71.38 3.29 ;
      RECT 71.355 2.984 71.36 3.238 ;
      RECT 71.345 2.983 71.355 3.205 ;
      RECT 71.295 2.981 71.345 3.19 ;
      RECT 71.27 2.979 71.295 3.185 ;
      RECT 71.227 2.977 71.27 3.181 ;
      RECT 71.141 2.973 71.227 3.169 ;
      RECT 71.055 2.968 71.141 3.153 ;
      RECT 71.025 2.965 71.055 3.14 ;
      RECT 71 2.964 71.025 3.128 ;
      RECT 70.995 2.964 71 3.118 ;
      RECT 70.955 2.963 70.995 3.11 ;
      RECT 70.94 2.962 70.955 3.103 ;
      RECT 70.89 2.961 70.94 3.095 ;
      RECT 70.888 2.96 70.89 3.09 ;
      RECT 70.802 2.958 70.888 3.09 ;
      RECT 70.716 2.953 70.802 3.09 ;
      RECT 70.63 2.949 70.716 3.09 ;
      RECT 70.581 2.945 70.63 3.088 ;
      RECT 70.495 2.942 70.581 3.083 ;
      RECT 70.472 2.939 70.495 3.079 ;
      RECT 70.386 2.936 70.472 3.074 ;
      RECT 70.3 2.932 70.386 3.065 ;
      RECT 70.275 2.925 70.3 3.06 ;
      RECT 70.215 2.89 70.275 3.057 ;
      RECT 70.195 2.815 70.215 3.054 ;
      RECT 70.19 2.757 70.195 3.053 ;
      RECT 70.165 2.697 70.19 3.052 ;
      RECT 70.09 2.575 70.165 3.048 ;
      RECT 70.08 2.575 70.09 3.04 ;
      RECT 70.065 2.575 70.08 3.03 ;
      RECT 70.05 2.575 70.065 3 ;
      RECT 70.035 2.575 70.05 2.945 ;
      RECT 70.02 2.575 70.035 2.883 ;
      RECT 69.995 2.575 70.02 2.808 ;
      RECT 69.99 2.575 69.995 2.758 ;
      RECT 71.335 2.12 71.355 2.429 ;
      RECT 71.321 2.122 71.37 2.426 ;
      RECT 71.321 2.127 71.39 2.417 ;
      RECT 71.235 2.125 71.37 2.411 ;
      RECT 71.235 2.133 71.425 2.394 ;
      RECT 71.2 2.135 71.425 2.393 ;
      RECT 71.17 2.143 71.425 2.384 ;
      RECT 71.16 2.148 71.445 2.37 ;
      RECT 71.2 2.138 71.445 2.37 ;
      RECT 71.2 2.141 71.455 2.358 ;
      RECT 71.17 2.143 71.465 2.345 ;
      RECT 71.17 2.147 71.475 2.288 ;
      RECT 71.16 2.152 71.48 2.203 ;
      RECT 71.321 2.12 71.355 2.426 ;
      RECT 71.2 7.855 71.37 8.305 ;
      RECT 71.255 6.075 71.425 8.025 ;
      RECT 71.2 5.015 71.37 6.245 ;
      RECT 70.76 2.223 70.765 2.435 ;
      RECT 70.635 2.22 70.65 2.435 ;
      RECT 70.1 2.25 70.17 2.435 ;
      RECT 69.985 2.25 70.02 2.43 ;
      RECT 71.106 2.552 71.125 2.746 ;
      RECT 71.02 2.507 71.106 2.747 ;
      RECT 71.01 2.46 71.02 2.749 ;
      RECT 71.005 2.44 71.01 2.75 ;
      RECT 70.985 2.405 71.005 2.751 ;
      RECT 70.97 2.355 70.985 2.752 ;
      RECT 70.95 2.292 70.97 2.753 ;
      RECT 70.94 2.255 70.95 2.754 ;
      RECT 70.925 2.244 70.94 2.755 ;
      RECT 70.92 2.236 70.925 2.753 ;
      RECT 70.91 2.235 70.92 2.745 ;
      RECT 70.88 2.232 70.91 2.724 ;
      RECT 70.805 2.227 70.88 2.669 ;
      RECT 70.79 2.223 70.805 2.615 ;
      RECT 70.78 2.223 70.79 2.51 ;
      RECT 70.765 2.223 70.78 2.443 ;
      RECT 70.75 2.223 70.76 2.433 ;
      RECT 70.695 2.222 70.75 2.43 ;
      RECT 70.65 2.22 70.695 2.433 ;
      RECT 70.622 2.22 70.635 2.436 ;
      RECT 70.536 2.224 70.622 2.438 ;
      RECT 70.45 2.23 70.536 2.443 ;
      RECT 70.43 2.234 70.45 2.445 ;
      RECT 70.428 2.235 70.43 2.444 ;
      RECT 70.342 2.237 70.428 2.443 ;
      RECT 70.256 2.242 70.342 2.44 ;
      RECT 70.17 2.247 70.256 2.437 ;
      RECT 70.02 2.25 70.1 2.433 ;
      RECT 70.68 5.015 70.85 8.305 ;
      RECT 70.68 7.315 71.085 7.645 ;
      RECT 70.68 6.475 71.085 6.805 ;
      RECT 70.796 3.225 70.845 3.559 ;
      RECT 70.796 3.225 70.85 3.558 ;
      RECT 70.71 3.225 70.85 3.557 ;
      RECT 70.485 3.333 70.855 3.555 ;
      RECT 70.71 3.225 70.88 3.548 ;
      RECT 70.68 3.237 70.885 3.539 ;
      RECT 70.665 3.255 70.89 3.536 ;
      RECT 70.48 3.339 70.89 3.463 ;
      RECT 70.475 3.346 70.89 3.423 ;
      RECT 70.49 3.312 70.89 3.536 ;
      RECT 70.651 3.258 70.855 3.555 ;
      RECT 70.565 3.278 70.89 3.536 ;
      RECT 70.665 3.252 70.885 3.539 ;
      RECT 70.435 2.576 70.625 2.77 ;
      RECT 70.43 2.578 70.625 2.769 ;
      RECT 70.425 2.582 70.64 2.766 ;
      RECT 70.44 2.575 70.64 2.766 ;
      RECT 70.425 2.685 70.645 2.761 ;
      RECT 69.72 3.185 69.811 3.483 ;
      RECT 69.715 3.187 69.89 3.478 ;
      RECT 69.72 3.185 69.89 3.478 ;
      RECT 69.715 3.191 69.91 3.476 ;
      RECT 69.715 3.246 69.95 3.475 ;
      RECT 69.715 3.281 69.965 3.469 ;
      RECT 69.715 3.315 69.975 3.459 ;
      RECT 69.705 3.195 69.91 3.31 ;
      RECT 69.705 3.215 69.925 3.31 ;
      RECT 69.705 3.198 69.915 3.31 ;
      RECT 69.93 1.966 69.935 2.028 ;
      RECT 69.925 1.888 69.93 2.051 ;
      RECT 69.92 1.845 69.925 2.062 ;
      RECT 69.915 1.835 69.92 2.074 ;
      RECT 69.91 1.835 69.915 2.083 ;
      RECT 69.885 1.835 69.91 2.115 ;
      RECT 69.88 1.835 69.885 2.148 ;
      RECT 69.865 1.835 69.88 2.173 ;
      RECT 69.855 1.835 69.865 2.2 ;
      RECT 69.85 1.835 69.855 2.213 ;
      RECT 69.845 1.835 69.85 2.228 ;
      RECT 69.835 1.835 69.845 2.243 ;
      RECT 69.83 1.835 69.835 2.263 ;
      RECT 69.805 1.835 69.83 2.298 ;
      RECT 69.76 1.835 69.805 2.343 ;
      RECT 69.75 1.835 69.76 2.356 ;
      RECT 69.665 1.92 69.75 2.363 ;
      RECT 69.63 2.042 69.665 2.372 ;
      RECT 69.625 2.082 69.63 2.376 ;
      RECT 69.605 2.105 69.625 2.378 ;
      RECT 69.6 2.135 69.605 2.381 ;
      RECT 69.59 2.147 69.6 2.382 ;
      RECT 69.545 2.17 69.59 2.387 ;
      RECT 69.505 2.2 69.545 2.395 ;
      RECT 69.47 2.212 69.505 2.401 ;
      RECT 69.465 2.217 69.47 2.405 ;
      RECT 69.395 2.227 69.465 2.412 ;
      RECT 69.355 2.237 69.395 2.422 ;
      RECT 69.335 2.242 69.355 2.428 ;
      RECT 69.325 2.246 69.335 2.433 ;
      RECT 69.32 2.249 69.325 2.436 ;
      RECT 69.31 2.25 69.32 2.437 ;
      RECT 69.285 2.252 69.31 2.441 ;
      RECT 69.275 2.257 69.285 2.444 ;
      RECT 69.23 2.265 69.275 2.445 ;
      RECT 69.105 2.27 69.23 2.445 ;
      RECT 69.66 2.567 69.68 2.749 ;
      RECT 69.611 2.552 69.66 2.748 ;
      RECT 69.525 2.567 69.68 2.746 ;
      RECT 69.51 2.567 69.68 2.745 ;
      RECT 69.475 2.545 69.645 2.73 ;
      RECT 69.545 3.565 69.56 3.774 ;
      RECT 69.545 3.573 69.565 3.773 ;
      RECT 69.49 3.573 69.565 3.772 ;
      RECT 69.47 3.577 69.57 3.77 ;
      RECT 69.45 3.527 69.49 3.769 ;
      RECT 69.395 3.585 69.575 3.767 ;
      RECT 69.36 3.542 69.49 3.765 ;
      RECT 69.356 3.545 69.545 3.764 ;
      RECT 69.27 3.553 69.545 3.762 ;
      RECT 69.27 3.597 69.58 3.755 ;
      RECT 69.26 3.69 69.58 3.753 ;
      RECT 69.27 3.609 69.585 3.738 ;
      RECT 69.27 3.63 69.6 3.708 ;
      RECT 69.27 3.657 69.605 3.678 ;
      RECT 69.395 3.535 69.49 3.767 ;
      RECT 69.025 2.58 69.03 3.118 ;
      RECT 68.83 2.91 68.835 3.105 ;
      RECT 67.13 2.575 67.145 2.955 ;
      RECT 69.195 2.575 69.2 2.745 ;
      RECT 69.19 2.575 69.195 2.755 ;
      RECT 69.185 2.575 69.19 2.768 ;
      RECT 69.16 2.575 69.185 2.81 ;
      RECT 69.135 2.575 69.16 2.883 ;
      RECT 69.12 2.575 69.135 2.935 ;
      RECT 69.115 2.575 69.12 2.965 ;
      RECT 69.09 2.575 69.115 3.005 ;
      RECT 69.075 2.575 69.09 3.06 ;
      RECT 69.07 2.575 69.075 3.093 ;
      RECT 69.045 2.575 69.07 3.113 ;
      RECT 69.03 2.575 69.045 3.119 ;
      RECT 68.96 2.61 69.025 3.115 ;
      RECT 68.91 2.665 68.96 3.11 ;
      RECT 68.9 2.697 68.91 3.108 ;
      RECT 68.895 2.722 68.9 3.108 ;
      RECT 68.875 2.795 68.895 3.108 ;
      RECT 68.865 2.875 68.875 3.107 ;
      RECT 68.85 2.905 68.865 3.107 ;
      RECT 68.835 2.91 68.85 3.106 ;
      RECT 68.775 2.912 68.83 3.103 ;
      RECT 68.745 2.917 68.775 3.099 ;
      RECT 68.743 2.92 68.745 3.098 ;
      RECT 68.657 2.922 68.743 3.095 ;
      RECT 68.571 2.928 68.657 3.089 ;
      RECT 68.485 2.933 68.571 3.083 ;
      RECT 68.412 2.938 68.485 3.084 ;
      RECT 68.326 2.944 68.412 3.092 ;
      RECT 68.24 2.95 68.326 3.101 ;
      RECT 68.22 2.954 68.24 3.106 ;
      RECT 68.173 2.956 68.22 3.109 ;
      RECT 68.087 2.961 68.173 3.115 ;
      RECT 68.001 2.966 68.087 3.124 ;
      RECT 67.915 2.972 68.001 3.132 ;
      RECT 67.83 2.97 67.915 3.141 ;
      RECT 67.826 2.965 67.83 3.145 ;
      RECT 67.74 2.96 67.826 3.137 ;
      RECT 67.676 2.951 67.74 3.125 ;
      RECT 67.59 2.942 67.676 3.112 ;
      RECT 67.566 2.935 67.59 3.103 ;
      RECT 67.48 2.929 67.566 3.09 ;
      RECT 67.44 2.922 67.48 3.076 ;
      RECT 67.435 2.912 67.44 3.072 ;
      RECT 67.425 2.9 67.435 3.071 ;
      RECT 67.405 2.87 67.425 3.068 ;
      RECT 67.35 2.79 67.405 3.062 ;
      RECT 67.33 2.709 67.35 3.057 ;
      RECT 67.31 2.667 67.33 3.053 ;
      RECT 67.285 2.62 67.31 3.047 ;
      RECT 67.28 2.595 67.285 3.044 ;
      RECT 67.245 2.575 67.28 3.039 ;
      RECT 67.236 2.575 67.245 3.032 ;
      RECT 67.15 2.575 67.236 3.002 ;
      RECT 67.145 2.575 67.15 2.965 ;
      RECT 67.11 2.575 67.13 2.887 ;
      RECT 67.105 2.617 67.11 2.852 ;
      RECT 67.1 2.692 67.105 2.808 ;
      RECT 68.55 2.497 68.725 2.745 ;
      RECT 68.55 2.497 68.73 2.743 ;
      RECT 68.545 2.529 68.73 2.703 ;
      RECT 68.575 2.47 68.745 2.69 ;
      RECT 68.54 2.547 68.745 2.623 ;
      RECT 67.85 2.01 68.02 2.185 ;
      RECT 67.85 2.01 68.192 2.177 ;
      RECT 67.85 2.01 68.275 2.171 ;
      RECT 67.85 2.01 68.31 2.167 ;
      RECT 67.85 2.01 68.33 2.166 ;
      RECT 67.85 2.01 68.416 2.162 ;
      RECT 68.31 1.835 68.48 2.157 ;
      RECT 67.885 1.942 68.51 2.155 ;
      RECT 67.875 1.997 68.515 2.153 ;
      RECT 67.85 2.033 68.525 2.148 ;
      RECT 67.85 2.06 68.53 2.078 ;
      RECT 67.915 1.885 68.49 2.155 ;
      RECT 68.106 1.87 68.49 2.155 ;
      RECT 67.94 1.873 68.49 2.155 ;
      RECT 68.02 1.871 68.106 2.182 ;
      RECT 68.106 1.868 68.485 2.155 ;
      RECT 68.29 1.845 68.485 2.155 ;
      RECT 68.192 1.866 68.485 2.155 ;
      RECT 68.275 1.86 68.29 2.168 ;
      RECT 68.425 3.225 68.43 3.425 ;
      RECT 67.89 3.29 67.935 3.425 ;
      RECT 68.46 3.225 68.48 3.398 ;
      RECT 68.43 3.225 68.46 3.413 ;
      RECT 68.365 3.225 68.425 3.45 ;
      RECT 68.35 3.225 68.365 3.48 ;
      RECT 68.335 3.225 68.35 3.493 ;
      RECT 68.315 3.225 68.335 3.508 ;
      RECT 68.31 3.225 68.315 3.517 ;
      RECT 68.3 3.229 68.31 3.522 ;
      RECT 68.285 3.239 68.3 3.533 ;
      RECT 68.26 3.255 68.285 3.543 ;
      RECT 68.25 3.269 68.26 3.545 ;
      RECT 68.23 3.281 68.25 3.542 ;
      RECT 68.2 3.302 68.23 3.536 ;
      RECT 68.19 3.314 68.2 3.531 ;
      RECT 68.18 3.312 68.19 3.528 ;
      RECT 68.165 3.311 68.18 3.523 ;
      RECT 68.16 3.31 68.165 3.518 ;
      RECT 68.125 3.308 68.16 3.508 ;
      RECT 68.105 3.305 68.125 3.49 ;
      RECT 68.095 3.303 68.105 3.485 ;
      RECT 68.085 3.302 68.095 3.48 ;
      RECT 68.05 3.3 68.085 3.468 ;
      RECT 67.995 3.296 68.05 3.448 ;
      RECT 67.985 3.294 67.995 3.433 ;
      RECT 67.98 3.294 67.985 3.428 ;
      RECT 67.935 3.292 67.98 3.425 ;
      RECT 67.84 3.29 67.89 3.429 ;
      RECT 67.83 3.291 67.84 3.434 ;
      RECT 67.77 3.298 67.83 3.448 ;
      RECT 67.745 3.306 67.77 3.468 ;
      RECT 67.735 3.31 67.745 3.48 ;
      RECT 67.73 3.311 67.735 3.485 ;
      RECT 67.715 3.313 67.73 3.488 ;
      RECT 67.7 3.315 67.715 3.493 ;
      RECT 67.695 3.315 67.7 3.496 ;
      RECT 67.65 3.32 67.695 3.507 ;
      RECT 67.645 3.324 67.65 3.519 ;
      RECT 67.62 3.32 67.645 3.523 ;
      RECT 67.61 3.316 67.62 3.527 ;
      RECT 67.6 3.315 67.61 3.531 ;
      RECT 67.585 3.305 67.6 3.537 ;
      RECT 67.58 3.293 67.585 3.541 ;
      RECT 67.575 3.29 67.58 3.542 ;
      RECT 67.57 3.287 67.575 3.544 ;
      RECT 67.555 3.275 67.57 3.543 ;
      RECT 67.54 3.257 67.555 3.54 ;
      RECT 67.52 3.236 67.54 3.533 ;
      RECT 67.455 3.225 67.52 3.505 ;
      RECT 67.451 3.225 67.455 3.484 ;
      RECT 67.365 3.225 67.451 3.454 ;
      RECT 67.35 3.225 67.365 3.41 ;
      RECT 67.925 2.325 67.93 2.56 ;
      RECT 67.055 2.241 67.06 2.445 ;
      RECT 67.635 2.27 67.64 2.425 ;
      RECT 67.555 2.25 67.56 2.425 ;
      RECT 68.225 2.392 68.24 2.745 ;
      RECT 68.151 2.377 68.225 2.745 ;
      RECT 68.065 2.36 68.151 2.745 ;
      RECT 68.055 2.35 68.065 2.743 ;
      RECT 68.05 2.348 68.055 2.738 ;
      RECT 68.035 2.346 68.05 2.724 ;
      RECT 67.965 2.338 68.035 2.664 ;
      RECT 67.945 2.329 67.965 2.598 ;
      RECT 67.94 2.326 67.945 2.578 ;
      RECT 67.93 2.325 67.94 2.568 ;
      RECT 67.92 2.325 67.925 2.552 ;
      RECT 67.91 2.324 67.92 2.542 ;
      RECT 67.9 2.322 67.91 2.53 ;
      RECT 67.885 2.319 67.9 2.51 ;
      RECT 67.875 2.317 67.885 2.495 ;
      RECT 67.855 2.314 67.875 2.483 ;
      RECT 67.85 2.312 67.855 2.473 ;
      RECT 67.825 2.31 67.85 2.46 ;
      RECT 67.795 2.305 67.825 2.445 ;
      RECT 67.715 2.296 67.795 2.436 ;
      RECT 67.67 2.285 67.715 2.429 ;
      RECT 67.65 2.276 67.67 2.426 ;
      RECT 67.64 2.271 67.65 2.425 ;
      RECT 67.595 2.265 67.635 2.425 ;
      RECT 67.58 2.257 67.595 2.425 ;
      RECT 67.56 2.252 67.58 2.425 ;
      RECT 67.54 2.249 67.555 2.425 ;
      RECT 67.457 2.248 67.54 2.424 ;
      RECT 67.371 2.247 67.457 2.42 ;
      RECT 67.285 2.245 67.371 2.417 ;
      RECT 67.232 2.244 67.285 2.419 ;
      RECT 67.146 2.243 67.232 2.428 ;
      RECT 67.06 2.242 67.146 2.44 ;
      RECT 67.04 2.241 67.055 2.448 ;
      RECT 66.96 2.24 67.04 2.46 ;
      RECT 66.935 2.24 66.96 2.473 ;
      RECT 66.91 2.24 66.935 2.488 ;
      RECT 66.905 2.24 66.91 2.51 ;
      RECT 66.9 2.24 66.905 2.528 ;
      RECT 66.895 2.24 66.9 2.545 ;
      RECT 66.89 2.24 66.895 2.558 ;
      RECT 66.885 2.24 66.89 2.568 ;
      RECT 66.845 2.24 66.885 2.653 ;
      RECT 66.83 2.24 66.845 2.738 ;
      RECT 66.82 2.241 66.83 2.75 ;
      RECT 66.785 2.246 66.82 2.755 ;
      RECT 66.745 2.255 66.785 2.755 ;
      RECT 66.73 2.265 66.745 2.755 ;
      RECT 66.725 2.275 66.73 2.755 ;
      RECT 66.705 2.302 66.725 2.755 ;
      RECT 66.655 2.385 66.705 2.755 ;
      RECT 66.65 2.447 66.655 2.755 ;
      RECT 66.64 2.46 66.65 2.755 ;
      RECT 66.63 2.482 66.64 2.755 ;
      RECT 66.62 2.507 66.63 2.75 ;
      RECT 66.615 2.545 66.62 2.743 ;
      RECT 66.605 2.655 66.615 2.738 ;
      RECT 68 3.576 68.015 3.835 ;
      RECT 68 3.591 68.02 3.834 ;
      RECT 67.916 3.591 68.02 3.832 ;
      RECT 67.916 3.605 68.025 3.831 ;
      RECT 67.83 3.647 68.03 3.828 ;
      RECT 67.825 3.59 68.015 3.823 ;
      RECT 67.825 3.661 68.035 3.82 ;
      RECT 67.82 3.692 68.035 3.818 ;
      RECT 67.825 3.689 68.05 3.808 ;
      RECT 67.82 3.735 68.065 3.793 ;
      RECT 67.82 3.763 68.07 3.778 ;
      RECT 67.83 3.565 68 3.828 ;
      RECT 67.59 2.575 67.76 2.745 ;
      RECT 67.555 2.575 67.76 2.74 ;
      RECT 67.545 2.575 67.76 2.733 ;
      RECT 67.54 2.56 67.71 2.73 ;
      RECT 66.37 3.097 66.635 3.54 ;
      RECT 66.365 3.068 66.58 3.538 ;
      RECT 66.36 3.222 66.64 3.533 ;
      RECT 66.365 3.117 66.64 3.533 ;
      RECT 66.365 3.128 66.65 3.52 ;
      RECT 66.365 3.075 66.61 3.538 ;
      RECT 66.37 3.062 66.58 3.54 ;
      RECT 66.37 3.06 66.53 3.54 ;
      RECT 66.471 3.052 66.53 3.54 ;
      RECT 66.385 3.053 66.53 3.54 ;
      RECT 66.471 3.051 66.52 3.54 ;
      RECT 66.275 1.866 66.45 2.165 ;
      RECT 66.325 1.828 66.45 2.165 ;
      RECT 66.31 1.83 66.536 2.157 ;
      RECT 66.31 1.833 66.575 2.144 ;
      RECT 66.31 1.834 66.585 2.13 ;
      RECT 66.265 1.885 66.585 2.12 ;
      RECT 66.31 1.835 66.59 2.115 ;
      RECT 66.265 2.045 66.595 2.105 ;
      RECT 66.25 1.905 66.59 2.045 ;
      RECT 66.245 1.921 66.59 1.985 ;
      RECT 66.29 1.845 66.59 2.115 ;
      RECT 66.325 1.826 66.411 2.165 ;
      RECT 64.785 5.02 64.955 6.49 ;
      RECT 64.785 6.315 64.96 6.485 ;
      RECT 64.415 1.74 64.585 2.93 ;
      RECT 64.415 1.74 64.885 1.91 ;
      RECT 64.415 6.97 64.885 7.14 ;
      RECT 64.415 5.95 64.585 7.14 ;
      RECT 63.425 1.74 63.595 2.93 ;
      RECT 63.425 1.74 63.895 1.91 ;
      RECT 63.425 6.97 63.895 7.14 ;
      RECT 63.425 5.95 63.595 7.14 ;
      RECT 61.575 2.635 61.745 3.865 ;
      RECT 61.63 0.855 61.8 2.805 ;
      RECT 61.575 0.575 61.745 1.025 ;
      RECT 61.575 7.855 61.745 8.305 ;
      RECT 61.63 6.075 61.8 8.025 ;
      RECT 61.575 5.015 61.745 6.245 ;
      RECT 61.055 0.575 61.225 3.865 ;
      RECT 61.055 2.075 61.46 2.405 ;
      RECT 61.055 1.235 61.46 1.565 ;
      RECT 61.055 5.015 61.225 8.305 ;
      RECT 61.055 7.315 61.46 7.645 ;
      RECT 61.055 6.475 61.46 6.805 ;
      RECT 58.98 3.126 58.985 3.298 ;
      RECT 58.975 3.119 58.98 3.388 ;
      RECT 58.97 3.113 58.975 3.407 ;
      RECT 58.95 3.107 58.97 3.417 ;
      RECT 58.935 3.102 58.95 3.425 ;
      RECT 58.898 3.096 58.935 3.423 ;
      RECT 58.812 3.082 58.898 3.419 ;
      RECT 58.726 3.064 58.812 3.414 ;
      RECT 58.64 3.045 58.726 3.408 ;
      RECT 58.61 3.033 58.64 3.404 ;
      RECT 58.59 3.027 58.61 3.403 ;
      RECT 58.525 3.025 58.59 3.401 ;
      RECT 58.51 3.025 58.525 3.393 ;
      RECT 58.495 3.025 58.51 3.38 ;
      RECT 58.49 3.025 58.495 3.37 ;
      RECT 58.475 3.025 58.49 3.348 ;
      RECT 58.46 3.025 58.475 3.315 ;
      RECT 58.455 3.025 58.46 3.293 ;
      RECT 58.445 3.025 58.455 3.275 ;
      RECT 58.43 3.025 58.445 3.253 ;
      RECT 58.41 3.025 58.43 3.215 ;
      RECT 58.76 2.31 58.795 2.749 ;
      RECT 58.76 2.31 58.8 2.748 ;
      RECT 58.705 2.37 58.8 2.747 ;
      RECT 58.57 2.542 58.8 2.746 ;
      RECT 58.68 2.42 58.8 2.746 ;
      RECT 58.57 2.542 58.825 2.736 ;
      RECT 58.625 2.487 58.905 2.653 ;
      RECT 58.8 2.281 58.805 2.744 ;
      RECT 58.655 2.457 58.945 2.53 ;
      RECT 58.67 2.44 58.8 2.746 ;
      RECT 58.805 2.28 58.975 2.468 ;
      RECT 58.795 2.283 58.975 2.468 ;
      RECT 58.3 2.16 58.47 2.47 ;
      RECT 58.3 2.16 58.475 2.443 ;
      RECT 58.3 2.16 58.48 2.42 ;
      RECT 58.3 2.16 58.49 2.37 ;
      RECT 58.295 2.265 58.49 2.34 ;
      RECT 58.33 1.835 58.5 2.313 ;
      RECT 58.33 1.835 58.515 2.234 ;
      RECT 58.32 2.045 58.515 2.234 ;
      RECT 58.33 1.845 58.525 2.149 ;
      RECT 58.26 2.587 58.265 2.79 ;
      RECT 58.25 2.575 58.26 2.9 ;
      RECT 58.225 2.575 58.25 2.94 ;
      RECT 58.145 2.575 58.225 3.025 ;
      RECT 58.135 2.575 58.145 3.095 ;
      RECT 58.11 2.575 58.135 3.118 ;
      RECT 58.09 2.575 58.11 3.153 ;
      RECT 58.045 2.585 58.09 3.196 ;
      RECT 58.035 2.597 58.045 3.233 ;
      RECT 58.015 2.611 58.035 3.253 ;
      RECT 58.005 2.629 58.015 3.269 ;
      RECT 57.99 2.655 58.005 3.279 ;
      RECT 57.975 2.696 57.99 3.293 ;
      RECT 57.965 2.731 57.975 3.303 ;
      RECT 57.96 2.747 57.965 3.308 ;
      RECT 57.95 2.762 57.96 3.313 ;
      RECT 57.93 2.805 57.95 3.323 ;
      RECT 57.91 2.842 57.93 3.336 ;
      RECT 57.875 2.865 57.91 3.354 ;
      RECT 57.865 2.879 57.875 3.37 ;
      RECT 57.845 2.889 57.865 3.38 ;
      RECT 57.84 2.898 57.845 3.388 ;
      RECT 57.83 2.905 57.84 3.395 ;
      RECT 57.82 2.912 57.83 3.403 ;
      RECT 57.805 2.922 57.82 3.411 ;
      RECT 57.795 2.936 57.805 3.421 ;
      RECT 57.785 2.948 57.795 3.433 ;
      RECT 57.77 2.97 57.785 3.446 ;
      RECT 57.76 2.992 57.77 3.457 ;
      RECT 57.75 3.012 57.76 3.466 ;
      RECT 57.745 3.027 57.75 3.473 ;
      RECT 57.715 3.06 57.745 3.487 ;
      RECT 57.705 3.095 57.715 3.502 ;
      RECT 57.7 3.102 57.705 3.508 ;
      RECT 57.68 3.117 57.7 3.515 ;
      RECT 57.675 3.132 57.68 3.523 ;
      RECT 57.67 3.141 57.675 3.528 ;
      RECT 57.655 3.147 57.67 3.535 ;
      RECT 57.65 3.153 57.655 3.543 ;
      RECT 57.645 3.157 57.65 3.55 ;
      RECT 57.64 3.161 57.645 3.56 ;
      RECT 57.63 3.166 57.64 3.57 ;
      RECT 57.61 3.177 57.63 3.598 ;
      RECT 57.595 3.189 57.61 3.625 ;
      RECT 57.575 3.202 57.595 3.65 ;
      RECT 57.555 3.217 57.575 3.674 ;
      RECT 57.54 3.232 57.555 3.689 ;
      RECT 57.535 3.243 57.54 3.698 ;
      RECT 57.47 3.288 57.535 3.708 ;
      RECT 57.435 3.347 57.47 3.721 ;
      RECT 57.43 3.37 57.435 3.727 ;
      RECT 57.425 3.377 57.43 3.729 ;
      RECT 57.41 3.387 57.425 3.732 ;
      RECT 57.38 3.412 57.41 3.736 ;
      RECT 57.375 3.43 57.38 3.74 ;
      RECT 57.37 3.437 57.375 3.741 ;
      RECT 57.35 3.445 57.37 3.745 ;
      RECT 57.34 3.452 57.35 3.749 ;
      RECT 57.296 3.463 57.34 3.756 ;
      RECT 57.21 3.491 57.296 3.772 ;
      RECT 57.15 3.515 57.21 3.79 ;
      RECT 57.105 3.525 57.15 3.804 ;
      RECT 57.046 3.533 57.105 3.818 ;
      RECT 56.96 3.54 57.046 3.837 ;
      RECT 56.935 3.545 56.96 3.852 ;
      RECT 56.855 3.548 56.935 3.855 ;
      RECT 56.775 3.552 56.855 3.842 ;
      RECT 56.766 3.555 56.775 3.827 ;
      RECT 56.68 3.555 56.766 3.812 ;
      RECT 56.62 3.557 56.68 3.789 ;
      RECT 56.616 3.56 56.62 3.779 ;
      RECT 56.53 3.56 56.616 3.764 ;
      RECT 56.455 3.56 56.53 3.74 ;
      RECT 57.77 2.569 57.78 2.745 ;
      RECT 57.725 2.536 57.77 2.745 ;
      RECT 57.68 2.487 57.725 2.745 ;
      RECT 57.65 2.457 57.68 2.746 ;
      RECT 57.645 2.44 57.65 2.747 ;
      RECT 57.62 2.42 57.645 2.748 ;
      RECT 57.605 2.395 57.62 2.749 ;
      RECT 57.6 2.382 57.605 2.75 ;
      RECT 57.595 2.376 57.6 2.748 ;
      RECT 57.59 2.368 57.595 2.742 ;
      RECT 57.565 2.36 57.59 2.722 ;
      RECT 57.545 2.349 57.565 2.693 ;
      RECT 57.515 2.334 57.545 2.664 ;
      RECT 57.495 2.32 57.515 2.636 ;
      RECT 57.485 2.314 57.495 2.615 ;
      RECT 57.48 2.311 57.485 2.598 ;
      RECT 57.475 2.308 57.48 2.583 ;
      RECT 57.46 2.303 57.475 2.548 ;
      RECT 57.455 2.299 57.46 2.515 ;
      RECT 57.435 2.294 57.455 2.491 ;
      RECT 57.405 2.286 57.435 2.456 ;
      RECT 57.39 2.28 57.405 2.433 ;
      RECT 57.35 2.273 57.39 2.418 ;
      RECT 57.325 2.265 57.35 2.398 ;
      RECT 57.305 2.26 57.325 2.388 ;
      RECT 57.27 2.254 57.305 2.383 ;
      RECT 57.225 2.245 57.27 2.382 ;
      RECT 57.195 2.241 57.225 2.384 ;
      RECT 57.11 2.249 57.195 2.388 ;
      RECT 57.04 2.26 57.11 2.41 ;
      RECT 57.027 2.266 57.04 2.433 ;
      RECT 56.941 2.273 57.027 2.455 ;
      RECT 56.855 2.285 56.941 2.492 ;
      RECT 56.855 2.662 56.865 2.9 ;
      RECT 56.85 2.291 56.855 2.515 ;
      RECT 56.845 2.547 56.855 2.9 ;
      RECT 56.845 2.292 56.85 2.52 ;
      RECT 56.84 2.293 56.845 2.9 ;
      RECT 56.816 2.295 56.84 2.901 ;
      RECT 56.73 2.303 56.816 2.903 ;
      RECT 56.71 2.317 56.73 2.906 ;
      RECT 56.705 2.345 56.71 2.907 ;
      RECT 56.7 2.357 56.705 2.908 ;
      RECT 56.695 2.372 56.7 2.909 ;
      RECT 56.685 2.402 56.695 2.91 ;
      RECT 56.68 2.44 56.685 2.908 ;
      RECT 56.675 2.46 56.68 2.903 ;
      RECT 56.66 2.495 56.675 2.888 ;
      RECT 56.65 2.547 56.66 2.868 ;
      RECT 56.645 2.577 56.65 2.856 ;
      RECT 56.63 2.59 56.645 2.839 ;
      RECT 56.605 2.594 56.63 2.806 ;
      RECT 56.59 2.592 56.605 2.783 ;
      RECT 56.575 2.591 56.59 2.78 ;
      RECT 56.515 2.589 56.575 2.778 ;
      RECT 56.505 2.587 56.515 2.773 ;
      RECT 56.465 2.586 56.505 2.77 ;
      RECT 56.395 2.583 56.465 2.768 ;
      RECT 56.34 2.581 56.395 2.763 ;
      RECT 56.27 2.575 56.34 2.758 ;
      RECT 56.261 2.575 56.27 2.755 ;
      RECT 56.175 2.575 56.261 2.75 ;
      RECT 56.17 2.575 56.175 2.745 ;
      RECT 57.475 1.81 57.65 2.16 ;
      RECT 57.475 1.825 57.66 2.158 ;
      RECT 57.45 1.775 57.595 2.155 ;
      RECT 57.43 1.776 57.595 2.148 ;
      RECT 57.42 1.777 57.605 2.143 ;
      RECT 57.39 1.778 57.605 2.13 ;
      RECT 57.34 1.779 57.605 2.106 ;
      RECT 57.335 1.781 57.605 2.091 ;
      RECT 57.335 1.847 57.665 2.085 ;
      RECT 57.315 1.788 57.62 2.065 ;
      RECT 57.305 1.797 57.63 1.92 ;
      RECT 57.315 1.792 57.63 2.065 ;
      RECT 57.335 1.782 57.62 2.091 ;
      RECT 56.92 3.107 57.09 3.395 ;
      RECT 56.915 3.125 57.1 3.39 ;
      RECT 56.88 3.133 57.165 3.31 ;
      RECT 56.88 3.133 57.251 3.3 ;
      RECT 56.88 3.133 57.305 3.246 ;
      RECT 57.165 3.03 57.335 3.214 ;
      RECT 56.88 3.185 57.34 3.202 ;
      RECT 56.865 3.155 57.335 3.198 ;
      RECT 57.125 3.037 57.165 3.349 ;
      RECT 57.005 3.074 57.335 3.214 ;
      RECT 57.1 3.049 57.125 3.375 ;
      RECT 57.09 3.056 57.335 3.214 ;
      RECT 57.221 2.52 57.29 2.779 ;
      RECT 57.221 2.575 57.295 2.778 ;
      RECT 57.135 2.575 57.295 2.777 ;
      RECT 57.13 2.575 57.3 2.77 ;
      RECT 57.12 2.52 57.29 2.765 ;
      RECT 56.5 1.819 56.675 2.12 ;
      RECT 56.485 1.807 56.5 2.105 ;
      RECT 56.455 1.806 56.485 2.058 ;
      RECT 56.455 1.824 56.68 2.053 ;
      RECT 56.44 1.808 56.5 2.018 ;
      RECT 56.435 1.83 56.69 1.918 ;
      RECT 56.435 1.813 56.586 1.918 ;
      RECT 56.435 1.815 56.59 1.918 ;
      RECT 56.44 1.811 56.586 2.018 ;
      RECT 56.545 3.047 56.55 3.395 ;
      RECT 56.535 3.037 56.545 3.401 ;
      RECT 56.5 3.027 56.535 3.403 ;
      RECT 56.462 3.022 56.5 3.407 ;
      RECT 56.376 3.015 56.462 3.414 ;
      RECT 56.29 3.005 56.376 3.424 ;
      RECT 56.245 3 56.29 3.432 ;
      RECT 56.241 3 56.245 3.436 ;
      RECT 56.155 3 56.241 3.443 ;
      RECT 56.14 3 56.155 3.443 ;
      RECT 56.13 2.998 56.14 3.415 ;
      RECT 56.12 2.994 56.13 3.358 ;
      RECT 56.1 2.988 56.12 3.29 ;
      RECT 56.095 2.984 56.1 3.238 ;
      RECT 56.085 2.983 56.095 3.205 ;
      RECT 56.035 2.981 56.085 3.19 ;
      RECT 56.01 2.979 56.035 3.185 ;
      RECT 55.967 2.977 56.01 3.181 ;
      RECT 55.881 2.973 55.967 3.169 ;
      RECT 55.795 2.968 55.881 3.153 ;
      RECT 55.765 2.965 55.795 3.14 ;
      RECT 55.74 2.964 55.765 3.128 ;
      RECT 55.735 2.964 55.74 3.118 ;
      RECT 55.695 2.963 55.735 3.11 ;
      RECT 55.68 2.962 55.695 3.103 ;
      RECT 55.63 2.961 55.68 3.095 ;
      RECT 55.628 2.96 55.63 3.09 ;
      RECT 55.542 2.958 55.628 3.09 ;
      RECT 55.456 2.953 55.542 3.09 ;
      RECT 55.37 2.949 55.456 3.09 ;
      RECT 55.321 2.945 55.37 3.088 ;
      RECT 55.235 2.942 55.321 3.083 ;
      RECT 55.212 2.939 55.235 3.079 ;
      RECT 55.126 2.936 55.212 3.074 ;
      RECT 55.04 2.932 55.126 3.065 ;
      RECT 55.015 2.925 55.04 3.06 ;
      RECT 54.955 2.89 55.015 3.057 ;
      RECT 54.935 2.815 54.955 3.054 ;
      RECT 54.93 2.757 54.935 3.053 ;
      RECT 54.905 2.697 54.93 3.052 ;
      RECT 54.83 2.575 54.905 3.048 ;
      RECT 54.82 2.575 54.83 3.04 ;
      RECT 54.805 2.575 54.82 3.03 ;
      RECT 54.79 2.575 54.805 3 ;
      RECT 54.775 2.575 54.79 2.945 ;
      RECT 54.76 2.575 54.775 2.883 ;
      RECT 54.735 2.575 54.76 2.808 ;
      RECT 54.73 2.575 54.735 2.758 ;
      RECT 56.075 2.12 56.095 2.429 ;
      RECT 56.061 2.122 56.11 2.426 ;
      RECT 56.061 2.127 56.13 2.417 ;
      RECT 55.975 2.125 56.11 2.411 ;
      RECT 55.975 2.133 56.165 2.394 ;
      RECT 55.94 2.135 56.165 2.393 ;
      RECT 55.91 2.143 56.165 2.384 ;
      RECT 55.9 2.148 56.185 2.37 ;
      RECT 55.94 2.138 56.185 2.37 ;
      RECT 55.94 2.141 56.195 2.358 ;
      RECT 55.91 2.143 56.205 2.345 ;
      RECT 55.91 2.147 56.215 2.288 ;
      RECT 55.9 2.152 56.22 2.203 ;
      RECT 56.061 2.12 56.095 2.426 ;
      RECT 55.94 7.855 56.11 8.305 ;
      RECT 55.995 6.075 56.165 8.025 ;
      RECT 55.94 5.015 56.11 6.245 ;
      RECT 55.5 2.223 55.505 2.435 ;
      RECT 55.375 2.22 55.39 2.435 ;
      RECT 54.84 2.25 54.91 2.435 ;
      RECT 54.725 2.25 54.76 2.43 ;
      RECT 55.846 2.552 55.865 2.746 ;
      RECT 55.76 2.507 55.846 2.747 ;
      RECT 55.75 2.46 55.76 2.749 ;
      RECT 55.745 2.44 55.75 2.75 ;
      RECT 55.725 2.405 55.745 2.751 ;
      RECT 55.71 2.355 55.725 2.752 ;
      RECT 55.69 2.292 55.71 2.753 ;
      RECT 55.68 2.255 55.69 2.754 ;
      RECT 55.665 2.244 55.68 2.755 ;
      RECT 55.66 2.236 55.665 2.753 ;
      RECT 55.65 2.235 55.66 2.745 ;
      RECT 55.62 2.232 55.65 2.724 ;
      RECT 55.545 2.227 55.62 2.669 ;
      RECT 55.53 2.223 55.545 2.615 ;
      RECT 55.52 2.223 55.53 2.51 ;
      RECT 55.505 2.223 55.52 2.443 ;
      RECT 55.49 2.223 55.5 2.433 ;
      RECT 55.435 2.222 55.49 2.43 ;
      RECT 55.39 2.22 55.435 2.433 ;
      RECT 55.362 2.22 55.375 2.436 ;
      RECT 55.276 2.224 55.362 2.438 ;
      RECT 55.19 2.23 55.276 2.443 ;
      RECT 55.17 2.234 55.19 2.445 ;
      RECT 55.168 2.235 55.17 2.444 ;
      RECT 55.082 2.237 55.168 2.443 ;
      RECT 54.996 2.242 55.082 2.44 ;
      RECT 54.91 2.247 54.996 2.437 ;
      RECT 54.76 2.25 54.84 2.433 ;
      RECT 55.42 5.015 55.59 8.305 ;
      RECT 55.42 7.315 55.825 7.645 ;
      RECT 55.42 6.475 55.825 6.805 ;
      RECT 55.536 3.225 55.585 3.559 ;
      RECT 55.536 3.225 55.59 3.558 ;
      RECT 55.45 3.225 55.59 3.557 ;
      RECT 55.225 3.333 55.595 3.555 ;
      RECT 55.45 3.225 55.62 3.548 ;
      RECT 55.42 3.237 55.625 3.539 ;
      RECT 55.405 3.255 55.63 3.536 ;
      RECT 55.22 3.339 55.63 3.463 ;
      RECT 55.215 3.346 55.63 3.423 ;
      RECT 55.23 3.312 55.63 3.536 ;
      RECT 55.391 3.258 55.595 3.555 ;
      RECT 55.305 3.278 55.63 3.536 ;
      RECT 55.405 3.252 55.625 3.539 ;
      RECT 55.175 2.576 55.365 2.77 ;
      RECT 55.17 2.578 55.365 2.769 ;
      RECT 55.165 2.582 55.38 2.766 ;
      RECT 55.18 2.575 55.38 2.766 ;
      RECT 55.165 2.685 55.385 2.761 ;
      RECT 54.46 3.185 54.551 3.483 ;
      RECT 54.455 3.187 54.63 3.478 ;
      RECT 54.46 3.185 54.63 3.478 ;
      RECT 54.455 3.191 54.65 3.476 ;
      RECT 54.455 3.246 54.69 3.475 ;
      RECT 54.455 3.281 54.705 3.469 ;
      RECT 54.455 3.315 54.715 3.459 ;
      RECT 54.445 3.195 54.65 3.31 ;
      RECT 54.445 3.215 54.665 3.31 ;
      RECT 54.445 3.198 54.655 3.31 ;
      RECT 54.67 1.966 54.675 2.028 ;
      RECT 54.665 1.888 54.67 2.051 ;
      RECT 54.66 1.845 54.665 2.062 ;
      RECT 54.655 1.835 54.66 2.074 ;
      RECT 54.65 1.835 54.655 2.083 ;
      RECT 54.625 1.835 54.65 2.115 ;
      RECT 54.62 1.835 54.625 2.148 ;
      RECT 54.605 1.835 54.62 2.173 ;
      RECT 54.595 1.835 54.605 2.2 ;
      RECT 54.59 1.835 54.595 2.213 ;
      RECT 54.585 1.835 54.59 2.228 ;
      RECT 54.575 1.835 54.585 2.243 ;
      RECT 54.57 1.835 54.575 2.263 ;
      RECT 54.545 1.835 54.57 2.298 ;
      RECT 54.5 1.835 54.545 2.343 ;
      RECT 54.49 1.835 54.5 2.356 ;
      RECT 54.405 1.92 54.49 2.363 ;
      RECT 54.37 2.042 54.405 2.372 ;
      RECT 54.365 2.082 54.37 2.376 ;
      RECT 54.345 2.105 54.365 2.378 ;
      RECT 54.34 2.135 54.345 2.381 ;
      RECT 54.33 2.147 54.34 2.382 ;
      RECT 54.285 2.17 54.33 2.387 ;
      RECT 54.245 2.2 54.285 2.395 ;
      RECT 54.21 2.212 54.245 2.401 ;
      RECT 54.205 2.217 54.21 2.405 ;
      RECT 54.135 2.227 54.205 2.412 ;
      RECT 54.095 2.237 54.135 2.422 ;
      RECT 54.075 2.242 54.095 2.428 ;
      RECT 54.065 2.246 54.075 2.433 ;
      RECT 54.06 2.249 54.065 2.436 ;
      RECT 54.05 2.25 54.06 2.437 ;
      RECT 54.025 2.252 54.05 2.441 ;
      RECT 54.015 2.257 54.025 2.444 ;
      RECT 53.97 2.265 54.015 2.445 ;
      RECT 53.845 2.27 53.97 2.445 ;
      RECT 54.4 2.567 54.42 2.749 ;
      RECT 54.351 2.552 54.4 2.748 ;
      RECT 54.265 2.567 54.42 2.746 ;
      RECT 54.25 2.567 54.42 2.745 ;
      RECT 54.215 2.545 54.385 2.73 ;
      RECT 54.285 3.565 54.3 3.774 ;
      RECT 54.285 3.573 54.305 3.773 ;
      RECT 54.23 3.573 54.305 3.772 ;
      RECT 54.21 3.577 54.31 3.77 ;
      RECT 54.19 3.527 54.23 3.769 ;
      RECT 54.135 3.585 54.315 3.767 ;
      RECT 54.1 3.542 54.23 3.765 ;
      RECT 54.096 3.545 54.285 3.764 ;
      RECT 54.01 3.553 54.285 3.762 ;
      RECT 54.01 3.597 54.32 3.755 ;
      RECT 54 3.69 54.32 3.753 ;
      RECT 54.01 3.609 54.325 3.738 ;
      RECT 54.01 3.63 54.34 3.708 ;
      RECT 54.01 3.657 54.345 3.678 ;
      RECT 54.135 3.535 54.23 3.767 ;
      RECT 53.765 2.58 53.77 3.118 ;
      RECT 53.57 2.91 53.575 3.105 ;
      RECT 51.87 2.575 51.885 2.955 ;
      RECT 53.935 2.575 53.94 2.745 ;
      RECT 53.93 2.575 53.935 2.755 ;
      RECT 53.925 2.575 53.93 2.768 ;
      RECT 53.9 2.575 53.925 2.81 ;
      RECT 53.875 2.575 53.9 2.883 ;
      RECT 53.86 2.575 53.875 2.935 ;
      RECT 53.855 2.575 53.86 2.965 ;
      RECT 53.83 2.575 53.855 3.005 ;
      RECT 53.815 2.575 53.83 3.06 ;
      RECT 53.81 2.575 53.815 3.093 ;
      RECT 53.785 2.575 53.81 3.113 ;
      RECT 53.77 2.575 53.785 3.119 ;
      RECT 53.7 2.61 53.765 3.115 ;
      RECT 53.65 2.665 53.7 3.11 ;
      RECT 53.64 2.697 53.65 3.108 ;
      RECT 53.635 2.722 53.64 3.108 ;
      RECT 53.615 2.795 53.635 3.108 ;
      RECT 53.605 2.875 53.615 3.107 ;
      RECT 53.59 2.905 53.605 3.107 ;
      RECT 53.575 2.91 53.59 3.106 ;
      RECT 53.515 2.912 53.57 3.103 ;
      RECT 53.485 2.917 53.515 3.099 ;
      RECT 53.483 2.92 53.485 3.098 ;
      RECT 53.397 2.922 53.483 3.095 ;
      RECT 53.311 2.928 53.397 3.089 ;
      RECT 53.225 2.933 53.311 3.083 ;
      RECT 53.152 2.938 53.225 3.084 ;
      RECT 53.066 2.944 53.152 3.092 ;
      RECT 52.98 2.95 53.066 3.101 ;
      RECT 52.96 2.954 52.98 3.106 ;
      RECT 52.913 2.956 52.96 3.109 ;
      RECT 52.827 2.961 52.913 3.115 ;
      RECT 52.741 2.966 52.827 3.124 ;
      RECT 52.655 2.972 52.741 3.132 ;
      RECT 52.57 2.97 52.655 3.141 ;
      RECT 52.566 2.965 52.57 3.145 ;
      RECT 52.48 2.96 52.566 3.137 ;
      RECT 52.416 2.951 52.48 3.125 ;
      RECT 52.33 2.942 52.416 3.112 ;
      RECT 52.306 2.935 52.33 3.103 ;
      RECT 52.22 2.929 52.306 3.09 ;
      RECT 52.18 2.922 52.22 3.076 ;
      RECT 52.175 2.912 52.18 3.072 ;
      RECT 52.165 2.9 52.175 3.071 ;
      RECT 52.145 2.87 52.165 3.068 ;
      RECT 52.09 2.79 52.145 3.062 ;
      RECT 52.07 2.709 52.09 3.057 ;
      RECT 52.05 2.667 52.07 3.053 ;
      RECT 52.025 2.62 52.05 3.047 ;
      RECT 52.02 2.595 52.025 3.044 ;
      RECT 51.985 2.575 52.02 3.039 ;
      RECT 51.976 2.575 51.985 3.032 ;
      RECT 51.89 2.575 51.976 3.002 ;
      RECT 51.885 2.575 51.89 2.965 ;
      RECT 51.85 2.575 51.87 2.887 ;
      RECT 51.845 2.617 51.85 2.852 ;
      RECT 51.84 2.692 51.845 2.808 ;
      RECT 53.29 2.497 53.465 2.745 ;
      RECT 53.29 2.497 53.47 2.743 ;
      RECT 53.285 2.529 53.47 2.703 ;
      RECT 53.315 2.47 53.485 2.69 ;
      RECT 53.28 2.547 53.485 2.623 ;
      RECT 52.59 2.01 52.76 2.185 ;
      RECT 52.59 2.01 52.932 2.177 ;
      RECT 52.59 2.01 53.015 2.171 ;
      RECT 52.59 2.01 53.05 2.167 ;
      RECT 52.59 2.01 53.07 2.166 ;
      RECT 52.59 2.01 53.156 2.162 ;
      RECT 53.05 1.835 53.22 2.157 ;
      RECT 52.625 1.942 53.25 2.155 ;
      RECT 52.615 1.997 53.255 2.153 ;
      RECT 52.59 2.033 53.265 2.148 ;
      RECT 52.59 2.06 53.27 2.078 ;
      RECT 52.655 1.885 53.23 2.155 ;
      RECT 52.846 1.87 53.23 2.155 ;
      RECT 52.68 1.873 53.23 2.155 ;
      RECT 52.76 1.871 52.846 2.182 ;
      RECT 52.846 1.868 53.225 2.155 ;
      RECT 53.03 1.845 53.225 2.155 ;
      RECT 52.932 1.866 53.225 2.155 ;
      RECT 53.015 1.86 53.03 2.168 ;
      RECT 53.165 3.225 53.17 3.425 ;
      RECT 52.63 3.29 52.675 3.425 ;
      RECT 53.2 3.225 53.22 3.398 ;
      RECT 53.17 3.225 53.2 3.413 ;
      RECT 53.105 3.225 53.165 3.45 ;
      RECT 53.09 3.225 53.105 3.48 ;
      RECT 53.075 3.225 53.09 3.493 ;
      RECT 53.055 3.225 53.075 3.508 ;
      RECT 53.05 3.225 53.055 3.517 ;
      RECT 53.04 3.229 53.05 3.522 ;
      RECT 53.025 3.239 53.04 3.533 ;
      RECT 53 3.255 53.025 3.543 ;
      RECT 52.99 3.269 53 3.545 ;
      RECT 52.97 3.281 52.99 3.542 ;
      RECT 52.94 3.302 52.97 3.536 ;
      RECT 52.93 3.314 52.94 3.531 ;
      RECT 52.92 3.312 52.93 3.528 ;
      RECT 52.905 3.311 52.92 3.523 ;
      RECT 52.9 3.31 52.905 3.518 ;
      RECT 52.865 3.308 52.9 3.508 ;
      RECT 52.845 3.305 52.865 3.49 ;
      RECT 52.835 3.303 52.845 3.485 ;
      RECT 52.825 3.302 52.835 3.48 ;
      RECT 52.79 3.3 52.825 3.468 ;
      RECT 52.735 3.296 52.79 3.448 ;
      RECT 52.725 3.294 52.735 3.433 ;
      RECT 52.72 3.294 52.725 3.428 ;
      RECT 52.675 3.292 52.72 3.425 ;
      RECT 52.58 3.29 52.63 3.429 ;
      RECT 52.57 3.291 52.58 3.434 ;
      RECT 52.51 3.298 52.57 3.448 ;
      RECT 52.485 3.306 52.51 3.468 ;
      RECT 52.475 3.31 52.485 3.48 ;
      RECT 52.47 3.311 52.475 3.485 ;
      RECT 52.455 3.313 52.47 3.488 ;
      RECT 52.44 3.315 52.455 3.493 ;
      RECT 52.435 3.315 52.44 3.496 ;
      RECT 52.39 3.32 52.435 3.507 ;
      RECT 52.385 3.324 52.39 3.519 ;
      RECT 52.36 3.32 52.385 3.523 ;
      RECT 52.35 3.316 52.36 3.527 ;
      RECT 52.34 3.315 52.35 3.531 ;
      RECT 52.325 3.305 52.34 3.537 ;
      RECT 52.32 3.293 52.325 3.541 ;
      RECT 52.315 3.29 52.32 3.542 ;
      RECT 52.31 3.287 52.315 3.544 ;
      RECT 52.295 3.275 52.31 3.543 ;
      RECT 52.28 3.257 52.295 3.54 ;
      RECT 52.26 3.236 52.28 3.533 ;
      RECT 52.195 3.225 52.26 3.505 ;
      RECT 52.191 3.225 52.195 3.484 ;
      RECT 52.105 3.225 52.191 3.454 ;
      RECT 52.09 3.225 52.105 3.41 ;
      RECT 52.665 2.325 52.67 2.56 ;
      RECT 51.795 2.241 51.8 2.445 ;
      RECT 52.375 2.27 52.38 2.425 ;
      RECT 52.295 2.25 52.3 2.425 ;
      RECT 52.965 2.392 52.98 2.745 ;
      RECT 52.891 2.377 52.965 2.745 ;
      RECT 52.805 2.36 52.891 2.745 ;
      RECT 52.795 2.35 52.805 2.743 ;
      RECT 52.79 2.348 52.795 2.738 ;
      RECT 52.775 2.346 52.79 2.724 ;
      RECT 52.705 2.338 52.775 2.664 ;
      RECT 52.685 2.329 52.705 2.598 ;
      RECT 52.68 2.326 52.685 2.578 ;
      RECT 52.67 2.325 52.68 2.568 ;
      RECT 52.66 2.325 52.665 2.552 ;
      RECT 52.65 2.324 52.66 2.542 ;
      RECT 52.64 2.322 52.65 2.53 ;
      RECT 52.625 2.319 52.64 2.51 ;
      RECT 52.615 2.317 52.625 2.495 ;
      RECT 52.595 2.314 52.615 2.483 ;
      RECT 52.59 2.312 52.595 2.473 ;
      RECT 52.565 2.31 52.59 2.46 ;
      RECT 52.535 2.305 52.565 2.445 ;
      RECT 52.455 2.296 52.535 2.436 ;
      RECT 52.41 2.285 52.455 2.429 ;
      RECT 52.39 2.276 52.41 2.426 ;
      RECT 52.38 2.271 52.39 2.425 ;
      RECT 52.335 2.265 52.375 2.425 ;
      RECT 52.32 2.257 52.335 2.425 ;
      RECT 52.3 2.252 52.32 2.425 ;
      RECT 52.28 2.249 52.295 2.425 ;
      RECT 52.197 2.248 52.28 2.424 ;
      RECT 52.111 2.247 52.197 2.42 ;
      RECT 52.025 2.245 52.111 2.417 ;
      RECT 51.972 2.244 52.025 2.419 ;
      RECT 51.886 2.243 51.972 2.428 ;
      RECT 51.8 2.242 51.886 2.44 ;
      RECT 51.78 2.241 51.795 2.448 ;
      RECT 51.7 2.24 51.78 2.46 ;
      RECT 51.675 2.24 51.7 2.473 ;
      RECT 51.65 2.24 51.675 2.488 ;
      RECT 51.645 2.24 51.65 2.51 ;
      RECT 51.64 2.24 51.645 2.528 ;
      RECT 51.635 2.24 51.64 2.545 ;
      RECT 51.63 2.24 51.635 2.558 ;
      RECT 51.625 2.24 51.63 2.568 ;
      RECT 51.585 2.24 51.625 2.653 ;
      RECT 51.57 2.24 51.585 2.738 ;
      RECT 51.56 2.241 51.57 2.75 ;
      RECT 51.525 2.246 51.56 2.755 ;
      RECT 51.485 2.255 51.525 2.755 ;
      RECT 51.47 2.265 51.485 2.755 ;
      RECT 51.465 2.275 51.47 2.755 ;
      RECT 51.445 2.302 51.465 2.755 ;
      RECT 51.395 2.385 51.445 2.755 ;
      RECT 51.39 2.447 51.395 2.755 ;
      RECT 51.38 2.46 51.39 2.755 ;
      RECT 51.37 2.482 51.38 2.755 ;
      RECT 51.36 2.507 51.37 2.75 ;
      RECT 51.355 2.545 51.36 2.743 ;
      RECT 51.345 2.655 51.355 2.738 ;
      RECT 52.74 3.576 52.755 3.835 ;
      RECT 52.74 3.591 52.76 3.834 ;
      RECT 52.656 3.591 52.76 3.832 ;
      RECT 52.656 3.605 52.765 3.831 ;
      RECT 52.57 3.647 52.77 3.828 ;
      RECT 52.565 3.59 52.755 3.823 ;
      RECT 52.565 3.661 52.775 3.82 ;
      RECT 52.56 3.692 52.775 3.818 ;
      RECT 52.565 3.689 52.79 3.808 ;
      RECT 52.56 3.735 52.805 3.793 ;
      RECT 52.56 3.763 52.81 3.778 ;
      RECT 52.57 3.565 52.74 3.828 ;
      RECT 52.33 2.575 52.5 2.745 ;
      RECT 52.295 2.575 52.5 2.74 ;
      RECT 52.285 2.575 52.5 2.733 ;
      RECT 52.28 2.56 52.45 2.73 ;
      RECT 51.11 3.097 51.375 3.54 ;
      RECT 51.105 3.068 51.32 3.538 ;
      RECT 51.1 3.222 51.38 3.533 ;
      RECT 51.105 3.117 51.38 3.533 ;
      RECT 51.105 3.128 51.39 3.52 ;
      RECT 51.105 3.075 51.35 3.538 ;
      RECT 51.11 3.062 51.32 3.54 ;
      RECT 51.11 3.06 51.27 3.54 ;
      RECT 51.211 3.052 51.27 3.54 ;
      RECT 51.125 3.053 51.27 3.54 ;
      RECT 51.211 3.051 51.26 3.54 ;
      RECT 51.015 1.866 51.19 2.165 ;
      RECT 51.065 1.828 51.19 2.165 ;
      RECT 51.05 1.83 51.276 2.157 ;
      RECT 51.05 1.833 51.315 2.144 ;
      RECT 51.05 1.834 51.325 2.13 ;
      RECT 51.005 1.885 51.325 2.12 ;
      RECT 51.05 1.835 51.33 2.115 ;
      RECT 51.005 2.045 51.335 2.105 ;
      RECT 50.99 1.905 51.33 2.045 ;
      RECT 50.985 1.921 51.33 1.985 ;
      RECT 51.03 1.845 51.33 2.115 ;
      RECT 51.065 1.826 51.151 2.165 ;
      RECT 49.525 5.02 49.695 6.49 ;
      RECT 49.525 6.315 49.7 6.485 ;
      RECT 49.155 1.74 49.325 2.93 ;
      RECT 49.155 1.74 49.625 1.91 ;
      RECT 49.155 6.97 49.625 7.14 ;
      RECT 49.155 5.95 49.325 7.14 ;
      RECT 48.165 1.74 48.335 2.93 ;
      RECT 48.165 1.74 48.635 1.91 ;
      RECT 48.165 6.97 48.635 7.14 ;
      RECT 48.165 5.95 48.335 7.14 ;
      RECT 46.315 2.635 46.485 3.865 ;
      RECT 46.37 0.855 46.54 2.805 ;
      RECT 46.315 0.575 46.485 1.025 ;
      RECT 46.315 7.855 46.485 8.305 ;
      RECT 46.37 6.075 46.54 8.025 ;
      RECT 46.315 5.015 46.485 6.245 ;
      RECT 45.795 0.575 45.965 3.865 ;
      RECT 45.795 2.075 46.2 2.405 ;
      RECT 45.795 1.235 46.2 1.565 ;
      RECT 45.795 5.015 45.965 8.305 ;
      RECT 45.795 7.315 46.2 7.645 ;
      RECT 45.795 6.475 46.2 6.805 ;
      RECT 43.72 3.126 43.725 3.298 ;
      RECT 43.715 3.119 43.72 3.388 ;
      RECT 43.71 3.113 43.715 3.407 ;
      RECT 43.69 3.107 43.71 3.417 ;
      RECT 43.675 3.102 43.69 3.425 ;
      RECT 43.638 3.096 43.675 3.423 ;
      RECT 43.552 3.082 43.638 3.419 ;
      RECT 43.466 3.064 43.552 3.414 ;
      RECT 43.38 3.045 43.466 3.408 ;
      RECT 43.35 3.033 43.38 3.404 ;
      RECT 43.33 3.027 43.35 3.403 ;
      RECT 43.265 3.025 43.33 3.401 ;
      RECT 43.25 3.025 43.265 3.393 ;
      RECT 43.235 3.025 43.25 3.38 ;
      RECT 43.23 3.025 43.235 3.37 ;
      RECT 43.215 3.025 43.23 3.348 ;
      RECT 43.2 3.025 43.215 3.315 ;
      RECT 43.195 3.025 43.2 3.293 ;
      RECT 43.185 3.025 43.195 3.275 ;
      RECT 43.17 3.025 43.185 3.253 ;
      RECT 43.15 3.025 43.17 3.215 ;
      RECT 43.5 2.31 43.535 2.749 ;
      RECT 43.5 2.31 43.54 2.748 ;
      RECT 43.445 2.37 43.54 2.747 ;
      RECT 43.31 2.542 43.54 2.746 ;
      RECT 43.42 2.42 43.54 2.746 ;
      RECT 43.31 2.542 43.565 2.736 ;
      RECT 43.365 2.487 43.645 2.653 ;
      RECT 43.54 2.281 43.545 2.744 ;
      RECT 43.395 2.457 43.685 2.53 ;
      RECT 43.41 2.44 43.54 2.746 ;
      RECT 43.545 2.28 43.715 2.468 ;
      RECT 43.535 2.283 43.715 2.468 ;
      RECT 43.04 2.16 43.21 2.47 ;
      RECT 43.04 2.16 43.215 2.443 ;
      RECT 43.04 2.16 43.22 2.42 ;
      RECT 43.04 2.16 43.23 2.37 ;
      RECT 43.035 2.265 43.23 2.34 ;
      RECT 43.07 1.835 43.24 2.313 ;
      RECT 43.07 1.835 43.255 2.234 ;
      RECT 43.06 2.045 43.255 2.234 ;
      RECT 43.07 1.845 43.265 2.149 ;
      RECT 43 2.587 43.005 2.79 ;
      RECT 42.99 2.575 43 2.9 ;
      RECT 42.965 2.575 42.99 2.94 ;
      RECT 42.885 2.575 42.965 3.025 ;
      RECT 42.875 2.575 42.885 3.095 ;
      RECT 42.85 2.575 42.875 3.118 ;
      RECT 42.83 2.575 42.85 3.153 ;
      RECT 42.785 2.585 42.83 3.196 ;
      RECT 42.775 2.597 42.785 3.233 ;
      RECT 42.755 2.611 42.775 3.253 ;
      RECT 42.745 2.629 42.755 3.269 ;
      RECT 42.73 2.655 42.745 3.279 ;
      RECT 42.715 2.696 42.73 3.293 ;
      RECT 42.705 2.731 42.715 3.303 ;
      RECT 42.7 2.747 42.705 3.308 ;
      RECT 42.69 2.762 42.7 3.313 ;
      RECT 42.67 2.805 42.69 3.323 ;
      RECT 42.65 2.842 42.67 3.336 ;
      RECT 42.615 2.865 42.65 3.354 ;
      RECT 42.605 2.879 42.615 3.37 ;
      RECT 42.585 2.889 42.605 3.38 ;
      RECT 42.58 2.898 42.585 3.388 ;
      RECT 42.57 2.905 42.58 3.395 ;
      RECT 42.56 2.912 42.57 3.403 ;
      RECT 42.545 2.922 42.56 3.411 ;
      RECT 42.535 2.936 42.545 3.421 ;
      RECT 42.525 2.948 42.535 3.433 ;
      RECT 42.51 2.97 42.525 3.446 ;
      RECT 42.5 2.992 42.51 3.457 ;
      RECT 42.49 3.012 42.5 3.466 ;
      RECT 42.485 3.027 42.49 3.473 ;
      RECT 42.455 3.06 42.485 3.487 ;
      RECT 42.445 3.095 42.455 3.502 ;
      RECT 42.44 3.102 42.445 3.508 ;
      RECT 42.42 3.117 42.44 3.515 ;
      RECT 42.415 3.132 42.42 3.523 ;
      RECT 42.41 3.141 42.415 3.528 ;
      RECT 42.395 3.147 42.41 3.535 ;
      RECT 42.39 3.153 42.395 3.543 ;
      RECT 42.385 3.157 42.39 3.55 ;
      RECT 42.38 3.161 42.385 3.56 ;
      RECT 42.37 3.166 42.38 3.57 ;
      RECT 42.35 3.177 42.37 3.598 ;
      RECT 42.335 3.189 42.35 3.625 ;
      RECT 42.315 3.202 42.335 3.65 ;
      RECT 42.295 3.217 42.315 3.674 ;
      RECT 42.28 3.232 42.295 3.689 ;
      RECT 42.275 3.243 42.28 3.698 ;
      RECT 42.21 3.288 42.275 3.708 ;
      RECT 42.175 3.347 42.21 3.721 ;
      RECT 42.17 3.37 42.175 3.727 ;
      RECT 42.165 3.377 42.17 3.729 ;
      RECT 42.15 3.387 42.165 3.732 ;
      RECT 42.12 3.412 42.15 3.736 ;
      RECT 42.115 3.43 42.12 3.74 ;
      RECT 42.11 3.437 42.115 3.741 ;
      RECT 42.09 3.445 42.11 3.745 ;
      RECT 42.08 3.452 42.09 3.749 ;
      RECT 42.036 3.463 42.08 3.756 ;
      RECT 41.95 3.491 42.036 3.772 ;
      RECT 41.89 3.515 41.95 3.79 ;
      RECT 41.845 3.525 41.89 3.804 ;
      RECT 41.786 3.533 41.845 3.818 ;
      RECT 41.7 3.54 41.786 3.837 ;
      RECT 41.675 3.545 41.7 3.852 ;
      RECT 41.595 3.548 41.675 3.855 ;
      RECT 41.515 3.552 41.595 3.842 ;
      RECT 41.506 3.555 41.515 3.827 ;
      RECT 41.42 3.555 41.506 3.812 ;
      RECT 41.36 3.557 41.42 3.789 ;
      RECT 41.356 3.56 41.36 3.779 ;
      RECT 41.27 3.56 41.356 3.764 ;
      RECT 41.195 3.56 41.27 3.74 ;
      RECT 42.51 2.569 42.52 2.745 ;
      RECT 42.465 2.536 42.51 2.745 ;
      RECT 42.42 2.487 42.465 2.745 ;
      RECT 42.39 2.457 42.42 2.746 ;
      RECT 42.385 2.44 42.39 2.747 ;
      RECT 42.36 2.42 42.385 2.748 ;
      RECT 42.345 2.395 42.36 2.749 ;
      RECT 42.34 2.382 42.345 2.75 ;
      RECT 42.335 2.376 42.34 2.748 ;
      RECT 42.33 2.368 42.335 2.742 ;
      RECT 42.305 2.36 42.33 2.722 ;
      RECT 42.285 2.349 42.305 2.693 ;
      RECT 42.255 2.334 42.285 2.664 ;
      RECT 42.235 2.32 42.255 2.636 ;
      RECT 42.225 2.314 42.235 2.615 ;
      RECT 42.22 2.311 42.225 2.598 ;
      RECT 42.215 2.308 42.22 2.583 ;
      RECT 42.2 2.303 42.215 2.548 ;
      RECT 42.195 2.299 42.2 2.515 ;
      RECT 42.175 2.294 42.195 2.491 ;
      RECT 42.145 2.286 42.175 2.456 ;
      RECT 42.13 2.28 42.145 2.433 ;
      RECT 42.09 2.273 42.13 2.418 ;
      RECT 42.065 2.265 42.09 2.398 ;
      RECT 42.045 2.26 42.065 2.388 ;
      RECT 42.01 2.254 42.045 2.383 ;
      RECT 41.965 2.245 42.01 2.382 ;
      RECT 41.935 2.241 41.965 2.384 ;
      RECT 41.85 2.249 41.935 2.388 ;
      RECT 41.78 2.26 41.85 2.41 ;
      RECT 41.767 2.266 41.78 2.433 ;
      RECT 41.681 2.273 41.767 2.455 ;
      RECT 41.595 2.285 41.681 2.492 ;
      RECT 41.595 2.662 41.605 2.9 ;
      RECT 41.59 2.291 41.595 2.515 ;
      RECT 41.585 2.547 41.595 2.9 ;
      RECT 41.585 2.292 41.59 2.52 ;
      RECT 41.58 2.293 41.585 2.9 ;
      RECT 41.556 2.295 41.58 2.901 ;
      RECT 41.47 2.303 41.556 2.903 ;
      RECT 41.45 2.317 41.47 2.906 ;
      RECT 41.445 2.345 41.45 2.907 ;
      RECT 41.44 2.357 41.445 2.908 ;
      RECT 41.435 2.372 41.44 2.909 ;
      RECT 41.425 2.402 41.435 2.91 ;
      RECT 41.42 2.44 41.425 2.908 ;
      RECT 41.415 2.46 41.42 2.903 ;
      RECT 41.4 2.495 41.415 2.888 ;
      RECT 41.39 2.547 41.4 2.868 ;
      RECT 41.385 2.577 41.39 2.856 ;
      RECT 41.37 2.59 41.385 2.839 ;
      RECT 41.345 2.594 41.37 2.806 ;
      RECT 41.33 2.592 41.345 2.783 ;
      RECT 41.315 2.591 41.33 2.78 ;
      RECT 41.255 2.589 41.315 2.778 ;
      RECT 41.245 2.587 41.255 2.773 ;
      RECT 41.205 2.586 41.245 2.77 ;
      RECT 41.135 2.583 41.205 2.768 ;
      RECT 41.08 2.581 41.135 2.763 ;
      RECT 41.01 2.575 41.08 2.758 ;
      RECT 41.001 2.575 41.01 2.755 ;
      RECT 40.915 2.575 41.001 2.75 ;
      RECT 40.91 2.575 40.915 2.745 ;
      RECT 42.215 1.81 42.39 2.16 ;
      RECT 42.215 1.825 42.4 2.158 ;
      RECT 42.19 1.775 42.335 2.155 ;
      RECT 42.17 1.776 42.335 2.148 ;
      RECT 42.16 1.777 42.345 2.143 ;
      RECT 42.13 1.778 42.345 2.13 ;
      RECT 42.08 1.779 42.345 2.106 ;
      RECT 42.075 1.781 42.345 2.091 ;
      RECT 42.075 1.847 42.405 2.085 ;
      RECT 42.055 1.788 42.36 2.065 ;
      RECT 42.045 1.797 42.37 1.92 ;
      RECT 42.055 1.792 42.37 2.065 ;
      RECT 42.075 1.782 42.36 2.091 ;
      RECT 41.66 3.107 41.83 3.395 ;
      RECT 41.655 3.125 41.84 3.39 ;
      RECT 41.62 3.133 41.905 3.31 ;
      RECT 41.62 3.133 41.991 3.3 ;
      RECT 41.62 3.133 42.045 3.246 ;
      RECT 41.905 3.03 42.075 3.214 ;
      RECT 41.62 3.185 42.08 3.202 ;
      RECT 41.605 3.155 42.075 3.198 ;
      RECT 41.865 3.037 41.905 3.349 ;
      RECT 41.745 3.074 42.075 3.214 ;
      RECT 41.84 3.049 41.865 3.375 ;
      RECT 41.83 3.056 42.075 3.214 ;
      RECT 41.961 2.52 42.03 2.779 ;
      RECT 41.961 2.575 42.035 2.778 ;
      RECT 41.875 2.575 42.035 2.777 ;
      RECT 41.87 2.575 42.04 2.77 ;
      RECT 41.86 2.52 42.03 2.765 ;
      RECT 41.24 1.819 41.415 2.12 ;
      RECT 41.225 1.807 41.24 2.105 ;
      RECT 41.195 1.806 41.225 2.058 ;
      RECT 41.195 1.824 41.42 2.053 ;
      RECT 41.18 1.808 41.24 2.018 ;
      RECT 41.175 1.83 41.43 1.918 ;
      RECT 41.175 1.813 41.326 1.918 ;
      RECT 41.175 1.815 41.33 1.918 ;
      RECT 41.18 1.811 41.326 2.018 ;
      RECT 41.285 3.047 41.29 3.395 ;
      RECT 41.275 3.037 41.285 3.401 ;
      RECT 41.24 3.027 41.275 3.403 ;
      RECT 41.202 3.022 41.24 3.407 ;
      RECT 41.116 3.015 41.202 3.414 ;
      RECT 41.03 3.005 41.116 3.424 ;
      RECT 40.985 3 41.03 3.432 ;
      RECT 40.981 3 40.985 3.436 ;
      RECT 40.895 3 40.981 3.443 ;
      RECT 40.88 3 40.895 3.443 ;
      RECT 40.87 2.998 40.88 3.415 ;
      RECT 40.86 2.994 40.87 3.358 ;
      RECT 40.84 2.988 40.86 3.29 ;
      RECT 40.835 2.984 40.84 3.238 ;
      RECT 40.825 2.983 40.835 3.205 ;
      RECT 40.775 2.981 40.825 3.19 ;
      RECT 40.75 2.979 40.775 3.185 ;
      RECT 40.707 2.977 40.75 3.181 ;
      RECT 40.621 2.973 40.707 3.169 ;
      RECT 40.535 2.968 40.621 3.153 ;
      RECT 40.505 2.965 40.535 3.14 ;
      RECT 40.48 2.964 40.505 3.128 ;
      RECT 40.475 2.964 40.48 3.118 ;
      RECT 40.435 2.963 40.475 3.11 ;
      RECT 40.42 2.962 40.435 3.103 ;
      RECT 40.37 2.961 40.42 3.095 ;
      RECT 40.368 2.96 40.37 3.09 ;
      RECT 40.282 2.958 40.368 3.09 ;
      RECT 40.196 2.953 40.282 3.09 ;
      RECT 40.11 2.949 40.196 3.09 ;
      RECT 40.061 2.945 40.11 3.088 ;
      RECT 39.975 2.942 40.061 3.083 ;
      RECT 39.952 2.939 39.975 3.079 ;
      RECT 39.866 2.936 39.952 3.074 ;
      RECT 39.78 2.932 39.866 3.065 ;
      RECT 39.755 2.925 39.78 3.06 ;
      RECT 39.695 2.89 39.755 3.057 ;
      RECT 39.675 2.815 39.695 3.054 ;
      RECT 39.67 2.757 39.675 3.053 ;
      RECT 39.645 2.697 39.67 3.052 ;
      RECT 39.57 2.575 39.645 3.048 ;
      RECT 39.56 2.575 39.57 3.04 ;
      RECT 39.545 2.575 39.56 3.03 ;
      RECT 39.53 2.575 39.545 3 ;
      RECT 39.515 2.575 39.53 2.945 ;
      RECT 39.5 2.575 39.515 2.883 ;
      RECT 39.475 2.575 39.5 2.808 ;
      RECT 39.47 2.575 39.475 2.758 ;
      RECT 40.815 2.12 40.835 2.429 ;
      RECT 40.801 2.122 40.85 2.426 ;
      RECT 40.801 2.127 40.87 2.417 ;
      RECT 40.715 2.125 40.85 2.411 ;
      RECT 40.715 2.133 40.905 2.394 ;
      RECT 40.68 2.135 40.905 2.393 ;
      RECT 40.65 2.143 40.905 2.384 ;
      RECT 40.64 2.148 40.925 2.37 ;
      RECT 40.68 2.138 40.925 2.37 ;
      RECT 40.68 2.141 40.935 2.358 ;
      RECT 40.65 2.143 40.945 2.345 ;
      RECT 40.65 2.147 40.955 2.288 ;
      RECT 40.64 2.152 40.96 2.203 ;
      RECT 40.801 2.12 40.835 2.426 ;
      RECT 40.68 7.855 40.85 8.305 ;
      RECT 40.735 6.075 40.905 8.025 ;
      RECT 40.68 5.015 40.85 6.245 ;
      RECT 40.24 2.223 40.245 2.435 ;
      RECT 40.115 2.22 40.13 2.435 ;
      RECT 39.58 2.25 39.65 2.435 ;
      RECT 39.465 2.25 39.5 2.43 ;
      RECT 40.586 2.552 40.605 2.746 ;
      RECT 40.5 2.507 40.586 2.747 ;
      RECT 40.49 2.46 40.5 2.749 ;
      RECT 40.485 2.44 40.49 2.75 ;
      RECT 40.465 2.405 40.485 2.751 ;
      RECT 40.45 2.355 40.465 2.752 ;
      RECT 40.43 2.292 40.45 2.753 ;
      RECT 40.42 2.255 40.43 2.754 ;
      RECT 40.405 2.244 40.42 2.755 ;
      RECT 40.4 2.236 40.405 2.753 ;
      RECT 40.39 2.235 40.4 2.745 ;
      RECT 40.36 2.232 40.39 2.724 ;
      RECT 40.285 2.227 40.36 2.669 ;
      RECT 40.27 2.223 40.285 2.615 ;
      RECT 40.26 2.223 40.27 2.51 ;
      RECT 40.245 2.223 40.26 2.443 ;
      RECT 40.23 2.223 40.24 2.433 ;
      RECT 40.175 2.222 40.23 2.43 ;
      RECT 40.13 2.22 40.175 2.433 ;
      RECT 40.102 2.22 40.115 2.436 ;
      RECT 40.016 2.224 40.102 2.438 ;
      RECT 39.93 2.23 40.016 2.443 ;
      RECT 39.91 2.234 39.93 2.445 ;
      RECT 39.908 2.235 39.91 2.444 ;
      RECT 39.822 2.237 39.908 2.443 ;
      RECT 39.736 2.242 39.822 2.44 ;
      RECT 39.65 2.247 39.736 2.437 ;
      RECT 39.5 2.25 39.58 2.433 ;
      RECT 40.16 5.015 40.33 8.305 ;
      RECT 40.16 7.315 40.565 7.645 ;
      RECT 40.16 6.475 40.565 6.805 ;
      RECT 40.276 3.225 40.325 3.559 ;
      RECT 40.276 3.225 40.33 3.558 ;
      RECT 40.19 3.225 40.33 3.557 ;
      RECT 39.965 3.333 40.335 3.555 ;
      RECT 40.19 3.225 40.36 3.548 ;
      RECT 40.16 3.237 40.365 3.539 ;
      RECT 40.145 3.255 40.37 3.536 ;
      RECT 39.96 3.339 40.37 3.463 ;
      RECT 39.955 3.346 40.37 3.423 ;
      RECT 39.97 3.312 40.37 3.536 ;
      RECT 40.131 3.258 40.335 3.555 ;
      RECT 40.045 3.278 40.37 3.536 ;
      RECT 40.145 3.252 40.365 3.539 ;
      RECT 39.915 2.576 40.105 2.77 ;
      RECT 39.91 2.578 40.105 2.769 ;
      RECT 39.905 2.582 40.12 2.766 ;
      RECT 39.92 2.575 40.12 2.766 ;
      RECT 39.905 2.685 40.125 2.761 ;
      RECT 39.2 3.185 39.291 3.483 ;
      RECT 39.195 3.187 39.37 3.478 ;
      RECT 39.2 3.185 39.37 3.478 ;
      RECT 39.195 3.191 39.39 3.476 ;
      RECT 39.195 3.246 39.43 3.475 ;
      RECT 39.195 3.281 39.445 3.469 ;
      RECT 39.195 3.315 39.455 3.459 ;
      RECT 39.185 3.195 39.39 3.31 ;
      RECT 39.185 3.215 39.405 3.31 ;
      RECT 39.185 3.198 39.395 3.31 ;
      RECT 39.41 1.966 39.415 2.028 ;
      RECT 39.405 1.888 39.41 2.051 ;
      RECT 39.4 1.845 39.405 2.062 ;
      RECT 39.395 1.835 39.4 2.074 ;
      RECT 39.39 1.835 39.395 2.083 ;
      RECT 39.365 1.835 39.39 2.115 ;
      RECT 39.36 1.835 39.365 2.148 ;
      RECT 39.345 1.835 39.36 2.173 ;
      RECT 39.335 1.835 39.345 2.2 ;
      RECT 39.33 1.835 39.335 2.213 ;
      RECT 39.325 1.835 39.33 2.228 ;
      RECT 39.315 1.835 39.325 2.243 ;
      RECT 39.31 1.835 39.315 2.263 ;
      RECT 39.285 1.835 39.31 2.298 ;
      RECT 39.24 1.835 39.285 2.343 ;
      RECT 39.23 1.835 39.24 2.356 ;
      RECT 39.145 1.92 39.23 2.363 ;
      RECT 39.11 2.042 39.145 2.372 ;
      RECT 39.105 2.082 39.11 2.376 ;
      RECT 39.085 2.105 39.105 2.378 ;
      RECT 39.08 2.135 39.085 2.381 ;
      RECT 39.07 2.147 39.08 2.382 ;
      RECT 39.025 2.17 39.07 2.387 ;
      RECT 38.985 2.2 39.025 2.395 ;
      RECT 38.95 2.212 38.985 2.401 ;
      RECT 38.945 2.217 38.95 2.405 ;
      RECT 38.875 2.227 38.945 2.412 ;
      RECT 38.835 2.237 38.875 2.422 ;
      RECT 38.815 2.242 38.835 2.428 ;
      RECT 38.805 2.246 38.815 2.433 ;
      RECT 38.8 2.249 38.805 2.436 ;
      RECT 38.79 2.25 38.8 2.437 ;
      RECT 38.765 2.252 38.79 2.441 ;
      RECT 38.755 2.257 38.765 2.444 ;
      RECT 38.71 2.265 38.755 2.445 ;
      RECT 38.585 2.27 38.71 2.445 ;
      RECT 39.14 2.567 39.16 2.749 ;
      RECT 39.091 2.552 39.14 2.748 ;
      RECT 39.005 2.567 39.16 2.746 ;
      RECT 38.99 2.567 39.16 2.745 ;
      RECT 38.955 2.545 39.125 2.73 ;
      RECT 39.025 3.565 39.04 3.774 ;
      RECT 39.025 3.573 39.045 3.773 ;
      RECT 38.97 3.573 39.045 3.772 ;
      RECT 38.95 3.577 39.05 3.77 ;
      RECT 38.93 3.527 38.97 3.769 ;
      RECT 38.875 3.585 39.055 3.767 ;
      RECT 38.84 3.542 38.97 3.765 ;
      RECT 38.836 3.545 39.025 3.764 ;
      RECT 38.75 3.553 39.025 3.762 ;
      RECT 38.75 3.597 39.06 3.755 ;
      RECT 38.74 3.69 39.06 3.753 ;
      RECT 38.75 3.609 39.065 3.738 ;
      RECT 38.75 3.63 39.08 3.708 ;
      RECT 38.75 3.657 39.085 3.678 ;
      RECT 38.875 3.535 38.97 3.767 ;
      RECT 38.505 2.58 38.51 3.118 ;
      RECT 38.31 2.91 38.315 3.105 ;
      RECT 36.61 2.575 36.625 2.955 ;
      RECT 38.675 2.575 38.68 2.745 ;
      RECT 38.67 2.575 38.675 2.755 ;
      RECT 38.665 2.575 38.67 2.768 ;
      RECT 38.64 2.575 38.665 2.81 ;
      RECT 38.615 2.575 38.64 2.883 ;
      RECT 38.6 2.575 38.615 2.935 ;
      RECT 38.595 2.575 38.6 2.965 ;
      RECT 38.57 2.575 38.595 3.005 ;
      RECT 38.555 2.575 38.57 3.06 ;
      RECT 38.55 2.575 38.555 3.093 ;
      RECT 38.525 2.575 38.55 3.113 ;
      RECT 38.51 2.575 38.525 3.119 ;
      RECT 38.44 2.61 38.505 3.115 ;
      RECT 38.39 2.665 38.44 3.11 ;
      RECT 38.38 2.697 38.39 3.108 ;
      RECT 38.375 2.722 38.38 3.108 ;
      RECT 38.355 2.795 38.375 3.108 ;
      RECT 38.345 2.875 38.355 3.107 ;
      RECT 38.33 2.905 38.345 3.107 ;
      RECT 38.315 2.91 38.33 3.106 ;
      RECT 38.255 2.912 38.31 3.103 ;
      RECT 38.225 2.917 38.255 3.099 ;
      RECT 38.223 2.92 38.225 3.098 ;
      RECT 38.137 2.922 38.223 3.095 ;
      RECT 38.051 2.928 38.137 3.089 ;
      RECT 37.965 2.933 38.051 3.083 ;
      RECT 37.892 2.938 37.965 3.084 ;
      RECT 37.806 2.944 37.892 3.092 ;
      RECT 37.72 2.95 37.806 3.101 ;
      RECT 37.7 2.954 37.72 3.106 ;
      RECT 37.653 2.956 37.7 3.109 ;
      RECT 37.567 2.961 37.653 3.115 ;
      RECT 37.481 2.966 37.567 3.124 ;
      RECT 37.395 2.972 37.481 3.132 ;
      RECT 37.31 2.97 37.395 3.141 ;
      RECT 37.306 2.965 37.31 3.145 ;
      RECT 37.22 2.96 37.306 3.137 ;
      RECT 37.156 2.951 37.22 3.125 ;
      RECT 37.07 2.942 37.156 3.112 ;
      RECT 37.046 2.935 37.07 3.103 ;
      RECT 36.96 2.929 37.046 3.09 ;
      RECT 36.92 2.922 36.96 3.076 ;
      RECT 36.915 2.912 36.92 3.072 ;
      RECT 36.905 2.9 36.915 3.071 ;
      RECT 36.885 2.87 36.905 3.068 ;
      RECT 36.83 2.79 36.885 3.062 ;
      RECT 36.81 2.709 36.83 3.057 ;
      RECT 36.79 2.667 36.81 3.053 ;
      RECT 36.765 2.62 36.79 3.047 ;
      RECT 36.76 2.595 36.765 3.044 ;
      RECT 36.725 2.575 36.76 3.039 ;
      RECT 36.716 2.575 36.725 3.032 ;
      RECT 36.63 2.575 36.716 3.002 ;
      RECT 36.625 2.575 36.63 2.965 ;
      RECT 36.59 2.575 36.61 2.887 ;
      RECT 36.585 2.617 36.59 2.852 ;
      RECT 36.58 2.692 36.585 2.808 ;
      RECT 38.03 2.497 38.205 2.745 ;
      RECT 38.03 2.497 38.21 2.743 ;
      RECT 38.025 2.529 38.21 2.703 ;
      RECT 38.055 2.47 38.225 2.69 ;
      RECT 38.02 2.547 38.225 2.623 ;
      RECT 37.33 2.01 37.5 2.185 ;
      RECT 37.33 2.01 37.672 2.177 ;
      RECT 37.33 2.01 37.755 2.171 ;
      RECT 37.33 2.01 37.79 2.167 ;
      RECT 37.33 2.01 37.81 2.166 ;
      RECT 37.33 2.01 37.896 2.162 ;
      RECT 37.79 1.835 37.96 2.157 ;
      RECT 37.365 1.942 37.99 2.155 ;
      RECT 37.355 1.997 37.995 2.153 ;
      RECT 37.33 2.033 38.005 2.148 ;
      RECT 37.33 2.06 38.01 2.078 ;
      RECT 37.395 1.885 37.97 2.155 ;
      RECT 37.586 1.87 37.97 2.155 ;
      RECT 37.42 1.873 37.97 2.155 ;
      RECT 37.5 1.871 37.586 2.182 ;
      RECT 37.586 1.868 37.965 2.155 ;
      RECT 37.77 1.845 37.965 2.155 ;
      RECT 37.672 1.866 37.965 2.155 ;
      RECT 37.755 1.86 37.77 2.168 ;
      RECT 37.905 3.225 37.91 3.425 ;
      RECT 37.37 3.29 37.415 3.425 ;
      RECT 37.94 3.225 37.96 3.398 ;
      RECT 37.91 3.225 37.94 3.413 ;
      RECT 37.845 3.225 37.905 3.45 ;
      RECT 37.83 3.225 37.845 3.48 ;
      RECT 37.815 3.225 37.83 3.493 ;
      RECT 37.795 3.225 37.815 3.508 ;
      RECT 37.79 3.225 37.795 3.517 ;
      RECT 37.78 3.229 37.79 3.522 ;
      RECT 37.765 3.239 37.78 3.533 ;
      RECT 37.74 3.255 37.765 3.543 ;
      RECT 37.73 3.269 37.74 3.545 ;
      RECT 37.71 3.281 37.73 3.542 ;
      RECT 37.68 3.302 37.71 3.536 ;
      RECT 37.67 3.314 37.68 3.531 ;
      RECT 37.66 3.312 37.67 3.528 ;
      RECT 37.645 3.311 37.66 3.523 ;
      RECT 37.64 3.31 37.645 3.518 ;
      RECT 37.605 3.308 37.64 3.508 ;
      RECT 37.585 3.305 37.605 3.49 ;
      RECT 37.575 3.303 37.585 3.485 ;
      RECT 37.565 3.302 37.575 3.48 ;
      RECT 37.53 3.3 37.565 3.468 ;
      RECT 37.475 3.296 37.53 3.448 ;
      RECT 37.465 3.294 37.475 3.433 ;
      RECT 37.46 3.294 37.465 3.428 ;
      RECT 37.415 3.292 37.46 3.425 ;
      RECT 37.32 3.29 37.37 3.429 ;
      RECT 37.31 3.291 37.32 3.434 ;
      RECT 37.25 3.298 37.31 3.448 ;
      RECT 37.225 3.306 37.25 3.468 ;
      RECT 37.215 3.31 37.225 3.48 ;
      RECT 37.21 3.311 37.215 3.485 ;
      RECT 37.195 3.313 37.21 3.488 ;
      RECT 37.18 3.315 37.195 3.493 ;
      RECT 37.175 3.315 37.18 3.496 ;
      RECT 37.13 3.32 37.175 3.507 ;
      RECT 37.125 3.324 37.13 3.519 ;
      RECT 37.1 3.32 37.125 3.523 ;
      RECT 37.09 3.316 37.1 3.527 ;
      RECT 37.08 3.315 37.09 3.531 ;
      RECT 37.065 3.305 37.08 3.537 ;
      RECT 37.06 3.293 37.065 3.541 ;
      RECT 37.055 3.29 37.06 3.542 ;
      RECT 37.05 3.287 37.055 3.544 ;
      RECT 37.035 3.275 37.05 3.543 ;
      RECT 37.02 3.257 37.035 3.54 ;
      RECT 37 3.236 37.02 3.533 ;
      RECT 36.935 3.225 37 3.505 ;
      RECT 36.931 3.225 36.935 3.484 ;
      RECT 36.845 3.225 36.931 3.454 ;
      RECT 36.83 3.225 36.845 3.41 ;
      RECT 37.405 2.325 37.41 2.56 ;
      RECT 36.535 2.241 36.54 2.445 ;
      RECT 37.115 2.27 37.12 2.425 ;
      RECT 37.035 2.25 37.04 2.425 ;
      RECT 37.705 2.392 37.72 2.745 ;
      RECT 37.631 2.377 37.705 2.745 ;
      RECT 37.545 2.36 37.631 2.745 ;
      RECT 37.535 2.35 37.545 2.743 ;
      RECT 37.53 2.348 37.535 2.738 ;
      RECT 37.515 2.346 37.53 2.724 ;
      RECT 37.445 2.338 37.515 2.664 ;
      RECT 37.425 2.329 37.445 2.598 ;
      RECT 37.42 2.326 37.425 2.578 ;
      RECT 37.41 2.325 37.42 2.568 ;
      RECT 37.4 2.325 37.405 2.552 ;
      RECT 37.39 2.324 37.4 2.542 ;
      RECT 37.38 2.322 37.39 2.53 ;
      RECT 37.365 2.319 37.38 2.51 ;
      RECT 37.355 2.317 37.365 2.495 ;
      RECT 37.335 2.314 37.355 2.483 ;
      RECT 37.33 2.312 37.335 2.473 ;
      RECT 37.305 2.31 37.33 2.46 ;
      RECT 37.275 2.305 37.305 2.445 ;
      RECT 37.195 2.296 37.275 2.436 ;
      RECT 37.15 2.285 37.195 2.429 ;
      RECT 37.13 2.276 37.15 2.426 ;
      RECT 37.12 2.271 37.13 2.425 ;
      RECT 37.075 2.265 37.115 2.425 ;
      RECT 37.06 2.257 37.075 2.425 ;
      RECT 37.04 2.252 37.06 2.425 ;
      RECT 37.02 2.249 37.035 2.425 ;
      RECT 36.937 2.248 37.02 2.424 ;
      RECT 36.851 2.247 36.937 2.42 ;
      RECT 36.765 2.245 36.851 2.417 ;
      RECT 36.712 2.244 36.765 2.419 ;
      RECT 36.626 2.243 36.712 2.428 ;
      RECT 36.54 2.242 36.626 2.44 ;
      RECT 36.52 2.241 36.535 2.448 ;
      RECT 36.44 2.24 36.52 2.46 ;
      RECT 36.415 2.24 36.44 2.473 ;
      RECT 36.39 2.24 36.415 2.488 ;
      RECT 36.385 2.24 36.39 2.51 ;
      RECT 36.38 2.24 36.385 2.528 ;
      RECT 36.375 2.24 36.38 2.545 ;
      RECT 36.37 2.24 36.375 2.558 ;
      RECT 36.365 2.24 36.37 2.568 ;
      RECT 36.325 2.24 36.365 2.653 ;
      RECT 36.31 2.24 36.325 2.738 ;
      RECT 36.3 2.241 36.31 2.75 ;
      RECT 36.265 2.246 36.3 2.755 ;
      RECT 36.225 2.255 36.265 2.755 ;
      RECT 36.21 2.265 36.225 2.755 ;
      RECT 36.205 2.275 36.21 2.755 ;
      RECT 36.185 2.302 36.205 2.755 ;
      RECT 36.135 2.385 36.185 2.755 ;
      RECT 36.13 2.447 36.135 2.755 ;
      RECT 36.12 2.46 36.13 2.755 ;
      RECT 36.11 2.482 36.12 2.755 ;
      RECT 36.1 2.507 36.11 2.75 ;
      RECT 36.095 2.545 36.1 2.743 ;
      RECT 36.085 2.655 36.095 2.738 ;
      RECT 37.48 3.576 37.495 3.835 ;
      RECT 37.48 3.591 37.5 3.834 ;
      RECT 37.396 3.591 37.5 3.832 ;
      RECT 37.396 3.605 37.505 3.831 ;
      RECT 37.31 3.647 37.51 3.828 ;
      RECT 37.305 3.59 37.495 3.823 ;
      RECT 37.305 3.661 37.515 3.82 ;
      RECT 37.3 3.692 37.515 3.818 ;
      RECT 37.305 3.689 37.53 3.808 ;
      RECT 37.3 3.735 37.545 3.793 ;
      RECT 37.3 3.763 37.55 3.778 ;
      RECT 37.31 3.565 37.48 3.828 ;
      RECT 37.07 2.575 37.24 2.745 ;
      RECT 37.035 2.575 37.24 2.74 ;
      RECT 37.025 2.575 37.24 2.733 ;
      RECT 37.02 2.56 37.19 2.73 ;
      RECT 35.85 3.097 36.115 3.54 ;
      RECT 35.845 3.068 36.06 3.538 ;
      RECT 35.84 3.222 36.12 3.533 ;
      RECT 35.845 3.117 36.12 3.533 ;
      RECT 35.845 3.128 36.13 3.52 ;
      RECT 35.845 3.075 36.09 3.538 ;
      RECT 35.85 3.062 36.06 3.54 ;
      RECT 35.85 3.06 36.01 3.54 ;
      RECT 35.951 3.052 36.01 3.54 ;
      RECT 35.865 3.053 36.01 3.54 ;
      RECT 35.951 3.051 36 3.54 ;
      RECT 35.755 1.866 35.93 2.165 ;
      RECT 35.805 1.828 35.93 2.165 ;
      RECT 35.79 1.83 36.016 2.157 ;
      RECT 35.79 1.833 36.055 2.144 ;
      RECT 35.79 1.834 36.065 2.13 ;
      RECT 35.745 1.885 36.065 2.12 ;
      RECT 35.79 1.835 36.07 2.115 ;
      RECT 35.745 2.045 36.075 2.105 ;
      RECT 35.73 1.905 36.07 2.045 ;
      RECT 35.725 1.921 36.07 1.985 ;
      RECT 35.77 1.845 36.07 2.115 ;
      RECT 35.805 1.826 35.891 2.165 ;
      RECT 34.265 5.02 34.435 6.49 ;
      RECT 34.265 6.315 34.44 6.485 ;
      RECT 33.895 1.74 34.065 2.93 ;
      RECT 33.895 1.74 34.365 1.91 ;
      RECT 33.895 6.97 34.365 7.14 ;
      RECT 33.895 5.95 34.065 7.14 ;
      RECT 32.905 1.74 33.075 2.93 ;
      RECT 32.905 1.74 33.375 1.91 ;
      RECT 32.905 6.97 33.375 7.14 ;
      RECT 32.905 5.95 33.075 7.14 ;
      RECT 31.055 2.635 31.225 3.865 ;
      RECT 31.11 0.855 31.28 2.805 ;
      RECT 31.055 0.575 31.225 1.025 ;
      RECT 31.055 7.855 31.225 8.305 ;
      RECT 31.11 6.075 31.28 8.025 ;
      RECT 31.055 5.015 31.225 6.245 ;
      RECT 30.535 0.575 30.705 3.865 ;
      RECT 30.535 2.075 30.94 2.405 ;
      RECT 30.535 1.235 30.94 1.565 ;
      RECT 30.535 5.015 30.705 8.305 ;
      RECT 30.535 7.315 30.94 7.645 ;
      RECT 30.535 6.475 30.94 6.805 ;
      RECT 28.46 3.126 28.465 3.298 ;
      RECT 28.455 3.119 28.46 3.388 ;
      RECT 28.45 3.113 28.455 3.407 ;
      RECT 28.43 3.107 28.45 3.417 ;
      RECT 28.415 3.102 28.43 3.425 ;
      RECT 28.378 3.096 28.415 3.423 ;
      RECT 28.292 3.082 28.378 3.419 ;
      RECT 28.206 3.064 28.292 3.414 ;
      RECT 28.12 3.045 28.206 3.408 ;
      RECT 28.09 3.033 28.12 3.404 ;
      RECT 28.07 3.027 28.09 3.403 ;
      RECT 28.005 3.025 28.07 3.401 ;
      RECT 27.99 3.025 28.005 3.393 ;
      RECT 27.975 3.025 27.99 3.38 ;
      RECT 27.97 3.025 27.975 3.37 ;
      RECT 27.955 3.025 27.97 3.348 ;
      RECT 27.94 3.025 27.955 3.315 ;
      RECT 27.935 3.025 27.94 3.293 ;
      RECT 27.925 3.025 27.935 3.275 ;
      RECT 27.91 3.025 27.925 3.253 ;
      RECT 27.89 3.025 27.91 3.215 ;
      RECT 28.24 2.31 28.275 2.749 ;
      RECT 28.24 2.31 28.28 2.748 ;
      RECT 28.185 2.37 28.28 2.747 ;
      RECT 28.05 2.542 28.28 2.746 ;
      RECT 28.16 2.42 28.28 2.746 ;
      RECT 28.05 2.542 28.305 2.736 ;
      RECT 28.105 2.487 28.385 2.653 ;
      RECT 28.28 2.281 28.285 2.744 ;
      RECT 28.135 2.457 28.425 2.53 ;
      RECT 28.15 2.44 28.28 2.746 ;
      RECT 28.285 2.28 28.455 2.468 ;
      RECT 28.275 2.283 28.455 2.468 ;
      RECT 27.78 2.16 27.95 2.47 ;
      RECT 27.78 2.16 27.955 2.443 ;
      RECT 27.78 2.16 27.96 2.42 ;
      RECT 27.78 2.16 27.97 2.37 ;
      RECT 27.775 2.265 27.97 2.34 ;
      RECT 27.81 1.835 27.98 2.313 ;
      RECT 27.81 1.835 27.995 2.234 ;
      RECT 27.8 2.045 27.995 2.234 ;
      RECT 27.81 1.845 28.005 2.149 ;
      RECT 27.74 2.587 27.745 2.79 ;
      RECT 27.73 2.575 27.74 2.9 ;
      RECT 27.705 2.575 27.73 2.94 ;
      RECT 27.625 2.575 27.705 3.025 ;
      RECT 27.615 2.575 27.625 3.095 ;
      RECT 27.59 2.575 27.615 3.118 ;
      RECT 27.57 2.575 27.59 3.153 ;
      RECT 27.525 2.585 27.57 3.196 ;
      RECT 27.515 2.597 27.525 3.233 ;
      RECT 27.495 2.611 27.515 3.253 ;
      RECT 27.485 2.629 27.495 3.269 ;
      RECT 27.47 2.655 27.485 3.279 ;
      RECT 27.455 2.696 27.47 3.293 ;
      RECT 27.445 2.731 27.455 3.303 ;
      RECT 27.44 2.747 27.445 3.308 ;
      RECT 27.43 2.762 27.44 3.313 ;
      RECT 27.41 2.805 27.43 3.323 ;
      RECT 27.39 2.842 27.41 3.336 ;
      RECT 27.355 2.865 27.39 3.354 ;
      RECT 27.345 2.879 27.355 3.37 ;
      RECT 27.325 2.889 27.345 3.38 ;
      RECT 27.32 2.898 27.325 3.388 ;
      RECT 27.31 2.905 27.32 3.395 ;
      RECT 27.3 2.912 27.31 3.403 ;
      RECT 27.285 2.922 27.3 3.411 ;
      RECT 27.275 2.936 27.285 3.421 ;
      RECT 27.265 2.948 27.275 3.433 ;
      RECT 27.25 2.97 27.265 3.446 ;
      RECT 27.24 2.992 27.25 3.457 ;
      RECT 27.23 3.012 27.24 3.466 ;
      RECT 27.225 3.027 27.23 3.473 ;
      RECT 27.195 3.06 27.225 3.487 ;
      RECT 27.185 3.095 27.195 3.502 ;
      RECT 27.18 3.102 27.185 3.508 ;
      RECT 27.16 3.117 27.18 3.515 ;
      RECT 27.155 3.132 27.16 3.523 ;
      RECT 27.15 3.141 27.155 3.528 ;
      RECT 27.135 3.147 27.15 3.535 ;
      RECT 27.13 3.153 27.135 3.543 ;
      RECT 27.125 3.157 27.13 3.55 ;
      RECT 27.12 3.161 27.125 3.56 ;
      RECT 27.11 3.166 27.12 3.57 ;
      RECT 27.09 3.177 27.11 3.598 ;
      RECT 27.075 3.189 27.09 3.625 ;
      RECT 27.055 3.202 27.075 3.65 ;
      RECT 27.035 3.217 27.055 3.674 ;
      RECT 27.02 3.232 27.035 3.689 ;
      RECT 27.015 3.243 27.02 3.698 ;
      RECT 26.95 3.288 27.015 3.708 ;
      RECT 26.915 3.347 26.95 3.721 ;
      RECT 26.91 3.37 26.915 3.727 ;
      RECT 26.905 3.377 26.91 3.729 ;
      RECT 26.89 3.387 26.905 3.732 ;
      RECT 26.86 3.412 26.89 3.736 ;
      RECT 26.855 3.43 26.86 3.74 ;
      RECT 26.85 3.437 26.855 3.741 ;
      RECT 26.83 3.445 26.85 3.745 ;
      RECT 26.82 3.452 26.83 3.749 ;
      RECT 26.776 3.463 26.82 3.756 ;
      RECT 26.69 3.491 26.776 3.772 ;
      RECT 26.63 3.515 26.69 3.79 ;
      RECT 26.585 3.525 26.63 3.804 ;
      RECT 26.526 3.533 26.585 3.818 ;
      RECT 26.44 3.54 26.526 3.837 ;
      RECT 26.415 3.545 26.44 3.852 ;
      RECT 26.335 3.548 26.415 3.855 ;
      RECT 26.255 3.552 26.335 3.842 ;
      RECT 26.246 3.555 26.255 3.827 ;
      RECT 26.16 3.555 26.246 3.812 ;
      RECT 26.1 3.557 26.16 3.789 ;
      RECT 26.096 3.56 26.1 3.779 ;
      RECT 26.01 3.56 26.096 3.764 ;
      RECT 25.935 3.56 26.01 3.74 ;
      RECT 27.25 2.569 27.26 2.745 ;
      RECT 27.205 2.536 27.25 2.745 ;
      RECT 27.16 2.487 27.205 2.745 ;
      RECT 27.13 2.457 27.16 2.746 ;
      RECT 27.125 2.44 27.13 2.747 ;
      RECT 27.1 2.42 27.125 2.748 ;
      RECT 27.085 2.395 27.1 2.749 ;
      RECT 27.08 2.382 27.085 2.75 ;
      RECT 27.075 2.376 27.08 2.748 ;
      RECT 27.07 2.368 27.075 2.742 ;
      RECT 27.045 2.36 27.07 2.722 ;
      RECT 27.025 2.349 27.045 2.693 ;
      RECT 26.995 2.334 27.025 2.664 ;
      RECT 26.975 2.32 26.995 2.636 ;
      RECT 26.965 2.314 26.975 2.615 ;
      RECT 26.96 2.311 26.965 2.598 ;
      RECT 26.955 2.308 26.96 2.583 ;
      RECT 26.94 2.303 26.955 2.548 ;
      RECT 26.935 2.299 26.94 2.515 ;
      RECT 26.915 2.294 26.935 2.491 ;
      RECT 26.885 2.286 26.915 2.456 ;
      RECT 26.87 2.28 26.885 2.433 ;
      RECT 26.83 2.273 26.87 2.418 ;
      RECT 26.805 2.265 26.83 2.398 ;
      RECT 26.785 2.26 26.805 2.388 ;
      RECT 26.75 2.254 26.785 2.383 ;
      RECT 26.705 2.245 26.75 2.382 ;
      RECT 26.675 2.241 26.705 2.384 ;
      RECT 26.59 2.249 26.675 2.388 ;
      RECT 26.52 2.26 26.59 2.41 ;
      RECT 26.507 2.266 26.52 2.433 ;
      RECT 26.421 2.273 26.507 2.455 ;
      RECT 26.335 2.285 26.421 2.492 ;
      RECT 26.335 2.662 26.345 2.9 ;
      RECT 26.33 2.291 26.335 2.515 ;
      RECT 26.325 2.547 26.335 2.9 ;
      RECT 26.325 2.292 26.33 2.52 ;
      RECT 26.32 2.293 26.325 2.9 ;
      RECT 26.296 2.295 26.32 2.901 ;
      RECT 26.21 2.303 26.296 2.903 ;
      RECT 26.19 2.317 26.21 2.906 ;
      RECT 26.185 2.345 26.19 2.907 ;
      RECT 26.18 2.357 26.185 2.908 ;
      RECT 26.175 2.372 26.18 2.909 ;
      RECT 26.165 2.402 26.175 2.91 ;
      RECT 26.16 2.44 26.165 2.908 ;
      RECT 26.155 2.46 26.16 2.903 ;
      RECT 26.14 2.495 26.155 2.888 ;
      RECT 26.13 2.547 26.14 2.868 ;
      RECT 26.125 2.577 26.13 2.856 ;
      RECT 26.11 2.59 26.125 2.839 ;
      RECT 26.085 2.594 26.11 2.806 ;
      RECT 26.07 2.592 26.085 2.783 ;
      RECT 26.055 2.591 26.07 2.78 ;
      RECT 25.995 2.589 26.055 2.778 ;
      RECT 25.985 2.587 25.995 2.773 ;
      RECT 25.945 2.586 25.985 2.77 ;
      RECT 25.875 2.583 25.945 2.768 ;
      RECT 25.82 2.581 25.875 2.763 ;
      RECT 25.75 2.575 25.82 2.758 ;
      RECT 25.741 2.575 25.75 2.755 ;
      RECT 25.655 2.575 25.741 2.75 ;
      RECT 25.65 2.575 25.655 2.745 ;
      RECT 26.955 1.81 27.13 2.16 ;
      RECT 26.955 1.825 27.14 2.158 ;
      RECT 26.93 1.775 27.075 2.155 ;
      RECT 26.91 1.776 27.075 2.148 ;
      RECT 26.9 1.777 27.085 2.143 ;
      RECT 26.87 1.778 27.085 2.13 ;
      RECT 26.82 1.779 27.085 2.106 ;
      RECT 26.815 1.781 27.085 2.091 ;
      RECT 26.815 1.847 27.145 2.085 ;
      RECT 26.795 1.788 27.1 2.065 ;
      RECT 26.785 1.797 27.11 1.92 ;
      RECT 26.795 1.792 27.11 2.065 ;
      RECT 26.815 1.782 27.1 2.091 ;
      RECT 26.4 3.107 26.57 3.395 ;
      RECT 26.395 3.125 26.58 3.39 ;
      RECT 26.36 3.133 26.645 3.31 ;
      RECT 26.36 3.133 26.731 3.3 ;
      RECT 26.36 3.133 26.785 3.246 ;
      RECT 26.645 3.03 26.815 3.214 ;
      RECT 26.36 3.185 26.82 3.202 ;
      RECT 26.345 3.155 26.815 3.198 ;
      RECT 26.605 3.037 26.645 3.349 ;
      RECT 26.485 3.074 26.815 3.214 ;
      RECT 26.58 3.049 26.605 3.375 ;
      RECT 26.57 3.056 26.815 3.214 ;
      RECT 26.701 2.52 26.77 2.779 ;
      RECT 26.701 2.575 26.775 2.778 ;
      RECT 26.615 2.575 26.775 2.777 ;
      RECT 26.61 2.575 26.78 2.77 ;
      RECT 26.6 2.52 26.77 2.765 ;
      RECT 25.98 1.819 26.155 2.12 ;
      RECT 25.965 1.807 25.98 2.105 ;
      RECT 25.935 1.806 25.965 2.058 ;
      RECT 25.935 1.824 26.16 2.053 ;
      RECT 25.92 1.808 25.98 2.018 ;
      RECT 25.915 1.83 26.17 1.918 ;
      RECT 25.915 1.813 26.066 1.918 ;
      RECT 25.915 1.815 26.07 1.918 ;
      RECT 25.92 1.811 26.066 2.018 ;
      RECT 26.025 3.047 26.03 3.395 ;
      RECT 26.015 3.037 26.025 3.401 ;
      RECT 25.98 3.027 26.015 3.403 ;
      RECT 25.942 3.022 25.98 3.407 ;
      RECT 25.856 3.015 25.942 3.414 ;
      RECT 25.77 3.005 25.856 3.424 ;
      RECT 25.725 3 25.77 3.432 ;
      RECT 25.721 3 25.725 3.436 ;
      RECT 25.635 3 25.721 3.443 ;
      RECT 25.62 3 25.635 3.443 ;
      RECT 25.61 2.998 25.62 3.415 ;
      RECT 25.6 2.994 25.61 3.358 ;
      RECT 25.58 2.988 25.6 3.29 ;
      RECT 25.575 2.984 25.58 3.238 ;
      RECT 25.565 2.983 25.575 3.205 ;
      RECT 25.515 2.981 25.565 3.19 ;
      RECT 25.49 2.979 25.515 3.185 ;
      RECT 25.447 2.977 25.49 3.181 ;
      RECT 25.361 2.973 25.447 3.169 ;
      RECT 25.275 2.968 25.361 3.153 ;
      RECT 25.245 2.965 25.275 3.14 ;
      RECT 25.22 2.964 25.245 3.128 ;
      RECT 25.215 2.964 25.22 3.118 ;
      RECT 25.175 2.963 25.215 3.11 ;
      RECT 25.16 2.962 25.175 3.103 ;
      RECT 25.11 2.961 25.16 3.095 ;
      RECT 25.108 2.96 25.11 3.09 ;
      RECT 25.022 2.958 25.108 3.09 ;
      RECT 24.936 2.953 25.022 3.09 ;
      RECT 24.85 2.949 24.936 3.09 ;
      RECT 24.801 2.945 24.85 3.088 ;
      RECT 24.715 2.942 24.801 3.083 ;
      RECT 24.692 2.939 24.715 3.079 ;
      RECT 24.606 2.936 24.692 3.074 ;
      RECT 24.52 2.932 24.606 3.065 ;
      RECT 24.495 2.925 24.52 3.06 ;
      RECT 24.435 2.89 24.495 3.057 ;
      RECT 24.415 2.815 24.435 3.054 ;
      RECT 24.41 2.757 24.415 3.053 ;
      RECT 24.385 2.697 24.41 3.052 ;
      RECT 24.31 2.575 24.385 3.048 ;
      RECT 24.3 2.575 24.31 3.04 ;
      RECT 24.285 2.575 24.3 3.03 ;
      RECT 24.27 2.575 24.285 3 ;
      RECT 24.255 2.575 24.27 2.945 ;
      RECT 24.24 2.575 24.255 2.883 ;
      RECT 24.215 2.575 24.24 2.808 ;
      RECT 24.21 2.575 24.215 2.758 ;
      RECT 25.555 2.12 25.575 2.429 ;
      RECT 25.541 2.122 25.59 2.426 ;
      RECT 25.541 2.127 25.61 2.417 ;
      RECT 25.455 2.125 25.59 2.411 ;
      RECT 25.455 2.133 25.645 2.394 ;
      RECT 25.42 2.135 25.645 2.393 ;
      RECT 25.39 2.143 25.645 2.384 ;
      RECT 25.38 2.148 25.665 2.37 ;
      RECT 25.42 2.138 25.665 2.37 ;
      RECT 25.42 2.141 25.675 2.358 ;
      RECT 25.39 2.143 25.685 2.345 ;
      RECT 25.39 2.147 25.695 2.288 ;
      RECT 25.38 2.152 25.7 2.203 ;
      RECT 25.541 2.12 25.575 2.426 ;
      RECT 25.42 7.855 25.59 8.305 ;
      RECT 25.475 6.075 25.645 8.025 ;
      RECT 25.42 5.015 25.59 6.245 ;
      RECT 24.98 2.223 24.985 2.435 ;
      RECT 24.855 2.22 24.87 2.435 ;
      RECT 24.32 2.25 24.39 2.435 ;
      RECT 24.205 2.25 24.24 2.43 ;
      RECT 25.326 2.552 25.345 2.746 ;
      RECT 25.24 2.507 25.326 2.747 ;
      RECT 25.23 2.46 25.24 2.749 ;
      RECT 25.225 2.44 25.23 2.75 ;
      RECT 25.205 2.405 25.225 2.751 ;
      RECT 25.19 2.355 25.205 2.752 ;
      RECT 25.17 2.292 25.19 2.753 ;
      RECT 25.16 2.255 25.17 2.754 ;
      RECT 25.145 2.244 25.16 2.755 ;
      RECT 25.14 2.236 25.145 2.753 ;
      RECT 25.13 2.235 25.14 2.745 ;
      RECT 25.1 2.232 25.13 2.724 ;
      RECT 25.025 2.227 25.1 2.669 ;
      RECT 25.01 2.223 25.025 2.615 ;
      RECT 25 2.223 25.01 2.51 ;
      RECT 24.985 2.223 25 2.443 ;
      RECT 24.97 2.223 24.98 2.433 ;
      RECT 24.915 2.222 24.97 2.43 ;
      RECT 24.87 2.22 24.915 2.433 ;
      RECT 24.842 2.22 24.855 2.436 ;
      RECT 24.756 2.224 24.842 2.438 ;
      RECT 24.67 2.23 24.756 2.443 ;
      RECT 24.65 2.234 24.67 2.445 ;
      RECT 24.648 2.235 24.65 2.444 ;
      RECT 24.562 2.237 24.648 2.443 ;
      RECT 24.476 2.242 24.562 2.44 ;
      RECT 24.39 2.247 24.476 2.437 ;
      RECT 24.24 2.25 24.32 2.433 ;
      RECT 24.9 5.015 25.07 8.305 ;
      RECT 24.9 7.315 25.305 7.645 ;
      RECT 24.9 6.475 25.305 6.805 ;
      RECT 25.016 3.225 25.065 3.559 ;
      RECT 25.016 3.225 25.07 3.558 ;
      RECT 24.93 3.225 25.07 3.557 ;
      RECT 24.705 3.333 25.075 3.555 ;
      RECT 24.93 3.225 25.1 3.548 ;
      RECT 24.9 3.237 25.105 3.539 ;
      RECT 24.885 3.255 25.11 3.536 ;
      RECT 24.7 3.339 25.11 3.463 ;
      RECT 24.695 3.346 25.11 3.423 ;
      RECT 24.71 3.312 25.11 3.536 ;
      RECT 24.871 3.258 25.075 3.555 ;
      RECT 24.785 3.278 25.11 3.536 ;
      RECT 24.885 3.252 25.105 3.539 ;
      RECT 24.655 2.576 24.845 2.77 ;
      RECT 24.65 2.578 24.845 2.769 ;
      RECT 24.645 2.582 24.86 2.766 ;
      RECT 24.66 2.575 24.86 2.766 ;
      RECT 24.645 2.685 24.865 2.761 ;
      RECT 23.94 3.185 24.031 3.483 ;
      RECT 23.935 3.187 24.11 3.478 ;
      RECT 23.94 3.185 24.11 3.478 ;
      RECT 23.935 3.191 24.13 3.476 ;
      RECT 23.935 3.246 24.17 3.475 ;
      RECT 23.935 3.281 24.185 3.469 ;
      RECT 23.935 3.315 24.195 3.459 ;
      RECT 23.925 3.195 24.13 3.31 ;
      RECT 23.925 3.215 24.145 3.31 ;
      RECT 23.925 3.198 24.135 3.31 ;
      RECT 24.15 1.966 24.155 2.028 ;
      RECT 24.145 1.888 24.15 2.051 ;
      RECT 24.14 1.845 24.145 2.062 ;
      RECT 24.135 1.835 24.14 2.074 ;
      RECT 24.13 1.835 24.135 2.083 ;
      RECT 24.105 1.835 24.13 2.115 ;
      RECT 24.1 1.835 24.105 2.148 ;
      RECT 24.085 1.835 24.1 2.173 ;
      RECT 24.075 1.835 24.085 2.2 ;
      RECT 24.07 1.835 24.075 2.213 ;
      RECT 24.065 1.835 24.07 2.228 ;
      RECT 24.055 1.835 24.065 2.243 ;
      RECT 24.05 1.835 24.055 2.263 ;
      RECT 24.025 1.835 24.05 2.298 ;
      RECT 23.98 1.835 24.025 2.343 ;
      RECT 23.97 1.835 23.98 2.356 ;
      RECT 23.885 1.92 23.97 2.363 ;
      RECT 23.85 2.042 23.885 2.372 ;
      RECT 23.845 2.082 23.85 2.376 ;
      RECT 23.825 2.105 23.845 2.378 ;
      RECT 23.82 2.135 23.825 2.381 ;
      RECT 23.81 2.147 23.82 2.382 ;
      RECT 23.765 2.17 23.81 2.387 ;
      RECT 23.725 2.2 23.765 2.395 ;
      RECT 23.69 2.212 23.725 2.401 ;
      RECT 23.685 2.217 23.69 2.405 ;
      RECT 23.615 2.227 23.685 2.412 ;
      RECT 23.575 2.237 23.615 2.422 ;
      RECT 23.555 2.242 23.575 2.428 ;
      RECT 23.545 2.246 23.555 2.433 ;
      RECT 23.54 2.249 23.545 2.436 ;
      RECT 23.53 2.25 23.54 2.437 ;
      RECT 23.505 2.252 23.53 2.441 ;
      RECT 23.495 2.257 23.505 2.444 ;
      RECT 23.45 2.265 23.495 2.445 ;
      RECT 23.325 2.27 23.45 2.445 ;
      RECT 23.88 2.567 23.9 2.749 ;
      RECT 23.831 2.552 23.88 2.748 ;
      RECT 23.745 2.567 23.9 2.746 ;
      RECT 23.73 2.567 23.9 2.745 ;
      RECT 23.695 2.545 23.865 2.73 ;
      RECT 23.765 3.565 23.78 3.774 ;
      RECT 23.765 3.573 23.785 3.773 ;
      RECT 23.71 3.573 23.785 3.772 ;
      RECT 23.69 3.577 23.79 3.77 ;
      RECT 23.67 3.527 23.71 3.769 ;
      RECT 23.615 3.585 23.795 3.767 ;
      RECT 23.58 3.542 23.71 3.765 ;
      RECT 23.576 3.545 23.765 3.764 ;
      RECT 23.49 3.553 23.765 3.762 ;
      RECT 23.49 3.597 23.8 3.755 ;
      RECT 23.48 3.69 23.8 3.753 ;
      RECT 23.49 3.609 23.805 3.738 ;
      RECT 23.49 3.63 23.82 3.708 ;
      RECT 23.49 3.657 23.825 3.678 ;
      RECT 23.615 3.535 23.71 3.767 ;
      RECT 23.245 2.58 23.25 3.118 ;
      RECT 23.05 2.91 23.055 3.105 ;
      RECT 21.35 2.575 21.365 2.955 ;
      RECT 23.415 2.575 23.42 2.745 ;
      RECT 23.41 2.575 23.415 2.755 ;
      RECT 23.405 2.575 23.41 2.768 ;
      RECT 23.38 2.575 23.405 2.81 ;
      RECT 23.355 2.575 23.38 2.883 ;
      RECT 23.34 2.575 23.355 2.935 ;
      RECT 23.335 2.575 23.34 2.965 ;
      RECT 23.31 2.575 23.335 3.005 ;
      RECT 23.295 2.575 23.31 3.06 ;
      RECT 23.29 2.575 23.295 3.093 ;
      RECT 23.265 2.575 23.29 3.113 ;
      RECT 23.25 2.575 23.265 3.119 ;
      RECT 23.18 2.61 23.245 3.115 ;
      RECT 23.13 2.665 23.18 3.11 ;
      RECT 23.12 2.697 23.13 3.108 ;
      RECT 23.115 2.722 23.12 3.108 ;
      RECT 23.095 2.795 23.115 3.108 ;
      RECT 23.085 2.875 23.095 3.107 ;
      RECT 23.07 2.905 23.085 3.107 ;
      RECT 23.055 2.91 23.07 3.106 ;
      RECT 22.995 2.912 23.05 3.103 ;
      RECT 22.965 2.917 22.995 3.099 ;
      RECT 22.963 2.92 22.965 3.098 ;
      RECT 22.877 2.922 22.963 3.095 ;
      RECT 22.791 2.928 22.877 3.089 ;
      RECT 22.705 2.933 22.791 3.083 ;
      RECT 22.632 2.938 22.705 3.084 ;
      RECT 22.546 2.944 22.632 3.092 ;
      RECT 22.46 2.95 22.546 3.101 ;
      RECT 22.44 2.954 22.46 3.106 ;
      RECT 22.393 2.956 22.44 3.109 ;
      RECT 22.307 2.961 22.393 3.115 ;
      RECT 22.221 2.966 22.307 3.124 ;
      RECT 22.135 2.972 22.221 3.132 ;
      RECT 22.05 2.97 22.135 3.141 ;
      RECT 22.046 2.965 22.05 3.145 ;
      RECT 21.96 2.96 22.046 3.137 ;
      RECT 21.896 2.951 21.96 3.125 ;
      RECT 21.81 2.942 21.896 3.112 ;
      RECT 21.786 2.935 21.81 3.103 ;
      RECT 21.7 2.929 21.786 3.09 ;
      RECT 21.66 2.922 21.7 3.076 ;
      RECT 21.655 2.912 21.66 3.072 ;
      RECT 21.645 2.9 21.655 3.071 ;
      RECT 21.625 2.87 21.645 3.068 ;
      RECT 21.57 2.79 21.625 3.062 ;
      RECT 21.55 2.709 21.57 3.057 ;
      RECT 21.53 2.667 21.55 3.053 ;
      RECT 21.505 2.62 21.53 3.047 ;
      RECT 21.5 2.595 21.505 3.044 ;
      RECT 21.465 2.575 21.5 3.039 ;
      RECT 21.456 2.575 21.465 3.032 ;
      RECT 21.37 2.575 21.456 3.002 ;
      RECT 21.365 2.575 21.37 2.965 ;
      RECT 21.33 2.575 21.35 2.887 ;
      RECT 21.325 2.617 21.33 2.852 ;
      RECT 21.32 2.692 21.325 2.808 ;
      RECT 22.77 2.497 22.945 2.745 ;
      RECT 22.77 2.497 22.95 2.743 ;
      RECT 22.765 2.529 22.95 2.703 ;
      RECT 22.795 2.47 22.965 2.69 ;
      RECT 22.76 2.547 22.965 2.623 ;
      RECT 22.07 2.01 22.24 2.185 ;
      RECT 22.07 2.01 22.412 2.177 ;
      RECT 22.07 2.01 22.495 2.171 ;
      RECT 22.07 2.01 22.53 2.167 ;
      RECT 22.07 2.01 22.55 2.166 ;
      RECT 22.07 2.01 22.636 2.162 ;
      RECT 22.53 1.835 22.7 2.157 ;
      RECT 22.105 1.942 22.73 2.155 ;
      RECT 22.095 1.997 22.735 2.153 ;
      RECT 22.07 2.033 22.745 2.148 ;
      RECT 22.07 2.06 22.75 2.078 ;
      RECT 22.135 1.885 22.71 2.155 ;
      RECT 22.326 1.87 22.71 2.155 ;
      RECT 22.16 1.873 22.71 2.155 ;
      RECT 22.24 1.871 22.326 2.182 ;
      RECT 22.326 1.868 22.705 2.155 ;
      RECT 22.51 1.845 22.705 2.155 ;
      RECT 22.412 1.866 22.705 2.155 ;
      RECT 22.495 1.86 22.51 2.168 ;
      RECT 22.645 3.225 22.65 3.425 ;
      RECT 22.11 3.29 22.155 3.425 ;
      RECT 22.68 3.225 22.7 3.398 ;
      RECT 22.65 3.225 22.68 3.413 ;
      RECT 22.585 3.225 22.645 3.45 ;
      RECT 22.57 3.225 22.585 3.48 ;
      RECT 22.555 3.225 22.57 3.493 ;
      RECT 22.535 3.225 22.555 3.508 ;
      RECT 22.53 3.225 22.535 3.517 ;
      RECT 22.52 3.229 22.53 3.522 ;
      RECT 22.505 3.239 22.52 3.533 ;
      RECT 22.48 3.255 22.505 3.543 ;
      RECT 22.47 3.269 22.48 3.545 ;
      RECT 22.45 3.281 22.47 3.542 ;
      RECT 22.42 3.302 22.45 3.536 ;
      RECT 22.41 3.314 22.42 3.531 ;
      RECT 22.4 3.312 22.41 3.528 ;
      RECT 22.385 3.311 22.4 3.523 ;
      RECT 22.38 3.31 22.385 3.518 ;
      RECT 22.345 3.308 22.38 3.508 ;
      RECT 22.325 3.305 22.345 3.49 ;
      RECT 22.315 3.303 22.325 3.485 ;
      RECT 22.305 3.302 22.315 3.48 ;
      RECT 22.27 3.3 22.305 3.468 ;
      RECT 22.215 3.296 22.27 3.448 ;
      RECT 22.205 3.294 22.215 3.433 ;
      RECT 22.2 3.294 22.205 3.428 ;
      RECT 22.155 3.292 22.2 3.425 ;
      RECT 22.06 3.29 22.11 3.429 ;
      RECT 22.05 3.291 22.06 3.434 ;
      RECT 21.99 3.298 22.05 3.448 ;
      RECT 21.965 3.306 21.99 3.468 ;
      RECT 21.955 3.31 21.965 3.48 ;
      RECT 21.95 3.311 21.955 3.485 ;
      RECT 21.935 3.313 21.95 3.488 ;
      RECT 21.92 3.315 21.935 3.493 ;
      RECT 21.915 3.315 21.92 3.496 ;
      RECT 21.87 3.32 21.915 3.507 ;
      RECT 21.865 3.324 21.87 3.519 ;
      RECT 21.84 3.32 21.865 3.523 ;
      RECT 21.83 3.316 21.84 3.527 ;
      RECT 21.82 3.315 21.83 3.531 ;
      RECT 21.805 3.305 21.82 3.537 ;
      RECT 21.8 3.293 21.805 3.541 ;
      RECT 21.795 3.29 21.8 3.542 ;
      RECT 21.79 3.287 21.795 3.544 ;
      RECT 21.775 3.275 21.79 3.543 ;
      RECT 21.76 3.257 21.775 3.54 ;
      RECT 21.74 3.236 21.76 3.533 ;
      RECT 21.675 3.225 21.74 3.505 ;
      RECT 21.671 3.225 21.675 3.484 ;
      RECT 21.585 3.225 21.671 3.454 ;
      RECT 21.57 3.225 21.585 3.41 ;
      RECT 22.145 2.325 22.15 2.56 ;
      RECT 21.275 2.241 21.28 2.445 ;
      RECT 21.855 2.27 21.86 2.425 ;
      RECT 21.775 2.25 21.78 2.425 ;
      RECT 22.445 2.392 22.46 2.745 ;
      RECT 22.371 2.377 22.445 2.745 ;
      RECT 22.285 2.36 22.371 2.745 ;
      RECT 22.275 2.35 22.285 2.743 ;
      RECT 22.27 2.348 22.275 2.738 ;
      RECT 22.255 2.346 22.27 2.724 ;
      RECT 22.185 2.338 22.255 2.664 ;
      RECT 22.165 2.329 22.185 2.598 ;
      RECT 22.16 2.326 22.165 2.578 ;
      RECT 22.15 2.325 22.16 2.568 ;
      RECT 22.14 2.325 22.145 2.552 ;
      RECT 22.13 2.324 22.14 2.542 ;
      RECT 22.12 2.322 22.13 2.53 ;
      RECT 22.105 2.319 22.12 2.51 ;
      RECT 22.095 2.317 22.105 2.495 ;
      RECT 22.075 2.314 22.095 2.483 ;
      RECT 22.07 2.312 22.075 2.473 ;
      RECT 22.045 2.31 22.07 2.46 ;
      RECT 22.015 2.305 22.045 2.445 ;
      RECT 21.935 2.296 22.015 2.436 ;
      RECT 21.89 2.285 21.935 2.429 ;
      RECT 21.87 2.276 21.89 2.426 ;
      RECT 21.86 2.271 21.87 2.425 ;
      RECT 21.815 2.265 21.855 2.425 ;
      RECT 21.8 2.257 21.815 2.425 ;
      RECT 21.78 2.252 21.8 2.425 ;
      RECT 21.76 2.249 21.775 2.425 ;
      RECT 21.677 2.248 21.76 2.424 ;
      RECT 21.591 2.247 21.677 2.42 ;
      RECT 21.505 2.245 21.591 2.417 ;
      RECT 21.452 2.244 21.505 2.419 ;
      RECT 21.366 2.243 21.452 2.428 ;
      RECT 21.28 2.242 21.366 2.44 ;
      RECT 21.26 2.241 21.275 2.448 ;
      RECT 21.18 2.24 21.26 2.46 ;
      RECT 21.155 2.24 21.18 2.473 ;
      RECT 21.13 2.24 21.155 2.488 ;
      RECT 21.125 2.24 21.13 2.51 ;
      RECT 21.12 2.24 21.125 2.528 ;
      RECT 21.115 2.24 21.12 2.545 ;
      RECT 21.11 2.24 21.115 2.558 ;
      RECT 21.105 2.24 21.11 2.568 ;
      RECT 21.065 2.24 21.105 2.653 ;
      RECT 21.05 2.24 21.065 2.738 ;
      RECT 21.04 2.241 21.05 2.75 ;
      RECT 21.005 2.246 21.04 2.755 ;
      RECT 20.965 2.255 21.005 2.755 ;
      RECT 20.95 2.265 20.965 2.755 ;
      RECT 20.945 2.275 20.95 2.755 ;
      RECT 20.925 2.302 20.945 2.755 ;
      RECT 20.875 2.385 20.925 2.755 ;
      RECT 20.87 2.447 20.875 2.755 ;
      RECT 20.86 2.46 20.87 2.755 ;
      RECT 20.85 2.482 20.86 2.755 ;
      RECT 20.84 2.507 20.85 2.75 ;
      RECT 20.835 2.545 20.84 2.743 ;
      RECT 20.825 2.655 20.835 2.738 ;
      RECT 22.22 3.576 22.235 3.835 ;
      RECT 22.22 3.591 22.24 3.834 ;
      RECT 22.136 3.591 22.24 3.832 ;
      RECT 22.136 3.605 22.245 3.831 ;
      RECT 22.05 3.647 22.25 3.828 ;
      RECT 22.045 3.59 22.235 3.823 ;
      RECT 22.045 3.661 22.255 3.82 ;
      RECT 22.04 3.692 22.255 3.818 ;
      RECT 22.045 3.689 22.27 3.808 ;
      RECT 22.04 3.735 22.285 3.793 ;
      RECT 22.04 3.763 22.29 3.778 ;
      RECT 22.05 3.565 22.22 3.828 ;
      RECT 21.81 2.575 21.98 2.745 ;
      RECT 21.775 2.575 21.98 2.74 ;
      RECT 21.765 2.575 21.98 2.733 ;
      RECT 21.76 2.56 21.93 2.73 ;
      RECT 20.59 3.097 20.855 3.54 ;
      RECT 20.585 3.068 20.8 3.538 ;
      RECT 20.58 3.222 20.86 3.533 ;
      RECT 20.585 3.117 20.86 3.533 ;
      RECT 20.585 3.128 20.87 3.52 ;
      RECT 20.585 3.075 20.83 3.538 ;
      RECT 20.59 3.062 20.8 3.54 ;
      RECT 20.59 3.06 20.75 3.54 ;
      RECT 20.691 3.052 20.75 3.54 ;
      RECT 20.605 3.053 20.75 3.54 ;
      RECT 20.691 3.051 20.74 3.54 ;
      RECT 20.495 1.866 20.67 2.165 ;
      RECT 20.545 1.828 20.67 2.165 ;
      RECT 20.53 1.83 20.756 2.157 ;
      RECT 20.53 1.833 20.795 2.144 ;
      RECT 20.53 1.834 20.805 2.13 ;
      RECT 20.485 1.885 20.805 2.12 ;
      RECT 20.53 1.835 20.81 2.115 ;
      RECT 20.485 2.045 20.815 2.105 ;
      RECT 20.47 1.905 20.81 2.045 ;
      RECT 20.465 1.921 20.81 1.985 ;
      RECT 20.51 1.845 20.81 2.115 ;
      RECT 20.545 1.826 20.631 2.165 ;
      RECT 19.005 5.02 19.175 6.49 ;
      RECT 19.005 6.315 19.18 6.485 ;
      RECT 18.635 1.74 18.805 2.93 ;
      RECT 18.635 1.74 19.105 1.91 ;
      RECT 18.635 6.97 19.105 7.14 ;
      RECT 18.635 5.95 18.805 7.14 ;
      RECT 17.645 1.74 17.815 2.93 ;
      RECT 17.645 1.74 18.115 1.91 ;
      RECT 17.645 6.97 18.115 7.14 ;
      RECT 17.645 5.95 17.815 7.14 ;
      RECT 15.795 2.635 15.965 3.865 ;
      RECT 15.85 0.855 16.02 2.805 ;
      RECT 15.795 0.575 15.965 1.025 ;
      RECT 15.795 7.855 15.965 8.305 ;
      RECT 15.85 6.075 16.02 8.025 ;
      RECT 15.795 5.015 15.965 6.245 ;
      RECT 15.275 0.575 15.445 3.865 ;
      RECT 15.275 2.075 15.68 2.405 ;
      RECT 15.275 1.235 15.68 1.565 ;
      RECT 15.275 5.015 15.445 8.305 ;
      RECT 15.275 7.315 15.68 7.645 ;
      RECT 15.275 6.475 15.68 6.805 ;
      RECT 13.2 3.126 13.205 3.298 ;
      RECT 13.195 3.119 13.2 3.388 ;
      RECT 13.19 3.113 13.195 3.407 ;
      RECT 13.17 3.107 13.19 3.417 ;
      RECT 13.155 3.102 13.17 3.425 ;
      RECT 13.118 3.096 13.155 3.423 ;
      RECT 13.032 3.082 13.118 3.419 ;
      RECT 12.946 3.064 13.032 3.414 ;
      RECT 12.86 3.045 12.946 3.408 ;
      RECT 12.83 3.033 12.86 3.404 ;
      RECT 12.81 3.027 12.83 3.403 ;
      RECT 12.745 3.025 12.81 3.401 ;
      RECT 12.73 3.025 12.745 3.393 ;
      RECT 12.715 3.025 12.73 3.38 ;
      RECT 12.71 3.025 12.715 3.37 ;
      RECT 12.695 3.025 12.71 3.348 ;
      RECT 12.68 3.025 12.695 3.315 ;
      RECT 12.675 3.025 12.68 3.293 ;
      RECT 12.665 3.025 12.675 3.275 ;
      RECT 12.65 3.025 12.665 3.253 ;
      RECT 12.63 3.025 12.65 3.215 ;
      RECT 12.98 2.31 13.015 2.749 ;
      RECT 12.98 2.31 13.02 2.748 ;
      RECT 12.925 2.37 13.02 2.747 ;
      RECT 12.79 2.542 13.02 2.746 ;
      RECT 12.9 2.42 13.02 2.746 ;
      RECT 12.79 2.542 13.045 2.736 ;
      RECT 12.845 2.487 13.125 2.653 ;
      RECT 13.02 2.281 13.025 2.744 ;
      RECT 12.875 2.457 13.165 2.53 ;
      RECT 12.89 2.44 13.02 2.746 ;
      RECT 13.025 2.28 13.195 2.468 ;
      RECT 13.015 2.283 13.195 2.468 ;
      RECT 12.52 2.16 12.69 2.47 ;
      RECT 12.52 2.16 12.695 2.443 ;
      RECT 12.52 2.16 12.7 2.42 ;
      RECT 12.52 2.16 12.71 2.37 ;
      RECT 12.515 2.265 12.71 2.34 ;
      RECT 12.55 1.835 12.72 2.313 ;
      RECT 12.55 1.835 12.735 2.234 ;
      RECT 12.54 2.045 12.735 2.234 ;
      RECT 12.55 1.845 12.745 2.149 ;
      RECT 12.48 2.587 12.485 2.79 ;
      RECT 12.47 2.575 12.48 2.9 ;
      RECT 12.445 2.575 12.47 2.94 ;
      RECT 12.365 2.575 12.445 3.025 ;
      RECT 12.355 2.575 12.365 3.095 ;
      RECT 12.33 2.575 12.355 3.118 ;
      RECT 12.31 2.575 12.33 3.153 ;
      RECT 12.265 2.585 12.31 3.196 ;
      RECT 12.255 2.597 12.265 3.233 ;
      RECT 12.235 2.611 12.255 3.253 ;
      RECT 12.225 2.629 12.235 3.269 ;
      RECT 12.21 2.655 12.225 3.279 ;
      RECT 12.195 2.696 12.21 3.293 ;
      RECT 12.185 2.731 12.195 3.303 ;
      RECT 12.18 2.747 12.185 3.308 ;
      RECT 12.17 2.762 12.18 3.313 ;
      RECT 12.15 2.805 12.17 3.323 ;
      RECT 12.13 2.842 12.15 3.336 ;
      RECT 12.095 2.865 12.13 3.354 ;
      RECT 12.085 2.879 12.095 3.37 ;
      RECT 12.065 2.889 12.085 3.38 ;
      RECT 12.06 2.898 12.065 3.388 ;
      RECT 12.05 2.905 12.06 3.395 ;
      RECT 12.04 2.912 12.05 3.403 ;
      RECT 12.025 2.922 12.04 3.411 ;
      RECT 12.015 2.936 12.025 3.421 ;
      RECT 12.005 2.948 12.015 3.433 ;
      RECT 11.99 2.97 12.005 3.446 ;
      RECT 11.98 2.992 11.99 3.457 ;
      RECT 11.97 3.012 11.98 3.466 ;
      RECT 11.965 3.027 11.97 3.473 ;
      RECT 11.935 3.06 11.965 3.487 ;
      RECT 11.925 3.095 11.935 3.502 ;
      RECT 11.92 3.102 11.925 3.508 ;
      RECT 11.9 3.117 11.92 3.515 ;
      RECT 11.895 3.132 11.9 3.523 ;
      RECT 11.89 3.141 11.895 3.528 ;
      RECT 11.875 3.147 11.89 3.535 ;
      RECT 11.87 3.153 11.875 3.543 ;
      RECT 11.865 3.157 11.87 3.55 ;
      RECT 11.86 3.161 11.865 3.56 ;
      RECT 11.85 3.166 11.86 3.57 ;
      RECT 11.83 3.177 11.85 3.598 ;
      RECT 11.815 3.189 11.83 3.625 ;
      RECT 11.795 3.202 11.815 3.65 ;
      RECT 11.775 3.217 11.795 3.674 ;
      RECT 11.76 3.232 11.775 3.689 ;
      RECT 11.755 3.243 11.76 3.698 ;
      RECT 11.69 3.288 11.755 3.708 ;
      RECT 11.655 3.347 11.69 3.721 ;
      RECT 11.65 3.37 11.655 3.727 ;
      RECT 11.645 3.377 11.65 3.729 ;
      RECT 11.63 3.387 11.645 3.732 ;
      RECT 11.6 3.412 11.63 3.736 ;
      RECT 11.595 3.43 11.6 3.74 ;
      RECT 11.59 3.437 11.595 3.741 ;
      RECT 11.57 3.445 11.59 3.745 ;
      RECT 11.56 3.452 11.57 3.749 ;
      RECT 11.516 3.463 11.56 3.756 ;
      RECT 11.43 3.491 11.516 3.772 ;
      RECT 11.37 3.515 11.43 3.79 ;
      RECT 11.325 3.525 11.37 3.804 ;
      RECT 11.266 3.533 11.325 3.818 ;
      RECT 11.18 3.54 11.266 3.837 ;
      RECT 11.155 3.545 11.18 3.852 ;
      RECT 11.075 3.548 11.155 3.855 ;
      RECT 10.995 3.552 11.075 3.842 ;
      RECT 10.986 3.555 10.995 3.827 ;
      RECT 10.9 3.555 10.986 3.812 ;
      RECT 10.84 3.557 10.9 3.789 ;
      RECT 10.836 3.56 10.84 3.779 ;
      RECT 10.75 3.56 10.836 3.764 ;
      RECT 10.675 3.56 10.75 3.74 ;
      RECT 11.99 2.569 12 2.745 ;
      RECT 11.945 2.536 11.99 2.745 ;
      RECT 11.9 2.487 11.945 2.745 ;
      RECT 11.87 2.457 11.9 2.746 ;
      RECT 11.865 2.44 11.87 2.747 ;
      RECT 11.84 2.42 11.865 2.748 ;
      RECT 11.825 2.395 11.84 2.749 ;
      RECT 11.82 2.382 11.825 2.75 ;
      RECT 11.815 2.376 11.82 2.748 ;
      RECT 11.81 2.368 11.815 2.742 ;
      RECT 11.785 2.36 11.81 2.722 ;
      RECT 11.765 2.349 11.785 2.693 ;
      RECT 11.735 2.334 11.765 2.664 ;
      RECT 11.715 2.32 11.735 2.636 ;
      RECT 11.705 2.314 11.715 2.615 ;
      RECT 11.7 2.311 11.705 2.598 ;
      RECT 11.695 2.308 11.7 2.583 ;
      RECT 11.68 2.303 11.695 2.548 ;
      RECT 11.675 2.299 11.68 2.515 ;
      RECT 11.655 2.294 11.675 2.491 ;
      RECT 11.625 2.286 11.655 2.456 ;
      RECT 11.61 2.28 11.625 2.433 ;
      RECT 11.57 2.273 11.61 2.418 ;
      RECT 11.545 2.265 11.57 2.398 ;
      RECT 11.525 2.26 11.545 2.388 ;
      RECT 11.49 2.254 11.525 2.383 ;
      RECT 11.445 2.245 11.49 2.382 ;
      RECT 11.415 2.241 11.445 2.384 ;
      RECT 11.33 2.249 11.415 2.388 ;
      RECT 11.26 2.26 11.33 2.41 ;
      RECT 11.247 2.266 11.26 2.433 ;
      RECT 11.161 2.273 11.247 2.455 ;
      RECT 11.075 2.285 11.161 2.492 ;
      RECT 11.075 2.662 11.085 2.9 ;
      RECT 11.07 2.291 11.075 2.515 ;
      RECT 11.065 2.547 11.075 2.9 ;
      RECT 11.065 2.292 11.07 2.52 ;
      RECT 11.06 2.293 11.065 2.9 ;
      RECT 11.036 2.295 11.06 2.901 ;
      RECT 10.95 2.303 11.036 2.903 ;
      RECT 10.93 2.317 10.95 2.906 ;
      RECT 10.925 2.345 10.93 2.907 ;
      RECT 10.92 2.357 10.925 2.908 ;
      RECT 10.915 2.372 10.92 2.909 ;
      RECT 10.905 2.402 10.915 2.91 ;
      RECT 10.9 2.44 10.905 2.908 ;
      RECT 10.895 2.46 10.9 2.903 ;
      RECT 10.88 2.495 10.895 2.888 ;
      RECT 10.87 2.547 10.88 2.868 ;
      RECT 10.865 2.577 10.87 2.856 ;
      RECT 10.85 2.59 10.865 2.839 ;
      RECT 10.825 2.594 10.85 2.806 ;
      RECT 10.81 2.592 10.825 2.783 ;
      RECT 10.795 2.591 10.81 2.78 ;
      RECT 10.735 2.589 10.795 2.778 ;
      RECT 10.725 2.587 10.735 2.773 ;
      RECT 10.685 2.586 10.725 2.77 ;
      RECT 10.615 2.583 10.685 2.768 ;
      RECT 10.56 2.581 10.615 2.763 ;
      RECT 10.49 2.575 10.56 2.758 ;
      RECT 10.481 2.575 10.49 2.755 ;
      RECT 10.395 2.575 10.481 2.75 ;
      RECT 10.39 2.575 10.395 2.745 ;
      RECT 11.695 1.81 11.87 2.16 ;
      RECT 11.695 1.825 11.88 2.158 ;
      RECT 11.67 1.775 11.815 2.155 ;
      RECT 11.65 1.776 11.815 2.148 ;
      RECT 11.64 1.777 11.825 2.143 ;
      RECT 11.61 1.778 11.825 2.13 ;
      RECT 11.56 1.779 11.825 2.106 ;
      RECT 11.555 1.781 11.825 2.091 ;
      RECT 11.555 1.847 11.885 2.085 ;
      RECT 11.535 1.788 11.84 2.065 ;
      RECT 11.525 1.797 11.85 1.92 ;
      RECT 11.535 1.792 11.85 2.065 ;
      RECT 11.555 1.782 11.84 2.091 ;
      RECT 11.14 3.107 11.31 3.395 ;
      RECT 11.135 3.125 11.32 3.39 ;
      RECT 11.1 3.133 11.385 3.31 ;
      RECT 11.1 3.133 11.471 3.3 ;
      RECT 11.1 3.133 11.525 3.246 ;
      RECT 11.385 3.03 11.555 3.214 ;
      RECT 11.1 3.185 11.56 3.202 ;
      RECT 11.085 3.155 11.555 3.198 ;
      RECT 11.345 3.037 11.385 3.349 ;
      RECT 11.225 3.074 11.555 3.214 ;
      RECT 11.32 3.049 11.345 3.375 ;
      RECT 11.31 3.056 11.555 3.214 ;
      RECT 11.441 2.52 11.51 2.779 ;
      RECT 11.441 2.575 11.515 2.778 ;
      RECT 11.355 2.575 11.515 2.777 ;
      RECT 11.35 2.575 11.52 2.77 ;
      RECT 11.34 2.52 11.51 2.765 ;
      RECT 10.72 1.819 10.895 2.12 ;
      RECT 10.705 1.807 10.72 2.105 ;
      RECT 10.675 1.806 10.705 2.058 ;
      RECT 10.675 1.824 10.9 2.053 ;
      RECT 10.66 1.808 10.72 2.018 ;
      RECT 10.655 1.83 10.91 1.918 ;
      RECT 10.655 1.813 10.806 1.918 ;
      RECT 10.655 1.815 10.81 1.918 ;
      RECT 10.66 1.811 10.806 2.018 ;
      RECT 10.765 3.047 10.77 3.395 ;
      RECT 10.755 3.037 10.765 3.401 ;
      RECT 10.72 3.027 10.755 3.403 ;
      RECT 10.682 3.022 10.72 3.407 ;
      RECT 10.596 3.015 10.682 3.414 ;
      RECT 10.51 3.005 10.596 3.424 ;
      RECT 10.465 3 10.51 3.432 ;
      RECT 10.461 3 10.465 3.436 ;
      RECT 10.375 3 10.461 3.443 ;
      RECT 10.36 3 10.375 3.443 ;
      RECT 10.35 2.998 10.36 3.415 ;
      RECT 10.34 2.994 10.35 3.358 ;
      RECT 10.32 2.988 10.34 3.29 ;
      RECT 10.315 2.984 10.32 3.238 ;
      RECT 10.305 2.983 10.315 3.205 ;
      RECT 10.255 2.981 10.305 3.19 ;
      RECT 10.23 2.979 10.255 3.185 ;
      RECT 10.187 2.977 10.23 3.181 ;
      RECT 10.101 2.973 10.187 3.169 ;
      RECT 10.015 2.968 10.101 3.153 ;
      RECT 9.985 2.965 10.015 3.14 ;
      RECT 9.96 2.964 9.985 3.128 ;
      RECT 9.955 2.964 9.96 3.118 ;
      RECT 9.915 2.963 9.955 3.11 ;
      RECT 9.9 2.962 9.915 3.103 ;
      RECT 9.85 2.961 9.9 3.095 ;
      RECT 9.848 2.96 9.85 3.09 ;
      RECT 9.762 2.958 9.848 3.09 ;
      RECT 9.676 2.953 9.762 3.09 ;
      RECT 9.59 2.949 9.676 3.09 ;
      RECT 9.541 2.945 9.59 3.088 ;
      RECT 9.455 2.942 9.541 3.083 ;
      RECT 9.432 2.939 9.455 3.079 ;
      RECT 9.346 2.936 9.432 3.074 ;
      RECT 9.26 2.932 9.346 3.065 ;
      RECT 9.235 2.925 9.26 3.06 ;
      RECT 9.175 2.89 9.235 3.057 ;
      RECT 9.155 2.815 9.175 3.054 ;
      RECT 9.15 2.757 9.155 3.053 ;
      RECT 9.125 2.697 9.15 3.052 ;
      RECT 9.05 2.575 9.125 3.048 ;
      RECT 9.04 2.575 9.05 3.04 ;
      RECT 9.025 2.575 9.04 3.03 ;
      RECT 9.01 2.575 9.025 3 ;
      RECT 8.995 2.575 9.01 2.945 ;
      RECT 8.98 2.575 8.995 2.883 ;
      RECT 8.955 2.575 8.98 2.808 ;
      RECT 8.95 2.575 8.955 2.758 ;
      RECT 10.295 2.12 10.315 2.429 ;
      RECT 10.281 2.122 10.33 2.426 ;
      RECT 10.281 2.127 10.35 2.417 ;
      RECT 10.195 2.125 10.33 2.411 ;
      RECT 10.195 2.133 10.385 2.394 ;
      RECT 10.16 2.135 10.385 2.393 ;
      RECT 10.13 2.143 10.385 2.384 ;
      RECT 10.12 2.148 10.405 2.37 ;
      RECT 10.16 2.138 10.405 2.37 ;
      RECT 10.16 2.141 10.415 2.358 ;
      RECT 10.13 2.143 10.425 2.345 ;
      RECT 10.13 2.147 10.435 2.288 ;
      RECT 10.12 2.152 10.44 2.203 ;
      RECT 10.281 2.12 10.315 2.426 ;
      RECT 10.16 7.855 10.33 8.305 ;
      RECT 10.215 6.075 10.385 8.025 ;
      RECT 10.16 5.015 10.33 6.245 ;
      RECT 9.72 2.223 9.725 2.435 ;
      RECT 9.595 2.22 9.61 2.435 ;
      RECT 9.06 2.25 9.13 2.435 ;
      RECT 8.945 2.25 8.98 2.43 ;
      RECT 10.066 2.552 10.085 2.746 ;
      RECT 9.98 2.507 10.066 2.747 ;
      RECT 9.97 2.46 9.98 2.749 ;
      RECT 9.965 2.44 9.97 2.75 ;
      RECT 9.945 2.405 9.965 2.751 ;
      RECT 9.93 2.355 9.945 2.752 ;
      RECT 9.91 2.292 9.93 2.753 ;
      RECT 9.9 2.255 9.91 2.754 ;
      RECT 9.885 2.244 9.9 2.755 ;
      RECT 9.88 2.236 9.885 2.753 ;
      RECT 9.87 2.235 9.88 2.745 ;
      RECT 9.84 2.232 9.87 2.724 ;
      RECT 9.765 2.227 9.84 2.669 ;
      RECT 9.75 2.223 9.765 2.615 ;
      RECT 9.74 2.223 9.75 2.51 ;
      RECT 9.725 2.223 9.74 2.443 ;
      RECT 9.71 2.223 9.72 2.433 ;
      RECT 9.655 2.222 9.71 2.43 ;
      RECT 9.61 2.22 9.655 2.433 ;
      RECT 9.582 2.22 9.595 2.436 ;
      RECT 9.496 2.224 9.582 2.438 ;
      RECT 9.41 2.23 9.496 2.443 ;
      RECT 9.39 2.234 9.41 2.445 ;
      RECT 9.388 2.235 9.39 2.444 ;
      RECT 9.302 2.237 9.388 2.443 ;
      RECT 9.216 2.242 9.302 2.44 ;
      RECT 9.13 2.247 9.216 2.437 ;
      RECT 8.98 2.25 9.06 2.433 ;
      RECT 9.64 5.015 9.81 8.305 ;
      RECT 9.64 7.315 10.045 7.645 ;
      RECT 9.64 6.475 10.045 6.805 ;
      RECT 9.756 3.225 9.805 3.559 ;
      RECT 9.756 3.225 9.81 3.558 ;
      RECT 9.67 3.225 9.81 3.557 ;
      RECT 9.445 3.333 9.815 3.555 ;
      RECT 9.67 3.225 9.84 3.548 ;
      RECT 9.64 3.237 9.845 3.539 ;
      RECT 9.625 3.255 9.85 3.536 ;
      RECT 9.44 3.339 9.85 3.463 ;
      RECT 9.435 3.346 9.85 3.423 ;
      RECT 9.45 3.312 9.85 3.536 ;
      RECT 9.611 3.258 9.815 3.555 ;
      RECT 9.525 3.278 9.85 3.536 ;
      RECT 9.625 3.252 9.845 3.539 ;
      RECT 9.395 2.576 9.585 2.77 ;
      RECT 9.39 2.578 9.585 2.769 ;
      RECT 9.385 2.582 9.6 2.766 ;
      RECT 9.4 2.575 9.6 2.766 ;
      RECT 9.385 2.685 9.605 2.761 ;
      RECT 8.68 3.185 8.771 3.483 ;
      RECT 8.675 3.187 8.85 3.478 ;
      RECT 8.68 3.185 8.85 3.478 ;
      RECT 8.675 3.191 8.87 3.476 ;
      RECT 8.675 3.246 8.91 3.475 ;
      RECT 8.675 3.281 8.925 3.469 ;
      RECT 8.675 3.315 8.935 3.459 ;
      RECT 8.665 3.195 8.87 3.31 ;
      RECT 8.665 3.215 8.885 3.31 ;
      RECT 8.665 3.198 8.875 3.31 ;
      RECT 8.89 1.966 8.895 2.028 ;
      RECT 8.885 1.888 8.89 2.051 ;
      RECT 8.88 1.845 8.885 2.062 ;
      RECT 8.875 1.835 8.88 2.074 ;
      RECT 8.87 1.835 8.875 2.083 ;
      RECT 8.845 1.835 8.87 2.115 ;
      RECT 8.84 1.835 8.845 2.148 ;
      RECT 8.825 1.835 8.84 2.173 ;
      RECT 8.815 1.835 8.825 2.2 ;
      RECT 8.81 1.835 8.815 2.213 ;
      RECT 8.805 1.835 8.81 2.228 ;
      RECT 8.795 1.835 8.805 2.243 ;
      RECT 8.79 1.835 8.795 2.263 ;
      RECT 8.765 1.835 8.79 2.298 ;
      RECT 8.72 1.835 8.765 2.343 ;
      RECT 8.71 1.835 8.72 2.356 ;
      RECT 8.625 1.92 8.71 2.363 ;
      RECT 8.59 2.042 8.625 2.372 ;
      RECT 8.585 2.082 8.59 2.376 ;
      RECT 8.565 2.105 8.585 2.378 ;
      RECT 8.56 2.135 8.565 2.381 ;
      RECT 8.55 2.147 8.56 2.382 ;
      RECT 8.505 2.17 8.55 2.387 ;
      RECT 8.465 2.2 8.505 2.395 ;
      RECT 8.43 2.212 8.465 2.401 ;
      RECT 8.425 2.217 8.43 2.405 ;
      RECT 8.355 2.227 8.425 2.412 ;
      RECT 8.315 2.237 8.355 2.422 ;
      RECT 8.295 2.242 8.315 2.428 ;
      RECT 8.285 2.246 8.295 2.433 ;
      RECT 8.28 2.249 8.285 2.436 ;
      RECT 8.27 2.25 8.28 2.437 ;
      RECT 8.245 2.252 8.27 2.441 ;
      RECT 8.235 2.257 8.245 2.444 ;
      RECT 8.19 2.265 8.235 2.445 ;
      RECT 8.065 2.27 8.19 2.445 ;
      RECT 8.62 2.567 8.64 2.749 ;
      RECT 8.571 2.552 8.62 2.748 ;
      RECT 8.485 2.567 8.64 2.746 ;
      RECT 8.47 2.567 8.64 2.745 ;
      RECT 8.435 2.545 8.605 2.73 ;
      RECT 8.505 3.565 8.52 3.774 ;
      RECT 8.505 3.573 8.525 3.773 ;
      RECT 8.45 3.573 8.525 3.772 ;
      RECT 8.43 3.577 8.53 3.77 ;
      RECT 8.41 3.527 8.45 3.769 ;
      RECT 8.355 3.585 8.535 3.767 ;
      RECT 8.32 3.542 8.45 3.765 ;
      RECT 8.316 3.545 8.505 3.764 ;
      RECT 8.23 3.553 8.505 3.762 ;
      RECT 8.23 3.597 8.54 3.755 ;
      RECT 8.22 3.69 8.54 3.753 ;
      RECT 8.23 3.609 8.545 3.738 ;
      RECT 8.23 3.63 8.56 3.708 ;
      RECT 8.23 3.657 8.565 3.678 ;
      RECT 8.355 3.535 8.45 3.767 ;
      RECT 7.985 2.58 7.99 3.118 ;
      RECT 7.79 2.91 7.795 3.105 ;
      RECT 6.09 2.575 6.105 2.955 ;
      RECT 8.155 2.575 8.16 2.745 ;
      RECT 8.15 2.575 8.155 2.755 ;
      RECT 8.145 2.575 8.15 2.768 ;
      RECT 8.12 2.575 8.145 2.81 ;
      RECT 8.095 2.575 8.12 2.883 ;
      RECT 8.08 2.575 8.095 2.935 ;
      RECT 8.075 2.575 8.08 2.965 ;
      RECT 8.05 2.575 8.075 3.005 ;
      RECT 8.035 2.575 8.05 3.06 ;
      RECT 8.03 2.575 8.035 3.093 ;
      RECT 8.005 2.575 8.03 3.113 ;
      RECT 7.99 2.575 8.005 3.119 ;
      RECT 7.92 2.61 7.985 3.115 ;
      RECT 7.87 2.665 7.92 3.11 ;
      RECT 7.86 2.697 7.87 3.108 ;
      RECT 7.855 2.722 7.86 3.108 ;
      RECT 7.835 2.795 7.855 3.108 ;
      RECT 7.825 2.875 7.835 3.107 ;
      RECT 7.81 2.905 7.825 3.107 ;
      RECT 7.795 2.91 7.81 3.106 ;
      RECT 7.735 2.912 7.79 3.103 ;
      RECT 7.705 2.917 7.735 3.099 ;
      RECT 7.703 2.92 7.705 3.098 ;
      RECT 7.617 2.922 7.703 3.095 ;
      RECT 7.531 2.928 7.617 3.089 ;
      RECT 7.445 2.933 7.531 3.083 ;
      RECT 7.372 2.938 7.445 3.084 ;
      RECT 7.286 2.944 7.372 3.092 ;
      RECT 7.2 2.95 7.286 3.101 ;
      RECT 7.18 2.954 7.2 3.106 ;
      RECT 7.133 2.956 7.18 3.109 ;
      RECT 7.047 2.961 7.133 3.115 ;
      RECT 6.961 2.966 7.047 3.124 ;
      RECT 6.875 2.972 6.961 3.132 ;
      RECT 6.79 2.97 6.875 3.141 ;
      RECT 6.786 2.965 6.79 3.145 ;
      RECT 6.7 2.96 6.786 3.137 ;
      RECT 6.636 2.951 6.7 3.125 ;
      RECT 6.55 2.942 6.636 3.112 ;
      RECT 6.526 2.935 6.55 3.103 ;
      RECT 6.44 2.929 6.526 3.09 ;
      RECT 6.4 2.922 6.44 3.076 ;
      RECT 6.395 2.912 6.4 3.072 ;
      RECT 6.385 2.9 6.395 3.071 ;
      RECT 6.365 2.87 6.385 3.068 ;
      RECT 6.31 2.79 6.365 3.062 ;
      RECT 6.29 2.709 6.31 3.057 ;
      RECT 6.27 2.667 6.29 3.053 ;
      RECT 6.245 2.62 6.27 3.047 ;
      RECT 6.24 2.595 6.245 3.044 ;
      RECT 6.205 2.575 6.24 3.039 ;
      RECT 6.196 2.575 6.205 3.032 ;
      RECT 6.11 2.575 6.196 3.002 ;
      RECT 6.105 2.575 6.11 2.965 ;
      RECT 6.07 2.575 6.09 2.887 ;
      RECT 6.065 2.617 6.07 2.852 ;
      RECT 6.06 2.692 6.065 2.808 ;
      RECT 7.51 2.497 7.685 2.745 ;
      RECT 7.51 2.497 7.69 2.743 ;
      RECT 7.505 2.529 7.69 2.703 ;
      RECT 7.535 2.47 7.705 2.69 ;
      RECT 7.5 2.547 7.705 2.623 ;
      RECT 6.81 2.01 6.98 2.185 ;
      RECT 6.81 2.01 7.152 2.177 ;
      RECT 6.81 2.01 7.235 2.171 ;
      RECT 6.81 2.01 7.27 2.167 ;
      RECT 6.81 2.01 7.29 2.166 ;
      RECT 6.81 2.01 7.376 2.162 ;
      RECT 7.27 1.835 7.44 2.157 ;
      RECT 6.845 1.942 7.47 2.155 ;
      RECT 6.835 1.997 7.475 2.153 ;
      RECT 6.81 2.033 7.485 2.148 ;
      RECT 6.81 2.06 7.49 2.078 ;
      RECT 6.875 1.885 7.45 2.155 ;
      RECT 7.066 1.87 7.45 2.155 ;
      RECT 6.9 1.873 7.45 2.155 ;
      RECT 6.98 1.871 7.066 2.182 ;
      RECT 7.066 1.868 7.445 2.155 ;
      RECT 7.25 1.845 7.445 2.155 ;
      RECT 7.152 1.866 7.445 2.155 ;
      RECT 7.235 1.86 7.25 2.168 ;
      RECT 7.385 3.225 7.39 3.425 ;
      RECT 6.85 3.29 6.895 3.425 ;
      RECT 7.42 3.225 7.44 3.398 ;
      RECT 7.39 3.225 7.42 3.413 ;
      RECT 7.325 3.225 7.385 3.45 ;
      RECT 7.31 3.225 7.325 3.48 ;
      RECT 7.295 3.225 7.31 3.493 ;
      RECT 7.275 3.225 7.295 3.508 ;
      RECT 7.27 3.225 7.275 3.517 ;
      RECT 7.26 3.229 7.27 3.522 ;
      RECT 7.245 3.239 7.26 3.533 ;
      RECT 7.22 3.255 7.245 3.543 ;
      RECT 7.21 3.269 7.22 3.545 ;
      RECT 7.19 3.281 7.21 3.542 ;
      RECT 7.16 3.302 7.19 3.536 ;
      RECT 7.15 3.314 7.16 3.531 ;
      RECT 7.14 3.312 7.15 3.528 ;
      RECT 7.125 3.311 7.14 3.523 ;
      RECT 7.12 3.31 7.125 3.518 ;
      RECT 7.085 3.308 7.12 3.508 ;
      RECT 7.065 3.305 7.085 3.49 ;
      RECT 7.055 3.303 7.065 3.485 ;
      RECT 7.045 3.302 7.055 3.48 ;
      RECT 7.01 3.3 7.045 3.468 ;
      RECT 6.955 3.296 7.01 3.448 ;
      RECT 6.945 3.294 6.955 3.433 ;
      RECT 6.94 3.294 6.945 3.428 ;
      RECT 6.895 3.292 6.94 3.425 ;
      RECT 6.8 3.29 6.85 3.429 ;
      RECT 6.79 3.291 6.8 3.434 ;
      RECT 6.73 3.298 6.79 3.448 ;
      RECT 6.705 3.306 6.73 3.468 ;
      RECT 6.695 3.31 6.705 3.48 ;
      RECT 6.69 3.311 6.695 3.485 ;
      RECT 6.675 3.313 6.69 3.488 ;
      RECT 6.66 3.315 6.675 3.493 ;
      RECT 6.655 3.315 6.66 3.496 ;
      RECT 6.61 3.32 6.655 3.507 ;
      RECT 6.605 3.324 6.61 3.519 ;
      RECT 6.58 3.32 6.605 3.523 ;
      RECT 6.57 3.316 6.58 3.527 ;
      RECT 6.56 3.315 6.57 3.531 ;
      RECT 6.545 3.305 6.56 3.537 ;
      RECT 6.54 3.293 6.545 3.541 ;
      RECT 6.535 3.29 6.54 3.542 ;
      RECT 6.53 3.287 6.535 3.544 ;
      RECT 6.515 3.275 6.53 3.543 ;
      RECT 6.5 3.257 6.515 3.54 ;
      RECT 6.48 3.236 6.5 3.533 ;
      RECT 6.415 3.225 6.48 3.505 ;
      RECT 6.411 3.225 6.415 3.484 ;
      RECT 6.325 3.225 6.411 3.454 ;
      RECT 6.31 3.225 6.325 3.41 ;
      RECT 6.885 2.325 6.89 2.56 ;
      RECT 6.015 2.241 6.02 2.445 ;
      RECT 6.595 2.27 6.6 2.425 ;
      RECT 6.515 2.25 6.52 2.425 ;
      RECT 7.185 2.392 7.2 2.745 ;
      RECT 7.111 2.377 7.185 2.745 ;
      RECT 7.025 2.36 7.111 2.745 ;
      RECT 7.015 2.35 7.025 2.743 ;
      RECT 7.01 2.348 7.015 2.738 ;
      RECT 6.995 2.346 7.01 2.724 ;
      RECT 6.925 2.338 6.995 2.664 ;
      RECT 6.905 2.329 6.925 2.598 ;
      RECT 6.9 2.326 6.905 2.578 ;
      RECT 6.89 2.325 6.9 2.568 ;
      RECT 6.88 2.325 6.885 2.552 ;
      RECT 6.87 2.324 6.88 2.542 ;
      RECT 6.86 2.322 6.87 2.53 ;
      RECT 6.845 2.319 6.86 2.51 ;
      RECT 6.835 2.317 6.845 2.495 ;
      RECT 6.815 2.314 6.835 2.483 ;
      RECT 6.81 2.312 6.815 2.473 ;
      RECT 6.785 2.31 6.81 2.46 ;
      RECT 6.755 2.305 6.785 2.445 ;
      RECT 6.675 2.296 6.755 2.436 ;
      RECT 6.63 2.285 6.675 2.429 ;
      RECT 6.61 2.276 6.63 2.426 ;
      RECT 6.6 2.271 6.61 2.425 ;
      RECT 6.555 2.265 6.595 2.425 ;
      RECT 6.54 2.257 6.555 2.425 ;
      RECT 6.52 2.252 6.54 2.425 ;
      RECT 6.5 2.249 6.515 2.425 ;
      RECT 6.417 2.248 6.5 2.424 ;
      RECT 6.331 2.247 6.417 2.42 ;
      RECT 6.245 2.245 6.331 2.417 ;
      RECT 6.192 2.244 6.245 2.419 ;
      RECT 6.106 2.243 6.192 2.428 ;
      RECT 6.02 2.242 6.106 2.44 ;
      RECT 6 2.241 6.015 2.448 ;
      RECT 5.92 2.24 6 2.46 ;
      RECT 5.895 2.24 5.92 2.473 ;
      RECT 5.87 2.24 5.895 2.488 ;
      RECT 5.865 2.24 5.87 2.51 ;
      RECT 5.86 2.24 5.865 2.528 ;
      RECT 5.855 2.24 5.86 2.545 ;
      RECT 5.85 2.24 5.855 2.558 ;
      RECT 5.845 2.24 5.85 2.568 ;
      RECT 5.805 2.24 5.845 2.653 ;
      RECT 5.79 2.24 5.805 2.738 ;
      RECT 5.78 2.241 5.79 2.75 ;
      RECT 5.745 2.246 5.78 2.755 ;
      RECT 5.705 2.255 5.745 2.755 ;
      RECT 5.69 2.265 5.705 2.755 ;
      RECT 5.685 2.275 5.69 2.755 ;
      RECT 5.665 2.302 5.685 2.755 ;
      RECT 5.615 2.385 5.665 2.755 ;
      RECT 5.61 2.447 5.615 2.755 ;
      RECT 5.6 2.46 5.61 2.755 ;
      RECT 5.59 2.482 5.6 2.755 ;
      RECT 5.58 2.507 5.59 2.75 ;
      RECT 5.575 2.545 5.58 2.743 ;
      RECT 5.565 2.655 5.575 2.738 ;
      RECT 6.96 3.576 6.975 3.835 ;
      RECT 6.96 3.591 6.98 3.834 ;
      RECT 6.876 3.591 6.98 3.832 ;
      RECT 6.876 3.605 6.985 3.831 ;
      RECT 6.79 3.647 6.99 3.828 ;
      RECT 6.785 3.59 6.975 3.823 ;
      RECT 6.785 3.661 6.995 3.82 ;
      RECT 6.78 3.692 6.995 3.818 ;
      RECT 6.785 3.689 7.01 3.808 ;
      RECT 6.78 3.735 7.025 3.793 ;
      RECT 6.78 3.763 7.03 3.778 ;
      RECT 6.79 3.565 6.96 3.828 ;
      RECT 6.55 2.575 6.72 2.745 ;
      RECT 6.515 2.575 6.72 2.74 ;
      RECT 6.505 2.575 6.72 2.733 ;
      RECT 6.5 2.56 6.67 2.73 ;
      RECT 5.33 3.097 5.595 3.54 ;
      RECT 5.325 3.068 5.54 3.538 ;
      RECT 5.32 3.222 5.6 3.533 ;
      RECT 5.325 3.117 5.6 3.533 ;
      RECT 5.325 3.128 5.61 3.52 ;
      RECT 5.325 3.075 5.57 3.538 ;
      RECT 5.33 3.062 5.54 3.54 ;
      RECT 5.33 3.06 5.49 3.54 ;
      RECT 5.431 3.052 5.49 3.54 ;
      RECT 5.345 3.053 5.49 3.54 ;
      RECT 5.431 3.051 5.48 3.54 ;
      RECT 5.235 1.866 5.41 2.165 ;
      RECT 5.285 1.828 5.41 2.165 ;
      RECT 5.27 1.83 5.496 2.157 ;
      RECT 5.27 1.833 5.535 2.144 ;
      RECT 5.27 1.834 5.545 2.13 ;
      RECT 5.225 1.885 5.545 2.12 ;
      RECT 5.27 1.835 5.55 2.115 ;
      RECT 5.225 2.045 5.555 2.105 ;
      RECT 5.21 1.905 5.55 2.045 ;
      RECT 5.205 1.921 5.55 1.985 ;
      RECT 5.25 1.845 5.55 2.115 ;
      RECT 5.285 1.826 5.371 2.165 ;
      RECT 2.665 7.855 2.835 8.305 ;
      RECT 2.72 6.075 2.89 8.025 ;
      RECT 2.665 5.015 2.835 6.245 ;
      RECT 2.145 5.015 2.315 8.305 ;
      RECT 2.145 7.315 2.55 7.645 ;
      RECT 2.145 6.475 2.55 6.805 ;
      RECT 80.045 7.8 80.215 8.31 ;
      RECT 79.055 0.57 79.225 1.08 ;
      RECT 79.055 2.39 79.225 3.86 ;
      RECT 79.055 5.02 79.225 6.49 ;
      RECT 79.055 7.8 79.225 8.31 ;
      RECT 77.695 0.575 77.865 3.865 ;
      RECT 77.695 5.015 77.865 8.305 ;
      RECT 77.265 0.575 77.435 1.085 ;
      RECT 77.265 1.655 77.435 3.865 ;
      RECT 77.265 5.015 77.435 7.225 ;
      RECT 77.265 7.795 77.435 8.305 ;
      RECT 72.06 5.015 72.23 8.305 ;
      RECT 71.63 5.015 71.8 7.225 ;
      RECT 71.63 7.795 71.8 8.305 ;
      RECT 64.785 7.8 64.955 8.31 ;
      RECT 63.795 0.57 63.965 1.08 ;
      RECT 63.795 2.39 63.965 3.86 ;
      RECT 63.795 5.02 63.965 6.49 ;
      RECT 63.795 7.8 63.965 8.31 ;
      RECT 62.435 0.575 62.605 3.865 ;
      RECT 62.435 5.015 62.605 8.305 ;
      RECT 62.005 0.575 62.175 1.085 ;
      RECT 62.005 1.655 62.175 3.865 ;
      RECT 62.005 5.015 62.175 7.225 ;
      RECT 62.005 7.795 62.175 8.305 ;
      RECT 56.8 5.015 56.97 8.305 ;
      RECT 56.37 5.015 56.54 7.225 ;
      RECT 56.37 7.795 56.54 8.305 ;
      RECT 49.525 7.8 49.695 8.31 ;
      RECT 48.535 0.57 48.705 1.08 ;
      RECT 48.535 2.39 48.705 3.86 ;
      RECT 48.535 5.02 48.705 6.49 ;
      RECT 48.535 7.8 48.705 8.31 ;
      RECT 47.175 0.575 47.345 3.865 ;
      RECT 47.175 5.015 47.345 8.305 ;
      RECT 46.745 0.575 46.915 1.085 ;
      RECT 46.745 1.655 46.915 3.865 ;
      RECT 46.745 5.015 46.915 7.225 ;
      RECT 46.745 7.795 46.915 8.305 ;
      RECT 41.54 5.015 41.71 8.305 ;
      RECT 41.11 5.015 41.28 7.225 ;
      RECT 41.11 7.795 41.28 8.305 ;
      RECT 34.265 7.8 34.435 8.31 ;
      RECT 33.275 0.57 33.445 1.08 ;
      RECT 33.275 2.39 33.445 3.86 ;
      RECT 33.275 5.02 33.445 6.49 ;
      RECT 33.275 7.8 33.445 8.31 ;
      RECT 31.915 0.575 32.085 3.865 ;
      RECT 31.915 5.015 32.085 8.305 ;
      RECT 31.485 0.575 31.655 1.085 ;
      RECT 31.485 1.655 31.655 3.865 ;
      RECT 31.485 5.015 31.655 7.225 ;
      RECT 31.485 7.795 31.655 8.305 ;
      RECT 26.28 5.015 26.45 8.305 ;
      RECT 25.85 5.015 26.02 7.225 ;
      RECT 25.85 7.795 26.02 8.305 ;
      RECT 19.005 7.8 19.175 8.31 ;
      RECT 18.015 0.57 18.185 1.08 ;
      RECT 18.015 2.39 18.185 3.86 ;
      RECT 18.015 5.02 18.185 6.49 ;
      RECT 18.015 7.8 18.185 8.31 ;
      RECT 16.655 0.575 16.825 3.865 ;
      RECT 16.655 5.015 16.825 8.305 ;
      RECT 16.225 0.575 16.395 1.085 ;
      RECT 16.225 1.655 16.395 3.865 ;
      RECT 16.225 5.015 16.395 7.225 ;
      RECT 16.225 7.795 16.395 8.305 ;
      RECT 11.02 5.015 11.19 8.305 ;
      RECT 10.59 5.015 10.76 7.225 ;
      RECT 10.59 7.795 10.76 8.305 ;
      RECT 3.095 5.015 3.265 7.225 ;
      RECT 3.095 7.795 3.265 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2ya_8_b0r1

MACRO sky130_osu_ring_oscillator_mpr2ya_8_b0r2
  CLASS BLOCK ;
  ORIGIN -1.48 0 ;
  FOREIGN sky130_osu_ring_oscillator_mpr2ya_8_b0r2 ;
  SIZE 79.095 BY 8.88 ;
  PIN X1_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 18.995 0.915 19.165 1.085 ;
        RECT 18.99 0.91 19.16 1.08 ;
        RECT 18.99 2.39 19.16 2.56 ;
      LAYER li1 ;
        RECT 18.995 0.915 19.165 1.085 ;
        RECT 18.99 0.57 19.16 1.08 ;
        RECT 18.99 2.39 19.16 3.86 ;
      LAYER met1 ;
        RECT 18.93 2.36 19.22 2.59 ;
        RECT 18.93 0.88 19.22 1.11 ;
        RECT 18.99 0.88 19.16 2.59 ;
    END
  END X1_Y1
  PIN X2_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 34.255 0.915 34.425 1.085 ;
        RECT 34.25 0.91 34.42 1.08 ;
        RECT 34.25 2.39 34.42 2.56 ;
      LAYER li1 ;
        RECT 34.255 0.915 34.425 1.085 ;
        RECT 34.25 0.57 34.42 1.08 ;
        RECT 34.25 2.39 34.42 3.86 ;
      LAYER met1 ;
        RECT 34.19 2.36 34.48 2.59 ;
        RECT 34.19 0.88 34.48 1.11 ;
        RECT 34.25 0.88 34.42 2.59 ;
    END
  END X2_Y1
  PIN X3_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 49.515 0.915 49.685 1.085 ;
        RECT 49.51 0.91 49.68 1.08 ;
        RECT 49.51 2.39 49.68 2.56 ;
      LAYER li1 ;
        RECT 49.515 0.915 49.685 1.085 ;
        RECT 49.51 0.57 49.68 1.08 ;
        RECT 49.51 2.39 49.68 3.86 ;
      LAYER met1 ;
        RECT 49.45 2.36 49.74 2.59 ;
        RECT 49.45 0.88 49.74 1.11 ;
        RECT 49.51 0.88 49.68 2.59 ;
    END
  END X3_Y1
  PIN X4_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 64.775 0.915 64.945 1.085 ;
        RECT 64.77 0.91 64.94 1.08 ;
        RECT 64.77 2.39 64.94 2.56 ;
      LAYER li1 ;
        RECT 64.775 0.915 64.945 1.085 ;
        RECT 64.77 0.57 64.94 1.08 ;
        RECT 64.77 2.39 64.94 3.86 ;
      LAYER met1 ;
        RECT 64.71 2.36 65 2.59 ;
        RECT 64.71 0.88 65 1.11 ;
        RECT 64.77 0.88 64.94 2.59 ;
    END
  END X4_Y1
  PIN X5_Y1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.143 ;
    PORT
      LAYER mcon ;
        RECT 80.035 0.915 80.205 1.085 ;
        RECT 80.03 0.91 80.2 1.08 ;
        RECT 80.03 2.39 80.2 2.56 ;
      LAYER li1 ;
        RECT 80.035 0.915 80.205 1.085 ;
        RECT 80.03 0.57 80.2 1.08 ;
        RECT 80.03 2.39 80.2 3.86 ;
      LAYER met1 ;
        RECT 79.97 2.36 80.26 2.59 ;
        RECT 79.97 0.88 80.26 1.11 ;
        RECT 80.03 0.88 80.2 2.59 ;
    END
  END X5_Y1
  PIN s1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 14.76 2.705 15.1 3.055 ;
        RECT 14.755 5.86 15.095 6.21 ;
        RECT 14.835 2.705 15.01 6.21 ;
      LAYER li1 ;
        RECT 14.84 1.66 15.01 2.935 ;
        RECT 14.84 5.945 15.01 7.22 ;
        RECT 9.205 5.945 9.375 7.22 ;
      LAYER met1 ;
        RECT 14.76 2.765 15.24 2.935 ;
        RECT 14.76 2.705 15.1 3.055 ;
        RECT 9.145 5.945 15.24 6.115 ;
        RECT 14.755 5.86 15.095 6.21 ;
        RECT 9.145 5.915 9.435 6.145 ;
      LAYER via1 ;
        RECT 14.855 5.96 15.005 6.11 ;
        RECT 14.86 2.805 15.01 2.955 ;
      LAYER mcon ;
        RECT 9.205 5.945 9.375 6.115 ;
        RECT 14.84 5.945 15.01 6.115 ;
        RECT 14.84 2.765 15.01 2.935 ;
    END
  END s1
  PIN s2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 30.02 2.705 30.36 3.055 ;
        RECT 30.015 5.86 30.355 6.21 ;
        RECT 30.095 2.705 30.27 6.21 ;
      LAYER li1 ;
        RECT 30.1 1.66 30.27 2.935 ;
        RECT 30.1 5.945 30.27 7.22 ;
        RECT 24.465 5.945 24.635 7.22 ;
      LAYER met1 ;
        RECT 30.02 2.765 30.5 2.935 ;
        RECT 30.02 2.705 30.36 3.055 ;
        RECT 24.405 5.945 30.5 6.115 ;
        RECT 30.015 5.86 30.355 6.21 ;
        RECT 24.405 5.915 24.695 6.145 ;
      LAYER via1 ;
        RECT 30.115 5.96 30.265 6.11 ;
        RECT 30.12 2.805 30.27 2.955 ;
      LAYER mcon ;
        RECT 24.465 5.945 24.635 6.115 ;
        RECT 30.1 5.945 30.27 6.115 ;
        RECT 30.1 2.765 30.27 2.935 ;
    END
  END s2
  PIN s3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 45.28 2.705 45.62 3.055 ;
        RECT 45.275 5.86 45.615 6.21 ;
        RECT 45.355 2.705 45.53 6.21 ;
      LAYER li1 ;
        RECT 45.36 1.66 45.53 2.935 ;
        RECT 45.36 5.945 45.53 7.22 ;
        RECT 39.725 5.945 39.895 7.22 ;
      LAYER met1 ;
        RECT 45.28 2.765 45.76 2.935 ;
        RECT 45.28 2.705 45.62 3.055 ;
        RECT 39.665 5.945 45.76 6.115 ;
        RECT 45.275 5.86 45.615 6.21 ;
        RECT 39.665 5.915 39.955 6.145 ;
      LAYER via1 ;
        RECT 45.375 5.96 45.525 6.11 ;
        RECT 45.38 2.805 45.53 2.955 ;
      LAYER mcon ;
        RECT 39.725 5.945 39.895 6.115 ;
        RECT 45.36 5.945 45.53 6.115 ;
        RECT 45.36 2.765 45.53 2.935 ;
    END
  END s3
  PIN s4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 60.54 2.705 60.88 3.055 ;
        RECT 60.535 5.86 60.875 6.21 ;
        RECT 60.615 2.705 60.79 6.21 ;
      LAYER li1 ;
        RECT 60.62 1.66 60.79 2.935 ;
        RECT 60.62 5.945 60.79 7.22 ;
        RECT 54.985 5.945 55.155 7.22 ;
      LAYER met1 ;
        RECT 60.54 2.765 61.02 2.935 ;
        RECT 60.54 2.705 60.88 3.055 ;
        RECT 54.925 5.945 61.02 6.115 ;
        RECT 60.535 5.86 60.875 6.21 ;
        RECT 54.925 5.915 55.215 6.145 ;
      LAYER via1 ;
        RECT 60.635 5.96 60.785 6.11 ;
        RECT 60.64 2.805 60.79 2.955 ;
      LAYER mcon ;
        RECT 54.985 5.945 55.155 6.115 ;
        RECT 60.62 5.945 60.79 6.115 ;
        RECT 60.62 2.765 60.79 2.935 ;
    END
  END s4
  PIN s5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.629 ;
    PORT
      LAYER met2 ;
        RECT 75.8 2.705 76.14 3.055 ;
        RECT 75.795 5.86 76.135 6.21 ;
        RECT 75.875 2.705 76.05 6.21 ;
      LAYER li1 ;
        RECT 75.88 1.66 76.05 2.935 ;
        RECT 75.88 5.945 76.05 7.22 ;
        RECT 70.245 5.945 70.415 7.22 ;
      LAYER met1 ;
        RECT 75.8 2.765 76.28 2.935 ;
        RECT 75.8 2.705 76.14 3.055 ;
        RECT 70.185 5.945 76.28 6.115 ;
        RECT 75.795 5.86 76.135 6.21 ;
        RECT 70.185 5.915 70.475 6.145 ;
      LAYER via1 ;
        RECT 75.895 5.96 76.045 6.11 ;
        RECT 75.9 2.805 76.05 2.955 ;
      LAYER mcon ;
        RECT 70.245 5.945 70.415 6.115 ;
        RECT 75.88 5.945 76.05 6.115 ;
        RECT 75.88 2.765 76.05 2.935 ;
    END
  END s5
  PIN start
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.543 ;
    PORT
      LAYER li1 ;
        RECT 1.71 5.945 1.88 7.22 ;
      LAYER met1 ;
        RECT 1.65 5.945 2.11 6.115 ;
        RECT 1.65 5.915 1.94 6.145 ;
      LAYER mcon ;
        RECT 1.71 5.945 1.88 6.115 ;
    END
  END start
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 1.48 4.14 80.575 4.745 ;
        RECT 66.065 4.135 80.575 4.745 ;
        RECT 78.44 4.13 80.42 4.75 ;
        RECT 79.6 3.4 79.77 5.48 ;
        RECT 78.61 3.4 78.78 5.48 ;
        RECT 75.87 3.405 76.04 5.475 ;
        RECT 73.095 3.635 73.265 4.745 ;
        RECT 71.175 3.635 71.345 4.745 ;
        RECT 70.235 3.635 70.405 5.475 ;
        RECT 68.775 3.635 68.945 4.745 ;
        RECT 66.855 3.635 67.025 4.745 ;
        RECT 50.805 4.135 65.315 4.745 ;
        RECT 63.18 4.13 65.16 4.75 ;
        RECT 64.34 3.4 64.51 5.48 ;
        RECT 63.35 3.4 63.52 5.48 ;
        RECT 60.61 3.405 60.78 5.475 ;
        RECT 57.835 3.635 58.005 4.745 ;
        RECT 55.915 3.635 56.085 4.745 ;
        RECT 54.975 3.635 55.145 5.475 ;
        RECT 53.515 3.635 53.685 4.745 ;
        RECT 51.595 3.635 51.765 4.745 ;
        RECT 35.545 4.135 50.055 4.745 ;
        RECT 47.92 4.13 49.9 4.75 ;
        RECT 49.08 3.4 49.25 5.48 ;
        RECT 48.09 3.4 48.26 5.48 ;
        RECT 45.35 3.405 45.52 5.475 ;
        RECT 42.575 3.635 42.745 4.745 ;
        RECT 40.655 3.635 40.825 4.745 ;
        RECT 39.715 3.635 39.885 5.475 ;
        RECT 38.255 3.635 38.425 4.745 ;
        RECT 36.335 3.635 36.505 4.745 ;
        RECT 20.285 4.135 34.795 4.745 ;
        RECT 32.66 4.13 34.64 4.75 ;
        RECT 33.82 3.4 33.99 5.48 ;
        RECT 32.83 3.4 33 5.48 ;
        RECT 30.09 3.405 30.26 5.475 ;
        RECT 27.315 3.635 27.485 4.745 ;
        RECT 25.395 3.635 25.565 4.745 ;
        RECT 24.455 3.635 24.625 5.475 ;
        RECT 22.995 3.635 23.165 4.745 ;
        RECT 21.075 3.635 21.245 4.745 ;
        RECT 5.025 4.135 19.535 4.745 ;
        RECT 17.4 4.13 19.38 4.75 ;
        RECT 18.56 3.4 18.73 5.48 ;
        RECT 17.57 3.4 17.74 5.48 ;
        RECT 14.83 3.405 15 5.475 ;
        RECT 12.055 3.635 12.225 4.745 ;
        RECT 10.135 3.635 10.305 4.745 ;
        RECT 9.195 3.635 9.365 5.475 ;
        RECT 7.735 3.635 7.905 4.745 ;
        RECT 5.815 3.635 5.985 4.745 ;
        RECT 3.51 4.14 3.68 8.305 ;
        RECT 1.7 4.14 1.87 5.475 ;
      LAYER met1 ;
        RECT 1.48 4.14 80.575 4.745 ;
        RECT 66.065 4.135 80.575 4.745 ;
        RECT 78.44 4.13 80.42 4.75 ;
        RECT 66.065 3.98 74.805 4.745 ;
        RECT 50.805 4.135 65.315 4.745 ;
        RECT 63.18 4.13 65.16 4.75 ;
        RECT 50.805 3.98 59.545 4.745 ;
        RECT 35.545 4.135 50.055 4.745 ;
        RECT 47.92 4.13 49.9 4.75 ;
        RECT 35.545 3.98 44.285 4.745 ;
        RECT 20.285 4.135 34.795 4.745 ;
        RECT 32.66 4.13 34.64 4.75 ;
        RECT 20.285 3.98 29.025 4.745 ;
        RECT 5.025 4.135 19.535 4.745 ;
        RECT 17.4 4.13 19.38 4.75 ;
        RECT 5.025 3.98 13.765 4.745 ;
        RECT 3.45 6.655 3.74 6.885 ;
        RECT 3.28 6.685 3.74 6.855 ;
      LAYER mcon ;
        RECT 3.51 6.685 3.68 6.855 ;
        RECT 3.82 4.545 3.99 4.715 ;
        RECT 5.17 4.135 5.34 4.305 ;
        RECT 5.63 4.135 5.8 4.305 ;
        RECT 6.09 4.135 6.26 4.305 ;
        RECT 6.55 4.135 6.72 4.305 ;
        RECT 7.01 4.135 7.18 4.305 ;
        RECT 7.47 4.135 7.64 4.305 ;
        RECT 7.93 4.135 8.1 4.305 ;
        RECT 8.39 4.135 8.56 4.305 ;
        RECT 8.85 4.135 9.02 4.305 ;
        RECT 9.31 4.135 9.48 4.305 ;
        RECT 9.77 4.135 9.94 4.305 ;
        RECT 10.23 4.135 10.4 4.305 ;
        RECT 10.69 4.135 10.86 4.305 ;
        RECT 11.15 4.135 11.32 4.305 ;
        RECT 11.315 4.545 11.485 4.715 ;
        RECT 11.61 4.135 11.78 4.305 ;
        RECT 12.07 4.135 12.24 4.305 ;
        RECT 12.53 4.135 12.7 4.305 ;
        RECT 12.99 4.135 13.16 4.305 ;
        RECT 13.45 4.135 13.62 4.305 ;
        RECT 16.95 4.545 17.12 4.715 ;
        RECT 16.95 4.165 17.12 4.335 ;
        RECT 17.65 4.55 17.82 4.72 ;
        RECT 17.65 4.16 17.82 4.33 ;
        RECT 18.64 4.55 18.81 4.72 ;
        RECT 18.64 4.16 18.81 4.33 ;
        RECT 20.43 4.135 20.6 4.305 ;
        RECT 20.89 4.135 21.06 4.305 ;
        RECT 21.35 4.135 21.52 4.305 ;
        RECT 21.81 4.135 21.98 4.305 ;
        RECT 22.27 4.135 22.44 4.305 ;
        RECT 22.73 4.135 22.9 4.305 ;
        RECT 23.19 4.135 23.36 4.305 ;
        RECT 23.65 4.135 23.82 4.305 ;
        RECT 24.11 4.135 24.28 4.305 ;
        RECT 24.57 4.135 24.74 4.305 ;
        RECT 25.03 4.135 25.2 4.305 ;
        RECT 25.49 4.135 25.66 4.305 ;
        RECT 25.95 4.135 26.12 4.305 ;
        RECT 26.41 4.135 26.58 4.305 ;
        RECT 26.575 4.545 26.745 4.715 ;
        RECT 26.87 4.135 27.04 4.305 ;
        RECT 27.33 4.135 27.5 4.305 ;
        RECT 27.79 4.135 27.96 4.305 ;
        RECT 28.25 4.135 28.42 4.305 ;
        RECT 28.71 4.135 28.88 4.305 ;
        RECT 32.21 4.545 32.38 4.715 ;
        RECT 32.21 4.165 32.38 4.335 ;
        RECT 32.91 4.55 33.08 4.72 ;
        RECT 32.91 4.16 33.08 4.33 ;
        RECT 33.9 4.55 34.07 4.72 ;
        RECT 33.9 4.16 34.07 4.33 ;
        RECT 35.69 4.135 35.86 4.305 ;
        RECT 36.15 4.135 36.32 4.305 ;
        RECT 36.61 4.135 36.78 4.305 ;
        RECT 37.07 4.135 37.24 4.305 ;
        RECT 37.53 4.135 37.7 4.305 ;
        RECT 37.99 4.135 38.16 4.305 ;
        RECT 38.45 4.135 38.62 4.305 ;
        RECT 38.91 4.135 39.08 4.305 ;
        RECT 39.37 4.135 39.54 4.305 ;
        RECT 39.83 4.135 40 4.305 ;
        RECT 40.29 4.135 40.46 4.305 ;
        RECT 40.75 4.135 40.92 4.305 ;
        RECT 41.21 4.135 41.38 4.305 ;
        RECT 41.67 4.135 41.84 4.305 ;
        RECT 41.835 4.545 42.005 4.715 ;
        RECT 42.13 4.135 42.3 4.305 ;
        RECT 42.59 4.135 42.76 4.305 ;
        RECT 43.05 4.135 43.22 4.305 ;
        RECT 43.51 4.135 43.68 4.305 ;
        RECT 43.97 4.135 44.14 4.305 ;
        RECT 47.47 4.545 47.64 4.715 ;
        RECT 47.47 4.165 47.64 4.335 ;
        RECT 48.17 4.55 48.34 4.72 ;
        RECT 48.17 4.16 48.34 4.33 ;
        RECT 49.16 4.55 49.33 4.72 ;
        RECT 49.16 4.16 49.33 4.33 ;
        RECT 50.95 4.135 51.12 4.305 ;
        RECT 51.41 4.135 51.58 4.305 ;
        RECT 51.87 4.135 52.04 4.305 ;
        RECT 52.33 4.135 52.5 4.305 ;
        RECT 52.79 4.135 52.96 4.305 ;
        RECT 53.25 4.135 53.42 4.305 ;
        RECT 53.71 4.135 53.88 4.305 ;
        RECT 54.17 4.135 54.34 4.305 ;
        RECT 54.63 4.135 54.8 4.305 ;
        RECT 55.09 4.135 55.26 4.305 ;
        RECT 55.55 4.135 55.72 4.305 ;
        RECT 56.01 4.135 56.18 4.305 ;
        RECT 56.47 4.135 56.64 4.305 ;
        RECT 56.93 4.135 57.1 4.305 ;
        RECT 57.095 4.545 57.265 4.715 ;
        RECT 57.39 4.135 57.56 4.305 ;
        RECT 57.85 4.135 58.02 4.305 ;
        RECT 58.31 4.135 58.48 4.305 ;
        RECT 58.77 4.135 58.94 4.305 ;
        RECT 59.23 4.135 59.4 4.305 ;
        RECT 62.73 4.545 62.9 4.715 ;
        RECT 62.73 4.165 62.9 4.335 ;
        RECT 63.43 4.55 63.6 4.72 ;
        RECT 63.43 4.16 63.6 4.33 ;
        RECT 64.42 4.55 64.59 4.72 ;
        RECT 64.42 4.16 64.59 4.33 ;
        RECT 66.21 4.135 66.38 4.305 ;
        RECT 66.67 4.135 66.84 4.305 ;
        RECT 67.13 4.135 67.3 4.305 ;
        RECT 67.59 4.135 67.76 4.305 ;
        RECT 68.05 4.135 68.22 4.305 ;
        RECT 68.51 4.135 68.68 4.305 ;
        RECT 68.97 4.135 69.14 4.305 ;
        RECT 69.43 4.135 69.6 4.305 ;
        RECT 69.89 4.135 70.06 4.305 ;
        RECT 70.35 4.135 70.52 4.305 ;
        RECT 70.81 4.135 70.98 4.305 ;
        RECT 71.27 4.135 71.44 4.305 ;
        RECT 71.73 4.135 71.9 4.305 ;
        RECT 72.19 4.135 72.36 4.305 ;
        RECT 72.355 4.545 72.525 4.715 ;
        RECT 72.65 4.135 72.82 4.305 ;
        RECT 73.11 4.135 73.28 4.305 ;
        RECT 73.57 4.135 73.74 4.305 ;
        RECT 74.03 4.135 74.2 4.305 ;
        RECT 74.49 4.135 74.66 4.305 ;
        RECT 77.99 4.545 78.16 4.715 ;
        RECT 77.99 4.165 78.16 4.335 ;
        RECT 78.69 4.55 78.86 4.72 ;
        RECT 78.69 4.16 78.86 4.33 ;
        RECT 79.68 4.55 79.85 4.72 ;
        RECT 79.68 4.16 79.85 4.33 ;
    END
  END vccd1
  OBS
    LAYER met3 ;
      RECT 75.185 0.95 75.515 3.055 ;
      RECT 75.185 2.735 75.53 3.025 ;
      RECT 69.175 0.95 69.505 2.585 ;
      RECT 69.175 0.95 75.515 1.28 ;
      RECT 71.515 7.055 71.885 7.425 ;
      RECT 71.55 4.27 71.85 7.425 ;
      RECT 67.36 4.27 71.85 4.57 ;
      RECT 70.54 1.855 70.84 4.57 ;
      RECT 67.36 2.435 67.66 4.57 ;
      RECT 70.495 2.76 70.84 3.49 ;
      RECT 67.255 2.015 67.585 2.745 ;
      RECT 70.135 1.855 70.865 2.185 ;
      RECT 59.925 0.95 60.255 3.055 ;
      RECT 59.925 2.735 60.27 3.025 ;
      RECT 53.915 0.95 54.245 2.585 ;
      RECT 53.915 0.95 60.255 1.28 ;
      RECT 56.255 7.055 56.625 7.425 ;
      RECT 56.29 4.27 56.59 7.425 ;
      RECT 52.1 4.27 56.59 4.57 ;
      RECT 55.28 1.855 55.58 4.57 ;
      RECT 52.1 2.435 52.4 4.57 ;
      RECT 55.235 2.76 55.58 3.49 ;
      RECT 51.995 2.015 52.325 2.745 ;
      RECT 54.875 1.855 55.605 2.185 ;
      RECT 44.665 0.95 44.995 3.055 ;
      RECT 44.665 2.735 45.01 3.025 ;
      RECT 38.655 0.95 38.985 2.585 ;
      RECT 38.655 0.95 44.995 1.28 ;
      RECT 40.995 7.055 41.365 7.425 ;
      RECT 41.03 4.27 41.33 7.425 ;
      RECT 36.84 4.27 41.33 4.57 ;
      RECT 40.02 1.855 40.32 4.57 ;
      RECT 36.84 2.435 37.14 4.57 ;
      RECT 39.975 2.76 40.32 3.49 ;
      RECT 36.735 2.015 37.065 2.745 ;
      RECT 39.615 1.855 40.345 2.185 ;
      RECT 29.405 0.95 29.735 3.055 ;
      RECT 29.405 2.735 29.75 3.025 ;
      RECT 23.395 0.95 23.725 2.585 ;
      RECT 23.395 0.95 29.735 1.28 ;
      RECT 25.735 7.055 26.105 7.425 ;
      RECT 25.77 4.27 26.07 7.425 ;
      RECT 21.58 4.27 26.07 4.57 ;
      RECT 24.76 1.855 25.06 4.57 ;
      RECT 21.58 2.435 21.88 4.57 ;
      RECT 24.715 2.76 25.06 3.49 ;
      RECT 21.475 2.015 21.805 2.745 ;
      RECT 24.355 1.855 25.085 2.185 ;
      RECT 14.145 0.95 14.475 3.055 ;
      RECT 14.145 2.735 14.49 3.025 ;
      RECT 8.135 0.95 8.465 2.585 ;
      RECT 8.135 0.95 14.475 1.28 ;
      RECT 10.475 7.055 10.845 7.425 ;
      RECT 10.51 4.27 10.81 7.425 ;
      RECT 6.32 4.27 10.81 4.57 ;
      RECT 9.5 1.855 9.8 4.57 ;
      RECT 6.32 2.435 6.62 4.57 ;
      RECT 9.455 2.76 9.8 3.49 ;
      RECT 6.215 2.015 6.545 2.745 ;
      RECT 9.095 1.855 9.825 2.185 ;
      RECT 73.615 2.015 73.945 2.745 ;
      RECT 72.415 2.88 72.745 3.61 ;
      RECT 71.575 1.855 72.305 2.185 ;
      RECT 67.975 2.015 68.305 2.745 ;
      RECT 58.355 2.015 58.685 2.745 ;
      RECT 57.155 2.88 57.485 3.61 ;
      RECT 56.315 1.855 57.045 2.185 ;
      RECT 52.715 2.015 53.045 2.745 ;
      RECT 43.095 2.015 43.425 2.745 ;
      RECT 41.895 2.88 42.225 3.61 ;
      RECT 41.055 1.855 41.785 2.185 ;
      RECT 37.455 2.015 37.785 2.745 ;
      RECT 27.835 2.015 28.165 2.745 ;
      RECT 26.635 2.88 26.965 3.61 ;
      RECT 25.795 1.855 26.525 2.185 ;
      RECT 22.195 2.015 22.525 2.745 ;
      RECT 12.575 2.015 12.905 2.745 ;
      RECT 11.375 2.88 11.705 3.61 ;
      RECT 10.535 1.855 11.265 2.185 ;
      RECT 6.935 2.015 7.265 2.745 ;
    LAYER via2 ;
      RECT 75.285 2.78 75.485 2.98 ;
      RECT 73.68 2.48 73.88 2.68 ;
      RECT 72.48 3.04 72.68 3.24 ;
      RECT 71.64 1.92 71.84 2.12 ;
      RECT 71.6 7.14 71.8 7.34 ;
      RECT 70.56 2.825 70.76 3.025 ;
      RECT 70.2 1.92 70.4 2.12 ;
      RECT 69.24 1.92 69.44 2.12 ;
      RECT 68.04 2.48 68.24 2.68 ;
      RECT 67.32 2.48 67.52 2.68 ;
      RECT 60.025 2.78 60.225 2.98 ;
      RECT 58.42 2.48 58.62 2.68 ;
      RECT 57.22 3.04 57.42 3.24 ;
      RECT 56.38 1.92 56.58 2.12 ;
      RECT 56.34 7.14 56.54 7.34 ;
      RECT 55.3 2.825 55.5 3.025 ;
      RECT 54.94 1.92 55.14 2.12 ;
      RECT 53.98 1.92 54.18 2.12 ;
      RECT 52.78 2.48 52.98 2.68 ;
      RECT 52.06 2.48 52.26 2.68 ;
      RECT 44.765 2.78 44.965 2.98 ;
      RECT 43.16 2.48 43.36 2.68 ;
      RECT 41.96 3.04 42.16 3.24 ;
      RECT 41.12 1.92 41.32 2.12 ;
      RECT 41.08 7.14 41.28 7.34 ;
      RECT 40.04 2.825 40.24 3.025 ;
      RECT 39.68 1.92 39.88 2.12 ;
      RECT 38.72 1.92 38.92 2.12 ;
      RECT 37.52 2.48 37.72 2.68 ;
      RECT 36.8 2.48 37 2.68 ;
      RECT 29.505 2.78 29.705 2.98 ;
      RECT 27.9 2.48 28.1 2.68 ;
      RECT 26.7 3.04 26.9 3.24 ;
      RECT 25.86 1.92 26.06 2.12 ;
      RECT 25.82 7.14 26.02 7.34 ;
      RECT 24.78 2.825 24.98 3.025 ;
      RECT 24.42 1.92 24.62 2.12 ;
      RECT 23.46 1.92 23.66 2.12 ;
      RECT 22.26 2.48 22.46 2.68 ;
      RECT 21.54 2.48 21.74 2.68 ;
      RECT 14.245 2.78 14.445 2.98 ;
      RECT 12.64 2.48 12.84 2.68 ;
      RECT 11.44 3.04 11.64 3.24 ;
      RECT 10.6 1.92 10.8 2.12 ;
      RECT 10.56 7.14 10.76 7.34 ;
      RECT 9.52 2.825 9.72 3.025 ;
      RECT 9.16 1.92 9.36 2.12 ;
      RECT 8.2 1.92 8.4 2.12 ;
      RECT 7 2.48 7.2 2.68 ;
      RECT 6.28 2.48 6.48 2.68 ;
    LAYER met2 ;
      RECT 2.705 8.4 80.205 8.57 ;
      RECT 80.035 7.275 80.205 8.57 ;
      RECT 2.705 6.255 2.875 8.57 ;
      RECT 80.005 7.275 80.355 7.625 ;
      RECT 2.645 6.255 2.935 6.605 ;
      RECT 76.845 6.22 77.165 6.545 ;
      RECT 76.875 5.695 77.045 6.545 ;
      RECT 76.875 5.695 77.05 6.045 ;
      RECT 76.875 5.695 77.85 5.87 ;
      RECT 77.675 1.965 77.85 5.87 ;
      RECT 77.62 1.965 77.97 2.315 ;
      RECT 77.645 6.655 77.97 6.98 ;
      RECT 76.53 6.745 77.97 6.915 ;
      RECT 76.53 2.395 76.69 6.915 ;
      RECT 76.845 2.365 77.165 2.685 ;
      RECT 76.53 2.395 77.165 2.565 ;
      RECT 75.195 2.705 75.58 3.055 ;
      RECT 75.185 2.77 75.58 2.97 ;
      RECT 75.33 2.7 75.5 3.055 ;
      RECT 73.64 2.44 73.92 2.72 ;
      RECT 73.635 2.44 73.92 2.673 ;
      RECT 73.615 2.44 73.92 2.65 ;
      RECT 73.605 2.44 73.92 2.63 ;
      RECT 73.595 2.44 73.92 2.615 ;
      RECT 73.57 2.44 73.92 2.588 ;
      RECT 73.56 2.44 73.92 2.563 ;
      RECT 73.515 2.295 73.795 2.555 ;
      RECT 73.515 2.39 73.895 2.555 ;
      RECT 73.515 2.335 73.84 2.555 ;
      RECT 73.515 2.327 73.835 2.555 ;
      RECT 73.515 2.317 73.83 2.555 ;
      RECT 73.515 2.305 73.825 2.555 ;
      RECT 72.44 3 72.72 3.28 ;
      RECT 72.44 3 72.755 3.26 ;
      RECT 64.72 6.655 65.07 7.005 ;
      RECT 72.185 6.61 72.535 6.96 ;
      RECT 64.72 6.685 72.535 6.885 ;
      RECT 72.475 2.42 72.525 2.68 ;
      RECT 72.265 2.42 72.27 2.68 ;
      RECT 71.46 1.975 71.49 2.235 ;
      RECT 71.23 1.975 71.305 2.235 ;
      RECT 72.45 2.37 72.475 2.68 ;
      RECT 72.445 2.327 72.45 2.68 ;
      RECT 72.44 2.31 72.445 2.68 ;
      RECT 72.435 2.297 72.44 2.68 ;
      RECT 72.36 2.18 72.435 2.68 ;
      RECT 72.315 1.997 72.36 2.68 ;
      RECT 72.31 1.925 72.315 2.68 ;
      RECT 72.295 1.9 72.31 2.68 ;
      RECT 72.27 1.862 72.295 2.68 ;
      RECT 72.26 1.842 72.27 2.402 ;
      RECT 72.245 1.834 72.26 2.357 ;
      RECT 72.24 1.826 72.245 2.328 ;
      RECT 72.235 1.823 72.24 2.308 ;
      RECT 72.23 1.82 72.235 2.288 ;
      RECT 72.225 1.817 72.23 2.268 ;
      RECT 72.195 1.806 72.225 2.205 ;
      RECT 72.175 1.791 72.195 2.12 ;
      RECT 72.17 1.783 72.175 2.083 ;
      RECT 72.16 1.777 72.17 2.05 ;
      RECT 72.145 1.769 72.16 2.01 ;
      RECT 72.14 1.762 72.145 1.97 ;
      RECT 72.135 1.759 72.14 1.948 ;
      RECT 72.13 1.756 72.135 1.935 ;
      RECT 72.125 1.755 72.13 1.925 ;
      RECT 72.11 1.749 72.125 1.915 ;
      RECT 72.085 1.736 72.11 1.9 ;
      RECT 72.035 1.711 72.085 1.871 ;
      RECT 72.02 1.69 72.035 1.846 ;
      RECT 72.01 1.683 72.02 1.835 ;
      RECT 71.955 1.664 72.01 1.808 ;
      RECT 71.93 1.642 71.955 1.781 ;
      RECT 71.925 1.635 71.93 1.776 ;
      RECT 71.91 1.635 71.925 1.774 ;
      RECT 71.885 1.627 71.91 1.77 ;
      RECT 71.87 1.625 71.885 1.766 ;
      RECT 71.84 1.625 71.87 1.763 ;
      RECT 71.83 1.625 71.84 1.758 ;
      RECT 71.785 1.625 71.83 1.756 ;
      RECT 71.756 1.625 71.785 1.757 ;
      RECT 71.67 1.625 71.756 1.759 ;
      RECT 71.656 1.626 71.67 1.761 ;
      RECT 71.57 1.627 71.656 1.763 ;
      RECT 71.555 1.628 71.57 1.773 ;
      RECT 71.55 1.629 71.555 1.782 ;
      RECT 71.53 1.632 71.55 1.792 ;
      RECT 71.515 1.64 71.53 1.807 ;
      RECT 71.495 1.658 71.515 1.822 ;
      RECT 71.485 1.67 71.495 1.845 ;
      RECT 71.475 1.679 71.485 1.875 ;
      RECT 71.46 1.691 71.475 1.92 ;
      RECT 71.405 1.724 71.46 2.235 ;
      RECT 71.4 1.752 71.405 2.235 ;
      RECT 71.38 1.767 71.4 2.235 ;
      RECT 71.345 1.827 71.38 2.235 ;
      RECT 71.343 1.877 71.345 2.235 ;
      RECT 71.34 1.885 71.343 2.235 ;
      RECT 71.33 1.9 71.34 2.235 ;
      RECT 71.325 1.912 71.33 2.235 ;
      RECT 71.315 1.937 71.325 2.235 ;
      RECT 71.305 1.965 71.315 2.235 ;
      RECT 69.21 3.47 69.26 3.73 ;
      RECT 72.12 3.02 72.18 3.28 ;
      RECT 72.105 3.02 72.12 3.29 ;
      RECT 72.086 3.02 72.105 3.323 ;
      RECT 72 3.02 72.086 3.448 ;
      RECT 71.92 3.02 72 3.63 ;
      RECT 71.915 3.257 71.92 3.715 ;
      RECT 71.89 3.327 71.915 3.743 ;
      RECT 71.885 3.397 71.89 3.77 ;
      RECT 71.865 3.469 71.885 3.792 ;
      RECT 71.86 3.536 71.865 3.815 ;
      RECT 71.85 3.565 71.86 3.83 ;
      RECT 71.84 3.587 71.85 3.847 ;
      RECT 71.835 3.597 71.84 3.858 ;
      RECT 71.83 3.605 71.835 3.866 ;
      RECT 71.82 3.613 71.83 3.878 ;
      RECT 71.815 3.625 71.82 3.888 ;
      RECT 71.81 3.633 71.815 3.893 ;
      RECT 71.79 3.651 71.81 3.903 ;
      RECT 71.785 3.668 71.79 3.91 ;
      RECT 71.78 3.676 71.785 3.911 ;
      RECT 71.775 3.687 71.78 3.913 ;
      RECT 71.735 3.725 71.775 3.923 ;
      RECT 71.73 3.76 71.735 3.934 ;
      RECT 71.725 3.765 71.73 3.937 ;
      RECT 71.7 3.775 71.725 3.944 ;
      RECT 71.69 3.789 71.7 3.953 ;
      RECT 71.67 3.801 71.69 3.956 ;
      RECT 71.62 3.82 71.67 3.96 ;
      RECT 71.575 3.835 71.62 3.965 ;
      RECT 71.51 3.838 71.575 3.971 ;
      RECT 71.495 3.836 71.51 3.978 ;
      RECT 71.465 3.835 71.495 3.978 ;
      RECT 71.426 3.834 71.465 3.974 ;
      RECT 71.34 3.831 71.426 3.97 ;
      RECT 71.323 3.829 71.34 3.967 ;
      RECT 71.237 3.827 71.323 3.964 ;
      RECT 71.151 3.824 71.237 3.958 ;
      RECT 71.065 3.82 71.151 3.953 ;
      RECT 70.987 3.817 71.065 3.949 ;
      RECT 70.901 3.814 70.987 3.947 ;
      RECT 70.815 3.811 70.901 3.944 ;
      RECT 70.757 3.809 70.815 3.941 ;
      RECT 70.671 3.806 70.757 3.939 ;
      RECT 70.585 3.802 70.671 3.937 ;
      RECT 70.499 3.799 70.585 3.934 ;
      RECT 70.413 3.795 70.499 3.932 ;
      RECT 70.327 3.791 70.413 3.929 ;
      RECT 70.241 3.788 70.327 3.927 ;
      RECT 70.155 3.784 70.241 3.924 ;
      RECT 70.069 3.781 70.155 3.922 ;
      RECT 69.983 3.777 70.069 3.919 ;
      RECT 69.897 3.774 69.983 3.917 ;
      RECT 69.811 3.77 69.897 3.914 ;
      RECT 69.725 3.767 69.811 3.912 ;
      RECT 69.715 3.765 69.725 3.908 ;
      RECT 69.71 3.765 69.715 3.906 ;
      RECT 69.67 3.76 69.71 3.9 ;
      RECT 69.656 3.751 69.67 3.893 ;
      RECT 69.57 3.721 69.656 3.878 ;
      RECT 69.55 3.687 69.57 3.863 ;
      RECT 69.48 3.656 69.55 3.85 ;
      RECT 69.475 3.631 69.48 3.839 ;
      RECT 69.47 3.625 69.475 3.837 ;
      RECT 69.401 3.47 69.47 3.825 ;
      RECT 69.315 3.47 69.401 3.799 ;
      RECT 69.29 3.47 69.315 3.778 ;
      RECT 69.285 3.47 69.29 3.768 ;
      RECT 69.28 3.47 69.285 3.76 ;
      RECT 69.26 3.47 69.28 3.743 ;
      RECT 71.68 2.04 71.94 2.3 ;
      RECT 71.665 2.04 71.94 2.203 ;
      RECT 71.635 2.04 71.94 2.178 ;
      RECT 71.6 1.88 71.88 2.16 ;
      RECT 71.57 3.37 71.63 3.63 ;
      RECT 70.595 2.06 70.65 2.32 ;
      RECT 71.53 3.327 71.57 3.63 ;
      RECT 71.501 3.248 71.53 3.63 ;
      RECT 71.415 3.12 71.501 3.63 ;
      RECT 71.395 3 71.415 3.63 ;
      RECT 71.37 2.951 71.395 3.63 ;
      RECT 71.365 2.916 71.37 3.48 ;
      RECT 71.335 2.876 71.365 3.418 ;
      RECT 71.31 2.813 71.335 3.333 ;
      RECT 71.3 2.775 71.31 3.27 ;
      RECT 71.285 2.75 71.3 3.231 ;
      RECT 71.242 2.708 71.285 3.137 ;
      RECT 71.24 2.681 71.242 3.064 ;
      RECT 71.235 2.676 71.24 3.055 ;
      RECT 71.23 2.669 71.235 3.03 ;
      RECT 71.225 2.663 71.23 3.015 ;
      RECT 71.22 2.657 71.225 3.003 ;
      RECT 71.21 2.648 71.22 2.985 ;
      RECT 71.205 2.639 71.21 2.963 ;
      RECT 71.18 2.62 71.205 2.913 ;
      RECT 71.175 2.601 71.18 2.863 ;
      RECT 71.16 2.587 71.175 2.823 ;
      RECT 71.155 2.573 71.16 2.79 ;
      RECT 71.15 2.566 71.155 2.783 ;
      RECT 71.135 2.553 71.15 2.775 ;
      RECT 71.09 2.515 71.135 2.748 ;
      RECT 71.06 2.468 71.09 2.713 ;
      RECT 71.04 2.437 71.06 2.69 ;
      RECT 70.96 2.37 71.04 2.643 ;
      RECT 70.93 2.3 70.96 2.59 ;
      RECT 70.925 2.277 70.93 2.573 ;
      RECT 70.895 2.255 70.925 2.558 ;
      RECT 70.865 2.214 70.895 2.53 ;
      RECT 70.86 2.189 70.865 2.515 ;
      RECT 70.855 2.183 70.86 2.508 ;
      RECT 70.845 2.06 70.855 2.5 ;
      RECT 70.835 2.06 70.845 2.493 ;
      RECT 70.83 2.06 70.835 2.485 ;
      RECT 70.81 2.06 70.83 2.473 ;
      RECT 70.76 2.06 70.81 2.443 ;
      RECT 70.705 2.06 70.76 2.393 ;
      RECT 70.675 2.06 70.705 2.353 ;
      RECT 70.65 2.06 70.675 2.33 ;
      RECT 70.52 2.785 70.8 3.065 ;
      RECT 70.485 2.7 70.745 2.96 ;
      RECT 70.485 2.782 70.755 2.96 ;
      RECT 68.685 2.155 68.69 2.64 ;
      RECT 68.575 2.34 68.58 2.64 ;
      RECT 68.485 2.38 68.55 2.64 ;
      RECT 70.16 1.88 70.25 2.51 ;
      RECT 70.125 1.93 70.13 2.51 ;
      RECT 70.07 1.955 70.08 2.51 ;
      RECT 70.025 1.955 70.035 2.51 ;
      RECT 70.395 1.88 70.44 2.16 ;
      RECT 69.245 1.61 69.445 1.75 ;
      RECT 70.361 1.88 70.395 2.172 ;
      RECT 70.275 1.88 70.361 2.212 ;
      RECT 70.26 1.88 70.275 2.253 ;
      RECT 70.255 1.88 70.26 2.273 ;
      RECT 70.25 1.88 70.255 2.293 ;
      RECT 70.13 1.922 70.16 2.51 ;
      RECT 70.08 1.942 70.125 2.51 ;
      RECT 70.065 1.957 70.07 2.51 ;
      RECT 70.035 1.957 70.065 2.51 ;
      RECT 69.99 1.942 70.025 2.51 ;
      RECT 69.985 1.93 69.99 2.29 ;
      RECT 69.98 1.927 69.985 2.27 ;
      RECT 69.965 1.917 69.98 2.223 ;
      RECT 69.96 1.91 69.965 2.186 ;
      RECT 69.955 1.907 69.96 2.169 ;
      RECT 69.94 1.897 69.955 2.125 ;
      RECT 69.935 1.888 69.94 2.085 ;
      RECT 69.93 1.884 69.935 2.07 ;
      RECT 69.92 1.878 69.93 2.053 ;
      RECT 69.88 1.859 69.92 2.028 ;
      RECT 69.875 1.841 69.88 2.008 ;
      RECT 69.865 1.835 69.875 2.003 ;
      RECT 69.835 1.819 69.865 1.99 ;
      RECT 69.82 1.801 69.835 1.973 ;
      RECT 69.805 1.789 69.82 1.96 ;
      RECT 69.8 1.781 69.805 1.953 ;
      RECT 69.77 1.767 69.8 1.94 ;
      RECT 69.765 1.752 69.77 1.928 ;
      RECT 69.755 1.746 69.765 1.92 ;
      RECT 69.735 1.734 69.755 1.908 ;
      RECT 69.725 1.722 69.735 1.895 ;
      RECT 69.695 1.706 69.725 1.88 ;
      RECT 69.675 1.686 69.695 1.863 ;
      RECT 69.67 1.676 69.675 1.853 ;
      RECT 69.645 1.664 69.67 1.84 ;
      RECT 69.64 1.652 69.645 1.828 ;
      RECT 69.635 1.647 69.64 1.824 ;
      RECT 69.62 1.64 69.635 1.816 ;
      RECT 69.61 1.627 69.62 1.806 ;
      RECT 69.605 1.625 69.61 1.8 ;
      RECT 69.58 1.618 69.605 1.789 ;
      RECT 69.575 1.611 69.58 1.778 ;
      RECT 69.55 1.61 69.575 1.765 ;
      RECT 69.531 1.61 69.55 1.755 ;
      RECT 69.445 1.61 69.531 1.752 ;
      RECT 69.215 1.61 69.245 1.755 ;
      RECT 69.175 1.617 69.215 1.768 ;
      RECT 69.15 1.627 69.175 1.781 ;
      RECT 69.135 1.636 69.15 1.791 ;
      RECT 69.105 1.641 69.135 1.81 ;
      RECT 69.1 1.647 69.105 1.828 ;
      RECT 69.08 1.657 69.1 1.843 ;
      RECT 69.07 1.67 69.08 1.863 ;
      RECT 69.055 1.682 69.07 1.88 ;
      RECT 69.05 1.692 69.055 1.89 ;
      RECT 69.045 1.697 69.05 1.895 ;
      RECT 69.035 1.705 69.045 1.908 ;
      RECT 68.985 1.737 69.035 1.945 ;
      RECT 68.97 1.772 68.985 1.986 ;
      RECT 68.965 1.782 68.97 2.001 ;
      RECT 68.96 1.787 68.965 2.008 ;
      RECT 68.935 1.803 68.96 2.028 ;
      RECT 68.92 1.824 68.935 2.053 ;
      RECT 68.895 1.845 68.92 2.078 ;
      RECT 68.885 1.864 68.895 2.101 ;
      RECT 68.86 1.882 68.885 2.124 ;
      RECT 68.845 1.902 68.86 2.148 ;
      RECT 68.84 1.912 68.845 2.16 ;
      RECT 68.825 1.924 68.84 2.18 ;
      RECT 68.815 1.939 68.825 2.22 ;
      RECT 68.81 1.947 68.815 2.248 ;
      RECT 68.8 1.957 68.81 2.268 ;
      RECT 68.795 1.97 68.8 2.293 ;
      RECT 68.79 1.983 68.795 2.313 ;
      RECT 68.785 1.989 68.79 2.335 ;
      RECT 68.775 1.998 68.785 2.355 ;
      RECT 68.77 2.018 68.775 2.378 ;
      RECT 68.765 2.024 68.77 2.398 ;
      RECT 68.76 2.031 68.765 2.42 ;
      RECT 68.755 2.042 68.76 2.433 ;
      RECT 68.745 2.052 68.755 2.458 ;
      RECT 68.725 2.077 68.745 2.64 ;
      RECT 68.695 2.117 68.725 2.64 ;
      RECT 68.69 2.147 68.695 2.64 ;
      RECT 68.665 2.175 68.685 2.64 ;
      RECT 68.635 2.22 68.665 2.64 ;
      RECT 68.63 2.247 68.635 2.64 ;
      RECT 68.61 2.265 68.63 2.64 ;
      RECT 68.6 2.29 68.61 2.64 ;
      RECT 68.595 2.302 68.6 2.64 ;
      RECT 68.58 2.325 68.595 2.64 ;
      RECT 68.56 2.352 68.575 2.64 ;
      RECT 68.55 2.375 68.56 2.64 ;
      RECT 70.34 3.26 70.42 3.52 ;
      RECT 69.575 2.48 69.645 2.74 ;
      RECT 70.306 3.227 70.34 3.52 ;
      RECT 70.22 3.13 70.306 3.52 ;
      RECT 70.2 3.042 70.22 3.52 ;
      RECT 70.19 3.012 70.2 3.52 ;
      RECT 70.18 2.992 70.19 3.52 ;
      RECT 70.16 2.979 70.18 3.52 ;
      RECT 70.145 2.969 70.16 3.348 ;
      RECT 70.14 2.962 70.145 3.303 ;
      RECT 70.13 2.956 70.14 3.293 ;
      RECT 70.12 2.948 70.13 3.275 ;
      RECT 70.115 2.942 70.12 3.263 ;
      RECT 70.105 2.937 70.115 3.25 ;
      RECT 70.085 2.927 70.105 3.223 ;
      RECT 70.045 2.906 70.085 3.175 ;
      RECT 70.03 2.887 70.045 3.133 ;
      RECT 70.005 2.873 70.03 3.103 ;
      RECT 69.995 2.861 70.005 3.07 ;
      RECT 69.99 2.856 69.995 3.06 ;
      RECT 69.96 2.842 69.99 3.04 ;
      RECT 69.95 2.826 69.96 3.013 ;
      RECT 69.945 2.821 69.95 3.003 ;
      RECT 69.92 2.812 69.945 2.983 ;
      RECT 69.91 2.8 69.92 2.963 ;
      RECT 69.84 2.768 69.91 2.938 ;
      RECT 69.835 2.737 69.84 2.915 ;
      RECT 69.786 2.48 69.835 2.898 ;
      RECT 69.7 2.48 69.786 2.857 ;
      RECT 69.645 2.48 69.7 2.785 ;
      RECT 69.735 3.265 69.895 3.525 ;
      RECT 69.26 1.88 69.31 2.565 ;
      RECT 69.05 2.305 69.085 2.565 ;
      RECT 69.365 1.88 69.37 2.34 ;
      RECT 69.455 1.88 69.48 2.16 ;
      RECT 69.73 3.262 69.735 3.525 ;
      RECT 69.695 3.25 69.73 3.525 ;
      RECT 69.635 3.223 69.695 3.525 ;
      RECT 69.63 3.206 69.635 3.379 ;
      RECT 69.625 3.203 69.63 3.366 ;
      RECT 69.605 3.196 69.625 3.353 ;
      RECT 69.57 3.179 69.605 3.335 ;
      RECT 69.53 3.158 69.57 3.315 ;
      RECT 69.525 3.146 69.53 3.303 ;
      RECT 69.485 3.132 69.525 3.289 ;
      RECT 69.465 3.115 69.485 3.271 ;
      RECT 69.455 3.107 69.465 3.263 ;
      RECT 69.44 1.88 69.455 2.178 ;
      RECT 69.425 3.097 69.455 3.25 ;
      RECT 69.41 1.88 69.44 2.223 ;
      RECT 69.415 3.087 69.425 3.237 ;
      RECT 69.385 3.072 69.415 3.224 ;
      RECT 69.37 1.88 69.41 2.29 ;
      RECT 69.37 3.04 69.385 3.21 ;
      RECT 69.365 3.012 69.37 3.204 ;
      RECT 69.36 1.88 69.365 2.345 ;
      RECT 69.35 2.982 69.365 3.198 ;
      RECT 69.355 1.88 69.36 2.358 ;
      RECT 69.345 1.88 69.355 2.378 ;
      RECT 69.31 2.895 69.35 3.183 ;
      RECT 69.31 1.88 69.345 2.418 ;
      RECT 69.305 2.827 69.31 3.171 ;
      RECT 69.29 2.782 69.305 3.166 ;
      RECT 69.285 2.72 69.29 3.161 ;
      RECT 69.26 2.627 69.285 3.154 ;
      RECT 69.255 1.88 69.26 3.146 ;
      RECT 69.24 1.88 69.255 3.133 ;
      RECT 69.22 1.88 69.24 3.09 ;
      RECT 69.21 1.88 69.22 3.04 ;
      RECT 69.205 1.88 69.21 3.013 ;
      RECT 69.2 1.88 69.205 2.991 ;
      RECT 69.195 2.106 69.2 2.974 ;
      RECT 69.19 2.128 69.195 2.952 ;
      RECT 69.185 2.17 69.19 2.935 ;
      RECT 69.155 2.22 69.185 2.879 ;
      RECT 69.15 2.247 69.155 2.821 ;
      RECT 69.135 2.265 69.15 2.785 ;
      RECT 69.13 2.283 69.135 2.749 ;
      RECT 69.124 2.29 69.13 2.73 ;
      RECT 69.12 2.297 69.124 2.713 ;
      RECT 69.115 2.302 69.12 2.682 ;
      RECT 69.105 2.305 69.115 2.657 ;
      RECT 69.095 2.305 69.105 2.623 ;
      RECT 69.09 2.305 69.095 2.6 ;
      RECT 69.085 2.305 69.09 2.58 ;
      RECT 68 2.44 68.28 2.72 ;
      RECT 68 2.44 68.3 2.615 ;
      RECT 68.09 2.33 68.35 2.59 ;
      RECT 68.055 2.425 68.35 2.59 ;
      RECT 68.18 0.945 68.345 2.59 ;
      RECT 68.08 0.945 68.45 1.315 ;
      RECT 67.705 3.47 67.965 3.73 ;
      RECT 67.725 3.397 67.905 3.73 ;
      RECT 67.725 3.14 67.9 3.73 ;
      RECT 67.725 2.932 67.89 3.73 ;
      RECT 67.73 2.85 67.89 3.73 ;
      RECT 67.73 2.615 67.88 3.73 ;
      RECT 67.73 2.462 67.875 3.73 ;
      RECT 67.735 2.447 67.875 3.73 ;
      RECT 67.785 2.162 67.875 3.73 ;
      RECT 67.74 2.397 67.875 3.73 ;
      RECT 67.77 2.215 67.875 3.73 ;
      RECT 67.755 2.327 67.875 3.73 ;
      RECT 67.76 2.285 67.875 3.73 ;
      RECT 67.755 2.327 67.89 2.39 ;
      RECT 67.79 1.915 67.895 2.335 ;
      RECT 67.79 1.915 67.91 2.318 ;
      RECT 67.79 1.915 67.945 2.28 ;
      RECT 67.785 2.162 67.995 2.213 ;
      RECT 67.79 1.915 68.05 2.175 ;
      RECT 67.05 2.62 67.31 2.88 ;
      RECT 67.05 2.62 67.32 2.838 ;
      RECT 67.05 2.62 67.406 2.809 ;
      RECT 67.05 2.62 67.475 2.761 ;
      RECT 67.05 2.62 67.51 2.73 ;
      RECT 67.28 2.44 67.56 2.72 ;
      RECT 67.115 2.605 67.56 2.72 ;
      RECT 67.205 2.482 67.31 2.88 ;
      RECT 67.135 2.545 67.56 2.72 ;
      RECT 61.585 6.22 61.905 6.545 ;
      RECT 61.615 5.695 61.785 6.545 ;
      RECT 61.615 5.695 61.79 6.045 ;
      RECT 61.615 5.695 62.59 5.87 ;
      RECT 62.415 1.965 62.59 5.87 ;
      RECT 62.36 1.965 62.71 2.315 ;
      RECT 62.385 6.655 62.71 6.98 ;
      RECT 61.27 6.745 62.71 6.915 ;
      RECT 61.27 2.395 61.43 6.915 ;
      RECT 61.585 2.365 61.905 2.685 ;
      RECT 61.27 2.395 61.905 2.565 ;
      RECT 59.935 2.705 60.32 3.055 ;
      RECT 59.925 2.77 60.32 2.97 ;
      RECT 60.07 2.7 60.24 3.055 ;
      RECT 58.38 2.44 58.66 2.72 ;
      RECT 58.375 2.44 58.66 2.673 ;
      RECT 58.355 2.44 58.66 2.65 ;
      RECT 58.345 2.44 58.66 2.63 ;
      RECT 58.335 2.44 58.66 2.615 ;
      RECT 58.31 2.44 58.66 2.588 ;
      RECT 58.3 2.44 58.66 2.563 ;
      RECT 58.255 2.295 58.535 2.555 ;
      RECT 58.255 2.39 58.635 2.555 ;
      RECT 58.255 2.335 58.58 2.555 ;
      RECT 58.255 2.327 58.575 2.555 ;
      RECT 58.255 2.317 58.57 2.555 ;
      RECT 58.255 2.305 58.565 2.555 ;
      RECT 57.18 3 57.46 3.28 ;
      RECT 57.18 3 57.495 3.26 ;
      RECT 49.46 6.655 49.81 7.005 ;
      RECT 56.925 6.61 57.275 6.96 ;
      RECT 49.46 6.685 57.275 6.885 ;
      RECT 57.215 2.42 57.265 2.68 ;
      RECT 57.005 2.42 57.01 2.68 ;
      RECT 56.2 1.975 56.23 2.235 ;
      RECT 55.97 1.975 56.045 2.235 ;
      RECT 57.19 2.37 57.215 2.68 ;
      RECT 57.185 2.327 57.19 2.68 ;
      RECT 57.18 2.31 57.185 2.68 ;
      RECT 57.175 2.297 57.18 2.68 ;
      RECT 57.1 2.18 57.175 2.68 ;
      RECT 57.055 1.997 57.1 2.68 ;
      RECT 57.05 1.925 57.055 2.68 ;
      RECT 57.035 1.9 57.05 2.68 ;
      RECT 57.01 1.862 57.035 2.68 ;
      RECT 57 1.842 57.01 2.402 ;
      RECT 56.985 1.834 57 2.357 ;
      RECT 56.98 1.826 56.985 2.328 ;
      RECT 56.975 1.823 56.98 2.308 ;
      RECT 56.97 1.82 56.975 2.288 ;
      RECT 56.965 1.817 56.97 2.268 ;
      RECT 56.935 1.806 56.965 2.205 ;
      RECT 56.915 1.791 56.935 2.12 ;
      RECT 56.91 1.783 56.915 2.083 ;
      RECT 56.9 1.777 56.91 2.05 ;
      RECT 56.885 1.769 56.9 2.01 ;
      RECT 56.88 1.762 56.885 1.97 ;
      RECT 56.875 1.759 56.88 1.948 ;
      RECT 56.87 1.756 56.875 1.935 ;
      RECT 56.865 1.755 56.87 1.925 ;
      RECT 56.85 1.749 56.865 1.915 ;
      RECT 56.825 1.736 56.85 1.9 ;
      RECT 56.775 1.711 56.825 1.871 ;
      RECT 56.76 1.69 56.775 1.846 ;
      RECT 56.75 1.683 56.76 1.835 ;
      RECT 56.695 1.664 56.75 1.808 ;
      RECT 56.67 1.642 56.695 1.781 ;
      RECT 56.665 1.635 56.67 1.776 ;
      RECT 56.65 1.635 56.665 1.774 ;
      RECT 56.625 1.627 56.65 1.77 ;
      RECT 56.61 1.625 56.625 1.766 ;
      RECT 56.58 1.625 56.61 1.763 ;
      RECT 56.57 1.625 56.58 1.758 ;
      RECT 56.525 1.625 56.57 1.756 ;
      RECT 56.496 1.625 56.525 1.757 ;
      RECT 56.41 1.625 56.496 1.759 ;
      RECT 56.396 1.626 56.41 1.761 ;
      RECT 56.31 1.627 56.396 1.763 ;
      RECT 56.295 1.628 56.31 1.773 ;
      RECT 56.29 1.629 56.295 1.782 ;
      RECT 56.27 1.632 56.29 1.792 ;
      RECT 56.255 1.64 56.27 1.807 ;
      RECT 56.235 1.658 56.255 1.822 ;
      RECT 56.225 1.67 56.235 1.845 ;
      RECT 56.215 1.679 56.225 1.875 ;
      RECT 56.2 1.691 56.215 1.92 ;
      RECT 56.145 1.724 56.2 2.235 ;
      RECT 56.14 1.752 56.145 2.235 ;
      RECT 56.12 1.767 56.14 2.235 ;
      RECT 56.085 1.827 56.12 2.235 ;
      RECT 56.083 1.877 56.085 2.235 ;
      RECT 56.08 1.885 56.083 2.235 ;
      RECT 56.07 1.9 56.08 2.235 ;
      RECT 56.065 1.912 56.07 2.235 ;
      RECT 56.055 1.937 56.065 2.235 ;
      RECT 56.045 1.965 56.055 2.235 ;
      RECT 53.95 3.47 54 3.73 ;
      RECT 56.86 3.02 56.92 3.28 ;
      RECT 56.845 3.02 56.86 3.29 ;
      RECT 56.826 3.02 56.845 3.323 ;
      RECT 56.74 3.02 56.826 3.448 ;
      RECT 56.66 3.02 56.74 3.63 ;
      RECT 56.655 3.257 56.66 3.715 ;
      RECT 56.63 3.327 56.655 3.743 ;
      RECT 56.625 3.397 56.63 3.77 ;
      RECT 56.605 3.469 56.625 3.792 ;
      RECT 56.6 3.536 56.605 3.815 ;
      RECT 56.59 3.565 56.6 3.83 ;
      RECT 56.58 3.587 56.59 3.847 ;
      RECT 56.575 3.597 56.58 3.858 ;
      RECT 56.57 3.605 56.575 3.866 ;
      RECT 56.56 3.613 56.57 3.878 ;
      RECT 56.555 3.625 56.56 3.888 ;
      RECT 56.55 3.633 56.555 3.893 ;
      RECT 56.53 3.651 56.55 3.903 ;
      RECT 56.525 3.668 56.53 3.91 ;
      RECT 56.52 3.676 56.525 3.911 ;
      RECT 56.515 3.687 56.52 3.913 ;
      RECT 56.475 3.725 56.515 3.923 ;
      RECT 56.47 3.76 56.475 3.934 ;
      RECT 56.465 3.765 56.47 3.937 ;
      RECT 56.44 3.775 56.465 3.944 ;
      RECT 56.43 3.789 56.44 3.953 ;
      RECT 56.41 3.801 56.43 3.956 ;
      RECT 56.36 3.82 56.41 3.96 ;
      RECT 56.315 3.835 56.36 3.965 ;
      RECT 56.25 3.838 56.315 3.971 ;
      RECT 56.235 3.836 56.25 3.978 ;
      RECT 56.205 3.835 56.235 3.978 ;
      RECT 56.166 3.834 56.205 3.974 ;
      RECT 56.08 3.831 56.166 3.97 ;
      RECT 56.063 3.829 56.08 3.967 ;
      RECT 55.977 3.827 56.063 3.964 ;
      RECT 55.891 3.824 55.977 3.958 ;
      RECT 55.805 3.82 55.891 3.953 ;
      RECT 55.727 3.817 55.805 3.949 ;
      RECT 55.641 3.814 55.727 3.947 ;
      RECT 55.555 3.811 55.641 3.944 ;
      RECT 55.497 3.809 55.555 3.941 ;
      RECT 55.411 3.806 55.497 3.939 ;
      RECT 55.325 3.802 55.411 3.937 ;
      RECT 55.239 3.799 55.325 3.934 ;
      RECT 55.153 3.795 55.239 3.932 ;
      RECT 55.067 3.791 55.153 3.929 ;
      RECT 54.981 3.788 55.067 3.927 ;
      RECT 54.895 3.784 54.981 3.924 ;
      RECT 54.809 3.781 54.895 3.922 ;
      RECT 54.723 3.777 54.809 3.919 ;
      RECT 54.637 3.774 54.723 3.917 ;
      RECT 54.551 3.77 54.637 3.914 ;
      RECT 54.465 3.767 54.551 3.912 ;
      RECT 54.455 3.765 54.465 3.908 ;
      RECT 54.45 3.765 54.455 3.906 ;
      RECT 54.41 3.76 54.45 3.9 ;
      RECT 54.396 3.751 54.41 3.893 ;
      RECT 54.31 3.721 54.396 3.878 ;
      RECT 54.29 3.687 54.31 3.863 ;
      RECT 54.22 3.656 54.29 3.85 ;
      RECT 54.215 3.631 54.22 3.839 ;
      RECT 54.21 3.625 54.215 3.837 ;
      RECT 54.141 3.47 54.21 3.825 ;
      RECT 54.055 3.47 54.141 3.799 ;
      RECT 54.03 3.47 54.055 3.778 ;
      RECT 54.025 3.47 54.03 3.768 ;
      RECT 54.02 3.47 54.025 3.76 ;
      RECT 54 3.47 54.02 3.743 ;
      RECT 56.42 2.04 56.68 2.3 ;
      RECT 56.405 2.04 56.68 2.203 ;
      RECT 56.375 2.04 56.68 2.178 ;
      RECT 56.34 1.88 56.62 2.16 ;
      RECT 56.31 3.37 56.37 3.63 ;
      RECT 55.335 2.06 55.39 2.32 ;
      RECT 56.27 3.327 56.31 3.63 ;
      RECT 56.241 3.248 56.27 3.63 ;
      RECT 56.155 3.12 56.241 3.63 ;
      RECT 56.135 3 56.155 3.63 ;
      RECT 56.11 2.951 56.135 3.63 ;
      RECT 56.105 2.916 56.11 3.48 ;
      RECT 56.075 2.876 56.105 3.418 ;
      RECT 56.05 2.813 56.075 3.333 ;
      RECT 56.04 2.775 56.05 3.27 ;
      RECT 56.025 2.75 56.04 3.231 ;
      RECT 55.982 2.708 56.025 3.137 ;
      RECT 55.98 2.681 55.982 3.064 ;
      RECT 55.975 2.676 55.98 3.055 ;
      RECT 55.97 2.669 55.975 3.03 ;
      RECT 55.965 2.663 55.97 3.015 ;
      RECT 55.96 2.657 55.965 3.003 ;
      RECT 55.95 2.648 55.96 2.985 ;
      RECT 55.945 2.639 55.95 2.963 ;
      RECT 55.92 2.62 55.945 2.913 ;
      RECT 55.915 2.601 55.92 2.863 ;
      RECT 55.9 2.587 55.915 2.823 ;
      RECT 55.895 2.573 55.9 2.79 ;
      RECT 55.89 2.566 55.895 2.783 ;
      RECT 55.875 2.553 55.89 2.775 ;
      RECT 55.83 2.515 55.875 2.748 ;
      RECT 55.8 2.468 55.83 2.713 ;
      RECT 55.78 2.437 55.8 2.69 ;
      RECT 55.7 2.37 55.78 2.643 ;
      RECT 55.67 2.3 55.7 2.59 ;
      RECT 55.665 2.277 55.67 2.573 ;
      RECT 55.635 2.255 55.665 2.558 ;
      RECT 55.605 2.214 55.635 2.53 ;
      RECT 55.6 2.189 55.605 2.515 ;
      RECT 55.595 2.183 55.6 2.508 ;
      RECT 55.585 2.06 55.595 2.5 ;
      RECT 55.575 2.06 55.585 2.493 ;
      RECT 55.57 2.06 55.575 2.485 ;
      RECT 55.55 2.06 55.57 2.473 ;
      RECT 55.5 2.06 55.55 2.443 ;
      RECT 55.445 2.06 55.5 2.393 ;
      RECT 55.415 2.06 55.445 2.353 ;
      RECT 55.39 2.06 55.415 2.33 ;
      RECT 55.26 2.785 55.54 3.065 ;
      RECT 55.225 2.7 55.485 2.96 ;
      RECT 55.225 2.782 55.495 2.96 ;
      RECT 53.425 2.155 53.43 2.64 ;
      RECT 53.315 2.34 53.32 2.64 ;
      RECT 53.225 2.38 53.29 2.64 ;
      RECT 54.9 1.88 54.99 2.51 ;
      RECT 54.865 1.93 54.87 2.51 ;
      RECT 54.81 1.955 54.82 2.51 ;
      RECT 54.765 1.955 54.775 2.51 ;
      RECT 55.135 1.88 55.18 2.16 ;
      RECT 53.985 1.61 54.185 1.75 ;
      RECT 55.101 1.88 55.135 2.172 ;
      RECT 55.015 1.88 55.101 2.212 ;
      RECT 55 1.88 55.015 2.253 ;
      RECT 54.995 1.88 55 2.273 ;
      RECT 54.99 1.88 54.995 2.293 ;
      RECT 54.87 1.922 54.9 2.51 ;
      RECT 54.82 1.942 54.865 2.51 ;
      RECT 54.805 1.957 54.81 2.51 ;
      RECT 54.775 1.957 54.805 2.51 ;
      RECT 54.73 1.942 54.765 2.51 ;
      RECT 54.725 1.93 54.73 2.29 ;
      RECT 54.72 1.927 54.725 2.27 ;
      RECT 54.705 1.917 54.72 2.223 ;
      RECT 54.7 1.91 54.705 2.186 ;
      RECT 54.695 1.907 54.7 2.169 ;
      RECT 54.68 1.897 54.695 2.125 ;
      RECT 54.675 1.888 54.68 2.085 ;
      RECT 54.67 1.884 54.675 2.07 ;
      RECT 54.66 1.878 54.67 2.053 ;
      RECT 54.62 1.859 54.66 2.028 ;
      RECT 54.615 1.841 54.62 2.008 ;
      RECT 54.605 1.835 54.615 2.003 ;
      RECT 54.575 1.819 54.605 1.99 ;
      RECT 54.56 1.801 54.575 1.973 ;
      RECT 54.545 1.789 54.56 1.96 ;
      RECT 54.54 1.781 54.545 1.953 ;
      RECT 54.51 1.767 54.54 1.94 ;
      RECT 54.505 1.752 54.51 1.928 ;
      RECT 54.495 1.746 54.505 1.92 ;
      RECT 54.475 1.734 54.495 1.908 ;
      RECT 54.465 1.722 54.475 1.895 ;
      RECT 54.435 1.706 54.465 1.88 ;
      RECT 54.415 1.686 54.435 1.863 ;
      RECT 54.41 1.676 54.415 1.853 ;
      RECT 54.385 1.664 54.41 1.84 ;
      RECT 54.38 1.652 54.385 1.828 ;
      RECT 54.375 1.647 54.38 1.824 ;
      RECT 54.36 1.64 54.375 1.816 ;
      RECT 54.35 1.627 54.36 1.806 ;
      RECT 54.345 1.625 54.35 1.8 ;
      RECT 54.32 1.618 54.345 1.789 ;
      RECT 54.315 1.611 54.32 1.778 ;
      RECT 54.29 1.61 54.315 1.765 ;
      RECT 54.271 1.61 54.29 1.755 ;
      RECT 54.185 1.61 54.271 1.752 ;
      RECT 53.955 1.61 53.985 1.755 ;
      RECT 53.915 1.617 53.955 1.768 ;
      RECT 53.89 1.627 53.915 1.781 ;
      RECT 53.875 1.636 53.89 1.791 ;
      RECT 53.845 1.641 53.875 1.81 ;
      RECT 53.84 1.647 53.845 1.828 ;
      RECT 53.82 1.657 53.84 1.843 ;
      RECT 53.81 1.67 53.82 1.863 ;
      RECT 53.795 1.682 53.81 1.88 ;
      RECT 53.79 1.692 53.795 1.89 ;
      RECT 53.785 1.697 53.79 1.895 ;
      RECT 53.775 1.705 53.785 1.908 ;
      RECT 53.725 1.737 53.775 1.945 ;
      RECT 53.71 1.772 53.725 1.986 ;
      RECT 53.705 1.782 53.71 2.001 ;
      RECT 53.7 1.787 53.705 2.008 ;
      RECT 53.675 1.803 53.7 2.028 ;
      RECT 53.66 1.824 53.675 2.053 ;
      RECT 53.635 1.845 53.66 2.078 ;
      RECT 53.625 1.864 53.635 2.101 ;
      RECT 53.6 1.882 53.625 2.124 ;
      RECT 53.585 1.902 53.6 2.148 ;
      RECT 53.58 1.912 53.585 2.16 ;
      RECT 53.565 1.924 53.58 2.18 ;
      RECT 53.555 1.939 53.565 2.22 ;
      RECT 53.55 1.947 53.555 2.248 ;
      RECT 53.54 1.957 53.55 2.268 ;
      RECT 53.535 1.97 53.54 2.293 ;
      RECT 53.53 1.983 53.535 2.313 ;
      RECT 53.525 1.989 53.53 2.335 ;
      RECT 53.515 1.998 53.525 2.355 ;
      RECT 53.51 2.018 53.515 2.378 ;
      RECT 53.505 2.024 53.51 2.398 ;
      RECT 53.5 2.031 53.505 2.42 ;
      RECT 53.495 2.042 53.5 2.433 ;
      RECT 53.485 2.052 53.495 2.458 ;
      RECT 53.465 2.077 53.485 2.64 ;
      RECT 53.435 2.117 53.465 2.64 ;
      RECT 53.43 2.147 53.435 2.64 ;
      RECT 53.405 2.175 53.425 2.64 ;
      RECT 53.375 2.22 53.405 2.64 ;
      RECT 53.37 2.247 53.375 2.64 ;
      RECT 53.35 2.265 53.37 2.64 ;
      RECT 53.34 2.29 53.35 2.64 ;
      RECT 53.335 2.302 53.34 2.64 ;
      RECT 53.32 2.325 53.335 2.64 ;
      RECT 53.3 2.352 53.315 2.64 ;
      RECT 53.29 2.375 53.3 2.64 ;
      RECT 55.08 3.26 55.16 3.52 ;
      RECT 54.315 2.48 54.385 2.74 ;
      RECT 55.046 3.227 55.08 3.52 ;
      RECT 54.96 3.13 55.046 3.52 ;
      RECT 54.94 3.042 54.96 3.52 ;
      RECT 54.93 3.012 54.94 3.52 ;
      RECT 54.92 2.992 54.93 3.52 ;
      RECT 54.9 2.979 54.92 3.52 ;
      RECT 54.885 2.969 54.9 3.348 ;
      RECT 54.88 2.962 54.885 3.303 ;
      RECT 54.87 2.956 54.88 3.293 ;
      RECT 54.86 2.948 54.87 3.275 ;
      RECT 54.855 2.942 54.86 3.263 ;
      RECT 54.845 2.937 54.855 3.25 ;
      RECT 54.825 2.927 54.845 3.223 ;
      RECT 54.785 2.906 54.825 3.175 ;
      RECT 54.77 2.887 54.785 3.133 ;
      RECT 54.745 2.873 54.77 3.103 ;
      RECT 54.735 2.861 54.745 3.07 ;
      RECT 54.73 2.856 54.735 3.06 ;
      RECT 54.7 2.842 54.73 3.04 ;
      RECT 54.69 2.826 54.7 3.013 ;
      RECT 54.685 2.821 54.69 3.003 ;
      RECT 54.66 2.812 54.685 2.983 ;
      RECT 54.65 2.8 54.66 2.963 ;
      RECT 54.58 2.768 54.65 2.938 ;
      RECT 54.575 2.737 54.58 2.915 ;
      RECT 54.526 2.48 54.575 2.898 ;
      RECT 54.44 2.48 54.526 2.857 ;
      RECT 54.385 2.48 54.44 2.785 ;
      RECT 54.475 3.265 54.635 3.525 ;
      RECT 54 1.88 54.05 2.565 ;
      RECT 53.79 2.305 53.825 2.565 ;
      RECT 54.105 1.88 54.11 2.34 ;
      RECT 54.195 1.88 54.22 2.16 ;
      RECT 54.47 3.262 54.475 3.525 ;
      RECT 54.435 3.25 54.47 3.525 ;
      RECT 54.375 3.223 54.435 3.525 ;
      RECT 54.37 3.206 54.375 3.379 ;
      RECT 54.365 3.203 54.37 3.366 ;
      RECT 54.345 3.196 54.365 3.353 ;
      RECT 54.31 3.179 54.345 3.335 ;
      RECT 54.27 3.158 54.31 3.315 ;
      RECT 54.265 3.146 54.27 3.303 ;
      RECT 54.225 3.132 54.265 3.289 ;
      RECT 54.205 3.115 54.225 3.271 ;
      RECT 54.195 3.107 54.205 3.263 ;
      RECT 54.18 1.88 54.195 2.178 ;
      RECT 54.165 3.097 54.195 3.25 ;
      RECT 54.15 1.88 54.18 2.223 ;
      RECT 54.155 3.087 54.165 3.237 ;
      RECT 54.125 3.072 54.155 3.224 ;
      RECT 54.11 1.88 54.15 2.29 ;
      RECT 54.11 3.04 54.125 3.21 ;
      RECT 54.105 3.012 54.11 3.204 ;
      RECT 54.1 1.88 54.105 2.345 ;
      RECT 54.09 2.982 54.105 3.198 ;
      RECT 54.095 1.88 54.1 2.358 ;
      RECT 54.085 1.88 54.095 2.378 ;
      RECT 54.05 2.895 54.09 3.183 ;
      RECT 54.05 1.88 54.085 2.418 ;
      RECT 54.045 2.827 54.05 3.171 ;
      RECT 54.03 2.782 54.045 3.166 ;
      RECT 54.025 2.72 54.03 3.161 ;
      RECT 54 2.627 54.025 3.154 ;
      RECT 53.995 1.88 54 3.146 ;
      RECT 53.98 1.88 53.995 3.133 ;
      RECT 53.96 1.88 53.98 3.09 ;
      RECT 53.95 1.88 53.96 3.04 ;
      RECT 53.945 1.88 53.95 3.013 ;
      RECT 53.94 1.88 53.945 2.991 ;
      RECT 53.935 2.106 53.94 2.974 ;
      RECT 53.93 2.128 53.935 2.952 ;
      RECT 53.925 2.17 53.93 2.935 ;
      RECT 53.895 2.22 53.925 2.879 ;
      RECT 53.89 2.247 53.895 2.821 ;
      RECT 53.875 2.265 53.89 2.785 ;
      RECT 53.87 2.283 53.875 2.749 ;
      RECT 53.864 2.29 53.87 2.73 ;
      RECT 53.86 2.297 53.864 2.713 ;
      RECT 53.855 2.302 53.86 2.682 ;
      RECT 53.845 2.305 53.855 2.657 ;
      RECT 53.835 2.305 53.845 2.623 ;
      RECT 53.83 2.305 53.835 2.6 ;
      RECT 53.825 2.305 53.83 2.58 ;
      RECT 52.74 2.44 53.02 2.72 ;
      RECT 52.74 2.44 53.04 2.615 ;
      RECT 52.83 2.33 53.09 2.59 ;
      RECT 52.795 2.425 53.09 2.59 ;
      RECT 52.92 0.945 53.085 2.59 ;
      RECT 52.82 0.945 53.19 1.315 ;
      RECT 52.445 3.47 52.705 3.73 ;
      RECT 52.465 3.397 52.645 3.73 ;
      RECT 52.465 3.14 52.64 3.73 ;
      RECT 52.465 2.932 52.63 3.73 ;
      RECT 52.47 2.85 52.63 3.73 ;
      RECT 52.47 2.615 52.62 3.73 ;
      RECT 52.47 2.462 52.615 3.73 ;
      RECT 52.475 2.447 52.615 3.73 ;
      RECT 52.525 2.162 52.615 3.73 ;
      RECT 52.48 2.397 52.615 3.73 ;
      RECT 52.51 2.215 52.615 3.73 ;
      RECT 52.495 2.327 52.615 3.73 ;
      RECT 52.5 2.285 52.615 3.73 ;
      RECT 52.495 2.327 52.63 2.39 ;
      RECT 52.53 1.915 52.635 2.335 ;
      RECT 52.53 1.915 52.65 2.318 ;
      RECT 52.53 1.915 52.685 2.28 ;
      RECT 52.525 2.162 52.735 2.213 ;
      RECT 52.53 1.915 52.79 2.175 ;
      RECT 51.79 2.62 52.05 2.88 ;
      RECT 51.79 2.62 52.06 2.838 ;
      RECT 51.79 2.62 52.146 2.809 ;
      RECT 51.79 2.62 52.215 2.761 ;
      RECT 51.79 2.62 52.25 2.73 ;
      RECT 52.02 2.44 52.3 2.72 ;
      RECT 51.855 2.605 52.3 2.72 ;
      RECT 51.945 2.482 52.05 2.88 ;
      RECT 51.875 2.545 52.3 2.72 ;
      RECT 46.325 6.22 46.645 6.545 ;
      RECT 46.355 5.695 46.525 6.545 ;
      RECT 46.355 5.695 46.53 6.045 ;
      RECT 46.355 5.695 47.33 5.87 ;
      RECT 47.155 1.965 47.33 5.87 ;
      RECT 47.1 1.965 47.45 2.315 ;
      RECT 47.125 6.655 47.45 6.98 ;
      RECT 46.01 6.745 47.45 6.915 ;
      RECT 46.01 2.395 46.17 6.915 ;
      RECT 46.325 2.365 46.645 2.685 ;
      RECT 46.01 2.395 46.645 2.565 ;
      RECT 44.675 2.705 45.06 3.055 ;
      RECT 44.665 2.77 45.06 2.97 ;
      RECT 44.81 2.7 44.98 3.055 ;
      RECT 43.12 2.44 43.4 2.72 ;
      RECT 43.115 2.44 43.4 2.673 ;
      RECT 43.095 2.44 43.4 2.65 ;
      RECT 43.085 2.44 43.4 2.63 ;
      RECT 43.075 2.44 43.4 2.615 ;
      RECT 43.05 2.44 43.4 2.588 ;
      RECT 43.04 2.44 43.4 2.563 ;
      RECT 42.995 2.295 43.275 2.555 ;
      RECT 42.995 2.39 43.375 2.555 ;
      RECT 42.995 2.335 43.32 2.555 ;
      RECT 42.995 2.327 43.315 2.555 ;
      RECT 42.995 2.317 43.31 2.555 ;
      RECT 42.995 2.305 43.305 2.555 ;
      RECT 41.92 3 42.2 3.28 ;
      RECT 41.92 3 42.235 3.26 ;
      RECT 34.245 6.66 34.595 7.01 ;
      RECT 41.665 6.615 42.015 6.965 ;
      RECT 34.245 6.69 42.015 6.89 ;
      RECT 41.955 2.42 42.005 2.68 ;
      RECT 41.745 2.42 41.75 2.68 ;
      RECT 40.94 1.975 40.97 2.235 ;
      RECT 40.71 1.975 40.785 2.235 ;
      RECT 41.93 2.37 41.955 2.68 ;
      RECT 41.925 2.327 41.93 2.68 ;
      RECT 41.92 2.31 41.925 2.68 ;
      RECT 41.915 2.297 41.92 2.68 ;
      RECT 41.84 2.18 41.915 2.68 ;
      RECT 41.795 1.997 41.84 2.68 ;
      RECT 41.79 1.925 41.795 2.68 ;
      RECT 41.775 1.9 41.79 2.68 ;
      RECT 41.75 1.862 41.775 2.68 ;
      RECT 41.74 1.842 41.75 2.402 ;
      RECT 41.725 1.834 41.74 2.357 ;
      RECT 41.72 1.826 41.725 2.328 ;
      RECT 41.715 1.823 41.72 2.308 ;
      RECT 41.71 1.82 41.715 2.288 ;
      RECT 41.705 1.817 41.71 2.268 ;
      RECT 41.675 1.806 41.705 2.205 ;
      RECT 41.655 1.791 41.675 2.12 ;
      RECT 41.65 1.783 41.655 2.083 ;
      RECT 41.64 1.777 41.65 2.05 ;
      RECT 41.625 1.769 41.64 2.01 ;
      RECT 41.62 1.762 41.625 1.97 ;
      RECT 41.615 1.759 41.62 1.948 ;
      RECT 41.61 1.756 41.615 1.935 ;
      RECT 41.605 1.755 41.61 1.925 ;
      RECT 41.59 1.749 41.605 1.915 ;
      RECT 41.565 1.736 41.59 1.9 ;
      RECT 41.515 1.711 41.565 1.871 ;
      RECT 41.5 1.69 41.515 1.846 ;
      RECT 41.49 1.683 41.5 1.835 ;
      RECT 41.435 1.664 41.49 1.808 ;
      RECT 41.41 1.642 41.435 1.781 ;
      RECT 41.405 1.635 41.41 1.776 ;
      RECT 41.39 1.635 41.405 1.774 ;
      RECT 41.365 1.627 41.39 1.77 ;
      RECT 41.35 1.625 41.365 1.766 ;
      RECT 41.32 1.625 41.35 1.763 ;
      RECT 41.31 1.625 41.32 1.758 ;
      RECT 41.265 1.625 41.31 1.756 ;
      RECT 41.236 1.625 41.265 1.757 ;
      RECT 41.15 1.625 41.236 1.759 ;
      RECT 41.136 1.626 41.15 1.761 ;
      RECT 41.05 1.627 41.136 1.763 ;
      RECT 41.035 1.628 41.05 1.773 ;
      RECT 41.03 1.629 41.035 1.782 ;
      RECT 41.01 1.632 41.03 1.792 ;
      RECT 40.995 1.64 41.01 1.807 ;
      RECT 40.975 1.658 40.995 1.822 ;
      RECT 40.965 1.67 40.975 1.845 ;
      RECT 40.955 1.679 40.965 1.875 ;
      RECT 40.94 1.691 40.955 1.92 ;
      RECT 40.885 1.724 40.94 2.235 ;
      RECT 40.88 1.752 40.885 2.235 ;
      RECT 40.86 1.767 40.88 2.235 ;
      RECT 40.825 1.827 40.86 2.235 ;
      RECT 40.823 1.877 40.825 2.235 ;
      RECT 40.82 1.885 40.823 2.235 ;
      RECT 40.81 1.9 40.82 2.235 ;
      RECT 40.805 1.912 40.81 2.235 ;
      RECT 40.795 1.937 40.805 2.235 ;
      RECT 40.785 1.965 40.795 2.235 ;
      RECT 38.69 3.47 38.74 3.73 ;
      RECT 41.6 3.02 41.66 3.28 ;
      RECT 41.585 3.02 41.6 3.29 ;
      RECT 41.566 3.02 41.585 3.323 ;
      RECT 41.48 3.02 41.566 3.448 ;
      RECT 41.4 3.02 41.48 3.63 ;
      RECT 41.395 3.257 41.4 3.715 ;
      RECT 41.37 3.327 41.395 3.743 ;
      RECT 41.365 3.397 41.37 3.77 ;
      RECT 41.345 3.469 41.365 3.792 ;
      RECT 41.34 3.536 41.345 3.815 ;
      RECT 41.33 3.565 41.34 3.83 ;
      RECT 41.32 3.587 41.33 3.847 ;
      RECT 41.315 3.597 41.32 3.858 ;
      RECT 41.31 3.605 41.315 3.866 ;
      RECT 41.3 3.613 41.31 3.878 ;
      RECT 41.295 3.625 41.3 3.888 ;
      RECT 41.29 3.633 41.295 3.893 ;
      RECT 41.27 3.651 41.29 3.903 ;
      RECT 41.265 3.668 41.27 3.91 ;
      RECT 41.26 3.676 41.265 3.911 ;
      RECT 41.255 3.687 41.26 3.913 ;
      RECT 41.215 3.725 41.255 3.923 ;
      RECT 41.21 3.76 41.215 3.934 ;
      RECT 41.205 3.765 41.21 3.937 ;
      RECT 41.18 3.775 41.205 3.944 ;
      RECT 41.17 3.789 41.18 3.953 ;
      RECT 41.15 3.801 41.17 3.956 ;
      RECT 41.1 3.82 41.15 3.96 ;
      RECT 41.055 3.835 41.1 3.965 ;
      RECT 40.99 3.838 41.055 3.971 ;
      RECT 40.975 3.836 40.99 3.978 ;
      RECT 40.945 3.835 40.975 3.978 ;
      RECT 40.906 3.834 40.945 3.974 ;
      RECT 40.82 3.831 40.906 3.97 ;
      RECT 40.803 3.829 40.82 3.967 ;
      RECT 40.717 3.827 40.803 3.964 ;
      RECT 40.631 3.824 40.717 3.958 ;
      RECT 40.545 3.82 40.631 3.953 ;
      RECT 40.467 3.817 40.545 3.949 ;
      RECT 40.381 3.814 40.467 3.947 ;
      RECT 40.295 3.811 40.381 3.944 ;
      RECT 40.237 3.809 40.295 3.941 ;
      RECT 40.151 3.806 40.237 3.939 ;
      RECT 40.065 3.802 40.151 3.937 ;
      RECT 39.979 3.799 40.065 3.934 ;
      RECT 39.893 3.795 39.979 3.932 ;
      RECT 39.807 3.791 39.893 3.929 ;
      RECT 39.721 3.788 39.807 3.927 ;
      RECT 39.635 3.784 39.721 3.924 ;
      RECT 39.549 3.781 39.635 3.922 ;
      RECT 39.463 3.777 39.549 3.919 ;
      RECT 39.377 3.774 39.463 3.917 ;
      RECT 39.291 3.77 39.377 3.914 ;
      RECT 39.205 3.767 39.291 3.912 ;
      RECT 39.195 3.765 39.205 3.908 ;
      RECT 39.19 3.765 39.195 3.906 ;
      RECT 39.15 3.76 39.19 3.9 ;
      RECT 39.136 3.751 39.15 3.893 ;
      RECT 39.05 3.721 39.136 3.878 ;
      RECT 39.03 3.687 39.05 3.863 ;
      RECT 38.96 3.656 39.03 3.85 ;
      RECT 38.955 3.631 38.96 3.839 ;
      RECT 38.95 3.625 38.955 3.837 ;
      RECT 38.881 3.47 38.95 3.825 ;
      RECT 38.795 3.47 38.881 3.799 ;
      RECT 38.77 3.47 38.795 3.778 ;
      RECT 38.765 3.47 38.77 3.768 ;
      RECT 38.76 3.47 38.765 3.76 ;
      RECT 38.74 3.47 38.76 3.743 ;
      RECT 41.16 2.04 41.42 2.3 ;
      RECT 41.145 2.04 41.42 2.203 ;
      RECT 41.115 2.04 41.42 2.178 ;
      RECT 41.08 1.88 41.36 2.16 ;
      RECT 41.05 3.37 41.11 3.63 ;
      RECT 40.075 2.06 40.13 2.32 ;
      RECT 41.01 3.327 41.05 3.63 ;
      RECT 40.981 3.248 41.01 3.63 ;
      RECT 40.895 3.12 40.981 3.63 ;
      RECT 40.875 3 40.895 3.63 ;
      RECT 40.85 2.951 40.875 3.63 ;
      RECT 40.845 2.916 40.85 3.48 ;
      RECT 40.815 2.876 40.845 3.418 ;
      RECT 40.79 2.813 40.815 3.333 ;
      RECT 40.78 2.775 40.79 3.27 ;
      RECT 40.765 2.75 40.78 3.231 ;
      RECT 40.722 2.708 40.765 3.137 ;
      RECT 40.72 2.681 40.722 3.064 ;
      RECT 40.715 2.676 40.72 3.055 ;
      RECT 40.71 2.669 40.715 3.03 ;
      RECT 40.705 2.663 40.71 3.015 ;
      RECT 40.7 2.657 40.705 3.003 ;
      RECT 40.69 2.648 40.7 2.985 ;
      RECT 40.685 2.639 40.69 2.963 ;
      RECT 40.66 2.62 40.685 2.913 ;
      RECT 40.655 2.601 40.66 2.863 ;
      RECT 40.64 2.587 40.655 2.823 ;
      RECT 40.635 2.573 40.64 2.79 ;
      RECT 40.63 2.566 40.635 2.783 ;
      RECT 40.615 2.553 40.63 2.775 ;
      RECT 40.57 2.515 40.615 2.748 ;
      RECT 40.54 2.468 40.57 2.713 ;
      RECT 40.52 2.437 40.54 2.69 ;
      RECT 40.44 2.37 40.52 2.643 ;
      RECT 40.41 2.3 40.44 2.59 ;
      RECT 40.405 2.277 40.41 2.573 ;
      RECT 40.375 2.255 40.405 2.558 ;
      RECT 40.345 2.214 40.375 2.53 ;
      RECT 40.34 2.189 40.345 2.515 ;
      RECT 40.335 2.183 40.34 2.508 ;
      RECT 40.325 2.06 40.335 2.5 ;
      RECT 40.315 2.06 40.325 2.493 ;
      RECT 40.31 2.06 40.315 2.485 ;
      RECT 40.29 2.06 40.31 2.473 ;
      RECT 40.24 2.06 40.29 2.443 ;
      RECT 40.185 2.06 40.24 2.393 ;
      RECT 40.155 2.06 40.185 2.353 ;
      RECT 40.13 2.06 40.155 2.33 ;
      RECT 40 2.785 40.28 3.065 ;
      RECT 39.965 2.7 40.225 2.96 ;
      RECT 39.965 2.782 40.235 2.96 ;
      RECT 38.165 2.155 38.17 2.64 ;
      RECT 38.055 2.34 38.06 2.64 ;
      RECT 37.965 2.38 38.03 2.64 ;
      RECT 39.64 1.88 39.73 2.51 ;
      RECT 39.605 1.93 39.61 2.51 ;
      RECT 39.55 1.955 39.56 2.51 ;
      RECT 39.505 1.955 39.515 2.51 ;
      RECT 39.875 1.88 39.92 2.16 ;
      RECT 38.725 1.61 38.925 1.75 ;
      RECT 39.841 1.88 39.875 2.172 ;
      RECT 39.755 1.88 39.841 2.212 ;
      RECT 39.74 1.88 39.755 2.253 ;
      RECT 39.735 1.88 39.74 2.273 ;
      RECT 39.73 1.88 39.735 2.293 ;
      RECT 39.61 1.922 39.64 2.51 ;
      RECT 39.56 1.942 39.605 2.51 ;
      RECT 39.545 1.957 39.55 2.51 ;
      RECT 39.515 1.957 39.545 2.51 ;
      RECT 39.47 1.942 39.505 2.51 ;
      RECT 39.465 1.93 39.47 2.29 ;
      RECT 39.46 1.927 39.465 2.27 ;
      RECT 39.445 1.917 39.46 2.223 ;
      RECT 39.44 1.91 39.445 2.186 ;
      RECT 39.435 1.907 39.44 2.169 ;
      RECT 39.42 1.897 39.435 2.125 ;
      RECT 39.415 1.888 39.42 2.085 ;
      RECT 39.41 1.884 39.415 2.07 ;
      RECT 39.4 1.878 39.41 2.053 ;
      RECT 39.36 1.859 39.4 2.028 ;
      RECT 39.355 1.841 39.36 2.008 ;
      RECT 39.345 1.835 39.355 2.003 ;
      RECT 39.315 1.819 39.345 1.99 ;
      RECT 39.3 1.801 39.315 1.973 ;
      RECT 39.285 1.789 39.3 1.96 ;
      RECT 39.28 1.781 39.285 1.953 ;
      RECT 39.25 1.767 39.28 1.94 ;
      RECT 39.245 1.752 39.25 1.928 ;
      RECT 39.235 1.746 39.245 1.92 ;
      RECT 39.215 1.734 39.235 1.908 ;
      RECT 39.205 1.722 39.215 1.895 ;
      RECT 39.175 1.706 39.205 1.88 ;
      RECT 39.155 1.686 39.175 1.863 ;
      RECT 39.15 1.676 39.155 1.853 ;
      RECT 39.125 1.664 39.15 1.84 ;
      RECT 39.12 1.652 39.125 1.828 ;
      RECT 39.115 1.647 39.12 1.824 ;
      RECT 39.1 1.64 39.115 1.816 ;
      RECT 39.09 1.627 39.1 1.806 ;
      RECT 39.085 1.625 39.09 1.8 ;
      RECT 39.06 1.618 39.085 1.789 ;
      RECT 39.055 1.611 39.06 1.778 ;
      RECT 39.03 1.61 39.055 1.765 ;
      RECT 39.011 1.61 39.03 1.755 ;
      RECT 38.925 1.61 39.011 1.752 ;
      RECT 38.695 1.61 38.725 1.755 ;
      RECT 38.655 1.617 38.695 1.768 ;
      RECT 38.63 1.627 38.655 1.781 ;
      RECT 38.615 1.636 38.63 1.791 ;
      RECT 38.585 1.641 38.615 1.81 ;
      RECT 38.58 1.647 38.585 1.828 ;
      RECT 38.56 1.657 38.58 1.843 ;
      RECT 38.55 1.67 38.56 1.863 ;
      RECT 38.535 1.682 38.55 1.88 ;
      RECT 38.53 1.692 38.535 1.89 ;
      RECT 38.525 1.697 38.53 1.895 ;
      RECT 38.515 1.705 38.525 1.908 ;
      RECT 38.465 1.737 38.515 1.945 ;
      RECT 38.45 1.772 38.465 1.986 ;
      RECT 38.445 1.782 38.45 2.001 ;
      RECT 38.44 1.787 38.445 2.008 ;
      RECT 38.415 1.803 38.44 2.028 ;
      RECT 38.4 1.824 38.415 2.053 ;
      RECT 38.375 1.845 38.4 2.078 ;
      RECT 38.365 1.864 38.375 2.101 ;
      RECT 38.34 1.882 38.365 2.124 ;
      RECT 38.325 1.902 38.34 2.148 ;
      RECT 38.32 1.912 38.325 2.16 ;
      RECT 38.305 1.924 38.32 2.18 ;
      RECT 38.295 1.939 38.305 2.22 ;
      RECT 38.29 1.947 38.295 2.248 ;
      RECT 38.28 1.957 38.29 2.268 ;
      RECT 38.275 1.97 38.28 2.293 ;
      RECT 38.27 1.983 38.275 2.313 ;
      RECT 38.265 1.989 38.27 2.335 ;
      RECT 38.255 1.998 38.265 2.355 ;
      RECT 38.25 2.018 38.255 2.378 ;
      RECT 38.245 2.024 38.25 2.398 ;
      RECT 38.24 2.031 38.245 2.42 ;
      RECT 38.235 2.042 38.24 2.433 ;
      RECT 38.225 2.052 38.235 2.458 ;
      RECT 38.205 2.077 38.225 2.64 ;
      RECT 38.175 2.117 38.205 2.64 ;
      RECT 38.17 2.147 38.175 2.64 ;
      RECT 38.145 2.175 38.165 2.64 ;
      RECT 38.115 2.22 38.145 2.64 ;
      RECT 38.11 2.247 38.115 2.64 ;
      RECT 38.09 2.265 38.11 2.64 ;
      RECT 38.08 2.29 38.09 2.64 ;
      RECT 38.075 2.302 38.08 2.64 ;
      RECT 38.06 2.325 38.075 2.64 ;
      RECT 38.04 2.352 38.055 2.64 ;
      RECT 38.03 2.375 38.04 2.64 ;
      RECT 39.82 3.26 39.9 3.52 ;
      RECT 39.055 2.48 39.125 2.74 ;
      RECT 39.786 3.227 39.82 3.52 ;
      RECT 39.7 3.13 39.786 3.52 ;
      RECT 39.68 3.042 39.7 3.52 ;
      RECT 39.67 3.012 39.68 3.52 ;
      RECT 39.66 2.992 39.67 3.52 ;
      RECT 39.64 2.979 39.66 3.52 ;
      RECT 39.625 2.969 39.64 3.348 ;
      RECT 39.62 2.962 39.625 3.303 ;
      RECT 39.61 2.956 39.62 3.293 ;
      RECT 39.6 2.948 39.61 3.275 ;
      RECT 39.595 2.942 39.6 3.263 ;
      RECT 39.585 2.937 39.595 3.25 ;
      RECT 39.565 2.927 39.585 3.223 ;
      RECT 39.525 2.906 39.565 3.175 ;
      RECT 39.51 2.887 39.525 3.133 ;
      RECT 39.485 2.873 39.51 3.103 ;
      RECT 39.475 2.861 39.485 3.07 ;
      RECT 39.47 2.856 39.475 3.06 ;
      RECT 39.44 2.842 39.47 3.04 ;
      RECT 39.43 2.826 39.44 3.013 ;
      RECT 39.425 2.821 39.43 3.003 ;
      RECT 39.4 2.812 39.425 2.983 ;
      RECT 39.39 2.8 39.4 2.963 ;
      RECT 39.32 2.768 39.39 2.938 ;
      RECT 39.315 2.737 39.32 2.915 ;
      RECT 39.266 2.48 39.315 2.898 ;
      RECT 39.18 2.48 39.266 2.857 ;
      RECT 39.125 2.48 39.18 2.785 ;
      RECT 39.215 3.265 39.375 3.525 ;
      RECT 38.74 1.88 38.79 2.565 ;
      RECT 38.53 2.305 38.565 2.565 ;
      RECT 38.845 1.88 38.85 2.34 ;
      RECT 38.935 1.88 38.96 2.16 ;
      RECT 39.21 3.262 39.215 3.525 ;
      RECT 39.175 3.25 39.21 3.525 ;
      RECT 39.115 3.223 39.175 3.525 ;
      RECT 39.11 3.206 39.115 3.379 ;
      RECT 39.105 3.203 39.11 3.366 ;
      RECT 39.085 3.196 39.105 3.353 ;
      RECT 39.05 3.179 39.085 3.335 ;
      RECT 39.01 3.158 39.05 3.315 ;
      RECT 39.005 3.146 39.01 3.303 ;
      RECT 38.965 3.132 39.005 3.289 ;
      RECT 38.945 3.115 38.965 3.271 ;
      RECT 38.935 3.107 38.945 3.263 ;
      RECT 38.92 1.88 38.935 2.178 ;
      RECT 38.905 3.097 38.935 3.25 ;
      RECT 38.89 1.88 38.92 2.223 ;
      RECT 38.895 3.087 38.905 3.237 ;
      RECT 38.865 3.072 38.895 3.224 ;
      RECT 38.85 1.88 38.89 2.29 ;
      RECT 38.85 3.04 38.865 3.21 ;
      RECT 38.845 3.012 38.85 3.204 ;
      RECT 38.84 1.88 38.845 2.345 ;
      RECT 38.83 2.982 38.845 3.198 ;
      RECT 38.835 1.88 38.84 2.358 ;
      RECT 38.825 1.88 38.835 2.378 ;
      RECT 38.79 2.895 38.83 3.183 ;
      RECT 38.79 1.88 38.825 2.418 ;
      RECT 38.785 2.827 38.79 3.171 ;
      RECT 38.77 2.782 38.785 3.166 ;
      RECT 38.765 2.72 38.77 3.161 ;
      RECT 38.74 2.627 38.765 3.154 ;
      RECT 38.735 1.88 38.74 3.146 ;
      RECT 38.72 1.88 38.735 3.133 ;
      RECT 38.7 1.88 38.72 3.09 ;
      RECT 38.69 1.88 38.7 3.04 ;
      RECT 38.685 1.88 38.69 3.013 ;
      RECT 38.68 1.88 38.685 2.991 ;
      RECT 38.675 2.106 38.68 2.974 ;
      RECT 38.67 2.128 38.675 2.952 ;
      RECT 38.665 2.17 38.67 2.935 ;
      RECT 38.635 2.22 38.665 2.879 ;
      RECT 38.63 2.247 38.635 2.821 ;
      RECT 38.615 2.265 38.63 2.785 ;
      RECT 38.61 2.283 38.615 2.749 ;
      RECT 38.604 2.29 38.61 2.73 ;
      RECT 38.6 2.297 38.604 2.713 ;
      RECT 38.595 2.302 38.6 2.682 ;
      RECT 38.585 2.305 38.595 2.657 ;
      RECT 38.575 2.305 38.585 2.623 ;
      RECT 38.57 2.305 38.575 2.6 ;
      RECT 38.565 2.305 38.57 2.58 ;
      RECT 37.48 2.44 37.76 2.72 ;
      RECT 37.48 2.44 37.78 2.615 ;
      RECT 37.57 2.33 37.83 2.59 ;
      RECT 37.535 2.425 37.83 2.59 ;
      RECT 37.66 0.945 37.825 2.59 ;
      RECT 37.56 0.945 37.93 1.315 ;
      RECT 37.185 3.47 37.445 3.73 ;
      RECT 37.205 3.397 37.385 3.73 ;
      RECT 37.205 3.14 37.38 3.73 ;
      RECT 37.205 2.932 37.37 3.73 ;
      RECT 37.21 2.85 37.37 3.73 ;
      RECT 37.21 2.615 37.36 3.73 ;
      RECT 37.21 2.462 37.355 3.73 ;
      RECT 37.215 2.447 37.355 3.73 ;
      RECT 37.265 2.162 37.355 3.73 ;
      RECT 37.22 2.397 37.355 3.73 ;
      RECT 37.25 2.215 37.355 3.73 ;
      RECT 37.235 2.327 37.355 3.73 ;
      RECT 37.24 2.285 37.355 3.73 ;
      RECT 37.235 2.327 37.37 2.39 ;
      RECT 37.27 1.915 37.375 2.335 ;
      RECT 37.27 1.915 37.39 2.318 ;
      RECT 37.27 1.915 37.425 2.28 ;
      RECT 37.265 2.162 37.475 2.213 ;
      RECT 37.27 1.915 37.53 2.175 ;
      RECT 36.53 2.62 36.79 2.88 ;
      RECT 36.53 2.62 36.8 2.838 ;
      RECT 36.53 2.62 36.886 2.809 ;
      RECT 36.53 2.62 36.955 2.761 ;
      RECT 36.53 2.62 36.99 2.73 ;
      RECT 36.76 2.44 37.04 2.72 ;
      RECT 36.595 2.605 37.04 2.72 ;
      RECT 36.685 2.482 36.79 2.88 ;
      RECT 36.615 2.545 37.04 2.72 ;
      RECT 31.065 6.22 31.385 6.545 ;
      RECT 31.095 5.695 31.265 6.545 ;
      RECT 31.095 5.695 31.27 6.045 ;
      RECT 31.095 5.695 32.07 5.87 ;
      RECT 31.895 1.965 32.07 5.87 ;
      RECT 31.84 1.965 32.19 2.315 ;
      RECT 31.865 6.655 32.19 6.98 ;
      RECT 30.75 6.745 32.19 6.915 ;
      RECT 30.75 2.395 30.91 6.915 ;
      RECT 31.065 2.365 31.385 2.685 ;
      RECT 30.75 2.395 31.385 2.565 ;
      RECT 29.415 2.705 29.8 3.055 ;
      RECT 29.405 2.77 29.8 2.97 ;
      RECT 29.55 2.7 29.72 3.055 ;
      RECT 27.86 2.44 28.14 2.72 ;
      RECT 27.855 2.44 28.14 2.673 ;
      RECT 27.835 2.44 28.14 2.65 ;
      RECT 27.825 2.44 28.14 2.63 ;
      RECT 27.815 2.44 28.14 2.615 ;
      RECT 27.79 2.44 28.14 2.588 ;
      RECT 27.78 2.44 28.14 2.563 ;
      RECT 27.735 2.295 28.015 2.555 ;
      RECT 27.735 2.39 28.115 2.555 ;
      RECT 27.735 2.335 28.06 2.555 ;
      RECT 27.735 2.327 28.055 2.555 ;
      RECT 27.735 2.317 28.05 2.555 ;
      RECT 27.735 2.305 28.045 2.555 ;
      RECT 26.66 3 26.94 3.28 ;
      RECT 26.66 3 26.975 3.26 ;
      RECT 18.985 6.655 19.335 7.005 ;
      RECT 26.405 6.61 26.755 6.96 ;
      RECT 18.985 6.685 26.755 6.885 ;
      RECT 26.695 2.42 26.745 2.68 ;
      RECT 26.485 2.42 26.49 2.68 ;
      RECT 25.68 1.975 25.71 2.235 ;
      RECT 25.45 1.975 25.525 2.235 ;
      RECT 26.67 2.37 26.695 2.68 ;
      RECT 26.665 2.327 26.67 2.68 ;
      RECT 26.66 2.31 26.665 2.68 ;
      RECT 26.655 2.297 26.66 2.68 ;
      RECT 26.58 2.18 26.655 2.68 ;
      RECT 26.535 1.997 26.58 2.68 ;
      RECT 26.53 1.925 26.535 2.68 ;
      RECT 26.515 1.9 26.53 2.68 ;
      RECT 26.49 1.862 26.515 2.68 ;
      RECT 26.48 1.842 26.49 2.402 ;
      RECT 26.465 1.834 26.48 2.357 ;
      RECT 26.46 1.826 26.465 2.328 ;
      RECT 26.455 1.823 26.46 2.308 ;
      RECT 26.45 1.82 26.455 2.288 ;
      RECT 26.445 1.817 26.45 2.268 ;
      RECT 26.415 1.806 26.445 2.205 ;
      RECT 26.395 1.791 26.415 2.12 ;
      RECT 26.39 1.783 26.395 2.083 ;
      RECT 26.38 1.777 26.39 2.05 ;
      RECT 26.365 1.769 26.38 2.01 ;
      RECT 26.36 1.762 26.365 1.97 ;
      RECT 26.355 1.759 26.36 1.948 ;
      RECT 26.35 1.756 26.355 1.935 ;
      RECT 26.345 1.755 26.35 1.925 ;
      RECT 26.33 1.749 26.345 1.915 ;
      RECT 26.305 1.736 26.33 1.9 ;
      RECT 26.255 1.711 26.305 1.871 ;
      RECT 26.24 1.69 26.255 1.846 ;
      RECT 26.23 1.683 26.24 1.835 ;
      RECT 26.175 1.664 26.23 1.808 ;
      RECT 26.15 1.642 26.175 1.781 ;
      RECT 26.145 1.635 26.15 1.776 ;
      RECT 26.13 1.635 26.145 1.774 ;
      RECT 26.105 1.627 26.13 1.77 ;
      RECT 26.09 1.625 26.105 1.766 ;
      RECT 26.06 1.625 26.09 1.763 ;
      RECT 26.05 1.625 26.06 1.758 ;
      RECT 26.005 1.625 26.05 1.756 ;
      RECT 25.976 1.625 26.005 1.757 ;
      RECT 25.89 1.625 25.976 1.759 ;
      RECT 25.876 1.626 25.89 1.761 ;
      RECT 25.79 1.627 25.876 1.763 ;
      RECT 25.775 1.628 25.79 1.773 ;
      RECT 25.77 1.629 25.775 1.782 ;
      RECT 25.75 1.632 25.77 1.792 ;
      RECT 25.735 1.64 25.75 1.807 ;
      RECT 25.715 1.658 25.735 1.822 ;
      RECT 25.705 1.67 25.715 1.845 ;
      RECT 25.695 1.679 25.705 1.875 ;
      RECT 25.68 1.691 25.695 1.92 ;
      RECT 25.625 1.724 25.68 2.235 ;
      RECT 25.62 1.752 25.625 2.235 ;
      RECT 25.6 1.767 25.62 2.235 ;
      RECT 25.565 1.827 25.6 2.235 ;
      RECT 25.563 1.877 25.565 2.235 ;
      RECT 25.56 1.885 25.563 2.235 ;
      RECT 25.55 1.9 25.56 2.235 ;
      RECT 25.545 1.912 25.55 2.235 ;
      RECT 25.535 1.937 25.545 2.235 ;
      RECT 25.525 1.965 25.535 2.235 ;
      RECT 23.43 3.47 23.48 3.73 ;
      RECT 26.34 3.02 26.4 3.28 ;
      RECT 26.325 3.02 26.34 3.29 ;
      RECT 26.306 3.02 26.325 3.323 ;
      RECT 26.22 3.02 26.306 3.448 ;
      RECT 26.14 3.02 26.22 3.63 ;
      RECT 26.135 3.257 26.14 3.715 ;
      RECT 26.11 3.327 26.135 3.743 ;
      RECT 26.105 3.397 26.11 3.77 ;
      RECT 26.085 3.469 26.105 3.792 ;
      RECT 26.08 3.536 26.085 3.815 ;
      RECT 26.07 3.565 26.08 3.83 ;
      RECT 26.06 3.587 26.07 3.847 ;
      RECT 26.055 3.597 26.06 3.858 ;
      RECT 26.05 3.605 26.055 3.866 ;
      RECT 26.04 3.613 26.05 3.878 ;
      RECT 26.035 3.625 26.04 3.888 ;
      RECT 26.03 3.633 26.035 3.893 ;
      RECT 26.01 3.651 26.03 3.903 ;
      RECT 26.005 3.668 26.01 3.91 ;
      RECT 26 3.676 26.005 3.911 ;
      RECT 25.995 3.687 26 3.913 ;
      RECT 25.955 3.725 25.995 3.923 ;
      RECT 25.95 3.76 25.955 3.934 ;
      RECT 25.945 3.765 25.95 3.937 ;
      RECT 25.92 3.775 25.945 3.944 ;
      RECT 25.91 3.789 25.92 3.953 ;
      RECT 25.89 3.801 25.91 3.956 ;
      RECT 25.84 3.82 25.89 3.96 ;
      RECT 25.795 3.835 25.84 3.965 ;
      RECT 25.73 3.838 25.795 3.971 ;
      RECT 25.715 3.836 25.73 3.978 ;
      RECT 25.685 3.835 25.715 3.978 ;
      RECT 25.646 3.834 25.685 3.974 ;
      RECT 25.56 3.831 25.646 3.97 ;
      RECT 25.543 3.829 25.56 3.967 ;
      RECT 25.457 3.827 25.543 3.964 ;
      RECT 25.371 3.824 25.457 3.958 ;
      RECT 25.285 3.82 25.371 3.953 ;
      RECT 25.207 3.817 25.285 3.949 ;
      RECT 25.121 3.814 25.207 3.947 ;
      RECT 25.035 3.811 25.121 3.944 ;
      RECT 24.977 3.809 25.035 3.941 ;
      RECT 24.891 3.806 24.977 3.939 ;
      RECT 24.805 3.802 24.891 3.937 ;
      RECT 24.719 3.799 24.805 3.934 ;
      RECT 24.633 3.795 24.719 3.932 ;
      RECT 24.547 3.791 24.633 3.929 ;
      RECT 24.461 3.788 24.547 3.927 ;
      RECT 24.375 3.784 24.461 3.924 ;
      RECT 24.289 3.781 24.375 3.922 ;
      RECT 24.203 3.777 24.289 3.919 ;
      RECT 24.117 3.774 24.203 3.917 ;
      RECT 24.031 3.77 24.117 3.914 ;
      RECT 23.945 3.767 24.031 3.912 ;
      RECT 23.935 3.765 23.945 3.908 ;
      RECT 23.93 3.765 23.935 3.906 ;
      RECT 23.89 3.76 23.93 3.9 ;
      RECT 23.876 3.751 23.89 3.893 ;
      RECT 23.79 3.721 23.876 3.878 ;
      RECT 23.77 3.687 23.79 3.863 ;
      RECT 23.7 3.656 23.77 3.85 ;
      RECT 23.695 3.631 23.7 3.839 ;
      RECT 23.69 3.625 23.695 3.837 ;
      RECT 23.621 3.47 23.69 3.825 ;
      RECT 23.535 3.47 23.621 3.799 ;
      RECT 23.51 3.47 23.535 3.778 ;
      RECT 23.505 3.47 23.51 3.768 ;
      RECT 23.5 3.47 23.505 3.76 ;
      RECT 23.48 3.47 23.5 3.743 ;
      RECT 25.9 2.04 26.16 2.3 ;
      RECT 25.885 2.04 26.16 2.203 ;
      RECT 25.855 2.04 26.16 2.178 ;
      RECT 25.82 1.88 26.1 2.16 ;
      RECT 25.79 3.37 25.85 3.63 ;
      RECT 24.815 2.06 24.87 2.32 ;
      RECT 25.75 3.327 25.79 3.63 ;
      RECT 25.721 3.248 25.75 3.63 ;
      RECT 25.635 3.12 25.721 3.63 ;
      RECT 25.615 3 25.635 3.63 ;
      RECT 25.59 2.951 25.615 3.63 ;
      RECT 25.585 2.916 25.59 3.48 ;
      RECT 25.555 2.876 25.585 3.418 ;
      RECT 25.53 2.813 25.555 3.333 ;
      RECT 25.52 2.775 25.53 3.27 ;
      RECT 25.505 2.75 25.52 3.231 ;
      RECT 25.462 2.708 25.505 3.137 ;
      RECT 25.46 2.681 25.462 3.064 ;
      RECT 25.455 2.676 25.46 3.055 ;
      RECT 25.45 2.669 25.455 3.03 ;
      RECT 25.445 2.663 25.45 3.015 ;
      RECT 25.44 2.657 25.445 3.003 ;
      RECT 25.43 2.648 25.44 2.985 ;
      RECT 25.425 2.639 25.43 2.963 ;
      RECT 25.4 2.62 25.425 2.913 ;
      RECT 25.395 2.601 25.4 2.863 ;
      RECT 25.38 2.587 25.395 2.823 ;
      RECT 25.375 2.573 25.38 2.79 ;
      RECT 25.37 2.566 25.375 2.783 ;
      RECT 25.355 2.553 25.37 2.775 ;
      RECT 25.31 2.515 25.355 2.748 ;
      RECT 25.28 2.468 25.31 2.713 ;
      RECT 25.26 2.437 25.28 2.69 ;
      RECT 25.18 2.37 25.26 2.643 ;
      RECT 25.15 2.3 25.18 2.59 ;
      RECT 25.145 2.277 25.15 2.573 ;
      RECT 25.115 2.255 25.145 2.558 ;
      RECT 25.085 2.214 25.115 2.53 ;
      RECT 25.08 2.189 25.085 2.515 ;
      RECT 25.075 2.183 25.08 2.508 ;
      RECT 25.065 2.06 25.075 2.5 ;
      RECT 25.055 2.06 25.065 2.493 ;
      RECT 25.05 2.06 25.055 2.485 ;
      RECT 25.03 2.06 25.05 2.473 ;
      RECT 24.98 2.06 25.03 2.443 ;
      RECT 24.925 2.06 24.98 2.393 ;
      RECT 24.895 2.06 24.925 2.353 ;
      RECT 24.87 2.06 24.895 2.33 ;
      RECT 24.74 2.785 25.02 3.065 ;
      RECT 24.705 2.7 24.965 2.96 ;
      RECT 24.705 2.782 24.975 2.96 ;
      RECT 22.905 2.155 22.91 2.64 ;
      RECT 22.795 2.34 22.8 2.64 ;
      RECT 22.705 2.38 22.77 2.64 ;
      RECT 24.38 1.88 24.47 2.51 ;
      RECT 24.345 1.93 24.35 2.51 ;
      RECT 24.29 1.955 24.3 2.51 ;
      RECT 24.245 1.955 24.255 2.51 ;
      RECT 24.615 1.88 24.66 2.16 ;
      RECT 23.465 1.61 23.665 1.75 ;
      RECT 24.581 1.88 24.615 2.172 ;
      RECT 24.495 1.88 24.581 2.212 ;
      RECT 24.48 1.88 24.495 2.253 ;
      RECT 24.475 1.88 24.48 2.273 ;
      RECT 24.47 1.88 24.475 2.293 ;
      RECT 24.35 1.922 24.38 2.51 ;
      RECT 24.3 1.942 24.345 2.51 ;
      RECT 24.285 1.957 24.29 2.51 ;
      RECT 24.255 1.957 24.285 2.51 ;
      RECT 24.21 1.942 24.245 2.51 ;
      RECT 24.205 1.93 24.21 2.29 ;
      RECT 24.2 1.927 24.205 2.27 ;
      RECT 24.185 1.917 24.2 2.223 ;
      RECT 24.18 1.91 24.185 2.186 ;
      RECT 24.175 1.907 24.18 2.169 ;
      RECT 24.16 1.897 24.175 2.125 ;
      RECT 24.155 1.888 24.16 2.085 ;
      RECT 24.15 1.884 24.155 2.07 ;
      RECT 24.14 1.878 24.15 2.053 ;
      RECT 24.1 1.859 24.14 2.028 ;
      RECT 24.095 1.841 24.1 2.008 ;
      RECT 24.085 1.835 24.095 2.003 ;
      RECT 24.055 1.819 24.085 1.99 ;
      RECT 24.04 1.801 24.055 1.973 ;
      RECT 24.025 1.789 24.04 1.96 ;
      RECT 24.02 1.781 24.025 1.953 ;
      RECT 23.99 1.767 24.02 1.94 ;
      RECT 23.985 1.752 23.99 1.928 ;
      RECT 23.975 1.746 23.985 1.92 ;
      RECT 23.955 1.734 23.975 1.908 ;
      RECT 23.945 1.722 23.955 1.895 ;
      RECT 23.915 1.706 23.945 1.88 ;
      RECT 23.895 1.686 23.915 1.863 ;
      RECT 23.89 1.676 23.895 1.853 ;
      RECT 23.865 1.664 23.89 1.84 ;
      RECT 23.86 1.652 23.865 1.828 ;
      RECT 23.855 1.647 23.86 1.824 ;
      RECT 23.84 1.64 23.855 1.816 ;
      RECT 23.83 1.627 23.84 1.806 ;
      RECT 23.825 1.625 23.83 1.8 ;
      RECT 23.8 1.618 23.825 1.789 ;
      RECT 23.795 1.611 23.8 1.778 ;
      RECT 23.77 1.61 23.795 1.765 ;
      RECT 23.751 1.61 23.77 1.755 ;
      RECT 23.665 1.61 23.751 1.752 ;
      RECT 23.435 1.61 23.465 1.755 ;
      RECT 23.395 1.617 23.435 1.768 ;
      RECT 23.37 1.627 23.395 1.781 ;
      RECT 23.355 1.636 23.37 1.791 ;
      RECT 23.325 1.641 23.355 1.81 ;
      RECT 23.32 1.647 23.325 1.828 ;
      RECT 23.3 1.657 23.32 1.843 ;
      RECT 23.29 1.67 23.3 1.863 ;
      RECT 23.275 1.682 23.29 1.88 ;
      RECT 23.27 1.692 23.275 1.89 ;
      RECT 23.265 1.697 23.27 1.895 ;
      RECT 23.255 1.705 23.265 1.908 ;
      RECT 23.205 1.737 23.255 1.945 ;
      RECT 23.19 1.772 23.205 1.986 ;
      RECT 23.185 1.782 23.19 2.001 ;
      RECT 23.18 1.787 23.185 2.008 ;
      RECT 23.155 1.803 23.18 2.028 ;
      RECT 23.14 1.824 23.155 2.053 ;
      RECT 23.115 1.845 23.14 2.078 ;
      RECT 23.105 1.864 23.115 2.101 ;
      RECT 23.08 1.882 23.105 2.124 ;
      RECT 23.065 1.902 23.08 2.148 ;
      RECT 23.06 1.912 23.065 2.16 ;
      RECT 23.045 1.924 23.06 2.18 ;
      RECT 23.035 1.939 23.045 2.22 ;
      RECT 23.03 1.947 23.035 2.248 ;
      RECT 23.02 1.957 23.03 2.268 ;
      RECT 23.015 1.97 23.02 2.293 ;
      RECT 23.01 1.983 23.015 2.313 ;
      RECT 23.005 1.989 23.01 2.335 ;
      RECT 22.995 1.998 23.005 2.355 ;
      RECT 22.99 2.018 22.995 2.378 ;
      RECT 22.985 2.024 22.99 2.398 ;
      RECT 22.98 2.031 22.985 2.42 ;
      RECT 22.975 2.042 22.98 2.433 ;
      RECT 22.965 2.052 22.975 2.458 ;
      RECT 22.945 2.077 22.965 2.64 ;
      RECT 22.915 2.117 22.945 2.64 ;
      RECT 22.91 2.147 22.915 2.64 ;
      RECT 22.885 2.175 22.905 2.64 ;
      RECT 22.855 2.22 22.885 2.64 ;
      RECT 22.85 2.247 22.855 2.64 ;
      RECT 22.83 2.265 22.85 2.64 ;
      RECT 22.82 2.29 22.83 2.64 ;
      RECT 22.815 2.302 22.82 2.64 ;
      RECT 22.8 2.325 22.815 2.64 ;
      RECT 22.78 2.352 22.795 2.64 ;
      RECT 22.77 2.375 22.78 2.64 ;
      RECT 24.56 3.26 24.64 3.52 ;
      RECT 23.795 2.48 23.865 2.74 ;
      RECT 24.526 3.227 24.56 3.52 ;
      RECT 24.44 3.13 24.526 3.52 ;
      RECT 24.42 3.042 24.44 3.52 ;
      RECT 24.41 3.012 24.42 3.52 ;
      RECT 24.4 2.992 24.41 3.52 ;
      RECT 24.38 2.979 24.4 3.52 ;
      RECT 24.365 2.969 24.38 3.348 ;
      RECT 24.36 2.962 24.365 3.303 ;
      RECT 24.35 2.956 24.36 3.293 ;
      RECT 24.34 2.948 24.35 3.275 ;
      RECT 24.335 2.942 24.34 3.263 ;
      RECT 24.325 2.937 24.335 3.25 ;
      RECT 24.305 2.927 24.325 3.223 ;
      RECT 24.265 2.906 24.305 3.175 ;
      RECT 24.25 2.887 24.265 3.133 ;
      RECT 24.225 2.873 24.25 3.103 ;
      RECT 24.215 2.861 24.225 3.07 ;
      RECT 24.21 2.856 24.215 3.06 ;
      RECT 24.18 2.842 24.21 3.04 ;
      RECT 24.17 2.826 24.18 3.013 ;
      RECT 24.165 2.821 24.17 3.003 ;
      RECT 24.14 2.812 24.165 2.983 ;
      RECT 24.13 2.8 24.14 2.963 ;
      RECT 24.06 2.768 24.13 2.938 ;
      RECT 24.055 2.737 24.06 2.915 ;
      RECT 24.006 2.48 24.055 2.898 ;
      RECT 23.92 2.48 24.006 2.857 ;
      RECT 23.865 2.48 23.92 2.785 ;
      RECT 23.955 3.265 24.115 3.525 ;
      RECT 23.48 1.88 23.53 2.565 ;
      RECT 23.27 2.305 23.305 2.565 ;
      RECT 23.585 1.88 23.59 2.34 ;
      RECT 23.675 1.88 23.7 2.16 ;
      RECT 23.95 3.262 23.955 3.525 ;
      RECT 23.915 3.25 23.95 3.525 ;
      RECT 23.855 3.223 23.915 3.525 ;
      RECT 23.85 3.206 23.855 3.379 ;
      RECT 23.845 3.203 23.85 3.366 ;
      RECT 23.825 3.196 23.845 3.353 ;
      RECT 23.79 3.179 23.825 3.335 ;
      RECT 23.75 3.158 23.79 3.315 ;
      RECT 23.745 3.146 23.75 3.303 ;
      RECT 23.705 3.132 23.745 3.289 ;
      RECT 23.685 3.115 23.705 3.271 ;
      RECT 23.675 3.107 23.685 3.263 ;
      RECT 23.66 1.88 23.675 2.178 ;
      RECT 23.645 3.097 23.675 3.25 ;
      RECT 23.63 1.88 23.66 2.223 ;
      RECT 23.635 3.087 23.645 3.237 ;
      RECT 23.605 3.072 23.635 3.224 ;
      RECT 23.59 1.88 23.63 2.29 ;
      RECT 23.59 3.04 23.605 3.21 ;
      RECT 23.585 3.012 23.59 3.204 ;
      RECT 23.58 1.88 23.585 2.345 ;
      RECT 23.57 2.982 23.585 3.198 ;
      RECT 23.575 1.88 23.58 2.358 ;
      RECT 23.565 1.88 23.575 2.378 ;
      RECT 23.53 2.895 23.57 3.183 ;
      RECT 23.53 1.88 23.565 2.418 ;
      RECT 23.525 2.827 23.53 3.171 ;
      RECT 23.51 2.782 23.525 3.166 ;
      RECT 23.505 2.72 23.51 3.161 ;
      RECT 23.48 2.627 23.505 3.154 ;
      RECT 23.475 1.88 23.48 3.146 ;
      RECT 23.46 1.88 23.475 3.133 ;
      RECT 23.44 1.88 23.46 3.09 ;
      RECT 23.43 1.88 23.44 3.04 ;
      RECT 23.425 1.88 23.43 3.013 ;
      RECT 23.42 1.88 23.425 2.991 ;
      RECT 23.415 2.106 23.42 2.974 ;
      RECT 23.41 2.128 23.415 2.952 ;
      RECT 23.405 2.17 23.41 2.935 ;
      RECT 23.375 2.22 23.405 2.879 ;
      RECT 23.37 2.247 23.375 2.821 ;
      RECT 23.355 2.265 23.37 2.785 ;
      RECT 23.35 2.283 23.355 2.749 ;
      RECT 23.344 2.29 23.35 2.73 ;
      RECT 23.34 2.297 23.344 2.713 ;
      RECT 23.335 2.302 23.34 2.682 ;
      RECT 23.325 2.305 23.335 2.657 ;
      RECT 23.315 2.305 23.325 2.623 ;
      RECT 23.31 2.305 23.315 2.6 ;
      RECT 23.305 2.305 23.31 2.58 ;
      RECT 22.22 2.44 22.5 2.72 ;
      RECT 22.22 2.44 22.52 2.615 ;
      RECT 22.31 2.33 22.57 2.59 ;
      RECT 22.275 2.425 22.57 2.59 ;
      RECT 22.4 0.945 22.565 2.59 ;
      RECT 22.3 0.945 22.67 1.315 ;
      RECT 21.925 3.47 22.185 3.73 ;
      RECT 21.945 3.397 22.125 3.73 ;
      RECT 21.945 3.14 22.12 3.73 ;
      RECT 21.945 2.932 22.11 3.73 ;
      RECT 21.95 2.85 22.11 3.73 ;
      RECT 21.95 2.615 22.1 3.73 ;
      RECT 21.95 2.462 22.095 3.73 ;
      RECT 21.955 2.447 22.095 3.73 ;
      RECT 22.005 2.162 22.095 3.73 ;
      RECT 21.96 2.397 22.095 3.73 ;
      RECT 21.99 2.215 22.095 3.73 ;
      RECT 21.975 2.327 22.095 3.73 ;
      RECT 21.98 2.285 22.095 3.73 ;
      RECT 21.975 2.327 22.11 2.39 ;
      RECT 22.01 1.915 22.115 2.335 ;
      RECT 22.01 1.915 22.13 2.318 ;
      RECT 22.01 1.915 22.165 2.28 ;
      RECT 22.005 2.162 22.215 2.213 ;
      RECT 22.01 1.915 22.27 2.175 ;
      RECT 21.27 2.62 21.53 2.88 ;
      RECT 21.27 2.62 21.54 2.838 ;
      RECT 21.27 2.62 21.626 2.809 ;
      RECT 21.27 2.62 21.695 2.761 ;
      RECT 21.27 2.62 21.73 2.73 ;
      RECT 21.5 2.44 21.78 2.72 ;
      RECT 21.335 2.605 21.78 2.72 ;
      RECT 21.425 2.482 21.53 2.88 ;
      RECT 21.355 2.545 21.78 2.72 ;
      RECT 15.805 6.22 16.125 6.545 ;
      RECT 15.835 5.695 16.005 6.545 ;
      RECT 15.835 5.695 16.01 6.045 ;
      RECT 15.835 5.695 16.81 5.87 ;
      RECT 16.635 1.965 16.81 5.87 ;
      RECT 16.58 1.965 16.93 2.315 ;
      RECT 16.605 6.655 16.93 6.98 ;
      RECT 15.49 6.745 16.93 6.915 ;
      RECT 15.49 2.395 15.65 6.915 ;
      RECT 15.805 2.365 16.125 2.685 ;
      RECT 15.49 2.395 16.125 2.565 ;
      RECT 14.155 2.705 14.54 3.055 ;
      RECT 14.145 2.77 14.54 2.97 ;
      RECT 14.29 2.7 14.46 3.055 ;
      RECT 12.6 2.44 12.88 2.72 ;
      RECT 12.595 2.44 12.88 2.673 ;
      RECT 12.575 2.44 12.88 2.65 ;
      RECT 12.565 2.44 12.88 2.63 ;
      RECT 12.555 2.44 12.88 2.615 ;
      RECT 12.53 2.44 12.88 2.588 ;
      RECT 12.52 2.44 12.88 2.563 ;
      RECT 12.475 2.295 12.755 2.555 ;
      RECT 12.475 2.39 12.855 2.555 ;
      RECT 12.475 2.335 12.8 2.555 ;
      RECT 12.475 2.327 12.795 2.555 ;
      RECT 12.475 2.317 12.79 2.555 ;
      RECT 12.475 2.305 12.785 2.555 ;
      RECT 11.4 3 11.68 3.28 ;
      RECT 11.4 3 11.715 3.26 ;
      RECT 3.02 6.995 3.31 7.345 ;
      RECT 3.02 7.07 4.385 7.24 ;
      RECT 4.215 6.685 4.385 7.24 ;
      RECT 11.145 6.605 11.495 6.955 ;
      RECT 4.215 6.685 11.495 6.855 ;
      RECT 11.435 2.42 11.485 2.68 ;
      RECT 11.225 2.42 11.23 2.68 ;
      RECT 10.42 1.975 10.45 2.235 ;
      RECT 10.19 1.975 10.265 2.235 ;
      RECT 11.41 2.37 11.435 2.68 ;
      RECT 11.405 2.327 11.41 2.68 ;
      RECT 11.4 2.31 11.405 2.68 ;
      RECT 11.395 2.297 11.4 2.68 ;
      RECT 11.32 2.18 11.395 2.68 ;
      RECT 11.275 1.997 11.32 2.68 ;
      RECT 11.27 1.925 11.275 2.68 ;
      RECT 11.255 1.9 11.27 2.68 ;
      RECT 11.23 1.862 11.255 2.68 ;
      RECT 11.22 1.842 11.23 2.402 ;
      RECT 11.205 1.834 11.22 2.357 ;
      RECT 11.2 1.826 11.205 2.328 ;
      RECT 11.195 1.823 11.2 2.308 ;
      RECT 11.19 1.82 11.195 2.288 ;
      RECT 11.185 1.817 11.19 2.268 ;
      RECT 11.155 1.806 11.185 2.205 ;
      RECT 11.135 1.791 11.155 2.12 ;
      RECT 11.13 1.783 11.135 2.083 ;
      RECT 11.12 1.777 11.13 2.05 ;
      RECT 11.105 1.769 11.12 2.01 ;
      RECT 11.1 1.762 11.105 1.97 ;
      RECT 11.095 1.759 11.1 1.948 ;
      RECT 11.09 1.756 11.095 1.935 ;
      RECT 11.085 1.755 11.09 1.925 ;
      RECT 11.07 1.749 11.085 1.915 ;
      RECT 11.045 1.736 11.07 1.9 ;
      RECT 10.995 1.711 11.045 1.871 ;
      RECT 10.98 1.69 10.995 1.846 ;
      RECT 10.97 1.683 10.98 1.835 ;
      RECT 10.915 1.664 10.97 1.808 ;
      RECT 10.89 1.642 10.915 1.781 ;
      RECT 10.885 1.635 10.89 1.776 ;
      RECT 10.87 1.635 10.885 1.774 ;
      RECT 10.845 1.627 10.87 1.77 ;
      RECT 10.83 1.625 10.845 1.766 ;
      RECT 10.8 1.625 10.83 1.763 ;
      RECT 10.79 1.625 10.8 1.758 ;
      RECT 10.745 1.625 10.79 1.756 ;
      RECT 10.716 1.625 10.745 1.757 ;
      RECT 10.63 1.625 10.716 1.759 ;
      RECT 10.616 1.626 10.63 1.761 ;
      RECT 10.53 1.627 10.616 1.763 ;
      RECT 10.515 1.628 10.53 1.773 ;
      RECT 10.51 1.629 10.515 1.782 ;
      RECT 10.49 1.632 10.51 1.792 ;
      RECT 10.475 1.64 10.49 1.807 ;
      RECT 10.455 1.658 10.475 1.822 ;
      RECT 10.445 1.67 10.455 1.845 ;
      RECT 10.435 1.679 10.445 1.875 ;
      RECT 10.42 1.691 10.435 1.92 ;
      RECT 10.365 1.724 10.42 2.235 ;
      RECT 10.36 1.752 10.365 2.235 ;
      RECT 10.34 1.767 10.36 2.235 ;
      RECT 10.305 1.827 10.34 2.235 ;
      RECT 10.303 1.877 10.305 2.235 ;
      RECT 10.3 1.885 10.303 2.235 ;
      RECT 10.29 1.9 10.3 2.235 ;
      RECT 10.285 1.912 10.29 2.235 ;
      RECT 10.275 1.937 10.285 2.235 ;
      RECT 10.265 1.965 10.275 2.235 ;
      RECT 8.17 3.47 8.22 3.73 ;
      RECT 11.08 3.02 11.14 3.28 ;
      RECT 11.065 3.02 11.08 3.29 ;
      RECT 11.046 3.02 11.065 3.323 ;
      RECT 10.96 3.02 11.046 3.448 ;
      RECT 10.88 3.02 10.96 3.63 ;
      RECT 10.875 3.257 10.88 3.715 ;
      RECT 10.85 3.327 10.875 3.743 ;
      RECT 10.845 3.397 10.85 3.77 ;
      RECT 10.825 3.469 10.845 3.792 ;
      RECT 10.82 3.536 10.825 3.815 ;
      RECT 10.81 3.565 10.82 3.83 ;
      RECT 10.8 3.587 10.81 3.847 ;
      RECT 10.795 3.597 10.8 3.858 ;
      RECT 10.79 3.605 10.795 3.866 ;
      RECT 10.78 3.613 10.79 3.878 ;
      RECT 10.775 3.625 10.78 3.888 ;
      RECT 10.77 3.633 10.775 3.893 ;
      RECT 10.75 3.651 10.77 3.903 ;
      RECT 10.745 3.668 10.75 3.91 ;
      RECT 10.74 3.676 10.745 3.911 ;
      RECT 10.735 3.687 10.74 3.913 ;
      RECT 10.695 3.725 10.735 3.923 ;
      RECT 10.69 3.76 10.695 3.934 ;
      RECT 10.685 3.765 10.69 3.937 ;
      RECT 10.66 3.775 10.685 3.944 ;
      RECT 10.65 3.789 10.66 3.953 ;
      RECT 10.63 3.801 10.65 3.956 ;
      RECT 10.58 3.82 10.63 3.96 ;
      RECT 10.535 3.835 10.58 3.965 ;
      RECT 10.47 3.838 10.535 3.971 ;
      RECT 10.455 3.836 10.47 3.978 ;
      RECT 10.425 3.835 10.455 3.978 ;
      RECT 10.386 3.834 10.425 3.974 ;
      RECT 10.3 3.831 10.386 3.97 ;
      RECT 10.283 3.829 10.3 3.967 ;
      RECT 10.197 3.827 10.283 3.964 ;
      RECT 10.111 3.824 10.197 3.958 ;
      RECT 10.025 3.82 10.111 3.953 ;
      RECT 9.947 3.817 10.025 3.949 ;
      RECT 9.861 3.814 9.947 3.947 ;
      RECT 9.775 3.811 9.861 3.944 ;
      RECT 9.717 3.809 9.775 3.941 ;
      RECT 9.631 3.806 9.717 3.939 ;
      RECT 9.545 3.802 9.631 3.937 ;
      RECT 9.459 3.799 9.545 3.934 ;
      RECT 9.373 3.795 9.459 3.932 ;
      RECT 9.287 3.791 9.373 3.929 ;
      RECT 9.201 3.788 9.287 3.927 ;
      RECT 9.115 3.784 9.201 3.924 ;
      RECT 9.029 3.781 9.115 3.922 ;
      RECT 8.943 3.777 9.029 3.919 ;
      RECT 8.857 3.774 8.943 3.917 ;
      RECT 8.771 3.77 8.857 3.914 ;
      RECT 8.685 3.767 8.771 3.912 ;
      RECT 8.675 3.765 8.685 3.908 ;
      RECT 8.67 3.765 8.675 3.906 ;
      RECT 8.63 3.76 8.67 3.9 ;
      RECT 8.616 3.751 8.63 3.893 ;
      RECT 8.53 3.721 8.616 3.878 ;
      RECT 8.51 3.687 8.53 3.863 ;
      RECT 8.44 3.656 8.51 3.85 ;
      RECT 8.435 3.631 8.44 3.839 ;
      RECT 8.43 3.625 8.435 3.837 ;
      RECT 8.361 3.47 8.43 3.825 ;
      RECT 8.275 3.47 8.361 3.799 ;
      RECT 8.25 3.47 8.275 3.778 ;
      RECT 8.245 3.47 8.25 3.768 ;
      RECT 8.24 3.47 8.245 3.76 ;
      RECT 8.22 3.47 8.24 3.743 ;
      RECT 10.64 2.04 10.9 2.3 ;
      RECT 10.625 2.04 10.9 2.203 ;
      RECT 10.595 2.04 10.9 2.178 ;
      RECT 10.56 1.88 10.84 2.16 ;
      RECT 10.53 3.37 10.59 3.63 ;
      RECT 9.555 2.06 9.61 2.32 ;
      RECT 10.49 3.327 10.53 3.63 ;
      RECT 10.461 3.248 10.49 3.63 ;
      RECT 10.375 3.12 10.461 3.63 ;
      RECT 10.355 3 10.375 3.63 ;
      RECT 10.33 2.951 10.355 3.63 ;
      RECT 10.325 2.916 10.33 3.48 ;
      RECT 10.295 2.876 10.325 3.418 ;
      RECT 10.27 2.813 10.295 3.333 ;
      RECT 10.26 2.775 10.27 3.27 ;
      RECT 10.245 2.75 10.26 3.231 ;
      RECT 10.202 2.708 10.245 3.137 ;
      RECT 10.2 2.681 10.202 3.064 ;
      RECT 10.195 2.676 10.2 3.055 ;
      RECT 10.19 2.669 10.195 3.03 ;
      RECT 10.185 2.663 10.19 3.015 ;
      RECT 10.18 2.657 10.185 3.003 ;
      RECT 10.17 2.648 10.18 2.985 ;
      RECT 10.165 2.639 10.17 2.963 ;
      RECT 10.14 2.62 10.165 2.913 ;
      RECT 10.135 2.601 10.14 2.863 ;
      RECT 10.12 2.587 10.135 2.823 ;
      RECT 10.115 2.573 10.12 2.79 ;
      RECT 10.11 2.566 10.115 2.783 ;
      RECT 10.095 2.553 10.11 2.775 ;
      RECT 10.05 2.515 10.095 2.748 ;
      RECT 10.02 2.468 10.05 2.713 ;
      RECT 10 2.437 10.02 2.69 ;
      RECT 9.92 2.37 10 2.643 ;
      RECT 9.89 2.3 9.92 2.59 ;
      RECT 9.885 2.277 9.89 2.573 ;
      RECT 9.855 2.255 9.885 2.558 ;
      RECT 9.825 2.214 9.855 2.53 ;
      RECT 9.82 2.189 9.825 2.515 ;
      RECT 9.815 2.183 9.82 2.508 ;
      RECT 9.805 2.06 9.815 2.5 ;
      RECT 9.795 2.06 9.805 2.493 ;
      RECT 9.79 2.06 9.795 2.485 ;
      RECT 9.77 2.06 9.79 2.473 ;
      RECT 9.72 2.06 9.77 2.443 ;
      RECT 9.665 2.06 9.72 2.393 ;
      RECT 9.635 2.06 9.665 2.353 ;
      RECT 9.61 2.06 9.635 2.33 ;
      RECT 9.48 2.785 9.76 3.065 ;
      RECT 9.445 2.7 9.705 2.96 ;
      RECT 9.445 2.782 9.715 2.96 ;
      RECT 7.645 2.155 7.65 2.64 ;
      RECT 7.535 2.34 7.54 2.64 ;
      RECT 7.445 2.38 7.51 2.64 ;
      RECT 9.12 1.88 9.21 2.51 ;
      RECT 9.085 1.93 9.09 2.51 ;
      RECT 9.03 1.955 9.04 2.51 ;
      RECT 8.985 1.955 8.995 2.51 ;
      RECT 9.355 1.88 9.4 2.16 ;
      RECT 8.205 1.61 8.405 1.75 ;
      RECT 9.321 1.88 9.355 2.172 ;
      RECT 9.235 1.88 9.321 2.212 ;
      RECT 9.22 1.88 9.235 2.253 ;
      RECT 9.215 1.88 9.22 2.273 ;
      RECT 9.21 1.88 9.215 2.293 ;
      RECT 9.09 1.922 9.12 2.51 ;
      RECT 9.04 1.942 9.085 2.51 ;
      RECT 9.025 1.957 9.03 2.51 ;
      RECT 8.995 1.957 9.025 2.51 ;
      RECT 8.95 1.942 8.985 2.51 ;
      RECT 8.945 1.93 8.95 2.29 ;
      RECT 8.94 1.927 8.945 2.27 ;
      RECT 8.925 1.917 8.94 2.223 ;
      RECT 8.92 1.91 8.925 2.186 ;
      RECT 8.915 1.907 8.92 2.169 ;
      RECT 8.9 1.897 8.915 2.125 ;
      RECT 8.895 1.888 8.9 2.085 ;
      RECT 8.89 1.884 8.895 2.07 ;
      RECT 8.88 1.878 8.89 2.053 ;
      RECT 8.84 1.859 8.88 2.028 ;
      RECT 8.835 1.841 8.84 2.008 ;
      RECT 8.825 1.835 8.835 2.003 ;
      RECT 8.795 1.819 8.825 1.99 ;
      RECT 8.78 1.801 8.795 1.973 ;
      RECT 8.765 1.789 8.78 1.96 ;
      RECT 8.76 1.781 8.765 1.953 ;
      RECT 8.73 1.767 8.76 1.94 ;
      RECT 8.725 1.752 8.73 1.928 ;
      RECT 8.715 1.746 8.725 1.92 ;
      RECT 8.695 1.734 8.715 1.908 ;
      RECT 8.685 1.722 8.695 1.895 ;
      RECT 8.655 1.706 8.685 1.88 ;
      RECT 8.635 1.686 8.655 1.863 ;
      RECT 8.63 1.676 8.635 1.853 ;
      RECT 8.605 1.664 8.63 1.84 ;
      RECT 8.6 1.652 8.605 1.828 ;
      RECT 8.595 1.647 8.6 1.824 ;
      RECT 8.58 1.64 8.595 1.816 ;
      RECT 8.57 1.627 8.58 1.806 ;
      RECT 8.565 1.625 8.57 1.8 ;
      RECT 8.54 1.618 8.565 1.789 ;
      RECT 8.535 1.611 8.54 1.778 ;
      RECT 8.51 1.61 8.535 1.765 ;
      RECT 8.491 1.61 8.51 1.755 ;
      RECT 8.405 1.61 8.491 1.752 ;
      RECT 8.175 1.61 8.205 1.755 ;
      RECT 8.135 1.617 8.175 1.768 ;
      RECT 8.11 1.627 8.135 1.781 ;
      RECT 8.095 1.636 8.11 1.791 ;
      RECT 8.065 1.641 8.095 1.81 ;
      RECT 8.06 1.647 8.065 1.828 ;
      RECT 8.04 1.657 8.06 1.843 ;
      RECT 8.03 1.67 8.04 1.863 ;
      RECT 8.015 1.682 8.03 1.88 ;
      RECT 8.01 1.692 8.015 1.89 ;
      RECT 8.005 1.697 8.01 1.895 ;
      RECT 7.995 1.705 8.005 1.908 ;
      RECT 7.945 1.737 7.995 1.945 ;
      RECT 7.93 1.772 7.945 1.986 ;
      RECT 7.925 1.782 7.93 2.001 ;
      RECT 7.92 1.787 7.925 2.008 ;
      RECT 7.895 1.803 7.92 2.028 ;
      RECT 7.88 1.824 7.895 2.053 ;
      RECT 7.855 1.845 7.88 2.078 ;
      RECT 7.845 1.864 7.855 2.101 ;
      RECT 7.82 1.882 7.845 2.124 ;
      RECT 7.805 1.902 7.82 2.148 ;
      RECT 7.8 1.912 7.805 2.16 ;
      RECT 7.785 1.924 7.8 2.18 ;
      RECT 7.775 1.939 7.785 2.22 ;
      RECT 7.77 1.947 7.775 2.248 ;
      RECT 7.76 1.957 7.77 2.268 ;
      RECT 7.755 1.97 7.76 2.293 ;
      RECT 7.75 1.983 7.755 2.313 ;
      RECT 7.745 1.989 7.75 2.335 ;
      RECT 7.735 1.998 7.745 2.355 ;
      RECT 7.73 2.018 7.735 2.378 ;
      RECT 7.725 2.024 7.73 2.398 ;
      RECT 7.72 2.031 7.725 2.42 ;
      RECT 7.715 2.042 7.72 2.433 ;
      RECT 7.705 2.052 7.715 2.458 ;
      RECT 7.685 2.077 7.705 2.64 ;
      RECT 7.655 2.117 7.685 2.64 ;
      RECT 7.65 2.147 7.655 2.64 ;
      RECT 7.625 2.175 7.645 2.64 ;
      RECT 7.595 2.22 7.625 2.64 ;
      RECT 7.59 2.247 7.595 2.64 ;
      RECT 7.57 2.265 7.59 2.64 ;
      RECT 7.56 2.29 7.57 2.64 ;
      RECT 7.555 2.302 7.56 2.64 ;
      RECT 7.54 2.325 7.555 2.64 ;
      RECT 7.52 2.352 7.535 2.64 ;
      RECT 7.51 2.375 7.52 2.64 ;
      RECT 9.3 3.26 9.38 3.52 ;
      RECT 8.535 2.48 8.605 2.74 ;
      RECT 9.266 3.227 9.3 3.52 ;
      RECT 9.18 3.13 9.266 3.52 ;
      RECT 9.16 3.042 9.18 3.52 ;
      RECT 9.15 3.012 9.16 3.52 ;
      RECT 9.14 2.992 9.15 3.52 ;
      RECT 9.12 2.979 9.14 3.52 ;
      RECT 9.105 2.969 9.12 3.348 ;
      RECT 9.1 2.962 9.105 3.303 ;
      RECT 9.09 2.956 9.1 3.293 ;
      RECT 9.08 2.948 9.09 3.275 ;
      RECT 9.075 2.942 9.08 3.263 ;
      RECT 9.065 2.937 9.075 3.25 ;
      RECT 9.045 2.927 9.065 3.223 ;
      RECT 9.005 2.906 9.045 3.175 ;
      RECT 8.99 2.887 9.005 3.133 ;
      RECT 8.965 2.873 8.99 3.103 ;
      RECT 8.955 2.861 8.965 3.07 ;
      RECT 8.95 2.856 8.955 3.06 ;
      RECT 8.92 2.842 8.95 3.04 ;
      RECT 8.91 2.826 8.92 3.013 ;
      RECT 8.905 2.821 8.91 3.003 ;
      RECT 8.88 2.812 8.905 2.983 ;
      RECT 8.87 2.8 8.88 2.963 ;
      RECT 8.8 2.768 8.87 2.938 ;
      RECT 8.795 2.737 8.8 2.915 ;
      RECT 8.746 2.48 8.795 2.898 ;
      RECT 8.66 2.48 8.746 2.857 ;
      RECT 8.605 2.48 8.66 2.785 ;
      RECT 8.695 3.265 8.855 3.525 ;
      RECT 8.22 1.88 8.27 2.565 ;
      RECT 8.01 2.305 8.045 2.565 ;
      RECT 8.325 1.88 8.33 2.34 ;
      RECT 8.415 1.88 8.44 2.16 ;
      RECT 8.69 3.262 8.695 3.525 ;
      RECT 8.655 3.25 8.69 3.525 ;
      RECT 8.595 3.223 8.655 3.525 ;
      RECT 8.59 3.206 8.595 3.379 ;
      RECT 8.585 3.203 8.59 3.366 ;
      RECT 8.565 3.196 8.585 3.353 ;
      RECT 8.53 3.179 8.565 3.335 ;
      RECT 8.49 3.158 8.53 3.315 ;
      RECT 8.485 3.146 8.49 3.303 ;
      RECT 8.445 3.132 8.485 3.289 ;
      RECT 8.425 3.115 8.445 3.271 ;
      RECT 8.415 3.107 8.425 3.263 ;
      RECT 8.4 1.88 8.415 2.178 ;
      RECT 8.385 3.097 8.415 3.25 ;
      RECT 8.37 1.88 8.4 2.223 ;
      RECT 8.375 3.087 8.385 3.237 ;
      RECT 8.345 3.072 8.375 3.224 ;
      RECT 8.33 1.88 8.37 2.29 ;
      RECT 8.33 3.04 8.345 3.21 ;
      RECT 8.325 3.012 8.33 3.204 ;
      RECT 8.32 1.88 8.325 2.345 ;
      RECT 8.31 2.982 8.325 3.198 ;
      RECT 8.315 1.88 8.32 2.358 ;
      RECT 8.305 1.88 8.315 2.378 ;
      RECT 8.27 2.895 8.31 3.183 ;
      RECT 8.27 1.88 8.305 2.418 ;
      RECT 8.265 2.827 8.27 3.171 ;
      RECT 8.25 2.782 8.265 3.166 ;
      RECT 8.245 2.72 8.25 3.161 ;
      RECT 8.22 2.627 8.245 3.154 ;
      RECT 8.215 1.88 8.22 3.146 ;
      RECT 8.2 1.88 8.215 3.133 ;
      RECT 8.18 1.88 8.2 3.09 ;
      RECT 8.17 1.88 8.18 3.04 ;
      RECT 8.165 1.88 8.17 3.013 ;
      RECT 8.16 1.88 8.165 2.991 ;
      RECT 8.155 2.106 8.16 2.974 ;
      RECT 8.15 2.128 8.155 2.952 ;
      RECT 8.145 2.17 8.15 2.935 ;
      RECT 8.115 2.22 8.145 2.879 ;
      RECT 8.11 2.247 8.115 2.821 ;
      RECT 8.095 2.265 8.11 2.785 ;
      RECT 8.09 2.283 8.095 2.749 ;
      RECT 8.084 2.29 8.09 2.73 ;
      RECT 8.08 2.297 8.084 2.713 ;
      RECT 8.075 2.302 8.08 2.682 ;
      RECT 8.065 2.305 8.075 2.657 ;
      RECT 8.055 2.305 8.065 2.623 ;
      RECT 8.05 2.305 8.055 2.6 ;
      RECT 8.045 2.305 8.05 2.58 ;
      RECT 6.96 2.44 7.24 2.72 ;
      RECT 6.96 2.44 7.26 2.615 ;
      RECT 7.05 2.33 7.31 2.59 ;
      RECT 7.015 2.425 7.31 2.59 ;
      RECT 7.14 0.945 7.305 2.59 ;
      RECT 7.04 0.945 7.41 1.315 ;
      RECT 6.665 3.47 6.925 3.73 ;
      RECT 6.685 3.397 6.865 3.73 ;
      RECT 6.685 3.14 6.86 3.73 ;
      RECT 6.685 2.932 6.85 3.73 ;
      RECT 6.69 2.85 6.85 3.73 ;
      RECT 6.69 2.615 6.84 3.73 ;
      RECT 6.69 2.462 6.835 3.73 ;
      RECT 6.695 2.447 6.835 3.73 ;
      RECT 6.745 2.162 6.835 3.73 ;
      RECT 6.7 2.397 6.835 3.73 ;
      RECT 6.73 2.215 6.835 3.73 ;
      RECT 6.715 2.327 6.835 3.73 ;
      RECT 6.72 2.285 6.835 3.73 ;
      RECT 6.715 2.327 6.85 2.39 ;
      RECT 6.75 1.915 6.855 2.335 ;
      RECT 6.75 1.915 6.87 2.318 ;
      RECT 6.75 1.915 6.905 2.28 ;
      RECT 6.745 2.162 6.955 2.213 ;
      RECT 6.75 1.915 7.01 2.175 ;
      RECT 6.01 2.62 6.27 2.88 ;
      RECT 6.01 2.62 6.28 2.838 ;
      RECT 6.01 2.62 6.366 2.809 ;
      RECT 6.01 2.62 6.435 2.761 ;
      RECT 6.01 2.62 6.47 2.73 ;
      RECT 6.24 2.44 6.52 2.72 ;
      RECT 6.075 2.605 6.52 2.72 ;
      RECT 6.165 2.482 6.27 2.88 ;
      RECT 6.095 2.545 6.52 2.72 ;
      RECT 71.515 7.055 71.885 7.425 ;
      RECT 56.255 7.055 56.625 7.425 ;
      RECT 40.995 7.055 41.365 7.425 ;
      RECT 25.735 7.055 26.105 7.425 ;
      RECT 10.475 7.055 10.845 7.425 ;
    LAYER via1 ;
      RECT 80.105 7.375 80.255 7.525 ;
      RECT 77.735 6.74 77.885 6.89 ;
      RECT 77.72 2.065 77.87 2.215 ;
      RECT 76.93 2.45 77.08 2.6 ;
      RECT 76.93 6.325 77.08 6.475 ;
      RECT 75.34 2.805 75.49 2.955 ;
      RECT 73.57 2.35 73.72 2.5 ;
      RECT 72.55 3.055 72.7 3.205 ;
      RECT 72.32 2.475 72.47 2.625 ;
      RECT 72.285 6.71 72.435 6.86 ;
      RECT 71.975 3.075 72.125 3.225 ;
      RECT 71.735 2.095 71.885 2.245 ;
      RECT 71.625 7.165 71.775 7.315 ;
      RECT 71.425 3.425 71.575 3.575 ;
      RECT 71.285 2.03 71.435 2.18 ;
      RECT 70.65 2.115 70.8 2.265 ;
      RECT 70.54 2.755 70.69 2.905 ;
      RECT 70.215 3.315 70.365 3.465 ;
      RECT 70.045 2.305 70.195 2.455 ;
      RECT 69.69 3.32 69.84 3.47 ;
      RECT 69.63 2.535 69.78 2.685 ;
      RECT 69.265 3.525 69.415 3.675 ;
      RECT 69.105 2.36 69.255 2.51 ;
      RECT 68.54 2.435 68.69 2.585 ;
      RECT 68.19 1.055 68.34 1.205 ;
      RECT 68.145 2.385 68.295 2.535 ;
      RECT 67.845 1.97 67.995 2.12 ;
      RECT 67.76 3.525 67.91 3.675 ;
      RECT 67.105 2.675 67.255 2.825 ;
      RECT 64.82 6.755 64.97 6.905 ;
      RECT 62.475 6.74 62.625 6.89 ;
      RECT 62.46 2.065 62.61 2.215 ;
      RECT 61.67 2.45 61.82 2.6 ;
      RECT 61.67 6.325 61.82 6.475 ;
      RECT 60.08 2.805 60.23 2.955 ;
      RECT 58.31 2.35 58.46 2.5 ;
      RECT 57.29 3.055 57.44 3.205 ;
      RECT 57.06 2.475 57.21 2.625 ;
      RECT 57.025 6.71 57.175 6.86 ;
      RECT 56.715 3.075 56.865 3.225 ;
      RECT 56.475 2.095 56.625 2.245 ;
      RECT 56.365 7.165 56.515 7.315 ;
      RECT 56.165 3.425 56.315 3.575 ;
      RECT 56.025 2.03 56.175 2.18 ;
      RECT 55.39 2.115 55.54 2.265 ;
      RECT 55.28 2.755 55.43 2.905 ;
      RECT 54.955 3.315 55.105 3.465 ;
      RECT 54.785 2.305 54.935 2.455 ;
      RECT 54.43 3.32 54.58 3.47 ;
      RECT 54.37 2.535 54.52 2.685 ;
      RECT 54.005 3.525 54.155 3.675 ;
      RECT 53.845 2.36 53.995 2.51 ;
      RECT 53.28 2.435 53.43 2.585 ;
      RECT 52.93 1.055 53.08 1.205 ;
      RECT 52.885 2.385 53.035 2.535 ;
      RECT 52.585 1.97 52.735 2.12 ;
      RECT 52.5 3.525 52.65 3.675 ;
      RECT 51.845 2.675 51.995 2.825 ;
      RECT 49.56 6.755 49.71 6.905 ;
      RECT 47.215 6.74 47.365 6.89 ;
      RECT 47.2 2.065 47.35 2.215 ;
      RECT 46.41 2.45 46.56 2.6 ;
      RECT 46.41 6.325 46.56 6.475 ;
      RECT 44.82 2.805 44.97 2.955 ;
      RECT 43.05 2.35 43.2 2.5 ;
      RECT 42.03 3.055 42.18 3.205 ;
      RECT 41.8 2.475 41.95 2.625 ;
      RECT 41.765 6.715 41.915 6.865 ;
      RECT 41.455 3.075 41.605 3.225 ;
      RECT 41.215 2.095 41.365 2.245 ;
      RECT 41.105 7.165 41.255 7.315 ;
      RECT 40.905 3.425 41.055 3.575 ;
      RECT 40.765 2.03 40.915 2.18 ;
      RECT 40.13 2.115 40.28 2.265 ;
      RECT 40.02 2.755 40.17 2.905 ;
      RECT 39.695 3.315 39.845 3.465 ;
      RECT 39.525 2.305 39.675 2.455 ;
      RECT 39.17 3.32 39.32 3.47 ;
      RECT 39.11 2.535 39.26 2.685 ;
      RECT 38.745 3.525 38.895 3.675 ;
      RECT 38.585 2.36 38.735 2.51 ;
      RECT 38.02 2.435 38.17 2.585 ;
      RECT 37.67 1.055 37.82 1.205 ;
      RECT 37.625 2.385 37.775 2.535 ;
      RECT 37.325 1.97 37.475 2.12 ;
      RECT 37.24 3.525 37.39 3.675 ;
      RECT 36.585 2.675 36.735 2.825 ;
      RECT 34.345 6.76 34.495 6.91 ;
      RECT 31.955 6.74 32.105 6.89 ;
      RECT 31.94 2.065 32.09 2.215 ;
      RECT 31.15 2.45 31.3 2.6 ;
      RECT 31.15 6.325 31.3 6.475 ;
      RECT 29.56 2.805 29.71 2.955 ;
      RECT 27.79 2.35 27.94 2.5 ;
      RECT 26.77 3.055 26.92 3.205 ;
      RECT 26.54 2.475 26.69 2.625 ;
      RECT 26.505 6.71 26.655 6.86 ;
      RECT 26.195 3.075 26.345 3.225 ;
      RECT 25.955 2.095 26.105 2.245 ;
      RECT 25.845 7.165 25.995 7.315 ;
      RECT 25.645 3.425 25.795 3.575 ;
      RECT 25.505 2.03 25.655 2.18 ;
      RECT 24.87 2.115 25.02 2.265 ;
      RECT 24.76 2.755 24.91 2.905 ;
      RECT 24.435 3.315 24.585 3.465 ;
      RECT 24.265 2.305 24.415 2.455 ;
      RECT 23.91 3.32 24.06 3.47 ;
      RECT 23.85 2.535 24 2.685 ;
      RECT 23.485 3.525 23.635 3.675 ;
      RECT 23.325 2.36 23.475 2.51 ;
      RECT 22.76 2.435 22.91 2.585 ;
      RECT 22.41 1.055 22.56 1.205 ;
      RECT 22.365 2.385 22.515 2.535 ;
      RECT 22.065 1.97 22.215 2.12 ;
      RECT 21.98 3.525 22.13 3.675 ;
      RECT 21.325 2.675 21.475 2.825 ;
      RECT 19.085 6.755 19.235 6.905 ;
      RECT 16.695 6.74 16.845 6.89 ;
      RECT 16.68 2.065 16.83 2.215 ;
      RECT 15.89 2.45 16.04 2.6 ;
      RECT 15.89 6.325 16.04 6.475 ;
      RECT 14.3 2.805 14.45 2.955 ;
      RECT 12.53 2.35 12.68 2.5 ;
      RECT 11.51 3.055 11.66 3.205 ;
      RECT 11.28 2.475 11.43 2.625 ;
      RECT 11.245 6.705 11.395 6.855 ;
      RECT 10.935 3.075 11.085 3.225 ;
      RECT 10.695 2.095 10.845 2.245 ;
      RECT 10.585 7.165 10.735 7.315 ;
      RECT 10.385 3.425 10.535 3.575 ;
      RECT 10.245 2.03 10.395 2.18 ;
      RECT 9.61 2.115 9.76 2.265 ;
      RECT 9.5 2.755 9.65 2.905 ;
      RECT 9.175 3.315 9.325 3.465 ;
      RECT 9.005 2.305 9.155 2.455 ;
      RECT 8.65 3.32 8.8 3.47 ;
      RECT 8.59 2.535 8.74 2.685 ;
      RECT 8.225 3.525 8.375 3.675 ;
      RECT 8.065 2.36 8.215 2.51 ;
      RECT 7.5 2.435 7.65 2.585 ;
      RECT 7.15 1.055 7.3 1.205 ;
      RECT 7.105 2.385 7.255 2.535 ;
      RECT 6.805 1.97 6.955 2.12 ;
      RECT 6.72 3.525 6.87 3.675 ;
      RECT 6.065 2.675 6.215 2.825 ;
      RECT 3.09 7.095 3.24 7.245 ;
      RECT 2.715 6.355 2.865 6.505 ;
    LAYER met1 ;
      RECT 66.065 0 74.805 1.74 ;
      RECT 50.805 0 59.545 1.74 ;
      RECT 35.545 0 44.285 1.74 ;
      RECT 20.285 0 29.025 1.74 ;
      RECT 5.025 0 13.765 1.74 ;
      RECT 80.395 0 80.575 0.305 ;
      RECT 65.135 0 78.445 0.305 ;
      RECT 49.875 0 63.185 0.305 ;
      RECT 34.615 0 47.925 0.305 ;
      RECT 19.355 0 32.665 0.305 ;
      RECT 1.48 0 17.405 0.305 ;
      RECT 1.48 0 80.575 0.3 ;
      RECT 1.48 8.58 80.575 8.88 ;
      RECT 80.395 8.575 80.575 8.88 ;
      RECT 65.135 8.575 78.445 8.88 ;
      RECT 49.875 8.575 63.185 8.88 ;
      RECT 34.615 8.575 47.925 8.88 ;
      RECT 19.355 8.575 32.665 8.88 ;
      RECT 1.48 8.575 17.405 8.88 ;
      RECT 71.01 6.315 71.18 8.88 ;
      RECT 55.75 6.315 55.92 8.88 ;
      RECT 40.49 6.315 40.66 8.88 ;
      RECT 25.23 6.315 25.4 8.88 ;
      RECT 9.97 6.315 10.14 8.88 ;
      RECT 71.18 6.285 71.47 6.515 ;
      RECT 55.92 6.285 56.21 6.515 ;
      RECT 40.66 6.285 40.95 6.515 ;
      RECT 25.4 6.285 25.69 6.515 ;
      RECT 10.14 6.285 10.43 6.515 ;
      RECT 79.97 7.77 80.26 8 ;
      RECT 80.03 6.29 80.2 8 ;
      RECT 80.005 7.275 80.355 7.625 ;
      RECT 79.97 6.29 80.26 6.52 ;
      RECT 79.565 2.395 79.67 2.965 ;
      RECT 79.565 2.73 79.89 2.96 ;
      RECT 79.565 2.76 80.06 2.93 ;
      RECT 79.565 2.395 79.755 2.96 ;
      RECT 78.98 2.36 79.27 2.59 ;
      RECT 78.98 2.395 79.755 2.565 ;
      RECT 79.04 0.88 79.21 2.59 ;
      RECT 78.98 0.88 79.27 1.11 ;
      RECT 78.98 7.77 79.27 8 ;
      RECT 79.04 6.29 79.21 8 ;
      RECT 78.98 6.29 79.27 6.52 ;
      RECT 78.98 6.325 79.835 6.485 ;
      RECT 79.665 5.92 79.835 6.485 ;
      RECT 78.98 6.32 79.375 6.485 ;
      RECT 79.6 5.92 79.89 6.15 ;
      RECT 79.6 5.95 80.06 6.12 ;
      RECT 78.61 2.73 78.9 2.96 ;
      RECT 78.61 2.76 79.07 2.93 ;
      RECT 78.675 1.655 78.84 2.96 ;
      RECT 77.19 1.625 77.48 1.855 ;
      RECT 77.19 1.655 78.84 1.825 ;
      RECT 77.25 0.885 77.42 1.855 ;
      RECT 77.19 0.885 77.48 1.115 ;
      RECT 77.19 7.765 77.48 7.995 ;
      RECT 77.25 7.025 77.42 7.995 ;
      RECT 77.25 7.12 78.84 7.29 ;
      RECT 78.67 5.92 78.84 7.29 ;
      RECT 77.19 7.025 77.48 7.255 ;
      RECT 78.61 5.92 78.9 6.15 ;
      RECT 78.61 5.95 79.07 6.12 ;
      RECT 75.24 2.705 75.58 3.055 ;
      RECT 75.33 2.025 75.5 3.055 ;
      RECT 77.62 1.965 77.97 2.315 ;
      RECT 75.33 2.025 77.97 2.195 ;
      RECT 77.645 6.655 77.97 6.98 ;
      RECT 72.185 6.61 72.535 6.96 ;
      RECT 77.62 6.655 77.97 6.885 ;
      RECT 71.985 6.655 72.535 6.885 ;
      RECT 71.815 6.685 77.97 6.855 ;
      RECT 76.845 2.365 77.165 2.685 ;
      RECT 76.815 2.365 77.165 2.595 ;
      RECT 76.645 2.395 77.165 2.565 ;
      RECT 76.845 6.255 77.165 6.545 ;
      RECT 76.815 6.285 77.165 6.515 ;
      RECT 76.645 6.315 77.165 6.485 ;
      RECT 72.535 2.985 72.685 3.26 ;
      RECT 73.075 2.065 73.08 2.285 ;
      RECT 74.225 2.265 74.24 2.463 ;
      RECT 74.19 2.257 74.225 2.47 ;
      RECT 74.16 2.25 74.19 2.47 ;
      RECT 74.105 2.215 74.16 2.47 ;
      RECT 74.04 2.152 74.105 2.47 ;
      RECT 74.035 2.117 74.04 2.468 ;
      RECT 74.03 2.112 74.035 2.46 ;
      RECT 74.025 2.107 74.03 2.446 ;
      RECT 74.02 2.104 74.025 2.439 ;
      RECT 73.975 2.094 74.02 2.39 ;
      RECT 73.955 2.081 73.975 2.325 ;
      RECT 73.95 2.076 73.955 2.298 ;
      RECT 73.945 2.075 73.95 2.291 ;
      RECT 73.94 2.074 73.945 2.284 ;
      RECT 73.855 2.059 73.94 2.23 ;
      RECT 73.825 2.04 73.855 2.18 ;
      RECT 73.745 2.023 73.825 2.165 ;
      RECT 73.71 2.01 73.745 2.15 ;
      RECT 73.702 2.01 73.71 2.145 ;
      RECT 73.616 2.011 73.702 2.145 ;
      RECT 73.53 2.013 73.616 2.145 ;
      RECT 73.505 2.014 73.53 2.149 ;
      RECT 73.43 2.02 73.505 2.164 ;
      RECT 73.347 2.032 73.43 2.188 ;
      RECT 73.261 2.045 73.347 2.214 ;
      RECT 73.175 2.058 73.261 2.24 ;
      RECT 73.14 2.067 73.175 2.259 ;
      RECT 73.09 2.067 73.14 2.272 ;
      RECT 73.08 2.065 73.09 2.283 ;
      RECT 73.065 2.062 73.075 2.285 ;
      RECT 73.05 2.054 73.065 2.293 ;
      RECT 73.035 2.046 73.05 2.313 ;
      RECT 73.03 2.041 73.035 2.37 ;
      RECT 73.015 2.036 73.03 2.443 ;
      RECT 73.01 2.031 73.015 2.485 ;
      RECT 73.005 2.029 73.01 2.513 ;
      RECT 73 2.027 73.005 2.535 ;
      RECT 72.99 2.023 73 2.578 ;
      RECT 72.985 2.02 72.99 2.603 ;
      RECT 72.98 2.018 72.985 2.623 ;
      RECT 72.975 2.016 72.98 2.647 ;
      RECT 72.97 2.012 72.975 2.67 ;
      RECT 72.965 2.008 72.97 2.693 ;
      RECT 72.93 1.998 72.965 2.8 ;
      RECT 72.925 1.988 72.93 2.898 ;
      RECT 72.92 1.986 72.925 2.925 ;
      RECT 72.915 1.985 72.92 2.945 ;
      RECT 72.91 1.977 72.915 2.965 ;
      RECT 72.905 1.972 72.91 3 ;
      RECT 72.9 1.97 72.905 3.018 ;
      RECT 72.895 1.97 72.9 3.043 ;
      RECT 72.89 1.97 72.895 3.065 ;
      RECT 72.855 1.97 72.89 3.108 ;
      RECT 72.83 1.97 72.855 3.137 ;
      RECT 72.82 1.97 72.83 2.323 ;
      RECT 72.823 2.38 72.83 3.147 ;
      RECT 72.82 2.437 72.823 3.15 ;
      RECT 72.815 1.97 72.82 2.295 ;
      RECT 72.815 2.487 72.82 3.153 ;
      RECT 72.805 1.97 72.815 2.285 ;
      RECT 72.81 2.54 72.815 3.156 ;
      RECT 72.805 2.625 72.81 3.16 ;
      RECT 72.795 1.97 72.805 2.273 ;
      RECT 72.8 2.672 72.805 3.164 ;
      RECT 72.795 2.747 72.8 3.168 ;
      RECT 72.76 1.97 72.795 2.248 ;
      RECT 72.785 2.83 72.795 3.173 ;
      RECT 72.775 2.897 72.785 3.18 ;
      RECT 72.77 2.925 72.775 3.185 ;
      RECT 72.76 2.938 72.77 3.191 ;
      RECT 72.715 1.97 72.76 2.205 ;
      RECT 72.755 2.943 72.76 3.198 ;
      RECT 72.715 2.96 72.755 3.26 ;
      RECT 72.71 1.972 72.715 2.178 ;
      RECT 72.685 2.98 72.715 3.26 ;
      RECT 72.705 1.977 72.71 2.15 ;
      RECT 72.495 2.989 72.535 3.26 ;
      RECT 72.47 2.997 72.495 3.23 ;
      RECT 72.425 3.005 72.47 3.23 ;
      RECT 72.41 3.01 72.425 3.225 ;
      RECT 72.4 3.01 72.41 3.219 ;
      RECT 72.39 3.017 72.4 3.216 ;
      RECT 72.385 3.055 72.39 3.205 ;
      RECT 72.38 3.117 72.385 3.183 ;
      RECT 73.65 2.992 73.835 3.215 ;
      RECT 73.65 3.007 73.84 3.211 ;
      RECT 73.64 2.28 73.725 3.21 ;
      RECT 73.64 3.007 73.845 3.204 ;
      RECT 73.635 3.015 73.845 3.203 ;
      RECT 73.84 2.735 74.16 3.055 ;
      RECT 73.635 2.907 73.805 2.998 ;
      RECT 73.63 2.907 73.805 2.98 ;
      RECT 73.62 2.715 73.755 2.955 ;
      RECT 73.615 2.715 73.755 2.9 ;
      RECT 73.575 2.295 73.745 2.8 ;
      RECT 73.56 2.295 73.745 2.67 ;
      RECT 73.555 2.295 73.745 2.623 ;
      RECT 73.55 2.295 73.745 2.603 ;
      RECT 73.545 2.295 73.745 2.578 ;
      RECT 73.515 2.295 73.775 2.555 ;
      RECT 73.525 2.292 73.735 2.555 ;
      RECT 73.65 2.287 73.735 3.215 ;
      RECT 73.535 2.28 73.725 2.555 ;
      RECT 73.53 2.285 73.725 2.555 ;
      RECT 72.36 2.497 72.545 2.71 ;
      RECT 72.36 2.505 72.555 2.703 ;
      RECT 72.34 2.505 72.555 2.7 ;
      RECT 72.335 2.505 72.555 2.685 ;
      RECT 72.265 2.42 72.525 2.68 ;
      RECT 72.265 2.565 72.56 2.593 ;
      RECT 71.92 3.02 72.18 3.28 ;
      RECT 71.945 2.965 72.14 3.28 ;
      RECT 71.94 2.714 72.12 3.008 ;
      RECT 71.94 2.72 72.13 3.008 ;
      RECT 71.92 2.722 72.13 2.953 ;
      RECT 71.915 2.732 72.13 2.82 ;
      RECT 71.945 2.712 72.12 3.28 ;
      RECT 72.031 2.71 72.12 3.28 ;
      RECT 71.89 1.93 71.925 2.3 ;
      RECT 71.68 2.04 71.685 2.3 ;
      RECT 71.925 1.937 71.94 2.3 ;
      RECT 71.815 1.93 71.89 2.378 ;
      RECT 71.805 1.93 71.815 2.463 ;
      RECT 71.78 1.93 71.805 2.498 ;
      RECT 71.74 1.93 71.78 2.566 ;
      RECT 71.73 1.937 71.74 2.618 ;
      RECT 71.7 2.04 71.73 2.659 ;
      RECT 71.695 2.04 71.7 2.698 ;
      RECT 71.685 2.04 71.695 2.718 ;
      RECT 71.68 2.335 71.685 2.755 ;
      RECT 71.675 2.352 71.68 2.775 ;
      RECT 71.66 2.415 71.675 2.815 ;
      RECT 71.655 2.458 71.66 2.85 ;
      RECT 71.65 2.466 71.655 2.863 ;
      RECT 71.64 2.48 71.65 2.885 ;
      RECT 71.615 2.515 71.64 2.95 ;
      RECT 71.605 2.55 71.615 3.013 ;
      RECT 71.585 2.58 71.605 3.074 ;
      RECT 71.57 2.616 71.585 3.141 ;
      RECT 71.56 2.644 71.57 3.18 ;
      RECT 71.55 2.666 71.56 3.2 ;
      RECT 71.545 2.676 71.55 3.211 ;
      RECT 71.54 2.685 71.545 3.214 ;
      RECT 71.53 2.703 71.54 3.218 ;
      RECT 71.52 2.721 71.53 3.219 ;
      RECT 71.495 2.76 71.52 3.216 ;
      RECT 71.475 2.802 71.495 3.213 ;
      RECT 71.46 2.84 71.475 3.212 ;
      RECT 71.425 2.875 71.46 3.209 ;
      RECT 71.42 2.897 71.425 3.207 ;
      RECT 71.355 2.937 71.42 3.204 ;
      RECT 71.35 2.977 71.355 3.2 ;
      RECT 71.335 2.987 71.35 3.191 ;
      RECT 71.325 3.107 71.335 3.176 ;
      RECT 71.805 3.52 71.815 3.78 ;
      RECT 71.805 3.523 71.825 3.779 ;
      RECT 71.795 3.513 71.805 3.778 ;
      RECT 71.785 3.528 71.865 3.774 ;
      RECT 71.77 3.507 71.785 3.772 ;
      RECT 71.745 3.532 71.87 3.768 ;
      RECT 71.73 3.492 71.745 3.763 ;
      RECT 71.73 3.534 71.88 3.762 ;
      RECT 71.73 3.542 71.895 3.755 ;
      RECT 71.67 3.479 71.73 3.745 ;
      RECT 71.66 3.466 71.67 3.727 ;
      RECT 71.635 3.456 71.66 3.717 ;
      RECT 71.63 3.446 71.635 3.709 ;
      RECT 71.565 3.542 71.895 3.691 ;
      RECT 71.48 3.542 71.895 3.653 ;
      RECT 71.37 3.37 71.63 3.63 ;
      RECT 71.745 3.5 71.77 3.768 ;
      RECT 71.785 3.51 71.795 3.774 ;
      RECT 71.37 3.518 71.81 3.63 ;
      RECT 71.555 7.765 71.845 7.995 ;
      RECT 71.615 7.025 71.785 7.995 ;
      RECT 71.515 7.055 71.885 7.425 ;
      RECT 71.555 7.025 71.845 7.425 ;
      RECT 70.585 3.275 70.615 3.575 ;
      RECT 70.36 3.26 70.365 3.535 ;
      RECT 70.16 3.26 70.315 3.52 ;
      RECT 71.46 1.975 71.49 2.235 ;
      RECT 71.45 1.975 71.46 2.343 ;
      RECT 71.43 1.975 71.45 2.353 ;
      RECT 71.415 1.975 71.43 2.365 ;
      RECT 71.36 1.975 71.415 2.415 ;
      RECT 71.345 1.975 71.36 2.463 ;
      RECT 71.315 1.975 71.345 2.498 ;
      RECT 71.26 1.975 71.315 2.56 ;
      RECT 71.24 1.975 71.26 2.628 ;
      RECT 71.235 1.975 71.24 2.658 ;
      RECT 71.23 1.975 71.235 2.67 ;
      RECT 71.225 2.092 71.23 2.688 ;
      RECT 71.205 2.11 71.225 2.713 ;
      RECT 71.185 2.137 71.205 2.763 ;
      RECT 71.18 2.157 71.185 2.794 ;
      RECT 71.175 2.165 71.18 2.811 ;
      RECT 71.16 2.191 71.175 2.84 ;
      RECT 71.145 2.233 71.16 2.875 ;
      RECT 71.14 2.262 71.145 2.898 ;
      RECT 71.135 2.277 71.14 2.911 ;
      RECT 71.13 2.3 71.135 2.922 ;
      RECT 71.12 2.32 71.13 2.94 ;
      RECT 71.11 2.35 71.12 2.963 ;
      RECT 71.105 2.372 71.11 2.983 ;
      RECT 71.1 2.387 71.105 2.998 ;
      RECT 71.085 2.417 71.1 3.025 ;
      RECT 71.08 2.447 71.085 3.051 ;
      RECT 71.075 2.465 71.08 3.063 ;
      RECT 71.065 2.495 71.075 3.082 ;
      RECT 71.055 2.52 71.065 3.107 ;
      RECT 71.05 2.54 71.055 3.126 ;
      RECT 71.045 2.557 71.05 3.139 ;
      RECT 71.035 2.583 71.045 3.158 ;
      RECT 71.025 2.621 71.035 3.185 ;
      RECT 71.02 2.647 71.025 3.205 ;
      RECT 71.015 2.657 71.02 3.215 ;
      RECT 71.01 2.67 71.015 3.23 ;
      RECT 71.005 2.685 71.01 3.24 ;
      RECT 71 2.707 71.005 3.255 ;
      RECT 70.995 2.725 71 3.266 ;
      RECT 70.99 2.735 70.995 3.277 ;
      RECT 70.985 2.743 70.99 3.289 ;
      RECT 70.98 2.751 70.985 3.3 ;
      RECT 70.975 2.777 70.98 3.313 ;
      RECT 70.965 2.805 70.975 3.326 ;
      RECT 70.96 2.835 70.965 3.335 ;
      RECT 70.955 2.85 70.96 3.342 ;
      RECT 70.94 2.875 70.955 3.349 ;
      RECT 70.935 2.897 70.94 3.355 ;
      RECT 70.93 2.922 70.935 3.358 ;
      RECT 70.921 2.95 70.93 3.362 ;
      RECT 70.915 2.967 70.921 3.367 ;
      RECT 70.91 2.985 70.915 3.371 ;
      RECT 70.905 2.997 70.91 3.374 ;
      RECT 70.9 3.018 70.905 3.378 ;
      RECT 70.895 3.036 70.9 3.381 ;
      RECT 70.89 3.05 70.895 3.384 ;
      RECT 70.885 3.067 70.89 3.387 ;
      RECT 70.88 3.08 70.885 3.39 ;
      RECT 70.855 3.117 70.88 3.398 ;
      RECT 70.85 3.162 70.855 3.407 ;
      RECT 70.845 3.19 70.85 3.41 ;
      RECT 70.835 3.21 70.845 3.414 ;
      RECT 70.83 3.23 70.835 3.419 ;
      RECT 70.825 3.245 70.83 3.422 ;
      RECT 70.805 3.255 70.825 3.429 ;
      RECT 70.74 3.262 70.805 3.455 ;
      RECT 70.705 3.265 70.74 3.483 ;
      RECT 70.69 3.268 70.705 3.498 ;
      RECT 70.68 3.269 70.69 3.513 ;
      RECT 70.67 3.27 70.68 3.53 ;
      RECT 70.665 3.27 70.67 3.545 ;
      RECT 70.66 3.27 70.665 3.553 ;
      RECT 70.645 3.271 70.66 3.568 ;
      RECT 70.615 3.273 70.645 3.575 ;
      RECT 70.505 3.28 70.585 3.575 ;
      RECT 70.46 3.285 70.505 3.575 ;
      RECT 70.45 3.286 70.46 3.565 ;
      RECT 70.44 3.287 70.45 3.558 ;
      RECT 70.42 3.289 70.44 3.553 ;
      RECT 70.41 3.26 70.42 3.548 ;
      RECT 70.365 3.26 70.41 3.54 ;
      RECT 70.335 3.26 70.36 3.53 ;
      RECT 70.315 3.26 70.335 3.523 ;
      RECT 70.595 2.06 70.855 2.32 ;
      RECT 70.475 2.075 70.485 2.24 ;
      RECT 70.46 2.075 70.465 2.235 ;
      RECT 67.825 1.915 68.01 2.205 ;
      RECT 69.64 2.04 69.655 2.195 ;
      RECT 67.79 1.915 67.815 2.175 ;
      RECT 70.205 1.965 70.21 2.107 ;
      RECT 70.12 1.96 70.145 2.1 ;
      RECT 70.52 2.077 70.595 2.27 ;
      RECT 70.505 2.075 70.52 2.253 ;
      RECT 70.485 2.075 70.505 2.245 ;
      RECT 70.465 2.075 70.475 2.238 ;
      RECT 70.42 2.07 70.46 2.228 ;
      RECT 70.38 2.045 70.42 2.213 ;
      RECT 70.365 2.02 70.38 2.203 ;
      RECT 70.36 2.014 70.365 2.201 ;
      RECT 70.325 2.006 70.36 2.184 ;
      RECT 70.32 1.999 70.325 2.172 ;
      RECT 70.3 1.994 70.32 2.16 ;
      RECT 70.29 1.988 70.3 2.145 ;
      RECT 70.27 1.983 70.29 2.13 ;
      RECT 70.26 1.978 70.27 2.123 ;
      RECT 70.255 1.976 70.26 2.118 ;
      RECT 70.25 1.975 70.255 2.115 ;
      RECT 70.21 1.97 70.25 2.111 ;
      RECT 70.19 1.964 70.205 2.106 ;
      RECT 70.155 1.961 70.19 2.103 ;
      RECT 70.145 1.96 70.155 2.101 ;
      RECT 70.085 1.96 70.12 2.098 ;
      RECT 70.04 1.96 70.085 2.098 ;
      RECT 69.99 1.96 70.04 2.101 ;
      RECT 69.975 1.962 69.99 2.103 ;
      RECT 69.96 1.965 69.975 2.104 ;
      RECT 69.95 1.97 69.96 2.105 ;
      RECT 69.92 1.975 69.95 2.11 ;
      RECT 69.91 1.981 69.92 2.118 ;
      RECT 69.9 1.983 69.91 2.122 ;
      RECT 69.89 1.987 69.9 2.126 ;
      RECT 69.865 1.993 69.89 2.134 ;
      RECT 69.855 1.998 69.865 2.142 ;
      RECT 69.84 2.002 69.855 2.146 ;
      RECT 69.805 2.008 69.84 2.154 ;
      RECT 69.785 2.013 69.805 2.164 ;
      RECT 69.755 2.02 69.785 2.173 ;
      RECT 69.71 2.029 69.755 2.187 ;
      RECT 69.705 2.034 69.71 2.198 ;
      RECT 69.685 2.037 69.705 2.199 ;
      RECT 69.655 2.04 69.685 2.197 ;
      RECT 69.62 2.04 69.64 2.193 ;
      RECT 69.55 2.04 69.62 2.184 ;
      RECT 69.535 2.037 69.55 2.176 ;
      RECT 69.495 2.03 69.535 2.171 ;
      RECT 69.47 2.02 69.495 2.164 ;
      RECT 69.465 2.014 69.47 2.161 ;
      RECT 69.425 2.008 69.465 2.158 ;
      RECT 69.41 2.001 69.425 2.153 ;
      RECT 69.39 1.997 69.41 2.148 ;
      RECT 69.375 1.992 69.39 2.144 ;
      RECT 69.36 1.987 69.375 2.142 ;
      RECT 69.345 1.983 69.36 2.141 ;
      RECT 69.33 1.981 69.345 2.137 ;
      RECT 69.32 1.979 69.33 2.132 ;
      RECT 69.305 1.976 69.32 2.128 ;
      RECT 69.295 1.974 69.305 2.123 ;
      RECT 69.275 1.971 69.295 2.119 ;
      RECT 69.23 1.97 69.275 2.117 ;
      RECT 69.17 1.972 69.23 2.118 ;
      RECT 69.15 1.974 69.17 2.12 ;
      RECT 69.12 1.977 69.15 2.121 ;
      RECT 69.07 1.982 69.12 2.123 ;
      RECT 69.065 1.985 69.07 2.125 ;
      RECT 69.055 1.987 69.065 2.128 ;
      RECT 69.05 1.989 69.055 2.131 ;
      RECT 69 1.992 69.05 2.138 ;
      RECT 68.98 1.996 69 2.15 ;
      RECT 68.97 1.999 68.98 2.156 ;
      RECT 68.96 2 68.97 2.159 ;
      RECT 68.921 2.003 68.96 2.161 ;
      RECT 68.835 2.01 68.921 2.164 ;
      RECT 68.761 2.02 68.835 2.168 ;
      RECT 68.675 2.031 68.761 2.173 ;
      RECT 68.66 2.038 68.675 2.175 ;
      RECT 68.605 2.042 68.66 2.176 ;
      RECT 68.591 2.045 68.605 2.178 ;
      RECT 68.505 2.045 68.591 2.18 ;
      RECT 68.465 2.042 68.505 2.183 ;
      RECT 68.441 2.038 68.465 2.185 ;
      RECT 68.355 2.028 68.441 2.188 ;
      RECT 68.325 2.017 68.355 2.189 ;
      RECT 68.306 2.013 68.325 2.188 ;
      RECT 68.22 2.006 68.306 2.185 ;
      RECT 68.16 1.995 68.22 2.182 ;
      RECT 68.14 1.987 68.16 2.18 ;
      RECT 68.105 1.982 68.14 2.179 ;
      RECT 68.08 1.977 68.105 2.178 ;
      RECT 68.05 1.972 68.08 2.177 ;
      RECT 68.025 1.915 68.05 2.176 ;
      RECT 68.01 1.915 68.025 2.2 ;
      RECT 67.815 1.915 67.825 2.2 ;
      RECT 69.59 2.935 69.595 3.075 ;
      RECT 69.25 2.935 69.285 3.073 ;
      RECT 68.825 2.92 68.84 3.065 ;
      RECT 70.655 2.7 70.745 2.96 ;
      RECT 70.485 2.565 70.585 2.96 ;
      RECT 67.52 2.54 67.6 2.75 ;
      RECT 70.61 2.677 70.655 2.96 ;
      RECT 70.6 2.647 70.61 2.96 ;
      RECT 70.585 2.57 70.6 2.96 ;
      RECT 70.4 2.565 70.485 2.925 ;
      RECT 70.395 2.567 70.4 2.92 ;
      RECT 70.39 2.572 70.395 2.92 ;
      RECT 70.355 2.672 70.39 2.92 ;
      RECT 70.345 2.7 70.355 2.92 ;
      RECT 70.335 2.715 70.345 2.92 ;
      RECT 70.325 2.727 70.335 2.92 ;
      RECT 70.32 2.737 70.325 2.92 ;
      RECT 70.305 2.747 70.32 2.922 ;
      RECT 70.3 2.762 70.305 2.924 ;
      RECT 70.285 2.775 70.3 2.926 ;
      RECT 70.28 2.79 70.285 2.929 ;
      RECT 70.26 2.8 70.28 2.933 ;
      RECT 70.245 2.81 70.26 2.936 ;
      RECT 70.21 2.817 70.245 2.941 ;
      RECT 70.166 2.824 70.21 2.949 ;
      RECT 70.08 2.836 70.166 2.962 ;
      RECT 70.055 2.847 70.08 2.973 ;
      RECT 70.025 2.852 70.055 2.978 ;
      RECT 69.99 2.857 70.025 2.986 ;
      RECT 69.96 2.862 69.99 2.993 ;
      RECT 69.935 2.867 69.96 2.998 ;
      RECT 69.87 2.874 69.935 3.007 ;
      RECT 69.8 2.887 69.87 3.023 ;
      RECT 69.77 2.897 69.8 3.035 ;
      RECT 69.745 2.902 69.77 3.042 ;
      RECT 69.69 2.909 69.745 3.05 ;
      RECT 69.685 2.916 69.69 3.055 ;
      RECT 69.68 2.918 69.685 3.056 ;
      RECT 69.665 2.92 69.68 3.058 ;
      RECT 69.66 2.92 69.665 3.061 ;
      RECT 69.595 2.927 69.66 3.068 ;
      RECT 69.56 2.937 69.59 3.078 ;
      RECT 69.543 2.94 69.56 3.08 ;
      RECT 69.457 2.939 69.543 3.079 ;
      RECT 69.371 2.937 69.457 3.076 ;
      RECT 69.285 2.936 69.371 3.074 ;
      RECT 69.184 2.934 69.25 3.073 ;
      RECT 69.098 2.931 69.184 3.071 ;
      RECT 69.012 2.927 69.098 3.069 ;
      RECT 68.926 2.924 69.012 3.068 ;
      RECT 68.84 2.921 68.926 3.066 ;
      RECT 68.74 2.92 68.825 3.063 ;
      RECT 68.69 2.918 68.74 3.061 ;
      RECT 68.67 2.915 68.69 3.059 ;
      RECT 68.65 2.913 68.67 3.056 ;
      RECT 68.625 2.909 68.65 3.053 ;
      RECT 68.58 2.903 68.625 3.048 ;
      RECT 68.54 2.897 68.58 3.04 ;
      RECT 68.515 2.892 68.54 3.033 ;
      RECT 68.46 2.885 68.515 3.025 ;
      RECT 68.436 2.878 68.46 3.018 ;
      RECT 68.35 2.869 68.436 3.008 ;
      RECT 68.32 2.861 68.35 2.998 ;
      RECT 68.29 2.857 68.32 2.993 ;
      RECT 68.285 2.854 68.29 2.99 ;
      RECT 68.28 2.853 68.285 2.99 ;
      RECT 68.205 2.846 68.28 2.983 ;
      RECT 68.166 2.837 68.205 2.972 ;
      RECT 68.08 2.827 68.166 2.96 ;
      RECT 68.04 2.817 68.08 2.948 ;
      RECT 68.001 2.812 68.04 2.941 ;
      RECT 67.915 2.802 68.001 2.93 ;
      RECT 67.875 2.79 67.915 2.919 ;
      RECT 67.84 2.775 67.875 2.912 ;
      RECT 67.83 2.765 67.84 2.909 ;
      RECT 67.81 2.75 67.83 2.907 ;
      RECT 67.78 2.72 67.81 2.903 ;
      RECT 67.77 2.7 67.78 2.898 ;
      RECT 67.765 2.692 67.77 2.895 ;
      RECT 67.76 2.685 67.765 2.893 ;
      RECT 67.745 2.672 67.76 2.886 ;
      RECT 67.74 2.662 67.745 2.878 ;
      RECT 67.735 2.655 67.74 2.873 ;
      RECT 67.73 2.65 67.735 2.869 ;
      RECT 67.715 2.637 67.73 2.861 ;
      RECT 67.71 2.547 67.715 2.85 ;
      RECT 67.705 2.542 67.71 2.843 ;
      RECT 67.63 2.54 67.705 2.803 ;
      RECT 67.6 2.54 67.63 2.758 ;
      RECT 67.505 2.545 67.52 2.745 ;
      RECT 69.99 2.25 70.25 2.51 ;
      RECT 69.975 2.238 70.155 2.475 ;
      RECT 69.97 2.239 70.155 2.473 ;
      RECT 69.955 2.243 70.165 2.463 ;
      RECT 69.95 2.248 70.17 2.433 ;
      RECT 69.955 2.245 70.17 2.463 ;
      RECT 69.97 2.24 70.165 2.473 ;
      RECT 69.99 2.237 70.155 2.51 ;
      RECT 69.99 2.236 70.145 2.51 ;
      RECT 70.015 2.235 70.145 2.51 ;
      RECT 69.575 2.48 69.835 2.74 ;
      RECT 69.45 2.525 69.835 2.735 ;
      RECT 69.44 2.53 69.835 2.73 ;
      RECT 69.455 3.47 69.47 3.78 ;
      RECT 68.05 3.24 68.06 3.37 ;
      RECT 67.83 3.235 67.935 3.37 ;
      RECT 67.745 3.24 67.795 3.37 ;
      RECT 66.295 1.975 66.3 3.08 ;
      RECT 69.55 3.562 69.555 3.698 ;
      RECT 69.545 3.557 69.55 3.758 ;
      RECT 69.54 3.555 69.545 3.771 ;
      RECT 69.525 3.552 69.54 3.773 ;
      RECT 69.52 3.547 69.525 3.775 ;
      RECT 69.515 3.543 69.52 3.778 ;
      RECT 69.5 3.538 69.515 3.78 ;
      RECT 69.47 3.53 69.5 3.78 ;
      RECT 69.431 3.47 69.455 3.78 ;
      RECT 69.345 3.47 69.431 3.777 ;
      RECT 69.315 3.47 69.345 3.77 ;
      RECT 69.29 3.47 69.315 3.763 ;
      RECT 69.265 3.47 69.29 3.755 ;
      RECT 69.25 3.47 69.265 3.748 ;
      RECT 69.225 3.47 69.25 3.74 ;
      RECT 69.21 3.47 69.225 3.733 ;
      RECT 69.17 3.48 69.21 3.722 ;
      RECT 69.16 3.475 69.17 3.712 ;
      RECT 69.156 3.474 69.16 3.709 ;
      RECT 69.07 3.466 69.156 3.692 ;
      RECT 69.037 3.455 69.07 3.669 ;
      RECT 68.951 3.444 69.037 3.647 ;
      RECT 68.865 3.428 68.951 3.616 ;
      RECT 68.795 3.413 68.865 3.588 ;
      RECT 68.785 3.406 68.795 3.575 ;
      RECT 68.755 3.403 68.785 3.565 ;
      RECT 68.73 3.399 68.755 3.558 ;
      RECT 68.715 3.396 68.73 3.553 ;
      RECT 68.71 3.395 68.715 3.548 ;
      RECT 68.68 3.39 68.71 3.541 ;
      RECT 68.675 3.385 68.68 3.536 ;
      RECT 68.66 3.382 68.675 3.531 ;
      RECT 68.655 3.377 68.66 3.526 ;
      RECT 68.635 3.372 68.655 3.523 ;
      RECT 68.62 3.367 68.635 3.515 ;
      RECT 68.605 3.361 68.62 3.51 ;
      RECT 68.575 3.352 68.605 3.503 ;
      RECT 68.57 3.345 68.575 3.495 ;
      RECT 68.565 3.343 68.57 3.493 ;
      RECT 68.56 3.342 68.565 3.49 ;
      RECT 68.52 3.335 68.56 3.483 ;
      RECT 68.506 3.325 68.52 3.473 ;
      RECT 68.455 3.314 68.506 3.461 ;
      RECT 68.43 3.3 68.455 3.447 ;
      RECT 68.405 3.289 68.43 3.439 ;
      RECT 68.385 3.278 68.405 3.433 ;
      RECT 68.375 3.272 68.385 3.428 ;
      RECT 68.37 3.27 68.375 3.424 ;
      RECT 68.35 3.265 68.37 3.419 ;
      RECT 68.32 3.255 68.35 3.409 ;
      RECT 68.315 3.247 68.32 3.402 ;
      RECT 68.3 3.245 68.315 3.398 ;
      RECT 68.28 3.245 68.3 3.393 ;
      RECT 68.275 3.244 68.28 3.391 ;
      RECT 68.27 3.244 68.275 3.388 ;
      RECT 68.23 3.243 68.27 3.383 ;
      RECT 68.205 3.242 68.23 3.378 ;
      RECT 68.145 3.241 68.205 3.375 ;
      RECT 68.06 3.24 68.145 3.373 ;
      RECT 68.021 3.239 68.05 3.37 ;
      RECT 67.935 3.237 68.021 3.37 ;
      RECT 67.795 3.237 67.83 3.37 ;
      RECT 67.705 3.241 67.745 3.373 ;
      RECT 67.69 3.244 67.705 3.38 ;
      RECT 67.68 3.245 67.69 3.387 ;
      RECT 67.655 3.248 67.68 3.392 ;
      RECT 67.65 3.25 67.655 3.395 ;
      RECT 67.6 3.252 67.65 3.396 ;
      RECT 67.561 3.256 67.6 3.398 ;
      RECT 67.475 3.258 67.561 3.401 ;
      RECT 67.457 3.26 67.475 3.403 ;
      RECT 67.371 3.263 67.457 3.405 ;
      RECT 67.285 3.267 67.371 3.408 ;
      RECT 67.248 3.271 67.285 3.411 ;
      RECT 67.162 3.274 67.248 3.414 ;
      RECT 67.076 3.278 67.162 3.417 ;
      RECT 66.99 3.283 67.076 3.421 ;
      RECT 66.97 3.285 66.99 3.424 ;
      RECT 66.95 3.284 66.97 3.425 ;
      RECT 66.901 3.281 66.95 3.426 ;
      RECT 66.815 3.276 66.901 3.429 ;
      RECT 66.765 3.271 66.815 3.431 ;
      RECT 66.741 3.269 66.765 3.432 ;
      RECT 66.655 3.264 66.741 3.434 ;
      RECT 66.63 3.26 66.655 3.433 ;
      RECT 66.62 3.257 66.63 3.431 ;
      RECT 66.61 3.25 66.62 3.428 ;
      RECT 66.605 3.23 66.61 3.423 ;
      RECT 66.595 3.2 66.605 3.418 ;
      RECT 66.58 3.07 66.595 3.409 ;
      RECT 66.575 3.062 66.58 3.402 ;
      RECT 66.555 3.055 66.575 3.394 ;
      RECT 66.55 3.037 66.555 3.386 ;
      RECT 66.54 3.017 66.55 3.381 ;
      RECT 66.535 2.99 66.54 3.377 ;
      RECT 66.53 2.967 66.535 3.374 ;
      RECT 66.51 2.925 66.53 3.366 ;
      RECT 66.475 2.84 66.51 3.35 ;
      RECT 66.47 2.772 66.475 3.338 ;
      RECT 66.455 2.742 66.47 3.332 ;
      RECT 66.45 1.987 66.455 2.233 ;
      RECT 66.44 2.712 66.455 3.323 ;
      RECT 66.445 1.982 66.45 2.265 ;
      RECT 66.44 1.977 66.445 2.308 ;
      RECT 66.435 1.975 66.44 2.343 ;
      RECT 66.42 2.675 66.44 3.313 ;
      RECT 66.43 1.975 66.435 2.38 ;
      RECT 66.415 1.975 66.43 2.478 ;
      RECT 66.415 2.648 66.42 3.306 ;
      RECT 66.41 1.975 66.415 2.553 ;
      RECT 66.41 2.636 66.415 3.303 ;
      RECT 66.405 1.975 66.41 2.585 ;
      RECT 66.405 2.615 66.41 3.3 ;
      RECT 66.4 1.975 66.405 3.297 ;
      RECT 66.365 1.975 66.4 3.283 ;
      RECT 66.35 1.975 66.365 3.265 ;
      RECT 66.33 1.975 66.35 3.255 ;
      RECT 66.305 1.975 66.33 3.238 ;
      RECT 66.3 1.975 66.305 3.188 ;
      RECT 66.29 1.975 66.295 3.018 ;
      RECT 66.285 1.975 66.29 2.925 ;
      RECT 66.28 1.975 66.285 2.838 ;
      RECT 66.275 1.975 66.28 2.77 ;
      RECT 66.27 1.975 66.275 2.713 ;
      RECT 66.26 1.975 66.27 2.608 ;
      RECT 66.255 1.975 66.26 2.48 ;
      RECT 66.25 1.975 66.255 2.398 ;
      RECT 66.245 1.977 66.25 2.315 ;
      RECT 66.24 1.982 66.245 2.248 ;
      RECT 66.235 1.987 66.24 2.175 ;
      RECT 69.05 2.305 69.31 2.565 ;
      RECT 69.07 2.272 69.28 2.565 ;
      RECT 69.07 2.27 69.27 2.565 ;
      RECT 69.08 2.257 69.27 2.565 ;
      RECT 69.08 2.255 69.195 2.565 ;
      RECT 68.555 2.38 68.73 2.66 ;
      RECT 68.55 2.38 68.73 2.658 ;
      RECT 68.55 2.38 68.745 2.655 ;
      RECT 68.54 2.38 68.745 2.653 ;
      RECT 68.485 2.38 68.745 2.64 ;
      RECT 68.485 2.455 68.75 2.618 ;
      RECT 68.03 2.392 68.05 2.635 ;
      RECT 68.03 2.392 68.09 2.634 ;
      RECT 68.025 2.394 68.09 2.633 ;
      RECT 68.025 2.394 68.176 2.632 ;
      RECT 68.025 2.394 68.245 2.631 ;
      RECT 68.025 2.394 68.265 2.623 ;
      RECT 68.005 2.397 68.265 2.621 ;
      RECT 67.99 2.407 68.265 2.606 ;
      RECT 67.99 2.407 68.28 2.605 ;
      RECT 67.985 2.416 68.28 2.597 ;
      RECT 67.985 2.416 68.285 2.593 ;
      RECT 68.09 2.33 68.35 2.59 ;
      RECT 67.98 2.418 68.35 2.475 ;
      RECT 68.05 2.385 68.35 2.59 ;
      RECT 68.015 3.578 68.02 3.785 ;
      RECT 67.965 3.572 68.015 3.784 ;
      RECT 67.932 3.586 68.025 3.783 ;
      RECT 67.846 3.586 68.025 3.782 ;
      RECT 67.76 3.586 68.025 3.781 ;
      RECT 67.76 3.685 68.03 3.778 ;
      RECT 67.755 3.685 68.03 3.773 ;
      RECT 67.75 3.685 68.03 3.755 ;
      RECT 67.745 3.685 68.03 3.738 ;
      RECT 67.705 3.47 67.965 3.73 ;
      RECT 67.165 2.62 67.251 3.034 ;
      RECT 67.165 2.62 67.29 3.031 ;
      RECT 67.165 2.62 67.31 3.021 ;
      RECT 67.12 2.62 67.31 3.018 ;
      RECT 67.12 2.772 67.32 3.008 ;
      RECT 67.12 2.793 67.325 3.002 ;
      RECT 67.12 2.811 67.33 2.998 ;
      RECT 67.12 2.831 67.34 2.993 ;
      RECT 67.095 2.831 67.34 2.99 ;
      RECT 67.085 2.831 67.34 2.968 ;
      RECT 67.085 2.847 67.345 2.938 ;
      RECT 67.05 2.62 67.31 2.925 ;
      RECT 67.05 2.859 67.35 2.88 ;
      RECT 64.71 7.77 65 8 ;
      RECT 64.77 6.29 64.94 8 ;
      RECT 64.72 6.655 65.07 7.005 ;
      RECT 64.71 6.29 65 6.52 ;
      RECT 64.305 2.395 64.41 2.965 ;
      RECT 64.305 2.73 64.63 2.96 ;
      RECT 64.305 2.76 64.8 2.93 ;
      RECT 64.305 2.395 64.495 2.96 ;
      RECT 63.72 2.36 64.01 2.59 ;
      RECT 63.72 2.395 64.495 2.565 ;
      RECT 63.78 0.88 63.95 2.59 ;
      RECT 63.72 0.88 64.01 1.11 ;
      RECT 63.72 7.77 64.01 8 ;
      RECT 63.78 6.29 63.95 8 ;
      RECT 63.72 6.29 64.01 6.52 ;
      RECT 63.72 6.325 64.575 6.485 ;
      RECT 64.405 5.92 64.575 6.485 ;
      RECT 63.72 6.32 64.115 6.485 ;
      RECT 64.34 5.92 64.63 6.15 ;
      RECT 64.34 5.95 64.8 6.12 ;
      RECT 63.35 2.73 63.64 2.96 ;
      RECT 63.35 2.76 63.81 2.93 ;
      RECT 63.415 1.655 63.58 2.96 ;
      RECT 61.93 1.625 62.22 1.855 ;
      RECT 61.93 1.655 63.58 1.825 ;
      RECT 61.99 0.885 62.16 1.855 ;
      RECT 61.93 0.885 62.22 1.115 ;
      RECT 61.93 7.765 62.22 7.995 ;
      RECT 61.99 7.025 62.16 7.995 ;
      RECT 61.99 7.12 63.58 7.29 ;
      RECT 63.41 5.92 63.58 7.29 ;
      RECT 61.93 7.025 62.22 7.255 ;
      RECT 63.35 5.92 63.64 6.15 ;
      RECT 63.35 5.95 63.81 6.12 ;
      RECT 59.98 2.705 60.32 3.055 ;
      RECT 60.07 2.025 60.24 3.055 ;
      RECT 62.36 1.965 62.71 2.315 ;
      RECT 60.07 2.025 62.71 2.195 ;
      RECT 62.385 6.655 62.71 6.98 ;
      RECT 56.925 6.61 57.275 6.96 ;
      RECT 62.36 6.655 62.71 6.885 ;
      RECT 56.725 6.655 57.275 6.885 ;
      RECT 56.555 6.685 62.71 6.855 ;
      RECT 61.585 2.365 61.905 2.685 ;
      RECT 61.555 2.365 61.905 2.595 ;
      RECT 61.385 2.395 61.905 2.565 ;
      RECT 61.585 6.255 61.905 6.545 ;
      RECT 61.555 6.285 61.905 6.515 ;
      RECT 61.385 6.315 61.905 6.485 ;
      RECT 57.275 2.985 57.425 3.26 ;
      RECT 57.815 2.065 57.82 2.285 ;
      RECT 58.965 2.265 58.98 2.463 ;
      RECT 58.93 2.257 58.965 2.47 ;
      RECT 58.9 2.25 58.93 2.47 ;
      RECT 58.845 2.215 58.9 2.47 ;
      RECT 58.78 2.152 58.845 2.47 ;
      RECT 58.775 2.117 58.78 2.468 ;
      RECT 58.77 2.112 58.775 2.46 ;
      RECT 58.765 2.107 58.77 2.446 ;
      RECT 58.76 2.104 58.765 2.439 ;
      RECT 58.715 2.094 58.76 2.39 ;
      RECT 58.695 2.081 58.715 2.325 ;
      RECT 58.69 2.076 58.695 2.298 ;
      RECT 58.685 2.075 58.69 2.291 ;
      RECT 58.68 2.074 58.685 2.284 ;
      RECT 58.595 2.059 58.68 2.23 ;
      RECT 58.565 2.04 58.595 2.18 ;
      RECT 58.485 2.023 58.565 2.165 ;
      RECT 58.45 2.01 58.485 2.15 ;
      RECT 58.442 2.01 58.45 2.145 ;
      RECT 58.356 2.011 58.442 2.145 ;
      RECT 58.27 2.013 58.356 2.145 ;
      RECT 58.245 2.014 58.27 2.149 ;
      RECT 58.17 2.02 58.245 2.164 ;
      RECT 58.087 2.032 58.17 2.188 ;
      RECT 58.001 2.045 58.087 2.214 ;
      RECT 57.915 2.058 58.001 2.24 ;
      RECT 57.88 2.067 57.915 2.259 ;
      RECT 57.83 2.067 57.88 2.272 ;
      RECT 57.82 2.065 57.83 2.283 ;
      RECT 57.805 2.062 57.815 2.285 ;
      RECT 57.79 2.054 57.805 2.293 ;
      RECT 57.775 2.046 57.79 2.313 ;
      RECT 57.77 2.041 57.775 2.37 ;
      RECT 57.755 2.036 57.77 2.443 ;
      RECT 57.75 2.031 57.755 2.485 ;
      RECT 57.745 2.029 57.75 2.513 ;
      RECT 57.74 2.027 57.745 2.535 ;
      RECT 57.73 2.023 57.74 2.578 ;
      RECT 57.725 2.02 57.73 2.603 ;
      RECT 57.72 2.018 57.725 2.623 ;
      RECT 57.715 2.016 57.72 2.647 ;
      RECT 57.71 2.012 57.715 2.67 ;
      RECT 57.705 2.008 57.71 2.693 ;
      RECT 57.67 1.998 57.705 2.8 ;
      RECT 57.665 1.988 57.67 2.898 ;
      RECT 57.66 1.986 57.665 2.925 ;
      RECT 57.655 1.985 57.66 2.945 ;
      RECT 57.65 1.977 57.655 2.965 ;
      RECT 57.645 1.972 57.65 3 ;
      RECT 57.64 1.97 57.645 3.018 ;
      RECT 57.635 1.97 57.64 3.043 ;
      RECT 57.63 1.97 57.635 3.065 ;
      RECT 57.595 1.97 57.63 3.108 ;
      RECT 57.57 1.97 57.595 3.137 ;
      RECT 57.56 1.97 57.57 2.323 ;
      RECT 57.563 2.38 57.57 3.147 ;
      RECT 57.56 2.437 57.563 3.15 ;
      RECT 57.555 1.97 57.56 2.295 ;
      RECT 57.555 2.487 57.56 3.153 ;
      RECT 57.545 1.97 57.555 2.285 ;
      RECT 57.55 2.54 57.555 3.156 ;
      RECT 57.545 2.625 57.55 3.16 ;
      RECT 57.535 1.97 57.545 2.273 ;
      RECT 57.54 2.672 57.545 3.164 ;
      RECT 57.535 2.747 57.54 3.168 ;
      RECT 57.5 1.97 57.535 2.248 ;
      RECT 57.525 2.83 57.535 3.173 ;
      RECT 57.515 2.897 57.525 3.18 ;
      RECT 57.51 2.925 57.515 3.185 ;
      RECT 57.5 2.938 57.51 3.191 ;
      RECT 57.455 1.97 57.5 2.205 ;
      RECT 57.495 2.943 57.5 3.198 ;
      RECT 57.455 2.96 57.495 3.26 ;
      RECT 57.45 1.972 57.455 2.178 ;
      RECT 57.425 2.98 57.455 3.26 ;
      RECT 57.445 1.977 57.45 2.15 ;
      RECT 57.235 2.989 57.275 3.26 ;
      RECT 57.21 2.997 57.235 3.23 ;
      RECT 57.165 3.005 57.21 3.23 ;
      RECT 57.15 3.01 57.165 3.225 ;
      RECT 57.14 3.01 57.15 3.219 ;
      RECT 57.13 3.017 57.14 3.216 ;
      RECT 57.125 3.055 57.13 3.205 ;
      RECT 57.12 3.117 57.125 3.183 ;
      RECT 58.39 2.992 58.575 3.215 ;
      RECT 58.39 3.007 58.58 3.211 ;
      RECT 58.38 2.28 58.465 3.21 ;
      RECT 58.38 3.007 58.585 3.204 ;
      RECT 58.375 3.015 58.585 3.203 ;
      RECT 58.58 2.735 58.9 3.055 ;
      RECT 58.375 2.907 58.545 2.998 ;
      RECT 58.37 2.907 58.545 2.98 ;
      RECT 58.36 2.715 58.495 2.955 ;
      RECT 58.355 2.715 58.495 2.9 ;
      RECT 58.315 2.295 58.485 2.8 ;
      RECT 58.3 2.295 58.485 2.67 ;
      RECT 58.295 2.295 58.485 2.623 ;
      RECT 58.29 2.295 58.485 2.603 ;
      RECT 58.285 2.295 58.485 2.578 ;
      RECT 58.255 2.295 58.515 2.555 ;
      RECT 58.265 2.292 58.475 2.555 ;
      RECT 58.39 2.287 58.475 3.215 ;
      RECT 58.275 2.28 58.465 2.555 ;
      RECT 58.27 2.285 58.465 2.555 ;
      RECT 57.1 2.497 57.285 2.71 ;
      RECT 57.1 2.505 57.295 2.703 ;
      RECT 57.08 2.505 57.295 2.7 ;
      RECT 57.075 2.505 57.295 2.685 ;
      RECT 57.005 2.42 57.265 2.68 ;
      RECT 57.005 2.565 57.3 2.593 ;
      RECT 56.66 3.02 56.92 3.28 ;
      RECT 56.685 2.965 56.88 3.28 ;
      RECT 56.68 2.714 56.86 3.008 ;
      RECT 56.68 2.72 56.87 3.008 ;
      RECT 56.66 2.722 56.87 2.953 ;
      RECT 56.655 2.732 56.87 2.82 ;
      RECT 56.685 2.712 56.86 3.28 ;
      RECT 56.771 2.71 56.86 3.28 ;
      RECT 56.63 1.93 56.665 2.3 ;
      RECT 56.42 2.04 56.425 2.3 ;
      RECT 56.665 1.937 56.68 2.3 ;
      RECT 56.555 1.93 56.63 2.378 ;
      RECT 56.545 1.93 56.555 2.463 ;
      RECT 56.52 1.93 56.545 2.498 ;
      RECT 56.48 1.93 56.52 2.566 ;
      RECT 56.47 1.937 56.48 2.618 ;
      RECT 56.44 2.04 56.47 2.659 ;
      RECT 56.435 2.04 56.44 2.698 ;
      RECT 56.425 2.04 56.435 2.718 ;
      RECT 56.42 2.335 56.425 2.755 ;
      RECT 56.415 2.352 56.42 2.775 ;
      RECT 56.4 2.415 56.415 2.815 ;
      RECT 56.395 2.458 56.4 2.85 ;
      RECT 56.39 2.466 56.395 2.863 ;
      RECT 56.38 2.48 56.39 2.885 ;
      RECT 56.355 2.515 56.38 2.95 ;
      RECT 56.345 2.55 56.355 3.013 ;
      RECT 56.325 2.58 56.345 3.074 ;
      RECT 56.31 2.616 56.325 3.141 ;
      RECT 56.3 2.644 56.31 3.18 ;
      RECT 56.29 2.666 56.3 3.2 ;
      RECT 56.285 2.676 56.29 3.211 ;
      RECT 56.28 2.685 56.285 3.214 ;
      RECT 56.27 2.703 56.28 3.218 ;
      RECT 56.26 2.721 56.27 3.219 ;
      RECT 56.235 2.76 56.26 3.216 ;
      RECT 56.215 2.802 56.235 3.213 ;
      RECT 56.2 2.84 56.215 3.212 ;
      RECT 56.165 2.875 56.2 3.209 ;
      RECT 56.16 2.897 56.165 3.207 ;
      RECT 56.095 2.937 56.16 3.204 ;
      RECT 56.09 2.977 56.095 3.2 ;
      RECT 56.075 2.987 56.09 3.191 ;
      RECT 56.065 3.107 56.075 3.176 ;
      RECT 56.545 3.52 56.555 3.78 ;
      RECT 56.545 3.523 56.565 3.779 ;
      RECT 56.535 3.513 56.545 3.778 ;
      RECT 56.525 3.528 56.605 3.774 ;
      RECT 56.51 3.507 56.525 3.772 ;
      RECT 56.485 3.532 56.61 3.768 ;
      RECT 56.47 3.492 56.485 3.763 ;
      RECT 56.47 3.534 56.62 3.762 ;
      RECT 56.47 3.542 56.635 3.755 ;
      RECT 56.41 3.479 56.47 3.745 ;
      RECT 56.4 3.466 56.41 3.727 ;
      RECT 56.375 3.456 56.4 3.717 ;
      RECT 56.37 3.446 56.375 3.709 ;
      RECT 56.305 3.542 56.635 3.691 ;
      RECT 56.22 3.542 56.635 3.653 ;
      RECT 56.11 3.37 56.37 3.63 ;
      RECT 56.485 3.5 56.51 3.768 ;
      RECT 56.525 3.51 56.535 3.774 ;
      RECT 56.11 3.518 56.55 3.63 ;
      RECT 56.295 7.765 56.585 7.995 ;
      RECT 56.355 7.025 56.525 7.995 ;
      RECT 56.255 7.055 56.625 7.425 ;
      RECT 56.295 7.025 56.585 7.425 ;
      RECT 55.325 3.275 55.355 3.575 ;
      RECT 55.1 3.26 55.105 3.535 ;
      RECT 54.9 3.26 55.055 3.52 ;
      RECT 56.2 1.975 56.23 2.235 ;
      RECT 56.19 1.975 56.2 2.343 ;
      RECT 56.17 1.975 56.19 2.353 ;
      RECT 56.155 1.975 56.17 2.365 ;
      RECT 56.1 1.975 56.155 2.415 ;
      RECT 56.085 1.975 56.1 2.463 ;
      RECT 56.055 1.975 56.085 2.498 ;
      RECT 56 1.975 56.055 2.56 ;
      RECT 55.98 1.975 56 2.628 ;
      RECT 55.975 1.975 55.98 2.658 ;
      RECT 55.97 1.975 55.975 2.67 ;
      RECT 55.965 2.092 55.97 2.688 ;
      RECT 55.945 2.11 55.965 2.713 ;
      RECT 55.925 2.137 55.945 2.763 ;
      RECT 55.92 2.157 55.925 2.794 ;
      RECT 55.915 2.165 55.92 2.811 ;
      RECT 55.9 2.191 55.915 2.84 ;
      RECT 55.885 2.233 55.9 2.875 ;
      RECT 55.88 2.262 55.885 2.898 ;
      RECT 55.875 2.277 55.88 2.911 ;
      RECT 55.87 2.3 55.875 2.922 ;
      RECT 55.86 2.32 55.87 2.94 ;
      RECT 55.85 2.35 55.86 2.963 ;
      RECT 55.845 2.372 55.85 2.983 ;
      RECT 55.84 2.387 55.845 2.998 ;
      RECT 55.825 2.417 55.84 3.025 ;
      RECT 55.82 2.447 55.825 3.051 ;
      RECT 55.815 2.465 55.82 3.063 ;
      RECT 55.805 2.495 55.815 3.082 ;
      RECT 55.795 2.52 55.805 3.107 ;
      RECT 55.79 2.54 55.795 3.126 ;
      RECT 55.785 2.557 55.79 3.139 ;
      RECT 55.775 2.583 55.785 3.158 ;
      RECT 55.765 2.621 55.775 3.185 ;
      RECT 55.76 2.647 55.765 3.205 ;
      RECT 55.755 2.657 55.76 3.215 ;
      RECT 55.75 2.67 55.755 3.23 ;
      RECT 55.745 2.685 55.75 3.24 ;
      RECT 55.74 2.707 55.745 3.255 ;
      RECT 55.735 2.725 55.74 3.266 ;
      RECT 55.73 2.735 55.735 3.277 ;
      RECT 55.725 2.743 55.73 3.289 ;
      RECT 55.72 2.751 55.725 3.3 ;
      RECT 55.715 2.777 55.72 3.313 ;
      RECT 55.705 2.805 55.715 3.326 ;
      RECT 55.7 2.835 55.705 3.335 ;
      RECT 55.695 2.85 55.7 3.342 ;
      RECT 55.68 2.875 55.695 3.349 ;
      RECT 55.675 2.897 55.68 3.355 ;
      RECT 55.67 2.922 55.675 3.358 ;
      RECT 55.661 2.95 55.67 3.362 ;
      RECT 55.655 2.967 55.661 3.367 ;
      RECT 55.65 2.985 55.655 3.371 ;
      RECT 55.645 2.997 55.65 3.374 ;
      RECT 55.64 3.018 55.645 3.378 ;
      RECT 55.635 3.036 55.64 3.381 ;
      RECT 55.63 3.05 55.635 3.384 ;
      RECT 55.625 3.067 55.63 3.387 ;
      RECT 55.62 3.08 55.625 3.39 ;
      RECT 55.595 3.117 55.62 3.398 ;
      RECT 55.59 3.162 55.595 3.407 ;
      RECT 55.585 3.19 55.59 3.41 ;
      RECT 55.575 3.21 55.585 3.414 ;
      RECT 55.57 3.23 55.575 3.419 ;
      RECT 55.565 3.245 55.57 3.422 ;
      RECT 55.545 3.255 55.565 3.429 ;
      RECT 55.48 3.262 55.545 3.455 ;
      RECT 55.445 3.265 55.48 3.483 ;
      RECT 55.43 3.268 55.445 3.498 ;
      RECT 55.42 3.269 55.43 3.513 ;
      RECT 55.41 3.27 55.42 3.53 ;
      RECT 55.405 3.27 55.41 3.545 ;
      RECT 55.4 3.27 55.405 3.553 ;
      RECT 55.385 3.271 55.4 3.568 ;
      RECT 55.355 3.273 55.385 3.575 ;
      RECT 55.245 3.28 55.325 3.575 ;
      RECT 55.2 3.285 55.245 3.575 ;
      RECT 55.19 3.286 55.2 3.565 ;
      RECT 55.18 3.287 55.19 3.558 ;
      RECT 55.16 3.289 55.18 3.553 ;
      RECT 55.15 3.26 55.16 3.548 ;
      RECT 55.105 3.26 55.15 3.54 ;
      RECT 55.075 3.26 55.1 3.53 ;
      RECT 55.055 3.26 55.075 3.523 ;
      RECT 55.335 2.06 55.595 2.32 ;
      RECT 55.215 2.075 55.225 2.24 ;
      RECT 55.2 2.075 55.205 2.235 ;
      RECT 52.565 1.915 52.75 2.205 ;
      RECT 54.38 2.04 54.395 2.195 ;
      RECT 52.53 1.915 52.555 2.175 ;
      RECT 54.945 1.965 54.95 2.107 ;
      RECT 54.86 1.96 54.885 2.1 ;
      RECT 55.26 2.077 55.335 2.27 ;
      RECT 55.245 2.075 55.26 2.253 ;
      RECT 55.225 2.075 55.245 2.245 ;
      RECT 55.205 2.075 55.215 2.238 ;
      RECT 55.16 2.07 55.2 2.228 ;
      RECT 55.12 2.045 55.16 2.213 ;
      RECT 55.105 2.02 55.12 2.203 ;
      RECT 55.1 2.014 55.105 2.201 ;
      RECT 55.065 2.006 55.1 2.184 ;
      RECT 55.06 1.999 55.065 2.172 ;
      RECT 55.04 1.994 55.06 2.16 ;
      RECT 55.03 1.988 55.04 2.145 ;
      RECT 55.01 1.983 55.03 2.13 ;
      RECT 55 1.978 55.01 2.123 ;
      RECT 54.995 1.976 55 2.118 ;
      RECT 54.99 1.975 54.995 2.115 ;
      RECT 54.95 1.97 54.99 2.111 ;
      RECT 54.93 1.964 54.945 2.106 ;
      RECT 54.895 1.961 54.93 2.103 ;
      RECT 54.885 1.96 54.895 2.101 ;
      RECT 54.825 1.96 54.86 2.098 ;
      RECT 54.78 1.96 54.825 2.098 ;
      RECT 54.73 1.96 54.78 2.101 ;
      RECT 54.715 1.962 54.73 2.103 ;
      RECT 54.7 1.965 54.715 2.104 ;
      RECT 54.69 1.97 54.7 2.105 ;
      RECT 54.66 1.975 54.69 2.11 ;
      RECT 54.65 1.981 54.66 2.118 ;
      RECT 54.64 1.983 54.65 2.122 ;
      RECT 54.63 1.987 54.64 2.126 ;
      RECT 54.605 1.993 54.63 2.134 ;
      RECT 54.595 1.998 54.605 2.142 ;
      RECT 54.58 2.002 54.595 2.146 ;
      RECT 54.545 2.008 54.58 2.154 ;
      RECT 54.525 2.013 54.545 2.164 ;
      RECT 54.495 2.02 54.525 2.173 ;
      RECT 54.45 2.029 54.495 2.187 ;
      RECT 54.445 2.034 54.45 2.198 ;
      RECT 54.425 2.037 54.445 2.199 ;
      RECT 54.395 2.04 54.425 2.197 ;
      RECT 54.36 2.04 54.38 2.193 ;
      RECT 54.29 2.04 54.36 2.184 ;
      RECT 54.275 2.037 54.29 2.176 ;
      RECT 54.235 2.03 54.275 2.171 ;
      RECT 54.21 2.02 54.235 2.164 ;
      RECT 54.205 2.014 54.21 2.161 ;
      RECT 54.165 2.008 54.205 2.158 ;
      RECT 54.15 2.001 54.165 2.153 ;
      RECT 54.13 1.997 54.15 2.148 ;
      RECT 54.115 1.992 54.13 2.144 ;
      RECT 54.1 1.987 54.115 2.142 ;
      RECT 54.085 1.983 54.1 2.141 ;
      RECT 54.07 1.981 54.085 2.137 ;
      RECT 54.06 1.979 54.07 2.132 ;
      RECT 54.045 1.976 54.06 2.128 ;
      RECT 54.035 1.974 54.045 2.123 ;
      RECT 54.015 1.971 54.035 2.119 ;
      RECT 53.97 1.97 54.015 2.117 ;
      RECT 53.91 1.972 53.97 2.118 ;
      RECT 53.89 1.974 53.91 2.12 ;
      RECT 53.86 1.977 53.89 2.121 ;
      RECT 53.81 1.982 53.86 2.123 ;
      RECT 53.805 1.985 53.81 2.125 ;
      RECT 53.795 1.987 53.805 2.128 ;
      RECT 53.79 1.989 53.795 2.131 ;
      RECT 53.74 1.992 53.79 2.138 ;
      RECT 53.72 1.996 53.74 2.15 ;
      RECT 53.71 1.999 53.72 2.156 ;
      RECT 53.7 2 53.71 2.159 ;
      RECT 53.661 2.003 53.7 2.161 ;
      RECT 53.575 2.01 53.661 2.164 ;
      RECT 53.501 2.02 53.575 2.168 ;
      RECT 53.415 2.031 53.501 2.173 ;
      RECT 53.4 2.038 53.415 2.175 ;
      RECT 53.345 2.042 53.4 2.176 ;
      RECT 53.331 2.045 53.345 2.178 ;
      RECT 53.245 2.045 53.331 2.18 ;
      RECT 53.205 2.042 53.245 2.183 ;
      RECT 53.181 2.038 53.205 2.185 ;
      RECT 53.095 2.028 53.181 2.188 ;
      RECT 53.065 2.017 53.095 2.189 ;
      RECT 53.046 2.013 53.065 2.188 ;
      RECT 52.96 2.006 53.046 2.185 ;
      RECT 52.9 1.995 52.96 2.182 ;
      RECT 52.88 1.987 52.9 2.18 ;
      RECT 52.845 1.982 52.88 2.179 ;
      RECT 52.82 1.977 52.845 2.178 ;
      RECT 52.79 1.972 52.82 2.177 ;
      RECT 52.765 1.915 52.79 2.176 ;
      RECT 52.75 1.915 52.765 2.2 ;
      RECT 52.555 1.915 52.565 2.2 ;
      RECT 54.33 2.935 54.335 3.075 ;
      RECT 53.99 2.935 54.025 3.073 ;
      RECT 53.565 2.92 53.58 3.065 ;
      RECT 55.395 2.7 55.485 2.96 ;
      RECT 55.225 2.565 55.325 2.96 ;
      RECT 52.26 2.54 52.34 2.75 ;
      RECT 55.35 2.677 55.395 2.96 ;
      RECT 55.34 2.647 55.35 2.96 ;
      RECT 55.325 2.57 55.34 2.96 ;
      RECT 55.14 2.565 55.225 2.925 ;
      RECT 55.135 2.567 55.14 2.92 ;
      RECT 55.13 2.572 55.135 2.92 ;
      RECT 55.095 2.672 55.13 2.92 ;
      RECT 55.085 2.7 55.095 2.92 ;
      RECT 55.075 2.715 55.085 2.92 ;
      RECT 55.065 2.727 55.075 2.92 ;
      RECT 55.06 2.737 55.065 2.92 ;
      RECT 55.045 2.747 55.06 2.922 ;
      RECT 55.04 2.762 55.045 2.924 ;
      RECT 55.025 2.775 55.04 2.926 ;
      RECT 55.02 2.79 55.025 2.929 ;
      RECT 55 2.8 55.02 2.933 ;
      RECT 54.985 2.81 55 2.936 ;
      RECT 54.95 2.817 54.985 2.941 ;
      RECT 54.906 2.824 54.95 2.949 ;
      RECT 54.82 2.836 54.906 2.962 ;
      RECT 54.795 2.847 54.82 2.973 ;
      RECT 54.765 2.852 54.795 2.978 ;
      RECT 54.73 2.857 54.765 2.986 ;
      RECT 54.7 2.862 54.73 2.993 ;
      RECT 54.675 2.867 54.7 2.998 ;
      RECT 54.61 2.874 54.675 3.007 ;
      RECT 54.54 2.887 54.61 3.023 ;
      RECT 54.51 2.897 54.54 3.035 ;
      RECT 54.485 2.902 54.51 3.042 ;
      RECT 54.43 2.909 54.485 3.05 ;
      RECT 54.425 2.916 54.43 3.055 ;
      RECT 54.42 2.918 54.425 3.056 ;
      RECT 54.405 2.92 54.42 3.058 ;
      RECT 54.4 2.92 54.405 3.061 ;
      RECT 54.335 2.927 54.4 3.068 ;
      RECT 54.3 2.937 54.33 3.078 ;
      RECT 54.283 2.94 54.3 3.08 ;
      RECT 54.197 2.939 54.283 3.079 ;
      RECT 54.111 2.937 54.197 3.076 ;
      RECT 54.025 2.936 54.111 3.074 ;
      RECT 53.924 2.934 53.99 3.073 ;
      RECT 53.838 2.931 53.924 3.071 ;
      RECT 53.752 2.927 53.838 3.069 ;
      RECT 53.666 2.924 53.752 3.068 ;
      RECT 53.58 2.921 53.666 3.066 ;
      RECT 53.48 2.92 53.565 3.063 ;
      RECT 53.43 2.918 53.48 3.061 ;
      RECT 53.41 2.915 53.43 3.059 ;
      RECT 53.39 2.913 53.41 3.056 ;
      RECT 53.365 2.909 53.39 3.053 ;
      RECT 53.32 2.903 53.365 3.048 ;
      RECT 53.28 2.897 53.32 3.04 ;
      RECT 53.255 2.892 53.28 3.033 ;
      RECT 53.2 2.885 53.255 3.025 ;
      RECT 53.176 2.878 53.2 3.018 ;
      RECT 53.09 2.869 53.176 3.008 ;
      RECT 53.06 2.861 53.09 2.998 ;
      RECT 53.03 2.857 53.06 2.993 ;
      RECT 53.025 2.854 53.03 2.99 ;
      RECT 53.02 2.853 53.025 2.99 ;
      RECT 52.945 2.846 53.02 2.983 ;
      RECT 52.906 2.837 52.945 2.972 ;
      RECT 52.82 2.827 52.906 2.96 ;
      RECT 52.78 2.817 52.82 2.948 ;
      RECT 52.741 2.812 52.78 2.941 ;
      RECT 52.655 2.802 52.741 2.93 ;
      RECT 52.615 2.79 52.655 2.919 ;
      RECT 52.58 2.775 52.615 2.912 ;
      RECT 52.57 2.765 52.58 2.909 ;
      RECT 52.55 2.75 52.57 2.907 ;
      RECT 52.52 2.72 52.55 2.903 ;
      RECT 52.51 2.7 52.52 2.898 ;
      RECT 52.505 2.692 52.51 2.895 ;
      RECT 52.5 2.685 52.505 2.893 ;
      RECT 52.485 2.672 52.5 2.886 ;
      RECT 52.48 2.662 52.485 2.878 ;
      RECT 52.475 2.655 52.48 2.873 ;
      RECT 52.47 2.65 52.475 2.869 ;
      RECT 52.455 2.637 52.47 2.861 ;
      RECT 52.45 2.547 52.455 2.85 ;
      RECT 52.445 2.542 52.45 2.843 ;
      RECT 52.37 2.54 52.445 2.803 ;
      RECT 52.34 2.54 52.37 2.758 ;
      RECT 52.245 2.545 52.26 2.745 ;
      RECT 54.73 2.25 54.99 2.51 ;
      RECT 54.715 2.238 54.895 2.475 ;
      RECT 54.71 2.239 54.895 2.473 ;
      RECT 54.695 2.243 54.905 2.463 ;
      RECT 54.69 2.248 54.91 2.433 ;
      RECT 54.695 2.245 54.91 2.463 ;
      RECT 54.71 2.24 54.905 2.473 ;
      RECT 54.73 2.237 54.895 2.51 ;
      RECT 54.73 2.236 54.885 2.51 ;
      RECT 54.755 2.235 54.885 2.51 ;
      RECT 54.315 2.48 54.575 2.74 ;
      RECT 54.19 2.525 54.575 2.735 ;
      RECT 54.18 2.53 54.575 2.73 ;
      RECT 54.195 3.47 54.21 3.78 ;
      RECT 52.79 3.24 52.8 3.37 ;
      RECT 52.57 3.235 52.675 3.37 ;
      RECT 52.485 3.24 52.535 3.37 ;
      RECT 51.035 1.975 51.04 3.08 ;
      RECT 54.29 3.562 54.295 3.698 ;
      RECT 54.285 3.557 54.29 3.758 ;
      RECT 54.28 3.555 54.285 3.771 ;
      RECT 54.265 3.552 54.28 3.773 ;
      RECT 54.26 3.547 54.265 3.775 ;
      RECT 54.255 3.543 54.26 3.778 ;
      RECT 54.24 3.538 54.255 3.78 ;
      RECT 54.21 3.53 54.24 3.78 ;
      RECT 54.171 3.47 54.195 3.78 ;
      RECT 54.085 3.47 54.171 3.777 ;
      RECT 54.055 3.47 54.085 3.77 ;
      RECT 54.03 3.47 54.055 3.763 ;
      RECT 54.005 3.47 54.03 3.755 ;
      RECT 53.99 3.47 54.005 3.748 ;
      RECT 53.965 3.47 53.99 3.74 ;
      RECT 53.95 3.47 53.965 3.733 ;
      RECT 53.91 3.48 53.95 3.722 ;
      RECT 53.9 3.475 53.91 3.712 ;
      RECT 53.896 3.474 53.9 3.709 ;
      RECT 53.81 3.466 53.896 3.692 ;
      RECT 53.777 3.455 53.81 3.669 ;
      RECT 53.691 3.444 53.777 3.647 ;
      RECT 53.605 3.428 53.691 3.616 ;
      RECT 53.535 3.413 53.605 3.588 ;
      RECT 53.525 3.406 53.535 3.575 ;
      RECT 53.495 3.403 53.525 3.565 ;
      RECT 53.47 3.399 53.495 3.558 ;
      RECT 53.455 3.396 53.47 3.553 ;
      RECT 53.45 3.395 53.455 3.548 ;
      RECT 53.42 3.39 53.45 3.541 ;
      RECT 53.415 3.385 53.42 3.536 ;
      RECT 53.4 3.382 53.415 3.531 ;
      RECT 53.395 3.377 53.4 3.526 ;
      RECT 53.375 3.372 53.395 3.523 ;
      RECT 53.36 3.367 53.375 3.515 ;
      RECT 53.345 3.361 53.36 3.51 ;
      RECT 53.315 3.352 53.345 3.503 ;
      RECT 53.31 3.345 53.315 3.495 ;
      RECT 53.305 3.343 53.31 3.493 ;
      RECT 53.3 3.342 53.305 3.49 ;
      RECT 53.26 3.335 53.3 3.483 ;
      RECT 53.246 3.325 53.26 3.473 ;
      RECT 53.195 3.314 53.246 3.461 ;
      RECT 53.17 3.3 53.195 3.447 ;
      RECT 53.145 3.289 53.17 3.439 ;
      RECT 53.125 3.278 53.145 3.433 ;
      RECT 53.115 3.272 53.125 3.428 ;
      RECT 53.11 3.27 53.115 3.424 ;
      RECT 53.09 3.265 53.11 3.419 ;
      RECT 53.06 3.255 53.09 3.409 ;
      RECT 53.055 3.247 53.06 3.402 ;
      RECT 53.04 3.245 53.055 3.398 ;
      RECT 53.02 3.245 53.04 3.393 ;
      RECT 53.015 3.244 53.02 3.391 ;
      RECT 53.01 3.244 53.015 3.388 ;
      RECT 52.97 3.243 53.01 3.383 ;
      RECT 52.945 3.242 52.97 3.378 ;
      RECT 52.885 3.241 52.945 3.375 ;
      RECT 52.8 3.24 52.885 3.373 ;
      RECT 52.761 3.239 52.79 3.37 ;
      RECT 52.675 3.237 52.761 3.37 ;
      RECT 52.535 3.237 52.57 3.37 ;
      RECT 52.445 3.241 52.485 3.373 ;
      RECT 52.43 3.244 52.445 3.38 ;
      RECT 52.42 3.245 52.43 3.387 ;
      RECT 52.395 3.248 52.42 3.392 ;
      RECT 52.39 3.25 52.395 3.395 ;
      RECT 52.34 3.252 52.39 3.396 ;
      RECT 52.301 3.256 52.34 3.398 ;
      RECT 52.215 3.258 52.301 3.401 ;
      RECT 52.197 3.26 52.215 3.403 ;
      RECT 52.111 3.263 52.197 3.405 ;
      RECT 52.025 3.267 52.111 3.408 ;
      RECT 51.988 3.271 52.025 3.411 ;
      RECT 51.902 3.274 51.988 3.414 ;
      RECT 51.816 3.278 51.902 3.417 ;
      RECT 51.73 3.283 51.816 3.421 ;
      RECT 51.71 3.285 51.73 3.424 ;
      RECT 51.69 3.284 51.71 3.425 ;
      RECT 51.641 3.281 51.69 3.426 ;
      RECT 51.555 3.276 51.641 3.429 ;
      RECT 51.505 3.271 51.555 3.431 ;
      RECT 51.481 3.269 51.505 3.432 ;
      RECT 51.395 3.264 51.481 3.434 ;
      RECT 51.37 3.26 51.395 3.433 ;
      RECT 51.36 3.257 51.37 3.431 ;
      RECT 51.35 3.25 51.36 3.428 ;
      RECT 51.345 3.23 51.35 3.423 ;
      RECT 51.335 3.2 51.345 3.418 ;
      RECT 51.32 3.07 51.335 3.409 ;
      RECT 51.315 3.062 51.32 3.402 ;
      RECT 51.295 3.055 51.315 3.394 ;
      RECT 51.29 3.037 51.295 3.386 ;
      RECT 51.28 3.017 51.29 3.381 ;
      RECT 51.275 2.99 51.28 3.377 ;
      RECT 51.27 2.967 51.275 3.374 ;
      RECT 51.25 2.925 51.27 3.366 ;
      RECT 51.215 2.84 51.25 3.35 ;
      RECT 51.21 2.772 51.215 3.338 ;
      RECT 51.195 2.742 51.21 3.332 ;
      RECT 51.19 1.987 51.195 2.233 ;
      RECT 51.18 2.712 51.195 3.323 ;
      RECT 51.185 1.982 51.19 2.265 ;
      RECT 51.18 1.977 51.185 2.308 ;
      RECT 51.175 1.975 51.18 2.343 ;
      RECT 51.16 2.675 51.18 3.313 ;
      RECT 51.17 1.975 51.175 2.38 ;
      RECT 51.155 1.975 51.17 2.478 ;
      RECT 51.155 2.648 51.16 3.306 ;
      RECT 51.15 1.975 51.155 2.553 ;
      RECT 51.15 2.636 51.155 3.303 ;
      RECT 51.145 1.975 51.15 2.585 ;
      RECT 51.145 2.615 51.15 3.3 ;
      RECT 51.14 1.975 51.145 3.297 ;
      RECT 51.105 1.975 51.14 3.283 ;
      RECT 51.09 1.975 51.105 3.265 ;
      RECT 51.07 1.975 51.09 3.255 ;
      RECT 51.045 1.975 51.07 3.238 ;
      RECT 51.04 1.975 51.045 3.188 ;
      RECT 51.03 1.975 51.035 3.018 ;
      RECT 51.025 1.975 51.03 2.925 ;
      RECT 51.02 1.975 51.025 2.838 ;
      RECT 51.015 1.975 51.02 2.77 ;
      RECT 51.01 1.975 51.015 2.713 ;
      RECT 51 1.975 51.01 2.608 ;
      RECT 50.995 1.975 51 2.48 ;
      RECT 50.99 1.975 50.995 2.398 ;
      RECT 50.985 1.977 50.99 2.315 ;
      RECT 50.98 1.982 50.985 2.248 ;
      RECT 50.975 1.987 50.98 2.175 ;
      RECT 53.79 2.305 54.05 2.565 ;
      RECT 53.81 2.272 54.02 2.565 ;
      RECT 53.81 2.27 54.01 2.565 ;
      RECT 53.82 2.257 54.01 2.565 ;
      RECT 53.82 2.255 53.935 2.565 ;
      RECT 53.295 2.38 53.47 2.66 ;
      RECT 53.29 2.38 53.47 2.658 ;
      RECT 53.29 2.38 53.485 2.655 ;
      RECT 53.28 2.38 53.485 2.653 ;
      RECT 53.225 2.38 53.485 2.64 ;
      RECT 53.225 2.455 53.49 2.618 ;
      RECT 52.77 2.392 52.79 2.635 ;
      RECT 52.77 2.392 52.83 2.634 ;
      RECT 52.765 2.394 52.83 2.633 ;
      RECT 52.765 2.394 52.916 2.632 ;
      RECT 52.765 2.394 52.985 2.631 ;
      RECT 52.765 2.394 53.005 2.623 ;
      RECT 52.745 2.397 53.005 2.621 ;
      RECT 52.73 2.407 53.005 2.606 ;
      RECT 52.73 2.407 53.02 2.605 ;
      RECT 52.725 2.416 53.02 2.597 ;
      RECT 52.725 2.416 53.025 2.593 ;
      RECT 52.83 2.33 53.09 2.59 ;
      RECT 52.72 2.418 53.09 2.475 ;
      RECT 52.79 2.385 53.09 2.59 ;
      RECT 52.755 3.578 52.76 3.785 ;
      RECT 52.705 3.572 52.755 3.784 ;
      RECT 52.672 3.586 52.765 3.783 ;
      RECT 52.586 3.586 52.765 3.782 ;
      RECT 52.5 3.586 52.765 3.781 ;
      RECT 52.5 3.685 52.77 3.778 ;
      RECT 52.495 3.685 52.77 3.773 ;
      RECT 52.49 3.685 52.77 3.755 ;
      RECT 52.485 3.685 52.77 3.738 ;
      RECT 52.445 3.47 52.705 3.73 ;
      RECT 51.905 2.62 51.991 3.034 ;
      RECT 51.905 2.62 52.03 3.031 ;
      RECT 51.905 2.62 52.05 3.021 ;
      RECT 51.86 2.62 52.05 3.018 ;
      RECT 51.86 2.772 52.06 3.008 ;
      RECT 51.86 2.793 52.065 3.002 ;
      RECT 51.86 2.811 52.07 2.998 ;
      RECT 51.86 2.831 52.08 2.993 ;
      RECT 51.835 2.831 52.08 2.99 ;
      RECT 51.825 2.831 52.08 2.968 ;
      RECT 51.825 2.847 52.085 2.938 ;
      RECT 51.79 2.62 52.05 2.925 ;
      RECT 51.79 2.859 52.09 2.88 ;
      RECT 49.45 7.77 49.74 8 ;
      RECT 49.51 6.29 49.68 8 ;
      RECT 49.46 6.655 49.81 7.005 ;
      RECT 49.45 6.29 49.74 6.52 ;
      RECT 49.045 2.395 49.15 2.965 ;
      RECT 49.045 2.73 49.37 2.96 ;
      RECT 49.045 2.76 49.54 2.93 ;
      RECT 49.045 2.395 49.235 2.96 ;
      RECT 48.46 2.36 48.75 2.59 ;
      RECT 48.46 2.395 49.235 2.565 ;
      RECT 48.52 0.88 48.69 2.59 ;
      RECT 48.46 0.88 48.75 1.11 ;
      RECT 48.46 7.77 48.75 8 ;
      RECT 48.52 6.29 48.69 8 ;
      RECT 48.46 6.29 48.75 6.52 ;
      RECT 48.46 6.325 49.315 6.485 ;
      RECT 49.145 5.92 49.315 6.485 ;
      RECT 48.46 6.32 48.855 6.485 ;
      RECT 49.08 5.92 49.37 6.15 ;
      RECT 49.08 5.95 49.54 6.12 ;
      RECT 48.09 2.73 48.38 2.96 ;
      RECT 48.09 2.76 48.55 2.93 ;
      RECT 48.155 1.655 48.32 2.96 ;
      RECT 46.67 1.625 46.96 1.855 ;
      RECT 46.67 1.655 48.32 1.825 ;
      RECT 46.73 0.885 46.9 1.855 ;
      RECT 46.67 0.885 46.96 1.115 ;
      RECT 46.67 7.765 46.96 7.995 ;
      RECT 46.73 7.025 46.9 7.995 ;
      RECT 46.73 7.12 48.32 7.29 ;
      RECT 48.15 5.92 48.32 7.29 ;
      RECT 46.67 7.025 46.96 7.255 ;
      RECT 48.09 5.92 48.38 6.15 ;
      RECT 48.09 5.95 48.55 6.12 ;
      RECT 44.72 2.705 45.06 3.055 ;
      RECT 44.81 2.025 44.98 3.055 ;
      RECT 47.1 1.965 47.45 2.315 ;
      RECT 44.81 2.025 47.45 2.195 ;
      RECT 47.125 6.655 47.45 6.98 ;
      RECT 41.665 6.615 42.015 6.965 ;
      RECT 47.1 6.655 47.45 6.885 ;
      RECT 41.465 6.655 42.015 6.885 ;
      RECT 41.295 6.685 47.45 6.855 ;
      RECT 46.325 2.365 46.645 2.685 ;
      RECT 46.295 2.365 46.645 2.595 ;
      RECT 46.125 2.395 46.645 2.565 ;
      RECT 46.325 6.255 46.645 6.545 ;
      RECT 46.295 6.285 46.645 6.515 ;
      RECT 46.125 6.315 46.645 6.485 ;
      RECT 42.015 2.985 42.165 3.26 ;
      RECT 42.555 2.065 42.56 2.285 ;
      RECT 43.705 2.265 43.72 2.463 ;
      RECT 43.67 2.257 43.705 2.47 ;
      RECT 43.64 2.25 43.67 2.47 ;
      RECT 43.585 2.215 43.64 2.47 ;
      RECT 43.52 2.152 43.585 2.47 ;
      RECT 43.515 2.117 43.52 2.468 ;
      RECT 43.51 2.112 43.515 2.46 ;
      RECT 43.505 2.107 43.51 2.446 ;
      RECT 43.5 2.104 43.505 2.439 ;
      RECT 43.455 2.094 43.5 2.39 ;
      RECT 43.435 2.081 43.455 2.325 ;
      RECT 43.43 2.076 43.435 2.298 ;
      RECT 43.425 2.075 43.43 2.291 ;
      RECT 43.42 2.074 43.425 2.284 ;
      RECT 43.335 2.059 43.42 2.23 ;
      RECT 43.305 2.04 43.335 2.18 ;
      RECT 43.225 2.023 43.305 2.165 ;
      RECT 43.19 2.01 43.225 2.15 ;
      RECT 43.182 2.01 43.19 2.145 ;
      RECT 43.096 2.011 43.182 2.145 ;
      RECT 43.01 2.013 43.096 2.145 ;
      RECT 42.985 2.014 43.01 2.149 ;
      RECT 42.91 2.02 42.985 2.164 ;
      RECT 42.827 2.032 42.91 2.188 ;
      RECT 42.741 2.045 42.827 2.214 ;
      RECT 42.655 2.058 42.741 2.24 ;
      RECT 42.62 2.067 42.655 2.259 ;
      RECT 42.57 2.067 42.62 2.272 ;
      RECT 42.56 2.065 42.57 2.283 ;
      RECT 42.545 2.062 42.555 2.285 ;
      RECT 42.53 2.054 42.545 2.293 ;
      RECT 42.515 2.046 42.53 2.313 ;
      RECT 42.51 2.041 42.515 2.37 ;
      RECT 42.495 2.036 42.51 2.443 ;
      RECT 42.49 2.031 42.495 2.485 ;
      RECT 42.485 2.029 42.49 2.513 ;
      RECT 42.48 2.027 42.485 2.535 ;
      RECT 42.47 2.023 42.48 2.578 ;
      RECT 42.465 2.02 42.47 2.603 ;
      RECT 42.46 2.018 42.465 2.623 ;
      RECT 42.455 2.016 42.46 2.647 ;
      RECT 42.45 2.012 42.455 2.67 ;
      RECT 42.445 2.008 42.45 2.693 ;
      RECT 42.41 1.998 42.445 2.8 ;
      RECT 42.405 1.988 42.41 2.898 ;
      RECT 42.4 1.986 42.405 2.925 ;
      RECT 42.395 1.985 42.4 2.945 ;
      RECT 42.39 1.977 42.395 2.965 ;
      RECT 42.385 1.972 42.39 3 ;
      RECT 42.38 1.97 42.385 3.018 ;
      RECT 42.375 1.97 42.38 3.043 ;
      RECT 42.37 1.97 42.375 3.065 ;
      RECT 42.335 1.97 42.37 3.108 ;
      RECT 42.31 1.97 42.335 3.137 ;
      RECT 42.3 1.97 42.31 2.323 ;
      RECT 42.303 2.38 42.31 3.147 ;
      RECT 42.3 2.437 42.303 3.15 ;
      RECT 42.295 1.97 42.3 2.295 ;
      RECT 42.295 2.487 42.3 3.153 ;
      RECT 42.285 1.97 42.295 2.285 ;
      RECT 42.29 2.54 42.295 3.156 ;
      RECT 42.285 2.625 42.29 3.16 ;
      RECT 42.275 1.97 42.285 2.273 ;
      RECT 42.28 2.672 42.285 3.164 ;
      RECT 42.275 2.747 42.28 3.168 ;
      RECT 42.24 1.97 42.275 2.248 ;
      RECT 42.265 2.83 42.275 3.173 ;
      RECT 42.255 2.897 42.265 3.18 ;
      RECT 42.25 2.925 42.255 3.185 ;
      RECT 42.24 2.938 42.25 3.191 ;
      RECT 42.195 1.97 42.24 2.205 ;
      RECT 42.235 2.943 42.24 3.198 ;
      RECT 42.195 2.96 42.235 3.26 ;
      RECT 42.19 1.972 42.195 2.178 ;
      RECT 42.165 2.98 42.195 3.26 ;
      RECT 42.185 1.977 42.19 2.15 ;
      RECT 41.975 2.989 42.015 3.26 ;
      RECT 41.95 2.997 41.975 3.23 ;
      RECT 41.905 3.005 41.95 3.23 ;
      RECT 41.89 3.01 41.905 3.225 ;
      RECT 41.88 3.01 41.89 3.219 ;
      RECT 41.87 3.017 41.88 3.216 ;
      RECT 41.865 3.055 41.87 3.205 ;
      RECT 41.86 3.117 41.865 3.183 ;
      RECT 43.13 2.992 43.315 3.215 ;
      RECT 43.13 3.007 43.32 3.211 ;
      RECT 43.12 2.28 43.205 3.21 ;
      RECT 43.12 3.007 43.325 3.204 ;
      RECT 43.115 3.015 43.325 3.203 ;
      RECT 43.32 2.735 43.64 3.055 ;
      RECT 43.115 2.907 43.285 2.998 ;
      RECT 43.11 2.907 43.285 2.98 ;
      RECT 43.1 2.715 43.235 2.955 ;
      RECT 43.095 2.715 43.235 2.9 ;
      RECT 43.055 2.295 43.225 2.8 ;
      RECT 43.04 2.295 43.225 2.67 ;
      RECT 43.035 2.295 43.225 2.623 ;
      RECT 43.03 2.295 43.225 2.603 ;
      RECT 43.025 2.295 43.225 2.578 ;
      RECT 42.995 2.295 43.255 2.555 ;
      RECT 43.005 2.292 43.215 2.555 ;
      RECT 43.13 2.287 43.215 3.215 ;
      RECT 43.015 2.28 43.205 2.555 ;
      RECT 43.01 2.285 43.205 2.555 ;
      RECT 41.84 2.497 42.025 2.71 ;
      RECT 41.84 2.505 42.035 2.703 ;
      RECT 41.82 2.505 42.035 2.7 ;
      RECT 41.815 2.505 42.035 2.685 ;
      RECT 41.745 2.42 42.005 2.68 ;
      RECT 41.745 2.565 42.04 2.593 ;
      RECT 41.4 3.02 41.66 3.28 ;
      RECT 41.425 2.965 41.62 3.28 ;
      RECT 41.42 2.714 41.6 3.008 ;
      RECT 41.42 2.72 41.61 3.008 ;
      RECT 41.4 2.722 41.61 2.953 ;
      RECT 41.395 2.732 41.61 2.82 ;
      RECT 41.425 2.712 41.6 3.28 ;
      RECT 41.511 2.71 41.6 3.28 ;
      RECT 41.37 1.93 41.405 2.3 ;
      RECT 41.16 2.04 41.165 2.3 ;
      RECT 41.405 1.937 41.42 2.3 ;
      RECT 41.295 1.93 41.37 2.378 ;
      RECT 41.285 1.93 41.295 2.463 ;
      RECT 41.26 1.93 41.285 2.498 ;
      RECT 41.22 1.93 41.26 2.566 ;
      RECT 41.21 1.937 41.22 2.618 ;
      RECT 41.18 2.04 41.21 2.659 ;
      RECT 41.175 2.04 41.18 2.698 ;
      RECT 41.165 2.04 41.175 2.718 ;
      RECT 41.16 2.335 41.165 2.755 ;
      RECT 41.155 2.352 41.16 2.775 ;
      RECT 41.14 2.415 41.155 2.815 ;
      RECT 41.135 2.458 41.14 2.85 ;
      RECT 41.13 2.466 41.135 2.863 ;
      RECT 41.12 2.48 41.13 2.885 ;
      RECT 41.095 2.515 41.12 2.95 ;
      RECT 41.085 2.55 41.095 3.013 ;
      RECT 41.065 2.58 41.085 3.074 ;
      RECT 41.05 2.616 41.065 3.141 ;
      RECT 41.04 2.644 41.05 3.18 ;
      RECT 41.03 2.666 41.04 3.2 ;
      RECT 41.025 2.676 41.03 3.211 ;
      RECT 41.02 2.685 41.025 3.214 ;
      RECT 41.01 2.703 41.02 3.218 ;
      RECT 41 2.721 41.01 3.219 ;
      RECT 40.975 2.76 41 3.216 ;
      RECT 40.955 2.802 40.975 3.213 ;
      RECT 40.94 2.84 40.955 3.212 ;
      RECT 40.905 2.875 40.94 3.209 ;
      RECT 40.9 2.897 40.905 3.207 ;
      RECT 40.835 2.937 40.9 3.204 ;
      RECT 40.83 2.977 40.835 3.2 ;
      RECT 40.815 2.987 40.83 3.191 ;
      RECT 40.805 3.107 40.815 3.176 ;
      RECT 41.285 3.52 41.295 3.78 ;
      RECT 41.285 3.523 41.305 3.779 ;
      RECT 41.275 3.513 41.285 3.778 ;
      RECT 41.265 3.528 41.345 3.774 ;
      RECT 41.25 3.507 41.265 3.772 ;
      RECT 41.225 3.532 41.35 3.768 ;
      RECT 41.21 3.492 41.225 3.763 ;
      RECT 41.21 3.534 41.36 3.762 ;
      RECT 41.21 3.542 41.375 3.755 ;
      RECT 41.15 3.479 41.21 3.745 ;
      RECT 41.14 3.466 41.15 3.727 ;
      RECT 41.115 3.456 41.14 3.717 ;
      RECT 41.11 3.446 41.115 3.709 ;
      RECT 41.045 3.542 41.375 3.691 ;
      RECT 40.96 3.542 41.375 3.653 ;
      RECT 40.85 3.37 41.11 3.63 ;
      RECT 41.225 3.5 41.25 3.768 ;
      RECT 41.265 3.51 41.275 3.774 ;
      RECT 40.85 3.518 41.29 3.63 ;
      RECT 41.035 7.765 41.325 7.995 ;
      RECT 41.095 7.025 41.265 7.995 ;
      RECT 40.995 7.055 41.365 7.425 ;
      RECT 41.035 7.025 41.325 7.425 ;
      RECT 40.065 3.275 40.095 3.575 ;
      RECT 39.84 3.26 39.845 3.535 ;
      RECT 39.64 3.26 39.795 3.52 ;
      RECT 40.94 1.975 40.97 2.235 ;
      RECT 40.93 1.975 40.94 2.343 ;
      RECT 40.91 1.975 40.93 2.353 ;
      RECT 40.895 1.975 40.91 2.365 ;
      RECT 40.84 1.975 40.895 2.415 ;
      RECT 40.825 1.975 40.84 2.463 ;
      RECT 40.795 1.975 40.825 2.498 ;
      RECT 40.74 1.975 40.795 2.56 ;
      RECT 40.72 1.975 40.74 2.628 ;
      RECT 40.715 1.975 40.72 2.658 ;
      RECT 40.71 1.975 40.715 2.67 ;
      RECT 40.705 2.092 40.71 2.688 ;
      RECT 40.685 2.11 40.705 2.713 ;
      RECT 40.665 2.137 40.685 2.763 ;
      RECT 40.66 2.157 40.665 2.794 ;
      RECT 40.655 2.165 40.66 2.811 ;
      RECT 40.64 2.191 40.655 2.84 ;
      RECT 40.625 2.233 40.64 2.875 ;
      RECT 40.62 2.262 40.625 2.898 ;
      RECT 40.615 2.277 40.62 2.911 ;
      RECT 40.61 2.3 40.615 2.922 ;
      RECT 40.6 2.32 40.61 2.94 ;
      RECT 40.59 2.35 40.6 2.963 ;
      RECT 40.585 2.372 40.59 2.983 ;
      RECT 40.58 2.387 40.585 2.998 ;
      RECT 40.565 2.417 40.58 3.025 ;
      RECT 40.56 2.447 40.565 3.051 ;
      RECT 40.555 2.465 40.56 3.063 ;
      RECT 40.545 2.495 40.555 3.082 ;
      RECT 40.535 2.52 40.545 3.107 ;
      RECT 40.53 2.54 40.535 3.126 ;
      RECT 40.525 2.557 40.53 3.139 ;
      RECT 40.515 2.583 40.525 3.158 ;
      RECT 40.505 2.621 40.515 3.185 ;
      RECT 40.5 2.647 40.505 3.205 ;
      RECT 40.495 2.657 40.5 3.215 ;
      RECT 40.49 2.67 40.495 3.23 ;
      RECT 40.485 2.685 40.49 3.24 ;
      RECT 40.48 2.707 40.485 3.255 ;
      RECT 40.475 2.725 40.48 3.266 ;
      RECT 40.47 2.735 40.475 3.277 ;
      RECT 40.465 2.743 40.47 3.289 ;
      RECT 40.46 2.751 40.465 3.3 ;
      RECT 40.455 2.777 40.46 3.313 ;
      RECT 40.445 2.805 40.455 3.326 ;
      RECT 40.44 2.835 40.445 3.335 ;
      RECT 40.435 2.85 40.44 3.342 ;
      RECT 40.42 2.875 40.435 3.349 ;
      RECT 40.415 2.897 40.42 3.355 ;
      RECT 40.41 2.922 40.415 3.358 ;
      RECT 40.401 2.95 40.41 3.362 ;
      RECT 40.395 2.967 40.401 3.367 ;
      RECT 40.39 2.985 40.395 3.371 ;
      RECT 40.385 2.997 40.39 3.374 ;
      RECT 40.38 3.018 40.385 3.378 ;
      RECT 40.375 3.036 40.38 3.381 ;
      RECT 40.37 3.05 40.375 3.384 ;
      RECT 40.365 3.067 40.37 3.387 ;
      RECT 40.36 3.08 40.365 3.39 ;
      RECT 40.335 3.117 40.36 3.398 ;
      RECT 40.33 3.162 40.335 3.407 ;
      RECT 40.325 3.19 40.33 3.41 ;
      RECT 40.315 3.21 40.325 3.414 ;
      RECT 40.31 3.23 40.315 3.419 ;
      RECT 40.305 3.245 40.31 3.422 ;
      RECT 40.285 3.255 40.305 3.429 ;
      RECT 40.22 3.262 40.285 3.455 ;
      RECT 40.185 3.265 40.22 3.483 ;
      RECT 40.17 3.268 40.185 3.498 ;
      RECT 40.16 3.269 40.17 3.513 ;
      RECT 40.15 3.27 40.16 3.53 ;
      RECT 40.145 3.27 40.15 3.545 ;
      RECT 40.14 3.27 40.145 3.553 ;
      RECT 40.125 3.271 40.14 3.568 ;
      RECT 40.095 3.273 40.125 3.575 ;
      RECT 39.985 3.28 40.065 3.575 ;
      RECT 39.94 3.285 39.985 3.575 ;
      RECT 39.93 3.286 39.94 3.565 ;
      RECT 39.92 3.287 39.93 3.558 ;
      RECT 39.9 3.289 39.92 3.553 ;
      RECT 39.89 3.26 39.9 3.548 ;
      RECT 39.845 3.26 39.89 3.54 ;
      RECT 39.815 3.26 39.84 3.53 ;
      RECT 39.795 3.26 39.815 3.523 ;
      RECT 40.075 2.06 40.335 2.32 ;
      RECT 39.955 2.075 39.965 2.24 ;
      RECT 39.94 2.075 39.945 2.235 ;
      RECT 37.305 1.915 37.49 2.205 ;
      RECT 39.12 2.04 39.135 2.195 ;
      RECT 37.27 1.915 37.295 2.175 ;
      RECT 39.685 1.965 39.69 2.107 ;
      RECT 39.6 1.96 39.625 2.1 ;
      RECT 40 2.077 40.075 2.27 ;
      RECT 39.985 2.075 40 2.253 ;
      RECT 39.965 2.075 39.985 2.245 ;
      RECT 39.945 2.075 39.955 2.238 ;
      RECT 39.9 2.07 39.94 2.228 ;
      RECT 39.86 2.045 39.9 2.213 ;
      RECT 39.845 2.02 39.86 2.203 ;
      RECT 39.84 2.014 39.845 2.201 ;
      RECT 39.805 2.006 39.84 2.184 ;
      RECT 39.8 1.999 39.805 2.172 ;
      RECT 39.78 1.994 39.8 2.16 ;
      RECT 39.77 1.988 39.78 2.145 ;
      RECT 39.75 1.983 39.77 2.13 ;
      RECT 39.74 1.978 39.75 2.123 ;
      RECT 39.735 1.976 39.74 2.118 ;
      RECT 39.73 1.975 39.735 2.115 ;
      RECT 39.69 1.97 39.73 2.111 ;
      RECT 39.67 1.964 39.685 2.106 ;
      RECT 39.635 1.961 39.67 2.103 ;
      RECT 39.625 1.96 39.635 2.101 ;
      RECT 39.565 1.96 39.6 2.098 ;
      RECT 39.52 1.96 39.565 2.098 ;
      RECT 39.47 1.96 39.52 2.101 ;
      RECT 39.455 1.962 39.47 2.103 ;
      RECT 39.44 1.965 39.455 2.104 ;
      RECT 39.43 1.97 39.44 2.105 ;
      RECT 39.4 1.975 39.43 2.11 ;
      RECT 39.39 1.981 39.4 2.118 ;
      RECT 39.38 1.983 39.39 2.122 ;
      RECT 39.37 1.987 39.38 2.126 ;
      RECT 39.345 1.993 39.37 2.134 ;
      RECT 39.335 1.998 39.345 2.142 ;
      RECT 39.32 2.002 39.335 2.146 ;
      RECT 39.285 2.008 39.32 2.154 ;
      RECT 39.265 2.013 39.285 2.164 ;
      RECT 39.235 2.02 39.265 2.173 ;
      RECT 39.19 2.029 39.235 2.187 ;
      RECT 39.185 2.034 39.19 2.198 ;
      RECT 39.165 2.037 39.185 2.199 ;
      RECT 39.135 2.04 39.165 2.197 ;
      RECT 39.1 2.04 39.12 2.193 ;
      RECT 39.03 2.04 39.1 2.184 ;
      RECT 39.015 2.037 39.03 2.176 ;
      RECT 38.975 2.03 39.015 2.171 ;
      RECT 38.95 2.02 38.975 2.164 ;
      RECT 38.945 2.014 38.95 2.161 ;
      RECT 38.905 2.008 38.945 2.158 ;
      RECT 38.89 2.001 38.905 2.153 ;
      RECT 38.87 1.997 38.89 2.148 ;
      RECT 38.855 1.992 38.87 2.144 ;
      RECT 38.84 1.987 38.855 2.142 ;
      RECT 38.825 1.983 38.84 2.141 ;
      RECT 38.81 1.981 38.825 2.137 ;
      RECT 38.8 1.979 38.81 2.132 ;
      RECT 38.785 1.976 38.8 2.128 ;
      RECT 38.775 1.974 38.785 2.123 ;
      RECT 38.755 1.971 38.775 2.119 ;
      RECT 38.71 1.97 38.755 2.117 ;
      RECT 38.65 1.972 38.71 2.118 ;
      RECT 38.63 1.974 38.65 2.12 ;
      RECT 38.6 1.977 38.63 2.121 ;
      RECT 38.55 1.982 38.6 2.123 ;
      RECT 38.545 1.985 38.55 2.125 ;
      RECT 38.535 1.987 38.545 2.128 ;
      RECT 38.53 1.989 38.535 2.131 ;
      RECT 38.48 1.992 38.53 2.138 ;
      RECT 38.46 1.996 38.48 2.15 ;
      RECT 38.45 1.999 38.46 2.156 ;
      RECT 38.44 2 38.45 2.159 ;
      RECT 38.401 2.003 38.44 2.161 ;
      RECT 38.315 2.01 38.401 2.164 ;
      RECT 38.241 2.02 38.315 2.168 ;
      RECT 38.155 2.031 38.241 2.173 ;
      RECT 38.14 2.038 38.155 2.175 ;
      RECT 38.085 2.042 38.14 2.176 ;
      RECT 38.071 2.045 38.085 2.178 ;
      RECT 37.985 2.045 38.071 2.18 ;
      RECT 37.945 2.042 37.985 2.183 ;
      RECT 37.921 2.038 37.945 2.185 ;
      RECT 37.835 2.028 37.921 2.188 ;
      RECT 37.805 2.017 37.835 2.189 ;
      RECT 37.786 2.013 37.805 2.188 ;
      RECT 37.7 2.006 37.786 2.185 ;
      RECT 37.64 1.995 37.7 2.182 ;
      RECT 37.62 1.987 37.64 2.18 ;
      RECT 37.585 1.982 37.62 2.179 ;
      RECT 37.56 1.977 37.585 2.178 ;
      RECT 37.53 1.972 37.56 2.177 ;
      RECT 37.505 1.915 37.53 2.176 ;
      RECT 37.49 1.915 37.505 2.2 ;
      RECT 37.295 1.915 37.305 2.2 ;
      RECT 39.07 2.935 39.075 3.075 ;
      RECT 38.73 2.935 38.765 3.073 ;
      RECT 38.305 2.92 38.32 3.065 ;
      RECT 40.135 2.7 40.225 2.96 ;
      RECT 39.965 2.565 40.065 2.96 ;
      RECT 37 2.54 37.08 2.75 ;
      RECT 40.09 2.677 40.135 2.96 ;
      RECT 40.08 2.647 40.09 2.96 ;
      RECT 40.065 2.57 40.08 2.96 ;
      RECT 39.88 2.565 39.965 2.925 ;
      RECT 39.875 2.567 39.88 2.92 ;
      RECT 39.87 2.572 39.875 2.92 ;
      RECT 39.835 2.672 39.87 2.92 ;
      RECT 39.825 2.7 39.835 2.92 ;
      RECT 39.815 2.715 39.825 2.92 ;
      RECT 39.805 2.727 39.815 2.92 ;
      RECT 39.8 2.737 39.805 2.92 ;
      RECT 39.785 2.747 39.8 2.922 ;
      RECT 39.78 2.762 39.785 2.924 ;
      RECT 39.765 2.775 39.78 2.926 ;
      RECT 39.76 2.79 39.765 2.929 ;
      RECT 39.74 2.8 39.76 2.933 ;
      RECT 39.725 2.81 39.74 2.936 ;
      RECT 39.69 2.817 39.725 2.941 ;
      RECT 39.646 2.824 39.69 2.949 ;
      RECT 39.56 2.836 39.646 2.962 ;
      RECT 39.535 2.847 39.56 2.973 ;
      RECT 39.505 2.852 39.535 2.978 ;
      RECT 39.47 2.857 39.505 2.986 ;
      RECT 39.44 2.862 39.47 2.993 ;
      RECT 39.415 2.867 39.44 2.998 ;
      RECT 39.35 2.874 39.415 3.007 ;
      RECT 39.28 2.887 39.35 3.023 ;
      RECT 39.25 2.897 39.28 3.035 ;
      RECT 39.225 2.902 39.25 3.042 ;
      RECT 39.17 2.909 39.225 3.05 ;
      RECT 39.165 2.916 39.17 3.055 ;
      RECT 39.16 2.918 39.165 3.056 ;
      RECT 39.145 2.92 39.16 3.058 ;
      RECT 39.14 2.92 39.145 3.061 ;
      RECT 39.075 2.927 39.14 3.068 ;
      RECT 39.04 2.937 39.07 3.078 ;
      RECT 39.023 2.94 39.04 3.08 ;
      RECT 38.937 2.939 39.023 3.079 ;
      RECT 38.851 2.937 38.937 3.076 ;
      RECT 38.765 2.936 38.851 3.074 ;
      RECT 38.664 2.934 38.73 3.073 ;
      RECT 38.578 2.931 38.664 3.071 ;
      RECT 38.492 2.927 38.578 3.069 ;
      RECT 38.406 2.924 38.492 3.068 ;
      RECT 38.32 2.921 38.406 3.066 ;
      RECT 38.22 2.92 38.305 3.063 ;
      RECT 38.17 2.918 38.22 3.061 ;
      RECT 38.15 2.915 38.17 3.059 ;
      RECT 38.13 2.913 38.15 3.056 ;
      RECT 38.105 2.909 38.13 3.053 ;
      RECT 38.06 2.903 38.105 3.048 ;
      RECT 38.02 2.897 38.06 3.04 ;
      RECT 37.995 2.892 38.02 3.033 ;
      RECT 37.94 2.885 37.995 3.025 ;
      RECT 37.916 2.878 37.94 3.018 ;
      RECT 37.83 2.869 37.916 3.008 ;
      RECT 37.8 2.861 37.83 2.998 ;
      RECT 37.77 2.857 37.8 2.993 ;
      RECT 37.765 2.854 37.77 2.99 ;
      RECT 37.76 2.853 37.765 2.99 ;
      RECT 37.685 2.846 37.76 2.983 ;
      RECT 37.646 2.837 37.685 2.972 ;
      RECT 37.56 2.827 37.646 2.96 ;
      RECT 37.52 2.817 37.56 2.948 ;
      RECT 37.481 2.812 37.52 2.941 ;
      RECT 37.395 2.802 37.481 2.93 ;
      RECT 37.355 2.79 37.395 2.919 ;
      RECT 37.32 2.775 37.355 2.912 ;
      RECT 37.31 2.765 37.32 2.909 ;
      RECT 37.29 2.75 37.31 2.907 ;
      RECT 37.26 2.72 37.29 2.903 ;
      RECT 37.25 2.7 37.26 2.898 ;
      RECT 37.245 2.692 37.25 2.895 ;
      RECT 37.24 2.685 37.245 2.893 ;
      RECT 37.225 2.672 37.24 2.886 ;
      RECT 37.22 2.662 37.225 2.878 ;
      RECT 37.215 2.655 37.22 2.873 ;
      RECT 37.21 2.65 37.215 2.869 ;
      RECT 37.195 2.637 37.21 2.861 ;
      RECT 37.19 2.547 37.195 2.85 ;
      RECT 37.185 2.542 37.19 2.843 ;
      RECT 37.11 2.54 37.185 2.803 ;
      RECT 37.08 2.54 37.11 2.758 ;
      RECT 36.985 2.545 37 2.745 ;
      RECT 39.47 2.25 39.73 2.51 ;
      RECT 39.455 2.238 39.635 2.475 ;
      RECT 39.45 2.239 39.635 2.473 ;
      RECT 39.435 2.243 39.645 2.463 ;
      RECT 39.43 2.248 39.65 2.433 ;
      RECT 39.435 2.245 39.65 2.463 ;
      RECT 39.45 2.24 39.645 2.473 ;
      RECT 39.47 2.237 39.635 2.51 ;
      RECT 39.47 2.236 39.625 2.51 ;
      RECT 39.495 2.235 39.625 2.51 ;
      RECT 39.055 2.48 39.315 2.74 ;
      RECT 38.93 2.525 39.315 2.735 ;
      RECT 38.92 2.53 39.315 2.73 ;
      RECT 38.935 3.47 38.95 3.78 ;
      RECT 37.53 3.24 37.54 3.37 ;
      RECT 37.31 3.235 37.415 3.37 ;
      RECT 37.225 3.24 37.275 3.37 ;
      RECT 35.775 1.975 35.78 3.08 ;
      RECT 39.03 3.562 39.035 3.698 ;
      RECT 39.025 3.557 39.03 3.758 ;
      RECT 39.02 3.555 39.025 3.771 ;
      RECT 39.005 3.552 39.02 3.773 ;
      RECT 39 3.547 39.005 3.775 ;
      RECT 38.995 3.543 39 3.778 ;
      RECT 38.98 3.538 38.995 3.78 ;
      RECT 38.95 3.53 38.98 3.78 ;
      RECT 38.911 3.47 38.935 3.78 ;
      RECT 38.825 3.47 38.911 3.777 ;
      RECT 38.795 3.47 38.825 3.77 ;
      RECT 38.77 3.47 38.795 3.763 ;
      RECT 38.745 3.47 38.77 3.755 ;
      RECT 38.73 3.47 38.745 3.748 ;
      RECT 38.705 3.47 38.73 3.74 ;
      RECT 38.69 3.47 38.705 3.733 ;
      RECT 38.65 3.48 38.69 3.722 ;
      RECT 38.64 3.475 38.65 3.712 ;
      RECT 38.636 3.474 38.64 3.709 ;
      RECT 38.55 3.466 38.636 3.692 ;
      RECT 38.517 3.455 38.55 3.669 ;
      RECT 38.431 3.444 38.517 3.647 ;
      RECT 38.345 3.428 38.431 3.616 ;
      RECT 38.275 3.413 38.345 3.588 ;
      RECT 38.265 3.406 38.275 3.575 ;
      RECT 38.235 3.403 38.265 3.565 ;
      RECT 38.21 3.399 38.235 3.558 ;
      RECT 38.195 3.396 38.21 3.553 ;
      RECT 38.19 3.395 38.195 3.548 ;
      RECT 38.16 3.39 38.19 3.541 ;
      RECT 38.155 3.385 38.16 3.536 ;
      RECT 38.14 3.382 38.155 3.531 ;
      RECT 38.135 3.377 38.14 3.526 ;
      RECT 38.115 3.372 38.135 3.523 ;
      RECT 38.1 3.367 38.115 3.515 ;
      RECT 38.085 3.361 38.1 3.51 ;
      RECT 38.055 3.352 38.085 3.503 ;
      RECT 38.05 3.345 38.055 3.495 ;
      RECT 38.045 3.343 38.05 3.493 ;
      RECT 38.04 3.342 38.045 3.49 ;
      RECT 38 3.335 38.04 3.483 ;
      RECT 37.986 3.325 38 3.473 ;
      RECT 37.935 3.314 37.986 3.461 ;
      RECT 37.91 3.3 37.935 3.447 ;
      RECT 37.885 3.289 37.91 3.439 ;
      RECT 37.865 3.278 37.885 3.433 ;
      RECT 37.855 3.272 37.865 3.428 ;
      RECT 37.85 3.27 37.855 3.424 ;
      RECT 37.83 3.265 37.85 3.419 ;
      RECT 37.8 3.255 37.83 3.409 ;
      RECT 37.795 3.247 37.8 3.402 ;
      RECT 37.78 3.245 37.795 3.398 ;
      RECT 37.76 3.245 37.78 3.393 ;
      RECT 37.755 3.244 37.76 3.391 ;
      RECT 37.75 3.244 37.755 3.388 ;
      RECT 37.71 3.243 37.75 3.383 ;
      RECT 37.685 3.242 37.71 3.378 ;
      RECT 37.625 3.241 37.685 3.375 ;
      RECT 37.54 3.24 37.625 3.373 ;
      RECT 37.501 3.239 37.53 3.37 ;
      RECT 37.415 3.237 37.501 3.37 ;
      RECT 37.275 3.237 37.31 3.37 ;
      RECT 37.185 3.241 37.225 3.373 ;
      RECT 37.17 3.244 37.185 3.38 ;
      RECT 37.16 3.245 37.17 3.387 ;
      RECT 37.135 3.248 37.16 3.392 ;
      RECT 37.13 3.25 37.135 3.395 ;
      RECT 37.08 3.252 37.13 3.396 ;
      RECT 37.041 3.256 37.08 3.398 ;
      RECT 36.955 3.258 37.041 3.401 ;
      RECT 36.937 3.26 36.955 3.403 ;
      RECT 36.851 3.263 36.937 3.405 ;
      RECT 36.765 3.267 36.851 3.408 ;
      RECT 36.728 3.271 36.765 3.411 ;
      RECT 36.642 3.274 36.728 3.414 ;
      RECT 36.556 3.278 36.642 3.417 ;
      RECT 36.47 3.283 36.556 3.421 ;
      RECT 36.45 3.285 36.47 3.424 ;
      RECT 36.43 3.284 36.45 3.425 ;
      RECT 36.381 3.281 36.43 3.426 ;
      RECT 36.295 3.276 36.381 3.429 ;
      RECT 36.245 3.271 36.295 3.431 ;
      RECT 36.221 3.269 36.245 3.432 ;
      RECT 36.135 3.264 36.221 3.434 ;
      RECT 36.11 3.26 36.135 3.433 ;
      RECT 36.1 3.257 36.11 3.431 ;
      RECT 36.09 3.25 36.1 3.428 ;
      RECT 36.085 3.23 36.09 3.423 ;
      RECT 36.075 3.2 36.085 3.418 ;
      RECT 36.06 3.07 36.075 3.409 ;
      RECT 36.055 3.062 36.06 3.402 ;
      RECT 36.035 3.055 36.055 3.394 ;
      RECT 36.03 3.037 36.035 3.386 ;
      RECT 36.02 3.017 36.03 3.381 ;
      RECT 36.015 2.99 36.02 3.377 ;
      RECT 36.01 2.967 36.015 3.374 ;
      RECT 35.99 2.925 36.01 3.366 ;
      RECT 35.955 2.84 35.99 3.35 ;
      RECT 35.95 2.772 35.955 3.338 ;
      RECT 35.935 2.742 35.95 3.332 ;
      RECT 35.93 1.987 35.935 2.233 ;
      RECT 35.92 2.712 35.935 3.323 ;
      RECT 35.925 1.982 35.93 2.265 ;
      RECT 35.92 1.977 35.925 2.308 ;
      RECT 35.915 1.975 35.92 2.343 ;
      RECT 35.9 2.675 35.92 3.313 ;
      RECT 35.91 1.975 35.915 2.38 ;
      RECT 35.895 1.975 35.91 2.478 ;
      RECT 35.895 2.648 35.9 3.306 ;
      RECT 35.89 1.975 35.895 2.553 ;
      RECT 35.89 2.636 35.895 3.303 ;
      RECT 35.885 1.975 35.89 2.585 ;
      RECT 35.885 2.615 35.89 3.3 ;
      RECT 35.88 1.975 35.885 3.297 ;
      RECT 35.845 1.975 35.88 3.283 ;
      RECT 35.83 1.975 35.845 3.265 ;
      RECT 35.81 1.975 35.83 3.255 ;
      RECT 35.785 1.975 35.81 3.238 ;
      RECT 35.78 1.975 35.785 3.188 ;
      RECT 35.77 1.975 35.775 3.018 ;
      RECT 35.765 1.975 35.77 2.925 ;
      RECT 35.76 1.975 35.765 2.838 ;
      RECT 35.755 1.975 35.76 2.77 ;
      RECT 35.75 1.975 35.755 2.713 ;
      RECT 35.74 1.975 35.75 2.608 ;
      RECT 35.735 1.975 35.74 2.48 ;
      RECT 35.73 1.975 35.735 2.398 ;
      RECT 35.725 1.977 35.73 2.315 ;
      RECT 35.72 1.982 35.725 2.248 ;
      RECT 35.715 1.987 35.72 2.175 ;
      RECT 38.53 2.305 38.79 2.565 ;
      RECT 38.55 2.272 38.76 2.565 ;
      RECT 38.55 2.27 38.75 2.565 ;
      RECT 38.56 2.257 38.75 2.565 ;
      RECT 38.56 2.255 38.675 2.565 ;
      RECT 38.035 2.38 38.21 2.66 ;
      RECT 38.03 2.38 38.21 2.658 ;
      RECT 38.03 2.38 38.225 2.655 ;
      RECT 38.02 2.38 38.225 2.653 ;
      RECT 37.965 2.38 38.225 2.64 ;
      RECT 37.965 2.455 38.23 2.618 ;
      RECT 37.51 2.392 37.53 2.635 ;
      RECT 37.51 2.392 37.57 2.634 ;
      RECT 37.505 2.394 37.57 2.633 ;
      RECT 37.505 2.394 37.656 2.632 ;
      RECT 37.505 2.394 37.725 2.631 ;
      RECT 37.505 2.394 37.745 2.623 ;
      RECT 37.485 2.397 37.745 2.621 ;
      RECT 37.47 2.407 37.745 2.606 ;
      RECT 37.47 2.407 37.76 2.605 ;
      RECT 37.465 2.416 37.76 2.597 ;
      RECT 37.465 2.416 37.765 2.593 ;
      RECT 37.57 2.33 37.83 2.59 ;
      RECT 37.46 2.418 37.83 2.475 ;
      RECT 37.53 2.385 37.83 2.59 ;
      RECT 37.495 3.578 37.5 3.785 ;
      RECT 37.445 3.572 37.495 3.784 ;
      RECT 37.412 3.586 37.505 3.783 ;
      RECT 37.326 3.586 37.505 3.782 ;
      RECT 37.24 3.586 37.505 3.781 ;
      RECT 37.24 3.685 37.51 3.778 ;
      RECT 37.235 3.685 37.51 3.773 ;
      RECT 37.23 3.685 37.51 3.755 ;
      RECT 37.225 3.685 37.51 3.738 ;
      RECT 37.185 3.47 37.445 3.73 ;
      RECT 36.645 2.62 36.731 3.034 ;
      RECT 36.645 2.62 36.77 3.031 ;
      RECT 36.645 2.62 36.79 3.021 ;
      RECT 36.6 2.62 36.79 3.018 ;
      RECT 36.6 2.772 36.8 3.008 ;
      RECT 36.6 2.793 36.805 3.002 ;
      RECT 36.6 2.811 36.81 2.998 ;
      RECT 36.6 2.831 36.82 2.993 ;
      RECT 36.575 2.831 36.82 2.99 ;
      RECT 36.565 2.831 36.82 2.968 ;
      RECT 36.565 2.847 36.825 2.938 ;
      RECT 36.53 2.62 36.79 2.925 ;
      RECT 36.53 2.859 36.83 2.88 ;
      RECT 34.19 7.77 34.48 8 ;
      RECT 34.25 6.29 34.42 8 ;
      RECT 34.24 6.66 34.595 7.015 ;
      RECT 34.19 6.29 34.48 6.52 ;
      RECT 33.785 2.395 33.89 2.965 ;
      RECT 33.785 2.73 34.11 2.96 ;
      RECT 33.785 2.76 34.28 2.93 ;
      RECT 33.785 2.395 33.975 2.96 ;
      RECT 33.2 2.36 33.49 2.59 ;
      RECT 33.2 2.395 33.975 2.565 ;
      RECT 33.26 0.88 33.43 2.59 ;
      RECT 33.2 0.88 33.49 1.11 ;
      RECT 33.2 7.77 33.49 8 ;
      RECT 33.26 6.29 33.43 8 ;
      RECT 33.2 6.29 33.49 6.52 ;
      RECT 33.2 6.325 34.055 6.485 ;
      RECT 33.885 5.92 34.055 6.485 ;
      RECT 33.2 6.32 33.595 6.485 ;
      RECT 33.82 5.92 34.11 6.15 ;
      RECT 33.82 5.95 34.28 6.12 ;
      RECT 32.83 2.73 33.12 2.96 ;
      RECT 32.83 2.76 33.29 2.93 ;
      RECT 32.895 1.655 33.06 2.96 ;
      RECT 31.41 1.625 31.7 1.855 ;
      RECT 31.41 1.655 33.06 1.825 ;
      RECT 31.47 0.885 31.64 1.855 ;
      RECT 31.41 0.885 31.7 1.115 ;
      RECT 31.41 7.765 31.7 7.995 ;
      RECT 31.47 7.025 31.64 7.995 ;
      RECT 31.47 7.12 33.06 7.29 ;
      RECT 32.89 5.92 33.06 7.29 ;
      RECT 31.41 7.025 31.7 7.255 ;
      RECT 32.83 5.92 33.12 6.15 ;
      RECT 32.83 5.95 33.29 6.12 ;
      RECT 29.46 2.705 29.8 3.055 ;
      RECT 29.55 2.025 29.72 3.055 ;
      RECT 31.84 1.965 32.19 2.315 ;
      RECT 29.55 2.025 32.19 2.195 ;
      RECT 31.865 6.655 32.19 6.98 ;
      RECT 26.405 6.61 26.755 6.96 ;
      RECT 31.84 6.655 32.19 6.885 ;
      RECT 26.205 6.655 26.755 6.885 ;
      RECT 26.035 6.685 32.19 6.855 ;
      RECT 31.065 2.365 31.385 2.685 ;
      RECT 31.035 2.365 31.385 2.595 ;
      RECT 30.865 2.395 31.385 2.565 ;
      RECT 31.065 6.255 31.385 6.545 ;
      RECT 31.035 6.285 31.385 6.515 ;
      RECT 30.865 6.315 31.385 6.485 ;
      RECT 26.755 2.985 26.905 3.26 ;
      RECT 27.295 2.065 27.3 2.285 ;
      RECT 28.445 2.265 28.46 2.463 ;
      RECT 28.41 2.257 28.445 2.47 ;
      RECT 28.38 2.25 28.41 2.47 ;
      RECT 28.325 2.215 28.38 2.47 ;
      RECT 28.26 2.152 28.325 2.47 ;
      RECT 28.255 2.117 28.26 2.468 ;
      RECT 28.25 2.112 28.255 2.46 ;
      RECT 28.245 2.107 28.25 2.446 ;
      RECT 28.24 2.104 28.245 2.439 ;
      RECT 28.195 2.094 28.24 2.39 ;
      RECT 28.175 2.081 28.195 2.325 ;
      RECT 28.17 2.076 28.175 2.298 ;
      RECT 28.165 2.075 28.17 2.291 ;
      RECT 28.16 2.074 28.165 2.284 ;
      RECT 28.075 2.059 28.16 2.23 ;
      RECT 28.045 2.04 28.075 2.18 ;
      RECT 27.965 2.023 28.045 2.165 ;
      RECT 27.93 2.01 27.965 2.15 ;
      RECT 27.922 2.01 27.93 2.145 ;
      RECT 27.836 2.011 27.922 2.145 ;
      RECT 27.75 2.013 27.836 2.145 ;
      RECT 27.725 2.014 27.75 2.149 ;
      RECT 27.65 2.02 27.725 2.164 ;
      RECT 27.567 2.032 27.65 2.188 ;
      RECT 27.481 2.045 27.567 2.214 ;
      RECT 27.395 2.058 27.481 2.24 ;
      RECT 27.36 2.067 27.395 2.259 ;
      RECT 27.31 2.067 27.36 2.272 ;
      RECT 27.3 2.065 27.31 2.283 ;
      RECT 27.285 2.062 27.295 2.285 ;
      RECT 27.27 2.054 27.285 2.293 ;
      RECT 27.255 2.046 27.27 2.313 ;
      RECT 27.25 2.041 27.255 2.37 ;
      RECT 27.235 2.036 27.25 2.443 ;
      RECT 27.23 2.031 27.235 2.485 ;
      RECT 27.225 2.029 27.23 2.513 ;
      RECT 27.22 2.027 27.225 2.535 ;
      RECT 27.21 2.023 27.22 2.578 ;
      RECT 27.205 2.02 27.21 2.603 ;
      RECT 27.2 2.018 27.205 2.623 ;
      RECT 27.195 2.016 27.2 2.647 ;
      RECT 27.19 2.012 27.195 2.67 ;
      RECT 27.185 2.008 27.19 2.693 ;
      RECT 27.15 1.998 27.185 2.8 ;
      RECT 27.145 1.988 27.15 2.898 ;
      RECT 27.14 1.986 27.145 2.925 ;
      RECT 27.135 1.985 27.14 2.945 ;
      RECT 27.13 1.977 27.135 2.965 ;
      RECT 27.125 1.972 27.13 3 ;
      RECT 27.12 1.97 27.125 3.018 ;
      RECT 27.115 1.97 27.12 3.043 ;
      RECT 27.11 1.97 27.115 3.065 ;
      RECT 27.075 1.97 27.11 3.108 ;
      RECT 27.05 1.97 27.075 3.137 ;
      RECT 27.04 1.97 27.05 2.323 ;
      RECT 27.043 2.38 27.05 3.147 ;
      RECT 27.04 2.437 27.043 3.15 ;
      RECT 27.035 1.97 27.04 2.295 ;
      RECT 27.035 2.487 27.04 3.153 ;
      RECT 27.025 1.97 27.035 2.285 ;
      RECT 27.03 2.54 27.035 3.156 ;
      RECT 27.025 2.625 27.03 3.16 ;
      RECT 27.015 1.97 27.025 2.273 ;
      RECT 27.02 2.672 27.025 3.164 ;
      RECT 27.015 2.747 27.02 3.168 ;
      RECT 26.98 1.97 27.015 2.248 ;
      RECT 27.005 2.83 27.015 3.173 ;
      RECT 26.995 2.897 27.005 3.18 ;
      RECT 26.99 2.925 26.995 3.185 ;
      RECT 26.98 2.938 26.99 3.191 ;
      RECT 26.935 1.97 26.98 2.205 ;
      RECT 26.975 2.943 26.98 3.198 ;
      RECT 26.935 2.96 26.975 3.26 ;
      RECT 26.93 1.972 26.935 2.178 ;
      RECT 26.905 2.98 26.935 3.26 ;
      RECT 26.925 1.977 26.93 2.15 ;
      RECT 26.715 2.989 26.755 3.26 ;
      RECT 26.69 2.997 26.715 3.23 ;
      RECT 26.645 3.005 26.69 3.23 ;
      RECT 26.63 3.01 26.645 3.225 ;
      RECT 26.62 3.01 26.63 3.219 ;
      RECT 26.61 3.017 26.62 3.216 ;
      RECT 26.605 3.055 26.61 3.205 ;
      RECT 26.6 3.117 26.605 3.183 ;
      RECT 27.87 2.992 28.055 3.215 ;
      RECT 27.87 3.007 28.06 3.211 ;
      RECT 27.86 2.28 27.945 3.21 ;
      RECT 27.86 3.007 28.065 3.204 ;
      RECT 27.855 3.015 28.065 3.203 ;
      RECT 28.06 2.735 28.38 3.055 ;
      RECT 27.855 2.907 28.025 2.998 ;
      RECT 27.85 2.907 28.025 2.98 ;
      RECT 27.84 2.715 27.975 2.955 ;
      RECT 27.835 2.715 27.975 2.9 ;
      RECT 27.795 2.295 27.965 2.8 ;
      RECT 27.78 2.295 27.965 2.67 ;
      RECT 27.775 2.295 27.965 2.623 ;
      RECT 27.77 2.295 27.965 2.603 ;
      RECT 27.765 2.295 27.965 2.578 ;
      RECT 27.735 2.295 27.995 2.555 ;
      RECT 27.745 2.292 27.955 2.555 ;
      RECT 27.87 2.287 27.955 3.215 ;
      RECT 27.755 2.28 27.945 2.555 ;
      RECT 27.75 2.285 27.945 2.555 ;
      RECT 26.58 2.497 26.765 2.71 ;
      RECT 26.58 2.505 26.775 2.703 ;
      RECT 26.56 2.505 26.775 2.7 ;
      RECT 26.555 2.505 26.775 2.685 ;
      RECT 26.485 2.42 26.745 2.68 ;
      RECT 26.485 2.565 26.78 2.593 ;
      RECT 26.14 3.02 26.4 3.28 ;
      RECT 26.165 2.965 26.36 3.28 ;
      RECT 26.16 2.714 26.34 3.008 ;
      RECT 26.16 2.72 26.35 3.008 ;
      RECT 26.14 2.722 26.35 2.953 ;
      RECT 26.135 2.732 26.35 2.82 ;
      RECT 26.165 2.712 26.34 3.28 ;
      RECT 26.251 2.71 26.34 3.28 ;
      RECT 26.11 1.93 26.145 2.3 ;
      RECT 25.9 2.04 25.905 2.3 ;
      RECT 26.145 1.937 26.16 2.3 ;
      RECT 26.035 1.93 26.11 2.378 ;
      RECT 26.025 1.93 26.035 2.463 ;
      RECT 26 1.93 26.025 2.498 ;
      RECT 25.96 1.93 26 2.566 ;
      RECT 25.95 1.937 25.96 2.618 ;
      RECT 25.92 2.04 25.95 2.659 ;
      RECT 25.915 2.04 25.92 2.698 ;
      RECT 25.905 2.04 25.915 2.718 ;
      RECT 25.9 2.335 25.905 2.755 ;
      RECT 25.895 2.352 25.9 2.775 ;
      RECT 25.88 2.415 25.895 2.815 ;
      RECT 25.875 2.458 25.88 2.85 ;
      RECT 25.87 2.466 25.875 2.863 ;
      RECT 25.86 2.48 25.87 2.885 ;
      RECT 25.835 2.515 25.86 2.95 ;
      RECT 25.825 2.55 25.835 3.013 ;
      RECT 25.805 2.58 25.825 3.074 ;
      RECT 25.79 2.616 25.805 3.141 ;
      RECT 25.78 2.644 25.79 3.18 ;
      RECT 25.77 2.666 25.78 3.2 ;
      RECT 25.765 2.676 25.77 3.211 ;
      RECT 25.76 2.685 25.765 3.214 ;
      RECT 25.75 2.703 25.76 3.218 ;
      RECT 25.74 2.721 25.75 3.219 ;
      RECT 25.715 2.76 25.74 3.216 ;
      RECT 25.695 2.802 25.715 3.213 ;
      RECT 25.68 2.84 25.695 3.212 ;
      RECT 25.645 2.875 25.68 3.209 ;
      RECT 25.64 2.897 25.645 3.207 ;
      RECT 25.575 2.937 25.64 3.204 ;
      RECT 25.57 2.977 25.575 3.2 ;
      RECT 25.555 2.987 25.57 3.191 ;
      RECT 25.545 3.107 25.555 3.176 ;
      RECT 26.025 3.52 26.035 3.78 ;
      RECT 26.025 3.523 26.045 3.779 ;
      RECT 26.015 3.513 26.025 3.778 ;
      RECT 26.005 3.528 26.085 3.774 ;
      RECT 25.99 3.507 26.005 3.772 ;
      RECT 25.965 3.532 26.09 3.768 ;
      RECT 25.95 3.492 25.965 3.763 ;
      RECT 25.95 3.534 26.1 3.762 ;
      RECT 25.95 3.542 26.115 3.755 ;
      RECT 25.89 3.479 25.95 3.745 ;
      RECT 25.88 3.466 25.89 3.727 ;
      RECT 25.855 3.456 25.88 3.717 ;
      RECT 25.85 3.446 25.855 3.709 ;
      RECT 25.785 3.542 26.115 3.691 ;
      RECT 25.7 3.542 26.115 3.653 ;
      RECT 25.59 3.37 25.85 3.63 ;
      RECT 25.965 3.5 25.99 3.768 ;
      RECT 26.005 3.51 26.015 3.774 ;
      RECT 25.59 3.518 26.03 3.63 ;
      RECT 25.775 7.765 26.065 7.995 ;
      RECT 25.835 7.025 26.005 7.995 ;
      RECT 25.735 7.055 26.105 7.425 ;
      RECT 25.775 7.025 26.065 7.425 ;
      RECT 24.805 3.275 24.835 3.575 ;
      RECT 24.58 3.26 24.585 3.535 ;
      RECT 24.38 3.26 24.535 3.52 ;
      RECT 25.68 1.975 25.71 2.235 ;
      RECT 25.67 1.975 25.68 2.343 ;
      RECT 25.65 1.975 25.67 2.353 ;
      RECT 25.635 1.975 25.65 2.365 ;
      RECT 25.58 1.975 25.635 2.415 ;
      RECT 25.565 1.975 25.58 2.463 ;
      RECT 25.535 1.975 25.565 2.498 ;
      RECT 25.48 1.975 25.535 2.56 ;
      RECT 25.46 1.975 25.48 2.628 ;
      RECT 25.455 1.975 25.46 2.658 ;
      RECT 25.45 1.975 25.455 2.67 ;
      RECT 25.445 2.092 25.45 2.688 ;
      RECT 25.425 2.11 25.445 2.713 ;
      RECT 25.405 2.137 25.425 2.763 ;
      RECT 25.4 2.157 25.405 2.794 ;
      RECT 25.395 2.165 25.4 2.811 ;
      RECT 25.38 2.191 25.395 2.84 ;
      RECT 25.365 2.233 25.38 2.875 ;
      RECT 25.36 2.262 25.365 2.898 ;
      RECT 25.355 2.277 25.36 2.911 ;
      RECT 25.35 2.3 25.355 2.922 ;
      RECT 25.34 2.32 25.35 2.94 ;
      RECT 25.33 2.35 25.34 2.963 ;
      RECT 25.325 2.372 25.33 2.983 ;
      RECT 25.32 2.387 25.325 2.998 ;
      RECT 25.305 2.417 25.32 3.025 ;
      RECT 25.3 2.447 25.305 3.051 ;
      RECT 25.295 2.465 25.3 3.063 ;
      RECT 25.285 2.495 25.295 3.082 ;
      RECT 25.275 2.52 25.285 3.107 ;
      RECT 25.27 2.54 25.275 3.126 ;
      RECT 25.265 2.557 25.27 3.139 ;
      RECT 25.255 2.583 25.265 3.158 ;
      RECT 25.245 2.621 25.255 3.185 ;
      RECT 25.24 2.647 25.245 3.205 ;
      RECT 25.235 2.657 25.24 3.215 ;
      RECT 25.23 2.67 25.235 3.23 ;
      RECT 25.225 2.685 25.23 3.24 ;
      RECT 25.22 2.707 25.225 3.255 ;
      RECT 25.215 2.725 25.22 3.266 ;
      RECT 25.21 2.735 25.215 3.277 ;
      RECT 25.205 2.743 25.21 3.289 ;
      RECT 25.2 2.751 25.205 3.3 ;
      RECT 25.195 2.777 25.2 3.313 ;
      RECT 25.185 2.805 25.195 3.326 ;
      RECT 25.18 2.835 25.185 3.335 ;
      RECT 25.175 2.85 25.18 3.342 ;
      RECT 25.16 2.875 25.175 3.349 ;
      RECT 25.155 2.897 25.16 3.355 ;
      RECT 25.15 2.922 25.155 3.358 ;
      RECT 25.141 2.95 25.15 3.362 ;
      RECT 25.135 2.967 25.141 3.367 ;
      RECT 25.13 2.985 25.135 3.371 ;
      RECT 25.125 2.997 25.13 3.374 ;
      RECT 25.12 3.018 25.125 3.378 ;
      RECT 25.115 3.036 25.12 3.381 ;
      RECT 25.11 3.05 25.115 3.384 ;
      RECT 25.105 3.067 25.11 3.387 ;
      RECT 25.1 3.08 25.105 3.39 ;
      RECT 25.075 3.117 25.1 3.398 ;
      RECT 25.07 3.162 25.075 3.407 ;
      RECT 25.065 3.19 25.07 3.41 ;
      RECT 25.055 3.21 25.065 3.414 ;
      RECT 25.05 3.23 25.055 3.419 ;
      RECT 25.045 3.245 25.05 3.422 ;
      RECT 25.025 3.255 25.045 3.429 ;
      RECT 24.96 3.262 25.025 3.455 ;
      RECT 24.925 3.265 24.96 3.483 ;
      RECT 24.91 3.268 24.925 3.498 ;
      RECT 24.9 3.269 24.91 3.513 ;
      RECT 24.89 3.27 24.9 3.53 ;
      RECT 24.885 3.27 24.89 3.545 ;
      RECT 24.88 3.27 24.885 3.553 ;
      RECT 24.865 3.271 24.88 3.568 ;
      RECT 24.835 3.273 24.865 3.575 ;
      RECT 24.725 3.28 24.805 3.575 ;
      RECT 24.68 3.285 24.725 3.575 ;
      RECT 24.67 3.286 24.68 3.565 ;
      RECT 24.66 3.287 24.67 3.558 ;
      RECT 24.64 3.289 24.66 3.553 ;
      RECT 24.63 3.26 24.64 3.548 ;
      RECT 24.585 3.26 24.63 3.54 ;
      RECT 24.555 3.26 24.58 3.53 ;
      RECT 24.535 3.26 24.555 3.523 ;
      RECT 24.815 2.06 25.075 2.32 ;
      RECT 24.695 2.075 24.705 2.24 ;
      RECT 24.68 2.075 24.685 2.235 ;
      RECT 22.045 1.915 22.23 2.205 ;
      RECT 23.86 2.04 23.875 2.195 ;
      RECT 22.01 1.915 22.035 2.175 ;
      RECT 24.425 1.965 24.43 2.107 ;
      RECT 24.34 1.96 24.365 2.1 ;
      RECT 24.74 2.077 24.815 2.27 ;
      RECT 24.725 2.075 24.74 2.253 ;
      RECT 24.705 2.075 24.725 2.245 ;
      RECT 24.685 2.075 24.695 2.238 ;
      RECT 24.64 2.07 24.68 2.228 ;
      RECT 24.6 2.045 24.64 2.213 ;
      RECT 24.585 2.02 24.6 2.203 ;
      RECT 24.58 2.014 24.585 2.201 ;
      RECT 24.545 2.006 24.58 2.184 ;
      RECT 24.54 1.999 24.545 2.172 ;
      RECT 24.52 1.994 24.54 2.16 ;
      RECT 24.51 1.988 24.52 2.145 ;
      RECT 24.49 1.983 24.51 2.13 ;
      RECT 24.48 1.978 24.49 2.123 ;
      RECT 24.475 1.976 24.48 2.118 ;
      RECT 24.47 1.975 24.475 2.115 ;
      RECT 24.43 1.97 24.47 2.111 ;
      RECT 24.41 1.964 24.425 2.106 ;
      RECT 24.375 1.961 24.41 2.103 ;
      RECT 24.365 1.96 24.375 2.101 ;
      RECT 24.305 1.96 24.34 2.098 ;
      RECT 24.26 1.96 24.305 2.098 ;
      RECT 24.21 1.96 24.26 2.101 ;
      RECT 24.195 1.962 24.21 2.103 ;
      RECT 24.18 1.965 24.195 2.104 ;
      RECT 24.17 1.97 24.18 2.105 ;
      RECT 24.14 1.975 24.17 2.11 ;
      RECT 24.13 1.981 24.14 2.118 ;
      RECT 24.12 1.983 24.13 2.122 ;
      RECT 24.11 1.987 24.12 2.126 ;
      RECT 24.085 1.993 24.11 2.134 ;
      RECT 24.075 1.998 24.085 2.142 ;
      RECT 24.06 2.002 24.075 2.146 ;
      RECT 24.025 2.008 24.06 2.154 ;
      RECT 24.005 2.013 24.025 2.164 ;
      RECT 23.975 2.02 24.005 2.173 ;
      RECT 23.93 2.029 23.975 2.187 ;
      RECT 23.925 2.034 23.93 2.198 ;
      RECT 23.905 2.037 23.925 2.199 ;
      RECT 23.875 2.04 23.905 2.197 ;
      RECT 23.84 2.04 23.86 2.193 ;
      RECT 23.77 2.04 23.84 2.184 ;
      RECT 23.755 2.037 23.77 2.176 ;
      RECT 23.715 2.03 23.755 2.171 ;
      RECT 23.69 2.02 23.715 2.164 ;
      RECT 23.685 2.014 23.69 2.161 ;
      RECT 23.645 2.008 23.685 2.158 ;
      RECT 23.63 2.001 23.645 2.153 ;
      RECT 23.61 1.997 23.63 2.148 ;
      RECT 23.595 1.992 23.61 2.144 ;
      RECT 23.58 1.987 23.595 2.142 ;
      RECT 23.565 1.983 23.58 2.141 ;
      RECT 23.55 1.981 23.565 2.137 ;
      RECT 23.54 1.979 23.55 2.132 ;
      RECT 23.525 1.976 23.54 2.128 ;
      RECT 23.515 1.974 23.525 2.123 ;
      RECT 23.495 1.971 23.515 2.119 ;
      RECT 23.45 1.97 23.495 2.117 ;
      RECT 23.39 1.972 23.45 2.118 ;
      RECT 23.37 1.974 23.39 2.12 ;
      RECT 23.34 1.977 23.37 2.121 ;
      RECT 23.29 1.982 23.34 2.123 ;
      RECT 23.285 1.985 23.29 2.125 ;
      RECT 23.275 1.987 23.285 2.128 ;
      RECT 23.27 1.989 23.275 2.131 ;
      RECT 23.22 1.992 23.27 2.138 ;
      RECT 23.2 1.996 23.22 2.15 ;
      RECT 23.19 1.999 23.2 2.156 ;
      RECT 23.18 2 23.19 2.159 ;
      RECT 23.141 2.003 23.18 2.161 ;
      RECT 23.055 2.01 23.141 2.164 ;
      RECT 22.981 2.02 23.055 2.168 ;
      RECT 22.895 2.031 22.981 2.173 ;
      RECT 22.88 2.038 22.895 2.175 ;
      RECT 22.825 2.042 22.88 2.176 ;
      RECT 22.811 2.045 22.825 2.178 ;
      RECT 22.725 2.045 22.811 2.18 ;
      RECT 22.685 2.042 22.725 2.183 ;
      RECT 22.661 2.038 22.685 2.185 ;
      RECT 22.575 2.028 22.661 2.188 ;
      RECT 22.545 2.017 22.575 2.189 ;
      RECT 22.526 2.013 22.545 2.188 ;
      RECT 22.44 2.006 22.526 2.185 ;
      RECT 22.38 1.995 22.44 2.182 ;
      RECT 22.36 1.987 22.38 2.18 ;
      RECT 22.325 1.982 22.36 2.179 ;
      RECT 22.3 1.977 22.325 2.178 ;
      RECT 22.27 1.972 22.3 2.177 ;
      RECT 22.245 1.915 22.27 2.176 ;
      RECT 22.23 1.915 22.245 2.2 ;
      RECT 22.035 1.915 22.045 2.2 ;
      RECT 23.81 2.935 23.815 3.075 ;
      RECT 23.47 2.935 23.505 3.073 ;
      RECT 23.045 2.92 23.06 3.065 ;
      RECT 24.875 2.7 24.965 2.96 ;
      RECT 24.705 2.565 24.805 2.96 ;
      RECT 21.74 2.54 21.82 2.75 ;
      RECT 24.83 2.677 24.875 2.96 ;
      RECT 24.82 2.647 24.83 2.96 ;
      RECT 24.805 2.57 24.82 2.96 ;
      RECT 24.62 2.565 24.705 2.925 ;
      RECT 24.615 2.567 24.62 2.92 ;
      RECT 24.61 2.572 24.615 2.92 ;
      RECT 24.575 2.672 24.61 2.92 ;
      RECT 24.565 2.7 24.575 2.92 ;
      RECT 24.555 2.715 24.565 2.92 ;
      RECT 24.545 2.727 24.555 2.92 ;
      RECT 24.54 2.737 24.545 2.92 ;
      RECT 24.525 2.747 24.54 2.922 ;
      RECT 24.52 2.762 24.525 2.924 ;
      RECT 24.505 2.775 24.52 2.926 ;
      RECT 24.5 2.79 24.505 2.929 ;
      RECT 24.48 2.8 24.5 2.933 ;
      RECT 24.465 2.81 24.48 2.936 ;
      RECT 24.43 2.817 24.465 2.941 ;
      RECT 24.386 2.824 24.43 2.949 ;
      RECT 24.3 2.836 24.386 2.962 ;
      RECT 24.275 2.847 24.3 2.973 ;
      RECT 24.245 2.852 24.275 2.978 ;
      RECT 24.21 2.857 24.245 2.986 ;
      RECT 24.18 2.862 24.21 2.993 ;
      RECT 24.155 2.867 24.18 2.998 ;
      RECT 24.09 2.874 24.155 3.007 ;
      RECT 24.02 2.887 24.09 3.023 ;
      RECT 23.99 2.897 24.02 3.035 ;
      RECT 23.965 2.902 23.99 3.042 ;
      RECT 23.91 2.909 23.965 3.05 ;
      RECT 23.905 2.916 23.91 3.055 ;
      RECT 23.9 2.918 23.905 3.056 ;
      RECT 23.885 2.92 23.9 3.058 ;
      RECT 23.88 2.92 23.885 3.061 ;
      RECT 23.815 2.927 23.88 3.068 ;
      RECT 23.78 2.937 23.81 3.078 ;
      RECT 23.763 2.94 23.78 3.08 ;
      RECT 23.677 2.939 23.763 3.079 ;
      RECT 23.591 2.937 23.677 3.076 ;
      RECT 23.505 2.936 23.591 3.074 ;
      RECT 23.404 2.934 23.47 3.073 ;
      RECT 23.318 2.931 23.404 3.071 ;
      RECT 23.232 2.927 23.318 3.069 ;
      RECT 23.146 2.924 23.232 3.068 ;
      RECT 23.06 2.921 23.146 3.066 ;
      RECT 22.96 2.92 23.045 3.063 ;
      RECT 22.91 2.918 22.96 3.061 ;
      RECT 22.89 2.915 22.91 3.059 ;
      RECT 22.87 2.913 22.89 3.056 ;
      RECT 22.845 2.909 22.87 3.053 ;
      RECT 22.8 2.903 22.845 3.048 ;
      RECT 22.76 2.897 22.8 3.04 ;
      RECT 22.735 2.892 22.76 3.033 ;
      RECT 22.68 2.885 22.735 3.025 ;
      RECT 22.656 2.878 22.68 3.018 ;
      RECT 22.57 2.869 22.656 3.008 ;
      RECT 22.54 2.861 22.57 2.998 ;
      RECT 22.51 2.857 22.54 2.993 ;
      RECT 22.505 2.854 22.51 2.99 ;
      RECT 22.5 2.853 22.505 2.99 ;
      RECT 22.425 2.846 22.5 2.983 ;
      RECT 22.386 2.837 22.425 2.972 ;
      RECT 22.3 2.827 22.386 2.96 ;
      RECT 22.26 2.817 22.3 2.948 ;
      RECT 22.221 2.812 22.26 2.941 ;
      RECT 22.135 2.802 22.221 2.93 ;
      RECT 22.095 2.79 22.135 2.919 ;
      RECT 22.06 2.775 22.095 2.912 ;
      RECT 22.05 2.765 22.06 2.909 ;
      RECT 22.03 2.75 22.05 2.907 ;
      RECT 22 2.72 22.03 2.903 ;
      RECT 21.99 2.7 22 2.898 ;
      RECT 21.985 2.692 21.99 2.895 ;
      RECT 21.98 2.685 21.985 2.893 ;
      RECT 21.965 2.672 21.98 2.886 ;
      RECT 21.96 2.662 21.965 2.878 ;
      RECT 21.955 2.655 21.96 2.873 ;
      RECT 21.95 2.65 21.955 2.869 ;
      RECT 21.935 2.637 21.95 2.861 ;
      RECT 21.93 2.547 21.935 2.85 ;
      RECT 21.925 2.542 21.93 2.843 ;
      RECT 21.85 2.54 21.925 2.803 ;
      RECT 21.82 2.54 21.85 2.758 ;
      RECT 21.725 2.545 21.74 2.745 ;
      RECT 24.21 2.25 24.47 2.51 ;
      RECT 24.195 2.238 24.375 2.475 ;
      RECT 24.19 2.239 24.375 2.473 ;
      RECT 24.175 2.243 24.385 2.463 ;
      RECT 24.17 2.248 24.39 2.433 ;
      RECT 24.175 2.245 24.39 2.463 ;
      RECT 24.19 2.24 24.385 2.473 ;
      RECT 24.21 2.237 24.375 2.51 ;
      RECT 24.21 2.236 24.365 2.51 ;
      RECT 24.235 2.235 24.365 2.51 ;
      RECT 23.795 2.48 24.055 2.74 ;
      RECT 23.67 2.525 24.055 2.735 ;
      RECT 23.66 2.53 24.055 2.73 ;
      RECT 23.675 3.47 23.69 3.78 ;
      RECT 22.27 3.24 22.28 3.37 ;
      RECT 22.05 3.235 22.155 3.37 ;
      RECT 21.965 3.24 22.015 3.37 ;
      RECT 20.515 1.975 20.52 3.08 ;
      RECT 23.77 3.562 23.775 3.698 ;
      RECT 23.765 3.557 23.77 3.758 ;
      RECT 23.76 3.555 23.765 3.771 ;
      RECT 23.745 3.552 23.76 3.773 ;
      RECT 23.74 3.547 23.745 3.775 ;
      RECT 23.735 3.543 23.74 3.778 ;
      RECT 23.72 3.538 23.735 3.78 ;
      RECT 23.69 3.53 23.72 3.78 ;
      RECT 23.651 3.47 23.675 3.78 ;
      RECT 23.565 3.47 23.651 3.777 ;
      RECT 23.535 3.47 23.565 3.77 ;
      RECT 23.51 3.47 23.535 3.763 ;
      RECT 23.485 3.47 23.51 3.755 ;
      RECT 23.47 3.47 23.485 3.748 ;
      RECT 23.445 3.47 23.47 3.74 ;
      RECT 23.43 3.47 23.445 3.733 ;
      RECT 23.39 3.48 23.43 3.722 ;
      RECT 23.38 3.475 23.39 3.712 ;
      RECT 23.376 3.474 23.38 3.709 ;
      RECT 23.29 3.466 23.376 3.692 ;
      RECT 23.257 3.455 23.29 3.669 ;
      RECT 23.171 3.444 23.257 3.647 ;
      RECT 23.085 3.428 23.171 3.616 ;
      RECT 23.015 3.413 23.085 3.588 ;
      RECT 23.005 3.406 23.015 3.575 ;
      RECT 22.975 3.403 23.005 3.565 ;
      RECT 22.95 3.399 22.975 3.558 ;
      RECT 22.935 3.396 22.95 3.553 ;
      RECT 22.93 3.395 22.935 3.548 ;
      RECT 22.9 3.39 22.93 3.541 ;
      RECT 22.895 3.385 22.9 3.536 ;
      RECT 22.88 3.382 22.895 3.531 ;
      RECT 22.875 3.377 22.88 3.526 ;
      RECT 22.855 3.372 22.875 3.523 ;
      RECT 22.84 3.367 22.855 3.515 ;
      RECT 22.825 3.361 22.84 3.51 ;
      RECT 22.795 3.352 22.825 3.503 ;
      RECT 22.79 3.345 22.795 3.495 ;
      RECT 22.785 3.343 22.79 3.493 ;
      RECT 22.78 3.342 22.785 3.49 ;
      RECT 22.74 3.335 22.78 3.483 ;
      RECT 22.726 3.325 22.74 3.473 ;
      RECT 22.675 3.314 22.726 3.461 ;
      RECT 22.65 3.3 22.675 3.447 ;
      RECT 22.625 3.289 22.65 3.439 ;
      RECT 22.605 3.278 22.625 3.433 ;
      RECT 22.595 3.272 22.605 3.428 ;
      RECT 22.59 3.27 22.595 3.424 ;
      RECT 22.57 3.265 22.59 3.419 ;
      RECT 22.54 3.255 22.57 3.409 ;
      RECT 22.535 3.247 22.54 3.402 ;
      RECT 22.52 3.245 22.535 3.398 ;
      RECT 22.5 3.245 22.52 3.393 ;
      RECT 22.495 3.244 22.5 3.391 ;
      RECT 22.49 3.244 22.495 3.388 ;
      RECT 22.45 3.243 22.49 3.383 ;
      RECT 22.425 3.242 22.45 3.378 ;
      RECT 22.365 3.241 22.425 3.375 ;
      RECT 22.28 3.24 22.365 3.373 ;
      RECT 22.241 3.239 22.27 3.37 ;
      RECT 22.155 3.237 22.241 3.37 ;
      RECT 22.015 3.237 22.05 3.37 ;
      RECT 21.925 3.241 21.965 3.373 ;
      RECT 21.91 3.244 21.925 3.38 ;
      RECT 21.9 3.245 21.91 3.387 ;
      RECT 21.875 3.248 21.9 3.392 ;
      RECT 21.87 3.25 21.875 3.395 ;
      RECT 21.82 3.252 21.87 3.396 ;
      RECT 21.781 3.256 21.82 3.398 ;
      RECT 21.695 3.258 21.781 3.401 ;
      RECT 21.677 3.26 21.695 3.403 ;
      RECT 21.591 3.263 21.677 3.405 ;
      RECT 21.505 3.267 21.591 3.408 ;
      RECT 21.468 3.271 21.505 3.411 ;
      RECT 21.382 3.274 21.468 3.414 ;
      RECT 21.296 3.278 21.382 3.417 ;
      RECT 21.21 3.283 21.296 3.421 ;
      RECT 21.19 3.285 21.21 3.424 ;
      RECT 21.17 3.284 21.19 3.425 ;
      RECT 21.121 3.281 21.17 3.426 ;
      RECT 21.035 3.276 21.121 3.429 ;
      RECT 20.985 3.271 21.035 3.431 ;
      RECT 20.961 3.269 20.985 3.432 ;
      RECT 20.875 3.264 20.961 3.434 ;
      RECT 20.85 3.26 20.875 3.433 ;
      RECT 20.84 3.257 20.85 3.431 ;
      RECT 20.83 3.25 20.84 3.428 ;
      RECT 20.825 3.23 20.83 3.423 ;
      RECT 20.815 3.2 20.825 3.418 ;
      RECT 20.8 3.07 20.815 3.409 ;
      RECT 20.795 3.062 20.8 3.402 ;
      RECT 20.775 3.055 20.795 3.394 ;
      RECT 20.77 3.037 20.775 3.386 ;
      RECT 20.76 3.017 20.77 3.381 ;
      RECT 20.755 2.99 20.76 3.377 ;
      RECT 20.75 2.967 20.755 3.374 ;
      RECT 20.73 2.925 20.75 3.366 ;
      RECT 20.695 2.84 20.73 3.35 ;
      RECT 20.69 2.772 20.695 3.338 ;
      RECT 20.675 2.742 20.69 3.332 ;
      RECT 20.67 1.987 20.675 2.233 ;
      RECT 20.66 2.712 20.675 3.323 ;
      RECT 20.665 1.982 20.67 2.265 ;
      RECT 20.66 1.977 20.665 2.308 ;
      RECT 20.655 1.975 20.66 2.343 ;
      RECT 20.64 2.675 20.66 3.313 ;
      RECT 20.65 1.975 20.655 2.38 ;
      RECT 20.635 1.975 20.65 2.478 ;
      RECT 20.635 2.648 20.64 3.306 ;
      RECT 20.63 1.975 20.635 2.553 ;
      RECT 20.63 2.636 20.635 3.303 ;
      RECT 20.625 1.975 20.63 2.585 ;
      RECT 20.625 2.615 20.63 3.3 ;
      RECT 20.62 1.975 20.625 3.297 ;
      RECT 20.585 1.975 20.62 3.283 ;
      RECT 20.57 1.975 20.585 3.265 ;
      RECT 20.55 1.975 20.57 3.255 ;
      RECT 20.525 1.975 20.55 3.238 ;
      RECT 20.52 1.975 20.525 3.188 ;
      RECT 20.51 1.975 20.515 3.018 ;
      RECT 20.505 1.975 20.51 2.925 ;
      RECT 20.5 1.975 20.505 2.838 ;
      RECT 20.495 1.975 20.5 2.77 ;
      RECT 20.49 1.975 20.495 2.713 ;
      RECT 20.48 1.975 20.49 2.608 ;
      RECT 20.475 1.975 20.48 2.48 ;
      RECT 20.47 1.975 20.475 2.398 ;
      RECT 20.465 1.977 20.47 2.315 ;
      RECT 20.46 1.982 20.465 2.248 ;
      RECT 20.455 1.987 20.46 2.175 ;
      RECT 23.27 2.305 23.53 2.565 ;
      RECT 23.29 2.272 23.5 2.565 ;
      RECT 23.29 2.27 23.49 2.565 ;
      RECT 23.3 2.257 23.49 2.565 ;
      RECT 23.3 2.255 23.415 2.565 ;
      RECT 22.775 2.38 22.95 2.66 ;
      RECT 22.77 2.38 22.95 2.658 ;
      RECT 22.77 2.38 22.965 2.655 ;
      RECT 22.76 2.38 22.965 2.653 ;
      RECT 22.705 2.38 22.965 2.64 ;
      RECT 22.705 2.455 22.97 2.618 ;
      RECT 22.25 2.392 22.27 2.635 ;
      RECT 22.25 2.392 22.31 2.634 ;
      RECT 22.245 2.394 22.31 2.633 ;
      RECT 22.245 2.394 22.396 2.632 ;
      RECT 22.245 2.394 22.465 2.631 ;
      RECT 22.245 2.394 22.485 2.623 ;
      RECT 22.225 2.397 22.485 2.621 ;
      RECT 22.21 2.407 22.485 2.606 ;
      RECT 22.21 2.407 22.5 2.605 ;
      RECT 22.205 2.416 22.5 2.597 ;
      RECT 22.205 2.416 22.505 2.593 ;
      RECT 22.31 2.33 22.57 2.59 ;
      RECT 22.2 2.418 22.57 2.475 ;
      RECT 22.27 2.385 22.57 2.59 ;
      RECT 22.235 3.578 22.24 3.785 ;
      RECT 22.185 3.572 22.235 3.784 ;
      RECT 22.152 3.586 22.245 3.783 ;
      RECT 22.066 3.586 22.245 3.782 ;
      RECT 21.98 3.586 22.245 3.781 ;
      RECT 21.98 3.685 22.25 3.778 ;
      RECT 21.975 3.685 22.25 3.773 ;
      RECT 21.97 3.685 22.25 3.755 ;
      RECT 21.965 3.685 22.25 3.738 ;
      RECT 21.925 3.47 22.185 3.73 ;
      RECT 21.385 2.62 21.471 3.034 ;
      RECT 21.385 2.62 21.51 3.031 ;
      RECT 21.385 2.62 21.53 3.021 ;
      RECT 21.34 2.62 21.53 3.018 ;
      RECT 21.34 2.772 21.54 3.008 ;
      RECT 21.34 2.793 21.545 3.002 ;
      RECT 21.34 2.811 21.55 2.998 ;
      RECT 21.34 2.831 21.56 2.993 ;
      RECT 21.315 2.831 21.56 2.99 ;
      RECT 21.305 2.831 21.56 2.968 ;
      RECT 21.305 2.847 21.565 2.938 ;
      RECT 21.27 2.62 21.53 2.925 ;
      RECT 21.27 2.859 21.57 2.88 ;
      RECT 18.93 7.77 19.22 8 ;
      RECT 18.99 6.29 19.16 8 ;
      RECT 18.985 6.655 19.335 7.005 ;
      RECT 18.93 6.29 19.22 6.52 ;
      RECT 18.525 2.395 18.63 2.965 ;
      RECT 18.525 2.73 18.85 2.96 ;
      RECT 18.525 2.76 19.02 2.93 ;
      RECT 18.525 2.395 18.715 2.96 ;
      RECT 17.94 2.36 18.23 2.59 ;
      RECT 17.94 2.395 18.715 2.565 ;
      RECT 18 0.88 18.17 2.59 ;
      RECT 17.94 0.88 18.23 1.11 ;
      RECT 17.94 7.77 18.23 8 ;
      RECT 18 6.29 18.17 8 ;
      RECT 17.94 6.29 18.23 6.52 ;
      RECT 17.94 6.325 18.795 6.485 ;
      RECT 18.625 5.92 18.795 6.485 ;
      RECT 17.94 6.32 18.335 6.485 ;
      RECT 18.56 5.92 18.85 6.15 ;
      RECT 18.56 5.95 19.02 6.12 ;
      RECT 17.57 2.73 17.86 2.96 ;
      RECT 17.57 2.76 18.03 2.93 ;
      RECT 17.635 1.655 17.8 2.96 ;
      RECT 16.15 1.625 16.44 1.855 ;
      RECT 16.15 1.655 17.8 1.825 ;
      RECT 16.21 0.885 16.38 1.855 ;
      RECT 16.15 0.885 16.44 1.115 ;
      RECT 16.15 7.765 16.44 7.995 ;
      RECT 16.21 7.025 16.38 7.995 ;
      RECT 16.21 7.12 17.8 7.29 ;
      RECT 17.63 5.92 17.8 7.29 ;
      RECT 16.15 7.025 16.44 7.255 ;
      RECT 17.57 5.92 17.86 6.15 ;
      RECT 17.57 5.95 18.03 6.12 ;
      RECT 14.2 2.705 14.54 3.055 ;
      RECT 14.29 2.025 14.46 3.055 ;
      RECT 16.58 1.965 16.93 2.315 ;
      RECT 14.29 2.025 16.93 2.195 ;
      RECT 16.605 6.655 16.93 6.98 ;
      RECT 11.145 6.605 11.495 6.955 ;
      RECT 16.58 6.655 16.93 6.885 ;
      RECT 10.945 6.655 11.495 6.885 ;
      RECT 10.775 6.685 16.93 6.855 ;
      RECT 15.805 2.365 16.125 2.685 ;
      RECT 15.775 2.365 16.125 2.595 ;
      RECT 15.605 2.395 16.125 2.565 ;
      RECT 15.805 6.255 16.125 6.545 ;
      RECT 15.775 6.285 16.125 6.515 ;
      RECT 15.605 6.315 16.125 6.485 ;
      RECT 11.495 2.985 11.645 3.26 ;
      RECT 12.035 2.065 12.04 2.285 ;
      RECT 13.185 2.265 13.2 2.463 ;
      RECT 13.15 2.257 13.185 2.47 ;
      RECT 13.12 2.25 13.15 2.47 ;
      RECT 13.065 2.215 13.12 2.47 ;
      RECT 13 2.152 13.065 2.47 ;
      RECT 12.995 2.117 13 2.468 ;
      RECT 12.99 2.112 12.995 2.46 ;
      RECT 12.985 2.107 12.99 2.446 ;
      RECT 12.98 2.104 12.985 2.439 ;
      RECT 12.935 2.094 12.98 2.39 ;
      RECT 12.915 2.081 12.935 2.325 ;
      RECT 12.91 2.076 12.915 2.298 ;
      RECT 12.905 2.075 12.91 2.291 ;
      RECT 12.9 2.074 12.905 2.284 ;
      RECT 12.815 2.059 12.9 2.23 ;
      RECT 12.785 2.04 12.815 2.18 ;
      RECT 12.705 2.023 12.785 2.165 ;
      RECT 12.67 2.01 12.705 2.15 ;
      RECT 12.662 2.01 12.67 2.145 ;
      RECT 12.576 2.011 12.662 2.145 ;
      RECT 12.49 2.013 12.576 2.145 ;
      RECT 12.465 2.014 12.49 2.149 ;
      RECT 12.39 2.02 12.465 2.164 ;
      RECT 12.307 2.032 12.39 2.188 ;
      RECT 12.221 2.045 12.307 2.214 ;
      RECT 12.135 2.058 12.221 2.24 ;
      RECT 12.1 2.067 12.135 2.259 ;
      RECT 12.05 2.067 12.1 2.272 ;
      RECT 12.04 2.065 12.05 2.283 ;
      RECT 12.025 2.062 12.035 2.285 ;
      RECT 12.01 2.054 12.025 2.293 ;
      RECT 11.995 2.046 12.01 2.313 ;
      RECT 11.99 2.041 11.995 2.37 ;
      RECT 11.975 2.036 11.99 2.443 ;
      RECT 11.97 2.031 11.975 2.485 ;
      RECT 11.965 2.029 11.97 2.513 ;
      RECT 11.96 2.027 11.965 2.535 ;
      RECT 11.95 2.023 11.96 2.578 ;
      RECT 11.945 2.02 11.95 2.603 ;
      RECT 11.94 2.018 11.945 2.623 ;
      RECT 11.935 2.016 11.94 2.647 ;
      RECT 11.93 2.012 11.935 2.67 ;
      RECT 11.925 2.008 11.93 2.693 ;
      RECT 11.89 1.998 11.925 2.8 ;
      RECT 11.885 1.988 11.89 2.898 ;
      RECT 11.88 1.986 11.885 2.925 ;
      RECT 11.875 1.985 11.88 2.945 ;
      RECT 11.87 1.977 11.875 2.965 ;
      RECT 11.865 1.972 11.87 3 ;
      RECT 11.86 1.97 11.865 3.018 ;
      RECT 11.855 1.97 11.86 3.043 ;
      RECT 11.85 1.97 11.855 3.065 ;
      RECT 11.815 1.97 11.85 3.108 ;
      RECT 11.79 1.97 11.815 3.137 ;
      RECT 11.78 1.97 11.79 2.323 ;
      RECT 11.783 2.38 11.79 3.147 ;
      RECT 11.78 2.437 11.783 3.15 ;
      RECT 11.775 1.97 11.78 2.295 ;
      RECT 11.775 2.487 11.78 3.153 ;
      RECT 11.765 1.97 11.775 2.285 ;
      RECT 11.77 2.54 11.775 3.156 ;
      RECT 11.765 2.625 11.77 3.16 ;
      RECT 11.755 1.97 11.765 2.273 ;
      RECT 11.76 2.672 11.765 3.164 ;
      RECT 11.755 2.747 11.76 3.168 ;
      RECT 11.72 1.97 11.755 2.248 ;
      RECT 11.745 2.83 11.755 3.173 ;
      RECT 11.735 2.897 11.745 3.18 ;
      RECT 11.73 2.925 11.735 3.185 ;
      RECT 11.72 2.938 11.73 3.191 ;
      RECT 11.675 1.97 11.72 2.205 ;
      RECT 11.715 2.943 11.72 3.198 ;
      RECT 11.675 2.96 11.715 3.26 ;
      RECT 11.67 1.972 11.675 2.178 ;
      RECT 11.645 2.98 11.675 3.26 ;
      RECT 11.665 1.977 11.67 2.15 ;
      RECT 11.455 2.989 11.495 3.26 ;
      RECT 11.43 2.997 11.455 3.23 ;
      RECT 11.385 3.005 11.43 3.23 ;
      RECT 11.37 3.01 11.385 3.225 ;
      RECT 11.36 3.01 11.37 3.219 ;
      RECT 11.35 3.017 11.36 3.216 ;
      RECT 11.345 3.055 11.35 3.205 ;
      RECT 11.34 3.117 11.345 3.183 ;
      RECT 12.61 2.992 12.795 3.215 ;
      RECT 12.61 3.007 12.8 3.211 ;
      RECT 12.6 2.28 12.685 3.21 ;
      RECT 12.6 3.007 12.805 3.204 ;
      RECT 12.595 3.015 12.805 3.203 ;
      RECT 12.8 2.735 13.12 3.055 ;
      RECT 12.595 2.907 12.765 2.998 ;
      RECT 12.59 2.907 12.765 2.98 ;
      RECT 12.58 2.715 12.715 2.955 ;
      RECT 12.575 2.715 12.715 2.9 ;
      RECT 12.535 2.295 12.705 2.8 ;
      RECT 12.52 2.295 12.705 2.67 ;
      RECT 12.515 2.295 12.705 2.623 ;
      RECT 12.51 2.295 12.705 2.603 ;
      RECT 12.505 2.295 12.705 2.578 ;
      RECT 12.475 2.295 12.735 2.555 ;
      RECT 12.485 2.292 12.695 2.555 ;
      RECT 12.61 2.287 12.695 3.215 ;
      RECT 12.495 2.28 12.685 2.555 ;
      RECT 12.49 2.285 12.685 2.555 ;
      RECT 11.32 2.497 11.505 2.71 ;
      RECT 11.32 2.505 11.515 2.703 ;
      RECT 11.3 2.505 11.515 2.7 ;
      RECT 11.295 2.505 11.515 2.685 ;
      RECT 11.225 2.42 11.485 2.68 ;
      RECT 11.225 2.565 11.52 2.593 ;
      RECT 10.88 3.02 11.14 3.28 ;
      RECT 10.905 2.965 11.1 3.28 ;
      RECT 10.9 2.714 11.08 3.008 ;
      RECT 10.9 2.72 11.09 3.008 ;
      RECT 10.88 2.722 11.09 2.953 ;
      RECT 10.875 2.732 11.09 2.82 ;
      RECT 10.905 2.712 11.08 3.28 ;
      RECT 10.991 2.71 11.08 3.28 ;
      RECT 10.85 1.93 10.885 2.3 ;
      RECT 10.64 2.04 10.645 2.3 ;
      RECT 10.885 1.937 10.9 2.3 ;
      RECT 10.775 1.93 10.85 2.378 ;
      RECT 10.765 1.93 10.775 2.463 ;
      RECT 10.74 1.93 10.765 2.498 ;
      RECT 10.7 1.93 10.74 2.566 ;
      RECT 10.69 1.937 10.7 2.618 ;
      RECT 10.66 2.04 10.69 2.659 ;
      RECT 10.655 2.04 10.66 2.698 ;
      RECT 10.645 2.04 10.655 2.718 ;
      RECT 10.64 2.335 10.645 2.755 ;
      RECT 10.635 2.352 10.64 2.775 ;
      RECT 10.62 2.415 10.635 2.815 ;
      RECT 10.615 2.458 10.62 2.85 ;
      RECT 10.61 2.466 10.615 2.863 ;
      RECT 10.6 2.48 10.61 2.885 ;
      RECT 10.575 2.515 10.6 2.95 ;
      RECT 10.565 2.55 10.575 3.013 ;
      RECT 10.545 2.58 10.565 3.074 ;
      RECT 10.53 2.616 10.545 3.141 ;
      RECT 10.52 2.644 10.53 3.18 ;
      RECT 10.51 2.666 10.52 3.2 ;
      RECT 10.505 2.676 10.51 3.211 ;
      RECT 10.5 2.685 10.505 3.214 ;
      RECT 10.49 2.703 10.5 3.218 ;
      RECT 10.48 2.721 10.49 3.219 ;
      RECT 10.455 2.76 10.48 3.216 ;
      RECT 10.435 2.802 10.455 3.213 ;
      RECT 10.42 2.84 10.435 3.212 ;
      RECT 10.385 2.875 10.42 3.209 ;
      RECT 10.38 2.897 10.385 3.207 ;
      RECT 10.315 2.937 10.38 3.204 ;
      RECT 10.31 2.977 10.315 3.2 ;
      RECT 10.295 2.987 10.31 3.191 ;
      RECT 10.285 3.107 10.295 3.176 ;
      RECT 10.765 3.52 10.775 3.78 ;
      RECT 10.765 3.523 10.785 3.779 ;
      RECT 10.755 3.513 10.765 3.778 ;
      RECT 10.745 3.528 10.825 3.774 ;
      RECT 10.73 3.507 10.745 3.772 ;
      RECT 10.705 3.532 10.83 3.768 ;
      RECT 10.69 3.492 10.705 3.763 ;
      RECT 10.69 3.534 10.84 3.762 ;
      RECT 10.69 3.542 10.855 3.755 ;
      RECT 10.63 3.479 10.69 3.745 ;
      RECT 10.62 3.466 10.63 3.727 ;
      RECT 10.595 3.456 10.62 3.717 ;
      RECT 10.59 3.446 10.595 3.709 ;
      RECT 10.525 3.542 10.855 3.691 ;
      RECT 10.44 3.542 10.855 3.653 ;
      RECT 10.33 3.37 10.59 3.63 ;
      RECT 10.705 3.5 10.73 3.768 ;
      RECT 10.745 3.51 10.755 3.774 ;
      RECT 10.33 3.518 10.77 3.63 ;
      RECT 10.515 7.765 10.805 7.995 ;
      RECT 10.575 7.025 10.745 7.995 ;
      RECT 10.475 7.055 10.845 7.425 ;
      RECT 10.515 7.025 10.805 7.425 ;
      RECT 9.545 3.275 9.575 3.575 ;
      RECT 9.32 3.26 9.325 3.535 ;
      RECT 9.12 3.26 9.275 3.52 ;
      RECT 10.42 1.975 10.45 2.235 ;
      RECT 10.41 1.975 10.42 2.343 ;
      RECT 10.39 1.975 10.41 2.353 ;
      RECT 10.375 1.975 10.39 2.365 ;
      RECT 10.32 1.975 10.375 2.415 ;
      RECT 10.305 1.975 10.32 2.463 ;
      RECT 10.275 1.975 10.305 2.498 ;
      RECT 10.22 1.975 10.275 2.56 ;
      RECT 10.2 1.975 10.22 2.628 ;
      RECT 10.195 1.975 10.2 2.658 ;
      RECT 10.19 1.975 10.195 2.67 ;
      RECT 10.185 2.092 10.19 2.688 ;
      RECT 10.165 2.11 10.185 2.713 ;
      RECT 10.145 2.137 10.165 2.763 ;
      RECT 10.14 2.157 10.145 2.794 ;
      RECT 10.135 2.165 10.14 2.811 ;
      RECT 10.12 2.191 10.135 2.84 ;
      RECT 10.105 2.233 10.12 2.875 ;
      RECT 10.1 2.262 10.105 2.898 ;
      RECT 10.095 2.277 10.1 2.911 ;
      RECT 10.09 2.3 10.095 2.922 ;
      RECT 10.08 2.32 10.09 2.94 ;
      RECT 10.07 2.35 10.08 2.963 ;
      RECT 10.065 2.372 10.07 2.983 ;
      RECT 10.06 2.387 10.065 2.998 ;
      RECT 10.045 2.417 10.06 3.025 ;
      RECT 10.04 2.447 10.045 3.051 ;
      RECT 10.035 2.465 10.04 3.063 ;
      RECT 10.025 2.495 10.035 3.082 ;
      RECT 10.015 2.52 10.025 3.107 ;
      RECT 10.01 2.54 10.015 3.126 ;
      RECT 10.005 2.557 10.01 3.139 ;
      RECT 9.995 2.583 10.005 3.158 ;
      RECT 9.985 2.621 9.995 3.185 ;
      RECT 9.98 2.647 9.985 3.205 ;
      RECT 9.975 2.657 9.98 3.215 ;
      RECT 9.97 2.67 9.975 3.23 ;
      RECT 9.965 2.685 9.97 3.24 ;
      RECT 9.96 2.707 9.965 3.255 ;
      RECT 9.955 2.725 9.96 3.266 ;
      RECT 9.95 2.735 9.955 3.277 ;
      RECT 9.945 2.743 9.95 3.289 ;
      RECT 9.94 2.751 9.945 3.3 ;
      RECT 9.935 2.777 9.94 3.313 ;
      RECT 9.925 2.805 9.935 3.326 ;
      RECT 9.92 2.835 9.925 3.335 ;
      RECT 9.915 2.85 9.92 3.342 ;
      RECT 9.9 2.875 9.915 3.349 ;
      RECT 9.895 2.897 9.9 3.355 ;
      RECT 9.89 2.922 9.895 3.358 ;
      RECT 9.881 2.95 9.89 3.362 ;
      RECT 9.875 2.967 9.881 3.367 ;
      RECT 9.87 2.985 9.875 3.371 ;
      RECT 9.865 2.997 9.87 3.374 ;
      RECT 9.86 3.018 9.865 3.378 ;
      RECT 9.855 3.036 9.86 3.381 ;
      RECT 9.85 3.05 9.855 3.384 ;
      RECT 9.845 3.067 9.85 3.387 ;
      RECT 9.84 3.08 9.845 3.39 ;
      RECT 9.815 3.117 9.84 3.398 ;
      RECT 9.81 3.162 9.815 3.407 ;
      RECT 9.805 3.19 9.81 3.41 ;
      RECT 9.795 3.21 9.805 3.414 ;
      RECT 9.79 3.23 9.795 3.419 ;
      RECT 9.785 3.245 9.79 3.422 ;
      RECT 9.765 3.255 9.785 3.429 ;
      RECT 9.7 3.262 9.765 3.455 ;
      RECT 9.665 3.265 9.7 3.483 ;
      RECT 9.65 3.268 9.665 3.498 ;
      RECT 9.64 3.269 9.65 3.513 ;
      RECT 9.63 3.27 9.64 3.53 ;
      RECT 9.625 3.27 9.63 3.545 ;
      RECT 9.62 3.27 9.625 3.553 ;
      RECT 9.605 3.271 9.62 3.568 ;
      RECT 9.575 3.273 9.605 3.575 ;
      RECT 9.465 3.28 9.545 3.575 ;
      RECT 9.42 3.285 9.465 3.575 ;
      RECT 9.41 3.286 9.42 3.565 ;
      RECT 9.4 3.287 9.41 3.558 ;
      RECT 9.38 3.289 9.4 3.553 ;
      RECT 9.37 3.26 9.38 3.548 ;
      RECT 9.325 3.26 9.37 3.54 ;
      RECT 9.295 3.26 9.32 3.53 ;
      RECT 9.275 3.26 9.295 3.523 ;
      RECT 9.555 2.06 9.815 2.32 ;
      RECT 9.435 2.075 9.445 2.24 ;
      RECT 9.42 2.075 9.425 2.235 ;
      RECT 6.785 1.915 6.97 2.205 ;
      RECT 8.6 2.04 8.615 2.195 ;
      RECT 6.75 1.915 6.775 2.175 ;
      RECT 9.165 1.965 9.17 2.107 ;
      RECT 9.08 1.96 9.105 2.1 ;
      RECT 9.48 2.077 9.555 2.27 ;
      RECT 9.465 2.075 9.48 2.253 ;
      RECT 9.445 2.075 9.465 2.245 ;
      RECT 9.425 2.075 9.435 2.238 ;
      RECT 9.38 2.07 9.42 2.228 ;
      RECT 9.34 2.045 9.38 2.213 ;
      RECT 9.325 2.02 9.34 2.203 ;
      RECT 9.32 2.014 9.325 2.201 ;
      RECT 9.285 2.006 9.32 2.184 ;
      RECT 9.28 1.999 9.285 2.172 ;
      RECT 9.26 1.994 9.28 2.16 ;
      RECT 9.25 1.988 9.26 2.145 ;
      RECT 9.23 1.983 9.25 2.13 ;
      RECT 9.22 1.978 9.23 2.123 ;
      RECT 9.215 1.976 9.22 2.118 ;
      RECT 9.21 1.975 9.215 2.115 ;
      RECT 9.17 1.97 9.21 2.111 ;
      RECT 9.15 1.964 9.165 2.106 ;
      RECT 9.115 1.961 9.15 2.103 ;
      RECT 9.105 1.96 9.115 2.101 ;
      RECT 9.045 1.96 9.08 2.098 ;
      RECT 9 1.96 9.045 2.098 ;
      RECT 8.95 1.96 9 2.101 ;
      RECT 8.935 1.962 8.95 2.103 ;
      RECT 8.92 1.965 8.935 2.104 ;
      RECT 8.91 1.97 8.92 2.105 ;
      RECT 8.88 1.975 8.91 2.11 ;
      RECT 8.87 1.981 8.88 2.118 ;
      RECT 8.86 1.983 8.87 2.122 ;
      RECT 8.85 1.987 8.86 2.126 ;
      RECT 8.825 1.993 8.85 2.134 ;
      RECT 8.815 1.998 8.825 2.142 ;
      RECT 8.8 2.002 8.815 2.146 ;
      RECT 8.765 2.008 8.8 2.154 ;
      RECT 8.745 2.013 8.765 2.164 ;
      RECT 8.715 2.02 8.745 2.173 ;
      RECT 8.67 2.029 8.715 2.187 ;
      RECT 8.665 2.034 8.67 2.198 ;
      RECT 8.645 2.037 8.665 2.199 ;
      RECT 8.615 2.04 8.645 2.197 ;
      RECT 8.58 2.04 8.6 2.193 ;
      RECT 8.51 2.04 8.58 2.184 ;
      RECT 8.495 2.037 8.51 2.176 ;
      RECT 8.455 2.03 8.495 2.171 ;
      RECT 8.43 2.02 8.455 2.164 ;
      RECT 8.425 2.014 8.43 2.161 ;
      RECT 8.385 2.008 8.425 2.158 ;
      RECT 8.37 2.001 8.385 2.153 ;
      RECT 8.35 1.997 8.37 2.148 ;
      RECT 8.335 1.992 8.35 2.144 ;
      RECT 8.32 1.987 8.335 2.142 ;
      RECT 8.305 1.983 8.32 2.141 ;
      RECT 8.29 1.981 8.305 2.137 ;
      RECT 8.28 1.979 8.29 2.132 ;
      RECT 8.265 1.976 8.28 2.128 ;
      RECT 8.255 1.974 8.265 2.123 ;
      RECT 8.235 1.971 8.255 2.119 ;
      RECT 8.19 1.97 8.235 2.117 ;
      RECT 8.13 1.972 8.19 2.118 ;
      RECT 8.11 1.974 8.13 2.12 ;
      RECT 8.08 1.977 8.11 2.121 ;
      RECT 8.03 1.982 8.08 2.123 ;
      RECT 8.025 1.985 8.03 2.125 ;
      RECT 8.015 1.987 8.025 2.128 ;
      RECT 8.01 1.989 8.015 2.131 ;
      RECT 7.96 1.992 8.01 2.138 ;
      RECT 7.94 1.996 7.96 2.15 ;
      RECT 7.93 1.999 7.94 2.156 ;
      RECT 7.92 2 7.93 2.159 ;
      RECT 7.881 2.003 7.92 2.161 ;
      RECT 7.795 2.01 7.881 2.164 ;
      RECT 7.721 2.02 7.795 2.168 ;
      RECT 7.635 2.031 7.721 2.173 ;
      RECT 7.62 2.038 7.635 2.175 ;
      RECT 7.565 2.042 7.62 2.176 ;
      RECT 7.551 2.045 7.565 2.178 ;
      RECT 7.465 2.045 7.551 2.18 ;
      RECT 7.425 2.042 7.465 2.183 ;
      RECT 7.401 2.038 7.425 2.185 ;
      RECT 7.315 2.028 7.401 2.188 ;
      RECT 7.285 2.017 7.315 2.189 ;
      RECT 7.266 2.013 7.285 2.188 ;
      RECT 7.18 2.006 7.266 2.185 ;
      RECT 7.12 1.995 7.18 2.182 ;
      RECT 7.1 1.987 7.12 2.18 ;
      RECT 7.065 1.982 7.1 2.179 ;
      RECT 7.04 1.977 7.065 2.178 ;
      RECT 7.01 1.972 7.04 2.177 ;
      RECT 6.985 1.915 7.01 2.176 ;
      RECT 6.97 1.915 6.985 2.2 ;
      RECT 6.775 1.915 6.785 2.2 ;
      RECT 8.55 2.935 8.555 3.075 ;
      RECT 8.21 2.935 8.245 3.073 ;
      RECT 7.785 2.92 7.8 3.065 ;
      RECT 9.615 2.7 9.705 2.96 ;
      RECT 9.445 2.565 9.545 2.96 ;
      RECT 6.48 2.54 6.56 2.75 ;
      RECT 9.57 2.677 9.615 2.96 ;
      RECT 9.56 2.647 9.57 2.96 ;
      RECT 9.545 2.57 9.56 2.96 ;
      RECT 9.36 2.565 9.445 2.925 ;
      RECT 9.355 2.567 9.36 2.92 ;
      RECT 9.35 2.572 9.355 2.92 ;
      RECT 9.315 2.672 9.35 2.92 ;
      RECT 9.305 2.7 9.315 2.92 ;
      RECT 9.295 2.715 9.305 2.92 ;
      RECT 9.285 2.727 9.295 2.92 ;
      RECT 9.28 2.737 9.285 2.92 ;
      RECT 9.265 2.747 9.28 2.922 ;
      RECT 9.26 2.762 9.265 2.924 ;
      RECT 9.245 2.775 9.26 2.926 ;
      RECT 9.24 2.79 9.245 2.929 ;
      RECT 9.22 2.8 9.24 2.933 ;
      RECT 9.205 2.81 9.22 2.936 ;
      RECT 9.17 2.817 9.205 2.941 ;
      RECT 9.126 2.824 9.17 2.949 ;
      RECT 9.04 2.836 9.126 2.962 ;
      RECT 9.015 2.847 9.04 2.973 ;
      RECT 8.985 2.852 9.015 2.978 ;
      RECT 8.95 2.857 8.985 2.986 ;
      RECT 8.92 2.862 8.95 2.993 ;
      RECT 8.895 2.867 8.92 2.998 ;
      RECT 8.83 2.874 8.895 3.007 ;
      RECT 8.76 2.887 8.83 3.023 ;
      RECT 8.73 2.897 8.76 3.035 ;
      RECT 8.705 2.902 8.73 3.042 ;
      RECT 8.65 2.909 8.705 3.05 ;
      RECT 8.645 2.916 8.65 3.055 ;
      RECT 8.64 2.918 8.645 3.056 ;
      RECT 8.625 2.92 8.64 3.058 ;
      RECT 8.62 2.92 8.625 3.061 ;
      RECT 8.555 2.927 8.62 3.068 ;
      RECT 8.52 2.937 8.55 3.078 ;
      RECT 8.503 2.94 8.52 3.08 ;
      RECT 8.417 2.939 8.503 3.079 ;
      RECT 8.331 2.937 8.417 3.076 ;
      RECT 8.245 2.936 8.331 3.074 ;
      RECT 8.144 2.934 8.21 3.073 ;
      RECT 8.058 2.931 8.144 3.071 ;
      RECT 7.972 2.927 8.058 3.069 ;
      RECT 7.886 2.924 7.972 3.068 ;
      RECT 7.8 2.921 7.886 3.066 ;
      RECT 7.7 2.92 7.785 3.063 ;
      RECT 7.65 2.918 7.7 3.061 ;
      RECT 7.63 2.915 7.65 3.059 ;
      RECT 7.61 2.913 7.63 3.056 ;
      RECT 7.585 2.909 7.61 3.053 ;
      RECT 7.54 2.903 7.585 3.048 ;
      RECT 7.5 2.897 7.54 3.04 ;
      RECT 7.475 2.892 7.5 3.033 ;
      RECT 7.42 2.885 7.475 3.025 ;
      RECT 7.396 2.878 7.42 3.018 ;
      RECT 7.31 2.869 7.396 3.008 ;
      RECT 7.28 2.861 7.31 2.998 ;
      RECT 7.25 2.857 7.28 2.993 ;
      RECT 7.245 2.854 7.25 2.99 ;
      RECT 7.24 2.853 7.245 2.99 ;
      RECT 7.165 2.846 7.24 2.983 ;
      RECT 7.126 2.837 7.165 2.972 ;
      RECT 7.04 2.827 7.126 2.96 ;
      RECT 7 2.817 7.04 2.948 ;
      RECT 6.961 2.812 7 2.941 ;
      RECT 6.875 2.802 6.961 2.93 ;
      RECT 6.835 2.79 6.875 2.919 ;
      RECT 6.8 2.775 6.835 2.912 ;
      RECT 6.79 2.765 6.8 2.909 ;
      RECT 6.77 2.75 6.79 2.907 ;
      RECT 6.74 2.72 6.77 2.903 ;
      RECT 6.73 2.7 6.74 2.898 ;
      RECT 6.725 2.692 6.73 2.895 ;
      RECT 6.72 2.685 6.725 2.893 ;
      RECT 6.705 2.672 6.72 2.886 ;
      RECT 6.7 2.662 6.705 2.878 ;
      RECT 6.695 2.655 6.7 2.873 ;
      RECT 6.69 2.65 6.695 2.869 ;
      RECT 6.675 2.637 6.69 2.861 ;
      RECT 6.67 2.547 6.675 2.85 ;
      RECT 6.665 2.542 6.67 2.843 ;
      RECT 6.59 2.54 6.665 2.803 ;
      RECT 6.56 2.54 6.59 2.758 ;
      RECT 6.465 2.545 6.48 2.745 ;
      RECT 8.95 2.25 9.21 2.51 ;
      RECT 8.935 2.238 9.115 2.475 ;
      RECT 8.93 2.239 9.115 2.473 ;
      RECT 8.915 2.243 9.125 2.463 ;
      RECT 8.91 2.248 9.13 2.433 ;
      RECT 8.915 2.245 9.13 2.463 ;
      RECT 8.93 2.24 9.125 2.473 ;
      RECT 8.95 2.237 9.115 2.51 ;
      RECT 8.95 2.236 9.105 2.51 ;
      RECT 8.975 2.235 9.105 2.51 ;
      RECT 8.535 2.48 8.795 2.74 ;
      RECT 8.41 2.525 8.795 2.735 ;
      RECT 8.4 2.53 8.795 2.73 ;
      RECT 8.415 3.47 8.43 3.78 ;
      RECT 7.01 3.24 7.02 3.37 ;
      RECT 6.79 3.235 6.895 3.37 ;
      RECT 6.705 3.24 6.755 3.37 ;
      RECT 5.255 1.975 5.26 3.08 ;
      RECT 8.51 3.562 8.515 3.698 ;
      RECT 8.505 3.557 8.51 3.758 ;
      RECT 8.5 3.555 8.505 3.771 ;
      RECT 8.485 3.552 8.5 3.773 ;
      RECT 8.48 3.547 8.485 3.775 ;
      RECT 8.475 3.543 8.48 3.778 ;
      RECT 8.46 3.538 8.475 3.78 ;
      RECT 8.43 3.53 8.46 3.78 ;
      RECT 8.391 3.47 8.415 3.78 ;
      RECT 8.305 3.47 8.391 3.777 ;
      RECT 8.275 3.47 8.305 3.77 ;
      RECT 8.25 3.47 8.275 3.763 ;
      RECT 8.225 3.47 8.25 3.755 ;
      RECT 8.21 3.47 8.225 3.748 ;
      RECT 8.185 3.47 8.21 3.74 ;
      RECT 8.17 3.47 8.185 3.733 ;
      RECT 8.13 3.48 8.17 3.722 ;
      RECT 8.12 3.475 8.13 3.712 ;
      RECT 8.116 3.474 8.12 3.709 ;
      RECT 8.03 3.466 8.116 3.692 ;
      RECT 7.997 3.455 8.03 3.669 ;
      RECT 7.911 3.444 7.997 3.647 ;
      RECT 7.825 3.428 7.911 3.616 ;
      RECT 7.755 3.413 7.825 3.588 ;
      RECT 7.745 3.406 7.755 3.575 ;
      RECT 7.715 3.403 7.745 3.565 ;
      RECT 7.69 3.399 7.715 3.558 ;
      RECT 7.675 3.396 7.69 3.553 ;
      RECT 7.67 3.395 7.675 3.548 ;
      RECT 7.64 3.39 7.67 3.541 ;
      RECT 7.635 3.385 7.64 3.536 ;
      RECT 7.62 3.382 7.635 3.531 ;
      RECT 7.615 3.377 7.62 3.526 ;
      RECT 7.595 3.372 7.615 3.523 ;
      RECT 7.58 3.367 7.595 3.515 ;
      RECT 7.565 3.361 7.58 3.51 ;
      RECT 7.535 3.352 7.565 3.503 ;
      RECT 7.53 3.345 7.535 3.495 ;
      RECT 7.525 3.343 7.53 3.493 ;
      RECT 7.52 3.342 7.525 3.49 ;
      RECT 7.48 3.335 7.52 3.483 ;
      RECT 7.466 3.325 7.48 3.473 ;
      RECT 7.415 3.314 7.466 3.461 ;
      RECT 7.39 3.3 7.415 3.447 ;
      RECT 7.365 3.289 7.39 3.439 ;
      RECT 7.345 3.278 7.365 3.433 ;
      RECT 7.335 3.272 7.345 3.428 ;
      RECT 7.33 3.27 7.335 3.424 ;
      RECT 7.31 3.265 7.33 3.419 ;
      RECT 7.28 3.255 7.31 3.409 ;
      RECT 7.275 3.247 7.28 3.402 ;
      RECT 7.26 3.245 7.275 3.398 ;
      RECT 7.24 3.245 7.26 3.393 ;
      RECT 7.235 3.244 7.24 3.391 ;
      RECT 7.23 3.244 7.235 3.388 ;
      RECT 7.19 3.243 7.23 3.383 ;
      RECT 7.165 3.242 7.19 3.378 ;
      RECT 7.105 3.241 7.165 3.375 ;
      RECT 7.02 3.24 7.105 3.373 ;
      RECT 6.981 3.239 7.01 3.37 ;
      RECT 6.895 3.237 6.981 3.37 ;
      RECT 6.755 3.237 6.79 3.37 ;
      RECT 6.665 3.241 6.705 3.373 ;
      RECT 6.65 3.244 6.665 3.38 ;
      RECT 6.64 3.245 6.65 3.387 ;
      RECT 6.615 3.248 6.64 3.392 ;
      RECT 6.61 3.25 6.615 3.395 ;
      RECT 6.56 3.252 6.61 3.396 ;
      RECT 6.521 3.256 6.56 3.398 ;
      RECT 6.435 3.258 6.521 3.401 ;
      RECT 6.417 3.26 6.435 3.403 ;
      RECT 6.331 3.263 6.417 3.405 ;
      RECT 6.245 3.267 6.331 3.408 ;
      RECT 6.208 3.271 6.245 3.411 ;
      RECT 6.122 3.274 6.208 3.414 ;
      RECT 6.036 3.278 6.122 3.417 ;
      RECT 5.95 3.283 6.036 3.421 ;
      RECT 5.93 3.285 5.95 3.424 ;
      RECT 5.91 3.284 5.93 3.425 ;
      RECT 5.861 3.281 5.91 3.426 ;
      RECT 5.775 3.276 5.861 3.429 ;
      RECT 5.725 3.271 5.775 3.431 ;
      RECT 5.701 3.269 5.725 3.432 ;
      RECT 5.615 3.264 5.701 3.434 ;
      RECT 5.59 3.26 5.615 3.433 ;
      RECT 5.58 3.257 5.59 3.431 ;
      RECT 5.57 3.25 5.58 3.428 ;
      RECT 5.565 3.23 5.57 3.423 ;
      RECT 5.555 3.2 5.565 3.418 ;
      RECT 5.54 3.07 5.555 3.409 ;
      RECT 5.535 3.062 5.54 3.402 ;
      RECT 5.515 3.055 5.535 3.394 ;
      RECT 5.51 3.037 5.515 3.386 ;
      RECT 5.5 3.017 5.51 3.381 ;
      RECT 5.495 2.99 5.5 3.377 ;
      RECT 5.49 2.967 5.495 3.374 ;
      RECT 5.47 2.925 5.49 3.366 ;
      RECT 5.435 2.84 5.47 3.35 ;
      RECT 5.43 2.772 5.435 3.338 ;
      RECT 5.415 2.742 5.43 3.332 ;
      RECT 5.41 1.987 5.415 2.233 ;
      RECT 5.4 2.712 5.415 3.323 ;
      RECT 5.405 1.982 5.41 2.265 ;
      RECT 5.4 1.977 5.405 2.308 ;
      RECT 5.395 1.975 5.4 2.343 ;
      RECT 5.38 2.675 5.4 3.313 ;
      RECT 5.39 1.975 5.395 2.38 ;
      RECT 5.375 1.975 5.39 2.478 ;
      RECT 5.375 2.648 5.38 3.306 ;
      RECT 5.37 1.975 5.375 2.553 ;
      RECT 5.37 2.636 5.375 3.303 ;
      RECT 5.365 1.975 5.37 2.585 ;
      RECT 5.365 2.615 5.37 3.3 ;
      RECT 5.36 1.975 5.365 3.297 ;
      RECT 5.325 1.975 5.36 3.283 ;
      RECT 5.31 1.975 5.325 3.265 ;
      RECT 5.29 1.975 5.31 3.255 ;
      RECT 5.265 1.975 5.29 3.238 ;
      RECT 5.26 1.975 5.265 3.188 ;
      RECT 5.25 1.975 5.255 3.018 ;
      RECT 5.245 1.975 5.25 2.925 ;
      RECT 5.24 1.975 5.245 2.838 ;
      RECT 5.235 1.975 5.24 2.77 ;
      RECT 5.23 1.975 5.235 2.713 ;
      RECT 5.22 1.975 5.23 2.608 ;
      RECT 5.215 1.975 5.22 2.48 ;
      RECT 5.21 1.975 5.215 2.398 ;
      RECT 5.205 1.977 5.21 2.315 ;
      RECT 5.2 1.982 5.205 2.248 ;
      RECT 5.195 1.987 5.2 2.175 ;
      RECT 8.01 2.305 8.27 2.565 ;
      RECT 8.03 2.272 8.24 2.565 ;
      RECT 8.03 2.27 8.23 2.565 ;
      RECT 8.04 2.257 8.23 2.565 ;
      RECT 8.04 2.255 8.155 2.565 ;
      RECT 7.515 2.38 7.69 2.66 ;
      RECT 7.51 2.38 7.69 2.658 ;
      RECT 7.51 2.38 7.705 2.655 ;
      RECT 7.5 2.38 7.705 2.653 ;
      RECT 7.445 2.38 7.705 2.64 ;
      RECT 7.445 2.455 7.71 2.618 ;
      RECT 6.99 2.392 7.01 2.635 ;
      RECT 6.99 2.392 7.05 2.634 ;
      RECT 6.985 2.394 7.05 2.633 ;
      RECT 6.985 2.394 7.136 2.632 ;
      RECT 6.985 2.394 7.205 2.631 ;
      RECT 6.985 2.394 7.225 2.623 ;
      RECT 6.965 2.397 7.225 2.621 ;
      RECT 6.95 2.407 7.225 2.606 ;
      RECT 6.95 2.407 7.24 2.605 ;
      RECT 6.945 2.416 7.24 2.597 ;
      RECT 6.945 2.416 7.245 2.593 ;
      RECT 7.05 2.33 7.31 2.59 ;
      RECT 6.94 2.418 7.31 2.475 ;
      RECT 7.01 2.385 7.31 2.59 ;
      RECT 6.975 3.578 6.98 3.785 ;
      RECT 6.925 3.572 6.975 3.784 ;
      RECT 6.892 3.586 6.985 3.783 ;
      RECT 6.806 3.586 6.985 3.782 ;
      RECT 6.72 3.586 6.985 3.781 ;
      RECT 6.72 3.685 6.99 3.778 ;
      RECT 6.715 3.685 6.99 3.773 ;
      RECT 6.71 3.685 6.99 3.755 ;
      RECT 6.705 3.685 6.99 3.738 ;
      RECT 6.665 3.47 6.925 3.73 ;
      RECT 6.125 2.62 6.211 3.034 ;
      RECT 6.125 2.62 6.25 3.031 ;
      RECT 6.125 2.62 6.27 3.021 ;
      RECT 6.08 2.62 6.27 3.018 ;
      RECT 6.08 2.772 6.28 3.008 ;
      RECT 6.08 2.793 6.285 3.002 ;
      RECT 6.08 2.811 6.29 2.998 ;
      RECT 6.08 2.831 6.3 2.993 ;
      RECT 6.055 2.831 6.3 2.99 ;
      RECT 6.045 2.831 6.3 2.968 ;
      RECT 6.045 2.847 6.305 2.938 ;
      RECT 6.01 2.62 6.27 2.925 ;
      RECT 6.01 2.859 6.31 2.88 ;
      RECT 3.02 7.765 3.31 7.995 ;
      RECT 3.08 7.025 3.25 7.995 ;
      RECT 2.99 7.025 3.34 7.315 ;
      RECT 2.615 6.285 2.965 6.575 ;
      RECT 2.475 6.315 2.965 6.485 ;
      RECT 69.635 3.265 69.895 3.525 ;
      RECT 54.375 3.265 54.635 3.525 ;
      RECT 39.115 3.265 39.375 3.525 ;
      RECT 23.855 3.265 24.115 3.525 ;
      RECT 8.595 3.265 8.855 3.525 ;
    LAYER mcon ;
      RECT 80.03 6.32 80.2 6.49 ;
      RECT 80.035 6.315 80.205 6.485 ;
      RECT 64.77 6.32 64.94 6.49 ;
      RECT 64.775 6.315 64.945 6.485 ;
      RECT 49.51 6.32 49.68 6.49 ;
      RECT 49.515 6.315 49.685 6.485 ;
      RECT 34.25 6.32 34.42 6.49 ;
      RECT 34.255 6.315 34.425 6.485 ;
      RECT 18.99 6.32 19.16 6.49 ;
      RECT 18.995 6.315 19.165 6.485 ;
      RECT 80.03 7.8 80.2 7.97 ;
      RECT 79.68 0.1 79.85 0.27 ;
      RECT 79.68 8.61 79.85 8.78 ;
      RECT 79.66 2.76 79.83 2.93 ;
      RECT 79.66 5.95 79.83 6.12 ;
      RECT 79.04 0.91 79.21 1.08 ;
      RECT 79.04 2.39 79.21 2.56 ;
      RECT 79.04 6.32 79.21 6.49 ;
      RECT 79.04 7.8 79.21 7.97 ;
      RECT 78.69 0.1 78.86 0.27 ;
      RECT 78.69 8.61 78.86 8.78 ;
      RECT 78.67 2.76 78.84 2.93 ;
      RECT 78.67 5.95 78.84 6.12 ;
      RECT 77.99 0.105 78.16 0.275 ;
      RECT 77.99 8.605 78.16 8.775 ;
      RECT 77.68 2.025 77.85 2.195 ;
      RECT 77.68 6.685 77.85 6.855 ;
      RECT 77.31 0.105 77.48 0.275 ;
      RECT 77.31 8.605 77.48 8.775 ;
      RECT 77.25 0.915 77.42 1.085 ;
      RECT 77.25 1.655 77.42 1.825 ;
      RECT 77.25 7.055 77.42 7.225 ;
      RECT 77.25 7.795 77.42 7.965 ;
      RECT 76.875 2.395 77.045 2.565 ;
      RECT 76.875 6.315 77.045 6.485 ;
      RECT 76.63 0.105 76.8 0.275 ;
      RECT 76.63 8.605 76.8 8.775 ;
      RECT 75.95 0.105 76.12 0.275 ;
      RECT 75.95 8.605 76.12 8.775 ;
      RECT 74.49 1.415 74.66 1.585 ;
      RECT 74.05 2.28 74.22 2.45 ;
      RECT 74.03 1.415 74.2 1.585 ;
      RECT 73.655 3.025 73.825 3.195 ;
      RECT 73.57 1.415 73.74 1.585 ;
      RECT 73.545 2.3 73.715 2.47 ;
      RECT 73.11 1.415 73.28 1.585 ;
      RECT 72.725 1.99 72.895 2.16 ;
      RECT 72.65 1.415 72.82 1.585 ;
      RECT 72.41 3.03 72.58 3.2 ;
      RECT 72.365 2.52 72.535 2.69 ;
      RECT 72.355 8.605 72.525 8.775 ;
      RECT 72.19 1.415 72.36 1.585 ;
      RECT 72.045 6.685 72.215 6.855 ;
      RECT 71.94 2.73 72.11 2.9 ;
      RECT 71.75 1.95 71.92 2.12 ;
      RECT 71.73 1.415 71.9 1.585 ;
      RECT 71.7 3.56 71.87 3.73 ;
      RECT 71.675 8.605 71.845 8.775 ;
      RECT 71.615 7.055 71.785 7.225 ;
      RECT 71.615 7.795 71.785 7.965 ;
      RECT 71.365 3 71.535 3.17 ;
      RECT 71.27 1.415 71.44 1.585 ;
      RECT 71.27 2.16 71.44 2.33 ;
      RECT 71.24 6.315 71.41 6.485 ;
      RECT 70.995 8.605 71.165 8.775 ;
      RECT 70.81 1.415 70.98 1.585 ;
      RECT 70.47 3.385 70.64 3.555 ;
      RECT 70.41 2.585 70.58 2.755 ;
      RECT 70.35 1.415 70.52 1.585 ;
      RECT 70.315 8.605 70.485 8.775 ;
      RECT 69.97 2.255 70.14 2.425 ;
      RECT 69.89 1.415 70.06 1.585 ;
      RECT 69.705 3.305 69.875 3.475 ;
      RECT 69.46 2.545 69.63 2.715 ;
      RECT 69.43 1.415 69.6 1.585 ;
      RECT 69.365 3.575 69.535 3.745 ;
      RECT 69.09 2.27 69.26 2.44 ;
      RECT 68.97 1.415 69.14 1.585 ;
      RECT 68.56 2.47 68.73 2.64 ;
      RECT 68.51 1.415 68.68 1.585 ;
      RECT 68.05 1.415 68.22 1.585 ;
      RECT 68.04 2.415 68.21 2.585 ;
      RECT 67.835 2.015 68.005 2.185 ;
      RECT 67.835 3.595 68.005 3.765 ;
      RECT 67.59 1.415 67.76 1.585 ;
      RECT 67.525 2.56 67.695 2.73 ;
      RECT 67.13 1.415 67.3 1.585 ;
      RECT 67.115 2.785 67.285 2.955 ;
      RECT 66.67 1.415 66.84 1.585 ;
      RECT 66.405 3.085 66.575 3.255 ;
      RECT 66.26 1.995 66.43 2.165 ;
      RECT 66.21 1.415 66.38 1.585 ;
      RECT 64.77 7.8 64.94 7.97 ;
      RECT 64.42 0.1 64.59 0.27 ;
      RECT 64.42 8.61 64.59 8.78 ;
      RECT 64.4 2.76 64.57 2.93 ;
      RECT 64.4 5.95 64.57 6.12 ;
      RECT 63.78 0.91 63.95 1.08 ;
      RECT 63.78 2.39 63.95 2.56 ;
      RECT 63.78 6.32 63.95 6.49 ;
      RECT 63.78 7.8 63.95 7.97 ;
      RECT 63.43 0.1 63.6 0.27 ;
      RECT 63.43 8.61 63.6 8.78 ;
      RECT 63.41 2.76 63.58 2.93 ;
      RECT 63.41 5.95 63.58 6.12 ;
      RECT 62.73 0.105 62.9 0.275 ;
      RECT 62.73 8.605 62.9 8.775 ;
      RECT 62.42 2.025 62.59 2.195 ;
      RECT 62.42 6.685 62.59 6.855 ;
      RECT 62.05 0.105 62.22 0.275 ;
      RECT 62.05 8.605 62.22 8.775 ;
      RECT 61.99 0.915 62.16 1.085 ;
      RECT 61.99 1.655 62.16 1.825 ;
      RECT 61.99 7.055 62.16 7.225 ;
      RECT 61.99 7.795 62.16 7.965 ;
      RECT 61.615 2.395 61.785 2.565 ;
      RECT 61.615 6.315 61.785 6.485 ;
      RECT 61.37 0.105 61.54 0.275 ;
      RECT 61.37 8.605 61.54 8.775 ;
      RECT 60.69 0.105 60.86 0.275 ;
      RECT 60.69 8.605 60.86 8.775 ;
      RECT 59.23 1.415 59.4 1.585 ;
      RECT 58.79 2.28 58.96 2.45 ;
      RECT 58.77 1.415 58.94 1.585 ;
      RECT 58.395 3.025 58.565 3.195 ;
      RECT 58.31 1.415 58.48 1.585 ;
      RECT 58.285 2.3 58.455 2.47 ;
      RECT 57.85 1.415 58.02 1.585 ;
      RECT 57.465 1.99 57.635 2.16 ;
      RECT 57.39 1.415 57.56 1.585 ;
      RECT 57.15 3.03 57.32 3.2 ;
      RECT 57.105 2.52 57.275 2.69 ;
      RECT 57.095 8.605 57.265 8.775 ;
      RECT 56.93 1.415 57.1 1.585 ;
      RECT 56.785 6.685 56.955 6.855 ;
      RECT 56.68 2.73 56.85 2.9 ;
      RECT 56.49 1.95 56.66 2.12 ;
      RECT 56.47 1.415 56.64 1.585 ;
      RECT 56.44 3.56 56.61 3.73 ;
      RECT 56.415 8.605 56.585 8.775 ;
      RECT 56.355 7.055 56.525 7.225 ;
      RECT 56.355 7.795 56.525 7.965 ;
      RECT 56.105 3 56.275 3.17 ;
      RECT 56.01 1.415 56.18 1.585 ;
      RECT 56.01 2.16 56.18 2.33 ;
      RECT 55.98 6.315 56.15 6.485 ;
      RECT 55.735 8.605 55.905 8.775 ;
      RECT 55.55 1.415 55.72 1.585 ;
      RECT 55.21 3.385 55.38 3.555 ;
      RECT 55.15 2.585 55.32 2.755 ;
      RECT 55.09 1.415 55.26 1.585 ;
      RECT 55.055 8.605 55.225 8.775 ;
      RECT 54.71 2.255 54.88 2.425 ;
      RECT 54.63 1.415 54.8 1.585 ;
      RECT 54.445 3.305 54.615 3.475 ;
      RECT 54.2 2.545 54.37 2.715 ;
      RECT 54.17 1.415 54.34 1.585 ;
      RECT 54.105 3.575 54.275 3.745 ;
      RECT 53.83 2.27 54 2.44 ;
      RECT 53.71 1.415 53.88 1.585 ;
      RECT 53.3 2.47 53.47 2.64 ;
      RECT 53.25 1.415 53.42 1.585 ;
      RECT 52.79 1.415 52.96 1.585 ;
      RECT 52.78 2.415 52.95 2.585 ;
      RECT 52.575 2.015 52.745 2.185 ;
      RECT 52.575 3.595 52.745 3.765 ;
      RECT 52.33 1.415 52.5 1.585 ;
      RECT 52.265 2.56 52.435 2.73 ;
      RECT 51.87 1.415 52.04 1.585 ;
      RECT 51.855 2.785 52.025 2.955 ;
      RECT 51.41 1.415 51.58 1.585 ;
      RECT 51.145 3.085 51.315 3.255 ;
      RECT 51 1.995 51.17 2.165 ;
      RECT 50.95 1.415 51.12 1.585 ;
      RECT 49.51 7.8 49.68 7.97 ;
      RECT 49.16 0.1 49.33 0.27 ;
      RECT 49.16 8.61 49.33 8.78 ;
      RECT 49.14 2.76 49.31 2.93 ;
      RECT 49.14 5.95 49.31 6.12 ;
      RECT 48.52 0.91 48.69 1.08 ;
      RECT 48.52 2.39 48.69 2.56 ;
      RECT 48.52 6.32 48.69 6.49 ;
      RECT 48.52 7.8 48.69 7.97 ;
      RECT 48.17 0.1 48.34 0.27 ;
      RECT 48.17 8.61 48.34 8.78 ;
      RECT 48.15 2.76 48.32 2.93 ;
      RECT 48.15 5.95 48.32 6.12 ;
      RECT 47.47 0.105 47.64 0.275 ;
      RECT 47.47 8.605 47.64 8.775 ;
      RECT 47.16 2.025 47.33 2.195 ;
      RECT 47.16 6.685 47.33 6.855 ;
      RECT 46.79 0.105 46.96 0.275 ;
      RECT 46.79 8.605 46.96 8.775 ;
      RECT 46.73 0.915 46.9 1.085 ;
      RECT 46.73 1.655 46.9 1.825 ;
      RECT 46.73 7.055 46.9 7.225 ;
      RECT 46.73 7.795 46.9 7.965 ;
      RECT 46.355 2.395 46.525 2.565 ;
      RECT 46.355 6.315 46.525 6.485 ;
      RECT 46.11 0.105 46.28 0.275 ;
      RECT 46.11 8.605 46.28 8.775 ;
      RECT 45.43 0.105 45.6 0.275 ;
      RECT 45.43 8.605 45.6 8.775 ;
      RECT 43.97 1.415 44.14 1.585 ;
      RECT 43.53 2.28 43.7 2.45 ;
      RECT 43.51 1.415 43.68 1.585 ;
      RECT 43.135 3.025 43.305 3.195 ;
      RECT 43.05 1.415 43.22 1.585 ;
      RECT 43.025 2.3 43.195 2.47 ;
      RECT 42.59 1.415 42.76 1.585 ;
      RECT 42.205 1.99 42.375 2.16 ;
      RECT 42.13 1.415 42.3 1.585 ;
      RECT 41.89 3.03 42.06 3.2 ;
      RECT 41.845 2.52 42.015 2.69 ;
      RECT 41.835 8.605 42.005 8.775 ;
      RECT 41.67 1.415 41.84 1.585 ;
      RECT 41.525 6.685 41.695 6.855 ;
      RECT 41.42 2.73 41.59 2.9 ;
      RECT 41.23 1.95 41.4 2.12 ;
      RECT 41.21 1.415 41.38 1.585 ;
      RECT 41.18 3.56 41.35 3.73 ;
      RECT 41.155 8.605 41.325 8.775 ;
      RECT 41.095 7.055 41.265 7.225 ;
      RECT 41.095 7.795 41.265 7.965 ;
      RECT 40.845 3 41.015 3.17 ;
      RECT 40.75 1.415 40.92 1.585 ;
      RECT 40.75 2.16 40.92 2.33 ;
      RECT 40.72 6.315 40.89 6.485 ;
      RECT 40.475 8.605 40.645 8.775 ;
      RECT 40.29 1.415 40.46 1.585 ;
      RECT 39.95 3.385 40.12 3.555 ;
      RECT 39.89 2.585 40.06 2.755 ;
      RECT 39.83 1.415 40 1.585 ;
      RECT 39.795 8.605 39.965 8.775 ;
      RECT 39.45 2.255 39.62 2.425 ;
      RECT 39.37 1.415 39.54 1.585 ;
      RECT 39.185 3.305 39.355 3.475 ;
      RECT 38.94 2.545 39.11 2.715 ;
      RECT 38.91 1.415 39.08 1.585 ;
      RECT 38.845 3.575 39.015 3.745 ;
      RECT 38.57 2.27 38.74 2.44 ;
      RECT 38.45 1.415 38.62 1.585 ;
      RECT 38.04 2.47 38.21 2.64 ;
      RECT 37.99 1.415 38.16 1.585 ;
      RECT 37.53 1.415 37.7 1.585 ;
      RECT 37.52 2.415 37.69 2.585 ;
      RECT 37.315 2.015 37.485 2.185 ;
      RECT 37.315 3.595 37.485 3.765 ;
      RECT 37.07 1.415 37.24 1.585 ;
      RECT 37.005 2.56 37.175 2.73 ;
      RECT 36.61 1.415 36.78 1.585 ;
      RECT 36.595 2.785 36.765 2.955 ;
      RECT 36.15 1.415 36.32 1.585 ;
      RECT 35.885 3.085 36.055 3.255 ;
      RECT 35.74 1.995 35.91 2.165 ;
      RECT 35.69 1.415 35.86 1.585 ;
      RECT 34.25 7.8 34.42 7.97 ;
      RECT 33.9 0.1 34.07 0.27 ;
      RECT 33.9 8.61 34.07 8.78 ;
      RECT 33.88 2.76 34.05 2.93 ;
      RECT 33.88 5.95 34.05 6.12 ;
      RECT 33.26 0.91 33.43 1.08 ;
      RECT 33.26 2.39 33.43 2.56 ;
      RECT 33.26 6.32 33.43 6.49 ;
      RECT 33.26 7.8 33.43 7.97 ;
      RECT 32.91 0.1 33.08 0.27 ;
      RECT 32.91 8.61 33.08 8.78 ;
      RECT 32.89 2.76 33.06 2.93 ;
      RECT 32.89 5.95 33.06 6.12 ;
      RECT 32.21 0.105 32.38 0.275 ;
      RECT 32.21 8.605 32.38 8.775 ;
      RECT 31.9 2.025 32.07 2.195 ;
      RECT 31.9 6.685 32.07 6.855 ;
      RECT 31.53 0.105 31.7 0.275 ;
      RECT 31.53 8.605 31.7 8.775 ;
      RECT 31.47 0.915 31.64 1.085 ;
      RECT 31.47 1.655 31.64 1.825 ;
      RECT 31.47 7.055 31.64 7.225 ;
      RECT 31.47 7.795 31.64 7.965 ;
      RECT 31.095 2.395 31.265 2.565 ;
      RECT 31.095 6.315 31.265 6.485 ;
      RECT 30.85 0.105 31.02 0.275 ;
      RECT 30.85 8.605 31.02 8.775 ;
      RECT 30.17 0.105 30.34 0.275 ;
      RECT 30.17 8.605 30.34 8.775 ;
      RECT 28.71 1.415 28.88 1.585 ;
      RECT 28.27 2.28 28.44 2.45 ;
      RECT 28.25 1.415 28.42 1.585 ;
      RECT 27.875 3.025 28.045 3.195 ;
      RECT 27.79 1.415 27.96 1.585 ;
      RECT 27.765 2.3 27.935 2.47 ;
      RECT 27.33 1.415 27.5 1.585 ;
      RECT 26.945 1.99 27.115 2.16 ;
      RECT 26.87 1.415 27.04 1.585 ;
      RECT 26.63 3.03 26.8 3.2 ;
      RECT 26.585 2.52 26.755 2.69 ;
      RECT 26.575 8.605 26.745 8.775 ;
      RECT 26.41 1.415 26.58 1.585 ;
      RECT 26.265 6.685 26.435 6.855 ;
      RECT 26.16 2.73 26.33 2.9 ;
      RECT 25.97 1.95 26.14 2.12 ;
      RECT 25.95 1.415 26.12 1.585 ;
      RECT 25.92 3.56 26.09 3.73 ;
      RECT 25.895 8.605 26.065 8.775 ;
      RECT 25.835 7.055 26.005 7.225 ;
      RECT 25.835 7.795 26.005 7.965 ;
      RECT 25.585 3 25.755 3.17 ;
      RECT 25.49 1.415 25.66 1.585 ;
      RECT 25.49 2.16 25.66 2.33 ;
      RECT 25.46 6.315 25.63 6.485 ;
      RECT 25.215 8.605 25.385 8.775 ;
      RECT 25.03 1.415 25.2 1.585 ;
      RECT 24.69 3.385 24.86 3.555 ;
      RECT 24.63 2.585 24.8 2.755 ;
      RECT 24.57 1.415 24.74 1.585 ;
      RECT 24.535 8.605 24.705 8.775 ;
      RECT 24.19 2.255 24.36 2.425 ;
      RECT 24.11 1.415 24.28 1.585 ;
      RECT 23.925 3.305 24.095 3.475 ;
      RECT 23.68 2.545 23.85 2.715 ;
      RECT 23.65 1.415 23.82 1.585 ;
      RECT 23.585 3.575 23.755 3.745 ;
      RECT 23.31 2.27 23.48 2.44 ;
      RECT 23.19 1.415 23.36 1.585 ;
      RECT 22.78 2.47 22.95 2.64 ;
      RECT 22.73 1.415 22.9 1.585 ;
      RECT 22.27 1.415 22.44 1.585 ;
      RECT 22.26 2.415 22.43 2.585 ;
      RECT 22.055 2.015 22.225 2.185 ;
      RECT 22.055 3.595 22.225 3.765 ;
      RECT 21.81 1.415 21.98 1.585 ;
      RECT 21.745 2.56 21.915 2.73 ;
      RECT 21.35 1.415 21.52 1.585 ;
      RECT 21.335 2.785 21.505 2.955 ;
      RECT 20.89 1.415 21.06 1.585 ;
      RECT 20.625 3.085 20.795 3.255 ;
      RECT 20.48 1.995 20.65 2.165 ;
      RECT 20.43 1.415 20.6 1.585 ;
      RECT 18.99 7.8 19.16 7.97 ;
      RECT 18.64 0.1 18.81 0.27 ;
      RECT 18.64 8.61 18.81 8.78 ;
      RECT 18.62 2.76 18.79 2.93 ;
      RECT 18.62 5.95 18.79 6.12 ;
      RECT 18 0.91 18.17 1.08 ;
      RECT 18 2.39 18.17 2.56 ;
      RECT 18 6.32 18.17 6.49 ;
      RECT 18 7.8 18.17 7.97 ;
      RECT 17.65 0.1 17.82 0.27 ;
      RECT 17.65 8.61 17.82 8.78 ;
      RECT 17.63 2.76 17.8 2.93 ;
      RECT 17.63 5.95 17.8 6.12 ;
      RECT 16.95 0.105 17.12 0.275 ;
      RECT 16.95 8.605 17.12 8.775 ;
      RECT 16.64 2.025 16.81 2.195 ;
      RECT 16.64 6.685 16.81 6.855 ;
      RECT 16.27 0.105 16.44 0.275 ;
      RECT 16.27 8.605 16.44 8.775 ;
      RECT 16.21 0.915 16.38 1.085 ;
      RECT 16.21 1.655 16.38 1.825 ;
      RECT 16.21 7.055 16.38 7.225 ;
      RECT 16.21 7.795 16.38 7.965 ;
      RECT 15.835 2.395 16.005 2.565 ;
      RECT 15.835 6.315 16.005 6.485 ;
      RECT 15.59 0.105 15.76 0.275 ;
      RECT 15.59 8.605 15.76 8.775 ;
      RECT 14.91 0.105 15.08 0.275 ;
      RECT 14.91 8.605 15.08 8.775 ;
      RECT 13.45 1.415 13.62 1.585 ;
      RECT 13.01 2.28 13.18 2.45 ;
      RECT 12.99 1.415 13.16 1.585 ;
      RECT 12.615 3.025 12.785 3.195 ;
      RECT 12.53 1.415 12.7 1.585 ;
      RECT 12.505 2.3 12.675 2.47 ;
      RECT 12.07 1.415 12.24 1.585 ;
      RECT 11.685 1.99 11.855 2.16 ;
      RECT 11.61 1.415 11.78 1.585 ;
      RECT 11.37 3.03 11.54 3.2 ;
      RECT 11.325 2.52 11.495 2.69 ;
      RECT 11.315 8.605 11.485 8.775 ;
      RECT 11.15 1.415 11.32 1.585 ;
      RECT 11.005 6.685 11.175 6.855 ;
      RECT 10.9 2.73 11.07 2.9 ;
      RECT 10.71 1.95 10.88 2.12 ;
      RECT 10.69 1.415 10.86 1.585 ;
      RECT 10.66 3.56 10.83 3.73 ;
      RECT 10.635 8.605 10.805 8.775 ;
      RECT 10.575 7.055 10.745 7.225 ;
      RECT 10.575 7.795 10.745 7.965 ;
      RECT 10.325 3 10.495 3.17 ;
      RECT 10.23 1.415 10.4 1.585 ;
      RECT 10.23 2.16 10.4 2.33 ;
      RECT 10.2 6.315 10.37 6.485 ;
      RECT 9.955 8.605 10.125 8.775 ;
      RECT 9.77 1.415 9.94 1.585 ;
      RECT 9.43 3.385 9.6 3.555 ;
      RECT 9.37 2.585 9.54 2.755 ;
      RECT 9.31 1.415 9.48 1.585 ;
      RECT 9.275 8.605 9.445 8.775 ;
      RECT 8.93 2.255 9.1 2.425 ;
      RECT 8.85 1.415 9.02 1.585 ;
      RECT 8.665 3.305 8.835 3.475 ;
      RECT 8.42 2.545 8.59 2.715 ;
      RECT 8.39 1.415 8.56 1.585 ;
      RECT 8.325 3.575 8.495 3.745 ;
      RECT 8.05 2.27 8.22 2.44 ;
      RECT 7.93 1.415 8.1 1.585 ;
      RECT 7.52 2.47 7.69 2.64 ;
      RECT 7.47 1.415 7.64 1.585 ;
      RECT 7.01 1.415 7.18 1.585 ;
      RECT 7 2.415 7.17 2.585 ;
      RECT 6.795 2.015 6.965 2.185 ;
      RECT 6.795 3.595 6.965 3.765 ;
      RECT 6.55 1.415 6.72 1.585 ;
      RECT 6.485 2.56 6.655 2.73 ;
      RECT 6.09 1.415 6.26 1.585 ;
      RECT 6.075 2.785 6.245 2.955 ;
      RECT 5.63 1.415 5.8 1.585 ;
      RECT 5.365 3.085 5.535 3.255 ;
      RECT 5.22 1.995 5.39 2.165 ;
      RECT 5.17 1.415 5.34 1.585 ;
      RECT 3.82 8.605 3.99 8.775 ;
      RECT 3.14 8.605 3.31 8.775 ;
      RECT 3.08 7.055 3.25 7.225 ;
      RECT 3.08 7.795 3.25 7.965 ;
      RECT 2.705 6.315 2.875 6.485 ;
      RECT 2.46 8.605 2.63 8.775 ;
      RECT 1.78 8.605 1.95 8.775 ;
    LAYER li1 ;
      RECT 74.035 0 74.205 2.085 ;
      RECT 73.095 0 73.265 2.085 ;
      RECT 72.135 0 72.305 2.085 ;
      RECT 70.215 0 70.385 2.085 ;
      RECT 69.255 0 69.425 2.085 ;
      RECT 67.335 0 67.505 2.085 ;
      RECT 58.775 0 58.945 2.085 ;
      RECT 57.835 0 58.005 2.085 ;
      RECT 56.875 0 57.045 2.085 ;
      RECT 54.955 0 55.125 2.085 ;
      RECT 53.995 0 54.165 2.085 ;
      RECT 52.075 0 52.245 2.085 ;
      RECT 43.515 0 43.685 2.085 ;
      RECT 42.575 0 42.745 2.085 ;
      RECT 41.615 0 41.785 2.085 ;
      RECT 39.695 0 39.865 2.085 ;
      RECT 38.735 0 38.905 2.085 ;
      RECT 36.815 0 36.985 2.085 ;
      RECT 28.255 0 28.425 2.085 ;
      RECT 27.315 0 27.485 2.085 ;
      RECT 26.355 0 26.525 2.085 ;
      RECT 24.435 0 24.605 2.085 ;
      RECT 23.475 0 23.645 2.085 ;
      RECT 21.555 0 21.725 2.085 ;
      RECT 12.995 0 13.165 2.085 ;
      RECT 12.055 0 12.225 2.085 ;
      RECT 11.095 0 11.265 2.085 ;
      RECT 9.175 0 9.345 2.085 ;
      RECT 8.215 0 8.385 2.085 ;
      RECT 6.295 0 6.465 2.085 ;
      RECT 71.09 0 71.285 1.595 ;
      RECT 67.335 0 67.61 1.595 ;
      RECT 55.83 0 56.025 1.595 ;
      RECT 52.075 0 52.35 1.595 ;
      RECT 40.57 0 40.765 1.595 ;
      RECT 36.815 0 37.09 1.595 ;
      RECT 25.31 0 25.505 1.595 ;
      RECT 21.555 0 21.83 1.595 ;
      RECT 10.05 0 10.245 1.595 ;
      RECT 6.295 0 6.57 1.595 ;
      RECT 66.065 0 74.805 1.585 ;
      RECT 50.805 0 59.545 1.585 ;
      RECT 35.545 0 44.285 1.585 ;
      RECT 20.285 0 29.025 1.585 ;
      RECT 5.025 0 13.765 1.585 ;
      RECT 75.87 0 76.04 0.935 ;
      RECT 60.61 0 60.78 0.935 ;
      RECT 45.35 0 45.52 0.935 ;
      RECT 30.09 0 30.26 0.935 ;
      RECT 14.83 0 15 0.935 ;
      RECT 79.6 0 79.77 0.93 ;
      RECT 78.61 0 78.78 0.93 ;
      RECT 64.34 0 64.51 0.93 ;
      RECT 63.35 0 63.52 0.93 ;
      RECT 49.08 0 49.25 0.93 ;
      RECT 48.09 0 48.26 0.93 ;
      RECT 33.82 0 33.99 0.93 ;
      RECT 32.83 0 33 0.93 ;
      RECT 18.56 0 18.73 0.93 ;
      RECT 17.57 0 17.74 0.93 ;
      RECT 80.395 0 80.575 0.305 ;
      RECT 65.135 0 78.445 0.305 ;
      RECT 49.875 0 63.185 0.305 ;
      RECT 34.615 0 47.925 0.305 ;
      RECT 19.355 0 32.665 0.305 ;
      RECT 1.48 0 17.405 0.305 ;
      RECT 1.48 0 80.575 0.3 ;
      RECT 1.48 8.58 80.575 8.88 ;
      RECT 80.395 8.575 80.575 8.88 ;
      RECT 79.6 7.95 79.77 8.88 ;
      RECT 78.61 7.95 78.78 8.88 ;
      RECT 65.135 8.575 78.445 8.88 ;
      RECT 64.34 7.95 64.51 8.88 ;
      RECT 63.35 7.95 63.52 8.88 ;
      RECT 49.875 8.575 63.185 8.88 ;
      RECT 49.08 7.95 49.25 8.88 ;
      RECT 48.09 7.95 48.26 8.88 ;
      RECT 34.615 8.575 47.925 8.88 ;
      RECT 33.82 7.95 33.99 8.88 ;
      RECT 32.83 7.95 33 8.88 ;
      RECT 19.355 8.575 32.665 8.88 ;
      RECT 18.56 7.95 18.73 8.88 ;
      RECT 17.57 7.95 17.74 8.88 ;
      RECT 1.48 8.575 17.405 8.88 ;
      RECT 75.87 7.945 76.04 8.88 ;
      RECT 70.235 7.945 70.405 8.88 ;
      RECT 60.61 7.945 60.78 8.88 ;
      RECT 54.975 7.945 55.145 8.88 ;
      RECT 45.35 7.945 45.52 8.88 ;
      RECT 39.715 7.945 39.885 8.88 ;
      RECT 30.09 7.945 30.26 8.88 ;
      RECT 24.455 7.945 24.625 8.88 ;
      RECT 14.83 7.945 15 8.88 ;
      RECT 9.195 7.945 9.365 8.88 ;
      RECT 1.7 7.945 1.87 8.88 ;
      RECT 80.03 5.02 80.2 6.49 ;
      RECT 80.03 6.315 80.205 6.485 ;
      RECT 79.66 1.74 79.83 2.93 ;
      RECT 79.66 1.74 80.13 1.91 ;
      RECT 79.66 6.97 80.13 7.14 ;
      RECT 79.66 5.95 79.83 7.14 ;
      RECT 78.67 1.74 78.84 2.93 ;
      RECT 78.67 1.74 79.14 1.91 ;
      RECT 78.67 6.97 79.14 7.14 ;
      RECT 78.67 5.95 78.84 7.14 ;
      RECT 76.82 2.635 76.99 3.865 ;
      RECT 76.875 0.855 77.045 2.805 ;
      RECT 76.82 0.575 76.99 1.025 ;
      RECT 76.82 7.855 76.99 8.305 ;
      RECT 76.875 6.075 77.045 8.025 ;
      RECT 76.82 5.015 76.99 6.245 ;
      RECT 76.3 0.575 76.47 3.865 ;
      RECT 76.3 2.075 76.705 2.405 ;
      RECT 76.3 1.235 76.705 1.565 ;
      RECT 76.3 5.015 76.47 8.305 ;
      RECT 76.3 7.315 76.705 7.645 ;
      RECT 76.3 6.475 76.705 6.805 ;
      RECT 74.225 3.126 74.23 3.298 ;
      RECT 74.22 3.119 74.225 3.388 ;
      RECT 74.215 3.113 74.22 3.407 ;
      RECT 74.195 3.107 74.215 3.417 ;
      RECT 74.18 3.102 74.195 3.425 ;
      RECT 74.143 3.096 74.18 3.423 ;
      RECT 74.057 3.082 74.143 3.419 ;
      RECT 73.971 3.064 74.057 3.414 ;
      RECT 73.885 3.045 73.971 3.408 ;
      RECT 73.855 3.033 73.885 3.404 ;
      RECT 73.835 3.027 73.855 3.403 ;
      RECT 73.77 3.025 73.835 3.401 ;
      RECT 73.755 3.025 73.77 3.393 ;
      RECT 73.74 3.025 73.755 3.38 ;
      RECT 73.735 3.025 73.74 3.37 ;
      RECT 73.72 3.025 73.735 3.348 ;
      RECT 73.705 3.025 73.72 3.315 ;
      RECT 73.7 3.025 73.705 3.293 ;
      RECT 73.69 3.025 73.7 3.275 ;
      RECT 73.675 3.025 73.69 3.253 ;
      RECT 73.655 3.025 73.675 3.215 ;
      RECT 74.005 2.31 74.04 2.749 ;
      RECT 74.005 2.31 74.045 2.748 ;
      RECT 73.95 2.37 74.045 2.747 ;
      RECT 73.815 2.542 74.045 2.746 ;
      RECT 73.925 2.42 74.045 2.746 ;
      RECT 73.815 2.542 74.07 2.736 ;
      RECT 73.87 2.487 74.15 2.653 ;
      RECT 74.045 2.281 74.05 2.744 ;
      RECT 73.9 2.457 74.19 2.53 ;
      RECT 73.915 2.44 74.045 2.746 ;
      RECT 74.05 2.28 74.22 2.468 ;
      RECT 74.04 2.283 74.22 2.468 ;
      RECT 73.545 2.16 73.715 2.47 ;
      RECT 73.545 2.16 73.72 2.443 ;
      RECT 73.545 2.16 73.725 2.42 ;
      RECT 73.545 2.16 73.735 2.37 ;
      RECT 73.54 2.265 73.735 2.34 ;
      RECT 73.575 1.835 73.745 2.313 ;
      RECT 73.575 1.835 73.76 2.234 ;
      RECT 73.565 2.045 73.76 2.234 ;
      RECT 73.575 1.845 73.77 2.149 ;
      RECT 73.505 2.587 73.51 2.79 ;
      RECT 73.495 2.575 73.505 2.9 ;
      RECT 73.47 2.575 73.495 2.94 ;
      RECT 73.39 2.575 73.47 3.025 ;
      RECT 73.38 2.575 73.39 3.095 ;
      RECT 73.355 2.575 73.38 3.118 ;
      RECT 73.335 2.575 73.355 3.153 ;
      RECT 73.29 2.585 73.335 3.196 ;
      RECT 73.28 2.597 73.29 3.233 ;
      RECT 73.26 2.611 73.28 3.253 ;
      RECT 73.25 2.629 73.26 3.269 ;
      RECT 73.235 2.655 73.25 3.279 ;
      RECT 73.22 2.696 73.235 3.293 ;
      RECT 73.21 2.731 73.22 3.303 ;
      RECT 73.205 2.747 73.21 3.308 ;
      RECT 73.195 2.762 73.205 3.313 ;
      RECT 73.175 2.805 73.195 3.323 ;
      RECT 73.155 2.842 73.175 3.336 ;
      RECT 73.12 2.865 73.155 3.354 ;
      RECT 73.11 2.879 73.12 3.37 ;
      RECT 73.09 2.889 73.11 3.38 ;
      RECT 73.085 2.898 73.09 3.388 ;
      RECT 73.075 2.905 73.085 3.395 ;
      RECT 73.065 2.912 73.075 3.403 ;
      RECT 73.05 2.922 73.065 3.411 ;
      RECT 73.04 2.936 73.05 3.421 ;
      RECT 73.03 2.948 73.04 3.433 ;
      RECT 73.015 2.97 73.03 3.446 ;
      RECT 73.005 2.992 73.015 3.457 ;
      RECT 72.995 3.012 73.005 3.466 ;
      RECT 72.99 3.027 72.995 3.473 ;
      RECT 72.96 3.06 72.99 3.487 ;
      RECT 72.95 3.095 72.96 3.502 ;
      RECT 72.945 3.102 72.95 3.508 ;
      RECT 72.925 3.117 72.945 3.515 ;
      RECT 72.92 3.132 72.925 3.523 ;
      RECT 72.915 3.141 72.92 3.528 ;
      RECT 72.9 3.147 72.915 3.535 ;
      RECT 72.895 3.153 72.9 3.543 ;
      RECT 72.89 3.157 72.895 3.55 ;
      RECT 72.885 3.161 72.89 3.56 ;
      RECT 72.875 3.166 72.885 3.57 ;
      RECT 72.855 3.177 72.875 3.598 ;
      RECT 72.84 3.189 72.855 3.625 ;
      RECT 72.82 3.202 72.84 3.65 ;
      RECT 72.8 3.217 72.82 3.674 ;
      RECT 72.785 3.232 72.8 3.689 ;
      RECT 72.78 3.243 72.785 3.698 ;
      RECT 72.715 3.288 72.78 3.708 ;
      RECT 72.68 3.347 72.715 3.721 ;
      RECT 72.675 3.37 72.68 3.727 ;
      RECT 72.67 3.377 72.675 3.729 ;
      RECT 72.655 3.387 72.67 3.732 ;
      RECT 72.625 3.412 72.655 3.736 ;
      RECT 72.62 3.43 72.625 3.74 ;
      RECT 72.615 3.437 72.62 3.741 ;
      RECT 72.595 3.445 72.615 3.745 ;
      RECT 72.585 3.452 72.595 3.749 ;
      RECT 72.541 3.463 72.585 3.756 ;
      RECT 72.455 3.491 72.541 3.772 ;
      RECT 72.395 3.515 72.455 3.79 ;
      RECT 72.35 3.525 72.395 3.804 ;
      RECT 72.291 3.533 72.35 3.818 ;
      RECT 72.205 3.54 72.291 3.837 ;
      RECT 72.18 3.545 72.205 3.852 ;
      RECT 72.1 3.548 72.18 3.855 ;
      RECT 72.02 3.552 72.1 3.842 ;
      RECT 72.011 3.555 72.02 3.827 ;
      RECT 71.925 3.555 72.011 3.812 ;
      RECT 71.865 3.557 71.925 3.789 ;
      RECT 71.861 3.56 71.865 3.779 ;
      RECT 71.775 3.56 71.861 3.764 ;
      RECT 71.7 3.56 71.775 3.74 ;
      RECT 73.015 2.569 73.025 2.745 ;
      RECT 72.97 2.536 73.015 2.745 ;
      RECT 72.925 2.487 72.97 2.745 ;
      RECT 72.895 2.457 72.925 2.746 ;
      RECT 72.89 2.44 72.895 2.747 ;
      RECT 72.865 2.42 72.89 2.748 ;
      RECT 72.85 2.395 72.865 2.749 ;
      RECT 72.845 2.382 72.85 2.75 ;
      RECT 72.84 2.376 72.845 2.748 ;
      RECT 72.835 2.368 72.84 2.742 ;
      RECT 72.81 2.36 72.835 2.722 ;
      RECT 72.79 2.349 72.81 2.693 ;
      RECT 72.76 2.334 72.79 2.664 ;
      RECT 72.74 2.32 72.76 2.636 ;
      RECT 72.73 2.314 72.74 2.615 ;
      RECT 72.725 2.311 72.73 2.598 ;
      RECT 72.72 2.308 72.725 2.583 ;
      RECT 72.705 2.303 72.72 2.548 ;
      RECT 72.7 2.299 72.705 2.515 ;
      RECT 72.68 2.294 72.7 2.491 ;
      RECT 72.65 2.286 72.68 2.456 ;
      RECT 72.635 2.28 72.65 2.433 ;
      RECT 72.595 2.273 72.635 2.418 ;
      RECT 72.57 2.265 72.595 2.398 ;
      RECT 72.55 2.26 72.57 2.388 ;
      RECT 72.515 2.254 72.55 2.383 ;
      RECT 72.47 2.245 72.515 2.382 ;
      RECT 72.44 2.241 72.47 2.384 ;
      RECT 72.355 2.249 72.44 2.388 ;
      RECT 72.285 2.26 72.355 2.41 ;
      RECT 72.272 2.266 72.285 2.433 ;
      RECT 72.186 2.273 72.272 2.455 ;
      RECT 72.1 2.285 72.186 2.492 ;
      RECT 72.1 2.662 72.11 2.9 ;
      RECT 72.095 2.291 72.1 2.515 ;
      RECT 72.09 2.547 72.1 2.9 ;
      RECT 72.09 2.292 72.095 2.52 ;
      RECT 72.085 2.293 72.09 2.9 ;
      RECT 72.061 2.295 72.085 2.901 ;
      RECT 71.975 2.303 72.061 2.903 ;
      RECT 71.955 2.317 71.975 2.906 ;
      RECT 71.95 2.345 71.955 2.907 ;
      RECT 71.945 2.357 71.95 2.908 ;
      RECT 71.94 2.372 71.945 2.909 ;
      RECT 71.93 2.402 71.94 2.91 ;
      RECT 71.925 2.44 71.93 2.908 ;
      RECT 71.92 2.46 71.925 2.903 ;
      RECT 71.905 2.495 71.92 2.888 ;
      RECT 71.895 2.547 71.905 2.868 ;
      RECT 71.89 2.577 71.895 2.856 ;
      RECT 71.875 2.59 71.89 2.839 ;
      RECT 71.85 2.594 71.875 2.806 ;
      RECT 71.835 2.592 71.85 2.783 ;
      RECT 71.82 2.591 71.835 2.78 ;
      RECT 71.76 2.589 71.82 2.778 ;
      RECT 71.75 2.587 71.76 2.773 ;
      RECT 71.71 2.586 71.75 2.77 ;
      RECT 71.64 2.583 71.71 2.768 ;
      RECT 71.585 2.581 71.64 2.763 ;
      RECT 71.515 2.575 71.585 2.758 ;
      RECT 71.506 2.575 71.515 2.755 ;
      RECT 71.42 2.575 71.506 2.75 ;
      RECT 71.415 2.575 71.42 2.745 ;
      RECT 72.72 1.81 72.895 2.16 ;
      RECT 72.72 1.825 72.905 2.158 ;
      RECT 72.695 1.775 72.84 2.155 ;
      RECT 72.675 1.776 72.84 2.148 ;
      RECT 72.665 1.777 72.85 2.143 ;
      RECT 72.635 1.778 72.85 2.13 ;
      RECT 72.585 1.779 72.85 2.106 ;
      RECT 72.58 1.781 72.85 2.091 ;
      RECT 72.58 1.847 72.91 2.085 ;
      RECT 72.56 1.788 72.865 2.065 ;
      RECT 72.55 1.797 72.875 1.92 ;
      RECT 72.56 1.792 72.875 2.065 ;
      RECT 72.58 1.782 72.865 2.091 ;
      RECT 72.165 3.107 72.335 3.395 ;
      RECT 72.16 3.125 72.345 3.39 ;
      RECT 72.125 3.133 72.41 3.31 ;
      RECT 72.125 3.133 72.496 3.3 ;
      RECT 72.125 3.133 72.55 3.246 ;
      RECT 72.41 3.03 72.58 3.214 ;
      RECT 72.125 3.185 72.585 3.202 ;
      RECT 72.11 3.155 72.58 3.198 ;
      RECT 72.37 3.037 72.41 3.349 ;
      RECT 72.25 3.074 72.58 3.214 ;
      RECT 72.345 3.049 72.37 3.375 ;
      RECT 72.335 3.056 72.58 3.214 ;
      RECT 72.466 2.52 72.535 2.779 ;
      RECT 72.466 2.575 72.54 2.778 ;
      RECT 72.38 2.575 72.54 2.777 ;
      RECT 72.375 2.575 72.545 2.77 ;
      RECT 72.365 2.52 72.535 2.765 ;
      RECT 71.745 1.819 71.92 2.12 ;
      RECT 71.73 1.807 71.745 2.105 ;
      RECT 71.7 1.806 71.73 2.058 ;
      RECT 71.7 1.824 71.925 2.053 ;
      RECT 71.685 1.808 71.745 2.018 ;
      RECT 71.68 1.83 71.935 1.918 ;
      RECT 71.68 1.813 71.831 1.918 ;
      RECT 71.68 1.815 71.835 1.918 ;
      RECT 71.685 1.811 71.831 2.018 ;
      RECT 71.79 3.047 71.795 3.395 ;
      RECT 71.78 3.037 71.79 3.401 ;
      RECT 71.745 3.027 71.78 3.403 ;
      RECT 71.707 3.022 71.745 3.407 ;
      RECT 71.621 3.015 71.707 3.414 ;
      RECT 71.535 3.005 71.621 3.424 ;
      RECT 71.49 3 71.535 3.432 ;
      RECT 71.486 3 71.49 3.436 ;
      RECT 71.4 3 71.486 3.443 ;
      RECT 71.385 3 71.4 3.443 ;
      RECT 71.375 2.998 71.385 3.415 ;
      RECT 71.365 2.994 71.375 3.358 ;
      RECT 71.345 2.988 71.365 3.29 ;
      RECT 71.34 2.984 71.345 3.238 ;
      RECT 71.33 2.983 71.34 3.205 ;
      RECT 71.28 2.981 71.33 3.19 ;
      RECT 71.255 2.979 71.28 3.185 ;
      RECT 71.212 2.977 71.255 3.181 ;
      RECT 71.126 2.973 71.212 3.169 ;
      RECT 71.04 2.968 71.126 3.153 ;
      RECT 71.01 2.965 71.04 3.14 ;
      RECT 70.985 2.964 71.01 3.128 ;
      RECT 70.98 2.964 70.985 3.118 ;
      RECT 70.94 2.963 70.98 3.11 ;
      RECT 70.925 2.962 70.94 3.103 ;
      RECT 70.875 2.961 70.925 3.095 ;
      RECT 70.873 2.96 70.875 3.09 ;
      RECT 70.787 2.958 70.873 3.09 ;
      RECT 70.701 2.953 70.787 3.09 ;
      RECT 70.615 2.949 70.701 3.09 ;
      RECT 70.566 2.945 70.615 3.088 ;
      RECT 70.48 2.942 70.566 3.083 ;
      RECT 70.457 2.939 70.48 3.079 ;
      RECT 70.371 2.936 70.457 3.074 ;
      RECT 70.285 2.932 70.371 3.065 ;
      RECT 70.26 2.925 70.285 3.06 ;
      RECT 70.2 2.89 70.26 3.057 ;
      RECT 70.18 2.815 70.2 3.054 ;
      RECT 70.175 2.757 70.18 3.053 ;
      RECT 70.15 2.697 70.175 3.052 ;
      RECT 70.075 2.575 70.15 3.048 ;
      RECT 70.065 2.575 70.075 3.04 ;
      RECT 70.05 2.575 70.065 3.03 ;
      RECT 70.035 2.575 70.05 3 ;
      RECT 70.02 2.575 70.035 2.945 ;
      RECT 70.005 2.575 70.02 2.883 ;
      RECT 69.98 2.575 70.005 2.808 ;
      RECT 69.975 2.575 69.98 2.758 ;
      RECT 71.32 2.12 71.34 2.429 ;
      RECT 71.306 2.122 71.355 2.426 ;
      RECT 71.306 2.127 71.375 2.417 ;
      RECT 71.22 2.125 71.355 2.411 ;
      RECT 71.22 2.133 71.41 2.394 ;
      RECT 71.185 2.135 71.41 2.393 ;
      RECT 71.155 2.143 71.41 2.384 ;
      RECT 71.145 2.148 71.43 2.37 ;
      RECT 71.185 2.138 71.43 2.37 ;
      RECT 71.185 2.141 71.44 2.358 ;
      RECT 71.155 2.143 71.45 2.345 ;
      RECT 71.155 2.147 71.46 2.288 ;
      RECT 71.145 2.152 71.465 2.203 ;
      RECT 71.306 2.12 71.34 2.426 ;
      RECT 71.185 7.855 71.355 8.305 ;
      RECT 71.24 6.075 71.41 8.025 ;
      RECT 71.185 5.015 71.355 6.245 ;
      RECT 70.745 2.223 70.75 2.435 ;
      RECT 70.62 2.22 70.635 2.435 ;
      RECT 70.085 2.25 70.155 2.435 ;
      RECT 69.97 2.25 70.005 2.43 ;
      RECT 71.091 2.552 71.11 2.746 ;
      RECT 71.005 2.507 71.091 2.747 ;
      RECT 70.995 2.46 71.005 2.749 ;
      RECT 70.99 2.44 70.995 2.75 ;
      RECT 70.97 2.405 70.99 2.751 ;
      RECT 70.955 2.355 70.97 2.752 ;
      RECT 70.935 2.292 70.955 2.753 ;
      RECT 70.925 2.255 70.935 2.754 ;
      RECT 70.91 2.244 70.925 2.755 ;
      RECT 70.905 2.236 70.91 2.753 ;
      RECT 70.895 2.235 70.905 2.745 ;
      RECT 70.865 2.232 70.895 2.724 ;
      RECT 70.79 2.227 70.865 2.669 ;
      RECT 70.775 2.223 70.79 2.615 ;
      RECT 70.765 2.223 70.775 2.51 ;
      RECT 70.75 2.223 70.765 2.443 ;
      RECT 70.735 2.223 70.745 2.433 ;
      RECT 70.68 2.222 70.735 2.43 ;
      RECT 70.635 2.22 70.68 2.433 ;
      RECT 70.607 2.22 70.62 2.436 ;
      RECT 70.521 2.224 70.607 2.438 ;
      RECT 70.435 2.23 70.521 2.443 ;
      RECT 70.415 2.234 70.435 2.445 ;
      RECT 70.413 2.235 70.415 2.444 ;
      RECT 70.327 2.237 70.413 2.443 ;
      RECT 70.241 2.242 70.327 2.44 ;
      RECT 70.155 2.247 70.241 2.437 ;
      RECT 70.005 2.25 70.085 2.433 ;
      RECT 70.665 5.015 70.835 8.305 ;
      RECT 70.665 7.315 71.07 7.645 ;
      RECT 70.665 6.475 71.07 6.805 ;
      RECT 70.781 3.225 70.83 3.559 ;
      RECT 70.781 3.225 70.835 3.558 ;
      RECT 70.695 3.225 70.835 3.557 ;
      RECT 70.47 3.333 70.84 3.555 ;
      RECT 70.695 3.225 70.865 3.548 ;
      RECT 70.665 3.237 70.87 3.539 ;
      RECT 70.65 3.255 70.875 3.536 ;
      RECT 70.465 3.339 70.875 3.463 ;
      RECT 70.46 3.346 70.875 3.423 ;
      RECT 70.475 3.312 70.875 3.536 ;
      RECT 70.636 3.258 70.84 3.555 ;
      RECT 70.55 3.278 70.875 3.536 ;
      RECT 70.65 3.252 70.87 3.539 ;
      RECT 70.42 2.576 70.61 2.77 ;
      RECT 70.415 2.578 70.61 2.769 ;
      RECT 70.41 2.582 70.625 2.766 ;
      RECT 70.425 2.575 70.625 2.766 ;
      RECT 70.41 2.685 70.63 2.761 ;
      RECT 69.705 3.185 69.796 3.483 ;
      RECT 69.7 3.187 69.875 3.478 ;
      RECT 69.705 3.185 69.875 3.478 ;
      RECT 69.7 3.191 69.895 3.476 ;
      RECT 69.7 3.246 69.935 3.475 ;
      RECT 69.7 3.281 69.95 3.469 ;
      RECT 69.7 3.315 69.96 3.459 ;
      RECT 69.69 3.195 69.895 3.31 ;
      RECT 69.69 3.215 69.91 3.31 ;
      RECT 69.69 3.198 69.9 3.31 ;
      RECT 69.915 1.966 69.92 2.028 ;
      RECT 69.91 1.888 69.915 2.051 ;
      RECT 69.905 1.845 69.91 2.062 ;
      RECT 69.9 1.835 69.905 2.074 ;
      RECT 69.895 1.835 69.9 2.083 ;
      RECT 69.87 1.835 69.895 2.115 ;
      RECT 69.865 1.835 69.87 2.148 ;
      RECT 69.85 1.835 69.865 2.173 ;
      RECT 69.84 1.835 69.85 2.2 ;
      RECT 69.835 1.835 69.84 2.213 ;
      RECT 69.83 1.835 69.835 2.228 ;
      RECT 69.82 1.835 69.83 2.243 ;
      RECT 69.815 1.835 69.82 2.263 ;
      RECT 69.79 1.835 69.815 2.298 ;
      RECT 69.745 1.835 69.79 2.343 ;
      RECT 69.735 1.835 69.745 2.356 ;
      RECT 69.65 1.92 69.735 2.363 ;
      RECT 69.615 2.042 69.65 2.372 ;
      RECT 69.61 2.082 69.615 2.376 ;
      RECT 69.59 2.105 69.61 2.378 ;
      RECT 69.585 2.135 69.59 2.381 ;
      RECT 69.575 2.147 69.585 2.382 ;
      RECT 69.53 2.17 69.575 2.387 ;
      RECT 69.49 2.2 69.53 2.395 ;
      RECT 69.455 2.212 69.49 2.401 ;
      RECT 69.45 2.217 69.455 2.405 ;
      RECT 69.38 2.227 69.45 2.412 ;
      RECT 69.34 2.237 69.38 2.422 ;
      RECT 69.32 2.242 69.34 2.428 ;
      RECT 69.31 2.246 69.32 2.433 ;
      RECT 69.305 2.249 69.31 2.436 ;
      RECT 69.295 2.25 69.305 2.437 ;
      RECT 69.27 2.252 69.295 2.441 ;
      RECT 69.26 2.257 69.27 2.444 ;
      RECT 69.215 2.265 69.26 2.445 ;
      RECT 69.09 2.27 69.215 2.445 ;
      RECT 69.645 2.567 69.665 2.749 ;
      RECT 69.596 2.552 69.645 2.748 ;
      RECT 69.51 2.567 69.665 2.746 ;
      RECT 69.495 2.567 69.665 2.745 ;
      RECT 69.46 2.545 69.63 2.73 ;
      RECT 69.53 3.565 69.545 3.774 ;
      RECT 69.53 3.573 69.55 3.773 ;
      RECT 69.475 3.573 69.55 3.772 ;
      RECT 69.455 3.577 69.555 3.77 ;
      RECT 69.435 3.527 69.475 3.769 ;
      RECT 69.38 3.585 69.56 3.767 ;
      RECT 69.345 3.542 69.475 3.765 ;
      RECT 69.341 3.545 69.53 3.764 ;
      RECT 69.255 3.553 69.53 3.762 ;
      RECT 69.255 3.597 69.565 3.755 ;
      RECT 69.245 3.69 69.565 3.753 ;
      RECT 69.255 3.609 69.57 3.738 ;
      RECT 69.255 3.63 69.585 3.708 ;
      RECT 69.255 3.657 69.59 3.678 ;
      RECT 69.38 3.535 69.475 3.767 ;
      RECT 69.01 2.58 69.015 3.118 ;
      RECT 68.815 2.91 68.82 3.105 ;
      RECT 67.115 2.575 67.13 2.955 ;
      RECT 69.18 2.575 69.185 2.745 ;
      RECT 69.175 2.575 69.18 2.755 ;
      RECT 69.17 2.575 69.175 2.768 ;
      RECT 69.145 2.575 69.17 2.81 ;
      RECT 69.12 2.575 69.145 2.883 ;
      RECT 69.105 2.575 69.12 2.935 ;
      RECT 69.1 2.575 69.105 2.965 ;
      RECT 69.075 2.575 69.1 3.005 ;
      RECT 69.06 2.575 69.075 3.06 ;
      RECT 69.055 2.575 69.06 3.093 ;
      RECT 69.03 2.575 69.055 3.113 ;
      RECT 69.015 2.575 69.03 3.119 ;
      RECT 68.945 2.61 69.01 3.115 ;
      RECT 68.895 2.665 68.945 3.11 ;
      RECT 68.885 2.697 68.895 3.108 ;
      RECT 68.88 2.722 68.885 3.108 ;
      RECT 68.86 2.795 68.88 3.108 ;
      RECT 68.85 2.875 68.86 3.107 ;
      RECT 68.835 2.905 68.85 3.107 ;
      RECT 68.82 2.91 68.835 3.106 ;
      RECT 68.76 2.912 68.815 3.103 ;
      RECT 68.73 2.917 68.76 3.099 ;
      RECT 68.728 2.92 68.73 3.098 ;
      RECT 68.642 2.922 68.728 3.095 ;
      RECT 68.556 2.928 68.642 3.089 ;
      RECT 68.47 2.933 68.556 3.083 ;
      RECT 68.397 2.938 68.47 3.084 ;
      RECT 68.311 2.944 68.397 3.092 ;
      RECT 68.225 2.95 68.311 3.101 ;
      RECT 68.205 2.954 68.225 3.106 ;
      RECT 68.158 2.956 68.205 3.109 ;
      RECT 68.072 2.961 68.158 3.115 ;
      RECT 67.986 2.966 68.072 3.124 ;
      RECT 67.9 2.972 67.986 3.132 ;
      RECT 67.815 2.97 67.9 3.141 ;
      RECT 67.811 2.965 67.815 3.145 ;
      RECT 67.725 2.96 67.811 3.137 ;
      RECT 67.661 2.951 67.725 3.125 ;
      RECT 67.575 2.942 67.661 3.112 ;
      RECT 67.551 2.935 67.575 3.103 ;
      RECT 67.465 2.929 67.551 3.09 ;
      RECT 67.425 2.922 67.465 3.076 ;
      RECT 67.42 2.912 67.425 3.072 ;
      RECT 67.41 2.9 67.42 3.071 ;
      RECT 67.39 2.87 67.41 3.068 ;
      RECT 67.335 2.79 67.39 3.062 ;
      RECT 67.315 2.709 67.335 3.057 ;
      RECT 67.295 2.667 67.315 3.053 ;
      RECT 67.27 2.62 67.295 3.047 ;
      RECT 67.265 2.595 67.27 3.044 ;
      RECT 67.23 2.575 67.265 3.039 ;
      RECT 67.221 2.575 67.23 3.032 ;
      RECT 67.135 2.575 67.221 3.002 ;
      RECT 67.13 2.575 67.135 2.965 ;
      RECT 67.095 2.575 67.115 2.887 ;
      RECT 67.09 2.617 67.095 2.852 ;
      RECT 67.085 2.692 67.09 2.808 ;
      RECT 68.535 2.497 68.71 2.745 ;
      RECT 68.535 2.497 68.715 2.743 ;
      RECT 68.53 2.529 68.715 2.703 ;
      RECT 68.56 2.47 68.73 2.69 ;
      RECT 68.525 2.547 68.73 2.623 ;
      RECT 67.835 2.01 68.005 2.185 ;
      RECT 67.835 2.01 68.177 2.177 ;
      RECT 67.835 2.01 68.26 2.171 ;
      RECT 67.835 2.01 68.295 2.167 ;
      RECT 67.835 2.01 68.315 2.166 ;
      RECT 67.835 2.01 68.401 2.162 ;
      RECT 68.295 1.835 68.465 2.157 ;
      RECT 67.87 1.942 68.495 2.155 ;
      RECT 67.86 1.997 68.5 2.153 ;
      RECT 67.835 2.033 68.51 2.148 ;
      RECT 67.835 2.06 68.515 2.078 ;
      RECT 67.9 1.885 68.475 2.155 ;
      RECT 68.091 1.87 68.475 2.155 ;
      RECT 67.925 1.873 68.475 2.155 ;
      RECT 68.005 1.871 68.091 2.182 ;
      RECT 68.091 1.868 68.47 2.155 ;
      RECT 68.275 1.845 68.47 2.155 ;
      RECT 68.177 1.866 68.47 2.155 ;
      RECT 68.26 1.86 68.275 2.168 ;
      RECT 68.41 3.225 68.415 3.425 ;
      RECT 67.875 3.29 67.92 3.425 ;
      RECT 68.445 3.225 68.465 3.398 ;
      RECT 68.415 3.225 68.445 3.413 ;
      RECT 68.35 3.225 68.41 3.45 ;
      RECT 68.335 3.225 68.35 3.48 ;
      RECT 68.32 3.225 68.335 3.493 ;
      RECT 68.3 3.225 68.32 3.508 ;
      RECT 68.295 3.225 68.3 3.517 ;
      RECT 68.285 3.229 68.295 3.522 ;
      RECT 68.27 3.239 68.285 3.533 ;
      RECT 68.245 3.255 68.27 3.543 ;
      RECT 68.235 3.269 68.245 3.545 ;
      RECT 68.215 3.281 68.235 3.542 ;
      RECT 68.185 3.302 68.215 3.536 ;
      RECT 68.175 3.314 68.185 3.531 ;
      RECT 68.165 3.312 68.175 3.528 ;
      RECT 68.15 3.311 68.165 3.523 ;
      RECT 68.145 3.31 68.15 3.518 ;
      RECT 68.11 3.308 68.145 3.508 ;
      RECT 68.09 3.305 68.11 3.49 ;
      RECT 68.08 3.303 68.09 3.485 ;
      RECT 68.07 3.302 68.08 3.48 ;
      RECT 68.035 3.3 68.07 3.468 ;
      RECT 67.98 3.296 68.035 3.448 ;
      RECT 67.97 3.294 67.98 3.433 ;
      RECT 67.965 3.294 67.97 3.428 ;
      RECT 67.92 3.292 67.965 3.425 ;
      RECT 67.825 3.29 67.875 3.429 ;
      RECT 67.815 3.291 67.825 3.434 ;
      RECT 67.755 3.298 67.815 3.448 ;
      RECT 67.73 3.306 67.755 3.468 ;
      RECT 67.72 3.31 67.73 3.48 ;
      RECT 67.715 3.311 67.72 3.485 ;
      RECT 67.7 3.313 67.715 3.488 ;
      RECT 67.685 3.315 67.7 3.493 ;
      RECT 67.68 3.315 67.685 3.496 ;
      RECT 67.635 3.32 67.68 3.507 ;
      RECT 67.63 3.324 67.635 3.519 ;
      RECT 67.605 3.32 67.63 3.523 ;
      RECT 67.595 3.316 67.605 3.527 ;
      RECT 67.585 3.315 67.595 3.531 ;
      RECT 67.57 3.305 67.585 3.537 ;
      RECT 67.565 3.293 67.57 3.541 ;
      RECT 67.56 3.29 67.565 3.542 ;
      RECT 67.555 3.287 67.56 3.544 ;
      RECT 67.54 3.275 67.555 3.543 ;
      RECT 67.525 3.257 67.54 3.54 ;
      RECT 67.505 3.236 67.525 3.533 ;
      RECT 67.44 3.225 67.505 3.505 ;
      RECT 67.436 3.225 67.44 3.484 ;
      RECT 67.35 3.225 67.436 3.454 ;
      RECT 67.335 3.225 67.35 3.41 ;
      RECT 67.91 2.325 67.915 2.56 ;
      RECT 67.04 2.241 67.045 2.445 ;
      RECT 67.62 2.27 67.625 2.425 ;
      RECT 67.54 2.25 67.545 2.425 ;
      RECT 68.21 2.392 68.225 2.745 ;
      RECT 68.136 2.377 68.21 2.745 ;
      RECT 68.05 2.36 68.136 2.745 ;
      RECT 68.04 2.35 68.05 2.743 ;
      RECT 68.035 2.348 68.04 2.738 ;
      RECT 68.02 2.346 68.035 2.724 ;
      RECT 67.95 2.338 68.02 2.664 ;
      RECT 67.93 2.329 67.95 2.598 ;
      RECT 67.925 2.326 67.93 2.578 ;
      RECT 67.915 2.325 67.925 2.568 ;
      RECT 67.905 2.325 67.91 2.552 ;
      RECT 67.895 2.324 67.905 2.542 ;
      RECT 67.885 2.322 67.895 2.53 ;
      RECT 67.87 2.319 67.885 2.51 ;
      RECT 67.86 2.317 67.87 2.495 ;
      RECT 67.84 2.314 67.86 2.483 ;
      RECT 67.835 2.312 67.84 2.473 ;
      RECT 67.81 2.31 67.835 2.46 ;
      RECT 67.78 2.305 67.81 2.445 ;
      RECT 67.7 2.296 67.78 2.436 ;
      RECT 67.655 2.285 67.7 2.429 ;
      RECT 67.635 2.276 67.655 2.426 ;
      RECT 67.625 2.271 67.635 2.425 ;
      RECT 67.58 2.265 67.62 2.425 ;
      RECT 67.565 2.257 67.58 2.425 ;
      RECT 67.545 2.252 67.565 2.425 ;
      RECT 67.525 2.249 67.54 2.425 ;
      RECT 67.442 2.248 67.525 2.424 ;
      RECT 67.356 2.247 67.442 2.42 ;
      RECT 67.27 2.245 67.356 2.417 ;
      RECT 67.217 2.244 67.27 2.419 ;
      RECT 67.131 2.243 67.217 2.428 ;
      RECT 67.045 2.242 67.131 2.44 ;
      RECT 67.025 2.241 67.04 2.448 ;
      RECT 66.945 2.24 67.025 2.46 ;
      RECT 66.92 2.24 66.945 2.473 ;
      RECT 66.895 2.24 66.92 2.488 ;
      RECT 66.89 2.24 66.895 2.51 ;
      RECT 66.885 2.24 66.89 2.528 ;
      RECT 66.88 2.24 66.885 2.545 ;
      RECT 66.875 2.24 66.88 2.558 ;
      RECT 66.87 2.24 66.875 2.568 ;
      RECT 66.83 2.24 66.87 2.653 ;
      RECT 66.815 2.24 66.83 2.738 ;
      RECT 66.805 2.241 66.815 2.75 ;
      RECT 66.77 2.246 66.805 2.755 ;
      RECT 66.73 2.255 66.77 2.755 ;
      RECT 66.715 2.265 66.73 2.755 ;
      RECT 66.71 2.275 66.715 2.755 ;
      RECT 66.69 2.302 66.71 2.755 ;
      RECT 66.64 2.385 66.69 2.755 ;
      RECT 66.635 2.447 66.64 2.755 ;
      RECT 66.625 2.46 66.635 2.755 ;
      RECT 66.615 2.482 66.625 2.755 ;
      RECT 66.605 2.507 66.615 2.75 ;
      RECT 66.6 2.545 66.605 2.743 ;
      RECT 66.59 2.655 66.6 2.738 ;
      RECT 67.985 3.576 68 3.835 ;
      RECT 67.985 3.591 68.005 3.834 ;
      RECT 67.901 3.591 68.005 3.832 ;
      RECT 67.901 3.605 68.01 3.831 ;
      RECT 67.815 3.647 68.015 3.828 ;
      RECT 67.81 3.59 68 3.823 ;
      RECT 67.81 3.661 68.02 3.82 ;
      RECT 67.805 3.692 68.02 3.818 ;
      RECT 67.81 3.689 68.035 3.808 ;
      RECT 67.805 3.735 68.05 3.793 ;
      RECT 67.805 3.763 68.055 3.778 ;
      RECT 67.815 3.565 67.985 3.828 ;
      RECT 67.575 2.575 67.745 2.745 ;
      RECT 67.54 2.575 67.745 2.74 ;
      RECT 67.53 2.575 67.745 2.733 ;
      RECT 67.525 2.56 67.695 2.73 ;
      RECT 66.355 3.097 66.62 3.54 ;
      RECT 66.35 3.068 66.565 3.538 ;
      RECT 66.345 3.222 66.625 3.533 ;
      RECT 66.35 3.117 66.625 3.533 ;
      RECT 66.35 3.128 66.635 3.52 ;
      RECT 66.35 3.075 66.595 3.538 ;
      RECT 66.355 3.062 66.565 3.54 ;
      RECT 66.355 3.06 66.515 3.54 ;
      RECT 66.456 3.052 66.515 3.54 ;
      RECT 66.37 3.053 66.515 3.54 ;
      RECT 66.456 3.051 66.505 3.54 ;
      RECT 66.26 1.866 66.435 2.165 ;
      RECT 66.31 1.828 66.435 2.165 ;
      RECT 66.295 1.83 66.521 2.157 ;
      RECT 66.295 1.833 66.56 2.144 ;
      RECT 66.295 1.834 66.57 2.13 ;
      RECT 66.25 1.885 66.57 2.12 ;
      RECT 66.295 1.835 66.575 2.115 ;
      RECT 66.25 2.045 66.58 2.105 ;
      RECT 66.235 1.905 66.575 2.045 ;
      RECT 66.23 1.921 66.575 1.985 ;
      RECT 66.275 1.845 66.575 2.115 ;
      RECT 66.31 1.826 66.396 2.165 ;
      RECT 64.77 5.02 64.94 6.49 ;
      RECT 64.77 6.315 64.945 6.485 ;
      RECT 64.4 1.74 64.57 2.93 ;
      RECT 64.4 1.74 64.87 1.91 ;
      RECT 64.4 6.97 64.87 7.14 ;
      RECT 64.4 5.95 64.57 7.14 ;
      RECT 63.41 1.74 63.58 2.93 ;
      RECT 63.41 1.74 63.88 1.91 ;
      RECT 63.41 6.97 63.88 7.14 ;
      RECT 63.41 5.95 63.58 7.14 ;
      RECT 61.56 2.635 61.73 3.865 ;
      RECT 61.615 0.855 61.785 2.805 ;
      RECT 61.56 0.575 61.73 1.025 ;
      RECT 61.56 7.855 61.73 8.305 ;
      RECT 61.615 6.075 61.785 8.025 ;
      RECT 61.56 5.015 61.73 6.245 ;
      RECT 61.04 0.575 61.21 3.865 ;
      RECT 61.04 2.075 61.445 2.405 ;
      RECT 61.04 1.235 61.445 1.565 ;
      RECT 61.04 5.015 61.21 8.305 ;
      RECT 61.04 7.315 61.445 7.645 ;
      RECT 61.04 6.475 61.445 6.805 ;
      RECT 58.965 3.126 58.97 3.298 ;
      RECT 58.96 3.119 58.965 3.388 ;
      RECT 58.955 3.113 58.96 3.407 ;
      RECT 58.935 3.107 58.955 3.417 ;
      RECT 58.92 3.102 58.935 3.425 ;
      RECT 58.883 3.096 58.92 3.423 ;
      RECT 58.797 3.082 58.883 3.419 ;
      RECT 58.711 3.064 58.797 3.414 ;
      RECT 58.625 3.045 58.711 3.408 ;
      RECT 58.595 3.033 58.625 3.404 ;
      RECT 58.575 3.027 58.595 3.403 ;
      RECT 58.51 3.025 58.575 3.401 ;
      RECT 58.495 3.025 58.51 3.393 ;
      RECT 58.48 3.025 58.495 3.38 ;
      RECT 58.475 3.025 58.48 3.37 ;
      RECT 58.46 3.025 58.475 3.348 ;
      RECT 58.445 3.025 58.46 3.315 ;
      RECT 58.44 3.025 58.445 3.293 ;
      RECT 58.43 3.025 58.44 3.275 ;
      RECT 58.415 3.025 58.43 3.253 ;
      RECT 58.395 3.025 58.415 3.215 ;
      RECT 58.745 2.31 58.78 2.749 ;
      RECT 58.745 2.31 58.785 2.748 ;
      RECT 58.69 2.37 58.785 2.747 ;
      RECT 58.555 2.542 58.785 2.746 ;
      RECT 58.665 2.42 58.785 2.746 ;
      RECT 58.555 2.542 58.81 2.736 ;
      RECT 58.61 2.487 58.89 2.653 ;
      RECT 58.785 2.281 58.79 2.744 ;
      RECT 58.64 2.457 58.93 2.53 ;
      RECT 58.655 2.44 58.785 2.746 ;
      RECT 58.79 2.28 58.96 2.468 ;
      RECT 58.78 2.283 58.96 2.468 ;
      RECT 58.285 2.16 58.455 2.47 ;
      RECT 58.285 2.16 58.46 2.443 ;
      RECT 58.285 2.16 58.465 2.42 ;
      RECT 58.285 2.16 58.475 2.37 ;
      RECT 58.28 2.265 58.475 2.34 ;
      RECT 58.315 1.835 58.485 2.313 ;
      RECT 58.315 1.835 58.5 2.234 ;
      RECT 58.305 2.045 58.5 2.234 ;
      RECT 58.315 1.845 58.51 2.149 ;
      RECT 58.245 2.587 58.25 2.79 ;
      RECT 58.235 2.575 58.245 2.9 ;
      RECT 58.21 2.575 58.235 2.94 ;
      RECT 58.13 2.575 58.21 3.025 ;
      RECT 58.12 2.575 58.13 3.095 ;
      RECT 58.095 2.575 58.12 3.118 ;
      RECT 58.075 2.575 58.095 3.153 ;
      RECT 58.03 2.585 58.075 3.196 ;
      RECT 58.02 2.597 58.03 3.233 ;
      RECT 58 2.611 58.02 3.253 ;
      RECT 57.99 2.629 58 3.269 ;
      RECT 57.975 2.655 57.99 3.279 ;
      RECT 57.96 2.696 57.975 3.293 ;
      RECT 57.95 2.731 57.96 3.303 ;
      RECT 57.945 2.747 57.95 3.308 ;
      RECT 57.935 2.762 57.945 3.313 ;
      RECT 57.915 2.805 57.935 3.323 ;
      RECT 57.895 2.842 57.915 3.336 ;
      RECT 57.86 2.865 57.895 3.354 ;
      RECT 57.85 2.879 57.86 3.37 ;
      RECT 57.83 2.889 57.85 3.38 ;
      RECT 57.825 2.898 57.83 3.388 ;
      RECT 57.815 2.905 57.825 3.395 ;
      RECT 57.805 2.912 57.815 3.403 ;
      RECT 57.79 2.922 57.805 3.411 ;
      RECT 57.78 2.936 57.79 3.421 ;
      RECT 57.77 2.948 57.78 3.433 ;
      RECT 57.755 2.97 57.77 3.446 ;
      RECT 57.745 2.992 57.755 3.457 ;
      RECT 57.735 3.012 57.745 3.466 ;
      RECT 57.73 3.027 57.735 3.473 ;
      RECT 57.7 3.06 57.73 3.487 ;
      RECT 57.69 3.095 57.7 3.502 ;
      RECT 57.685 3.102 57.69 3.508 ;
      RECT 57.665 3.117 57.685 3.515 ;
      RECT 57.66 3.132 57.665 3.523 ;
      RECT 57.655 3.141 57.66 3.528 ;
      RECT 57.64 3.147 57.655 3.535 ;
      RECT 57.635 3.153 57.64 3.543 ;
      RECT 57.63 3.157 57.635 3.55 ;
      RECT 57.625 3.161 57.63 3.56 ;
      RECT 57.615 3.166 57.625 3.57 ;
      RECT 57.595 3.177 57.615 3.598 ;
      RECT 57.58 3.189 57.595 3.625 ;
      RECT 57.56 3.202 57.58 3.65 ;
      RECT 57.54 3.217 57.56 3.674 ;
      RECT 57.525 3.232 57.54 3.689 ;
      RECT 57.52 3.243 57.525 3.698 ;
      RECT 57.455 3.288 57.52 3.708 ;
      RECT 57.42 3.347 57.455 3.721 ;
      RECT 57.415 3.37 57.42 3.727 ;
      RECT 57.41 3.377 57.415 3.729 ;
      RECT 57.395 3.387 57.41 3.732 ;
      RECT 57.365 3.412 57.395 3.736 ;
      RECT 57.36 3.43 57.365 3.74 ;
      RECT 57.355 3.437 57.36 3.741 ;
      RECT 57.335 3.445 57.355 3.745 ;
      RECT 57.325 3.452 57.335 3.749 ;
      RECT 57.281 3.463 57.325 3.756 ;
      RECT 57.195 3.491 57.281 3.772 ;
      RECT 57.135 3.515 57.195 3.79 ;
      RECT 57.09 3.525 57.135 3.804 ;
      RECT 57.031 3.533 57.09 3.818 ;
      RECT 56.945 3.54 57.031 3.837 ;
      RECT 56.92 3.545 56.945 3.852 ;
      RECT 56.84 3.548 56.92 3.855 ;
      RECT 56.76 3.552 56.84 3.842 ;
      RECT 56.751 3.555 56.76 3.827 ;
      RECT 56.665 3.555 56.751 3.812 ;
      RECT 56.605 3.557 56.665 3.789 ;
      RECT 56.601 3.56 56.605 3.779 ;
      RECT 56.515 3.56 56.601 3.764 ;
      RECT 56.44 3.56 56.515 3.74 ;
      RECT 57.755 2.569 57.765 2.745 ;
      RECT 57.71 2.536 57.755 2.745 ;
      RECT 57.665 2.487 57.71 2.745 ;
      RECT 57.635 2.457 57.665 2.746 ;
      RECT 57.63 2.44 57.635 2.747 ;
      RECT 57.605 2.42 57.63 2.748 ;
      RECT 57.59 2.395 57.605 2.749 ;
      RECT 57.585 2.382 57.59 2.75 ;
      RECT 57.58 2.376 57.585 2.748 ;
      RECT 57.575 2.368 57.58 2.742 ;
      RECT 57.55 2.36 57.575 2.722 ;
      RECT 57.53 2.349 57.55 2.693 ;
      RECT 57.5 2.334 57.53 2.664 ;
      RECT 57.48 2.32 57.5 2.636 ;
      RECT 57.47 2.314 57.48 2.615 ;
      RECT 57.465 2.311 57.47 2.598 ;
      RECT 57.46 2.308 57.465 2.583 ;
      RECT 57.445 2.303 57.46 2.548 ;
      RECT 57.44 2.299 57.445 2.515 ;
      RECT 57.42 2.294 57.44 2.491 ;
      RECT 57.39 2.286 57.42 2.456 ;
      RECT 57.375 2.28 57.39 2.433 ;
      RECT 57.335 2.273 57.375 2.418 ;
      RECT 57.31 2.265 57.335 2.398 ;
      RECT 57.29 2.26 57.31 2.388 ;
      RECT 57.255 2.254 57.29 2.383 ;
      RECT 57.21 2.245 57.255 2.382 ;
      RECT 57.18 2.241 57.21 2.384 ;
      RECT 57.095 2.249 57.18 2.388 ;
      RECT 57.025 2.26 57.095 2.41 ;
      RECT 57.012 2.266 57.025 2.433 ;
      RECT 56.926 2.273 57.012 2.455 ;
      RECT 56.84 2.285 56.926 2.492 ;
      RECT 56.84 2.662 56.85 2.9 ;
      RECT 56.835 2.291 56.84 2.515 ;
      RECT 56.83 2.547 56.84 2.9 ;
      RECT 56.83 2.292 56.835 2.52 ;
      RECT 56.825 2.293 56.83 2.9 ;
      RECT 56.801 2.295 56.825 2.901 ;
      RECT 56.715 2.303 56.801 2.903 ;
      RECT 56.695 2.317 56.715 2.906 ;
      RECT 56.69 2.345 56.695 2.907 ;
      RECT 56.685 2.357 56.69 2.908 ;
      RECT 56.68 2.372 56.685 2.909 ;
      RECT 56.67 2.402 56.68 2.91 ;
      RECT 56.665 2.44 56.67 2.908 ;
      RECT 56.66 2.46 56.665 2.903 ;
      RECT 56.645 2.495 56.66 2.888 ;
      RECT 56.635 2.547 56.645 2.868 ;
      RECT 56.63 2.577 56.635 2.856 ;
      RECT 56.615 2.59 56.63 2.839 ;
      RECT 56.59 2.594 56.615 2.806 ;
      RECT 56.575 2.592 56.59 2.783 ;
      RECT 56.56 2.591 56.575 2.78 ;
      RECT 56.5 2.589 56.56 2.778 ;
      RECT 56.49 2.587 56.5 2.773 ;
      RECT 56.45 2.586 56.49 2.77 ;
      RECT 56.38 2.583 56.45 2.768 ;
      RECT 56.325 2.581 56.38 2.763 ;
      RECT 56.255 2.575 56.325 2.758 ;
      RECT 56.246 2.575 56.255 2.755 ;
      RECT 56.16 2.575 56.246 2.75 ;
      RECT 56.155 2.575 56.16 2.745 ;
      RECT 57.46 1.81 57.635 2.16 ;
      RECT 57.46 1.825 57.645 2.158 ;
      RECT 57.435 1.775 57.58 2.155 ;
      RECT 57.415 1.776 57.58 2.148 ;
      RECT 57.405 1.777 57.59 2.143 ;
      RECT 57.375 1.778 57.59 2.13 ;
      RECT 57.325 1.779 57.59 2.106 ;
      RECT 57.32 1.781 57.59 2.091 ;
      RECT 57.32 1.847 57.65 2.085 ;
      RECT 57.3 1.788 57.605 2.065 ;
      RECT 57.29 1.797 57.615 1.92 ;
      RECT 57.3 1.792 57.615 2.065 ;
      RECT 57.32 1.782 57.605 2.091 ;
      RECT 56.905 3.107 57.075 3.395 ;
      RECT 56.9 3.125 57.085 3.39 ;
      RECT 56.865 3.133 57.15 3.31 ;
      RECT 56.865 3.133 57.236 3.3 ;
      RECT 56.865 3.133 57.29 3.246 ;
      RECT 57.15 3.03 57.32 3.214 ;
      RECT 56.865 3.185 57.325 3.202 ;
      RECT 56.85 3.155 57.32 3.198 ;
      RECT 57.11 3.037 57.15 3.349 ;
      RECT 56.99 3.074 57.32 3.214 ;
      RECT 57.085 3.049 57.11 3.375 ;
      RECT 57.075 3.056 57.32 3.214 ;
      RECT 57.206 2.52 57.275 2.779 ;
      RECT 57.206 2.575 57.28 2.778 ;
      RECT 57.12 2.575 57.28 2.777 ;
      RECT 57.115 2.575 57.285 2.77 ;
      RECT 57.105 2.52 57.275 2.765 ;
      RECT 56.485 1.819 56.66 2.12 ;
      RECT 56.47 1.807 56.485 2.105 ;
      RECT 56.44 1.806 56.47 2.058 ;
      RECT 56.44 1.824 56.665 2.053 ;
      RECT 56.425 1.808 56.485 2.018 ;
      RECT 56.42 1.83 56.675 1.918 ;
      RECT 56.42 1.813 56.571 1.918 ;
      RECT 56.42 1.815 56.575 1.918 ;
      RECT 56.425 1.811 56.571 2.018 ;
      RECT 56.53 3.047 56.535 3.395 ;
      RECT 56.52 3.037 56.53 3.401 ;
      RECT 56.485 3.027 56.52 3.403 ;
      RECT 56.447 3.022 56.485 3.407 ;
      RECT 56.361 3.015 56.447 3.414 ;
      RECT 56.275 3.005 56.361 3.424 ;
      RECT 56.23 3 56.275 3.432 ;
      RECT 56.226 3 56.23 3.436 ;
      RECT 56.14 3 56.226 3.443 ;
      RECT 56.125 3 56.14 3.443 ;
      RECT 56.115 2.998 56.125 3.415 ;
      RECT 56.105 2.994 56.115 3.358 ;
      RECT 56.085 2.988 56.105 3.29 ;
      RECT 56.08 2.984 56.085 3.238 ;
      RECT 56.07 2.983 56.08 3.205 ;
      RECT 56.02 2.981 56.07 3.19 ;
      RECT 55.995 2.979 56.02 3.185 ;
      RECT 55.952 2.977 55.995 3.181 ;
      RECT 55.866 2.973 55.952 3.169 ;
      RECT 55.78 2.968 55.866 3.153 ;
      RECT 55.75 2.965 55.78 3.14 ;
      RECT 55.725 2.964 55.75 3.128 ;
      RECT 55.72 2.964 55.725 3.118 ;
      RECT 55.68 2.963 55.72 3.11 ;
      RECT 55.665 2.962 55.68 3.103 ;
      RECT 55.615 2.961 55.665 3.095 ;
      RECT 55.613 2.96 55.615 3.09 ;
      RECT 55.527 2.958 55.613 3.09 ;
      RECT 55.441 2.953 55.527 3.09 ;
      RECT 55.355 2.949 55.441 3.09 ;
      RECT 55.306 2.945 55.355 3.088 ;
      RECT 55.22 2.942 55.306 3.083 ;
      RECT 55.197 2.939 55.22 3.079 ;
      RECT 55.111 2.936 55.197 3.074 ;
      RECT 55.025 2.932 55.111 3.065 ;
      RECT 55 2.925 55.025 3.06 ;
      RECT 54.94 2.89 55 3.057 ;
      RECT 54.92 2.815 54.94 3.054 ;
      RECT 54.915 2.757 54.92 3.053 ;
      RECT 54.89 2.697 54.915 3.052 ;
      RECT 54.815 2.575 54.89 3.048 ;
      RECT 54.805 2.575 54.815 3.04 ;
      RECT 54.79 2.575 54.805 3.03 ;
      RECT 54.775 2.575 54.79 3 ;
      RECT 54.76 2.575 54.775 2.945 ;
      RECT 54.745 2.575 54.76 2.883 ;
      RECT 54.72 2.575 54.745 2.808 ;
      RECT 54.715 2.575 54.72 2.758 ;
      RECT 56.06 2.12 56.08 2.429 ;
      RECT 56.046 2.122 56.095 2.426 ;
      RECT 56.046 2.127 56.115 2.417 ;
      RECT 55.96 2.125 56.095 2.411 ;
      RECT 55.96 2.133 56.15 2.394 ;
      RECT 55.925 2.135 56.15 2.393 ;
      RECT 55.895 2.143 56.15 2.384 ;
      RECT 55.885 2.148 56.17 2.37 ;
      RECT 55.925 2.138 56.17 2.37 ;
      RECT 55.925 2.141 56.18 2.358 ;
      RECT 55.895 2.143 56.19 2.345 ;
      RECT 55.895 2.147 56.2 2.288 ;
      RECT 55.885 2.152 56.205 2.203 ;
      RECT 56.046 2.12 56.08 2.426 ;
      RECT 55.925 7.855 56.095 8.305 ;
      RECT 55.98 6.075 56.15 8.025 ;
      RECT 55.925 5.015 56.095 6.245 ;
      RECT 55.485 2.223 55.49 2.435 ;
      RECT 55.36 2.22 55.375 2.435 ;
      RECT 54.825 2.25 54.895 2.435 ;
      RECT 54.71 2.25 54.745 2.43 ;
      RECT 55.831 2.552 55.85 2.746 ;
      RECT 55.745 2.507 55.831 2.747 ;
      RECT 55.735 2.46 55.745 2.749 ;
      RECT 55.73 2.44 55.735 2.75 ;
      RECT 55.71 2.405 55.73 2.751 ;
      RECT 55.695 2.355 55.71 2.752 ;
      RECT 55.675 2.292 55.695 2.753 ;
      RECT 55.665 2.255 55.675 2.754 ;
      RECT 55.65 2.244 55.665 2.755 ;
      RECT 55.645 2.236 55.65 2.753 ;
      RECT 55.635 2.235 55.645 2.745 ;
      RECT 55.605 2.232 55.635 2.724 ;
      RECT 55.53 2.227 55.605 2.669 ;
      RECT 55.515 2.223 55.53 2.615 ;
      RECT 55.505 2.223 55.515 2.51 ;
      RECT 55.49 2.223 55.505 2.443 ;
      RECT 55.475 2.223 55.485 2.433 ;
      RECT 55.42 2.222 55.475 2.43 ;
      RECT 55.375 2.22 55.42 2.433 ;
      RECT 55.347 2.22 55.36 2.436 ;
      RECT 55.261 2.224 55.347 2.438 ;
      RECT 55.175 2.23 55.261 2.443 ;
      RECT 55.155 2.234 55.175 2.445 ;
      RECT 55.153 2.235 55.155 2.444 ;
      RECT 55.067 2.237 55.153 2.443 ;
      RECT 54.981 2.242 55.067 2.44 ;
      RECT 54.895 2.247 54.981 2.437 ;
      RECT 54.745 2.25 54.825 2.433 ;
      RECT 55.405 5.015 55.575 8.305 ;
      RECT 55.405 7.315 55.81 7.645 ;
      RECT 55.405 6.475 55.81 6.805 ;
      RECT 55.521 3.225 55.57 3.559 ;
      RECT 55.521 3.225 55.575 3.558 ;
      RECT 55.435 3.225 55.575 3.557 ;
      RECT 55.21 3.333 55.58 3.555 ;
      RECT 55.435 3.225 55.605 3.548 ;
      RECT 55.405 3.237 55.61 3.539 ;
      RECT 55.39 3.255 55.615 3.536 ;
      RECT 55.205 3.339 55.615 3.463 ;
      RECT 55.2 3.346 55.615 3.423 ;
      RECT 55.215 3.312 55.615 3.536 ;
      RECT 55.376 3.258 55.58 3.555 ;
      RECT 55.29 3.278 55.615 3.536 ;
      RECT 55.39 3.252 55.61 3.539 ;
      RECT 55.16 2.576 55.35 2.77 ;
      RECT 55.155 2.578 55.35 2.769 ;
      RECT 55.15 2.582 55.365 2.766 ;
      RECT 55.165 2.575 55.365 2.766 ;
      RECT 55.15 2.685 55.37 2.761 ;
      RECT 54.445 3.185 54.536 3.483 ;
      RECT 54.44 3.187 54.615 3.478 ;
      RECT 54.445 3.185 54.615 3.478 ;
      RECT 54.44 3.191 54.635 3.476 ;
      RECT 54.44 3.246 54.675 3.475 ;
      RECT 54.44 3.281 54.69 3.469 ;
      RECT 54.44 3.315 54.7 3.459 ;
      RECT 54.43 3.195 54.635 3.31 ;
      RECT 54.43 3.215 54.65 3.31 ;
      RECT 54.43 3.198 54.64 3.31 ;
      RECT 54.655 1.966 54.66 2.028 ;
      RECT 54.65 1.888 54.655 2.051 ;
      RECT 54.645 1.845 54.65 2.062 ;
      RECT 54.64 1.835 54.645 2.074 ;
      RECT 54.635 1.835 54.64 2.083 ;
      RECT 54.61 1.835 54.635 2.115 ;
      RECT 54.605 1.835 54.61 2.148 ;
      RECT 54.59 1.835 54.605 2.173 ;
      RECT 54.58 1.835 54.59 2.2 ;
      RECT 54.575 1.835 54.58 2.213 ;
      RECT 54.57 1.835 54.575 2.228 ;
      RECT 54.56 1.835 54.57 2.243 ;
      RECT 54.555 1.835 54.56 2.263 ;
      RECT 54.53 1.835 54.555 2.298 ;
      RECT 54.485 1.835 54.53 2.343 ;
      RECT 54.475 1.835 54.485 2.356 ;
      RECT 54.39 1.92 54.475 2.363 ;
      RECT 54.355 2.042 54.39 2.372 ;
      RECT 54.35 2.082 54.355 2.376 ;
      RECT 54.33 2.105 54.35 2.378 ;
      RECT 54.325 2.135 54.33 2.381 ;
      RECT 54.315 2.147 54.325 2.382 ;
      RECT 54.27 2.17 54.315 2.387 ;
      RECT 54.23 2.2 54.27 2.395 ;
      RECT 54.195 2.212 54.23 2.401 ;
      RECT 54.19 2.217 54.195 2.405 ;
      RECT 54.12 2.227 54.19 2.412 ;
      RECT 54.08 2.237 54.12 2.422 ;
      RECT 54.06 2.242 54.08 2.428 ;
      RECT 54.05 2.246 54.06 2.433 ;
      RECT 54.045 2.249 54.05 2.436 ;
      RECT 54.035 2.25 54.045 2.437 ;
      RECT 54.01 2.252 54.035 2.441 ;
      RECT 54 2.257 54.01 2.444 ;
      RECT 53.955 2.265 54 2.445 ;
      RECT 53.83 2.27 53.955 2.445 ;
      RECT 54.385 2.567 54.405 2.749 ;
      RECT 54.336 2.552 54.385 2.748 ;
      RECT 54.25 2.567 54.405 2.746 ;
      RECT 54.235 2.567 54.405 2.745 ;
      RECT 54.2 2.545 54.37 2.73 ;
      RECT 54.27 3.565 54.285 3.774 ;
      RECT 54.27 3.573 54.29 3.773 ;
      RECT 54.215 3.573 54.29 3.772 ;
      RECT 54.195 3.577 54.295 3.77 ;
      RECT 54.175 3.527 54.215 3.769 ;
      RECT 54.12 3.585 54.3 3.767 ;
      RECT 54.085 3.542 54.215 3.765 ;
      RECT 54.081 3.545 54.27 3.764 ;
      RECT 53.995 3.553 54.27 3.762 ;
      RECT 53.995 3.597 54.305 3.755 ;
      RECT 53.985 3.69 54.305 3.753 ;
      RECT 53.995 3.609 54.31 3.738 ;
      RECT 53.995 3.63 54.325 3.708 ;
      RECT 53.995 3.657 54.33 3.678 ;
      RECT 54.12 3.535 54.215 3.767 ;
      RECT 53.75 2.58 53.755 3.118 ;
      RECT 53.555 2.91 53.56 3.105 ;
      RECT 51.855 2.575 51.87 2.955 ;
      RECT 53.92 2.575 53.925 2.745 ;
      RECT 53.915 2.575 53.92 2.755 ;
      RECT 53.91 2.575 53.915 2.768 ;
      RECT 53.885 2.575 53.91 2.81 ;
      RECT 53.86 2.575 53.885 2.883 ;
      RECT 53.845 2.575 53.86 2.935 ;
      RECT 53.84 2.575 53.845 2.965 ;
      RECT 53.815 2.575 53.84 3.005 ;
      RECT 53.8 2.575 53.815 3.06 ;
      RECT 53.795 2.575 53.8 3.093 ;
      RECT 53.77 2.575 53.795 3.113 ;
      RECT 53.755 2.575 53.77 3.119 ;
      RECT 53.685 2.61 53.75 3.115 ;
      RECT 53.635 2.665 53.685 3.11 ;
      RECT 53.625 2.697 53.635 3.108 ;
      RECT 53.62 2.722 53.625 3.108 ;
      RECT 53.6 2.795 53.62 3.108 ;
      RECT 53.59 2.875 53.6 3.107 ;
      RECT 53.575 2.905 53.59 3.107 ;
      RECT 53.56 2.91 53.575 3.106 ;
      RECT 53.5 2.912 53.555 3.103 ;
      RECT 53.47 2.917 53.5 3.099 ;
      RECT 53.468 2.92 53.47 3.098 ;
      RECT 53.382 2.922 53.468 3.095 ;
      RECT 53.296 2.928 53.382 3.089 ;
      RECT 53.21 2.933 53.296 3.083 ;
      RECT 53.137 2.938 53.21 3.084 ;
      RECT 53.051 2.944 53.137 3.092 ;
      RECT 52.965 2.95 53.051 3.101 ;
      RECT 52.945 2.954 52.965 3.106 ;
      RECT 52.898 2.956 52.945 3.109 ;
      RECT 52.812 2.961 52.898 3.115 ;
      RECT 52.726 2.966 52.812 3.124 ;
      RECT 52.64 2.972 52.726 3.132 ;
      RECT 52.555 2.97 52.64 3.141 ;
      RECT 52.551 2.965 52.555 3.145 ;
      RECT 52.465 2.96 52.551 3.137 ;
      RECT 52.401 2.951 52.465 3.125 ;
      RECT 52.315 2.942 52.401 3.112 ;
      RECT 52.291 2.935 52.315 3.103 ;
      RECT 52.205 2.929 52.291 3.09 ;
      RECT 52.165 2.922 52.205 3.076 ;
      RECT 52.16 2.912 52.165 3.072 ;
      RECT 52.15 2.9 52.16 3.071 ;
      RECT 52.13 2.87 52.15 3.068 ;
      RECT 52.075 2.79 52.13 3.062 ;
      RECT 52.055 2.709 52.075 3.057 ;
      RECT 52.035 2.667 52.055 3.053 ;
      RECT 52.01 2.62 52.035 3.047 ;
      RECT 52.005 2.595 52.01 3.044 ;
      RECT 51.97 2.575 52.005 3.039 ;
      RECT 51.961 2.575 51.97 3.032 ;
      RECT 51.875 2.575 51.961 3.002 ;
      RECT 51.87 2.575 51.875 2.965 ;
      RECT 51.835 2.575 51.855 2.887 ;
      RECT 51.83 2.617 51.835 2.852 ;
      RECT 51.825 2.692 51.83 2.808 ;
      RECT 53.275 2.497 53.45 2.745 ;
      RECT 53.275 2.497 53.455 2.743 ;
      RECT 53.27 2.529 53.455 2.703 ;
      RECT 53.3 2.47 53.47 2.69 ;
      RECT 53.265 2.547 53.47 2.623 ;
      RECT 52.575 2.01 52.745 2.185 ;
      RECT 52.575 2.01 52.917 2.177 ;
      RECT 52.575 2.01 53 2.171 ;
      RECT 52.575 2.01 53.035 2.167 ;
      RECT 52.575 2.01 53.055 2.166 ;
      RECT 52.575 2.01 53.141 2.162 ;
      RECT 53.035 1.835 53.205 2.157 ;
      RECT 52.61 1.942 53.235 2.155 ;
      RECT 52.6 1.997 53.24 2.153 ;
      RECT 52.575 2.033 53.25 2.148 ;
      RECT 52.575 2.06 53.255 2.078 ;
      RECT 52.64 1.885 53.215 2.155 ;
      RECT 52.831 1.87 53.215 2.155 ;
      RECT 52.665 1.873 53.215 2.155 ;
      RECT 52.745 1.871 52.831 2.182 ;
      RECT 52.831 1.868 53.21 2.155 ;
      RECT 53.015 1.845 53.21 2.155 ;
      RECT 52.917 1.866 53.21 2.155 ;
      RECT 53 1.86 53.015 2.168 ;
      RECT 53.15 3.225 53.155 3.425 ;
      RECT 52.615 3.29 52.66 3.425 ;
      RECT 53.185 3.225 53.205 3.398 ;
      RECT 53.155 3.225 53.185 3.413 ;
      RECT 53.09 3.225 53.15 3.45 ;
      RECT 53.075 3.225 53.09 3.48 ;
      RECT 53.06 3.225 53.075 3.493 ;
      RECT 53.04 3.225 53.06 3.508 ;
      RECT 53.035 3.225 53.04 3.517 ;
      RECT 53.025 3.229 53.035 3.522 ;
      RECT 53.01 3.239 53.025 3.533 ;
      RECT 52.985 3.255 53.01 3.543 ;
      RECT 52.975 3.269 52.985 3.545 ;
      RECT 52.955 3.281 52.975 3.542 ;
      RECT 52.925 3.302 52.955 3.536 ;
      RECT 52.915 3.314 52.925 3.531 ;
      RECT 52.905 3.312 52.915 3.528 ;
      RECT 52.89 3.311 52.905 3.523 ;
      RECT 52.885 3.31 52.89 3.518 ;
      RECT 52.85 3.308 52.885 3.508 ;
      RECT 52.83 3.305 52.85 3.49 ;
      RECT 52.82 3.303 52.83 3.485 ;
      RECT 52.81 3.302 52.82 3.48 ;
      RECT 52.775 3.3 52.81 3.468 ;
      RECT 52.72 3.296 52.775 3.448 ;
      RECT 52.71 3.294 52.72 3.433 ;
      RECT 52.705 3.294 52.71 3.428 ;
      RECT 52.66 3.292 52.705 3.425 ;
      RECT 52.565 3.29 52.615 3.429 ;
      RECT 52.555 3.291 52.565 3.434 ;
      RECT 52.495 3.298 52.555 3.448 ;
      RECT 52.47 3.306 52.495 3.468 ;
      RECT 52.46 3.31 52.47 3.48 ;
      RECT 52.455 3.311 52.46 3.485 ;
      RECT 52.44 3.313 52.455 3.488 ;
      RECT 52.425 3.315 52.44 3.493 ;
      RECT 52.42 3.315 52.425 3.496 ;
      RECT 52.375 3.32 52.42 3.507 ;
      RECT 52.37 3.324 52.375 3.519 ;
      RECT 52.345 3.32 52.37 3.523 ;
      RECT 52.335 3.316 52.345 3.527 ;
      RECT 52.325 3.315 52.335 3.531 ;
      RECT 52.31 3.305 52.325 3.537 ;
      RECT 52.305 3.293 52.31 3.541 ;
      RECT 52.3 3.29 52.305 3.542 ;
      RECT 52.295 3.287 52.3 3.544 ;
      RECT 52.28 3.275 52.295 3.543 ;
      RECT 52.265 3.257 52.28 3.54 ;
      RECT 52.245 3.236 52.265 3.533 ;
      RECT 52.18 3.225 52.245 3.505 ;
      RECT 52.176 3.225 52.18 3.484 ;
      RECT 52.09 3.225 52.176 3.454 ;
      RECT 52.075 3.225 52.09 3.41 ;
      RECT 52.65 2.325 52.655 2.56 ;
      RECT 51.78 2.241 51.785 2.445 ;
      RECT 52.36 2.27 52.365 2.425 ;
      RECT 52.28 2.25 52.285 2.425 ;
      RECT 52.95 2.392 52.965 2.745 ;
      RECT 52.876 2.377 52.95 2.745 ;
      RECT 52.79 2.36 52.876 2.745 ;
      RECT 52.78 2.35 52.79 2.743 ;
      RECT 52.775 2.348 52.78 2.738 ;
      RECT 52.76 2.346 52.775 2.724 ;
      RECT 52.69 2.338 52.76 2.664 ;
      RECT 52.67 2.329 52.69 2.598 ;
      RECT 52.665 2.326 52.67 2.578 ;
      RECT 52.655 2.325 52.665 2.568 ;
      RECT 52.645 2.325 52.65 2.552 ;
      RECT 52.635 2.324 52.645 2.542 ;
      RECT 52.625 2.322 52.635 2.53 ;
      RECT 52.61 2.319 52.625 2.51 ;
      RECT 52.6 2.317 52.61 2.495 ;
      RECT 52.58 2.314 52.6 2.483 ;
      RECT 52.575 2.312 52.58 2.473 ;
      RECT 52.55 2.31 52.575 2.46 ;
      RECT 52.52 2.305 52.55 2.445 ;
      RECT 52.44 2.296 52.52 2.436 ;
      RECT 52.395 2.285 52.44 2.429 ;
      RECT 52.375 2.276 52.395 2.426 ;
      RECT 52.365 2.271 52.375 2.425 ;
      RECT 52.32 2.265 52.36 2.425 ;
      RECT 52.305 2.257 52.32 2.425 ;
      RECT 52.285 2.252 52.305 2.425 ;
      RECT 52.265 2.249 52.28 2.425 ;
      RECT 52.182 2.248 52.265 2.424 ;
      RECT 52.096 2.247 52.182 2.42 ;
      RECT 52.01 2.245 52.096 2.417 ;
      RECT 51.957 2.244 52.01 2.419 ;
      RECT 51.871 2.243 51.957 2.428 ;
      RECT 51.785 2.242 51.871 2.44 ;
      RECT 51.765 2.241 51.78 2.448 ;
      RECT 51.685 2.24 51.765 2.46 ;
      RECT 51.66 2.24 51.685 2.473 ;
      RECT 51.635 2.24 51.66 2.488 ;
      RECT 51.63 2.24 51.635 2.51 ;
      RECT 51.625 2.24 51.63 2.528 ;
      RECT 51.62 2.24 51.625 2.545 ;
      RECT 51.615 2.24 51.62 2.558 ;
      RECT 51.61 2.24 51.615 2.568 ;
      RECT 51.57 2.24 51.61 2.653 ;
      RECT 51.555 2.24 51.57 2.738 ;
      RECT 51.545 2.241 51.555 2.75 ;
      RECT 51.51 2.246 51.545 2.755 ;
      RECT 51.47 2.255 51.51 2.755 ;
      RECT 51.455 2.265 51.47 2.755 ;
      RECT 51.45 2.275 51.455 2.755 ;
      RECT 51.43 2.302 51.45 2.755 ;
      RECT 51.38 2.385 51.43 2.755 ;
      RECT 51.375 2.447 51.38 2.755 ;
      RECT 51.365 2.46 51.375 2.755 ;
      RECT 51.355 2.482 51.365 2.755 ;
      RECT 51.345 2.507 51.355 2.75 ;
      RECT 51.34 2.545 51.345 2.743 ;
      RECT 51.33 2.655 51.34 2.738 ;
      RECT 52.725 3.576 52.74 3.835 ;
      RECT 52.725 3.591 52.745 3.834 ;
      RECT 52.641 3.591 52.745 3.832 ;
      RECT 52.641 3.605 52.75 3.831 ;
      RECT 52.555 3.647 52.755 3.828 ;
      RECT 52.55 3.59 52.74 3.823 ;
      RECT 52.55 3.661 52.76 3.82 ;
      RECT 52.545 3.692 52.76 3.818 ;
      RECT 52.55 3.689 52.775 3.808 ;
      RECT 52.545 3.735 52.79 3.793 ;
      RECT 52.545 3.763 52.795 3.778 ;
      RECT 52.555 3.565 52.725 3.828 ;
      RECT 52.315 2.575 52.485 2.745 ;
      RECT 52.28 2.575 52.485 2.74 ;
      RECT 52.27 2.575 52.485 2.733 ;
      RECT 52.265 2.56 52.435 2.73 ;
      RECT 51.095 3.097 51.36 3.54 ;
      RECT 51.09 3.068 51.305 3.538 ;
      RECT 51.085 3.222 51.365 3.533 ;
      RECT 51.09 3.117 51.365 3.533 ;
      RECT 51.09 3.128 51.375 3.52 ;
      RECT 51.09 3.075 51.335 3.538 ;
      RECT 51.095 3.062 51.305 3.54 ;
      RECT 51.095 3.06 51.255 3.54 ;
      RECT 51.196 3.052 51.255 3.54 ;
      RECT 51.11 3.053 51.255 3.54 ;
      RECT 51.196 3.051 51.245 3.54 ;
      RECT 51 1.866 51.175 2.165 ;
      RECT 51.05 1.828 51.175 2.165 ;
      RECT 51.035 1.83 51.261 2.157 ;
      RECT 51.035 1.833 51.3 2.144 ;
      RECT 51.035 1.834 51.31 2.13 ;
      RECT 50.99 1.885 51.31 2.12 ;
      RECT 51.035 1.835 51.315 2.115 ;
      RECT 50.99 2.045 51.32 2.105 ;
      RECT 50.975 1.905 51.315 2.045 ;
      RECT 50.97 1.921 51.315 1.985 ;
      RECT 51.015 1.845 51.315 2.115 ;
      RECT 51.05 1.826 51.136 2.165 ;
      RECT 49.51 5.02 49.68 6.49 ;
      RECT 49.51 6.315 49.685 6.485 ;
      RECT 49.14 1.74 49.31 2.93 ;
      RECT 49.14 1.74 49.61 1.91 ;
      RECT 49.14 6.97 49.61 7.14 ;
      RECT 49.14 5.95 49.31 7.14 ;
      RECT 48.15 1.74 48.32 2.93 ;
      RECT 48.15 1.74 48.62 1.91 ;
      RECT 48.15 6.97 48.62 7.14 ;
      RECT 48.15 5.95 48.32 7.14 ;
      RECT 46.3 2.635 46.47 3.865 ;
      RECT 46.355 0.855 46.525 2.805 ;
      RECT 46.3 0.575 46.47 1.025 ;
      RECT 46.3 7.855 46.47 8.305 ;
      RECT 46.355 6.075 46.525 8.025 ;
      RECT 46.3 5.015 46.47 6.245 ;
      RECT 45.78 0.575 45.95 3.865 ;
      RECT 45.78 2.075 46.185 2.405 ;
      RECT 45.78 1.235 46.185 1.565 ;
      RECT 45.78 5.015 45.95 8.305 ;
      RECT 45.78 7.315 46.185 7.645 ;
      RECT 45.78 6.475 46.185 6.805 ;
      RECT 43.705 3.126 43.71 3.298 ;
      RECT 43.7 3.119 43.705 3.388 ;
      RECT 43.695 3.113 43.7 3.407 ;
      RECT 43.675 3.107 43.695 3.417 ;
      RECT 43.66 3.102 43.675 3.425 ;
      RECT 43.623 3.096 43.66 3.423 ;
      RECT 43.537 3.082 43.623 3.419 ;
      RECT 43.451 3.064 43.537 3.414 ;
      RECT 43.365 3.045 43.451 3.408 ;
      RECT 43.335 3.033 43.365 3.404 ;
      RECT 43.315 3.027 43.335 3.403 ;
      RECT 43.25 3.025 43.315 3.401 ;
      RECT 43.235 3.025 43.25 3.393 ;
      RECT 43.22 3.025 43.235 3.38 ;
      RECT 43.215 3.025 43.22 3.37 ;
      RECT 43.2 3.025 43.215 3.348 ;
      RECT 43.185 3.025 43.2 3.315 ;
      RECT 43.18 3.025 43.185 3.293 ;
      RECT 43.17 3.025 43.18 3.275 ;
      RECT 43.155 3.025 43.17 3.253 ;
      RECT 43.135 3.025 43.155 3.215 ;
      RECT 43.485 2.31 43.52 2.749 ;
      RECT 43.485 2.31 43.525 2.748 ;
      RECT 43.43 2.37 43.525 2.747 ;
      RECT 43.295 2.542 43.525 2.746 ;
      RECT 43.405 2.42 43.525 2.746 ;
      RECT 43.295 2.542 43.55 2.736 ;
      RECT 43.35 2.487 43.63 2.653 ;
      RECT 43.525 2.281 43.53 2.744 ;
      RECT 43.38 2.457 43.67 2.53 ;
      RECT 43.395 2.44 43.525 2.746 ;
      RECT 43.53 2.28 43.7 2.468 ;
      RECT 43.52 2.283 43.7 2.468 ;
      RECT 43.025 2.16 43.195 2.47 ;
      RECT 43.025 2.16 43.2 2.443 ;
      RECT 43.025 2.16 43.205 2.42 ;
      RECT 43.025 2.16 43.215 2.37 ;
      RECT 43.02 2.265 43.215 2.34 ;
      RECT 43.055 1.835 43.225 2.313 ;
      RECT 43.055 1.835 43.24 2.234 ;
      RECT 43.045 2.045 43.24 2.234 ;
      RECT 43.055 1.845 43.25 2.149 ;
      RECT 42.985 2.587 42.99 2.79 ;
      RECT 42.975 2.575 42.985 2.9 ;
      RECT 42.95 2.575 42.975 2.94 ;
      RECT 42.87 2.575 42.95 3.025 ;
      RECT 42.86 2.575 42.87 3.095 ;
      RECT 42.835 2.575 42.86 3.118 ;
      RECT 42.815 2.575 42.835 3.153 ;
      RECT 42.77 2.585 42.815 3.196 ;
      RECT 42.76 2.597 42.77 3.233 ;
      RECT 42.74 2.611 42.76 3.253 ;
      RECT 42.73 2.629 42.74 3.269 ;
      RECT 42.715 2.655 42.73 3.279 ;
      RECT 42.7 2.696 42.715 3.293 ;
      RECT 42.69 2.731 42.7 3.303 ;
      RECT 42.685 2.747 42.69 3.308 ;
      RECT 42.675 2.762 42.685 3.313 ;
      RECT 42.655 2.805 42.675 3.323 ;
      RECT 42.635 2.842 42.655 3.336 ;
      RECT 42.6 2.865 42.635 3.354 ;
      RECT 42.59 2.879 42.6 3.37 ;
      RECT 42.57 2.889 42.59 3.38 ;
      RECT 42.565 2.898 42.57 3.388 ;
      RECT 42.555 2.905 42.565 3.395 ;
      RECT 42.545 2.912 42.555 3.403 ;
      RECT 42.53 2.922 42.545 3.411 ;
      RECT 42.52 2.936 42.53 3.421 ;
      RECT 42.51 2.948 42.52 3.433 ;
      RECT 42.495 2.97 42.51 3.446 ;
      RECT 42.485 2.992 42.495 3.457 ;
      RECT 42.475 3.012 42.485 3.466 ;
      RECT 42.47 3.027 42.475 3.473 ;
      RECT 42.44 3.06 42.47 3.487 ;
      RECT 42.43 3.095 42.44 3.502 ;
      RECT 42.425 3.102 42.43 3.508 ;
      RECT 42.405 3.117 42.425 3.515 ;
      RECT 42.4 3.132 42.405 3.523 ;
      RECT 42.395 3.141 42.4 3.528 ;
      RECT 42.38 3.147 42.395 3.535 ;
      RECT 42.375 3.153 42.38 3.543 ;
      RECT 42.37 3.157 42.375 3.55 ;
      RECT 42.365 3.161 42.37 3.56 ;
      RECT 42.355 3.166 42.365 3.57 ;
      RECT 42.335 3.177 42.355 3.598 ;
      RECT 42.32 3.189 42.335 3.625 ;
      RECT 42.3 3.202 42.32 3.65 ;
      RECT 42.28 3.217 42.3 3.674 ;
      RECT 42.265 3.232 42.28 3.689 ;
      RECT 42.26 3.243 42.265 3.698 ;
      RECT 42.195 3.288 42.26 3.708 ;
      RECT 42.16 3.347 42.195 3.721 ;
      RECT 42.155 3.37 42.16 3.727 ;
      RECT 42.15 3.377 42.155 3.729 ;
      RECT 42.135 3.387 42.15 3.732 ;
      RECT 42.105 3.412 42.135 3.736 ;
      RECT 42.1 3.43 42.105 3.74 ;
      RECT 42.095 3.437 42.1 3.741 ;
      RECT 42.075 3.445 42.095 3.745 ;
      RECT 42.065 3.452 42.075 3.749 ;
      RECT 42.021 3.463 42.065 3.756 ;
      RECT 41.935 3.491 42.021 3.772 ;
      RECT 41.875 3.515 41.935 3.79 ;
      RECT 41.83 3.525 41.875 3.804 ;
      RECT 41.771 3.533 41.83 3.818 ;
      RECT 41.685 3.54 41.771 3.837 ;
      RECT 41.66 3.545 41.685 3.852 ;
      RECT 41.58 3.548 41.66 3.855 ;
      RECT 41.5 3.552 41.58 3.842 ;
      RECT 41.491 3.555 41.5 3.827 ;
      RECT 41.405 3.555 41.491 3.812 ;
      RECT 41.345 3.557 41.405 3.789 ;
      RECT 41.341 3.56 41.345 3.779 ;
      RECT 41.255 3.56 41.341 3.764 ;
      RECT 41.18 3.56 41.255 3.74 ;
      RECT 42.495 2.569 42.505 2.745 ;
      RECT 42.45 2.536 42.495 2.745 ;
      RECT 42.405 2.487 42.45 2.745 ;
      RECT 42.375 2.457 42.405 2.746 ;
      RECT 42.37 2.44 42.375 2.747 ;
      RECT 42.345 2.42 42.37 2.748 ;
      RECT 42.33 2.395 42.345 2.749 ;
      RECT 42.325 2.382 42.33 2.75 ;
      RECT 42.32 2.376 42.325 2.748 ;
      RECT 42.315 2.368 42.32 2.742 ;
      RECT 42.29 2.36 42.315 2.722 ;
      RECT 42.27 2.349 42.29 2.693 ;
      RECT 42.24 2.334 42.27 2.664 ;
      RECT 42.22 2.32 42.24 2.636 ;
      RECT 42.21 2.314 42.22 2.615 ;
      RECT 42.205 2.311 42.21 2.598 ;
      RECT 42.2 2.308 42.205 2.583 ;
      RECT 42.185 2.303 42.2 2.548 ;
      RECT 42.18 2.299 42.185 2.515 ;
      RECT 42.16 2.294 42.18 2.491 ;
      RECT 42.13 2.286 42.16 2.456 ;
      RECT 42.115 2.28 42.13 2.433 ;
      RECT 42.075 2.273 42.115 2.418 ;
      RECT 42.05 2.265 42.075 2.398 ;
      RECT 42.03 2.26 42.05 2.388 ;
      RECT 41.995 2.254 42.03 2.383 ;
      RECT 41.95 2.245 41.995 2.382 ;
      RECT 41.92 2.241 41.95 2.384 ;
      RECT 41.835 2.249 41.92 2.388 ;
      RECT 41.765 2.26 41.835 2.41 ;
      RECT 41.752 2.266 41.765 2.433 ;
      RECT 41.666 2.273 41.752 2.455 ;
      RECT 41.58 2.285 41.666 2.492 ;
      RECT 41.58 2.662 41.59 2.9 ;
      RECT 41.575 2.291 41.58 2.515 ;
      RECT 41.57 2.547 41.58 2.9 ;
      RECT 41.57 2.292 41.575 2.52 ;
      RECT 41.565 2.293 41.57 2.9 ;
      RECT 41.541 2.295 41.565 2.901 ;
      RECT 41.455 2.303 41.541 2.903 ;
      RECT 41.435 2.317 41.455 2.906 ;
      RECT 41.43 2.345 41.435 2.907 ;
      RECT 41.425 2.357 41.43 2.908 ;
      RECT 41.42 2.372 41.425 2.909 ;
      RECT 41.41 2.402 41.42 2.91 ;
      RECT 41.405 2.44 41.41 2.908 ;
      RECT 41.4 2.46 41.405 2.903 ;
      RECT 41.385 2.495 41.4 2.888 ;
      RECT 41.375 2.547 41.385 2.868 ;
      RECT 41.37 2.577 41.375 2.856 ;
      RECT 41.355 2.59 41.37 2.839 ;
      RECT 41.33 2.594 41.355 2.806 ;
      RECT 41.315 2.592 41.33 2.783 ;
      RECT 41.3 2.591 41.315 2.78 ;
      RECT 41.24 2.589 41.3 2.778 ;
      RECT 41.23 2.587 41.24 2.773 ;
      RECT 41.19 2.586 41.23 2.77 ;
      RECT 41.12 2.583 41.19 2.768 ;
      RECT 41.065 2.581 41.12 2.763 ;
      RECT 40.995 2.575 41.065 2.758 ;
      RECT 40.986 2.575 40.995 2.755 ;
      RECT 40.9 2.575 40.986 2.75 ;
      RECT 40.895 2.575 40.9 2.745 ;
      RECT 42.2 1.81 42.375 2.16 ;
      RECT 42.2 1.825 42.385 2.158 ;
      RECT 42.175 1.775 42.32 2.155 ;
      RECT 42.155 1.776 42.32 2.148 ;
      RECT 42.145 1.777 42.33 2.143 ;
      RECT 42.115 1.778 42.33 2.13 ;
      RECT 42.065 1.779 42.33 2.106 ;
      RECT 42.06 1.781 42.33 2.091 ;
      RECT 42.06 1.847 42.39 2.085 ;
      RECT 42.04 1.788 42.345 2.065 ;
      RECT 42.03 1.797 42.355 1.92 ;
      RECT 42.04 1.792 42.355 2.065 ;
      RECT 42.06 1.782 42.345 2.091 ;
      RECT 41.645 3.107 41.815 3.395 ;
      RECT 41.64 3.125 41.825 3.39 ;
      RECT 41.605 3.133 41.89 3.31 ;
      RECT 41.605 3.133 41.976 3.3 ;
      RECT 41.605 3.133 42.03 3.246 ;
      RECT 41.89 3.03 42.06 3.214 ;
      RECT 41.605 3.185 42.065 3.202 ;
      RECT 41.59 3.155 42.06 3.198 ;
      RECT 41.85 3.037 41.89 3.349 ;
      RECT 41.73 3.074 42.06 3.214 ;
      RECT 41.825 3.049 41.85 3.375 ;
      RECT 41.815 3.056 42.06 3.214 ;
      RECT 41.946 2.52 42.015 2.779 ;
      RECT 41.946 2.575 42.02 2.778 ;
      RECT 41.86 2.575 42.02 2.777 ;
      RECT 41.855 2.575 42.025 2.77 ;
      RECT 41.845 2.52 42.015 2.765 ;
      RECT 41.225 1.819 41.4 2.12 ;
      RECT 41.21 1.807 41.225 2.105 ;
      RECT 41.18 1.806 41.21 2.058 ;
      RECT 41.18 1.824 41.405 2.053 ;
      RECT 41.165 1.808 41.225 2.018 ;
      RECT 41.16 1.83 41.415 1.918 ;
      RECT 41.16 1.813 41.311 1.918 ;
      RECT 41.16 1.815 41.315 1.918 ;
      RECT 41.165 1.811 41.311 2.018 ;
      RECT 41.27 3.047 41.275 3.395 ;
      RECT 41.26 3.037 41.27 3.401 ;
      RECT 41.225 3.027 41.26 3.403 ;
      RECT 41.187 3.022 41.225 3.407 ;
      RECT 41.101 3.015 41.187 3.414 ;
      RECT 41.015 3.005 41.101 3.424 ;
      RECT 40.97 3 41.015 3.432 ;
      RECT 40.966 3 40.97 3.436 ;
      RECT 40.88 3 40.966 3.443 ;
      RECT 40.865 3 40.88 3.443 ;
      RECT 40.855 2.998 40.865 3.415 ;
      RECT 40.845 2.994 40.855 3.358 ;
      RECT 40.825 2.988 40.845 3.29 ;
      RECT 40.82 2.984 40.825 3.238 ;
      RECT 40.81 2.983 40.82 3.205 ;
      RECT 40.76 2.981 40.81 3.19 ;
      RECT 40.735 2.979 40.76 3.185 ;
      RECT 40.692 2.977 40.735 3.181 ;
      RECT 40.606 2.973 40.692 3.169 ;
      RECT 40.52 2.968 40.606 3.153 ;
      RECT 40.49 2.965 40.52 3.14 ;
      RECT 40.465 2.964 40.49 3.128 ;
      RECT 40.46 2.964 40.465 3.118 ;
      RECT 40.42 2.963 40.46 3.11 ;
      RECT 40.405 2.962 40.42 3.103 ;
      RECT 40.355 2.961 40.405 3.095 ;
      RECT 40.353 2.96 40.355 3.09 ;
      RECT 40.267 2.958 40.353 3.09 ;
      RECT 40.181 2.953 40.267 3.09 ;
      RECT 40.095 2.949 40.181 3.09 ;
      RECT 40.046 2.945 40.095 3.088 ;
      RECT 39.96 2.942 40.046 3.083 ;
      RECT 39.937 2.939 39.96 3.079 ;
      RECT 39.851 2.936 39.937 3.074 ;
      RECT 39.765 2.932 39.851 3.065 ;
      RECT 39.74 2.925 39.765 3.06 ;
      RECT 39.68 2.89 39.74 3.057 ;
      RECT 39.66 2.815 39.68 3.054 ;
      RECT 39.655 2.757 39.66 3.053 ;
      RECT 39.63 2.697 39.655 3.052 ;
      RECT 39.555 2.575 39.63 3.048 ;
      RECT 39.545 2.575 39.555 3.04 ;
      RECT 39.53 2.575 39.545 3.03 ;
      RECT 39.515 2.575 39.53 3 ;
      RECT 39.5 2.575 39.515 2.945 ;
      RECT 39.485 2.575 39.5 2.883 ;
      RECT 39.46 2.575 39.485 2.808 ;
      RECT 39.455 2.575 39.46 2.758 ;
      RECT 40.8 2.12 40.82 2.429 ;
      RECT 40.786 2.122 40.835 2.426 ;
      RECT 40.786 2.127 40.855 2.417 ;
      RECT 40.7 2.125 40.835 2.411 ;
      RECT 40.7 2.133 40.89 2.394 ;
      RECT 40.665 2.135 40.89 2.393 ;
      RECT 40.635 2.143 40.89 2.384 ;
      RECT 40.625 2.148 40.91 2.37 ;
      RECT 40.665 2.138 40.91 2.37 ;
      RECT 40.665 2.141 40.92 2.358 ;
      RECT 40.635 2.143 40.93 2.345 ;
      RECT 40.635 2.147 40.94 2.288 ;
      RECT 40.625 2.152 40.945 2.203 ;
      RECT 40.786 2.12 40.82 2.426 ;
      RECT 40.665 7.855 40.835 8.305 ;
      RECT 40.72 6.075 40.89 8.025 ;
      RECT 40.665 5.015 40.835 6.245 ;
      RECT 40.225 2.223 40.23 2.435 ;
      RECT 40.1 2.22 40.115 2.435 ;
      RECT 39.565 2.25 39.635 2.435 ;
      RECT 39.45 2.25 39.485 2.43 ;
      RECT 40.571 2.552 40.59 2.746 ;
      RECT 40.485 2.507 40.571 2.747 ;
      RECT 40.475 2.46 40.485 2.749 ;
      RECT 40.47 2.44 40.475 2.75 ;
      RECT 40.45 2.405 40.47 2.751 ;
      RECT 40.435 2.355 40.45 2.752 ;
      RECT 40.415 2.292 40.435 2.753 ;
      RECT 40.405 2.255 40.415 2.754 ;
      RECT 40.39 2.244 40.405 2.755 ;
      RECT 40.385 2.236 40.39 2.753 ;
      RECT 40.375 2.235 40.385 2.745 ;
      RECT 40.345 2.232 40.375 2.724 ;
      RECT 40.27 2.227 40.345 2.669 ;
      RECT 40.255 2.223 40.27 2.615 ;
      RECT 40.245 2.223 40.255 2.51 ;
      RECT 40.23 2.223 40.245 2.443 ;
      RECT 40.215 2.223 40.225 2.433 ;
      RECT 40.16 2.222 40.215 2.43 ;
      RECT 40.115 2.22 40.16 2.433 ;
      RECT 40.087 2.22 40.1 2.436 ;
      RECT 40.001 2.224 40.087 2.438 ;
      RECT 39.915 2.23 40.001 2.443 ;
      RECT 39.895 2.234 39.915 2.445 ;
      RECT 39.893 2.235 39.895 2.444 ;
      RECT 39.807 2.237 39.893 2.443 ;
      RECT 39.721 2.242 39.807 2.44 ;
      RECT 39.635 2.247 39.721 2.437 ;
      RECT 39.485 2.25 39.565 2.433 ;
      RECT 40.145 5.015 40.315 8.305 ;
      RECT 40.145 7.315 40.55 7.645 ;
      RECT 40.145 6.475 40.55 6.805 ;
      RECT 40.261 3.225 40.31 3.559 ;
      RECT 40.261 3.225 40.315 3.558 ;
      RECT 40.175 3.225 40.315 3.557 ;
      RECT 39.95 3.333 40.32 3.555 ;
      RECT 40.175 3.225 40.345 3.548 ;
      RECT 40.145 3.237 40.35 3.539 ;
      RECT 40.13 3.255 40.355 3.536 ;
      RECT 39.945 3.339 40.355 3.463 ;
      RECT 39.94 3.346 40.355 3.423 ;
      RECT 39.955 3.312 40.355 3.536 ;
      RECT 40.116 3.258 40.32 3.555 ;
      RECT 40.03 3.278 40.355 3.536 ;
      RECT 40.13 3.252 40.35 3.539 ;
      RECT 39.9 2.576 40.09 2.77 ;
      RECT 39.895 2.578 40.09 2.769 ;
      RECT 39.89 2.582 40.105 2.766 ;
      RECT 39.905 2.575 40.105 2.766 ;
      RECT 39.89 2.685 40.11 2.761 ;
      RECT 39.185 3.185 39.276 3.483 ;
      RECT 39.18 3.187 39.355 3.478 ;
      RECT 39.185 3.185 39.355 3.478 ;
      RECT 39.18 3.191 39.375 3.476 ;
      RECT 39.18 3.246 39.415 3.475 ;
      RECT 39.18 3.281 39.43 3.469 ;
      RECT 39.18 3.315 39.44 3.459 ;
      RECT 39.17 3.195 39.375 3.31 ;
      RECT 39.17 3.215 39.39 3.31 ;
      RECT 39.17 3.198 39.38 3.31 ;
      RECT 39.395 1.966 39.4 2.028 ;
      RECT 39.39 1.888 39.395 2.051 ;
      RECT 39.385 1.845 39.39 2.062 ;
      RECT 39.38 1.835 39.385 2.074 ;
      RECT 39.375 1.835 39.38 2.083 ;
      RECT 39.35 1.835 39.375 2.115 ;
      RECT 39.345 1.835 39.35 2.148 ;
      RECT 39.33 1.835 39.345 2.173 ;
      RECT 39.32 1.835 39.33 2.2 ;
      RECT 39.315 1.835 39.32 2.213 ;
      RECT 39.31 1.835 39.315 2.228 ;
      RECT 39.3 1.835 39.31 2.243 ;
      RECT 39.295 1.835 39.3 2.263 ;
      RECT 39.27 1.835 39.295 2.298 ;
      RECT 39.225 1.835 39.27 2.343 ;
      RECT 39.215 1.835 39.225 2.356 ;
      RECT 39.13 1.92 39.215 2.363 ;
      RECT 39.095 2.042 39.13 2.372 ;
      RECT 39.09 2.082 39.095 2.376 ;
      RECT 39.07 2.105 39.09 2.378 ;
      RECT 39.065 2.135 39.07 2.381 ;
      RECT 39.055 2.147 39.065 2.382 ;
      RECT 39.01 2.17 39.055 2.387 ;
      RECT 38.97 2.2 39.01 2.395 ;
      RECT 38.935 2.212 38.97 2.401 ;
      RECT 38.93 2.217 38.935 2.405 ;
      RECT 38.86 2.227 38.93 2.412 ;
      RECT 38.82 2.237 38.86 2.422 ;
      RECT 38.8 2.242 38.82 2.428 ;
      RECT 38.79 2.246 38.8 2.433 ;
      RECT 38.785 2.249 38.79 2.436 ;
      RECT 38.775 2.25 38.785 2.437 ;
      RECT 38.75 2.252 38.775 2.441 ;
      RECT 38.74 2.257 38.75 2.444 ;
      RECT 38.695 2.265 38.74 2.445 ;
      RECT 38.57 2.27 38.695 2.445 ;
      RECT 39.125 2.567 39.145 2.749 ;
      RECT 39.076 2.552 39.125 2.748 ;
      RECT 38.99 2.567 39.145 2.746 ;
      RECT 38.975 2.567 39.145 2.745 ;
      RECT 38.94 2.545 39.11 2.73 ;
      RECT 39.01 3.565 39.025 3.774 ;
      RECT 39.01 3.573 39.03 3.773 ;
      RECT 38.955 3.573 39.03 3.772 ;
      RECT 38.935 3.577 39.035 3.77 ;
      RECT 38.915 3.527 38.955 3.769 ;
      RECT 38.86 3.585 39.04 3.767 ;
      RECT 38.825 3.542 38.955 3.765 ;
      RECT 38.821 3.545 39.01 3.764 ;
      RECT 38.735 3.553 39.01 3.762 ;
      RECT 38.735 3.597 39.045 3.755 ;
      RECT 38.725 3.69 39.045 3.753 ;
      RECT 38.735 3.609 39.05 3.738 ;
      RECT 38.735 3.63 39.065 3.708 ;
      RECT 38.735 3.657 39.07 3.678 ;
      RECT 38.86 3.535 38.955 3.767 ;
      RECT 38.49 2.58 38.495 3.118 ;
      RECT 38.295 2.91 38.3 3.105 ;
      RECT 36.595 2.575 36.61 2.955 ;
      RECT 38.66 2.575 38.665 2.745 ;
      RECT 38.655 2.575 38.66 2.755 ;
      RECT 38.65 2.575 38.655 2.768 ;
      RECT 38.625 2.575 38.65 2.81 ;
      RECT 38.6 2.575 38.625 2.883 ;
      RECT 38.585 2.575 38.6 2.935 ;
      RECT 38.58 2.575 38.585 2.965 ;
      RECT 38.555 2.575 38.58 3.005 ;
      RECT 38.54 2.575 38.555 3.06 ;
      RECT 38.535 2.575 38.54 3.093 ;
      RECT 38.51 2.575 38.535 3.113 ;
      RECT 38.495 2.575 38.51 3.119 ;
      RECT 38.425 2.61 38.49 3.115 ;
      RECT 38.375 2.665 38.425 3.11 ;
      RECT 38.365 2.697 38.375 3.108 ;
      RECT 38.36 2.722 38.365 3.108 ;
      RECT 38.34 2.795 38.36 3.108 ;
      RECT 38.33 2.875 38.34 3.107 ;
      RECT 38.315 2.905 38.33 3.107 ;
      RECT 38.3 2.91 38.315 3.106 ;
      RECT 38.24 2.912 38.295 3.103 ;
      RECT 38.21 2.917 38.24 3.099 ;
      RECT 38.208 2.92 38.21 3.098 ;
      RECT 38.122 2.922 38.208 3.095 ;
      RECT 38.036 2.928 38.122 3.089 ;
      RECT 37.95 2.933 38.036 3.083 ;
      RECT 37.877 2.938 37.95 3.084 ;
      RECT 37.791 2.944 37.877 3.092 ;
      RECT 37.705 2.95 37.791 3.101 ;
      RECT 37.685 2.954 37.705 3.106 ;
      RECT 37.638 2.956 37.685 3.109 ;
      RECT 37.552 2.961 37.638 3.115 ;
      RECT 37.466 2.966 37.552 3.124 ;
      RECT 37.38 2.972 37.466 3.132 ;
      RECT 37.295 2.97 37.38 3.141 ;
      RECT 37.291 2.965 37.295 3.145 ;
      RECT 37.205 2.96 37.291 3.137 ;
      RECT 37.141 2.951 37.205 3.125 ;
      RECT 37.055 2.942 37.141 3.112 ;
      RECT 37.031 2.935 37.055 3.103 ;
      RECT 36.945 2.929 37.031 3.09 ;
      RECT 36.905 2.922 36.945 3.076 ;
      RECT 36.9 2.912 36.905 3.072 ;
      RECT 36.89 2.9 36.9 3.071 ;
      RECT 36.87 2.87 36.89 3.068 ;
      RECT 36.815 2.79 36.87 3.062 ;
      RECT 36.795 2.709 36.815 3.057 ;
      RECT 36.775 2.667 36.795 3.053 ;
      RECT 36.75 2.62 36.775 3.047 ;
      RECT 36.745 2.595 36.75 3.044 ;
      RECT 36.71 2.575 36.745 3.039 ;
      RECT 36.701 2.575 36.71 3.032 ;
      RECT 36.615 2.575 36.701 3.002 ;
      RECT 36.61 2.575 36.615 2.965 ;
      RECT 36.575 2.575 36.595 2.887 ;
      RECT 36.57 2.617 36.575 2.852 ;
      RECT 36.565 2.692 36.57 2.808 ;
      RECT 38.015 2.497 38.19 2.745 ;
      RECT 38.015 2.497 38.195 2.743 ;
      RECT 38.01 2.529 38.195 2.703 ;
      RECT 38.04 2.47 38.21 2.69 ;
      RECT 38.005 2.547 38.21 2.623 ;
      RECT 37.315 2.01 37.485 2.185 ;
      RECT 37.315 2.01 37.657 2.177 ;
      RECT 37.315 2.01 37.74 2.171 ;
      RECT 37.315 2.01 37.775 2.167 ;
      RECT 37.315 2.01 37.795 2.166 ;
      RECT 37.315 2.01 37.881 2.162 ;
      RECT 37.775 1.835 37.945 2.157 ;
      RECT 37.35 1.942 37.975 2.155 ;
      RECT 37.34 1.997 37.98 2.153 ;
      RECT 37.315 2.033 37.99 2.148 ;
      RECT 37.315 2.06 37.995 2.078 ;
      RECT 37.38 1.885 37.955 2.155 ;
      RECT 37.571 1.87 37.955 2.155 ;
      RECT 37.405 1.873 37.955 2.155 ;
      RECT 37.485 1.871 37.571 2.182 ;
      RECT 37.571 1.868 37.95 2.155 ;
      RECT 37.755 1.845 37.95 2.155 ;
      RECT 37.657 1.866 37.95 2.155 ;
      RECT 37.74 1.86 37.755 2.168 ;
      RECT 37.89 3.225 37.895 3.425 ;
      RECT 37.355 3.29 37.4 3.425 ;
      RECT 37.925 3.225 37.945 3.398 ;
      RECT 37.895 3.225 37.925 3.413 ;
      RECT 37.83 3.225 37.89 3.45 ;
      RECT 37.815 3.225 37.83 3.48 ;
      RECT 37.8 3.225 37.815 3.493 ;
      RECT 37.78 3.225 37.8 3.508 ;
      RECT 37.775 3.225 37.78 3.517 ;
      RECT 37.765 3.229 37.775 3.522 ;
      RECT 37.75 3.239 37.765 3.533 ;
      RECT 37.725 3.255 37.75 3.543 ;
      RECT 37.715 3.269 37.725 3.545 ;
      RECT 37.695 3.281 37.715 3.542 ;
      RECT 37.665 3.302 37.695 3.536 ;
      RECT 37.655 3.314 37.665 3.531 ;
      RECT 37.645 3.312 37.655 3.528 ;
      RECT 37.63 3.311 37.645 3.523 ;
      RECT 37.625 3.31 37.63 3.518 ;
      RECT 37.59 3.308 37.625 3.508 ;
      RECT 37.57 3.305 37.59 3.49 ;
      RECT 37.56 3.303 37.57 3.485 ;
      RECT 37.55 3.302 37.56 3.48 ;
      RECT 37.515 3.3 37.55 3.468 ;
      RECT 37.46 3.296 37.515 3.448 ;
      RECT 37.45 3.294 37.46 3.433 ;
      RECT 37.445 3.294 37.45 3.428 ;
      RECT 37.4 3.292 37.445 3.425 ;
      RECT 37.305 3.29 37.355 3.429 ;
      RECT 37.295 3.291 37.305 3.434 ;
      RECT 37.235 3.298 37.295 3.448 ;
      RECT 37.21 3.306 37.235 3.468 ;
      RECT 37.2 3.31 37.21 3.48 ;
      RECT 37.195 3.311 37.2 3.485 ;
      RECT 37.18 3.313 37.195 3.488 ;
      RECT 37.165 3.315 37.18 3.493 ;
      RECT 37.16 3.315 37.165 3.496 ;
      RECT 37.115 3.32 37.16 3.507 ;
      RECT 37.11 3.324 37.115 3.519 ;
      RECT 37.085 3.32 37.11 3.523 ;
      RECT 37.075 3.316 37.085 3.527 ;
      RECT 37.065 3.315 37.075 3.531 ;
      RECT 37.05 3.305 37.065 3.537 ;
      RECT 37.045 3.293 37.05 3.541 ;
      RECT 37.04 3.29 37.045 3.542 ;
      RECT 37.035 3.287 37.04 3.544 ;
      RECT 37.02 3.275 37.035 3.543 ;
      RECT 37.005 3.257 37.02 3.54 ;
      RECT 36.985 3.236 37.005 3.533 ;
      RECT 36.92 3.225 36.985 3.505 ;
      RECT 36.916 3.225 36.92 3.484 ;
      RECT 36.83 3.225 36.916 3.454 ;
      RECT 36.815 3.225 36.83 3.41 ;
      RECT 37.39 2.325 37.395 2.56 ;
      RECT 36.52 2.241 36.525 2.445 ;
      RECT 37.1 2.27 37.105 2.425 ;
      RECT 37.02 2.25 37.025 2.425 ;
      RECT 37.69 2.392 37.705 2.745 ;
      RECT 37.616 2.377 37.69 2.745 ;
      RECT 37.53 2.36 37.616 2.745 ;
      RECT 37.52 2.35 37.53 2.743 ;
      RECT 37.515 2.348 37.52 2.738 ;
      RECT 37.5 2.346 37.515 2.724 ;
      RECT 37.43 2.338 37.5 2.664 ;
      RECT 37.41 2.329 37.43 2.598 ;
      RECT 37.405 2.326 37.41 2.578 ;
      RECT 37.395 2.325 37.405 2.568 ;
      RECT 37.385 2.325 37.39 2.552 ;
      RECT 37.375 2.324 37.385 2.542 ;
      RECT 37.365 2.322 37.375 2.53 ;
      RECT 37.35 2.319 37.365 2.51 ;
      RECT 37.34 2.317 37.35 2.495 ;
      RECT 37.32 2.314 37.34 2.483 ;
      RECT 37.315 2.312 37.32 2.473 ;
      RECT 37.29 2.31 37.315 2.46 ;
      RECT 37.26 2.305 37.29 2.445 ;
      RECT 37.18 2.296 37.26 2.436 ;
      RECT 37.135 2.285 37.18 2.429 ;
      RECT 37.115 2.276 37.135 2.426 ;
      RECT 37.105 2.271 37.115 2.425 ;
      RECT 37.06 2.265 37.1 2.425 ;
      RECT 37.045 2.257 37.06 2.425 ;
      RECT 37.025 2.252 37.045 2.425 ;
      RECT 37.005 2.249 37.02 2.425 ;
      RECT 36.922 2.248 37.005 2.424 ;
      RECT 36.836 2.247 36.922 2.42 ;
      RECT 36.75 2.245 36.836 2.417 ;
      RECT 36.697 2.244 36.75 2.419 ;
      RECT 36.611 2.243 36.697 2.428 ;
      RECT 36.525 2.242 36.611 2.44 ;
      RECT 36.505 2.241 36.52 2.448 ;
      RECT 36.425 2.24 36.505 2.46 ;
      RECT 36.4 2.24 36.425 2.473 ;
      RECT 36.375 2.24 36.4 2.488 ;
      RECT 36.37 2.24 36.375 2.51 ;
      RECT 36.365 2.24 36.37 2.528 ;
      RECT 36.36 2.24 36.365 2.545 ;
      RECT 36.355 2.24 36.36 2.558 ;
      RECT 36.35 2.24 36.355 2.568 ;
      RECT 36.31 2.24 36.35 2.653 ;
      RECT 36.295 2.24 36.31 2.738 ;
      RECT 36.285 2.241 36.295 2.75 ;
      RECT 36.25 2.246 36.285 2.755 ;
      RECT 36.21 2.255 36.25 2.755 ;
      RECT 36.195 2.265 36.21 2.755 ;
      RECT 36.19 2.275 36.195 2.755 ;
      RECT 36.17 2.302 36.19 2.755 ;
      RECT 36.12 2.385 36.17 2.755 ;
      RECT 36.115 2.447 36.12 2.755 ;
      RECT 36.105 2.46 36.115 2.755 ;
      RECT 36.095 2.482 36.105 2.755 ;
      RECT 36.085 2.507 36.095 2.75 ;
      RECT 36.08 2.545 36.085 2.743 ;
      RECT 36.07 2.655 36.08 2.738 ;
      RECT 37.465 3.576 37.48 3.835 ;
      RECT 37.465 3.591 37.485 3.834 ;
      RECT 37.381 3.591 37.485 3.832 ;
      RECT 37.381 3.605 37.49 3.831 ;
      RECT 37.295 3.647 37.495 3.828 ;
      RECT 37.29 3.59 37.48 3.823 ;
      RECT 37.29 3.661 37.5 3.82 ;
      RECT 37.285 3.692 37.5 3.818 ;
      RECT 37.29 3.689 37.515 3.808 ;
      RECT 37.285 3.735 37.53 3.793 ;
      RECT 37.285 3.763 37.535 3.778 ;
      RECT 37.295 3.565 37.465 3.828 ;
      RECT 37.055 2.575 37.225 2.745 ;
      RECT 37.02 2.575 37.225 2.74 ;
      RECT 37.01 2.575 37.225 2.733 ;
      RECT 37.005 2.56 37.175 2.73 ;
      RECT 35.835 3.097 36.1 3.54 ;
      RECT 35.83 3.068 36.045 3.538 ;
      RECT 35.825 3.222 36.105 3.533 ;
      RECT 35.83 3.117 36.105 3.533 ;
      RECT 35.83 3.128 36.115 3.52 ;
      RECT 35.83 3.075 36.075 3.538 ;
      RECT 35.835 3.062 36.045 3.54 ;
      RECT 35.835 3.06 35.995 3.54 ;
      RECT 35.936 3.052 35.995 3.54 ;
      RECT 35.85 3.053 35.995 3.54 ;
      RECT 35.936 3.051 35.985 3.54 ;
      RECT 35.74 1.866 35.915 2.165 ;
      RECT 35.79 1.828 35.915 2.165 ;
      RECT 35.775 1.83 36.001 2.157 ;
      RECT 35.775 1.833 36.04 2.144 ;
      RECT 35.775 1.834 36.05 2.13 ;
      RECT 35.73 1.885 36.05 2.12 ;
      RECT 35.775 1.835 36.055 2.115 ;
      RECT 35.73 2.045 36.06 2.105 ;
      RECT 35.715 1.905 36.055 2.045 ;
      RECT 35.71 1.921 36.055 1.985 ;
      RECT 35.755 1.845 36.055 2.115 ;
      RECT 35.79 1.826 35.876 2.165 ;
      RECT 34.25 5.02 34.42 6.49 ;
      RECT 34.25 6.315 34.425 6.485 ;
      RECT 33.88 1.74 34.05 2.93 ;
      RECT 33.88 1.74 34.35 1.91 ;
      RECT 33.88 6.97 34.35 7.14 ;
      RECT 33.88 5.95 34.05 7.14 ;
      RECT 32.89 1.74 33.06 2.93 ;
      RECT 32.89 1.74 33.36 1.91 ;
      RECT 32.89 6.97 33.36 7.14 ;
      RECT 32.89 5.95 33.06 7.14 ;
      RECT 31.04 2.635 31.21 3.865 ;
      RECT 31.095 0.855 31.265 2.805 ;
      RECT 31.04 0.575 31.21 1.025 ;
      RECT 31.04 7.855 31.21 8.305 ;
      RECT 31.095 6.075 31.265 8.025 ;
      RECT 31.04 5.015 31.21 6.245 ;
      RECT 30.52 0.575 30.69 3.865 ;
      RECT 30.52 2.075 30.925 2.405 ;
      RECT 30.52 1.235 30.925 1.565 ;
      RECT 30.52 5.015 30.69 8.305 ;
      RECT 30.52 7.315 30.925 7.645 ;
      RECT 30.52 6.475 30.925 6.805 ;
      RECT 28.445 3.126 28.45 3.298 ;
      RECT 28.44 3.119 28.445 3.388 ;
      RECT 28.435 3.113 28.44 3.407 ;
      RECT 28.415 3.107 28.435 3.417 ;
      RECT 28.4 3.102 28.415 3.425 ;
      RECT 28.363 3.096 28.4 3.423 ;
      RECT 28.277 3.082 28.363 3.419 ;
      RECT 28.191 3.064 28.277 3.414 ;
      RECT 28.105 3.045 28.191 3.408 ;
      RECT 28.075 3.033 28.105 3.404 ;
      RECT 28.055 3.027 28.075 3.403 ;
      RECT 27.99 3.025 28.055 3.401 ;
      RECT 27.975 3.025 27.99 3.393 ;
      RECT 27.96 3.025 27.975 3.38 ;
      RECT 27.955 3.025 27.96 3.37 ;
      RECT 27.94 3.025 27.955 3.348 ;
      RECT 27.925 3.025 27.94 3.315 ;
      RECT 27.92 3.025 27.925 3.293 ;
      RECT 27.91 3.025 27.92 3.275 ;
      RECT 27.895 3.025 27.91 3.253 ;
      RECT 27.875 3.025 27.895 3.215 ;
      RECT 28.225 2.31 28.26 2.749 ;
      RECT 28.225 2.31 28.265 2.748 ;
      RECT 28.17 2.37 28.265 2.747 ;
      RECT 28.035 2.542 28.265 2.746 ;
      RECT 28.145 2.42 28.265 2.746 ;
      RECT 28.035 2.542 28.29 2.736 ;
      RECT 28.09 2.487 28.37 2.653 ;
      RECT 28.265 2.281 28.27 2.744 ;
      RECT 28.12 2.457 28.41 2.53 ;
      RECT 28.135 2.44 28.265 2.746 ;
      RECT 28.27 2.28 28.44 2.468 ;
      RECT 28.26 2.283 28.44 2.468 ;
      RECT 27.765 2.16 27.935 2.47 ;
      RECT 27.765 2.16 27.94 2.443 ;
      RECT 27.765 2.16 27.945 2.42 ;
      RECT 27.765 2.16 27.955 2.37 ;
      RECT 27.76 2.265 27.955 2.34 ;
      RECT 27.795 1.835 27.965 2.313 ;
      RECT 27.795 1.835 27.98 2.234 ;
      RECT 27.785 2.045 27.98 2.234 ;
      RECT 27.795 1.845 27.99 2.149 ;
      RECT 27.725 2.587 27.73 2.79 ;
      RECT 27.715 2.575 27.725 2.9 ;
      RECT 27.69 2.575 27.715 2.94 ;
      RECT 27.61 2.575 27.69 3.025 ;
      RECT 27.6 2.575 27.61 3.095 ;
      RECT 27.575 2.575 27.6 3.118 ;
      RECT 27.555 2.575 27.575 3.153 ;
      RECT 27.51 2.585 27.555 3.196 ;
      RECT 27.5 2.597 27.51 3.233 ;
      RECT 27.48 2.611 27.5 3.253 ;
      RECT 27.47 2.629 27.48 3.269 ;
      RECT 27.455 2.655 27.47 3.279 ;
      RECT 27.44 2.696 27.455 3.293 ;
      RECT 27.43 2.731 27.44 3.303 ;
      RECT 27.425 2.747 27.43 3.308 ;
      RECT 27.415 2.762 27.425 3.313 ;
      RECT 27.395 2.805 27.415 3.323 ;
      RECT 27.375 2.842 27.395 3.336 ;
      RECT 27.34 2.865 27.375 3.354 ;
      RECT 27.33 2.879 27.34 3.37 ;
      RECT 27.31 2.889 27.33 3.38 ;
      RECT 27.305 2.898 27.31 3.388 ;
      RECT 27.295 2.905 27.305 3.395 ;
      RECT 27.285 2.912 27.295 3.403 ;
      RECT 27.27 2.922 27.285 3.411 ;
      RECT 27.26 2.936 27.27 3.421 ;
      RECT 27.25 2.948 27.26 3.433 ;
      RECT 27.235 2.97 27.25 3.446 ;
      RECT 27.225 2.992 27.235 3.457 ;
      RECT 27.215 3.012 27.225 3.466 ;
      RECT 27.21 3.027 27.215 3.473 ;
      RECT 27.18 3.06 27.21 3.487 ;
      RECT 27.17 3.095 27.18 3.502 ;
      RECT 27.165 3.102 27.17 3.508 ;
      RECT 27.145 3.117 27.165 3.515 ;
      RECT 27.14 3.132 27.145 3.523 ;
      RECT 27.135 3.141 27.14 3.528 ;
      RECT 27.12 3.147 27.135 3.535 ;
      RECT 27.115 3.153 27.12 3.543 ;
      RECT 27.11 3.157 27.115 3.55 ;
      RECT 27.105 3.161 27.11 3.56 ;
      RECT 27.095 3.166 27.105 3.57 ;
      RECT 27.075 3.177 27.095 3.598 ;
      RECT 27.06 3.189 27.075 3.625 ;
      RECT 27.04 3.202 27.06 3.65 ;
      RECT 27.02 3.217 27.04 3.674 ;
      RECT 27.005 3.232 27.02 3.689 ;
      RECT 27 3.243 27.005 3.698 ;
      RECT 26.935 3.288 27 3.708 ;
      RECT 26.9 3.347 26.935 3.721 ;
      RECT 26.895 3.37 26.9 3.727 ;
      RECT 26.89 3.377 26.895 3.729 ;
      RECT 26.875 3.387 26.89 3.732 ;
      RECT 26.845 3.412 26.875 3.736 ;
      RECT 26.84 3.43 26.845 3.74 ;
      RECT 26.835 3.437 26.84 3.741 ;
      RECT 26.815 3.445 26.835 3.745 ;
      RECT 26.805 3.452 26.815 3.749 ;
      RECT 26.761 3.463 26.805 3.756 ;
      RECT 26.675 3.491 26.761 3.772 ;
      RECT 26.615 3.515 26.675 3.79 ;
      RECT 26.57 3.525 26.615 3.804 ;
      RECT 26.511 3.533 26.57 3.818 ;
      RECT 26.425 3.54 26.511 3.837 ;
      RECT 26.4 3.545 26.425 3.852 ;
      RECT 26.32 3.548 26.4 3.855 ;
      RECT 26.24 3.552 26.32 3.842 ;
      RECT 26.231 3.555 26.24 3.827 ;
      RECT 26.145 3.555 26.231 3.812 ;
      RECT 26.085 3.557 26.145 3.789 ;
      RECT 26.081 3.56 26.085 3.779 ;
      RECT 25.995 3.56 26.081 3.764 ;
      RECT 25.92 3.56 25.995 3.74 ;
      RECT 27.235 2.569 27.245 2.745 ;
      RECT 27.19 2.536 27.235 2.745 ;
      RECT 27.145 2.487 27.19 2.745 ;
      RECT 27.115 2.457 27.145 2.746 ;
      RECT 27.11 2.44 27.115 2.747 ;
      RECT 27.085 2.42 27.11 2.748 ;
      RECT 27.07 2.395 27.085 2.749 ;
      RECT 27.065 2.382 27.07 2.75 ;
      RECT 27.06 2.376 27.065 2.748 ;
      RECT 27.055 2.368 27.06 2.742 ;
      RECT 27.03 2.36 27.055 2.722 ;
      RECT 27.01 2.349 27.03 2.693 ;
      RECT 26.98 2.334 27.01 2.664 ;
      RECT 26.96 2.32 26.98 2.636 ;
      RECT 26.95 2.314 26.96 2.615 ;
      RECT 26.945 2.311 26.95 2.598 ;
      RECT 26.94 2.308 26.945 2.583 ;
      RECT 26.925 2.303 26.94 2.548 ;
      RECT 26.92 2.299 26.925 2.515 ;
      RECT 26.9 2.294 26.92 2.491 ;
      RECT 26.87 2.286 26.9 2.456 ;
      RECT 26.855 2.28 26.87 2.433 ;
      RECT 26.815 2.273 26.855 2.418 ;
      RECT 26.79 2.265 26.815 2.398 ;
      RECT 26.77 2.26 26.79 2.388 ;
      RECT 26.735 2.254 26.77 2.383 ;
      RECT 26.69 2.245 26.735 2.382 ;
      RECT 26.66 2.241 26.69 2.384 ;
      RECT 26.575 2.249 26.66 2.388 ;
      RECT 26.505 2.26 26.575 2.41 ;
      RECT 26.492 2.266 26.505 2.433 ;
      RECT 26.406 2.273 26.492 2.455 ;
      RECT 26.32 2.285 26.406 2.492 ;
      RECT 26.32 2.662 26.33 2.9 ;
      RECT 26.315 2.291 26.32 2.515 ;
      RECT 26.31 2.547 26.32 2.9 ;
      RECT 26.31 2.292 26.315 2.52 ;
      RECT 26.305 2.293 26.31 2.9 ;
      RECT 26.281 2.295 26.305 2.901 ;
      RECT 26.195 2.303 26.281 2.903 ;
      RECT 26.175 2.317 26.195 2.906 ;
      RECT 26.17 2.345 26.175 2.907 ;
      RECT 26.165 2.357 26.17 2.908 ;
      RECT 26.16 2.372 26.165 2.909 ;
      RECT 26.15 2.402 26.16 2.91 ;
      RECT 26.145 2.44 26.15 2.908 ;
      RECT 26.14 2.46 26.145 2.903 ;
      RECT 26.125 2.495 26.14 2.888 ;
      RECT 26.115 2.547 26.125 2.868 ;
      RECT 26.11 2.577 26.115 2.856 ;
      RECT 26.095 2.59 26.11 2.839 ;
      RECT 26.07 2.594 26.095 2.806 ;
      RECT 26.055 2.592 26.07 2.783 ;
      RECT 26.04 2.591 26.055 2.78 ;
      RECT 25.98 2.589 26.04 2.778 ;
      RECT 25.97 2.587 25.98 2.773 ;
      RECT 25.93 2.586 25.97 2.77 ;
      RECT 25.86 2.583 25.93 2.768 ;
      RECT 25.805 2.581 25.86 2.763 ;
      RECT 25.735 2.575 25.805 2.758 ;
      RECT 25.726 2.575 25.735 2.755 ;
      RECT 25.64 2.575 25.726 2.75 ;
      RECT 25.635 2.575 25.64 2.745 ;
      RECT 26.94 1.81 27.115 2.16 ;
      RECT 26.94 1.825 27.125 2.158 ;
      RECT 26.915 1.775 27.06 2.155 ;
      RECT 26.895 1.776 27.06 2.148 ;
      RECT 26.885 1.777 27.07 2.143 ;
      RECT 26.855 1.778 27.07 2.13 ;
      RECT 26.805 1.779 27.07 2.106 ;
      RECT 26.8 1.781 27.07 2.091 ;
      RECT 26.8 1.847 27.13 2.085 ;
      RECT 26.78 1.788 27.085 2.065 ;
      RECT 26.77 1.797 27.095 1.92 ;
      RECT 26.78 1.792 27.095 2.065 ;
      RECT 26.8 1.782 27.085 2.091 ;
      RECT 26.385 3.107 26.555 3.395 ;
      RECT 26.38 3.125 26.565 3.39 ;
      RECT 26.345 3.133 26.63 3.31 ;
      RECT 26.345 3.133 26.716 3.3 ;
      RECT 26.345 3.133 26.77 3.246 ;
      RECT 26.63 3.03 26.8 3.214 ;
      RECT 26.345 3.185 26.805 3.202 ;
      RECT 26.33 3.155 26.8 3.198 ;
      RECT 26.59 3.037 26.63 3.349 ;
      RECT 26.47 3.074 26.8 3.214 ;
      RECT 26.565 3.049 26.59 3.375 ;
      RECT 26.555 3.056 26.8 3.214 ;
      RECT 26.686 2.52 26.755 2.779 ;
      RECT 26.686 2.575 26.76 2.778 ;
      RECT 26.6 2.575 26.76 2.777 ;
      RECT 26.595 2.575 26.765 2.77 ;
      RECT 26.585 2.52 26.755 2.765 ;
      RECT 25.965 1.819 26.14 2.12 ;
      RECT 25.95 1.807 25.965 2.105 ;
      RECT 25.92 1.806 25.95 2.058 ;
      RECT 25.92 1.824 26.145 2.053 ;
      RECT 25.905 1.808 25.965 2.018 ;
      RECT 25.9 1.83 26.155 1.918 ;
      RECT 25.9 1.813 26.051 1.918 ;
      RECT 25.9 1.815 26.055 1.918 ;
      RECT 25.905 1.811 26.051 2.018 ;
      RECT 26.01 3.047 26.015 3.395 ;
      RECT 26 3.037 26.01 3.401 ;
      RECT 25.965 3.027 26 3.403 ;
      RECT 25.927 3.022 25.965 3.407 ;
      RECT 25.841 3.015 25.927 3.414 ;
      RECT 25.755 3.005 25.841 3.424 ;
      RECT 25.71 3 25.755 3.432 ;
      RECT 25.706 3 25.71 3.436 ;
      RECT 25.62 3 25.706 3.443 ;
      RECT 25.605 3 25.62 3.443 ;
      RECT 25.595 2.998 25.605 3.415 ;
      RECT 25.585 2.994 25.595 3.358 ;
      RECT 25.565 2.988 25.585 3.29 ;
      RECT 25.56 2.984 25.565 3.238 ;
      RECT 25.55 2.983 25.56 3.205 ;
      RECT 25.5 2.981 25.55 3.19 ;
      RECT 25.475 2.979 25.5 3.185 ;
      RECT 25.432 2.977 25.475 3.181 ;
      RECT 25.346 2.973 25.432 3.169 ;
      RECT 25.26 2.968 25.346 3.153 ;
      RECT 25.23 2.965 25.26 3.14 ;
      RECT 25.205 2.964 25.23 3.128 ;
      RECT 25.2 2.964 25.205 3.118 ;
      RECT 25.16 2.963 25.2 3.11 ;
      RECT 25.145 2.962 25.16 3.103 ;
      RECT 25.095 2.961 25.145 3.095 ;
      RECT 25.093 2.96 25.095 3.09 ;
      RECT 25.007 2.958 25.093 3.09 ;
      RECT 24.921 2.953 25.007 3.09 ;
      RECT 24.835 2.949 24.921 3.09 ;
      RECT 24.786 2.945 24.835 3.088 ;
      RECT 24.7 2.942 24.786 3.083 ;
      RECT 24.677 2.939 24.7 3.079 ;
      RECT 24.591 2.936 24.677 3.074 ;
      RECT 24.505 2.932 24.591 3.065 ;
      RECT 24.48 2.925 24.505 3.06 ;
      RECT 24.42 2.89 24.48 3.057 ;
      RECT 24.4 2.815 24.42 3.054 ;
      RECT 24.395 2.757 24.4 3.053 ;
      RECT 24.37 2.697 24.395 3.052 ;
      RECT 24.295 2.575 24.37 3.048 ;
      RECT 24.285 2.575 24.295 3.04 ;
      RECT 24.27 2.575 24.285 3.03 ;
      RECT 24.255 2.575 24.27 3 ;
      RECT 24.24 2.575 24.255 2.945 ;
      RECT 24.225 2.575 24.24 2.883 ;
      RECT 24.2 2.575 24.225 2.808 ;
      RECT 24.195 2.575 24.2 2.758 ;
      RECT 25.54 2.12 25.56 2.429 ;
      RECT 25.526 2.122 25.575 2.426 ;
      RECT 25.526 2.127 25.595 2.417 ;
      RECT 25.44 2.125 25.575 2.411 ;
      RECT 25.44 2.133 25.63 2.394 ;
      RECT 25.405 2.135 25.63 2.393 ;
      RECT 25.375 2.143 25.63 2.384 ;
      RECT 25.365 2.148 25.65 2.37 ;
      RECT 25.405 2.138 25.65 2.37 ;
      RECT 25.405 2.141 25.66 2.358 ;
      RECT 25.375 2.143 25.67 2.345 ;
      RECT 25.375 2.147 25.68 2.288 ;
      RECT 25.365 2.152 25.685 2.203 ;
      RECT 25.526 2.12 25.56 2.426 ;
      RECT 25.405 7.855 25.575 8.305 ;
      RECT 25.46 6.075 25.63 8.025 ;
      RECT 25.405 5.015 25.575 6.245 ;
      RECT 24.965 2.223 24.97 2.435 ;
      RECT 24.84 2.22 24.855 2.435 ;
      RECT 24.305 2.25 24.375 2.435 ;
      RECT 24.19 2.25 24.225 2.43 ;
      RECT 25.311 2.552 25.33 2.746 ;
      RECT 25.225 2.507 25.311 2.747 ;
      RECT 25.215 2.46 25.225 2.749 ;
      RECT 25.21 2.44 25.215 2.75 ;
      RECT 25.19 2.405 25.21 2.751 ;
      RECT 25.175 2.355 25.19 2.752 ;
      RECT 25.155 2.292 25.175 2.753 ;
      RECT 25.145 2.255 25.155 2.754 ;
      RECT 25.13 2.244 25.145 2.755 ;
      RECT 25.125 2.236 25.13 2.753 ;
      RECT 25.115 2.235 25.125 2.745 ;
      RECT 25.085 2.232 25.115 2.724 ;
      RECT 25.01 2.227 25.085 2.669 ;
      RECT 24.995 2.223 25.01 2.615 ;
      RECT 24.985 2.223 24.995 2.51 ;
      RECT 24.97 2.223 24.985 2.443 ;
      RECT 24.955 2.223 24.965 2.433 ;
      RECT 24.9 2.222 24.955 2.43 ;
      RECT 24.855 2.22 24.9 2.433 ;
      RECT 24.827 2.22 24.84 2.436 ;
      RECT 24.741 2.224 24.827 2.438 ;
      RECT 24.655 2.23 24.741 2.443 ;
      RECT 24.635 2.234 24.655 2.445 ;
      RECT 24.633 2.235 24.635 2.444 ;
      RECT 24.547 2.237 24.633 2.443 ;
      RECT 24.461 2.242 24.547 2.44 ;
      RECT 24.375 2.247 24.461 2.437 ;
      RECT 24.225 2.25 24.305 2.433 ;
      RECT 24.885 5.015 25.055 8.305 ;
      RECT 24.885 7.315 25.29 7.645 ;
      RECT 24.885 6.475 25.29 6.805 ;
      RECT 25.001 3.225 25.05 3.559 ;
      RECT 25.001 3.225 25.055 3.558 ;
      RECT 24.915 3.225 25.055 3.557 ;
      RECT 24.69 3.333 25.06 3.555 ;
      RECT 24.915 3.225 25.085 3.548 ;
      RECT 24.885 3.237 25.09 3.539 ;
      RECT 24.87 3.255 25.095 3.536 ;
      RECT 24.685 3.339 25.095 3.463 ;
      RECT 24.68 3.346 25.095 3.423 ;
      RECT 24.695 3.312 25.095 3.536 ;
      RECT 24.856 3.258 25.06 3.555 ;
      RECT 24.77 3.278 25.095 3.536 ;
      RECT 24.87 3.252 25.09 3.539 ;
      RECT 24.64 2.576 24.83 2.77 ;
      RECT 24.635 2.578 24.83 2.769 ;
      RECT 24.63 2.582 24.845 2.766 ;
      RECT 24.645 2.575 24.845 2.766 ;
      RECT 24.63 2.685 24.85 2.761 ;
      RECT 23.925 3.185 24.016 3.483 ;
      RECT 23.92 3.187 24.095 3.478 ;
      RECT 23.925 3.185 24.095 3.478 ;
      RECT 23.92 3.191 24.115 3.476 ;
      RECT 23.92 3.246 24.155 3.475 ;
      RECT 23.92 3.281 24.17 3.469 ;
      RECT 23.92 3.315 24.18 3.459 ;
      RECT 23.91 3.195 24.115 3.31 ;
      RECT 23.91 3.215 24.13 3.31 ;
      RECT 23.91 3.198 24.12 3.31 ;
      RECT 24.135 1.966 24.14 2.028 ;
      RECT 24.13 1.888 24.135 2.051 ;
      RECT 24.125 1.845 24.13 2.062 ;
      RECT 24.12 1.835 24.125 2.074 ;
      RECT 24.115 1.835 24.12 2.083 ;
      RECT 24.09 1.835 24.115 2.115 ;
      RECT 24.085 1.835 24.09 2.148 ;
      RECT 24.07 1.835 24.085 2.173 ;
      RECT 24.06 1.835 24.07 2.2 ;
      RECT 24.055 1.835 24.06 2.213 ;
      RECT 24.05 1.835 24.055 2.228 ;
      RECT 24.04 1.835 24.05 2.243 ;
      RECT 24.035 1.835 24.04 2.263 ;
      RECT 24.01 1.835 24.035 2.298 ;
      RECT 23.965 1.835 24.01 2.343 ;
      RECT 23.955 1.835 23.965 2.356 ;
      RECT 23.87 1.92 23.955 2.363 ;
      RECT 23.835 2.042 23.87 2.372 ;
      RECT 23.83 2.082 23.835 2.376 ;
      RECT 23.81 2.105 23.83 2.378 ;
      RECT 23.805 2.135 23.81 2.381 ;
      RECT 23.795 2.147 23.805 2.382 ;
      RECT 23.75 2.17 23.795 2.387 ;
      RECT 23.71 2.2 23.75 2.395 ;
      RECT 23.675 2.212 23.71 2.401 ;
      RECT 23.67 2.217 23.675 2.405 ;
      RECT 23.6 2.227 23.67 2.412 ;
      RECT 23.56 2.237 23.6 2.422 ;
      RECT 23.54 2.242 23.56 2.428 ;
      RECT 23.53 2.246 23.54 2.433 ;
      RECT 23.525 2.249 23.53 2.436 ;
      RECT 23.515 2.25 23.525 2.437 ;
      RECT 23.49 2.252 23.515 2.441 ;
      RECT 23.48 2.257 23.49 2.444 ;
      RECT 23.435 2.265 23.48 2.445 ;
      RECT 23.31 2.27 23.435 2.445 ;
      RECT 23.865 2.567 23.885 2.749 ;
      RECT 23.816 2.552 23.865 2.748 ;
      RECT 23.73 2.567 23.885 2.746 ;
      RECT 23.715 2.567 23.885 2.745 ;
      RECT 23.68 2.545 23.85 2.73 ;
      RECT 23.75 3.565 23.765 3.774 ;
      RECT 23.75 3.573 23.77 3.773 ;
      RECT 23.695 3.573 23.77 3.772 ;
      RECT 23.675 3.577 23.775 3.77 ;
      RECT 23.655 3.527 23.695 3.769 ;
      RECT 23.6 3.585 23.78 3.767 ;
      RECT 23.565 3.542 23.695 3.765 ;
      RECT 23.561 3.545 23.75 3.764 ;
      RECT 23.475 3.553 23.75 3.762 ;
      RECT 23.475 3.597 23.785 3.755 ;
      RECT 23.465 3.69 23.785 3.753 ;
      RECT 23.475 3.609 23.79 3.738 ;
      RECT 23.475 3.63 23.805 3.708 ;
      RECT 23.475 3.657 23.81 3.678 ;
      RECT 23.6 3.535 23.695 3.767 ;
      RECT 23.23 2.58 23.235 3.118 ;
      RECT 23.035 2.91 23.04 3.105 ;
      RECT 21.335 2.575 21.35 2.955 ;
      RECT 23.4 2.575 23.405 2.745 ;
      RECT 23.395 2.575 23.4 2.755 ;
      RECT 23.39 2.575 23.395 2.768 ;
      RECT 23.365 2.575 23.39 2.81 ;
      RECT 23.34 2.575 23.365 2.883 ;
      RECT 23.325 2.575 23.34 2.935 ;
      RECT 23.32 2.575 23.325 2.965 ;
      RECT 23.295 2.575 23.32 3.005 ;
      RECT 23.28 2.575 23.295 3.06 ;
      RECT 23.275 2.575 23.28 3.093 ;
      RECT 23.25 2.575 23.275 3.113 ;
      RECT 23.235 2.575 23.25 3.119 ;
      RECT 23.165 2.61 23.23 3.115 ;
      RECT 23.115 2.665 23.165 3.11 ;
      RECT 23.105 2.697 23.115 3.108 ;
      RECT 23.1 2.722 23.105 3.108 ;
      RECT 23.08 2.795 23.1 3.108 ;
      RECT 23.07 2.875 23.08 3.107 ;
      RECT 23.055 2.905 23.07 3.107 ;
      RECT 23.04 2.91 23.055 3.106 ;
      RECT 22.98 2.912 23.035 3.103 ;
      RECT 22.95 2.917 22.98 3.099 ;
      RECT 22.948 2.92 22.95 3.098 ;
      RECT 22.862 2.922 22.948 3.095 ;
      RECT 22.776 2.928 22.862 3.089 ;
      RECT 22.69 2.933 22.776 3.083 ;
      RECT 22.617 2.938 22.69 3.084 ;
      RECT 22.531 2.944 22.617 3.092 ;
      RECT 22.445 2.95 22.531 3.101 ;
      RECT 22.425 2.954 22.445 3.106 ;
      RECT 22.378 2.956 22.425 3.109 ;
      RECT 22.292 2.961 22.378 3.115 ;
      RECT 22.206 2.966 22.292 3.124 ;
      RECT 22.12 2.972 22.206 3.132 ;
      RECT 22.035 2.97 22.12 3.141 ;
      RECT 22.031 2.965 22.035 3.145 ;
      RECT 21.945 2.96 22.031 3.137 ;
      RECT 21.881 2.951 21.945 3.125 ;
      RECT 21.795 2.942 21.881 3.112 ;
      RECT 21.771 2.935 21.795 3.103 ;
      RECT 21.685 2.929 21.771 3.09 ;
      RECT 21.645 2.922 21.685 3.076 ;
      RECT 21.64 2.912 21.645 3.072 ;
      RECT 21.63 2.9 21.64 3.071 ;
      RECT 21.61 2.87 21.63 3.068 ;
      RECT 21.555 2.79 21.61 3.062 ;
      RECT 21.535 2.709 21.555 3.057 ;
      RECT 21.515 2.667 21.535 3.053 ;
      RECT 21.49 2.62 21.515 3.047 ;
      RECT 21.485 2.595 21.49 3.044 ;
      RECT 21.45 2.575 21.485 3.039 ;
      RECT 21.441 2.575 21.45 3.032 ;
      RECT 21.355 2.575 21.441 3.002 ;
      RECT 21.35 2.575 21.355 2.965 ;
      RECT 21.315 2.575 21.335 2.887 ;
      RECT 21.31 2.617 21.315 2.852 ;
      RECT 21.305 2.692 21.31 2.808 ;
      RECT 22.755 2.497 22.93 2.745 ;
      RECT 22.755 2.497 22.935 2.743 ;
      RECT 22.75 2.529 22.935 2.703 ;
      RECT 22.78 2.47 22.95 2.69 ;
      RECT 22.745 2.547 22.95 2.623 ;
      RECT 22.055 2.01 22.225 2.185 ;
      RECT 22.055 2.01 22.397 2.177 ;
      RECT 22.055 2.01 22.48 2.171 ;
      RECT 22.055 2.01 22.515 2.167 ;
      RECT 22.055 2.01 22.535 2.166 ;
      RECT 22.055 2.01 22.621 2.162 ;
      RECT 22.515 1.835 22.685 2.157 ;
      RECT 22.09 1.942 22.715 2.155 ;
      RECT 22.08 1.997 22.72 2.153 ;
      RECT 22.055 2.033 22.73 2.148 ;
      RECT 22.055 2.06 22.735 2.078 ;
      RECT 22.12 1.885 22.695 2.155 ;
      RECT 22.311 1.87 22.695 2.155 ;
      RECT 22.145 1.873 22.695 2.155 ;
      RECT 22.225 1.871 22.311 2.182 ;
      RECT 22.311 1.868 22.69 2.155 ;
      RECT 22.495 1.845 22.69 2.155 ;
      RECT 22.397 1.866 22.69 2.155 ;
      RECT 22.48 1.86 22.495 2.168 ;
      RECT 22.63 3.225 22.635 3.425 ;
      RECT 22.095 3.29 22.14 3.425 ;
      RECT 22.665 3.225 22.685 3.398 ;
      RECT 22.635 3.225 22.665 3.413 ;
      RECT 22.57 3.225 22.63 3.45 ;
      RECT 22.555 3.225 22.57 3.48 ;
      RECT 22.54 3.225 22.555 3.493 ;
      RECT 22.52 3.225 22.54 3.508 ;
      RECT 22.515 3.225 22.52 3.517 ;
      RECT 22.505 3.229 22.515 3.522 ;
      RECT 22.49 3.239 22.505 3.533 ;
      RECT 22.465 3.255 22.49 3.543 ;
      RECT 22.455 3.269 22.465 3.545 ;
      RECT 22.435 3.281 22.455 3.542 ;
      RECT 22.405 3.302 22.435 3.536 ;
      RECT 22.395 3.314 22.405 3.531 ;
      RECT 22.385 3.312 22.395 3.528 ;
      RECT 22.37 3.311 22.385 3.523 ;
      RECT 22.365 3.31 22.37 3.518 ;
      RECT 22.33 3.308 22.365 3.508 ;
      RECT 22.31 3.305 22.33 3.49 ;
      RECT 22.3 3.303 22.31 3.485 ;
      RECT 22.29 3.302 22.3 3.48 ;
      RECT 22.255 3.3 22.29 3.468 ;
      RECT 22.2 3.296 22.255 3.448 ;
      RECT 22.19 3.294 22.2 3.433 ;
      RECT 22.185 3.294 22.19 3.428 ;
      RECT 22.14 3.292 22.185 3.425 ;
      RECT 22.045 3.29 22.095 3.429 ;
      RECT 22.035 3.291 22.045 3.434 ;
      RECT 21.975 3.298 22.035 3.448 ;
      RECT 21.95 3.306 21.975 3.468 ;
      RECT 21.94 3.31 21.95 3.48 ;
      RECT 21.935 3.311 21.94 3.485 ;
      RECT 21.92 3.313 21.935 3.488 ;
      RECT 21.905 3.315 21.92 3.493 ;
      RECT 21.9 3.315 21.905 3.496 ;
      RECT 21.855 3.32 21.9 3.507 ;
      RECT 21.85 3.324 21.855 3.519 ;
      RECT 21.825 3.32 21.85 3.523 ;
      RECT 21.815 3.316 21.825 3.527 ;
      RECT 21.805 3.315 21.815 3.531 ;
      RECT 21.79 3.305 21.805 3.537 ;
      RECT 21.785 3.293 21.79 3.541 ;
      RECT 21.78 3.29 21.785 3.542 ;
      RECT 21.775 3.287 21.78 3.544 ;
      RECT 21.76 3.275 21.775 3.543 ;
      RECT 21.745 3.257 21.76 3.54 ;
      RECT 21.725 3.236 21.745 3.533 ;
      RECT 21.66 3.225 21.725 3.505 ;
      RECT 21.656 3.225 21.66 3.484 ;
      RECT 21.57 3.225 21.656 3.454 ;
      RECT 21.555 3.225 21.57 3.41 ;
      RECT 22.13 2.325 22.135 2.56 ;
      RECT 21.26 2.241 21.265 2.445 ;
      RECT 21.84 2.27 21.845 2.425 ;
      RECT 21.76 2.25 21.765 2.425 ;
      RECT 22.43 2.392 22.445 2.745 ;
      RECT 22.356 2.377 22.43 2.745 ;
      RECT 22.27 2.36 22.356 2.745 ;
      RECT 22.26 2.35 22.27 2.743 ;
      RECT 22.255 2.348 22.26 2.738 ;
      RECT 22.24 2.346 22.255 2.724 ;
      RECT 22.17 2.338 22.24 2.664 ;
      RECT 22.15 2.329 22.17 2.598 ;
      RECT 22.145 2.326 22.15 2.578 ;
      RECT 22.135 2.325 22.145 2.568 ;
      RECT 22.125 2.325 22.13 2.552 ;
      RECT 22.115 2.324 22.125 2.542 ;
      RECT 22.105 2.322 22.115 2.53 ;
      RECT 22.09 2.319 22.105 2.51 ;
      RECT 22.08 2.317 22.09 2.495 ;
      RECT 22.06 2.314 22.08 2.483 ;
      RECT 22.055 2.312 22.06 2.473 ;
      RECT 22.03 2.31 22.055 2.46 ;
      RECT 22 2.305 22.03 2.445 ;
      RECT 21.92 2.296 22 2.436 ;
      RECT 21.875 2.285 21.92 2.429 ;
      RECT 21.855 2.276 21.875 2.426 ;
      RECT 21.845 2.271 21.855 2.425 ;
      RECT 21.8 2.265 21.84 2.425 ;
      RECT 21.785 2.257 21.8 2.425 ;
      RECT 21.765 2.252 21.785 2.425 ;
      RECT 21.745 2.249 21.76 2.425 ;
      RECT 21.662 2.248 21.745 2.424 ;
      RECT 21.576 2.247 21.662 2.42 ;
      RECT 21.49 2.245 21.576 2.417 ;
      RECT 21.437 2.244 21.49 2.419 ;
      RECT 21.351 2.243 21.437 2.428 ;
      RECT 21.265 2.242 21.351 2.44 ;
      RECT 21.245 2.241 21.26 2.448 ;
      RECT 21.165 2.24 21.245 2.46 ;
      RECT 21.14 2.24 21.165 2.473 ;
      RECT 21.115 2.24 21.14 2.488 ;
      RECT 21.11 2.24 21.115 2.51 ;
      RECT 21.105 2.24 21.11 2.528 ;
      RECT 21.1 2.24 21.105 2.545 ;
      RECT 21.095 2.24 21.1 2.558 ;
      RECT 21.09 2.24 21.095 2.568 ;
      RECT 21.05 2.24 21.09 2.653 ;
      RECT 21.035 2.24 21.05 2.738 ;
      RECT 21.025 2.241 21.035 2.75 ;
      RECT 20.99 2.246 21.025 2.755 ;
      RECT 20.95 2.255 20.99 2.755 ;
      RECT 20.935 2.265 20.95 2.755 ;
      RECT 20.93 2.275 20.935 2.755 ;
      RECT 20.91 2.302 20.93 2.755 ;
      RECT 20.86 2.385 20.91 2.755 ;
      RECT 20.855 2.447 20.86 2.755 ;
      RECT 20.845 2.46 20.855 2.755 ;
      RECT 20.835 2.482 20.845 2.755 ;
      RECT 20.825 2.507 20.835 2.75 ;
      RECT 20.82 2.545 20.825 2.743 ;
      RECT 20.81 2.655 20.82 2.738 ;
      RECT 22.205 3.576 22.22 3.835 ;
      RECT 22.205 3.591 22.225 3.834 ;
      RECT 22.121 3.591 22.225 3.832 ;
      RECT 22.121 3.605 22.23 3.831 ;
      RECT 22.035 3.647 22.235 3.828 ;
      RECT 22.03 3.59 22.22 3.823 ;
      RECT 22.03 3.661 22.24 3.82 ;
      RECT 22.025 3.692 22.24 3.818 ;
      RECT 22.03 3.689 22.255 3.808 ;
      RECT 22.025 3.735 22.27 3.793 ;
      RECT 22.025 3.763 22.275 3.778 ;
      RECT 22.035 3.565 22.205 3.828 ;
      RECT 21.795 2.575 21.965 2.745 ;
      RECT 21.76 2.575 21.965 2.74 ;
      RECT 21.75 2.575 21.965 2.733 ;
      RECT 21.745 2.56 21.915 2.73 ;
      RECT 20.575 3.097 20.84 3.54 ;
      RECT 20.57 3.068 20.785 3.538 ;
      RECT 20.565 3.222 20.845 3.533 ;
      RECT 20.57 3.117 20.845 3.533 ;
      RECT 20.57 3.128 20.855 3.52 ;
      RECT 20.57 3.075 20.815 3.538 ;
      RECT 20.575 3.062 20.785 3.54 ;
      RECT 20.575 3.06 20.735 3.54 ;
      RECT 20.676 3.052 20.735 3.54 ;
      RECT 20.59 3.053 20.735 3.54 ;
      RECT 20.676 3.051 20.725 3.54 ;
      RECT 20.48 1.866 20.655 2.165 ;
      RECT 20.53 1.828 20.655 2.165 ;
      RECT 20.515 1.83 20.741 2.157 ;
      RECT 20.515 1.833 20.78 2.144 ;
      RECT 20.515 1.834 20.79 2.13 ;
      RECT 20.47 1.885 20.79 2.12 ;
      RECT 20.515 1.835 20.795 2.115 ;
      RECT 20.47 2.045 20.8 2.105 ;
      RECT 20.455 1.905 20.795 2.045 ;
      RECT 20.45 1.921 20.795 1.985 ;
      RECT 20.495 1.845 20.795 2.115 ;
      RECT 20.53 1.826 20.616 2.165 ;
      RECT 18.99 5.02 19.16 6.49 ;
      RECT 18.99 6.315 19.165 6.485 ;
      RECT 18.62 1.74 18.79 2.93 ;
      RECT 18.62 1.74 19.09 1.91 ;
      RECT 18.62 6.97 19.09 7.14 ;
      RECT 18.62 5.95 18.79 7.14 ;
      RECT 17.63 1.74 17.8 2.93 ;
      RECT 17.63 1.74 18.1 1.91 ;
      RECT 17.63 6.97 18.1 7.14 ;
      RECT 17.63 5.95 17.8 7.14 ;
      RECT 15.78 2.635 15.95 3.865 ;
      RECT 15.835 0.855 16.005 2.805 ;
      RECT 15.78 0.575 15.95 1.025 ;
      RECT 15.78 7.855 15.95 8.305 ;
      RECT 15.835 6.075 16.005 8.025 ;
      RECT 15.78 5.015 15.95 6.245 ;
      RECT 15.26 0.575 15.43 3.865 ;
      RECT 15.26 2.075 15.665 2.405 ;
      RECT 15.26 1.235 15.665 1.565 ;
      RECT 15.26 5.015 15.43 8.305 ;
      RECT 15.26 7.315 15.665 7.645 ;
      RECT 15.26 6.475 15.665 6.805 ;
      RECT 13.185 3.126 13.19 3.298 ;
      RECT 13.18 3.119 13.185 3.388 ;
      RECT 13.175 3.113 13.18 3.407 ;
      RECT 13.155 3.107 13.175 3.417 ;
      RECT 13.14 3.102 13.155 3.425 ;
      RECT 13.103 3.096 13.14 3.423 ;
      RECT 13.017 3.082 13.103 3.419 ;
      RECT 12.931 3.064 13.017 3.414 ;
      RECT 12.845 3.045 12.931 3.408 ;
      RECT 12.815 3.033 12.845 3.404 ;
      RECT 12.795 3.027 12.815 3.403 ;
      RECT 12.73 3.025 12.795 3.401 ;
      RECT 12.715 3.025 12.73 3.393 ;
      RECT 12.7 3.025 12.715 3.38 ;
      RECT 12.695 3.025 12.7 3.37 ;
      RECT 12.68 3.025 12.695 3.348 ;
      RECT 12.665 3.025 12.68 3.315 ;
      RECT 12.66 3.025 12.665 3.293 ;
      RECT 12.65 3.025 12.66 3.275 ;
      RECT 12.635 3.025 12.65 3.253 ;
      RECT 12.615 3.025 12.635 3.215 ;
      RECT 12.965 2.31 13 2.749 ;
      RECT 12.965 2.31 13.005 2.748 ;
      RECT 12.91 2.37 13.005 2.747 ;
      RECT 12.775 2.542 13.005 2.746 ;
      RECT 12.885 2.42 13.005 2.746 ;
      RECT 12.775 2.542 13.03 2.736 ;
      RECT 12.83 2.487 13.11 2.653 ;
      RECT 13.005 2.281 13.01 2.744 ;
      RECT 12.86 2.457 13.15 2.53 ;
      RECT 12.875 2.44 13.005 2.746 ;
      RECT 13.01 2.28 13.18 2.468 ;
      RECT 13 2.283 13.18 2.468 ;
      RECT 12.505 2.16 12.675 2.47 ;
      RECT 12.505 2.16 12.68 2.443 ;
      RECT 12.505 2.16 12.685 2.42 ;
      RECT 12.505 2.16 12.695 2.37 ;
      RECT 12.5 2.265 12.695 2.34 ;
      RECT 12.535 1.835 12.705 2.313 ;
      RECT 12.535 1.835 12.72 2.234 ;
      RECT 12.525 2.045 12.72 2.234 ;
      RECT 12.535 1.845 12.73 2.149 ;
      RECT 12.465 2.587 12.47 2.79 ;
      RECT 12.455 2.575 12.465 2.9 ;
      RECT 12.43 2.575 12.455 2.94 ;
      RECT 12.35 2.575 12.43 3.025 ;
      RECT 12.34 2.575 12.35 3.095 ;
      RECT 12.315 2.575 12.34 3.118 ;
      RECT 12.295 2.575 12.315 3.153 ;
      RECT 12.25 2.585 12.295 3.196 ;
      RECT 12.24 2.597 12.25 3.233 ;
      RECT 12.22 2.611 12.24 3.253 ;
      RECT 12.21 2.629 12.22 3.269 ;
      RECT 12.195 2.655 12.21 3.279 ;
      RECT 12.18 2.696 12.195 3.293 ;
      RECT 12.17 2.731 12.18 3.303 ;
      RECT 12.165 2.747 12.17 3.308 ;
      RECT 12.155 2.762 12.165 3.313 ;
      RECT 12.135 2.805 12.155 3.323 ;
      RECT 12.115 2.842 12.135 3.336 ;
      RECT 12.08 2.865 12.115 3.354 ;
      RECT 12.07 2.879 12.08 3.37 ;
      RECT 12.05 2.889 12.07 3.38 ;
      RECT 12.045 2.898 12.05 3.388 ;
      RECT 12.035 2.905 12.045 3.395 ;
      RECT 12.025 2.912 12.035 3.403 ;
      RECT 12.01 2.922 12.025 3.411 ;
      RECT 12 2.936 12.01 3.421 ;
      RECT 11.99 2.948 12 3.433 ;
      RECT 11.975 2.97 11.99 3.446 ;
      RECT 11.965 2.992 11.975 3.457 ;
      RECT 11.955 3.012 11.965 3.466 ;
      RECT 11.95 3.027 11.955 3.473 ;
      RECT 11.92 3.06 11.95 3.487 ;
      RECT 11.91 3.095 11.92 3.502 ;
      RECT 11.905 3.102 11.91 3.508 ;
      RECT 11.885 3.117 11.905 3.515 ;
      RECT 11.88 3.132 11.885 3.523 ;
      RECT 11.875 3.141 11.88 3.528 ;
      RECT 11.86 3.147 11.875 3.535 ;
      RECT 11.855 3.153 11.86 3.543 ;
      RECT 11.85 3.157 11.855 3.55 ;
      RECT 11.845 3.161 11.85 3.56 ;
      RECT 11.835 3.166 11.845 3.57 ;
      RECT 11.815 3.177 11.835 3.598 ;
      RECT 11.8 3.189 11.815 3.625 ;
      RECT 11.78 3.202 11.8 3.65 ;
      RECT 11.76 3.217 11.78 3.674 ;
      RECT 11.745 3.232 11.76 3.689 ;
      RECT 11.74 3.243 11.745 3.698 ;
      RECT 11.675 3.288 11.74 3.708 ;
      RECT 11.64 3.347 11.675 3.721 ;
      RECT 11.635 3.37 11.64 3.727 ;
      RECT 11.63 3.377 11.635 3.729 ;
      RECT 11.615 3.387 11.63 3.732 ;
      RECT 11.585 3.412 11.615 3.736 ;
      RECT 11.58 3.43 11.585 3.74 ;
      RECT 11.575 3.437 11.58 3.741 ;
      RECT 11.555 3.445 11.575 3.745 ;
      RECT 11.545 3.452 11.555 3.749 ;
      RECT 11.501 3.463 11.545 3.756 ;
      RECT 11.415 3.491 11.501 3.772 ;
      RECT 11.355 3.515 11.415 3.79 ;
      RECT 11.31 3.525 11.355 3.804 ;
      RECT 11.251 3.533 11.31 3.818 ;
      RECT 11.165 3.54 11.251 3.837 ;
      RECT 11.14 3.545 11.165 3.852 ;
      RECT 11.06 3.548 11.14 3.855 ;
      RECT 10.98 3.552 11.06 3.842 ;
      RECT 10.971 3.555 10.98 3.827 ;
      RECT 10.885 3.555 10.971 3.812 ;
      RECT 10.825 3.557 10.885 3.789 ;
      RECT 10.821 3.56 10.825 3.779 ;
      RECT 10.735 3.56 10.821 3.764 ;
      RECT 10.66 3.56 10.735 3.74 ;
      RECT 11.975 2.569 11.985 2.745 ;
      RECT 11.93 2.536 11.975 2.745 ;
      RECT 11.885 2.487 11.93 2.745 ;
      RECT 11.855 2.457 11.885 2.746 ;
      RECT 11.85 2.44 11.855 2.747 ;
      RECT 11.825 2.42 11.85 2.748 ;
      RECT 11.81 2.395 11.825 2.749 ;
      RECT 11.805 2.382 11.81 2.75 ;
      RECT 11.8 2.376 11.805 2.748 ;
      RECT 11.795 2.368 11.8 2.742 ;
      RECT 11.77 2.36 11.795 2.722 ;
      RECT 11.75 2.349 11.77 2.693 ;
      RECT 11.72 2.334 11.75 2.664 ;
      RECT 11.7 2.32 11.72 2.636 ;
      RECT 11.69 2.314 11.7 2.615 ;
      RECT 11.685 2.311 11.69 2.598 ;
      RECT 11.68 2.308 11.685 2.583 ;
      RECT 11.665 2.303 11.68 2.548 ;
      RECT 11.66 2.299 11.665 2.515 ;
      RECT 11.64 2.294 11.66 2.491 ;
      RECT 11.61 2.286 11.64 2.456 ;
      RECT 11.595 2.28 11.61 2.433 ;
      RECT 11.555 2.273 11.595 2.418 ;
      RECT 11.53 2.265 11.555 2.398 ;
      RECT 11.51 2.26 11.53 2.388 ;
      RECT 11.475 2.254 11.51 2.383 ;
      RECT 11.43 2.245 11.475 2.382 ;
      RECT 11.4 2.241 11.43 2.384 ;
      RECT 11.315 2.249 11.4 2.388 ;
      RECT 11.245 2.26 11.315 2.41 ;
      RECT 11.232 2.266 11.245 2.433 ;
      RECT 11.146 2.273 11.232 2.455 ;
      RECT 11.06 2.285 11.146 2.492 ;
      RECT 11.06 2.662 11.07 2.9 ;
      RECT 11.055 2.291 11.06 2.515 ;
      RECT 11.05 2.547 11.06 2.9 ;
      RECT 11.05 2.292 11.055 2.52 ;
      RECT 11.045 2.293 11.05 2.9 ;
      RECT 11.021 2.295 11.045 2.901 ;
      RECT 10.935 2.303 11.021 2.903 ;
      RECT 10.915 2.317 10.935 2.906 ;
      RECT 10.91 2.345 10.915 2.907 ;
      RECT 10.905 2.357 10.91 2.908 ;
      RECT 10.9 2.372 10.905 2.909 ;
      RECT 10.89 2.402 10.9 2.91 ;
      RECT 10.885 2.44 10.89 2.908 ;
      RECT 10.88 2.46 10.885 2.903 ;
      RECT 10.865 2.495 10.88 2.888 ;
      RECT 10.855 2.547 10.865 2.868 ;
      RECT 10.85 2.577 10.855 2.856 ;
      RECT 10.835 2.59 10.85 2.839 ;
      RECT 10.81 2.594 10.835 2.806 ;
      RECT 10.795 2.592 10.81 2.783 ;
      RECT 10.78 2.591 10.795 2.78 ;
      RECT 10.72 2.589 10.78 2.778 ;
      RECT 10.71 2.587 10.72 2.773 ;
      RECT 10.67 2.586 10.71 2.77 ;
      RECT 10.6 2.583 10.67 2.768 ;
      RECT 10.545 2.581 10.6 2.763 ;
      RECT 10.475 2.575 10.545 2.758 ;
      RECT 10.466 2.575 10.475 2.755 ;
      RECT 10.38 2.575 10.466 2.75 ;
      RECT 10.375 2.575 10.38 2.745 ;
      RECT 11.68 1.81 11.855 2.16 ;
      RECT 11.68 1.825 11.865 2.158 ;
      RECT 11.655 1.775 11.8 2.155 ;
      RECT 11.635 1.776 11.8 2.148 ;
      RECT 11.625 1.777 11.81 2.143 ;
      RECT 11.595 1.778 11.81 2.13 ;
      RECT 11.545 1.779 11.81 2.106 ;
      RECT 11.54 1.781 11.81 2.091 ;
      RECT 11.54 1.847 11.87 2.085 ;
      RECT 11.52 1.788 11.825 2.065 ;
      RECT 11.51 1.797 11.835 1.92 ;
      RECT 11.52 1.792 11.835 2.065 ;
      RECT 11.54 1.782 11.825 2.091 ;
      RECT 11.125 3.107 11.295 3.395 ;
      RECT 11.12 3.125 11.305 3.39 ;
      RECT 11.085 3.133 11.37 3.31 ;
      RECT 11.085 3.133 11.456 3.3 ;
      RECT 11.085 3.133 11.51 3.246 ;
      RECT 11.37 3.03 11.54 3.214 ;
      RECT 11.085 3.185 11.545 3.202 ;
      RECT 11.07 3.155 11.54 3.198 ;
      RECT 11.33 3.037 11.37 3.349 ;
      RECT 11.21 3.074 11.54 3.214 ;
      RECT 11.305 3.049 11.33 3.375 ;
      RECT 11.295 3.056 11.54 3.214 ;
      RECT 11.426 2.52 11.495 2.779 ;
      RECT 11.426 2.575 11.5 2.778 ;
      RECT 11.34 2.575 11.5 2.777 ;
      RECT 11.335 2.575 11.505 2.77 ;
      RECT 11.325 2.52 11.495 2.765 ;
      RECT 10.705 1.819 10.88 2.12 ;
      RECT 10.69 1.807 10.705 2.105 ;
      RECT 10.66 1.806 10.69 2.058 ;
      RECT 10.66 1.824 10.885 2.053 ;
      RECT 10.645 1.808 10.705 2.018 ;
      RECT 10.64 1.83 10.895 1.918 ;
      RECT 10.64 1.813 10.791 1.918 ;
      RECT 10.64 1.815 10.795 1.918 ;
      RECT 10.645 1.811 10.791 2.018 ;
      RECT 10.75 3.047 10.755 3.395 ;
      RECT 10.74 3.037 10.75 3.401 ;
      RECT 10.705 3.027 10.74 3.403 ;
      RECT 10.667 3.022 10.705 3.407 ;
      RECT 10.581 3.015 10.667 3.414 ;
      RECT 10.495 3.005 10.581 3.424 ;
      RECT 10.45 3 10.495 3.432 ;
      RECT 10.446 3 10.45 3.436 ;
      RECT 10.36 3 10.446 3.443 ;
      RECT 10.345 3 10.36 3.443 ;
      RECT 10.335 2.998 10.345 3.415 ;
      RECT 10.325 2.994 10.335 3.358 ;
      RECT 10.305 2.988 10.325 3.29 ;
      RECT 10.3 2.984 10.305 3.238 ;
      RECT 10.29 2.983 10.3 3.205 ;
      RECT 10.24 2.981 10.29 3.19 ;
      RECT 10.215 2.979 10.24 3.185 ;
      RECT 10.172 2.977 10.215 3.181 ;
      RECT 10.086 2.973 10.172 3.169 ;
      RECT 10 2.968 10.086 3.153 ;
      RECT 9.97 2.965 10 3.14 ;
      RECT 9.945 2.964 9.97 3.128 ;
      RECT 9.94 2.964 9.945 3.118 ;
      RECT 9.9 2.963 9.94 3.11 ;
      RECT 9.885 2.962 9.9 3.103 ;
      RECT 9.835 2.961 9.885 3.095 ;
      RECT 9.833 2.96 9.835 3.09 ;
      RECT 9.747 2.958 9.833 3.09 ;
      RECT 9.661 2.953 9.747 3.09 ;
      RECT 9.575 2.949 9.661 3.09 ;
      RECT 9.526 2.945 9.575 3.088 ;
      RECT 9.44 2.942 9.526 3.083 ;
      RECT 9.417 2.939 9.44 3.079 ;
      RECT 9.331 2.936 9.417 3.074 ;
      RECT 9.245 2.932 9.331 3.065 ;
      RECT 9.22 2.925 9.245 3.06 ;
      RECT 9.16 2.89 9.22 3.057 ;
      RECT 9.14 2.815 9.16 3.054 ;
      RECT 9.135 2.757 9.14 3.053 ;
      RECT 9.11 2.697 9.135 3.052 ;
      RECT 9.035 2.575 9.11 3.048 ;
      RECT 9.025 2.575 9.035 3.04 ;
      RECT 9.01 2.575 9.025 3.03 ;
      RECT 8.995 2.575 9.01 3 ;
      RECT 8.98 2.575 8.995 2.945 ;
      RECT 8.965 2.575 8.98 2.883 ;
      RECT 8.94 2.575 8.965 2.808 ;
      RECT 8.935 2.575 8.94 2.758 ;
      RECT 10.28 2.12 10.3 2.429 ;
      RECT 10.266 2.122 10.315 2.426 ;
      RECT 10.266 2.127 10.335 2.417 ;
      RECT 10.18 2.125 10.315 2.411 ;
      RECT 10.18 2.133 10.37 2.394 ;
      RECT 10.145 2.135 10.37 2.393 ;
      RECT 10.115 2.143 10.37 2.384 ;
      RECT 10.105 2.148 10.39 2.37 ;
      RECT 10.145 2.138 10.39 2.37 ;
      RECT 10.145 2.141 10.4 2.358 ;
      RECT 10.115 2.143 10.41 2.345 ;
      RECT 10.115 2.147 10.42 2.288 ;
      RECT 10.105 2.152 10.425 2.203 ;
      RECT 10.266 2.12 10.3 2.426 ;
      RECT 10.145 7.855 10.315 8.305 ;
      RECT 10.2 6.075 10.37 8.025 ;
      RECT 10.145 5.015 10.315 6.245 ;
      RECT 9.705 2.223 9.71 2.435 ;
      RECT 9.58 2.22 9.595 2.435 ;
      RECT 9.045 2.25 9.115 2.435 ;
      RECT 8.93 2.25 8.965 2.43 ;
      RECT 10.051 2.552 10.07 2.746 ;
      RECT 9.965 2.507 10.051 2.747 ;
      RECT 9.955 2.46 9.965 2.749 ;
      RECT 9.95 2.44 9.955 2.75 ;
      RECT 9.93 2.405 9.95 2.751 ;
      RECT 9.915 2.355 9.93 2.752 ;
      RECT 9.895 2.292 9.915 2.753 ;
      RECT 9.885 2.255 9.895 2.754 ;
      RECT 9.87 2.244 9.885 2.755 ;
      RECT 9.865 2.236 9.87 2.753 ;
      RECT 9.855 2.235 9.865 2.745 ;
      RECT 9.825 2.232 9.855 2.724 ;
      RECT 9.75 2.227 9.825 2.669 ;
      RECT 9.735 2.223 9.75 2.615 ;
      RECT 9.725 2.223 9.735 2.51 ;
      RECT 9.71 2.223 9.725 2.443 ;
      RECT 9.695 2.223 9.705 2.433 ;
      RECT 9.64 2.222 9.695 2.43 ;
      RECT 9.595 2.22 9.64 2.433 ;
      RECT 9.567 2.22 9.58 2.436 ;
      RECT 9.481 2.224 9.567 2.438 ;
      RECT 9.395 2.23 9.481 2.443 ;
      RECT 9.375 2.234 9.395 2.445 ;
      RECT 9.373 2.235 9.375 2.444 ;
      RECT 9.287 2.237 9.373 2.443 ;
      RECT 9.201 2.242 9.287 2.44 ;
      RECT 9.115 2.247 9.201 2.437 ;
      RECT 8.965 2.25 9.045 2.433 ;
      RECT 9.625 5.015 9.795 8.305 ;
      RECT 9.625 7.315 10.03 7.645 ;
      RECT 9.625 6.475 10.03 6.805 ;
      RECT 9.741 3.225 9.79 3.559 ;
      RECT 9.741 3.225 9.795 3.558 ;
      RECT 9.655 3.225 9.795 3.557 ;
      RECT 9.43 3.333 9.8 3.555 ;
      RECT 9.655 3.225 9.825 3.548 ;
      RECT 9.625 3.237 9.83 3.539 ;
      RECT 9.61 3.255 9.835 3.536 ;
      RECT 9.425 3.339 9.835 3.463 ;
      RECT 9.42 3.346 9.835 3.423 ;
      RECT 9.435 3.312 9.835 3.536 ;
      RECT 9.596 3.258 9.8 3.555 ;
      RECT 9.51 3.278 9.835 3.536 ;
      RECT 9.61 3.252 9.83 3.539 ;
      RECT 9.38 2.576 9.57 2.77 ;
      RECT 9.375 2.578 9.57 2.769 ;
      RECT 9.37 2.582 9.585 2.766 ;
      RECT 9.385 2.575 9.585 2.766 ;
      RECT 9.37 2.685 9.59 2.761 ;
      RECT 8.665 3.185 8.756 3.483 ;
      RECT 8.66 3.187 8.835 3.478 ;
      RECT 8.665 3.185 8.835 3.478 ;
      RECT 8.66 3.191 8.855 3.476 ;
      RECT 8.66 3.246 8.895 3.475 ;
      RECT 8.66 3.281 8.91 3.469 ;
      RECT 8.66 3.315 8.92 3.459 ;
      RECT 8.65 3.195 8.855 3.31 ;
      RECT 8.65 3.215 8.87 3.31 ;
      RECT 8.65 3.198 8.86 3.31 ;
      RECT 8.875 1.966 8.88 2.028 ;
      RECT 8.87 1.888 8.875 2.051 ;
      RECT 8.865 1.845 8.87 2.062 ;
      RECT 8.86 1.835 8.865 2.074 ;
      RECT 8.855 1.835 8.86 2.083 ;
      RECT 8.83 1.835 8.855 2.115 ;
      RECT 8.825 1.835 8.83 2.148 ;
      RECT 8.81 1.835 8.825 2.173 ;
      RECT 8.8 1.835 8.81 2.2 ;
      RECT 8.795 1.835 8.8 2.213 ;
      RECT 8.79 1.835 8.795 2.228 ;
      RECT 8.78 1.835 8.79 2.243 ;
      RECT 8.775 1.835 8.78 2.263 ;
      RECT 8.75 1.835 8.775 2.298 ;
      RECT 8.705 1.835 8.75 2.343 ;
      RECT 8.695 1.835 8.705 2.356 ;
      RECT 8.61 1.92 8.695 2.363 ;
      RECT 8.575 2.042 8.61 2.372 ;
      RECT 8.57 2.082 8.575 2.376 ;
      RECT 8.55 2.105 8.57 2.378 ;
      RECT 8.545 2.135 8.55 2.381 ;
      RECT 8.535 2.147 8.545 2.382 ;
      RECT 8.49 2.17 8.535 2.387 ;
      RECT 8.45 2.2 8.49 2.395 ;
      RECT 8.415 2.212 8.45 2.401 ;
      RECT 8.41 2.217 8.415 2.405 ;
      RECT 8.34 2.227 8.41 2.412 ;
      RECT 8.3 2.237 8.34 2.422 ;
      RECT 8.28 2.242 8.3 2.428 ;
      RECT 8.27 2.246 8.28 2.433 ;
      RECT 8.265 2.249 8.27 2.436 ;
      RECT 8.255 2.25 8.265 2.437 ;
      RECT 8.23 2.252 8.255 2.441 ;
      RECT 8.22 2.257 8.23 2.444 ;
      RECT 8.175 2.265 8.22 2.445 ;
      RECT 8.05 2.27 8.175 2.445 ;
      RECT 8.605 2.567 8.625 2.749 ;
      RECT 8.556 2.552 8.605 2.748 ;
      RECT 8.47 2.567 8.625 2.746 ;
      RECT 8.455 2.567 8.625 2.745 ;
      RECT 8.42 2.545 8.59 2.73 ;
      RECT 8.49 3.565 8.505 3.774 ;
      RECT 8.49 3.573 8.51 3.773 ;
      RECT 8.435 3.573 8.51 3.772 ;
      RECT 8.415 3.577 8.515 3.77 ;
      RECT 8.395 3.527 8.435 3.769 ;
      RECT 8.34 3.585 8.52 3.767 ;
      RECT 8.305 3.542 8.435 3.765 ;
      RECT 8.301 3.545 8.49 3.764 ;
      RECT 8.215 3.553 8.49 3.762 ;
      RECT 8.215 3.597 8.525 3.755 ;
      RECT 8.205 3.69 8.525 3.753 ;
      RECT 8.215 3.609 8.53 3.738 ;
      RECT 8.215 3.63 8.545 3.708 ;
      RECT 8.215 3.657 8.55 3.678 ;
      RECT 8.34 3.535 8.435 3.767 ;
      RECT 7.97 2.58 7.975 3.118 ;
      RECT 7.775 2.91 7.78 3.105 ;
      RECT 6.075 2.575 6.09 2.955 ;
      RECT 8.14 2.575 8.145 2.745 ;
      RECT 8.135 2.575 8.14 2.755 ;
      RECT 8.13 2.575 8.135 2.768 ;
      RECT 8.105 2.575 8.13 2.81 ;
      RECT 8.08 2.575 8.105 2.883 ;
      RECT 8.065 2.575 8.08 2.935 ;
      RECT 8.06 2.575 8.065 2.965 ;
      RECT 8.035 2.575 8.06 3.005 ;
      RECT 8.02 2.575 8.035 3.06 ;
      RECT 8.015 2.575 8.02 3.093 ;
      RECT 7.99 2.575 8.015 3.113 ;
      RECT 7.975 2.575 7.99 3.119 ;
      RECT 7.905 2.61 7.97 3.115 ;
      RECT 7.855 2.665 7.905 3.11 ;
      RECT 7.845 2.697 7.855 3.108 ;
      RECT 7.84 2.722 7.845 3.108 ;
      RECT 7.82 2.795 7.84 3.108 ;
      RECT 7.81 2.875 7.82 3.107 ;
      RECT 7.795 2.905 7.81 3.107 ;
      RECT 7.78 2.91 7.795 3.106 ;
      RECT 7.72 2.912 7.775 3.103 ;
      RECT 7.69 2.917 7.72 3.099 ;
      RECT 7.688 2.92 7.69 3.098 ;
      RECT 7.602 2.922 7.688 3.095 ;
      RECT 7.516 2.928 7.602 3.089 ;
      RECT 7.43 2.933 7.516 3.083 ;
      RECT 7.357 2.938 7.43 3.084 ;
      RECT 7.271 2.944 7.357 3.092 ;
      RECT 7.185 2.95 7.271 3.101 ;
      RECT 7.165 2.954 7.185 3.106 ;
      RECT 7.118 2.956 7.165 3.109 ;
      RECT 7.032 2.961 7.118 3.115 ;
      RECT 6.946 2.966 7.032 3.124 ;
      RECT 6.86 2.972 6.946 3.132 ;
      RECT 6.775 2.97 6.86 3.141 ;
      RECT 6.771 2.965 6.775 3.145 ;
      RECT 6.685 2.96 6.771 3.137 ;
      RECT 6.621 2.951 6.685 3.125 ;
      RECT 6.535 2.942 6.621 3.112 ;
      RECT 6.511 2.935 6.535 3.103 ;
      RECT 6.425 2.929 6.511 3.09 ;
      RECT 6.385 2.922 6.425 3.076 ;
      RECT 6.38 2.912 6.385 3.072 ;
      RECT 6.37 2.9 6.38 3.071 ;
      RECT 6.35 2.87 6.37 3.068 ;
      RECT 6.295 2.79 6.35 3.062 ;
      RECT 6.275 2.709 6.295 3.057 ;
      RECT 6.255 2.667 6.275 3.053 ;
      RECT 6.23 2.62 6.255 3.047 ;
      RECT 6.225 2.595 6.23 3.044 ;
      RECT 6.19 2.575 6.225 3.039 ;
      RECT 6.181 2.575 6.19 3.032 ;
      RECT 6.095 2.575 6.181 3.002 ;
      RECT 6.09 2.575 6.095 2.965 ;
      RECT 6.055 2.575 6.075 2.887 ;
      RECT 6.05 2.617 6.055 2.852 ;
      RECT 6.045 2.692 6.05 2.808 ;
      RECT 7.495 2.497 7.67 2.745 ;
      RECT 7.495 2.497 7.675 2.743 ;
      RECT 7.49 2.529 7.675 2.703 ;
      RECT 7.52 2.47 7.69 2.69 ;
      RECT 7.485 2.547 7.69 2.623 ;
      RECT 6.795 2.01 6.965 2.185 ;
      RECT 6.795 2.01 7.137 2.177 ;
      RECT 6.795 2.01 7.22 2.171 ;
      RECT 6.795 2.01 7.255 2.167 ;
      RECT 6.795 2.01 7.275 2.166 ;
      RECT 6.795 2.01 7.361 2.162 ;
      RECT 7.255 1.835 7.425 2.157 ;
      RECT 6.83 1.942 7.455 2.155 ;
      RECT 6.82 1.997 7.46 2.153 ;
      RECT 6.795 2.033 7.47 2.148 ;
      RECT 6.795 2.06 7.475 2.078 ;
      RECT 6.86 1.885 7.435 2.155 ;
      RECT 7.051 1.87 7.435 2.155 ;
      RECT 6.885 1.873 7.435 2.155 ;
      RECT 6.965 1.871 7.051 2.182 ;
      RECT 7.051 1.868 7.43 2.155 ;
      RECT 7.235 1.845 7.43 2.155 ;
      RECT 7.137 1.866 7.43 2.155 ;
      RECT 7.22 1.86 7.235 2.168 ;
      RECT 7.37 3.225 7.375 3.425 ;
      RECT 6.835 3.29 6.88 3.425 ;
      RECT 7.405 3.225 7.425 3.398 ;
      RECT 7.375 3.225 7.405 3.413 ;
      RECT 7.31 3.225 7.37 3.45 ;
      RECT 7.295 3.225 7.31 3.48 ;
      RECT 7.28 3.225 7.295 3.493 ;
      RECT 7.26 3.225 7.28 3.508 ;
      RECT 7.255 3.225 7.26 3.517 ;
      RECT 7.245 3.229 7.255 3.522 ;
      RECT 7.23 3.239 7.245 3.533 ;
      RECT 7.205 3.255 7.23 3.543 ;
      RECT 7.195 3.269 7.205 3.545 ;
      RECT 7.175 3.281 7.195 3.542 ;
      RECT 7.145 3.302 7.175 3.536 ;
      RECT 7.135 3.314 7.145 3.531 ;
      RECT 7.125 3.312 7.135 3.528 ;
      RECT 7.11 3.311 7.125 3.523 ;
      RECT 7.105 3.31 7.11 3.518 ;
      RECT 7.07 3.308 7.105 3.508 ;
      RECT 7.05 3.305 7.07 3.49 ;
      RECT 7.04 3.303 7.05 3.485 ;
      RECT 7.03 3.302 7.04 3.48 ;
      RECT 6.995 3.3 7.03 3.468 ;
      RECT 6.94 3.296 6.995 3.448 ;
      RECT 6.93 3.294 6.94 3.433 ;
      RECT 6.925 3.294 6.93 3.428 ;
      RECT 6.88 3.292 6.925 3.425 ;
      RECT 6.785 3.29 6.835 3.429 ;
      RECT 6.775 3.291 6.785 3.434 ;
      RECT 6.715 3.298 6.775 3.448 ;
      RECT 6.69 3.306 6.715 3.468 ;
      RECT 6.68 3.31 6.69 3.48 ;
      RECT 6.675 3.311 6.68 3.485 ;
      RECT 6.66 3.313 6.675 3.488 ;
      RECT 6.645 3.315 6.66 3.493 ;
      RECT 6.64 3.315 6.645 3.496 ;
      RECT 6.595 3.32 6.64 3.507 ;
      RECT 6.59 3.324 6.595 3.519 ;
      RECT 6.565 3.32 6.59 3.523 ;
      RECT 6.555 3.316 6.565 3.527 ;
      RECT 6.545 3.315 6.555 3.531 ;
      RECT 6.53 3.305 6.545 3.537 ;
      RECT 6.525 3.293 6.53 3.541 ;
      RECT 6.52 3.29 6.525 3.542 ;
      RECT 6.515 3.287 6.52 3.544 ;
      RECT 6.5 3.275 6.515 3.543 ;
      RECT 6.485 3.257 6.5 3.54 ;
      RECT 6.465 3.236 6.485 3.533 ;
      RECT 6.4 3.225 6.465 3.505 ;
      RECT 6.396 3.225 6.4 3.484 ;
      RECT 6.31 3.225 6.396 3.454 ;
      RECT 6.295 3.225 6.31 3.41 ;
      RECT 6.87 2.325 6.875 2.56 ;
      RECT 6 2.241 6.005 2.445 ;
      RECT 6.58 2.27 6.585 2.425 ;
      RECT 6.5 2.25 6.505 2.425 ;
      RECT 7.17 2.392 7.185 2.745 ;
      RECT 7.096 2.377 7.17 2.745 ;
      RECT 7.01 2.36 7.096 2.745 ;
      RECT 7 2.35 7.01 2.743 ;
      RECT 6.995 2.348 7 2.738 ;
      RECT 6.98 2.346 6.995 2.724 ;
      RECT 6.91 2.338 6.98 2.664 ;
      RECT 6.89 2.329 6.91 2.598 ;
      RECT 6.885 2.326 6.89 2.578 ;
      RECT 6.875 2.325 6.885 2.568 ;
      RECT 6.865 2.325 6.87 2.552 ;
      RECT 6.855 2.324 6.865 2.542 ;
      RECT 6.845 2.322 6.855 2.53 ;
      RECT 6.83 2.319 6.845 2.51 ;
      RECT 6.82 2.317 6.83 2.495 ;
      RECT 6.8 2.314 6.82 2.483 ;
      RECT 6.795 2.312 6.8 2.473 ;
      RECT 6.77 2.31 6.795 2.46 ;
      RECT 6.74 2.305 6.77 2.445 ;
      RECT 6.66 2.296 6.74 2.436 ;
      RECT 6.615 2.285 6.66 2.429 ;
      RECT 6.595 2.276 6.615 2.426 ;
      RECT 6.585 2.271 6.595 2.425 ;
      RECT 6.54 2.265 6.58 2.425 ;
      RECT 6.525 2.257 6.54 2.425 ;
      RECT 6.505 2.252 6.525 2.425 ;
      RECT 6.485 2.249 6.5 2.425 ;
      RECT 6.402 2.248 6.485 2.424 ;
      RECT 6.316 2.247 6.402 2.42 ;
      RECT 6.23 2.245 6.316 2.417 ;
      RECT 6.177 2.244 6.23 2.419 ;
      RECT 6.091 2.243 6.177 2.428 ;
      RECT 6.005 2.242 6.091 2.44 ;
      RECT 5.985 2.241 6 2.448 ;
      RECT 5.905 2.24 5.985 2.46 ;
      RECT 5.88 2.24 5.905 2.473 ;
      RECT 5.855 2.24 5.88 2.488 ;
      RECT 5.85 2.24 5.855 2.51 ;
      RECT 5.845 2.24 5.85 2.528 ;
      RECT 5.84 2.24 5.845 2.545 ;
      RECT 5.835 2.24 5.84 2.558 ;
      RECT 5.83 2.24 5.835 2.568 ;
      RECT 5.79 2.24 5.83 2.653 ;
      RECT 5.775 2.24 5.79 2.738 ;
      RECT 5.765 2.241 5.775 2.75 ;
      RECT 5.73 2.246 5.765 2.755 ;
      RECT 5.69 2.255 5.73 2.755 ;
      RECT 5.675 2.265 5.69 2.755 ;
      RECT 5.67 2.275 5.675 2.755 ;
      RECT 5.65 2.302 5.67 2.755 ;
      RECT 5.6 2.385 5.65 2.755 ;
      RECT 5.595 2.447 5.6 2.755 ;
      RECT 5.585 2.46 5.595 2.755 ;
      RECT 5.575 2.482 5.585 2.755 ;
      RECT 5.565 2.507 5.575 2.75 ;
      RECT 5.56 2.545 5.565 2.743 ;
      RECT 5.55 2.655 5.56 2.738 ;
      RECT 6.945 3.576 6.96 3.835 ;
      RECT 6.945 3.591 6.965 3.834 ;
      RECT 6.861 3.591 6.965 3.832 ;
      RECT 6.861 3.605 6.97 3.831 ;
      RECT 6.775 3.647 6.975 3.828 ;
      RECT 6.77 3.59 6.96 3.823 ;
      RECT 6.77 3.661 6.98 3.82 ;
      RECT 6.765 3.692 6.98 3.818 ;
      RECT 6.77 3.689 6.995 3.808 ;
      RECT 6.765 3.735 7.01 3.793 ;
      RECT 6.765 3.763 7.015 3.778 ;
      RECT 6.775 3.565 6.945 3.828 ;
      RECT 6.535 2.575 6.705 2.745 ;
      RECT 6.5 2.575 6.705 2.74 ;
      RECT 6.49 2.575 6.705 2.733 ;
      RECT 6.485 2.56 6.655 2.73 ;
      RECT 5.315 3.097 5.58 3.54 ;
      RECT 5.31 3.068 5.525 3.538 ;
      RECT 5.305 3.222 5.585 3.533 ;
      RECT 5.31 3.117 5.585 3.533 ;
      RECT 5.31 3.128 5.595 3.52 ;
      RECT 5.31 3.075 5.555 3.538 ;
      RECT 5.315 3.062 5.525 3.54 ;
      RECT 5.315 3.06 5.475 3.54 ;
      RECT 5.416 3.052 5.475 3.54 ;
      RECT 5.33 3.053 5.475 3.54 ;
      RECT 5.416 3.051 5.465 3.54 ;
      RECT 5.22 1.866 5.395 2.165 ;
      RECT 5.27 1.828 5.395 2.165 ;
      RECT 5.255 1.83 5.481 2.157 ;
      RECT 5.255 1.833 5.52 2.144 ;
      RECT 5.255 1.834 5.53 2.13 ;
      RECT 5.21 1.885 5.53 2.12 ;
      RECT 5.255 1.835 5.535 2.115 ;
      RECT 5.21 2.045 5.54 2.105 ;
      RECT 5.195 1.905 5.535 2.045 ;
      RECT 5.19 1.921 5.535 1.985 ;
      RECT 5.235 1.845 5.535 2.115 ;
      RECT 5.27 1.826 5.356 2.165 ;
      RECT 2.65 7.855 2.82 8.305 ;
      RECT 2.705 6.075 2.875 8.025 ;
      RECT 2.65 5.015 2.82 6.245 ;
      RECT 2.13 5.015 2.3 8.305 ;
      RECT 2.13 7.315 2.535 7.645 ;
      RECT 2.13 6.475 2.535 6.805 ;
      RECT 80.03 7.8 80.2 8.31 ;
      RECT 79.04 0.57 79.21 1.08 ;
      RECT 79.04 2.39 79.21 3.86 ;
      RECT 79.04 5.02 79.21 6.49 ;
      RECT 79.04 7.8 79.21 8.31 ;
      RECT 77.68 0.575 77.85 3.865 ;
      RECT 77.68 5.015 77.85 8.305 ;
      RECT 77.25 0.575 77.42 1.085 ;
      RECT 77.25 1.655 77.42 3.865 ;
      RECT 77.25 5.015 77.42 7.225 ;
      RECT 77.25 7.795 77.42 8.305 ;
      RECT 72.045 5.015 72.215 8.305 ;
      RECT 71.615 5.015 71.785 7.225 ;
      RECT 71.615 7.795 71.785 8.305 ;
      RECT 64.77 7.8 64.94 8.31 ;
      RECT 63.78 0.57 63.95 1.08 ;
      RECT 63.78 2.39 63.95 3.86 ;
      RECT 63.78 5.02 63.95 6.49 ;
      RECT 63.78 7.8 63.95 8.31 ;
      RECT 62.42 0.575 62.59 3.865 ;
      RECT 62.42 5.015 62.59 8.305 ;
      RECT 61.99 0.575 62.16 1.085 ;
      RECT 61.99 1.655 62.16 3.865 ;
      RECT 61.99 5.015 62.16 7.225 ;
      RECT 61.99 7.795 62.16 8.305 ;
      RECT 56.785 5.015 56.955 8.305 ;
      RECT 56.355 5.015 56.525 7.225 ;
      RECT 56.355 7.795 56.525 8.305 ;
      RECT 49.51 7.8 49.68 8.31 ;
      RECT 48.52 0.57 48.69 1.08 ;
      RECT 48.52 2.39 48.69 3.86 ;
      RECT 48.52 5.02 48.69 6.49 ;
      RECT 48.52 7.8 48.69 8.31 ;
      RECT 47.16 0.575 47.33 3.865 ;
      RECT 47.16 5.015 47.33 8.305 ;
      RECT 46.73 0.575 46.9 1.085 ;
      RECT 46.73 1.655 46.9 3.865 ;
      RECT 46.73 5.015 46.9 7.225 ;
      RECT 46.73 7.795 46.9 8.305 ;
      RECT 41.525 5.015 41.695 8.305 ;
      RECT 41.095 5.015 41.265 7.225 ;
      RECT 41.095 7.795 41.265 8.305 ;
      RECT 34.25 7.8 34.42 8.31 ;
      RECT 33.26 0.57 33.43 1.08 ;
      RECT 33.26 2.39 33.43 3.86 ;
      RECT 33.26 5.02 33.43 6.49 ;
      RECT 33.26 7.8 33.43 8.31 ;
      RECT 31.9 0.575 32.07 3.865 ;
      RECT 31.9 5.015 32.07 8.305 ;
      RECT 31.47 0.575 31.64 1.085 ;
      RECT 31.47 1.655 31.64 3.865 ;
      RECT 31.47 5.015 31.64 7.225 ;
      RECT 31.47 7.795 31.64 8.305 ;
      RECT 26.265 5.015 26.435 8.305 ;
      RECT 25.835 5.015 26.005 7.225 ;
      RECT 25.835 7.795 26.005 8.305 ;
      RECT 18.99 7.8 19.16 8.31 ;
      RECT 18 0.57 18.17 1.08 ;
      RECT 18 2.39 18.17 3.86 ;
      RECT 18 5.02 18.17 6.49 ;
      RECT 18 7.8 18.17 8.31 ;
      RECT 16.64 0.575 16.81 3.865 ;
      RECT 16.64 5.015 16.81 8.305 ;
      RECT 16.21 0.575 16.38 1.085 ;
      RECT 16.21 1.655 16.38 3.865 ;
      RECT 16.21 5.015 16.38 7.225 ;
      RECT 16.21 7.795 16.38 8.305 ;
      RECT 11.005 5.015 11.175 8.305 ;
      RECT 10.575 5.015 10.745 7.225 ;
      RECT 10.575 7.795 10.745 8.305 ;
      RECT 3.08 5.015 3.25 7.225 ;
      RECT 3.08 7.795 3.25 8.305 ;
  END
END sky130_osu_ring_oscillator_mpr2ya_8_b0r2

END LIBRARY
