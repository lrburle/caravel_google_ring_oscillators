magic
tech sky130A
magscale 1 2
timestamp 1713455822
<< nwell >>
rect 5002 1407 7635 1749
rect 9588 1636 9646 1694
rect 12640 1636 12698 1694
rect 15692 1636 15750 1694
rect 18744 1636 18802 1694
rect 5000 1087 20819 1407
rect 5000 1019 7635 1087
rect 5002 820 7635 1019
rect 8490 985 8548 1043
rect 11542 985 11600 1043
rect 14594 985 14652 1043
rect 17646 985 17704 1043
rect 20698 985 20756 1043
<< ndiff >>
rect 8501 441 8536 475
rect 11553 441 11588 475
rect 14605 441 14640 475
rect 17657 441 17692 475
rect 20709 441 20744 475
<< pdiff >>
rect 5045 1648 5079 1682
rect 6536 1636 6594 1694
rect 9588 1636 9646 1694
rect 12640 1636 12698 1694
rect 15692 1636 15750 1694
rect 18744 1636 18802 1694
<< locali >>
rect 0 2173 20819 2493
rect 5406 1407 5440 1477
rect 0 1087 20819 1407
rect 0 0 20819 320
<< viali >>
rect 5045 1648 5079 1682
rect 8502 441 8536 475
rect 11554 441 11588 475
rect 14606 441 14640 475
rect 17658 441 17692 475
rect 20710 441 20744 475
<< metal1 >>
rect 0 2173 20819 2493
rect 20741 1983 20745 2012
rect 20705 1977 20775 1983
rect 5302 1863 5308 1921
rect 5366 1863 5372 1921
rect 20705 1919 20711 1977
rect 20769 1919 20775 1977
rect 20705 1913 20775 1919
rect 8501 1854 8571 1860
rect 6937 1843 7007 1849
rect 6937 1785 6943 1843
rect 7001 1785 7007 1843
rect 8501 1796 8507 1854
rect 8565 1796 8571 1854
rect 11552 1854 11623 1861
rect 8501 1790 8571 1796
rect 9989 1845 10059 1851
rect 6937 1779 7007 1785
rect 9989 1787 9995 1845
rect 10053 1787 10059 1845
rect 11552 1796 11559 1854
rect 11617 1796 11623 1854
rect 14596 1854 14666 1860
rect 11552 1790 11623 1796
rect 13041 1845 13111 1851
rect 9989 1781 10059 1787
rect 13041 1787 13047 1845
rect 13105 1787 13111 1845
rect 14596 1796 14602 1854
rect 14660 1796 14666 1854
rect 17648 1854 17718 1860
rect 14596 1790 14666 1796
rect 16094 1845 16164 1851
rect 13041 1781 13111 1787
rect 16094 1787 16100 1845
rect 16158 1787 16164 1845
rect 17648 1796 17654 1854
rect 17712 1796 17718 1854
rect 17648 1790 17718 1796
rect 19145 1845 19215 1851
rect 16094 1781 16164 1787
rect 19145 1787 19151 1845
rect 19209 1787 19215 1845
rect 19145 1781 19215 1787
rect 5227 1715 5233 1773
rect 5291 1715 5297 1773
rect 5034 1682 5092 1687
rect 5034 1648 5045 1682
rect 5079 1648 5092 1682
rect 5034 1641 5092 1648
rect 0 1087 20819 1407
rect 0 0 20819 320
<< via1 >>
rect 5308 1863 5366 1921
rect 20711 1919 20769 1977
rect 6943 1785 7001 1843
rect 8507 1796 8565 1854
rect 9995 1787 10053 1845
rect 11559 1796 11617 1854
rect 13047 1787 13105 1845
rect 14602 1796 14660 1854
rect 16100 1787 16158 1845
rect 17654 1796 17712 1854
rect 19151 1787 19209 1845
rect 5233 1715 5291 1773
rect 6536 1636 6594 1694
rect 9588 1636 9646 1694
rect 12640 1636 12698 1694
rect 15692 1636 15750 1694
rect 18744 1636 18802 1694
rect 8490 985 8548 1043
rect 11542 985 11600 1043
rect 14594 985 14652 1043
rect 17646 985 17704 1043
rect 20698 985 20756 1043
<< metal2 >>
rect 5246 2138 20745 2172
rect 5246 1779 5280 2138
rect 20711 1983 20745 2138
rect 20705 1977 20775 1983
rect 5308 1921 5366 1927
rect 20705 1919 20711 1977
rect 20769 1919 20775 1977
rect 20705 1913 20775 1919
rect 5366 1868 5559 1902
rect 5308 1857 5366 1863
rect 5525 1829 5559 1868
rect 8501 1854 8571 1860
rect 6937 1843 7007 1849
rect 6937 1829 6943 1843
rect 5525 1795 6943 1829
rect 6937 1785 6943 1795
rect 7001 1785 7007 1843
rect 8501 1796 8507 1854
rect 8565 1836 8571 1854
rect 11553 1854 11623 1860
rect 9989 1845 10059 1851
rect 9989 1836 9995 1845
rect 8565 1796 9995 1836
rect 8501 1790 8571 1796
rect 6937 1779 7007 1785
rect 9989 1787 9995 1796
rect 10053 1787 10059 1845
rect 11553 1796 11559 1854
rect 11617 1836 11623 1854
rect 14596 1854 14666 1860
rect 13041 1845 13111 1851
rect 13041 1836 13047 1845
rect 11617 1796 13047 1836
rect 11553 1790 11623 1796
rect 9989 1781 10059 1787
rect 13041 1787 13047 1796
rect 13105 1787 13111 1845
rect 14596 1796 14602 1854
rect 14660 1836 14666 1854
rect 17648 1854 17718 1860
rect 16094 1845 16164 1851
rect 16094 1836 16100 1845
rect 14660 1796 16100 1836
rect 14596 1790 14666 1796
rect 13041 1781 13111 1787
rect 16094 1787 16100 1796
rect 16158 1787 16164 1845
rect 17648 1796 17654 1854
rect 17712 1836 17718 1854
rect 19145 1845 19215 1851
rect 19145 1836 19151 1845
rect 17712 1796 19151 1836
rect 17648 1790 17718 1796
rect 16094 1781 16164 1787
rect 19145 1787 19151 1796
rect 19209 1787 19215 1845
rect 19145 1781 19215 1787
rect 5233 1773 5291 1779
rect 5233 1709 5291 1715
<< via2 >>
rect 6536 1636 6594 1694
rect 9588 1636 9646 1694
rect 12640 1636 12698 1694
rect 15692 1636 15750 1694
rect 18744 1636 18802 1694
rect 8490 985 8548 1043
rect 11542 985 11600 1043
rect 14594 985 14652 1043
rect 17646 985 17704 1043
rect 20698 985 20756 1043
<< metal3 >>
rect 6530 1694 6600 2493
rect 9582 1694 9652 2493
rect 12634 1694 12704 2493
rect 15686 1694 15756 2493
rect 18738 1694 18808 2493
rect 8481 0 8557 985
rect 11533 0 11609 985
rect 14585 0 14661 985
rect 17637 0 17713 985
rect 20689 0 20765 985
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_0
timestamp 1713287902
transform 1 0 5009 0 -1 2234
box -10 0 552 902
use sky130_osu_single_mpr2xa_8_b0r2  sky130_osu_single_mpr2xa_8_b0r2_0
timestamp 1713454888
transform 1 0 17767 0 1 0
box 0 0 3052 2493
use sky130_osu_single_mpr2xa_8_b0r2  sky130_osu_single_mpr2xa_8_b0r2_1
timestamp 1713454888
transform 1 0 5559 0 1 0
box 0 0 3052 2493
use sky130_osu_single_mpr2xa_8_b0r2  sky130_osu_single_mpr2xa_8_b0r2_2
timestamp 1713454888
transform 1 0 8611 0 1 0
box 0 0 3052 2493
use sky130_osu_single_mpr2xa_8_b0r2  sky130_osu_single_mpr2xa_8_b0r2_3
timestamp 1713454888
transform 1 0 11663 0 1 0
box 0 0 3052 2493
use sky130_osu_single_mpr2xa_8_b0r2  sky130_osu_single_mpr2xa_8_b0r2_4
timestamp 1713454888
transform 1 0 14715 0 1 0
box 0 0 3052 2493
<< labels >>
flabel metal1 s 5034 1641 5092 1687 0 FreeSans 100 0 0 0 start
port 13 nsew signal input
flabel metal3 s 8502 441 8536 475 0 FreeSans 100 0 0 0 X1_Y1
port 6 se signal output
flabel metal3 s 11554 441 11588 475 0 FreeSans 100 0 0 0 X2_Y1
port 7 se signal output
flabel metal3 s 14606 441 14640 475 0 FreeSans 100 0 0 0 X3_Y1
port 8 se signal output
flabel metal3 s 17658 441 17692 475 0 FreeSans 100 0 0 0 X4_Y1
port 9 se signal output
flabel metal3 s 20710 441 20744 475 0 FreeSans 100 0 0 0 X5_Y1
port 10 se signal output
flabel metal1 s 0 2173 20819 2493 0 FreeSans 100 0 0 0 vssd1
port 14 nsew ground bidirectional
flabel metal1 s 0 1087 20819 1407 0 FreeSans 100 0 0 0 vccd1
port 15 nsew power bidirectional
flabel metal1 s 0 0 20819 320 0 FreeSans 100 0 0 0 vssd1
port 14 nsew ground bidirectional
flabel metal1 s 6548 1648 6582 1682 0 FreeSans 100 0 0 0 s1
port 1 nw signal input
flabel metal1 s 9600 1648 9634 1682 0 FreeSans 100 0 0 0 s2
port 2 nw signal input
flabel metal1 s 12652 1648 12686 1682 0 FreeSans 100 0 0 0 s3
port 3 nw signal input
flabel metal1 s 15704 1648 15738 1682 0 FreeSans 100 0 0 0 s4
port 4 nw signal input
flabel metal1 s 18756 1648 18790 1682 0 FreeSans 100 0 0 0 s5
port 5 nw signal input
<< end >>
