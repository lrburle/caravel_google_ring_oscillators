magic
tech sky130A
magscale 1 2
timestamp 1708619673
<< error_s >>
rect 3118 2103 3119 2114
rect 3308 2103 3309 2114
rect 3394 2103 3395 2114
rect 4896 2103 4897 2114
rect 5086 2103 5087 2114
rect 5172 2103 5173 2114
rect 5852 2103 5853 2114
rect 6042 2103 6043 2114
rect 6128 2103 6129 2114
rect 6401 2103 6402 2114
rect 3129 2063 3130 2103
rect 3319 2063 3320 2103
rect 3405 2063 3406 2103
rect 4907 2063 4908 2103
rect 5097 2063 5098 2103
rect 5183 2063 5184 2103
rect 5863 2063 5864 2103
rect 6053 2063 6054 2103
rect 6139 2063 6140 2103
rect 6412 2063 6413 2103
rect 6600 2102 6601 2113
rect 8052 2103 8053 2114
rect 8242 2103 8243 2114
rect 8328 2103 8329 2114
rect 9008 2103 9009 2114
rect 9198 2103 9199 2114
rect 9284 2103 9285 2114
rect 9557 2103 9558 2114
rect 6611 2062 6612 2102
rect 8063 2063 8064 2103
rect 8253 2063 8254 2103
rect 8339 2063 8340 2103
rect 9019 2063 9020 2103
rect 9209 2063 9210 2103
rect 9295 2063 9296 2103
rect 9568 2063 9569 2103
rect 9756 2102 9757 2113
rect 11207 2103 11208 2114
rect 11397 2103 11398 2114
rect 11483 2103 11484 2114
rect 12163 2103 12164 2114
rect 12353 2103 12354 2114
rect 12439 2103 12440 2114
rect 12712 2103 12713 2114
rect 9767 2062 9768 2102
rect 11218 2063 11219 2103
rect 11408 2063 11409 2103
rect 11494 2063 11495 2103
rect 12174 2063 12175 2103
rect 12364 2063 12365 2103
rect 12450 2063 12451 2103
rect 12723 2063 12724 2103
rect 12911 2102 12912 2113
rect 14364 2103 14365 2114
rect 14554 2103 14555 2114
rect 14640 2103 14641 2114
rect 15320 2103 15321 2114
rect 15510 2103 15511 2114
rect 15596 2103 15597 2114
rect 15869 2103 15870 2114
rect 12922 2062 12923 2102
rect 14375 2063 14376 2103
rect 14565 2063 14566 2103
rect 14651 2063 14652 2103
rect 15331 2063 15332 2103
rect 15521 2063 15522 2103
rect 15607 2063 15608 2103
rect 15880 2063 15881 2103
rect 16068 2102 16069 2113
rect 17521 2103 17522 2114
rect 17711 2103 17712 2114
rect 17797 2103 17798 2114
rect 18477 2103 18478 2114
rect 18667 2103 18668 2114
rect 18753 2103 18754 2114
rect 19026 2103 19027 2114
rect 16079 2062 16080 2102
rect 17532 2063 17533 2103
rect 17722 2063 17723 2103
rect 17808 2063 17809 2103
rect 18488 2063 18489 2103
rect 18678 2063 18679 2103
rect 18764 2063 18765 2103
rect 19037 2063 19038 2103
rect 19225 2102 19226 2113
rect 19236 2062 19237 2102
rect 6060 1936 6087 1943
rect 9216 1936 9243 1943
rect 12371 1936 12398 1943
rect 15528 1936 15555 1943
rect 18685 1936 18712 1943
rect 6060 1915 6128 1936
rect 9216 1915 9284 1936
rect 12371 1915 12439 1936
rect 15528 1915 15596 1936
rect 18685 1915 18753 1936
rect 6060 1909 6115 1915
rect 9216 1909 9271 1915
rect 12371 1909 12426 1915
rect 15528 1909 15583 1915
rect 18685 1909 18740 1915
rect 6099 1908 6100 1909
rect 9255 1908 9256 1909
rect 12410 1908 12411 1909
rect 15567 1908 15568 1909
rect 18724 1908 18725 1909
rect 6072 1902 6127 1908
rect 9228 1902 9283 1908
rect 12383 1902 12438 1908
rect 15540 1902 15595 1908
rect 18697 1902 18752 1908
rect 6099 1880 6100 1902
rect 9255 1880 9256 1902
rect 12410 1880 12411 1902
rect 15567 1880 15568 1902
rect 18724 1880 18725 1902
rect 4949 1754 4971 1783
rect 4977 1754 4999 1755
rect 8105 1754 8127 1783
rect 8133 1754 8155 1755
rect 11260 1754 11282 1783
rect 11288 1754 11310 1755
rect 14417 1754 14439 1783
rect 14445 1754 14467 1755
rect 17574 1754 17596 1783
rect 17602 1754 17624 1755
rect 2999 1470 3001 1749
rect 2999 1425 3000 1470
rect 3035 1461 3037 1713
rect 3118 1673 3119 1684
rect 3308 1673 3309 1684
rect 3394 1673 3395 1684
rect 4896 1673 4897 1684
rect 5086 1673 5087 1684
rect 5172 1673 5173 1684
rect 5852 1673 5853 1684
rect 6042 1673 6043 1684
rect 6128 1673 6129 1684
rect 6401 1673 6402 1684
rect 3129 1477 3130 1673
rect 3319 1477 3320 1673
rect 3405 1477 3406 1673
rect 4842 1641 4869 1647
rect 4870 1646 4897 1647
rect 3439 1466 3440 1495
rect 4907 1477 4908 1673
rect 5097 1477 5098 1673
rect 5183 1477 5184 1673
rect 5863 1477 5864 1673
rect 6053 1477 6054 1673
rect 6139 1477 6140 1673
rect 6412 1477 6413 1673
rect 6600 1672 6601 1683
rect 8052 1673 8053 1684
rect 8242 1673 8243 1684
rect 8328 1673 8329 1684
rect 9008 1673 9009 1684
rect 9198 1673 9199 1684
rect 9284 1673 9285 1684
rect 9557 1673 9558 1684
rect 6611 1476 6612 1672
rect 7998 1641 8025 1647
rect 8026 1646 8053 1647
rect 8063 1477 8064 1673
rect 8253 1477 8254 1673
rect 8339 1477 8340 1673
rect 9019 1477 9020 1673
rect 9209 1477 9210 1673
rect 9295 1477 9296 1673
rect 9568 1477 9569 1673
rect 9756 1672 9757 1683
rect 11207 1673 11208 1684
rect 11397 1673 11398 1684
rect 11483 1673 11484 1684
rect 12163 1673 12164 1684
rect 12353 1673 12354 1684
rect 12439 1673 12440 1684
rect 12712 1673 12713 1684
rect 9767 1476 9768 1672
rect 11153 1641 11180 1647
rect 11181 1646 11208 1647
rect 11218 1477 11219 1673
rect 11408 1477 11409 1673
rect 11494 1477 11495 1673
rect 12174 1477 12175 1673
rect 12364 1477 12365 1673
rect 12450 1477 12451 1673
rect 12723 1477 12724 1673
rect 12911 1672 12912 1683
rect 14364 1673 14365 1684
rect 14554 1673 14555 1684
rect 14640 1673 14641 1684
rect 15320 1673 15321 1684
rect 15510 1673 15511 1684
rect 15596 1673 15597 1684
rect 15869 1673 15870 1684
rect 12922 1476 12923 1672
rect 14310 1641 14337 1647
rect 14338 1646 14365 1647
rect 14375 1477 14376 1673
rect 14565 1477 14566 1673
rect 14651 1477 14652 1673
rect 15331 1477 15332 1673
rect 15521 1477 15522 1673
rect 15607 1477 15608 1673
rect 15880 1477 15881 1673
rect 16068 1672 16069 1683
rect 17521 1673 17522 1684
rect 17711 1673 17712 1684
rect 17797 1673 17798 1684
rect 18477 1673 18478 1684
rect 18667 1673 18668 1684
rect 18753 1673 18754 1684
rect 19026 1673 19027 1684
rect 16079 1476 16080 1672
rect 17467 1641 17494 1647
rect 17495 1646 17522 1647
rect 17532 1477 17533 1673
rect 17722 1477 17723 1673
rect 17808 1477 17809 1673
rect 18488 1477 18489 1673
rect 18678 1477 18679 1673
rect 18764 1477 18765 1673
rect 19037 1477 19038 1673
rect 19225 1672 19226 1683
rect 19236 1476 19237 1672
rect 3443 1373 3467 1407
rect 5221 1373 5245 1407
rect 6177 1373 6201 1407
rect 8377 1373 8401 1407
rect 9333 1373 9357 1407
rect 11532 1373 11556 1407
rect 12488 1373 12512 1407
rect 14689 1373 14713 1407
rect 15645 1373 15669 1407
rect 17846 1373 17870 1407
rect 18802 1373 18826 1407
rect 6177 1085 6201 1119
rect 6672 1085 6703 1086
rect 6706 1085 6737 1086
rect 9333 1085 9357 1119
rect 9827 1085 9859 1086
rect 9861 1085 9893 1086
rect 12488 1085 12512 1119
rect 12984 1085 13017 1086
rect 13018 1085 13048 1086
rect 15645 1085 15669 1119
rect 16141 1085 16174 1086
rect 16175 1085 16205 1086
rect 18802 1085 18826 1119
rect 4929 1037 5072 1039
rect 8085 1037 8228 1039
rect 11240 1037 11383 1039
rect 14397 1037 14540 1039
rect 17554 1037 17697 1039
rect 3870 1023 3971 1034
rect 4157 1033 4421 1034
rect 4421 1023 4476 1033
rect 4579 1027 4588 1036
rect 4626 1027 4635 1036
rect 4929 1034 5051 1037
rect 4901 1033 4918 1034
rect 4731 1027 4901 1033
rect 3855 1021 3870 1023
rect 3849 1019 3855 1021
rect 4478 1019 4483 1021
rect 3845 1014 3849 1019
rect 4483 1014 4490 1019
rect 4570 1018 4579 1027
rect 4635 1024 4731 1027
rect 5072 1023 5180 1037
rect 4930 1015 4946 1022
rect 4948 1015 4964 1022
rect 4490 1007 4502 1014
rect 4920 1013 4932 1015
rect 4942 1013 4954 1015
rect 4960 1013 4964 1015
rect 5148 1013 5164 1022
rect 5180 1021 5198 1023
rect 5199 1017 5206 1020
rect 5206 1013 5212 1017
rect 5852 1015 5853 1026
rect 6042 1015 6043 1026
rect 6128 1015 6129 1026
rect 6401 1015 6402 1026
rect 6599 1016 6600 1027
rect 7026 1023 7127 1034
rect 7313 1033 7577 1034
rect 7577 1023 7632 1033
rect 7735 1027 7744 1036
rect 7782 1027 7791 1036
rect 8085 1034 8207 1037
rect 8057 1033 8074 1034
rect 7887 1027 8057 1033
rect 7011 1021 7026 1023
rect 7005 1019 7011 1021
rect 7634 1019 7639 1021
rect 4920 1008 4964 1013
rect 5107 1008 5144 1009
rect 5212 1008 5215 1013
rect 4916 1006 4918 1008
rect 4920 1006 5052 1008
rect 3971 1005 4325 1006
rect 3951 1003 3969 1005
rect 4411 1003 4424 1005
rect 4503 1003 4506 1005
rect 4914 1003 5052 1006
rect 3895 1000 3951 1003
rect 3769 992 3781 1000
rect 3791 992 3803 1000
rect 3867 994 3951 1000
rect 4424 994 4434 1003
rect 3867 993 3895 994
rect 3765 989 3767 992
rect 3867 991 3886 993
rect 4435 991 4438 993
rect 3807 988 3811 989
rect 3757 977 3765 988
rect 3768 986 3803 988
rect 3766 977 3768 983
rect 3757 976 3766 977
rect 3765 972 3766 976
rect 3764 971 3765 972
rect 3762 966 3764 969
rect 3637 964 3702 965
rect 3629 956 3637 964
rect 3702 956 3706 964
rect 3628 950 3629 956
rect 3757 954 3765 966
rect 3769 956 3771 986
rect 3800 985 3803 986
rect 3802 979 3803 985
rect 3807 981 3815 988
rect 3811 980 3819 981
rect 3843 980 3844 990
rect 3867 980 3882 991
rect 4141 981 4178 983
rect 3819 979 3825 980
rect 3842 979 3843 980
rect 3867 979 3874 980
rect 3825 969 3887 979
rect 3895 972 3901 978
rect 3941 972 3947 978
rect 4141 977 4167 981
rect 4178 977 4183 981
rect 4438 980 4451 991
rect 4414 979 4428 980
rect 4135 972 4141 977
rect 4183 972 4192 977
rect 4396 972 4414 979
rect 4428 977 4435 979
rect 4506 977 4527 1003
rect 4908 996 5052 1003
rect 5068 1006 5169 1008
rect 5068 996 5180 1006
rect 4869 990 4930 996
rect 4834 987 4869 990
rect 4647 981 4834 987
rect 4920 986 4930 990
rect 4435 972 4450 977
rect 3889 969 3895 972
rect 3896 970 3953 972
rect 4192 971 4193 972
rect 4030 970 4033 971
rect 4051 970 4054 971
rect 4133 970 4134 971
rect 4193 970 4196 971
rect 3896 969 3904 970
rect 3867 968 3904 969
rect 3769 954 3803 956
rect 3758 951 3760 954
rect 3754 939 3758 950
rect 3769 942 3781 950
rect 3794 945 3803 954
rect 3841 952 3842 955
rect 3867 951 3872 968
rect 3889 966 3904 968
rect 3947 966 3953 970
rect 4026 967 4030 970
rect 4054 967 4059 970
rect 4196 968 4197 970
rect 4388 969 4396 972
rect 4425 971 4450 972
rect 4459 971 4463 972
rect 4421 970 4425 971
rect 4435 970 4472 971
rect 4197 967 4200 968
rect 3895 964 3904 966
rect 3895 951 3900 964
rect 3948 955 3967 958
rect 4002 955 4026 967
rect 4059 959 4077 967
rect 4132 959 4133 967
rect 3804 948 3814 950
rect 3814 947 3817 948
rect 3819 945 3828 947
rect 3792 942 3794 945
rect 3828 943 3839 945
rect 3840 943 3841 951
rect 3867 943 3873 951
rect 3791 939 3792 942
rect 3839 938 3873 943
rect 3705 924 3706 938
rect 3655 915 3664 924
rect 3702 920 3711 924
rect 3702 915 3716 920
rect 3646 912 3655 915
rect 3646 911 3649 912
rect 3639 908 3648 911
rect 3627 907 3648 908
rect 3627 905 3645 907
rect 3685 905 3691 911
rect 3705 906 3720 915
rect 3745 908 3754 937
rect 3627 900 3639 905
rect 3623 898 3626 900
rect 3627 899 3628 900
rect 3633 899 3639 900
rect 3691 899 3697 905
rect 3704 904 3716 906
rect 3743 904 3745 908
rect 3783 907 3791 938
rect 3840 926 3841 938
rect 3867 935 3895 938
rect 3867 931 3897 935
rect 3899 931 3900 951
rect 3967 946 4029 955
rect 4077 952 4085 959
rect 4131 951 4132 958
rect 4200 954 4204 967
rect 4380 966 4388 969
rect 4418 968 4421 970
rect 4414 967 4418 968
rect 4409 965 4414 967
rect 4435 965 4450 970
rect 4459 969 4463 970
rect 4472 969 4473 970
rect 4529 969 4534 975
rect 4570 971 4579 980
rect 4635 978 4647 981
rect 4635 971 4644 978
rect 4914 972 4930 986
rect 4953 972 4954 996
rect 4959 991 4980 996
rect 4964 990 4980 991
rect 5097 989 5103 996
rect 5149 989 5155 996
rect 5169 990 5180 996
rect 5215 990 5224 1008
rect 4964 972 4980 988
rect 5097 985 5105 989
rect 5103 983 5105 985
rect 5013 974 5041 978
rect 5043 974 5054 978
rect 4463 965 4468 969
rect 4473 965 4475 968
rect 4534 965 4537 969
rect 4375 964 4379 965
rect 4450 964 4453 965
rect 4475 964 4476 965
rect 4371 962 4375 964
rect 4340 950 4371 962
rect 4455 959 4459 962
rect 4470 960 4474 963
rect 4579 962 4588 971
rect 4612 961 4615 963
rect 4626 962 4635 971
rect 4920 970 4954 972
rect 4963 971 4964 972
rect 5010 971 5013 974
rect 4959 970 4964 971
rect 5009 970 5010 971
rect 4920 968 4964 970
rect 5007 969 5009 970
rect 4916 965 4917 967
rect 4690 961 4699 963
rect 4607 959 4612 961
rect 3985 945 3995 946
rect 4017 945 4018 946
rect 3981 943 3985 945
rect 4029 943 4049 946
rect 4130 943 4131 950
rect 4203 943 4204 950
rect 4252 943 4258 949
rect 4298 948 4304 949
rect 4335 948 4340 950
rect 4298 947 4335 948
rect 4298 943 4304 947
rect 4390 946 4396 952
rect 4436 946 4442 952
rect 4458 950 4459 959
rect 4605 958 4607 959
rect 4701 958 4707 961
rect 4476 955 4480 958
rect 4544 955 4546 958
rect 4480 946 4490 955
rect 3969 931 3977 943
rect 3981 941 4015 943
rect 3867 928 3928 931
rect 3867 917 3873 928
rect 3895 926 3928 928
rect 3889 925 3928 926
rect 3947 925 3953 926
rect 3889 921 3953 925
rect 3889 920 3975 921
rect 3867 915 3874 917
rect 3867 913 3876 915
rect 3895 914 3901 920
rect 3941 914 3947 920
rect 3950 917 3975 920
rect 3959 915 3975 917
rect 3964 913 3975 915
rect 3981 913 3983 941
rect 4012 939 4015 941
rect 3867 909 3882 913
rect 3969 909 3983 913
rect 4013 909 4015 939
rect 4019 931 4027 943
rect 4049 934 4112 943
rect 4246 938 4252 943
rect 4264 941 4300 943
rect 4264 939 4269 941
rect 4205 937 4252 938
rect 4266 937 4269 939
rect 4304 937 4310 943
rect 4384 940 4390 946
rect 4442 940 4448 946
rect 4457 938 4458 943
rect 4490 942 4495 946
rect 4546 942 4558 955
rect 4707 951 4720 958
rect 4930 956 4946 968
rect 4948 956 4964 968
rect 5003 965 5007 968
rect 5001 963 5003 965
rect 4999 961 5001 963
rect 5054 961 5067 974
rect 5103 967 5106 983
rect 5105 961 5106 967
rect 5109 967 5110 989
rect 5148 985 5155 989
rect 5176 987 5178 990
rect 5148 983 5149 985
rect 5169 984 5170 986
rect 5109 963 5111 967
rect 5142 963 5143 966
rect 5147 965 5149 983
rect 5178 981 5181 987
rect 5181 979 5182 981
rect 5183 975 5184 977
rect 5184 972 5185 975
rect 5224 973 5232 990
rect 5186 965 5189 969
rect 5109 961 5113 963
rect 5147 962 5148 965
rect 5189 963 5190 965
rect 4995 958 4998 961
rect 5067 959 5070 961
rect 4993 953 4995 958
rect 5070 957 5072 959
rect 4828 952 4865 953
rect 4992 952 4993 953
rect 5072 952 5074 957
rect 5100 955 5106 961
rect 5113 959 5119 961
rect 5120 957 5126 959
rect 5146 957 5152 961
rect 5190 960 5191 963
rect 5191 958 5192 960
rect 5126 956 5152 957
rect 4828 951 4853 952
rect 4865 951 4866 952
rect 4991 951 4992 952
rect 4722 948 4726 951
rect 4793 948 4820 951
rect 4868 948 4875 951
rect 4989 948 4991 951
rect 4875 943 4886 948
rect 4922 945 4923 947
rect 4987 943 4989 948
rect 5074 944 5077 951
rect 5094 949 5100 955
rect 5126 951 5170 956
rect 5192 955 5194 958
rect 5152 949 5158 951
rect 5194 948 5197 955
rect 4886 942 4890 943
rect 4558 939 4559 942
rect 4890 939 4895 942
rect 4895 938 4897 939
rect 4923 938 4926 943
rect 4957 941 4958 943
rect 4986 942 4987 943
rect 5197 942 5200 948
rect 5232 943 5233 973
rect 5340 951 5356 954
rect 5268 943 5291 951
rect 5356 943 5363 951
rect 4985 940 4986 942
rect 4984 939 4985 940
rect 5200 939 5201 942
rect 4205 936 4248 937
rect 4129 934 4130 936
rect 4151 934 4205 936
rect 4085 922 4100 934
rect 4112 933 4151 934
rect 4129 929 4130 933
rect 4261 929 4264 936
rect 4388 933 4390 934
rect 3782 904 3783 906
rect 3842 905 3843 909
rect 3848 903 3854 909
rect 3867 903 3886 909
rect 3894 903 3900 909
rect 3702 899 3704 903
rect 3742 899 3743 903
rect 3701 897 3702 899
rect 3741 897 3742 899
rect 3615 884 3623 896
rect 3627 894 3645 896
rect 3700 895 3701 896
rect 3780 895 3782 903
rect 3842 897 3848 903
rect 3867 897 3906 903
rect 3908 897 3920 905
rect 3981 904 3998 909
rect 4085 904 4100 920
rect 4127 906 4129 928
rect 3989 903 3990 904
rect 3998 903 4002 904
rect 4017 903 4019 904
rect 3979 901 3980 903
rect 3990 899 3996 903
rect 4002 900 4021 903
rect 4126 900 4138 905
rect 4148 900 4160 905
rect 4201 904 4203 928
rect 4252 904 4261 928
rect 4384 925 4388 933
rect 4297 904 4300 909
rect 4338 908 4373 910
rect 4333 907 4338 908
rect 4373 907 4381 908
rect 4384 907 4386 915
rect 4408 909 4409 929
rect 4456 928 4457 936
rect 4453 917 4455 920
rect 4450 915 4452 916
rect 4447 913 4450 915
rect 4444 911 4447 913
rect 4442 910 4444 911
rect 4328 906 4333 907
rect 4381 906 4390 907
rect 4317 904 4328 906
rect 4251 900 4252 903
rect 4295 900 4297 903
rect 4305 901 4317 904
rect 4384 900 4386 906
rect 4408 904 4409 906
rect 4476 904 4492 920
rect 4500 915 4526 938
rect 4560 931 4566 938
rect 4897 937 4899 938
rect 4899 933 4915 937
rect 4915 932 4920 933
rect 4926 932 4931 938
rect 4570 920 4578 927
rect 4578 918 4585 920
rect 4585 915 4597 918
rect 4526 910 4532 915
rect 4597 914 4601 915
rect 4604 914 4605 929
rect 4920 927 4936 932
rect 4958 929 4961 938
rect 4983 937 4984 938
rect 4980 933 4983 937
rect 4978 932 4980 933
rect 5201 932 5202 938
rect 5230 932 5232 942
rect 5262 939 5268 943
rect 5363 939 5367 943
rect 5260 938 5262 939
rect 5367 938 5370 939
rect 5250 932 5260 938
rect 5367 936 5372 938
rect 4961 927 4962 928
rect 4975 927 4978 932
rect 5099 927 5100 929
rect 4931 923 4932 926
rect 4936 924 4973 927
rect 4663 921 4694 922
rect 4654 920 4663 921
rect 4694 920 4701 921
rect 4961 920 4962 924
rect 4625 917 4654 920
rect 4701 917 4716 920
rect 4623 916 4625 917
rect 4620 915 4623 916
rect 4716 915 4724 917
rect 4933 915 4934 917
rect 4962 915 4963 920
rect 4967 915 4976 924
rect 5014 915 5023 924
rect 5098 922 5099 927
rect 5097 920 5098 922
rect 5096 918 5097 920
rect 5095 916 5096 918
rect 4613 914 4620 915
rect 4724 914 4733 915
rect 4958 914 4967 915
rect 4601 911 4967 914
rect 4604 910 4605 911
rect 4607 910 4609 911
rect 4743 910 4751 911
rect 4532 909 4534 910
rect 4409 903 4410 904
rect 4473 903 4476 904
rect 4534 903 4542 909
rect 4603 908 4607 910
rect 4751 907 4764 910
rect 4764 906 4769 907
rect 4596 904 4601 906
rect 4769 904 4779 906
rect 4410 900 4413 903
rect 4463 900 4476 903
rect 3867 895 3922 897
rect 3996 895 4002 899
rect 4016 898 4017 900
rect 3615 862 3623 874
rect 3627 864 3629 894
rect 3699 893 3700 894
rect 3740 893 3741 894
rect 3867 893 3924 895
rect 4002 893 4003 895
rect 4015 894 4016 897
rect 4021 896 4190 900
rect 4249 897 4251 900
rect 4246 896 4252 897
rect 4292 896 4295 900
rect 4122 894 4124 896
rect 4126 895 4127 896
rect 4190 895 4252 896
rect 3694 889 3700 893
rect 3739 889 3740 893
rect 3779 889 3780 893
rect 3835 889 3842 893
rect 3867 892 3932 893
rect 3680 888 3700 889
rect 3680 878 3694 888
rect 3736 879 3739 889
rect 3777 878 3779 889
rect 3832 879 3835 889
rect 3667 868 3680 878
rect 3733 869 3736 878
rect 3776 875 3777 878
rect 3831 875 3832 878
rect 3774 868 3776 875
rect 3829 869 3831 875
rect 3664 866 3667 868
rect 3627 862 3630 864
rect 3661 862 3664 866
rect 3711 859 3720 868
rect 3732 866 3733 868
rect 3731 862 3732 866
rect 3626 857 3628 858
rect 3633 857 3639 859
rect 3627 853 3639 857
rect 3691 853 3697 859
rect 3703 857 3711 859
rect 3730 858 3731 862
rect 3772 859 3774 867
rect 3826 859 3829 868
rect 3844 864 3847 892
rect 3894 891 3920 892
rect 3918 861 3920 891
rect 3924 881 3932 892
rect 4003 879 4023 893
rect 4071 879 4085 894
rect 4114 881 4122 893
rect 4126 891 4160 893
rect 3979 876 3980 879
rect 4009 876 4010 879
rect 4023 877 4035 879
rect 4069 877 4071 879
rect 4023 875 4069 877
rect 3894 859 3920 861
rect 3924 859 3932 871
rect 3977 869 3978 871
rect 4006 868 4007 870
rect 3974 860 3976 866
rect 4003 860 4006 867
rect 4126 859 4128 891
rect 4158 873 4160 891
rect 4164 881 4172 893
rect 4246 891 4252 895
rect 4290 891 4292 895
rect 4304 891 4310 897
rect 4384 894 4390 900
rect 4413 896 4428 900
rect 4428 895 4429 896
rect 4442 895 4476 900
rect 4542 899 4548 903
rect 4592 901 4596 904
rect 4200 881 4201 889
rect 4244 881 4247 891
rect 4252 885 4258 891
rect 4284 881 4290 891
rect 4298 885 4304 891
rect 4387 883 4388 891
rect 4390 888 4396 894
rect 4429 893 4448 895
rect 4159 865 4160 872
rect 4194 870 4200 880
rect 4239 870 4244 881
rect 4188 868 4194 870
rect 4238 868 4239 870
rect 4278 869 4284 881
rect 4427 872 4430 892
rect 4436 888 4442 893
rect 4460 888 4476 895
rect 4548 894 4559 899
rect 4587 898 4591 900
rect 4584 897 4587 898
rect 4580 894 4584 897
rect 4604 895 4607 900
rect 4779 897 4814 904
rect 4860 902 4873 903
rect 4839 900 4857 902
rect 4878 900 4901 902
rect 4837 899 4849 900
rect 4901 899 4910 900
rect 4910 898 4911 899
rect 4935 898 4936 904
rect 4830 897 4837 898
rect 4559 886 4590 894
rect 4607 893 4609 895
rect 4609 891 4611 893
rect 4814 891 4837 897
rect 4911 894 4918 898
rect 4918 891 4924 894
rect 4936 891 4937 897
rect 4549 880 4590 886
rect 4611 886 4684 891
rect 4814 889 4836 891
rect 4611 881 4761 886
rect 4822 882 4830 889
rect 4836 887 4841 889
rect 4841 886 4843 887
rect 4924 886 4937 891
rect 4965 887 4968 903
rect 5023 901 5032 915
rect 5093 911 5094 914
rect 5120 909 5152 914
rect 5087 903 5091 906
rect 5094 903 5100 909
rect 5120 904 5158 909
rect 5189 904 5250 932
rect 5369 931 5372 936
rect 5368 922 5372 931
rect 5117 903 5158 904
rect 5187 903 5189 904
rect 5197 903 5198 904
rect 5074 901 5086 902
rect 5032 899 5036 901
rect 5054 900 5074 901
rect 5048 899 5054 900
rect 5074 895 5076 900
rect 5100 897 5106 903
rect 5134 899 5135 901
rect 5072 892 5074 895
rect 5071 891 5072 892
rect 4549 876 4566 880
rect 4590 876 4608 880
rect 4611 876 4631 881
rect 4683 876 4774 881
rect 4608 875 4774 876
rect 4815 875 4822 882
rect 4843 876 4867 886
rect 4924 882 4938 886
rect 4937 881 4940 882
rect 4937 878 4938 881
rect 4940 880 4941 881
rect 4867 875 4870 876
rect 4546 874 4548 875
rect 4607 874 4777 875
rect 4544 873 4546 874
rect 4605 873 4607 874
rect 4603 872 4605 873
rect 4608 872 4774 874
rect 4777 873 4785 874
rect 4785 872 4793 873
rect 4812 872 4815 875
rect 4870 874 4872 875
rect 4872 873 4875 874
rect 4875 872 4877 873
rect 4886 872 4898 878
rect 4941 875 4950 880
rect 4968 876 4970 886
rect 5059 882 5071 891
rect 5053 881 5059 882
rect 5025 880 5041 881
rect 5049 880 5053 881
rect 5118 880 5133 899
rect 5146 897 5152 903
rect 5183 901 5187 903
rect 5172 895 5183 901
rect 5196 899 5197 901
rect 5169 892 5172 895
rect 5168 891 5169 892
rect 5160 886 5168 891
rect 4997 875 5020 880
rect 5148 876 5180 886
rect 5193 880 5196 898
rect 5192 876 5193 880
rect 5228 878 5230 904
rect 5368 903 5369 922
rect 5383 915 5392 924
rect 5430 915 5439 924
rect 5374 906 5379 915
rect 5444 906 5448 915
rect 5349 881 5368 901
rect 4182 866 4188 868
rect 4277 867 4278 868
rect 4276 866 4277 867
rect 4181 865 4182 866
rect 4159 860 4181 865
rect 4235 862 4238 866
rect 4160 859 4181 860
rect 4232 859 4238 862
rect 3702 855 3711 857
rect 3627 850 3636 853
rect 3639 850 3645 853
rect 3690 852 3691 853
rect 3700 852 3711 855
rect 3647 851 3695 852
rect 3698 851 3700 852
rect 3647 850 3698 851
rect 3702 850 3711 852
rect 3637 847 3645 850
rect 3637 842 3641 847
rect 3690 840 3691 850
rect 3726 845 3730 858
rect 3769 846 3772 858
rect 3822 846 3826 858
rect 3842 851 3848 857
rect 3871 856 3875 859
rect 4165 858 4166 859
rect 3848 845 3854 851
rect 3866 845 3871 856
rect 3900 851 3906 857
rect 3973 855 3974 858
rect 4002 855 4003 858
rect 4232 857 4235 859
rect 4234 856 4235 857
rect 4230 855 4234 856
rect 3894 845 3900 851
rect 3908 847 3920 855
rect 4124 853 4125 855
rect 3971 851 3972 853
rect 3722 841 3726 845
rect 3768 841 3769 845
rect 3820 842 3822 845
rect 3720 840 3722 841
rect 3864 840 3866 845
rect 3968 841 3971 850
rect 3998 841 4001 850
rect 4125 841 4127 849
rect 4166 842 4167 849
rect 4227 847 4234 855
rect 4224 842 4227 847
rect 4230 845 4234 847
rect 4264 845 4276 865
rect 4388 859 4390 872
rect 4541 871 4543 872
rect 4601 871 4603 872
rect 4224 841 4226 842
rect 4221 840 4224 841
rect 4228 840 4230 845
rect 4261 844 4268 845
rect 4423 844 4427 870
rect 4536 868 4541 871
rect 4596 869 4600 871
rect 4684 869 4908 872
rect 4950 871 4956 875
rect 4987 871 4997 875
rect 5111 872 5114 876
rect 5145 875 5180 876
rect 4956 869 4962 871
rect 4969 869 4997 871
rect 4593 867 4595 868
rect 4533 866 4535 867
rect 4591 866 4593 867
rect 4700 866 4908 869
rect 4962 868 4963 869
rect 4969 868 4987 869
rect 4963 867 4967 868
rect 4982 867 4985 868
rect 4523 860 4533 866
rect 4581 862 4591 866
rect 4700 863 4910 866
rect 4813 862 4822 863
rect 4896 862 4918 863
rect 4939 862 4940 867
rect 5103 863 5111 872
rect 5158 869 5159 874
rect 5278 873 5289 874
rect 5306 873 5317 874
rect 5278 872 5286 873
rect 5310 872 5317 873
rect 4822 860 4825 862
rect 4518 857 4523 860
rect 4509 852 4518 857
rect 4825 852 4840 860
rect 4896 854 4910 862
rect 4918 856 4951 862
rect 5099 857 5103 862
rect 5026 856 5038 857
rect 4951 855 4957 856
rect 4975 855 4997 856
rect 4957 854 4997 855
rect 5018 854 5038 856
rect 4507 851 4509 852
rect 4840 851 4842 852
rect 4504 850 4507 851
rect 4842 850 4844 851
rect 4469 849 4475 850
rect 4502 849 4504 850
rect 4451 844 4502 849
rect 4515 844 4521 850
rect 4565 845 4568 849
rect 4845 845 4853 849
rect 4896 846 4908 854
rect 5026 851 5058 854
rect 5027 847 5058 851
rect 5096 849 5098 856
rect 5096 847 5097 849
rect 4261 840 4265 844
rect 3642 836 3643 840
rect 3643 833 3644 836
rect 3690 832 3692 840
rect 3708 832 3720 840
rect 3767 838 3768 840
rect 3819 838 3820 840
rect 3766 832 3767 838
rect 3818 833 3819 838
rect 3861 832 3864 840
rect 3967 837 3968 840
rect 3966 833 3967 836
rect 3995 834 3997 840
rect 4167 837 4168 840
rect 4128 832 4132 837
rect 4219 832 4228 840
rect 4257 834 4265 840
rect 4257 832 4261 834
rect 3644 817 3652 832
rect 3690 825 3694 832
rect 3707 830 3708 832
rect 3860 830 3861 832
rect 3706 828 3707 830
rect 3765 828 3766 830
rect 3816 828 3817 830
rect 3705 825 3706 828
rect 3692 817 3694 825
rect 3764 824 3765 828
rect 3815 824 3816 827
rect 3858 824 3860 829
rect 3703 819 3705 824
rect 3763 819 3764 824
rect 3810 820 3815 824
rect 3652 809 3656 817
rect 3694 811 3695 817
rect 3702 815 3703 819
rect 3762 815 3763 819
rect 3810 815 3814 820
rect 3856 819 3858 824
rect 3701 809 3702 814
rect 3760 809 3762 814
rect 3810 809 3812 815
rect 3853 814 3856 818
rect 3906 814 3922 824
rect 3924 814 3940 824
rect 3960 817 3966 832
rect 3849 809 3853 814
rect 3893 809 3900 814
rect 3945 808 3953 814
rect 3958 811 3960 817
rect 3988 811 3995 832
rect 4129 827 4133 832
rect 4168 827 4174 832
rect 4217 830 4219 832
rect 4256 830 4257 832
rect 3987 809 3988 811
rect 4002 808 4018 824
rect 4118 822 4184 827
rect 4210 824 4217 830
rect 4253 825 4256 830
rect 4259 828 4261 832
rect 4390 832 4392 844
rect 4402 840 4414 844
rect 4430 842 4451 844
rect 4421 841 4430 842
rect 4416 840 4423 841
rect 4402 836 4416 840
rect 4118 821 4174 822
rect 4109 814 4118 821
rect 4129 818 4133 821
rect 4107 811 4109 814
rect 4132 811 4133 817
rect 4168 811 4174 821
rect 4184 814 4188 821
rect 4202 819 4210 824
rect 4250 819 4253 824
rect 4202 818 4204 819
rect 4202 815 4203 818
rect 4248 817 4250 819
rect 4247 816 4248 817
rect 4188 811 4189 814
rect 4201 812 4202 813
rect 4247 812 4250 816
rect 4280 812 4292 815
rect 4190 811 4199 812
rect 4025 808 4044 809
rect 4050 808 4052 809
rect 3657 804 3658 807
rect 3658 799 3660 803
rect 3695 799 3696 803
rect 3698 800 3701 808
rect 3758 800 3760 808
rect 3660 794 3662 798
rect 3698 794 3700 800
rect 3756 794 3758 798
rect 3663 785 3666 793
rect 3697 790 3699 793
rect 3700 790 3714 794
rect 3697 786 3714 790
rect 3666 775 3671 785
rect 3671 771 3672 775
rect 3698 774 3714 786
rect 3748 790 3756 794
rect 3794 792 3810 808
rect 3844 801 3849 808
rect 3889 801 3893 808
rect 3945 807 3956 808
rect 3986 807 4002 808
rect 4052 807 4053 808
rect 4101 807 4107 810
rect 4174 809 4175 811
rect 4129 808 4131 809
rect 4189 808 4199 811
rect 4246 808 4247 812
rect 4280 808 4296 812
rect 4298 808 4314 824
rect 4316 808 4332 824
rect 4390 820 4398 832
rect 4402 831 4418 832
rect 4402 830 4412 831
rect 4334 808 4343 812
rect 4393 810 4394 811
rect 4118 807 4128 808
rect 3945 806 3957 807
rect 3952 804 3957 806
rect 3844 792 3847 801
rect 3748 774 3764 790
rect 3794 774 3810 790
rect 3844 787 3860 790
rect 3839 781 3860 787
rect 3880 787 3889 801
rect 3952 792 3956 804
rect 3985 803 4002 807
rect 4053 806 4056 807
rect 3984 799 3985 803
rect 3982 794 3984 798
rect 3986 792 4002 803
rect 4025 798 4037 806
rect 4056 803 4059 806
rect 4079 803 4118 807
rect 4175 803 4176 807
rect 4186 803 4201 808
rect 4280 807 4297 808
rect 4302 807 4314 808
rect 4040 799 4079 803
rect 4090 799 4096 803
rect 4101 799 4107 803
rect 4176 799 4177 803
rect 3880 785 3891 787
rect 3900 785 3912 791
rect 3952 785 3953 792
rect 3980 788 3982 792
rect 3869 783 3891 785
rect 3901 783 3912 785
rect 3951 783 3956 785
rect 3863 781 3868 783
rect 3833 775 3839 781
rect 3844 774 3860 781
rect 3878 779 3880 783
rect 3885 781 3891 783
rect 3912 781 3916 783
rect 3891 775 3897 781
rect 3900 778 3912 779
rect 3700 771 3704 774
rect 3672 754 3680 771
rect 3704 754 3711 771
rect 3714 758 3730 774
rect 3732 758 3748 774
rect 3810 772 3818 774
rect 3836 772 3844 774
rect 3910 772 3912 778
rect 3916 772 3924 779
rect 3949 778 3951 783
rect 3952 778 3956 783
rect 3949 774 3956 778
rect 3949 772 3951 774
rect 3810 758 3826 772
rect 3828 758 3844 772
rect 3891 757 3954 772
rect 3978 760 3980 786
rect 3986 774 4002 790
rect 4013 782 4021 794
rect 4025 793 4046 794
rect 4084 793 4090 799
rect 4025 792 4043 793
rect 4002 763 4006 767
rect 4013 763 4021 772
rect 4025 763 4027 792
rect 4178 788 4180 796
rect 4186 794 4208 803
rect 4186 792 4201 794
rect 4238 790 4246 806
rect 4276 804 4278 807
rect 4282 806 4296 807
rect 4280 803 4296 806
rect 4332 805 4348 808
rect 4330 803 4348 805
rect 4268 791 4276 803
rect 4278 801 4314 803
rect 4278 793 4298 801
rect 4311 800 4314 801
rect 4312 793 4314 800
rect 4318 799 4326 803
rect 4330 799 4352 803
rect 4332 794 4352 799
rect 4390 798 4398 810
rect 4402 800 4404 830
rect 4421 826 4423 840
rect 4463 838 4469 844
rect 4521 838 4527 844
rect 4560 841 4565 845
rect 4853 841 4858 845
rect 4852 832 4860 841
rect 4864 834 4866 839
rect 4896 834 4898 846
rect 5156 845 5158 865
rect 5190 863 5192 872
rect 5227 863 5228 872
rect 5278 871 5280 872
rect 5316 871 5317 872
rect 5349 868 5363 881
rect 5342 866 5355 868
rect 5342 865 5354 866
rect 5383 865 5388 866
rect 5189 857 5190 862
rect 5187 849 5188 855
rect 4908 844 4911 845
rect 4864 832 4898 834
rect 4902 840 4911 844
rect 4902 832 4910 840
rect 4911 832 4915 840
rect 4915 830 4916 832
rect 4436 826 4437 830
rect 4547 829 4550 830
rect 4523 827 4558 829
rect 4421 818 4422 826
rect 4519 825 4523 827
rect 4517 824 4519 825
rect 4437 812 4439 824
rect 4422 800 4425 811
rect 4490 808 4517 824
rect 4521 812 4525 817
rect 4531 812 4547 827
rect 4558 824 4583 827
rect 4526 811 4547 812
rect 4402 798 4436 800
rect 4422 795 4425 798
rect 4180 778 4183 788
rect 4183 769 4185 778
rect 4186 774 4201 790
rect 4238 774 4252 790
rect 4275 781 4276 788
rect 4185 765 4186 769
rect 4002 762 4027 763
rect 4056 762 4059 763
rect 4002 760 4059 762
rect 4002 758 4018 760
rect 4186 759 4187 763
rect 3680 746 3683 754
rect 3711 748 3716 754
rect 3716 745 3720 748
rect 3910 745 3912 757
rect 3915 745 3949 757
rect 3954 756 3956 757
rect 4063 756 4090 759
rect 4187 757 4188 759
rect 4202 758 4218 772
rect 4220 758 4236 772
rect 4268 769 4276 781
rect 4280 774 4298 793
rect 4332 792 4348 794
rect 4332 774 4348 790
rect 4378 774 4393 790
rect 4395 775 4397 792
rect 4402 786 4414 794
rect 4424 786 4436 794
rect 4438 790 4439 808
rect 4525 805 4535 811
rect 4583 808 4724 824
rect 4786 808 4802 824
rect 4804 808 4820 824
rect 4864 820 4876 828
rect 4886 820 4898 828
rect 4916 826 4917 830
rect 4942 828 4944 845
rect 4864 810 4866 820
rect 4917 816 4920 824
rect 4944 819 4945 828
rect 4972 819 4975 845
rect 5014 833 5020 845
rect 5061 843 5063 844
rect 5186 843 5187 847
rect 5097 838 5098 843
rect 5064 827 5065 836
rect 5098 827 5099 836
rect 5154 825 5156 840
rect 5185 837 5186 843
rect 5183 827 5185 836
rect 5225 829 5227 862
rect 5338 855 5354 865
rect 5391 864 5395 868
rect 5275 845 5338 855
rect 5383 851 5391 864
rect 5266 844 5275 845
rect 5260 842 5266 844
rect 5258 840 5260 842
rect 5014 811 5020 823
rect 5182 821 5183 826
rect 5223 820 5225 827
rect 5239 825 5258 840
rect 5238 824 5239 825
rect 5066 817 5067 820
rect 5099 816 5100 820
rect 5067 811 5072 816
rect 5100 811 5101 816
rect 5153 811 5154 818
rect 5167 811 5173 817
rect 5181 816 5182 820
rect 5222 818 5223 820
rect 5230 818 5238 824
rect 5179 812 5181 816
rect 5213 811 5219 817
rect 5221 816 5230 818
rect 5220 811 5230 816
rect 4976 808 4977 810
rect 5068 808 5069 810
rect 4530 803 4535 805
rect 4655 803 4664 808
rect 4702 803 4711 808
rect 4442 802 4451 803
rect 4440 798 4448 802
rect 4451 799 4466 802
rect 4466 798 4469 799
rect 4463 792 4469 798
rect 4521 792 4527 798
rect 4535 794 4544 803
rect 4646 794 4655 803
rect 4711 794 4720 803
rect 4637 792 4644 793
rect 4469 790 4475 792
rect 4280 772 4314 774
rect 4327 772 4332 774
rect 4425 772 4428 786
rect 4438 774 4444 790
rect 4469 786 4490 790
rect 4515 786 4521 792
rect 4631 791 4637 792
rect 4688 791 4692 793
rect 4724 792 4740 808
rect 4770 792 4786 808
rect 4797 803 4803 808
rect 4797 802 4812 803
rect 4791 796 4797 802
rect 4820 798 4836 808
rect 4843 802 4849 808
rect 4796 791 4797 793
rect 4829 791 4834 798
rect 4849 796 4855 802
rect 4867 800 4868 808
rect 4629 790 4631 791
rect 4628 787 4629 790
rect 4693 789 4695 790
rect 4474 774 4490 786
rect 4541 778 4568 781
rect 4524 774 4541 778
rect 4568 774 4576 778
rect 4280 769 4332 772
rect 4393 769 4399 772
rect 4428 771 4432 772
rect 4280 757 4284 765
rect 4316 758 4332 769
rect 4394 762 4411 769
rect 4428 762 4438 771
rect 4394 758 4410 762
rect 4411 760 4416 762
rect 4420 760 4432 762
rect 4416 759 4432 760
rect 4412 758 4432 759
rect 4490 758 4506 774
rect 4576 772 4579 774
rect 4644 772 4650 778
rect 4653 772 4655 779
rect 4695 772 4696 778
rect 4724 774 4740 790
rect 4770 774 4786 790
rect 4788 779 4797 791
rect 4579 763 4599 772
rect 4628 767 4629 769
rect 4638 766 4644 772
rect 4696 766 4702 772
rect 4717 763 4724 774
rect 4599 762 4601 763
rect 4601 759 4607 762
rect 3956 751 3977 756
rect 3977 747 3993 751
rect 4025 748 4037 756
rect 4188 754 4189 756
rect 4084 747 4090 753
rect 4115 747 4170 753
rect 4189 750 4190 754
rect 4190 747 4192 748
rect 4199 747 4208 756
rect 4278 747 4284 756
rect 4336 747 4342 753
rect 4343 747 4352 756
rect 4397 751 4400 758
rect 3683 741 3685 745
rect 3720 740 3728 745
rect 3946 742 3947 745
rect 3993 742 4013 747
rect 4013 741 4018 742
rect 4090 741 4096 747
rect 4136 741 4142 747
rect 3912 740 3914 741
rect 3685 737 3687 740
rect 3728 737 3733 740
rect 3902 739 3912 740
rect 3891 738 3912 739
rect 4018 738 4022 741
rect 4143 738 4152 747
rect 4190 745 4199 747
rect 4190 742 4205 745
rect 4190 738 4199 742
rect 4205 740 4209 742
rect 4284 741 4296 747
rect 4330 741 4343 747
rect 4399 744 4400 751
rect 4209 739 4212 740
rect 3733 736 3735 737
rect 3900 736 3919 738
rect 3688 733 3689 736
rect 3735 733 3739 736
rect 3689 727 3692 733
rect 3739 731 3743 733
rect 3743 729 3746 731
rect 3833 729 3839 735
rect 3891 729 3897 735
rect 3900 733 3937 736
rect 3944 733 3945 736
rect 3911 729 3937 733
rect 3940 729 3944 731
rect 3976 729 3977 730
rect 3746 726 3750 729
rect 3692 720 3696 726
rect 3750 720 3760 726
rect 3763 720 3775 724
rect 3839 723 3845 729
rect 3885 723 3891 729
rect 3937 726 3977 729
rect 3937 723 3976 726
rect 4022 725 4039 738
rect 4143 737 4144 738
rect 4212 736 4219 739
rect 4287 738 4296 741
rect 4334 738 4343 741
rect 4393 739 4400 744
rect 4428 742 4432 758
rect 4470 747 4479 756
rect 4535 747 4544 756
rect 4607 754 4618 759
rect 4711 758 4724 763
rect 4786 769 4795 774
rect 4796 769 4797 779
rect 4786 763 4797 769
rect 4800 763 4802 791
rect 4868 790 4870 791
rect 4866 785 4870 790
rect 4919 790 4920 808
rect 5026 799 5038 803
rect 5048 799 5060 803
rect 5070 796 5071 799
rect 5101 796 5102 805
rect 5152 799 5153 808
rect 5161 805 5167 811
rect 5219 808 5225 811
rect 5274 808 5290 824
rect 5863 819 5864 1015
rect 6053 819 6054 1015
rect 6139 819 6140 1015
rect 6412 819 6413 1015
rect 6610 820 6611 1016
rect 7001 1014 7005 1019
rect 7639 1014 7646 1019
rect 7726 1018 7735 1027
rect 7791 1024 7887 1027
rect 8228 1023 8336 1037
rect 8086 1015 8102 1022
rect 8104 1015 8120 1022
rect 7646 1007 7658 1014
rect 8076 1013 8088 1015
rect 8098 1013 8110 1015
rect 8116 1013 8120 1015
rect 8304 1013 8320 1022
rect 8336 1021 8354 1023
rect 8355 1017 8362 1020
rect 8362 1013 8368 1017
rect 9008 1015 9009 1026
rect 9198 1015 9199 1026
rect 9284 1015 9285 1026
rect 9557 1015 9558 1026
rect 9755 1016 9756 1027
rect 10181 1023 10282 1034
rect 10468 1033 10732 1034
rect 10732 1023 10787 1033
rect 10890 1027 10899 1036
rect 10937 1027 10946 1036
rect 11240 1034 11362 1037
rect 11212 1033 11229 1034
rect 11042 1027 11212 1033
rect 10166 1021 10181 1023
rect 10160 1019 10166 1021
rect 10789 1019 10794 1021
rect 8076 1008 8120 1013
rect 8263 1008 8300 1009
rect 8368 1008 8371 1013
rect 8072 1006 8074 1008
rect 8076 1006 8208 1008
rect 7127 1005 7481 1006
rect 7107 1003 7125 1005
rect 7567 1003 7580 1005
rect 7659 1003 7662 1005
rect 8070 1003 8208 1006
rect 7051 1000 7107 1003
rect 6925 992 6937 1000
rect 6947 992 6959 1000
rect 7023 994 7107 1000
rect 7580 994 7590 1003
rect 7023 993 7051 994
rect 6921 989 6923 992
rect 7023 991 7042 993
rect 7591 991 7594 993
rect 6963 988 6967 989
rect 6913 977 6921 988
rect 6924 986 6959 988
rect 6922 977 6924 983
rect 6913 976 6922 977
rect 6921 972 6922 976
rect 6920 971 6921 972
rect 6918 966 6920 969
rect 6793 964 6858 965
rect 6785 956 6793 964
rect 6858 956 6862 964
rect 6784 950 6785 956
rect 6913 954 6921 966
rect 6925 956 6927 986
rect 6956 985 6959 986
rect 6958 979 6959 985
rect 6963 981 6971 988
rect 6967 980 6975 981
rect 6999 980 7000 990
rect 7023 980 7038 991
rect 7297 981 7334 983
rect 6975 979 6981 980
rect 6998 979 6999 980
rect 7023 979 7030 980
rect 6981 969 7043 979
rect 7051 972 7057 978
rect 7097 972 7103 978
rect 7297 977 7323 981
rect 7334 977 7339 981
rect 7594 980 7607 991
rect 7570 979 7584 980
rect 7291 972 7297 977
rect 7339 972 7348 977
rect 7552 972 7570 979
rect 7584 977 7591 979
rect 7662 977 7683 1003
rect 8064 996 8208 1003
rect 8224 1006 8325 1008
rect 8224 996 8336 1006
rect 8025 990 8086 996
rect 7990 987 8025 990
rect 7803 981 7990 987
rect 8076 986 8086 990
rect 7591 972 7606 977
rect 7045 969 7051 972
rect 7052 970 7109 972
rect 7348 971 7349 972
rect 7186 970 7189 971
rect 7207 970 7210 971
rect 7289 970 7290 971
rect 7349 970 7352 971
rect 7052 969 7060 970
rect 7023 968 7060 969
rect 6925 954 6959 956
rect 6914 951 6916 954
rect 6910 939 6914 950
rect 6925 942 6937 950
rect 6950 945 6959 954
rect 6997 952 6998 955
rect 7023 951 7028 968
rect 7045 966 7060 968
rect 7103 966 7109 970
rect 7182 967 7186 970
rect 7210 967 7215 970
rect 7352 968 7353 970
rect 7544 969 7552 972
rect 7581 971 7606 972
rect 7615 971 7619 972
rect 7577 970 7581 971
rect 7591 970 7628 971
rect 7353 967 7356 968
rect 7051 964 7060 966
rect 7051 951 7056 964
rect 7104 955 7123 958
rect 7158 955 7182 967
rect 7215 959 7233 967
rect 7288 959 7289 967
rect 6960 948 6970 950
rect 6970 947 6973 948
rect 6975 945 6984 947
rect 6948 942 6950 945
rect 6984 943 6995 945
rect 6996 943 6997 951
rect 7023 943 7029 951
rect 6947 939 6948 942
rect 6995 938 7029 943
rect 6861 924 6862 938
rect 6811 915 6820 924
rect 6858 920 6867 924
rect 6858 915 6872 920
rect 6802 912 6811 915
rect 6802 911 6805 912
rect 6795 908 6804 911
rect 6783 907 6804 908
rect 6783 905 6801 907
rect 6841 905 6847 911
rect 6861 906 6876 915
rect 6901 908 6910 937
rect 6783 900 6795 905
rect 6779 898 6782 900
rect 6783 899 6784 900
rect 6789 899 6795 900
rect 6847 899 6853 905
rect 6860 904 6872 906
rect 6899 904 6901 908
rect 6939 907 6947 938
rect 6996 926 6997 938
rect 7023 935 7051 938
rect 7023 931 7053 935
rect 7055 931 7056 951
rect 7123 946 7185 955
rect 7233 952 7241 959
rect 7287 951 7288 958
rect 7356 954 7360 967
rect 7536 966 7544 969
rect 7574 968 7577 970
rect 7570 967 7574 968
rect 7565 965 7570 967
rect 7591 965 7606 970
rect 7615 969 7619 970
rect 7628 969 7629 970
rect 7685 969 7690 975
rect 7726 971 7735 980
rect 7791 978 7803 981
rect 7791 971 7800 978
rect 8070 972 8086 986
rect 8109 972 8110 996
rect 8115 991 8136 996
rect 8120 990 8136 991
rect 8253 989 8259 996
rect 8305 989 8311 996
rect 8325 990 8336 996
rect 8371 990 8380 1008
rect 8120 972 8136 988
rect 8253 985 8261 989
rect 8259 983 8261 985
rect 8169 974 8197 978
rect 8199 974 8210 978
rect 7619 965 7624 969
rect 7629 965 7631 968
rect 7690 965 7693 969
rect 7531 964 7535 965
rect 7606 964 7609 965
rect 7631 964 7632 965
rect 7527 962 7531 964
rect 7496 950 7527 962
rect 7611 959 7615 962
rect 7626 960 7630 963
rect 7735 962 7744 971
rect 7768 961 7771 963
rect 7782 962 7791 971
rect 8076 970 8110 972
rect 8119 971 8120 972
rect 8166 971 8169 974
rect 8115 970 8120 971
rect 8165 970 8166 971
rect 8076 968 8120 970
rect 8163 969 8165 970
rect 8072 965 8073 967
rect 7846 961 7855 963
rect 7763 959 7768 961
rect 7141 945 7151 946
rect 7173 945 7174 946
rect 7137 943 7141 945
rect 7185 943 7205 946
rect 7286 943 7287 950
rect 7359 943 7360 950
rect 7408 943 7414 949
rect 7454 948 7460 949
rect 7491 948 7496 950
rect 7454 947 7491 948
rect 7454 943 7460 947
rect 7546 946 7552 952
rect 7592 946 7598 952
rect 7614 950 7615 959
rect 7761 958 7763 959
rect 7857 958 7863 961
rect 7632 955 7636 958
rect 7700 955 7702 958
rect 7636 946 7646 955
rect 7125 931 7133 943
rect 7137 941 7171 943
rect 7023 928 7084 931
rect 7023 917 7029 928
rect 7051 926 7084 928
rect 7045 925 7084 926
rect 7103 925 7109 926
rect 7045 921 7109 925
rect 7045 920 7131 921
rect 7023 915 7030 917
rect 7023 913 7032 915
rect 7051 914 7057 920
rect 7097 914 7103 920
rect 7106 917 7131 920
rect 7115 915 7131 917
rect 7120 913 7131 915
rect 7137 913 7139 941
rect 7168 939 7171 941
rect 7023 909 7038 913
rect 7125 909 7139 913
rect 7169 909 7171 939
rect 7175 931 7183 943
rect 7205 934 7268 943
rect 7402 938 7408 943
rect 7420 941 7456 943
rect 7420 939 7425 941
rect 7361 937 7408 938
rect 7422 937 7425 939
rect 7460 937 7466 943
rect 7540 940 7546 946
rect 7598 940 7604 946
rect 7613 938 7614 943
rect 7646 942 7651 946
rect 7702 942 7714 955
rect 7863 951 7876 958
rect 8086 956 8102 968
rect 8104 956 8120 968
rect 8159 965 8163 968
rect 8157 963 8159 965
rect 8155 961 8157 963
rect 8210 961 8223 974
rect 8259 967 8262 983
rect 8261 961 8262 967
rect 8265 967 8266 989
rect 8304 985 8311 989
rect 8332 987 8334 990
rect 8304 983 8305 985
rect 8325 984 8326 986
rect 8265 963 8267 967
rect 8298 963 8299 966
rect 8303 965 8305 983
rect 8334 981 8337 987
rect 8337 979 8338 981
rect 8339 975 8340 977
rect 8340 972 8341 975
rect 8380 973 8388 990
rect 8342 965 8345 969
rect 8265 961 8269 963
rect 8303 962 8304 965
rect 8345 963 8346 965
rect 8151 958 8154 961
rect 8223 959 8226 961
rect 8149 953 8151 958
rect 8226 957 8228 959
rect 7984 952 8021 953
rect 8148 952 8149 953
rect 8228 952 8230 957
rect 8256 955 8262 961
rect 8269 959 8275 961
rect 8276 957 8282 959
rect 8302 957 8308 961
rect 8346 960 8347 963
rect 8347 958 8348 960
rect 8282 956 8308 957
rect 7984 951 8009 952
rect 8021 951 8022 952
rect 8147 951 8148 952
rect 7878 948 7882 951
rect 7949 948 7976 951
rect 8024 948 8031 951
rect 8145 948 8147 951
rect 8031 943 8042 948
rect 8078 945 8079 947
rect 8143 943 8145 948
rect 8230 944 8233 951
rect 8250 949 8256 955
rect 8282 951 8326 956
rect 8348 955 8350 958
rect 8308 949 8314 951
rect 8350 948 8353 955
rect 8042 942 8046 943
rect 7714 939 7715 942
rect 8046 939 8051 942
rect 8051 938 8053 939
rect 8079 938 8082 943
rect 8113 941 8114 943
rect 8142 942 8143 943
rect 8353 942 8356 948
rect 8388 943 8389 973
rect 8496 951 8512 954
rect 8424 943 8447 951
rect 8512 943 8519 951
rect 8141 940 8142 942
rect 8140 939 8141 940
rect 8356 939 8357 942
rect 7361 936 7404 937
rect 7285 934 7286 936
rect 7307 934 7361 936
rect 7241 922 7256 934
rect 7268 933 7307 934
rect 7285 929 7286 933
rect 7417 929 7420 936
rect 7544 933 7546 934
rect 6938 904 6939 906
rect 6998 905 6999 909
rect 7004 903 7010 909
rect 7023 903 7042 909
rect 7050 903 7056 909
rect 6858 899 6860 903
rect 6898 899 6899 903
rect 6857 897 6858 899
rect 6897 897 6898 899
rect 6771 884 6779 896
rect 6783 894 6801 896
rect 6856 895 6857 896
rect 6936 895 6938 903
rect 6998 897 7004 903
rect 7023 897 7062 903
rect 7064 897 7076 905
rect 7137 904 7154 909
rect 7241 904 7256 920
rect 7283 906 7285 928
rect 7145 903 7146 904
rect 7154 903 7158 904
rect 7173 903 7175 904
rect 7135 901 7136 903
rect 7146 899 7152 903
rect 7158 900 7177 903
rect 7282 900 7294 905
rect 7304 900 7316 905
rect 7357 904 7359 928
rect 7408 904 7417 928
rect 7540 925 7544 933
rect 7453 904 7456 909
rect 7494 908 7529 910
rect 7489 907 7494 908
rect 7529 907 7537 908
rect 7540 907 7542 915
rect 7564 909 7565 929
rect 7612 928 7613 936
rect 7609 917 7611 920
rect 7606 915 7608 916
rect 7603 913 7606 915
rect 7600 911 7603 913
rect 7598 910 7600 911
rect 7484 906 7489 907
rect 7537 906 7546 907
rect 7473 904 7484 906
rect 7407 900 7408 903
rect 7451 900 7453 903
rect 7461 901 7473 904
rect 7540 900 7542 906
rect 7564 904 7565 906
rect 7632 904 7648 920
rect 7656 915 7682 938
rect 7716 931 7722 938
rect 8053 937 8055 938
rect 8055 933 8071 937
rect 8071 932 8076 933
rect 8082 932 8087 938
rect 7726 920 7734 927
rect 7734 918 7741 920
rect 7741 915 7753 918
rect 7682 910 7688 915
rect 7753 914 7757 915
rect 7760 914 7761 929
rect 8076 927 8092 932
rect 8114 929 8117 938
rect 8139 937 8140 938
rect 8136 933 8139 937
rect 8134 932 8136 933
rect 8357 932 8358 938
rect 8386 932 8388 942
rect 8418 939 8424 943
rect 8519 939 8523 943
rect 8416 938 8418 939
rect 8523 938 8526 939
rect 8406 932 8416 938
rect 8523 936 8528 938
rect 8117 927 8118 928
rect 8131 927 8134 932
rect 8255 927 8256 929
rect 8087 923 8088 926
rect 8092 924 8129 927
rect 7819 921 7850 922
rect 7810 920 7819 921
rect 7850 920 7857 921
rect 8117 920 8118 924
rect 7781 917 7810 920
rect 7857 917 7872 920
rect 7779 916 7781 917
rect 7776 915 7779 916
rect 7872 915 7880 917
rect 8089 915 8090 917
rect 8118 915 8119 920
rect 8123 915 8132 924
rect 8170 915 8179 924
rect 8254 922 8255 927
rect 8253 920 8254 922
rect 8252 918 8253 920
rect 8251 916 8252 918
rect 7769 914 7776 915
rect 7880 914 7889 915
rect 8114 914 8123 915
rect 7757 911 8123 914
rect 7760 910 7761 911
rect 7763 910 7765 911
rect 7899 910 7907 911
rect 7688 909 7690 910
rect 7565 903 7566 904
rect 7629 903 7632 904
rect 7690 903 7698 909
rect 7759 908 7763 910
rect 7907 907 7920 910
rect 7920 906 7925 907
rect 7752 904 7757 906
rect 7925 904 7935 906
rect 7566 900 7569 903
rect 7619 900 7632 903
rect 7023 895 7078 897
rect 7152 895 7158 899
rect 7172 898 7173 900
rect 6771 862 6779 874
rect 6783 864 6785 894
rect 6855 893 6856 894
rect 6896 893 6897 894
rect 7023 893 7080 895
rect 7158 893 7159 895
rect 7171 894 7172 897
rect 7177 896 7346 900
rect 7405 897 7407 900
rect 7402 896 7408 897
rect 7448 896 7451 900
rect 7278 894 7280 896
rect 7282 895 7283 896
rect 7346 895 7408 896
rect 6850 889 6856 893
rect 6895 889 6896 893
rect 6935 889 6936 893
rect 6991 889 6998 893
rect 7023 892 7088 893
rect 6836 888 6856 889
rect 6836 878 6850 888
rect 6892 879 6895 889
rect 6933 878 6935 889
rect 6988 879 6991 889
rect 6823 868 6836 878
rect 6889 869 6892 878
rect 6932 875 6933 878
rect 6987 875 6988 878
rect 6930 868 6932 875
rect 6985 869 6987 875
rect 6820 866 6823 868
rect 6783 862 6786 864
rect 6817 862 6820 866
rect 6867 859 6876 868
rect 6888 866 6889 868
rect 6887 862 6888 866
rect 6782 857 6784 858
rect 6789 857 6795 859
rect 6783 853 6795 857
rect 6847 853 6853 859
rect 6859 857 6867 859
rect 6886 858 6887 862
rect 6928 859 6930 867
rect 6982 859 6985 868
rect 7000 864 7003 892
rect 7050 891 7076 892
rect 7074 861 7076 891
rect 7080 881 7088 892
rect 7159 879 7179 893
rect 7227 879 7241 894
rect 7270 881 7278 893
rect 7282 891 7316 893
rect 7135 876 7136 879
rect 7165 876 7166 879
rect 7179 877 7191 879
rect 7225 877 7227 879
rect 7179 875 7225 877
rect 7050 859 7076 861
rect 7080 859 7088 871
rect 7133 869 7134 871
rect 7162 868 7163 870
rect 7130 860 7132 866
rect 7159 860 7162 867
rect 7282 859 7284 891
rect 7314 873 7316 891
rect 7320 881 7328 893
rect 7402 891 7408 895
rect 7446 891 7448 895
rect 7460 891 7466 897
rect 7540 894 7546 900
rect 7569 896 7584 900
rect 7584 895 7585 896
rect 7598 895 7632 900
rect 7698 899 7704 903
rect 7748 901 7752 904
rect 7356 881 7357 889
rect 7400 881 7403 891
rect 7408 885 7414 891
rect 7440 881 7446 891
rect 7454 885 7460 891
rect 7543 883 7544 891
rect 7546 888 7552 894
rect 7585 893 7604 895
rect 7315 865 7316 872
rect 7350 870 7356 880
rect 7395 870 7400 881
rect 7344 868 7350 870
rect 7394 868 7395 870
rect 7434 869 7440 881
rect 7583 872 7586 892
rect 7592 888 7598 893
rect 7616 888 7632 895
rect 7704 894 7715 899
rect 7743 898 7747 900
rect 7740 897 7743 898
rect 7736 894 7740 897
rect 7760 895 7763 900
rect 7935 897 7970 904
rect 8016 902 8029 903
rect 7995 900 8013 902
rect 8034 900 8057 902
rect 7993 899 8005 900
rect 8057 899 8066 900
rect 8066 898 8067 899
rect 8091 898 8092 904
rect 7986 897 7993 898
rect 7715 886 7746 894
rect 7763 893 7765 895
rect 7765 891 7767 893
rect 7970 891 7993 897
rect 8067 894 8074 898
rect 8074 891 8080 894
rect 8092 891 8093 897
rect 7705 880 7746 886
rect 7767 886 7840 891
rect 7970 889 7992 891
rect 7767 881 7917 886
rect 7978 882 7986 889
rect 7992 887 7997 889
rect 7997 886 7999 887
rect 8080 886 8093 891
rect 8121 887 8124 903
rect 8179 901 8188 915
rect 8249 911 8250 914
rect 8276 909 8308 914
rect 8243 903 8247 906
rect 8250 903 8256 909
rect 8276 904 8314 909
rect 8345 904 8406 932
rect 8525 931 8528 936
rect 8524 922 8528 931
rect 8273 903 8314 904
rect 8343 903 8345 904
rect 8353 903 8354 904
rect 8230 901 8242 902
rect 8188 899 8192 901
rect 8210 900 8230 901
rect 8204 899 8210 900
rect 8230 895 8232 900
rect 8256 897 8262 903
rect 8290 899 8291 901
rect 8228 892 8230 895
rect 8227 891 8228 892
rect 7705 876 7722 880
rect 7746 876 7764 880
rect 7767 876 7787 881
rect 7839 876 7930 881
rect 7764 875 7930 876
rect 7971 875 7978 882
rect 7999 876 8023 886
rect 8080 882 8094 886
rect 8093 881 8096 882
rect 8093 878 8094 881
rect 8096 880 8097 881
rect 8023 875 8026 876
rect 7702 874 7704 875
rect 7763 874 7933 875
rect 7700 873 7702 874
rect 7761 873 7763 874
rect 7759 872 7761 873
rect 7764 872 7930 874
rect 7933 873 7941 874
rect 7941 872 7949 873
rect 7968 872 7971 875
rect 8026 874 8028 875
rect 8028 873 8031 874
rect 8031 872 8033 873
rect 8042 872 8054 878
rect 8097 875 8106 880
rect 8124 876 8126 886
rect 8215 882 8227 891
rect 8209 881 8215 882
rect 8181 880 8197 881
rect 8205 880 8209 881
rect 8274 880 8289 899
rect 8302 897 8308 903
rect 8339 901 8343 903
rect 8328 895 8339 901
rect 8352 899 8353 901
rect 8325 892 8328 895
rect 8324 891 8325 892
rect 8316 886 8324 891
rect 8153 875 8176 880
rect 8304 876 8336 886
rect 8349 880 8352 898
rect 8348 876 8349 880
rect 8384 878 8386 904
rect 8524 903 8525 922
rect 8539 915 8548 924
rect 8586 915 8595 924
rect 8530 906 8535 915
rect 8600 906 8604 915
rect 8505 881 8524 901
rect 7338 866 7344 868
rect 7433 867 7434 868
rect 7432 866 7433 867
rect 7337 865 7338 866
rect 7315 860 7337 865
rect 7391 862 7394 866
rect 7316 859 7337 860
rect 7388 859 7394 862
rect 6858 855 6867 857
rect 6783 850 6792 853
rect 6795 850 6801 853
rect 6846 852 6847 853
rect 6856 852 6867 855
rect 6803 851 6851 852
rect 6854 851 6856 852
rect 6803 850 6854 851
rect 6858 850 6867 852
rect 6793 847 6801 850
rect 6793 842 6797 847
rect 6846 840 6847 850
rect 6882 845 6886 858
rect 6925 846 6928 858
rect 6978 846 6982 858
rect 6998 851 7004 857
rect 7027 856 7031 859
rect 7321 858 7322 859
rect 7004 845 7010 851
rect 7022 845 7027 856
rect 7056 851 7062 857
rect 7129 855 7130 858
rect 7158 855 7159 858
rect 7388 857 7391 859
rect 7390 856 7391 857
rect 7386 855 7390 856
rect 7050 845 7056 851
rect 7064 847 7076 855
rect 7280 853 7281 855
rect 7127 851 7128 853
rect 6878 841 6882 845
rect 6924 841 6925 845
rect 6976 842 6978 845
rect 6876 840 6878 841
rect 7020 840 7022 845
rect 7124 841 7127 850
rect 7154 841 7157 850
rect 7281 841 7283 849
rect 7322 842 7323 849
rect 7383 847 7390 855
rect 7380 842 7383 847
rect 7386 845 7390 847
rect 7420 845 7432 865
rect 7544 859 7546 872
rect 7697 871 7699 872
rect 7757 871 7759 872
rect 7380 841 7382 842
rect 7377 840 7380 841
rect 7384 840 7386 845
rect 7417 844 7424 845
rect 7579 844 7583 870
rect 7692 868 7697 871
rect 7752 869 7756 871
rect 7840 869 8064 872
rect 8106 871 8112 875
rect 8143 871 8153 875
rect 8267 872 8270 876
rect 8301 875 8336 876
rect 8112 869 8118 871
rect 8125 869 8153 871
rect 7749 867 7751 868
rect 7689 866 7691 867
rect 7747 866 7749 867
rect 7856 866 8064 869
rect 8118 868 8119 869
rect 8125 868 8143 869
rect 8119 867 8123 868
rect 8138 867 8141 868
rect 7679 860 7689 866
rect 7737 862 7747 866
rect 7856 863 8066 866
rect 7969 862 7978 863
rect 8052 862 8074 863
rect 8095 862 8096 867
rect 8259 863 8267 872
rect 8314 869 8315 874
rect 8434 873 8445 874
rect 8462 873 8473 874
rect 8434 872 8442 873
rect 8466 872 8473 873
rect 7978 860 7981 862
rect 7674 857 7679 860
rect 7665 852 7674 857
rect 7981 852 7996 860
rect 8052 854 8066 862
rect 8074 856 8107 862
rect 8255 857 8259 862
rect 8182 856 8194 857
rect 8107 855 8113 856
rect 8131 855 8153 856
rect 8113 854 8153 855
rect 8174 854 8194 856
rect 7663 851 7665 852
rect 7996 851 7998 852
rect 7660 850 7663 851
rect 7998 850 8000 851
rect 7625 849 7631 850
rect 7658 849 7660 850
rect 7607 844 7658 849
rect 7671 844 7677 850
rect 7721 845 7724 849
rect 8001 845 8009 849
rect 8052 846 8064 854
rect 8182 851 8214 854
rect 8183 847 8214 851
rect 8252 849 8254 856
rect 8252 847 8253 849
rect 7417 840 7421 844
rect 6798 836 6799 840
rect 6799 833 6800 836
rect 6846 832 6848 840
rect 6864 832 6876 840
rect 6923 838 6924 840
rect 6975 838 6976 840
rect 6922 832 6923 838
rect 6974 833 6975 838
rect 7017 832 7020 840
rect 7123 837 7124 840
rect 7122 833 7123 836
rect 7151 834 7153 840
rect 7323 837 7324 840
rect 7284 832 7288 837
rect 7375 832 7384 840
rect 7413 834 7421 840
rect 7413 832 7417 834
rect 6800 817 6808 832
rect 6846 825 6850 832
rect 6863 830 6864 832
rect 7016 830 7017 832
rect 6862 828 6863 830
rect 6921 828 6922 830
rect 6972 828 6973 830
rect 6861 825 6862 828
rect 6848 817 6850 825
rect 6920 824 6921 828
rect 6971 824 6972 827
rect 7014 824 7016 829
rect 6859 819 6861 824
rect 6919 819 6920 824
rect 6966 820 6971 824
rect 5217 805 5225 808
rect 5217 804 5219 805
rect 5220 800 5221 802
rect 5221 797 5223 800
rect 4978 790 4980 793
rect 4786 758 4802 763
rect 4851 773 4912 785
rect 4919 779 4932 790
rect 4918 774 4932 779
rect 4962 777 4980 790
rect 5071 789 5072 793
rect 5102 789 5103 795
rect 4962 774 4978 777
rect 4851 759 4916 773
rect 4882 758 4898 759
rect 4900 758 4916 759
rect 4943 758 4944 760
rect 4978 758 4994 774
rect 5072 767 5076 785
rect 5103 779 5104 788
rect 5152 787 5154 794
rect 5217 790 5218 794
rect 5223 791 5226 797
rect 5258 792 5274 808
rect 5308 802 5336 808
rect 5372 806 5392 816
rect 6808 809 6812 817
rect 6850 811 6851 817
rect 6858 815 6859 819
rect 6918 815 6919 819
rect 6966 815 6970 820
rect 7012 819 7014 824
rect 6857 809 6858 814
rect 6916 809 6918 814
rect 6966 809 6968 815
rect 7009 814 7012 818
rect 7062 814 7078 824
rect 7080 814 7096 824
rect 7116 817 7122 832
rect 7005 809 7009 814
rect 7049 809 7056 814
rect 7101 808 7109 814
rect 7114 811 7116 817
rect 7144 811 7151 832
rect 7285 827 7289 832
rect 7324 827 7330 832
rect 7373 830 7375 832
rect 7412 830 7413 832
rect 7143 809 7144 811
rect 7158 808 7174 824
rect 7274 822 7340 827
rect 7366 824 7373 830
rect 7409 825 7412 830
rect 7415 828 7417 832
rect 7546 832 7548 844
rect 7558 840 7570 844
rect 7586 842 7607 844
rect 7577 841 7586 842
rect 7572 840 7579 841
rect 7558 836 7572 840
rect 7274 821 7330 822
rect 7265 814 7274 821
rect 7285 818 7289 821
rect 7263 811 7265 814
rect 7288 811 7289 817
rect 7324 811 7330 821
rect 7340 814 7344 821
rect 7358 819 7366 824
rect 7406 819 7409 824
rect 7358 818 7360 819
rect 7358 815 7359 818
rect 7404 817 7406 819
rect 7403 816 7404 817
rect 7344 811 7345 814
rect 7357 812 7358 813
rect 7403 812 7406 816
rect 7436 812 7448 815
rect 7346 811 7355 812
rect 7181 808 7200 809
rect 7206 808 7208 809
rect 6813 804 6814 807
rect 5302 794 5336 802
rect 6814 799 6816 803
rect 6851 799 6852 803
rect 6854 800 6857 808
rect 6914 800 6916 808
rect 6816 794 6818 798
rect 6854 794 6856 800
rect 6912 794 6914 798
rect 5298 791 5300 794
rect 5308 790 5336 794
rect 5154 781 5155 787
rect 5217 782 5234 790
rect 5104 766 5109 779
rect 5156 774 5164 780
rect 5218 776 5234 782
rect 5290 779 5298 790
rect 5287 778 5298 779
rect 5302 788 5336 790
rect 5218 774 5228 776
rect 5164 773 5166 774
rect 5076 760 5077 766
rect 5109 759 5111 766
rect 5166 765 5180 773
rect 5218 766 5219 774
rect 5234 768 5239 776
rect 5287 770 5296 778
rect 5215 765 5219 766
rect 5161 764 5194 765
rect 5215 764 5225 765
rect 5161 759 5167 764
rect 4711 756 4717 758
rect 4788 757 4802 758
rect 4914 757 4917 758
rect 4796 756 4849 757
rect 4629 754 4630 756
rect 4711 754 4720 756
rect 4393 738 4399 739
rect 4439 738 4445 744
rect 4479 738 4488 747
rect 4526 738 4535 747
rect 4618 746 4632 754
rect 4706 747 4720 754
rect 4791 750 4855 756
rect 4918 750 4933 756
rect 4940 754 4941 756
rect 4982 752 4983 753
rect 4706 746 4711 747
rect 4632 745 4635 746
rect 4145 734 4146 736
rect 4147 727 4150 733
rect 4219 731 4234 736
rect 4387 732 4393 738
rect 4445 733 4451 738
rect 4499 734 4511 738
rect 4552 734 4568 744
rect 4630 742 4631 745
rect 4635 742 4674 745
rect 4704 743 4711 746
rect 4797 745 4812 750
rect 4843 747 4852 750
rect 4797 744 4803 745
rect 4843 744 4849 747
rect 4631 740 4674 742
rect 4635 737 4674 740
rect 4697 739 4704 743
rect 4706 739 4711 743
rect 4852 742 4866 747
rect 4933 745 4946 750
rect 4982 747 4990 752
rect 5078 751 5079 756
rect 5112 750 5115 756
rect 5167 753 5173 759
rect 5178 758 5194 764
rect 5196 758 5212 764
rect 5219 759 5225 764
rect 5239 762 5242 768
rect 5278 761 5287 770
rect 5213 753 5219 759
rect 5244 756 5246 760
rect 5274 757 5275 758
rect 4932 742 4934 745
rect 4946 742 4952 745
rect 4983 744 4990 747
rect 5079 746 5080 750
rect 5115 744 5117 750
rect 5201 745 5204 747
rect 4992 742 4993 744
rect 5246 743 5254 756
rect 5275 754 5278 757
rect 5290 756 5298 768
rect 5302 758 5304 788
rect 5333 787 5336 788
rect 5340 779 5383 791
rect 6819 785 6822 793
rect 6853 790 6855 793
rect 6856 790 6870 794
rect 6853 786 6870 790
rect 5334 776 5383 779
rect 5334 770 5343 776
rect 5354 774 5370 776
rect 5383 774 5404 776
rect 6822 775 6827 785
rect 5343 764 5352 770
rect 5346 763 5352 764
rect 5370 768 5404 774
rect 6827 771 6828 775
rect 6854 774 6870 786
rect 6904 790 6912 794
rect 6950 792 6966 808
rect 7000 801 7005 808
rect 7045 801 7049 808
rect 7101 807 7112 808
rect 7142 807 7158 808
rect 7208 807 7209 808
rect 7257 807 7263 810
rect 7330 809 7331 811
rect 7285 808 7287 809
rect 7345 808 7355 811
rect 7402 808 7403 812
rect 7436 808 7452 812
rect 7454 808 7470 824
rect 7472 808 7488 824
rect 7546 820 7554 832
rect 7558 831 7574 832
rect 7558 830 7568 831
rect 7490 808 7499 812
rect 7549 810 7550 811
rect 7274 807 7284 808
rect 7101 806 7113 807
rect 7108 804 7113 806
rect 7000 792 7003 801
rect 6904 774 6920 790
rect 6950 774 6966 790
rect 7000 787 7016 790
rect 6995 781 7016 787
rect 7036 787 7045 801
rect 7108 792 7112 804
rect 7141 803 7158 807
rect 7209 806 7212 807
rect 7140 799 7141 803
rect 7138 794 7140 798
rect 7142 792 7158 803
rect 7181 798 7193 806
rect 7212 803 7215 806
rect 7235 803 7274 807
rect 7331 803 7332 807
rect 7342 803 7357 808
rect 7436 807 7453 808
rect 7458 807 7470 808
rect 7196 799 7235 803
rect 7246 799 7252 803
rect 7257 799 7263 803
rect 7332 799 7333 803
rect 7036 785 7047 787
rect 7056 785 7068 791
rect 7108 785 7109 792
rect 7136 788 7138 792
rect 7025 783 7047 785
rect 7057 783 7068 785
rect 7107 783 7112 785
rect 7019 781 7024 783
rect 6989 775 6995 781
rect 7000 774 7016 781
rect 7034 779 7036 783
rect 7041 781 7047 783
rect 7068 781 7072 783
rect 7047 775 7053 781
rect 7056 778 7068 779
rect 6856 771 6860 774
rect 5347 759 5350 763
rect 5370 758 5386 768
rect 5404 762 5421 768
rect 5407 758 5413 762
rect 5421 760 5427 762
rect 5427 758 5431 760
rect 5453 758 5459 764
rect 5302 757 5317 758
rect 5302 756 5321 757
rect 5278 750 5283 754
rect 5318 752 5336 756
rect 5353 753 5359 756
rect 5401 753 5407 758
rect 5302 750 5336 752
rect 5359 751 5407 753
rect 5459 752 5465 758
rect 6828 754 6836 771
rect 6860 754 6867 771
rect 6870 758 6886 774
rect 6888 758 6904 774
rect 6966 772 6974 774
rect 6992 772 7000 774
rect 7066 772 7068 778
rect 7072 772 7080 779
rect 7105 778 7107 783
rect 7108 778 7112 783
rect 7105 774 7112 778
rect 7105 772 7107 774
rect 6966 758 6982 772
rect 6984 758 7000 772
rect 7047 757 7110 772
rect 7134 760 7136 786
rect 7142 774 7158 790
rect 7169 782 7177 794
rect 7181 793 7202 794
rect 7240 793 7246 799
rect 7181 792 7199 793
rect 7158 763 7162 767
rect 7169 763 7177 772
rect 7181 763 7183 792
rect 7334 788 7336 796
rect 7342 794 7364 803
rect 7342 792 7357 794
rect 7394 790 7402 806
rect 7432 804 7434 807
rect 7438 806 7452 807
rect 7436 803 7452 806
rect 7488 805 7504 808
rect 7486 803 7504 805
rect 7424 791 7432 803
rect 7434 801 7470 803
rect 7434 793 7454 801
rect 7467 800 7470 801
rect 7468 793 7470 800
rect 7474 799 7482 803
rect 7486 799 7508 803
rect 7488 794 7508 799
rect 7546 798 7554 810
rect 7558 800 7560 830
rect 7577 826 7579 840
rect 7619 838 7625 844
rect 7677 838 7683 844
rect 7716 841 7721 845
rect 8009 841 8014 845
rect 8008 832 8016 841
rect 8020 834 8022 839
rect 8052 834 8054 846
rect 8312 845 8314 865
rect 8346 863 8348 872
rect 8383 863 8384 872
rect 8434 871 8436 872
rect 8472 871 8473 872
rect 8505 868 8519 881
rect 8498 866 8511 868
rect 8498 865 8510 866
rect 8539 865 8544 866
rect 8345 857 8346 862
rect 8343 849 8344 855
rect 8064 844 8067 845
rect 8020 832 8054 834
rect 8058 840 8067 844
rect 8058 832 8066 840
rect 8067 832 8071 840
rect 8071 830 8072 832
rect 7592 826 7593 830
rect 7703 829 7706 830
rect 7679 827 7714 829
rect 7577 818 7578 826
rect 7675 825 7679 827
rect 7673 824 7675 825
rect 7593 812 7595 824
rect 7578 800 7581 811
rect 7646 808 7673 824
rect 7677 812 7681 817
rect 7687 812 7703 827
rect 7714 824 7739 827
rect 7682 811 7703 812
rect 7558 798 7592 800
rect 7578 795 7581 798
rect 7336 778 7339 788
rect 7339 769 7341 778
rect 7342 774 7357 790
rect 7394 774 7408 790
rect 7431 781 7432 788
rect 7341 765 7342 769
rect 7158 762 7183 763
rect 7212 762 7215 763
rect 7158 760 7215 762
rect 7158 758 7174 760
rect 7342 759 7343 763
rect 5283 749 5319 750
rect 5302 744 5314 749
rect 5369 744 5380 749
rect 6836 746 6839 754
rect 6867 748 6872 754
rect 6872 745 6876 748
rect 7066 745 7068 757
rect 7071 745 7105 757
rect 7110 756 7112 757
rect 7219 756 7246 759
rect 7343 757 7344 759
rect 7358 758 7374 772
rect 7376 758 7392 772
rect 7424 769 7432 781
rect 7436 774 7454 793
rect 7488 792 7504 794
rect 7488 774 7504 790
rect 7534 774 7549 790
rect 7551 775 7553 792
rect 7558 786 7570 794
rect 7580 786 7592 794
rect 7594 790 7595 808
rect 7681 805 7691 811
rect 7739 808 7880 824
rect 7942 808 7958 824
rect 7960 808 7976 824
rect 8020 820 8032 828
rect 8042 820 8054 828
rect 8072 826 8073 830
rect 8098 828 8100 845
rect 8020 810 8022 820
rect 8073 816 8076 824
rect 8100 819 8101 828
rect 8128 819 8131 845
rect 8170 833 8176 845
rect 8217 843 8219 844
rect 8342 843 8343 847
rect 8253 838 8254 843
rect 8220 827 8221 836
rect 8254 827 8255 836
rect 8310 825 8312 840
rect 8341 837 8342 843
rect 8339 827 8341 836
rect 8381 829 8383 862
rect 8494 855 8510 865
rect 8547 864 8551 868
rect 8431 845 8494 855
rect 8539 851 8547 864
rect 8422 844 8431 845
rect 8416 842 8422 844
rect 8414 840 8416 842
rect 8170 811 8176 823
rect 8338 821 8339 826
rect 8379 820 8381 827
rect 8395 825 8414 840
rect 8394 824 8395 825
rect 8222 817 8223 820
rect 8255 816 8256 820
rect 8223 811 8228 816
rect 8256 811 8257 816
rect 8309 811 8310 818
rect 8323 811 8329 817
rect 8337 816 8338 820
rect 8378 818 8379 820
rect 8386 818 8394 824
rect 8335 812 8337 816
rect 8369 811 8375 817
rect 8377 816 8386 818
rect 8376 811 8386 816
rect 8132 808 8133 810
rect 8224 808 8225 810
rect 7686 803 7691 805
rect 7811 803 7820 808
rect 7858 803 7867 808
rect 7598 802 7607 803
rect 7596 798 7604 802
rect 7607 799 7622 802
rect 7622 798 7625 799
rect 7619 792 7625 798
rect 7677 792 7683 798
rect 7691 794 7700 803
rect 7802 794 7811 803
rect 7867 794 7876 803
rect 7793 792 7800 793
rect 7625 790 7631 792
rect 7436 772 7470 774
rect 7483 772 7488 774
rect 7581 772 7584 786
rect 7594 774 7600 790
rect 7625 786 7646 790
rect 7671 786 7677 792
rect 7787 791 7793 792
rect 7844 791 7848 793
rect 7880 792 7896 808
rect 7926 792 7942 808
rect 7953 803 7959 808
rect 7953 802 7968 803
rect 7947 796 7953 802
rect 7976 798 7992 808
rect 7999 802 8005 808
rect 7952 791 7953 793
rect 7985 791 7990 798
rect 8005 796 8011 802
rect 8023 800 8024 808
rect 7785 790 7787 791
rect 7784 787 7785 790
rect 7849 789 7851 790
rect 7630 774 7646 786
rect 7697 778 7724 781
rect 7680 774 7697 778
rect 7724 774 7732 778
rect 7436 769 7488 772
rect 7549 769 7555 772
rect 7584 771 7588 772
rect 7436 757 7440 765
rect 7472 758 7488 769
rect 7550 762 7567 769
rect 7584 762 7594 771
rect 7550 758 7566 762
rect 7567 760 7572 762
rect 7576 760 7588 762
rect 7572 759 7588 760
rect 7568 758 7588 759
rect 7646 758 7662 774
rect 7732 772 7735 774
rect 7800 772 7806 778
rect 7809 772 7811 779
rect 7851 772 7852 778
rect 7880 774 7896 790
rect 7926 774 7942 790
rect 7944 779 7953 791
rect 7735 763 7755 772
rect 7784 767 7785 769
rect 7794 766 7800 772
rect 7852 766 7858 772
rect 7873 763 7880 774
rect 7755 762 7757 763
rect 7757 759 7763 762
rect 7112 751 7133 756
rect 7133 747 7149 751
rect 7181 748 7193 756
rect 7344 754 7345 756
rect 7240 747 7246 753
rect 7271 747 7326 753
rect 7345 750 7346 754
rect 7346 747 7348 748
rect 7355 747 7364 756
rect 7434 747 7440 756
rect 7492 747 7498 753
rect 7499 747 7508 756
rect 7553 751 7556 758
rect 5380 743 5382 744
rect 4866 739 4875 742
rect 4952 741 4954 742
rect 5254 741 5255 743
rect 6839 741 6841 745
rect 4697 738 4711 739
rect 4684 737 4697 738
rect 4704 735 4706 738
rect 4875 735 4886 739
rect 4929 737 4930 739
rect 4886 734 4889 735
rect 4495 733 4577 734
rect 4445 732 4511 733
rect 4488 731 4511 732
rect 4234 726 4246 731
rect 4488 729 4495 731
rect 4499 730 4511 731
rect 4577 729 4580 732
rect 4696 731 4703 734
rect 4889 731 4898 734
rect 4926 733 4928 736
rect 4898 729 4905 731
rect 4921 729 4925 731
rect 4484 728 4488 729
rect 4477 726 4484 728
rect 4514 727 4515 729
rect 4580 728 4582 729
rect 3936 721 4007 723
rect 3760 719 3775 720
rect 3937 719 4007 721
rect 4039 719 4043 725
rect 4150 723 4152 726
rect 3763 716 3775 719
rect 3699 712 3704 716
rect 3776 714 3779 716
rect 3928 712 3936 719
rect 3938 717 3948 719
rect 3938 712 3942 717
rect 3704 696 3725 712
rect 3769 710 3793 712
rect 3773 705 3793 710
rect 3928 707 3938 712
rect 3935 705 3938 707
rect 3725 695 3727 696
rect 3731 689 3732 692
rect 3729 678 3736 687
rect 3773 680 3775 705
rect 3779 700 3787 705
rect 3793 699 3799 705
rect 3933 701 3935 705
rect 3927 699 3935 701
rect 3799 694 3805 699
rect 3927 695 3933 699
rect 3805 692 3808 694
rect 3741 678 3775 680
rect 3779 678 3787 690
rect 3808 688 3809 692
rect 3921 689 3927 695
rect 3931 692 3932 694
rect 3930 688 3931 691
rect 3940 689 3942 712
rect 3972 715 4027 719
rect 3972 701 3995 715
rect 4003 713 4027 715
rect 4047 713 4048 715
rect 4008 708 4027 713
rect 4048 708 4052 713
rect 4152 710 4159 723
rect 4246 722 4276 726
rect 4495 724 4511 726
rect 4246 714 4288 722
rect 4015 701 4027 708
rect 4052 706 4053 708
rect 4159 705 4162 710
rect 4240 709 4289 710
rect 3972 695 3979 701
rect 3972 693 3985 695
rect 3972 689 3974 693
rect 3979 689 3985 693
rect 3990 691 3999 700
rect 4018 696 4027 701
rect 4058 696 4061 701
rect 4021 691 4027 696
rect 3929 685 3930 687
rect 3973 685 3974 689
rect 3991 687 4008 691
rect 4024 689 4027 691
rect 4061 689 4067 696
rect 4162 695 4199 705
rect 4240 702 4254 709
rect 4270 708 4289 709
rect 4286 703 4289 708
rect 4239 699 4240 701
rect 4199 693 4205 695
rect 4237 694 4239 699
rect 4205 692 4210 693
rect 4236 692 4237 694
rect 4026 687 4027 689
rect 3992 686 4008 687
rect 4067 686 4069 689
rect 4210 688 4226 692
rect 4226 687 4228 688
rect 3809 680 3811 685
rect 3928 680 3929 685
rect 3994 682 3997 686
rect 3999 682 4008 686
rect 4000 680 4001 682
rect 3736 676 3737 678
rect 3740 676 3741 678
rect 3927 676 3928 678
rect 4001 677 4002 680
rect 3736 660 3740 676
rect 3776 674 3779 676
rect 3741 666 3753 674
rect 3763 666 3775 674
rect 3811 660 3815 676
rect 3735 654 3736 658
rect 3815 657 3816 660
rect 3735 630 3737 654
rect 3815 630 3816 654
rect 3927 649 3979 663
rect 4000 662 4002 675
rect 4029 672 4041 685
rect 4069 672 4081 686
rect 4231 685 4237 687
rect 4237 683 4245 685
rect 4242 681 4246 683
rect 4242 676 4249 681
rect 4286 678 4288 703
rect 4289 697 4290 702
rect 4292 698 4300 710
rect 4445 694 4473 695
rect 4509 694 4511 724
rect 4515 714 4523 726
rect 4582 712 4584 728
rect 4905 727 4911 729
rect 4918 727 4921 729
rect 4638 720 4644 726
rect 4696 720 4702 726
rect 4902 723 4922 727
rect 4954 723 4975 741
rect 4980 738 4991 740
rect 4902 721 4918 723
rect 4897 720 4902 721
rect 4922 720 4930 723
rect 4644 714 4650 720
rect 4690 714 4696 720
rect 4890 717 4897 720
rect 4930 719 4933 720
rect 4975 719 4980 723
rect 4885 716 4890 717
rect 4933 716 4939 719
rect 4980 716 4984 719
rect 4988 716 4990 738
rect 4991 737 4992 738
rect 4994 737 5002 740
rect 4992 734 5002 737
rect 4994 729 5002 734
rect 5081 733 5082 741
rect 5118 737 5121 741
rect 5082 729 5083 733
rect 5111 729 5123 737
rect 5133 729 5145 737
rect 5208 729 5221 741
rect 4994 728 5003 729
rect 4999 726 5003 728
rect 4994 716 5002 718
rect 4876 713 4885 716
rect 4871 711 4876 713
rect 4290 693 4291 694
rect 4465 692 4473 694
rect 4477 692 4511 694
rect 4515 692 4523 704
rect 4582 694 4584 710
rect 4855 706 4871 711
rect 4939 706 4950 716
rect 4984 707 5002 716
rect 4966 706 5002 707
rect 5003 706 5026 726
rect 5083 724 5090 729
rect 5107 727 5110 729
rect 5123 725 5124 729
rect 5130 725 5136 729
rect 5084 723 5090 724
rect 5099 723 5107 725
rect 5111 723 5157 725
rect 5078 717 5084 723
rect 5111 717 5113 723
rect 5136 717 5142 723
rect 5143 717 5157 723
rect 5082 713 5084 714
rect 5080 709 5082 713
rect 4839 701 4855 706
rect 4950 705 4957 706
rect 4995 705 5028 706
rect 4950 702 4958 705
rect 4932 701 4966 702
rect 4992 701 5053 705
rect 5143 702 5145 717
rect 5149 713 5164 717
rect 5152 705 5164 713
rect 5221 712 5240 729
rect 5255 715 5289 741
rect 5384 723 5407 741
rect 6876 740 6884 745
rect 7102 742 7103 745
rect 7149 742 7169 747
rect 7169 741 7174 742
rect 7246 741 7252 747
rect 7292 741 7298 747
rect 7068 740 7070 741
rect 6841 737 6843 740
rect 6884 737 6889 740
rect 7058 739 7068 740
rect 7047 738 7068 739
rect 7174 738 7178 741
rect 7299 738 7308 747
rect 7346 745 7355 747
rect 7346 742 7361 745
rect 7346 738 7355 742
rect 7361 740 7365 742
rect 7440 741 7452 747
rect 7486 741 7499 747
rect 7555 744 7556 751
rect 7365 739 7368 740
rect 6889 736 6891 737
rect 7056 736 7075 738
rect 6844 733 6845 736
rect 6891 733 6895 736
rect 6845 727 6848 733
rect 6895 731 6899 733
rect 6899 729 6902 731
rect 6989 729 6995 735
rect 7047 729 7053 735
rect 7056 733 7093 736
rect 7100 733 7101 736
rect 7067 729 7093 733
rect 7096 729 7100 731
rect 7132 729 7133 730
rect 6902 726 6906 729
rect 6848 720 6852 726
rect 6906 720 6916 726
rect 6919 720 6931 724
rect 6995 723 7001 729
rect 7041 723 7047 729
rect 7093 726 7133 729
rect 7093 723 7132 726
rect 7178 725 7195 738
rect 7299 737 7300 738
rect 7368 736 7375 739
rect 7443 738 7452 741
rect 7490 738 7499 741
rect 7549 739 7556 744
rect 7584 742 7588 758
rect 7626 747 7635 756
rect 7691 747 7700 756
rect 7763 754 7774 759
rect 7867 758 7880 763
rect 7942 769 7951 774
rect 7952 769 7953 779
rect 7942 763 7953 769
rect 7956 763 7958 791
rect 8024 790 8026 791
rect 8022 785 8026 790
rect 8075 790 8076 808
rect 8182 799 8194 803
rect 8204 799 8216 803
rect 8226 796 8227 799
rect 8257 796 8258 805
rect 8308 799 8309 808
rect 8317 805 8323 811
rect 8375 808 8381 811
rect 8430 808 8446 824
rect 9019 819 9020 1015
rect 9209 819 9210 1015
rect 9295 819 9296 1015
rect 9568 819 9569 1015
rect 9766 820 9767 1016
rect 10156 1014 10160 1019
rect 10794 1014 10801 1019
rect 10881 1018 10890 1027
rect 10946 1024 11042 1027
rect 11383 1023 11491 1037
rect 11241 1015 11257 1022
rect 11259 1015 11275 1022
rect 10801 1007 10813 1014
rect 11231 1013 11243 1015
rect 11253 1013 11265 1015
rect 11271 1013 11275 1015
rect 11459 1013 11475 1022
rect 11491 1021 11509 1023
rect 11510 1017 11517 1020
rect 11517 1013 11523 1017
rect 12163 1015 12164 1026
rect 12353 1015 12354 1026
rect 12439 1015 12440 1026
rect 12712 1015 12713 1026
rect 12910 1016 12911 1027
rect 13338 1023 13439 1034
rect 13625 1033 13889 1034
rect 13889 1023 13944 1033
rect 14047 1027 14056 1036
rect 14094 1027 14103 1036
rect 14397 1034 14519 1037
rect 14369 1033 14386 1034
rect 14199 1027 14369 1033
rect 13323 1021 13338 1023
rect 13317 1019 13323 1021
rect 13946 1019 13951 1021
rect 11231 1008 11275 1013
rect 11418 1008 11455 1009
rect 11523 1008 11526 1013
rect 11227 1006 11229 1008
rect 11231 1006 11363 1008
rect 10282 1005 10636 1006
rect 10262 1003 10280 1005
rect 10722 1003 10735 1005
rect 10814 1003 10817 1005
rect 11225 1003 11363 1006
rect 10206 1000 10262 1003
rect 10080 992 10092 1000
rect 10102 992 10114 1000
rect 10178 994 10262 1000
rect 10735 994 10745 1003
rect 10178 993 10206 994
rect 10076 989 10078 992
rect 10178 991 10197 993
rect 10746 991 10749 993
rect 10118 988 10122 989
rect 10068 977 10076 988
rect 10079 986 10114 988
rect 10077 977 10079 983
rect 10068 976 10077 977
rect 10076 972 10077 976
rect 10075 971 10076 972
rect 10073 966 10075 969
rect 9948 964 10013 965
rect 9940 956 9948 964
rect 10013 956 10017 964
rect 9939 950 9940 956
rect 10068 954 10076 966
rect 10080 956 10082 986
rect 10111 985 10114 986
rect 10113 979 10114 985
rect 10118 981 10126 988
rect 10122 980 10130 981
rect 10154 980 10155 990
rect 10178 980 10193 991
rect 10452 981 10489 983
rect 10130 979 10136 980
rect 10153 979 10154 980
rect 10178 979 10185 980
rect 10136 969 10198 979
rect 10206 972 10212 978
rect 10252 972 10258 978
rect 10452 977 10478 981
rect 10489 977 10494 981
rect 10749 980 10762 991
rect 10725 979 10739 980
rect 10446 972 10452 977
rect 10494 972 10503 977
rect 10707 972 10725 979
rect 10739 977 10746 979
rect 10817 977 10838 1003
rect 11219 996 11363 1003
rect 11379 1006 11480 1008
rect 11379 996 11491 1006
rect 11180 990 11241 996
rect 11145 987 11180 990
rect 10958 981 11145 987
rect 11231 986 11241 990
rect 10746 972 10761 977
rect 10200 969 10206 972
rect 10207 970 10264 972
rect 10503 971 10504 972
rect 10341 970 10344 971
rect 10362 970 10365 971
rect 10444 970 10445 971
rect 10504 970 10507 971
rect 10207 969 10215 970
rect 10178 968 10215 969
rect 10080 954 10114 956
rect 10069 951 10071 954
rect 10065 939 10069 950
rect 10080 942 10092 950
rect 10105 945 10114 954
rect 10152 952 10153 955
rect 10178 951 10183 968
rect 10200 966 10215 968
rect 10258 966 10264 970
rect 10337 967 10341 970
rect 10365 967 10370 970
rect 10507 968 10508 970
rect 10699 969 10707 972
rect 10736 971 10761 972
rect 10770 971 10774 972
rect 10732 970 10736 971
rect 10746 970 10783 971
rect 10508 967 10511 968
rect 10206 964 10215 966
rect 10206 951 10211 964
rect 10259 955 10278 958
rect 10313 955 10337 967
rect 10370 959 10388 967
rect 10443 959 10444 967
rect 10115 948 10125 950
rect 10125 947 10128 948
rect 10130 945 10139 947
rect 10103 942 10105 945
rect 10139 943 10150 945
rect 10151 943 10152 951
rect 10178 943 10184 951
rect 10102 939 10103 942
rect 10150 938 10184 943
rect 10016 924 10017 938
rect 9966 915 9975 924
rect 10013 920 10022 924
rect 10013 915 10027 920
rect 9957 912 9966 915
rect 9957 911 9960 912
rect 9950 908 9959 911
rect 9938 907 9959 908
rect 9938 905 9956 907
rect 9996 905 10002 911
rect 10016 906 10031 915
rect 10056 908 10065 937
rect 9938 900 9950 905
rect 9934 898 9937 900
rect 9938 899 9939 900
rect 9944 899 9950 900
rect 10002 899 10008 905
rect 10015 904 10027 906
rect 10054 904 10056 908
rect 10094 907 10102 938
rect 10151 926 10152 938
rect 10178 935 10206 938
rect 10178 931 10208 935
rect 10210 931 10211 951
rect 10278 946 10340 955
rect 10388 952 10396 959
rect 10442 951 10443 958
rect 10511 954 10515 967
rect 10691 966 10699 969
rect 10729 968 10732 970
rect 10725 967 10729 968
rect 10720 965 10725 967
rect 10746 965 10761 970
rect 10770 969 10774 970
rect 10783 969 10784 970
rect 10840 969 10845 975
rect 10881 971 10890 980
rect 10946 978 10958 981
rect 10946 971 10955 978
rect 11225 972 11241 986
rect 11264 972 11265 996
rect 11270 991 11291 996
rect 11275 990 11291 991
rect 11408 989 11414 996
rect 11460 989 11466 996
rect 11480 990 11491 996
rect 11526 990 11535 1008
rect 11275 972 11291 988
rect 11408 985 11416 989
rect 11414 983 11416 985
rect 11324 974 11352 978
rect 11354 974 11365 978
rect 10774 965 10779 969
rect 10784 965 10786 968
rect 10845 965 10848 969
rect 10686 964 10690 965
rect 10761 964 10764 965
rect 10786 964 10787 965
rect 10682 962 10686 964
rect 10651 950 10682 962
rect 10766 959 10770 962
rect 10781 960 10785 963
rect 10890 962 10899 971
rect 10923 961 10926 963
rect 10937 962 10946 971
rect 11231 970 11265 972
rect 11274 971 11275 972
rect 11321 971 11324 974
rect 11270 970 11275 971
rect 11320 970 11321 971
rect 11231 968 11275 970
rect 11318 969 11320 970
rect 11227 965 11228 967
rect 11001 961 11010 963
rect 10918 959 10923 961
rect 10296 945 10306 946
rect 10328 945 10329 946
rect 10292 943 10296 945
rect 10340 943 10360 946
rect 10441 943 10442 950
rect 10514 943 10515 950
rect 10563 943 10569 949
rect 10609 948 10615 949
rect 10646 948 10651 950
rect 10609 947 10646 948
rect 10609 943 10615 947
rect 10701 946 10707 952
rect 10747 946 10753 952
rect 10769 950 10770 959
rect 10916 958 10918 959
rect 11012 958 11018 961
rect 10787 955 10791 958
rect 10855 955 10857 958
rect 10791 946 10801 955
rect 10280 931 10288 943
rect 10292 941 10326 943
rect 10178 928 10239 931
rect 10178 917 10184 928
rect 10206 926 10239 928
rect 10200 925 10239 926
rect 10258 925 10264 926
rect 10200 921 10264 925
rect 10200 920 10286 921
rect 10178 915 10185 917
rect 10178 913 10187 915
rect 10206 914 10212 920
rect 10252 914 10258 920
rect 10261 917 10286 920
rect 10270 915 10286 917
rect 10275 913 10286 915
rect 10292 913 10294 941
rect 10323 939 10326 941
rect 10178 909 10193 913
rect 10280 909 10294 913
rect 10324 909 10326 939
rect 10330 931 10338 943
rect 10360 934 10423 943
rect 10557 938 10563 943
rect 10575 941 10611 943
rect 10575 939 10580 941
rect 10516 937 10563 938
rect 10577 937 10580 939
rect 10615 937 10621 943
rect 10695 940 10701 946
rect 10753 940 10759 946
rect 10768 938 10769 943
rect 10801 942 10806 946
rect 10857 942 10869 955
rect 11018 951 11031 958
rect 11241 956 11257 968
rect 11259 956 11275 968
rect 11314 965 11318 968
rect 11312 963 11314 965
rect 11310 961 11312 963
rect 11365 961 11378 974
rect 11414 967 11417 983
rect 11416 961 11417 967
rect 11420 967 11421 989
rect 11459 985 11466 989
rect 11487 987 11489 990
rect 11459 983 11460 985
rect 11480 984 11481 986
rect 11420 963 11422 967
rect 11453 963 11454 966
rect 11458 965 11460 983
rect 11489 981 11492 987
rect 11492 979 11493 981
rect 11494 975 11495 977
rect 11495 972 11496 975
rect 11535 973 11543 990
rect 11497 965 11500 969
rect 11420 961 11424 963
rect 11458 962 11459 965
rect 11500 963 11501 965
rect 11306 958 11309 961
rect 11378 959 11381 961
rect 11304 953 11306 958
rect 11381 957 11383 959
rect 11139 952 11176 953
rect 11303 952 11304 953
rect 11383 952 11385 957
rect 11411 955 11417 961
rect 11424 959 11430 961
rect 11431 957 11437 959
rect 11457 957 11463 961
rect 11501 960 11502 963
rect 11502 958 11503 960
rect 11437 956 11463 957
rect 11139 951 11164 952
rect 11176 951 11177 952
rect 11302 951 11303 952
rect 11033 948 11037 951
rect 11104 948 11131 951
rect 11179 948 11186 951
rect 11300 948 11302 951
rect 11186 943 11197 948
rect 11233 945 11234 947
rect 11298 943 11300 948
rect 11385 944 11388 951
rect 11405 949 11411 955
rect 11437 951 11481 956
rect 11503 955 11505 958
rect 11463 949 11469 951
rect 11505 948 11508 955
rect 11197 942 11201 943
rect 10869 939 10870 942
rect 11201 939 11206 942
rect 11206 938 11208 939
rect 11234 938 11237 943
rect 11268 941 11269 943
rect 11297 942 11298 943
rect 11508 942 11511 948
rect 11543 943 11544 973
rect 11651 951 11667 954
rect 11579 943 11602 951
rect 11667 943 11674 951
rect 11296 940 11297 942
rect 11295 939 11296 940
rect 11511 939 11512 942
rect 10516 936 10559 937
rect 10440 934 10441 936
rect 10462 934 10516 936
rect 10396 922 10411 934
rect 10423 933 10462 934
rect 10440 929 10441 933
rect 10572 929 10575 936
rect 10699 933 10701 934
rect 10093 904 10094 906
rect 10153 905 10154 909
rect 10159 903 10165 909
rect 10178 903 10197 909
rect 10205 903 10211 909
rect 10013 899 10015 903
rect 10053 899 10054 903
rect 10012 897 10013 899
rect 10052 897 10053 899
rect 9926 884 9934 896
rect 9938 894 9956 896
rect 10011 895 10012 896
rect 10091 895 10093 903
rect 10153 897 10159 903
rect 10178 897 10217 903
rect 10219 897 10231 905
rect 10292 904 10309 909
rect 10396 904 10411 920
rect 10438 906 10440 928
rect 10300 903 10301 904
rect 10309 903 10313 904
rect 10328 903 10330 904
rect 10290 901 10291 903
rect 10301 899 10307 903
rect 10313 900 10332 903
rect 10437 900 10449 905
rect 10459 900 10471 905
rect 10512 904 10514 928
rect 10563 904 10572 928
rect 10695 925 10699 933
rect 10608 904 10611 909
rect 10649 908 10684 910
rect 10644 907 10649 908
rect 10684 907 10692 908
rect 10695 907 10697 915
rect 10719 909 10720 929
rect 10767 928 10768 936
rect 10764 917 10766 920
rect 10761 915 10763 916
rect 10758 913 10761 915
rect 10755 911 10758 913
rect 10753 910 10755 911
rect 10639 906 10644 907
rect 10692 906 10701 907
rect 10628 904 10639 906
rect 10562 900 10563 903
rect 10606 900 10608 903
rect 10616 901 10628 904
rect 10695 900 10697 906
rect 10719 904 10720 906
rect 10787 904 10803 920
rect 10811 915 10837 938
rect 10871 931 10877 938
rect 11208 937 11210 938
rect 11210 933 11226 937
rect 11226 932 11231 933
rect 11237 932 11242 938
rect 10881 920 10889 927
rect 10889 918 10896 920
rect 10896 915 10908 918
rect 10837 910 10843 915
rect 10908 914 10912 915
rect 10915 914 10916 929
rect 11231 927 11247 932
rect 11269 929 11272 938
rect 11294 937 11295 938
rect 11291 933 11294 937
rect 11289 932 11291 933
rect 11512 932 11513 938
rect 11541 932 11543 942
rect 11573 939 11579 943
rect 11674 939 11678 943
rect 11571 938 11573 939
rect 11678 938 11681 939
rect 11561 932 11571 938
rect 11678 936 11683 938
rect 11272 927 11273 928
rect 11286 927 11289 932
rect 11410 927 11411 929
rect 11242 923 11243 926
rect 11247 924 11284 927
rect 10974 921 11005 922
rect 10965 920 10974 921
rect 11005 920 11012 921
rect 11272 920 11273 924
rect 10936 917 10965 920
rect 11012 917 11027 920
rect 10934 916 10936 917
rect 10931 915 10934 916
rect 11027 915 11035 917
rect 11244 915 11245 917
rect 11273 915 11274 920
rect 11278 915 11287 924
rect 11325 915 11334 924
rect 11409 922 11410 927
rect 11408 920 11409 922
rect 11407 918 11408 920
rect 11406 916 11407 918
rect 10924 914 10931 915
rect 11035 914 11044 915
rect 11269 914 11278 915
rect 10912 911 11278 914
rect 10915 910 10916 911
rect 10918 910 10920 911
rect 11054 910 11062 911
rect 10843 909 10845 910
rect 10720 903 10721 904
rect 10784 903 10787 904
rect 10845 903 10853 909
rect 10914 908 10918 910
rect 11062 907 11075 910
rect 11075 906 11080 907
rect 10907 904 10912 906
rect 11080 904 11090 906
rect 10721 900 10724 903
rect 10774 900 10787 903
rect 10178 895 10233 897
rect 10307 895 10313 899
rect 10327 898 10328 900
rect 9926 862 9934 874
rect 9938 864 9940 894
rect 10010 893 10011 894
rect 10051 893 10052 894
rect 10178 893 10235 895
rect 10313 893 10314 895
rect 10326 894 10327 897
rect 10332 896 10501 900
rect 10560 897 10562 900
rect 10557 896 10563 897
rect 10603 896 10606 900
rect 10433 894 10435 896
rect 10437 895 10438 896
rect 10501 895 10563 896
rect 10005 889 10011 893
rect 10050 889 10051 893
rect 10090 889 10091 893
rect 10146 889 10153 893
rect 10178 892 10243 893
rect 9991 888 10011 889
rect 9991 878 10005 888
rect 10047 879 10050 889
rect 10088 878 10090 889
rect 10143 879 10146 889
rect 9978 868 9991 878
rect 10044 869 10047 878
rect 10087 875 10088 878
rect 10142 875 10143 878
rect 10085 868 10087 875
rect 10140 869 10142 875
rect 9975 866 9978 868
rect 9938 862 9941 864
rect 9972 862 9975 866
rect 10022 859 10031 868
rect 10043 866 10044 868
rect 10042 862 10043 866
rect 9937 857 9939 858
rect 9944 857 9950 859
rect 9938 853 9950 857
rect 10002 853 10008 859
rect 10014 857 10022 859
rect 10041 858 10042 862
rect 10083 859 10085 867
rect 10137 859 10140 868
rect 10155 864 10158 892
rect 10205 891 10231 892
rect 10229 861 10231 891
rect 10235 881 10243 892
rect 10314 879 10334 893
rect 10382 879 10396 894
rect 10425 881 10433 893
rect 10437 891 10471 893
rect 10290 876 10291 879
rect 10320 876 10321 879
rect 10334 877 10346 879
rect 10380 877 10382 879
rect 10334 875 10380 877
rect 10205 859 10231 861
rect 10235 859 10243 871
rect 10288 869 10289 871
rect 10317 868 10318 870
rect 10285 860 10287 866
rect 10314 860 10317 867
rect 10437 859 10439 891
rect 10469 873 10471 891
rect 10475 881 10483 893
rect 10557 891 10563 895
rect 10601 891 10603 895
rect 10615 891 10621 897
rect 10695 894 10701 900
rect 10724 896 10739 900
rect 10739 895 10740 896
rect 10753 895 10787 900
rect 10853 899 10859 903
rect 10903 901 10907 904
rect 10511 881 10512 889
rect 10555 881 10558 891
rect 10563 885 10569 891
rect 10595 881 10601 891
rect 10609 885 10615 891
rect 10698 883 10699 891
rect 10701 888 10707 894
rect 10740 893 10759 895
rect 10470 865 10471 872
rect 10505 870 10511 880
rect 10550 870 10555 881
rect 10499 868 10505 870
rect 10549 868 10550 870
rect 10589 869 10595 881
rect 10738 872 10741 892
rect 10747 888 10753 893
rect 10771 888 10787 895
rect 10859 894 10870 899
rect 10898 898 10902 900
rect 10895 897 10898 898
rect 10891 894 10895 897
rect 10915 895 10918 900
rect 11090 897 11125 904
rect 11171 902 11184 903
rect 11150 900 11168 902
rect 11189 900 11212 902
rect 11148 899 11160 900
rect 11212 899 11221 900
rect 11221 898 11222 899
rect 11246 898 11247 904
rect 11141 897 11148 898
rect 10870 886 10901 894
rect 10918 893 10920 895
rect 10920 891 10922 893
rect 11125 891 11148 897
rect 11222 894 11229 898
rect 11229 891 11235 894
rect 11247 891 11248 897
rect 10860 880 10901 886
rect 10922 886 10995 891
rect 11125 889 11147 891
rect 10922 881 11072 886
rect 11133 882 11141 889
rect 11147 887 11152 889
rect 11152 886 11154 887
rect 11235 886 11248 891
rect 11276 887 11279 903
rect 11334 901 11343 915
rect 11404 911 11405 914
rect 11431 909 11463 914
rect 11398 903 11402 906
rect 11405 903 11411 909
rect 11431 904 11469 909
rect 11500 904 11561 932
rect 11680 931 11683 936
rect 11679 922 11683 931
rect 11428 903 11469 904
rect 11498 903 11500 904
rect 11508 903 11509 904
rect 11385 901 11397 902
rect 11343 899 11347 901
rect 11365 900 11385 901
rect 11359 899 11365 900
rect 11385 895 11387 900
rect 11411 897 11417 903
rect 11445 899 11446 901
rect 11383 892 11385 895
rect 11382 891 11383 892
rect 10860 876 10877 880
rect 10901 876 10919 880
rect 10922 876 10942 881
rect 10994 876 11085 881
rect 10919 875 11085 876
rect 11126 875 11133 882
rect 11154 876 11178 886
rect 11235 882 11249 886
rect 11248 881 11251 882
rect 11248 878 11249 881
rect 11251 880 11252 881
rect 11178 875 11181 876
rect 10857 874 10859 875
rect 10918 874 11088 875
rect 10855 873 10857 874
rect 10916 873 10918 874
rect 10914 872 10916 873
rect 10919 872 11085 874
rect 11088 873 11096 874
rect 11096 872 11104 873
rect 11123 872 11126 875
rect 11181 874 11183 875
rect 11183 873 11186 874
rect 11186 872 11188 873
rect 11197 872 11209 878
rect 11252 875 11261 880
rect 11279 876 11281 886
rect 11370 882 11382 891
rect 11364 881 11370 882
rect 11336 880 11352 881
rect 11360 880 11364 881
rect 11429 880 11444 899
rect 11457 897 11463 903
rect 11494 901 11498 903
rect 11483 895 11494 901
rect 11507 899 11508 901
rect 11480 892 11483 895
rect 11479 891 11480 892
rect 11471 886 11479 891
rect 11308 875 11331 880
rect 11459 876 11491 886
rect 11504 880 11507 898
rect 11503 876 11504 880
rect 11539 878 11541 904
rect 11679 903 11680 922
rect 11694 915 11703 924
rect 11741 915 11750 924
rect 11685 906 11690 915
rect 11755 906 11759 915
rect 11660 881 11679 901
rect 10493 866 10499 868
rect 10588 867 10589 868
rect 10587 866 10588 867
rect 10492 865 10493 866
rect 10470 860 10492 865
rect 10546 862 10549 866
rect 10471 859 10492 860
rect 10543 859 10549 862
rect 10013 855 10022 857
rect 9938 850 9947 853
rect 9950 850 9956 853
rect 10001 852 10002 853
rect 10011 852 10022 855
rect 9958 851 10006 852
rect 10009 851 10011 852
rect 9958 850 10009 851
rect 10013 850 10022 852
rect 9948 847 9956 850
rect 9948 842 9952 847
rect 10001 840 10002 850
rect 10037 845 10041 858
rect 10080 846 10083 858
rect 10133 846 10137 858
rect 10153 851 10159 857
rect 10182 856 10186 859
rect 10476 858 10477 859
rect 10159 845 10165 851
rect 10177 845 10182 856
rect 10211 851 10217 857
rect 10284 855 10285 858
rect 10313 855 10314 858
rect 10543 857 10546 859
rect 10545 856 10546 857
rect 10541 855 10545 856
rect 10205 845 10211 851
rect 10219 847 10231 855
rect 10435 853 10436 855
rect 10282 851 10283 853
rect 10033 841 10037 845
rect 10079 841 10080 845
rect 10131 842 10133 845
rect 10031 840 10033 841
rect 10175 840 10177 845
rect 10279 841 10282 850
rect 10309 841 10312 850
rect 10436 841 10438 849
rect 10477 842 10478 849
rect 10538 847 10545 855
rect 10535 842 10538 847
rect 10541 845 10545 847
rect 10575 845 10587 865
rect 10699 859 10701 872
rect 10852 871 10854 872
rect 10912 871 10914 872
rect 10535 841 10537 842
rect 10532 840 10535 841
rect 10539 840 10541 845
rect 10572 844 10579 845
rect 10734 844 10738 870
rect 10847 868 10852 871
rect 10907 869 10911 871
rect 10995 869 11219 872
rect 11261 871 11267 875
rect 11298 871 11308 875
rect 11422 872 11425 876
rect 11456 875 11491 876
rect 11267 869 11273 871
rect 11280 869 11308 871
rect 10904 867 10906 868
rect 10844 866 10846 867
rect 10902 866 10904 867
rect 11011 866 11219 869
rect 11273 868 11274 869
rect 11280 868 11298 869
rect 11274 867 11278 868
rect 11293 867 11296 868
rect 10834 860 10844 866
rect 10892 862 10902 866
rect 11011 863 11221 866
rect 11124 862 11133 863
rect 11207 862 11229 863
rect 11250 862 11251 867
rect 11414 863 11422 872
rect 11469 869 11470 874
rect 11589 873 11600 874
rect 11617 873 11628 874
rect 11589 872 11597 873
rect 11621 872 11628 873
rect 11133 860 11136 862
rect 10829 857 10834 860
rect 10820 852 10829 857
rect 11136 852 11151 860
rect 11207 854 11221 862
rect 11229 856 11262 862
rect 11410 857 11414 862
rect 11337 856 11349 857
rect 11262 855 11268 856
rect 11286 855 11308 856
rect 11268 854 11308 855
rect 11329 854 11349 856
rect 10818 851 10820 852
rect 11151 851 11153 852
rect 10815 850 10818 851
rect 11153 850 11155 851
rect 10780 849 10786 850
rect 10813 849 10815 850
rect 10762 844 10813 849
rect 10826 844 10832 850
rect 10876 845 10879 849
rect 11156 845 11164 849
rect 11207 846 11219 854
rect 11337 851 11369 854
rect 11338 847 11369 851
rect 11407 849 11409 856
rect 11407 847 11408 849
rect 10572 840 10576 844
rect 9953 836 9954 840
rect 9954 833 9955 836
rect 10001 832 10003 840
rect 10019 832 10031 840
rect 10078 838 10079 840
rect 10130 838 10131 840
rect 10077 832 10078 838
rect 10129 833 10130 838
rect 10172 832 10175 840
rect 10278 837 10279 840
rect 10277 833 10278 836
rect 10306 834 10308 840
rect 10478 837 10479 840
rect 10439 832 10443 837
rect 10530 832 10539 840
rect 10568 834 10576 840
rect 10568 832 10572 834
rect 9955 817 9963 832
rect 10001 825 10005 832
rect 10018 830 10019 832
rect 10171 830 10172 832
rect 10017 828 10018 830
rect 10076 828 10077 830
rect 10127 828 10128 830
rect 10016 825 10017 828
rect 10003 817 10005 825
rect 10075 824 10076 828
rect 10126 824 10127 827
rect 10169 824 10171 829
rect 10014 819 10016 824
rect 10074 819 10075 824
rect 10121 820 10126 824
rect 8373 805 8381 808
rect 8373 804 8375 805
rect 8376 800 8377 802
rect 8377 797 8379 800
rect 8134 790 8136 793
rect 7942 758 7958 763
rect 8007 773 8068 785
rect 8075 779 8088 790
rect 8074 774 8088 779
rect 8118 777 8136 790
rect 8227 789 8228 793
rect 8258 789 8259 795
rect 8118 774 8134 777
rect 8007 759 8072 773
rect 8038 758 8054 759
rect 8056 758 8072 759
rect 8099 758 8100 760
rect 8134 758 8150 774
rect 8228 767 8232 785
rect 8259 779 8260 788
rect 8308 787 8310 794
rect 8373 790 8374 794
rect 8379 791 8382 797
rect 8414 792 8430 808
rect 8464 802 8492 808
rect 8528 806 8548 816
rect 9963 809 9967 817
rect 10005 811 10006 817
rect 10013 815 10014 819
rect 10073 815 10074 819
rect 10121 815 10125 820
rect 10167 819 10169 824
rect 10012 809 10013 814
rect 10071 809 10073 814
rect 10121 809 10123 815
rect 10164 814 10167 818
rect 10217 814 10233 824
rect 10235 814 10251 824
rect 10271 817 10277 832
rect 10160 809 10164 814
rect 10204 809 10211 814
rect 10256 808 10264 814
rect 10269 811 10271 817
rect 10299 811 10306 832
rect 10440 827 10444 832
rect 10479 827 10485 832
rect 10528 830 10530 832
rect 10567 830 10568 832
rect 10298 809 10299 811
rect 10313 808 10329 824
rect 10429 822 10495 827
rect 10521 824 10528 830
rect 10564 825 10567 830
rect 10570 828 10572 832
rect 10701 832 10703 844
rect 10713 840 10725 844
rect 10741 842 10762 844
rect 10732 841 10741 842
rect 10727 840 10734 841
rect 10713 836 10727 840
rect 10429 821 10485 822
rect 10420 814 10429 821
rect 10440 818 10444 821
rect 10418 811 10420 814
rect 10443 811 10444 817
rect 10479 811 10485 821
rect 10495 814 10499 821
rect 10513 819 10521 824
rect 10561 819 10564 824
rect 10513 818 10515 819
rect 10513 815 10514 818
rect 10559 817 10561 819
rect 10558 816 10559 817
rect 10499 811 10500 814
rect 10512 812 10513 813
rect 10558 812 10561 816
rect 10591 812 10603 815
rect 10501 811 10510 812
rect 10336 808 10355 809
rect 10361 808 10363 809
rect 9968 804 9969 807
rect 8458 794 8492 802
rect 9969 799 9971 803
rect 10006 799 10007 803
rect 10009 800 10012 808
rect 10069 800 10071 808
rect 9971 794 9973 798
rect 10009 794 10011 800
rect 10067 794 10069 798
rect 8454 791 8456 794
rect 8464 790 8492 794
rect 8310 781 8311 787
rect 8373 782 8390 790
rect 8260 766 8265 779
rect 8312 774 8320 780
rect 8374 776 8390 782
rect 8446 779 8454 790
rect 8443 778 8454 779
rect 8458 788 8492 790
rect 8374 774 8384 776
rect 8320 773 8322 774
rect 8232 760 8233 766
rect 8265 759 8267 766
rect 8322 765 8336 773
rect 8374 766 8375 774
rect 8390 768 8395 776
rect 8443 770 8452 778
rect 8371 765 8375 766
rect 8317 764 8350 765
rect 8371 764 8381 765
rect 8317 759 8323 764
rect 7867 756 7873 758
rect 7944 757 7958 758
rect 8070 757 8073 758
rect 7952 756 8005 757
rect 7785 754 7786 756
rect 7867 754 7876 756
rect 7549 738 7555 739
rect 7595 738 7601 744
rect 7635 738 7644 747
rect 7682 738 7691 747
rect 7774 746 7788 754
rect 7862 747 7876 754
rect 7947 750 8011 756
rect 8074 750 8089 756
rect 8096 754 8097 756
rect 8138 752 8139 753
rect 7862 746 7867 747
rect 7788 745 7791 746
rect 7301 734 7302 736
rect 7303 727 7306 733
rect 7375 731 7390 736
rect 7543 732 7549 738
rect 7601 733 7607 738
rect 7655 734 7667 738
rect 7708 734 7724 744
rect 7786 742 7787 745
rect 7791 742 7830 745
rect 7860 743 7867 746
rect 7953 745 7968 750
rect 7999 747 8008 750
rect 7953 744 7959 745
rect 7999 744 8005 747
rect 7787 740 7830 742
rect 7791 737 7830 740
rect 7853 739 7860 743
rect 7862 739 7867 743
rect 8008 742 8022 747
rect 8089 745 8102 750
rect 8138 747 8146 752
rect 8234 751 8235 756
rect 8268 750 8271 756
rect 8323 753 8329 759
rect 8334 758 8350 764
rect 8352 758 8368 764
rect 8375 759 8381 764
rect 8395 762 8398 768
rect 8434 761 8443 770
rect 8369 753 8375 759
rect 8400 756 8402 760
rect 8430 757 8431 758
rect 8088 742 8090 745
rect 8102 742 8108 745
rect 8139 744 8146 747
rect 8235 746 8236 750
rect 8271 744 8273 750
rect 8357 745 8360 747
rect 8148 742 8149 744
rect 8402 743 8410 756
rect 8431 754 8434 757
rect 8446 756 8454 768
rect 8458 758 8460 788
rect 8489 787 8492 788
rect 8496 779 8539 791
rect 9974 785 9977 793
rect 10008 790 10010 793
rect 10011 790 10025 794
rect 10008 786 10025 790
rect 8490 776 8539 779
rect 8490 770 8499 776
rect 8510 774 8526 776
rect 8539 774 8560 776
rect 9977 775 9982 785
rect 8499 764 8508 770
rect 8502 763 8508 764
rect 8526 768 8560 774
rect 9982 771 9983 775
rect 10009 774 10025 786
rect 10059 790 10067 794
rect 10105 792 10121 808
rect 10155 801 10160 808
rect 10200 801 10204 808
rect 10256 807 10267 808
rect 10297 807 10313 808
rect 10363 807 10364 808
rect 10412 807 10418 810
rect 10485 809 10486 811
rect 10440 808 10442 809
rect 10500 808 10510 811
rect 10557 808 10558 812
rect 10591 808 10607 812
rect 10609 808 10625 824
rect 10627 808 10643 824
rect 10701 820 10709 832
rect 10713 831 10729 832
rect 10713 830 10723 831
rect 10645 808 10654 812
rect 10704 810 10705 811
rect 10429 807 10439 808
rect 10256 806 10268 807
rect 10263 804 10268 806
rect 10155 792 10158 801
rect 10059 774 10075 790
rect 10105 774 10121 790
rect 10155 787 10171 790
rect 10150 781 10171 787
rect 10191 787 10200 801
rect 10263 792 10267 804
rect 10296 803 10313 807
rect 10364 806 10367 807
rect 10295 799 10296 803
rect 10293 794 10295 798
rect 10297 792 10313 803
rect 10336 798 10348 806
rect 10367 803 10370 806
rect 10390 803 10429 807
rect 10486 803 10487 807
rect 10497 803 10512 808
rect 10591 807 10608 808
rect 10613 807 10625 808
rect 10351 799 10390 803
rect 10401 799 10407 803
rect 10412 799 10418 803
rect 10487 799 10488 803
rect 10191 785 10202 787
rect 10211 785 10223 791
rect 10263 785 10264 792
rect 10291 788 10293 792
rect 10180 783 10202 785
rect 10212 783 10223 785
rect 10262 783 10267 785
rect 10174 781 10179 783
rect 10144 775 10150 781
rect 10155 774 10171 781
rect 10189 779 10191 783
rect 10196 781 10202 783
rect 10223 781 10227 783
rect 10202 775 10208 781
rect 10211 778 10223 779
rect 10011 771 10015 774
rect 8503 759 8506 763
rect 8526 758 8542 768
rect 8560 762 8577 768
rect 8563 758 8569 762
rect 8577 760 8583 762
rect 8583 758 8587 760
rect 8609 758 8615 764
rect 8458 757 8473 758
rect 8458 756 8477 757
rect 8434 750 8439 754
rect 8474 752 8492 756
rect 8509 753 8515 756
rect 8557 753 8563 758
rect 8458 750 8492 752
rect 8515 751 8563 753
rect 8615 752 8621 758
rect 9983 754 9991 771
rect 10015 754 10022 771
rect 10025 758 10041 774
rect 10043 758 10059 774
rect 10121 772 10129 774
rect 10147 772 10155 774
rect 10221 772 10223 778
rect 10227 772 10235 779
rect 10260 778 10262 783
rect 10263 778 10267 783
rect 10260 774 10267 778
rect 10260 772 10262 774
rect 10121 758 10137 772
rect 10139 758 10155 772
rect 10202 757 10265 772
rect 10289 760 10291 786
rect 10297 774 10313 790
rect 10324 782 10332 794
rect 10336 793 10357 794
rect 10395 793 10401 799
rect 10336 792 10354 793
rect 10313 763 10317 767
rect 10324 763 10332 772
rect 10336 763 10338 792
rect 10489 788 10491 796
rect 10497 794 10519 803
rect 10497 792 10512 794
rect 10549 790 10557 806
rect 10587 804 10589 807
rect 10593 806 10607 807
rect 10591 803 10607 806
rect 10643 805 10659 808
rect 10641 803 10659 805
rect 10579 791 10587 803
rect 10589 801 10625 803
rect 10589 793 10609 801
rect 10622 800 10625 801
rect 10623 793 10625 800
rect 10629 799 10637 803
rect 10641 799 10663 803
rect 10643 794 10663 799
rect 10701 798 10709 810
rect 10713 800 10715 830
rect 10732 826 10734 840
rect 10774 838 10780 844
rect 10832 838 10838 844
rect 10871 841 10876 845
rect 11164 841 11169 845
rect 11163 832 11171 841
rect 11175 834 11177 839
rect 11207 834 11209 846
rect 11467 845 11469 865
rect 11501 863 11503 872
rect 11538 863 11539 872
rect 11589 871 11591 872
rect 11627 871 11628 872
rect 11660 868 11674 881
rect 11653 866 11666 868
rect 11653 865 11665 866
rect 11694 865 11699 866
rect 11500 857 11501 862
rect 11498 849 11499 855
rect 11219 844 11222 845
rect 11175 832 11209 834
rect 11213 840 11222 844
rect 11213 832 11221 840
rect 11222 832 11226 840
rect 11226 830 11227 832
rect 10747 826 10748 830
rect 10858 829 10861 830
rect 10834 827 10869 829
rect 10732 818 10733 826
rect 10830 825 10834 827
rect 10828 824 10830 825
rect 10748 812 10750 824
rect 10733 800 10736 811
rect 10801 808 10828 824
rect 10832 812 10836 817
rect 10842 812 10858 827
rect 10869 824 10894 827
rect 10837 811 10858 812
rect 10713 798 10747 800
rect 10733 795 10736 798
rect 10491 778 10494 788
rect 10494 769 10496 778
rect 10497 774 10512 790
rect 10549 774 10563 790
rect 10586 781 10587 788
rect 10496 765 10497 769
rect 10313 762 10338 763
rect 10367 762 10370 763
rect 10313 760 10370 762
rect 10313 758 10329 760
rect 10497 759 10498 763
rect 8439 749 8475 750
rect 8458 744 8470 749
rect 8525 744 8536 749
rect 9991 746 9994 754
rect 10022 748 10027 754
rect 10027 745 10031 748
rect 10221 745 10223 757
rect 10226 745 10260 757
rect 10265 756 10267 757
rect 10374 756 10401 759
rect 10498 757 10499 759
rect 10513 758 10529 772
rect 10531 758 10547 772
rect 10579 769 10587 781
rect 10591 774 10609 793
rect 10643 792 10659 794
rect 10643 774 10659 790
rect 10689 774 10704 790
rect 10706 775 10708 792
rect 10713 786 10725 794
rect 10735 786 10747 794
rect 10749 790 10750 808
rect 10836 805 10846 811
rect 10894 808 11035 824
rect 11097 808 11113 824
rect 11115 808 11131 824
rect 11175 820 11187 828
rect 11197 820 11209 828
rect 11227 826 11228 830
rect 11253 828 11255 845
rect 11175 810 11177 820
rect 11228 816 11231 824
rect 11255 819 11256 828
rect 11283 819 11286 845
rect 11325 833 11331 845
rect 11372 843 11374 844
rect 11497 843 11498 847
rect 11408 838 11409 843
rect 11375 827 11376 836
rect 11409 827 11410 836
rect 11465 825 11467 840
rect 11496 837 11497 843
rect 11494 827 11496 836
rect 11536 829 11538 862
rect 11649 855 11665 865
rect 11702 864 11706 868
rect 11586 845 11649 855
rect 11694 851 11702 864
rect 11577 844 11586 845
rect 11571 842 11577 844
rect 11569 840 11571 842
rect 11325 811 11331 823
rect 11493 821 11494 826
rect 11534 820 11536 827
rect 11550 825 11569 840
rect 11549 824 11550 825
rect 11377 817 11378 820
rect 11410 816 11411 820
rect 11378 811 11383 816
rect 11411 811 11412 816
rect 11464 811 11465 818
rect 11478 811 11484 817
rect 11492 816 11493 820
rect 11533 818 11534 820
rect 11541 818 11549 824
rect 11490 812 11492 816
rect 11524 811 11530 817
rect 11532 816 11541 818
rect 11531 811 11541 816
rect 11287 808 11288 810
rect 11379 808 11380 810
rect 10841 803 10846 805
rect 10966 803 10975 808
rect 11013 803 11022 808
rect 10753 802 10762 803
rect 10751 798 10759 802
rect 10762 799 10777 802
rect 10777 798 10780 799
rect 10774 792 10780 798
rect 10832 792 10838 798
rect 10846 794 10855 803
rect 10957 794 10966 803
rect 11022 794 11031 803
rect 10948 792 10955 793
rect 10780 790 10786 792
rect 10591 772 10625 774
rect 10638 772 10643 774
rect 10736 772 10739 786
rect 10749 774 10755 790
rect 10780 786 10801 790
rect 10826 786 10832 792
rect 10942 791 10948 792
rect 10999 791 11003 793
rect 11035 792 11051 808
rect 11081 792 11097 808
rect 11108 803 11114 808
rect 11108 802 11123 803
rect 11102 796 11108 802
rect 11131 798 11147 808
rect 11154 802 11160 808
rect 11107 791 11108 793
rect 11140 791 11145 798
rect 11160 796 11166 802
rect 11178 800 11179 808
rect 10940 790 10942 791
rect 10939 787 10940 790
rect 11004 789 11006 790
rect 10785 774 10801 786
rect 10852 778 10879 781
rect 10835 774 10852 778
rect 10879 774 10887 778
rect 10591 769 10643 772
rect 10704 769 10710 772
rect 10739 771 10743 772
rect 10591 757 10595 765
rect 10627 758 10643 769
rect 10705 762 10722 769
rect 10739 762 10749 771
rect 10705 758 10721 762
rect 10722 760 10727 762
rect 10731 760 10743 762
rect 10727 759 10743 760
rect 10723 758 10743 759
rect 10801 758 10817 774
rect 10887 772 10890 774
rect 10955 772 10961 778
rect 10964 772 10966 779
rect 11006 772 11007 778
rect 11035 774 11051 790
rect 11081 774 11097 790
rect 11099 779 11108 791
rect 10890 763 10910 772
rect 10939 767 10940 769
rect 10949 766 10955 772
rect 11007 766 11013 772
rect 11028 763 11035 774
rect 10910 762 10912 763
rect 10912 759 10918 762
rect 10267 751 10288 756
rect 10288 747 10304 751
rect 10336 748 10348 756
rect 10499 754 10500 756
rect 10395 747 10401 753
rect 10426 747 10481 753
rect 10500 750 10501 754
rect 10501 747 10503 748
rect 10510 747 10519 756
rect 10589 747 10595 756
rect 10647 747 10653 753
rect 10654 747 10663 756
rect 10708 751 10711 758
rect 8536 743 8538 744
rect 8022 739 8031 742
rect 8108 741 8110 742
rect 8410 741 8411 743
rect 9994 741 9996 745
rect 7853 738 7867 739
rect 7840 737 7853 738
rect 7860 735 7862 738
rect 8031 735 8042 739
rect 8085 737 8086 739
rect 8042 734 8045 735
rect 7651 733 7733 734
rect 7601 732 7667 733
rect 7644 731 7667 732
rect 7390 726 7402 731
rect 7644 729 7651 731
rect 7655 730 7667 731
rect 7733 729 7736 732
rect 7852 731 7859 734
rect 8045 731 8054 734
rect 8082 733 8084 736
rect 8054 729 8061 731
rect 8077 729 8081 731
rect 7640 728 7644 729
rect 7633 726 7640 728
rect 7670 727 7671 729
rect 7736 728 7738 729
rect 7092 721 7163 723
rect 6916 719 6931 720
rect 7093 719 7163 721
rect 7195 719 7199 725
rect 7306 723 7308 726
rect 6919 716 6931 719
rect 5243 706 5253 709
rect 5254 706 5266 715
rect 5289 714 5291 715
rect 5291 709 5331 714
rect 5353 709 5365 714
rect 6855 712 6860 716
rect 6932 714 6935 716
rect 7084 712 7092 719
rect 7094 717 7104 719
rect 7094 712 7098 717
rect 5331 707 5365 709
rect 5331 706 5379 707
rect 5401 706 5407 712
rect 5459 706 5465 712
rect 4828 698 4839 701
rect 4922 698 4930 701
rect 4950 700 4958 701
rect 4291 688 4292 692
rect 4254 676 4288 678
rect 4292 676 4300 688
rect 4387 686 4393 692
rect 4445 686 4451 692
rect 4477 688 4484 692
rect 4593 691 4599 697
rect 4639 691 4645 697
rect 4685 691 4828 698
rect 4900 691 4922 698
rect 4956 692 4958 700
rect 4959 693 4965 698
rect 4978 694 4990 701
rect 4580 688 4582 691
rect 4477 687 4489 688
rect 4393 680 4399 686
rect 4439 680 4445 686
rect 4477 685 4492 687
rect 4499 685 4511 688
rect 4579 687 4580 688
rect 4578 685 4579 687
rect 4587 685 4593 691
rect 4645 685 4651 691
rect 4652 689 4673 691
rect 4895 689 4900 691
rect 4889 687 4895 689
rect 4958 688 4959 692
rect 4967 689 4970 691
rect 4656 685 4691 687
rect 4477 680 4489 685
rect 4492 680 4514 685
rect 4576 683 4578 685
rect 4514 676 4527 680
rect 4527 675 4532 676
rect 4541 675 4591 683
rect 4644 682 4656 685
rect 4635 680 4644 682
rect 4696 680 4698 685
rect 4879 684 4887 687
rect 4959 686 4960 687
rect 4872 682 4879 684
rect 4634 676 4635 680
rect 4865 679 4872 682
rect 4960 680 4962 682
rect 4860 678 4865 679
rect 4854 676 4860 678
rect 4962 676 4964 680
rect 4976 678 4983 684
rect 4995 682 5053 701
rect 5080 692 5081 698
rect 5144 692 5145 701
rect 5149 693 5157 703
rect 5164 702 5168 705
rect 5229 702 5254 706
rect 5351 704 5364 706
rect 5152 691 5157 693
rect 5168 692 5179 702
rect 4995 678 5028 682
rect 4290 672 4292 675
rect 4532 674 4591 675
rect 4541 672 4591 674
rect 3997 656 4000 662
rect 3921 643 3985 649
rect 3995 648 3997 656
rect 4041 652 4058 672
rect 4081 666 4088 672
rect 4254 666 4266 672
rect 4276 666 4288 672
rect 4518 666 4541 672
rect 4088 664 4294 666
rect 4507 664 4518 666
rect 3927 637 3954 643
rect 3973 637 3979 643
rect 3989 642 3995 647
rect 3999 642 4008 644
rect 4058 643 4066 652
rect 4235 642 4236 660
rect 3737 626 3740 630
rect 3930 626 3954 637
rect 3989 635 4008 642
rect 4067 639 4071 642
rect 4071 636 4076 639
rect 4076 635 4084 636
rect 3989 630 4004 635
rect 4084 631 4120 635
rect 3988 626 4004 630
rect 4120 628 4140 631
rect 4234 630 4236 642
rect 4294 654 4453 664
rect 4465 654 4507 664
rect 4631 663 4634 674
rect 4698 663 4701 676
rect 4849 674 4854 676
rect 4846 673 4849 674
rect 4841 672 4846 673
rect 4835 670 4841 672
rect 4964 670 4967 676
rect 4983 671 4991 678
rect 5028 671 5036 678
rect 5053 676 5059 682
rect 5082 679 5083 682
rect 5084 677 5085 687
rect 5136 681 5149 682
rect 5136 679 5145 681
rect 5179 679 5184 692
rect 5229 688 5278 702
rect 5303 698 5349 704
rect 5367 703 5369 706
rect 5379 704 5399 706
rect 5407 704 5426 706
rect 5350 700 5365 702
rect 5295 694 5303 698
rect 5229 687 5254 688
rect 5278 687 5284 688
rect 5286 687 5295 694
rect 5211 678 5229 687
rect 5278 686 5286 687
rect 5284 685 5288 686
rect 5274 677 5281 683
rect 5288 682 5296 685
rect 5296 681 5301 682
rect 5301 680 5306 681
rect 5307 678 5310 679
rect 5078 676 5099 677
rect 5136 676 5142 677
rect 5059 673 5063 676
rect 4816 668 4835 670
rect 4779 664 4816 668
rect 4702 663 4779 664
rect 4593 655 4779 663
rect 4967 660 4980 670
rect 4991 660 5013 671
rect 5036 663 5046 671
rect 5063 663 5067 673
rect 5078 671 5084 676
rect 5085 672 5099 676
rect 5125 671 5142 676
rect 5183 671 5184 676
rect 5194 671 5209 677
rect 5084 665 5090 671
rect 5130 665 5136 671
rect 5174 663 5194 671
rect 5265 669 5274 677
rect 5313 676 5318 678
rect 5319 674 5325 676
rect 4294 652 4465 654
rect 4593 653 4708 655
rect 4294 642 4296 652
rect 4593 651 4705 653
rect 4593 649 4698 651
rect 4593 648 4661 649
rect 4593 645 4645 648
rect 4587 644 4651 645
rect 4565 643 4651 644
rect 4565 642 4583 643
rect 4294 634 4300 642
rect 4559 639 4576 642
rect 4587 639 4651 643
rect 4684 641 4696 649
rect 4701 643 4705 651
rect 4541 636 4559 639
rect 4295 630 4300 634
rect 4522 633 4541 636
rect 4593 633 4599 639
rect 4625 636 4631 639
rect 4639 633 4645 639
rect 4703 636 4705 643
rect 4980 642 5026 660
rect 5046 652 5076 663
rect 5056 647 5090 652
rect 5110 647 5111 660
rect 5147 652 5174 663
rect 5183 660 5184 663
rect 5056 646 5127 647
rect 5135 646 5164 652
rect 5056 643 5164 646
rect 5062 642 5067 643
rect 4980 641 5028 642
rect 4507 631 4522 633
rect 4311 630 4351 631
rect 4505 630 4507 631
rect 4150 628 4311 630
rect 4351 628 4380 630
rect 4234 626 4237 628
rect 4293 626 4300 628
rect 3740 618 3748 626
rect 3808 618 3815 625
rect 3748 617 3808 618
rect 3972 610 3988 626
rect 4237 615 4243 626
rect 4290 618 4293 625
rect 4380 622 4441 628
rect 4451 622 4501 630
rect 4701 627 4703 636
rect 4282 615 4290 618
rect 4243 613 4284 615
rect 4625 613 4638 624
rect 4679 616 4701 627
rect 4980 626 5026 641
rect 5030 637 5033 639
rect 5033 636 5035 637
rect 5035 633 5042 636
rect 5062 634 5076 642
rect 5110 634 5111 643
rect 5182 637 5183 653
rect 5224 652 5265 669
rect 5319 668 5327 674
rect 5331 670 5333 672
rect 5363 670 5365 700
rect 5369 690 5377 702
rect 5407 700 5413 704
rect 5453 700 5459 706
rect 5477 693 5488 702
rect 6860 696 6881 712
rect 6925 710 6949 712
rect 6929 705 6949 710
rect 7084 707 7094 712
rect 7091 705 7094 707
rect 6881 695 6883 696
rect 5331 668 5365 670
rect 5369 668 5377 680
rect 5488 678 5491 692
rect 6887 689 6888 692
rect 6885 678 6892 687
rect 6929 680 6931 705
rect 6935 700 6943 705
rect 6949 699 6955 705
rect 7089 701 7091 705
rect 7083 699 7091 701
rect 6955 694 6961 699
rect 7083 695 7089 699
rect 6961 692 6964 694
rect 6897 678 6931 680
rect 6935 678 6943 690
rect 6964 688 6965 692
rect 7077 689 7083 695
rect 7087 692 7088 694
rect 7086 688 7087 691
rect 7096 689 7098 712
rect 7128 715 7183 719
rect 7128 701 7151 715
rect 7159 713 7183 715
rect 7203 713 7204 715
rect 7164 708 7183 713
rect 7204 708 7208 713
rect 7308 710 7315 723
rect 7402 722 7432 726
rect 7651 724 7667 726
rect 7402 714 7444 722
rect 7171 701 7183 708
rect 7208 706 7209 708
rect 7315 705 7318 710
rect 7396 709 7445 710
rect 7128 695 7135 701
rect 7128 693 7141 695
rect 7128 689 7130 693
rect 7135 689 7141 693
rect 7146 691 7155 700
rect 7174 696 7183 701
rect 7214 696 7217 701
rect 7177 691 7183 696
rect 7085 685 7086 687
rect 7129 685 7130 689
rect 7147 687 7164 691
rect 7180 689 7183 691
rect 7217 689 7223 696
rect 7318 695 7355 705
rect 7396 702 7410 709
rect 7426 708 7445 709
rect 7442 703 7445 708
rect 7395 699 7396 701
rect 7355 693 7361 695
rect 7393 694 7395 699
rect 7361 692 7366 693
rect 7392 692 7393 694
rect 7182 687 7183 689
rect 7148 686 7164 687
rect 7223 686 7225 689
rect 7366 688 7382 692
rect 7382 687 7384 688
rect 6965 680 6967 685
rect 7084 680 7085 685
rect 7150 682 7153 686
rect 7155 682 7164 686
rect 7156 680 7157 682
rect 5491 676 5492 678
rect 6892 676 6893 678
rect 6896 676 6897 678
rect 7083 676 7084 678
rect 7157 677 7158 680
rect 5327 664 5330 666
rect 5331 656 5343 664
rect 5353 656 5365 664
rect 5492 661 5495 676
rect 5209 646 5224 652
rect 5331 648 5340 656
rect 5494 648 5495 661
rect 6892 660 6896 676
rect 6932 674 6935 676
rect 6897 666 6909 674
rect 6919 666 6931 674
rect 6967 660 6971 676
rect 6891 654 6892 658
rect 6971 657 6972 660
rect 5200 643 5207 646
rect 5195 641 5200 643
rect 5186 637 5195 641
rect 5042 631 5048 633
rect 5060 630 5076 634
rect 5051 626 5076 630
rect 5110 626 5112 630
rect 5044 622 5069 626
rect 4639 613 4679 616
rect 4250 610 4266 613
rect 4268 610 4284 613
rect 5044 610 5060 622
rect 5069 619 5077 622
rect 5077 618 5086 619
rect 5112 615 5117 626
rect 5144 620 5186 637
rect 5141 619 5144 620
rect 5135 618 5141 619
rect 5173 618 5180 620
rect 5169 615 5173 618
rect 5117 611 5138 615
rect 5160 611 5169 615
rect 5310 606 5334 629
rect 5340 626 5379 648
rect 5379 621 5388 626
rect 5485 622 5494 643
rect 6891 630 6893 654
rect 6971 630 6972 654
rect 7083 649 7135 663
rect 7156 662 7158 675
rect 7185 672 7197 685
rect 7225 672 7237 686
rect 7387 685 7393 687
rect 7393 683 7401 685
rect 7398 681 7402 683
rect 7398 676 7405 681
rect 7442 678 7444 703
rect 7445 697 7446 702
rect 7448 698 7456 710
rect 7601 694 7629 695
rect 7665 694 7667 724
rect 7671 714 7679 726
rect 7738 712 7740 728
rect 8061 727 8067 729
rect 8074 727 8077 729
rect 7794 720 7800 726
rect 7852 720 7858 726
rect 8058 723 8078 727
rect 8110 723 8131 741
rect 8136 738 8147 740
rect 8058 721 8074 723
rect 8053 720 8058 721
rect 8078 720 8086 723
rect 7800 714 7806 720
rect 7846 714 7852 720
rect 8046 717 8053 720
rect 8086 719 8089 720
rect 8131 719 8136 723
rect 8041 716 8046 717
rect 8089 716 8095 719
rect 8136 716 8140 719
rect 8144 716 8146 738
rect 8147 737 8148 738
rect 8150 737 8158 740
rect 8148 734 8158 737
rect 8150 729 8158 734
rect 8237 733 8238 741
rect 8274 737 8277 741
rect 8238 729 8239 733
rect 8267 729 8279 737
rect 8289 729 8301 737
rect 8364 729 8377 741
rect 8150 728 8159 729
rect 8155 726 8159 728
rect 8150 716 8158 718
rect 8032 713 8041 716
rect 8027 711 8032 713
rect 7446 693 7447 694
rect 7621 692 7629 694
rect 7633 692 7667 694
rect 7671 692 7679 704
rect 7738 694 7740 710
rect 8011 706 8027 711
rect 8095 706 8106 716
rect 8140 707 8158 716
rect 8122 706 8158 707
rect 8159 706 8182 726
rect 8239 724 8246 729
rect 8263 727 8266 729
rect 8279 725 8280 729
rect 8286 725 8292 729
rect 8240 723 8246 724
rect 8255 723 8263 725
rect 8267 723 8313 725
rect 8234 717 8240 723
rect 8267 717 8269 723
rect 8292 717 8298 723
rect 8299 717 8313 723
rect 8238 713 8240 714
rect 8236 709 8238 713
rect 7995 701 8011 706
rect 8106 705 8113 706
rect 8151 705 8184 706
rect 8106 702 8114 705
rect 8088 701 8122 702
rect 8148 701 8209 705
rect 8299 702 8301 717
rect 8305 713 8320 717
rect 8308 705 8320 713
rect 8377 712 8396 729
rect 8411 715 8445 741
rect 8540 723 8563 741
rect 10031 740 10039 745
rect 10257 742 10258 745
rect 10304 742 10324 747
rect 10324 741 10329 742
rect 10401 741 10407 747
rect 10447 741 10453 747
rect 10223 740 10225 741
rect 9996 737 9998 740
rect 10039 737 10044 740
rect 10213 739 10223 740
rect 10202 738 10223 739
rect 10329 738 10333 741
rect 10454 738 10463 747
rect 10501 745 10510 747
rect 10501 742 10516 745
rect 10501 738 10510 742
rect 10516 740 10520 742
rect 10595 741 10607 747
rect 10641 741 10654 747
rect 10710 744 10711 751
rect 10520 739 10523 740
rect 10044 736 10046 737
rect 10211 736 10230 738
rect 9999 733 10000 736
rect 10046 733 10050 736
rect 10000 727 10003 733
rect 10050 731 10054 733
rect 10054 729 10057 731
rect 10144 729 10150 735
rect 10202 729 10208 735
rect 10211 733 10248 736
rect 10255 733 10256 736
rect 10222 729 10248 733
rect 10251 729 10255 731
rect 10287 729 10288 730
rect 10057 726 10061 729
rect 10003 720 10007 726
rect 10061 720 10071 726
rect 10074 720 10086 724
rect 10150 723 10156 729
rect 10196 723 10202 729
rect 10248 726 10288 729
rect 10248 723 10287 726
rect 10333 725 10350 738
rect 10454 737 10455 738
rect 10523 736 10530 739
rect 10598 738 10607 741
rect 10645 738 10654 741
rect 10704 739 10711 744
rect 10739 742 10743 758
rect 10781 747 10790 756
rect 10846 747 10855 756
rect 10918 754 10929 759
rect 11022 758 11035 763
rect 11097 769 11106 774
rect 11107 769 11108 779
rect 11097 763 11108 769
rect 11111 763 11113 791
rect 11179 790 11181 791
rect 11177 785 11181 790
rect 11230 790 11231 808
rect 11337 799 11349 803
rect 11359 799 11371 803
rect 11381 796 11382 799
rect 11412 796 11413 805
rect 11463 799 11464 808
rect 11472 805 11478 811
rect 11530 808 11536 811
rect 11585 808 11601 824
rect 12174 819 12175 1015
rect 12364 819 12365 1015
rect 12450 819 12451 1015
rect 12723 819 12724 1015
rect 12921 820 12922 1016
rect 13313 1014 13317 1019
rect 13951 1014 13958 1019
rect 14038 1018 14047 1027
rect 14103 1024 14199 1027
rect 14540 1023 14648 1037
rect 14398 1015 14414 1022
rect 14416 1015 14432 1022
rect 13958 1007 13970 1014
rect 14388 1013 14400 1015
rect 14410 1013 14422 1015
rect 14428 1013 14432 1015
rect 14616 1013 14632 1022
rect 14648 1021 14666 1023
rect 14667 1017 14674 1020
rect 14674 1013 14680 1017
rect 15320 1015 15321 1026
rect 15510 1015 15511 1026
rect 15596 1015 15597 1026
rect 15869 1015 15870 1026
rect 16067 1016 16068 1027
rect 16495 1023 16596 1034
rect 16782 1033 17046 1034
rect 17046 1023 17101 1033
rect 17204 1027 17213 1036
rect 17251 1027 17260 1036
rect 17554 1034 17676 1037
rect 17526 1033 17543 1034
rect 17356 1027 17526 1033
rect 16480 1021 16495 1023
rect 16474 1019 16480 1021
rect 17103 1019 17108 1021
rect 14388 1008 14432 1013
rect 14575 1008 14612 1009
rect 14680 1008 14683 1013
rect 14384 1006 14386 1008
rect 14388 1006 14520 1008
rect 13439 1005 13793 1006
rect 13419 1003 13437 1005
rect 13879 1003 13892 1005
rect 13971 1003 13974 1005
rect 14382 1003 14520 1006
rect 13363 1000 13419 1003
rect 13237 992 13249 1000
rect 13259 992 13271 1000
rect 13335 994 13419 1000
rect 13892 994 13902 1003
rect 13335 993 13363 994
rect 13233 989 13235 992
rect 13335 991 13354 993
rect 13903 991 13906 993
rect 13275 988 13279 989
rect 13225 977 13233 988
rect 13236 986 13271 988
rect 13234 977 13236 983
rect 13225 976 13234 977
rect 13233 972 13234 976
rect 13232 971 13233 972
rect 13230 966 13232 969
rect 13105 964 13170 965
rect 13097 956 13105 964
rect 13170 956 13174 964
rect 13096 950 13097 956
rect 13225 954 13233 966
rect 13237 956 13239 986
rect 13268 985 13271 986
rect 13270 979 13271 985
rect 13275 981 13283 988
rect 13279 980 13287 981
rect 13311 980 13312 990
rect 13335 980 13350 991
rect 13609 981 13646 983
rect 13287 979 13293 980
rect 13310 979 13311 980
rect 13335 979 13342 980
rect 13293 969 13355 979
rect 13363 972 13369 978
rect 13409 972 13415 978
rect 13609 977 13635 981
rect 13646 977 13651 981
rect 13906 980 13919 991
rect 13882 979 13896 980
rect 13603 972 13609 977
rect 13651 972 13660 977
rect 13864 972 13882 979
rect 13896 977 13903 979
rect 13974 977 13995 1003
rect 14376 996 14520 1003
rect 14536 1006 14637 1008
rect 14536 996 14648 1006
rect 14337 990 14398 996
rect 14302 987 14337 990
rect 14115 981 14302 987
rect 14388 986 14398 990
rect 13903 972 13918 977
rect 13357 969 13363 972
rect 13364 970 13421 972
rect 13660 971 13661 972
rect 13498 970 13501 971
rect 13519 970 13522 971
rect 13601 970 13602 971
rect 13661 970 13664 971
rect 13364 969 13372 970
rect 13335 968 13372 969
rect 13237 954 13271 956
rect 13226 951 13228 954
rect 13222 939 13226 950
rect 13237 942 13249 950
rect 13262 945 13271 954
rect 13309 952 13310 955
rect 13335 951 13340 968
rect 13357 966 13372 968
rect 13415 966 13421 970
rect 13494 967 13498 970
rect 13522 967 13527 970
rect 13664 968 13665 970
rect 13856 969 13864 972
rect 13893 971 13918 972
rect 13927 971 13931 972
rect 13889 970 13893 971
rect 13903 970 13940 971
rect 13665 967 13668 968
rect 13363 964 13372 966
rect 13363 951 13368 964
rect 13416 955 13435 958
rect 13470 955 13494 967
rect 13527 959 13545 967
rect 13600 959 13601 967
rect 13272 948 13282 950
rect 13282 947 13285 948
rect 13287 945 13296 947
rect 13260 942 13262 945
rect 13296 943 13307 945
rect 13308 943 13309 951
rect 13335 943 13341 951
rect 13259 939 13260 942
rect 13307 938 13341 943
rect 13173 924 13174 938
rect 13123 915 13132 924
rect 13170 920 13179 924
rect 13170 915 13184 920
rect 13114 912 13123 915
rect 13114 911 13117 912
rect 13107 908 13116 911
rect 13095 907 13116 908
rect 13095 905 13113 907
rect 13153 905 13159 911
rect 13173 906 13188 915
rect 13213 908 13222 937
rect 13095 900 13107 905
rect 13091 898 13094 900
rect 13095 899 13096 900
rect 13101 899 13107 900
rect 13159 899 13165 905
rect 13172 904 13184 906
rect 13211 904 13213 908
rect 13251 907 13259 938
rect 13308 926 13309 938
rect 13335 935 13363 938
rect 13335 931 13365 935
rect 13367 931 13368 951
rect 13435 946 13497 955
rect 13545 952 13553 959
rect 13599 951 13600 958
rect 13668 954 13672 967
rect 13848 966 13856 969
rect 13886 968 13889 970
rect 13882 967 13886 968
rect 13877 965 13882 967
rect 13903 965 13918 970
rect 13927 969 13931 970
rect 13940 969 13941 970
rect 13997 969 14002 975
rect 14038 971 14047 980
rect 14103 978 14115 981
rect 14103 971 14112 978
rect 14382 972 14398 986
rect 14421 972 14422 996
rect 14427 991 14448 996
rect 14432 990 14448 991
rect 14565 989 14571 996
rect 14617 989 14623 996
rect 14637 990 14648 996
rect 14683 990 14692 1008
rect 14432 972 14448 988
rect 14565 985 14573 989
rect 14571 983 14573 985
rect 14481 974 14509 978
rect 14511 974 14522 978
rect 13931 965 13936 969
rect 13941 965 13943 968
rect 14002 965 14005 969
rect 13843 964 13847 965
rect 13918 964 13921 965
rect 13943 964 13944 965
rect 13839 962 13843 964
rect 13453 945 13463 946
rect 13485 945 13486 946
rect 13449 943 13453 945
rect 13497 943 13517 946
rect 13598 943 13599 950
rect 13671 943 13672 950
rect 13720 943 13726 949
rect 13766 948 13772 949
rect 13803 948 13839 962
rect 13923 959 13927 962
rect 13938 960 13942 963
rect 14047 962 14056 971
rect 14080 961 14083 963
rect 14094 962 14103 971
rect 14388 970 14422 972
rect 14431 971 14432 972
rect 14478 971 14481 974
rect 14427 970 14432 971
rect 14477 970 14478 971
rect 14388 968 14432 970
rect 14475 969 14477 970
rect 14384 965 14385 967
rect 14158 961 14167 963
rect 14075 959 14080 961
rect 13766 947 13803 948
rect 13766 943 13772 947
rect 13858 946 13864 952
rect 13904 946 13910 952
rect 13926 949 13927 959
rect 14073 958 14075 959
rect 14169 958 14175 961
rect 13944 955 13948 958
rect 14012 955 14014 958
rect 13948 946 13958 955
rect 13437 931 13445 943
rect 13449 941 13483 943
rect 13335 928 13396 931
rect 13335 917 13341 928
rect 13363 926 13396 928
rect 13357 925 13396 926
rect 13415 925 13421 926
rect 13357 921 13421 925
rect 13357 920 13443 921
rect 13335 915 13342 917
rect 13335 913 13344 915
rect 13363 914 13369 920
rect 13409 914 13415 920
rect 13418 917 13443 920
rect 13427 915 13443 917
rect 13432 913 13443 915
rect 13449 913 13451 941
rect 13480 939 13483 941
rect 13335 909 13350 913
rect 13437 909 13451 913
rect 13481 909 13483 939
rect 13487 931 13495 943
rect 13517 934 13580 943
rect 13714 938 13720 943
rect 13732 941 13768 943
rect 13732 939 13737 941
rect 13673 937 13720 938
rect 13734 937 13737 939
rect 13772 937 13778 943
rect 13852 940 13858 946
rect 13910 940 13916 946
rect 13673 936 13716 937
rect 13597 934 13598 936
rect 13619 934 13673 936
rect 13553 922 13568 934
rect 13580 933 13619 934
rect 13597 929 13598 933
rect 13729 929 13732 936
rect 13856 933 13858 934
rect 13250 904 13251 906
rect 13310 905 13311 909
rect 13316 903 13322 909
rect 13335 903 13354 909
rect 13362 903 13368 909
rect 13170 899 13172 903
rect 13210 899 13211 903
rect 13169 897 13170 899
rect 13209 897 13210 899
rect 13083 884 13091 896
rect 13095 894 13113 896
rect 13168 895 13169 896
rect 13248 895 13250 903
rect 13310 897 13316 903
rect 13335 897 13374 903
rect 13376 897 13388 905
rect 13449 904 13466 909
rect 13553 904 13568 920
rect 13595 906 13597 928
rect 13457 903 13458 904
rect 13466 903 13470 904
rect 13485 903 13487 904
rect 13447 901 13448 903
rect 13458 899 13464 903
rect 13470 900 13489 903
rect 13594 900 13606 905
rect 13616 900 13628 905
rect 13669 904 13671 928
rect 13720 904 13729 928
rect 13852 925 13856 933
rect 13765 904 13768 909
rect 13806 908 13841 910
rect 13801 907 13806 908
rect 13841 907 13849 908
rect 13852 907 13854 915
rect 13876 909 13877 929
rect 13924 928 13926 944
rect 13958 942 13963 946
rect 14014 942 14026 955
rect 14175 951 14188 958
rect 14398 956 14414 968
rect 14416 956 14432 968
rect 14471 965 14475 968
rect 14469 963 14471 965
rect 14467 961 14469 963
rect 14522 961 14535 974
rect 14571 967 14574 983
rect 14573 961 14574 967
rect 14577 967 14578 989
rect 14616 985 14623 989
rect 14644 987 14646 990
rect 14616 983 14617 985
rect 14637 984 14638 986
rect 14577 963 14579 967
rect 14610 963 14611 966
rect 14615 965 14617 983
rect 14646 981 14649 987
rect 14649 979 14650 981
rect 14651 975 14652 977
rect 14652 972 14653 975
rect 14692 973 14700 990
rect 14654 965 14657 969
rect 14577 961 14581 963
rect 14615 962 14616 965
rect 14657 963 14658 965
rect 14463 958 14466 961
rect 14535 959 14538 961
rect 14461 953 14463 958
rect 14538 957 14540 959
rect 14296 952 14333 953
rect 14460 952 14461 953
rect 14540 952 14542 957
rect 14568 955 14574 961
rect 14581 959 14587 961
rect 14588 957 14594 959
rect 14614 957 14620 961
rect 14658 960 14659 963
rect 14659 958 14660 960
rect 14594 956 14620 957
rect 14296 951 14321 952
rect 14333 951 14334 952
rect 14190 948 14194 951
rect 14261 948 14288 951
rect 14336 948 14343 951
rect 14388 949 14389 952
rect 14343 943 14354 948
rect 14389 945 14391 949
rect 14424 947 14425 952
rect 14459 951 14460 952
rect 14457 948 14459 951
rect 14354 942 14358 943
rect 14026 939 14027 942
rect 14358 939 14363 942
rect 14363 938 14365 939
rect 13921 917 13923 920
rect 13918 915 13920 916
rect 13915 913 13918 915
rect 13912 911 13915 913
rect 13910 910 13912 911
rect 13796 906 13801 907
rect 13849 906 13858 907
rect 13785 904 13796 906
rect 13719 900 13720 903
rect 13763 900 13765 903
rect 13773 901 13785 904
rect 13852 900 13854 906
rect 13876 904 13877 906
rect 13944 904 13960 920
rect 13968 915 13994 938
rect 14028 931 14034 938
rect 14365 937 14367 938
rect 14367 933 14383 937
rect 14383 932 14388 933
rect 14391 932 14399 944
rect 14038 920 14046 927
rect 14046 918 14053 920
rect 14053 915 14065 918
rect 13994 910 14000 915
rect 14065 914 14069 915
rect 14072 914 14073 929
rect 14388 927 14404 932
rect 14425 929 14429 945
rect 14455 943 14457 948
rect 14542 944 14545 951
rect 14562 949 14568 955
rect 14594 951 14638 956
rect 14660 955 14662 958
rect 14620 949 14626 951
rect 14662 948 14665 955
rect 14454 942 14455 943
rect 14665 942 14668 948
rect 14700 943 14701 973
rect 14808 951 14824 954
rect 14736 943 14759 951
rect 14824 943 14831 951
rect 14453 940 14454 942
rect 14452 939 14453 940
rect 14668 939 14669 942
rect 14451 937 14452 938
rect 14448 933 14451 937
rect 14446 932 14448 933
rect 14669 932 14670 938
rect 14698 932 14700 942
rect 14730 939 14736 943
rect 14831 939 14835 943
rect 14728 938 14730 939
rect 14835 938 14838 939
rect 14718 932 14728 938
rect 14835 936 14840 938
rect 14429 927 14430 928
rect 14443 927 14446 932
rect 14567 927 14568 929
rect 14399 923 14400 926
rect 14404 924 14441 927
rect 14131 921 14162 922
rect 14122 920 14131 921
rect 14162 920 14169 921
rect 14429 920 14430 924
rect 14093 917 14122 920
rect 14169 917 14184 920
rect 14091 916 14093 917
rect 14088 915 14091 916
rect 14184 915 14192 917
rect 14401 915 14402 917
rect 14430 915 14431 920
rect 14435 915 14444 924
rect 14482 915 14491 924
rect 14566 922 14567 927
rect 14565 920 14566 922
rect 14564 918 14565 920
rect 14563 916 14564 918
rect 14081 914 14088 915
rect 14192 914 14201 915
rect 14426 914 14435 915
rect 14069 911 14435 914
rect 14072 910 14073 911
rect 14075 910 14077 911
rect 14211 910 14219 911
rect 14000 909 14002 910
rect 13877 903 13878 904
rect 13941 903 13944 904
rect 14002 903 14010 909
rect 14071 908 14075 910
rect 14219 907 14232 910
rect 14232 906 14237 907
rect 14064 904 14069 906
rect 14237 904 14247 906
rect 13878 900 13881 903
rect 13931 900 13944 903
rect 13335 895 13390 897
rect 13464 895 13470 899
rect 13484 898 13485 900
rect 13083 862 13091 874
rect 13095 864 13097 894
rect 13167 893 13168 894
rect 13208 893 13209 894
rect 13335 893 13392 895
rect 13470 893 13471 895
rect 13483 894 13484 897
rect 13489 896 13658 900
rect 13717 897 13719 900
rect 13714 896 13720 897
rect 13760 896 13763 900
rect 13590 894 13592 896
rect 13594 895 13595 896
rect 13658 895 13720 896
rect 13162 889 13168 893
rect 13207 889 13208 893
rect 13247 889 13248 893
rect 13303 889 13310 893
rect 13335 892 13400 893
rect 13148 888 13168 889
rect 13148 878 13162 888
rect 13204 879 13207 889
rect 13245 878 13247 889
rect 13300 879 13303 889
rect 13135 868 13148 878
rect 13201 869 13204 878
rect 13244 875 13245 878
rect 13299 875 13300 878
rect 13242 868 13244 875
rect 13297 869 13299 875
rect 13132 866 13135 868
rect 13095 862 13098 864
rect 13129 862 13132 866
rect 13179 859 13188 868
rect 13200 866 13201 868
rect 13199 862 13200 866
rect 13094 857 13096 858
rect 13101 857 13107 859
rect 13095 853 13107 857
rect 13159 853 13165 859
rect 13171 857 13179 859
rect 13198 858 13199 862
rect 13240 859 13242 867
rect 13294 859 13297 868
rect 13312 864 13315 892
rect 13362 891 13388 892
rect 13386 861 13388 891
rect 13392 881 13400 892
rect 13471 879 13491 893
rect 13539 879 13553 894
rect 13582 881 13590 893
rect 13594 891 13628 893
rect 13447 876 13448 879
rect 13477 876 13478 879
rect 13491 877 13503 879
rect 13537 877 13539 879
rect 13491 875 13537 877
rect 13362 859 13388 861
rect 13392 859 13400 871
rect 13445 869 13446 871
rect 13474 868 13475 870
rect 13442 860 13444 866
rect 13471 860 13474 867
rect 13594 859 13596 891
rect 13626 873 13628 891
rect 13632 881 13640 893
rect 13714 891 13720 895
rect 13758 891 13760 895
rect 13772 891 13778 897
rect 13852 894 13858 900
rect 13881 896 13896 900
rect 13896 895 13897 896
rect 13910 895 13944 900
rect 14010 899 14016 903
rect 14060 901 14064 904
rect 13668 881 13669 889
rect 13712 881 13715 891
rect 13720 885 13726 891
rect 13752 881 13758 891
rect 13766 885 13772 891
rect 13855 883 13856 891
rect 13858 888 13864 894
rect 13897 893 13916 895
rect 13627 865 13628 872
rect 13662 870 13668 880
rect 13707 870 13712 881
rect 13656 868 13662 870
rect 13706 868 13707 870
rect 13746 869 13752 881
rect 13895 872 13898 892
rect 13904 888 13910 893
rect 13928 888 13944 895
rect 14016 894 14027 899
rect 14055 898 14059 900
rect 14052 897 14055 898
rect 14048 894 14052 897
rect 14072 895 14075 900
rect 14247 897 14282 904
rect 14328 902 14341 903
rect 14307 900 14325 902
rect 14346 900 14369 902
rect 14305 899 14317 900
rect 14369 899 14378 900
rect 14378 898 14379 899
rect 14403 898 14404 904
rect 14298 897 14305 898
rect 14027 886 14058 894
rect 14075 893 14077 895
rect 14077 891 14079 893
rect 14282 891 14305 897
rect 14379 894 14386 898
rect 14386 891 14392 894
rect 14404 891 14405 897
rect 14017 880 14058 886
rect 14079 886 14152 891
rect 14282 889 14304 891
rect 14079 881 14229 886
rect 14290 882 14298 889
rect 14304 887 14309 889
rect 14309 886 14311 887
rect 14392 886 14405 891
rect 14433 887 14436 903
rect 14491 901 14500 915
rect 14561 911 14562 914
rect 14588 909 14620 914
rect 14555 903 14559 906
rect 14562 903 14568 909
rect 14588 904 14626 909
rect 14657 904 14718 932
rect 14837 931 14840 936
rect 14836 922 14840 931
rect 14585 903 14626 904
rect 14655 903 14657 904
rect 14665 903 14666 904
rect 14542 901 14554 902
rect 14500 899 14504 901
rect 14522 900 14542 901
rect 14516 899 14522 900
rect 14542 895 14544 900
rect 14568 897 14574 903
rect 14602 899 14603 901
rect 14540 892 14542 895
rect 14539 891 14540 892
rect 14017 876 14034 880
rect 14058 876 14076 880
rect 14079 876 14099 881
rect 14151 876 14242 881
rect 14076 875 14242 876
rect 14283 875 14290 882
rect 14311 876 14335 886
rect 14392 882 14406 886
rect 14405 881 14408 882
rect 14405 878 14406 881
rect 14408 880 14409 881
rect 14335 875 14338 876
rect 14014 874 14016 875
rect 14075 874 14245 875
rect 14012 873 14014 874
rect 14073 873 14075 874
rect 14071 872 14073 873
rect 14076 872 14242 874
rect 14245 873 14253 874
rect 14253 872 14261 873
rect 14280 872 14283 875
rect 14338 874 14340 875
rect 14340 873 14343 874
rect 14343 872 14345 873
rect 14354 872 14366 878
rect 14409 875 14418 880
rect 14436 876 14438 886
rect 14527 882 14539 891
rect 14521 881 14527 882
rect 14493 880 14509 881
rect 14517 880 14521 881
rect 14586 880 14601 899
rect 14614 897 14620 903
rect 14651 901 14655 903
rect 14640 895 14651 901
rect 14664 899 14665 901
rect 14637 892 14640 895
rect 14636 891 14637 892
rect 14628 886 14636 891
rect 14465 875 14488 880
rect 14616 876 14648 886
rect 14661 880 14664 898
rect 14660 876 14661 880
rect 14696 878 14698 904
rect 14836 903 14837 922
rect 14851 915 14860 924
rect 14898 915 14907 924
rect 14842 906 14847 915
rect 14912 906 14916 915
rect 14817 881 14836 901
rect 13650 866 13656 868
rect 13745 867 13746 868
rect 13744 866 13745 867
rect 13649 865 13650 866
rect 13627 860 13649 865
rect 13703 862 13706 866
rect 13628 859 13649 860
rect 13700 859 13706 862
rect 13170 855 13179 857
rect 13095 850 13104 853
rect 13107 850 13113 853
rect 13158 852 13159 853
rect 13168 852 13179 855
rect 13115 851 13163 852
rect 13166 851 13168 852
rect 13115 850 13166 851
rect 13170 850 13179 852
rect 13105 847 13113 850
rect 13105 842 13109 847
rect 13158 840 13159 850
rect 13194 845 13198 858
rect 13237 846 13240 858
rect 13290 846 13294 858
rect 13310 851 13316 857
rect 13339 856 13343 859
rect 13633 858 13634 859
rect 13316 845 13322 851
rect 13334 845 13339 856
rect 13368 851 13374 857
rect 13441 855 13442 858
rect 13470 855 13471 858
rect 13700 857 13703 859
rect 13702 856 13703 857
rect 13698 855 13702 856
rect 13362 845 13368 851
rect 13376 847 13388 855
rect 13592 853 13593 855
rect 13439 851 13440 853
rect 13190 841 13194 845
rect 13236 841 13237 845
rect 13288 842 13290 845
rect 13188 840 13190 841
rect 13332 840 13334 845
rect 13436 841 13439 850
rect 13466 841 13469 850
rect 13593 841 13595 849
rect 13634 842 13635 849
rect 13695 847 13702 855
rect 13692 842 13695 847
rect 13698 845 13702 847
rect 13732 845 13744 865
rect 13856 859 13858 872
rect 14009 871 14011 872
rect 14069 871 14071 872
rect 13692 841 13694 842
rect 13689 840 13692 841
rect 13696 840 13698 845
rect 13729 844 13736 845
rect 13891 844 13895 870
rect 14004 868 14009 871
rect 14064 869 14068 871
rect 14152 869 14376 872
rect 14418 871 14424 875
rect 14455 871 14465 875
rect 14579 872 14582 876
rect 14613 875 14648 876
rect 14424 869 14430 871
rect 14437 869 14465 871
rect 14061 867 14063 868
rect 14001 866 14003 867
rect 14059 866 14061 867
rect 14168 866 14376 869
rect 14430 868 14431 869
rect 14437 868 14455 869
rect 14431 867 14435 868
rect 14450 867 14453 868
rect 13991 860 14001 866
rect 14049 862 14059 866
rect 14168 863 14378 866
rect 14281 862 14290 863
rect 14364 862 14386 863
rect 14407 862 14408 867
rect 14571 863 14579 872
rect 14626 869 14627 874
rect 14746 873 14757 874
rect 14774 873 14785 874
rect 14746 872 14754 873
rect 14778 872 14785 873
rect 14290 860 14293 862
rect 13986 857 13991 860
rect 13977 852 13986 857
rect 14293 852 14308 860
rect 14364 854 14378 862
rect 14386 856 14419 862
rect 14567 857 14571 862
rect 14494 856 14506 857
rect 14419 855 14425 856
rect 14443 855 14465 856
rect 14425 854 14465 855
rect 14486 854 14506 856
rect 13975 851 13977 852
rect 14308 851 14310 852
rect 13972 850 13975 851
rect 14310 850 14312 851
rect 13937 849 13943 850
rect 13970 849 13972 850
rect 13919 844 13970 849
rect 13983 844 13989 850
rect 14033 845 14036 849
rect 14313 845 14321 849
rect 14364 846 14376 854
rect 14494 851 14526 854
rect 14495 847 14526 851
rect 14564 849 14566 856
rect 14564 847 14565 849
rect 13729 840 13733 844
rect 13110 836 13111 840
rect 13111 833 13112 836
rect 13158 832 13160 840
rect 13176 832 13188 840
rect 13235 838 13236 840
rect 13287 838 13288 840
rect 13234 832 13235 838
rect 13286 833 13287 838
rect 13329 832 13332 840
rect 13435 837 13436 840
rect 13434 833 13435 836
rect 13463 834 13465 840
rect 13635 837 13636 840
rect 13596 832 13600 837
rect 13687 832 13696 840
rect 13725 834 13733 840
rect 13725 832 13729 834
rect 13112 817 13120 832
rect 13158 825 13162 832
rect 13175 830 13176 832
rect 13328 830 13329 832
rect 13174 828 13175 830
rect 13233 828 13234 830
rect 13284 828 13285 830
rect 13173 825 13174 828
rect 13160 817 13162 825
rect 13232 824 13233 828
rect 13283 824 13284 827
rect 13326 824 13328 829
rect 13171 819 13173 824
rect 13231 819 13232 824
rect 13278 820 13283 824
rect 11528 805 11536 808
rect 11528 804 11530 805
rect 11531 800 11532 802
rect 11532 797 11534 800
rect 11289 790 11291 793
rect 11097 758 11113 763
rect 11162 773 11223 785
rect 11230 779 11243 790
rect 11229 774 11243 779
rect 11273 777 11291 790
rect 11382 789 11383 793
rect 11413 789 11414 795
rect 11273 774 11289 777
rect 11162 759 11227 773
rect 11193 758 11209 759
rect 11211 758 11227 759
rect 11254 758 11255 760
rect 11289 758 11305 774
rect 11383 767 11387 785
rect 11414 779 11415 788
rect 11463 787 11465 794
rect 11528 790 11529 794
rect 11534 791 11537 797
rect 11569 792 11585 808
rect 11619 802 11647 808
rect 11683 806 11703 816
rect 13120 809 13124 817
rect 13162 811 13163 817
rect 13170 815 13171 819
rect 13230 815 13231 819
rect 13278 815 13282 820
rect 13324 819 13326 824
rect 13169 809 13170 814
rect 13228 809 13230 814
rect 13278 809 13280 815
rect 13321 814 13324 818
rect 13374 814 13390 824
rect 13392 814 13408 824
rect 13428 817 13434 832
rect 13317 809 13321 814
rect 13361 809 13368 814
rect 13413 808 13421 814
rect 13426 811 13428 817
rect 13456 811 13463 832
rect 13597 827 13601 832
rect 13636 827 13642 832
rect 13685 830 13687 832
rect 13724 830 13725 832
rect 13455 809 13456 811
rect 13470 808 13486 824
rect 13586 822 13652 827
rect 13678 824 13685 830
rect 13721 825 13724 830
rect 13727 828 13729 832
rect 13858 832 13860 844
rect 13870 840 13882 844
rect 13898 842 13919 844
rect 13889 841 13898 842
rect 13884 840 13891 841
rect 13870 836 13884 840
rect 13586 821 13642 822
rect 13577 814 13586 821
rect 13597 818 13601 821
rect 13575 811 13577 814
rect 13600 811 13601 817
rect 13636 811 13642 821
rect 13652 814 13656 821
rect 13670 819 13678 824
rect 13718 819 13721 824
rect 13670 818 13672 819
rect 13670 815 13671 818
rect 13716 817 13718 819
rect 13715 816 13716 817
rect 13656 811 13657 814
rect 13669 812 13670 813
rect 13715 812 13718 816
rect 13748 812 13760 815
rect 13658 811 13667 812
rect 13493 808 13512 809
rect 13518 808 13520 809
rect 13125 804 13126 807
rect 11613 794 11647 802
rect 13126 799 13128 803
rect 13163 799 13164 803
rect 13166 800 13169 808
rect 13226 800 13228 808
rect 13128 794 13130 798
rect 13166 794 13168 800
rect 13224 794 13226 798
rect 11609 791 11611 794
rect 11619 790 11647 794
rect 11465 781 11466 787
rect 11528 782 11545 790
rect 11415 766 11420 779
rect 11467 774 11475 780
rect 11529 776 11545 782
rect 11601 779 11609 790
rect 11598 778 11609 779
rect 11613 788 11647 790
rect 11529 774 11539 776
rect 11475 773 11477 774
rect 11387 760 11388 766
rect 11420 759 11422 766
rect 11477 765 11491 773
rect 11529 766 11530 774
rect 11545 768 11550 776
rect 11598 770 11607 778
rect 11526 765 11530 766
rect 11472 764 11505 765
rect 11526 764 11536 765
rect 11472 759 11478 764
rect 11022 756 11028 758
rect 11099 757 11113 758
rect 11225 757 11228 758
rect 11107 756 11160 757
rect 10940 754 10941 756
rect 11022 754 11031 756
rect 10704 738 10710 739
rect 10750 738 10756 744
rect 10790 738 10799 747
rect 10837 738 10846 747
rect 10929 746 10943 754
rect 11017 747 11031 754
rect 11102 750 11166 756
rect 11229 750 11244 756
rect 11251 754 11252 756
rect 11293 752 11294 753
rect 11017 746 11022 747
rect 10943 745 10946 746
rect 10456 734 10457 736
rect 10458 727 10461 733
rect 10530 731 10545 736
rect 10698 732 10704 738
rect 10756 733 10762 738
rect 10810 734 10822 738
rect 10863 734 10879 744
rect 10941 742 10942 745
rect 10946 742 10985 745
rect 11015 743 11022 746
rect 11108 745 11123 750
rect 11154 747 11163 750
rect 11108 744 11114 745
rect 11154 744 11160 747
rect 10942 740 10985 742
rect 10946 737 10985 740
rect 11008 739 11015 743
rect 11017 739 11022 743
rect 11163 742 11177 747
rect 11244 745 11257 750
rect 11293 747 11301 752
rect 11389 751 11390 756
rect 11423 750 11426 756
rect 11478 753 11484 759
rect 11489 758 11505 764
rect 11507 758 11523 764
rect 11530 759 11536 764
rect 11550 762 11553 768
rect 11589 761 11598 770
rect 11524 753 11530 759
rect 11555 756 11557 760
rect 11585 757 11586 758
rect 11243 742 11245 745
rect 11257 742 11263 745
rect 11294 744 11301 747
rect 11390 746 11391 750
rect 11426 744 11428 750
rect 11512 745 11515 747
rect 11303 742 11304 744
rect 11557 743 11565 756
rect 11586 754 11589 757
rect 11601 756 11609 768
rect 11613 758 11615 788
rect 11644 787 11647 788
rect 11651 779 11694 791
rect 13131 785 13134 793
rect 13165 790 13167 793
rect 13168 790 13182 794
rect 13165 786 13182 790
rect 11645 776 11694 779
rect 11645 770 11654 776
rect 11665 774 11681 776
rect 11694 774 11715 776
rect 13134 775 13139 785
rect 11654 764 11663 770
rect 11657 763 11663 764
rect 11681 768 11715 774
rect 13139 771 13140 775
rect 13166 774 13182 786
rect 13216 790 13224 794
rect 13262 792 13278 808
rect 13312 801 13317 808
rect 13357 801 13361 808
rect 13413 807 13424 808
rect 13454 807 13470 808
rect 13520 807 13521 808
rect 13569 807 13575 810
rect 13642 809 13643 811
rect 13597 808 13599 809
rect 13657 808 13667 811
rect 13714 808 13715 812
rect 13748 808 13764 812
rect 13766 808 13782 824
rect 13784 808 13800 824
rect 13858 820 13866 832
rect 13870 831 13886 832
rect 13870 830 13880 831
rect 13802 808 13811 812
rect 13861 810 13862 811
rect 13586 807 13596 808
rect 13413 806 13425 807
rect 13420 804 13425 806
rect 13312 792 13315 801
rect 13216 774 13232 790
rect 13262 774 13278 790
rect 13312 787 13328 790
rect 13307 781 13328 787
rect 13348 787 13357 801
rect 13420 792 13424 804
rect 13453 803 13470 807
rect 13521 806 13524 807
rect 13452 799 13453 803
rect 13450 794 13452 798
rect 13454 792 13470 803
rect 13493 798 13505 806
rect 13524 803 13527 806
rect 13547 803 13586 807
rect 13643 803 13644 807
rect 13654 803 13669 808
rect 13748 807 13765 808
rect 13770 807 13782 808
rect 13508 799 13547 803
rect 13558 799 13564 803
rect 13569 799 13575 803
rect 13644 799 13645 803
rect 13348 785 13359 787
rect 13368 785 13380 791
rect 13420 785 13421 792
rect 13448 788 13450 792
rect 13337 783 13359 785
rect 13369 783 13380 785
rect 13419 783 13424 785
rect 13331 781 13336 783
rect 13301 775 13307 781
rect 13312 774 13328 781
rect 13346 779 13348 783
rect 13353 781 13359 783
rect 13380 781 13384 783
rect 13359 775 13365 781
rect 13368 778 13380 779
rect 13168 771 13172 774
rect 11658 759 11661 763
rect 11681 758 11697 768
rect 11715 762 11732 768
rect 11718 758 11724 762
rect 11732 760 11738 762
rect 11738 758 11742 760
rect 11764 758 11770 764
rect 11613 757 11628 758
rect 11613 756 11632 757
rect 11589 750 11594 754
rect 11629 752 11647 756
rect 11664 753 11670 756
rect 11712 753 11718 758
rect 11613 750 11647 752
rect 11670 751 11718 753
rect 11770 752 11776 758
rect 13140 754 13148 771
rect 13172 754 13179 771
rect 13182 758 13198 774
rect 13200 758 13216 774
rect 13278 772 13286 774
rect 13304 772 13312 774
rect 13378 772 13380 778
rect 13384 772 13392 779
rect 13417 778 13419 783
rect 13420 778 13424 783
rect 13417 774 13424 778
rect 13417 772 13419 774
rect 13278 758 13294 772
rect 13296 758 13312 772
rect 13359 757 13422 772
rect 13446 760 13448 786
rect 13454 774 13470 790
rect 13481 782 13489 794
rect 13493 793 13514 794
rect 13552 793 13558 799
rect 13493 792 13511 793
rect 13470 763 13474 767
rect 13481 763 13489 772
rect 13493 763 13495 792
rect 13646 788 13648 796
rect 13654 794 13676 803
rect 13654 792 13669 794
rect 13706 790 13714 806
rect 13744 804 13746 807
rect 13750 806 13764 807
rect 13748 803 13764 806
rect 13800 805 13816 808
rect 13798 803 13816 805
rect 13736 791 13744 803
rect 13746 801 13782 803
rect 13746 793 13766 801
rect 13779 800 13782 801
rect 13780 793 13782 800
rect 13786 799 13794 803
rect 13798 799 13820 803
rect 13800 794 13820 799
rect 13858 798 13866 810
rect 13870 800 13872 830
rect 13889 826 13891 840
rect 13931 838 13937 844
rect 13989 838 13995 844
rect 14028 841 14033 845
rect 14321 841 14326 845
rect 14320 832 14328 841
rect 14332 834 14334 839
rect 14364 834 14366 846
rect 14624 845 14626 865
rect 14658 863 14660 872
rect 14695 863 14696 872
rect 14746 871 14748 872
rect 14784 871 14785 872
rect 14817 868 14831 881
rect 14810 866 14823 868
rect 14810 865 14822 866
rect 14851 865 14856 866
rect 14657 857 14658 862
rect 14655 849 14656 855
rect 14376 844 14379 845
rect 14332 832 14366 834
rect 14370 840 14379 844
rect 14370 832 14378 840
rect 14379 832 14383 840
rect 14383 830 14384 832
rect 13904 826 13905 830
rect 14015 829 14018 830
rect 13991 827 14026 829
rect 13889 818 13890 826
rect 13987 825 13991 827
rect 13985 824 13987 825
rect 13905 812 13907 824
rect 13890 800 13893 811
rect 13958 808 13985 824
rect 13989 812 13993 817
rect 13999 812 14015 827
rect 14026 824 14051 827
rect 13994 811 14015 812
rect 13870 798 13904 800
rect 13890 795 13893 798
rect 13648 778 13651 788
rect 13651 769 13653 778
rect 13654 774 13669 790
rect 13706 774 13720 790
rect 13743 781 13744 788
rect 13653 765 13654 769
rect 13470 762 13495 763
rect 13524 762 13527 763
rect 13470 760 13527 762
rect 13470 758 13486 760
rect 13654 759 13655 763
rect 11594 749 11630 750
rect 11613 744 11625 749
rect 11680 744 11691 749
rect 13148 746 13151 754
rect 13179 748 13184 754
rect 13184 745 13188 748
rect 13378 745 13380 757
rect 13383 745 13417 757
rect 13422 756 13424 757
rect 13531 756 13558 759
rect 13655 757 13656 759
rect 13670 758 13686 772
rect 13688 758 13704 772
rect 13736 769 13744 781
rect 13748 774 13766 793
rect 13800 792 13816 794
rect 13800 774 13816 790
rect 13846 774 13861 790
rect 13863 775 13865 792
rect 13870 786 13882 794
rect 13892 786 13904 794
rect 13906 790 13907 808
rect 13993 805 14003 811
rect 14051 808 14192 824
rect 14254 808 14270 824
rect 14272 808 14288 824
rect 14332 820 14344 828
rect 14354 820 14366 828
rect 14384 826 14385 830
rect 14410 828 14412 845
rect 14332 810 14334 820
rect 14385 816 14388 824
rect 14412 819 14413 828
rect 14440 819 14443 845
rect 14482 833 14488 845
rect 14529 843 14531 844
rect 14654 843 14655 847
rect 14565 838 14566 843
rect 14532 827 14533 836
rect 14566 827 14567 836
rect 14622 825 14624 840
rect 14653 837 14654 843
rect 14651 827 14653 836
rect 14693 829 14695 862
rect 14806 855 14822 865
rect 14859 864 14863 868
rect 14743 845 14806 855
rect 14851 851 14859 864
rect 14734 844 14743 845
rect 14728 842 14734 844
rect 14726 840 14728 842
rect 14482 811 14488 823
rect 14650 821 14651 826
rect 14691 820 14693 827
rect 14707 825 14726 840
rect 14706 824 14707 825
rect 14534 817 14535 820
rect 14567 816 14568 820
rect 14535 811 14540 816
rect 14568 811 14569 816
rect 14621 811 14622 818
rect 14635 811 14641 817
rect 14649 816 14650 820
rect 14690 818 14691 820
rect 14698 818 14706 824
rect 14647 812 14649 816
rect 14681 811 14687 817
rect 14689 816 14698 818
rect 14688 811 14698 816
rect 14444 808 14445 810
rect 14536 808 14537 810
rect 13998 803 14003 805
rect 14123 803 14132 808
rect 14170 803 14179 808
rect 13910 802 13919 803
rect 13908 798 13916 802
rect 13919 799 13934 802
rect 13934 798 13937 799
rect 13931 792 13937 798
rect 13989 792 13995 798
rect 14003 794 14012 803
rect 14114 794 14123 803
rect 14179 794 14188 803
rect 14105 792 14112 793
rect 13937 790 13943 792
rect 13748 772 13782 774
rect 13795 772 13800 774
rect 13893 772 13896 786
rect 13906 774 13912 790
rect 13937 786 13958 790
rect 13983 786 13989 792
rect 14099 791 14105 792
rect 14156 791 14160 793
rect 14192 792 14208 808
rect 14238 792 14254 808
rect 14265 803 14271 808
rect 14265 802 14280 803
rect 14259 796 14265 802
rect 14288 798 14304 808
rect 14311 802 14317 808
rect 14264 791 14265 793
rect 14297 791 14302 798
rect 14317 796 14323 802
rect 14335 800 14336 808
rect 14097 790 14099 791
rect 14096 787 14097 790
rect 14161 789 14163 790
rect 13942 774 13958 786
rect 14009 778 14036 781
rect 13992 774 14009 778
rect 14036 774 14044 778
rect 13748 769 13800 772
rect 13861 769 13867 772
rect 13896 771 13900 772
rect 13748 757 13752 765
rect 13784 758 13800 769
rect 13862 762 13879 769
rect 13896 762 13906 771
rect 13862 758 13878 762
rect 13879 760 13884 762
rect 13888 760 13900 762
rect 13884 759 13900 760
rect 13880 758 13900 759
rect 13958 758 13974 774
rect 14044 772 14047 774
rect 14112 772 14118 778
rect 14121 772 14123 779
rect 14163 772 14164 778
rect 14192 774 14208 790
rect 14238 774 14254 790
rect 14256 779 14265 791
rect 14047 763 14067 772
rect 14096 767 14097 769
rect 14106 766 14112 772
rect 14164 766 14170 772
rect 14185 763 14192 774
rect 14067 762 14069 763
rect 14069 759 14075 762
rect 13424 751 13445 756
rect 13445 747 13461 751
rect 13493 748 13505 756
rect 13656 754 13657 756
rect 13552 747 13558 753
rect 13583 747 13638 753
rect 13657 750 13658 754
rect 13658 747 13660 748
rect 13667 747 13676 756
rect 13746 747 13752 756
rect 13804 747 13810 753
rect 13811 747 13820 756
rect 13865 751 13868 758
rect 11691 743 11693 744
rect 11177 739 11186 742
rect 11263 741 11265 742
rect 11565 741 11566 743
rect 13151 741 13153 745
rect 11008 738 11022 739
rect 10995 737 11008 738
rect 11015 735 11017 738
rect 11186 735 11197 739
rect 11240 737 11241 739
rect 11197 734 11200 735
rect 10806 733 10888 734
rect 10756 732 10822 733
rect 10799 731 10822 732
rect 10545 726 10557 731
rect 10799 729 10806 731
rect 10810 730 10822 731
rect 10888 729 10891 732
rect 11007 731 11014 734
rect 11200 731 11209 734
rect 11237 733 11239 736
rect 11209 729 11216 731
rect 11232 729 11236 731
rect 10795 728 10799 729
rect 10788 726 10795 728
rect 10825 727 10826 729
rect 10891 728 10893 729
rect 10247 721 10318 723
rect 10071 719 10086 720
rect 10248 719 10318 721
rect 10350 719 10354 725
rect 10461 723 10463 726
rect 10074 716 10086 719
rect 8399 706 8409 709
rect 8410 706 8422 715
rect 8445 714 8447 715
rect 8447 709 8487 714
rect 8509 709 8521 714
rect 10010 712 10015 716
rect 10087 714 10090 716
rect 10239 712 10247 719
rect 10249 717 10259 719
rect 10249 712 10253 717
rect 8487 707 8521 709
rect 8487 706 8535 707
rect 8557 706 8563 712
rect 8615 706 8621 712
rect 7984 698 7995 701
rect 8078 698 8086 701
rect 8106 700 8114 701
rect 7447 688 7448 692
rect 7410 676 7444 678
rect 7448 676 7456 688
rect 7543 686 7549 692
rect 7601 686 7607 692
rect 7633 688 7640 692
rect 7749 691 7755 697
rect 7795 691 7801 697
rect 7841 691 7984 698
rect 8056 691 8078 698
rect 8112 692 8114 700
rect 8115 693 8121 698
rect 8134 694 8146 701
rect 7736 688 7738 691
rect 7633 687 7645 688
rect 7549 680 7555 686
rect 7595 680 7601 686
rect 7633 685 7648 687
rect 7655 685 7667 688
rect 7735 687 7736 688
rect 7734 685 7735 687
rect 7743 685 7749 691
rect 7801 685 7807 691
rect 7808 689 7829 691
rect 8051 689 8056 691
rect 8045 687 8051 689
rect 8114 688 8115 692
rect 8123 689 8126 691
rect 7812 685 7847 687
rect 7633 680 7645 685
rect 7648 680 7670 685
rect 7732 683 7734 685
rect 7670 676 7683 680
rect 7683 675 7688 676
rect 7697 675 7747 683
rect 7800 682 7812 685
rect 7791 680 7800 682
rect 7852 680 7854 685
rect 8035 684 8043 687
rect 8115 686 8116 687
rect 8028 682 8035 684
rect 7790 676 7791 680
rect 8021 679 8028 682
rect 8116 680 8118 682
rect 8016 678 8021 679
rect 8010 676 8016 678
rect 8118 676 8120 680
rect 8132 678 8139 684
rect 8151 682 8209 701
rect 8236 692 8237 698
rect 8300 692 8301 701
rect 8305 693 8313 703
rect 8320 702 8324 705
rect 8385 702 8410 706
rect 8507 704 8520 706
rect 8308 691 8313 693
rect 8324 692 8335 702
rect 8151 678 8184 682
rect 7446 672 7448 675
rect 7688 674 7747 675
rect 7697 672 7747 674
rect 7153 656 7156 662
rect 7077 643 7141 649
rect 7151 648 7153 656
rect 7197 652 7214 672
rect 7237 666 7244 672
rect 7410 666 7422 672
rect 7432 666 7444 672
rect 7674 666 7697 672
rect 7244 664 7450 666
rect 7663 664 7674 666
rect 7083 637 7110 643
rect 7129 637 7135 643
rect 7145 642 7151 647
rect 7155 642 7164 644
rect 7214 643 7222 652
rect 7391 642 7392 660
rect 6072 623 6099 629
rect 6893 626 6896 630
rect 7086 626 7110 637
rect 7145 635 7164 642
rect 7223 639 7227 642
rect 7227 636 7232 639
rect 7232 635 7240 636
rect 7145 630 7160 635
rect 7240 631 7276 635
rect 7144 626 7160 630
rect 7276 628 7296 631
rect 7390 630 7392 642
rect 7450 654 7609 664
rect 7621 654 7663 664
rect 7787 663 7790 674
rect 7854 663 7857 676
rect 8005 674 8010 676
rect 8002 673 8005 674
rect 7997 672 8002 673
rect 7991 670 7997 672
rect 8120 670 8123 676
rect 8139 671 8147 678
rect 8184 671 8192 678
rect 8209 676 8215 682
rect 8238 679 8239 682
rect 8240 677 8241 687
rect 8292 681 8305 682
rect 8292 679 8301 681
rect 8335 679 8340 692
rect 8385 688 8434 702
rect 8459 698 8505 704
rect 8523 703 8525 706
rect 8535 704 8555 706
rect 8563 704 8582 706
rect 8506 700 8521 702
rect 8451 694 8459 698
rect 8385 687 8410 688
rect 8434 687 8440 688
rect 8442 687 8451 694
rect 8367 678 8385 687
rect 8434 686 8442 687
rect 8440 685 8444 686
rect 8430 677 8437 683
rect 8444 682 8452 685
rect 8452 681 8457 682
rect 8457 680 8462 681
rect 8463 678 8466 679
rect 8234 676 8255 677
rect 8292 676 8298 677
rect 8215 673 8219 676
rect 7972 668 7991 670
rect 7935 664 7972 668
rect 7858 663 7935 664
rect 7749 655 7935 663
rect 8123 660 8136 670
rect 8147 660 8169 671
rect 8192 663 8202 671
rect 8219 663 8223 673
rect 8234 671 8240 676
rect 8241 672 8255 676
rect 8281 671 8298 676
rect 8339 671 8340 676
rect 8350 671 8365 677
rect 8240 665 8246 671
rect 8286 665 8292 671
rect 8330 663 8350 671
rect 8421 669 8430 677
rect 8469 676 8474 678
rect 8475 674 8481 676
rect 7450 652 7621 654
rect 7749 653 7864 655
rect 7450 642 7452 652
rect 7749 651 7861 653
rect 7749 649 7854 651
rect 7749 648 7817 649
rect 7749 645 7801 648
rect 7743 644 7807 645
rect 7721 643 7807 644
rect 7721 642 7739 643
rect 7450 634 7456 642
rect 7715 639 7732 642
rect 7743 639 7807 643
rect 7840 641 7852 649
rect 7857 643 7861 651
rect 7697 636 7715 639
rect 7451 630 7456 634
rect 7678 633 7697 636
rect 7749 633 7755 639
rect 7781 636 7787 639
rect 7795 633 7801 639
rect 7859 636 7861 643
rect 8136 642 8182 660
rect 8202 652 8232 663
rect 8212 647 8246 652
rect 8266 647 8267 660
rect 8303 652 8330 663
rect 8339 660 8340 663
rect 8212 646 8283 647
rect 8291 646 8320 652
rect 8212 643 8320 646
rect 8218 642 8223 643
rect 8136 641 8184 642
rect 7663 631 7678 633
rect 7467 630 7507 631
rect 7661 630 7663 631
rect 7306 628 7467 630
rect 7507 628 7536 630
rect 7390 626 7393 628
rect 7449 626 7456 628
rect 6100 623 6127 624
rect 5484 621 5485 622
rect 5388 615 5405 621
rect 5480 616 5484 621
rect 6896 618 6904 626
rect 6964 618 6971 625
rect 6904 617 6964 618
rect 5477 615 5480 616
rect 5405 611 5477 615
rect 7128 610 7144 626
rect 7393 615 7399 626
rect 7446 618 7449 625
rect 7536 622 7597 628
rect 7607 622 7657 630
rect 7857 627 7859 636
rect 7438 615 7446 618
rect 7399 613 7440 615
rect 7781 613 7794 624
rect 7835 616 7857 627
rect 8136 626 8182 641
rect 8186 637 8189 639
rect 8189 636 8191 637
rect 8191 633 8198 636
rect 8218 634 8232 642
rect 8266 634 8267 643
rect 8338 637 8339 653
rect 8380 652 8421 669
rect 8475 668 8483 674
rect 8487 670 8489 672
rect 8519 670 8521 700
rect 8525 690 8533 702
rect 8563 700 8569 704
rect 8609 700 8615 706
rect 8633 693 8644 702
rect 10015 696 10036 712
rect 10080 710 10104 712
rect 10084 705 10104 710
rect 10239 707 10249 712
rect 10246 705 10249 707
rect 10036 695 10038 696
rect 8487 668 8521 670
rect 8525 668 8533 680
rect 8644 678 8647 692
rect 10042 689 10043 692
rect 10040 678 10047 687
rect 10084 680 10086 705
rect 10090 700 10098 705
rect 10104 699 10110 705
rect 10244 701 10246 705
rect 10238 699 10246 701
rect 10110 694 10116 699
rect 10238 695 10244 699
rect 10116 692 10119 694
rect 10052 678 10086 680
rect 10090 678 10098 690
rect 10119 688 10120 692
rect 10232 689 10238 695
rect 10242 692 10243 694
rect 10241 688 10242 691
rect 10251 689 10253 712
rect 10283 715 10338 719
rect 10283 701 10306 715
rect 10314 713 10338 715
rect 10358 713 10359 715
rect 10319 708 10338 713
rect 10359 708 10363 713
rect 10463 710 10470 723
rect 10557 722 10587 726
rect 10806 724 10822 726
rect 10557 714 10599 722
rect 10326 701 10338 708
rect 10363 706 10364 708
rect 10470 705 10473 710
rect 10551 709 10600 710
rect 10283 695 10290 701
rect 10283 693 10296 695
rect 10283 689 10285 693
rect 10290 689 10296 693
rect 10301 691 10310 700
rect 10329 696 10338 701
rect 10369 696 10372 701
rect 10332 691 10338 696
rect 10240 685 10241 687
rect 10284 685 10285 689
rect 10302 687 10319 691
rect 10335 689 10338 691
rect 10372 689 10378 696
rect 10473 695 10510 705
rect 10551 702 10565 709
rect 10581 708 10600 709
rect 10597 703 10600 708
rect 10550 699 10551 701
rect 10510 693 10516 695
rect 10548 694 10550 699
rect 10516 692 10521 693
rect 10547 692 10548 694
rect 10337 687 10338 689
rect 10303 686 10319 687
rect 10378 686 10380 689
rect 10521 688 10537 692
rect 10537 687 10539 688
rect 10120 680 10122 685
rect 10239 680 10240 685
rect 10305 682 10308 686
rect 10310 682 10319 686
rect 10311 680 10312 682
rect 8647 676 8648 678
rect 10047 676 10048 678
rect 10051 676 10052 678
rect 10238 676 10239 678
rect 10312 677 10313 680
rect 8483 664 8486 666
rect 8487 656 8499 664
rect 8509 656 8521 664
rect 8648 661 8651 676
rect 8365 646 8380 652
rect 8487 648 8496 656
rect 8650 648 8651 661
rect 10047 660 10051 676
rect 10087 674 10090 676
rect 10052 666 10064 674
rect 10074 666 10086 674
rect 10122 660 10126 676
rect 10046 654 10047 658
rect 10126 657 10127 660
rect 8356 643 8363 646
rect 8351 641 8356 643
rect 8342 637 8351 641
rect 8198 631 8204 633
rect 8216 630 8232 634
rect 8207 626 8232 630
rect 8266 626 8268 630
rect 8200 622 8225 626
rect 7795 613 7835 616
rect 7406 610 7422 613
rect 7424 610 7440 613
rect 8200 610 8216 622
rect 8225 619 8233 622
rect 8233 618 8242 619
rect 8268 615 8273 626
rect 8300 620 8342 637
rect 8297 619 8300 620
rect 8291 618 8297 619
rect 8329 618 8336 620
rect 8325 615 8329 618
rect 8273 611 8294 615
rect 8316 611 8325 615
rect 8466 606 8490 629
rect 8496 626 8535 648
rect 8535 621 8544 626
rect 8641 622 8650 643
rect 10046 630 10048 654
rect 10126 630 10127 654
rect 10238 649 10290 663
rect 10311 662 10313 675
rect 10340 672 10352 685
rect 10380 672 10392 686
rect 10542 685 10548 687
rect 10548 683 10556 685
rect 10553 681 10557 683
rect 10553 676 10560 681
rect 10597 678 10599 703
rect 10600 697 10601 702
rect 10603 698 10611 710
rect 10756 694 10784 695
rect 10820 694 10822 724
rect 10826 714 10834 726
rect 10893 712 10895 728
rect 11216 727 11222 729
rect 11229 727 11232 729
rect 10949 720 10955 726
rect 11007 720 11013 726
rect 11213 723 11233 727
rect 11265 723 11286 741
rect 11291 738 11302 740
rect 11213 721 11229 723
rect 11208 720 11213 721
rect 11233 720 11241 723
rect 10955 714 10961 720
rect 11001 714 11007 720
rect 11201 717 11208 720
rect 11241 719 11244 720
rect 11286 719 11291 723
rect 11196 716 11201 717
rect 11244 716 11250 719
rect 11291 716 11295 719
rect 11299 716 11301 738
rect 11302 737 11303 738
rect 11305 737 11313 740
rect 11303 734 11313 737
rect 11305 729 11313 734
rect 11392 733 11393 741
rect 11429 737 11432 741
rect 11393 729 11394 733
rect 11422 729 11434 737
rect 11444 729 11456 737
rect 11519 729 11532 741
rect 11305 728 11314 729
rect 11310 726 11314 728
rect 11305 716 11313 718
rect 11187 713 11196 716
rect 11182 711 11187 713
rect 10601 693 10602 694
rect 10776 692 10784 694
rect 10788 692 10822 694
rect 10826 692 10834 704
rect 10893 694 10895 710
rect 11166 706 11182 711
rect 11250 706 11261 716
rect 11295 707 11313 716
rect 11277 706 11313 707
rect 11314 706 11337 726
rect 11394 724 11401 729
rect 11418 727 11421 729
rect 11434 725 11435 729
rect 11441 725 11447 729
rect 11395 723 11401 724
rect 11410 723 11418 725
rect 11422 723 11468 725
rect 11389 717 11395 723
rect 11422 717 11424 723
rect 11447 717 11453 723
rect 11454 717 11468 723
rect 11393 713 11395 714
rect 11391 709 11393 713
rect 11150 701 11166 706
rect 11261 705 11268 706
rect 11306 705 11339 706
rect 11261 702 11269 705
rect 11243 701 11277 702
rect 11303 701 11364 705
rect 11454 702 11456 717
rect 11460 713 11475 717
rect 11463 705 11475 713
rect 11532 712 11551 729
rect 11566 715 11600 741
rect 11695 723 11718 741
rect 13188 740 13196 745
rect 13414 742 13415 745
rect 13461 742 13481 747
rect 13481 741 13486 742
rect 13558 741 13564 747
rect 13604 741 13610 747
rect 13380 740 13382 741
rect 13153 737 13155 740
rect 13196 737 13201 740
rect 13370 739 13380 740
rect 13359 738 13380 739
rect 13486 738 13490 741
rect 13611 738 13620 747
rect 13658 745 13667 747
rect 13658 742 13673 745
rect 13658 738 13667 742
rect 13673 740 13677 742
rect 13752 741 13764 747
rect 13798 741 13811 747
rect 13867 744 13868 751
rect 13677 739 13680 740
rect 13201 736 13203 737
rect 13368 736 13387 738
rect 13156 733 13157 736
rect 13203 733 13207 736
rect 13157 727 13160 733
rect 13207 731 13211 733
rect 13211 729 13214 731
rect 13301 729 13307 735
rect 13359 729 13365 735
rect 13368 733 13405 736
rect 13412 733 13413 736
rect 13379 729 13405 733
rect 13408 729 13412 731
rect 13444 729 13445 730
rect 13214 726 13218 729
rect 13160 720 13164 726
rect 13218 720 13228 726
rect 13231 720 13243 724
rect 13307 723 13313 729
rect 13353 723 13359 729
rect 13405 726 13445 729
rect 13405 723 13444 726
rect 13490 725 13507 738
rect 13611 737 13612 738
rect 13680 736 13687 739
rect 13755 738 13764 741
rect 13802 738 13811 741
rect 13861 739 13868 744
rect 13896 742 13900 758
rect 13938 747 13947 756
rect 14003 747 14012 756
rect 14075 754 14086 759
rect 14179 758 14192 763
rect 14254 769 14263 774
rect 14264 769 14265 779
rect 14254 763 14265 769
rect 14268 763 14270 791
rect 14336 790 14338 791
rect 14334 785 14338 790
rect 14387 790 14388 808
rect 14494 799 14506 803
rect 14516 799 14528 803
rect 14538 796 14539 799
rect 14569 796 14570 805
rect 14620 799 14621 808
rect 14629 805 14635 811
rect 14687 808 14693 811
rect 14742 808 14758 824
rect 15331 819 15332 1015
rect 15521 819 15522 1015
rect 15607 819 15608 1015
rect 15880 819 15881 1015
rect 16078 820 16079 1016
rect 16470 1014 16474 1019
rect 17108 1014 17115 1019
rect 17195 1018 17204 1027
rect 17260 1024 17356 1027
rect 17697 1023 17805 1037
rect 17555 1015 17571 1022
rect 17573 1015 17589 1022
rect 17115 1007 17127 1014
rect 17545 1013 17557 1015
rect 17567 1013 17579 1015
rect 17585 1013 17589 1015
rect 17773 1013 17789 1022
rect 17805 1021 17823 1023
rect 17824 1017 17831 1020
rect 17831 1013 17837 1017
rect 18477 1015 18478 1026
rect 18667 1015 18668 1026
rect 18753 1015 18754 1026
rect 19026 1015 19027 1026
rect 19224 1016 19225 1027
rect 17545 1008 17589 1013
rect 17732 1008 17769 1009
rect 17837 1008 17840 1013
rect 17541 1006 17543 1008
rect 17545 1006 17677 1008
rect 16596 1005 16950 1006
rect 16576 1003 16594 1005
rect 17036 1003 17049 1005
rect 17128 1003 17131 1005
rect 17539 1003 17677 1006
rect 16520 1000 16576 1003
rect 16394 992 16406 1000
rect 16416 992 16428 1000
rect 16492 994 16576 1000
rect 17049 994 17059 1003
rect 16492 993 16520 994
rect 16390 989 16392 992
rect 16492 991 16511 993
rect 17060 991 17063 993
rect 16432 988 16436 989
rect 16382 977 16390 988
rect 16393 986 16428 988
rect 16391 977 16393 983
rect 16382 976 16391 977
rect 16390 972 16391 976
rect 16389 971 16390 972
rect 16387 966 16389 969
rect 16262 964 16327 965
rect 16254 956 16262 964
rect 16327 956 16331 964
rect 16253 950 16254 956
rect 16382 954 16390 966
rect 16394 956 16396 986
rect 16425 985 16428 986
rect 16427 979 16428 985
rect 16432 981 16440 988
rect 16436 980 16444 981
rect 16468 980 16469 990
rect 16492 980 16507 991
rect 16766 981 16803 983
rect 16444 979 16450 980
rect 16467 979 16468 980
rect 16492 979 16499 980
rect 16450 969 16512 979
rect 16520 972 16526 978
rect 16566 972 16572 978
rect 16766 977 16792 981
rect 16803 977 16808 981
rect 17063 980 17076 991
rect 17039 979 17053 980
rect 16760 972 16766 977
rect 16808 972 16817 977
rect 17021 972 17039 979
rect 17053 977 17060 979
rect 17131 977 17152 1003
rect 17533 996 17677 1003
rect 17693 1006 17794 1008
rect 17693 996 17805 1006
rect 17494 990 17555 996
rect 17459 987 17494 990
rect 17272 981 17459 987
rect 17545 986 17555 990
rect 17060 972 17075 977
rect 16514 969 16520 972
rect 16521 970 16578 972
rect 16817 971 16818 972
rect 16655 970 16658 971
rect 16676 970 16679 971
rect 16758 970 16759 971
rect 16818 970 16821 971
rect 16521 969 16529 970
rect 16492 968 16529 969
rect 16394 954 16428 956
rect 16383 951 16385 954
rect 16379 939 16383 950
rect 16394 942 16406 950
rect 16419 945 16428 954
rect 16466 952 16467 955
rect 16492 951 16497 968
rect 16514 966 16529 968
rect 16572 966 16578 970
rect 16651 967 16655 970
rect 16679 967 16684 970
rect 16821 968 16822 970
rect 17013 969 17021 972
rect 17050 971 17075 972
rect 17084 971 17088 972
rect 17046 970 17050 971
rect 17060 970 17097 971
rect 16822 967 16825 968
rect 16520 964 16529 966
rect 16520 951 16525 964
rect 16573 955 16592 958
rect 16627 955 16651 967
rect 16684 959 16702 967
rect 16757 959 16758 967
rect 16429 948 16439 950
rect 16439 947 16442 948
rect 16444 945 16453 947
rect 16417 942 16419 945
rect 16453 943 16464 945
rect 16465 943 16466 951
rect 16492 943 16498 951
rect 16416 939 16417 942
rect 16464 938 16498 943
rect 16330 924 16331 938
rect 16280 915 16289 924
rect 16327 920 16336 924
rect 16327 915 16341 920
rect 16271 912 16280 915
rect 16271 911 16274 912
rect 16264 908 16273 911
rect 16252 907 16273 908
rect 16252 905 16270 907
rect 16310 905 16316 911
rect 16330 906 16345 915
rect 16370 908 16379 937
rect 16252 900 16264 905
rect 16248 898 16251 900
rect 16252 899 16253 900
rect 16258 899 16264 900
rect 16316 899 16322 905
rect 16329 904 16341 906
rect 16368 904 16370 908
rect 16408 907 16416 938
rect 16465 926 16466 938
rect 16492 935 16520 938
rect 16492 931 16522 935
rect 16524 931 16525 951
rect 16592 946 16654 955
rect 16702 952 16710 959
rect 16756 951 16757 958
rect 16825 954 16829 967
rect 17005 966 17013 969
rect 17043 968 17046 970
rect 17039 967 17043 968
rect 17034 965 17039 967
rect 17060 965 17075 970
rect 17084 969 17088 970
rect 17097 969 17098 970
rect 17154 969 17159 975
rect 17195 971 17204 980
rect 17260 978 17272 981
rect 17260 971 17269 978
rect 17539 972 17555 986
rect 17578 972 17579 996
rect 17584 991 17605 996
rect 17589 990 17605 991
rect 17722 989 17728 996
rect 17774 989 17780 996
rect 17794 990 17805 996
rect 17840 990 17849 1008
rect 17589 972 17605 988
rect 17722 985 17730 989
rect 17728 983 17730 985
rect 17638 974 17666 978
rect 17668 974 17679 978
rect 17088 965 17093 969
rect 17098 965 17100 968
rect 17159 965 17162 969
rect 17000 964 17004 965
rect 17075 964 17078 965
rect 17100 964 17101 965
rect 16996 962 17000 964
rect 16610 945 16620 946
rect 16642 945 16643 946
rect 16606 943 16610 945
rect 16654 943 16674 946
rect 16755 943 16756 950
rect 16828 943 16829 950
rect 16877 943 16883 949
rect 16923 948 16929 949
rect 16960 948 16996 962
rect 17080 959 17084 962
rect 17095 960 17099 963
rect 17204 962 17213 971
rect 17237 961 17240 963
rect 17251 962 17260 971
rect 17545 970 17579 972
rect 17588 971 17589 972
rect 17635 971 17638 974
rect 17584 970 17589 971
rect 17634 970 17635 971
rect 17545 968 17589 970
rect 17632 969 17634 970
rect 17541 965 17542 967
rect 17315 961 17324 963
rect 17232 959 17237 961
rect 16923 947 16960 948
rect 16923 943 16929 947
rect 17015 946 17021 952
rect 17061 946 17067 952
rect 17083 949 17084 959
rect 17230 958 17232 959
rect 17326 958 17332 961
rect 17101 955 17105 958
rect 17169 955 17171 958
rect 17105 946 17115 955
rect 16594 931 16602 943
rect 16606 941 16640 943
rect 16492 928 16553 931
rect 16492 917 16498 928
rect 16520 926 16553 928
rect 16514 925 16553 926
rect 16572 925 16578 926
rect 16514 921 16578 925
rect 16514 920 16600 921
rect 16492 915 16499 917
rect 16492 913 16501 915
rect 16520 914 16526 920
rect 16566 914 16572 920
rect 16575 917 16600 920
rect 16584 915 16600 917
rect 16589 913 16600 915
rect 16606 913 16608 941
rect 16637 939 16640 941
rect 16492 909 16507 913
rect 16594 909 16608 913
rect 16638 909 16640 939
rect 16644 931 16652 943
rect 16674 934 16737 943
rect 16871 938 16877 943
rect 16889 941 16925 943
rect 16889 939 16894 941
rect 16830 937 16877 938
rect 16891 937 16894 939
rect 16929 937 16935 943
rect 17009 940 17015 946
rect 17067 940 17073 946
rect 16830 936 16873 937
rect 16754 934 16755 936
rect 16776 934 16830 936
rect 16710 922 16725 934
rect 16737 933 16776 934
rect 16754 929 16755 933
rect 16886 929 16889 936
rect 17013 933 17015 934
rect 16407 904 16408 906
rect 16467 905 16468 909
rect 16473 903 16479 909
rect 16492 903 16511 909
rect 16519 903 16525 909
rect 16327 899 16329 903
rect 16367 899 16368 903
rect 16326 897 16327 899
rect 16366 897 16367 899
rect 16240 884 16248 896
rect 16252 894 16270 896
rect 16325 895 16326 896
rect 16405 895 16407 903
rect 16467 897 16473 903
rect 16492 897 16531 903
rect 16533 897 16545 905
rect 16606 904 16623 909
rect 16710 904 16725 920
rect 16752 906 16754 928
rect 16614 903 16615 904
rect 16623 903 16627 904
rect 16642 903 16644 904
rect 16604 901 16605 903
rect 16615 899 16621 903
rect 16627 900 16646 903
rect 16751 900 16763 905
rect 16773 900 16785 905
rect 16826 904 16828 928
rect 16877 904 16886 928
rect 17009 925 17013 933
rect 16922 904 16925 909
rect 16963 908 16998 910
rect 16958 907 16963 908
rect 16998 907 17006 908
rect 17009 907 17011 915
rect 17033 909 17034 929
rect 17081 928 17083 944
rect 17115 942 17120 946
rect 17171 942 17183 955
rect 17332 951 17345 958
rect 17555 956 17571 968
rect 17573 956 17589 968
rect 17628 965 17632 968
rect 17626 963 17628 965
rect 17624 961 17626 963
rect 17679 961 17692 974
rect 17728 967 17731 983
rect 17730 961 17731 967
rect 17734 967 17735 989
rect 17773 985 17780 989
rect 17801 987 17803 990
rect 17773 983 17774 985
rect 17794 984 17795 986
rect 17734 963 17736 967
rect 17767 963 17768 966
rect 17772 965 17774 983
rect 17803 981 17806 987
rect 17806 979 17807 981
rect 17808 975 17809 977
rect 17809 972 17810 975
rect 17849 973 17857 990
rect 17811 965 17814 969
rect 17734 961 17738 963
rect 17772 962 17773 965
rect 17814 963 17815 965
rect 17620 958 17623 961
rect 17692 959 17695 961
rect 17618 953 17620 958
rect 17695 957 17697 959
rect 17453 952 17490 953
rect 17617 952 17618 953
rect 17697 952 17699 957
rect 17725 955 17731 961
rect 17738 959 17744 961
rect 17745 957 17751 959
rect 17771 957 17777 961
rect 17815 960 17816 963
rect 17816 958 17817 960
rect 17751 956 17777 957
rect 17453 951 17478 952
rect 17490 951 17491 952
rect 17347 948 17351 951
rect 17418 948 17445 951
rect 17493 948 17500 951
rect 17545 949 17546 952
rect 17500 943 17511 948
rect 17546 945 17548 949
rect 17581 947 17582 952
rect 17616 951 17617 952
rect 17614 948 17616 951
rect 17511 942 17515 943
rect 17183 939 17184 942
rect 17515 939 17520 942
rect 17520 938 17522 939
rect 17078 917 17080 920
rect 17075 915 17077 916
rect 17072 913 17075 915
rect 17069 911 17072 913
rect 17067 910 17069 911
rect 16953 906 16958 907
rect 17006 906 17015 907
rect 16942 904 16953 906
rect 16876 900 16877 903
rect 16920 900 16922 903
rect 16930 901 16942 904
rect 17009 900 17011 906
rect 17033 904 17034 906
rect 17101 904 17117 920
rect 17125 915 17151 938
rect 17185 931 17191 938
rect 17522 937 17524 938
rect 17524 933 17540 937
rect 17540 932 17545 933
rect 17548 932 17556 944
rect 17195 920 17203 927
rect 17203 918 17210 920
rect 17210 915 17222 918
rect 17151 910 17157 915
rect 17222 914 17226 915
rect 17229 914 17230 929
rect 17545 927 17561 932
rect 17582 929 17586 945
rect 17612 943 17614 948
rect 17699 944 17702 951
rect 17719 949 17725 955
rect 17751 951 17795 956
rect 17817 955 17819 958
rect 17777 949 17783 951
rect 17819 948 17822 955
rect 17611 942 17612 943
rect 17822 942 17825 948
rect 17857 943 17858 973
rect 17965 951 17981 954
rect 17893 943 17916 951
rect 17981 943 17988 951
rect 17610 940 17611 942
rect 17609 939 17610 940
rect 17825 939 17826 942
rect 17608 937 17609 938
rect 17605 933 17608 937
rect 17603 932 17605 933
rect 17826 932 17827 938
rect 17855 932 17857 942
rect 17887 939 17893 943
rect 17988 939 17992 943
rect 17885 938 17887 939
rect 17992 938 17995 939
rect 17875 932 17885 938
rect 17992 936 17997 938
rect 17586 927 17587 928
rect 17600 927 17603 932
rect 17724 927 17725 929
rect 17556 923 17557 926
rect 17561 924 17598 927
rect 17288 921 17319 922
rect 17279 920 17288 921
rect 17319 920 17326 921
rect 17586 920 17587 924
rect 17250 917 17279 920
rect 17326 917 17341 920
rect 17248 916 17250 917
rect 17245 915 17248 916
rect 17341 915 17349 917
rect 17558 915 17559 917
rect 17587 915 17588 920
rect 17592 915 17601 924
rect 17639 915 17648 924
rect 17723 922 17724 927
rect 17722 920 17723 922
rect 17721 918 17722 920
rect 17720 916 17721 918
rect 17238 914 17245 915
rect 17349 914 17358 915
rect 17583 914 17592 915
rect 17226 911 17592 914
rect 17229 910 17230 911
rect 17232 910 17234 911
rect 17368 910 17376 911
rect 17157 909 17159 910
rect 17034 903 17035 904
rect 17098 903 17101 904
rect 17159 903 17167 909
rect 17228 908 17232 910
rect 17376 907 17389 910
rect 17389 906 17394 907
rect 17221 904 17226 906
rect 17394 904 17404 906
rect 17035 900 17038 903
rect 17088 900 17101 903
rect 16492 895 16547 897
rect 16621 895 16627 899
rect 16641 898 16642 900
rect 16240 862 16248 874
rect 16252 864 16254 894
rect 16324 893 16325 894
rect 16365 893 16366 894
rect 16492 893 16549 895
rect 16627 893 16628 895
rect 16640 894 16641 897
rect 16646 896 16815 900
rect 16874 897 16876 900
rect 16871 896 16877 897
rect 16917 896 16920 900
rect 16747 894 16749 896
rect 16751 895 16752 896
rect 16815 895 16877 896
rect 16319 889 16325 893
rect 16364 889 16365 893
rect 16404 889 16405 893
rect 16460 889 16467 893
rect 16492 892 16557 893
rect 16305 888 16325 889
rect 16305 878 16319 888
rect 16361 879 16364 889
rect 16402 878 16404 889
rect 16457 879 16460 889
rect 16292 868 16305 878
rect 16358 869 16361 878
rect 16401 875 16402 878
rect 16456 875 16457 878
rect 16399 868 16401 875
rect 16454 869 16456 875
rect 16289 866 16292 868
rect 16252 862 16255 864
rect 16286 862 16289 866
rect 16336 859 16345 868
rect 16357 866 16358 868
rect 16356 862 16357 866
rect 16251 857 16253 858
rect 16258 857 16264 859
rect 16252 853 16264 857
rect 16316 853 16322 859
rect 16328 857 16336 859
rect 16355 858 16356 862
rect 16397 859 16399 867
rect 16451 859 16454 868
rect 16469 864 16472 892
rect 16519 891 16545 892
rect 16543 861 16545 891
rect 16549 881 16557 892
rect 16628 879 16648 893
rect 16696 879 16710 894
rect 16739 881 16747 893
rect 16751 891 16785 893
rect 16604 876 16605 879
rect 16634 876 16635 879
rect 16648 877 16660 879
rect 16694 877 16696 879
rect 16648 875 16694 877
rect 16519 859 16545 861
rect 16549 859 16557 871
rect 16602 869 16603 871
rect 16631 868 16632 870
rect 16599 860 16601 866
rect 16628 860 16631 867
rect 16751 859 16753 891
rect 16783 873 16785 891
rect 16789 881 16797 893
rect 16871 891 16877 895
rect 16915 891 16917 895
rect 16929 891 16935 897
rect 17009 894 17015 900
rect 17038 896 17053 900
rect 17053 895 17054 896
rect 17067 895 17101 900
rect 17167 899 17173 903
rect 17217 901 17221 904
rect 16825 881 16826 889
rect 16869 881 16872 891
rect 16877 885 16883 891
rect 16909 881 16915 891
rect 16923 885 16929 891
rect 17012 883 17013 891
rect 17015 888 17021 894
rect 17054 893 17073 895
rect 16784 865 16785 872
rect 16819 870 16825 880
rect 16864 870 16869 881
rect 16813 868 16819 870
rect 16863 868 16864 870
rect 16903 869 16909 881
rect 17052 872 17055 892
rect 17061 888 17067 893
rect 17085 888 17101 895
rect 17173 894 17184 899
rect 17212 898 17216 900
rect 17209 897 17212 898
rect 17205 894 17209 897
rect 17229 895 17232 900
rect 17404 897 17439 904
rect 17485 902 17498 903
rect 17464 900 17482 902
rect 17503 900 17526 902
rect 17462 899 17474 900
rect 17526 899 17535 900
rect 17535 898 17536 899
rect 17560 898 17561 904
rect 17455 897 17462 898
rect 17184 886 17215 894
rect 17232 893 17234 895
rect 17234 891 17236 893
rect 17439 891 17462 897
rect 17536 894 17543 898
rect 17543 891 17549 894
rect 17561 891 17562 897
rect 17174 880 17215 886
rect 17236 886 17309 891
rect 17439 889 17461 891
rect 17236 881 17386 886
rect 17447 882 17455 889
rect 17461 887 17466 889
rect 17466 886 17468 887
rect 17549 886 17562 891
rect 17590 887 17593 903
rect 17648 901 17657 915
rect 17718 911 17719 914
rect 17745 909 17777 914
rect 17712 903 17716 906
rect 17719 903 17725 909
rect 17745 904 17783 909
rect 17814 904 17875 932
rect 17994 931 17997 936
rect 17993 922 17997 931
rect 17742 903 17783 904
rect 17812 903 17814 904
rect 17822 903 17823 904
rect 17699 901 17711 902
rect 17657 899 17661 901
rect 17679 900 17699 901
rect 17673 899 17679 900
rect 17699 895 17701 900
rect 17725 897 17731 903
rect 17759 899 17760 901
rect 17697 892 17699 895
rect 17696 891 17697 892
rect 17174 876 17191 880
rect 17215 876 17233 880
rect 17236 876 17256 881
rect 17308 876 17399 881
rect 17233 875 17399 876
rect 17440 875 17447 882
rect 17468 876 17492 886
rect 17549 882 17563 886
rect 17562 881 17565 882
rect 17562 878 17563 881
rect 17565 880 17566 881
rect 17492 875 17495 876
rect 17171 874 17173 875
rect 17232 874 17402 875
rect 17169 873 17171 874
rect 17230 873 17232 874
rect 17228 872 17230 873
rect 17233 872 17399 874
rect 17402 873 17410 874
rect 17410 872 17418 873
rect 17437 872 17440 875
rect 17495 874 17497 875
rect 17497 873 17500 874
rect 17500 872 17502 873
rect 17511 872 17523 878
rect 17566 875 17575 880
rect 17593 876 17595 886
rect 17684 882 17696 891
rect 17678 881 17684 882
rect 17650 880 17666 881
rect 17674 880 17678 881
rect 17743 880 17758 899
rect 17771 897 17777 903
rect 17808 901 17812 903
rect 17797 895 17808 901
rect 17821 899 17822 901
rect 17794 892 17797 895
rect 17793 891 17794 892
rect 17785 886 17793 891
rect 17622 875 17645 880
rect 17773 876 17805 886
rect 17818 880 17821 898
rect 17817 876 17818 880
rect 17853 878 17855 904
rect 17993 903 17994 922
rect 18008 915 18017 924
rect 18055 915 18064 924
rect 17999 906 18004 915
rect 18069 906 18073 915
rect 17974 881 17993 901
rect 16807 866 16813 868
rect 16902 867 16903 868
rect 16901 866 16902 867
rect 16806 865 16807 866
rect 16784 860 16806 865
rect 16860 862 16863 866
rect 16785 859 16806 860
rect 16857 859 16863 862
rect 16327 855 16336 857
rect 16252 850 16261 853
rect 16264 850 16270 853
rect 16315 852 16316 853
rect 16325 852 16336 855
rect 16272 851 16320 852
rect 16323 851 16325 852
rect 16272 850 16323 851
rect 16327 850 16336 852
rect 16262 847 16270 850
rect 16262 846 16264 847
rect 16264 842 16266 846
rect 16315 840 16316 850
rect 16351 845 16355 858
rect 16394 846 16397 858
rect 16447 846 16451 858
rect 16467 851 16473 857
rect 16496 856 16500 859
rect 16790 858 16791 859
rect 16473 845 16479 851
rect 16491 845 16496 856
rect 16525 851 16531 857
rect 16598 855 16599 858
rect 16627 855 16628 858
rect 16857 857 16860 859
rect 16859 856 16860 857
rect 16855 855 16859 856
rect 16519 845 16525 851
rect 16533 847 16545 855
rect 16749 853 16750 855
rect 16596 851 16597 853
rect 16347 841 16351 845
rect 16393 841 16394 845
rect 16445 842 16447 845
rect 16345 840 16347 841
rect 16489 840 16491 845
rect 16593 841 16596 850
rect 16623 841 16626 850
rect 16750 841 16752 849
rect 16791 842 16792 849
rect 16852 847 16859 855
rect 16849 842 16852 847
rect 16855 845 16859 847
rect 16889 845 16901 865
rect 17013 859 17015 872
rect 17166 871 17168 872
rect 17226 871 17228 872
rect 16849 841 16851 842
rect 16846 840 16849 841
rect 16853 840 16855 845
rect 16886 844 16893 845
rect 17048 844 17052 870
rect 17161 868 17166 871
rect 17221 869 17225 871
rect 17309 869 17533 872
rect 17575 871 17581 875
rect 17612 871 17622 875
rect 17736 872 17739 876
rect 17770 875 17805 876
rect 17581 869 17587 871
rect 17594 869 17622 871
rect 17218 867 17220 868
rect 17158 866 17160 867
rect 17216 866 17218 867
rect 17325 866 17533 869
rect 17587 868 17588 869
rect 17594 868 17612 869
rect 17588 867 17592 868
rect 17607 867 17610 868
rect 17148 860 17158 866
rect 17206 862 17216 866
rect 17325 863 17535 866
rect 17438 862 17447 863
rect 17521 862 17543 863
rect 17564 862 17565 867
rect 17728 863 17736 872
rect 17783 869 17784 874
rect 17903 873 17914 874
rect 17931 873 17942 874
rect 17903 872 17911 873
rect 17935 872 17942 873
rect 17447 860 17450 862
rect 17143 857 17148 860
rect 17134 852 17143 857
rect 17450 852 17465 860
rect 17521 854 17535 862
rect 17543 856 17576 862
rect 17724 857 17728 862
rect 17651 856 17663 857
rect 17576 855 17582 856
rect 17600 855 17622 856
rect 17582 854 17622 855
rect 17643 854 17663 856
rect 17132 851 17134 852
rect 17465 851 17467 852
rect 17129 850 17132 851
rect 17467 850 17469 851
rect 17094 849 17100 850
rect 17127 849 17129 850
rect 17076 844 17127 849
rect 17140 844 17146 850
rect 17190 845 17193 849
rect 17470 845 17478 849
rect 17521 846 17533 854
rect 17651 851 17683 854
rect 17652 847 17683 851
rect 17721 849 17723 856
rect 17721 847 17722 849
rect 16886 840 16890 844
rect 16267 836 16268 840
rect 16268 833 16269 836
rect 16315 832 16317 840
rect 16333 832 16345 840
rect 16392 838 16393 840
rect 16444 838 16445 840
rect 16391 832 16392 838
rect 16443 833 16444 838
rect 16486 832 16489 840
rect 16592 837 16593 840
rect 16591 833 16592 836
rect 16620 834 16622 840
rect 16792 837 16793 840
rect 16753 832 16757 837
rect 16844 832 16853 840
rect 16882 834 16890 840
rect 16882 832 16886 834
rect 16269 817 16277 832
rect 16315 825 16319 832
rect 16332 830 16333 832
rect 16485 830 16486 832
rect 16331 828 16332 830
rect 16390 828 16391 830
rect 16441 828 16442 830
rect 16330 825 16331 828
rect 16317 817 16319 825
rect 16389 824 16390 828
rect 16440 824 16441 827
rect 16483 824 16485 829
rect 16328 819 16330 824
rect 16388 819 16389 824
rect 16435 820 16440 824
rect 14685 805 14693 808
rect 14685 804 14687 805
rect 14688 800 14689 802
rect 14689 797 14691 800
rect 14446 790 14448 793
rect 14254 758 14270 763
rect 14319 773 14380 785
rect 14387 779 14400 790
rect 14386 774 14400 779
rect 14430 777 14448 790
rect 14539 789 14540 793
rect 14570 789 14571 795
rect 14430 774 14446 777
rect 14319 759 14384 773
rect 14350 758 14366 759
rect 14368 758 14384 759
rect 14411 758 14412 760
rect 14446 758 14462 774
rect 14540 767 14544 785
rect 14571 779 14572 788
rect 14620 787 14622 794
rect 14685 790 14686 794
rect 14691 791 14694 797
rect 14726 792 14742 808
rect 14776 802 14804 808
rect 14840 806 14860 816
rect 16277 813 16279 817
rect 16279 809 16281 812
rect 16319 811 16320 817
rect 16327 815 16328 819
rect 16387 815 16388 819
rect 16435 815 16439 820
rect 16481 819 16483 824
rect 16326 809 16327 814
rect 16385 809 16387 814
rect 16435 809 16437 815
rect 16478 814 16481 818
rect 16531 814 16547 824
rect 16549 814 16565 824
rect 16585 817 16591 832
rect 16474 809 16478 814
rect 16518 809 16525 814
rect 16570 808 16578 814
rect 16583 811 16585 817
rect 16613 811 16620 832
rect 16754 827 16758 832
rect 16793 827 16799 832
rect 16842 830 16844 832
rect 16881 830 16882 832
rect 16612 809 16613 811
rect 16627 808 16643 824
rect 16743 822 16809 827
rect 16835 824 16842 830
rect 16878 825 16881 830
rect 16884 828 16886 832
rect 17015 832 17017 844
rect 17027 840 17039 844
rect 17055 842 17076 844
rect 17046 841 17055 842
rect 17041 840 17048 841
rect 17027 836 17041 840
rect 16743 821 16799 822
rect 16734 814 16743 821
rect 16754 818 16758 821
rect 16732 811 16734 814
rect 16757 811 16758 817
rect 16793 811 16799 821
rect 16809 814 16813 821
rect 16827 819 16835 824
rect 16875 819 16878 824
rect 16827 818 16829 819
rect 16827 815 16828 818
rect 16873 817 16875 819
rect 16872 816 16873 817
rect 16813 811 16814 814
rect 16826 812 16827 813
rect 16872 812 16875 816
rect 16905 812 16917 815
rect 16815 811 16824 812
rect 16650 808 16669 809
rect 16675 808 16677 809
rect 16282 804 16283 806
rect 14770 794 14804 802
rect 16283 799 16285 803
rect 16320 799 16321 803
rect 16323 800 16326 808
rect 16383 800 16385 808
rect 16285 794 16287 798
rect 16323 794 16325 800
rect 16381 794 16383 798
rect 14766 791 14768 794
rect 14776 790 14804 794
rect 14622 781 14623 787
rect 14685 782 14702 790
rect 14572 766 14577 779
rect 14624 774 14632 780
rect 14686 776 14702 782
rect 14758 779 14766 790
rect 14755 778 14766 779
rect 14770 788 14804 790
rect 14686 774 14696 776
rect 14632 773 14634 774
rect 14544 760 14545 766
rect 14577 759 14579 766
rect 14634 765 14648 773
rect 14686 766 14687 774
rect 14702 768 14707 776
rect 14755 770 14764 778
rect 14683 765 14687 766
rect 14629 764 14662 765
rect 14683 764 14693 765
rect 14629 759 14635 764
rect 14179 756 14185 758
rect 14256 757 14270 758
rect 14382 757 14385 758
rect 14264 756 14317 757
rect 14097 754 14098 756
rect 14179 754 14188 756
rect 13861 738 13867 739
rect 13907 738 13913 744
rect 13947 738 13956 747
rect 13994 738 14003 747
rect 14086 746 14100 754
rect 14174 747 14188 754
rect 14259 750 14323 756
rect 14386 750 14401 756
rect 14408 754 14409 756
rect 14450 752 14451 753
rect 14174 746 14179 747
rect 14100 745 14103 746
rect 13613 734 13614 736
rect 13615 727 13618 733
rect 13687 731 13702 736
rect 13855 732 13861 738
rect 13913 733 13919 738
rect 13967 734 13979 738
rect 14020 734 14036 744
rect 14098 742 14099 745
rect 14103 742 14142 745
rect 14172 743 14179 746
rect 14265 745 14280 750
rect 14311 747 14320 750
rect 14265 744 14271 745
rect 14311 744 14317 747
rect 14099 740 14142 742
rect 14103 737 14142 740
rect 14165 739 14172 743
rect 14174 739 14179 743
rect 14320 742 14334 747
rect 14401 745 14414 750
rect 14450 747 14458 752
rect 14546 751 14547 756
rect 14580 750 14583 756
rect 14635 753 14641 759
rect 14646 758 14662 764
rect 14664 758 14680 764
rect 14687 759 14693 764
rect 14707 762 14710 768
rect 14746 761 14755 770
rect 14681 753 14687 759
rect 14712 756 14714 760
rect 14742 757 14743 758
rect 14400 742 14402 745
rect 14414 742 14420 745
rect 14451 744 14458 747
rect 14547 746 14548 750
rect 14583 744 14585 750
rect 14669 745 14672 747
rect 14460 742 14461 744
rect 14714 743 14722 756
rect 14743 754 14746 757
rect 14758 756 14766 768
rect 14770 758 14772 788
rect 14801 787 14804 788
rect 14808 779 14851 791
rect 16288 785 16291 793
rect 16322 790 16324 793
rect 16325 790 16339 794
rect 16322 786 16339 790
rect 16291 779 16294 785
rect 14802 776 14851 779
rect 14802 770 14811 776
rect 14822 774 14838 776
rect 14851 774 14872 776
rect 16294 775 16296 778
rect 14811 764 14820 770
rect 14814 763 14820 764
rect 14838 768 14872 774
rect 16296 771 16297 775
rect 16323 774 16339 786
rect 16373 790 16381 794
rect 16419 792 16435 808
rect 16469 801 16474 808
rect 16514 801 16518 808
rect 16570 807 16581 808
rect 16611 807 16627 808
rect 16677 807 16678 808
rect 16726 807 16732 810
rect 16799 809 16800 811
rect 16754 808 16756 809
rect 16814 808 16824 811
rect 16871 808 16872 812
rect 16905 808 16921 812
rect 16923 808 16939 824
rect 16941 808 16957 824
rect 17015 820 17023 832
rect 17027 831 17043 832
rect 17027 830 17037 831
rect 16959 808 16968 812
rect 17018 810 17019 811
rect 16743 807 16753 808
rect 16570 806 16582 807
rect 16577 804 16582 806
rect 16469 792 16472 801
rect 16373 774 16389 790
rect 16419 774 16435 790
rect 16469 787 16485 790
rect 16464 781 16485 787
rect 16505 787 16514 801
rect 16577 792 16581 804
rect 16610 803 16627 807
rect 16678 806 16681 807
rect 16609 799 16610 803
rect 16607 794 16609 798
rect 16611 792 16627 803
rect 16650 798 16662 806
rect 16681 803 16684 806
rect 16704 803 16743 807
rect 16800 803 16801 807
rect 16811 803 16826 808
rect 16905 807 16922 808
rect 16927 807 16939 808
rect 16665 799 16704 803
rect 16715 799 16721 803
rect 16726 799 16732 803
rect 16801 799 16802 803
rect 16505 785 16516 787
rect 16525 785 16537 791
rect 16577 785 16578 792
rect 16605 788 16607 792
rect 16494 783 16516 785
rect 16526 783 16537 785
rect 16576 783 16581 785
rect 16488 781 16493 783
rect 16458 775 16464 781
rect 16469 774 16485 781
rect 16503 779 16505 783
rect 16510 781 16516 783
rect 16537 781 16541 783
rect 16516 775 16522 781
rect 16525 778 16537 779
rect 16325 771 16329 774
rect 14815 759 14818 763
rect 14838 758 14854 768
rect 14872 762 14889 768
rect 14875 758 14881 762
rect 14889 760 14895 762
rect 14895 758 14899 760
rect 14921 758 14927 764
rect 14770 757 14785 758
rect 14770 756 14789 757
rect 14746 750 14751 754
rect 14786 752 14804 756
rect 14821 753 14827 756
rect 14869 753 14875 758
rect 14770 750 14804 752
rect 14827 751 14875 753
rect 14927 752 14933 758
rect 16297 754 16305 771
rect 16329 754 16336 771
rect 16339 758 16355 774
rect 16357 758 16373 774
rect 16435 772 16443 774
rect 16461 772 16469 774
rect 16535 772 16537 778
rect 16541 772 16549 779
rect 16574 778 16576 783
rect 16577 778 16581 783
rect 16574 774 16581 778
rect 16574 772 16576 774
rect 16435 758 16451 772
rect 16453 758 16469 772
rect 16516 757 16579 772
rect 16603 760 16605 786
rect 16611 774 16627 790
rect 16638 782 16646 794
rect 16650 793 16671 794
rect 16709 793 16715 799
rect 16650 792 16668 793
rect 16627 763 16631 767
rect 16638 763 16646 772
rect 16650 763 16652 792
rect 16803 788 16805 796
rect 16811 794 16833 803
rect 16811 792 16826 794
rect 16863 790 16871 806
rect 16901 804 16903 807
rect 16907 806 16921 807
rect 16905 803 16921 806
rect 16957 805 16973 808
rect 16955 803 16973 805
rect 16893 791 16901 803
rect 16903 801 16939 803
rect 16903 793 16923 801
rect 16936 800 16939 801
rect 16937 793 16939 800
rect 16943 799 16951 803
rect 16955 799 16977 803
rect 16957 794 16977 799
rect 17015 798 17023 810
rect 17027 800 17029 830
rect 17046 826 17048 840
rect 17088 838 17094 844
rect 17146 838 17152 844
rect 17185 841 17190 845
rect 17478 841 17483 845
rect 17477 832 17485 841
rect 17489 834 17491 839
rect 17521 834 17523 846
rect 17781 845 17783 865
rect 17815 863 17817 872
rect 17852 863 17853 872
rect 17903 871 17905 872
rect 17941 871 17942 872
rect 17974 868 17988 881
rect 17967 866 17980 868
rect 17967 865 17979 866
rect 18008 865 18013 866
rect 17814 857 17815 862
rect 17812 849 17813 855
rect 17533 844 17536 845
rect 17489 832 17523 834
rect 17527 840 17536 844
rect 17527 832 17535 840
rect 17536 832 17540 840
rect 17540 830 17541 832
rect 17061 826 17062 830
rect 17172 829 17175 830
rect 17148 827 17183 829
rect 17046 818 17047 826
rect 17144 825 17148 827
rect 17142 824 17144 825
rect 17062 812 17064 824
rect 17047 800 17050 811
rect 17115 808 17142 824
rect 17146 812 17150 817
rect 17156 812 17172 827
rect 17183 824 17208 827
rect 17151 811 17172 812
rect 17027 798 17061 800
rect 17047 795 17050 798
rect 16805 778 16808 788
rect 16808 769 16810 778
rect 16811 774 16826 790
rect 16863 774 16877 790
rect 16900 781 16901 788
rect 16810 765 16811 769
rect 16627 762 16652 763
rect 16681 762 16684 763
rect 16627 760 16684 762
rect 16627 758 16643 760
rect 16811 759 16812 763
rect 14751 749 14787 750
rect 14770 744 14782 749
rect 14837 744 14848 749
rect 16305 746 16308 754
rect 16336 748 16341 754
rect 16341 745 16345 748
rect 16535 745 16537 757
rect 16540 745 16574 757
rect 16579 756 16581 757
rect 16688 756 16715 759
rect 16812 757 16813 759
rect 16827 758 16843 772
rect 16845 758 16861 772
rect 16893 769 16901 781
rect 16905 774 16923 793
rect 16957 792 16973 794
rect 16957 774 16973 790
rect 17003 774 17018 790
rect 17020 775 17022 792
rect 17027 786 17039 794
rect 17049 786 17061 794
rect 17063 790 17064 808
rect 17150 805 17160 811
rect 17208 808 17349 824
rect 17411 808 17427 824
rect 17429 808 17445 824
rect 17489 820 17501 828
rect 17511 820 17523 828
rect 17541 826 17542 830
rect 17567 828 17569 845
rect 17489 810 17491 820
rect 17542 816 17545 824
rect 17569 819 17570 828
rect 17597 819 17600 845
rect 17639 833 17645 845
rect 17686 843 17688 844
rect 17811 843 17812 847
rect 17722 838 17723 843
rect 17689 827 17690 836
rect 17723 827 17724 836
rect 17779 825 17781 840
rect 17810 837 17811 843
rect 17808 827 17810 836
rect 17850 829 17852 862
rect 17963 855 17979 865
rect 18016 864 18020 868
rect 17900 845 17963 855
rect 18008 851 18016 864
rect 17891 844 17900 845
rect 17885 842 17891 844
rect 17883 840 17885 842
rect 17639 811 17645 823
rect 17807 821 17808 826
rect 17848 820 17850 827
rect 17864 825 17883 840
rect 17863 824 17864 825
rect 17691 817 17692 820
rect 17724 816 17725 820
rect 17692 811 17697 816
rect 17725 811 17726 816
rect 17778 811 17779 818
rect 17792 811 17798 817
rect 17806 816 17807 820
rect 17847 818 17848 820
rect 17855 818 17863 824
rect 17804 812 17806 816
rect 17838 811 17844 817
rect 17846 816 17855 818
rect 17845 811 17855 816
rect 17601 808 17602 810
rect 17693 808 17694 810
rect 17155 803 17160 805
rect 17280 803 17289 808
rect 17327 803 17336 808
rect 17067 802 17076 803
rect 17065 798 17073 802
rect 17076 799 17091 802
rect 17091 798 17094 799
rect 17088 792 17094 798
rect 17146 792 17152 798
rect 17160 794 17169 803
rect 17271 794 17280 803
rect 17336 794 17345 803
rect 17262 792 17269 793
rect 17094 790 17100 792
rect 16905 772 16939 774
rect 16952 772 16957 774
rect 17050 772 17053 786
rect 17063 774 17069 790
rect 17094 786 17115 790
rect 17140 786 17146 792
rect 17256 791 17262 792
rect 17313 791 17317 793
rect 17349 792 17365 808
rect 17395 792 17411 808
rect 17422 803 17428 808
rect 17422 802 17437 803
rect 17416 796 17422 802
rect 17445 798 17461 808
rect 17468 802 17474 808
rect 17421 791 17422 793
rect 17454 791 17459 798
rect 17474 796 17480 802
rect 17492 800 17493 808
rect 17254 790 17256 791
rect 17253 787 17254 790
rect 17318 789 17320 790
rect 17099 774 17115 786
rect 17166 778 17193 781
rect 17149 774 17166 778
rect 17193 774 17201 778
rect 16905 769 16957 772
rect 17018 769 17024 772
rect 17053 771 17057 772
rect 16905 757 16909 765
rect 16941 758 16957 769
rect 17019 762 17036 769
rect 17053 762 17063 771
rect 17019 758 17035 762
rect 17036 760 17041 762
rect 17045 760 17057 762
rect 17041 759 17057 760
rect 17037 758 17057 759
rect 17115 758 17131 774
rect 17201 772 17204 774
rect 17269 772 17275 778
rect 17278 772 17280 779
rect 17320 772 17321 778
rect 17349 774 17365 790
rect 17395 774 17411 790
rect 17413 779 17422 791
rect 17204 763 17224 772
rect 17253 767 17254 769
rect 17263 766 17269 772
rect 17321 766 17327 772
rect 17342 763 17349 774
rect 17224 762 17226 763
rect 17226 759 17232 762
rect 16581 751 16602 756
rect 16602 747 16618 751
rect 16650 748 16662 756
rect 16813 754 16814 756
rect 16709 747 16715 753
rect 16740 747 16795 753
rect 16814 750 16815 754
rect 16815 747 16817 748
rect 16824 747 16833 756
rect 16903 747 16909 756
rect 16961 747 16967 753
rect 16968 747 16977 756
rect 17022 751 17025 758
rect 14848 743 14850 744
rect 14334 739 14343 742
rect 14420 741 14422 742
rect 14722 741 14723 743
rect 16308 741 16310 745
rect 14165 738 14179 739
rect 14152 737 14165 738
rect 14172 735 14174 738
rect 14343 735 14354 739
rect 14397 737 14398 739
rect 14354 734 14357 735
rect 13963 733 14045 734
rect 13913 732 13979 733
rect 13956 731 13979 732
rect 13702 726 13714 731
rect 13956 729 13963 731
rect 13967 730 13979 731
rect 14045 729 14048 732
rect 14164 731 14171 734
rect 14357 731 14366 734
rect 14394 733 14396 736
rect 14366 729 14373 731
rect 14389 729 14393 731
rect 13952 728 13956 729
rect 13945 726 13952 728
rect 13982 727 13983 729
rect 14048 728 14050 729
rect 13404 721 13475 723
rect 13228 719 13243 720
rect 13405 719 13475 721
rect 13507 719 13511 725
rect 13618 723 13620 726
rect 13231 716 13243 719
rect 11554 706 11564 709
rect 11565 706 11577 715
rect 11600 714 11602 715
rect 11602 709 11642 714
rect 11664 709 11676 714
rect 13167 712 13172 716
rect 13244 714 13247 716
rect 13396 712 13404 719
rect 13406 717 13416 719
rect 13406 712 13410 717
rect 11642 707 11676 709
rect 11642 706 11690 707
rect 11712 706 11718 712
rect 11770 706 11776 712
rect 11139 698 11150 701
rect 11233 698 11241 701
rect 11261 700 11269 701
rect 10602 688 10603 692
rect 10565 676 10599 678
rect 10603 676 10611 688
rect 10698 686 10704 692
rect 10756 686 10762 692
rect 10788 688 10795 692
rect 10904 691 10910 697
rect 10950 691 10956 697
rect 10996 691 11139 698
rect 11211 691 11233 698
rect 11267 692 11269 700
rect 11270 693 11276 698
rect 11289 694 11301 701
rect 10891 688 10893 691
rect 10788 687 10800 688
rect 10704 680 10710 686
rect 10750 680 10756 686
rect 10788 685 10803 687
rect 10810 685 10822 688
rect 10890 687 10891 688
rect 10889 685 10890 687
rect 10898 685 10904 691
rect 10956 685 10962 691
rect 10963 689 10984 691
rect 11206 689 11211 691
rect 11200 687 11206 689
rect 11269 688 11270 692
rect 11278 689 11281 691
rect 10967 685 11002 687
rect 10788 680 10800 685
rect 10803 680 10825 685
rect 10887 683 10889 685
rect 10825 676 10838 680
rect 10838 675 10843 676
rect 10852 675 10902 683
rect 10955 682 10967 685
rect 10946 680 10955 682
rect 11007 680 11009 685
rect 11190 684 11198 687
rect 11270 686 11271 687
rect 11183 682 11190 684
rect 10945 676 10946 680
rect 11176 679 11183 682
rect 11271 680 11273 682
rect 11171 678 11176 679
rect 11165 676 11171 678
rect 11273 676 11275 680
rect 11287 678 11294 684
rect 11306 682 11364 701
rect 11391 692 11392 698
rect 11455 692 11456 701
rect 11460 693 11468 703
rect 11475 702 11479 705
rect 11540 702 11565 706
rect 11662 704 11675 706
rect 11463 691 11468 693
rect 11479 692 11490 702
rect 11306 678 11339 682
rect 10601 672 10603 675
rect 10843 674 10902 675
rect 10852 672 10902 674
rect 10308 656 10311 662
rect 10232 643 10296 649
rect 10306 648 10308 656
rect 10352 652 10369 672
rect 10392 666 10399 672
rect 10565 666 10577 672
rect 10587 666 10599 672
rect 10829 666 10852 672
rect 10399 664 10605 666
rect 10818 664 10829 666
rect 10238 637 10265 643
rect 10284 637 10290 643
rect 10300 642 10306 647
rect 10310 642 10319 644
rect 10369 643 10377 652
rect 10546 642 10547 660
rect 9228 623 9255 629
rect 10048 626 10051 630
rect 10241 626 10265 637
rect 10300 635 10319 642
rect 10378 639 10382 642
rect 10382 636 10387 639
rect 10387 635 10395 636
rect 10300 630 10315 635
rect 10395 631 10431 635
rect 10299 626 10315 630
rect 10431 628 10451 631
rect 10545 630 10547 642
rect 10605 654 10764 664
rect 10776 654 10818 664
rect 10942 663 10945 674
rect 11009 663 11012 676
rect 11160 674 11165 676
rect 11157 673 11160 674
rect 11152 672 11157 673
rect 11146 670 11152 672
rect 11275 670 11278 676
rect 11294 671 11302 678
rect 11339 671 11347 678
rect 11364 676 11370 682
rect 11393 679 11394 682
rect 11395 677 11396 687
rect 11447 681 11460 682
rect 11447 679 11456 681
rect 11490 679 11495 692
rect 11540 688 11589 702
rect 11614 698 11660 704
rect 11678 703 11680 706
rect 11690 704 11710 706
rect 11718 704 11737 706
rect 11661 700 11676 702
rect 11606 694 11614 698
rect 11540 687 11565 688
rect 11589 687 11595 688
rect 11597 687 11606 694
rect 11522 678 11540 687
rect 11589 686 11597 687
rect 11595 685 11599 686
rect 11585 677 11592 683
rect 11599 682 11607 685
rect 11607 681 11612 682
rect 11612 680 11617 681
rect 11618 678 11621 679
rect 11389 676 11410 677
rect 11447 676 11453 677
rect 11370 673 11374 676
rect 11127 668 11146 670
rect 11090 664 11127 668
rect 11013 663 11090 664
rect 10904 655 11090 663
rect 11278 660 11291 670
rect 11302 660 11324 671
rect 11347 663 11357 671
rect 11374 663 11378 673
rect 11389 671 11395 676
rect 11396 672 11410 676
rect 11436 671 11453 676
rect 11494 671 11495 676
rect 11505 671 11520 677
rect 11395 665 11401 671
rect 11441 665 11447 671
rect 11485 663 11505 671
rect 11576 669 11585 677
rect 11624 676 11629 678
rect 11630 674 11636 676
rect 10605 652 10776 654
rect 10904 653 11019 655
rect 10605 642 10607 652
rect 10904 651 11016 653
rect 10904 649 11009 651
rect 10904 648 10972 649
rect 10904 645 10956 648
rect 10898 644 10962 645
rect 10876 643 10962 644
rect 10876 642 10894 643
rect 10605 634 10611 642
rect 10870 639 10887 642
rect 10898 639 10962 643
rect 10995 641 11007 649
rect 11012 643 11016 651
rect 10852 636 10870 639
rect 10606 630 10611 634
rect 10833 633 10852 636
rect 10904 633 10910 639
rect 10936 636 10942 639
rect 10950 633 10956 639
rect 11014 636 11016 643
rect 11291 642 11337 660
rect 11357 652 11387 663
rect 11367 647 11401 652
rect 11421 647 11422 660
rect 11458 652 11485 663
rect 11494 660 11495 663
rect 11367 646 11438 647
rect 11446 646 11475 652
rect 11367 643 11475 646
rect 11373 642 11378 643
rect 11291 641 11339 642
rect 10818 631 10833 633
rect 10622 630 10662 631
rect 10816 630 10818 631
rect 10461 628 10622 630
rect 10662 628 10691 630
rect 10545 626 10548 628
rect 10604 626 10611 628
rect 9256 623 9283 624
rect 8640 621 8641 622
rect 8544 615 8561 621
rect 8636 616 8640 621
rect 10051 618 10059 626
rect 10119 618 10126 625
rect 10059 617 10119 618
rect 8633 615 8636 616
rect 8561 611 8633 615
rect 10283 610 10299 626
rect 10548 615 10554 626
rect 10601 618 10604 625
rect 10691 622 10752 628
rect 10762 622 10812 630
rect 11012 627 11014 636
rect 10593 615 10601 618
rect 10554 613 10595 615
rect 10936 613 10949 624
rect 10990 616 11012 627
rect 11291 626 11337 641
rect 11341 637 11344 639
rect 11344 636 11346 637
rect 11346 633 11353 636
rect 11373 634 11387 642
rect 11421 634 11422 643
rect 11493 637 11494 653
rect 11535 652 11576 669
rect 11630 668 11638 674
rect 11642 670 11644 672
rect 11674 670 11676 700
rect 11680 690 11688 702
rect 11718 700 11724 704
rect 11764 700 11770 706
rect 11788 693 11799 702
rect 13172 696 13193 712
rect 13237 710 13261 712
rect 13241 705 13261 710
rect 13396 707 13406 712
rect 13403 705 13406 707
rect 13193 695 13195 696
rect 11642 668 11676 670
rect 11680 668 11688 680
rect 11799 678 11802 692
rect 13199 689 13200 692
rect 13197 678 13204 687
rect 13241 680 13243 705
rect 13247 700 13255 705
rect 13261 699 13267 705
rect 13401 701 13403 705
rect 13395 699 13403 701
rect 13267 694 13273 699
rect 13395 695 13401 699
rect 13273 692 13276 694
rect 13209 678 13243 680
rect 13247 678 13255 690
rect 13276 688 13277 692
rect 13389 689 13395 695
rect 13399 692 13400 694
rect 13398 688 13399 691
rect 13408 689 13410 712
rect 13440 715 13495 719
rect 13440 701 13463 715
rect 13471 713 13495 715
rect 13515 713 13516 715
rect 13476 708 13495 713
rect 13516 708 13520 713
rect 13620 710 13627 723
rect 13714 722 13744 726
rect 13963 724 13979 726
rect 13714 714 13756 722
rect 13483 701 13495 708
rect 13520 706 13521 708
rect 13627 705 13630 710
rect 13708 709 13757 710
rect 13440 695 13447 701
rect 13440 693 13453 695
rect 13440 689 13442 693
rect 13447 689 13453 693
rect 13458 691 13467 700
rect 13486 696 13495 701
rect 13526 696 13529 701
rect 13489 691 13495 696
rect 13397 685 13398 687
rect 13441 685 13442 689
rect 13459 687 13476 691
rect 13492 689 13495 691
rect 13529 689 13535 696
rect 13630 695 13667 705
rect 13708 702 13722 709
rect 13738 708 13757 709
rect 13754 703 13757 708
rect 13707 699 13708 701
rect 13667 693 13673 695
rect 13705 694 13707 699
rect 13673 692 13678 693
rect 13704 692 13705 694
rect 13494 687 13495 689
rect 13460 686 13476 687
rect 13535 686 13537 689
rect 13678 688 13694 692
rect 13694 687 13696 688
rect 13277 680 13279 685
rect 13396 680 13397 685
rect 13462 682 13465 686
rect 13467 682 13476 686
rect 13468 680 13469 682
rect 11802 676 11803 678
rect 13204 676 13205 678
rect 13208 676 13209 678
rect 13395 676 13396 678
rect 13469 677 13470 680
rect 11638 664 11641 666
rect 11642 656 11654 664
rect 11664 656 11676 664
rect 11803 661 11806 676
rect 11520 646 11535 652
rect 11642 648 11651 656
rect 11805 648 11806 661
rect 13204 660 13208 676
rect 13244 674 13247 676
rect 13209 666 13221 674
rect 13231 666 13243 674
rect 13279 660 13283 676
rect 13203 654 13204 658
rect 13283 657 13284 660
rect 11511 643 11518 646
rect 11506 641 11511 643
rect 11497 637 11506 641
rect 11353 631 11359 633
rect 11371 630 11387 634
rect 11362 626 11387 630
rect 11421 626 11423 630
rect 11355 622 11380 626
rect 10950 613 10990 616
rect 10561 610 10577 613
rect 10579 610 10595 613
rect 11355 610 11371 622
rect 11380 619 11388 622
rect 11388 618 11397 619
rect 11423 615 11428 626
rect 11455 620 11497 637
rect 11452 619 11455 620
rect 11446 618 11452 619
rect 11484 618 11491 620
rect 11480 615 11484 618
rect 11428 611 11449 615
rect 11471 611 11480 615
rect 11621 606 11645 629
rect 11651 626 11690 648
rect 11690 621 11699 626
rect 11796 622 11805 643
rect 13203 630 13205 654
rect 13283 630 13284 654
rect 13395 649 13447 663
rect 13468 662 13470 675
rect 13497 672 13509 685
rect 13537 672 13549 686
rect 13699 685 13705 687
rect 13705 683 13713 685
rect 13710 681 13714 683
rect 13710 676 13717 681
rect 13754 678 13756 703
rect 13757 697 13758 702
rect 13760 698 13768 710
rect 13913 694 13941 695
rect 13977 694 13979 724
rect 13983 714 13991 726
rect 14050 712 14052 728
rect 14373 727 14379 729
rect 14386 727 14389 729
rect 14106 720 14112 726
rect 14164 720 14170 726
rect 14370 723 14390 727
rect 14422 723 14443 741
rect 14448 738 14459 740
rect 14370 721 14386 723
rect 14365 720 14370 721
rect 14390 720 14398 723
rect 14112 714 14118 720
rect 14158 714 14164 720
rect 14358 717 14365 720
rect 14398 719 14401 720
rect 14443 719 14448 723
rect 14353 716 14358 717
rect 14401 716 14407 719
rect 14448 716 14452 719
rect 14456 716 14458 738
rect 14459 737 14460 738
rect 14462 737 14470 740
rect 14460 734 14470 737
rect 14462 729 14470 734
rect 14549 733 14550 741
rect 14586 737 14589 741
rect 14550 729 14551 733
rect 14579 729 14591 737
rect 14601 729 14613 737
rect 14676 729 14689 741
rect 14462 728 14471 729
rect 14467 726 14471 728
rect 14462 716 14470 718
rect 14344 713 14353 716
rect 14339 711 14344 713
rect 13758 693 13759 694
rect 13933 692 13941 694
rect 13945 692 13979 694
rect 13983 692 13991 704
rect 14050 694 14052 710
rect 14323 706 14339 711
rect 14407 706 14418 716
rect 14452 707 14470 716
rect 14434 706 14470 707
rect 14471 706 14494 726
rect 14551 724 14558 729
rect 14575 727 14578 729
rect 14591 725 14592 729
rect 14598 725 14604 729
rect 14552 723 14558 724
rect 14567 723 14575 725
rect 14579 723 14625 725
rect 14546 717 14552 723
rect 14579 717 14581 723
rect 14604 717 14610 723
rect 14611 717 14625 723
rect 14550 713 14552 714
rect 14548 709 14550 713
rect 14307 701 14323 706
rect 14418 705 14425 706
rect 14463 705 14496 706
rect 14418 702 14426 705
rect 14400 701 14434 702
rect 14460 701 14521 705
rect 14611 702 14613 717
rect 14617 713 14632 717
rect 14620 705 14632 713
rect 14689 712 14708 729
rect 14723 715 14757 741
rect 14852 723 14875 741
rect 16345 740 16353 745
rect 16571 742 16572 745
rect 16618 742 16638 747
rect 16638 741 16643 742
rect 16715 741 16721 747
rect 16761 741 16767 747
rect 16537 740 16539 741
rect 16310 737 16312 740
rect 16353 737 16358 740
rect 16527 739 16537 740
rect 16516 738 16537 739
rect 16643 738 16647 741
rect 16768 738 16777 747
rect 16815 745 16824 747
rect 16815 742 16830 745
rect 16815 738 16824 742
rect 16830 740 16834 742
rect 16909 741 16921 747
rect 16955 741 16968 747
rect 17024 744 17025 751
rect 16834 739 16837 740
rect 16358 736 16360 737
rect 16525 736 16544 738
rect 16313 733 16314 736
rect 16360 733 16364 736
rect 16314 727 16317 732
rect 16364 731 16368 733
rect 16368 729 16371 731
rect 16458 729 16464 735
rect 16516 729 16522 735
rect 16525 733 16562 736
rect 16569 733 16570 736
rect 16536 729 16562 733
rect 16565 729 16569 731
rect 16371 726 16375 729
rect 16317 720 16321 726
rect 16375 720 16385 726
rect 16388 720 16400 724
rect 16464 723 16470 729
rect 16510 723 16516 729
rect 16562 723 16589 729
rect 16601 726 16602 730
rect 16647 725 16664 738
rect 16768 737 16769 738
rect 16837 736 16844 739
rect 16912 738 16921 741
rect 16959 738 16968 741
rect 17018 739 17025 744
rect 17053 742 17057 758
rect 17095 747 17104 756
rect 17160 747 17169 756
rect 17232 754 17243 759
rect 17336 758 17349 763
rect 17411 769 17420 774
rect 17421 769 17422 779
rect 17411 763 17422 769
rect 17425 763 17427 791
rect 17493 790 17495 791
rect 17491 785 17495 790
rect 17544 790 17545 808
rect 17651 799 17663 803
rect 17673 799 17685 803
rect 17695 796 17696 799
rect 17726 796 17727 805
rect 17777 799 17778 808
rect 17786 805 17792 811
rect 17844 808 17850 811
rect 17899 808 17915 824
rect 18488 819 18489 1015
rect 18678 819 18679 1015
rect 18764 819 18765 1015
rect 19037 819 19038 1015
rect 19235 820 19236 1016
rect 17842 805 17850 808
rect 17842 804 17844 805
rect 17845 800 17846 802
rect 17846 797 17848 800
rect 17603 790 17605 793
rect 17411 758 17427 763
rect 17476 773 17537 785
rect 17544 779 17557 790
rect 17543 774 17557 779
rect 17587 777 17605 790
rect 17696 789 17697 793
rect 17727 789 17728 795
rect 17587 774 17603 777
rect 17476 759 17541 773
rect 17507 758 17523 759
rect 17525 758 17541 759
rect 17568 758 17569 760
rect 17603 758 17619 774
rect 17697 767 17701 785
rect 17728 779 17729 788
rect 17777 787 17779 794
rect 17842 790 17843 794
rect 17848 791 17851 797
rect 17883 792 17899 808
rect 17933 802 17961 808
rect 17997 806 18017 816
rect 17927 794 17961 802
rect 17923 791 17925 794
rect 17933 790 17961 794
rect 17779 781 17780 787
rect 17842 782 17859 790
rect 17729 766 17734 779
rect 17781 774 17789 780
rect 17843 776 17859 782
rect 17915 779 17923 790
rect 17912 778 17923 779
rect 17927 788 17961 790
rect 17843 774 17853 776
rect 17789 773 17791 774
rect 17701 760 17702 766
rect 17734 759 17736 766
rect 17791 765 17805 773
rect 17843 766 17844 774
rect 17859 768 17864 776
rect 17912 770 17921 778
rect 17840 765 17844 766
rect 17786 764 17819 765
rect 17840 764 17850 765
rect 17786 759 17792 764
rect 17336 756 17342 758
rect 17413 757 17427 758
rect 17539 757 17542 758
rect 17421 756 17474 757
rect 17254 754 17255 756
rect 17336 754 17345 756
rect 17018 738 17024 739
rect 17064 738 17070 744
rect 17104 738 17113 747
rect 17151 738 17160 747
rect 17243 746 17257 754
rect 17331 747 17345 754
rect 17416 750 17480 756
rect 17543 750 17558 756
rect 17565 754 17566 756
rect 17607 752 17608 753
rect 17331 746 17336 747
rect 17257 745 17260 746
rect 16770 734 16771 736
rect 16772 727 16775 733
rect 16844 731 16859 736
rect 17012 732 17018 738
rect 17070 733 17076 738
rect 17124 734 17136 738
rect 17177 734 17193 744
rect 17255 742 17256 745
rect 17260 742 17294 745
rect 17329 743 17336 746
rect 17422 745 17437 750
rect 17468 747 17477 750
rect 17422 744 17428 745
rect 17468 744 17474 747
rect 17256 740 17294 742
rect 17260 738 17294 740
rect 17322 739 17329 743
rect 17331 739 17336 743
rect 17477 742 17491 747
rect 17558 745 17571 750
rect 17607 747 17615 752
rect 17703 751 17704 756
rect 17737 750 17740 756
rect 17792 753 17798 759
rect 17803 758 17819 764
rect 17821 758 17837 764
rect 17844 759 17850 764
rect 17864 762 17867 768
rect 17903 761 17912 770
rect 17838 753 17844 759
rect 17869 756 17871 760
rect 17899 757 17900 758
rect 17557 742 17559 745
rect 17571 742 17577 745
rect 17608 744 17615 747
rect 17704 746 17705 750
rect 17740 744 17742 750
rect 17826 745 17829 747
rect 17617 742 17618 744
rect 17871 743 17879 756
rect 17900 754 17903 757
rect 17915 756 17923 768
rect 17927 758 17929 788
rect 17958 787 17961 788
rect 17965 779 18008 791
rect 17959 776 18008 779
rect 17959 770 17968 776
rect 17979 774 17995 776
rect 18008 774 18029 776
rect 17968 764 17977 770
rect 17971 763 17977 764
rect 17995 768 18029 774
rect 17972 759 17975 763
rect 17995 758 18011 768
rect 18029 762 18046 768
rect 18032 758 18038 762
rect 18046 760 18052 762
rect 18052 758 18056 760
rect 18078 758 18084 764
rect 17927 757 17942 758
rect 17927 756 17946 757
rect 17903 750 17908 754
rect 17943 752 17961 756
rect 17978 753 17984 756
rect 18026 753 18032 758
rect 17927 750 17961 752
rect 17984 751 18032 753
rect 18084 752 18090 758
rect 17908 749 17944 750
rect 17927 744 17939 749
rect 17994 744 18005 749
rect 18005 743 18007 744
rect 17491 739 17500 742
rect 17577 741 17579 742
rect 17879 741 17880 743
rect 17322 738 17336 739
rect 17265 737 17269 738
rect 17294 737 17299 738
rect 17309 737 17322 738
rect 17329 735 17331 738
rect 17500 735 17511 739
rect 17554 737 17555 739
rect 17511 734 17514 735
rect 17120 733 17202 734
rect 17070 732 17136 733
rect 17113 731 17136 732
rect 16859 726 16871 731
rect 17113 729 17120 731
rect 17124 730 17136 731
rect 17202 729 17205 732
rect 17321 731 17328 734
rect 17514 731 17523 734
rect 17551 733 17553 736
rect 17523 729 17530 731
rect 17546 729 17550 731
rect 17109 728 17113 729
rect 17102 726 17109 728
rect 17139 727 17140 729
rect 17205 728 17207 729
rect 16561 722 16632 723
rect 16561 721 16564 722
rect 16385 719 16400 720
rect 16589 719 16632 722
rect 16664 719 16668 725
rect 16775 723 16777 726
rect 16388 716 16400 719
rect 14711 706 14721 709
rect 14722 706 14734 715
rect 14757 714 14759 715
rect 14759 709 14799 714
rect 14821 709 14833 714
rect 16324 712 16329 716
rect 16401 714 16404 716
rect 16553 712 16561 719
rect 16563 717 16573 719
rect 16563 712 16567 717
rect 14799 707 14833 709
rect 14799 706 14847 707
rect 14869 706 14875 712
rect 14927 706 14933 712
rect 14296 698 14307 701
rect 14390 698 14398 701
rect 14418 700 14426 701
rect 13759 688 13760 692
rect 13722 676 13756 678
rect 13760 676 13768 688
rect 13855 686 13861 692
rect 13913 686 13919 692
rect 13945 688 13952 692
rect 14061 691 14067 697
rect 14107 691 14113 697
rect 14153 691 14296 698
rect 14368 691 14390 698
rect 14424 692 14426 700
rect 14427 693 14433 698
rect 14446 694 14458 701
rect 14048 688 14050 691
rect 13945 687 13957 688
rect 13861 680 13867 686
rect 13907 680 13913 686
rect 13945 685 13960 687
rect 13967 685 13979 688
rect 14047 687 14048 688
rect 14046 685 14047 687
rect 14055 685 14061 691
rect 14113 685 14119 691
rect 14120 689 14141 691
rect 14363 689 14368 691
rect 14357 687 14363 689
rect 14426 688 14427 692
rect 14435 689 14438 691
rect 14124 685 14159 687
rect 13945 680 13957 685
rect 13960 680 13982 685
rect 14044 683 14046 685
rect 13982 676 13995 680
rect 13995 675 14000 676
rect 14009 675 14059 683
rect 14112 682 14124 685
rect 14103 680 14112 682
rect 14164 680 14166 685
rect 14347 684 14355 687
rect 14427 686 14428 687
rect 14340 682 14347 684
rect 14102 676 14103 680
rect 14333 679 14340 682
rect 14428 680 14430 682
rect 14328 678 14333 679
rect 14322 676 14328 678
rect 14430 676 14432 680
rect 14444 678 14451 684
rect 14463 682 14521 701
rect 14548 692 14549 698
rect 14612 692 14613 701
rect 14617 693 14625 703
rect 14632 702 14636 705
rect 14697 702 14722 706
rect 14819 704 14832 706
rect 14620 691 14625 693
rect 14636 692 14647 702
rect 14463 678 14496 682
rect 13758 672 13760 675
rect 14000 674 14059 675
rect 14009 672 14059 674
rect 13465 656 13468 662
rect 13389 643 13453 649
rect 13463 648 13465 656
rect 13509 652 13526 672
rect 13549 666 13556 672
rect 13722 666 13734 672
rect 13744 666 13756 672
rect 13986 666 14009 672
rect 13556 664 13762 666
rect 13975 664 13986 666
rect 13395 637 13422 643
rect 13441 637 13447 643
rect 13457 642 13463 647
rect 13467 642 13476 644
rect 13526 643 13534 652
rect 13703 642 13704 660
rect 12383 623 12410 629
rect 13205 626 13208 630
rect 13398 626 13422 637
rect 13457 635 13476 642
rect 13535 639 13539 642
rect 13539 636 13544 639
rect 13544 635 13552 636
rect 13457 630 13472 635
rect 13552 631 13588 635
rect 13456 626 13472 630
rect 13588 628 13608 631
rect 13702 630 13704 642
rect 13762 654 13921 664
rect 13933 654 13975 664
rect 14099 663 14102 674
rect 14166 663 14169 676
rect 14317 674 14322 676
rect 14314 673 14317 674
rect 14309 672 14314 673
rect 14303 670 14309 672
rect 14432 670 14435 676
rect 14451 671 14459 678
rect 14496 671 14504 678
rect 14521 676 14527 682
rect 14550 679 14551 682
rect 14552 677 14553 687
rect 14604 681 14617 682
rect 14604 679 14613 681
rect 14647 679 14652 692
rect 14697 688 14746 702
rect 14771 698 14817 704
rect 14835 703 14837 706
rect 14847 704 14867 706
rect 14875 704 14894 706
rect 14818 700 14833 702
rect 14763 694 14771 698
rect 14697 687 14722 688
rect 14746 687 14752 688
rect 14754 687 14763 694
rect 14679 678 14697 687
rect 14746 686 14754 687
rect 14752 685 14756 686
rect 14742 677 14749 683
rect 14756 682 14764 685
rect 14764 681 14769 682
rect 14769 680 14774 681
rect 14775 678 14778 679
rect 14546 676 14567 677
rect 14604 676 14610 677
rect 14527 673 14531 676
rect 14284 668 14303 670
rect 14247 664 14284 668
rect 14170 663 14247 664
rect 14061 655 14247 663
rect 14435 660 14448 670
rect 14459 660 14481 671
rect 14504 663 14514 671
rect 14531 663 14535 673
rect 14546 671 14552 676
rect 14553 672 14567 676
rect 14593 671 14610 676
rect 14651 671 14652 676
rect 14662 671 14677 677
rect 14552 665 14558 671
rect 14598 665 14604 671
rect 14642 663 14662 671
rect 14733 669 14742 677
rect 14781 676 14786 678
rect 14787 674 14793 676
rect 13762 652 13933 654
rect 14061 653 14176 655
rect 13762 642 13764 652
rect 14061 651 14173 653
rect 14061 649 14166 651
rect 14061 648 14129 649
rect 14061 645 14113 648
rect 14055 644 14119 645
rect 14033 642 14119 644
rect 13762 634 13768 642
rect 14027 639 14044 642
rect 14055 639 14119 642
rect 14152 641 14164 649
rect 14169 643 14173 651
rect 14009 636 14027 639
rect 13763 630 13768 634
rect 13990 633 14009 636
rect 14061 633 14067 639
rect 14093 636 14099 639
rect 14107 633 14113 639
rect 14171 636 14173 643
rect 14448 642 14494 660
rect 14514 652 14544 663
rect 14524 647 14558 652
rect 14578 647 14579 660
rect 14615 652 14642 663
rect 14651 660 14652 663
rect 14524 646 14595 647
rect 14603 646 14632 652
rect 14524 643 14632 646
rect 14530 642 14535 643
rect 14448 641 14496 642
rect 13975 631 13990 633
rect 13779 630 13819 631
rect 13973 630 13975 631
rect 13618 628 13779 630
rect 13819 628 13848 630
rect 13702 626 13705 628
rect 13761 626 13768 628
rect 12411 623 12438 624
rect 11795 621 11796 622
rect 11699 615 11716 621
rect 11791 616 11795 621
rect 13208 618 13216 626
rect 13276 618 13283 625
rect 13216 617 13276 618
rect 11788 615 11791 616
rect 11716 611 11788 615
rect 13440 610 13456 626
rect 13705 615 13711 626
rect 13758 618 13761 625
rect 13848 622 13909 628
rect 13919 622 13969 630
rect 14169 627 14171 636
rect 13750 615 13758 618
rect 13711 613 13752 615
rect 14093 613 14106 624
rect 14147 616 14169 627
rect 14448 626 14494 641
rect 14498 637 14501 639
rect 14501 636 14503 637
rect 14503 633 14510 636
rect 14530 634 14544 642
rect 14578 634 14579 643
rect 14650 637 14651 653
rect 14692 652 14733 669
rect 14787 668 14795 674
rect 14799 670 14801 672
rect 14831 670 14833 700
rect 14837 690 14845 702
rect 14875 700 14881 704
rect 14921 700 14927 706
rect 14945 693 14956 702
rect 16329 696 16350 712
rect 16394 710 16418 712
rect 16398 705 16418 710
rect 16553 707 16563 712
rect 16560 705 16563 707
rect 16350 695 16352 696
rect 14799 668 14833 670
rect 14837 668 14845 680
rect 14956 678 14959 692
rect 16356 689 16357 692
rect 16354 678 16361 687
rect 16398 680 16400 705
rect 16404 700 16412 705
rect 16418 699 16424 705
rect 16558 701 16560 705
rect 16552 699 16560 701
rect 16424 694 16430 699
rect 16552 695 16558 699
rect 16430 692 16433 694
rect 16366 678 16400 680
rect 16404 678 16412 690
rect 16433 688 16434 692
rect 16546 689 16552 695
rect 16556 692 16557 694
rect 16555 688 16556 691
rect 16565 689 16567 712
rect 16597 715 16652 719
rect 16597 701 16620 715
rect 16628 713 16652 715
rect 16672 713 16673 715
rect 16633 708 16652 713
rect 16673 708 16677 713
rect 16777 710 16784 723
rect 16871 722 16901 726
rect 17120 724 17136 726
rect 16871 714 16913 722
rect 16640 701 16652 708
rect 16677 706 16678 708
rect 16784 705 16787 710
rect 16865 709 16914 710
rect 16597 695 16604 701
rect 16597 693 16610 695
rect 16597 689 16599 693
rect 16604 689 16610 693
rect 16615 691 16624 700
rect 16643 696 16652 701
rect 16683 696 16686 701
rect 16646 691 16652 696
rect 16554 685 16555 687
rect 16598 685 16599 689
rect 16616 687 16633 691
rect 16649 689 16652 691
rect 16686 689 16692 696
rect 16787 695 16824 705
rect 16865 702 16879 709
rect 16895 708 16914 709
rect 16911 703 16914 708
rect 16864 699 16865 701
rect 16824 693 16830 695
rect 16862 694 16864 699
rect 16830 692 16835 693
rect 16861 692 16862 694
rect 16651 687 16652 689
rect 16617 686 16633 687
rect 16692 686 16694 689
rect 16835 688 16851 692
rect 16851 687 16853 688
rect 16434 680 16436 685
rect 16553 680 16554 685
rect 16619 682 16622 686
rect 16624 682 16633 686
rect 16625 680 16626 682
rect 14959 676 14960 678
rect 16361 676 16362 678
rect 16365 676 16366 678
rect 16552 676 16553 678
rect 16626 677 16627 680
rect 14795 664 14798 666
rect 14799 656 14811 664
rect 14821 656 14833 664
rect 14960 661 14963 676
rect 14677 646 14692 652
rect 14799 648 14808 656
rect 14962 648 14963 661
rect 16361 660 16365 676
rect 16401 674 16404 676
rect 16366 666 16378 674
rect 16388 666 16400 674
rect 16436 660 16440 676
rect 16360 654 16361 658
rect 16440 657 16441 660
rect 14663 641 14675 646
rect 14654 637 14663 641
rect 14510 631 14516 633
rect 14528 630 14544 634
rect 14519 626 14544 630
rect 14578 626 14580 630
rect 14512 622 14537 626
rect 14107 613 14147 616
rect 13718 610 13734 613
rect 13736 610 13752 613
rect 14512 610 14528 622
rect 14537 619 14545 622
rect 14545 618 14554 619
rect 14580 615 14585 626
rect 14612 620 14654 637
rect 14609 619 14612 620
rect 14603 618 14609 619
rect 14641 618 14648 620
rect 14637 615 14641 618
rect 14585 611 14606 615
rect 14628 611 14637 615
rect 14778 606 14802 629
rect 14808 626 14847 648
rect 14847 621 14856 626
rect 14953 622 14962 643
rect 16360 630 16362 654
rect 16440 630 16441 654
rect 16552 649 16604 663
rect 16625 662 16627 675
rect 16654 672 16666 685
rect 16694 672 16706 686
rect 16856 685 16862 687
rect 16862 683 16870 685
rect 16867 681 16871 683
rect 16867 676 16874 681
rect 16911 678 16913 703
rect 16914 697 16915 702
rect 16917 698 16925 710
rect 17070 694 17098 695
rect 17134 694 17136 724
rect 17140 714 17148 726
rect 17207 712 17209 728
rect 17530 727 17536 729
rect 17543 727 17546 729
rect 17263 720 17269 726
rect 17321 720 17327 726
rect 17527 723 17547 727
rect 17579 723 17600 741
rect 17605 738 17616 740
rect 17527 721 17543 723
rect 17522 720 17527 721
rect 17547 720 17555 723
rect 17269 714 17275 720
rect 17315 714 17321 720
rect 17515 717 17522 720
rect 17555 719 17558 720
rect 17600 719 17605 723
rect 17510 716 17515 717
rect 17558 716 17564 719
rect 17605 716 17609 719
rect 17613 716 17615 738
rect 17616 737 17617 738
rect 17619 737 17627 740
rect 17617 734 17627 737
rect 17619 729 17627 734
rect 17706 733 17707 741
rect 17743 737 17746 741
rect 17707 729 17708 733
rect 17736 729 17748 737
rect 17758 729 17770 737
rect 17833 729 17846 741
rect 17619 728 17628 729
rect 17624 726 17628 728
rect 17619 716 17627 718
rect 17501 713 17510 716
rect 17496 711 17501 713
rect 16915 693 16916 694
rect 17090 692 17098 694
rect 17102 692 17136 694
rect 17140 692 17148 704
rect 17207 694 17209 710
rect 17480 706 17496 711
rect 17564 706 17575 716
rect 17609 707 17627 716
rect 17591 706 17627 707
rect 17628 706 17651 726
rect 17708 724 17715 729
rect 17732 727 17735 729
rect 17748 725 17749 729
rect 17755 725 17761 729
rect 17709 723 17715 724
rect 17724 723 17732 725
rect 17736 723 17782 725
rect 17703 717 17709 723
rect 17736 717 17738 723
rect 17761 717 17767 723
rect 17768 717 17782 723
rect 17707 713 17709 714
rect 17705 709 17707 713
rect 17464 701 17480 706
rect 17575 705 17582 706
rect 17620 705 17653 706
rect 17575 702 17583 705
rect 17557 701 17591 702
rect 17617 701 17678 705
rect 17768 702 17770 717
rect 17774 713 17789 717
rect 17777 705 17789 713
rect 17846 712 17865 729
rect 17880 715 17914 741
rect 18009 723 18032 741
rect 17868 706 17878 709
rect 17879 706 17891 715
rect 17914 714 17916 715
rect 17916 709 17956 714
rect 17978 709 17990 714
rect 17956 707 17990 709
rect 17956 706 18004 707
rect 18026 706 18032 712
rect 18084 706 18090 712
rect 17453 698 17464 701
rect 17547 698 17555 701
rect 17575 700 17583 701
rect 16916 688 16917 692
rect 16879 676 16913 678
rect 16917 676 16925 688
rect 17012 686 17018 692
rect 17070 686 17076 692
rect 17102 688 17109 692
rect 17218 691 17224 697
rect 17264 691 17270 697
rect 17310 691 17453 698
rect 17525 691 17547 698
rect 17581 692 17583 700
rect 17584 693 17590 698
rect 17603 694 17615 701
rect 17205 688 17207 691
rect 17102 687 17114 688
rect 17018 680 17024 686
rect 17064 680 17070 686
rect 17102 685 17117 687
rect 17124 685 17136 688
rect 17204 687 17205 688
rect 17203 685 17204 687
rect 17212 685 17218 691
rect 17270 685 17276 691
rect 17277 689 17298 691
rect 17520 689 17525 691
rect 17514 687 17520 689
rect 17583 688 17584 692
rect 17592 689 17595 691
rect 17281 685 17316 687
rect 17102 680 17114 685
rect 17117 680 17139 685
rect 17201 683 17203 685
rect 17139 676 17152 680
rect 17152 675 17157 676
rect 17166 675 17216 683
rect 17269 682 17281 685
rect 17260 680 17269 682
rect 17321 680 17323 685
rect 17504 684 17512 687
rect 17584 686 17585 687
rect 17497 682 17504 684
rect 17259 676 17260 680
rect 17490 679 17497 682
rect 17585 680 17587 682
rect 17485 678 17490 679
rect 17479 676 17485 678
rect 17587 676 17589 680
rect 17601 678 17608 684
rect 17620 682 17678 701
rect 17705 692 17706 698
rect 17769 692 17770 701
rect 17774 693 17782 703
rect 17789 702 17793 705
rect 17854 702 17879 706
rect 17976 704 17989 706
rect 17777 691 17782 693
rect 17793 692 17804 702
rect 17620 678 17653 682
rect 16915 672 16917 675
rect 17157 674 17216 675
rect 17166 672 17216 674
rect 16622 656 16625 662
rect 16546 643 16610 649
rect 16620 648 16622 656
rect 16666 652 16683 672
rect 16706 666 16713 672
rect 16879 666 16891 672
rect 16901 666 16913 672
rect 17143 666 17166 672
rect 16713 664 16919 666
rect 17132 664 17143 666
rect 16552 637 16579 643
rect 16598 637 16604 643
rect 16614 642 16620 647
rect 16624 642 16633 644
rect 16683 643 16691 652
rect 16860 642 16861 660
rect 15540 623 15567 629
rect 16362 626 16365 630
rect 16555 626 16579 637
rect 16614 635 16633 642
rect 16692 639 16696 642
rect 16696 636 16701 639
rect 16701 635 16709 636
rect 16614 630 16629 635
rect 16709 631 16745 635
rect 16613 626 16629 630
rect 16745 628 16765 631
rect 16859 630 16861 642
rect 16919 654 17078 664
rect 17090 654 17132 664
rect 17256 663 17259 674
rect 17323 663 17326 676
rect 17474 674 17479 676
rect 17471 673 17474 674
rect 17466 672 17471 673
rect 17460 670 17466 672
rect 17589 670 17592 676
rect 17608 671 17616 678
rect 17653 671 17661 678
rect 17678 676 17684 682
rect 17707 679 17708 682
rect 17709 677 17710 687
rect 17761 681 17774 682
rect 17761 679 17770 681
rect 17804 679 17809 692
rect 17854 688 17903 702
rect 17928 698 17974 704
rect 17992 703 17994 706
rect 18004 704 18024 706
rect 18032 704 18051 706
rect 17975 700 17990 702
rect 17920 694 17928 698
rect 17854 687 17879 688
rect 17903 687 17909 688
rect 17911 687 17920 694
rect 17836 678 17854 687
rect 17903 686 17911 687
rect 17909 685 17913 686
rect 17899 677 17906 683
rect 17913 682 17921 685
rect 17921 681 17926 682
rect 17926 680 17931 681
rect 17932 678 17935 679
rect 17703 676 17724 677
rect 17761 676 17767 677
rect 17684 673 17688 676
rect 17441 668 17460 670
rect 17404 664 17441 668
rect 17327 663 17404 664
rect 17218 655 17404 663
rect 17592 660 17605 670
rect 17616 660 17638 671
rect 17661 663 17671 671
rect 17688 663 17692 673
rect 17703 671 17709 676
rect 17710 672 17724 676
rect 17750 671 17767 676
rect 17808 671 17809 676
rect 17819 671 17834 677
rect 17709 665 17715 671
rect 17755 665 17761 671
rect 17799 663 17819 671
rect 17890 669 17899 677
rect 17938 676 17943 678
rect 17944 674 17950 676
rect 16919 652 17090 654
rect 17218 653 17333 655
rect 16919 642 16921 652
rect 17218 651 17330 653
rect 17218 649 17323 651
rect 17218 648 17286 649
rect 17218 645 17270 648
rect 17212 644 17276 645
rect 17190 642 17276 644
rect 16919 634 16925 642
rect 17184 639 17201 642
rect 17212 639 17276 642
rect 17309 641 17321 649
rect 17326 643 17330 651
rect 17166 636 17184 639
rect 16920 630 16925 634
rect 17147 633 17166 636
rect 17218 633 17224 639
rect 17250 636 17256 639
rect 17264 633 17270 639
rect 17328 636 17330 643
rect 17605 642 17651 660
rect 17671 652 17701 663
rect 17681 647 17715 652
rect 17735 647 17736 660
rect 17772 652 17799 663
rect 17808 660 17809 663
rect 17681 646 17752 647
rect 17760 646 17789 652
rect 17681 643 17789 646
rect 17687 642 17692 643
rect 17605 641 17653 642
rect 17132 631 17147 633
rect 16936 630 16976 631
rect 17130 630 17132 631
rect 16775 628 16936 630
rect 16976 628 17005 630
rect 16859 626 16862 628
rect 16918 626 16925 628
rect 15568 623 15595 624
rect 14952 621 14953 622
rect 14856 615 14873 621
rect 14948 616 14952 621
rect 16365 618 16373 626
rect 16433 618 16440 625
rect 16373 617 16433 618
rect 14945 615 14948 616
rect 14873 611 14945 615
rect 16597 610 16613 626
rect 16862 615 16868 626
rect 16915 618 16918 625
rect 17005 622 17066 628
rect 17076 622 17126 630
rect 17326 627 17328 636
rect 16907 615 16915 618
rect 16868 613 16909 615
rect 17250 613 17263 624
rect 17304 616 17326 627
rect 17605 626 17651 641
rect 17655 637 17658 639
rect 17658 636 17660 637
rect 17660 633 17667 636
rect 17687 634 17701 642
rect 17735 634 17736 643
rect 17807 637 17808 653
rect 17849 652 17890 669
rect 17944 668 17952 674
rect 17956 670 17958 672
rect 17988 670 17990 700
rect 17994 690 18002 702
rect 18032 700 18038 704
rect 18078 700 18084 706
rect 18102 693 18113 702
rect 17956 668 17990 670
rect 17994 668 18002 680
rect 18113 678 18116 692
rect 18116 676 18117 678
rect 17952 664 17955 666
rect 17956 656 17968 664
rect 17978 656 17990 664
rect 18117 661 18120 676
rect 17834 646 17849 652
rect 17956 648 17965 656
rect 18119 648 18120 661
rect 17820 641 17832 646
rect 17811 637 17820 641
rect 17667 631 17673 633
rect 17685 630 17701 634
rect 17676 626 17701 630
rect 17735 626 17737 630
rect 17669 622 17694 626
rect 17264 613 17304 616
rect 16875 610 16891 613
rect 16893 610 16909 613
rect 17669 610 17685 622
rect 17694 619 17702 622
rect 17702 618 17711 619
rect 17737 615 17742 626
rect 17769 620 17811 637
rect 17766 619 17769 620
rect 17760 618 17766 619
rect 17798 618 17805 620
rect 17794 615 17798 618
rect 17742 611 17763 615
rect 17785 611 17794 615
rect 17935 606 17959 629
rect 17965 626 18004 648
rect 18004 621 18013 626
rect 18110 622 18119 643
rect 18697 623 18724 629
rect 18725 623 18752 624
rect 18109 621 18110 622
rect 18013 615 18030 621
rect 18105 616 18109 621
rect 18102 615 18105 616
rect 18030 611 18102 615
rect 3666 557 3716 606
rect 3746 557 3812 606
rect 3842 557 3908 606
rect 3938 557 4004 606
rect 4034 557 4084 606
rect 4154 557 4204 606
rect 4234 557 4300 606
rect 4330 557 4396 606
rect 4426 557 4492 606
rect 4522 557 4572 606
rect 4642 557 4692 606
rect 4722 557 4788 606
rect 4818 557 4884 606
rect 4914 557 4980 606
rect 5010 557 5060 606
rect 5130 557 5180 606
rect 5210 557 5276 606
rect 5306 557 5372 606
rect 5402 557 5452 606
rect 6822 557 6872 606
rect 6902 557 6968 606
rect 6998 557 7064 606
rect 7094 557 7160 606
rect 7190 557 7240 606
rect 7310 557 7360 606
rect 7390 557 7456 606
rect 7486 557 7552 606
rect 7582 557 7648 606
rect 7678 557 7728 606
rect 7798 557 7848 606
rect 7878 557 7944 606
rect 7974 557 8040 606
rect 8070 557 8136 606
rect 8166 557 8216 606
rect 8286 557 8336 606
rect 8366 557 8432 606
rect 8462 557 8528 606
rect 8558 557 8608 606
rect 9977 557 10027 606
rect 10057 557 10123 606
rect 10153 557 10219 606
rect 10249 557 10315 606
rect 10345 557 10395 606
rect 10465 557 10515 606
rect 10545 557 10611 606
rect 10641 557 10707 606
rect 10737 557 10803 606
rect 10833 557 10883 606
rect 10953 557 11003 606
rect 11033 557 11099 606
rect 11129 557 11195 606
rect 11225 557 11291 606
rect 11321 557 11371 606
rect 11441 557 11491 606
rect 11521 557 11587 606
rect 11617 557 11683 606
rect 11713 557 11763 606
rect 13134 557 13184 606
rect 13214 557 13280 606
rect 13310 557 13376 606
rect 13406 557 13472 606
rect 13502 557 13552 606
rect 13622 557 13672 606
rect 13702 557 13768 606
rect 13798 557 13864 606
rect 13894 557 13960 606
rect 13990 557 14040 606
rect 14110 557 14160 606
rect 14190 557 14256 606
rect 14286 557 14352 606
rect 14382 557 14448 606
rect 14478 557 14528 606
rect 14598 557 14648 606
rect 14678 557 14744 606
rect 14774 557 14840 606
rect 14870 557 14920 606
rect 16291 557 16341 606
rect 16371 557 16437 606
rect 16467 557 16533 606
rect 16563 557 16629 606
rect 16659 557 16709 606
rect 16779 557 16829 606
rect 16859 557 16925 606
rect 16955 557 17021 606
rect 17051 557 17117 606
rect 17147 557 17197 606
rect 17267 557 17317 606
rect 17347 557 17413 606
rect 17443 557 17509 606
rect 17539 557 17605 606
rect 17635 557 17685 606
rect 17755 557 17805 606
rect 17835 557 17901 606
rect 17931 557 17997 606
rect 18027 557 18077 606
rect 6644 482 6645 488
rect 9800 482 9801 488
rect 12955 482 12956 488
rect 16112 482 16113 488
rect 19269 482 19270 488
rect 6610 442 6645 476
rect 6656 464 6657 476
rect 6656 442 6657 454
rect 9766 442 9801 476
rect 9812 464 9813 476
rect 9812 442 9813 454
rect 12921 442 12956 476
rect 12967 464 12968 476
rect 12967 442 12968 454
rect 16078 442 16113 476
rect 16124 464 16125 476
rect 16124 442 16125 454
rect 19235 442 19270 476
rect 19281 464 19282 476
rect 19281 442 19282 454
rect 5852 429 5853 440
rect 6042 429 6043 440
rect 6128 429 6129 440
rect 6401 429 6402 440
rect 6599 430 6600 441
rect 6633 430 6645 436
rect 5863 389 5864 429
rect 6053 389 6054 429
rect 6139 389 6140 429
rect 6412 389 6413 429
rect 6610 390 6611 430
rect 9008 429 9009 440
rect 9198 429 9199 440
rect 9284 429 9285 440
rect 9557 429 9558 440
rect 9755 430 9756 441
rect 9789 430 9801 436
rect 9019 389 9020 429
rect 9209 389 9210 429
rect 9295 389 9296 429
rect 9568 389 9569 429
rect 9766 390 9767 430
rect 12163 429 12164 440
rect 12353 429 12354 440
rect 12439 429 12440 440
rect 12712 429 12713 440
rect 12910 430 12911 441
rect 12944 430 12956 436
rect 12174 389 12175 429
rect 12364 389 12365 429
rect 12450 389 12451 429
rect 12723 389 12724 429
rect 12921 390 12922 430
rect 15320 429 15321 440
rect 15510 429 15511 440
rect 15596 429 15597 440
rect 15869 429 15870 440
rect 16067 430 16068 441
rect 16101 430 16113 436
rect 15331 389 15332 429
rect 15521 389 15522 429
rect 15607 389 15608 429
rect 15880 389 15881 429
rect 16078 390 16079 430
rect 18477 429 18478 440
rect 18667 429 18668 440
rect 18753 429 18754 440
rect 19026 429 19027 440
rect 19224 430 19225 441
rect 19258 430 19270 436
rect 18488 389 18489 429
rect 18678 389 18679 429
rect 18764 389 18765 429
rect 19037 389 19038 429
rect 19235 390 19236 430
<< nwell >>
rect 3009 1470 4458 1748
rect 4824 1646 4858 1680
rect 3000 840 4458 1470
rect 6097 1229 6131 1263
rect 12409 1229 12443 1263
rect 15566 1229 15600 1263
<< pdiff >>
rect 4824 1646 4858 1680
rect 15566 1229 15600 1263
<< locali >>
rect 4004 2492 19345 2493
rect 6 2172 19345 2492
rect 3406 1406 3440 1466
rect 0 1106 19340 1406
rect 0 0 19344 320
<< metal1 >>
rect 4004 2492 19345 2493
rect 6 2172 19345 2492
rect 19236 1982 19271 2010
rect 19230 1976 19300 1982
rect 3302 1862 3308 1920
rect 3366 1862 3372 1920
rect 19230 1918 19236 1976
rect 19294 1918 19300 1976
rect 19230 1912 19300 1918
rect 6609 1852 6679 1858
rect 5212 1842 5282 1848
rect 5212 1784 5218 1842
rect 5276 1784 5282 1842
rect 6609 1794 6615 1852
rect 6673 1794 6679 1852
rect 9764 1853 9835 1860
rect 6609 1788 6679 1794
rect 8374 1843 8444 1849
rect 5212 1778 5282 1784
rect 8374 1785 8380 1843
rect 8438 1785 8444 1843
rect 9764 1795 9771 1853
rect 9829 1795 9835 1853
rect 12911 1852 12981 1858
rect 9764 1789 9835 1795
rect 11530 1844 11600 1850
rect 8374 1779 8444 1785
rect 11530 1786 11536 1844
rect 11594 1786 11600 1844
rect 12911 1794 12917 1852
rect 12975 1794 12981 1852
rect 16068 1852 16138 1858
rect 12911 1788 12981 1794
rect 14676 1843 14746 1849
rect 11530 1780 11600 1786
rect 14676 1785 14682 1843
rect 14740 1785 14746 1843
rect 16068 1794 16074 1852
rect 16132 1794 16138 1852
rect 16068 1788 16138 1794
rect 17833 1843 17903 1849
rect 14676 1779 14746 1785
rect 17833 1785 17839 1843
rect 17897 1785 17903 1843
rect 17833 1779 17903 1785
rect 3227 1714 3233 1772
rect 3291 1714 3297 1772
rect 3034 1640 3092 1686
rect 4824 1646 4858 1680
rect 7980 1646 8014 1680
rect 11135 1646 11169 1680
rect 14292 1646 14326 1680
rect 17449 1646 17483 1680
rect 0 1106 19340 1406
rect 6610 441 6644 475
rect 9766 441 9800 475
rect 12921 441 12955 475
rect 16078 441 16112 475
rect 19235 441 19269 475
rect 0 0 19344 320
<< via1 >>
rect 3308 1862 3366 1920
rect 19236 1918 19294 1976
rect 5218 1784 5276 1842
rect 6615 1794 6673 1852
rect 8380 1785 8438 1843
rect 9771 1795 9829 1853
rect 11536 1786 11594 1844
rect 12917 1794 12975 1852
rect 14682 1785 14740 1843
rect 16074 1794 16132 1852
rect 17839 1785 17897 1843
rect 3233 1714 3291 1772
<< metal2 >>
rect 3246 2137 19270 2171
rect 3246 1778 3280 2137
rect 19236 1982 19270 2137
rect 19230 1976 19300 1982
rect 3308 1920 3366 1926
rect 19230 1918 19236 1976
rect 19294 1918 19300 1976
rect 19230 1912 19300 1918
rect 3366 1874 3589 1908
rect 3308 1856 3366 1862
rect 3555 1828 3589 1874
rect 6609 1852 6679 1858
rect 5212 1842 5282 1848
rect 5212 1828 5218 1842
rect 3555 1794 5218 1828
rect 5212 1784 5218 1794
rect 5276 1784 5282 1842
rect 6609 1794 6615 1852
rect 6673 1834 6679 1852
rect 9765 1853 9835 1859
rect 8374 1843 8444 1849
rect 8374 1834 8380 1843
rect 6673 1794 8380 1834
rect 6609 1788 6679 1794
rect 5212 1778 5282 1784
rect 8374 1785 8380 1794
rect 8438 1785 8444 1843
rect 9765 1795 9771 1853
rect 9829 1835 9835 1853
rect 12911 1852 12981 1858
rect 11530 1844 11600 1850
rect 11530 1835 11536 1844
rect 9829 1795 11536 1835
rect 9765 1789 9835 1795
rect 8374 1779 8444 1785
rect 11530 1786 11536 1795
rect 11594 1786 11600 1844
rect 12911 1794 12917 1852
rect 12975 1834 12981 1852
rect 16068 1852 16138 1858
rect 14676 1843 14746 1849
rect 14676 1834 14682 1843
rect 12975 1794 14682 1834
rect 12911 1788 12981 1794
rect 11530 1780 11600 1786
rect 14676 1785 14682 1794
rect 14740 1785 14746 1843
rect 16068 1794 16074 1852
rect 16132 1834 16138 1852
rect 17833 1843 17903 1849
rect 17833 1834 17839 1843
rect 16132 1794 17839 1834
rect 16068 1788 16138 1794
rect 14676 1779 14746 1785
rect 17833 1785 17839 1794
rect 17897 1785 17903 1843
rect 17833 1779 17903 1785
rect 3233 1772 3291 1778
rect 3233 1708 3291 1714
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_0
timestamp 1698882961
transform 1 0 3009 0 -1 2233
box -8 0 552 902
use sky130_osu_single_mpr2aa_8_b0r1  sky130_osu_single_mpr2aa_8_b0r1_0
timestamp 1707852425
transform 1 0 16174 0 1 0
box 0 0 3170 2492
use sky130_osu_single_mpr2aa_8_b0r1  sky130_osu_single_mpr2aa_8_b0r1_1
timestamp 1707852425
transform 1 0 3549 0 1 0
box 0 0 3170 2492
use sky130_osu_single_mpr2aa_8_b0r1  sky130_osu_single_mpr2aa_8_b0r1_2
timestamp 1707852425
transform 1 0 6705 0 1 0
box 0 0 3170 2492
use sky130_osu_single_mpr2aa_8_b0r1  sky130_osu_single_mpr2aa_8_b0r1_3
timestamp 1707852425
transform 1 0 9860 0 1 0
box 0 0 3170 2492
use sky130_osu_single_mpr2aa_8_b0r1  sky130_osu_single_mpr2aa_8_b0r1_4
timestamp 1707852425
transform 1 0 13017 0 1 0
box 0 0 3170 2492
<< labels >>
flabel metal1 s 3034 1640 3092 1686 0 FreeSans 100 0 0 0 start
port 13 nsew signal input
flabel metal1 s 4824 1646 4858 1680 0 FreeSans 100 0 0 0 s1
port 1 nsew signal input
flabel metal1 s 17449 1646 17483 1680 0 FreeSans 100 0 0 0 s5
port 5 nsew signal input
flabel metal1 s 14292 1646 14326 1680 0 FreeSans 100 0 0 0 s4
port 4 nsew signal input
flabel metal1 s 11135 1646 11169 1680 0 FreeSans 100 0 0 0 s3
port 3 nsew signal input
flabel metal1 s 7980 1646 8014 1680 0 FreeSans 100 0 0 0 s2
port 2 nsew signal input
flabel metal1 s 19235 441 19269 475 0 FreeSans 100 0 0 0 X5_Y1
port 10 nsew signal output
flabel metal1 s 9766 441 9800 475 0 FreeSans 100 0 0 0 X2_Y1
port 7 nsew signal output
flabel metal1 s 6610 441 6644 475 0 FreeSans 100 0 0 0 X1_Y1
port 6 nsew signal output
flabel metal1 s 12921 441 12955 475 0 FreeSans 100 0 0 0 X3_Y1
port 8 nsew signal output
flabel metal1 s 16078 441 16112 475 0 FreeSans 100 0 0 0 X4_Y1
port 9 nsew signal output
flabel metal1 s 3000 1106 19344 1406 0 FreeSans 100 0 0 0 vccd1
port 15 nsew power bidirectional
flabel metal1 s 6 2172 19345 2492 0 FreeSans 100 0 0 0 vssd1
port 16 nsew ground bidirectional
flabel metal1 s 0 1106 19340 1406 0 FreeSans 100 0 0 0 vccd1
port 15 nsew power bidirectional
flabel metal1 s 0 0 19344 320 0 FreeSans 100 0 0 0 vssd1
port 16 nsew ground bidirectional
<< end >>
