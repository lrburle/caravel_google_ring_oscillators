magic
tech sky130A
magscale 1 2
timestamp 1714073328
<< nwell >>
rect 3553 1747 4262 1748
rect 2997 1524 4262 1747
rect 6999 1634 7055 1690
rect 10316 1634 10372 1690
rect 13633 1634 13689 1690
rect 16949 1634 17005 1690
rect 2999 1446 4262 1524
rect 2999 1085 4263 1446
rect 5690 1086 7641 1406
rect 9007 1086 10958 1406
rect 12324 1086 14275 1406
rect 15641 1086 17592 1406
rect 18957 1086 20145 1406
rect 2997 861 4263 1085
rect 10075 985 10133 1043
rect 2997 743 4241 861
rect 6848 743 6880 745
rect 10162 742 10196 748
rect 13483 744 13513 747
rect 13481 742 13513 744
rect 16792 742 16862 760
<< ndiff >>
rect 6769 442 6804 476
rect 10086 442 10121 476
rect 13403 442 13438 476
rect 16720 442 16755 476
rect 20036 442 20071 476
rect 6772 441 6803 442
rect 10089 441 10120 442
rect 13406 441 13437 442
rect 16723 441 16754 442
rect 20039 441 20070 442
<< pdiff >>
rect 3047 1645 3081 1679
rect 3682 1634 3738 1690
rect 6999 1634 7055 1690
rect 10316 1634 10372 1690
rect 13633 1634 13689 1690
rect 16949 1634 17005 1690
<< locali >>
rect 11 2171 20145 2491
rect 3408 1405 3442 1470
rect 0 1085 4324 1405
rect 5690 1086 7641 1406
rect 9007 1086 10958 1406
rect 12324 1086 14275 1406
rect 15641 1086 17592 1406
rect 18957 1086 20145 1406
rect 6845 1085 6881 1086
rect 10161 1085 10200 1086
rect 13477 1085 13520 1086
rect 16793 1085 16834 1086
rect 0 0 20145 320
<< viali >>
rect 3047 1645 3081 1679
rect 6770 442 6804 476
rect 10087 442 10121 476
rect 13404 442 13438 476
rect 16721 442 16755 476
rect 20037 442 20071 476
<< metal1 >>
rect 11 2171 20145 2491
rect 20069 2007 20071 2012
rect 20030 1997 20083 2007
rect 20030 1975 20095 1997
rect 20030 1923 20037 1975
rect 20089 1923 20095 1975
rect 20030 1917 20095 1923
rect 3304 1861 3310 1917
rect 3366 1861 3372 1917
rect 6770 1847 6835 1854
rect 6770 1795 6777 1847
rect 6829 1795 6835 1847
rect 6770 1789 6835 1795
rect 10087 1847 10152 1854
rect 10087 1795 10094 1847
rect 10146 1795 10152 1847
rect 10087 1789 10152 1795
rect 13404 1847 13469 1854
rect 13404 1795 13411 1847
rect 13463 1795 13469 1847
rect 13404 1789 13469 1795
rect 16721 1847 16786 1854
rect 16721 1795 16728 1847
rect 16780 1795 16786 1847
rect 16721 1789 16786 1795
rect 3229 1713 3235 1769
rect 3291 1713 3297 1769
rect 6802 1759 6827 1789
rect 10117 1761 10144 1789
rect 13437 1761 13461 1789
rect 16753 1761 16778 1789
rect 3036 1679 3094 1685
rect 3036 1639 3041 1679
rect 3087 1639 3094 1679
rect 3743 1638 3763 1655
rect 7061 1638 7068 1653
rect 10377 1638 10404 1645
rect 13694 1638 13721 1645
rect 17008 1638 17020 1650
rect 0 1085 4324 1405
rect 5690 1086 7641 1406
rect 9007 1086 10958 1406
rect 12324 1086 14275 1406
rect 15641 1086 17592 1406
rect 18957 1086 20145 1406
rect 6845 1085 6881 1086
rect 10161 1085 10200 1086
rect 13477 1085 13520 1086
rect 16793 1085 16834 1086
rect 6769 441 6803 442
rect 10086 441 10120 442
rect 13403 441 13437 442
rect 16720 441 16754 442
rect 20036 441 20070 442
rect 0 0 20145 320
<< via1 >>
rect 20037 1923 20089 1975
rect 3310 1861 3366 1917
rect 6777 1795 6829 1847
rect 10094 1795 10146 1847
rect 13411 1795 13463 1847
rect 16728 1795 16780 1847
rect 3235 1713 3291 1769
rect 3682 1634 3738 1690
rect 6999 1634 7055 1690
rect 10316 1634 10372 1690
rect 13633 1634 13689 1690
rect 16949 1634 17005 1690
<< metal2 >>
rect 3553 2057 20071 2058
rect 3246 2024 20071 2057
rect 3246 2023 3553 2024
rect 3246 1775 3280 2023
rect 20037 1982 20071 2024
rect 20030 1975 20095 1982
rect 3310 1917 3366 1923
rect 3366 1868 3543 1902
rect 3310 1855 3366 1861
rect 3509 1829 3543 1868
rect 10582 1856 10656 1886
rect 13899 1856 13973 1886
rect 17289 1868 17290 1930
rect 20030 1923 20037 1975
rect 20089 1923 20095 1975
rect 20030 1917 20095 1923
rect 17216 1856 17290 1868
rect 6770 1847 6835 1854
rect 3509 1828 3573 1829
rect 3509 1794 4066 1828
rect 6770 1795 6777 1847
rect 6829 1829 6835 1847
rect 10087 1847 10152 1854
rect 6829 1828 6937 1829
rect 6829 1795 7383 1828
rect 6770 1789 6835 1795
rect 6937 1794 7383 1795
rect 10087 1795 10094 1847
rect 10146 1829 10152 1847
rect 13404 1847 13469 1854
rect 10146 1828 10210 1829
rect 10146 1795 10688 1828
rect 10087 1789 10152 1795
rect 10210 1794 10688 1795
rect 13404 1795 13411 1847
rect 13463 1829 13469 1847
rect 16721 1847 16786 1854
rect 13463 1828 13573 1829
rect 13463 1795 14005 1828
rect 13404 1789 13469 1795
rect 13573 1794 14005 1795
rect 16721 1795 16728 1847
rect 16780 1829 16786 1847
rect 16780 1828 16862 1829
rect 16780 1795 17322 1828
rect 16721 1789 16786 1795
rect 16862 1794 17322 1795
rect 10688 1782 10712 1783
rect 3235 1769 3291 1775
rect 3235 1707 3291 1713
<< via2 >>
rect 3682 1634 3738 1690
rect 6999 1634 7055 1690
rect 10316 1634 10372 1690
rect 13633 1634 13689 1690
rect 16949 1634 17005 1690
<< metal3 >>
rect 3676 1690 3744 2491
rect 6993 1690 7061 2491
rect 10310 1690 10378 2491
rect 13627 1690 13695 2491
rect 16943 1690 17011 2491
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_0
timestamp 1714057206
transform 1 0 3011 0 -1 2231
box -10 0 552 902
use sky130_osu_single_mpr2ca_8_b0r1  sky130_osu_single_mpr2ca_8_b0r1_0
timestamp 1714073328
transform 1 0 16827 0 1 0
box 0 0 3318 2491
use sky130_osu_single_mpr2ca_8_b0r1  sky130_osu_single_mpr2ca_8_b0r1_1
timestamp 1714073328
transform 1 0 3560 0 1 0
box 0 0 3318 2491
use sky130_osu_single_mpr2ca_8_b0r1  sky130_osu_single_mpr2ca_8_b0r1_2
timestamp 1714073328
transform 1 0 6877 0 1 0
box 0 0 3318 2491
use sky130_osu_single_mpr2ca_8_b0r1  sky130_osu_single_mpr2ca_8_b0r1_3
timestamp 1714073328
transform 1 0 10194 0 1 0
box 0 0 3318 2491
use sky130_osu_single_mpr2ca_8_b0r1  sky130_osu_single_mpr2ca_8_b0r1_4
timestamp 1714073328
transform 1 0 13511 0 1 0
box 0 0 3318 2491
<< labels >>
flabel metal1 s 3036 1639 3094 1685 0 FreeSans 100 0 0 0 start
port 13 nsew signal input
flabel metal1 s 0 1085 4324 1405 0 FreeSans 100 0 0 0 vccd1
port 15 nsew power bidirectional
flabel metal1 s 11 2171 20145 2491 0 FreeSans 100 0 0 0 vssd1
port 16 nsew ground bidirectional
flabel metal1 s 0 0 20145 320 0 FreeSans 100 0 0 0 vssd1
port 16 nsew ground bidirectional
flabel metal1 s 18957 1086 20145 1406 0 FreeSans 100 0 0 0 vccd1
port 15 nsew power bidirectional
flabel metal1 s 15641 1086 17592 1406 0 FreeSans 100 0 0 0 vccd1
port 15 nsew power bidirectional
flabel metal1 s 12324 1086 14275 1406 0 FreeSans 100 0 0 0 vccd1
port 15 nsew power bidirectional
flabel metal1 s 9007 1086 10958 1406 0 FreeSans 100 0 0 0 vccd1
port 15 nsew power bidirectional
flabel metal1 s 5690 1086 7641 1406 0 FreeSans 100 0 0 0 vccd1
port 15 nsew power bidirectional
flabel via2 s 3693 1645 3727 1679 0 FreeSans 100 0 0 0 s1
port 1 nw signal input
flabel via2 s 7010 1645 7044 1679 0 FreeSans 100 0 0 0 s2
port 2 nw signal input
flabel via2 s 10327 1645 10361 1679 0 FreeSans 100 0 0 0 s3
port 3 nw signal input
flabel via2 s 13644 1645 13678 1679 0 FreeSans 100 0 0 0 s4
port 4 nw signal input
flabel via2 s 16960 1645 16994 1679 0 FreeSans 100 0 0 0 s5
port 5 nw signal input
flabel viali s 16721 442 16755 476 0 FreeSans 100 0 0 0 X4_Y1
port 7 se signal output
flabel viali s 20037 442 20071 476 0 FreeSans 100 0 0 0 X5_Y1
port 6 se signal output
flabel viali s 10087 442 10121 476 0 FreeSans 100 0 0 0 X2_Y1
port 9 se signal output
flabel viali s 6770 442 6804 476 0 FreeSans 100 0 0 0 X1_Y1
port 10 se signal output
flabel viali s 13404 442 13438 476 0 FreeSans 100 0 0 0 X3_Y1
port 8 se signal output
<< end >>
