// Verilog for library /import/yukari1/brettcm/googleRO/char/liberate/VERILOG/b0r1_b0r2_MUX_IO_tt_1P8_25C.ccs created by Liberate 21.7.7.044.isr7 on Thu Nov  2 20:43:18 CDT 2023 for SDF version 2.1

// type:  
/// sta-blackbox
`timescale 1ns/10ps
`celldefine
module sky130_osu_ring_oscillator_mpr2aa_8_b0r1 (X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1, s1, s2, s3, s4, s5, start, vccd1, vssd1);
	output X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1;
	input s1, s2, s3, s4, s5, start;
	inout vccd1, vssd1;
endmodule
`endcelldefine

// type:  
/// sta-blackbox
`timescale 1ns/10ps
`celldefine
module sky130_osu_ring_oscillator_mpr2aa_8_b0r2 (X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1, s1, s2, s3, s4, s5, start, vccd1, vssd1);
	output X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1;
	input s1, s2, s3, s4, s5, start;
	inout vccd1, vssd1;
endmodule
`endcelldefine

/// sta-blackbox
`timescale 1ns/10ps
`celldefine
module sky130_osu_ring_oscillator_mpr2at_8_b0r1 (X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1, s1, s2, s3, s4, s5, start, vccd1, vssd1);
	output X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1;
	input s1, s2, s3, s4, s5, start;
	inout vccd1, vssd1;
endmodule
`endcelldefine

/// sta-blackbox
`timescale 1ns/10ps
`celldefine
module sky130_osu_ring_oscillator_mpr2at_8_b0r2 (X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1, s1, s2, s3, s4, s5, start, vccd1, vssd1);
	output X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1;
	input s1, s2, s3, s4, s5, start;
	inout vccd1, vssd1;
endmodule
`endcelldefine

/// sta-blackbox
`timescale 1ns/10ps
`celldefine
module sky130_osu_ring_oscillator_mpr2ca_8_b0r1 (X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1, s1, s2, s3, s4, s5, start, vccd1, vssd1);
	output X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1;
	input s1, s2, s3, s4, s5, start;
	inout vccd1, vssd1;
endmodule
`endcelldefine

/// sta-blackbox
`timescale 1ns/10ps
`celldefine
module sky130_osu_ring_oscillator_mpr2ca_8_b0r2 (X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1, s1, s2, s3, s4, s5, start, vccd1, vssd1);
	output X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1;
	input s1, s2, s3, s4, s5, start;
	inout vccd1, vssd1;
endmodule
`endcelldefine

/// sta-blackbox
`timescale 1ns/10ps
`celldefine
module sky130_osu_ring_oscillator_mpr2ct_8_b0r1 (X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1, s1, s2, s3, s4, s5, start, vccd1, vssd1);
	output X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1;
	input s1, s2, s3, s4, s5, start;
	inout vccd1, vssd1;
endmodule
`endcelldefine

/// sta-blackbox
`timescale 1ns/10ps
`celldefine
module sky130_osu_ring_oscillator_mpr2ct_8_b0r2 (X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1, s1, s2, s3, s4, s5, start, vccd1, vssd1);
	output X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1;
	input s1, s2, s3, s4, s5, start;
	inout vccd1, vssd1;
endmodule
`endcelldefine

/// sta-blackbox
`timescale 1ns/10ps
`celldefine
module sky130_osu_ring_oscillator_mpr2ea_8_b0r1 (X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1, s1, s2, s3, s4, s5, start, vccd1, vssd1);
	output X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1;
	input s1, s2, s3, s4, s5, start;
	inout vccd1, vssd1;
endmodule
`endcelldefine

/// sta-blackbox
`timescale 1ns/10ps
`celldefine
module sky130_osu_ring_oscillator_mpr2ea_8_b0r2 (X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1, s1, s2, s3, s4, s5, start, vccd1, vssd1);
	output X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1;
	input s1, s2, s3, s4, s5, start;
	inout vccd1, vssd1;
endmodule
`endcelldefine

/// sta-blackbox
`timescale 1ns/10ps
`celldefine
module sky130_osu_ring_oscillator_mpr2et_8_b0r1 (X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1, s1, s2, s3, s4, s5, start, vccd1, vssd1);
	output X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1;
	input s1, s2, s3, s4, s5, start;
	inout vccd1, vssd1;
endmodule
`endcelldefine

/// sta-blackbox
`timescale 1ns/10ps
`celldefine
module sky130_osu_ring_oscillator_mpr2et_8_b0r2 (X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1, s1, s2, s3, s4, s5, start, vccd1, vssd1);
	output X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1;
	input s1, s2, s3, s4, s5, start;
	inout vccd1, vssd1;
endmodule
`endcelldefine

/// sta-blackbox
`timescale 1ns/10ps
`celldefine
module sky130_osu_ring_oscillator_mpr2xa_8_b0r1 (X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1, s1, s2, s3, s4, s5, start, vccd1, vssd1);
	output X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1;
	input s1, s2, s3, s4, s5, start;
	inout vccd1, vssd1;
endmodule
`endcelldefine

/// sta-blackbox
`timescale 1ns/10ps
`celldefine
module sky130_osu_ring_oscillator_mpr2xa_8_b0r2 (X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1, s1, s2, s3, s4, s5, start, vccd1, vssd1);
	output X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1;
	input s1, s2, s3, s4, s5, start;
	inout vccd1, vssd1;
endmodule
`endcelldefine

/// sta-blackbox
`timescale 1ns/10ps
`celldefine
module sky130_osu_ring_oscillator_mpr2ya_8_b0r1 (X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1, s1, s2, s3, s4, s5, start, vccd1, vssd1);
	output X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1;
	input s1, s2, s3, s4, s5, start;
	inout vccd1, vssd1;
endmodule
`endcelldefine

/// sta-blackbox
`timescale 1ns/10ps
`celldefine
module sky130_osu_ring_oscillator_mpr2ya_8_b0r2 (X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1, s1, s2, s3, s4, s5, start, vccd1, vssd1);
	output X1_Y1, X2_Y1, X3_Y1, X4_Y1, X5_Y1;
	input s1, s2, s3, s4, s5, start;
	inout vccd1, vssd1;
endmodule
`endcelldefine
