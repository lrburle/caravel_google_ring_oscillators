magic
tech sky130A
magscale 1 2
timestamp 1699383188
<< viali >>
rect 295770 352665 295804 352699
rect 299087 352665 299121 352699
<< metal1 >>
rect 289722 352996 289728 353048
rect 289780 353036 289786 353048
rect 292040 353036 292068 353206
rect 289780 353008 292068 353036
rect 289780 352996 289786 353008
rect 295758 352699 295816 352705
rect 295758 352665 295770 352699
rect 295804 352696 295816 352699
rect 296530 352696 296536 352708
rect 295804 352668 296536 352696
rect 295804 352665 295816 352668
rect 295758 352659 295816 352665
rect 296530 352656 296536 352668
rect 296588 352656 296594 352708
rect 299075 352699 299133 352705
rect 299075 352665 299087 352699
rect 299121 352696 299133 352699
rect 299290 352696 299296 352708
rect 299121 352668 299296 352696
rect 299121 352665 299133 352668
rect 299075 352659 299133 352665
rect 299290 352656 299296 352668
rect 299348 352656 299354 352708
rect 302424 352226 302476 352232
rect 306282 352220 306288 352232
rect 305748 352192 306288 352220
rect 306282 352180 306288 352192
rect 306340 352180 306346 352232
rect 302424 352168 302476 352174
rect 309060 352152 309088 352200
rect 311158 352152 311164 352164
rect 309060 352124 311164 352152
rect 311158 352112 311164 352124
rect 311216 352112 311222 352164
rect 302418 349120 302424 349172
rect 302476 349160 302482 349172
rect 303522 349160 303528 349172
rect 302476 349132 303528 349160
rect 302476 349120 302482 349132
rect 303522 349120 303528 349132
rect 303580 349120 303586 349172
rect 296530 342184 296536 342236
rect 296588 342224 296594 342236
rect 517514 342224 517520 342236
rect 296588 342196 517520 342224
rect 296588 342184 296594 342196
rect 517514 342184 517520 342196
rect 517572 342184 517578 342236
rect 299290 340824 299296 340876
rect 299348 340864 299354 340876
rect 517514 340864 517520 340876
rect 299348 340836 517520 340864
rect 299348 340824 299354 340836
rect 517514 340824 517520 340836
rect 517572 340824 517578 340876
rect 303522 339396 303528 339448
rect 303580 339436 303586 339448
rect 517514 339436 517520 339448
rect 303580 339408 517520 339436
rect 303580 339396 303586 339408
rect 517514 339396 517520 339408
rect 517572 339396 517578 339448
rect 306282 338036 306288 338088
rect 306340 338076 306346 338088
rect 517514 338076 517520 338088
rect 306340 338048 517520 338076
rect 306340 338036 306346 338048
rect 517514 338036 517520 338048
rect 517572 338036 517578 338088
rect 311158 336676 311164 336728
rect 311216 336716 311222 336728
rect 517514 336716 517520 336728
rect 311216 336688 517520 336716
rect 311216 336676 311222 336688
rect 517514 336676 517520 336688
rect 517572 336676 517578 336728
rect 289722 206932 289728 206984
rect 289780 206972 289786 206984
rect 580166 206972 580172 206984
rect 289780 206944 580172 206972
rect 289780 206932 289786 206944
rect 580166 206932 580172 206944
rect 580224 206932 580230 206984
<< via1 >>
rect 289728 352996 289780 353048
rect 296536 352656 296588 352708
rect 299296 352656 299348 352708
rect 302424 352174 302476 352226
rect 306288 352180 306340 352232
rect 311164 352112 311216 352164
rect 302424 349120 302476 349172
rect 303528 349120 303580 349172
rect 296536 342184 296588 342236
rect 517520 342184 517572 342236
rect 299296 340824 299348 340876
rect 517520 340824 517572 340876
rect 303528 339396 303580 339448
rect 517520 339396 517572 339448
rect 306288 338036 306340 338088
rect 517520 338036 517572 338088
rect 311164 336676 311216 336728
rect 517520 336676 517572 336728
rect 289728 206932 289780 206984
rect 580172 206932 580224 206984
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 528650 404968 528706 404977
rect 528650 404903 528706 404912
rect 312542 354920 312598 354929
rect 312542 354855 312598 354864
rect 298243 353424 298299 353433
rect 298243 353359 298299 353368
rect 289728 353048 289780 353054
rect 289728 352990 289780 352996
rect 289740 206990 289768 352990
rect 294940 352594 294968 352852
rect 296536 352708 296588 352714
rect 296536 352650 296588 352656
rect 299296 352708 299348 352714
rect 299296 352650 299348 352656
rect 294940 352566 295012 352594
rect 294984 351937 295012 352566
rect 294970 351928 295026 351937
rect 294970 351863 295026 351872
rect 296548 342242 296576 352650
rect 296536 342236 296588 342242
rect 296536 342178 296588 342184
rect 299308 340882 299336 352650
rect 301574 352594 301602 352852
rect 304891 352594 304919 352852
rect 308184 352824 308193 352880
rect 308249 352824 308258 352880
rect 301574 352566 301636 352594
rect 304891 352566 304948 352594
rect 301608 351937 301636 352566
rect 302424 352226 302476 352232
rect 302424 352168 302476 352174
rect 301594 351928 301650 351937
rect 301594 351863 301650 351872
rect 302436 349178 302464 352168
rect 304920 351937 304948 352566
rect 306288 352232 306340 352238
rect 306288 352174 306340 352180
rect 304906 351928 304962 351937
rect 304906 351863 304962 351872
rect 302424 349172 302476 349178
rect 302424 349114 302476 349120
rect 303528 349172 303580 349178
rect 303528 349114 303580 349120
rect 299296 340876 299348 340882
rect 299296 340818 299348 340824
rect 303540 339454 303568 349114
rect 303528 339448 303580 339454
rect 303528 339390 303580 339396
rect 306300 338094 306328 352174
rect 311164 352164 311216 352170
rect 311164 352106 311216 352112
rect 306288 338088 306340 338094
rect 306288 338030 306340 338036
rect 311176 336734 311204 352106
rect 311164 336728 311216 336734
rect 311164 336670 311216 336676
rect 289728 206984 289780 206990
rect 289728 206926 289780 206932
rect 312556 46345 312584 354855
rect 526166 351928 526222 351937
rect 526166 351863 526222 351872
rect 523682 343768 523738 343777
rect 523682 343703 523738 343712
rect 517520 342236 517572 342242
rect 517520 342178 517572 342184
rect 517532 341057 517560 342178
rect 523696 341972 523724 343703
rect 526180 341972 526208 351863
rect 528664 341972 528692 404903
rect 530582 343768 530638 343777
rect 530582 343703 530638 343712
rect 520660 341414 521226 341442
rect 517518 341048 517574 341057
rect 517518 340983 517574 340992
rect 517520 340876 517572 340882
rect 517520 340818 517572 340824
rect 517532 339697 517560 340818
rect 517518 339688 517574 339697
rect 517518 339623 517574 339632
rect 517520 339448 517572 339454
rect 517520 339390 517572 339396
rect 517532 338337 517560 339390
rect 517518 338328 517574 338337
rect 517518 338263 517574 338272
rect 517520 338088 517572 338094
rect 517520 338030 517572 338036
rect 517532 336977 517560 338030
rect 517518 336968 517574 336977
rect 517518 336903 517574 336912
rect 517520 336728 517572 336734
rect 517520 336670 517572 336676
rect 517532 335617 517560 336670
rect 517518 335608 517574 335617
rect 517518 335543 517574 335552
rect 520660 245585 520688 341414
rect 530596 298761 530624 343703
rect 530582 298752 530638 298761
rect 530582 298687 530638 298696
rect 520646 245576 520702 245585
rect 520646 245511 520702 245520
rect 580172 206984 580224 206990
rect 580172 206926 580224 206932
rect 580184 205737 580212 206926
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 312542 46336 312598 46345
rect 312542 46271 312598 46280
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 528650 404912 528706 404968
rect 312542 354864 312598 354920
rect 298243 353368 298299 353424
rect 294970 351872 295026 351928
rect 308193 352824 308249 352880
rect 301594 351872 301650 351928
rect 304906 351872 304962 351928
rect 526166 351872 526222 351928
rect 523682 343712 523738 343768
rect 530582 343712 530638 343768
rect 517518 340992 517574 341048
rect 517518 339632 517574 339688
rect 517518 338272 517574 338328
rect 517518 336912 517574 336968
rect 517518 335552 517574 335608
rect 530582 298696 530638 298752
rect 520646 245520 520702 245576
rect 580170 205672 580226 205728
rect 312542 46280 312598 46336
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 528645 404970 528711 404973
rect 583520 404970 584960 405060
rect 528645 404968 584960 404970
rect 528645 404912 528650 404968
rect 528706 404912 584960 404968
rect 528645 404910 584960 404912
rect 528645 404907 528711 404910
rect 583520 404820 584960 404910
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 299238 354860 299244 354924
rect 299308 354922 299314 354924
rect 312537 354922 312603 354925
rect 299308 354920 312603 354922
rect 299308 354864 312542 354920
rect 312598 354864 312603 354920
rect 299308 354862 312603 354864
rect 299308 354860 299314 354862
rect 312537 354859 312603 354862
rect 298238 353426 298304 353429
rect 299238 353426 299244 353428
rect 298238 353424 299244 353426
rect 298238 353368 298243 353424
rect 298299 353368 299244 353424
rect 298238 353366 299244 353368
rect 298238 353363 298304 353366
rect 299238 353364 299244 353366
rect 299308 353364 299314 353428
rect 308188 352882 308254 352885
rect 308438 352882 308444 352884
rect 308188 352880 308444 352882
rect 308188 352824 308193 352880
rect 308249 352824 308444 352880
rect 308188 352822 308444 352824
rect 308188 352819 308254 352822
rect 308438 352820 308444 352822
rect 308508 352820 308514 352884
rect 294965 351932 295031 351933
rect 301589 351932 301655 351933
rect 294965 351928 295012 351932
rect 295076 351930 295082 351932
rect 294965 351872 294970 351928
rect 294965 351868 295012 351872
rect 295076 351870 295122 351930
rect 301589 351928 301636 351932
rect 301700 351930 301706 351932
rect 301589 351872 301594 351928
rect 295076 351868 295082 351870
rect 301589 351868 301636 351872
rect 301700 351870 301746 351930
rect 301700 351868 301706 351870
rect 304758 351868 304764 351932
rect 304828 351930 304834 351932
rect 304901 351930 304967 351933
rect 304828 351928 304967 351930
rect 304828 351872 304906 351928
rect 304962 351872 304967 351928
rect 304828 351870 304967 351872
rect 304828 351868 304834 351870
rect 294965 351867 295031 351868
rect 301589 351867 301655 351868
rect 304901 351867 304967 351870
rect 526161 351930 526227 351933
rect 583520 351930 584960 352020
rect 526161 351928 584960 351930
rect 526161 351872 526166 351928
rect 526222 351872 584960 351928
rect 526161 351870 584960 351872
rect 526161 351867 526227 351870
rect 583520 351780 584960 351870
rect -960 345252 480 345492
rect 523677 343770 523743 343773
rect 530577 343770 530643 343773
rect 523677 343768 530643 343770
rect 523677 343712 523682 343768
rect 523738 343712 530582 343768
rect 530638 343712 530643 343768
rect 523677 343710 530643 343712
rect 523677 343707 523743 343710
rect 530577 343707 530643 343710
rect 517513 341050 517579 341053
rect 517513 341048 520076 341050
rect 517513 340992 517518 341048
rect 517574 340992 520076 341048
rect 517513 340990 520076 340992
rect 517513 340987 517579 340990
rect 517513 339690 517579 339693
rect 517513 339688 520076 339690
rect 517513 339632 517518 339688
rect 517574 339632 520076 339688
rect 517513 339630 520076 339632
rect 517513 339627 517579 339630
rect 583520 338452 584960 338692
rect 517513 338330 517579 338333
rect 517513 338328 520076 338330
rect 517513 338272 517518 338328
rect 517574 338272 520076 338328
rect 517513 338270 520076 338272
rect 517513 338267 517579 338270
rect 517513 336970 517579 336973
rect 517513 336968 520076 336970
rect 517513 336912 517518 336968
rect 517574 336912 520076 336968
rect 517513 336910 520076 336912
rect 517513 336907 517579 336910
rect 517513 335610 517579 335613
rect 517513 335608 520076 335610
rect 517513 335552 517518 335608
rect 517574 335552 520076 335608
rect 517513 335550 520076 335552
rect 517513 335547 517579 335550
rect -960 332196 480 332436
rect 531814 330986 531820 330988
rect 529828 330926 531820 330986
rect 531814 330924 531820 330926
rect 531884 330924 531890 330988
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 530577 298754 530643 298757
rect 583520 298754 584960 298844
rect 530577 298752 584960 298754
rect 530577 298696 530582 298752
rect 530638 298696 584960 298752
rect 530577 298694 584960 298696
rect 530577 298691 530643 298694
rect 583520 298604 584960 298694
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 520641 245578 520707 245581
rect 583520 245578 584960 245668
rect 520641 245576 584960 245578
rect 520641 245520 520646 245576
rect 520702 245520 584960 245576
rect 520641 245518 584960 245520
rect 520641 245515 520707 245518
rect 583520 245428 584960 245518
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 308990 165820 308996 165884
rect 309060 165882 309066 165884
rect 583520 165882 584960 165972
rect 309060 165822 584960 165882
rect 309060 165820 309066 165822
rect 583520 165732 584960 165822
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 304758 125972 304764 126036
rect 304828 126034 304834 126036
rect 583520 126034 584960 126124
rect 304828 125974 584960 126034
rect 304828 125972 304834 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 301630 86124 301636 86188
rect 301700 86186 301706 86188
rect 583520 86186 584960 86276
rect 301700 86126 584960 86186
rect 301700 86124 301706 86126
rect 583520 86036 584960 86126
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 312537 46338 312603 46341
rect 583520 46338 584960 46428
rect 312537 46336 584960 46338
rect 312537 46280 312542 46336
rect 312598 46280 584960 46336
rect 312537 46278 584960 46280
rect 312537 46275 312603 46278
rect 583520 46188 584960 46278
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 531814 19756 531820 19820
rect 531884 19818 531890 19820
rect 583520 19818 584960 19908
rect 531884 19758 584960 19818
rect 531884 19756 531890 19758
rect 583520 19668 584960 19758
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 295190 6564 295196 6628
rect 295260 6626 295266 6628
rect 583520 6626 584960 6716
rect 295260 6566 584960 6626
rect 295260 6564 295266 6566
rect 583520 6476 584960 6566
<< via3 >>
rect 299244 354860 299308 354924
rect 299244 353364 299308 353428
rect 308444 352820 308508 352884
rect 295012 351928 295076 351932
rect 295012 351872 295026 351928
rect 295026 351872 295076 351928
rect 295012 351868 295076 351872
rect 301636 351928 301700 351932
rect 301636 351872 301650 351928
rect 301650 351872 301700 351928
rect 301636 351868 301700 351872
rect 304764 351868 304828 351932
rect 531820 330924 531884 330988
rect 308996 165820 309060 165884
rect 304764 125972 304828 126036
rect 301636 86124 301700 86188
rect 531820 19756 531884 19820
rect 295196 6564 295260 6628
<< metal4 >>
rect -3236 705918 -2636 706100
rect -3236 705682 -3054 705918
rect -2818 705682 -2636 705918
rect -3236 675494 -2636 705682
rect -3236 675258 -3054 675494
rect -2818 675258 -2636 675494
rect -3236 638294 -2636 675258
rect -3236 638058 -3054 638294
rect -2818 638058 -2636 638294
rect -3236 601094 -2636 638058
rect -3236 600858 -3054 601094
rect -2818 600858 -2636 601094
rect -3236 563894 -2636 600858
rect -3236 563658 -3054 563894
rect -2818 563658 -2636 563894
rect -3236 526694 -2636 563658
rect -3236 526458 -3054 526694
rect -2818 526458 -2636 526694
rect -3236 489494 -2636 526458
rect -3236 489258 -3054 489494
rect -2818 489258 -2636 489494
rect -3236 452294 -2636 489258
rect -3236 452058 -3054 452294
rect -2818 452058 -2636 452294
rect -3236 415094 -2636 452058
rect -3236 414858 -3054 415094
rect -2818 414858 -2636 415094
rect -3236 377894 -2636 414858
rect -3236 377658 -3054 377894
rect -2818 377658 -2636 377894
rect -3236 340694 -2636 377658
rect -3236 340458 -3054 340694
rect -2818 340458 -2636 340694
rect -3236 303494 -2636 340458
rect -3236 303258 -3054 303494
rect -2818 303258 -2636 303494
rect -3236 266294 -2636 303258
rect -3236 266058 -3054 266294
rect -2818 266058 -2636 266294
rect -3236 229094 -2636 266058
rect -3236 228858 -3054 229094
rect -2818 228858 -2636 229094
rect -3236 191894 -2636 228858
rect -3236 191658 -3054 191894
rect -2818 191658 -2636 191894
rect -3236 154694 -2636 191658
rect -3236 154458 -3054 154694
rect -2818 154458 -2636 154694
rect -3236 117494 -2636 154458
rect -3236 117258 -3054 117494
rect -2818 117258 -2636 117494
rect -3236 80294 -2636 117258
rect -3236 80058 -3054 80294
rect -2818 80058 -2636 80294
rect -3236 43094 -2636 80058
rect -3236 42858 -3054 43094
rect -2818 42858 -2636 43094
rect -3236 5894 -2636 42858
rect -3236 5658 -3054 5894
rect -2818 5658 -2636 5894
rect -3236 -1746 -2636 5658
rect -2296 704978 -1696 705160
rect -2296 704742 -2114 704978
rect -1878 704742 -1696 704978
rect -2296 671894 -1696 704742
rect -2296 671658 -2114 671894
rect -1878 671658 -1696 671894
rect -2296 634694 -1696 671658
rect -2296 634458 -2114 634694
rect -1878 634458 -1696 634694
rect -2296 597494 -1696 634458
rect -2296 597258 -2114 597494
rect -1878 597258 -1696 597494
rect -2296 560294 -1696 597258
rect -2296 560058 -2114 560294
rect -1878 560058 -1696 560294
rect -2296 523094 -1696 560058
rect -2296 522858 -2114 523094
rect -1878 522858 -1696 523094
rect -2296 485894 -1696 522858
rect -2296 485658 -2114 485894
rect -1878 485658 -1696 485894
rect -2296 448694 -1696 485658
rect -2296 448458 -2114 448694
rect -1878 448458 -1696 448694
rect -2296 411494 -1696 448458
rect -2296 411258 -2114 411494
rect -1878 411258 -1696 411494
rect -2296 374294 -1696 411258
rect -2296 374058 -2114 374294
rect -1878 374058 -1696 374294
rect -2296 337094 -1696 374058
rect -2296 336858 -2114 337094
rect -1878 336858 -1696 337094
rect -2296 299894 -1696 336858
rect -2296 299658 -2114 299894
rect -1878 299658 -1696 299894
rect -2296 262694 -1696 299658
rect -2296 262458 -2114 262694
rect -1878 262458 -1696 262694
rect -2296 225494 -1696 262458
rect -2296 225258 -2114 225494
rect -1878 225258 -1696 225494
rect -2296 188294 -1696 225258
rect -2296 188058 -2114 188294
rect -1878 188058 -1696 188294
rect -2296 151094 -1696 188058
rect -2296 150858 -2114 151094
rect -1878 150858 -1696 151094
rect -2296 113894 -1696 150858
rect -2296 113658 -2114 113894
rect -1878 113658 -1696 113894
rect -2296 76694 -1696 113658
rect -2296 76458 -2114 76694
rect -1878 76458 -1696 76694
rect -2296 39494 -1696 76458
rect -2296 39258 -2114 39494
rect -1878 39258 -1696 39494
rect -2296 2294 -1696 39258
rect -2296 2058 -2114 2294
rect -1878 2058 -1696 2294
rect -2296 -806 -1696 2058
rect -2296 -1042 -2114 -806
rect -1878 -1042 -1696 -806
rect -2296 -1224 -1696 -1042
rect 804 704978 1404 706100
rect 804 704742 986 704978
rect 1222 704742 1404 704978
rect 804 671894 1404 704742
rect 804 671658 986 671894
rect 1222 671658 1404 671894
rect 804 634694 1404 671658
rect 804 634458 986 634694
rect 1222 634458 1404 634694
rect 804 597494 1404 634458
rect 804 597258 986 597494
rect 1222 597258 1404 597494
rect 804 560294 1404 597258
rect 804 560058 986 560294
rect 1222 560058 1404 560294
rect 804 523094 1404 560058
rect 804 522858 986 523094
rect 1222 522858 1404 523094
rect 804 485894 1404 522858
rect 804 485658 986 485894
rect 1222 485658 1404 485894
rect 804 448694 1404 485658
rect 804 448458 986 448694
rect 1222 448458 1404 448694
rect 804 411494 1404 448458
rect 804 411258 986 411494
rect 1222 411258 1404 411494
rect 804 374294 1404 411258
rect 804 374058 986 374294
rect 1222 374058 1404 374294
rect 804 337094 1404 374058
rect 804 336858 986 337094
rect 1222 336858 1404 337094
rect 804 299894 1404 336858
rect 804 299658 986 299894
rect 1222 299658 1404 299894
rect 804 262694 1404 299658
rect 804 262458 986 262694
rect 1222 262458 1404 262694
rect 804 225494 1404 262458
rect 804 225258 986 225494
rect 1222 225258 1404 225494
rect 804 188294 1404 225258
rect 804 188058 986 188294
rect 1222 188058 1404 188294
rect 804 151094 1404 188058
rect 804 150858 986 151094
rect 1222 150858 1404 151094
rect 804 113894 1404 150858
rect 804 113658 986 113894
rect 1222 113658 1404 113894
rect 804 76694 1404 113658
rect 804 76458 986 76694
rect 1222 76458 1404 76694
rect 804 39494 1404 76458
rect 804 39258 986 39494
rect 1222 39258 1404 39494
rect 804 2294 1404 39258
rect 804 2058 986 2294
rect 1222 2058 1404 2294
rect 804 -806 1404 2058
rect 804 -1042 986 -806
rect 1222 -1042 1404 -806
rect -3236 -1982 -3054 -1746
rect -2818 -1982 -2636 -1746
rect -3236 -2164 -2636 -1982
rect 804 -2164 1404 -1042
rect 4404 705918 5004 706100
rect 4404 705682 4586 705918
rect 4822 705682 5004 705918
rect 4404 675494 5004 705682
rect 4404 675258 4586 675494
rect 4822 675258 5004 675494
rect 4404 638294 5004 675258
rect 4404 638058 4586 638294
rect 4822 638058 5004 638294
rect 4404 601094 5004 638058
rect 4404 600858 4586 601094
rect 4822 600858 5004 601094
rect 4404 563894 5004 600858
rect 4404 563658 4586 563894
rect 4822 563658 5004 563894
rect 4404 526694 5004 563658
rect 4404 526458 4586 526694
rect 4822 526458 5004 526694
rect 4404 489494 5004 526458
rect 4404 489258 4586 489494
rect 4822 489258 5004 489494
rect 4404 452294 5004 489258
rect 4404 452058 4586 452294
rect 4822 452058 5004 452294
rect 4404 415094 5004 452058
rect 4404 414858 4586 415094
rect 4822 414858 5004 415094
rect 4404 377894 5004 414858
rect 4404 377658 4586 377894
rect 4822 377658 5004 377894
rect 4404 340694 5004 377658
rect 4404 340458 4586 340694
rect 4822 340458 5004 340694
rect 4404 303494 5004 340458
rect 4404 303258 4586 303494
rect 4822 303258 5004 303494
rect 4404 266294 5004 303258
rect 4404 266058 4586 266294
rect 4822 266058 5004 266294
rect 4404 229094 5004 266058
rect 4404 228858 4586 229094
rect 4822 228858 5004 229094
rect 4404 191894 5004 228858
rect 4404 191658 4586 191894
rect 4822 191658 5004 191894
rect 4404 154694 5004 191658
rect 4404 154458 4586 154694
rect 4822 154458 5004 154694
rect 4404 117494 5004 154458
rect 4404 117258 4586 117494
rect 4822 117258 5004 117494
rect 4404 80294 5004 117258
rect 4404 80058 4586 80294
rect 4822 80058 5004 80294
rect 4404 43094 5004 80058
rect 4404 42858 4586 43094
rect 4822 42858 5004 43094
rect 4404 5894 5004 42858
rect 4404 5658 4586 5894
rect 4822 5658 5004 5894
rect 4404 -1746 5004 5658
rect 4404 -1982 4586 -1746
rect 4822 -1982 5004 -1746
rect 4404 -2164 5004 -1982
rect 38004 704978 38604 706100
rect 38004 704742 38186 704978
rect 38422 704742 38604 704978
rect 38004 671894 38604 704742
rect 38004 671658 38186 671894
rect 38422 671658 38604 671894
rect 38004 634694 38604 671658
rect 38004 634458 38186 634694
rect 38422 634458 38604 634694
rect 38004 597494 38604 634458
rect 38004 597258 38186 597494
rect 38422 597258 38604 597494
rect 38004 560294 38604 597258
rect 38004 560058 38186 560294
rect 38422 560058 38604 560294
rect 38004 523094 38604 560058
rect 38004 522858 38186 523094
rect 38422 522858 38604 523094
rect 38004 485894 38604 522858
rect 38004 485658 38186 485894
rect 38422 485658 38604 485894
rect 38004 448694 38604 485658
rect 38004 448458 38186 448694
rect 38422 448458 38604 448694
rect 38004 411494 38604 448458
rect 38004 411258 38186 411494
rect 38422 411258 38604 411494
rect 38004 374294 38604 411258
rect 38004 374058 38186 374294
rect 38422 374058 38604 374294
rect 38004 337094 38604 374058
rect 38004 336858 38186 337094
rect 38422 336858 38604 337094
rect 38004 299894 38604 336858
rect 38004 299658 38186 299894
rect 38422 299658 38604 299894
rect 38004 262694 38604 299658
rect 38004 262458 38186 262694
rect 38422 262458 38604 262694
rect 38004 225494 38604 262458
rect 38004 225258 38186 225494
rect 38422 225258 38604 225494
rect 38004 188294 38604 225258
rect 38004 188058 38186 188294
rect 38422 188058 38604 188294
rect 38004 151094 38604 188058
rect 38004 150858 38186 151094
rect 38422 150858 38604 151094
rect 38004 113894 38604 150858
rect 38004 113658 38186 113894
rect 38422 113658 38604 113894
rect 38004 76694 38604 113658
rect 38004 76458 38186 76694
rect 38422 76458 38604 76694
rect 38004 39494 38604 76458
rect 38004 39258 38186 39494
rect 38422 39258 38604 39494
rect 38004 2294 38604 39258
rect 38004 2058 38186 2294
rect 38422 2058 38604 2294
rect 38004 -806 38604 2058
rect 38004 -1042 38186 -806
rect 38422 -1042 38604 -806
rect 38004 -2164 38604 -1042
rect 41604 705918 42204 706100
rect 41604 705682 41786 705918
rect 42022 705682 42204 705918
rect 41604 675494 42204 705682
rect 41604 675258 41786 675494
rect 42022 675258 42204 675494
rect 41604 638294 42204 675258
rect 41604 638058 41786 638294
rect 42022 638058 42204 638294
rect 41604 601094 42204 638058
rect 41604 600858 41786 601094
rect 42022 600858 42204 601094
rect 41604 563894 42204 600858
rect 41604 563658 41786 563894
rect 42022 563658 42204 563894
rect 41604 526694 42204 563658
rect 41604 526458 41786 526694
rect 42022 526458 42204 526694
rect 41604 489494 42204 526458
rect 41604 489258 41786 489494
rect 42022 489258 42204 489494
rect 41604 452294 42204 489258
rect 41604 452058 41786 452294
rect 42022 452058 42204 452294
rect 41604 415094 42204 452058
rect 41604 414858 41786 415094
rect 42022 414858 42204 415094
rect 41604 377894 42204 414858
rect 41604 377658 41786 377894
rect 42022 377658 42204 377894
rect 41604 340694 42204 377658
rect 41604 340458 41786 340694
rect 42022 340458 42204 340694
rect 41604 303494 42204 340458
rect 41604 303258 41786 303494
rect 42022 303258 42204 303494
rect 41604 266294 42204 303258
rect 41604 266058 41786 266294
rect 42022 266058 42204 266294
rect 41604 229094 42204 266058
rect 41604 228858 41786 229094
rect 42022 228858 42204 229094
rect 41604 191894 42204 228858
rect 41604 191658 41786 191894
rect 42022 191658 42204 191894
rect 41604 154694 42204 191658
rect 41604 154458 41786 154694
rect 42022 154458 42204 154694
rect 41604 117494 42204 154458
rect 41604 117258 41786 117494
rect 42022 117258 42204 117494
rect 41604 80294 42204 117258
rect 41604 80058 41786 80294
rect 42022 80058 42204 80294
rect 41604 43094 42204 80058
rect 41604 42858 41786 43094
rect 42022 42858 42204 43094
rect 41604 5894 42204 42858
rect 41604 5658 41786 5894
rect 42022 5658 42204 5894
rect 41604 -1746 42204 5658
rect 41604 -1982 41786 -1746
rect 42022 -1982 42204 -1746
rect 41604 -2164 42204 -1982
rect 75204 704978 75804 706100
rect 75204 704742 75386 704978
rect 75622 704742 75804 704978
rect 75204 671894 75804 704742
rect 75204 671658 75386 671894
rect 75622 671658 75804 671894
rect 75204 634694 75804 671658
rect 75204 634458 75386 634694
rect 75622 634458 75804 634694
rect 75204 597494 75804 634458
rect 75204 597258 75386 597494
rect 75622 597258 75804 597494
rect 75204 560294 75804 597258
rect 75204 560058 75386 560294
rect 75622 560058 75804 560294
rect 75204 523094 75804 560058
rect 75204 522858 75386 523094
rect 75622 522858 75804 523094
rect 75204 485894 75804 522858
rect 75204 485658 75386 485894
rect 75622 485658 75804 485894
rect 75204 448694 75804 485658
rect 75204 448458 75386 448694
rect 75622 448458 75804 448694
rect 75204 411494 75804 448458
rect 75204 411258 75386 411494
rect 75622 411258 75804 411494
rect 75204 374294 75804 411258
rect 75204 374058 75386 374294
rect 75622 374058 75804 374294
rect 75204 337094 75804 374058
rect 75204 336858 75386 337094
rect 75622 336858 75804 337094
rect 75204 299894 75804 336858
rect 75204 299658 75386 299894
rect 75622 299658 75804 299894
rect 75204 262694 75804 299658
rect 75204 262458 75386 262694
rect 75622 262458 75804 262694
rect 75204 225494 75804 262458
rect 75204 225258 75386 225494
rect 75622 225258 75804 225494
rect 75204 188294 75804 225258
rect 75204 188058 75386 188294
rect 75622 188058 75804 188294
rect 75204 151094 75804 188058
rect 75204 150858 75386 151094
rect 75622 150858 75804 151094
rect 75204 113894 75804 150858
rect 75204 113658 75386 113894
rect 75622 113658 75804 113894
rect 75204 76694 75804 113658
rect 75204 76458 75386 76694
rect 75622 76458 75804 76694
rect 75204 39494 75804 76458
rect 75204 39258 75386 39494
rect 75622 39258 75804 39494
rect 75204 2294 75804 39258
rect 75204 2058 75386 2294
rect 75622 2058 75804 2294
rect 75204 -806 75804 2058
rect 75204 -1042 75386 -806
rect 75622 -1042 75804 -806
rect 75204 -2164 75804 -1042
rect 78804 705918 79404 706100
rect 78804 705682 78986 705918
rect 79222 705682 79404 705918
rect 78804 675494 79404 705682
rect 78804 675258 78986 675494
rect 79222 675258 79404 675494
rect 78804 638294 79404 675258
rect 78804 638058 78986 638294
rect 79222 638058 79404 638294
rect 78804 601094 79404 638058
rect 78804 600858 78986 601094
rect 79222 600858 79404 601094
rect 78804 563894 79404 600858
rect 78804 563658 78986 563894
rect 79222 563658 79404 563894
rect 78804 526694 79404 563658
rect 78804 526458 78986 526694
rect 79222 526458 79404 526694
rect 78804 489494 79404 526458
rect 78804 489258 78986 489494
rect 79222 489258 79404 489494
rect 78804 452294 79404 489258
rect 78804 452058 78986 452294
rect 79222 452058 79404 452294
rect 78804 415094 79404 452058
rect 78804 414858 78986 415094
rect 79222 414858 79404 415094
rect 78804 377894 79404 414858
rect 78804 377658 78986 377894
rect 79222 377658 79404 377894
rect 78804 340694 79404 377658
rect 78804 340458 78986 340694
rect 79222 340458 79404 340694
rect 78804 303494 79404 340458
rect 78804 303258 78986 303494
rect 79222 303258 79404 303494
rect 78804 266294 79404 303258
rect 78804 266058 78986 266294
rect 79222 266058 79404 266294
rect 78804 229094 79404 266058
rect 78804 228858 78986 229094
rect 79222 228858 79404 229094
rect 78804 191894 79404 228858
rect 78804 191658 78986 191894
rect 79222 191658 79404 191894
rect 78804 154694 79404 191658
rect 78804 154458 78986 154694
rect 79222 154458 79404 154694
rect 78804 117494 79404 154458
rect 78804 117258 78986 117494
rect 79222 117258 79404 117494
rect 78804 80294 79404 117258
rect 78804 80058 78986 80294
rect 79222 80058 79404 80294
rect 78804 43094 79404 80058
rect 78804 42858 78986 43094
rect 79222 42858 79404 43094
rect 78804 5894 79404 42858
rect 78804 5658 78986 5894
rect 79222 5658 79404 5894
rect 78804 -1746 79404 5658
rect 78804 -1982 78986 -1746
rect 79222 -1982 79404 -1746
rect 78804 -2164 79404 -1982
rect 112404 704978 113004 706100
rect 112404 704742 112586 704978
rect 112822 704742 113004 704978
rect 112404 671894 113004 704742
rect 112404 671658 112586 671894
rect 112822 671658 113004 671894
rect 112404 634694 113004 671658
rect 112404 634458 112586 634694
rect 112822 634458 113004 634694
rect 112404 597494 113004 634458
rect 112404 597258 112586 597494
rect 112822 597258 113004 597494
rect 112404 560294 113004 597258
rect 112404 560058 112586 560294
rect 112822 560058 113004 560294
rect 112404 523094 113004 560058
rect 112404 522858 112586 523094
rect 112822 522858 113004 523094
rect 112404 485894 113004 522858
rect 112404 485658 112586 485894
rect 112822 485658 113004 485894
rect 112404 448694 113004 485658
rect 112404 448458 112586 448694
rect 112822 448458 113004 448694
rect 112404 411494 113004 448458
rect 112404 411258 112586 411494
rect 112822 411258 113004 411494
rect 112404 374294 113004 411258
rect 112404 374058 112586 374294
rect 112822 374058 113004 374294
rect 112404 337094 113004 374058
rect 112404 336858 112586 337094
rect 112822 336858 113004 337094
rect 112404 299894 113004 336858
rect 112404 299658 112586 299894
rect 112822 299658 113004 299894
rect 112404 262694 113004 299658
rect 112404 262458 112586 262694
rect 112822 262458 113004 262694
rect 112404 225494 113004 262458
rect 112404 225258 112586 225494
rect 112822 225258 113004 225494
rect 112404 188294 113004 225258
rect 112404 188058 112586 188294
rect 112822 188058 113004 188294
rect 112404 151094 113004 188058
rect 112404 150858 112586 151094
rect 112822 150858 113004 151094
rect 112404 113894 113004 150858
rect 112404 113658 112586 113894
rect 112822 113658 113004 113894
rect 112404 76694 113004 113658
rect 112404 76458 112586 76694
rect 112822 76458 113004 76694
rect 112404 39494 113004 76458
rect 112404 39258 112586 39494
rect 112822 39258 113004 39494
rect 112404 2294 113004 39258
rect 112404 2058 112586 2294
rect 112822 2058 113004 2294
rect 112404 -806 113004 2058
rect 112404 -1042 112586 -806
rect 112822 -1042 113004 -806
rect 112404 -2164 113004 -1042
rect 116004 705918 116604 706100
rect 116004 705682 116186 705918
rect 116422 705682 116604 705918
rect 116004 675494 116604 705682
rect 116004 675258 116186 675494
rect 116422 675258 116604 675494
rect 116004 638294 116604 675258
rect 116004 638058 116186 638294
rect 116422 638058 116604 638294
rect 116004 601094 116604 638058
rect 116004 600858 116186 601094
rect 116422 600858 116604 601094
rect 116004 563894 116604 600858
rect 116004 563658 116186 563894
rect 116422 563658 116604 563894
rect 116004 526694 116604 563658
rect 116004 526458 116186 526694
rect 116422 526458 116604 526694
rect 116004 489494 116604 526458
rect 116004 489258 116186 489494
rect 116422 489258 116604 489494
rect 116004 452294 116604 489258
rect 116004 452058 116186 452294
rect 116422 452058 116604 452294
rect 116004 415094 116604 452058
rect 116004 414858 116186 415094
rect 116422 414858 116604 415094
rect 116004 377894 116604 414858
rect 116004 377658 116186 377894
rect 116422 377658 116604 377894
rect 116004 340694 116604 377658
rect 116004 340458 116186 340694
rect 116422 340458 116604 340694
rect 116004 303494 116604 340458
rect 116004 303258 116186 303494
rect 116422 303258 116604 303494
rect 116004 266294 116604 303258
rect 116004 266058 116186 266294
rect 116422 266058 116604 266294
rect 116004 229094 116604 266058
rect 116004 228858 116186 229094
rect 116422 228858 116604 229094
rect 116004 191894 116604 228858
rect 116004 191658 116186 191894
rect 116422 191658 116604 191894
rect 116004 154694 116604 191658
rect 116004 154458 116186 154694
rect 116422 154458 116604 154694
rect 116004 117494 116604 154458
rect 116004 117258 116186 117494
rect 116422 117258 116604 117494
rect 116004 80294 116604 117258
rect 116004 80058 116186 80294
rect 116422 80058 116604 80294
rect 116004 43094 116604 80058
rect 116004 42858 116186 43094
rect 116422 42858 116604 43094
rect 116004 5894 116604 42858
rect 116004 5658 116186 5894
rect 116422 5658 116604 5894
rect 116004 -1746 116604 5658
rect 116004 -1982 116186 -1746
rect 116422 -1982 116604 -1746
rect 116004 -2164 116604 -1982
rect 149604 704978 150204 706100
rect 149604 704742 149786 704978
rect 150022 704742 150204 704978
rect 149604 671894 150204 704742
rect 149604 671658 149786 671894
rect 150022 671658 150204 671894
rect 149604 634694 150204 671658
rect 149604 634458 149786 634694
rect 150022 634458 150204 634694
rect 149604 597494 150204 634458
rect 149604 597258 149786 597494
rect 150022 597258 150204 597494
rect 149604 560294 150204 597258
rect 149604 560058 149786 560294
rect 150022 560058 150204 560294
rect 149604 523094 150204 560058
rect 149604 522858 149786 523094
rect 150022 522858 150204 523094
rect 149604 485894 150204 522858
rect 149604 485658 149786 485894
rect 150022 485658 150204 485894
rect 149604 448694 150204 485658
rect 149604 448458 149786 448694
rect 150022 448458 150204 448694
rect 149604 411494 150204 448458
rect 149604 411258 149786 411494
rect 150022 411258 150204 411494
rect 149604 374294 150204 411258
rect 149604 374058 149786 374294
rect 150022 374058 150204 374294
rect 149604 337094 150204 374058
rect 149604 336858 149786 337094
rect 150022 336858 150204 337094
rect 149604 299894 150204 336858
rect 149604 299658 149786 299894
rect 150022 299658 150204 299894
rect 149604 262694 150204 299658
rect 149604 262458 149786 262694
rect 150022 262458 150204 262694
rect 149604 225494 150204 262458
rect 149604 225258 149786 225494
rect 150022 225258 150204 225494
rect 149604 188294 150204 225258
rect 149604 188058 149786 188294
rect 150022 188058 150204 188294
rect 149604 151094 150204 188058
rect 149604 150858 149786 151094
rect 150022 150858 150204 151094
rect 149604 113894 150204 150858
rect 149604 113658 149786 113894
rect 150022 113658 150204 113894
rect 149604 76694 150204 113658
rect 149604 76458 149786 76694
rect 150022 76458 150204 76694
rect 149604 39494 150204 76458
rect 149604 39258 149786 39494
rect 150022 39258 150204 39494
rect 149604 2294 150204 39258
rect 149604 2058 149786 2294
rect 150022 2058 150204 2294
rect 149604 -806 150204 2058
rect 149604 -1042 149786 -806
rect 150022 -1042 150204 -806
rect 149604 -2164 150204 -1042
rect 153204 705918 153804 706100
rect 153204 705682 153386 705918
rect 153622 705682 153804 705918
rect 153204 675494 153804 705682
rect 153204 675258 153386 675494
rect 153622 675258 153804 675494
rect 153204 638294 153804 675258
rect 153204 638058 153386 638294
rect 153622 638058 153804 638294
rect 153204 601094 153804 638058
rect 153204 600858 153386 601094
rect 153622 600858 153804 601094
rect 153204 563894 153804 600858
rect 153204 563658 153386 563894
rect 153622 563658 153804 563894
rect 153204 526694 153804 563658
rect 153204 526458 153386 526694
rect 153622 526458 153804 526694
rect 153204 489494 153804 526458
rect 153204 489258 153386 489494
rect 153622 489258 153804 489494
rect 153204 452294 153804 489258
rect 153204 452058 153386 452294
rect 153622 452058 153804 452294
rect 153204 415094 153804 452058
rect 153204 414858 153386 415094
rect 153622 414858 153804 415094
rect 153204 377894 153804 414858
rect 153204 377658 153386 377894
rect 153622 377658 153804 377894
rect 153204 340694 153804 377658
rect 153204 340458 153386 340694
rect 153622 340458 153804 340694
rect 153204 303494 153804 340458
rect 153204 303258 153386 303494
rect 153622 303258 153804 303494
rect 153204 266294 153804 303258
rect 153204 266058 153386 266294
rect 153622 266058 153804 266294
rect 153204 229094 153804 266058
rect 153204 228858 153386 229094
rect 153622 228858 153804 229094
rect 153204 191894 153804 228858
rect 153204 191658 153386 191894
rect 153622 191658 153804 191894
rect 153204 154694 153804 191658
rect 153204 154458 153386 154694
rect 153622 154458 153804 154694
rect 153204 117494 153804 154458
rect 153204 117258 153386 117494
rect 153622 117258 153804 117494
rect 153204 80294 153804 117258
rect 153204 80058 153386 80294
rect 153622 80058 153804 80294
rect 153204 43094 153804 80058
rect 153204 42858 153386 43094
rect 153622 42858 153804 43094
rect 153204 5894 153804 42858
rect 153204 5658 153386 5894
rect 153622 5658 153804 5894
rect 153204 -1746 153804 5658
rect 153204 -1982 153386 -1746
rect 153622 -1982 153804 -1746
rect 153204 -2164 153804 -1982
rect 186804 704978 187404 706100
rect 186804 704742 186986 704978
rect 187222 704742 187404 704978
rect 186804 671894 187404 704742
rect 186804 671658 186986 671894
rect 187222 671658 187404 671894
rect 186804 634694 187404 671658
rect 186804 634458 186986 634694
rect 187222 634458 187404 634694
rect 186804 597494 187404 634458
rect 186804 597258 186986 597494
rect 187222 597258 187404 597494
rect 186804 560294 187404 597258
rect 186804 560058 186986 560294
rect 187222 560058 187404 560294
rect 186804 523094 187404 560058
rect 186804 522858 186986 523094
rect 187222 522858 187404 523094
rect 186804 485894 187404 522858
rect 186804 485658 186986 485894
rect 187222 485658 187404 485894
rect 186804 448694 187404 485658
rect 186804 448458 186986 448694
rect 187222 448458 187404 448694
rect 186804 411494 187404 448458
rect 186804 411258 186986 411494
rect 187222 411258 187404 411494
rect 186804 374294 187404 411258
rect 186804 374058 186986 374294
rect 187222 374058 187404 374294
rect 186804 337094 187404 374058
rect 186804 336858 186986 337094
rect 187222 336858 187404 337094
rect 186804 299894 187404 336858
rect 186804 299658 186986 299894
rect 187222 299658 187404 299894
rect 186804 262694 187404 299658
rect 186804 262458 186986 262694
rect 187222 262458 187404 262694
rect 186804 225494 187404 262458
rect 186804 225258 186986 225494
rect 187222 225258 187404 225494
rect 186804 188294 187404 225258
rect 186804 188058 186986 188294
rect 187222 188058 187404 188294
rect 186804 151094 187404 188058
rect 186804 150858 186986 151094
rect 187222 150858 187404 151094
rect 186804 113894 187404 150858
rect 186804 113658 186986 113894
rect 187222 113658 187404 113894
rect 186804 76694 187404 113658
rect 186804 76458 186986 76694
rect 187222 76458 187404 76694
rect 186804 39494 187404 76458
rect 186804 39258 186986 39494
rect 187222 39258 187404 39494
rect 186804 2294 187404 39258
rect 186804 2058 186986 2294
rect 187222 2058 187404 2294
rect 186804 -806 187404 2058
rect 186804 -1042 186986 -806
rect 187222 -1042 187404 -806
rect 186804 -2164 187404 -1042
rect 190404 705918 191004 706100
rect 190404 705682 190586 705918
rect 190822 705682 191004 705918
rect 190404 675494 191004 705682
rect 190404 675258 190586 675494
rect 190822 675258 191004 675494
rect 190404 638294 191004 675258
rect 190404 638058 190586 638294
rect 190822 638058 191004 638294
rect 190404 601094 191004 638058
rect 190404 600858 190586 601094
rect 190822 600858 191004 601094
rect 190404 563894 191004 600858
rect 190404 563658 190586 563894
rect 190822 563658 191004 563894
rect 190404 526694 191004 563658
rect 190404 526458 190586 526694
rect 190822 526458 191004 526694
rect 190404 489494 191004 526458
rect 190404 489258 190586 489494
rect 190822 489258 191004 489494
rect 190404 452294 191004 489258
rect 190404 452058 190586 452294
rect 190822 452058 191004 452294
rect 190404 415094 191004 452058
rect 190404 414858 190586 415094
rect 190822 414858 191004 415094
rect 190404 377894 191004 414858
rect 190404 377658 190586 377894
rect 190822 377658 191004 377894
rect 190404 340694 191004 377658
rect 190404 340458 190586 340694
rect 190822 340458 191004 340694
rect 190404 303494 191004 340458
rect 190404 303258 190586 303494
rect 190822 303258 191004 303494
rect 190404 266294 191004 303258
rect 190404 266058 190586 266294
rect 190822 266058 191004 266294
rect 190404 229094 191004 266058
rect 190404 228858 190586 229094
rect 190822 228858 191004 229094
rect 190404 191894 191004 228858
rect 190404 191658 190586 191894
rect 190822 191658 191004 191894
rect 190404 154694 191004 191658
rect 190404 154458 190586 154694
rect 190822 154458 191004 154694
rect 190404 117494 191004 154458
rect 190404 117258 190586 117494
rect 190822 117258 191004 117494
rect 190404 80294 191004 117258
rect 190404 80058 190586 80294
rect 190822 80058 191004 80294
rect 190404 43094 191004 80058
rect 190404 42858 190586 43094
rect 190822 42858 191004 43094
rect 190404 5894 191004 42858
rect 190404 5658 190586 5894
rect 190822 5658 191004 5894
rect 190404 -1746 191004 5658
rect 190404 -1982 190586 -1746
rect 190822 -1982 191004 -1746
rect 190404 -2164 191004 -1982
rect 224004 704978 224604 706100
rect 224004 704742 224186 704978
rect 224422 704742 224604 704978
rect 224004 671894 224604 704742
rect 224004 671658 224186 671894
rect 224422 671658 224604 671894
rect 224004 634694 224604 671658
rect 224004 634458 224186 634694
rect 224422 634458 224604 634694
rect 224004 597494 224604 634458
rect 224004 597258 224186 597494
rect 224422 597258 224604 597494
rect 224004 560294 224604 597258
rect 224004 560058 224186 560294
rect 224422 560058 224604 560294
rect 224004 523094 224604 560058
rect 224004 522858 224186 523094
rect 224422 522858 224604 523094
rect 224004 485894 224604 522858
rect 224004 485658 224186 485894
rect 224422 485658 224604 485894
rect 224004 448694 224604 485658
rect 224004 448458 224186 448694
rect 224422 448458 224604 448694
rect 224004 411494 224604 448458
rect 224004 411258 224186 411494
rect 224422 411258 224604 411494
rect 224004 374294 224604 411258
rect 224004 374058 224186 374294
rect 224422 374058 224604 374294
rect 224004 337094 224604 374058
rect 224004 336858 224186 337094
rect 224422 336858 224604 337094
rect 224004 299894 224604 336858
rect 224004 299658 224186 299894
rect 224422 299658 224604 299894
rect 224004 262694 224604 299658
rect 224004 262458 224186 262694
rect 224422 262458 224604 262694
rect 224004 225494 224604 262458
rect 224004 225258 224186 225494
rect 224422 225258 224604 225494
rect 224004 188294 224604 225258
rect 224004 188058 224186 188294
rect 224422 188058 224604 188294
rect 224004 151094 224604 188058
rect 224004 150858 224186 151094
rect 224422 150858 224604 151094
rect 224004 113894 224604 150858
rect 224004 113658 224186 113894
rect 224422 113658 224604 113894
rect 224004 76694 224604 113658
rect 224004 76458 224186 76694
rect 224422 76458 224604 76694
rect 224004 39494 224604 76458
rect 224004 39258 224186 39494
rect 224422 39258 224604 39494
rect 224004 2294 224604 39258
rect 224004 2058 224186 2294
rect 224422 2058 224604 2294
rect 224004 -806 224604 2058
rect 224004 -1042 224186 -806
rect 224422 -1042 224604 -806
rect 224004 -2164 224604 -1042
rect 227604 705918 228204 706100
rect 227604 705682 227786 705918
rect 228022 705682 228204 705918
rect 227604 675494 228204 705682
rect 227604 675258 227786 675494
rect 228022 675258 228204 675494
rect 227604 638294 228204 675258
rect 227604 638058 227786 638294
rect 228022 638058 228204 638294
rect 227604 601094 228204 638058
rect 227604 600858 227786 601094
rect 228022 600858 228204 601094
rect 227604 563894 228204 600858
rect 227604 563658 227786 563894
rect 228022 563658 228204 563894
rect 227604 526694 228204 563658
rect 227604 526458 227786 526694
rect 228022 526458 228204 526694
rect 227604 489494 228204 526458
rect 227604 489258 227786 489494
rect 228022 489258 228204 489494
rect 227604 452294 228204 489258
rect 227604 452058 227786 452294
rect 228022 452058 228204 452294
rect 227604 415094 228204 452058
rect 227604 414858 227786 415094
rect 228022 414858 228204 415094
rect 227604 377894 228204 414858
rect 227604 377658 227786 377894
rect 228022 377658 228204 377894
rect 227604 340694 228204 377658
rect 227604 340458 227786 340694
rect 228022 340458 228204 340694
rect 227604 303494 228204 340458
rect 227604 303258 227786 303494
rect 228022 303258 228204 303494
rect 227604 266294 228204 303258
rect 227604 266058 227786 266294
rect 228022 266058 228204 266294
rect 227604 229094 228204 266058
rect 227604 228858 227786 229094
rect 228022 228858 228204 229094
rect 227604 191894 228204 228858
rect 227604 191658 227786 191894
rect 228022 191658 228204 191894
rect 227604 154694 228204 191658
rect 227604 154458 227786 154694
rect 228022 154458 228204 154694
rect 227604 117494 228204 154458
rect 227604 117258 227786 117494
rect 228022 117258 228204 117494
rect 227604 80294 228204 117258
rect 227604 80058 227786 80294
rect 228022 80058 228204 80294
rect 227604 43094 228204 80058
rect 227604 42858 227786 43094
rect 228022 42858 228204 43094
rect 227604 5894 228204 42858
rect 227604 5658 227786 5894
rect 228022 5658 228204 5894
rect 227604 -1746 228204 5658
rect 227604 -1982 227786 -1746
rect 228022 -1982 228204 -1746
rect 227604 -2164 228204 -1982
rect 261204 704978 261804 706100
rect 261204 704742 261386 704978
rect 261622 704742 261804 704978
rect 261204 671894 261804 704742
rect 261204 671658 261386 671894
rect 261622 671658 261804 671894
rect 261204 634694 261804 671658
rect 261204 634458 261386 634694
rect 261622 634458 261804 634694
rect 261204 597494 261804 634458
rect 261204 597258 261386 597494
rect 261622 597258 261804 597494
rect 261204 560294 261804 597258
rect 261204 560058 261386 560294
rect 261622 560058 261804 560294
rect 261204 523094 261804 560058
rect 261204 522858 261386 523094
rect 261622 522858 261804 523094
rect 261204 485894 261804 522858
rect 261204 485658 261386 485894
rect 261622 485658 261804 485894
rect 261204 448694 261804 485658
rect 261204 448458 261386 448694
rect 261622 448458 261804 448694
rect 261204 411494 261804 448458
rect 261204 411258 261386 411494
rect 261622 411258 261804 411494
rect 261204 374294 261804 411258
rect 261204 374058 261386 374294
rect 261622 374058 261804 374294
rect 261204 337094 261804 374058
rect 261204 336858 261386 337094
rect 261622 336858 261804 337094
rect 261204 299894 261804 336858
rect 261204 299658 261386 299894
rect 261622 299658 261804 299894
rect 261204 262694 261804 299658
rect 261204 262458 261386 262694
rect 261622 262458 261804 262694
rect 261204 225494 261804 262458
rect 261204 225258 261386 225494
rect 261622 225258 261804 225494
rect 261204 188294 261804 225258
rect 261204 188058 261386 188294
rect 261622 188058 261804 188294
rect 261204 151094 261804 188058
rect 261204 150858 261386 151094
rect 261622 150858 261804 151094
rect 261204 113894 261804 150858
rect 261204 113658 261386 113894
rect 261622 113658 261804 113894
rect 261204 76694 261804 113658
rect 261204 76458 261386 76694
rect 261622 76458 261804 76694
rect 261204 39494 261804 76458
rect 261204 39258 261386 39494
rect 261622 39258 261804 39494
rect 261204 2294 261804 39258
rect 261204 2058 261386 2294
rect 261622 2058 261804 2294
rect 261204 -806 261804 2058
rect 261204 -1042 261386 -806
rect 261622 -1042 261804 -806
rect 261204 -2164 261804 -1042
rect 264804 705918 265404 706100
rect 264804 705682 264986 705918
rect 265222 705682 265404 705918
rect 264804 675494 265404 705682
rect 264804 675258 264986 675494
rect 265222 675258 265404 675494
rect 264804 638294 265404 675258
rect 264804 638058 264986 638294
rect 265222 638058 265404 638294
rect 264804 601094 265404 638058
rect 264804 600858 264986 601094
rect 265222 600858 265404 601094
rect 264804 563894 265404 600858
rect 264804 563658 264986 563894
rect 265222 563658 265404 563894
rect 264804 526694 265404 563658
rect 264804 526458 264986 526694
rect 265222 526458 265404 526694
rect 264804 489494 265404 526458
rect 264804 489258 264986 489494
rect 265222 489258 265404 489494
rect 264804 452294 265404 489258
rect 264804 452058 264986 452294
rect 265222 452058 265404 452294
rect 264804 415094 265404 452058
rect 264804 414858 264986 415094
rect 265222 414858 265404 415094
rect 264804 377894 265404 414858
rect 264804 377658 264986 377894
rect 265222 377658 265404 377894
rect 264804 340694 265404 377658
rect 298404 704978 299004 706100
rect 298404 704742 298586 704978
rect 298822 704742 299004 704978
rect 298404 671894 299004 704742
rect 298404 671658 298586 671894
rect 298822 671658 299004 671894
rect 298404 634694 299004 671658
rect 298404 634458 298586 634694
rect 298822 634458 299004 634694
rect 298404 597494 299004 634458
rect 298404 597258 298586 597494
rect 298822 597258 299004 597494
rect 298404 560294 299004 597258
rect 298404 560058 298586 560294
rect 298822 560058 299004 560294
rect 298404 523094 299004 560058
rect 298404 522858 298586 523094
rect 298822 522858 299004 523094
rect 298404 485894 299004 522858
rect 298404 485658 298586 485894
rect 298822 485658 299004 485894
rect 298404 448694 299004 485658
rect 298404 448458 298586 448694
rect 298822 448458 299004 448694
rect 298404 411494 299004 448458
rect 298404 411258 298586 411494
rect 298822 411258 299004 411494
rect 298404 374294 299004 411258
rect 298404 374058 298586 374294
rect 298822 374058 299004 374294
rect 295011 351932 295077 351933
rect 295011 351868 295012 351932
rect 295076 351868 295077 351932
rect 295011 351867 295077 351868
rect 295014 345030 295074 351867
rect 295014 344970 295258 345030
rect 264804 340458 264986 340694
rect 265222 340458 265404 340694
rect 264804 303494 265404 340458
rect 264804 303258 264986 303494
rect 265222 303258 265404 303494
rect 264804 266294 265404 303258
rect 264804 266058 264986 266294
rect 265222 266058 265404 266294
rect 264804 229094 265404 266058
rect 264804 228858 264986 229094
rect 265222 228858 265404 229094
rect 264804 191894 265404 228858
rect 264804 191658 264986 191894
rect 265222 191658 265404 191894
rect 264804 154694 265404 191658
rect 264804 154458 264986 154694
rect 265222 154458 265404 154694
rect 264804 117494 265404 154458
rect 264804 117258 264986 117494
rect 265222 117258 265404 117494
rect 264804 80294 265404 117258
rect 264804 80058 264986 80294
rect 265222 80058 265404 80294
rect 264804 43094 265404 80058
rect 264804 42858 264986 43094
rect 265222 42858 265404 43094
rect 264804 5894 265404 42858
rect 295198 6629 295258 344970
rect 298404 337094 299004 374058
rect 302004 705918 302604 706100
rect 302004 705682 302186 705918
rect 302422 705682 302604 705918
rect 302004 675494 302604 705682
rect 302004 675258 302186 675494
rect 302422 675258 302604 675494
rect 302004 638294 302604 675258
rect 302004 638058 302186 638294
rect 302422 638058 302604 638294
rect 302004 601094 302604 638058
rect 302004 600858 302186 601094
rect 302422 600858 302604 601094
rect 302004 563894 302604 600858
rect 302004 563658 302186 563894
rect 302422 563658 302604 563894
rect 302004 526694 302604 563658
rect 302004 526458 302186 526694
rect 302422 526458 302604 526694
rect 302004 489494 302604 526458
rect 302004 489258 302186 489494
rect 302422 489258 302604 489494
rect 302004 452294 302604 489258
rect 302004 452058 302186 452294
rect 302422 452058 302604 452294
rect 302004 415094 302604 452058
rect 302004 414858 302186 415094
rect 302422 414858 302604 415094
rect 302004 377894 302604 414858
rect 302004 377658 302186 377894
rect 302422 377658 302604 377894
rect 299243 354924 299309 354925
rect 299243 354860 299244 354924
rect 299308 354860 299309 354924
rect 299243 354859 299309 354860
rect 299246 353429 299306 354859
rect 299243 353428 299309 353429
rect 299243 353364 299244 353428
rect 299308 353364 299309 353428
rect 299243 353363 299309 353364
rect 301635 351932 301701 351933
rect 301635 351868 301636 351932
rect 301700 351868 301701 351932
rect 301635 351867 301701 351868
rect 298404 336858 298586 337094
rect 298822 336858 299004 337094
rect 298404 299894 299004 336858
rect 298404 299658 298586 299894
rect 298822 299658 299004 299894
rect 298404 262694 299004 299658
rect 298404 262458 298586 262694
rect 298822 262458 299004 262694
rect 298404 225494 299004 262458
rect 298404 225258 298586 225494
rect 298822 225258 299004 225494
rect 298404 188294 299004 225258
rect 298404 188058 298586 188294
rect 298822 188058 299004 188294
rect 298404 151094 299004 188058
rect 298404 150858 298586 151094
rect 298822 150858 299004 151094
rect 298404 113894 299004 150858
rect 298404 113658 298586 113894
rect 298822 113658 299004 113894
rect 298404 76694 299004 113658
rect 301638 86189 301698 351867
rect 302004 340694 302604 377658
rect 335604 704978 336204 706100
rect 335604 704742 335786 704978
rect 336022 704742 336204 704978
rect 335604 671894 336204 704742
rect 335604 671658 335786 671894
rect 336022 671658 336204 671894
rect 335604 634694 336204 671658
rect 335604 634458 335786 634694
rect 336022 634458 336204 634694
rect 335604 597494 336204 634458
rect 335604 597258 335786 597494
rect 336022 597258 336204 597494
rect 335604 560294 336204 597258
rect 335604 560058 335786 560294
rect 336022 560058 336204 560294
rect 335604 523094 336204 560058
rect 335604 522858 335786 523094
rect 336022 522858 336204 523094
rect 335604 485894 336204 522858
rect 335604 485658 335786 485894
rect 336022 485658 336204 485894
rect 335604 448694 336204 485658
rect 335604 448458 335786 448694
rect 336022 448458 336204 448694
rect 335604 411494 336204 448458
rect 335604 411258 335786 411494
rect 336022 411258 336204 411494
rect 335604 374294 336204 411258
rect 335604 374058 335786 374294
rect 336022 374058 336204 374294
rect 308443 352884 308509 352885
rect 308443 352820 308444 352884
rect 308508 352820 308509 352884
rect 308443 352819 308509 352820
rect 308446 352610 308506 352819
rect 308446 352550 309058 352610
rect 304763 351932 304829 351933
rect 304763 351868 304764 351932
rect 304828 351868 304829 351932
rect 304763 351867 304829 351868
rect 302004 340458 302186 340694
rect 302422 340458 302604 340694
rect 302004 303494 302604 340458
rect 302004 303258 302186 303494
rect 302422 303258 302604 303494
rect 302004 266294 302604 303258
rect 302004 266058 302186 266294
rect 302422 266058 302604 266294
rect 302004 229094 302604 266058
rect 302004 228858 302186 229094
rect 302422 228858 302604 229094
rect 302004 191894 302604 228858
rect 302004 191658 302186 191894
rect 302422 191658 302604 191894
rect 302004 154694 302604 191658
rect 302004 154458 302186 154694
rect 302422 154458 302604 154694
rect 302004 117494 302604 154458
rect 304766 126037 304826 351867
rect 308998 165885 309058 352550
rect 335604 337094 336204 374058
rect 335604 336858 335786 337094
rect 336022 336858 336204 337094
rect 335604 299894 336204 336858
rect 335604 299658 335786 299894
rect 336022 299658 336204 299894
rect 335604 262694 336204 299658
rect 335604 262458 335786 262694
rect 336022 262458 336204 262694
rect 335604 225494 336204 262458
rect 335604 225258 335786 225494
rect 336022 225258 336204 225494
rect 335604 188294 336204 225258
rect 335604 188058 335786 188294
rect 336022 188058 336204 188294
rect 308995 165884 309061 165885
rect 308995 165820 308996 165884
rect 309060 165820 309061 165884
rect 308995 165819 309061 165820
rect 335604 151094 336204 188058
rect 335604 150858 335786 151094
rect 336022 150858 336204 151094
rect 304763 126036 304829 126037
rect 304763 125972 304764 126036
rect 304828 125972 304829 126036
rect 304763 125971 304829 125972
rect 302004 117258 302186 117494
rect 302422 117258 302604 117494
rect 301635 86188 301701 86189
rect 301635 86124 301636 86188
rect 301700 86124 301701 86188
rect 301635 86123 301701 86124
rect 298404 76458 298586 76694
rect 298822 76458 299004 76694
rect 298404 39494 299004 76458
rect 298404 39258 298586 39494
rect 298822 39258 299004 39494
rect 295195 6628 295261 6629
rect 295195 6564 295196 6628
rect 295260 6564 295261 6628
rect 295195 6563 295261 6564
rect 264804 5658 264986 5894
rect 265222 5658 265404 5894
rect 264804 -1746 265404 5658
rect 264804 -1982 264986 -1746
rect 265222 -1982 265404 -1746
rect 264804 -2164 265404 -1982
rect 298404 2294 299004 39258
rect 298404 2058 298586 2294
rect 298822 2058 299004 2294
rect 298404 -806 299004 2058
rect 298404 -1042 298586 -806
rect 298822 -1042 299004 -806
rect 298404 -2164 299004 -1042
rect 302004 80294 302604 117258
rect 302004 80058 302186 80294
rect 302422 80058 302604 80294
rect 302004 43094 302604 80058
rect 302004 42858 302186 43094
rect 302422 42858 302604 43094
rect 302004 5894 302604 42858
rect 302004 5658 302186 5894
rect 302422 5658 302604 5894
rect 302004 -1746 302604 5658
rect 302004 -1982 302186 -1746
rect 302422 -1982 302604 -1746
rect 302004 -2164 302604 -1982
rect 335604 113894 336204 150858
rect 335604 113658 335786 113894
rect 336022 113658 336204 113894
rect 335604 76694 336204 113658
rect 335604 76458 335786 76694
rect 336022 76458 336204 76694
rect 335604 39494 336204 76458
rect 335604 39258 335786 39494
rect 336022 39258 336204 39494
rect 335604 2294 336204 39258
rect 335604 2058 335786 2294
rect 336022 2058 336204 2294
rect 335604 -806 336204 2058
rect 335604 -1042 335786 -806
rect 336022 -1042 336204 -806
rect 335604 -2164 336204 -1042
rect 339204 705918 339804 706100
rect 339204 705682 339386 705918
rect 339622 705682 339804 705918
rect 339204 675494 339804 705682
rect 339204 675258 339386 675494
rect 339622 675258 339804 675494
rect 339204 638294 339804 675258
rect 339204 638058 339386 638294
rect 339622 638058 339804 638294
rect 339204 601094 339804 638058
rect 339204 600858 339386 601094
rect 339622 600858 339804 601094
rect 339204 563894 339804 600858
rect 339204 563658 339386 563894
rect 339622 563658 339804 563894
rect 339204 526694 339804 563658
rect 339204 526458 339386 526694
rect 339622 526458 339804 526694
rect 339204 489494 339804 526458
rect 339204 489258 339386 489494
rect 339622 489258 339804 489494
rect 339204 452294 339804 489258
rect 339204 452058 339386 452294
rect 339622 452058 339804 452294
rect 339204 415094 339804 452058
rect 339204 414858 339386 415094
rect 339622 414858 339804 415094
rect 339204 377894 339804 414858
rect 339204 377658 339386 377894
rect 339622 377658 339804 377894
rect 339204 340694 339804 377658
rect 339204 340458 339386 340694
rect 339622 340458 339804 340694
rect 339204 303494 339804 340458
rect 339204 303258 339386 303494
rect 339622 303258 339804 303494
rect 339204 266294 339804 303258
rect 339204 266058 339386 266294
rect 339622 266058 339804 266294
rect 339204 229094 339804 266058
rect 339204 228858 339386 229094
rect 339622 228858 339804 229094
rect 339204 191894 339804 228858
rect 339204 191658 339386 191894
rect 339622 191658 339804 191894
rect 339204 154694 339804 191658
rect 339204 154458 339386 154694
rect 339622 154458 339804 154694
rect 339204 117494 339804 154458
rect 339204 117258 339386 117494
rect 339622 117258 339804 117494
rect 339204 80294 339804 117258
rect 339204 80058 339386 80294
rect 339622 80058 339804 80294
rect 339204 43094 339804 80058
rect 339204 42858 339386 43094
rect 339622 42858 339804 43094
rect 339204 5894 339804 42858
rect 339204 5658 339386 5894
rect 339622 5658 339804 5894
rect 339204 -1746 339804 5658
rect 339204 -1982 339386 -1746
rect 339622 -1982 339804 -1746
rect 339204 -2164 339804 -1982
rect 372804 704978 373404 706100
rect 372804 704742 372986 704978
rect 373222 704742 373404 704978
rect 372804 671894 373404 704742
rect 372804 671658 372986 671894
rect 373222 671658 373404 671894
rect 372804 634694 373404 671658
rect 372804 634458 372986 634694
rect 373222 634458 373404 634694
rect 372804 597494 373404 634458
rect 372804 597258 372986 597494
rect 373222 597258 373404 597494
rect 372804 560294 373404 597258
rect 372804 560058 372986 560294
rect 373222 560058 373404 560294
rect 372804 523094 373404 560058
rect 372804 522858 372986 523094
rect 373222 522858 373404 523094
rect 372804 485894 373404 522858
rect 372804 485658 372986 485894
rect 373222 485658 373404 485894
rect 372804 448694 373404 485658
rect 372804 448458 372986 448694
rect 373222 448458 373404 448694
rect 372804 411494 373404 448458
rect 372804 411258 372986 411494
rect 373222 411258 373404 411494
rect 372804 374294 373404 411258
rect 372804 374058 372986 374294
rect 373222 374058 373404 374294
rect 372804 337094 373404 374058
rect 372804 336858 372986 337094
rect 373222 336858 373404 337094
rect 372804 299894 373404 336858
rect 372804 299658 372986 299894
rect 373222 299658 373404 299894
rect 372804 262694 373404 299658
rect 372804 262458 372986 262694
rect 373222 262458 373404 262694
rect 372804 225494 373404 262458
rect 372804 225258 372986 225494
rect 373222 225258 373404 225494
rect 372804 188294 373404 225258
rect 372804 188058 372986 188294
rect 373222 188058 373404 188294
rect 372804 151094 373404 188058
rect 372804 150858 372986 151094
rect 373222 150858 373404 151094
rect 372804 113894 373404 150858
rect 372804 113658 372986 113894
rect 373222 113658 373404 113894
rect 372804 76694 373404 113658
rect 372804 76458 372986 76694
rect 373222 76458 373404 76694
rect 372804 39494 373404 76458
rect 372804 39258 372986 39494
rect 373222 39258 373404 39494
rect 372804 2294 373404 39258
rect 372804 2058 372986 2294
rect 373222 2058 373404 2294
rect 372804 -806 373404 2058
rect 372804 -1042 372986 -806
rect 373222 -1042 373404 -806
rect 372804 -2164 373404 -1042
rect 376404 705918 377004 706100
rect 376404 705682 376586 705918
rect 376822 705682 377004 705918
rect 376404 675494 377004 705682
rect 376404 675258 376586 675494
rect 376822 675258 377004 675494
rect 376404 638294 377004 675258
rect 376404 638058 376586 638294
rect 376822 638058 377004 638294
rect 376404 601094 377004 638058
rect 376404 600858 376586 601094
rect 376822 600858 377004 601094
rect 376404 563894 377004 600858
rect 376404 563658 376586 563894
rect 376822 563658 377004 563894
rect 376404 526694 377004 563658
rect 376404 526458 376586 526694
rect 376822 526458 377004 526694
rect 376404 489494 377004 526458
rect 376404 489258 376586 489494
rect 376822 489258 377004 489494
rect 376404 452294 377004 489258
rect 376404 452058 376586 452294
rect 376822 452058 377004 452294
rect 376404 415094 377004 452058
rect 376404 414858 376586 415094
rect 376822 414858 377004 415094
rect 376404 377894 377004 414858
rect 376404 377658 376586 377894
rect 376822 377658 377004 377894
rect 376404 340694 377004 377658
rect 376404 340458 376586 340694
rect 376822 340458 377004 340694
rect 376404 303494 377004 340458
rect 376404 303258 376586 303494
rect 376822 303258 377004 303494
rect 376404 266294 377004 303258
rect 376404 266058 376586 266294
rect 376822 266058 377004 266294
rect 376404 229094 377004 266058
rect 376404 228858 376586 229094
rect 376822 228858 377004 229094
rect 376404 191894 377004 228858
rect 376404 191658 376586 191894
rect 376822 191658 377004 191894
rect 376404 154694 377004 191658
rect 376404 154458 376586 154694
rect 376822 154458 377004 154694
rect 376404 117494 377004 154458
rect 376404 117258 376586 117494
rect 376822 117258 377004 117494
rect 376404 80294 377004 117258
rect 376404 80058 376586 80294
rect 376822 80058 377004 80294
rect 376404 43094 377004 80058
rect 376404 42858 376586 43094
rect 376822 42858 377004 43094
rect 376404 5894 377004 42858
rect 376404 5658 376586 5894
rect 376822 5658 377004 5894
rect 376404 -1746 377004 5658
rect 376404 -1982 376586 -1746
rect 376822 -1982 377004 -1746
rect 376404 -2164 377004 -1982
rect 410004 704978 410604 706100
rect 410004 704742 410186 704978
rect 410422 704742 410604 704978
rect 410004 671894 410604 704742
rect 410004 671658 410186 671894
rect 410422 671658 410604 671894
rect 410004 634694 410604 671658
rect 410004 634458 410186 634694
rect 410422 634458 410604 634694
rect 410004 597494 410604 634458
rect 410004 597258 410186 597494
rect 410422 597258 410604 597494
rect 410004 560294 410604 597258
rect 410004 560058 410186 560294
rect 410422 560058 410604 560294
rect 410004 523094 410604 560058
rect 410004 522858 410186 523094
rect 410422 522858 410604 523094
rect 410004 485894 410604 522858
rect 410004 485658 410186 485894
rect 410422 485658 410604 485894
rect 410004 448694 410604 485658
rect 410004 448458 410186 448694
rect 410422 448458 410604 448694
rect 410004 411494 410604 448458
rect 410004 411258 410186 411494
rect 410422 411258 410604 411494
rect 410004 374294 410604 411258
rect 410004 374058 410186 374294
rect 410422 374058 410604 374294
rect 410004 337094 410604 374058
rect 410004 336858 410186 337094
rect 410422 336858 410604 337094
rect 410004 299894 410604 336858
rect 410004 299658 410186 299894
rect 410422 299658 410604 299894
rect 410004 262694 410604 299658
rect 410004 262458 410186 262694
rect 410422 262458 410604 262694
rect 410004 225494 410604 262458
rect 410004 225258 410186 225494
rect 410422 225258 410604 225494
rect 410004 188294 410604 225258
rect 410004 188058 410186 188294
rect 410422 188058 410604 188294
rect 410004 151094 410604 188058
rect 410004 150858 410186 151094
rect 410422 150858 410604 151094
rect 410004 113894 410604 150858
rect 410004 113658 410186 113894
rect 410422 113658 410604 113894
rect 410004 76694 410604 113658
rect 410004 76458 410186 76694
rect 410422 76458 410604 76694
rect 410004 39494 410604 76458
rect 410004 39258 410186 39494
rect 410422 39258 410604 39494
rect 410004 2294 410604 39258
rect 410004 2058 410186 2294
rect 410422 2058 410604 2294
rect 410004 -806 410604 2058
rect 410004 -1042 410186 -806
rect 410422 -1042 410604 -806
rect 410004 -2164 410604 -1042
rect 413604 705918 414204 706100
rect 413604 705682 413786 705918
rect 414022 705682 414204 705918
rect 413604 675494 414204 705682
rect 413604 675258 413786 675494
rect 414022 675258 414204 675494
rect 413604 638294 414204 675258
rect 413604 638058 413786 638294
rect 414022 638058 414204 638294
rect 413604 601094 414204 638058
rect 413604 600858 413786 601094
rect 414022 600858 414204 601094
rect 413604 563894 414204 600858
rect 413604 563658 413786 563894
rect 414022 563658 414204 563894
rect 413604 526694 414204 563658
rect 413604 526458 413786 526694
rect 414022 526458 414204 526694
rect 413604 489494 414204 526458
rect 413604 489258 413786 489494
rect 414022 489258 414204 489494
rect 413604 452294 414204 489258
rect 413604 452058 413786 452294
rect 414022 452058 414204 452294
rect 413604 415094 414204 452058
rect 413604 414858 413786 415094
rect 414022 414858 414204 415094
rect 413604 377894 414204 414858
rect 413604 377658 413786 377894
rect 414022 377658 414204 377894
rect 413604 340694 414204 377658
rect 413604 340458 413786 340694
rect 414022 340458 414204 340694
rect 413604 303494 414204 340458
rect 413604 303258 413786 303494
rect 414022 303258 414204 303494
rect 413604 266294 414204 303258
rect 413604 266058 413786 266294
rect 414022 266058 414204 266294
rect 413604 229094 414204 266058
rect 413604 228858 413786 229094
rect 414022 228858 414204 229094
rect 413604 191894 414204 228858
rect 413604 191658 413786 191894
rect 414022 191658 414204 191894
rect 413604 154694 414204 191658
rect 413604 154458 413786 154694
rect 414022 154458 414204 154694
rect 413604 117494 414204 154458
rect 413604 117258 413786 117494
rect 414022 117258 414204 117494
rect 413604 80294 414204 117258
rect 413604 80058 413786 80294
rect 414022 80058 414204 80294
rect 413604 43094 414204 80058
rect 413604 42858 413786 43094
rect 414022 42858 414204 43094
rect 413604 5894 414204 42858
rect 413604 5658 413786 5894
rect 414022 5658 414204 5894
rect 413604 -1746 414204 5658
rect 413604 -1982 413786 -1746
rect 414022 -1982 414204 -1746
rect 413604 -2164 414204 -1982
rect 447204 704978 447804 706100
rect 447204 704742 447386 704978
rect 447622 704742 447804 704978
rect 447204 671894 447804 704742
rect 447204 671658 447386 671894
rect 447622 671658 447804 671894
rect 447204 634694 447804 671658
rect 447204 634458 447386 634694
rect 447622 634458 447804 634694
rect 447204 597494 447804 634458
rect 447204 597258 447386 597494
rect 447622 597258 447804 597494
rect 447204 560294 447804 597258
rect 447204 560058 447386 560294
rect 447622 560058 447804 560294
rect 447204 523094 447804 560058
rect 447204 522858 447386 523094
rect 447622 522858 447804 523094
rect 447204 485894 447804 522858
rect 447204 485658 447386 485894
rect 447622 485658 447804 485894
rect 447204 448694 447804 485658
rect 447204 448458 447386 448694
rect 447622 448458 447804 448694
rect 447204 411494 447804 448458
rect 447204 411258 447386 411494
rect 447622 411258 447804 411494
rect 447204 374294 447804 411258
rect 447204 374058 447386 374294
rect 447622 374058 447804 374294
rect 447204 337094 447804 374058
rect 447204 336858 447386 337094
rect 447622 336858 447804 337094
rect 447204 299894 447804 336858
rect 447204 299658 447386 299894
rect 447622 299658 447804 299894
rect 447204 262694 447804 299658
rect 447204 262458 447386 262694
rect 447622 262458 447804 262694
rect 447204 225494 447804 262458
rect 447204 225258 447386 225494
rect 447622 225258 447804 225494
rect 447204 188294 447804 225258
rect 447204 188058 447386 188294
rect 447622 188058 447804 188294
rect 447204 151094 447804 188058
rect 447204 150858 447386 151094
rect 447622 150858 447804 151094
rect 447204 113894 447804 150858
rect 447204 113658 447386 113894
rect 447622 113658 447804 113894
rect 447204 76694 447804 113658
rect 447204 76458 447386 76694
rect 447622 76458 447804 76694
rect 447204 39494 447804 76458
rect 447204 39258 447386 39494
rect 447622 39258 447804 39494
rect 447204 2294 447804 39258
rect 447204 2058 447386 2294
rect 447622 2058 447804 2294
rect 447204 -806 447804 2058
rect 447204 -1042 447386 -806
rect 447622 -1042 447804 -806
rect 447204 -2164 447804 -1042
rect 450804 705918 451404 706100
rect 450804 705682 450986 705918
rect 451222 705682 451404 705918
rect 450804 675494 451404 705682
rect 450804 675258 450986 675494
rect 451222 675258 451404 675494
rect 450804 638294 451404 675258
rect 450804 638058 450986 638294
rect 451222 638058 451404 638294
rect 450804 601094 451404 638058
rect 450804 600858 450986 601094
rect 451222 600858 451404 601094
rect 450804 563894 451404 600858
rect 450804 563658 450986 563894
rect 451222 563658 451404 563894
rect 450804 526694 451404 563658
rect 450804 526458 450986 526694
rect 451222 526458 451404 526694
rect 450804 489494 451404 526458
rect 450804 489258 450986 489494
rect 451222 489258 451404 489494
rect 450804 452294 451404 489258
rect 450804 452058 450986 452294
rect 451222 452058 451404 452294
rect 450804 415094 451404 452058
rect 450804 414858 450986 415094
rect 451222 414858 451404 415094
rect 450804 377894 451404 414858
rect 450804 377658 450986 377894
rect 451222 377658 451404 377894
rect 450804 340694 451404 377658
rect 450804 340458 450986 340694
rect 451222 340458 451404 340694
rect 450804 303494 451404 340458
rect 450804 303258 450986 303494
rect 451222 303258 451404 303494
rect 450804 266294 451404 303258
rect 450804 266058 450986 266294
rect 451222 266058 451404 266294
rect 450804 229094 451404 266058
rect 450804 228858 450986 229094
rect 451222 228858 451404 229094
rect 450804 191894 451404 228858
rect 450804 191658 450986 191894
rect 451222 191658 451404 191894
rect 450804 154694 451404 191658
rect 450804 154458 450986 154694
rect 451222 154458 451404 154694
rect 450804 117494 451404 154458
rect 450804 117258 450986 117494
rect 451222 117258 451404 117494
rect 450804 80294 451404 117258
rect 450804 80058 450986 80294
rect 451222 80058 451404 80294
rect 450804 43094 451404 80058
rect 450804 42858 450986 43094
rect 451222 42858 451404 43094
rect 450804 5894 451404 42858
rect 450804 5658 450986 5894
rect 451222 5658 451404 5894
rect 450804 -1746 451404 5658
rect 450804 -1982 450986 -1746
rect 451222 -1982 451404 -1746
rect 450804 -2164 451404 -1982
rect 484404 704978 485004 706100
rect 484404 704742 484586 704978
rect 484822 704742 485004 704978
rect 484404 671894 485004 704742
rect 484404 671658 484586 671894
rect 484822 671658 485004 671894
rect 484404 634694 485004 671658
rect 484404 634458 484586 634694
rect 484822 634458 485004 634694
rect 484404 597494 485004 634458
rect 484404 597258 484586 597494
rect 484822 597258 485004 597494
rect 484404 560294 485004 597258
rect 484404 560058 484586 560294
rect 484822 560058 485004 560294
rect 484404 523094 485004 560058
rect 484404 522858 484586 523094
rect 484822 522858 485004 523094
rect 484404 485894 485004 522858
rect 484404 485658 484586 485894
rect 484822 485658 485004 485894
rect 484404 448694 485004 485658
rect 484404 448458 484586 448694
rect 484822 448458 485004 448694
rect 484404 411494 485004 448458
rect 484404 411258 484586 411494
rect 484822 411258 485004 411494
rect 484404 374294 485004 411258
rect 484404 374058 484586 374294
rect 484822 374058 485004 374294
rect 484404 337094 485004 374058
rect 484404 336858 484586 337094
rect 484822 336858 485004 337094
rect 484404 299894 485004 336858
rect 484404 299658 484586 299894
rect 484822 299658 485004 299894
rect 484404 262694 485004 299658
rect 484404 262458 484586 262694
rect 484822 262458 485004 262694
rect 484404 225494 485004 262458
rect 484404 225258 484586 225494
rect 484822 225258 485004 225494
rect 484404 188294 485004 225258
rect 484404 188058 484586 188294
rect 484822 188058 485004 188294
rect 484404 151094 485004 188058
rect 484404 150858 484586 151094
rect 484822 150858 485004 151094
rect 484404 113894 485004 150858
rect 484404 113658 484586 113894
rect 484822 113658 485004 113894
rect 484404 76694 485004 113658
rect 484404 76458 484586 76694
rect 484822 76458 485004 76694
rect 484404 39494 485004 76458
rect 484404 39258 484586 39494
rect 484822 39258 485004 39494
rect 484404 2294 485004 39258
rect 484404 2058 484586 2294
rect 484822 2058 485004 2294
rect 484404 -806 485004 2058
rect 484404 -1042 484586 -806
rect 484822 -1042 485004 -806
rect 484404 -2164 485004 -1042
rect 488004 705918 488604 706100
rect 488004 705682 488186 705918
rect 488422 705682 488604 705918
rect 488004 675494 488604 705682
rect 488004 675258 488186 675494
rect 488422 675258 488604 675494
rect 488004 638294 488604 675258
rect 488004 638058 488186 638294
rect 488422 638058 488604 638294
rect 488004 601094 488604 638058
rect 488004 600858 488186 601094
rect 488422 600858 488604 601094
rect 488004 563894 488604 600858
rect 488004 563658 488186 563894
rect 488422 563658 488604 563894
rect 488004 526694 488604 563658
rect 488004 526458 488186 526694
rect 488422 526458 488604 526694
rect 488004 489494 488604 526458
rect 488004 489258 488186 489494
rect 488422 489258 488604 489494
rect 488004 452294 488604 489258
rect 488004 452058 488186 452294
rect 488422 452058 488604 452294
rect 488004 415094 488604 452058
rect 488004 414858 488186 415094
rect 488422 414858 488604 415094
rect 488004 377894 488604 414858
rect 488004 377658 488186 377894
rect 488422 377658 488604 377894
rect 488004 340694 488604 377658
rect 521604 704978 522204 706100
rect 521604 704742 521786 704978
rect 522022 704742 522204 704978
rect 521604 671894 522204 704742
rect 521604 671658 521786 671894
rect 522022 671658 522204 671894
rect 521604 634694 522204 671658
rect 521604 634458 521786 634694
rect 522022 634458 522204 634694
rect 521604 597494 522204 634458
rect 521604 597258 521786 597494
rect 522022 597258 522204 597494
rect 521604 560294 522204 597258
rect 521604 560058 521786 560294
rect 522022 560058 522204 560294
rect 521604 523094 522204 560058
rect 521604 522858 521786 523094
rect 522022 522858 522204 523094
rect 521604 485894 522204 522858
rect 521604 485658 521786 485894
rect 522022 485658 522204 485894
rect 521604 448694 522204 485658
rect 521604 448458 521786 448694
rect 522022 448458 522204 448694
rect 521604 411494 522204 448458
rect 521604 411258 521786 411494
rect 522022 411258 522204 411494
rect 521604 374294 522204 411258
rect 521604 374058 521786 374294
rect 522022 374058 522204 374294
rect 521604 341752 522204 374058
rect 525204 705918 525804 706100
rect 525204 705682 525386 705918
rect 525622 705682 525804 705918
rect 525204 675494 525804 705682
rect 525204 675258 525386 675494
rect 525622 675258 525804 675494
rect 525204 638294 525804 675258
rect 525204 638058 525386 638294
rect 525622 638058 525804 638294
rect 525204 601094 525804 638058
rect 525204 600858 525386 601094
rect 525622 600858 525804 601094
rect 525204 563894 525804 600858
rect 525204 563658 525386 563894
rect 525622 563658 525804 563894
rect 525204 526694 525804 563658
rect 525204 526458 525386 526694
rect 525622 526458 525804 526694
rect 525204 489494 525804 526458
rect 525204 489258 525386 489494
rect 525622 489258 525804 489494
rect 525204 452294 525804 489258
rect 525204 452058 525386 452294
rect 525622 452058 525804 452294
rect 525204 415094 525804 452058
rect 525204 414858 525386 415094
rect 525622 414858 525804 415094
rect 525204 377894 525804 414858
rect 525204 377658 525386 377894
rect 525622 377658 525804 377894
rect 525204 341752 525804 377658
rect 558804 704978 559404 706100
rect 558804 704742 558986 704978
rect 559222 704742 559404 704978
rect 558804 671894 559404 704742
rect 558804 671658 558986 671894
rect 559222 671658 559404 671894
rect 558804 634694 559404 671658
rect 558804 634458 558986 634694
rect 559222 634458 559404 634694
rect 558804 597494 559404 634458
rect 558804 597258 558986 597494
rect 559222 597258 559404 597494
rect 558804 560294 559404 597258
rect 558804 560058 558986 560294
rect 559222 560058 559404 560294
rect 558804 523094 559404 560058
rect 558804 522858 558986 523094
rect 559222 522858 559404 523094
rect 558804 485894 559404 522858
rect 558804 485658 558986 485894
rect 559222 485658 559404 485894
rect 558804 448694 559404 485658
rect 558804 448458 558986 448694
rect 559222 448458 559404 448694
rect 558804 411494 559404 448458
rect 558804 411258 558986 411494
rect 559222 411258 559404 411494
rect 558804 374294 559404 411258
rect 558804 374058 558986 374294
rect 559222 374058 559404 374294
rect 488004 340458 488186 340694
rect 488422 340458 488604 340694
rect 488004 303494 488604 340458
rect 521910 337094 522230 337276
rect 521910 336858 521952 337094
rect 522188 336858 522230 337094
rect 521910 336676 522230 336858
rect 523842 337094 524162 337276
rect 523842 336858 523884 337094
rect 524120 336858 524162 337094
rect 523842 336676 524162 336858
rect 525774 337094 526094 337276
rect 525774 336858 525816 337094
rect 526052 336858 526094 337094
rect 525774 336676 526094 336858
rect 527706 337094 528026 337276
rect 527706 336858 527748 337094
rect 527984 336858 528026 337094
rect 527706 336676 528026 336858
rect 558804 337094 559404 374058
rect 558804 336858 558986 337094
rect 559222 336858 559404 337094
rect 531819 330988 531885 330989
rect 531819 330924 531820 330988
rect 531884 330924 531885 330988
rect 531819 330923 531885 330924
rect 488004 303258 488186 303494
rect 488422 303258 488604 303494
rect 488004 266294 488604 303258
rect 488004 266058 488186 266294
rect 488422 266058 488604 266294
rect 488004 229094 488604 266058
rect 488004 228858 488186 229094
rect 488422 228858 488604 229094
rect 488004 191894 488604 228858
rect 488004 191658 488186 191894
rect 488422 191658 488604 191894
rect 488004 154694 488604 191658
rect 488004 154458 488186 154694
rect 488422 154458 488604 154694
rect 488004 117494 488604 154458
rect 488004 117258 488186 117494
rect 488422 117258 488604 117494
rect 488004 80294 488604 117258
rect 488004 80058 488186 80294
rect 488422 80058 488604 80294
rect 488004 43094 488604 80058
rect 488004 42858 488186 43094
rect 488422 42858 488604 43094
rect 488004 5894 488604 42858
rect 488004 5658 488186 5894
rect 488422 5658 488604 5894
rect 488004 -1746 488604 5658
rect 488004 -1982 488186 -1746
rect 488422 -1982 488604 -1746
rect 488004 -2164 488604 -1982
rect 521604 299894 522204 320008
rect 521604 299658 521786 299894
rect 522022 299658 522204 299894
rect 521604 262694 522204 299658
rect 521604 262458 521786 262694
rect 522022 262458 522204 262694
rect 521604 225494 522204 262458
rect 521604 225258 521786 225494
rect 522022 225258 522204 225494
rect 521604 188294 522204 225258
rect 521604 188058 521786 188294
rect 522022 188058 522204 188294
rect 521604 151094 522204 188058
rect 521604 150858 521786 151094
rect 522022 150858 522204 151094
rect 521604 113894 522204 150858
rect 521604 113658 521786 113894
rect 522022 113658 522204 113894
rect 521604 76694 522204 113658
rect 521604 76458 521786 76694
rect 522022 76458 522204 76694
rect 521604 39494 522204 76458
rect 521604 39258 521786 39494
rect 522022 39258 522204 39494
rect 521604 2294 522204 39258
rect 521604 2058 521786 2294
rect 522022 2058 522204 2294
rect 521604 -806 522204 2058
rect 521604 -1042 521786 -806
rect 522022 -1042 522204 -806
rect 521604 -2164 522204 -1042
rect 525204 303494 525804 320008
rect 525204 303258 525386 303494
rect 525622 303258 525804 303494
rect 525204 266294 525804 303258
rect 525204 266058 525386 266294
rect 525622 266058 525804 266294
rect 525204 229094 525804 266058
rect 525204 228858 525386 229094
rect 525622 228858 525804 229094
rect 525204 191894 525804 228858
rect 525204 191658 525386 191894
rect 525622 191658 525804 191894
rect 525204 154694 525804 191658
rect 525204 154458 525386 154694
rect 525622 154458 525804 154694
rect 525204 117494 525804 154458
rect 525204 117258 525386 117494
rect 525622 117258 525804 117494
rect 525204 80294 525804 117258
rect 525204 80058 525386 80294
rect 525622 80058 525804 80294
rect 525204 43094 525804 80058
rect 525204 42858 525386 43094
rect 525622 42858 525804 43094
rect 525204 5894 525804 42858
rect 531822 19821 531882 330923
rect 558804 299894 559404 336858
rect 558804 299658 558986 299894
rect 559222 299658 559404 299894
rect 558804 262694 559404 299658
rect 558804 262458 558986 262694
rect 559222 262458 559404 262694
rect 558804 225494 559404 262458
rect 558804 225258 558986 225494
rect 559222 225258 559404 225494
rect 558804 188294 559404 225258
rect 558804 188058 558986 188294
rect 559222 188058 559404 188294
rect 558804 151094 559404 188058
rect 558804 150858 558986 151094
rect 559222 150858 559404 151094
rect 558804 113894 559404 150858
rect 558804 113658 558986 113894
rect 559222 113658 559404 113894
rect 558804 76694 559404 113658
rect 558804 76458 558986 76694
rect 559222 76458 559404 76694
rect 558804 39494 559404 76458
rect 558804 39258 558986 39494
rect 559222 39258 559404 39494
rect 531819 19820 531885 19821
rect 531819 19756 531820 19820
rect 531884 19756 531885 19820
rect 531819 19755 531885 19756
rect 525204 5658 525386 5894
rect 525622 5658 525804 5894
rect 525204 -1746 525804 5658
rect 525204 -1982 525386 -1746
rect 525622 -1982 525804 -1746
rect 525204 -2164 525804 -1982
rect 558804 2294 559404 39258
rect 558804 2058 558986 2294
rect 559222 2058 559404 2294
rect 558804 -806 559404 2058
rect 558804 -1042 558986 -806
rect 559222 -1042 559404 -806
rect 558804 -2164 559404 -1042
rect 562404 705918 563004 706100
rect 562404 705682 562586 705918
rect 562822 705682 563004 705918
rect 562404 675494 563004 705682
rect 586560 705918 587160 706100
rect 586560 705682 586742 705918
rect 586978 705682 587160 705918
rect 562404 675258 562586 675494
rect 562822 675258 563004 675494
rect 562404 638294 563004 675258
rect 562404 638058 562586 638294
rect 562822 638058 563004 638294
rect 562404 601094 563004 638058
rect 562404 600858 562586 601094
rect 562822 600858 563004 601094
rect 562404 563894 563004 600858
rect 562404 563658 562586 563894
rect 562822 563658 563004 563894
rect 562404 526694 563004 563658
rect 562404 526458 562586 526694
rect 562822 526458 563004 526694
rect 562404 489494 563004 526458
rect 562404 489258 562586 489494
rect 562822 489258 563004 489494
rect 562404 452294 563004 489258
rect 562404 452058 562586 452294
rect 562822 452058 563004 452294
rect 562404 415094 563004 452058
rect 562404 414858 562586 415094
rect 562822 414858 563004 415094
rect 562404 377894 563004 414858
rect 562404 377658 562586 377894
rect 562822 377658 563004 377894
rect 562404 340694 563004 377658
rect 562404 340458 562586 340694
rect 562822 340458 563004 340694
rect 562404 303494 563004 340458
rect 562404 303258 562586 303494
rect 562822 303258 563004 303494
rect 562404 266294 563004 303258
rect 562404 266058 562586 266294
rect 562822 266058 563004 266294
rect 562404 229094 563004 266058
rect 562404 228858 562586 229094
rect 562822 228858 563004 229094
rect 562404 191894 563004 228858
rect 562404 191658 562586 191894
rect 562822 191658 563004 191894
rect 562404 154694 563004 191658
rect 562404 154458 562586 154694
rect 562822 154458 563004 154694
rect 562404 117494 563004 154458
rect 562404 117258 562586 117494
rect 562822 117258 563004 117494
rect 562404 80294 563004 117258
rect 562404 80058 562586 80294
rect 562822 80058 563004 80294
rect 562404 43094 563004 80058
rect 562404 42858 562586 43094
rect 562822 42858 563004 43094
rect 562404 5894 563004 42858
rect 562404 5658 562586 5894
rect 562822 5658 563004 5894
rect 562404 -1746 563004 5658
rect 585620 704978 586220 705160
rect 585620 704742 585802 704978
rect 586038 704742 586220 704978
rect 585620 671894 586220 704742
rect 585620 671658 585802 671894
rect 586038 671658 586220 671894
rect 585620 634694 586220 671658
rect 585620 634458 585802 634694
rect 586038 634458 586220 634694
rect 585620 597494 586220 634458
rect 585620 597258 585802 597494
rect 586038 597258 586220 597494
rect 585620 560294 586220 597258
rect 585620 560058 585802 560294
rect 586038 560058 586220 560294
rect 585620 523094 586220 560058
rect 585620 522858 585802 523094
rect 586038 522858 586220 523094
rect 585620 485894 586220 522858
rect 585620 485658 585802 485894
rect 586038 485658 586220 485894
rect 585620 448694 586220 485658
rect 585620 448458 585802 448694
rect 586038 448458 586220 448694
rect 585620 411494 586220 448458
rect 585620 411258 585802 411494
rect 586038 411258 586220 411494
rect 585620 374294 586220 411258
rect 585620 374058 585802 374294
rect 586038 374058 586220 374294
rect 585620 337094 586220 374058
rect 585620 336858 585802 337094
rect 586038 336858 586220 337094
rect 585620 299894 586220 336858
rect 585620 299658 585802 299894
rect 586038 299658 586220 299894
rect 585620 262694 586220 299658
rect 585620 262458 585802 262694
rect 586038 262458 586220 262694
rect 585620 225494 586220 262458
rect 585620 225258 585802 225494
rect 586038 225258 586220 225494
rect 585620 188294 586220 225258
rect 585620 188058 585802 188294
rect 586038 188058 586220 188294
rect 585620 151094 586220 188058
rect 585620 150858 585802 151094
rect 586038 150858 586220 151094
rect 585620 113894 586220 150858
rect 585620 113658 585802 113894
rect 586038 113658 586220 113894
rect 585620 76694 586220 113658
rect 585620 76458 585802 76694
rect 586038 76458 586220 76694
rect 585620 39494 586220 76458
rect 585620 39258 585802 39494
rect 586038 39258 586220 39494
rect 585620 2294 586220 39258
rect 585620 2058 585802 2294
rect 586038 2058 586220 2294
rect 585620 -806 586220 2058
rect 585620 -1042 585802 -806
rect 586038 -1042 586220 -806
rect 585620 -1224 586220 -1042
rect 586560 675494 587160 705682
rect 586560 675258 586742 675494
rect 586978 675258 587160 675494
rect 586560 638294 587160 675258
rect 586560 638058 586742 638294
rect 586978 638058 587160 638294
rect 586560 601094 587160 638058
rect 586560 600858 586742 601094
rect 586978 600858 587160 601094
rect 586560 563894 587160 600858
rect 586560 563658 586742 563894
rect 586978 563658 587160 563894
rect 586560 526694 587160 563658
rect 586560 526458 586742 526694
rect 586978 526458 587160 526694
rect 586560 489494 587160 526458
rect 586560 489258 586742 489494
rect 586978 489258 587160 489494
rect 586560 452294 587160 489258
rect 586560 452058 586742 452294
rect 586978 452058 587160 452294
rect 586560 415094 587160 452058
rect 586560 414858 586742 415094
rect 586978 414858 587160 415094
rect 586560 377894 587160 414858
rect 586560 377658 586742 377894
rect 586978 377658 587160 377894
rect 586560 340694 587160 377658
rect 586560 340458 586742 340694
rect 586978 340458 587160 340694
rect 586560 303494 587160 340458
rect 586560 303258 586742 303494
rect 586978 303258 587160 303494
rect 586560 266294 587160 303258
rect 586560 266058 586742 266294
rect 586978 266058 587160 266294
rect 586560 229094 587160 266058
rect 586560 228858 586742 229094
rect 586978 228858 587160 229094
rect 586560 191894 587160 228858
rect 586560 191658 586742 191894
rect 586978 191658 587160 191894
rect 586560 154694 587160 191658
rect 586560 154458 586742 154694
rect 586978 154458 587160 154694
rect 586560 117494 587160 154458
rect 586560 117258 586742 117494
rect 586978 117258 587160 117494
rect 586560 80294 587160 117258
rect 586560 80058 586742 80294
rect 586978 80058 587160 80294
rect 586560 43094 587160 80058
rect 586560 42858 586742 43094
rect 586978 42858 587160 43094
rect 586560 5894 587160 42858
rect 586560 5658 586742 5894
rect 586978 5658 587160 5894
rect 562404 -1982 562586 -1746
rect 562822 -1982 563004 -1746
rect 562404 -2164 563004 -1982
rect 586560 -1746 587160 5658
rect 586560 -1982 586742 -1746
rect 586978 -1982 587160 -1746
rect 586560 -2164 587160 -1982
<< via4 >>
rect -3054 705682 -2818 705918
rect -3054 675258 -2818 675494
rect -3054 638058 -2818 638294
rect -3054 600858 -2818 601094
rect -3054 563658 -2818 563894
rect -3054 526458 -2818 526694
rect -3054 489258 -2818 489494
rect -3054 452058 -2818 452294
rect -3054 414858 -2818 415094
rect -3054 377658 -2818 377894
rect -3054 340458 -2818 340694
rect -3054 303258 -2818 303494
rect -3054 266058 -2818 266294
rect -3054 228858 -2818 229094
rect -3054 191658 -2818 191894
rect -3054 154458 -2818 154694
rect -3054 117258 -2818 117494
rect -3054 80058 -2818 80294
rect -3054 42858 -2818 43094
rect -3054 5658 -2818 5894
rect -2114 704742 -1878 704978
rect -2114 671658 -1878 671894
rect -2114 634458 -1878 634694
rect -2114 597258 -1878 597494
rect -2114 560058 -1878 560294
rect -2114 522858 -1878 523094
rect -2114 485658 -1878 485894
rect -2114 448458 -1878 448694
rect -2114 411258 -1878 411494
rect -2114 374058 -1878 374294
rect -2114 336858 -1878 337094
rect -2114 299658 -1878 299894
rect -2114 262458 -1878 262694
rect -2114 225258 -1878 225494
rect -2114 188058 -1878 188294
rect -2114 150858 -1878 151094
rect -2114 113658 -1878 113894
rect -2114 76458 -1878 76694
rect -2114 39258 -1878 39494
rect -2114 2058 -1878 2294
rect -2114 -1042 -1878 -806
rect 986 704742 1222 704978
rect 986 671658 1222 671894
rect 986 634458 1222 634694
rect 986 597258 1222 597494
rect 986 560058 1222 560294
rect 986 522858 1222 523094
rect 986 485658 1222 485894
rect 986 448458 1222 448694
rect 986 411258 1222 411494
rect 986 374058 1222 374294
rect 986 336858 1222 337094
rect 986 299658 1222 299894
rect 986 262458 1222 262694
rect 986 225258 1222 225494
rect 986 188058 1222 188294
rect 986 150858 1222 151094
rect 986 113658 1222 113894
rect 986 76458 1222 76694
rect 986 39258 1222 39494
rect 986 2058 1222 2294
rect 986 -1042 1222 -806
rect -3054 -1982 -2818 -1746
rect 4586 705682 4822 705918
rect 4586 675258 4822 675494
rect 4586 638058 4822 638294
rect 4586 600858 4822 601094
rect 4586 563658 4822 563894
rect 4586 526458 4822 526694
rect 4586 489258 4822 489494
rect 4586 452058 4822 452294
rect 4586 414858 4822 415094
rect 4586 377658 4822 377894
rect 4586 340458 4822 340694
rect 4586 303258 4822 303494
rect 4586 266058 4822 266294
rect 4586 228858 4822 229094
rect 4586 191658 4822 191894
rect 4586 154458 4822 154694
rect 4586 117258 4822 117494
rect 4586 80058 4822 80294
rect 4586 42858 4822 43094
rect 4586 5658 4822 5894
rect 4586 -1982 4822 -1746
rect 38186 704742 38422 704978
rect 38186 671658 38422 671894
rect 38186 634458 38422 634694
rect 38186 597258 38422 597494
rect 38186 560058 38422 560294
rect 38186 522858 38422 523094
rect 38186 485658 38422 485894
rect 38186 448458 38422 448694
rect 38186 411258 38422 411494
rect 38186 374058 38422 374294
rect 38186 336858 38422 337094
rect 38186 299658 38422 299894
rect 38186 262458 38422 262694
rect 38186 225258 38422 225494
rect 38186 188058 38422 188294
rect 38186 150858 38422 151094
rect 38186 113658 38422 113894
rect 38186 76458 38422 76694
rect 38186 39258 38422 39494
rect 38186 2058 38422 2294
rect 38186 -1042 38422 -806
rect 41786 705682 42022 705918
rect 41786 675258 42022 675494
rect 41786 638058 42022 638294
rect 41786 600858 42022 601094
rect 41786 563658 42022 563894
rect 41786 526458 42022 526694
rect 41786 489258 42022 489494
rect 41786 452058 42022 452294
rect 41786 414858 42022 415094
rect 41786 377658 42022 377894
rect 41786 340458 42022 340694
rect 41786 303258 42022 303494
rect 41786 266058 42022 266294
rect 41786 228858 42022 229094
rect 41786 191658 42022 191894
rect 41786 154458 42022 154694
rect 41786 117258 42022 117494
rect 41786 80058 42022 80294
rect 41786 42858 42022 43094
rect 41786 5658 42022 5894
rect 41786 -1982 42022 -1746
rect 75386 704742 75622 704978
rect 75386 671658 75622 671894
rect 75386 634458 75622 634694
rect 75386 597258 75622 597494
rect 75386 560058 75622 560294
rect 75386 522858 75622 523094
rect 75386 485658 75622 485894
rect 75386 448458 75622 448694
rect 75386 411258 75622 411494
rect 75386 374058 75622 374294
rect 75386 336858 75622 337094
rect 75386 299658 75622 299894
rect 75386 262458 75622 262694
rect 75386 225258 75622 225494
rect 75386 188058 75622 188294
rect 75386 150858 75622 151094
rect 75386 113658 75622 113894
rect 75386 76458 75622 76694
rect 75386 39258 75622 39494
rect 75386 2058 75622 2294
rect 75386 -1042 75622 -806
rect 78986 705682 79222 705918
rect 78986 675258 79222 675494
rect 78986 638058 79222 638294
rect 78986 600858 79222 601094
rect 78986 563658 79222 563894
rect 78986 526458 79222 526694
rect 78986 489258 79222 489494
rect 78986 452058 79222 452294
rect 78986 414858 79222 415094
rect 78986 377658 79222 377894
rect 78986 340458 79222 340694
rect 78986 303258 79222 303494
rect 78986 266058 79222 266294
rect 78986 228858 79222 229094
rect 78986 191658 79222 191894
rect 78986 154458 79222 154694
rect 78986 117258 79222 117494
rect 78986 80058 79222 80294
rect 78986 42858 79222 43094
rect 78986 5658 79222 5894
rect 78986 -1982 79222 -1746
rect 112586 704742 112822 704978
rect 112586 671658 112822 671894
rect 112586 634458 112822 634694
rect 112586 597258 112822 597494
rect 112586 560058 112822 560294
rect 112586 522858 112822 523094
rect 112586 485658 112822 485894
rect 112586 448458 112822 448694
rect 112586 411258 112822 411494
rect 112586 374058 112822 374294
rect 112586 336858 112822 337094
rect 112586 299658 112822 299894
rect 112586 262458 112822 262694
rect 112586 225258 112822 225494
rect 112586 188058 112822 188294
rect 112586 150858 112822 151094
rect 112586 113658 112822 113894
rect 112586 76458 112822 76694
rect 112586 39258 112822 39494
rect 112586 2058 112822 2294
rect 112586 -1042 112822 -806
rect 116186 705682 116422 705918
rect 116186 675258 116422 675494
rect 116186 638058 116422 638294
rect 116186 600858 116422 601094
rect 116186 563658 116422 563894
rect 116186 526458 116422 526694
rect 116186 489258 116422 489494
rect 116186 452058 116422 452294
rect 116186 414858 116422 415094
rect 116186 377658 116422 377894
rect 116186 340458 116422 340694
rect 116186 303258 116422 303494
rect 116186 266058 116422 266294
rect 116186 228858 116422 229094
rect 116186 191658 116422 191894
rect 116186 154458 116422 154694
rect 116186 117258 116422 117494
rect 116186 80058 116422 80294
rect 116186 42858 116422 43094
rect 116186 5658 116422 5894
rect 116186 -1982 116422 -1746
rect 149786 704742 150022 704978
rect 149786 671658 150022 671894
rect 149786 634458 150022 634694
rect 149786 597258 150022 597494
rect 149786 560058 150022 560294
rect 149786 522858 150022 523094
rect 149786 485658 150022 485894
rect 149786 448458 150022 448694
rect 149786 411258 150022 411494
rect 149786 374058 150022 374294
rect 149786 336858 150022 337094
rect 149786 299658 150022 299894
rect 149786 262458 150022 262694
rect 149786 225258 150022 225494
rect 149786 188058 150022 188294
rect 149786 150858 150022 151094
rect 149786 113658 150022 113894
rect 149786 76458 150022 76694
rect 149786 39258 150022 39494
rect 149786 2058 150022 2294
rect 149786 -1042 150022 -806
rect 153386 705682 153622 705918
rect 153386 675258 153622 675494
rect 153386 638058 153622 638294
rect 153386 600858 153622 601094
rect 153386 563658 153622 563894
rect 153386 526458 153622 526694
rect 153386 489258 153622 489494
rect 153386 452058 153622 452294
rect 153386 414858 153622 415094
rect 153386 377658 153622 377894
rect 153386 340458 153622 340694
rect 153386 303258 153622 303494
rect 153386 266058 153622 266294
rect 153386 228858 153622 229094
rect 153386 191658 153622 191894
rect 153386 154458 153622 154694
rect 153386 117258 153622 117494
rect 153386 80058 153622 80294
rect 153386 42858 153622 43094
rect 153386 5658 153622 5894
rect 153386 -1982 153622 -1746
rect 186986 704742 187222 704978
rect 186986 671658 187222 671894
rect 186986 634458 187222 634694
rect 186986 597258 187222 597494
rect 186986 560058 187222 560294
rect 186986 522858 187222 523094
rect 186986 485658 187222 485894
rect 186986 448458 187222 448694
rect 186986 411258 187222 411494
rect 186986 374058 187222 374294
rect 186986 336858 187222 337094
rect 186986 299658 187222 299894
rect 186986 262458 187222 262694
rect 186986 225258 187222 225494
rect 186986 188058 187222 188294
rect 186986 150858 187222 151094
rect 186986 113658 187222 113894
rect 186986 76458 187222 76694
rect 186986 39258 187222 39494
rect 186986 2058 187222 2294
rect 186986 -1042 187222 -806
rect 190586 705682 190822 705918
rect 190586 675258 190822 675494
rect 190586 638058 190822 638294
rect 190586 600858 190822 601094
rect 190586 563658 190822 563894
rect 190586 526458 190822 526694
rect 190586 489258 190822 489494
rect 190586 452058 190822 452294
rect 190586 414858 190822 415094
rect 190586 377658 190822 377894
rect 190586 340458 190822 340694
rect 190586 303258 190822 303494
rect 190586 266058 190822 266294
rect 190586 228858 190822 229094
rect 190586 191658 190822 191894
rect 190586 154458 190822 154694
rect 190586 117258 190822 117494
rect 190586 80058 190822 80294
rect 190586 42858 190822 43094
rect 190586 5658 190822 5894
rect 190586 -1982 190822 -1746
rect 224186 704742 224422 704978
rect 224186 671658 224422 671894
rect 224186 634458 224422 634694
rect 224186 597258 224422 597494
rect 224186 560058 224422 560294
rect 224186 522858 224422 523094
rect 224186 485658 224422 485894
rect 224186 448458 224422 448694
rect 224186 411258 224422 411494
rect 224186 374058 224422 374294
rect 224186 336858 224422 337094
rect 224186 299658 224422 299894
rect 224186 262458 224422 262694
rect 224186 225258 224422 225494
rect 224186 188058 224422 188294
rect 224186 150858 224422 151094
rect 224186 113658 224422 113894
rect 224186 76458 224422 76694
rect 224186 39258 224422 39494
rect 224186 2058 224422 2294
rect 224186 -1042 224422 -806
rect 227786 705682 228022 705918
rect 227786 675258 228022 675494
rect 227786 638058 228022 638294
rect 227786 600858 228022 601094
rect 227786 563658 228022 563894
rect 227786 526458 228022 526694
rect 227786 489258 228022 489494
rect 227786 452058 228022 452294
rect 227786 414858 228022 415094
rect 227786 377658 228022 377894
rect 227786 340458 228022 340694
rect 227786 303258 228022 303494
rect 227786 266058 228022 266294
rect 227786 228858 228022 229094
rect 227786 191658 228022 191894
rect 227786 154458 228022 154694
rect 227786 117258 228022 117494
rect 227786 80058 228022 80294
rect 227786 42858 228022 43094
rect 227786 5658 228022 5894
rect 227786 -1982 228022 -1746
rect 261386 704742 261622 704978
rect 261386 671658 261622 671894
rect 261386 634458 261622 634694
rect 261386 597258 261622 597494
rect 261386 560058 261622 560294
rect 261386 522858 261622 523094
rect 261386 485658 261622 485894
rect 261386 448458 261622 448694
rect 261386 411258 261622 411494
rect 261386 374058 261622 374294
rect 261386 336858 261622 337094
rect 261386 299658 261622 299894
rect 261386 262458 261622 262694
rect 261386 225258 261622 225494
rect 261386 188058 261622 188294
rect 261386 150858 261622 151094
rect 261386 113658 261622 113894
rect 261386 76458 261622 76694
rect 261386 39258 261622 39494
rect 261386 2058 261622 2294
rect 261386 -1042 261622 -806
rect 264986 705682 265222 705918
rect 264986 675258 265222 675494
rect 264986 638058 265222 638294
rect 264986 600858 265222 601094
rect 264986 563658 265222 563894
rect 264986 526458 265222 526694
rect 264986 489258 265222 489494
rect 264986 452058 265222 452294
rect 264986 414858 265222 415094
rect 264986 377658 265222 377894
rect 298586 704742 298822 704978
rect 298586 671658 298822 671894
rect 298586 634458 298822 634694
rect 298586 597258 298822 597494
rect 298586 560058 298822 560294
rect 298586 522858 298822 523094
rect 298586 485658 298822 485894
rect 298586 448458 298822 448694
rect 298586 411258 298822 411494
rect 298586 374058 298822 374294
rect 264986 340458 265222 340694
rect 264986 303258 265222 303494
rect 264986 266058 265222 266294
rect 264986 228858 265222 229094
rect 264986 191658 265222 191894
rect 264986 154458 265222 154694
rect 264986 117258 265222 117494
rect 264986 80058 265222 80294
rect 264986 42858 265222 43094
rect 302186 705682 302422 705918
rect 302186 675258 302422 675494
rect 302186 638058 302422 638294
rect 302186 600858 302422 601094
rect 302186 563658 302422 563894
rect 302186 526458 302422 526694
rect 302186 489258 302422 489494
rect 302186 452058 302422 452294
rect 302186 414858 302422 415094
rect 302186 377658 302422 377894
rect 298586 336858 298822 337094
rect 298586 299658 298822 299894
rect 298586 262458 298822 262694
rect 298586 225258 298822 225494
rect 298586 188058 298822 188294
rect 298586 150858 298822 151094
rect 298586 113658 298822 113894
rect 335786 704742 336022 704978
rect 335786 671658 336022 671894
rect 335786 634458 336022 634694
rect 335786 597258 336022 597494
rect 335786 560058 336022 560294
rect 335786 522858 336022 523094
rect 335786 485658 336022 485894
rect 335786 448458 336022 448694
rect 335786 411258 336022 411494
rect 335786 374058 336022 374294
rect 302186 340458 302422 340694
rect 302186 303258 302422 303494
rect 302186 266058 302422 266294
rect 302186 228858 302422 229094
rect 302186 191658 302422 191894
rect 302186 154458 302422 154694
rect 335786 336858 336022 337094
rect 335786 299658 336022 299894
rect 335786 262458 336022 262694
rect 335786 225258 336022 225494
rect 335786 188058 336022 188294
rect 335786 150858 336022 151094
rect 302186 117258 302422 117494
rect 298586 76458 298822 76694
rect 298586 39258 298822 39494
rect 264986 5658 265222 5894
rect 264986 -1982 265222 -1746
rect 298586 2058 298822 2294
rect 298586 -1042 298822 -806
rect 302186 80058 302422 80294
rect 302186 42858 302422 43094
rect 302186 5658 302422 5894
rect 302186 -1982 302422 -1746
rect 335786 113658 336022 113894
rect 335786 76458 336022 76694
rect 335786 39258 336022 39494
rect 335786 2058 336022 2294
rect 335786 -1042 336022 -806
rect 339386 705682 339622 705918
rect 339386 675258 339622 675494
rect 339386 638058 339622 638294
rect 339386 600858 339622 601094
rect 339386 563658 339622 563894
rect 339386 526458 339622 526694
rect 339386 489258 339622 489494
rect 339386 452058 339622 452294
rect 339386 414858 339622 415094
rect 339386 377658 339622 377894
rect 339386 340458 339622 340694
rect 339386 303258 339622 303494
rect 339386 266058 339622 266294
rect 339386 228858 339622 229094
rect 339386 191658 339622 191894
rect 339386 154458 339622 154694
rect 339386 117258 339622 117494
rect 339386 80058 339622 80294
rect 339386 42858 339622 43094
rect 339386 5658 339622 5894
rect 339386 -1982 339622 -1746
rect 372986 704742 373222 704978
rect 372986 671658 373222 671894
rect 372986 634458 373222 634694
rect 372986 597258 373222 597494
rect 372986 560058 373222 560294
rect 372986 522858 373222 523094
rect 372986 485658 373222 485894
rect 372986 448458 373222 448694
rect 372986 411258 373222 411494
rect 372986 374058 373222 374294
rect 372986 336858 373222 337094
rect 372986 299658 373222 299894
rect 372986 262458 373222 262694
rect 372986 225258 373222 225494
rect 372986 188058 373222 188294
rect 372986 150858 373222 151094
rect 372986 113658 373222 113894
rect 372986 76458 373222 76694
rect 372986 39258 373222 39494
rect 372986 2058 373222 2294
rect 372986 -1042 373222 -806
rect 376586 705682 376822 705918
rect 376586 675258 376822 675494
rect 376586 638058 376822 638294
rect 376586 600858 376822 601094
rect 376586 563658 376822 563894
rect 376586 526458 376822 526694
rect 376586 489258 376822 489494
rect 376586 452058 376822 452294
rect 376586 414858 376822 415094
rect 376586 377658 376822 377894
rect 376586 340458 376822 340694
rect 376586 303258 376822 303494
rect 376586 266058 376822 266294
rect 376586 228858 376822 229094
rect 376586 191658 376822 191894
rect 376586 154458 376822 154694
rect 376586 117258 376822 117494
rect 376586 80058 376822 80294
rect 376586 42858 376822 43094
rect 376586 5658 376822 5894
rect 376586 -1982 376822 -1746
rect 410186 704742 410422 704978
rect 410186 671658 410422 671894
rect 410186 634458 410422 634694
rect 410186 597258 410422 597494
rect 410186 560058 410422 560294
rect 410186 522858 410422 523094
rect 410186 485658 410422 485894
rect 410186 448458 410422 448694
rect 410186 411258 410422 411494
rect 410186 374058 410422 374294
rect 410186 336858 410422 337094
rect 410186 299658 410422 299894
rect 410186 262458 410422 262694
rect 410186 225258 410422 225494
rect 410186 188058 410422 188294
rect 410186 150858 410422 151094
rect 410186 113658 410422 113894
rect 410186 76458 410422 76694
rect 410186 39258 410422 39494
rect 410186 2058 410422 2294
rect 410186 -1042 410422 -806
rect 413786 705682 414022 705918
rect 413786 675258 414022 675494
rect 413786 638058 414022 638294
rect 413786 600858 414022 601094
rect 413786 563658 414022 563894
rect 413786 526458 414022 526694
rect 413786 489258 414022 489494
rect 413786 452058 414022 452294
rect 413786 414858 414022 415094
rect 413786 377658 414022 377894
rect 413786 340458 414022 340694
rect 413786 303258 414022 303494
rect 413786 266058 414022 266294
rect 413786 228858 414022 229094
rect 413786 191658 414022 191894
rect 413786 154458 414022 154694
rect 413786 117258 414022 117494
rect 413786 80058 414022 80294
rect 413786 42858 414022 43094
rect 413786 5658 414022 5894
rect 413786 -1982 414022 -1746
rect 447386 704742 447622 704978
rect 447386 671658 447622 671894
rect 447386 634458 447622 634694
rect 447386 597258 447622 597494
rect 447386 560058 447622 560294
rect 447386 522858 447622 523094
rect 447386 485658 447622 485894
rect 447386 448458 447622 448694
rect 447386 411258 447622 411494
rect 447386 374058 447622 374294
rect 447386 336858 447622 337094
rect 447386 299658 447622 299894
rect 447386 262458 447622 262694
rect 447386 225258 447622 225494
rect 447386 188058 447622 188294
rect 447386 150858 447622 151094
rect 447386 113658 447622 113894
rect 447386 76458 447622 76694
rect 447386 39258 447622 39494
rect 447386 2058 447622 2294
rect 447386 -1042 447622 -806
rect 450986 705682 451222 705918
rect 450986 675258 451222 675494
rect 450986 638058 451222 638294
rect 450986 600858 451222 601094
rect 450986 563658 451222 563894
rect 450986 526458 451222 526694
rect 450986 489258 451222 489494
rect 450986 452058 451222 452294
rect 450986 414858 451222 415094
rect 450986 377658 451222 377894
rect 450986 340458 451222 340694
rect 450986 303258 451222 303494
rect 450986 266058 451222 266294
rect 450986 228858 451222 229094
rect 450986 191658 451222 191894
rect 450986 154458 451222 154694
rect 450986 117258 451222 117494
rect 450986 80058 451222 80294
rect 450986 42858 451222 43094
rect 450986 5658 451222 5894
rect 450986 -1982 451222 -1746
rect 484586 704742 484822 704978
rect 484586 671658 484822 671894
rect 484586 634458 484822 634694
rect 484586 597258 484822 597494
rect 484586 560058 484822 560294
rect 484586 522858 484822 523094
rect 484586 485658 484822 485894
rect 484586 448458 484822 448694
rect 484586 411258 484822 411494
rect 484586 374058 484822 374294
rect 484586 336858 484822 337094
rect 484586 299658 484822 299894
rect 484586 262458 484822 262694
rect 484586 225258 484822 225494
rect 484586 188058 484822 188294
rect 484586 150858 484822 151094
rect 484586 113658 484822 113894
rect 484586 76458 484822 76694
rect 484586 39258 484822 39494
rect 484586 2058 484822 2294
rect 484586 -1042 484822 -806
rect 488186 705682 488422 705918
rect 488186 675258 488422 675494
rect 488186 638058 488422 638294
rect 488186 600858 488422 601094
rect 488186 563658 488422 563894
rect 488186 526458 488422 526694
rect 488186 489258 488422 489494
rect 488186 452058 488422 452294
rect 488186 414858 488422 415094
rect 488186 377658 488422 377894
rect 521786 704742 522022 704978
rect 521786 671658 522022 671894
rect 521786 634458 522022 634694
rect 521786 597258 522022 597494
rect 521786 560058 522022 560294
rect 521786 522858 522022 523094
rect 521786 485658 522022 485894
rect 521786 448458 522022 448694
rect 521786 411258 522022 411494
rect 521786 374058 522022 374294
rect 525386 705682 525622 705918
rect 525386 675258 525622 675494
rect 525386 638058 525622 638294
rect 525386 600858 525622 601094
rect 525386 563658 525622 563894
rect 525386 526458 525622 526694
rect 525386 489258 525622 489494
rect 525386 452058 525622 452294
rect 525386 414858 525622 415094
rect 525386 377658 525622 377894
rect 558986 704742 559222 704978
rect 558986 671658 559222 671894
rect 558986 634458 559222 634694
rect 558986 597258 559222 597494
rect 558986 560058 559222 560294
rect 558986 522858 559222 523094
rect 558986 485658 559222 485894
rect 558986 448458 559222 448694
rect 558986 411258 559222 411494
rect 558986 374058 559222 374294
rect 488186 340458 488422 340694
rect 521952 336858 522188 337094
rect 523884 336858 524120 337094
rect 525816 336858 526052 337094
rect 527748 336858 527984 337094
rect 558986 336858 559222 337094
rect 488186 303258 488422 303494
rect 488186 266058 488422 266294
rect 488186 228858 488422 229094
rect 488186 191658 488422 191894
rect 488186 154458 488422 154694
rect 488186 117258 488422 117494
rect 488186 80058 488422 80294
rect 488186 42858 488422 43094
rect 488186 5658 488422 5894
rect 488186 -1982 488422 -1746
rect 521786 299658 522022 299894
rect 521786 262458 522022 262694
rect 521786 225258 522022 225494
rect 521786 188058 522022 188294
rect 521786 150858 522022 151094
rect 521786 113658 522022 113894
rect 521786 76458 522022 76694
rect 521786 39258 522022 39494
rect 521786 2058 522022 2294
rect 521786 -1042 522022 -806
rect 525386 303258 525622 303494
rect 525386 266058 525622 266294
rect 525386 228858 525622 229094
rect 525386 191658 525622 191894
rect 525386 154458 525622 154694
rect 525386 117258 525622 117494
rect 525386 80058 525622 80294
rect 525386 42858 525622 43094
rect 558986 299658 559222 299894
rect 558986 262458 559222 262694
rect 558986 225258 559222 225494
rect 558986 188058 559222 188294
rect 558986 150858 559222 151094
rect 558986 113658 559222 113894
rect 558986 76458 559222 76694
rect 558986 39258 559222 39494
rect 525386 5658 525622 5894
rect 525386 -1982 525622 -1746
rect 558986 2058 559222 2294
rect 558986 -1042 559222 -806
rect 562586 705682 562822 705918
rect 586742 705682 586978 705918
rect 562586 675258 562822 675494
rect 562586 638058 562822 638294
rect 562586 600858 562822 601094
rect 562586 563658 562822 563894
rect 562586 526458 562822 526694
rect 562586 489258 562822 489494
rect 562586 452058 562822 452294
rect 562586 414858 562822 415094
rect 562586 377658 562822 377894
rect 562586 340458 562822 340694
rect 562586 303258 562822 303494
rect 562586 266058 562822 266294
rect 562586 228858 562822 229094
rect 562586 191658 562822 191894
rect 562586 154458 562822 154694
rect 562586 117258 562822 117494
rect 562586 80058 562822 80294
rect 562586 42858 562822 43094
rect 562586 5658 562822 5894
rect 585802 704742 586038 704978
rect 585802 671658 586038 671894
rect 585802 634458 586038 634694
rect 585802 597258 586038 597494
rect 585802 560058 586038 560294
rect 585802 522858 586038 523094
rect 585802 485658 586038 485894
rect 585802 448458 586038 448694
rect 585802 411258 586038 411494
rect 585802 374058 586038 374294
rect 585802 336858 586038 337094
rect 585802 299658 586038 299894
rect 585802 262458 586038 262694
rect 585802 225258 586038 225494
rect 585802 188058 586038 188294
rect 585802 150858 586038 151094
rect 585802 113658 586038 113894
rect 585802 76458 586038 76694
rect 585802 39258 586038 39494
rect 585802 2058 586038 2294
rect 585802 -1042 586038 -806
rect 586742 675258 586978 675494
rect 586742 638058 586978 638294
rect 586742 600858 586978 601094
rect 586742 563658 586978 563894
rect 586742 526458 586978 526694
rect 586742 489258 586978 489494
rect 586742 452058 586978 452294
rect 586742 414858 586978 415094
rect 586742 377658 586978 377894
rect 586742 340458 586978 340694
rect 586742 303258 586978 303494
rect 586742 266058 586978 266294
rect 586742 228858 586978 229094
rect 586742 191658 586978 191894
rect 586742 154458 586978 154694
rect 586742 117258 586978 117494
rect 586742 80058 586978 80294
rect 586742 42858 586978 43094
rect 586742 5658 586978 5894
rect 562586 -1982 562822 -1746
rect 586742 -1982 586978 -1746
<< metal5 >>
rect -3236 705918 587160 706100
rect -3236 705682 -3054 705918
rect -2818 705682 4586 705918
rect 4822 705682 41786 705918
rect 42022 705682 78986 705918
rect 79222 705682 116186 705918
rect 116422 705682 153386 705918
rect 153622 705682 190586 705918
rect 190822 705682 227786 705918
rect 228022 705682 264986 705918
rect 265222 705682 302186 705918
rect 302422 705682 339386 705918
rect 339622 705682 376586 705918
rect 376822 705682 413786 705918
rect 414022 705682 450986 705918
rect 451222 705682 488186 705918
rect 488422 705682 525386 705918
rect 525622 705682 562586 705918
rect 562822 705682 586742 705918
rect 586978 705682 587160 705918
rect -3236 705500 587160 705682
rect -2296 704978 586220 705160
rect -2296 704742 -2114 704978
rect -1878 704742 986 704978
rect 1222 704742 38186 704978
rect 38422 704742 75386 704978
rect 75622 704742 112586 704978
rect 112822 704742 149786 704978
rect 150022 704742 186986 704978
rect 187222 704742 224186 704978
rect 224422 704742 261386 704978
rect 261622 704742 298586 704978
rect 298822 704742 335786 704978
rect 336022 704742 372986 704978
rect 373222 704742 410186 704978
rect 410422 704742 447386 704978
rect 447622 704742 484586 704978
rect 484822 704742 521786 704978
rect 522022 704742 558986 704978
rect 559222 704742 585802 704978
rect 586038 704742 586220 704978
rect -2296 704560 586220 704742
rect -3236 675494 587160 675676
rect -3236 675258 -3054 675494
rect -2818 675258 4586 675494
rect 4822 675258 41786 675494
rect 42022 675258 78986 675494
rect 79222 675258 116186 675494
rect 116422 675258 153386 675494
rect 153622 675258 190586 675494
rect 190822 675258 227786 675494
rect 228022 675258 264986 675494
rect 265222 675258 302186 675494
rect 302422 675258 339386 675494
rect 339622 675258 376586 675494
rect 376822 675258 413786 675494
rect 414022 675258 450986 675494
rect 451222 675258 488186 675494
rect 488422 675258 525386 675494
rect 525622 675258 562586 675494
rect 562822 675258 586742 675494
rect 586978 675258 587160 675494
rect -3236 675076 587160 675258
rect -3236 671894 587160 672076
rect -3236 671658 -2114 671894
rect -1878 671658 986 671894
rect 1222 671658 38186 671894
rect 38422 671658 75386 671894
rect 75622 671658 112586 671894
rect 112822 671658 149786 671894
rect 150022 671658 186986 671894
rect 187222 671658 224186 671894
rect 224422 671658 261386 671894
rect 261622 671658 298586 671894
rect 298822 671658 335786 671894
rect 336022 671658 372986 671894
rect 373222 671658 410186 671894
rect 410422 671658 447386 671894
rect 447622 671658 484586 671894
rect 484822 671658 521786 671894
rect 522022 671658 558986 671894
rect 559222 671658 585802 671894
rect 586038 671658 587160 671894
rect -3236 671476 587160 671658
rect -3236 638294 587160 638476
rect -3236 638058 -3054 638294
rect -2818 638058 4586 638294
rect 4822 638058 41786 638294
rect 42022 638058 78986 638294
rect 79222 638058 116186 638294
rect 116422 638058 153386 638294
rect 153622 638058 190586 638294
rect 190822 638058 227786 638294
rect 228022 638058 264986 638294
rect 265222 638058 302186 638294
rect 302422 638058 339386 638294
rect 339622 638058 376586 638294
rect 376822 638058 413786 638294
rect 414022 638058 450986 638294
rect 451222 638058 488186 638294
rect 488422 638058 525386 638294
rect 525622 638058 562586 638294
rect 562822 638058 586742 638294
rect 586978 638058 587160 638294
rect -3236 637876 587160 638058
rect -3236 634694 587160 634876
rect -3236 634458 -2114 634694
rect -1878 634458 986 634694
rect 1222 634458 38186 634694
rect 38422 634458 75386 634694
rect 75622 634458 112586 634694
rect 112822 634458 149786 634694
rect 150022 634458 186986 634694
rect 187222 634458 224186 634694
rect 224422 634458 261386 634694
rect 261622 634458 298586 634694
rect 298822 634458 335786 634694
rect 336022 634458 372986 634694
rect 373222 634458 410186 634694
rect 410422 634458 447386 634694
rect 447622 634458 484586 634694
rect 484822 634458 521786 634694
rect 522022 634458 558986 634694
rect 559222 634458 585802 634694
rect 586038 634458 587160 634694
rect -3236 634276 587160 634458
rect -3236 601094 587160 601276
rect -3236 600858 -3054 601094
rect -2818 600858 4586 601094
rect 4822 600858 41786 601094
rect 42022 600858 78986 601094
rect 79222 600858 116186 601094
rect 116422 600858 153386 601094
rect 153622 600858 190586 601094
rect 190822 600858 227786 601094
rect 228022 600858 264986 601094
rect 265222 600858 302186 601094
rect 302422 600858 339386 601094
rect 339622 600858 376586 601094
rect 376822 600858 413786 601094
rect 414022 600858 450986 601094
rect 451222 600858 488186 601094
rect 488422 600858 525386 601094
rect 525622 600858 562586 601094
rect 562822 600858 586742 601094
rect 586978 600858 587160 601094
rect -3236 600676 587160 600858
rect -3236 597494 587160 597676
rect -3236 597258 -2114 597494
rect -1878 597258 986 597494
rect 1222 597258 38186 597494
rect 38422 597258 75386 597494
rect 75622 597258 112586 597494
rect 112822 597258 149786 597494
rect 150022 597258 186986 597494
rect 187222 597258 224186 597494
rect 224422 597258 261386 597494
rect 261622 597258 298586 597494
rect 298822 597258 335786 597494
rect 336022 597258 372986 597494
rect 373222 597258 410186 597494
rect 410422 597258 447386 597494
rect 447622 597258 484586 597494
rect 484822 597258 521786 597494
rect 522022 597258 558986 597494
rect 559222 597258 585802 597494
rect 586038 597258 587160 597494
rect -3236 597076 587160 597258
rect -3236 563894 587160 564076
rect -3236 563658 -3054 563894
rect -2818 563658 4586 563894
rect 4822 563658 41786 563894
rect 42022 563658 78986 563894
rect 79222 563658 116186 563894
rect 116422 563658 153386 563894
rect 153622 563658 190586 563894
rect 190822 563658 227786 563894
rect 228022 563658 264986 563894
rect 265222 563658 302186 563894
rect 302422 563658 339386 563894
rect 339622 563658 376586 563894
rect 376822 563658 413786 563894
rect 414022 563658 450986 563894
rect 451222 563658 488186 563894
rect 488422 563658 525386 563894
rect 525622 563658 562586 563894
rect 562822 563658 586742 563894
rect 586978 563658 587160 563894
rect -3236 563476 587160 563658
rect -3236 560294 587160 560476
rect -3236 560058 -2114 560294
rect -1878 560058 986 560294
rect 1222 560058 38186 560294
rect 38422 560058 75386 560294
rect 75622 560058 112586 560294
rect 112822 560058 149786 560294
rect 150022 560058 186986 560294
rect 187222 560058 224186 560294
rect 224422 560058 261386 560294
rect 261622 560058 298586 560294
rect 298822 560058 335786 560294
rect 336022 560058 372986 560294
rect 373222 560058 410186 560294
rect 410422 560058 447386 560294
rect 447622 560058 484586 560294
rect 484822 560058 521786 560294
rect 522022 560058 558986 560294
rect 559222 560058 585802 560294
rect 586038 560058 587160 560294
rect -3236 559876 587160 560058
rect -3236 526694 587160 526876
rect -3236 526458 -3054 526694
rect -2818 526458 4586 526694
rect 4822 526458 41786 526694
rect 42022 526458 78986 526694
rect 79222 526458 116186 526694
rect 116422 526458 153386 526694
rect 153622 526458 190586 526694
rect 190822 526458 227786 526694
rect 228022 526458 264986 526694
rect 265222 526458 302186 526694
rect 302422 526458 339386 526694
rect 339622 526458 376586 526694
rect 376822 526458 413786 526694
rect 414022 526458 450986 526694
rect 451222 526458 488186 526694
rect 488422 526458 525386 526694
rect 525622 526458 562586 526694
rect 562822 526458 586742 526694
rect 586978 526458 587160 526694
rect -3236 526276 587160 526458
rect -3236 523094 587160 523276
rect -3236 522858 -2114 523094
rect -1878 522858 986 523094
rect 1222 522858 38186 523094
rect 38422 522858 75386 523094
rect 75622 522858 112586 523094
rect 112822 522858 149786 523094
rect 150022 522858 186986 523094
rect 187222 522858 224186 523094
rect 224422 522858 261386 523094
rect 261622 522858 298586 523094
rect 298822 522858 335786 523094
rect 336022 522858 372986 523094
rect 373222 522858 410186 523094
rect 410422 522858 447386 523094
rect 447622 522858 484586 523094
rect 484822 522858 521786 523094
rect 522022 522858 558986 523094
rect 559222 522858 585802 523094
rect 586038 522858 587160 523094
rect -3236 522676 587160 522858
rect -3236 489494 587160 489676
rect -3236 489258 -3054 489494
rect -2818 489258 4586 489494
rect 4822 489258 41786 489494
rect 42022 489258 78986 489494
rect 79222 489258 116186 489494
rect 116422 489258 153386 489494
rect 153622 489258 190586 489494
rect 190822 489258 227786 489494
rect 228022 489258 264986 489494
rect 265222 489258 302186 489494
rect 302422 489258 339386 489494
rect 339622 489258 376586 489494
rect 376822 489258 413786 489494
rect 414022 489258 450986 489494
rect 451222 489258 488186 489494
rect 488422 489258 525386 489494
rect 525622 489258 562586 489494
rect 562822 489258 586742 489494
rect 586978 489258 587160 489494
rect -3236 489076 587160 489258
rect -3236 485894 587160 486076
rect -3236 485658 -2114 485894
rect -1878 485658 986 485894
rect 1222 485658 38186 485894
rect 38422 485658 75386 485894
rect 75622 485658 112586 485894
rect 112822 485658 149786 485894
rect 150022 485658 186986 485894
rect 187222 485658 224186 485894
rect 224422 485658 261386 485894
rect 261622 485658 298586 485894
rect 298822 485658 335786 485894
rect 336022 485658 372986 485894
rect 373222 485658 410186 485894
rect 410422 485658 447386 485894
rect 447622 485658 484586 485894
rect 484822 485658 521786 485894
rect 522022 485658 558986 485894
rect 559222 485658 585802 485894
rect 586038 485658 587160 485894
rect -3236 485476 587160 485658
rect -3236 452294 587160 452476
rect -3236 452058 -3054 452294
rect -2818 452058 4586 452294
rect 4822 452058 41786 452294
rect 42022 452058 78986 452294
rect 79222 452058 116186 452294
rect 116422 452058 153386 452294
rect 153622 452058 190586 452294
rect 190822 452058 227786 452294
rect 228022 452058 264986 452294
rect 265222 452058 302186 452294
rect 302422 452058 339386 452294
rect 339622 452058 376586 452294
rect 376822 452058 413786 452294
rect 414022 452058 450986 452294
rect 451222 452058 488186 452294
rect 488422 452058 525386 452294
rect 525622 452058 562586 452294
rect 562822 452058 586742 452294
rect 586978 452058 587160 452294
rect -3236 451876 587160 452058
rect -3236 448694 587160 448876
rect -3236 448458 -2114 448694
rect -1878 448458 986 448694
rect 1222 448458 38186 448694
rect 38422 448458 75386 448694
rect 75622 448458 112586 448694
rect 112822 448458 149786 448694
rect 150022 448458 186986 448694
rect 187222 448458 224186 448694
rect 224422 448458 261386 448694
rect 261622 448458 298586 448694
rect 298822 448458 335786 448694
rect 336022 448458 372986 448694
rect 373222 448458 410186 448694
rect 410422 448458 447386 448694
rect 447622 448458 484586 448694
rect 484822 448458 521786 448694
rect 522022 448458 558986 448694
rect 559222 448458 585802 448694
rect 586038 448458 587160 448694
rect -3236 448276 587160 448458
rect -3236 415094 587160 415276
rect -3236 414858 -3054 415094
rect -2818 414858 4586 415094
rect 4822 414858 41786 415094
rect 42022 414858 78986 415094
rect 79222 414858 116186 415094
rect 116422 414858 153386 415094
rect 153622 414858 190586 415094
rect 190822 414858 227786 415094
rect 228022 414858 264986 415094
rect 265222 414858 302186 415094
rect 302422 414858 339386 415094
rect 339622 414858 376586 415094
rect 376822 414858 413786 415094
rect 414022 414858 450986 415094
rect 451222 414858 488186 415094
rect 488422 414858 525386 415094
rect 525622 414858 562586 415094
rect 562822 414858 586742 415094
rect 586978 414858 587160 415094
rect -3236 414676 587160 414858
rect -3236 411494 587160 411676
rect -3236 411258 -2114 411494
rect -1878 411258 986 411494
rect 1222 411258 38186 411494
rect 38422 411258 75386 411494
rect 75622 411258 112586 411494
rect 112822 411258 149786 411494
rect 150022 411258 186986 411494
rect 187222 411258 224186 411494
rect 224422 411258 261386 411494
rect 261622 411258 298586 411494
rect 298822 411258 335786 411494
rect 336022 411258 372986 411494
rect 373222 411258 410186 411494
rect 410422 411258 447386 411494
rect 447622 411258 484586 411494
rect 484822 411258 521786 411494
rect 522022 411258 558986 411494
rect 559222 411258 585802 411494
rect 586038 411258 587160 411494
rect -3236 411076 587160 411258
rect -3236 377894 587160 378076
rect -3236 377658 -3054 377894
rect -2818 377658 4586 377894
rect 4822 377658 41786 377894
rect 42022 377658 78986 377894
rect 79222 377658 116186 377894
rect 116422 377658 153386 377894
rect 153622 377658 190586 377894
rect 190822 377658 227786 377894
rect 228022 377658 264986 377894
rect 265222 377658 302186 377894
rect 302422 377658 339386 377894
rect 339622 377658 376586 377894
rect 376822 377658 413786 377894
rect 414022 377658 450986 377894
rect 451222 377658 488186 377894
rect 488422 377658 525386 377894
rect 525622 377658 562586 377894
rect 562822 377658 586742 377894
rect 586978 377658 587160 377894
rect -3236 377476 587160 377658
rect -3236 374294 587160 374476
rect -3236 374058 -2114 374294
rect -1878 374058 986 374294
rect 1222 374058 38186 374294
rect 38422 374058 75386 374294
rect 75622 374058 112586 374294
rect 112822 374058 149786 374294
rect 150022 374058 186986 374294
rect 187222 374058 224186 374294
rect 224422 374058 261386 374294
rect 261622 374058 298586 374294
rect 298822 374058 335786 374294
rect 336022 374058 372986 374294
rect 373222 374058 410186 374294
rect 410422 374058 447386 374294
rect 447622 374058 484586 374294
rect 484822 374058 521786 374294
rect 522022 374058 558986 374294
rect 559222 374058 585802 374294
rect 586038 374058 587160 374294
rect -3236 373876 587160 374058
rect -3236 340694 587160 340876
rect -3236 340458 -3054 340694
rect -2818 340458 4586 340694
rect 4822 340458 41786 340694
rect 42022 340458 78986 340694
rect 79222 340458 116186 340694
rect 116422 340458 153386 340694
rect 153622 340458 190586 340694
rect 190822 340458 227786 340694
rect 228022 340458 264986 340694
rect 265222 340458 302186 340694
rect 302422 340458 339386 340694
rect 339622 340458 376586 340694
rect 376822 340458 413786 340694
rect 414022 340458 450986 340694
rect 451222 340458 488186 340694
rect 488422 340458 562586 340694
rect 562822 340458 586742 340694
rect 586978 340458 587160 340694
rect -3236 340276 587160 340458
rect -3236 337094 587160 337276
rect -3236 336858 -2114 337094
rect -1878 336858 986 337094
rect 1222 336858 38186 337094
rect 38422 336858 75386 337094
rect 75622 336858 112586 337094
rect 112822 336858 149786 337094
rect 150022 336858 186986 337094
rect 187222 336858 224186 337094
rect 224422 336858 261386 337094
rect 261622 336858 298586 337094
rect 298822 336858 335786 337094
rect 336022 336858 372986 337094
rect 373222 336858 410186 337094
rect 410422 336858 447386 337094
rect 447622 336858 484586 337094
rect 484822 336858 521952 337094
rect 522188 336858 523884 337094
rect 524120 336858 525816 337094
rect 526052 336858 527748 337094
rect 527984 336858 558986 337094
rect 559222 336858 585802 337094
rect 586038 336858 587160 337094
rect -3236 336676 587160 336858
rect -3236 303494 587160 303676
rect -3236 303258 -3054 303494
rect -2818 303258 4586 303494
rect 4822 303258 41786 303494
rect 42022 303258 78986 303494
rect 79222 303258 116186 303494
rect 116422 303258 153386 303494
rect 153622 303258 190586 303494
rect 190822 303258 227786 303494
rect 228022 303258 264986 303494
rect 265222 303258 302186 303494
rect 302422 303258 339386 303494
rect 339622 303258 376586 303494
rect 376822 303258 413786 303494
rect 414022 303258 450986 303494
rect 451222 303258 488186 303494
rect 488422 303258 525386 303494
rect 525622 303258 562586 303494
rect 562822 303258 586742 303494
rect 586978 303258 587160 303494
rect -3236 303076 587160 303258
rect -3236 299894 587160 300076
rect -3236 299658 -2114 299894
rect -1878 299658 986 299894
rect 1222 299658 38186 299894
rect 38422 299658 75386 299894
rect 75622 299658 112586 299894
rect 112822 299658 149786 299894
rect 150022 299658 186986 299894
rect 187222 299658 224186 299894
rect 224422 299658 261386 299894
rect 261622 299658 298586 299894
rect 298822 299658 335786 299894
rect 336022 299658 372986 299894
rect 373222 299658 410186 299894
rect 410422 299658 447386 299894
rect 447622 299658 484586 299894
rect 484822 299658 521786 299894
rect 522022 299658 558986 299894
rect 559222 299658 585802 299894
rect 586038 299658 587160 299894
rect -3236 299476 587160 299658
rect -3236 266294 587160 266476
rect -3236 266058 -3054 266294
rect -2818 266058 4586 266294
rect 4822 266058 41786 266294
rect 42022 266058 78986 266294
rect 79222 266058 116186 266294
rect 116422 266058 153386 266294
rect 153622 266058 190586 266294
rect 190822 266058 227786 266294
rect 228022 266058 264986 266294
rect 265222 266058 302186 266294
rect 302422 266058 339386 266294
rect 339622 266058 376586 266294
rect 376822 266058 413786 266294
rect 414022 266058 450986 266294
rect 451222 266058 488186 266294
rect 488422 266058 525386 266294
rect 525622 266058 562586 266294
rect 562822 266058 586742 266294
rect 586978 266058 587160 266294
rect -3236 265876 587160 266058
rect -3236 262694 587160 262876
rect -3236 262458 -2114 262694
rect -1878 262458 986 262694
rect 1222 262458 38186 262694
rect 38422 262458 75386 262694
rect 75622 262458 112586 262694
rect 112822 262458 149786 262694
rect 150022 262458 186986 262694
rect 187222 262458 224186 262694
rect 224422 262458 261386 262694
rect 261622 262458 298586 262694
rect 298822 262458 335786 262694
rect 336022 262458 372986 262694
rect 373222 262458 410186 262694
rect 410422 262458 447386 262694
rect 447622 262458 484586 262694
rect 484822 262458 521786 262694
rect 522022 262458 558986 262694
rect 559222 262458 585802 262694
rect 586038 262458 587160 262694
rect -3236 262276 587160 262458
rect -3236 229094 587160 229276
rect -3236 228858 -3054 229094
rect -2818 228858 4586 229094
rect 4822 228858 41786 229094
rect 42022 228858 78986 229094
rect 79222 228858 116186 229094
rect 116422 228858 153386 229094
rect 153622 228858 190586 229094
rect 190822 228858 227786 229094
rect 228022 228858 264986 229094
rect 265222 228858 302186 229094
rect 302422 228858 339386 229094
rect 339622 228858 376586 229094
rect 376822 228858 413786 229094
rect 414022 228858 450986 229094
rect 451222 228858 488186 229094
rect 488422 228858 525386 229094
rect 525622 228858 562586 229094
rect 562822 228858 586742 229094
rect 586978 228858 587160 229094
rect -3236 228676 587160 228858
rect -3236 225494 587160 225676
rect -3236 225258 -2114 225494
rect -1878 225258 986 225494
rect 1222 225258 38186 225494
rect 38422 225258 75386 225494
rect 75622 225258 112586 225494
rect 112822 225258 149786 225494
rect 150022 225258 186986 225494
rect 187222 225258 224186 225494
rect 224422 225258 261386 225494
rect 261622 225258 298586 225494
rect 298822 225258 335786 225494
rect 336022 225258 372986 225494
rect 373222 225258 410186 225494
rect 410422 225258 447386 225494
rect 447622 225258 484586 225494
rect 484822 225258 521786 225494
rect 522022 225258 558986 225494
rect 559222 225258 585802 225494
rect 586038 225258 587160 225494
rect -3236 225076 587160 225258
rect -3236 191894 587160 192076
rect -3236 191658 -3054 191894
rect -2818 191658 4586 191894
rect 4822 191658 41786 191894
rect 42022 191658 78986 191894
rect 79222 191658 116186 191894
rect 116422 191658 153386 191894
rect 153622 191658 190586 191894
rect 190822 191658 227786 191894
rect 228022 191658 264986 191894
rect 265222 191658 302186 191894
rect 302422 191658 339386 191894
rect 339622 191658 376586 191894
rect 376822 191658 413786 191894
rect 414022 191658 450986 191894
rect 451222 191658 488186 191894
rect 488422 191658 525386 191894
rect 525622 191658 562586 191894
rect 562822 191658 586742 191894
rect 586978 191658 587160 191894
rect -3236 191476 587160 191658
rect -3236 188294 587160 188476
rect -3236 188058 -2114 188294
rect -1878 188058 986 188294
rect 1222 188058 38186 188294
rect 38422 188058 75386 188294
rect 75622 188058 112586 188294
rect 112822 188058 149786 188294
rect 150022 188058 186986 188294
rect 187222 188058 224186 188294
rect 224422 188058 261386 188294
rect 261622 188058 298586 188294
rect 298822 188058 335786 188294
rect 336022 188058 372986 188294
rect 373222 188058 410186 188294
rect 410422 188058 447386 188294
rect 447622 188058 484586 188294
rect 484822 188058 521786 188294
rect 522022 188058 558986 188294
rect 559222 188058 585802 188294
rect 586038 188058 587160 188294
rect -3236 187876 587160 188058
rect -3236 154694 587160 154876
rect -3236 154458 -3054 154694
rect -2818 154458 4586 154694
rect 4822 154458 41786 154694
rect 42022 154458 78986 154694
rect 79222 154458 116186 154694
rect 116422 154458 153386 154694
rect 153622 154458 190586 154694
rect 190822 154458 227786 154694
rect 228022 154458 264986 154694
rect 265222 154458 302186 154694
rect 302422 154458 339386 154694
rect 339622 154458 376586 154694
rect 376822 154458 413786 154694
rect 414022 154458 450986 154694
rect 451222 154458 488186 154694
rect 488422 154458 525386 154694
rect 525622 154458 562586 154694
rect 562822 154458 586742 154694
rect 586978 154458 587160 154694
rect -3236 154276 587160 154458
rect -3236 151094 587160 151276
rect -3236 150858 -2114 151094
rect -1878 150858 986 151094
rect 1222 150858 38186 151094
rect 38422 150858 75386 151094
rect 75622 150858 112586 151094
rect 112822 150858 149786 151094
rect 150022 150858 186986 151094
rect 187222 150858 224186 151094
rect 224422 150858 261386 151094
rect 261622 150858 298586 151094
rect 298822 150858 335786 151094
rect 336022 150858 372986 151094
rect 373222 150858 410186 151094
rect 410422 150858 447386 151094
rect 447622 150858 484586 151094
rect 484822 150858 521786 151094
rect 522022 150858 558986 151094
rect 559222 150858 585802 151094
rect 586038 150858 587160 151094
rect -3236 150676 587160 150858
rect -3236 117494 587160 117676
rect -3236 117258 -3054 117494
rect -2818 117258 4586 117494
rect 4822 117258 41786 117494
rect 42022 117258 78986 117494
rect 79222 117258 116186 117494
rect 116422 117258 153386 117494
rect 153622 117258 190586 117494
rect 190822 117258 227786 117494
rect 228022 117258 264986 117494
rect 265222 117258 302186 117494
rect 302422 117258 339386 117494
rect 339622 117258 376586 117494
rect 376822 117258 413786 117494
rect 414022 117258 450986 117494
rect 451222 117258 488186 117494
rect 488422 117258 525386 117494
rect 525622 117258 562586 117494
rect 562822 117258 586742 117494
rect 586978 117258 587160 117494
rect -3236 117076 587160 117258
rect -3236 113894 587160 114076
rect -3236 113658 -2114 113894
rect -1878 113658 986 113894
rect 1222 113658 38186 113894
rect 38422 113658 75386 113894
rect 75622 113658 112586 113894
rect 112822 113658 149786 113894
rect 150022 113658 186986 113894
rect 187222 113658 224186 113894
rect 224422 113658 261386 113894
rect 261622 113658 298586 113894
rect 298822 113658 335786 113894
rect 336022 113658 372986 113894
rect 373222 113658 410186 113894
rect 410422 113658 447386 113894
rect 447622 113658 484586 113894
rect 484822 113658 521786 113894
rect 522022 113658 558986 113894
rect 559222 113658 585802 113894
rect 586038 113658 587160 113894
rect -3236 113476 587160 113658
rect -3236 80294 587160 80476
rect -3236 80058 -3054 80294
rect -2818 80058 4586 80294
rect 4822 80058 41786 80294
rect 42022 80058 78986 80294
rect 79222 80058 116186 80294
rect 116422 80058 153386 80294
rect 153622 80058 190586 80294
rect 190822 80058 227786 80294
rect 228022 80058 264986 80294
rect 265222 80058 302186 80294
rect 302422 80058 339386 80294
rect 339622 80058 376586 80294
rect 376822 80058 413786 80294
rect 414022 80058 450986 80294
rect 451222 80058 488186 80294
rect 488422 80058 525386 80294
rect 525622 80058 562586 80294
rect 562822 80058 586742 80294
rect 586978 80058 587160 80294
rect -3236 79876 587160 80058
rect -3236 76694 587160 76876
rect -3236 76458 -2114 76694
rect -1878 76458 986 76694
rect 1222 76458 38186 76694
rect 38422 76458 75386 76694
rect 75622 76458 112586 76694
rect 112822 76458 149786 76694
rect 150022 76458 186986 76694
rect 187222 76458 224186 76694
rect 224422 76458 261386 76694
rect 261622 76458 298586 76694
rect 298822 76458 335786 76694
rect 336022 76458 372986 76694
rect 373222 76458 410186 76694
rect 410422 76458 447386 76694
rect 447622 76458 484586 76694
rect 484822 76458 521786 76694
rect 522022 76458 558986 76694
rect 559222 76458 585802 76694
rect 586038 76458 587160 76694
rect -3236 76276 587160 76458
rect -3236 43094 587160 43276
rect -3236 42858 -3054 43094
rect -2818 42858 4586 43094
rect 4822 42858 41786 43094
rect 42022 42858 78986 43094
rect 79222 42858 116186 43094
rect 116422 42858 153386 43094
rect 153622 42858 190586 43094
rect 190822 42858 227786 43094
rect 228022 42858 264986 43094
rect 265222 42858 302186 43094
rect 302422 42858 339386 43094
rect 339622 42858 376586 43094
rect 376822 42858 413786 43094
rect 414022 42858 450986 43094
rect 451222 42858 488186 43094
rect 488422 42858 525386 43094
rect 525622 42858 562586 43094
rect 562822 42858 586742 43094
rect 586978 42858 587160 43094
rect -3236 42676 587160 42858
rect -3236 39494 587160 39676
rect -3236 39258 -2114 39494
rect -1878 39258 986 39494
rect 1222 39258 38186 39494
rect 38422 39258 75386 39494
rect 75622 39258 112586 39494
rect 112822 39258 149786 39494
rect 150022 39258 186986 39494
rect 187222 39258 224186 39494
rect 224422 39258 261386 39494
rect 261622 39258 298586 39494
rect 298822 39258 335786 39494
rect 336022 39258 372986 39494
rect 373222 39258 410186 39494
rect 410422 39258 447386 39494
rect 447622 39258 484586 39494
rect 484822 39258 521786 39494
rect 522022 39258 558986 39494
rect 559222 39258 585802 39494
rect 586038 39258 587160 39494
rect -3236 39076 587160 39258
rect -3236 5894 587160 6076
rect -3236 5658 -3054 5894
rect -2818 5658 4586 5894
rect 4822 5658 41786 5894
rect 42022 5658 78986 5894
rect 79222 5658 116186 5894
rect 116422 5658 153386 5894
rect 153622 5658 190586 5894
rect 190822 5658 227786 5894
rect 228022 5658 264986 5894
rect 265222 5658 302186 5894
rect 302422 5658 339386 5894
rect 339622 5658 376586 5894
rect 376822 5658 413786 5894
rect 414022 5658 450986 5894
rect 451222 5658 488186 5894
rect 488422 5658 525386 5894
rect 525622 5658 562586 5894
rect 562822 5658 586742 5894
rect 586978 5658 587160 5894
rect -3236 5476 587160 5658
rect -3236 2294 587160 2476
rect -3236 2058 -2114 2294
rect -1878 2058 986 2294
rect 1222 2058 38186 2294
rect 38422 2058 75386 2294
rect 75622 2058 112586 2294
rect 112822 2058 149786 2294
rect 150022 2058 186986 2294
rect 187222 2058 224186 2294
rect 224422 2058 261386 2294
rect 261622 2058 298586 2294
rect 298822 2058 335786 2294
rect 336022 2058 372986 2294
rect 373222 2058 410186 2294
rect 410422 2058 447386 2294
rect 447622 2058 484586 2294
rect 484822 2058 521786 2294
rect 522022 2058 558986 2294
rect 559222 2058 585802 2294
rect 586038 2058 587160 2294
rect -3236 1876 587160 2058
rect -2296 -806 586220 -624
rect -2296 -1042 -2114 -806
rect -1878 -1042 986 -806
rect 1222 -1042 38186 -806
rect 38422 -1042 75386 -806
rect 75622 -1042 112586 -806
rect 112822 -1042 149786 -806
rect 150022 -1042 186986 -806
rect 187222 -1042 224186 -806
rect 224422 -1042 261386 -806
rect 261622 -1042 298586 -806
rect 298822 -1042 335786 -806
rect 336022 -1042 372986 -806
rect 373222 -1042 410186 -806
rect 410422 -1042 447386 -806
rect 447622 -1042 484586 -806
rect 484822 -1042 521786 -806
rect 522022 -1042 558986 -806
rect 559222 -1042 585802 -806
rect 586038 -1042 586220 -806
rect -2296 -1224 586220 -1042
rect -3236 -1746 587160 -1564
rect -3236 -1982 -3054 -1746
rect -2818 -1982 4586 -1746
rect 4822 -1982 41786 -1746
rect 42022 -1982 78986 -1746
rect 79222 -1982 116186 -1746
rect 116422 -1982 153386 -1746
rect 153622 -1982 190586 -1746
rect 190822 -1982 227786 -1746
rect 228022 -1982 264986 -1746
rect 265222 -1982 302186 -1746
rect 302422 -1982 339386 -1746
rect 339622 -1982 376586 -1746
rect 376822 -1982 413786 -1746
rect 414022 -1982 450986 -1746
rect 451222 -1982 488186 -1746
rect 488422 -1982 525386 -1746
rect 525622 -1982 562586 -1746
rect 562822 -1982 586742 -1746
rect 586978 -1982 587160 -1746
rect -3236 -2164 587160 -1982
use mux16x1_project  mprj
timestamp 0
transform 1 0 520000 0 1 320000
box 0 552 10000 22000
use sky130_osu_ring_oscillator_mpr2ca_8_b0r1  ro1
timestamp 0
transform 1 0 292005 0 1 352000
box -5 0 17146 1776
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2296 -1224 -1696 705160 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2296 -1224 586220 -624 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2296 704560 586220 705160 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585620 -1224 586220 705160 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 804 -2164 1404 706100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 38004 -2164 38604 706100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 75204 -2164 75804 706100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 112404 -2164 113004 706100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 149604 -2164 150204 706100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 186804 -2164 187404 706100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 224004 -2164 224604 706100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 261204 -2164 261804 706100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 298404 -2164 299004 706100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 335604 -2164 336204 706100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 372804 -2164 373404 706100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 410004 -2164 410604 706100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 447204 -2164 447804 706100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 484404 -2164 485004 706100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 521604 -2164 522204 320008 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 521604 341752 522204 706100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 558804 -2164 559404 706100 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -3236 1876 587160 2476 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -3236 39076 587160 39676 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -3236 76276 587160 76876 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -3236 113476 587160 114076 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -3236 150676 587160 151276 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -3236 187876 587160 188476 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -3236 225076 587160 225676 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -3236 262276 587160 262876 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -3236 299476 587160 300076 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -3236 336676 587160 337276 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -3236 373876 587160 374476 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -3236 411076 587160 411676 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -3236 448276 587160 448876 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -3236 485476 587160 486076 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -3236 522676 587160 523276 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -3236 559876 587160 560476 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -3236 597076 587160 597676 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -3236 634276 587160 634876 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -3236 671476 587160 672076 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3236 -2164 -2636 706100 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -3236 -2164 587160 -1564 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -3236 705500 587160 706100 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 586560 -2164 587160 706100 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 4404 -2164 5004 706100 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 41604 -2164 42204 706100 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 78804 -2164 79404 706100 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 116004 -2164 116604 706100 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 153204 -2164 153804 706100 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 190404 -2164 191004 706100 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 227604 -2164 228204 706100 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 264804 -2164 265404 706100 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 302004 -2164 302604 706100 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 339204 -2164 339804 706100 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 376404 -2164 377004 706100 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 413604 -2164 414204 706100 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 450804 -2164 451404 706100 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 488004 -2164 488604 706100 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 525204 -2164 525804 320008 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 525204 341752 525804 706100 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal4 s 562404 -2164 563004 706100 0 FreeSans 3840 90 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -3236 5476 587160 6076 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -3236 42676 587160 43276 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -3236 79876 587160 80476 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -3236 117076 587160 117676 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -3236 154276 587160 154876 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -3236 191476 587160 192076 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -3236 228676 587160 229276 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -3236 265876 587160 266476 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -3236 303076 587160 303676 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -3236 340276 587160 340876 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -3236 377476 587160 378076 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -3236 414676 587160 415276 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -3236 451876 587160 452476 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -3236 489076 587160 489676 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -3236 526276 587160 526876 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -3236 563476 587160 564076 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -3236 600676 587160 601276 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -3236 637876 587160 638476 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal5 s -3236 675076 587160 675676 0 FreeSans 2560 0 0 0 vssd1
port 532 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 533 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 534 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 535 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 536 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 537 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 538 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 539 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 540 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 541 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 542 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 543 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 544 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 545 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 546 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 547 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 548 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 549 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 550 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 551 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 552 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 553 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 554 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 555 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 556 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 557 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 558 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 559 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 560 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 561 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 562 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 563 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 564 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 565 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 566 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 567 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 568 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 569 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 570 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 571 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 572 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 573 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 574 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 575 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 576 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 577 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 578 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 579 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 580 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 581 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 582 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 583 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 584 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 585 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 586 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 587 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 588 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 589 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 590 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 591 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 592 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 593 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 594 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 595 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 596 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 597 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 598 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 599 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 600 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 601 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 602 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 603 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 604 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 605 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 606 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 607 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 608 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 609 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 610 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 611 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 612 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 613 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 614 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 615 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 616 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 617 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 618 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 619 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 620 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 621 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 622 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 623 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 624 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 625 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 626 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 627 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 628 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 629 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 630 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 631 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 632 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 633 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 634 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 635 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 636 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 637 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 638 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
