magic
tech sky130A
magscale 1 2
timestamp 1710280277
<< nwell >>
rect -48 261 2440 582
<< pwell >>
rect 33 -17 67 17
rect 425 -17 459 17
rect 913 -17 947 17
rect 1401 -17 1435 17
rect 1793 -17 1827 17
<< nmos >>
rect 116 47 146 177
rect 212 47 242 177
rect 308 47 338 177
rect 508 47 538 177
rect 604 47 634 177
rect 700 47 730 177
rect 796 47 826 177
rect 996 47 1026 177
rect 1092 47 1122 177
rect 1188 47 1218 177
rect 1284 47 1314 177
rect 1484 47 1514 177
rect 1580 47 1610 177
rect 1676 47 1706 177
rect 1876 47 1906 177
rect 1972 47 2002 177
rect 2068 47 2098 177
rect 2164 47 2194 177
<< pmos >>
rect 116 297 146 497
rect 212 297 242 497
rect 308 297 338 497
rect 508 297 538 497
rect 604 297 634 497
rect 700 297 730 497
rect 796 297 826 497
rect 996 297 1026 497
rect 1092 297 1122 497
rect 1188 297 1218 497
rect 1284 297 1314 497
rect 1484 297 1514 497
rect 1580 297 1610 497
rect 1676 297 1706 497
rect 1876 297 1906 497
rect 1972 297 2002 497
rect 2068 297 2098 497
rect 2164 297 2194 497
<< ndiff >>
rect 58 101 116 177
rect 58 67 66 101
rect 100 67 116 101
rect 58 47 116 67
rect 146 101 212 177
rect 146 67 162 101
rect 196 67 212 101
rect 146 47 212 67
rect 242 47 308 177
rect 338 101 396 177
rect 338 67 354 101
rect 388 67 396 101
rect 338 47 396 67
rect 450 101 508 177
rect 450 67 458 101
rect 492 67 508 101
rect 450 47 508 67
rect 538 47 604 177
rect 634 101 700 177
rect 634 67 650 101
rect 684 67 700 101
rect 634 47 700 67
rect 730 47 796 177
rect 826 101 884 177
rect 826 67 842 101
rect 876 67 884 101
rect 826 47 884 67
rect 938 101 996 177
rect 938 67 946 101
rect 980 67 996 101
rect 938 47 996 67
rect 1026 47 1092 177
rect 1122 101 1188 177
rect 1122 67 1138 101
rect 1172 67 1188 101
rect 1122 47 1188 67
rect 1218 101 1284 177
rect 1218 67 1234 101
rect 1268 67 1284 101
rect 1218 47 1284 67
rect 1314 101 1372 177
rect 1314 67 1330 101
rect 1364 67 1372 101
rect 1314 47 1372 67
rect 1426 101 1484 177
rect 1426 67 1434 101
rect 1468 67 1484 101
rect 1426 47 1484 67
rect 1514 101 1580 177
rect 1514 67 1530 101
rect 1564 67 1580 101
rect 1514 47 1580 67
rect 1610 101 1676 177
rect 1610 67 1626 101
rect 1660 67 1676 101
rect 1610 47 1676 67
rect 1706 101 1764 177
rect 1706 67 1722 101
rect 1756 67 1764 101
rect 1706 47 1764 67
rect 1818 101 1876 177
rect 1818 67 1826 101
rect 1860 67 1876 101
rect 1818 47 1876 67
rect 1906 101 1972 177
rect 1906 67 1922 101
rect 1956 67 1972 101
rect 1906 47 1972 67
rect 2002 101 2068 177
rect 2002 67 2018 101
rect 2052 67 2068 101
rect 2002 47 2068 67
rect 2098 101 2164 177
rect 2098 67 2114 101
rect 2148 67 2164 101
rect 2098 47 2164 67
rect 2194 101 2252 177
rect 2194 67 2210 101
rect 2244 67 2252 101
rect 2194 47 2252 67
<< pdiff >>
rect 58 407 116 497
rect 58 373 66 407
rect 100 373 116 407
rect 58 297 116 373
rect 146 477 212 497
rect 146 443 162 477
rect 196 443 212 477
rect 146 297 212 443
rect 242 379 308 497
rect 242 345 258 379
rect 292 345 308 379
rect 242 297 308 345
rect 338 477 396 497
rect 338 443 354 477
rect 388 443 396 477
rect 338 297 396 443
rect 450 379 508 497
rect 450 345 458 379
rect 492 345 508 379
rect 450 297 508 345
rect 538 477 604 497
rect 538 443 554 477
rect 588 443 604 477
rect 538 297 604 443
rect 634 379 700 497
rect 634 345 650 379
rect 684 345 700 379
rect 634 297 700 345
rect 730 379 796 497
rect 730 345 746 379
rect 780 345 796 379
rect 730 297 796 345
rect 826 379 884 497
rect 826 345 842 379
rect 876 345 884 379
rect 826 297 884 345
rect 938 477 996 497
rect 938 443 946 477
rect 980 443 996 477
rect 938 297 996 443
rect 1026 379 1092 497
rect 1026 345 1042 379
rect 1076 345 1092 379
rect 1026 297 1092 345
rect 1122 477 1188 497
rect 1122 443 1138 477
rect 1172 443 1188 477
rect 1122 297 1188 443
rect 1218 297 1284 497
rect 1314 379 1372 497
rect 1314 345 1330 379
rect 1364 345 1372 379
rect 1314 297 1372 345
rect 1426 447 1484 497
rect 1426 413 1434 447
rect 1468 413 1484 447
rect 1426 297 1484 413
rect 1514 477 1580 497
rect 1514 443 1530 477
rect 1564 443 1580 477
rect 1514 297 1580 443
rect 1610 297 1676 497
rect 1706 379 1764 497
rect 1706 345 1722 379
rect 1756 345 1764 379
rect 1706 297 1764 345
rect 1818 379 1876 497
rect 1818 345 1826 379
rect 1860 345 1876 379
rect 1818 297 1876 345
rect 1906 297 1972 497
rect 2002 477 2068 497
rect 2002 443 2018 477
rect 2052 443 2068 477
rect 2002 297 2068 443
rect 2098 297 2164 497
rect 2194 379 2252 497
rect 2194 345 2210 379
rect 2244 345 2252 379
rect 2194 297 2252 345
<< ndiffc >>
rect 66 67 100 101
rect 162 67 196 101
rect 354 67 388 101
rect 458 67 492 101
rect 650 67 684 101
rect 842 67 876 101
rect 946 67 980 101
rect 1138 67 1172 101
rect 1234 67 1268 101
rect 1330 67 1364 101
rect 1434 67 1468 101
rect 1530 67 1564 101
rect 1626 67 1660 101
rect 1722 67 1756 101
rect 1826 67 1860 101
rect 1922 67 1956 101
rect 2018 67 2052 101
rect 2114 67 2148 101
rect 2210 67 2244 101
<< pdiffc >>
rect 66 373 100 407
rect 162 443 196 477
rect 258 345 292 379
rect 354 443 388 477
rect 458 345 492 379
rect 554 443 588 477
rect 650 345 684 379
rect 746 345 780 379
rect 842 345 876 379
rect 946 443 980 477
rect 1042 345 1076 379
rect 1138 443 1172 477
rect 1330 345 1364 379
rect 1434 413 1468 447
rect 1530 443 1564 477
rect 1722 345 1756 379
rect 1826 345 1860 379
rect 2018 443 2052 477
rect 2210 345 2244 379
<< poly >>
rect 116 497 146 523
rect 212 497 242 523
rect 308 497 338 523
rect 508 497 538 523
rect 604 497 634 523
rect 700 497 730 523
rect 796 497 826 523
rect 996 497 1026 523
rect 1092 497 1122 523
rect 1188 497 1218 523
rect 1284 497 1314 523
rect 1484 497 1514 523
rect 1580 497 1610 523
rect 1676 497 1706 523
rect 1876 497 1906 523
rect 1972 497 2002 523
rect 2068 497 2098 523
rect 2164 497 2194 523
rect 116 265 146 297
rect 212 265 242 297
rect 308 265 338 297
rect 508 265 538 297
rect 604 265 634 297
rect 700 265 730 297
rect 796 265 826 297
rect 996 265 1026 297
rect 1092 265 1122 297
rect 1188 265 1218 297
rect 1284 265 1314 297
rect 1484 265 1514 297
rect 1580 265 1610 297
rect 1676 265 1706 297
rect 1876 265 1906 297
rect 1972 265 2002 297
rect 2068 265 2098 297
rect 2164 265 2194 297
rect 104 249 158 265
rect 104 215 114 249
rect 148 215 158 249
rect 104 199 158 215
rect 200 249 254 265
rect 200 215 210 249
rect 244 215 254 249
rect 200 199 254 215
rect 296 249 350 265
rect 296 215 306 249
rect 340 215 350 249
rect 296 199 350 215
rect 496 249 550 265
rect 496 215 506 249
rect 540 215 550 249
rect 496 199 550 215
rect 592 249 646 265
rect 592 215 602 249
rect 636 215 646 249
rect 592 199 646 215
rect 688 249 742 265
rect 688 215 698 249
rect 732 215 742 249
rect 688 199 742 215
rect 784 249 838 265
rect 784 215 794 249
rect 828 215 838 249
rect 784 199 838 215
rect 984 249 1038 265
rect 984 215 994 249
rect 1028 215 1038 249
rect 984 199 1038 215
rect 1080 249 1134 265
rect 1080 215 1090 249
rect 1124 215 1134 249
rect 1080 199 1134 215
rect 1176 249 1230 265
rect 1176 215 1186 249
rect 1220 215 1230 249
rect 1176 199 1230 215
rect 1272 249 1326 265
rect 1272 215 1282 249
rect 1316 215 1326 249
rect 1272 199 1326 215
rect 1472 249 1526 265
rect 1472 215 1482 249
rect 1516 215 1526 249
rect 1472 199 1526 215
rect 1568 249 1622 265
rect 1568 215 1578 249
rect 1612 215 1622 249
rect 1568 199 1622 215
rect 1664 249 1718 265
rect 1664 215 1674 249
rect 1708 215 1718 249
rect 1664 199 1718 215
rect 1864 249 1918 265
rect 1864 215 1874 249
rect 1908 215 1918 249
rect 1864 199 1918 215
rect 1960 249 2014 265
rect 1960 215 1970 249
rect 2004 215 2014 249
rect 1960 199 2014 215
rect 2056 249 2110 265
rect 2056 215 2066 249
rect 2100 215 2110 249
rect 2056 199 2110 215
rect 2152 249 2206 265
rect 2152 215 2162 249
rect 2196 215 2206 249
rect 2152 199 2206 215
rect 116 177 146 199
rect 212 177 242 199
rect 308 177 338 199
rect 508 177 538 199
rect 604 177 634 199
rect 700 177 730 199
rect 796 177 826 199
rect 996 177 1026 199
rect 1092 177 1122 199
rect 1188 177 1218 199
rect 1284 177 1314 199
rect 1484 177 1514 199
rect 1580 177 1610 199
rect 1676 177 1706 199
rect 1876 177 1906 199
rect 1972 177 2002 199
rect 2068 177 2098 199
rect 2164 177 2194 199
rect 116 21 146 47
rect 212 21 242 47
rect 308 21 338 47
rect 508 21 538 47
rect 604 21 634 47
rect 700 21 730 47
rect 796 21 826 47
rect 996 21 1026 47
rect 1092 21 1122 47
rect 1188 21 1218 47
rect 1284 21 1314 47
rect 1484 21 1514 47
rect 1580 21 1610 47
rect 1676 21 1706 47
rect 1876 21 1906 47
rect 1972 21 2002 47
rect 2068 21 2098 47
rect 2164 21 2194 47
<< polycont >>
rect 114 215 148 249
rect 210 215 244 249
rect 306 215 340 249
rect 506 215 540 249
rect 602 215 636 249
rect 698 215 732 249
rect 794 215 828 249
rect 994 215 1028 249
rect 1090 215 1124 249
rect 1186 215 1220 249
rect 1282 215 1316 249
rect 1482 215 1516 249
rect 1578 215 1612 249
rect 1674 215 1708 249
rect 1874 215 1908 249
rect 1970 215 2004 249
rect 2066 215 2100 249
rect 2162 215 2196 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 162 477 196 527
rect 162 427 196 443
rect 354 477 388 527
rect 354 427 388 443
rect 554 477 588 527
rect 554 427 588 443
rect 946 477 980 527
rect 946 427 980 443
rect 1138 477 1172 527
rect 1530 477 1564 527
rect 1434 457 1468 463
rect 1138 427 1172 443
rect 66 357 100 373
rect 258 379 292 395
rect 746 379 780 395
rect 134 328 258 362
rect 442 345 458 379
rect 492 345 650 379
rect 684 345 700 379
rect 134 317 168 328
rect 114 283 168 317
rect 330 311 354 345
rect 1330 379 1364 423
rect 2018 477 2052 527
rect 1530 427 1564 443
rect 1660 423 1722 457
rect 1434 397 1468 413
rect 1026 345 1042 379
rect 1076 345 1124 379
rect 1698 379 1756 423
rect 1898 423 1922 457
rect 2018 427 2052 443
rect 1698 345 1722 379
rect 842 329 876 345
rect 1124 311 1292 345
rect 1330 329 1364 345
rect 114 269 148 283
rect 66 249 148 269
rect 66 215 114 249
rect 114 199 148 215
rect 210 249 244 265
rect 330 249 364 311
rect 602 249 636 255
rect 290 215 306 249
rect 340 215 364 249
rect 441 233 506 249
rect 475 215 506 233
rect 540 215 556 249
rect 602 199 636 215
rect 698 249 732 265
rect 946 249 980 311
rect 1258 265 1292 311
rect 1722 329 1756 345
rect 1826 379 1860 395
rect 1468 311 1612 317
rect 1898 345 1932 423
rect 2066 345 2210 379
rect 2244 345 2260 379
rect 1898 311 1922 345
rect 1434 283 1612 311
rect 1090 249 1124 265
rect 778 215 794 249
rect 828 233 876 249
rect 828 215 842 233
rect 946 215 994 249
rect 1028 215 1044 249
rect 1186 249 1220 265
rect 1258 249 1316 265
rect 1578 249 1612 283
rect 1674 255 1722 269
rect 1674 249 1756 255
rect 1898 249 1932 311
rect 1258 215 1282 249
rect 1282 199 1316 215
rect 1434 233 1482 249
rect 1468 215 1482 233
rect 1516 215 1532 249
rect 1658 215 1674 249
rect 1708 235 1756 249
rect 1708 215 1724 235
rect 1858 215 1874 249
rect 1908 215 1932 249
rect 1970 249 2004 265
rect 2162 249 2196 255
rect 2004 215 2066 249
rect 2100 215 2116 249
rect 1578 199 1612 215
rect 2162 199 2196 215
rect 66 51 100 67
rect 162 101 196 117
rect 458 101 492 117
rect 292 87 354 101
rect 258 67 354 87
rect 388 67 404 101
rect 634 67 650 101
rect 684 87 746 101
rect 684 67 780 87
rect 842 101 876 117
rect 930 67 946 101
rect 980 87 1042 101
rect 980 67 1076 87
rect 1138 101 1172 117
rect 162 17 196 67
rect 458 17 492 67
rect 842 17 876 67
rect 1138 17 1172 67
rect 1234 51 1268 67
rect 1330 101 1364 117
rect 1330 17 1364 67
rect 1434 51 1468 67
rect 1530 101 1564 117
rect 1530 17 1564 67
rect 1626 51 1660 67
rect 1722 101 1756 117
rect 1722 17 1756 67
rect 1826 101 1860 117
rect 1826 17 1860 67
rect 1922 51 1956 67
rect 2018 101 2052 117
rect 2018 17 2052 67
rect 2114 51 2148 67
rect 2210 101 2244 117
rect 2210 17 2244 67
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 66 407 100 429
rect 66 395 100 407
rect 1330 423 1364 457
rect 650 379 684 401
rect 650 367 684 379
rect 258 311 292 345
rect 354 311 388 345
rect 746 311 780 345
rect 842 379 876 401
rect 1434 447 1468 457
rect 1434 423 1468 447
rect 1626 423 1660 457
rect 1722 423 1756 457
rect 842 367 876 379
rect 1922 423 1956 457
rect 946 311 980 345
rect 1090 311 1124 345
rect 602 255 636 289
rect 210 215 244 233
rect 210 199 244 215
rect 441 199 475 233
rect 1434 311 1468 345
rect 1826 311 1860 345
rect 1922 311 1956 345
rect 2066 311 2100 345
rect 698 215 732 233
rect 698 199 732 215
rect 842 199 876 233
rect 1090 215 1124 233
rect 1090 199 1124 215
rect 1186 215 1220 233
rect 1722 255 1756 289
rect 1186 199 1220 215
rect 1434 199 1468 233
rect 2162 255 2196 289
rect 1970 215 2004 233
rect 1970 199 2004 215
rect 66 101 100 121
rect 66 87 100 101
rect 258 87 292 121
rect 746 87 780 121
rect 1042 87 1076 121
rect 1234 101 1268 121
rect 1234 87 1268 101
rect 1434 101 1468 121
rect 1434 87 1468 101
rect 1626 101 1660 121
rect 1626 87 1660 101
rect 1922 101 1956 121
rect 1922 87 1956 101
rect 2114 101 2148 121
rect 2114 87 2148 101
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
<< metal1 >>
rect 0 561 2392 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 0 521 2392 527
rect 51 429 115 435
rect 51 410 66 429
rect 100 410 115 429
rect 51 358 57 410
rect 109 358 115 410
rect 653 407 873 421
rect 1003 414 1009 466
rect 1061 454 1067 466
rect 1061 426 1217 454
rect 1061 414 1067 426
rect 638 401 888 407
rect 638 367 650 401
rect 684 393 842 401
rect 684 367 696 393
rect 638 361 696 367
rect 830 367 842 393
rect 876 367 888 401
rect 830 361 888 367
rect 51 352 115 358
rect 67 127 98 352
rect 243 302 249 354
rect 301 302 307 354
rect 339 302 345 354
rect 397 302 403 354
rect 467 302 473 354
rect 525 330 531 354
rect 734 345 792 351
rect 525 302 633 330
rect 734 311 746 345
rect 780 342 792 345
rect 780 311 801 342
rect 734 305 801 311
rect 590 295 633 302
rect 590 289 648 295
rect 590 255 602 289
rect 636 255 648 289
rect 590 249 648 255
rect 686 242 744 248
rect 147 190 153 242
rect 205 239 211 242
rect 205 238 256 239
rect 205 233 337 238
rect 205 199 210 233
rect 244 210 337 233
rect 429 233 487 239
rect 429 230 441 233
rect 244 199 256 210
rect 205 193 256 199
rect 309 202 337 210
rect 409 202 441 230
rect 309 199 441 202
rect 475 199 487 233
rect 686 202 689 242
rect 309 193 487 199
rect 205 190 211 193
rect 309 174 437 193
rect 533 190 689 202
rect 741 190 744 242
rect 533 174 744 190
rect 54 121 112 127
rect 54 87 66 121
rect 100 87 112 121
rect 54 81 112 87
rect 243 78 249 130
rect 301 118 307 130
rect 635 118 641 130
rect 301 90 641 118
rect 301 78 307 90
rect 635 78 641 90
rect 693 78 699 130
rect 773 127 801 305
rect 931 302 937 354
rect 989 302 995 354
rect 1075 302 1081 354
rect 1133 302 1139 354
rect 1189 342 1217 426
rect 1315 414 1321 466
rect 1373 414 1379 466
rect 1422 457 1480 463
rect 1422 423 1434 457
rect 1468 454 1480 457
rect 1515 454 1521 466
rect 1468 426 1521 454
rect 1468 423 1480 426
rect 1422 417 1480 423
rect 1515 414 1521 426
rect 1573 414 1579 466
rect 1611 414 1617 466
rect 1669 414 1675 466
rect 1707 414 1713 466
rect 1765 414 1771 466
rect 1907 414 1913 466
rect 1965 421 1971 466
rect 1965 414 2193 421
rect 1925 393 2193 414
rect 1422 345 1480 351
rect 1422 342 1434 345
rect 1189 314 1434 342
rect 1422 311 1434 314
rect 1468 311 1480 345
rect 1422 305 1480 311
rect 1811 302 1817 354
rect 1869 302 1875 354
rect 1925 351 1953 393
rect 1910 345 1968 351
rect 1910 311 1922 345
rect 1956 311 1968 345
rect 1910 305 1968 311
rect 2054 345 2112 351
rect 2054 311 2066 345
rect 2100 342 2112 345
rect 2100 311 2121 342
rect 2054 305 2121 311
rect 1710 289 1768 295
rect 1710 255 1722 289
rect 1756 286 1768 289
rect 1811 286 1857 302
rect 1756 258 1857 286
rect 1756 255 1768 258
rect 1710 249 1768 255
rect 879 239 885 242
rect 830 233 885 239
rect 830 199 842 233
rect 876 199 885 233
rect 830 193 885 199
rect 879 190 885 193
rect 937 230 943 242
rect 1078 233 1136 239
rect 1078 230 1090 233
rect 937 202 1090 230
rect 937 190 943 202
rect 1078 199 1090 202
rect 1124 199 1136 233
rect 1078 193 1136 199
rect 1174 233 1232 239
rect 1174 199 1186 233
rect 1220 230 1232 233
rect 1220 202 1361 230
rect 1220 199 1232 202
rect 1174 193 1232 199
rect 734 121 801 127
rect 734 87 746 121
rect 780 118 801 121
rect 931 118 937 130
rect 780 90 937 118
rect 780 87 792 90
rect 734 81 792 87
rect 931 78 937 90
rect 989 78 995 130
rect 1075 127 1081 130
rect 1030 121 1081 127
rect 1030 87 1042 121
rect 1076 87 1081 121
rect 1030 81 1081 87
rect 1075 78 1081 81
rect 1133 78 1139 130
rect 1219 78 1225 130
rect 1277 78 1283 130
rect 1333 118 1361 202
rect 1419 190 1425 242
rect 1477 202 1483 242
rect 1958 233 2016 239
rect 1958 202 1970 233
rect 1477 199 1970 202
rect 2004 199 2016 233
rect 1477 193 2016 199
rect 1477 190 2001 193
rect 1437 174 2001 190
rect 2093 130 2121 305
rect 2165 295 2193 393
rect 2150 289 2208 295
rect 2150 255 2162 289
rect 2196 255 2208 289
rect 2150 249 2208 255
rect 1467 127 1473 130
rect 1422 121 1473 127
rect 1422 118 1434 121
rect 1333 90 1434 118
rect 1422 87 1434 90
rect 1468 87 1473 121
rect 1422 81 1473 87
rect 1467 78 1473 81
rect 1525 78 1531 130
rect 1587 78 1593 130
rect 1645 121 1723 130
rect 1660 87 1723 121
rect 1645 78 1723 87
rect 1811 78 1817 130
rect 1869 118 1875 130
rect 1910 121 1968 127
rect 1910 118 1922 121
rect 1869 90 1922 118
rect 1869 78 1875 90
rect 1910 87 1922 90
rect 1956 87 1968 121
rect 2093 90 2105 130
rect 1910 81 1968 87
rect 2099 78 2105 90
rect 2157 78 2163 130
rect 0 17 2392 23
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
rect 0 -48 2392 -17
<< via1 >>
rect 57 395 66 410
rect 66 395 100 410
rect 100 395 109 410
rect 57 358 109 395
rect 1009 414 1061 466
rect 249 345 301 354
rect 249 311 258 345
rect 258 311 292 345
rect 292 311 301 345
rect 249 302 301 311
rect 345 345 397 354
rect 345 311 354 345
rect 354 311 388 345
rect 388 311 397 345
rect 345 302 397 311
rect 473 302 525 354
rect 153 190 205 242
rect 689 233 741 242
rect 689 199 698 233
rect 698 199 732 233
rect 732 199 741 233
rect 689 190 741 199
rect 249 121 301 130
rect 249 87 258 121
rect 258 87 292 121
rect 292 87 301 121
rect 249 78 301 87
rect 641 78 693 130
rect 937 345 989 354
rect 937 311 946 345
rect 946 311 980 345
rect 980 311 989 345
rect 937 302 989 311
rect 1081 345 1133 354
rect 1081 311 1090 345
rect 1090 311 1124 345
rect 1124 311 1133 345
rect 1081 302 1133 311
rect 1321 457 1373 466
rect 1321 423 1330 457
rect 1330 423 1364 457
rect 1364 423 1373 457
rect 1321 414 1373 423
rect 1521 414 1573 466
rect 1617 457 1669 466
rect 1617 423 1626 457
rect 1626 423 1660 457
rect 1660 423 1669 457
rect 1617 414 1669 423
rect 1713 457 1765 466
rect 1713 423 1722 457
rect 1722 423 1756 457
rect 1756 423 1765 457
rect 1713 414 1765 423
rect 1913 457 1965 466
rect 1913 423 1922 457
rect 1922 423 1956 457
rect 1956 423 1965 457
rect 1913 414 1965 423
rect 1817 345 1869 354
rect 1817 311 1826 345
rect 1826 311 1860 345
rect 1860 311 1869 345
rect 1817 302 1869 311
rect 885 190 937 242
rect 937 78 989 130
rect 1081 78 1133 130
rect 1225 121 1277 130
rect 1225 87 1234 121
rect 1234 87 1268 121
rect 1268 87 1277 121
rect 1225 78 1277 87
rect 1425 233 1477 242
rect 1425 199 1434 233
rect 1434 199 1468 233
rect 1468 199 1477 233
rect 1425 190 1477 199
rect 1473 78 1525 130
rect 1593 121 1645 130
rect 1593 87 1626 121
rect 1626 87 1645 121
rect 1593 78 1645 87
rect 1817 78 1869 130
rect 2105 121 2157 130
rect 2105 87 2114 121
rect 2114 87 2148 121
rect 2148 87 2157 121
rect 2105 78 2157 87
<< metal2 >>
rect 55 468 111 477
rect 55 410 111 412
rect 55 403 57 410
rect 109 403 111 410
rect 1009 466 1061 472
rect 1009 408 1061 414
rect 1319 468 1375 477
rect 543 360 599 365
rect 57 352 109 358
rect 249 354 301 360
rect 345 354 397 360
rect 249 296 301 302
rect 333 302 345 342
rect 333 296 397 302
rect 473 356 599 360
rect 473 354 543 356
rect 525 302 543 354
rect 473 300 543 302
rect 937 354 989 360
rect 599 314 937 342
rect 473 296 599 300
rect 937 296 989 302
rect 151 244 207 253
rect 151 179 207 188
rect 261 136 289 296
rect 333 230 361 296
rect 543 291 599 296
rect 395 244 451 253
rect 831 248 887 253
rect 333 202 395 230
rect 689 242 741 248
rect 451 202 689 230
rect 395 179 451 188
rect 689 184 741 190
rect 831 244 937 248
rect 887 242 937 244
rect 887 188 937 190
rect 831 184 937 188
rect 831 179 887 184
rect 249 130 301 136
rect 249 72 301 78
rect 641 130 693 136
rect 937 130 989 136
rect 693 90 849 118
rect 641 72 693 78
rect 821 42 849 90
rect 1021 118 1049 408
rect 1319 403 1375 412
rect 1521 466 1573 472
rect 1521 408 1573 414
rect 1617 466 1669 472
rect 1617 408 1669 414
rect 1711 468 1767 477
rect 1333 365 1361 403
rect 1079 356 1135 365
rect 1295 342 1361 365
rect 1079 291 1135 300
rect 1237 314 1361 342
rect 1093 136 1121 291
rect 1237 136 1265 314
rect 1295 291 1351 314
rect 1425 242 1477 248
rect 1309 202 1425 230
rect 989 90 1049 118
rect 1081 130 1133 136
rect 937 72 989 78
rect 1081 72 1133 78
rect 1225 130 1277 136
rect 1225 72 1277 78
rect 1309 42 1337 202
rect 1425 184 1477 190
rect 1533 136 1561 408
rect 1617 398 1657 408
rect 1711 403 1767 412
rect 1911 468 1967 477
rect 1911 403 1967 412
rect 1605 365 1657 398
rect 1605 291 1705 365
rect 1817 354 1869 360
rect 1817 296 1869 302
rect 1605 136 1633 291
rect 1829 136 1857 296
rect 1473 130 1561 136
rect 1525 90 1561 130
rect 1593 130 1645 136
rect 1473 72 1525 78
rect 1593 72 1645 78
rect 1817 130 1869 136
rect 1817 72 1869 78
rect 2103 132 2159 141
rect 2103 67 2159 76
rect 821 14 1337 42
<< via2 >>
rect 55 412 111 468
rect 1319 466 1375 468
rect 1319 414 1321 466
rect 1321 414 1373 466
rect 1373 414 1375 466
rect 1319 412 1375 414
rect 543 300 599 356
rect 151 242 207 244
rect 151 190 153 242
rect 153 190 205 242
rect 205 190 207 242
rect 151 188 207 190
rect 395 188 451 244
rect 831 242 887 244
rect 831 190 885 242
rect 885 190 887 242
rect 831 188 887 190
rect 1711 466 1767 468
rect 1711 414 1713 466
rect 1713 414 1765 466
rect 1765 414 1767 466
rect 1711 412 1767 414
rect 1079 354 1135 356
rect 1079 302 1081 354
rect 1081 302 1133 354
rect 1133 302 1135 354
rect 1079 300 1135 302
rect 1911 466 1967 468
rect 1911 414 1913 466
rect 1913 414 1965 466
rect 1965 414 1967 466
rect 1911 412 1967 414
rect 2103 130 2159 132
rect 2103 78 2105 130
rect 2105 78 2157 130
rect 2157 78 2159 130
rect 2103 76 2159 78
<< metal3 >>
rect 50 468 196 473
rect 50 412 55 468
rect 111 412 196 468
rect 50 407 196 412
rect 1314 468 1460 473
rect 1314 412 1319 468
rect 1375 412 1460 468
rect 1314 407 1460 412
rect 1654 468 1800 473
rect 1654 412 1711 468
rect 1767 412 1800 468
rect 1654 407 1800 412
rect 1861 468 1972 473
rect 1861 412 1911 468
rect 1967 412 1972 468
rect 1861 407 1972 412
rect 538 356 684 361
rect 538 300 543 356
rect 599 300 684 356
rect 538 295 684 300
rect 1074 356 1185 361
rect 1074 300 1079 356
rect 1135 300 1185 356
rect 1074 295 1185 300
rect 116 244 262 249
rect 116 188 151 244
rect 207 188 262 244
rect 116 183 262 188
rect 323 244 469 249
rect 323 188 395 244
rect 451 188 469 244
rect 323 183 469 188
rect 826 244 972 249
rect 826 188 831 244
rect 887 188 972 244
rect 826 183 972 188
rect 1125 134 1185 295
rect 1861 134 1921 407
rect 1125 74 1921 134
rect 2098 132 2244 137
rect 2098 76 2103 132
rect 2159 76 2244 132
rect 2098 71 2244 76
<< labels >>
flabel nwell s 1793 527 1827 561 0 FreeSans 100 0 0 0 VPB
port 1 nsew
flabel nwell s 1401 527 1435 561 0 FreeSans 100 0 0 0 VPB
port 1 nsew
flabel nwell s 913 527 947 561 0 FreeSans 100 0 0 0 VPB
port 1 nsew
flabel nwell s 425 527 459 561 0 FreeSans 100 0 0 0 VPB
port 1 nsew
flabel nwell s 33 527 67 561 0 FreeSans 100 0 0 0 VPB
port 1 nsew
flabel pwell s 1793 -17 1827 17 0 FreeSans 100 0 0 0 VNB
port 2 nsew
flabel pwell s 1401 -17 1435 17 0 FreeSans 100 0 0 0 VNB
port 2 nsew
flabel pwell s 913 -17 947 17 0 FreeSans 100 0 0 0 VNB
port 2 nsew
flabel pwell s 425 -17 459 17 0 FreeSans 100 0 0 0 VNB
port 2 nsew
flabel pwell s 33 -17 67 17 0 FreeSans 100 0 0 0 VNB
port 2 nsew
flabel comment s 0 0 0 0 0 FreeSans 100 0 0 0 mul2
rlabel metal3 s 323 183 469 249 4 B0
port 3 nsew
rlabel metal3 s 116 183 262 249 4 A0
port 4 nsew
rlabel metal3 s 538 295 684 361 4 B1
port 5 nsew
rlabel metal3 s 1654 407 1800 473 4 R1
port 6 nsew
rlabel metal3 s 1314 407 1460 473 4 R2
port 7 nsew
rlabel metal3 s 50 407 196 473 4 R0
port 8 nsew
rlabel metal3 s 2098 71 2244 137 4 R3
port 9 nsew
rlabel metal3 s 826 183 972 249 4 A1
port 10 nsew
flabel metal1 s 31 527 65 561 0 FreeSans 100 0 0 0 vpwr
port 11 nsew
flabel metal1 s 31 -17 65 17 0 FreeSans 100 0 0 0 vgnd
port 12 nsew
<< properties >>
string FIXED_BBOX 0 0 2392 544
<< end >>
