magic
tech sky130A
magscale 1 2
timestamp 1714079683
<< nwell >>
rect 0 1626 702 1748
rect 0 1406 706 1626
rect 2147 1645 2337 1748
rect 2147 1408 2342 1645
rect 2364 1630 2429 1695
rect 3045 1689 3046 1720
rect 3273 1408 3318 1748
rect 0 1391 716 1406
rect 0 1360 757 1391
rect 0 1128 759 1360
rect 2130 1193 3318 1408
rect 0 1097 757 1128
rect 0 1085 746 1097
rect 2104 1086 3318 1193
rect 0 866 706 1085
rect 2120 1058 2342 1086
rect 1697 1029 2342 1058
rect 2120 943 2342 1029
rect 2121 924 2342 943
rect 2101 921 2342 924
rect 2121 901 2342 921
rect 0 861 720 866
rect 2120 862 2342 901
rect 2161 861 2342 862
rect 0 742 640 861
rect 2179 744 2342 861
rect 3124 772 3154 807
rect 3273 744 3318 1086
<< pwell >>
rect 1229 1612 1280 1656
<< ndiff >>
rect 3209 442 3244 476
<< psubdiff >>
rect 2367 2172 2379 2206
rect 2505 2172 2580 2206
<< locali >>
rect 1 2182 3318 2492
rect 1 2172 802 2182
rect 646 2171 802 2172
rect 744 1700 802 2171
rect 858 1700 914 2182
rect 970 1700 1026 2182
rect 1082 1700 1138 2182
rect 1194 1700 1250 2182
rect 1306 1700 1362 2182
rect 1418 1700 1474 2182
rect 1530 1700 1586 2182
rect 1642 1700 1698 2182
rect 1754 1700 1810 2182
rect 1866 1700 1922 2182
rect 1978 1700 2034 2182
rect 2090 2172 3318 2182
rect 2090 1700 2125 2172
rect 2893 1868 2948 1884
rect 2847 1850 2948 1868
rect 3011 1720 3145 1754
rect 2124 1671 2125 1700
rect 3045 1689 3046 1720
rect 3210 1461 3244 1495
rect 1 1360 716 1405
rect 1 1128 759 1360
rect 2130 1193 3318 1408
rect 1 1127 750 1128
rect 1 1085 746 1127
rect 2104 1086 3318 1193
rect 3210 998 3244 1032
rect 3042 726 3158 760
rect 2847 624 2975 642
rect 693 600 759 619
rect 2124 618 2162 619
rect 2098 615 2162 618
rect 693 321 752 600
rect 2123 590 2162 615
rect 810 321 868 590
rect 926 321 984 590
rect 1042 321 1100 590
rect 1158 321 1216 590
rect 1274 321 1331 590
rect 1389 321 1447 590
rect 1505 321 1563 590
rect 1621 321 1679 590
rect 1737 321 1794 590
rect 1852 321 1910 590
rect 1968 321 2026 590
rect 2084 321 2162 590
rect 2893 608 2975 624
rect 693 320 2162 321
rect 1 0 3318 320
<< viali >>
rect 2847 1868 2893 1914
rect 3209 1742 3243 1776
rect 2847 578 2893 624
rect 3210 442 3244 476
<< metal1 >>
rect 1 2182 3318 2492
rect 1 2172 802 2182
rect 289 2170 324 2172
rect 646 2171 802 2172
rect 289 1720 323 2170
rect 388 1926 462 1935
rect 388 1870 397 1926
rect 453 1870 462 1926
rect 388 1861 462 1870
rect 488 1783 494 1839
rect 550 1783 556 1839
rect 744 1706 802 2171
rect 858 1706 914 2182
rect 970 1706 1026 2182
rect 1082 1706 1138 2182
rect 1194 1706 1250 2182
rect 1306 1706 1362 2182
rect 1418 1706 1474 2182
rect 1530 1706 1586 2182
rect 1642 1706 1698 2182
rect 1754 1706 1810 2182
rect 1866 1706 1922 2182
rect 1978 1706 2034 2182
rect 2090 2172 3318 2182
rect 2090 1706 2125 2172
rect 2835 1915 2905 1920
rect 2687 1914 2905 1915
rect 2687 1908 2847 1914
rect 2699 1902 2847 1908
rect 2653 1881 2847 1902
rect 2653 1868 2699 1881
rect 2835 1868 2847 1881
rect 2893 1868 2905 1914
rect 2835 1862 2905 1868
rect 2732 1846 2797 1853
rect 2732 1794 2739 1846
rect 2791 1794 2797 1846
rect 2732 1788 2797 1794
rect 2572 1772 2636 1778
rect 2572 1720 2578 1772
rect 2630 1720 2636 1772
rect 2572 1713 2636 1720
rect 116 1635 122 1691
rect 178 1673 184 1691
rect 578 1673 584 1691
rect 178 1639 584 1673
rect 178 1635 184 1639
rect 578 1635 584 1639
rect 640 1635 646 1691
rect 1229 1580 1281 1680
rect 2124 1665 2125 1706
rect 2364 1688 2429 1695
rect 2364 1636 2371 1688
rect 2423 1636 2429 1688
rect 2364 1630 2429 1636
rect 1 1391 716 1405
rect 1 1360 757 1391
rect 1 1128 759 1360
rect 2130 1193 3318 1408
rect 1 1097 757 1128
rect 1 1085 746 1097
rect 2104 1089 3318 1193
rect 2105 1086 3318 1089
rect 2363 1044 2428 1051
rect 2363 992 2370 1044
rect 2422 992 2428 1044
rect 2363 986 2428 992
rect 1933 893 2015 921
rect 2378 846 2414 986
rect 2572 790 2636 796
rect 2572 772 2578 790
rect 2509 738 2578 772
rect 2630 738 2636 790
rect 2572 732 2636 738
rect 2238 716 2303 723
rect 2238 664 2245 716
rect 2297 698 2303 716
rect 2727 716 2797 722
rect 2297 664 2722 698
rect 2238 658 2303 664
rect 2727 658 2733 716
rect 2791 658 2797 716
rect 2727 652 2797 658
rect 693 600 761 625
rect 2124 618 2162 625
rect 2835 624 2905 630
rect 693 321 752 600
rect 2123 590 2162 618
rect 2653 623 2687 624
rect 2699 623 2847 624
rect 2653 590 2847 623
rect 810 321 868 590
rect 926 321 984 590
rect 1042 321 1100 590
rect 1158 321 1216 590
rect 1274 321 1331 590
rect 1389 321 1447 590
rect 1505 321 1563 590
rect 1621 321 1679 590
rect 1737 321 1794 590
rect 1852 321 1910 590
rect 1968 321 2026 590
rect 2084 321 2162 590
rect 2835 578 2847 590
rect 2893 578 2905 624
rect 2835 572 2905 578
rect 693 320 2162 321
rect 1 0 3318 320
<< via1 >>
rect 397 1870 453 1926
rect 494 1783 550 1839
rect 2739 1794 2791 1846
rect 2578 1720 2630 1772
rect 122 1635 178 1691
rect 584 1635 640 1691
rect 2371 1636 2423 1688
rect 2370 992 2422 1044
rect 2578 738 2630 790
rect 2245 664 2297 716
rect 2733 658 2791 716
<< metal2 >>
rect 505 1941 2541 1975
rect 388 1926 462 1935
rect 388 1870 397 1926
rect 453 1870 462 1926
rect 388 1861 462 1870
rect 505 1845 539 1941
rect 595 1860 2412 1894
rect 494 1839 550 1845
rect 494 1777 550 1783
rect 122 1691 178 1700
rect 595 1697 629 1860
rect 122 1626 178 1635
rect 584 1691 640 1697
rect 2377 1695 2412 1860
rect 2509 1840 2541 1941
rect 2732 1846 2797 1853
rect 2732 1840 2739 1846
rect 2509 1806 2739 1840
rect 584 1629 640 1635
rect 2364 1688 2429 1695
rect 2364 1636 2371 1688
rect 2423 1636 2429 1688
rect 2364 1630 2429 1636
rect 2377 1051 2412 1630
rect 2363 1044 2428 1051
rect 2363 992 2370 1044
rect 2422 992 2428 1044
rect 2363 986 2428 992
rect 2509 772 2541 1806
rect 2732 1794 2739 1806
rect 2791 1794 2797 1846
rect 2732 1788 2797 1794
rect 2572 1772 2636 1778
rect 2572 1720 2578 1772
rect 2630 1720 2636 1772
rect 2572 1713 2636 1720
rect 2578 1666 2612 1713
rect 2578 1631 2613 1666
rect 2578 1596 2773 1631
rect 2572 790 2636 796
rect 2572 772 2578 790
rect 1305 614 1339 764
rect 2509 738 2578 772
rect 2630 738 2636 790
rect 2572 732 2636 738
rect 2238 716 2303 723
rect 2738 722 2773 1596
rect 2238 664 2245 716
rect 2297 664 2303 716
rect 2238 658 2303 664
rect 2727 716 2797 722
rect 2727 658 2733 716
rect 2791 658 2797 716
rect 2253 614 2287 658
rect 2727 652 2797 658
rect 1305 580 2287 614
<< via2 >>
rect 397 1870 453 1926
rect 122 1635 178 1691
<< metal3 >>
rect 116 1691 184 2492
rect 388 1926 462 1935
rect 388 1870 397 1926
rect 453 1923 462 1926
rect 453 1870 1419 1923
rect 388 1863 1419 1870
rect 388 1861 462 1863
rect 116 1635 122 1691
rect 178 1635 184 1691
rect 116 1626 184 1635
rect 1358 1484 1418 1863
rect 1232 1481 1420 1484
rect 1232 1478 1608 1481
rect 1232 1418 1621 1478
rect 1232 1416 1359 1418
rect 1232 1078 1292 1416
rect 1427 1276 1434 1280
rect 1427 1216 1493 1276
rect 1232 1012 1763 1078
rect 1703 1011 1763 1012
rect 1703 810 1763 872
rect 1699 805 1763 810
use scs130hd_mpr2ca_8  scs130hd_mpr2ca_8_0
timestamp 1714079683
transform 1 0 744 0 1 601
box -98 -60 1418 1148
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_1
timestamp 1714057206
transform 1 0 2891 0 1 260
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_2
timestamp 1714057206
transform 1 0 3089 0 1 260
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_3
timestamp 1714057206
transform 1 0 3089 0 -1 2232
box -10 0 199 902
use sky130_osu_sc_12T_hs__inv_1  sky130_osu_sc_12T_hs__inv_1_4
timestamp 1714057206
transform 1 0 2891 0 -1 2232
box -10 0 199 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_0
timestamp 1714057206
transform 1 0 2342 0 1 260
box -10 0 552 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_1
timestamp 1714057206
transform 1 0 97 0 -1 2231
box -10 0 552 902
use sky130_osu_sc_12T_hs__mux2_1  sky130_osu_sc_12T_hs__mux2_1_2
timestamp 1714057206
transform 1 0 2342 0 -1 2232
box -10 0 552 902
<< labels >>
rlabel via1 2397 1019 2397 1019 1 sel
port 8 n
rlabel metal1 63 1349 63 1349 1 vccd1
port 6 n
rlabel via1 536 1810 536 1810 1 in
port 9 n
rlabel viali 3210 442 3244 476 1 Y1
port 11 n
rlabel metal1 60 291 60 291 1 vssd1
port 5 n
rlabel viali 3209 1742 3243 1776 1 Y0
port 10 n
<< end >>
