magic
tech sky130A
magscale 1 2
timestamp 1713287902
<< nwell >>
rect -48 260 2440 582
<< pwell >>
rect 32 -12 66 16
rect 28 -16 66 -12
rect 28 -18 62 -16
rect 424 -18 458 16
rect 912 -18 946 16
rect 1400 -18 1434 16
rect 1792 -18 1826 16
<< nmos >>
rect 116 46 146 176
rect 212 46 242 176
rect 308 46 338 176
rect 508 46 538 176
rect 604 46 634 176
rect 700 46 730 176
rect 796 46 826 176
rect 996 46 1026 176
rect 1092 46 1122 176
rect 1188 46 1218 176
rect 1284 46 1314 176
rect 1484 46 1514 176
rect 1580 46 1610 176
rect 1676 46 1706 176
rect 1876 46 1906 176
rect 1972 46 2002 176
rect 2068 46 2098 176
rect 2164 46 2194 176
<< pmos >>
rect 116 296 146 496
rect 212 296 242 496
rect 308 296 338 496
rect 508 296 538 496
rect 604 296 634 496
rect 700 296 730 496
rect 796 296 826 496
rect 996 296 1026 496
rect 1092 296 1122 496
rect 1188 296 1218 496
rect 1284 296 1314 496
rect 1484 296 1514 496
rect 1580 296 1610 496
rect 1676 296 1706 496
rect 1876 296 1906 496
rect 1972 296 2002 496
rect 2068 296 2098 496
rect 2164 296 2194 496
<< ndiff >>
rect 58 100 116 176
rect 58 66 66 100
rect 100 66 116 100
rect 58 46 116 66
rect 146 100 212 176
rect 146 66 162 100
rect 196 66 212 100
rect 146 46 212 66
rect 242 46 308 176
rect 338 100 396 176
rect 338 66 354 100
rect 388 66 396 100
rect 338 46 396 66
rect 450 100 508 176
rect 450 66 458 100
rect 492 66 508 100
rect 450 46 508 66
rect 538 46 604 176
rect 634 100 700 176
rect 634 66 650 100
rect 684 66 700 100
rect 634 46 700 66
rect 730 46 796 176
rect 826 100 884 176
rect 826 66 842 100
rect 876 66 884 100
rect 826 46 884 66
rect 938 100 996 176
rect 938 66 946 100
rect 980 66 996 100
rect 938 46 996 66
rect 1026 46 1092 176
rect 1122 100 1188 176
rect 1122 66 1138 100
rect 1172 66 1188 100
rect 1122 46 1188 66
rect 1218 100 1284 176
rect 1218 66 1234 100
rect 1268 66 1284 100
rect 1218 46 1284 66
rect 1314 100 1372 176
rect 1314 66 1330 100
rect 1364 66 1372 100
rect 1314 46 1372 66
rect 1426 100 1484 176
rect 1426 66 1434 100
rect 1468 66 1484 100
rect 1426 46 1484 66
rect 1514 100 1580 176
rect 1514 66 1530 100
rect 1564 66 1580 100
rect 1514 46 1580 66
rect 1610 100 1676 176
rect 1610 66 1626 100
rect 1660 66 1676 100
rect 1610 46 1676 66
rect 1706 100 1764 176
rect 1706 66 1722 100
rect 1756 66 1764 100
rect 1706 46 1764 66
rect 1818 100 1876 176
rect 1818 66 1826 100
rect 1860 66 1876 100
rect 1818 46 1876 66
rect 1906 100 1972 176
rect 1906 66 1922 100
rect 1956 66 1972 100
rect 1906 46 1972 66
rect 2002 100 2068 176
rect 2002 66 2018 100
rect 2052 66 2068 100
rect 2002 46 2068 66
rect 2098 100 2164 176
rect 2098 66 2114 100
rect 2148 66 2164 100
rect 2098 46 2164 66
rect 2194 100 2252 176
rect 2194 66 2210 100
rect 2244 66 2252 100
rect 2194 46 2252 66
<< pdiff >>
rect 58 406 116 496
rect 58 372 66 406
rect 100 372 116 406
rect 58 296 116 372
rect 146 476 212 496
rect 146 442 162 476
rect 196 442 212 476
rect 146 296 212 442
rect 242 378 308 496
rect 242 344 258 378
rect 292 344 308 378
rect 242 296 308 344
rect 338 476 396 496
rect 338 442 354 476
rect 388 442 396 476
rect 338 296 396 442
rect 450 378 508 496
rect 450 344 458 378
rect 492 344 508 378
rect 450 296 508 344
rect 538 476 604 496
rect 538 442 554 476
rect 588 442 604 476
rect 538 296 604 442
rect 634 378 700 496
rect 634 344 650 378
rect 684 344 700 378
rect 634 296 700 344
rect 730 378 796 496
rect 730 344 746 378
rect 780 344 796 378
rect 730 296 796 344
rect 826 378 884 496
rect 826 344 842 378
rect 876 344 884 378
rect 826 296 884 344
rect 938 476 996 496
rect 938 442 946 476
rect 980 442 996 476
rect 938 296 996 442
rect 1026 378 1092 496
rect 1026 344 1042 378
rect 1076 344 1092 378
rect 1026 296 1092 344
rect 1122 476 1188 496
rect 1122 442 1138 476
rect 1172 442 1188 476
rect 1122 296 1188 442
rect 1218 296 1284 496
rect 1314 378 1372 496
rect 1314 344 1330 378
rect 1364 344 1372 378
rect 1314 296 1372 344
rect 1426 446 1484 496
rect 1426 412 1434 446
rect 1468 412 1484 446
rect 1426 296 1484 412
rect 1514 476 1580 496
rect 1514 442 1530 476
rect 1564 442 1580 476
rect 1514 296 1580 442
rect 1610 296 1676 496
rect 1706 378 1764 496
rect 1706 344 1722 378
rect 1756 344 1764 378
rect 1706 296 1764 344
rect 1818 378 1876 496
rect 1818 344 1826 378
rect 1860 344 1876 378
rect 1818 296 1876 344
rect 1906 296 1972 496
rect 2002 476 2068 496
rect 2002 442 2018 476
rect 2052 442 2068 476
rect 2002 296 2068 442
rect 2098 296 2164 496
rect 2194 378 2252 496
rect 2194 344 2210 378
rect 2244 344 2252 378
rect 2194 296 2252 344
<< ndiffc >>
rect 66 66 100 100
rect 162 66 196 100
rect 354 66 388 100
rect 458 66 492 100
rect 650 66 684 100
rect 842 66 876 100
rect 946 66 980 100
rect 1138 66 1172 100
rect 1234 66 1268 100
rect 1330 66 1364 100
rect 1434 66 1468 100
rect 1530 66 1564 100
rect 1626 66 1660 100
rect 1722 66 1756 100
rect 1826 66 1860 100
rect 1922 66 1956 100
rect 2018 66 2052 100
rect 2114 66 2148 100
rect 2210 66 2244 100
<< pdiffc >>
rect 66 372 100 406
rect 162 442 196 476
rect 258 344 292 378
rect 354 442 388 476
rect 458 344 492 378
rect 554 442 588 476
rect 650 344 684 378
rect 746 344 780 378
rect 842 344 876 378
rect 946 442 980 476
rect 1042 344 1076 378
rect 1138 442 1172 476
rect 1330 344 1364 378
rect 1434 412 1468 446
rect 1530 442 1564 476
rect 1722 344 1756 378
rect 1826 344 1860 378
rect 2018 442 2052 476
rect 2210 344 2244 378
<< poly >>
rect 116 496 146 522
rect 212 496 242 522
rect 308 496 338 522
rect 508 496 538 522
rect 604 496 634 522
rect 700 496 730 522
rect 796 496 826 522
rect 996 496 1026 522
rect 1092 496 1122 522
rect 1188 496 1218 522
rect 1284 496 1314 522
rect 1484 496 1514 522
rect 1580 496 1610 522
rect 1676 496 1706 522
rect 1876 496 1906 522
rect 1972 496 2002 522
rect 2068 496 2098 522
rect 2164 496 2194 522
rect 116 264 146 296
rect 212 264 242 296
rect 308 264 338 296
rect 508 264 538 296
rect 604 264 634 296
rect 700 264 730 296
rect 796 264 826 296
rect 996 264 1026 296
rect 1092 264 1122 296
rect 1188 264 1218 296
rect 1284 264 1314 296
rect 1484 264 1514 296
rect 1580 264 1610 296
rect 1676 264 1706 296
rect 1876 264 1906 296
rect 1972 264 2002 296
rect 2068 264 2098 296
rect 2164 264 2194 296
rect 104 248 158 264
rect 104 214 114 248
rect 148 214 158 248
rect 104 198 158 214
rect 200 248 254 264
rect 200 214 210 248
rect 244 214 254 248
rect 200 198 254 214
rect 296 248 350 264
rect 296 214 306 248
rect 340 214 350 248
rect 296 198 350 214
rect 496 248 550 264
rect 496 214 506 248
rect 540 214 550 248
rect 496 198 550 214
rect 592 248 646 264
rect 592 214 602 248
rect 636 214 646 248
rect 592 198 646 214
rect 688 248 742 264
rect 688 214 698 248
rect 732 214 742 248
rect 688 198 742 214
rect 784 248 838 264
rect 784 214 794 248
rect 828 214 838 248
rect 784 198 838 214
rect 984 248 1038 264
rect 984 214 994 248
rect 1028 214 1038 248
rect 984 198 1038 214
rect 1080 248 1134 264
rect 1080 214 1090 248
rect 1124 214 1134 248
rect 1080 198 1134 214
rect 1176 248 1230 264
rect 1176 214 1186 248
rect 1220 214 1230 248
rect 1176 198 1230 214
rect 1272 248 1326 264
rect 1272 214 1282 248
rect 1316 214 1326 248
rect 1272 198 1326 214
rect 1472 248 1526 264
rect 1472 214 1482 248
rect 1516 214 1526 248
rect 1472 198 1526 214
rect 1568 248 1622 264
rect 1568 214 1578 248
rect 1612 214 1622 248
rect 1568 198 1622 214
rect 1664 248 1718 264
rect 1664 214 1674 248
rect 1708 214 1718 248
rect 1664 198 1718 214
rect 1864 248 1918 264
rect 1864 214 1874 248
rect 1908 214 1918 248
rect 1864 198 1918 214
rect 1960 248 2014 264
rect 1960 214 1970 248
rect 2004 214 2014 248
rect 1960 198 2014 214
rect 2056 248 2110 264
rect 2056 214 2066 248
rect 2100 214 2110 248
rect 2056 198 2110 214
rect 2152 248 2206 264
rect 2152 214 2162 248
rect 2196 214 2206 248
rect 2152 198 2206 214
rect 116 176 146 198
rect 212 176 242 198
rect 308 176 338 198
rect 508 176 538 198
rect 604 176 634 198
rect 700 176 730 198
rect 796 176 826 198
rect 996 176 1026 198
rect 1092 176 1122 198
rect 1188 176 1218 198
rect 1284 176 1314 198
rect 1484 176 1514 198
rect 1580 176 1610 198
rect 1676 176 1706 198
rect 1876 176 1906 198
rect 1972 176 2002 198
rect 2068 176 2098 198
rect 2164 176 2194 198
rect 116 20 146 46
rect 212 20 242 46
rect 308 20 338 46
rect 508 20 538 46
rect 604 20 634 46
rect 700 20 730 46
rect 796 20 826 46
rect 996 20 1026 46
rect 1092 20 1122 46
rect 1188 20 1218 46
rect 1284 20 1314 46
rect 1484 20 1514 46
rect 1580 20 1610 46
rect 1676 20 1706 46
rect 1876 20 1906 46
rect 1972 20 2002 46
rect 2068 20 2098 46
rect 2164 20 2194 46
<< polycont >>
rect 114 214 148 248
rect 210 214 244 248
rect 306 214 340 248
rect 506 214 540 248
rect 602 214 636 248
rect 698 214 732 248
rect 794 214 828 248
rect 994 214 1028 248
rect 1090 214 1124 248
rect 1186 214 1220 248
rect 1282 214 1316 248
rect 1482 214 1516 248
rect 1578 214 1612 248
rect 1674 214 1708 248
rect 1874 214 1908 248
rect 1970 214 2004 248
rect 2066 214 2100 248
rect 2162 214 2196 248
<< locali >>
rect 0 526 28 560
rect 62 526 120 560
rect 154 526 212 560
rect 246 526 304 560
rect 338 526 396 560
rect 430 526 488 560
rect 522 526 580 560
rect 614 526 672 560
rect 706 526 764 560
rect 798 526 856 560
rect 890 526 948 560
rect 982 526 1040 560
rect 1074 526 1132 560
rect 1166 526 1224 560
rect 1258 526 1316 560
rect 1350 526 1408 560
rect 1442 526 1500 560
rect 1534 526 1592 560
rect 1626 526 1684 560
rect 1718 526 1776 560
rect 1810 526 1868 560
rect 1902 526 1960 560
rect 1994 526 2052 560
rect 2086 526 2144 560
rect 2178 526 2236 560
rect 2270 526 2328 560
rect 2362 526 2392 560
rect 162 476 196 526
rect 162 426 196 442
rect 354 476 388 526
rect 354 426 388 442
rect 554 476 588 526
rect 554 426 588 442
rect 946 476 980 526
rect 946 426 980 442
rect 1138 476 1172 526
rect 1530 476 1564 526
rect 1434 456 1468 462
rect 1138 426 1172 442
rect 66 356 100 372
rect 258 378 292 394
rect 746 378 780 394
rect 134 328 258 362
rect 442 344 458 378
rect 492 344 650 378
rect 684 344 700 378
rect 134 316 168 328
rect 114 282 168 316
rect 330 310 354 344
rect 1330 378 1364 422
rect 2018 476 2052 526
rect 1530 426 1564 442
rect 1660 422 1722 456
rect 1434 396 1468 412
rect 1026 344 1042 378
rect 1076 344 1124 378
rect 1698 378 1756 422
rect 1898 422 1922 456
rect 2018 426 2052 442
rect 1698 344 1722 378
rect 842 328 876 344
rect 1124 310 1292 344
rect 1330 328 1364 344
rect 114 268 148 282
rect 66 248 148 268
rect 66 214 114 248
rect 114 198 148 214
rect 210 248 244 264
rect 330 248 364 310
rect 602 248 636 254
rect 290 214 306 248
rect 340 214 364 248
rect 440 232 506 248
rect 474 214 506 232
rect 540 214 556 248
rect 602 198 636 214
rect 698 248 732 264
rect 946 248 980 310
rect 1258 264 1292 310
rect 1722 328 1756 344
rect 1826 378 1860 394
rect 1468 310 1612 316
rect 1898 344 1932 422
rect 2066 344 2210 378
rect 2244 344 2260 378
rect 1898 310 1922 344
rect 1434 282 1612 310
rect 1090 248 1124 264
rect 778 214 794 248
rect 828 232 876 248
rect 828 214 842 232
rect 946 214 994 248
rect 1028 214 1044 248
rect 1186 248 1220 264
rect 1258 248 1316 264
rect 1578 248 1612 282
rect 1674 254 1722 268
rect 1674 248 1756 254
rect 1898 248 1932 310
rect 1258 214 1282 248
rect 1282 198 1316 214
rect 1434 232 1482 248
rect 1468 214 1482 232
rect 1516 214 1532 248
rect 1658 214 1674 248
rect 1708 234 1756 248
rect 1708 214 1724 234
rect 1858 214 1874 248
rect 1908 214 1932 248
rect 1970 248 2004 264
rect 2162 248 2196 254
rect 2004 214 2066 248
rect 2100 214 2116 248
rect 1578 198 1612 214
rect 2162 198 2196 214
rect 66 50 100 66
rect 162 100 196 116
rect 458 100 492 116
rect 292 86 354 100
rect 258 66 354 86
rect 388 66 404 100
rect 634 66 650 100
rect 684 86 746 100
rect 684 66 780 86
rect 842 100 876 116
rect 930 66 946 100
rect 980 86 1042 100
rect 980 66 1076 86
rect 1138 100 1172 116
rect 162 16 196 66
rect 458 16 492 66
rect 842 16 876 66
rect 1138 16 1172 66
rect 1234 50 1268 66
rect 1330 100 1364 116
rect 1330 16 1364 66
rect 1434 50 1468 66
rect 1530 100 1564 116
rect 1530 16 1564 66
rect 1626 50 1660 66
rect 1722 100 1756 116
rect 1722 16 1756 66
rect 1826 100 1860 116
rect 1826 16 1860 66
rect 1922 50 1956 66
rect 2018 100 2052 116
rect 2018 16 2052 66
rect 2114 50 2148 66
rect 2210 100 2244 116
rect 2210 16 2244 66
rect 0 -18 28 16
rect 62 -18 120 16
rect 154 -18 212 16
rect 246 -18 304 16
rect 338 -18 396 16
rect 430 -18 488 16
rect 522 -18 580 16
rect 614 -18 672 16
rect 706 -18 764 16
rect 798 -18 856 16
rect 890 -18 948 16
rect 982 -18 1040 16
rect 1074 -18 1132 16
rect 1166 -18 1224 16
rect 1258 -18 1316 16
rect 1350 -18 1408 16
rect 1442 -18 1500 16
rect 1534 -18 1592 16
rect 1626 -18 1684 16
rect 1718 -18 1776 16
rect 1810 -18 1868 16
rect 1902 -18 1960 16
rect 1994 -18 2052 16
rect 2086 -18 2144 16
rect 2178 -18 2236 16
rect 2270 -18 2328 16
rect 2362 -18 2392 16
<< viali >>
rect 28 526 62 560
rect 120 526 154 560
rect 212 526 246 560
rect 304 526 338 560
rect 396 526 430 560
rect 488 526 522 560
rect 580 526 614 560
rect 672 526 706 560
rect 764 526 798 560
rect 856 526 890 560
rect 948 526 982 560
rect 1040 526 1074 560
rect 1132 526 1166 560
rect 1224 526 1258 560
rect 1316 526 1350 560
rect 1408 526 1442 560
rect 1500 526 1534 560
rect 1592 526 1626 560
rect 1684 526 1718 560
rect 1776 526 1810 560
rect 1868 526 1902 560
rect 1960 526 1994 560
rect 2052 526 2086 560
rect 2144 526 2178 560
rect 2236 526 2270 560
rect 2328 526 2362 560
rect 66 406 100 428
rect 66 394 100 406
rect 1330 422 1364 456
rect 650 378 684 400
rect 650 366 684 378
rect 258 310 292 344
rect 354 310 388 344
rect 746 310 780 344
rect 842 378 876 400
rect 1434 446 1468 456
rect 1434 422 1468 446
rect 1626 422 1660 456
rect 1722 422 1756 456
rect 842 366 876 378
rect 1922 422 1956 456
rect 946 310 980 344
rect 1090 310 1124 344
rect 602 254 636 288
rect 210 214 244 232
rect 210 198 244 214
rect 440 198 474 232
rect 1434 310 1468 344
rect 1826 310 1860 344
rect 1922 310 1956 344
rect 2066 310 2100 344
rect 698 214 732 232
rect 698 198 732 214
rect 842 198 876 232
rect 1090 214 1124 232
rect 1090 198 1124 214
rect 1186 214 1220 232
rect 1722 254 1756 288
rect 1186 198 1220 214
rect 1434 198 1468 232
rect 2162 254 2196 288
rect 1970 214 2004 232
rect 1970 198 2004 214
rect 66 100 100 120
rect 66 86 100 100
rect 258 86 292 120
rect 746 86 780 120
rect 1042 86 1076 120
rect 1234 100 1268 120
rect 1234 86 1268 100
rect 1434 100 1468 120
rect 1434 86 1468 100
rect 1626 100 1660 120
rect 1626 86 1660 100
rect 1922 100 1956 120
rect 1922 86 1956 100
rect 2114 100 2148 120
rect 2114 86 2148 100
rect 28 -18 62 16
rect 120 -18 154 16
rect 212 -18 246 16
rect 304 -18 338 16
rect 396 -18 430 16
rect 488 -18 522 16
rect 580 -18 614 16
rect 672 -18 706 16
rect 764 -18 798 16
rect 856 -18 890 16
rect 948 -18 982 16
rect 1040 -18 1074 16
rect 1132 -18 1166 16
rect 1224 -18 1258 16
rect 1316 -18 1350 16
rect 1408 -18 1442 16
rect 1500 -18 1534 16
rect 1592 -18 1626 16
rect 1684 -18 1718 16
rect 1776 -18 1810 16
rect 1868 -18 1902 16
rect 1960 -18 1994 16
rect 2052 -18 2086 16
rect 2144 -18 2178 16
rect 2236 -18 2270 16
rect 2328 -18 2362 16
<< metal1 >>
rect 0 560 2392 592
rect 0 526 28 560
rect 62 526 120 560
rect 154 526 212 560
rect 246 526 304 560
rect 338 526 396 560
rect 430 526 488 560
rect 522 526 580 560
rect 614 526 672 560
rect 706 526 764 560
rect 798 526 856 560
rect 890 526 948 560
rect 982 526 1040 560
rect 1074 526 1132 560
rect 1166 526 1224 560
rect 1258 526 1316 560
rect 1350 526 1408 560
rect 1442 526 1500 560
rect 1534 526 1592 560
rect 1626 526 1684 560
rect 1718 526 1776 560
rect 1810 526 1868 560
rect 1902 526 1960 560
rect 1994 526 2052 560
rect 2086 526 2144 560
rect 2178 526 2236 560
rect 2270 526 2328 560
rect 2362 526 2392 560
rect 0 520 2392 526
rect 50 428 114 434
rect 50 410 66 428
rect 100 410 114 428
rect 50 358 56 410
rect 108 358 114 410
rect 652 406 872 420
rect 1002 414 1008 466
rect 1060 454 1066 466
rect 1060 426 1216 454
rect 1060 414 1066 426
rect 638 400 888 406
rect 638 366 650 400
rect 684 392 842 400
rect 684 366 696 392
rect 638 360 696 366
rect 830 366 842 392
rect 876 366 888 400
rect 830 360 888 366
rect 50 352 114 358
rect 66 126 98 352
rect 242 302 248 354
rect 300 302 306 354
rect 338 302 344 354
rect 396 302 402 354
rect 466 302 472 354
rect 524 330 530 354
rect 734 344 792 350
rect 524 302 632 330
rect 734 310 746 344
rect 780 342 792 344
rect 780 310 800 342
rect 734 304 800 310
rect 590 294 632 302
rect 590 288 648 294
rect 590 254 602 288
rect 636 254 648 288
rect 590 248 648 254
rect 686 242 744 248
rect 146 190 152 242
rect 204 238 210 242
rect 204 232 336 238
rect 204 198 210 232
rect 244 210 336 232
rect 428 232 486 238
rect 428 230 440 232
rect 244 198 256 210
rect 204 192 256 198
rect 308 202 336 210
rect 408 202 440 230
rect 308 198 440 202
rect 474 198 486 232
rect 686 202 688 242
rect 308 192 486 198
rect 204 190 210 192
rect 308 174 436 192
rect 532 190 688 202
rect 740 190 744 242
rect 532 174 744 190
rect 54 120 112 126
rect 54 86 66 120
rect 100 86 112 120
rect 54 80 112 86
rect 242 78 248 130
rect 300 118 306 130
rect 634 118 640 130
rect 300 90 640 118
rect 300 78 306 90
rect 634 78 640 90
rect 692 78 698 130
rect 772 126 800 304
rect 930 302 936 354
rect 988 302 994 354
rect 1074 302 1080 354
rect 1132 302 1138 354
rect 1188 342 1216 426
rect 1314 414 1320 466
rect 1372 414 1378 466
rect 1422 456 1480 462
rect 1422 422 1434 456
rect 1468 454 1480 456
rect 1514 454 1520 466
rect 1468 426 1520 454
rect 1468 422 1480 426
rect 1422 416 1480 422
rect 1514 414 1520 426
rect 1572 414 1578 466
rect 1610 414 1616 466
rect 1668 414 1674 466
rect 1706 414 1712 466
rect 1764 414 1770 466
rect 1906 414 1912 466
rect 1964 420 1970 466
rect 1964 414 2192 420
rect 1924 392 2192 414
rect 1422 344 1480 350
rect 1422 342 1434 344
rect 1188 314 1434 342
rect 1422 310 1434 314
rect 1468 310 1480 344
rect 1422 304 1480 310
rect 1810 302 1816 354
rect 1868 302 1874 354
rect 1924 350 1952 392
rect 1910 344 1968 350
rect 1910 310 1922 344
rect 1956 310 1968 344
rect 1910 304 1968 310
rect 2054 344 2112 350
rect 2054 310 2066 344
rect 2100 342 2112 344
rect 2100 310 2120 342
rect 2054 304 2120 310
rect 1710 288 1768 294
rect 1710 254 1722 288
rect 1756 286 1768 288
rect 1810 286 1856 302
rect 1756 258 1856 286
rect 1756 254 1768 258
rect 1710 248 1768 254
rect 878 238 884 242
rect 830 232 884 238
rect 830 198 842 232
rect 876 198 884 232
rect 830 192 884 198
rect 878 190 884 192
rect 936 230 942 242
rect 1078 232 1136 238
rect 1078 230 1090 232
rect 936 202 1090 230
rect 936 190 942 202
rect 1078 198 1090 202
rect 1124 198 1136 232
rect 1078 192 1136 198
rect 1174 232 1232 238
rect 1174 198 1186 232
rect 1220 230 1232 232
rect 1220 202 1360 230
rect 1220 198 1232 202
rect 1174 192 1232 198
rect 734 120 800 126
rect 734 86 746 120
rect 780 118 800 120
rect 930 118 936 130
rect 780 90 936 118
rect 780 86 792 90
rect 734 80 792 86
rect 930 78 936 90
rect 988 78 994 130
rect 1074 126 1080 130
rect 1030 120 1080 126
rect 1030 86 1042 120
rect 1076 86 1080 120
rect 1030 80 1080 86
rect 1074 78 1080 80
rect 1132 78 1138 130
rect 1218 78 1224 130
rect 1276 78 1282 130
rect 1332 118 1360 202
rect 1418 190 1424 242
rect 1476 202 1482 242
rect 1958 232 2016 238
rect 1958 202 1970 232
rect 1476 198 1970 202
rect 2004 198 2016 232
rect 1476 192 2016 198
rect 1476 190 2000 192
rect 1436 174 2000 190
rect 2092 130 2120 304
rect 2164 294 2192 392
rect 2150 288 2208 294
rect 2150 254 2162 288
rect 2196 254 2208 288
rect 2150 248 2208 254
rect 1466 126 1472 130
rect 1422 120 1472 126
rect 1422 118 1434 120
rect 1332 90 1434 118
rect 1422 86 1434 90
rect 1468 86 1472 120
rect 1422 80 1472 86
rect 1466 78 1472 80
rect 1524 78 1530 130
rect 1586 78 1592 130
rect 1644 120 1722 130
rect 1660 86 1722 120
rect 1644 78 1722 86
rect 1810 78 1816 130
rect 1868 118 1874 130
rect 1910 120 1968 126
rect 1910 118 1922 120
rect 1868 90 1922 118
rect 1868 78 1874 90
rect 1910 86 1922 90
rect 1956 86 1968 120
rect 2092 90 2104 130
rect 1910 80 1968 86
rect 2098 78 2104 90
rect 2156 78 2162 130
rect 0 16 2392 22
rect 0 -18 28 16
rect 62 -18 120 16
rect 154 -18 212 16
rect 246 -18 304 16
rect 338 -18 396 16
rect 430 -18 488 16
rect 522 -18 580 16
rect 614 -18 672 16
rect 706 -18 764 16
rect 798 -18 856 16
rect 890 -18 948 16
rect 982 -18 1040 16
rect 1074 -18 1132 16
rect 1166 -18 1224 16
rect 1258 -18 1316 16
rect 1350 -18 1408 16
rect 1442 -18 1500 16
rect 1534 -18 1592 16
rect 1626 -18 1684 16
rect 1718 -18 1776 16
rect 1810 -18 1868 16
rect 1902 -18 1960 16
rect 1994 -18 2052 16
rect 2086 -18 2144 16
rect 2178 -18 2236 16
rect 2270 -18 2328 16
rect 2362 -18 2392 16
rect 0 -48 2392 -18
<< via1 >>
rect 56 394 66 410
rect 66 394 100 410
rect 100 394 108 410
rect 56 358 108 394
rect 1008 414 1060 466
rect 248 344 300 354
rect 248 310 258 344
rect 258 310 292 344
rect 292 310 300 344
rect 248 302 300 310
rect 344 344 396 354
rect 344 310 354 344
rect 354 310 388 344
rect 388 310 396 344
rect 344 302 396 310
rect 472 302 524 354
rect 152 190 204 242
rect 688 232 740 242
rect 688 198 698 232
rect 698 198 732 232
rect 732 198 740 232
rect 688 190 740 198
rect 248 120 300 130
rect 248 86 258 120
rect 258 86 292 120
rect 292 86 300 120
rect 248 78 300 86
rect 640 78 692 130
rect 936 344 988 354
rect 936 310 946 344
rect 946 310 980 344
rect 980 310 988 344
rect 936 302 988 310
rect 1080 344 1132 354
rect 1080 310 1090 344
rect 1090 310 1124 344
rect 1124 310 1132 344
rect 1080 302 1132 310
rect 1320 456 1372 466
rect 1320 422 1330 456
rect 1330 422 1364 456
rect 1364 422 1372 456
rect 1320 414 1372 422
rect 1520 414 1572 466
rect 1616 456 1668 466
rect 1616 422 1626 456
rect 1626 422 1660 456
rect 1660 422 1668 456
rect 1616 414 1668 422
rect 1712 456 1764 466
rect 1712 422 1722 456
rect 1722 422 1756 456
rect 1756 422 1764 456
rect 1712 414 1764 422
rect 1912 456 1964 466
rect 1912 422 1922 456
rect 1922 422 1956 456
rect 1956 422 1964 456
rect 1912 414 1964 422
rect 1816 344 1868 354
rect 1816 310 1826 344
rect 1826 310 1860 344
rect 1860 310 1868 344
rect 1816 302 1868 310
rect 884 190 936 242
rect 936 78 988 130
rect 1080 78 1132 130
rect 1224 120 1276 130
rect 1224 86 1234 120
rect 1234 86 1268 120
rect 1268 86 1276 120
rect 1224 78 1276 86
rect 1424 232 1476 242
rect 1424 198 1434 232
rect 1434 198 1468 232
rect 1468 198 1476 232
rect 1424 190 1476 198
rect 1472 78 1524 130
rect 1592 120 1644 130
rect 1592 86 1626 120
rect 1626 86 1644 120
rect 1592 78 1644 86
rect 1816 78 1868 130
rect 2104 120 2156 130
rect 2104 86 2114 120
rect 2114 86 2148 120
rect 2148 86 2156 120
rect 2104 78 2156 86
<< metal2 >>
rect 54 468 110 477
rect 54 410 110 412
rect 54 402 56 410
rect 108 402 110 410
rect 1008 466 1060 472
rect 1008 408 1060 414
rect 1318 468 1374 477
rect 542 360 598 365
rect 56 352 108 358
rect 248 354 300 360
rect 344 354 396 360
rect 248 296 300 302
rect 332 302 344 342
rect 332 296 396 302
rect 472 356 598 360
rect 472 354 542 356
rect 524 302 542 354
rect 472 300 542 302
rect 936 354 988 360
rect 598 314 936 342
rect 472 296 598 300
rect 936 296 988 302
rect 150 244 206 253
rect 150 178 206 188
rect 260 136 288 296
rect 332 230 360 296
rect 542 290 598 296
rect 394 244 450 253
rect 830 248 886 253
rect 332 202 394 230
rect 688 242 740 248
rect 450 202 688 230
rect 394 178 450 188
rect 688 184 740 190
rect 830 244 936 248
rect 886 242 936 244
rect 886 188 936 190
rect 830 184 936 188
rect 830 178 886 184
rect 248 130 300 136
rect 248 72 300 78
rect 640 130 692 136
rect 936 130 988 136
rect 692 90 848 118
rect 640 72 692 78
rect 820 42 848 90
rect 1020 118 1048 408
rect 1318 402 1374 412
rect 1520 466 1572 472
rect 1520 408 1572 414
rect 1616 466 1668 472
rect 1616 408 1668 414
rect 1710 468 1766 477
rect 1078 356 1134 365
rect 1332 364 1360 402
rect 1294 342 1360 364
rect 1078 290 1134 300
rect 1236 314 1360 342
rect 1092 136 1120 290
rect 1236 136 1264 314
rect 1294 290 1350 314
rect 1424 242 1476 248
rect 1308 202 1424 230
rect 988 90 1048 118
rect 1080 130 1132 136
rect 936 72 988 78
rect 1080 72 1132 78
rect 1224 130 1276 136
rect 1224 72 1276 78
rect 1308 42 1336 202
rect 1424 184 1476 190
rect 1532 136 1560 408
rect 1616 398 1656 408
rect 1710 402 1766 412
rect 1910 468 1966 477
rect 1910 402 1966 412
rect 1604 364 1656 398
rect 1604 290 1704 364
rect 1816 354 1868 360
rect 1816 296 1868 302
rect 1604 136 1632 290
rect 1828 136 1856 296
rect 1472 130 1560 136
rect 1524 90 1560 130
rect 1592 130 1644 136
rect 1472 72 1524 78
rect 1592 72 1644 78
rect 1816 130 1868 136
rect 1816 72 1868 78
rect 2102 132 2158 141
rect 2102 66 2158 76
rect 820 14 1336 42
<< via2 >>
rect 54 412 110 468
rect 1318 466 1374 468
rect 1318 414 1320 466
rect 1320 414 1372 466
rect 1372 414 1374 466
rect 1318 412 1374 414
rect 542 300 598 356
rect 150 242 206 244
rect 150 190 152 242
rect 152 190 204 242
rect 204 190 206 242
rect 150 188 206 190
rect 394 188 450 244
rect 830 242 886 244
rect 830 190 884 242
rect 884 190 886 242
rect 830 188 886 190
rect 1710 466 1766 468
rect 1710 414 1712 466
rect 1712 414 1764 466
rect 1764 414 1766 466
rect 1710 412 1766 414
rect 1078 354 1134 356
rect 1078 302 1080 354
rect 1080 302 1132 354
rect 1132 302 1134 354
rect 1078 300 1134 302
rect 1910 466 1966 468
rect 1910 414 1912 466
rect 1912 414 1964 466
rect 1964 414 1966 466
rect 1910 412 1966 414
rect 2102 130 2158 132
rect 2102 78 2104 130
rect 2104 78 2156 130
rect 2156 78 2158 130
rect 2102 76 2158 78
<< metal3 >>
rect 49 472 114 473
rect 1313 472 1379 473
rect 1706 472 1771 473
rect 1907 472 1971 473
rect 49 468 196 472
rect 49 412 54 468
rect 110 412 196 468
rect 49 406 196 412
rect 1313 468 1460 472
rect 1313 412 1318 468
rect 1374 412 1460 468
rect 1313 406 1460 412
rect 1654 468 1800 472
rect 1654 412 1710 468
rect 1766 412 1800 468
rect 1654 406 1800 412
rect 1860 468 1972 472
rect 1860 412 1910 468
rect 1966 412 1972 468
rect 1860 406 1972 412
rect 49 405 114 406
rect 1313 405 1379 406
rect 1706 405 1771 406
rect 537 360 603 361
rect 1073 360 1137 361
rect 537 356 684 360
rect 537 300 542 356
rect 598 300 684 356
rect 537 294 684 300
rect 1073 356 1184 360
rect 1073 300 1078 356
rect 1134 300 1184 356
rect 537 293 603 294
rect 1073 293 1184 300
rect 116 248 220 249
rect 390 248 455 249
rect 825 248 890 249
rect 116 244 262 248
rect 116 188 150 244
rect 206 188 262 244
rect 116 182 262 188
rect 322 244 468 248
rect 322 188 394 244
rect 450 188 468 244
rect 322 182 468 188
rect 825 244 972 248
rect 825 188 830 244
rect 886 188 972 244
rect 825 182 972 188
rect 390 181 455 182
rect 825 181 890 182
rect 1124 134 1184 293
rect 1860 134 1920 406
rect 1124 74 1920 134
rect 2097 136 2162 137
rect 2097 132 2244 136
rect 2097 76 2102 132
rect 2158 76 2244 132
rect 2097 70 2244 76
rect 2097 69 2162 70
<< labels >>
flabel nwell s 1792 526 1826 560 0 FreeSans 100 0 0 0 VPB
port 1 nsew
flabel nwell s 1400 526 1434 560 0 FreeSans 100 0 0 0 VPB
port 1 nsew
flabel nwell s 912 526 946 560 0 FreeSans 100 0 0 0 VPB
port 1 nsew
flabel nwell s 424 526 458 560 0 FreeSans 100 0 0 0 VPB
port 1 nsew
flabel nwell s 32 526 66 560 0 FreeSans 100 0 0 0 VPB
port 1 nsew
flabel pwell s 1792 -16 1826 16 0 FreeSans 100 0 0 0 VNB
port 2 nsew
flabel pwell s 1400 -16 1434 16 0 FreeSans 100 0 0 0 VNB
port 2 nsew
flabel pwell s 912 -16 946 16 0 FreeSans 100 0 0 0 VNB
port 2 nsew
flabel pwell s 424 -16 458 16 0 FreeSans 100 0 0 0 VNB
port 2 nsew
flabel pwell s 32 -16 66 16 0 FreeSans 100 0 0 0 VNB
port 2 nsew
flabel comment s 0 0 0 0 0 FreeSans 100 0 0 0 mul2
rlabel metal3 s 322 182 468 248 4 B0
port 3 nsew
rlabel metal3 s 116 182 262 248 4 A0
port 4 nsew
rlabel metal3 s 538 294 684 360 4 B1
port 5 nsew
rlabel metal3 s 1654 406 1800 472 4 R1
port 6 nsew
rlabel metal3 s 1314 406 1460 472 4 R2
port 7 nsew
rlabel metal3 s 50 406 196 472 4 R0
port 8 nsew
rlabel metal3 s 2098 70 2244 136 4 R3
port 9 nsew
rlabel metal3 s 826 182 972 248 4 A1
port 10 nsew
flabel metal1 s 30 526 64 560 0 FreeSans 100 0 0 0 vpwr
port 11 nsew
flabel metal1 s 30 -16 64 16 0 FreeSans 100 0 0 0 vgnd
port 12 nsew
<< properties >>
string FIXED_BBOX 0 0 2392 544
<< end >>
